module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(a[0], b[0], ha_xor0);
  and_gate and_gate_ha_and0(a[0], b[0], ha_and0);
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(a[0], b[0], fa_xor0);
  and_gate and_gate_fa_and0(a[0], b[0], fa_and0);
  xor_gate xor_gate_fa_xor1(fa_xor0[0], cin[0], fa_xor1);
  and_gate and_gate_fa_and1(fa_xor0[0], cin[0], fa_and1);
  or_gate or_gate_fa_or0(fa_and0[0], fa_and1[0], fa_or0);
endmodule

module pg_fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] pg_fa_xor0, output [0:0] pg_fa_and0, output [0:0] pg_fa_xor1);
  xor_gate xor_gate_pg_fa_xor0(a[0], b[0], pg_fa_xor0);
  and_gate and_gate_pg_fa_and0(a[0], b[0], pg_fa_and0);
  xor_gate xor_gate_pg_fa_xor1(pg_fa_xor0[0], cin[0], pg_fa_xor1);
endmodule

module u_pg_rca62(input [61:0] a, input [61:0] b, output [62:0] u_pg_rca62_out);
  wire [0:0] u_pg_rca62_pg_fa0_xor0;
  wire [0:0] u_pg_rca62_pg_fa0_and0;
  wire [0:0] u_pg_rca62_pg_fa1_xor0;
  wire [0:0] u_pg_rca62_pg_fa1_and0;
  wire [0:0] u_pg_rca62_pg_fa1_xor1;
  wire [0:0] u_pg_rca62_and1;
  wire [0:0] u_pg_rca62_or1;
  wire [0:0] u_pg_rca62_pg_fa2_xor0;
  wire [0:0] u_pg_rca62_pg_fa2_and0;
  wire [0:0] u_pg_rca62_pg_fa2_xor1;
  wire [0:0] u_pg_rca62_and2;
  wire [0:0] u_pg_rca62_or2;
  wire [0:0] u_pg_rca62_pg_fa3_xor0;
  wire [0:0] u_pg_rca62_pg_fa3_and0;
  wire [0:0] u_pg_rca62_pg_fa3_xor1;
  wire [0:0] u_pg_rca62_and3;
  wire [0:0] u_pg_rca62_or3;
  wire [0:0] u_pg_rca62_pg_fa4_xor0;
  wire [0:0] u_pg_rca62_pg_fa4_and0;
  wire [0:0] u_pg_rca62_pg_fa4_xor1;
  wire [0:0] u_pg_rca62_and4;
  wire [0:0] u_pg_rca62_or4;
  wire [0:0] u_pg_rca62_pg_fa5_xor0;
  wire [0:0] u_pg_rca62_pg_fa5_and0;
  wire [0:0] u_pg_rca62_pg_fa5_xor1;
  wire [0:0] u_pg_rca62_and5;
  wire [0:0] u_pg_rca62_or5;
  wire [0:0] u_pg_rca62_pg_fa6_xor0;
  wire [0:0] u_pg_rca62_pg_fa6_and0;
  wire [0:0] u_pg_rca62_pg_fa6_xor1;
  wire [0:0] u_pg_rca62_and6;
  wire [0:0] u_pg_rca62_or6;
  wire [0:0] u_pg_rca62_pg_fa7_xor0;
  wire [0:0] u_pg_rca62_pg_fa7_and0;
  wire [0:0] u_pg_rca62_pg_fa7_xor1;
  wire [0:0] u_pg_rca62_and7;
  wire [0:0] u_pg_rca62_or7;
  wire [0:0] u_pg_rca62_pg_fa8_xor0;
  wire [0:0] u_pg_rca62_pg_fa8_and0;
  wire [0:0] u_pg_rca62_pg_fa8_xor1;
  wire [0:0] u_pg_rca62_and8;
  wire [0:0] u_pg_rca62_or8;
  wire [0:0] u_pg_rca62_pg_fa9_xor0;
  wire [0:0] u_pg_rca62_pg_fa9_and0;
  wire [0:0] u_pg_rca62_pg_fa9_xor1;
  wire [0:0] u_pg_rca62_and9;
  wire [0:0] u_pg_rca62_or9;
  wire [0:0] u_pg_rca62_pg_fa10_xor0;
  wire [0:0] u_pg_rca62_pg_fa10_and0;
  wire [0:0] u_pg_rca62_pg_fa10_xor1;
  wire [0:0] u_pg_rca62_and10;
  wire [0:0] u_pg_rca62_or10;
  wire [0:0] u_pg_rca62_pg_fa11_xor0;
  wire [0:0] u_pg_rca62_pg_fa11_and0;
  wire [0:0] u_pg_rca62_pg_fa11_xor1;
  wire [0:0] u_pg_rca62_and11;
  wire [0:0] u_pg_rca62_or11;
  wire [0:0] u_pg_rca62_pg_fa12_xor0;
  wire [0:0] u_pg_rca62_pg_fa12_and0;
  wire [0:0] u_pg_rca62_pg_fa12_xor1;
  wire [0:0] u_pg_rca62_and12;
  wire [0:0] u_pg_rca62_or12;
  wire [0:0] u_pg_rca62_pg_fa13_xor0;
  wire [0:0] u_pg_rca62_pg_fa13_and0;
  wire [0:0] u_pg_rca62_pg_fa13_xor1;
  wire [0:0] u_pg_rca62_and13;
  wire [0:0] u_pg_rca62_or13;
  wire [0:0] u_pg_rca62_pg_fa14_xor0;
  wire [0:0] u_pg_rca62_pg_fa14_and0;
  wire [0:0] u_pg_rca62_pg_fa14_xor1;
  wire [0:0] u_pg_rca62_and14;
  wire [0:0] u_pg_rca62_or14;
  wire [0:0] u_pg_rca62_pg_fa15_xor0;
  wire [0:0] u_pg_rca62_pg_fa15_and0;
  wire [0:0] u_pg_rca62_pg_fa15_xor1;
  wire [0:0] u_pg_rca62_and15;
  wire [0:0] u_pg_rca62_or15;
  wire [0:0] u_pg_rca62_pg_fa16_xor0;
  wire [0:0] u_pg_rca62_pg_fa16_and0;
  wire [0:0] u_pg_rca62_pg_fa16_xor1;
  wire [0:0] u_pg_rca62_and16;
  wire [0:0] u_pg_rca62_or16;
  wire [0:0] u_pg_rca62_pg_fa17_xor0;
  wire [0:0] u_pg_rca62_pg_fa17_and0;
  wire [0:0] u_pg_rca62_pg_fa17_xor1;
  wire [0:0] u_pg_rca62_and17;
  wire [0:0] u_pg_rca62_or17;
  wire [0:0] u_pg_rca62_pg_fa18_xor0;
  wire [0:0] u_pg_rca62_pg_fa18_and0;
  wire [0:0] u_pg_rca62_pg_fa18_xor1;
  wire [0:0] u_pg_rca62_and18;
  wire [0:0] u_pg_rca62_or18;
  wire [0:0] u_pg_rca62_pg_fa19_xor0;
  wire [0:0] u_pg_rca62_pg_fa19_and0;
  wire [0:0] u_pg_rca62_pg_fa19_xor1;
  wire [0:0] u_pg_rca62_and19;
  wire [0:0] u_pg_rca62_or19;
  wire [0:0] u_pg_rca62_pg_fa20_xor0;
  wire [0:0] u_pg_rca62_pg_fa20_and0;
  wire [0:0] u_pg_rca62_pg_fa20_xor1;
  wire [0:0] u_pg_rca62_and20;
  wire [0:0] u_pg_rca62_or20;
  wire [0:0] u_pg_rca62_pg_fa21_xor0;
  wire [0:0] u_pg_rca62_pg_fa21_and0;
  wire [0:0] u_pg_rca62_pg_fa21_xor1;
  wire [0:0] u_pg_rca62_and21;
  wire [0:0] u_pg_rca62_or21;
  wire [0:0] u_pg_rca62_pg_fa22_xor0;
  wire [0:0] u_pg_rca62_pg_fa22_and0;
  wire [0:0] u_pg_rca62_pg_fa22_xor1;
  wire [0:0] u_pg_rca62_and22;
  wire [0:0] u_pg_rca62_or22;
  wire [0:0] u_pg_rca62_pg_fa23_xor0;
  wire [0:0] u_pg_rca62_pg_fa23_and0;
  wire [0:0] u_pg_rca62_pg_fa23_xor1;
  wire [0:0] u_pg_rca62_and23;
  wire [0:0] u_pg_rca62_or23;
  wire [0:0] u_pg_rca62_pg_fa24_xor0;
  wire [0:0] u_pg_rca62_pg_fa24_and0;
  wire [0:0] u_pg_rca62_pg_fa24_xor1;
  wire [0:0] u_pg_rca62_and24;
  wire [0:0] u_pg_rca62_or24;
  wire [0:0] u_pg_rca62_pg_fa25_xor0;
  wire [0:0] u_pg_rca62_pg_fa25_and0;
  wire [0:0] u_pg_rca62_pg_fa25_xor1;
  wire [0:0] u_pg_rca62_and25;
  wire [0:0] u_pg_rca62_or25;
  wire [0:0] u_pg_rca62_pg_fa26_xor0;
  wire [0:0] u_pg_rca62_pg_fa26_and0;
  wire [0:0] u_pg_rca62_pg_fa26_xor1;
  wire [0:0] u_pg_rca62_and26;
  wire [0:0] u_pg_rca62_or26;
  wire [0:0] u_pg_rca62_pg_fa27_xor0;
  wire [0:0] u_pg_rca62_pg_fa27_and0;
  wire [0:0] u_pg_rca62_pg_fa27_xor1;
  wire [0:0] u_pg_rca62_and27;
  wire [0:0] u_pg_rca62_or27;
  wire [0:0] u_pg_rca62_pg_fa28_xor0;
  wire [0:0] u_pg_rca62_pg_fa28_and0;
  wire [0:0] u_pg_rca62_pg_fa28_xor1;
  wire [0:0] u_pg_rca62_and28;
  wire [0:0] u_pg_rca62_or28;
  wire [0:0] u_pg_rca62_pg_fa29_xor0;
  wire [0:0] u_pg_rca62_pg_fa29_and0;
  wire [0:0] u_pg_rca62_pg_fa29_xor1;
  wire [0:0] u_pg_rca62_and29;
  wire [0:0] u_pg_rca62_or29;
  wire [0:0] u_pg_rca62_pg_fa30_xor0;
  wire [0:0] u_pg_rca62_pg_fa30_and0;
  wire [0:0] u_pg_rca62_pg_fa30_xor1;
  wire [0:0] u_pg_rca62_and30;
  wire [0:0] u_pg_rca62_or30;
  wire [0:0] u_pg_rca62_pg_fa31_xor0;
  wire [0:0] u_pg_rca62_pg_fa31_and0;
  wire [0:0] u_pg_rca62_pg_fa31_xor1;
  wire [0:0] u_pg_rca62_and31;
  wire [0:0] u_pg_rca62_or31;
  wire [0:0] u_pg_rca62_pg_fa32_xor0;
  wire [0:0] u_pg_rca62_pg_fa32_and0;
  wire [0:0] u_pg_rca62_pg_fa32_xor1;
  wire [0:0] u_pg_rca62_and32;
  wire [0:0] u_pg_rca62_or32;
  wire [0:0] u_pg_rca62_pg_fa33_xor0;
  wire [0:0] u_pg_rca62_pg_fa33_and0;
  wire [0:0] u_pg_rca62_pg_fa33_xor1;
  wire [0:0] u_pg_rca62_and33;
  wire [0:0] u_pg_rca62_or33;
  wire [0:0] u_pg_rca62_pg_fa34_xor0;
  wire [0:0] u_pg_rca62_pg_fa34_and0;
  wire [0:0] u_pg_rca62_pg_fa34_xor1;
  wire [0:0] u_pg_rca62_and34;
  wire [0:0] u_pg_rca62_or34;
  wire [0:0] u_pg_rca62_pg_fa35_xor0;
  wire [0:0] u_pg_rca62_pg_fa35_and0;
  wire [0:0] u_pg_rca62_pg_fa35_xor1;
  wire [0:0] u_pg_rca62_and35;
  wire [0:0] u_pg_rca62_or35;
  wire [0:0] u_pg_rca62_pg_fa36_xor0;
  wire [0:0] u_pg_rca62_pg_fa36_and0;
  wire [0:0] u_pg_rca62_pg_fa36_xor1;
  wire [0:0] u_pg_rca62_and36;
  wire [0:0] u_pg_rca62_or36;
  wire [0:0] u_pg_rca62_pg_fa37_xor0;
  wire [0:0] u_pg_rca62_pg_fa37_and0;
  wire [0:0] u_pg_rca62_pg_fa37_xor1;
  wire [0:0] u_pg_rca62_and37;
  wire [0:0] u_pg_rca62_or37;
  wire [0:0] u_pg_rca62_pg_fa38_xor0;
  wire [0:0] u_pg_rca62_pg_fa38_and0;
  wire [0:0] u_pg_rca62_pg_fa38_xor1;
  wire [0:0] u_pg_rca62_and38;
  wire [0:0] u_pg_rca62_or38;
  wire [0:0] u_pg_rca62_pg_fa39_xor0;
  wire [0:0] u_pg_rca62_pg_fa39_and0;
  wire [0:0] u_pg_rca62_pg_fa39_xor1;
  wire [0:0] u_pg_rca62_and39;
  wire [0:0] u_pg_rca62_or39;
  wire [0:0] u_pg_rca62_pg_fa40_xor0;
  wire [0:0] u_pg_rca62_pg_fa40_and0;
  wire [0:0] u_pg_rca62_pg_fa40_xor1;
  wire [0:0] u_pg_rca62_and40;
  wire [0:0] u_pg_rca62_or40;
  wire [0:0] u_pg_rca62_pg_fa41_xor0;
  wire [0:0] u_pg_rca62_pg_fa41_and0;
  wire [0:0] u_pg_rca62_pg_fa41_xor1;
  wire [0:0] u_pg_rca62_and41;
  wire [0:0] u_pg_rca62_or41;
  wire [0:0] u_pg_rca62_pg_fa42_xor0;
  wire [0:0] u_pg_rca62_pg_fa42_and0;
  wire [0:0] u_pg_rca62_pg_fa42_xor1;
  wire [0:0] u_pg_rca62_and42;
  wire [0:0] u_pg_rca62_or42;
  wire [0:0] u_pg_rca62_pg_fa43_xor0;
  wire [0:0] u_pg_rca62_pg_fa43_and0;
  wire [0:0] u_pg_rca62_pg_fa43_xor1;
  wire [0:0] u_pg_rca62_and43;
  wire [0:0] u_pg_rca62_or43;
  wire [0:0] u_pg_rca62_pg_fa44_xor0;
  wire [0:0] u_pg_rca62_pg_fa44_and0;
  wire [0:0] u_pg_rca62_pg_fa44_xor1;
  wire [0:0] u_pg_rca62_and44;
  wire [0:0] u_pg_rca62_or44;
  wire [0:0] u_pg_rca62_pg_fa45_xor0;
  wire [0:0] u_pg_rca62_pg_fa45_and0;
  wire [0:0] u_pg_rca62_pg_fa45_xor1;
  wire [0:0] u_pg_rca62_and45;
  wire [0:0] u_pg_rca62_or45;
  wire [0:0] u_pg_rca62_pg_fa46_xor0;
  wire [0:0] u_pg_rca62_pg_fa46_and0;
  wire [0:0] u_pg_rca62_pg_fa46_xor1;
  wire [0:0] u_pg_rca62_and46;
  wire [0:0] u_pg_rca62_or46;
  wire [0:0] u_pg_rca62_pg_fa47_xor0;
  wire [0:0] u_pg_rca62_pg_fa47_and0;
  wire [0:0] u_pg_rca62_pg_fa47_xor1;
  wire [0:0] u_pg_rca62_and47;
  wire [0:0] u_pg_rca62_or47;
  wire [0:0] u_pg_rca62_pg_fa48_xor0;
  wire [0:0] u_pg_rca62_pg_fa48_and0;
  wire [0:0] u_pg_rca62_pg_fa48_xor1;
  wire [0:0] u_pg_rca62_and48;
  wire [0:0] u_pg_rca62_or48;
  wire [0:0] u_pg_rca62_pg_fa49_xor0;
  wire [0:0] u_pg_rca62_pg_fa49_and0;
  wire [0:0] u_pg_rca62_pg_fa49_xor1;
  wire [0:0] u_pg_rca62_and49;
  wire [0:0] u_pg_rca62_or49;
  wire [0:0] u_pg_rca62_pg_fa50_xor0;
  wire [0:0] u_pg_rca62_pg_fa50_and0;
  wire [0:0] u_pg_rca62_pg_fa50_xor1;
  wire [0:0] u_pg_rca62_and50;
  wire [0:0] u_pg_rca62_or50;
  wire [0:0] u_pg_rca62_pg_fa51_xor0;
  wire [0:0] u_pg_rca62_pg_fa51_and0;
  wire [0:0] u_pg_rca62_pg_fa51_xor1;
  wire [0:0] u_pg_rca62_and51;
  wire [0:0] u_pg_rca62_or51;
  wire [0:0] u_pg_rca62_pg_fa52_xor0;
  wire [0:0] u_pg_rca62_pg_fa52_and0;
  wire [0:0] u_pg_rca62_pg_fa52_xor1;
  wire [0:0] u_pg_rca62_and52;
  wire [0:0] u_pg_rca62_or52;
  wire [0:0] u_pg_rca62_pg_fa53_xor0;
  wire [0:0] u_pg_rca62_pg_fa53_and0;
  wire [0:0] u_pg_rca62_pg_fa53_xor1;
  wire [0:0] u_pg_rca62_and53;
  wire [0:0] u_pg_rca62_or53;
  wire [0:0] u_pg_rca62_pg_fa54_xor0;
  wire [0:0] u_pg_rca62_pg_fa54_and0;
  wire [0:0] u_pg_rca62_pg_fa54_xor1;
  wire [0:0] u_pg_rca62_and54;
  wire [0:0] u_pg_rca62_or54;
  wire [0:0] u_pg_rca62_pg_fa55_xor0;
  wire [0:0] u_pg_rca62_pg_fa55_and0;
  wire [0:0] u_pg_rca62_pg_fa55_xor1;
  wire [0:0] u_pg_rca62_and55;
  wire [0:0] u_pg_rca62_or55;
  wire [0:0] u_pg_rca62_pg_fa56_xor0;
  wire [0:0] u_pg_rca62_pg_fa56_and0;
  wire [0:0] u_pg_rca62_pg_fa56_xor1;
  wire [0:0] u_pg_rca62_and56;
  wire [0:0] u_pg_rca62_or56;
  wire [0:0] u_pg_rca62_pg_fa57_xor0;
  wire [0:0] u_pg_rca62_pg_fa57_and0;
  wire [0:0] u_pg_rca62_pg_fa57_xor1;
  wire [0:0] u_pg_rca62_and57;
  wire [0:0] u_pg_rca62_or57;
  wire [0:0] u_pg_rca62_pg_fa58_xor0;
  wire [0:0] u_pg_rca62_pg_fa58_and0;
  wire [0:0] u_pg_rca62_pg_fa58_xor1;
  wire [0:0] u_pg_rca62_and58;
  wire [0:0] u_pg_rca62_or58;
  wire [0:0] u_pg_rca62_pg_fa59_xor0;
  wire [0:0] u_pg_rca62_pg_fa59_and0;
  wire [0:0] u_pg_rca62_pg_fa59_xor1;
  wire [0:0] u_pg_rca62_and59;
  wire [0:0] u_pg_rca62_or59;
  wire [0:0] u_pg_rca62_pg_fa60_xor0;
  wire [0:0] u_pg_rca62_pg_fa60_and0;
  wire [0:0] u_pg_rca62_pg_fa60_xor1;
  wire [0:0] u_pg_rca62_and60;
  wire [0:0] u_pg_rca62_or60;
  wire [0:0] u_pg_rca62_pg_fa61_xor0;
  wire [0:0] u_pg_rca62_pg_fa61_and0;
  wire [0:0] u_pg_rca62_pg_fa61_xor1;
  wire [0:0] u_pg_rca62_and61;
  wire [0:0] u_pg_rca62_or61;

  pg_fa pg_fa_u_pg_rca62_pg_fa0_out(a[0], b[0], 1'b0, u_pg_rca62_pg_fa0_xor0, u_pg_rca62_pg_fa0_and0);
  pg_fa pg_fa_u_pg_rca62_pg_fa1_out(a[1], b[1], u_pg_rca62_pg_fa0_and0[0], u_pg_rca62_pg_fa1_xor0, u_pg_rca62_pg_fa1_and0, u_pg_rca62_pg_fa1_xor1);
  and_gate and_gate_u_pg_rca62_and1(u_pg_rca62_pg_fa0_and0[0], u_pg_rca62_pg_fa1_xor0[0], u_pg_rca62_and1);
  or_gate or_gate_u_pg_rca62_or1(u_pg_rca62_and1[0], u_pg_rca62_pg_fa1_and0[0], u_pg_rca62_or1);
  pg_fa pg_fa_u_pg_rca62_pg_fa2_out(a[2], b[2], u_pg_rca62_or1[0], u_pg_rca62_pg_fa2_xor0, u_pg_rca62_pg_fa2_and0, u_pg_rca62_pg_fa2_xor1);
  and_gate and_gate_u_pg_rca62_and2(u_pg_rca62_or1[0], u_pg_rca62_pg_fa2_xor0[0], u_pg_rca62_and2);
  or_gate or_gate_u_pg_rca62_or2(u_pg_rca62_and2[0], u_pg_rca62_pg_fa2_and0[0], u_pg_rca62_or2);
  pg_fa pg_fa_u_pg_rca62_pg_fa3_out(a[3], b[3], u_pg_rca62_or2[0], u_pg_rca62_pg_fa3_xor0, u_pg_rca62_pg_fa3_and0, u_pg_rca62_pg_fa3_xor1);
  and_gate and_gate_u_pg_rca62_and3(u_pg_rca62_or2[0], u_pg_rca62_pg_fa3_xor0[0], u_pg_rca62_and3);
  or_gate or_gate_u_pg_rca62_or3(u_pg_rca62_and3[0], u_pg_rca62_pg_fa3_and0[0], u_pg_rca62_or3);
  pg_fa pg_fa_u_pg_rca62_pg_fa4_out(a[4], b[4], u_pg_rca62_or3[0], u_pg_rca62_pg_fa4_xor0, u_pg_rca62_pg_fa4_and0, u_pg_rca62_pg_fa4_xor1);
  and_gate and_gate_u_pg_rca62_and4(u_pg_rca62_or3[0], u_pg_rca62_pg_fa4_xor0[0], u_pg_rca62_and4);
  or_gate or_gate_u_pg_rca62_or4(u_pg_rca62_and4[0], u_pg_rca62_pg_fa4_and0[0], u_pg_rca62_or4);
  pg_fa pg_fa_u_pg_rca62_pg_fa5_out(a[5], b[5], u_pg_rca62_or4[0], u_pg_rca62_pg_fa5_xor0, u_pg_rca62_pg_fa5_and0, u_pg_rca62_pg_fa5_xor1);
  and_gate and_gate_u_pg_rca62_and5(u_pg_rca62_or4[0], u_pg_rca62_pg_fa5_xor0[0], u_pg_rca62_and5);
  or_gate or_gate_u_pg_rca62_or5(u_pg_rca62_and5[0], u_pg_rca62_pg_fa5_and0[0], u_pg_rca62_or5);
  pg_fa pg_fa_u_pg_rca62_pg_fa6_out(a[6], b[6], u_pg_rca62_or5[0], u_pg_rca62_pg_fa6_xor0, u_pg_rca62_pg_fa6_and0, u_pg_rca62_pg_fa6_xor1);
  and_gate and_gate_u_pg_rca62_and6(u_pg_rca62_or5[0], u_pg_rca62_pg_fa6_xor0[0], u_pg_rca62_and6);
  or_gate or_gate_u_pg_rca62_or6(u_pg_rca62_and6[0], u_pg_rca62_pg_fa6_and0[0], u_pg_rca62_or6);
  pg_fa pg_fa_u_pg_rca62_pg_fa7_out(a[7], b[7], u_pg_rca62_or6[0], u_pg_rca62_pg_fa7_xor0, u_pg_rca62_pg_fa7_and0, u_pg_rca62_pg_fa7_xor1);
  and_gate and_gate_u_pg_rca62_and7(u_pg_rca62_or6[0], u_pg_rca62_pg_fa7_xor0[0], u_pg_rca62_and7);
  or_gate or_gate_u_pg_rca62_or7(u_pg_rca62_and7[0], u_pg_rca62_pg_fa7_and0[0], u_pg_rca62_or7);
  pg_fa pg_fa_u_pg_rca62_pg_fa8_out(a[8], b[8], u_pg_rca62_or7[0], u_pg_rca62_pg_fa8_xor0, u_pg_rca62_pg_fa8_and0, u_pg_rca62_pg_fa8_xor1);
  and_gate and_gate_u_pg_rca62_and8(u_pg_rca62_or7[0], u_pg_rca62_pg_fa8_xor0[0], u_pg_rca62_and8);
  or_gate or_gate_u_pg_rca62_or8(u_pg_rca62_and8[0], u_pg_rca62_pg_fa8_and0[0], u_pg_rca62_or8);
  pg_fa pg_fa_u_pg_rca62_pg_fa9_out(a[9], b[9], u_pg_rca62_or8[0], u_pg_rca62_pg_fa9_xor0, u_pg_rca62_pg_fa9_and0, u_pg_rca62_pg_fa9_xor1);
  and_gate and_gate_u_pg_rca62_and9(u_pg_rca62_or8[0], u_pg_rca62_pg_fa9_xor0[0], u_pg_rca62_and9);
  or_gate or_gate_u_pg_rca62_or9(u_pg_rca62_and9[0], u_pg_rca62_pg_fa9_and0[0], u_pg_rca62_or9);
  pg_fa pg_fa_u_pg_rca62_pg_fa10_out(a[10], b[10], u_pg_rca62_or9[0], u_pg_rca62_pg_fa10_xor0, u_pg_rca62_pg_fa10_and0, u_pg_rca62_pg_fa10_xor1);
  and_gate and_gate_u_pg_rca62_and10(u_pg_rca62_or9[0], u_pg_rca62_pg_fa10_xor0[0], u_pg_rca62_and10);
  or_gate or_gate_u_pg_rca62_or10(u_pg_rca62_and10[0], u_pg_rca62_pg_fa10_and0[0], u_pg_rca62_or10);
  pg_fa pg_fa_u_pg_rca62_pg_fa11_out(a[11], b[11], u_pg_rca62_or10[0], u_pg_rca62_pg_fa11_xor0, u_pg_rca62_pg_fa11_and0, u_pg_rca62_pg_fa11_xor1);
  and_gate and_gate_u_pg_rca62_and11(u_pg_rca62_or10[0], u_pg_rca62_pg_fa11_xor0[0], u_pg_rca62_and11);
  or_gate or_gate_u_pg_rca62_or11(u_pg_rca62_and11[0], u_pg_rca62_pg_fa11_and0[0], u_pg_rca62_or11);
  pg_fa pg_fa_u_pg_rca62_pg_fa12_out(a[12], b[12], u_pg_rca62_or11[0], u_pg_rca62_pg_fa12_xor0, u_pg_rca62_pg_fa12_and0, u_pg_rca62_pg_fa12_xor1);
  and_gate and_gate_u_pg_rca62_and12(u_pg_rca62_or11[0], u_pg_rca62_pg_fa12_xor0[0], u_pg_rca62_and12);
  or_gate or_gate_u_pg_rca62_or12(u_pg_rca62_and12[0], u_pg_rca62_pg_fa12_and0[0], u_pg_rca62_or12);
  pg_fa pg_fa_u_pg_rca62_pg_fa13_out(a[13], b[13], u_pg_rca62_or12[0], u_pg_rca62_pg_fa13_xor0, u_pg_rca62_pg_fa13_and0, u_pg_rca62_pg_fa13_xor1);
  and_gate and_gate_u_pg_rca62_and13(u_pg_rca62_or12[0], u_pg_rca62_pg_fa13_xor0[0], u_pg_rca62_and13);
  or_gate or_gate_u_pg_rca62_or13(u_pg_rca62_and13[0], u_pg_rca62_pg_fa13_and0[0], u_pg_rca62_or13);
  pg_fa pg_fa_u_pg_rca62_pg_fa14_out(a[14], b[14], u_pg_rca62_or13[0], u_pg_rca62_pg_fa14_xor0, u_pg_rca62_pg_fa14_and0, u_pg_rca62_pg_fa14_xor1);
  and_gate and_gate_u_pg_rca62_and14(u_pg_rca62_or13[0], u_pg_rca62_pg_fa14_xor0[0], u_pg_rca62_and14);
  or_gate or_gate_u_pg_rca62_or14(u_pg_rca62_and14[0], u_pg_rca62_pg_fa14_and0[0], u_pg_rca62_or14);
  pg_fa pg_fa_u_pg_rca62_pg_fa15_out(a[15], b[15], u_pg_rca62_or14[0], u_pg_rca62_pg_fa15_xor0, u_pg_rca62_pg_fa15_and0, u_pg_rca62_pg_fa15_xor1);
  and_gate and_gate_u_pg_rca62_and15(u_pg_rca62_or14[0], u_pg_rca62_pg_fa15_xor0[0], u_pg_rca62_and15);
  or_gate or_gate_u_pg_rca62_or15(u_pg_rca62_and15[0], u_pg_rca62_pg_fa15_and0[0], u_pg_rca62_or15);
  pg_fa pg_fa_u_pg_rca62_pg_fa16_out(a[16], b[16], u_pg_rca62_or15[0], u_pg_rca62_pg_fa16_xor0, u_pg_rca62_pg_fa16_and0, u_pg_rca62_pg_fa16_xor1);
  and_gate and_gate_u_pg_rca62_and16(u_pg_rca62_or15[0], u_pg_rca62_pg_fa16_xor0[0], u_pg_rca62_and16);
  or_gate or_gate_u_pg_rca62_or16(u_pg_rca62_and16[0], u_pg_rca62_pg_fa16_and0[0], u_pg_rca62_or16);
  pg_fa pg_fa_u_pg_rca62_pg_fa17_out(a[17], b[17], u_pg_rca62_or16[0], u_pg_rca62_pg_fa17_xor0, u_pg_rca62_pg_fa17_and0, u_pg_rca62_pg_fa17_xor1);
  and_gate and_gate_u_pg_rca62_and17(u_pg_rca62_or16[0], u_pg_rca62_pg_fa17_xor0[0], u_pg_rca62_and17);
  or_gate or_gate_u_pg_rca62_or17(u_pg_rca62_and17[0], u_pg_rca62_pg_fa17_and0[0], u_pg_rca62_or17);
  pg_fa pg_fa_u_pg_rca62_pg_fa18_out(a[18], b[18], u_pg_rca62_or17[0], u_pg_rca62_pg_fa18_xor0, u_pg_rca62_pg_fa18_and0, u_pg_rca62_pg_fa18_xor1);
  and_gate and_gate_u_pg_rca62_and18(u_pg_rca62_or17[0], u_pg_rca62_pg_fa18_xor0[0], u_pg_rca62_and18);
  or_gate or_gate_u_pg_rca62_or18(u_pg_rca62_and18[0], u_pg_rca62_pg_fa18_and0[0], u_pg_rca62_or18);
  pg_fa pg_fa_u_pg_rca62_pg_fa19_out(a[19], b[19], u_pg_rca62_or18[0], u_pg_rca62_pg_fa19_xor0, u_pg_rca62_pg_fa19_and0, u_pg_rca62_pg_fa19_xor1);
  and_gate and_gate_u_pg_rca62_and19(u_pg_rca62_or18[0], u_pg_rca62_pg_fa19_xor0[0], u_pg_rca62_and19);
  or_gate or_gate_u_pg_rca62_or19(u_pg_rca62_and19[0], u_pg_rca62_pg_fa19_and0[0], u_pg_rca62_or19);
  pg_fa pg_fa_u_pg_rca62_pg_fa20_out(a[20], b[20], u_pg_rca62_or19[0], u_pg_rca62_pg_fa20_xor0, u_pg_rca62_pg_fa20_and0, u_pg_rca62_pg_fa20_xor1);
  and_gate and_gate_u_pg_rca62_and20(u_pg_rca62_or19[0], u_pg_rca62_pg_fa20_xor0[0], u_pg_rca62_and20);
  or_gate or_gate_u_pg_rca62_or20(u_pg_rca62_and20[0], u_pg_rca62_pg_fa20_and0[0], u_pg_rca62_or20);
  pg_fa pg_fa_u_pg_rca62_pg_fa21_out(a[21], b[21], u_pg_rca62_or20[0], u_pg_rca62_pg_fa21_xor0, u_pg_rca62_pg_fa21_and0, u_pg_rca62_pg_fa21_xor1);
  and_gate and_gate_u_pg_rca62_and21(u_pg_rca62_or20[0], u_pg_rca62_pg_fa21_xor0[0], u_pg_rca62_and21);
  or_gate or_gate_u_pg_rca62_or21(u_pg_rca62_and21[0], u_pg_rca62_pg_fa21_and0[0], u_pg_rca62_or21);
  pg_fa pg_fa_u_pg_rca62_pg_fa22_out(a[22], b[22], u_pg_rca62_or21[0], u_pg_rca62_pg_fa22_xor0, u_pg_rca62_pg_fa22_and0, u_pg_rca62_pg_fa22_xor1);
  and_gate and_gate_u_pg_rca62_and22(u_pg_rca62_or21[0], u_pg_rca62_pg_fa22_xor0[0], u_pg_rca62_and22);
  or_gate or_gate_u_pg_rca62_or22(u_pg_rca62_and22[0], u_pg_rca62_pg_fa22_and0[0], u_pg_rca62_or22);
  pg_fa pg_fa_u_pg_rca62_pg_fa23_out(a[23], b[23], u_pg_rca62_or22[0], u_pg_rca62_pg_fa23_xor0, u_pg_rca62_pg_fa23_and0, u_pg_rca62_pg_fa23_xor1);
  and_gate and_gate_u_pg_rca62_and23(u_pg_rca62_or22[0], u_pg_rca62_pg_fa23_xor0[0], u_pg_rca62_and23);
  or_gate or_gate_u_pg_rca62_or23(u_pg_rca62_and23[0], u_pg_rca62_pg_fa23_and0[0], u_pg_rca62_or23);
  pg_fa pg_fa_u_pg_rca62_pg_fa24_out(a[24], b[24], u_pg_rca62_or23[0], u_pg_rca62_pg_fa24_xor0, u_pg_rca62_pg_fa24_and0, u_pg_rca62_pg_fa24_xor1);
  and_gate and_gate_u_pg_rca62_and24(u_pg_rca62_or23[0], u_pg_rca62_pg_fa24_xor0[0], u_pg_rca62_and24);
  or_gate or_gate_u_pg_rca62_or24(u_pg_rca62_and24[0], u_pg_rca62_pg_fa24_and0[0], u_pg_rca62_or24);
  pg_fa pg_fa_u_pg_rca62_pg_fa25_out(a[25], b[25], u_pg_rca62_or24[0], u_pg_rca62_pg_fa25_xor0, u_pg_rca62_pg_fa25_and0, u_pg_rca62_pg_fa25_xor1);
  and_gate and_gate_u_pg_rca62_and25(u_pg_rca62_or24[0], u_pg_rca62_pg_fa25_xor0[0], u_pg_rca62_and25);
  or_gate or_gate_u_pg_rca62_or25(u_pg_rca62_and25[0], u_pg_rca62_pg_fa25_and0[0], u_pg_rca62_or25);
  pg_fa pg_fa_u_pg_rca62_pg_fa26_out(a[26], b[26], u_pg_rca62_or25[0], u_pg_rca62_pg_fa26_xor0, u_pg_rca62_pg_fa26_and0, u_pg_rca62_pg_fa26_xor1);
  and_gate and_gate_u_pg_rca62_and26(u_pg_rca62_or25[0], u_pg_rca62_pg_fa26_xor0[0], u_pg_rca62_and26);
  or_gate or_gate_u_pg_rca62_or26(u_pg_rca62_and26[0], u_pg_rca62_pg_fa26_and0[0], u_pg_rca62_or26);
  pg_fa pg_fa_u_pg_rca62_pg_fa27_out(a[27], b[27], u_pg_rca62_or26[0], u_pg_rca62_pg_fa27_xor0, u_pg_rca62_pg_fa27_and0, u_pg_rca62_pg_fa27_xor1);
  and_gate and_gate_u_pg_rca62_and27(u_pg_rca62_or26[0], u_pg_rca62_pg_fa27_xor0[0], u_pg_rca62_and27);
  or_gate or_gate_u_pg_rca62_or27(u_pg_rca62_and27[0], u_pg_rca62_pg_fa27_and0[0], u_pg_rca62_or27);
  pg_fa pg_fa_u_pg_rca62_pg_fa28_out(a[28], b[28], u_pg_rca62_or27[0], u_pg_rca62_pg_fa28_xor0, u_pg_rca62_pg_fa28_and0, u_pg_rca62_pg_fa28_xor1);
  and_gate and_gate_u_pg_rca62_and28(u_pg_rca62_or27[0], u_pg_rca62_pg_fa28_xor0[0], u_pg_rca62_and28);
  or_gate or_gate_u_pg_rca62_or28(u_pg_rca62_and28[0], u_pg_rca62_pg_fa28_and0[0], u_pg_rca62_or28);
  pg_fa pg_fa_u_pg_rca62_pg_fa29_out(a[29], b[29], u_pg_rca62_or28[0], u_pg_rca62_pg_fa29_xor0, u_pg_rca62_pg_fa29_and0, u_pg_rca62_pg_fa29_xor1);
  and_gate and_gate_u_pg_rca62_and29(u_pg_rca62_or28[0], u_pg_rca62_pg_fa29_xor0[0], u_pg_rca62_and29);
  or_gate or_gate_u_pg_rca62_or29(u_pg_rca62_and29[0], u_pg_rca62_pg_fa29_and0[0], u_pg_rca62_or29);
  pg_fa pg_fa_u_pg_rca62_pg_fa30_out(a[30], b[30], u_pg_rca62_or29[0], u_pg_rca62_pg_fa30_xor0, u_pg_rca62_pg_fa30_and0, u_pg_rca62_pg_fa30_xor1);
  and_gate and_gate_u_pg_rca62_and30(u_pg_rca62_or29[0], u_pg_rca62_pg_fa30_xor0[0], u_pg_rca62_and30);
  or_gate or_gate_u_pg_rca62_or30(u_pg_rca62_and30[0], u_pg_rca62_pg_fa30_and0[0], u_pg_rca62_or30);
  pg_fa pg_fa_u_pg_rca62_pg_fa31_out(a[31], b[31], u_pg_rca62_or30[0], u_pg_rca62_pg_fa31_xor0, u_pg_rca62_pg_fa31_and0, u_pg_rca62_pg_fa31_xor1);
  and_gate and_gate_u_pg_rca62_and31(u_pg_rca62_or30[0], u_pg_rca62_pg_fa31_xor0[0], u_pg_rca62_and31);
  or_gate or_gate_u_pg_rca62_or31(u_pg_rca62_and31[0], u_pg_rca62_pg_fa31_and0[0], u_pg_rca62_or31);
  pg_fa pg_fa_u_pg_rca62_pg_fa32_out(a[32], b[32], u_pg_rca62_or31[0], u_pg_rca62_pg_fa32_xor0, u_pg_rca62_pg_fa32_and0, u_pg_rca62_pg_fa32_xor1);
  and_gate and_gate_u_pg_rca62_and32(u_pg_rca62_or31[0], u_pg_rca62_pg_fa32_xor0[0], u_pg_rca62_and32);
  or_gate or_gate_u_pg_rca62_or32(u_pg_rca62_and32[0], u_pg_rca62_pg_fa32_and0[0], u_pg_rca62_or32);
  pg_fa pg_fa_u_pg_rca62_pg_fa33_out(a[33], b[33], u_pg_rca62_or32[0], u_pg_rca62_pg_fa33_xor0, u_pg_rca62_pg_fa33_and0, u_pg_rca62_pg_fa33_xor1);
  and_gate and_gate_u_pg_rca62_and33(u_pg_rca62_or32[0], u_pg_rca62_pg_fa33_xor0[0], u_pg_rca62_and33);
  or_gate or_gate_u_pg_rca62_or33(u_pg_rca62_and33[0], u_pg_rca62_pg_fa33_and0[0], u_pg_rca62_or33);
  pg_fa pg_fa_u_pg_rca62_pg_fa34_out(a[34], b[34], u_pg_rca62_or33[0], u_pg_rca62_pg_fa34_xor0, u_pg_rca62_pg_fa34_and0, u_pg_rca62_pg_fa34_xor1);
  and_gate and_gate_u_pg_rca62_and34(u_pg_rca62_or33[0], u_pg_rca62_pg_fa34_xor0[0], u_pg_rca62_and34);
  or_gate or_gate_u_pg_rca62_or34(u_pg_rca62_and34[0], u_pg_rca62_pg_fa34_and0[0], u_pg_rca62_or34);
  pg_fa pg_fa_u_pg_rca62_pg_fa35_out(a[35], b[35], u_pg_rca62_or34[0], u_pg_rca62_pg_fa35_xor0, u_pg_rca62_pg_fa35_and0, u_pg_rca62_pg_fa35_xor1);
  and_gate and_gate_u_pg_rca62_and35(u_pg_rca62_or34[0], u_pg_rca62_pg_fa35_xor0[0], u_pg_rca62_and35);
  or_gate or_gate_u_pg_rca62_or35(u_pg_rca62_and35[0], u_pg_rca62_pg_fa35_and0[0], u_pg_rca62_or35);
  pg_fa pg_fa_u_pg_rca62_pg_fa36_out(a[36], b[36], u_pg_rca62_or35[0], u_pg_rca62_pg_fa36_xor0, u_pg_rca62_pg_fa36_and0, u_pg_rca62_pg_fa36_xor1);
  and_gate and_gate_u_pg_rca62_and36(u_pg_rca62_or35[0], u_pg_rca62_pg_fa36_xor0[0], u_pg_rca62_and36);
  or_gate or_gate_u_pg_rca62_or36(u_pg_rca62_and36[0], u_pg_rca62_pg_fa36_and0[0], u_pg_rca62_or36);
  pg_fa pg_fa_u_pg_rca62_pg_fa37_out(a[37], b[37], u_pg_rca62_or36[0], u_pg_rca62_pg_fa37_xor0, u_pg_rca62_pg_fa37_and0, u_pg_rca62_pg_fa37_xor1);
  and_gate and_gate_u_pg_rca62_and37(u_pg_rca62_or36[0], u_pg_rca62_pg_fa37_xor0[0], u_pg_rca62_and37);
  or_gate or_gate_u_pg_rca62_or37(u_pg_rca62_and37[0], u_pg_rca62_pg_fa37_and0[0], u_pg_rca62_or37);
  pg_fa pg_fa_u_pg_rca62_pg_fa38_out(a[38], b[38], u_pg_rca62_or37[0], u_pg_rca62_pg_fa38_xor0, u_pg_rca62_pg_fa38_and0, u_pg_rca62_pg_fa38_xor1);
  and_gate and_gate_u_pg_rca62_and38(u_pg_rca62_or37[0], u_pg_rca62_pg_fa38_xor0[0], u_pg_rca62_and38);
  or_gate or_gate_u_pg_rca62_or38(u_pg_rca62_and38[0], u_pg_rca62_pg_fa38_and0[0], u_pg_rca62_or38);
  pg_fa pg_fa_u_pg_rca62_pg_fa39_out(a[39], b[39], u_pg_rca62_or38[0], u_pg_rca62_pg_fa39_xor0, u_pg_rca62_pg_fa39_and0, u_pg_rca62_pg_fa39_xor1);
  and_gate and_gate_u_pg_rca62_and39(u_pg_rca62_or38[0], u_pg_rca62_pg_fa39_xor0[0], u_pg_rca62_and39);
  or_gate or_gate_u_pg_rca62_or39(u_pg_rca62_and39[0], u_pg_rca62_pg_fa39_and0[0], u_pg_rca62_or39);
  pg_fa pg_fa_u_pg_rca62_pg_fa40_out(a[40], b[40], u_pg_rca62_or39[0], u_pg_rca62_pg_fa40_xor0, u_pg_rca62_pg_fa40_and0, u_pg_rca62_pg_fa40_xor1);
  and_gate and_gate_u_pg_rca62_and40(u_pg_rca62_or39[0], u_pg_rca62_pg_fa40_xor0[0], u_pg_rca62_and40);
  or_gate or_gate_u_pg_rca62_or40(u_pg_rca62_and40[0], u_pg_rca62_pg_fa40_and0[0], u_pg_rca62_or40);
  pg_fa pg_fa_u_pg_rca62_pg_fa41_out(a[41], b[41], u_pg_rca62_or40[0], u_pg_rca62_pg_fa41_xor0, u_pg_rca62_pg_fa41_and0, u_pg_rca62_pg_fa41_xor1);
  and_gate and_gate_u_pg_rca62_and41(u_pg_rca62_or40[0], u_pg_rca62_pg_fa41_xor0[0], u_pg_rca62_and41);
  or_gate or_gate_u_pg_rca62_or41(u_pg_rca62_and41[0], u_pg_rca62_pg_fa41_and0[0], u_pg_rca62_or41);
  pg_fa pg_fa_u_pg_rca62_pg_fa42_out(a[42], b[42], u_pg_rca62_or41[0], u_pg_rca62_pg_fa42_xor0, u_pg_rca62_pg_fa42_and0, u_pg_rca62_pg_fa42_xor1);
  and_gate and_gate_u_pg_rca62_and42(u_pg_rca62_or41[0], u_pg_rca62_pg_fa42_xor0[0], u_pg_rca62_and42);
  or_gate or_gate_u_pg_rca62_or42(u_pg_rca62_and42[0], u_pg_rca62_pg_fa42_and0[0], u_pg_rca62_or42);
  pg_fa pg_fa_u_pg_rca62_pg_fa43_out(a[43], b[43], u_pg_rca62_or42[0], u_pg_rca62_pg_fa43_xor0, u_pg_rca62_pg_fa43_and0, u_pg_rca62_pg_fa43_xor1);
  and_gate and_gate_u_pg_rca62_and43(u_pg_rca62_or42[0], u_pg_rca62_pg_fa43_xor0[0], u_pg_rca62_and43);
  or_gate or_gate_u_pg_rca62_or43(u_pg_rca62_and43[0], u_pg_rca62_pg_fa43_and0[0], u_pg_rca62_or43);
  pg_fa pg_fa_u_pg_rca62_pg_fa44_out(a[44], b[44], u_pg_rca62_or43[0], u_pg_rca62_pg_fa44_xor0, u_pg_rca62_pg_fa44_and0, u_pg_rca62_pg_fa44_xor1);
  and_gate and_gate_u_pg_rca62_and44(u_pg_rca62_or43[0], u_pg_rca62_pg_fa44_xor0[0], u_pg_rca62_and44);
  or_gate or_gate_u_pg_rca62_or44(u_pg_rca62_and44[0], u_pg_rca62_pg_fa44_and0[0], u_pg_rca62_or44);
  pg_fa pg_fa_u_pg_rca62_pg_fa45_out(a[45], b[45], u_pg_rca62_or44[0], u_pg_rca62_pg_fa45_xor0, u_pg_rca62_pg_fa45_and0, u_pg_rca62_pg_fa45_xor1);
  and_gate and_gate_u_pg_rca62_and45(u_pg_rca62_or44[0], u_pg_rca62_pg_fa45_xor0[0], u_pg_rca62_and45);
  or_gate or_gate_u_pg_rca62_or45(u_pg_rca62_and45[0], u_pg_rca62_pg_fa45_and0[0], u_pg_rca62_or45);
  pg_fa pg_fa_u_pg_rca62_pg_fa46_out(a[46], b[46], u_pg_rca62_or45[0], u_pg_rca62_pg_fa46_xor0, u_pg_rca62_pg_fa46_and0, u_pg_rca62_pg_fa46_xor1);
  and_gate and_gate_u_pg_rca62_and46(u_pg_rca62_or45[0], u_pg_rca62_pg_fa46_xor0[0], u_pg_rca62_and46);
  or_gate or_gate_u_pg_rca62_or46(u_pg_rca62_and46[0], u_pg_rca62_pg_fa46_and0[0], u_pg_rca62_or46);
  pg_fa pg_fa_u_pg_rca62_pg_fa47_out(a[47], b[47], u_pg_rca62_or46[0], u_pg_rca62_pg_fa47_xor0, u_pg_rca62_pg_fa47_and0, u_pg_rca62_pg_fa47_xor1);
  and_gate and_gate_u_pg_rca62_and47(u_pg_rca62_or46[0], u_pg_rca62_pg_fa47_xor0[0], u_pg_rca62_and47);
  or_gate or_gate_u_pg_rca62_or47(u_pg_rca62_and47[0], u_pg_rca62_pg_fa47_and0[0], u_pg_rca62_or47);
  pg_fa pg_fa_u_pg_rca62_pg_fa48_out(a[48], b[48], u_pg_rca62_or47[0], u_pg_rca62_pg_fa48_xor0, u_pg_rca62_pg_fa48_and0, u_pg_rca62_pg_fa48_xor1);
  and_gate and_gate_u_pg_rca62_and48(u_pg_rca62_or47[0], u_pg_rca62_pg_fa48_xor0[0], u_pg_rca62_and48);
  or_gate or_gate_u_pg_rca62_or48(u_pg_rca62_and48[0], u_pg_rca62_pg_fa48_and0[0], u_pg_rca62_or48);
  pg_fa pg_fa_u_pg_rca62_pg_fa49_out(a[49], b[49], u_pg_rca62_or48[0], u_pg_rca62_pg_fa49_xor0, u_pg_rca62_pg_fa49_and0, u_pg_rca62_pg_fa49_xor1);
  and_gate and_gate_u_pg_rca62_and49(u_pg_rca62_or48[0], u_pg_rca62_pg_fa49_xor0[0], u_pg_rca62_and49);
  or_gate or_gate_u_pg_rca62_or49(u_pg_rca62_and49[0], u_pg_rca62_pg_fa49_and0[0], u_pg_rca62_or49);
  pg_fa pg_fa_u_pg_rca62_pg_fa50_out(a[50], b[50], u_pg_rca62_or49[0], u_pg_rca62_pg_fa50_xor0, u_pg_rca62_pg_fa50_and0, u_pg_rca62_pg_fa50_xor1);
  and_gate and_gate_u_pg_rca62_and50(u_pg_rca62_or49[0], u_pg_rca62_pg_fa50_xor0[0], u_pg_rca62_and50);
  or_gate or_gate_u_pg_rca62_or50(u_pg_rca62_and50[0], u_pg_rca62_pg_fa50_and0[0], u_pg_rca62_or50);
  pg_fa pg_fa_u_pg_rca62_pg_fa51_out(a[51], b[51], u_pg_rca62_or50[0], u_pg_rca62_pg_fa51_xor0, u_pg_rca62_pg_fa51_and0, u_pg_rca62_pg_fa51_xor1);
  and_gate and_gate_u_pg_rca62_and51(u_pg_rca62_or50[0], u_pg_rca62_pg_fa51_xor0[0], u_pg_rca62_and51);
  or_gate or_gate_u_pg_rca62_or51(u_pg_rca62_and51[0], u_pg_rca62_pg_fa51_and0[0], u_pg_rca62_or51);
  pg_fa pg_fa_u_pg_rca62_pg_fa52_out(a[52], b[52], u_pg_rca62_or51[0], u_pg_rca62_pg_fa52_xor0, u_pg_rca62_pg_fa52_and0, u_pg_rca62_pg_fa52_xor1);
  and_gate and_gate_u_pg_rca62_and52(u_pg_rca62_or51[0], u_pg_rca62_pg_fa52_xor0[0], u_pg_rca62_and52);
  or_gate or_gate_u_pg_rca62_or52(u_pg_rca62_and52[0], u_pg_rca62_pg_fa52_and0[0], u_pg_rca62_or52);
  pg_fa pg_fa_u_pg_rca62_pg_fa53_out(a[53], b[53], u_pg_rca62_or52[0], u_pg_rca62_pg_fa53_xor0, u_pg_rca62_pg_fa53_and0, u_pg_rca62_pg_fa53_xor1);
  and_gate and_gate_u_pg_rca62_and53(u_pg_rca62_or52[0], u_pg_rca62_pg_fa53_xor0[0], u_pg_rca62_and53);
  or_gate or_gate_u_pg_rca62_or53(u_pg_rca62_and53[0], u_pg_rca62_pg_fa53_and0[0], u_pg_rca62_or53);
  pg_fa pg_fa_u_pg_rca62_pg_fa54_out(a[54], b[54], u_pg_rca62_or53[0], u_pg_rca62_pg_fa54_xor0, u_pg_rca62_pg_fa54_and0, u_pg_rca62_pg_fa54_xor1);
  and_gate and_gate_u_pg_rca62_and54(u_pg_rca62_or53[0], u_pg_rca62_pg_fa54_xor0[0], u_pg_rca62_and54);
  or_gate or_gate_u_pg_rca62_or54(u_pg_rca62_and54[0], u_pg_rca62_pg_fa54_and0[0], u_pg_rca62_or54);
  pg_fa pg_fa_u_pg_rca62_pg_fa55_out(a[55], b[55], u_pg_rca62_or54[0], u_pg_rca62_pg_fa55_xor0, u_pg_rca62_pg_fa55_and0, u_pg_rca62_pg_fa55_xor1);
  and_gate and_gate_u_pg_rca62_and55(u_pg_rca62_or54[0], u_pg_rca62_pg_fa55_xor0[0], u_pg_rca62_and55);
  or_gate or_gate_u_pg_rca62_or55(u_pg_rca62_and55[0], u_pg_rca62_pg_fa55_and0[0], u_pg_rca62_or55);
  pg_fa pg_fa_u_pg_rca62_pg_fa56_out(a[56], b[56], u_pg_rca62_or55[0], u_pg_rca62_pg_fa56_xor0, u_pg_rca62_pg_fa56_and0, u_pg_rca62_pg_fa56_xor1);
  and_gate and_gate_u_pg_rca62_and56(u_pg_rca62_or55[0], u_pg_rca62_pg_fa56_xor0[0], u_pg_rca62_and56);
  or_gate or_gate_u_pg_rca62_or56(u_pg_rca62_and56[0], u_pg_rca62_pg_fa56_and0[0], u_pg_rca62_or56);
  pg_fa pg_fa_u_pg_rca62_pg_fa57_out(a[57], b[57], u_pg_rca62_or56[0], u_pg_rca62_pg_fa57_xor0, u_pg_rca62_pg_fa57_and0, u_pg_rca62_pg_fa57_xor1);
  and_gate and_gate_u_pg_rca62_and57(u_pg_rca62_or56[0], u_pg_rca62_pg_fa57_xor0[0], u_pg_rca62_and57);
  or_gate or_gate_u_pg_rca62_or57(u_pg_rca62_and57[0], u_pg_rca62_pg_fa57_and0[0], u_pg_rca62_or57);
  pg_fa pg_fa_u_pg_rca62_pg_fa58_out(a[58], b[58], u_pg_rca62_or57[0], u_pg_rca62_pg_fa58_xor0, u_pg_rca62_pg_fa58_and0, u_pg_rca62_pg_fa58_xor1);
  and_gate and_gate_u_pg_rca62_and58(u_pg_rca62_or57[0], u_pg_rca62_pg_fa58_xor0[0], u_pg_rca62_and58);
  or_gate or_gate_u_pg_rca62_or58(u_pg_rca62_and58[0], u_pg_rca62_pg_fa58_and0[0], u_pg_rca62_or58);
  pg_fa pg_fa_u_pg_rca62_pg_fa59_out(a[59], b[59], u_pg_rca62_or58[0], u_pg_rca62_pg_fa59_xor0, u_pg_rca62_pg_fa59_and0, u_pg_rca62_pg_fa59_xor1);
  and_gate and_gate_u_pg_rca62_and59(u_pg_rca62_or58[0], u_pg_rca62_pg_fa59_xor0[0], u_pg_rca62_and59);
  or_gate or_gate_u_pg_rca62_or59(u_pg_rca62_and59[0], u_pg_rca62_pg_fa59_and0[0], u_pg_rca62_or59);
  pg_fa pg_fa_u_pg_rca62_pg_fa60_out(a[60], b[60], u_pg_rca62_or59[0], u_pg_rca62_pg_fa60_xor0, u_pg_rca62_pg_fa60_and0, u_pg_rca62_pg_fa60_xor1);
  and_gate and_gate_u_pg_rca62_and60(u_pg_rca62_or59[0], u_pg_rca62_pg_fa60_xor0[0], u_pg_rca62_and60);
  or_gate or_gate_u_pg_rca62_or60(u_pg_rca62_and60[0], u_pg_rca62_pg_fa60_and0[0], u_pg_rca62_or60);
  pg_fa pg_fa_u_pg_rca62_pg_fa61_out(a[61], b[61], u_pg_rca62_or60[0], u_pg_rca62_pg_fa61_xor0, u_pg_rca62_pg_fa61_and0, u_pg_rca62_pg_fa61_xor1);
  and_gate and_gate_u_pg_rca62_and61(u_pg_rca62_or60[0], u_pg_rca62_pg_fa61_xor0[0], u_pg_rca62_and61);
  or_gate or_gate_u_pg_rca62_or61(u_pg_rca62_and61[0], u_pg_rca62_pg_fa61_and0[0], u_pg_rca62_or61);

  assign u_pg_rca62_out[0] = u_pg_rca62_pg_fa0_xor0[0];
  assign u_pg_rca62_out[1] = u_pg_rca62_pg_fa1_xor1[0];
  assign u_pg_rca62_out[2] = u_pg_rca62_pg_fa2_xor1[0];
  assign u_pg_rca62_out[3] = u_pg_rca62_pg_fa3_xor1[0];
  assign u_pg_rca62_out[4] = u_pg_rca62_pg_fa4_xor1[0];
  assign u_pg_rca62_out[5] = u_pg_rca62_pg_fa5_xor1[0];
  assign u_pg_rca62_out[6] = u_pg_rca62_pg_fa6_xor1[0];
  assign u_pg_rca62_out[7] = u_pg_rca62_pg_fa7_xor1[0];
  assign u_pg_rca62_out[8] = u_pg_rca62_pg_fa8_xor1[0];
  assign u_pg_rca62_out[9] = u_pg_rca62_pg_fa9_xor1[0];
  assign u_pg_rca62_out[10] = u_pg_rca62_pg_fa10_xor1[0];
  assign u_pg_rca62_out[11] = u_pg_rca62_pg_fa11_xor1[0];
  assign u_pg_rca62_out[12] = u_pg_rca62_pg_fa12_xor1[0];
  assign u_pg_rca62_out[13] = u_pg_rca62_pg_fa13_xor1[0];
  assign u_pg_rca62_out[14] = u_pg_rca62_pg_fa14_xor1[0];
  assign u_pg_rca62_out[15] = u_pg_rca62_pg_fa15_xor1[0];
  assign u_pg_rca62_out[16] = u_pg_rca62_pg_fa16_xor1[0];
  assign u_pg_rca62_out[17] = u_pg_rca62_pg_fa17_xor1[0];
  assign u_pg_rca62_out[18] = u_pg_rca62_pg_fa18_xor1[0];
  assign u_pg_rca62_out[19] = u_pg_rca62_pg_fa19_xor1[0];
  assign u_pg_rca62_out[20] = u_pg_rca62_pg_fa20_xor1[0];
  assign u_pg_rca62_out[21] = u_pg_rca62_pg_fa21_xor1[0];
  assign u_pg_rca62_out[22] = u_pg_rca62_pg_fa22_xor1[0];
  assign u_pg_rca62_out[23] = u_pg_rca62_pg_fa23_xor1[0];
  assign u_pg_rca62_out[24] = u_pg_rca62_pg_fa24_xor1[0];
  assign u_pg_rca62_out[25] = u_pg_rca62_pg_fa25_xor1[0];
  assign u_pg_rca62_out[26] = u_pg_rca62_pg_fa26_xor1[0];
  assign u_pg_rca62_out[27] = u_pg_rca62_pg_fa27_xor1[0];
  assign u_pg_rca62_out[28] = u_pg_rca62_pg_fa28_xor1[0];
  assign u_pg_rca62_out[29] = u_pg_rca62_pg_fa29_xor1[0];
  assign u_pg_rca62_out[30] = u_pg_rca62_pg_fa30_xor1[0];
  assign u_pg_rca62_out[31] = u_pg_rca62_pg_fa31_xor1[0];
  assign u_pg_rca62_out[32] = u_pg_rca62_pg_fa32_xor1[0];
  assign u_pg_rca62_out[33] = u_pg_rca62_pg_fa33_xor1[0];
  assign u_pg_rca62_out[34] = u_pg_rca62_pg_fa34_xor1[0];
  assign u_pg_rca62_out[35] = u_pg_rca62_pg_fa35_xor1[0];
  assign u_pg_rca62_out[36] = u_pg_rca62_pg_fa36_xor1[0];
  assign u_pg_rca62_out[37] = u_pg_rca62_pg_fa37_xor1[0];
  assign u_pg_rca62_out[38] = u_pg_rca62_pg_fa38_xor1[0];
  assign u_pg_rca62_out[39] = u_pg_rca62_pg_fa39_xor1[0];
  assign u_pg_rca62_out[40] = u_pg_rca62_pg_fa40_xor1[0];
  assign u_pg_rca62_out[41] = u_pg_rca62_pg_fa41_xor1[0];
  assign u_pg_rca62_out[42] = u_pg_rca62_pg_fa42_xor1[0];
  assign u_pg_rca62_out[43] = u_pg_rca62_pg_fa43_xor1[0];
  assign u_pg_rca62_out[44] = u_pg_rca62_pg_fa44_xor1[0];
  assign u_pg_rca62_out[45] = u_pg_rca62_pg_fa45_xor1[0];
  assign u_pg_rca62_out[46] = u_pg_rca62_pg_fa46_xor1[0];
  assign u_pg_rca62_out[47] = u_pg_rca62_pg_fa47_xor1[0];
  assign u_pg_rca62_out[48] = u_pg_rca62_pg_fa48_xor1[0];
  assign u_pg_rca62_out[49] = u_pg_rca62_pg_fa49_xor1[0];
  assign u_pg_rca62_out[50] = u_pg_rca62_pg_fa50_xor1[0];
  assign u_pg_rca62_out[51] = u_pg_rca62_pg_fa51_xor1[0];
  assign u_pg_rca62_out[52] = u_pg_rca62_pg_fa52_xor1[0];
  assign u_pg_rca62_out[53] = u_pg_rca62_pg_fa53_xor1[0];
  assign u_pg_rca62_out[54] = u_pg_rca62_pg_fa54_xor1[0];
  assign u_pg_rca62_out[55] = u_pg_rca62_pg_fa55_xor1[0];
  assign u_pg_rca62_out[56] = u_pg_rca62_pg_fa56_xor1[0];
  assign u_pg_rca62_out[57] = u_pg_rca62_pg_fa57_xor1[0];
  assign u_pg_rca62_out[58] = u_pg_rca62_pg_fa58_xor1[0];
  assign u_pg_rca62_out[59] = u_pg_rca62_pg_fa59_xor1[0];
  assign u_pg_rca62_out[60] = u_pg_rca62_pg_fa60_xor1[0];
  assign u_pg_rca62_out[61] = u_pg_rca62_pg_fa61_xor1[0];
  assign u_pg_rca62_out[62] = u_pg_rca62_or61[0];
endmodule

module h_s_dadda_pg_rca32(input [31:0] a, input [31:0] b, output [63:0] h_s_dadda_pg_rca32_out);
  wire [0:0] h_s_dadda_pg_rca32_and_28_0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_1;
  wire [0:0] h_s_dadda_pg_rca32_ha0_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha0_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_1;
  wire [0:0] h_s_dadda_pg_rca32_fa0_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa0_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_2;
  wire [0:0] h_s_dadda_pg_rca32_and_26_3;
  wire [0:0] h_s_dadda_pg_rca32_ha1_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha1_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_0;
  wire [0:0] h_s_dadda_pg_rca32_fa1_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa1_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_1;
  wire [0:0] h_s_dadda_pg_rca32_and_28_2;
  wire [0:0] h_s_dadda_pg_rca32_and_27_3;
  wire [0:0] h_s_dadda_pg_rca32_fa2_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa2_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_4;
  wire [0:0] h_s_dadda_pg_rca32_and_25_5;
  wire [0:0] h_s_dadda_pg_rca32_ha2_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha2_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa3_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa3_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_1;
  wire [0:0] h_s_dadda_pg_rca32_and_29_2;
  wire [0:0] h_s_dadda_pg_rca32_fa4_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa4_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_3;
  wire [0:0] h_s_dadda_pg_rca32_and_27_4;
  wire [0:0] h_s_dadda_pg_rca32_and_26_5;
  wire [0:0] h_s_dadda_pg_rca32_fa5_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa5_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_6;
  wire [0:0] h_s_dadda_pg_rca32_and_24_7;
  wire [0:0] h_s_dadda_pg_rca32_ha3_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha3_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa6_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa6_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_1;
  wire [0:0] h_s_dadda_pg_rca32_fa7_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa7_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_2;
  wire [0:0] h_s_dadda_pg_rca32_and_29_3;
  wire [0:0] h_s_dadda_pg_rca32_and_28_4;
  wire [0:0] h_s_dadda_pg_rca32_fa8_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa8_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_5;
  wire [0:0] h_s_dadda_pg_rca32_and_26_6;
  wire [0:0] h_s_dadda_pg_rca32_and_25_7;
  wire [0:0] h_s_dadda_pg_rca32_fa9_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa9_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa10_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa10_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_2;
  wire [0:0] h_s_dadda_pg_rca32_and_30_3;
  wire [0:0] h_s_dadda_pg_rca32_fa11_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa11_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_4;
  wire [0:0] h_s_dadda_pg_rca32_and_28_5;
  wire [0:0] h_s_dadda_pg_rca32_and_27_6;
  wire [0:0] h_s_dadda_pg_rca32_fa12_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa12_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa13_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa13_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_3;
  wire [0:0] h_s_dadda_pg_rca32_and_30_4;
  wire [0:0] h_s_dadda_pg_rca32_and_29_5;
  wire [0:0] h_s_dadda_pg_rca32_fa14_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa14_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_4;
  wire [0:0] h_s_dadda_pg_rca32_fa15_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa15_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_1;
  wire [0:0] h_s_dadda_pg_rca32_ha4_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha4_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_1;
  wire [0:0] h_s_dadda_pg_rca32_fa16_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa16_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_2;
  wire [0:0] h_s_dadda_pg_rca32_and_4_3;
  wire [0:0] h_s_dadda_pg_rca32_ha5_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha5_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_0;
  wire [0:0] h_s_dadda_pg_rca32_fa17_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa17_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_1;
  wire [0:0] h_s_dadda_pg_rca32_and_6_2;
  wire [0:0] h_s_dadda_pg_rca32_and_5_3;
  wire [0:0] h_s_dadda_pg_rca32_fa18_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa18_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_4;
  wire [0:0] h_s_dadda_pg_rca32_and_3_5;
  wire [0:0] h_s_dadda_pg_rca32_ha6_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha6_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa19_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa19_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_1;
  wire [0:0] h_s_dadda_pg_rca32_and_7_2;
  wire [0:0] h_s_dadda_pg_rca32_fa20_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa20_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_3;
  wire [0:0] h_s_dadda_pg_rca32_and_5_4;
  wire [0:0] h_s_dadda_pg_rca32_and_4_5;
  wire [0:0] h_s_dadda_pg_rca32_fa21_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa21_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_6;
  wire [0:0] h_s_dadda_pg_rca32_and_2_7;
  wire [0:0] h_s_dadda_pg_rca32_ha7_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha7_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa22_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa22_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_1;
  wire [0:0] h_s_dadda_pg_rca32_fa23_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa23_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_2;
  wire [0:0] h_s_dadda_pg_rca32_and_7_3;
  wire [0:0] h_s_dadda_pg_rca32_and_6_4;
  wire [0:0] h_s_dadda_pg_rca32_fa24_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa24_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_5;
  wire [0:0] h_s_dadda_pg_rca32_and_4_6;
  wire [0:0] h_s_dadda_pg_rca32_and_3_7;
  wire [0:0] h_s_dadda_pg_rca32_fa25_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa25_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_8;
  wire [0:0] h_s_dadda_pg_rca32_and_1_9;
  wire [0:0] h_s_dadda_pg_rca32_ha8_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha8_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa26_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa26_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_0;
  wire [0:0] h_s_dadda_pg_rca32_fa27_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa27_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_1;
  wire [0:0] h_s_dadda_pg_rca32_and_9_2;
  wire [0:0] h_s_dadda_pg_rca32_and_8_3;
  wire [0:0] h_s_dadda_pg_rca32_fa28_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa28_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_4;
  wire [0:0] h_s_dadda_pg_rca32_and_6_5;
  wire [0:0] h_s_dadda_pg_rca32_and_5_6;
  wire [0:0] h_s_dadda_pg_rca32_fa29_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa29_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_7;
  wire [0:0] h_s_dadda_pg_rca32_and_3_8;
  wire [0:0] h_s_dadda_pg_rca32_and_2_9;
  wire [0:0] h_s_dadda_pg_rca32_fa30_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa30_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_10;
  wire [0:0] h_s_dadda_pg_rca32_and_0_11;
  wire [0:0] h_s_dadda_pg_rca32_ha9_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha9_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa31_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa31_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa32_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa32_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_1;
  wire [0:0] h_s_dadda_pg_rca32_and_10_2;
  wire [0:0] h_s_dadda_pg_rca32_fa33_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa33_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_3;
  wire [0:0] h_s_dadda_pg_rca32_and_8_4;
  wire [0:0] h_s_dadda_pg_rca32_and_7_5;
  wire [0:0] h_s_dadda_pg_rca32_fa34_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa34_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_6;
  wire [0:0] h_s_dadda_pg_rca32_and_5_7;
  wire [0:0] h_s_dadda_pg_rca32_and_4_8;
  wire [0:0] h_s_dadda_pg_rca32_fa35_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa35_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_9;
  wire [0:0] h_s_dadda_pg_rca32_and_2_10;
  wire [0:0] h_s_dadda_pg_rca32_and_1_11;
  wire [0:0] h_s_dadda_pg_rca32_fa36_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa36_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_12;
  wire [0:0] h_s_dadda_pg_rca32_ha10_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha10_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa37_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa37_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa38_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa38_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_1;
  wire [0:0] h_s_dadda_pg_rca32_fa39_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa39_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_2;
  wire [0:0] h_s_dadda_pg_rca32_and_10_3;
  wire [0:0] h_s_dadda_pg_rca32_and_9_4;
  wire [0:0] h_s_dadda_pg_rca32_fa40_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa40_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_5;
  wire [0:0] h_s_dadda_pg_rca32_and_7_6;
  wire [0:0] h_s_dadda_pg_rca32_and_6_7;
  wire [0:0] h_s_dadda_pg_rca32_fa41_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa41_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_8;
  wire [0:0] h_s_dadda_pg_rca32_and_4_9;
  wire [0:0] h_s_dadda_pg_rca32_and_3_10;
  wire [0:0] h_s_dadda_pg_rca32_fa42_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa42_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_11;
  wire [0:0] h_s_dadda_pg_rca32_and_1_12;
  wire [0:0] h_s_dadda_pg_rca32_and_0_13;
  wire [0:0] h_s_dadda_pg_rca32_fa43_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa43_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha11_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha11_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa44_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa44_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa45_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa45_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_0;
  wire [0:0] h_s_dadda_pg_rca32_fa46_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa46_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_1;
  wire [0:0] h_s_dadda_pg_rca32_and_12_2;
  wire [0:0] h_s_dadda_pg_rca32_and_11_3;
  wire [0:0] h_s_dadda_pg_rca32_fa47_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa47_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_4;
  wire [0:0] h_s_dadda_pg_rca32_and_9_5;
  wire [0:0] h_s_dadda_pg_rca32_and_8_6;
  wire [0:0] h_s_dadda_pg_rca32_fa48_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa48_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_7;
  wire [0:0] h_s_dadda_pg_rca32_and_6_8;
  wire [0:0] h_s_dadda_pg_rca32_and_5_9;
  wire [0:0] h_s_dadda_pg_rca32_fa49_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa49_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_10;
  wire [0:0] h_s_dadda_pg_rca32_and_3_11;
  wire [0:0] h_s_dadda_pg_rca32_and_2_12;
  wire [0:0] h_s_dadda_pg_rca32_fa50_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa50_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_13;
  wire [0:0] h_s_dadda_pg_rca32_and_0_14;
  wire [0:0] h_s_dadda_pg_rca32_fa51_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa51_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha12_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha12_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa52_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa52_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa53_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa53_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa54_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa54_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_1;
  wire [0:0] h_s_dadda_pg_rca32_and_13_2;
  wire [0:0] h_s_dadda_pg_rca32_fa55_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa55_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_3;
  wire [0:0] h_s_dadda_pg_rca32_and_11_4;
  wire [0:0] h_s_dadda_pg_rca32_and_10_5;
  wire [0:0] h_s_dadda_pg_rca32_fa56_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa56_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_6;
  wire [0:0] h_s_dadda_pg_rca32_and_8_7;
  wire [0:0] h_s_dadda_pg_rca32_and_7_8;
  wire [0:0] h_s_dadda_pg_rca32_fa57_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa57_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_9;
  wire [0:0] h_s_dadda_pg_rca32_and_5_10;
  wire [0:0] h_s_dadda_pg_rca32_and_4_11;
  wire [0:0] h_s_dadda_pg_rca32_fa58_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa58_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_12;
  wire [0:0] h_s_dadda_pg_rca32_and_2_13;
  wire [0:0] h_s_dadda_pg_rca32_and_1_14;
  wire [0:0] h_s_dadda_pg_rca32_fa59_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa59_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_15;
  wire [0:0] h_s_dadda_pg_rca32_fa60_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa60_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha13_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha13_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa61_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa61_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa62_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa62_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa63_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa63_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_1;
  wire [0:0] h_s_dadda_pg_rca32_fa64_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa64_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_2;
  wire [0:0] h_s_dadda_pg_rca32_and_13_3;
  wire [0:0] h_s_dadda_pg_rca32_and_12_4;
  wire [0:0] h_s_dadda_pg_rca32_fa65_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa65_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_5;
  wire [0:0] h_s_dadda_pg_rca32_and_10_6;
  wire [0:0] h_s_dadda_pg_rca32_and_9_7;
  wire [0:0] h_s_dadda_pg_rca32_fa66_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa66_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_8;
  wire [0:0] h_s_dadda_pg_rca32_and_7_9;
  wire [0:0] h_s_dadda_pg_rca32_and_6_10;
  wire [0:0] h_s_dadda_pg_rca32_fa67_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa67_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_11;
  wire [0:0] h_s_dadda_pg_rca32_and_4_12;
  wire [0:0] h_s_dadda_pg_rca32_and_3_13;
  wire [0:0] h_s_dadda_pg_rca32_fa68_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa68_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_14;
  wire [0:0] h_s_dadda_pg_rca32_and_1_15;
  wire [0:0] h_s_dadda_pg_rca32_and_0_16;
  wire [0:0] h_s_dadda_pg_rca32_fa69_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa69_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa70_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa70_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha14_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha14_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa71_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa71_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa72_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa72_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa73_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa73_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_0;
  wire [0:0] h_s_dadda_pg_rca32_fa74_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa74_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_1;
  wire [0:0] h_s_dadda_pg_rca32_and_15_2;
  wire [0:0] h_s_dadda_pg_rca32_and_14_3;
  wire [0:0] h_s_dadda_pg_rca32_fa75_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa75_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_4;
  wire [0:0] h_s_dadda_pg_rca32_and_12_5;
  wire [0:0] h_s_dadda_pg_rca32_and_11_6;
  wire [0:0] h_s_dadda_pg_rca32_fa76_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa76_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_7;
  wire [0:0] h_s_dadda_pg_rca32_and_9_8;
  wire [0:0] h_s_dadda_pg_rca32_and_8_9;
  wire [0:0] h_s_dadda_pg_rca32_fa77_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa77_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_10;
  wire [0:0] h_s_dadda_pg_rca32_and_6_11;
  wire [0:0] h_s_dadda_pg_rca32_and_5_12;
  wire [0:0] h_s_dadda_pg_rca32_fa78_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa78_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_13;
  wire [0:0] h_s_dadda_pg_rca32_and_3_14;
  wire [0:0] h_s_dadda_pg_rca32_and_2_15;
  wire [0:0] h_s_dadda_pg_rca32_fa79_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa79_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_16;
  wire [0:0] h_s_dadda_pg_rca32_and_0_17;
  wire [0:0] h_s_dadda_pg_rca32_fa80_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa80_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa81_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa81_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha15_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha15_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa82_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa82_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa83_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa83_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa84_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa84_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa85_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa85_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_1;
  wire [0:0] h_s_dadda_pg_rca32_and_16_2;
  wire [0:0] h_s_dadda_pg_rca32_fa86_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa86_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_3;
  wire [0:0] h_s_dadda_pg_rca32_and_14_4;
  wire [0:0] h_s_dadda_pg_rca32_and_13_5;
  wire [0:0] h_s_dadda_pg_rca32_fa87_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa87_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_6;
  wire [0:0] h_s_dadda_pg_rca32_and_11_7;
  wire [0:0] h_s_dadda_pg_rca32_and_10_8;
  wire [0:0] h_s_dadda_pg_rca32_fa88_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa88_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_9;
  wire [0:0] h_s_dadda_pg_rca32_and_8_10;
  wire [0:0] h_s_dadda_pg_rca32_and_7_11;
  wire [0:0] h_s_dadda_pg_rca32_fa89_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa89_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_12;
  wire [0:0] h_s_dadda_pg_rca32_and_5_13;
  wire [0:0] h_s_dadda_pg_rca32_and_4_14;
  wire [0:0] h_s_dadda_pg_rca32_fa90_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa90_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_15;
  wire [0:0] h_s_dadda_pg_rca32_and_2_16;
  wire [0:0] h_s_dadda_pg_rca32_and_1_17;
  wire [0:0] h_s_dadda_pg_rca32_fa91_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa91_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_18;
  wire [0:0] h_s_dadda_pg_rca32_fa92_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa92_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa93_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa93_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha16_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha16_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa94_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa94_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa95_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa95_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa96_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa96_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa97_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa97_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_1;
  wire [0:0] h_s_dadda_pg_rca32_fa98_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa98_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_2;
  wire [0:0] h_s_dadda_pg_rca32_and_16_3;
  wire [0:0] h_s_dadda_pg_rca32_and_15_4;
  wire [0:0] h_s_dadda_pg_rca32_fa99_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa99_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_5;
  wire [0:0] h_s_dadda_pg_rca32_and_13_6;
  wire [0:0] h_s_dadda_pg_rca32_and_12_7;
  wire [0:0] h_s_dadda_pg_rca32_fa100_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa100_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_8;
  wire [0:0] h_s_dadda_pg_rca32_and_10_9;
  wire [0:0] h_s_dadda_pg_rca32_and_9_10;
  wire [0:0] h_s_dadda_pg_rca32_fa101_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa101_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_11;
  wire [0:0] h_s_dadda_pg_rca32_and_7_12;
  wire [0:0] h_s_dadda_pg_rca32_and_6_13;
  wire [0:0] h_s_dadda_pg_rca32_fa102_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa102_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_14;
  wire [0:0] h_s_dadda_pg_rca32_and_4_15;
  wire [0:0] h_s_dadda_pg_rca32_and_3_16;
  wire [0:0] h_s_dadda_pg_rca32_fa103_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa103_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_17;
  wire [0:0] h_s_dadda_pg_rca32_and_1_18;
  wire [0:0] h_s_dadda_pg_rca32_and_0_19;
  wire [0:0] h_s_dadda_pg_rca32_fa104_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa104_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa105_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa105_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa106_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa106_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha17_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha17_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa107_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa107_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa108_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa108_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa109_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa109_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa110_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa110_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_0;
  wire [0:0] h_s_dadda_pg_rca32_fa111_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa111_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_1;
  wire [0:0] h_s_dadda_pg_rca32_and_18_2;
  wire [0:0] h_s_dadda_pg_rca32_and_17_3;
  wire [0:0] h_s_dadda_pg_rca32_fa112_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa112_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_4;
  wire [0:0] h_s_dadda_pg_rca32_and_15_5;
  wire [0:0] h_s_dadda_pg_rca32_and_14_6;
  wire [0:0] h_s_dadda_pg_rca32_fa113_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa113_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_7;
  wire [0:0] h_s_dadda_pg_rca32_and_12_8;
  wire [0:0] h_s_dadda_pg_rca32_and_11_9;
  wire [0:0] h_s_dadda_pg_rca32_fa114_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa114_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_10;
  wire [0:0] h_s_dadda_pg_rca32_and_9_11;
  wire [0:0] h_s_dadda_pg_rca32_and_8_12;
  wire [0:0] h_s_dadda_pg_rca32_fa115_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa115_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_13;
  wire [0:0] h_s_dadda_pg_rca32_and_6_14;
  wire [0:0] h_s_dadda_pg_rca32_and_5_15;
  wire [0:0] h_s_dadda_pg_rca32_fa116_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa116_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_16;
  wire [0:0] h_s_dadda_pg_rca32_and_3_17;
  wire [0:0] h_s_dadda_pg_rca32_and_2_18;
  wire [0:0] h_s_dadda_pg_rca32_fa117_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa117_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_19;
  wire [0:0] h_s_dadda_pg_rca32_and_0_20;
  wire [0:0] h_s_dadda_pg_rca32_fa118_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa118_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa119_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa119_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa120_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa120_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha18_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha18_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa121_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa121_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa122_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa122_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa123_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa123_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa124_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa124_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa125_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa125_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_1;
  wire [0:0] h_s_dadda_pg_rca32_and_19_2;
  wire [0:0] h_s_dadda_pg_rca32_fa126_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa126_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_3;
  wire [0:0] h_s_dadda_pg_rca32_and_17_4;
  wire [0:0] h_s_dadda_pg_rca32_and_16_5;
  wire [0:0] h_s_dadda_pg_rca32_fa127_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa127_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_6;
  wire [0:0] h_s_dadda_pg_rca32_and_14_7;
  wire [0:0] h_s_dadda_pg_rca32_and_13_8;
  wire [0:0] h_s_dadda_pg_rca32_fa128_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa128_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_9;
  wire [0:0] h_s_dadda_pg_rca32_and_11_10;
  wire [0:0] h_s_dadda_pg_rca32_and_10_11;
  wire [0:0] h_s_dadda_pg_rca32_fa129_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa129_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_12;
  wire [0:0] h_s_dadda_pg_rca32_and_8_13;
  wire [0:0] h_s_dadda_pg_rca32_and_7_14;
  wire [0:0] h_s_dadda_pg_rca32_fa130_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa130_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_15;
  wire [0:0] h_s_dadda_pg_rca32_and_5_16;
  wire [0:0] h_s_dadda_pg_rca32_and_4_17;
  wire [0:0] h_s_dadda_pg_rca32_fa131_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa131_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_18;
  wire [0:0] h_s_dadda_pg_rca32_and_2_19;
  wire [0:0] h_s_dadda_pg_rca32_and_1_20;
  wire [0:0] h_s_dadda_pg_rca32_fa132_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa132_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_21;
  wire [0:0] h_s_dadda_pg_rca32_fa133_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa133_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa134_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa134_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa135_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa135_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha19_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha19_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa136_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa136_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa137_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa137_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa138_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa138_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa139_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa139_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa140_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa140_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_1;
  wire [0:0] h_s_dadda_pg_rca32_fa141_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa141_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_2;
  wire [0:0] h_s_dadda_pg_rca32_and_19_3;
  wire [0:0] h_s_dadda_pg_rca32_and_18_4;
  wire [0:0] h_s_dadda_pg_rca32_fa142_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa142_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_5;
  wire [0:0] h_s_dadda_pg_rca32_and_16_6;
  wire [0:0] h_s_dadda_pg_rca32_and_15_7;
  wire [0:0] h_s_dadda_pg_rca32_fa143_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa143_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_8;
  wire [0:0] h_s_dadda_pg_rca32_and_13_9;
  wire [0:0] h_s_dadda_pg_rca32_and_12_10;
  wire [0:0] h_s_dadda_pg_rca32_fa144_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa144_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_11;
  wire [0:0] h_s_dadda_pg_rca32_and_10_12;
  wire [0:0] h_s_dadda_pg_rca32_and_9_13;
  wire [0:0] h_s_dadda_pg_rca32_fa145_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa145_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_14;
  wire [0:0] h_s_dadda_pg_rca32_and_7_15;
  wire [0:0] h_s_dadda_pg_rca32_and_6_16;
  wire [0:0] h_s_dadda_pg_rca32_fa146_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa146_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_17;
  wire [0:0] h_s_dadda_pg_rca32_and_4_18;
  wire [0:0] h_s_dadda_pg_rca32_and_3_19;
  wire [0:0] h_s_dadda_pg_rca32_fa147_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa147_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_20;
  wire [0:0] h_s_dadda_pg_rca32_and_1_21;
  wire [0:0] h_s_dadda_pg_rca32_and_0_22;
  wire [0:0] h_s_dadda_pg_rca32_fa148_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa148_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa149_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa149_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa150_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa150_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa151_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa151_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha20_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha20_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa152_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa152_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa153_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa153_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa154_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa154_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa155_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa155_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa156_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa156_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_0;
  wire [0:0] h_s_dadda_pg_rca32_fa157_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa157_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_1;
  wire [0:0] h_s_dadda_pg_rca32_and_21_2;
  wire [0:0] h_s_dadda_pg_rca32_and_20_3;
  wire [0:0] h_s_dadda_pg_rca32_fa158_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa158_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_4;
  wire [0:0] h_s_dadda_pg_rca32_and_18_5;
  wire [0:0] h_s_dadda_pg_rca32_and_17_6;
  wire [0:0] h_s_dadda_pg_rca32_fa159_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa159_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_7;
  wire [0:0] h_s_dadda_pg_rca32_and_15_8;
  wire [0:0] h_s_dadda_pg_rca32_and_14_9;
  wire [0:0] h_s_dadda_pg_rca32_fa160_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa160_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_10;
  wire [0:0] h_s_dadda_pg_rca32_and_12_11;
  wire [0:0] h_s_dadda_pg_rca32_and_11_12;
  wire [0:0] h_s_dadda_pg_rca32_fa161_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa161_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_13;
  wire [0:0] h_s_dadda_pg_rca32_and_9_14;
  wire [0:0] h_s_dadda_pg_rca32_and_8_15;
  wire [0:0] h_s_dadda_pg_rca32_fa162_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa162_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_16;
  wire [0:0] h_s_dadda_pg_rca32_and_6_17;
  wire [0:0] h_s_dadda_pg_rca32_and_5_18;
  wire [0:0] h_s_dadda_pg_rca32_fa163_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa163_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_19;
  wire [0:0] h_s_dadda_pg_rca32_and_3_20;
  wire [0:0] h_s_dadda_pg_rca32_and_2_21;
  wire [0:0] h_s_dadda_pg_rca32_fa164_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa164_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_22;
  wire [0:0] h_s_dadda_pg_rca32_and_0_23;
  wire [0:0] h_s_dadda_pg_rca32_fa165_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa165_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa166_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa166_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa167_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa167_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa168_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa168_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha21_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha21_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa169_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa169_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa170_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa170_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa171_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa171_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa172_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa172_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa173_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa173_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa174_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa174_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_1;
  wire [0:0] h_s_dadda_pg_rca32_and_22_2;
  wire [0:0] h_s_dadda_pg_rca32_fa175_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa175_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_3;
  wire [0:0] h_s_dadda_pg_rca32_and_20_4;
  wire [0:0] h_s_dadda_pg_rca32_and_19_5;
  wire [0:0] h_s_dadda_pg_rca32_fa176_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa176_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_6;
  wire [0:0] h_s_dadda_pg_rca32_and_17_7;
  wire [0:0] h_s_dadda_pg_rca32_and_16_8;
  wire [0:0] h_s_dadda_pg_rca32_fa177_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa177_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_9;
  wire [0:0] h_s_dadda_pg_rca32_and_14_10;
  wire [0:0] h_s_dadda_pg_rca32_and_13_11;
  wire [0:0] h_s_dadda_pg_rca32_fa178_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa178_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_12;
  wire [0:0] h_s_dadda_pg_rca32_and_11_13;
  wire [0:0] h_s_dadda_pg_rca32_and_10_14;
  wire [0:0] h_s_dadda_pg_rca32_fa179_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa179_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_15;
  wire [0:0] h_s_dadda_pg_rca32_and_8_16;
  wire [0:0] h_s_dadda_pg_rca32_and_7_17;
  wire [0:0] h_s_dadda_pg_rca32_fa180_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa180_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_18;
  wire [0:0] h_s_dadda_pg_rca32_and_5_19;
  wire [0:0] h_s_dadda_pg_rca32_and_4_20;
  wire [0:0] h_s_dadda_pg_rca32_fa181_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa181_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_21;
  wire [0:0] h_s_dadda_pg_rca32_and_2_22;
  wire [0:0] h_s_dadda_pg_rca32_and_1_23;
  wire [0:0] h_s_dadda_pg_rca32_fa182_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa182_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_24;
  wire [0:0] h_s_dadda_pg_rca32_fa183_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa183_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa184_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa184_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa185_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa185_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa186_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa186_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha22_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha22_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa187_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa187_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa188_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa188_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa189_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa189_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa190_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa190_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa191_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa191_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa192_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa192_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_1;
  wire [0:0] h_s_dadda_pg_rca32_fa193_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa193_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_2;
  wire [0:0] h_s_dadda_pg_rca32_and_22_3;
  wire [0:0] h_s_dadda_pg_rca32_and_21_4;
  wire [0:0] h_s_dadda_pg_rca32_fa194_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa194_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_5;
  wire [0:0] h_s_dadda_pg_rca32_and_19_6;
  wire [0:0] h_s_dadda_pg_rca32_and_18_7;
  wire [0:0] h_s_dadda_pg_rca32_fa195_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa195_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_8;
  wire [0:0] h_s_dadda_pg_rca32_and_16_9;
  wire [0:0] h_s_dadda_pg_rca32_and_15_10;
  wire [0:0] h_s_dadda_pg_rca32_fa196_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa196_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_11;
  wire [0:0] h_s_dadda_pg_rca32_and_13_12;
  wire [0:0] h_s_dadda_pg_rca32_and_12_13;
  wire [0:0] h_s_dadda_pg_rca32_fa197_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa197_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_14;
  wire [0:0] h_s_dadda_pg_rca32_and_10_15;
  wire [0:0] h_s_dadda_pg_rca32_and_9_16;
  wire [0:0] h_s_dadda_pg_rca32_fa198_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa198_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_17;
  wire [0:0] h_s_dadda_pg_rca32_and_7_18;
  wire [0:0] h_s_dadda_pg_rca32_and_6_19;
  wire [0:0] h_s_dadda_pg_rca32_fa199_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa199_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_20;
  wire [0:0] h_s_dadda_pg_rca32_and_4_21;
  wire [0:0] h_s_dadda_pg_rca32_and_3_22;
  wire [0:0] h_s_dadda_pg_rca32_fa200_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa200_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_23;
  wire [0:0] h_s_dadda_pg_rca32_and_1_24;
  wire [0:0] h_s_dadda_pg_rca32_and_0_25;
  wire [0:0] h_s_dadda_pg_rca32_fa201_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa201_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa202_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa202_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa203_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa203_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa204_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa204_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa205_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa205_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha23_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha23_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa206_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa206_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa207_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa207_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa208_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa208_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa209_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa209_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa210_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa210_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa211_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa211_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_0;
  wire [0:0] h_s_dadda_pg_rca32_fa212_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa212_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_1;
  wire [0:0] h_s_dadda_pg_rca32_and_24_2;
  wire [0:0] h_s_dadda_pg_rca32_and_23_3;
  wire [0:0] h_s_dadda_pg_rca32_fa213_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa213_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_4;
  wire [0:0] h_s_dadda_pg_rca32_and_21_5;
  wire [0:0] h_s_dadda_pg_rca32_and_20_6;
  wire [0:0] h_s_dadda_pg_rca32_fa214_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa214_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_7;
  wire [0:0] h_s_dadda_pg_rca32_and_18_8;
  wire [0:0] h_s_dadda_pg_rca32_and_17_9;
  wire [0:0] h_s_dadda_pg_rca32_fa215_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa215_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_10;
  wire [0:0] h_s_dadda_pg_rca32_and_15_11;
  wire [0:0] h_s_dadda_pg_rca32_and_14_12;
  wire [0:0] h_s_dadda_pg_rca32_fa216_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa216_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_13;
  wire [0:0] h_s_dadda_pg_rca32_and_12_14;
  wire [0:0] h_s_dadda_pg_rca32_and_11_15;
  wire [0:0] h_s_dadda_pg_rca32_fa217_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa217_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_16;
  wire [0:0] h_s_dadda_pg_rca32_and_9_17;
  wire [0:0] h_s_dadda_pg_rca32_and_8_18;
  wire [0:0] h_s_dadda_pg_rca32_fa218_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa218_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_19;
  wire [0:0] h_s_dadda_pg_rca32_and_6_20;
  wire [0:0] h_s_dadda_pg_rca32_and_5_21;
  wire [0:0] h_s_dadda_pg_rca32_fa219_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa219_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_22;
  wire [0:0] h_s_dadda_pg_rca32_and_3_23;
  wire [0:0] h_s_dadda_pg_rca32_and_2_24;
  wire [0:0] h_s_dadda_pg_rca32_fa220_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa220_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_25;
  wire [0:0] h_s_dadda_pg_rca32_and_0_26;
  wire [0:0] h_s_dadda_pg_rca32_fa221_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa221_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa222_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa222_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa223_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa223_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa224_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa224_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa225_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa225_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha24_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha24_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa226_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa226_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa227_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa227_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa228_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa228_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa229_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa229_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa230_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa230_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa231_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa231_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa232_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa232_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_1;
  wire [0:0] h_s_dadda_pg_rca32_and_25_2;
  wire [0:0] h_s_dadda_pg_rca32_fa233_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa233_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_3;
  wire [0:0] h_s_dadda_pg_rca32_and_23_4;
  wire [0:0] h_s_dadda_pg_rca32_and_22_5;
  wire [0:0] h_s_dadda_pg_rca32_fa234_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa234_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_6;
  wire [0:0] h_s_dadda_pg_rca32_and_20_7;
  wire [0:0] h_s_dadda_pg_rca32_and_19_8;
  wire [0:0] h_s_dadda_pg_rca32_fa235_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa235_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_9;
  wire [0:0] h_s_dadda_pg_rca32_and_17_10;
  wire [0:0] h_s_dadda_pg_rca32_and_16_11;
  wire [0:0] h_s_dadda_pg_rca32_fa236_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa236_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_12;
  wire [0:0] h_s_dadda_pg_rca32_and_14_13;
  wire [0:0] h_s_dadda_pg_rca32_and_13_14;
  wire [0:0] h_s_dadda_pg_rca32_fa237_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa237_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_15;
  wire [0:0] h_s_dadda_pg_rca32_and_11_16;
  wire [0:0] h_s_dadda_pg_rca32_and_10_17;
  wire [0:0] h_s_dadda_pg_rca32_fa238_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa238_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_18;
  wire [0:0] h_s_dadda_pg_rca32_and_8_19;
  wire [0:0] h_s_dadda_pg_rca32_and_7_20;
  wire [0:0] h_s_dadda_pg_rca32_fa239_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa239_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_21;
  wire [0:0] h_s_dadda_pg_rca32_and_5_22;
  wire [0:0] h_s_dadda_pg_rca32_and_4_23;
  wire [0:0] h_s_dadda_pg_rca32_fa240_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa240_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_24;
  wire [0:0] h_s_dadda_pg_rca32_and_2_25;
  wire [0:0] h_s_dadda_pg_rca32_and_1_26;
  wire [0:0] h_s_dadda_pg_rca32_fa241_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa241_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_27;
  wire [0:0] h_s_dadda_pg_rca32_fa242_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa242_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa243_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa243_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa244_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa244_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa245_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa245_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa246_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa246_or0;
  wire [0:0] h_s_dadda_pg_rca32_ha25_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha25_and0;
  wire [0:0] h_s_dadda_pg_rca32_fa247_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa247_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa248_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa248_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa249_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa249_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa250_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa250_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa251_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa251_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa252_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa252_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa253_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa253_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_2;
  wire [0:0] h_s_dadda_pg_rca32_and_25_3;
  wire [0:0] h_s_dadda_pg_rca32_fa254_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa254_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_4;
  wire [0:0] h_s_dadda_pg_rca32_and_23_5;
  wire [0:0] h_s_dadda_pg_rca32_and_22_6;
  wire [0:0] h_s_dadda_pg_rca32_fa255_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa255_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_7;
  wire [0:0] h_s_dadda_pg_rca32_and_20_8;
  wire [0:0] h_s_dadda_pg_rca32_and_19_9;
  wire [0:0] h_s_dadda_pg_rca32_fa256_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa256_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_10;
  wire [0:0] h_s_dadda_pg_rca32_and_17_11;
  wire [0:0] h_s_dadda_pg_rca32_and_16_12;
  wire [0:0] h_s_dadda_pg_rca32_fa257_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa257_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_13;
  wire [0:0] h_s_dadda_pg_rca32_and_14_14;
  wire [0:0] h_s_dadda_pg_rca32_and_13_15;
  wire [0:0] h_s_dadda_pg_rca32_fa258_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa258_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_16;
  wire [0:0] h_s_dadda_pg_rca32_and_11_17;
  wire [0:0] h_s_dadda_pg_rca32_and_10_18;
  wire [0:0] h_s_dadda_pg_rca32_fa259_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa259_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_19;
  wire [0:0] h_s_dadda_pg_rca32_and_8_20;
  wire [0:0] h_s_dadda_pg_rca32_and_7_21;
  wire [0:0] h_s_dadda_pg_rca32_fa260_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa260_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_22;
  wire [0:0] h_s_dadda_pg_rca32_and_5_23;
  wire [0:0] h_s_dadda_pg_rca32_and_4_24;
  wire [0:0] h_s_dadda_pg_rca32_fa261_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa261_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_25;
  wire [0:0] h_s_dadda_pg_rca32_and_2_26;
  wire [0:0] h_s_dadda_pg_rca32_and_1_27;
  wire [0:0] h_s_dadda_pg_rca32_fa262_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa262_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_28;
  wire [0:0] h_s_dadda_pg_rca32_fa263_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa263_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa264_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa264_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa265_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa265_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa266_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa266_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa267_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa267_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa268_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa268_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa269_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa269_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa270_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa270_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa271_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa271_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa272_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa272_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa273_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa273_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa274_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa274_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa275_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa275_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_4;
  wire [0:0] h_s_dadda_pg_rca32_and_24_5;
  wire [0:0] h_s_dadda_pg_rca32_fa276_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa276_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_6;
  wire [0:0] h_s_dadda_pg_rca32_and_22_7;
  wire [0:0] h_s_dadda_pg_rca32_and_21_8;
  wire [0:0] h_s_dadda_pg_rca32_fa277_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa277_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_9;
  wire [0:0] h_s_dadda_pg_rca32_and_19_10;
  wire [0:0] h_s_dadda_pg_rca32_and_18_11;
  wire [0:0] h_s_dadda_pg_rca32_fa278_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa278_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_12;
  wire [0:0] h_s_dadda_pg_rca32_and_16_13;
  wire [0:0] h_s_dadda_pg_rca32_and_15_14;
  wire [0:0] h_s_dadda_pg_rca32_fa279_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa279_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_15;
  wire [0:0] h_s_dadda_pg_rca32_and_13_16;
  wire [0:0] h_s_dadda_pg_rca32_and_12_17;
  wire [0:0] h_s_dadda_pg_rca32_fa280_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa280_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_18;
  wire [0:0] h_s_dadda_pg_rca32_and_10_19;
  wire [0:0] h_s_dadda_pg_rca32_and_9_20;
  wire [0:0] h_s_dadda_pg_rca32_fa281_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa281_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_21;
  wire [0:0] h_s_dadda_pg_rca32_and_7_22;
  wire [0:0] h_s_dadda_pg_rca32_and_6_23;
  wire [0:0] h_s_dadda_pg_rca32_fa282_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa282_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_24;
  wire [0:0] h_s_dadda_pg_rca32_and_4_25;
  wire [0:0] h_s_dadda_pg_rca32_and_3_26;
  wire [0:0] h_s_dadda_pg_rca32_fa283_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa283_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_27;
  wire [0:0] h_s_dadda_pg_rca32_and_1_28;
  wire [0:0] h_s_dadda_pg_rca32_and_0_29;
  wire [0:0] h_s_dadda_pg_rca32_fa284_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa284_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa285_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa285_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa286_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa286_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa287_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa287_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa288_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa288_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa289_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa289_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa290_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa290_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa291_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa291_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa292_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa292_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa293_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa293_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa294_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa294_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa295_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa295_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa296_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa296_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa297_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa297_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_6;
  wire [0:0] h_s_dadda_pg_rca32_and_23_7;
  wire [0:0] h_s_dadda_pg_rca32_fa298_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa298_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_8;
  wire [0:0] h_s_dadda_pg_rca32_and_21_9;
  wire [0:0] h_s_dadda_pg_rca32_and_20_10;
  wire [0:0] h_s_dadda_pg_rca32_fa299_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa299_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_11;
  wire [0:0] h_s_dadda_pg_rca32_and_18_12;
  wire [0:0] h_s_dadda_pg_rca32_and_17_13;
  wire [0:0] h_s_dadda_pg_rca32_fa300_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa300_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_14;
  wire [0:0] h_s_dadda_pg_rca32_and_15_15;
  wire [0:0] h_s_dadda_pg_rca32_and_14_16;
  wire [0:0] h_s_dadda_pg_rca32_fa301_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa301_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_17;
  wire [0:0] h_s_dadda_pg_rca32_and_12_18;
  wire [0:0] h_s_dadda_pg_rca32_and_11_19;
  wire [0:0] h_s_dadda_pg_rca32_fa302_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa302_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_20;
  wire [0:0] h_s_dadda_pg_rca32_and_9_21;
  wire [0:0] h_s_dadda_pg_rca32_and_8_22;
  wire [0:0] h_s_dadda_pg_rca32_fa303_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa303_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_23;
  wire [0:0] h_s_dadda_pg_rca32_and_6_24;
  wire [0:0] h_s_dadda_pg_rca32_and_5_25;
  wire [0:0] h_s_dadda_pg_rca32_fa304_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa304_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_26;
  wire [0:0] h_s_dadda_pg_rca32_and_3_27;
  wire [0:0] h_s_dadda_pg_rca32_and_2_28;
  wire [0:0] h_s_dadda_pg_rca32_fa305_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa305_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_29;
  wire [0:0] h_s_dadda_pg_rca32_and_0_30;
  wire [0:0] h_s_dadda_pg_rca32_fa306_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa306_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa307_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa307_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa308_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa308_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa309_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa309_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa310_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa310_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa311_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa311_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa312_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa312_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa313_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa313_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa314_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa314_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa315_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa315_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa316_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa316_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa317_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa317_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa318_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa318_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa319_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa319_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_8;
  wire [0:0] h_s_dadda_pg_rca32_and_22_9;
  wire [0:0] h_s_dadda_pg_rca32_fa320_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa320_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_10;
  wire [0:0] h_s_dadda_pg_rca32_and_20_11;
  wire [0:0] h_s_dadda_pg_rca32_and_19_12;
  wire [0:0] h_s_dadda_pg_rca32_fa321_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa321_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_13;
  wire [0:0] h_s_dadda_pg_rca32_and_17_14;
  wire [0:0] h_s_dadda_pg_rca32_and_16_15;
  wire [0:0] h_s_dadda_pg_rca32_fa322_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa322_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_16;
  wire [0:0] h_s_dadda_pg_rca32_and_14_17;
  wire [0:0] h_s_dadda_pg_rca32_and_13_18;
  wire [0:0] h_s_dadda_pg_rca32_fa323_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa323_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_19;
  wire [0:0] h_s_dadda_pg_rca32_and_11_20;
  wire [0:0] h_s_dadda_pg_rca32_and_10_21;
  wire [0:0] h_s_dadda_pg_rca32_fa324_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa324_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_22;
  wire [0:0] h_s_dadda_pg_rca32_and_8_23;
  wire [0:0] h_s_dadda_pg_rca32_and_7_24;
  wire [0:0] h_s_dadda_pg_rca32_fa325_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa325_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_25;
  wire [0:0] h_s_dadda_pg_rca32_and_5_26;
  wire [0:0] h_s_dadda_pg_rca32_and_4_27;
  wire [0:0] h_s_dadda_pg_rca32_fa326_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa326_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_28;
  wire [0:0] h_s_dadda_pg_rca32_and_2_29;
  wire [0:0] h_s_dadda_pg_rca32_and_1_30;
  wire [0:0] h_s_dadda_pg_rca32_fa327_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa327_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_0_31;
  wire [0:0] h_s_dadda_pg_rca32_fa328_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa328_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa329_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa329_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa330_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa330_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa331_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa331_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa332_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa332_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa333_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa333_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa334_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa334_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa335_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa335_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa336_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa336_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa337_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa337_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa338_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa338_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa339_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa339_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa340_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa340_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa341_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa341_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_8;
  wire [0:0] h_s_dadda_pg_rca32_and_23_9;
  wire [0:0] h_s_dadda_pg_rca32_fa342_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa342_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_10;
  wire [0:0] h_s_dadda_pg_rca32_and_21_11;
  wire [0:0] h_s_dadda_pg_rca32_and_20_12;
  wire [0:0] h_s_dadda_pg_rca32_fa343_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa343_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_13;
  wire [0:0] h_s_dadda_pg_rca32_and_18_14;
  wire [0:0] h_s_dadda_pg_rca32_and_17_15;
  wire [0:0] h_s_dadda_pg_rca32_fa344_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa344_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_16;
  wire [0:0] h_s_dadda_pg_rca32_and_15_17;
  wire [0:0] h_s_dadda_pg_rca32_and_14_18;
  wire [0:0] h_s_dadda_pg_rca32_fa345_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa345_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_19;
  wire [0:0] h_s_dadda_pg_rca32_and_12_20;
  wire [0:0] h_s_dadda_pg_rca32_and_11_21;
  wire [0:0] h_s_dadda_pg_rca32_fa346_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa346_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_22;
  wire [0:0] h_s_dadda_pg_rca32_and_9_23;
  wire [0:0] h_s_dadda_pg_rca32_and_8_24;
  wire [0:0] h_s_dadda_pg_rca32_fa347_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa347_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_25;
  wire [0:0] h_s_dadda_pg_rca32_and_6_26;
  wire [0:0] h_s_dadda_pg_rca32_and_5_27;
  wire [0:0] h_s_dadda_pg_rca32_fa348_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa348_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_28;
  wire [0:0] h_s_dadda_pg_rca32_and_3_29;
  wire [0:0] h_s_dadda_pg_rca32_and_2_30;
  wire [0:0] h_s_dadda_pg_rca32_fa349_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa349_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_1_31;
  wire [0:0] h_s_dadda_pg_rca32_fa350_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa350_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa351_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa351_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa352_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa352_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa353_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa353_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa354_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa354_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa355_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa355_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa356_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa356_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa357_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa357_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa358_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa358_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa359_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa359_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa360_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa360_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa361_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa361_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa362_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa362_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa363_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa363_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_7;
  wire [0:0] h_s_dadda_pg_rca32_and_25_8;
  wire [0:0] h_s_dadda_pg_rca32_fa364_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa364_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_9;
  wire [0:0] h_s_dadda_pg_rca32_and_23_10;
  wire [0:0] h_s_dadda_pg_rca32_and_22_11;
  wire [0:0] h_s_dadda_pg_rca32_fa365_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa365_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_12;
  wire [0:0] h_s_dadda_pg_rca32_and_20_13;
  wire [0:0] h_s_dadda_pg_rca32_and_19_14;
  wire [0:0] h_s_dadda_pg_rca32_fa366_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa366_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_15;
  wire [0:0] h_s_dadda_pg_rca32_and_17_16;
  wire [0:0] h_s_dadda_pg_rca32_and_16_17;
  wire [0:0] h_s_dadda_pg_rca32_fa367_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa367_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_18;
  wire [0:0] h_s_dadda_pg_rca32_and_14_19;
  wire [0:0] h_s_dadda_pg_rca32_and_13_20;
  wire [0:0] h_s_dadda_pg_rca32_fa368_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa368_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_21;
  wire [0:0] h_s_dadda_pg_rca32_and_11_22;
  wire [0:0] h_s_dadda_pg_rca32_and_10_23;
  wire [0:0] h_s_dadda_pg_rca32_fa369_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa369_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_24;
  wire [0:0] h_s_dadda_pg_rca32_and_8_25;
  wire [0:0] h_s_dadda_pg_rca32_and_7_26;
  wire [0:0] h_s_dadda_pg_rca32_fa370_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa370_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_27;
  wire [0:0] h_s_dadda_pg_rca32_and_5_28;
  wire [0:0] h_s_dadda_pg_rca32_and_4_29;
  wire [0:0] h_s_dadda_pg_rca32_fa371_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa371_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_2_31;
  wire [0:0] h_s_dadda_pg_rca32_fa372_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa372_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa373_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa373_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa374_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa374_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa375_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa375_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa376_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa376_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa377_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa377_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa378_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa378_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa379_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa379_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa380_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa380_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa381_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa381_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa382_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa382_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa383_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa383_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa384_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa384_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa385_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa385_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_6;
  wire [0:0] h_s_dadda_pg_rca32_and_27_7;
  wire [0:0] h_s_dadda_pg_rca32_fa386_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa386_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_8;
  wire [0:0] h_s_dadda_pg_rca32_and_25_9;
  wire [0:0] h_s_dadda_pg_rca32_and_24_10;
  wire [0:0] h_s_dadda_pg_rca32_fa387_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa387_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_11;
  wire [0:0] h_s_dadda_pg_rca32_and_22_12;
  wire [0:0] h_s_dadda_pg_rca32_and_21_13;
  wire [0:0] h_s_dadda_pg_rca32_fa388_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa388_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_14;
  wire [0:0] h_s_dadda_pg_rca32_and_19_15;
  wire [0:0] h_s_dadda_pg_rca32_and_18_16;
  wire [0:0] h_s_dadda_pg_rca32_fa389_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa389_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_17;
  wire [0:0] h_s_dadda_pg_rca32_and_16_18;
  wire [0:0] h_s_dadda_pg_rca32_and_15_19;
  wire [0:0] h_s_dadda_pg_rca32_fa390_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa390_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_20;
  wire [0:0] h_s_dadda_pg_rca32_and_13_21;
  wire [0:0] h_s_dadda_pg_rca32_and_12_22;
  wire [0:0] h_s_dadda_pg_rca32_fa391_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa391_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_23;
  wire [0:0] h_s_dadda_pg_rca32_and_10_24;
  wire [0:0] h_s_dadda_pg_rca32_and_9_25;
  wire [0:0] h_s_dadda_pg_rca32_fa392_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa392_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_26;
  wire [0:0] h_s_dadda_pg_rca32_and_7_27;
  wire [0:0] h_s_dadda_pg_rca32_and_6_28;
  wire [0:0] h_s_dadda_pg_rca32_fa393_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa393_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_29;
  wire [0:0] h_s_dadda_pg_rca32_and_4_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_3_31;
  wire [0:0] h_s_dadda_pg_rca32_fa394_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa394_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa395_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa395_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa396_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa396_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa397_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa397_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa398_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa398_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa399_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa399_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa400_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa400_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa401_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa401_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa402_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa402_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa403_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa403_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa404_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa404_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa405_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa405_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa406_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa406_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa407_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa407_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_5;
  wire [0:0] h_s_dadda_pg_rca32_and_29_6;
  wire [0:0] h_s_dadda_pg_rca32_fa408_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa408_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_7;
  wire [0:0] h_s_dadda_pg_rca32_and_27_8;
  wire [0:0] h_s_dadda_pg_rca32_and_26_9;
  wire [0:0] h_s_dadda_pg_rca32_fa409_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa409_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_10;
  wire [0:0] h_s_dadda_pg_rca32_and_24_11;
  wire [0:0] h_s_dadda_pg_rca32_and_23_12;
  wire [0:0] h_s_dadda_pg_rca32_fa410_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa410_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_13;
  wire [0:0] h_s_dadda_pg_rca32_and_21_14;
  wire [0:0] h_s_dadda_pg_rca32_and_20_15;
  wire [0:0] h_s_dadda_pg_rca32_fa411_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa411_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_16;
  wire [0:0] h_s_dadda_pg_rca32_and_18_17;
  wire [0:0] h_s_dadda_pg_rca32_and_17_18;
  wire [0:0] h_s_dadda_pg_rca32_fa412_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa412_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_19;
  wire [0:0] h_s_dadda_pg_rca32_and_15_20;
  wire [0:0] h_s_dadda_pg_rca32_and_14_21;
  wire [0:0] h_s_dadda_pg_rca32_fa413_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa413_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_22;
  wire [0:0] h_s_dadda_pg_rca32_and_12_23;
  wire [0:0] h_s_dadda_pg_rca32_and_11_24;
  wire [0:0] h_s_dadda_pg_rca32_fa414_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa414_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_25;
  wire [0:0] h_s_dadda_pg_rca32_and_9_26;
  wire [0:0] h_s_dadda_pg_rca32_and_8_27;
  wire [0:0] h_s_dadda_pg_rca32_fa415_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa415_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_7_28;
  wire [0:0] h_s_dadda_pg_rca32_and_6_29;
  wire [0:0] h_s_dadda_pg_rca32_and_5_30;
  wire [0:0] h_s_dadda_pg_rca32_fa416_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa416_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_4_31;
  wire [0:0] h_s_dadda_pg_rca32_fa417_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa417_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa418_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa418_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa419_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa419_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa420_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa420_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa421_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa421_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa422_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa422_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa423_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa423_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa424_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa424_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa425_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa425_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa426_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa426_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa427_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa427_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa428_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa428_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa429_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa429_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_5;
  wire [0:0] h_s_dadda_pg_rca32_fa430_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa430_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_6;
  wire [0:0] h_s_dadda_pg_rca32_and_29_7;
  wire [0:0] h_s_dadda_pg_rca32_and_28_8;
  wire [0:0] h_s_dadda_pg_rca32_fa431_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa431_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_9;
  wire [0:0] h_s_dadda_pg_rca32_and_26_10;
  wire [0:0] h_s_dadda_pg_rca32_and_25_11;
  wire [0:0] h_s_dadda_pg_rca32_fa432_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa432_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_12;
  wire [0:0] h_s_dadda_pg_rca32_and_23_13;
  wire [0:0] h_s_dadda_pg_rca32_and_22_14;
  wire [0:0] h_s_dadda_pg_rca32_fa433_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa433_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_15;
  wire [0:0] h_s_dadda_pg_rca32_and_20_16;
  wire [0:0] h_s_dadda_pg_rca32_and_19_17;
  wire [0:0] h_s_dadda_pg_rca32_fa434_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa434_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_18;
  wire [0:0] h_s_dadda_pg_rca32_and_17_19;
  wire [0:0] h_s_dadda_pg_rca32_and_16_20;
  wire [0:0] h_s_dadda_pg_rca32_fa435_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa435_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_21;
  wire [0:0] h_s_dadda_pg_rca32_and_14_22;
  wire [0:0] h_s_dadda_pg_rca32_and_13_23;
  wire [0:0] h_s_dadda_pg_rca32_fa436_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa436_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_24;
  wire [0:0] h_s_dadda_pg_rca32_and_11_25;
  wire [0:0] h_s_dadda_pg_rca32_and_10_26;
  wire [0:0] h_s_dadda_pg_rca32_fa437_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa437_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_27;
  wire [0:0] h_s_dadda_pg_rca32_and_8_28;
  wire [0:0] h_s_dadda_pg_rca32_and_7_29;
  wire [0:0] h_s_dadda_pg_rca32_fa438_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa438_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_6_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_5_31;
  wire [0:0] h_s_dadda_pg_rca32_fa439_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa439_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa440_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa440_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa441_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa441_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa442_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa442_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa443_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa443_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa444_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa444_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa445_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa445_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa446_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa446_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa447_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa447_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa448_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa448_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa449_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa449_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa450_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa450_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa451_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa451_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_6;
  wire [0:0] h_s_dadda_pg_rca32_and_30_7;
  wire [0:0] h_s_dadda_pg_rca32_fa452_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa452_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_8;
  wire [0:0] h_s_dadda_pg_rca32_and_28_9;
  wire [0:0] h_s_dadda_pg_rca32_and_27_10;
  wire [0:0] h_s_dadda_pg_rca32_fa453_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa453_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_11;
  wire [0:0] h_s_dadda_pg_rca32_and_25_12;
  wire [0:0] h_s_dadda_pg_rca32_and_24_13;
  wire [0:0] h_s_dadda_pg_rca32_fa454_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa454_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_14;
  wire [0:0] h_s_dadda_pg_rca32_and_22_15;
  wire [0:0] h_s_dadda_pg_rca32_and_21_16;
  wire [0:0] h_s_dadda_pg_rca32_fa455_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa455_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_17;
  wire [0:0] h_s_dadda_pg_rca32_and_19_18;
  wire [0:0] h_s_dadda_pg_rca32_and_18_19;
  wire [0:0] h_s_dadda_pg_rca32_fa456_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa456_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_20;
  wire [0:0] h_s_dadda_pg_rca32_and_16_21;
  wire [0:0] h_s_dadda_pg_rca32_and_15_22;
  wire [0:0] h_s_dadda_pg_rca32_fa457_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa457_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_23;
  wire [0:0] h_s_dadda_pg_rca32_and_13_24;
  wire [0:0] h_s_dadda_pg_rca32_and_12_25;
  wire [0:0] h_s_dadda_pg_rca32_fa458_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa458_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_26;
  wire [0:0] h_s_dadda_pg_rca32_and_10_27;
  wire [0:0] h_s_dadda_pg_rca32_and_9_28;
  wire [0:0] h_s_dadda_pg_rca32_fa459_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa459_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_8_29;
  wire [0:0] h_s_dadda_pg_rca32_and_7_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_6_31;
  wire [0:0] h_s_dadda_pg_rca32_fa460_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa460_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa461_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa461_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa462_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa462_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa463_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa463_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa464_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa464_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa465_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa465_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa466_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa466_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa467_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa467_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa468_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa468_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa469_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa469_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa470_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa470_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa471_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa471_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa472_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa472_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_7;
  wire [0:0] h_s_dadda_pg_rca32_and_30_8;
  wire [0:0] h_s_dadda_pg_rca32_and_29_9;
  wire [0:0] h_s_dadda_pg_rca32_fa473_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa473_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_10;
  wire [0:0] h_s_dadda_pg_rca32_and_27_11;
  wire [0:0] h_s_dadda_pg_rca32_and_26_12;
  wire [0:0] h_s_dadda_pg_rca32_fa474_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa474_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_13;
  wire [0:0] h_s_dadda_pg_rca32_and_24_14;
  wire [0:0] h_s_dadda_pg_rca32_and_23_15;
  wire [0:0] h_s_dadda_pg_rca32_fa475_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa475_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_16;
  wire [0:0] h_s_dadda_pg_rca32_and_21_17;
  wire [0:0] h_s_dadda_pg_rca32_and_20_18;
  wire [0:0] h_s_dadda_pg_rca32_fa476_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa476_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_19;
  wire [0:0] h_s_dadda_pg_rca32_and_18_20;
  wire [0:0] h_s_dadda_pg_rca32_and_17_21;
  wire [0:0] h_s_dadda_pg_rca32_fa477_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa477_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_22;
  wire [0:0] h_s_dadda_pg_rca32_and_15_23;
  wire [0:0] h_s_dadda_pg_rca32_and_14_24;
  wire [0:0] h_s_dadda_pg_rca32_fa478_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa478_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_25;
  wire [0:0] h_s_dadda_pg_rca32_and_12_26;
  wire [0:0] h_s_dadda_pg_rca32_and_11_27;
  wire [0:0] h_s_dadda_pg_rca32_fa479_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa479_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_10_28;
  wire [0:0] h_s_dadda_pg_rca32_and_9_29;
  wire [0:0] h_s_dadda_pg_rca32_and_8_30;
  wire [0:0] h_s_dadda_pg_rca32_fa480_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa480_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_7_31;
  wire [0:0] h_s_dadda_pg_rca32_fa481_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa481_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa482_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa482_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa483_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa483_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa484_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa484_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa485_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa485_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa486_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa486_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa487_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa487_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa488_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa488_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa489_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa489_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa490_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa490_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa491_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa491_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_8;
  wire [0:0] h_s_dadda_pg_rca32_fa492_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa492_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_9;
  wire [0:0] h_s_dadda_pg_rca32_and_29_10;
  wire [0:0] h_s_dadda_pg_rca32_and_28_11;
  wire [0:0] h_s_dadda_pg_rca32_fa493_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa493_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_12;
  wire [0:0] h_s_dadda_pg_rca32_and_26_13;
  wire [0:0] h_s_dadda_pg_rca32_and_25_14;
  wire [0:0] h_s_dadda_pg_rca32_fa494_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa494_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_15;
  wire [0:0] h_s_dadda_pg_rca32_and_23_16;
  wire [0:0] h_s_dadda_pg_rca32_and_22_17;
  wire [0:0] h_s_dadda_pg_rca32_fa495_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa495_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_18;
  wire [0:0] h_s_dadda_pg_rca32_and_20_19;
  wire [0:0] h_s_dadda_pg_rca32_and_19_20;
  wire [0:0] h_s_dadda_pg_rca32_fa496_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa496_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_21;
  wire [0:0] h_s_dadda_pg_rca32_and_17_22;
  wire [0:0] h_s_dadda_pg_rca32_and_16_23;
  wire [0:0] h_s_dadda_pg_rca32_fa497_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa497_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_24;
  wire [0:0] h_s_dadda_pg_rca32_and_14_25;
  wire [0:0] h_s_dadda_pg_rca32_and_13_26;
  wire [0:0] h_s_dadda_pg_rca32_fa498_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa498_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_27;
  wire [0:0] h_s_dadda_pg_rca32_and_11_28;
  wire [0:0] h_s_dadda_pg_rca32_and_10_29;
  wire [0:0] h_s_dadda_pg_rca32_fa499_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa499_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_9_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_8_31;
  wire [0:0] h_s_dadda_pg_rca32_fa500_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa500_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa501_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa501_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa502_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa502_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa503_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa503_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa504_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa504_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa505_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa505_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa506_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa506_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa507_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa507_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa508_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa508_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa509_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa509_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa510_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa510_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_9;
  wire [0:0] h_s_dadda_pg_rca32_and_30_10;
  wire [0:0] h_s_dadda_pg_rca32_fa511_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa511_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_11;
  wire [0:0] h_s_dadda_pg_rca32_and_28_12;
  wire [0:0] h_s_dadda_pg_rca32_and_27_13;
  wire [0:0] h_s_dadda_pg_rca32_fa512_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa512_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_14;
  wire [0:0] h_s_dadda_pg_rca32_and_25_15;
  wire [0:0] h_s_dadda_pg_rca32_and_24_16;
  wire [0:0] h_s_dadda_pg_rca32_fa513_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa513_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_17;
  wire [0:0] h_s_dadda_pg_rca32_and_22_18;
  wire [0:0] h_s_dadda_pg_rca32_and_21_19;
  wire [0:0] h_s_dadda_pg_rca32_fa514_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa514_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_20;
  wire [0:0] h_s_dadda_pg_rca32_and_19_21;
  wire [0:0] h_s_dadda_pg_rca32_and_18_22;
  wire [0:0] h_s_dadda_pg_rca32_fa515_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa515_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_23;
  wire [0:0] h_s_dadda_pg_rca32_and_16_24;
  wire [0:0] h_s_dadda_pg_rca32_and_15_25;
  wire [0:0] h_s_dadda_pg_rca32_fa516_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa516_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_26;
  wire [0:0] h_s_dadda_pg_rca32_and_13_27;
  wire [0:0] h_s_dadda_pg_rca32_and_12_28;
  wire [0:0] h_s_dadda_pg_rca32_fa517_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa517_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_11_29;
  wire [0:0] h_s_dadda_pg_rca32_and_10_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_9_31;
  wire [0:0] h_s_dadda_pg_rca32_fa518_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa518_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa519_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa519_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa520_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa520_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa521_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa521_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa522_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa522_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa523_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa523_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa524_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa524_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa525_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa525_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa526_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa526_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa527_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa527_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa528_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa528_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_10;
  wire [0:0] h_s_dadda_pg_rca32_and_30_11;
  wire [0:0] h_s_dadda_pg_rca32_and_29_12;
  wire [0:0] h_s_dadda_pg_rca32_fa529_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa529_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_13;
  wire [0:0] h_s_dadda_pg_rca32_and_27_14;
  wire [0:0] h_s_dadda_pg_rca32_and_26_15;
  wire [0:0] h_s_dadda_pg_rca32_fa530_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa530_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_16;
  wire [0:0] h_s_dadda_pg_rca32_and_24_17;
  wire [0:0] h_s_dadda_pg_rca32_and_23_18;
  wire [0:0] h_s_dadda_pg_rca32_fa531_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa531_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_19;
  wire [0:0] h_s_dadda_pg_rca32_and_21_20;
  wire [0:0] h_s_dadda_pg_rca32_and_20_21;
  wire [0:0] h_s_dadda_pg_rca32_fa532_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa532_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_22;
  wire [0:0] h_s_dadda_pg_rca32_and_18_23;
  wire [0:0] h_s_dadda_pg_rca32_and_17_24;
  wire [0:0] h_s_dadda_pg_rca32_fa533_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa533_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_25;
  wire [0:0] h_s_dadda_pg_rca32_and_15_26;
  wire [0:0] h_s_dadda_pg_rca32_and_14_27;
  wire [0:0] h_s_dadda_pg_rca32_fa534_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa534_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_13_28;
  wire [0:0] h_s_dadda_pg_rca32_and_12_29;
  wire [0:0] h_s_dadda_pg_rca32_and_11_30;
  wire [0:0] h_s_dadda_pg_rca32_fa535_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa535_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_10_31;
  wire [0:0] h_s_dadda_pg_rca32_fa536_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa536_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa537_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa537_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa538_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa538_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa539_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa539_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa540_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa540_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa541_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa541_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa542_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa542_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa543_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa543_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa544_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa544_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_11;
  wire [0:0] h_s_dadda_pg_rca32_fa545_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa545_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_12;
  wire [0:0] h_s_dadda_pg_rca32_and_29_13;
  wire [0:0] h_s_dadda_pg_rca32_and_28_14;
  wire [0:0] h_s_dadda_pg_rca32_fa546_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa546_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_15;
  wire [0:0] h_s_dadda_pg_rca32_and_26_16;
  wire [0:0] h_s_dadda_pg_rca32_and_25_17;
  wire [0:0] h_s_dadda_pg_rca32_fa547_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa547_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_18;
  wire [0:0] h_s_dadda_pg_rca32_and_23_19;
  wire [0:0] h_s_dadda_pg_rca32_and_22_20;
  wire [0:0] h_s_dadda_pg_rca32_fa548_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa548_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_21;
  wire [0:0] h_s_dadda_pg_rca32_and_20_22;
  wire [0:0] h_s_dadda_pg_rca32_and_19_23;
  wire [0:0] h_s_dadda_pg_rca32_fa549_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa549_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_24;
  wire [0:0] h_s_dadda_pg_rca32_and_17_25;
  wire [0:0] h_s_dadda_pg_rca32_and_16_26;
  wire [0:0] h_s_dadda_pg_rca32_fa550_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa550_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_27;
  wire [0:0] h_s_dadda_pg_rca32_and_14_28;
  wire [0:0] h_s_dadda_pg_rca32_and_13_29;
  wire [0:0] h_s_dadda_pg_rca32_fa551_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa551_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_12_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_11_31;
  wire [0:0] h_s_dadda_pg_rca32_fa552_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa552_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa553_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa553_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa554_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa554_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa555_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa555_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa556_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa556_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa557_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa557_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa558_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa558_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa559_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa559_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa560_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa560_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_12;
  wire [0:0] h_s_dadda_pg_rca32_and_30_13;
  wire [0:0] h_s_dadda_pg_rca32_fa561_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa561_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_14;
  wire [0:0] h_s_dadda_pg_rca32_and_28_15;
  wire [0:0] h_s_dadda_pg_rca32_and_27_16;
  wire [0:0] h_s_dadda_pg_rca32_fa562_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa562_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_17;
  wire [0:0] h_s_dadda_pg_rca32_and_25_18;
  wire [0:0] h_s_dadda_pg_rca32_and_24_19;
  wire [0:0] h_s_dadda_pg_rca32_fa563_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa563_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_20;
  wire [0:0] h_s_dadda_pg_rca32_and_22_21;
  wire [0:0] h_s_dadda_pg_rca32_and_21_22;
  wire [0:0] h_s_dadda_pg_rca32_fa564_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa564_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_23;
  wire [0:0] h_s_dadda_pg_rca32_and_19_24;
  wire [0:0] h_s_dadda_pg_rca32_and_18_25;
  wire [0:0] h_s_dadda_pg_rca32_fa565_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa565_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_26;
  wire [0:0] h_s_dadda_pg_rca32_and_16_27;
  wire [0:0] h_s_dadda_pg_rca32_and_15_28;
  wire [0:0] h_s_dadda_pg_rca32_fa566_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa566_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_14_29;
  wire [0:0] h_s_dadda_pg_rca32_and_13_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_12_31;
  wire [0:0] h_s_dadda_pg_rca32_fa567_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa567_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa568_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa568_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa569_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa569_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa570_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa570_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa571_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa571_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa572_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa572_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa573_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa573_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa574_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa574_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa575_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa575_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_13;
  wire [0:0] h_s_dadda_pg_rca32_and_30_14;
  wire [0:0] h_s_dadda_pg_rca32_and_29_15;
  wire [0:0] h_s_dadda_pg_rca32_fa576_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa576_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_16;
  wire [0:0] h_s_dadda_pg_rca32_and_27_17;
  wire [0:0] h_s_dadda_pg_rca32_and_26_18;
  wire [0:0] h_s_dadda_pg_rca32_fa577_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa577_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_19;
  wire [0:0] h_s_dadda_pg_rca32_and_24_20;
  wire [0:0] h_s_dadda_pg_rca32_and_23_21;
  wire [0:0] h_s_dadda_pg_rca32_fa578_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa578_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_22;
  wire [0:0] h_s_dadda_pg_rca32_and_21_23;
  wire [0:0] h_s_dadda_pg_rca32_and_20_24;
  wire [0:0] h_s_dadda_pg_rca32_fa579_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa579_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_25;
  wire [0:0] h_s_dadda_pg_rca32_and_18_26;
  wire [0:0] h_s_dadda_pg_rca32_and_17_27;
  wire [0:0] h_s_dadda_pg_rca32_fa580_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa580_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_16_28;
  wire [0:0] h_s_dadda_pg_rca32_and_15_29;
  wire [0:0] h_s_dadda_pg_rca32_and_14_30;
  wire [0:0] h_s_dadda_pg_rca32_fa581_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa581_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_13_31;
  wire [0:0] h_s_dadda_pg_rca32_fa582_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa582_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa583_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa583_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa584_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa584_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa585_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa585_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa586_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa586_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa587_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa587_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa588_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa588_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_14;
  wire [0:0] h_s_dadda_pg_rca32_fa589_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa589_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_15;
  wire [0:0] h_s_dadda_pg_rca32_and_29_16;
  wire [0:0] h_s_dadda_pg_rca32_and_28_17;
  wire [0:0] h_s_dadda_pg_rca32_fa590_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa590_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_18;
  wire [0:0] h_s_dadda_pg_rca32_and_26_19;
  wire [0:0] h_s_dadda_pg_rca32_and_25_20;
  wire [0:0] h_s_dadda_pg_rca32_fa591_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa591_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_21;
  wire [0:0] h_s_dadda_pg_rca32_and_23_22;
  wire [0:0] h_s_dadda_pg_rca32_and_22_23;
  wire [0:0] h_s_dadda_pg_rca32_fa592_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa592_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_24;
  wire [0:0] h_s_dadda_pg_rca32_and_20_25;
  wire [0:0] h_s_dadda_pg_rca32_and_19_26;
  wire [0:0] h_s_dadda_pg_rca32_fa593_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa593_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_27;
  wire [0:0] h_s_dadda_pg_rca32_and_17_28;
  wire [0:0] h_s_dadda_pg_rca32_and_16_29;
  wire [0:0] h_s_dadda_pg_rca32_fa594_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa594_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_15_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_14_31;
  wire [0:0] h_s_dadda_pg_rca32_fa595_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa595_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa596_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa596_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa597_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa597_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa598_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa598_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa599_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa599_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa600_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa600_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa601_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa601_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_15;
  wire [0:0] h_s_dadda_pg_rca32_and_30_16;
  wire [0:0] h_s_dadda_pg_rca32_fa602_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa602_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_17;
  wire [0:0] h_s_dadda_pg_rca32_and_28_18;
  wire [0:0] h_s_dadda_pg_rca32_and_27_19;
  wire [0:0] h_s_dadda_pg_rca32_fa603_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa603_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_20;
  wire [0:0] h_s_dadda_pg_rca32_and_25_21;
  wire [0:0] h_s_dadda_pg_rca32_and_24_22;
  wire [0:0] h_s_dadda_pg_rca32_fa604_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa604_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_23;
  wire [0:0] h_s_dadda_pg_rca32_and_22_24;
  wire [0:0] h_s_dadda_pg_rca32_and_21_25;
  wire [0:0] h_s_dadda_pg_rca32_fa605_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa605_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_26;
  wire [0:0] h_s_dadda_pg_rca32_and_19_27;
  wire [0:0] h_s_dadda_pg_rca32_and_18_28;
  wire [0:0] h_s_dadda_pg_rca32_fa606_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa606_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_17_29;
  wire [0:0] h_s_dadda_pg_rca32_and_16_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_15_31;
  wire [0:0] h_s_dadda_pg_rca32_fa607_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa607_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa608_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa608_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa609_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa609_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa610_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa610_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa611_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa611_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa612_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa612_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa613_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa613_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_16;
  wire [0:0] h_s_dadda_pg_rca32_and_30_17;
  wire [0:0] h_s_dadda_pg_rca32_and_29_18;
  wire [0:0] h_s_dadda_pg_rca32_fa614_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa614_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_19;
  wire [0:0] h_s_dadda_pg_rca32_and_27_20;
  wire [0:0] h_s_dadda_pg_rca32_and_26_21;
  wire [0:0] h_s_dadda_pg_rca32_fa615_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa615_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_22;
  wire [0:0] h_s_dadda_pg_rca32_and_24_23;
  wire [0:0] h_s_dadda_pg_rca32_and_23_24;
  wire [0:0] h_s_dadda_pg_rca32_fa616_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa616_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_25;
  wire [0:0] h_s_dadda_pg_rca32_and_21_26;
  wire [0:0] h_s_dadda_pg_rca32_and_20_27;
  wire [0:0] h_s_dadda_pg_rca32_fa617_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa617_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_19_28;
  wire [0:0] h_s_dadda_pg_rca32_and_18_29;
  wire [0:0] h_s_dadda_pg_rca32_and_17_30;
  wire [0:0] h_s_dadda_pg_rca32_fa618_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa618_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_16_31;
  wire [0:0] h_s_dadda_pg_rca32_fa619_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa619_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa620_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa620_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa621_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa621_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa622_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa622_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa623_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa623_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_17;
  wire [0:0] h_s_dadda_pg_rca32_fa624_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa624_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_18;
  wire [0:0] h_s_dadda_pg_rca32_and_29_19;
  wire [0:0] h_s_dadda_pg_rca32_and_28_20;
  wire [0:0] h_s_dadda_pg_rca32_fa625_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa625_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_21;
  wire [0:0] h_s_dadda_pg_rca32_and_26_22;
  wire [0:0] h_s_dadda_pg_rca32_and_25_23;
  wire [0:0] h_s_dadda_pg_rca32_fa626_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa626_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_24;
  wire [0:0] h_s_dadda_pg_rca32_and_23_25;
  wire [0:0] h_s_dadda_pg_rca32_and_22_26;
  wire [0:0] h_s_dadda_pg_rca32_fa627_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa627_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_27;
  wire [0:0] h_s_dadda_pg_rca32_and_20_28;
  wire [0:0] h_s_dadda_pg_rca32_and_19_29;
  wire [0:0] h_s_dadda_pg_rca32_fa628_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa628_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_18_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_17_31;
  wire [0:0] h_s_dadda_pg_rca32_fa629_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa629_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa630_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa630_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa631_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa631_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa632_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa632_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa633_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa633_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_18;
  wire [0:0] h_s_dadda_pg_rca32_and_30_19;
  wire [0:0] h_s_dadda_pg_rca32_fa634_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa634_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_20;
  wire [0:0] h_s_dadda_pg_rca32_and_28_21;
  wire [0:0] h_s_dadda_pg_rca32_and_27_22;
  wire [0:0] h_s_dadda_pg_rca32_fa635_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa635_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_23;
  wire [0:0] h_s_dadda_pg_rca32_and_25_24;
  wire [0:0] h_s_dadda_pg_rca32_and_24_25;
  wire [0:0] h_s_dadda_pg_rca32_fa636_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa636_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_26;
  wire [0:0] h_s_dadda_pg_rca32_and_22_27;
  wire [0:0] h_s_dadda_pg_rca32_and_21_28;
  wire [0:0] h_s_dadda_pg_rca32_fa637_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa637_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_20_29;
  wire [0:0] h_s_dadda_pg_rca32_and_19_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_18_31;
  wire [0:0] h_s_dadda_pg_rca32_fa638_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa638_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa639_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa639_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa640_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa640_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa641_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa641_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa642_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa642_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_19;
  wire [0:0] h_s_dadda_pg_rca32_and_30_20;
  wire [0:0] h_s_dadda_pg_rca32_and_29_21;
  wire [0:0] h_s_dadda_pg_rca32_fa643_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa643_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_22;
  wire [0:0] h_s_dadda_pg_rca32_and_27_23;
  wire [0:0] h_s_dadda_pg_rca32_and_26_24;
  wire [0:0] h_s_dadda_pg_rca32_fa644_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa644_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_25;
  wire [0:0] h_s_dadda_pg_rca32_and_24_26;
  wire [0:0] h_s_dadda_pg_rca32_and_23_27;
  wire [0:0] h_s_dadda_pg_rca32_fa645_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa645_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_22_28;
  wire [0:0] h_s_dadda_pg_rca32_and_21_29;
  wire [0:0] h_s_dadda_pg_rca32_and_20_30;
  wire [0:0] h_s_dadda_pg_rca32_fa646_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa646_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_19_31;
  wire [0:0] h_s_dadda_pg_rca32_fa647_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa647_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa648_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa648_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa649_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa649_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_20;
  wire [0:0] h_s_dadda_pg_rca32_fa650_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa650_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_21;
  wire [0:0] h_s_dadda_pg_rca32_and_29_22;
  wire [0:0] h_s_dadda_pg_rca32_and_28_23;
  wire [0:0] h_s_dadda_pg_rca32_fa651_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa651_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_24;
  wire [0:0] h_s_dadda_pg_rca32_and_26_25;
  wire [0:0] h_s_dadda_pg_rca32_and_25_26;
  wire [0:0] h_s_dadda_pg_rca32_fa652_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa652_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_27;
  wire [0:0] h_s_dadda_pg_rca32_and_23_28;
  wire [0:0] h_s_dadda_pg_rca32_and_22_29;
  wire [0:0] h_s_dadda_pg_rca32_fa653_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa653_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_21_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_20_31;
  wire [0:0] h_s_dadda_pg_rca32_fa654_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa654_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa655_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa655_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa656_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa656_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_21;
  wire [0:0] h_s_dadda_pg_rca32_and_30_22;
  wire [0:0] h_s_dadda_pg_rca32_fa657_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa657_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_23;
  wire [0:0] h_s_dadda_pg_rca32_and_28_24;
  wire [0:0] h_s_dadda_pg_rca32_and_27_25;
  wire [0:0] h_s_dadda_pg_rca32_fa658_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa658_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_26;
  wire [0:0] h_s_dadda_pg_rca32_and_25_27;
  wire [0:0] h_s_dadda_pg_rca32_and_24_28;
  wire [0:0] h_s_dadda_pg_rca32_fa659_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa659_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_23_29;
  wire [0:0] h_s_dadda_pg_rca32_and_22_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_21_31;
  wire [0:0] h_s_dadda_pg_rca32_fa660_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa660_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa661_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa661_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa662_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa662_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_22;
  wire [0:0] h_s_dadda_pg_rca32_and_30_23;
  wire [0:0] h_s_dadda_pg_rca32_and_29_24;
  wire [0:0] h_s_dadda_pg_rca32_fa663_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa663_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_25;
  wire [0:0] h_s_dadda_pg_rca32_and_27_26;
  wire [0:0] h_s_dadda_pg_rca32_and_26_27;
  wire [0:0] h_s_dadda_pg_rca32_fa664_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa664_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_28;
  wire [0:0] h_s_dadda_pg_rca32_and_24_29;
  wire [0:0] h_s_dadda_pg_rca32_and_23_30;
  wire [0:0] h_s_dadda_pg_rca32_fa665_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa665_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa666_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa666_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_23;
  wire [0:0] h_s_dadda_pg_rca32_fa667_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa667_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_24;
  wire [0:0] h_s_dadda_pg_rca32_and_29_25;
  wire [0:0] h_s_dadda_pg_rca32_and_28_26;
  wire [0:0] h_s_dadda_pg_rca32_fa668_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa668_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_27;
  wire [0:0] h_s_dadda_pg_rca32_and_26_28;
  wire [0:0] h_s_dadda_pg_rca32_and_25_29;
  wire [0:0] h_s_dadda_pg_rca32_fa669_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa669_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa670_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa670_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_24;
  wire [0:0] h_s_dadda_pg_rca32_and_30_25;
  wire [0:0] h_s_dadda_pg_rca32_fa671_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa671_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_26;
  wire [0:0] h_s_dadda_pg_rca32_and_28_27;
  wire [0:0] h_s_dadda_pg_rca32_and_27_28;
  wire [0:0] h_s_dadda_pg_rca32_fa672_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa672_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa673_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa673_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_25;
  wire [0:0] h_s_dadda_pg_rca32_and_30_26;
  wire [0:0] h_s_dadda_pg_rca32_and_29_27;
  wire [0:0] h_s_dadda_pg_rca32_fa674_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa674_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_26;
  wire [0:0] h_s_dadda_pg_rca32_fa675_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa675_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_1;
  wire [0:0] h_s_dadda_pg_rca32_ha26_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha26_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_5_0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_1;
  wire [0:0] h_s_dadda_pg_rca32_fa676_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa676_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_2;
  wire [0:0] h_s_dadda_pg_rca32_and_2_3;
  wire [0:0] h_s_dadda_pg_rca32_ha27_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha27_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_4_2;
  wire [0:0] h_s_dadda_pg_rca32_fa677_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa677_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_3;
  wire [0:0] h_s_dadda_pg_rca32_and_2_4;
  wire [0:0] h_s_dadda_pg_rca32_and_1_5;
  wire [0:0] h_s_dadda_pg_rca32_fa678_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa678_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_4;
  wire [0:0] h_s_dadda_pg_rca32_fa679_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa679_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_5;
  wire [0:0] h_s_dadda_pg_rca32_and_1_6;
  wire [0:0] h_s_dadda_pg_rca32_and_0_7;
  wire [0:0] h_s_dadda_pg_rca32_fa680_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa680_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_6;
  wire [0:0] h_s_dadda_pg_rca32_fa681_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa681_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_7;
  wire [0:0] h_s_dadda_pg_rca32_and_0_8;
  wire [0:0] h_s_dadda_pg_rca32_fa682_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa682_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_8;
  wire [0:0] h_s_dadda_pg_rca32_fa683_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa683_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_9;
  wire [0:0] h_s_dadda_pg_rca32_fa684_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa684_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_10;
  wire [0:0] h_s_dadda_pg_rca32_fa685_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa685_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa686_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa686_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa687_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa687_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa688_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa688_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa689_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa689_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa690_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa690_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa691_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa691_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa692_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa692_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa693_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa693_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa694_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa694_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa695_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa695_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa696_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa696_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa697_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa697_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa698_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa698_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa699_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa699_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa700_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa700_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa701_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa701_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa702_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa702_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa703_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa703_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa704_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa704_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa705_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa705_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa706_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa706_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa707_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa707_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa708_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa708_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa709_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa709_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa710_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa710_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa711_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa711_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa712_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa712_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa713_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa713_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa714_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa714_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa715_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa715_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa716_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa716_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa717_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa717_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa718_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa718_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa719_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa719_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa720_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa720_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa721_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa721_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa722_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa722_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa723_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa723_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa724_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa724_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa725_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa725_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa726_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa726_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa727_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa727_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa728_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa728_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa729_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa729_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa730_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa730_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa731_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa731_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa732_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa732_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa733_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa733_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa734_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa734_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa735_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa735_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa736_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa736_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa737_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa737_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa738_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa738_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa739_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa739_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa740_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa740_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa741_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa741_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa742_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa742_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa743_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa743_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa744_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa744_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa745_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa745_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa746_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa746_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa747_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa747_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa748_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa748_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa749_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa749_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa750_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa750_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa751_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa751_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa752_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa752_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa753_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa753_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa754_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa754_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa755_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa755_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa756_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa756_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa757_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa757_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa758_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa758_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa759_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa759_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa760_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa760_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa761_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa761_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa762_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa762_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa763_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa763_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa764_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa764_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa765_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa765_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa766_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa766_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa767_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa767_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa768_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa768_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa769_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa769_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa770_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa770_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_22_31;
  wire [0:0] h_s_dadda_pg_rca32_fa771_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa771_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa772_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa772_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_24_30;
  wire [0:0] h_s_dadda_pg_rca32_fa773_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa773_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_23_31;
  wire [0:0] h_s_dadda_pg_rca32_fa774_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa774_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_26_29;
  wire [0:0] h_s_dadda_pg_rca32_fa775_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa775_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_25_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_24_31;
  wire [0:0] h_s_dadda_pg_rca32_fa776_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa776_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_28;
  wire [0:0] h_s_dadda_pg_rca32_fa777_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa777_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_27_29;
  wire [0:0] h_s_dadda_pg_rca32_and_26_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_25_31;
  wire [0:0] h_s_dadda_pg_rca32_fa778_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa778_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_27;
  wire [0:0] h_s_dadda_pg_rca32_fa779_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa779_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_29_28;
  wire [0:0] h_s_dadda_pg_rca32_and_28_29;
  wire [0:0] h_s_dadda_pg_rca32_and_27_30;
  wire [0:0] h_s_dadda_pg_rca32_fa780_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa780_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa781_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa781_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_27;
  wire [0:0] h_s_dadda_pg_rca32_and_30_28;
  wire [0:0] h_s_dadda_pg_rca32_and_29_29;
  wire [0:0] h_s_dadda_pg_rca32_fa782_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa782_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_28;
  wire [0:0] h_s_dadda_pg_rca32_fa783_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa783_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_3_0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_1;
  wire [0:0] h_s_dadda_pg_rca32_ha28_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha28_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_2;
  wire [0:0] h_s_dadda_pg_rca32_and_1_3;
  wire [0:0] h_s_dadda_pg_rca32_fa784_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa784_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_4;
  wire [0:0] h_s_dadda_pg_rca32_and_0_5;
  wire [0:0] h_s_dadda_pg_rca32_fa785_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa785_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_6;
  wire [0:0] h_s_dadda_pg_rca32_fa786_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa786_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa787_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa787_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa788_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa788_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa789_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa789_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa790_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa790_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa791_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa791_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa792_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa792_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa793_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa793_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa794_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa794_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa795_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa795_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa796_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa796_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa797_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa797_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa798_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa798_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa799_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa799_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa800_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa800_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa801_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa801_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa802_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa802_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa803_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa803_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa804_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa804_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa805_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa805_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa806_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa806_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa807_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa807_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa808_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa808_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa809_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa809_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa810_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa810_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa811_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa811_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa812_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa812_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa813_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa813_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa814_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa814_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa815_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa815_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa816_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa816_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa817_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa817_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa818_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa818_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa819_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa819_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa820_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa820_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa821_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa821_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa822_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa822_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa823_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa823_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa824_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa824_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa825_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa825_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa826_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa826_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa827_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa827_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa828_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa828_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa829_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa829_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa830_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa830_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa831_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa831_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa832_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa832_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa833_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa833_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa834_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa834_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa835_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa835_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa836_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa836_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_26_31;
  wire [0:0] h_s_dadda_pg_rca32_fa837_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa837_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_28_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_27_31;
  wire [0:0] h_s_dadda_pg_rca32_fa838_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa838_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_29;
  wire [0:0] h_s_dadda_pg_rca32_and_29_30;
  wire [0:0] h_s_dadda_pg_rca32_fa839_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa839_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_29;
  wire [0:0] h_s_dadda_pg_rca32_fa840_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa840_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_2_0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_1;
  wire [0:0] h_s_dadda_pg_rca32_ha29_xor0;
  wire [0:0] h_s_dadda_pg_rca32_ha29_and0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_2;
  wire [0:0] h_s_dadda_pg_rca32_and_0_3;
  wire [0:0] h_s_dadda_pg_rca32_fa841_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa841_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_4;
  wire [0:0] h_s_dadda_pg_rca32_fa842_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa842_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa843_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa843_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa844_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa844_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa845_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa845_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa846_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa846_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa847_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa847_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa848_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa848_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa849_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa849_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa850_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa850_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa851_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa851_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa852_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa852_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa853_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa853_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa854_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa854_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa855_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa855_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa856_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa856_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa857_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa857_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa858_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa858_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa859_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa859_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa860_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa860_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa861_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa861_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa862_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa862_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa863_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa863_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa864_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa864_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa865_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa865_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa866_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa866_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa867_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa867_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa868_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa868_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa869_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa869_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa870_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa870_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa871_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa871_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa872_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa872_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa873_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa873_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa874_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa874_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa875_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa875_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa876_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa876_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa877_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa877_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa878_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa878_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa879_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa879_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa880_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa880_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa881_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa881_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa882_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa882_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa883_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa883_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa884_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa884_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa885_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa885_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa886_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa886_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa887_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa887_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa888_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa888_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa889_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa889_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa890_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa890_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa891_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa891_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa892_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa892_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa893_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa893_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa894_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa894_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa895_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa895_or0;
  wire [0:0] h_s_dadda_pg_rca32_fa896_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa896_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_28_31;
  wire [0:0] h_s_dadda_pg_rca32_fa897_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa897_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_30_30;
  wire [0:0] h_s_dadda_pg_rca32_nand_29_31;
  wire [0:0] h_s_dadda_pg_rca32_fa898_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa898_or0;
  wire [0:0] h_s_dadda_pg_rca32_nand_31_30;
  wire [0:0] h_s_dadda_pg_rca32_fa899_xor1;
  wire [0:0] h_s_dadda_pg_rca32_fa899_or0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_0;
  wire [0:0] h_s_dadda_pg_rca32_and_1_0;
  wire [0:0] h_s_dadda_pg_rca32_and_0_2;
  wire [0:0] h_s_dadda_pg_rca32_nand_30_31;
  wire [0:0] h_s_dadda_pg_rca32_and_0_1;
  wire [0:0] h_s_dadda_pg_rca32_and_31_31;
  wire [61:0] h_s_dadda_pg_rca32_u_pg_rca62_a;
  wire [61:0] h_s_dadda_pg_rca32_u_pg_rca62_b;
  wire [62:0] h_s_dadda_pg_rca32_u_pg_rca62_out;
  wire [0:0] h_s_dadda_pg_rca32_xor0;

  and_gate and_gate_h_s_dadda_pg_rca32_and_28_0(a[28], b[0], h_s_dadda_pg_rca32_and_28_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_1(a[27], b[1], h_s_dadda_pg_rca32_and_27_1);
  ha ha_h_s_dadda_pg_rca32_ha0_out(h_s_dadda_pg_rca32_and_28_0[0], h_s_dadda_pg_rca32_and_27_1[0], h_s_dadda_pg_rca32_ha0_xor0, h_s_dadda_pg_rca32_ha0_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_0(a[29], b[0], h_s_dadda_pg_rca32_and_29_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_1(a[28], b[1], h_s_dadda_pg_rca32_and_28_1);
  fa fa_h_s_dadda_pg_rca32_fa0_out(h_s_dadda_pg_rca32_ha0_and0[0], h_s_dadda_pg_rca32_and_29_0[0], h_s_dadda_pg_rca32_and_28_1[0], h_s_dadda_pg_rca32_fa0_xor1, h_s_dadda_pg_rca32_fa0_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_2(a[27], b[2], h_s_dadda_pg_rca32_and_27_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_3(a[26], b[3], h_s_dadda_pg_rca32_and_26_3);
  ha ha_h_s_dadda_pg_rca32_ha1_out(h_s_dadda_pg_rca32_and_27_2[0], h_s_dadda_pg_rca32_and_26_3[0], h_s_dadda_pg_rca32_ha1_xor0, h_s_dadda_pg_rca32_ha1_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_0(a[30], b[0], h_s_dadda_pg_rca32_and_30_0);
  fa fa_h_s_dadda_pg_rca32_fa1_out(h_s_dadda_pg_rca32_ha1_and0[0], h_s_dadda_pg_rca32_fa0_or0[0], h_s_dadda_pg_rca32_and_30_0[0], h_s_dadda_pg_rca32_fa1_xor1, h_s_dadda_pg_rca32_fa1_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_1(a[29], b[1], h_s_dadda_pg_rca32_and_29_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_2(a[28], b[2], h_s_dadda_pg_rca32_and_28_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_3(a[27], b[3], h_s_dadda_pg_rca32_and_27_3);
  fa fa_h_s_dadda_pg_rca32_fa2_out(h_s_dadda_pg_rca32_and_29_1[0], h_s_dadda_pg_rca32_and_28_2[0], h_s_dadda_pg_rca32_and_27_3[0], h_s_dadda_pg_rca32_fa2_xor1, h_s_dadda_pg_rca32_fa2_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_4(a[26], b[4], h_s_dadda_pg_rca32_and_26_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_5(a[25], b[5], h_s_dadda_pg_rca32_and_25_5);
  ha ha_h_s_dadda_pg_rca32_ha2_out(h_s_dadda_pg_rca32_and_26_4[0], h_s_dadda_pg_rca32_and_25_5[0], h_s_dadda_pg_rca32_ha2_xor0, h_s_dadda_pg_rca32_ha2_and0);
  fa fa_h_s_dadda_pg_rca32_fa3_out(h_s_dadda_pg_rca32_ha2_and0[0], h_s_dadda_pg_rca32_fa2_or0[0], h_s_dadda_pg_rca32_fa1_or0[0], h_s_dadda_pg_rca32_fa3_xor1, h_s_dadda_pg_rca32_fa3_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_0(a[31], b[0], h_s_dadda_pg_rca32_nand_31_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_1(a[30], b[1], h_s_dadda_pg_rca32_and_30_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_2(a[29], b[2], h_s_dadda_pg_rca32_and_29_2);
  fa fa_h_s_dadda_pg_rca32_fa4_out(h_s_dadda_pg_rca32_nand_31_0[0], h_s_dadda_pg_rca32_and_30_1[0], h_s_dadda_pg_rca32_and_29_2[0], h_s_dadda_pg_rca32_fa4_xor1, h_s_dadda_pg_rca32_fa4_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_3(a[28], b[3], h_s_dadda_pg_rca32_and_28_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_4(a[27], b[4], h_s_dadda_pg_rca32_and_27_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_5(a[26], b[5], h_s_dadda_pg_rca32_and_26_5);
  fa fa_h_s_dadda_pg_rca32_fa5_out(h_s_dadda_pg_rca32_and_28_3[0], h_s_dadda_pg_rca32_and_27_4[0], h_s_dadda_pg_rca32_and_26_5[0], h_s_dadda_pg_rca32_fa5_xor1, h_s_dadda_pg_rca32_fa5_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_6(a[25], b[6], h_s_dadda_pg_rca32_and_25_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_7(a[24], b[7], h_s_dadda_pg_rca32_and_24_7);
  ha ha_h_s_dadda_pg_rca32_ha3_out(h_s_dadda_pg_rca32_and_25_6[0], h_s_dadda_pg_rca32_and_24_7[0], h_s_dadda_pg_rca32_ha3_xor0, h_s_dadda_pg_rca32_ha3_and0);
  fa fa_h_s_dadda_pg_rca32_fa6_out(h_s_dadda_pg_rca32_ha3_and0[0], h_s_dadda_pg_rca32_fa5_or0[0], h_s_dadda_pg_rca32_fa4_or0[0], h_s_dadda_pg_rca32_fa6_xor1, h_s_dadda_pg_rca32_fa6_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_1(a[31], b[1], h_s_dadda_pg_rca32_nand_31_1);
  fa fa_h_s_dadda_pg_rca32_fa7_out(h_s_dadda_pg_rca32_fa3_or0[0], 1'b1, h_s_dadda_pg_rca32_nand_31_1[0], h_s_dadda_pg_rca32_fa7_xor1, h_s_dadda_pg_rca32_fa7_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_2(a[30], b[2], h_s_dadda_pg_rca32_and_30_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_3(a[29], b[3], h_s_dadda_pg_rca32_and_29_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_4(a[28], b[4], h_s_dadda_pg_rca32_and_28_4);
  fa fa_h_s_dadda_pg_rca32_fa8_out(h_s_dadda_pg_rca32_and_30_2[0], h_s_dadda_pg_rca32_and_29_3[0], h_s_dadda_pg_rca32_and_28_4[0], h_s_dadda_pg_rca32_fa8_xor1, h_s_dadda_pg_rca32_fa8_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_5(a[27], b[5], h_s_dadda_pg_rca32_and_27_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_6(a[26], b[6], h_s_dadda_pg_rca32_and_26_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_7(a[25], b[7], h_s_dadda_pg_rca32_and_25_7);
  fa fa_h_s_dadda_pg_rca32_fa9_out(h_s_dadda_pg_rca32_and_27_5[0], h_s_dadda_pg_rca32_and_26_6[0], h_s_dadda_pg_rca32_and_25_7[0], h_s_dadda_pg_rca32_fa9_xor1, h_s_dadda_pg_rca32_fa9_or0);
  fa fa_h_s_dadda_pg_rca32_fa10_out(h_s_dadda_pg_rca32_fa9_or0[0], h_s_dadda_pg_rca32_fa8_or0[0], h_s_dadda_pg_rca32_fa7_or0[0], h_s_dadda_pg_rca32_fa10_xor1, h_s_dadda_pg_rca32_fa10_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_2(a[31], b[2], h_s_dadda_pg_rca32_nand_31_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_3(a[30], b[3], h_s_dadda_pg_rca32_and_30_3);
  fa fa_h_s_dadda_pg_rca32_fa11_out(h_s_dadda_pg_rca32_fa6_or0[0], h_s_dadda_pg_rca32_nand_31_2[0], h_s_dadda_pg_rca32_and_30_3[0], h_s_dadda_pg_rca32_fa11_xor1, h_s_dadda_pg_rca32_fa11_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_4(a[29], b[4], h_s_dadda_pg_rca32_and_29_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_5(a[28], b[5], h_s_dadda_pg_rca32_and_28_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_6(a[27], b[6], h_s_dadda_pg_rca32_and_27_6);
  fa fa_h_s_dadda_pg_rca32_fa12_out(h_s_dadda_pg_rca32_and_29_4[0], h_s_dadda_pg_rca32_and_28_5[0], h_s_dadda_pg_rca32_and_27_6[0], h_s_dadda_pg_rca32_fa12_xor1, h_s_dadda_pg_rca32_fa12_or0);
  fa fa_h_s_dadda_pg_rca32_fa13_out(h_s_dadda_pg_rca32_fa12_or0[0], h_s_dadda_pg_rca32_fa11_or0[0], h_s_dadda_pg_rca32_fa10_or0[0], h_s_dadda_pg_rca32_fa13_xor1, h_s_dadda_pg_rca32_fa13_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_3(a[31], b[3], h_s_dadda_pg_rca32_nand_31_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_4(a[30], b[4], h_s_dadda_pg_rca32_and_30_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_5(a[29], b[5], h_s_dadda_pg_rca32_and_29_5);
  fa fa_h_s_dadda_pg_rca32_fa14_out(h_s_dadda_pg_rca32_nand_31_3[0], h_s_dadda_pg_rca32_and_30_4[0], h_s_dadda_pg_rca32_and_29_5[0], h_s_dadda_pg_rca32_fa14_xor1, h_s_dadda_pg_rca32_fa14_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_4(a[31], b[4], h_s_dadda_pg_rca32_nand_31_4);
  fa fa_h_s_dadda_pg_rca32_fa15_out(h_s_dadda_pg_rca32_fa14_or0[0], h_s_dadda_pg_rca32_fa13_or0[0], h_s_dadda_pg_rca32_nand_31_4[0], h_s_dadda_pg_rca32_fa15_xor1, h_s_dadda_pg_rca32_fa15_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_0(a[6], b[0], h_s_dadda_pg_rca32_and_6_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_1(a[5], b[1], h_s_dadda_pg_rca32_and_5_1);
  ha ha_h_s_dadda_pg_rca32_ha4_out(h_s_dadda_pg_rca32_and_6_0[0], h_s_dadda_pg_rca32_and_5_1[0], h_s_dadda_pg_rca32_ha4_xor0, h_s_dadda_pg_rca32_ha4_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_0(a[7], b[0], h_s_dadda_pg_rca32_and_7_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_1(a[6], b[1], h_s_dadda_pg_rca32_and_6_1);
  fa fa_h_s_dadda_pg_rca32_fa16_out(h_s_dadda_pg_rca32_ha4_and0[0], h_s_dadda_pg_rca32_and_7_0[0], h_s_dadda_pg_rca32_and_6_1[0], h_s_dadda_pg_rca32_fa16_xor1, h_s_dadda_pg_rca32_fa16_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_2(a[5], b[2], h_s_dadda_pg_rca32_and_5_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_3(a[4], b[3], h_s_dadda_pg_rca32_and_4_3);
  ha ha_h_s_dadda_pg_rca32_ha5_out(h_s_dadda_pg_rca32_and_5_2[0], h_s_dadda_pg_rca32_and_4_3[0], h_s_dadda_pg_rca32_ha5_xor0, h_s_dadda_pg_rca32_ha5_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_0(a[8], b[0], h_s_dadda_pg_rca32_and_8_0);
  fa fa_h_s_dadda_pg_rca32_fa17_out(h_s_dadda_pg_rca32_ha5_and0[0], h_s_dadda_pg_rca32_fa16_or0[0], h_s_dadda_pg_rca32_and_8_0[0], h_s_dadda_pg_rca32_fa17_xor1, h_s_dadda_pg_rca32_fa17_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_1(a[7], b[1], h_s_dadda_pg_rca32_and_7_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_2(a[6], b[2], h_s_dadda_pg_rca32_and_6_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_3(a[5], b[3], h_s_dadda_pg_rca32_and_5_3);
  fa fa_h_s_dadda_pg_rca32_fa18_out(h_s_dadda_pg_rca32_and_7_1[0], h_s_dadda_pg_rca32_and_6_2[0], h_s_dadda_pg_rca32_and_5_3[0], h_s_dadda_pg_rca32_fa18_xor1, h_s_dadda_pg_rca32_fa18_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_4(a[4], b[4], h_s_dadda_pg_rca32_and_4_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_5(a[3], b[5], h_s_dadda_pg_rca32_and_3_5);
  ha ha_h_s_dadda_pg_rca32_ha6_out(h_s_dadda_pg_rca32_and_4_4[0], h_s_dadda_pg_rca32_and_3_5[0], h_s_dadda_pg_rca32_ha6_xor0, h_s_dadda_pg_rca32_ha6_and0);
  fa fa_h_s_dadda_pg_rca32_fa19_out(h_s_dadda_pg_rca32_ha6_and0[0], h_s_dadda_pg_rca32_fa18_or0[0], h_s_dadda_pg_rca32_fa17_or0[0], h_s_dadda_pg_rca32_fa19_xor1, h_s_dadda_pg_rca32_fa19_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_0(a[9], b[0], h_s_dadda_pg_rca32_and_9_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_1(a[8], b[1], h_s_dadda_pg_rca32_and_8_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_2(a[7], b[2], h_s_dadda_pg_rca32_and_7_2);
  fa fa_h_s_dadda_pg_rca32_fa20_out(h_s_dadda_pg_rca32_and_9_0[0], h_s_dadda_pg_rca32_and_8_1[0], h_s_dadda_pg_rca32_and_7_2[0], h_s_dadda_pg_rca32_fa20_xor1, h_s_dadda_pg_rca32_fa20_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_3(a[6], b[3], h_s_dadda_pg_rca32_and_6_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_4(a[5], b[4], h_s_dadda_pg_rca32_and_5_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_5(a[4], b[5], h_s_dadda_pg_rca32_and_4_5);
  fa fa_h_s_dadda_pg_rca32_fa21_out(h_s_dadda_pg_rca32_and_6_3[0], h_s_dadda_pg_rca32_and_5_4[0], h_s_dadda_pg_rca32_and_4_5[0], h_s_dadda_pg_rca32_fa21_xor1, h_s_dadda_pg_rca32_fa21_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_6(a[3], b[6], h_s_dadda_pg_rca32_and_3_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_7(a[2], b[7], h_s_dadda_pg_rca32_and_2_7);
  ha ha_h_s_dadda_pg_rca32_ha7_out(h_s_dadda_pg_rca32_and_3_6[0], h_s_dadda_pg_rca32_and_2_7[0], h_s_dadda_pg_rca32_ha7_xor0, h_s_dadda_pg_rca32_ha7_and0);
  fa fa_h_s_dadda_pg_rca32_fa22_out(h_s_dadda_pg_rca32_ha7_and0[0], h_s_dadda_pg_rca32_fa21_or0[0], h_s_dadda_pg_rca32_fa20_or0[0], h_s_dadda_pg_rca32_fa22_xor1, h_s_dadda_pg_rca32_fa22_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_0(a[10], b[0], h_s_dadda_pg_rca32_and_10_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_1(a[9], b[1], h_s_dadda_pg_rca32_and_9_1);
  fa fa_h_s_dadda_pg_rca32_fa23_out(h_s_dadda_pg_rca32_fa19_or0[0], h_s_dadda_pg_rca32_and_10_0[0], h_s_dadda_pg_rca32_and_9_1[0], h_s_dadda_pg_rca32_fa23_xor1, h_s_dadda_pg_rca32_fa23_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_2(a[8], b[2], h_s_dadda_pg_rca32_and_8_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_3(a[7], b[3], h_s_dadda_pg_rca32_and_7_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_4(a[6], b[4], h_s_dadda_pg_rca32_and_6_4);
  fa fa_h_s_dadda_pg_rca32_fa24_out(h_s_dadda_pg_rca32_and_8_2[0], h_s_dadda_pg_rca32_and_7_3[0], h_s_dadda_pg_rca32_and_6_4[0], h_s_dadda_pg_rca32_fa24_xor1, h_s_dadda_pg_rca32_fa24_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_5(a[5], b[5], h_s_dadda_pg_rca32_and_5_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_6(a[4], b[6], h_s_dadda_pg_rca32_and_4_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_7(a[3], b[7], h_s_dadda_pg_rca32_and_3_7);
  fa fa_h_s_dadda_pg_rca32_fa25_out(h_s_dadda_pg_rca32_and_5_5[0], h_s_dadda_pg_rca32_and_4_6[0], h_s_dadda_pg_rca32_and_3_7[0], h_s_dadda_pg_rca32_fa25_xor1, h_s_dadda_pg_rca32_fa25_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_8(a[2], b[8], h_s_dadda_pg_rca32_and_2_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_9(a[1], b[9], h_s_dadda_pg_rca32_and_1_9);
  ha ha_h_s_dadda_pg_rca32_ha8_out(h_s_dadda_pg_rca32_and_2_8[0], h_s_dadda_pg_rca32_and_1_9[0], h_s_dadda_pg_rca32_ha8_xor0, h_s_dadda_pg_rca32_ha8_and0);
  fa fa_h_s_dadda_pg_rca32_fa26_out(h_s_dadda_pg_rca32_ha8_and0[0], h_s_dadda_pg_rca32_fa25_or0[0], h_s_dadda_pg_rca32_fa24_or0[0], h_s_dadda_pg_rca32_fa26_xor1, h_s_dadda_pg_rca32_fa26_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_0(a[11], b[0], h_s_dadda_pg_rca32_and_11_0);
  fa fa_h_s_dadda_pg_rca32_fa27_out(h_s_dadda_pg_rca32_fa23_or0[0], h_s_dadda_pg_rca32_fa22_or0[0], h_s_dadda_pg_rca32_and_11_0[0], h_s_dadda_pg_rca32_fa27_xor1, h_s_dadda_pg_rca32_fa27_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_1(a[10], b[1], h_s_dadda_pg_rca32_and_10_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_2(a[9], b[2], h_s_dadda_pg_rca32_and_9_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_3(a[8], b[3], h_s_dadda_pg_rca32_and_8_3);
  fa fa_h_s_dadda_pg_rca32_fa28_out(h_s_dadda_pg_rca32_and_10_1[0], h_s_dadda_pg_rca32_and_9_2[0], h_s_dadda_pg_rca32_and_8_3[0], h_s_dadda_pg_rca32_fa28_xor1, h_s_dadda_pg_rca32_fa28_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_4(a[7], b[4], h_s_dadda_pg_rca32_and_7_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_5(a[6], b[5], h_s_dadda_pg_rca32_and_6_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_6(a[5], b[6], h_s_dadda_pg_rca32_and_5_6);
  fa fa_h_s_dadda_pg_rca32_fa29_out(h_s_dadda_pg_rca32_and_7_4[0], h_s_dadda_pg_rca32_and_6_5[0], h_s_dadda_pg_rca32_and_5_6[0], h_s_dadda_pg_rca32_fa29_xor1, h_s_dadda_pg_rca32_fa29_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_7(a[4], b[7], h_s_dadda_pg_rca32_and_4_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_8(a[3], b[8], h_s_dadda_pg_rca32_and_3_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_9(a[2], b[9], h_s_dadda_pg_rca32_and_2_9);
  fa fa_h_s_dadda_pg_rca32_fa30_out(h_s_dadda_pg_rca32_and_4_7[0], h_s_dadda_pg_rca32_and_3_8[0], h_s_dadda_pg_rca32_and_2_9[0], h_s_dadda_pg_rca32_fa30_xor1, h_s_dadda_pg_rca32_fa30_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_10(a[1], b[10], h_s_dadda_pg_rca32_and_1_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_11(a[0], b[11], h_s_dadda_pg_rca32_and_0_11);
  ha ha_h_s_dadda_pg_rca32_ha9_out(h_s_dadda_pg_rca32_and_1_10[0], h_s_dadda_pg_rca32_and_0_11[0], h_s_dadda_pg_rca32_ha9_xor0, h_s_dadda_pg_rca32_ha9_and0);
  fa fa_h_s_dadda_pg_rca32_fa31_out(h_s_dadda_pg_rca32_ha9_and0[0], h_s_dadda_pg_rca32_fa30_or0[0], h_s_dadda_pg_rca32_fa29_or0[0], h_s_dadda_pg_rca32_fa31_xor1, h_s_dadda_pg_rca32_fa31_or0);
  fa fa_h_s_dadda_pg_rca32_fa32_out(h_s_dadda_pg_rca32_fa28_or0[0], h_s_dadda_pg_rca32_fa27_or0[0], h_s_dadda_pg_rca32_fa26_or0[0], h_s_dadda_pg_rca32_fa32_xor1, h_s_dadda_pg_rca32_fa32_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_0(a[12], b[0], h_s_dadda_pg_rca32_and_12_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_1(a[11], b[1], h_s_dadda_pg_rca32_and_11_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_2(a[10], b[2], h_s_dadda_pg_rca32_and_10_2);
  fa fa_h_s_dadda_pg_rca32_fa33_out(h_s_dadda_pg_rca32_and_12_0[0], h_s_dadda_pg_rca32_and_11_1[0], h_s_dadda_pg_rca32_and_10_2[0], h_s_dadda_pg_rca32_fa33_xor1, h_s_dadda_pg_rca32_fa33_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_3(a[9], b[3], h_s_dadda_pg_rca32_and_9_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_4(a[8], b[4], h_s_dadda_pg_rca32_and_8_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_5(a[7], b[5], h_s_dadda_pg_rca32_and_7_5);
  fa fa_h_s_dadda_pg_rca32_fa34_out(h_s_dadda_pg_rca32_and_9_3[0], h_s_dadda_pg_rca32_and_8_4[0], h_s_dadda_pg_rca32_and_7_5[0], h_s_dadda_pg_rca32_fa34_xor1, h_s_dadda_pg_rca32_fa34_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_6(a[6], b[6], h_s_dadda_pg_rca32_and_6_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_7(a[5], b[7], h_s_dadda_pg_rca32_and_5_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_8(a[4], b[8], h_s_dadda_pg_rca32_and_4_8);
  fa fa_h_s_dadda_pg_rca32_fa35_out(h_s_dadda_pg_rca32_and_6_6[0], h_s_dadda_pg_rca32_and_5_7[0], h_s_dadda_pg_rca32_and_4_8[0], h_s_dadda_pg_rca32_fa35_xor1, h_s_dadda_pg_rca32_fa35_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_9(a[3], b[9], h_s_dadda_pg_rca32_and_3_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_10(a[2], b[10], h_s_dadda_pg_rca32_and_2_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_11(a[1], b[11], h_s_dadda_pg_rca32_and_1_11);
  fa fa_h_s_dadda_pg_rca32_fa36_out(h_s_dadda_pg_rca32_and_3_9[0], h_s_dadda_pg_rca32_and_2_10[0], h_s_dadda_pg_rca32_and_1_11[0], h_s_dadda_pg_rca32_fa36_xor1, h_s_dadda_pg_rca32_fa36_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_12(a[0], b[12], h_s_dadda_pg_rca32_and_0_12);
  ha ha_h_s_dadda_pg_rca32_ha10_out(h_s_dadda_pg_rca32_and_0_12[0], h_s_dadda_pg_rca32_fa31_xor1[0], h_s_dadda_pg_rca32_ha10_xor0, h_s_dadda_pg_rca32_ha10_and0);
  fa fa_h_s_dadda_pg_rca32_fa37_out(h_s_dadda_pg_rca32_ha10_and0[0], h_s_dadda_pg_rca32_fa36_or0[0], h_s_dadda_pg_rca32_fa35_or0[0], h_s_dadda_pg_rca32_fa37_xor1, h_s_dadda_pg_rca32_fa37_or0);
  fa fa_h_s_dadda_pg_rca32_fa38_out(h_s_dadda_pg_rca32_fa34_or0[0], h_s_dadda_pg_rca32_fa33_or0[0], h_s_dadda_pg_rca32_fa32_or0[0], h_s_dadda_pg_rca32_fa38_xor1, h_s_dadda_pg_rca32_fa38_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_0(a[13], b[0], h_s_dadda_pg_rca32_and_13_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_1(a[12], b[1], h_s_dadda_pg_rca32_and_12_1);
  fa fa_h_s_dadda_pg_rca32_fa39_out(h_s_dadda_pg_rca32_fa31_or0[0], h_s_dadda_pg_rca32_and_13_0[0], h_s_dadda_pg_rca32_and_12_1[0], h_s_dadda_pg_rca32_fa39_xor1, h_s_dadda_pg_rca32_fa39_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_2(a[11], b[2], h_s_dadda_pg_rca32_and_11_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_3(a[10], b[3], h_s_dadda_pg_rca32_and_10_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_4(a[9], b[4], h_s_dadda_pg_rca32_and_9_4);
  fa fa_h_s_dadda_pg_rca32_fa40_out(h_s_dadda_pg_rca32_and_11_2[0], h_s_dadda_pg_rca32_and_10_3[0], h_s_dadda_pg_rca32_and_9_4[0], h_s_dadda_pg_rca32_fa40_xor1, h_s_dadda_pg_rca32_fa40_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_5(a[8], b[5], h_s_dadda_pg_rca32_and_8_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_6(a[7], b[6], h_s_dadda_pg_rca32_and_7_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_7(a[6], b[7], h_s_dadda_pg_rca32_and_6_7);
  fa fa_h_s_dadda_pg_rca32_fa41_out(h_s_dadda_pg_rca32_and_8_5[0], h_s_dadda_pg_rca32_and_7_6[0], h_s_dadda_pg_rca32_and_6_7[0], h_s_dadda_pg_rca32_fa41_xor1, h_s_dadda_pg_rca32_fa41_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_8(a[5], b[8], h_s_dadda_pg_rca32_and_5_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_9(a[4], b[9], h_s_dadda_pg_rca32_and_4_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_10(a[3], b[10], h_s_dadda_pg_rca32_and_3_10);
  fa fa_h_s_dadda_pg_rca32_fa42_out(h_s_dadda_pg_rca32_and_5_8[0], h_s_dadda_pg_rca32_and_4_9[0], h_s_dadda_pg_rca32_and_3_10[0], h_s_dadda_pg_rca32_fa42_xor1, h_s_dadda_pg_rca32_fa42_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_11(a[2], b[11], h_s_dadda_pg_rca32_and_2_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_12(a[1], b[12], h_s_dadda_pg_rca32_and_1_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_13(a[0], b[13], h_s_dadda_pg_rca32_and_0_13);
  fa fa_h_s_dadda_pg_rca32_fa43_out(h_s_dadda_pg_rca32_and_2_11[0], h_s_dadda_pg_rca32_and_1_12[0], h_s_dadda_pg_rca32_and_0_13[0], h_s_dadda_pg_rca32_fa43_xor1, h_s_dadda_pg_rca32_fa43_or0);
  ha ha_h_s_dadda_pg_rca32_ha11_out(h_s_dadda_pg_rca32_fa37_xor1[0], h_s_dadda_pg_rca32_fa38_xor1[0], h_s_dadda_pg_rca32_ha11_xor0, h_s_dadda_pg_rca32_ha11_and0);
  fa fa_h_s_dadda_pg_rca32_fa44_out(h_s_dadda_pg_rca32_ha11_and0[0], h_s_dadda_pg_rca32_fa43_or0[0], h_s_dadda_pg_rca32_fa42_or0[0], h_s_dadda_pg_rca32_fa44_xor1, h_s_dadda_pg_rca32_fa44_or0);
  fa fa_h_s_dadda_pg_rca32_fa45_out(h_s_dadda_pg_rca32_fa41_or0[0], h_s_dadda_pg_rca32_fa40_or0[0], h_s_dadda_pg_rca32_fa39_or0[0], h_s_dadda_pg_rca32_fa45_xor1, h_s_dadda_pg_rca32_fa45_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_0(a[14], b[0], h_s_dadda_pg_rca32_and_14_0);
  fa fa_h_s_dadda_pg_rca32_fa46_out(h_s_dadda_pg_rca32_fa38_or0[0], h_s_dadda_pg_rca32_fa37_or0[0], h_s_dadda_pg_rca32_and_14_0[0], h_s_dadda_pg_rca32_fa46_xor1, h_s_dadda_pg_rca32_fa46_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_1(a[13], b[1], h_s_dadda_pg_rca32_and_13_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_2(a[12], b[2], h_s_dadda_pg_rca32_and_12_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_3(a[11], b[3], h_s_dadda_pg_rca32_and_11_3);
  fa fa_h_s_dadda_pg_rca32_fa47_out(h_s_dadda_pg_rca32_and_13_1[0], h_s_dadda_pg_rca32_and_12_2[0], h_s_dadda_pg_rca32_and_11_3[0], h_s_dadda_pg_rca32_fa47_xor1, h_s_dadda_pg_rca32_fa47_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_4(a[10], b[4], h_s_dadda_pg_rca32_and_10_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_5(a[9], b[5], h_s_dadda_pg_rca32_and_9_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_6(a[8], b[6], h_s_dadda_pg_rca32_and_8_6);
  fa fa_h_s_dadda_pg_rca32_fa48_out(h_s_dadda_pg_rca32_and_10_4[0], h_s_dadda_pg_rca32_and_9_5[0], h_s_dadda_pg_rca32_and_8_6[0], h_s_dadda_pg_rca32_fa48_xor1, h_s_dadda_pg_rca32_fa48_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_7(a[7], b[7], h_s_dadda_pg_rca32_and_7_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_8(a[6], b[8], h_s_dadda_pg_rca32_and_6_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_9(a[5], b[9], h_s_dadda_pg_rca32_and_5_9);
  fa fa_h_s_dadda_pg_rca32_fa49_out(h_s_dadda_pg_rca32_and_7_7[0], h_s_dadda_pg_rca32_and_6_8[0], h_s_dadda_pg_rca32_and_5_9[0], h_s_dadda_pg_rca32_fa49_xor1, h_s_dadda_pg_rca32_fa49_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_10(a[4], b[10], h_s_dadda_pg_rca32_and_4_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_11(a[3], b[11], h_s_dadda_pg_rca32_and_3_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_12(a[2], b[12], h_s_dadda_pg_rca32_and_2_12);
  fa fa_h_s_dadda_pg_rca32_fa50_out(h_s_dadda_pg_rca32_and_4_10[0], h_s_dadda_pg_rca32_and_3_11[0], h_s_dadda_pg_rca32_and_2_12[0], h_s_dadda_pg_rca32_fa50_xor1, h_s_dadda_pg_rca32_fa50_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_13(a[1], b[13], h_s_dadda_pg_rca32_and_1_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_14(a[0], b[14], h_s_dadda_pg_rca32_and_0_14);
  fa fa_h_s_dadda_pg_rca32_fa51_out(h_s_dadda_pg_rca32_and_1_13[0], h_s_dadda_pg_rca32_and_0_14[0], h_s_dadda_pg_rca32_fa44_xor1[0], h_s_dadda_pg_rca32_fa51_xor1, h_s_dadda_pg_rca32_fa51_or0);
  ha ha_h_s_dadda_pg_rca32_ha12_out(h_s_dadda_pg_rca32_fa45_xor1[0], h_s_dadda_pg_rca32_fa46_xor1[0], h_s_dadda_pg_rca32_ha12_xor0, h_s_dadda_pg_rca32_ha12_and0);
  fa fa_h_s_dadda_pg_rca32_fa52_out(h_s_dadda_pg_rca32_ha12_and0[0], h_s_dadda_pg_rca32_fa51_or0[0], h_s_dadda_pg_rca32_fa50_or0[0], h_s_dadda_pg_rca32_fa52_xor1, h_s_dadda_pg_rca32_fa52_or0);
  fa fa_h_s_dadda_pg_rca32_fa53_out(h_s_dadda_pg_rca32_fa49_or0[0], h_s_dadda_pg_rca32_fa48_or0[0], h_s_dadda_pg_rca32_fa47_or0[0], h_s_dadda_pg_rca32_fa53_xor1, h_s_dadda_pg_rca32_fa53_or0);
  fa fa_h_s_dadda_pg_rca32_fa54_out(h_s_dadda_pg_rca32_fa46_or0[0], h_s_dadda_pg_rca32_fa45_or0[0], h_s_dadda_pg_rca32_fa44_or0[0], h_s_dadda_pg_rca32_fa54_xor1, h_s_dadda_pg_rca32_fa54_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_0(a[15], b[0], h_s_dadda_pg_rca32_and_15_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_1(a[14], b[1], h_s_dadda_pg_rca32_and_14_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_2(a[13], b[2], h_s_dadda_pg_rca32_and_13_2);
  fa fa_h_s_dadda_pg_rca32_fa55_out(h_s_dadda_pg_rca32_and_15_0[0], h_s_dadda_pg_rca32_and_14_1[0], h_s_dadda_pg_rca32_and_13_2[0], h_s_dadda_pg_rca32_fa55_xor1, h_s_dadda_pg_rca32_fa55_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_3(a[12], b[3], h_s_dadda_pg_rca32_and_12_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_4(a[11], b[4], h_s_dadda_pg_rca32_and_11_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_5(a[10], b[5], h_s_dadda_pg_rca32_and_10_5);
  fa fa_h_s_dadda_pg_rca32_fa56_out(h_s_dadda_pg_rca32_and_12_3[0], h_s_dadda_pg_rca32_and_11_4[0], h_s_dadda_pg_rca32_and_10_5[0], h_s_dadda_pg_rca32_fa56_xor1, h_s_dadda_pg_rca32_fa56_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_6(a[9], b[6], h_s_dadda_pg_rca32_and_9_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_7(a[8], b[7], h_s_dadda_pg_rca32_and_8_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_8(a[7], b[8], h_s_dadda_pg_rca32_and_7_8);
  fa fa_h_s_dadda_pg_rca32_fa57_out(h_s_dadda_pg_rca32_and_9_6[0], h_s_dadda_pg_rca32_and_8_7[0], h_s_dadda_pg_rca32_and_7_8[0], h_s_dadda_pg_rca32_fa57_xor1, h_s_dadda_pg_rca32_fa57_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_9(a[6], b[9], h_s_dadda_pg_rca32_and_6_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_10(a[5], b[10], h_s_dadda_pg_rca32_and_5_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_11(a[4], b[11], h_s_dadda_pg_rca32_and_4_11);
  fa fa_h_s_dadda_pg_rca32_fa58_out(h_s_dadda_pg_rca32_and_6_9[0], h_s_dadda_pg_rca32_and_5_10[0], h_s_dadda_pg_rca32_and_4_11[0], h_s_dadda_pg_rca32_fa58_xor1, h_s_dadda_pg_rca32_fa58_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_12(a[3], b[12], h_s_dadda_pg_rca32_and_3_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_13(a[2], b[13], h_s_dadda_pg_rca32_and_2_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_14(a[1], b[14], h_s_dadda_pg_rca32_and_1_14);
  fa fa_h_s_dadda_pg_rca32_fa59_out(h_s_dadda_pg_rca32_and_3_12[0], h_s_dadda_pg_rca32_and_2_13[0], h_s_dadda_pg_rca32_and_1_14[0], h_s_dadda_pg_rca32_fa59_xor1, h_s_dadda_pg_rca32_fa59_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_15(a[0], b[15], h_s_dadda_pg_rca32_and_0_15);
  fa fa_h_s_dadda_pg_rca32_fa60_out(h_s_dadda_pg_rca32_and_0_15[0], h_s_dadda_pg_rca32_fa52_xor1[0], h_s_dadda_pg_rca32_fa53_xor1[0], h_s_dadda_pg_rca32_fa60_xor1, h_s_dadda_pg_rca32_fa60_or0);
  ha ha_h_s_dadda_pg_rca32_ha13_out(h_s_dadda_pg_rca32_fa54_xor1[0], h_s_dadda_pg_rca32_fa55_xor1[0], h_s_dadda_pg_rca32_ha13_xor0, h_s_dadda_pg_rca32_ha13_and0);
  fa fa_h_s_dadda_pg_rca32_fa61_out(h_s_dadda_pg_rca32_ha13_and0[0], h_s_dadda_pg_rca32_fa60_or0[0], h_s_dadda_pg_rca32_fa59_or0[0], h_s_dadda_pg_rca32_fa61_xor1, h_s_dadda_pg_rca32_fa61_or0);
  fa fa_h_s_dadda_pg_rca32_fa62_out(h_s_dadda_pg_rca32_fa58_or0[0], h_s_dadda_pg_rca32_fa57_or0[0], h_s_dadda_pg_rca32_fa56_or0[0], h_s_dadda_pg_rca32_fa62_xor1, h_s_dadda_pg_rca32_fa62_or0);
  fa fa_h_s_dadda_pg_rca32_fa63_out(h_s_dadda_pg_rca32_fa55_or0[0], h_s_dadda_pg_rca32_fa54_or0[0], h_s_dadda_pg_rca32_fa53_or0[0], h_s_dadda_pg_rca32_fa63_xor1, h_s_dadda_pg_rca32_fa63_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_0(a[16], b[0], h_s_dadda_pg_rca32_and_16_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_1(a[15], b[1], h_s_dadda_pg_rca32_and_15_1);
  fa fa_h_s_dadda_pg_rca32_fa64_out(h_s_dadda_pg_rca32_fa52_or0[0], h_s_dadda_pg_rca32_and_16_0[0], h_s_dadda_pg_rca32_and_15_1[0], h_s_dadda_pg_rca32_fa64_xor1, h_s_dadda_pg_rca32_fa64_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_2(a[14], b[2], h_s_dadda_pg_rca32_and_14_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_3(a[13], b[3], h_s_dadda_pg_rca32_and_13_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_4(a[12], b[4], h_s_dadda_pg_rca32_and_12_4);
  fa fa_h_s_dadda_pg_rca32_fa65_out(h_s_dadda_pg_rca32_and_14_2[0], h_s_dadda_pg_rca32_and_13_3[0], h_s_dadda_pg_rca32_and_12_4[0], h_s_dadda_pg_rca32_fa65_xor1, h_s_dadda_pg_rca32_fa65_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_5(a[11], b[5], h_s_dadda_pg_rca32_and_11_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_6(a[10], b[6], h_s_dadda_pg_rca32_and_10_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_7(a[9], b[7], h_s_dadda_pg_rca32_and_9_7);
  fa fa_h_s_dadda_pg_rca32_fa66_out(h_s_dadda_pg_rca32_and_11_5[0], h_s_dadda_pg_rca32_and_10_6[0], h_s_dadda_pg_rca32_and_9_7[0], h_s_dadda_pg_rca32_fa66_xor1, h_s_dadda_pg_rca32_fa66_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_8(a[8], b[8], h_s_dadda_pg_rca32_and_8_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_9(a[7], b[9], h_s_dadda_pg_rca32_and_7_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_10(a[6], b[10], h_s_dadda_pg_rca32_and_6_10);
  fa fa_h_s_dadda_pg_rca32_fa67_out(h_s_dadda_pg_rca32_and_8_8[0], h_s_dadda_pg_rca32_and_7_9[0], h_s_dadda_pg_rca32_and_6_10[0], h_s_dadda_pg_rca32_fa67_xor1, h_s_dadda_pg_rca32_fa67_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_11(a[5], b[11], h_s_dadda_pg_rca32_and_5_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_12(a[4], b[12], h_s_dadda_pg_rca32_and_4_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_13(a[3], b[13], h_s_dadda_pg_rca32_and_3_13);
  fa fa_h_s_dadda_pg_rca32_fa68_out(h_s_dadda_pg_rca32_and_5_11[0], h_s_dadda_pg_rca32_and_4_12[0], h_s_dadda_pg_rca32_and_3_13[0], h_s_dadda_pg_rca32_fa68_xor1, h_s_dadda_pg_rca32_fa68_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_14(a[2], b[14], h_s_dadda_pg_rca32_and_2_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_15(a[1], b[15], h_s_dadda_pg_rca32_and_1_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_16(a[0], b[16], h_s_dadda_pg_rca32_and_0_16);
  fa fa_h_s_dadda_pg_rca32_fa69_out(h_s_dadda_pg_rca32_and_2_14[0], h_s_dadda_pg_rca32_and_1_15[0], h_s_dadda_pg_rca32_and_0_16[0], h_s_dadda_pg_rca32_fa69_xor1, h_s_dadda_pg_rca32_fa69_or0);
  fa fa_h_s_dadda_pg_rca32_fa70_out(h_s_dadda_pg_rca32_fa61_xor1[0], h_s_dadda_pg_rca32_fa62_xor1[0], h_s_dadda_pg_rca32_fa63_xor1[0], h_s_dadda_pg_rca32_fa70_xor1, h_s_dadda_pg_rca32_fa70_or0);
  ha ha_h_s_dadda_pg_rca32_ha14_out(h_s_dadda_pg_rca32_fa64_xor1[0], h_s_dadda_pg_rca32_fa65_xor1[0], h_s_dadda_pg_rca32_ha14_xor0, h_s_dadda_pg_rca32_ha14_and0);
  fa fa_h_s_dadda_pg_rca32_fa71_out(h_s_dadda_pg_rca32_ha14_and0[0], h_s_dadda_pg_rca32_fa70_or0[0], h_s_dadda_pg_rca32_fa69_or0[0], h_s_dadda_pg_rca32_fa71_xor1, h_s_dadda_pg_rca32_fa71_or0);
  fa fa_h_s_dadda_pg_rca32_fa72_out(h_s_dadda_pg_rca32_fa68_or0[0], h_s_dadda_pg_rca32_fa67_or0[0], h_s_dadda_pg_rca32_fa66_or0[0], h_s_dadda_pg_rca32_fa72_xor1, h_s_dadda_pg_rca32_fa72_or0);
  fa fa_h_s_dadda_pg_rca32_fa73_out(h_s_dadda_pg_rca32_fa65_or0[0], h_s_dadda_pg_rca32_fa64_or0[0], h_s_dadda_pg_rca32_fa63_or0[0], h_s_dadda_pg_rca32_fa73_xor1, h_s_dadda_pg_rca32_fa73_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_0(a[17], b[0], h_s_dadda_pg_rca32_and_17_0);
  fa fa_h_s_dadda_pg_rca32_fa74_out(h_s_dadda_pg_rca32_fa62_or0[0], h_s_dadda_pg_rca32_fa61_or0[0], h_s_dadda_pg_rca32_and_17_0[0], h_s_dadda_pg_rca32_fa74_xor1, h_s_dadda_pg_rca32_fa74_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_1(a[16], b[1], h_s_dadda_pg_rca32_and_16_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_2(a[15], b[2], h_s_dadda_pg_rca32_and_15_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_3(a[14], b[3], h_s_dadda_pg_rca32_and_14_3);
  fa fa_h_s_dadda_pg_rca32_fa75_out(h_s_dadda_pg_rca32_and_16_1[0], h_s_dadda_pg_rca32_and_15_2[0], h_s_dadda_pg_rca32_and_14_3[0], h_s_dadda_pg_rca32_fa75_xor1, h_s_dadda_pg_rca32_fa75_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_4(a[13], b[4], h_s_dadda_pg_rca32_and_13_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_5(a[12], b[5], h_s_dadda_pg_rca32_and_12_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_6(a[11], b[6], h_s_dadda_pg_rca32_and_11_6);
  fa fa_h_s_dadda_pg_rca32_fa76_out(h_s_dadda_pg_rca32_and_13_4[0], h_s_dadda_pg_rca32_and_12_5[0], h_s_dadda_pg_rca32_and_11_6[0], h_s_dadda_pg_rca32_fa76_xor1, h_s_dadda_pg_rca32_fa76_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_7(a[10], b[7], h_s_dadda_pg_rca32_and_10_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_8(a[9], b[8], h_s_dadda_pg_rca32_and_9_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_9(a[8], b[9], h_s_dadda_pg_rca32_and_8_9);
  fa fa_h_s_dadda_pg_rca32_fa77_out(h_s_dadda_pg_rca32_and_10_7[0], h_s_dadda_pg_rca32_and_9_8[0], h_s_dadda_pg_rca32_and_8_9[0], h_s_dadda_pg_rca32_fa77_xor1, h_s_dadda_pg_rca32_fa77_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_10(a[7], b[10], h_s_dadda_pg_rca32_and_7_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_11(a[6], b[11], h_s_dadda_pg_rca32_and_6_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_12(a[5], b[12], h_s_dadda_pg_rca32_and_5_12);
  fa fa_h_s_dadda_pg_rca32_fa78_out(h_s_dadda_pg_rca32_and_7_10[0], h_s_dadda_pg_rca32_and_6_11[0], h_s_dadda_pg_rca32_and_5_12[0], h_s_dadda_pg_rca32_fa78_xor1, h_s_dadda_pg_rca32_fa78_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_13(a[4], b[13], h_s_dadda_pg_rca32_and_4_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_14(a[3], b[14], h_s_dadda_pg_rca32_and_3_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_15(a[2], b[15], h_s_dadda_pg_rca32_and_2_15);
  fa fa_h_s_dadda_pg_rca32_fa79_out(h_s_dadda_pg_rca32_and_4_13[0], h_s_dadda_pg_rca32_and_3_14[0], h_s_dadda_pg_rca32_and_2_15[0], h_s_dadda_pg_rca32_fa79_xor1, h_s_dadda_pg_rca32_fa79_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_16(a[1], b[16], h_s_dadda_pg_rca32_and_1_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_17(a[0], b[17], h_s_dadda_pg_rca32_and_0_17);
  fa fa_h_s_dadda_pg_rca32_fa80_out(h_s_dadda_pg_rca32_and_1_16[0], h_s_dadda_pg_rca32_and_0_17[0], h_s_dadda_pg_rca32_fa71_xor1[0], h_s_dadda_pg_rca32_fa80_xor1, h_s_dadda_pg_rca32_fa80_or0);
  fa fa_h_s_dadda_pg_rca32_fa81_out(h_s_dadda_pg_rca32_fa72_xor1[0], h_s_dadda_pg_rca32_fa73_xor1[0], h_s_dadda_pg_rca32_fa74_xor1[0], h_s_dadda_pg_rca32_fa81_xor1, h_s_dadda_pg_rca32_fa81_or0);
  ha ha_h_s_dadda_pg_rca32_ha15_out(h_s_dadda_pg_rca32_fa75_xor1[0], h_s_dadda_pg_rca32_fa76_xor1[0], h_s_dadda_pg_rca32_ha15_xor0, h_s_dadda_pg_rca32_ha15_and0);
  fa fa_h_s_dadda_pg_rca32_fa82_out(h_s_dadda_pg_rca32_ha15_and0[0], h_s_dadda_pg_rca32_fa81_or0[0], h_s_dadda_pg_rca32_fa80_or0[0], h_s_dadda_pg_rca32_fa82_xor1, h_s_dadda_pg_rca32_fa82_or0);
  fa fa_h_s_dadda_pg_rca32_fa83_out(h_s_dadda_pg_rca32_fa79_or0[0], h_s_dadda_pg_rca32_fa78_or0[0], h_s_dadda_pg_rca32_fa77_or0[0], h_s_dadda_pg_rca32_fa83_xor1, h_s_dadda_pg_rca32_fa83_or0);
  fa fa_h_s_dadda_pg_rca32_fa84_out(h_s_dadda_pg_rca32_fa76_or0[0], h_s_dadda_pg_rca32_fa75_or0[0], h_s_dadda_pg_rca32_fa74_or0[0], h_s_dadda_pg_rca32_fa84_xor1, h_s_dadda_pg_rca32_fa84_or0);
  fa fa_h_s_dadda_pg_rca32_fa85_out(h_s_dadda_pg_rca32_fa73_or0[0], h_s_dadda_pg_rca32_fa72_or0[0], h_s_dadda_pg_rca32_fa71_or0[0], h_s_dadda_pg_rca32_fa85_xor1, h_s_dadda_pg_rca32_fa85_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_0(a[18], b[0], h_s_dadda_pg_rca32_and_18_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_1(a[17], b[1], h_s_dadda_pg_rca32_and_17_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_2(a[16], b[2], h_s_dadda_pg_rca32_and_16_2);
  fa fa_h_s_dadda_pg_rca32_fa86_out(h_s_dadda_pg_rca32_and_18_0[0], h_s_dadda_pg_rca32_and_17_1[0], h_s_dadda_pg_rca32_and_16_2[0], h_s_dadda_pg_rca32_fa86_xor1, h_s_dadda_pg_rca32_fa86_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_3(a[15], b[3], h_s_dadda_pg_rca32_and_15_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_4(a[14], b[4], h_s_dadda_pg_rca32_and_14_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_5(a[13], b[5], h_s_dadda_pg_rca32_and_13_5);
  fa fa_h_s_dadda_pg_rca32_fa87_out(h_s_dadda_pg_rca32_and_15_3[0], h_s_dadda_pg_rca32_and_14_4[0], h_s_dadda_pg_rca32_and_13_5[0], h_s_dadda_pg_rca32_fa87_xor1, h_s_dadda_pg_rca32_fa87_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_6(a[12], b[6], h_s_dadda_pg_rca32_and_12_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_7(a[11], b[7], h_s_dadda_pg_rca32_and_11_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_8(a[10], b[8], h_s_dadda_pg_rca32_and_10_8);
  fa fa_h_s_dadda_pg_rca32_fa88_out(h_s_dadda_pg_rca32_and_12_6[0], h_s_dadda_pg_rca32_and_11_7[0], h_s_dadda_pg_rca32_and_10_8[0], h_s_dadda_pg_rca32_fa88_xor1, h_s_dadda_pg_rca32_fa88_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_9(a[9], b[9], h_s_dadda_pg_rca32_and_9_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_10(a[8], b[10], h_s_dadda_pg_rca32_and_8_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_11(a[7], b[11], h_s_dadda_pg_rca32_and_7_11);
  fa fa_h_s_dadda_pg_rca32_fa89_out(h_s_dadda_pg_rca32_and_9_9[0], h_s_dadda_pg_rca32_and_8_10[0], h_s_dadda_pg_rca32_and_7_11[0], h_s_dadda_pg_rca32_fa89_xor1, h_s_dadda_pg_rca32_fa89_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_12(a[6], b[12], h_s_dadda_pg_rca32_and_6_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_13(a[5], b[13], h_s_dadda_pg_rca32_and_5_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_14(a[4], b[14], h_s_dadda_pg_rca32_and_4_14);
  fa fa_h_s_dadda_pg_rca32_fa90_out(h_s_dadda_pg_rca32_and_6_12[0], h_s_dadda_pg_rca32_and_5_13[0], h_s_dadda_pg_rca32_and_4_14[0], h_s_dadda_pg_rca32_fa90_xor1, h_s_dadda_pg_rca32_fa90_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_15(a[3], b[15], h_s_dadda_pg_rca32_and_3_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_16(a[2], b[16], h_s_dadda_pg_rca32_and_2_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_17(a[1], b[17], h_s_dadda_pg_rca32_and_1_17);
  fa fa_h_s_dadda_pg_rca32_fa91_out(h_s_dadda_pg_rca32_and_3_15[0], h_s_dadda_pg_rca32_and_2_16[0], h_s_dadda_pg_rca32_and_1_17[0], h_s_dadda_pg_rca32_fa91_xor1, h_s_dadda_pg_rca32_fa91_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_18(a[0], b[18], h_s_dadda_pg_rca32_and_0_18);
  fa fa_h_s_dadda_pg_rca32_fa92_out(h_s_dadda_pg_rca32_and_0_18[0], h_s_dadda_pg_rca32_fa82_xor1[0], h_s_dadda_pg_rca32_fa83_xor1[0], h_s_dadda_pg_rca32_fa92_xor1, h_s_dadda_pg_rca32_fa92_or0);
  fa fa_h_s_dadda_pg_rca32_fa93_out(h_s_dadda_pg_rca32_fa84_xor1[0], h_s_dadda_pg_rca32_fa85_xor1[0], h_s_dadda_pg_rca32_fa86_xor1[0], h_s_dadda_pg_rca32_fa93_xor1, h_s_dadda_pg_rca32_fa93_or0);
  ha ha_h_s_dadda_pg_rca32_ha16_out(h_s_dadda_pg_rca32_fa87_xor1[0], h_s_dadda_pg_rca32_fa88_xor1[0], h_s_dadda_pg_rca32_ha16_xor0, h_s_dadda_pg_rca32_ha16_and0);
  fa fa_h_s_dadda_pg_rca32_fa94_out(h_s_dadda_pg_rca32_ha16_and0[0], h_s_dadda_pg_rca32_fa93_or0[0], h_s_dadda_pg_rca32_fa92_or0[0], h_s_dadda_pg_rca32_fa94_xor1, h_s_dadda_pg_rca32_fa94_or0);
  fa fa_h_s_dadda_pg_rca32_fa95_out(h_s_dadda_pg_rca32_fa91_or0[0], h_s_dadda_pg_rca32_fa90_or0[0], h_s_dadda_pg_rca32_fa89_or0[0], h_s_dadda_pg_rca32_fa95_xor1, h_s_dadda_pg_rca32_fa95_or0);
  fa fa_h_s_dadda_pg_rca32_fa96_out(h_s_dadda_pg_rca32_fa88_or0[0], h_s_dadda_pg_rca32_fa87_or0[0], h_s_dadda_pg_rca32_fa86_or0[0], h_s_dadda_pg_rca32_fa96_xor1, h_s_dadda_pg_rca32_fa96_or0);
  fa fa_h_s_dadda_pg_rca32_fa97_out(h_s_dadda_pg_rca32_fa85_or0[0], h_s_dadda_pg_rca32_fa84_or0[0], h_s_dadda_pg_rca32_fa83_or0[0], h_s_dadda_pg_rca32_fa97_xor1, h_s_dadda_pg_rca32_fa97_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_0(a[19], b[0], h_s_dadda_pg_rca32_and_19_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_1(a[18], b[1], h_s_dadda_pg_rca32_and_18_1);
  fa fa_h_s_dadda_pg_rca32_fa98_out(h_s_dadda_pg_rca32_fa82_or0[0], h_s_dadda_pg_rca32_and_19_0[0], h_s_dadda_pg_rca32_and_18_1[0], h_s_dadda_pg_rca32_fa98_xor1, h_s_dadda_pg_rca32_fa98_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_2(a[17], b[2], h_s_dadda_pg_rca32_and_17_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_3(a[16], b[3], h_s_dadda_pg_rca32_and_16_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_4(a[15], b[4], h_s_dadda_pg_rca32_and_15_4);
  fa fa_h_s_dadda_pg_rca32_fa99_out(h_s_dadda_pg_rca32_and_17_2[0], h_s_dadda_pg_rca32_and_16_3[0], h_s_dadda_pg_rca32_and_15_4[0], h_s_dadda_pg_rca32_fa99_xor1, h_s_dadda_pg_rca32_fa99_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_5(a[14], b[5], h_s_dadda_pg_rca32_and_14_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_6(a[13], b[6], h_s_dadda_pg_rca32_and_13_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_7(a[12], b[7], h_s_dadda_pg_rca32_and_12_7);
  fa fa_h_s_dadda_pg_rca32_fa100_out(h_s_dadda_pg_rca32_and_14_5[0], h_s_dadda_pg_rca32_and_13_6[0], h_s_dadda_pg_rca32_and_12_7[0], h_s_dadda_pg_rca32_fa100_xor1, h_s_dadda_pg_rca32_fa100_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_8(a[11], b[8], h_s_dadda_pg_rca32_and_11_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_9(a[10], b[9], h_s_dadda_pg_rca32_and_10_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_10(a[9], b[10], h_s_dadda_pg_rca32_and_9_10);
  fa fa_h_s_dadda_pg_rca32_fa101_out(h_s_dadda_pg_rca32_and_11_8[0], h_s_dadda_pg_rca32_and_10_9[0], h_s_dadda_pg_rca32_and_9_10[0], h_s_dadda_pg_rca32_fa101_xor1, h_s_dadda_pg_rca32_fa101_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_11(a[8], b[11], h_s_dadda_pg_rca32_and_8_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_12(a[7], b[12], h_s_dadda_pg_rca32_and_7_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_13(a[6], b[13], h_s_dadda_pg_rca32_and_6_13);
  fa fa_h_s_dadda_pg_rca32_fa102_out(h_s_dadda_pg_rca32_and_8_11[0], h_s_dadda_pg_rca32_and_7_12[0], h_s_dadda_pg_rca32_and_6_13[0], h_s_dadda_pg_rca32_fa102_xor1, h_s_dadda_pg_rca32_fa102_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_14(a[5], b[14], h_s_dadda_pg_rca32_and_5_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_15(a[4], b[15], h_s_dadda_pg_rca32_and_4_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_16(a[3], b[16], h_s_dadda_pg_rca32_and_3_16);
  fa fa_h_s_dadda_pg_rca32_fa103_out(h_s_dadda_pg_rca32_and_5_14[0], h_s_dadda_pg_rca32_and_4_15[0], h_s_dadda_pg_rca32_and_3_16[0], h_s_dadda_pg_rca32_fa103_xor1, h_s_dadda_pg_rca32_fa103_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_17(a[2], b[17], h_s_dadda_pg_rca32_and_2_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_18(a[1], b[18], h_s_dadda_pg_rca32_and_1_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_19(a[0], b[19], h_s_dadda_pg_rca32_and_0_19);
  fa fa_h_s_dadda_pg_rca32_fa104_out(h_s_dadda_pg_rca32_and_2_17[0], h_s_dadda_pg_rca32_and_1_18[0], h_s_dadda_pg_rca32_and_0_19[0], h_s_dadda_pg_rca32_fa104_xor1, h_s_dadda_pg_rca32_fa104_or0);
  fa fa_h_s_dadda_pg_rca32_fa105_out(h_s_dadda_pg_rca32_fa94_xor1[0], h_s_dadda_pg_rca32_fa95_xor1[0], h_s_dadda_pg_rca32_fa96_xor1[0], h_s_dadda_pg_rca32_fa105_xor1, h_s_dadda_pg_rca32_fa105_or0);
  fa fa_h_s_dadda_pg_rca32_fa106_out(h_s_dadda_pg_rca32_fa97_xor1[0], h_s_dadda_pg_rca32_fa98_xor1[0], h_s_dadda_pg_rca32_fa99_xor1[0], h_s_dadda_pg_rca32_fa106_xor1, h_s_dadda_pg_rca32_fa106_or0);
  ha ha_h_s_dadda_pg_rca32_ha17_out(h_s_dadda_pg_rca32_fa100_xor1[0], h_s_dadda_pg_rca32_fa101_xor1[0], h_s_dadda_pg_rca32_ha17_xor0, h_s_dadda_pg_rca32_ha17_and0);
  fa fa_h_s_dadda_pg_rca32_fa107_out(h_s_dadda_pg_rca32_ha17_and0[0], h_s_dadda_pg_rca32_fa106_or0[0], h_s_dadda_pg_rca32_fa105_or0[0], h_s_dadda_pg_rca32_fa107_xor1, h_s_dadda_pg_rca32_fa107_or0);
  fa fa_h_s_dadda_pg_rca32_fa108_out(h_s_dadda_pg_rca32_fa104_or0[0], h_s_dadda_pg_rca32_fa103_or0[0], h_s_dadda_pg_rca32_fa102_or0[0], h_s_dadda_pg_rca32_fa108_xor1, h_s_dadda_pg_rca32_fa108_or0);
  fa fa_h_s_dadda_pg_rca32_fa109_out(h_s_dadda_pg_rca32_fa101_or0[0], h_s_dadda_pg_rca32_fa100_or0[0], h_s_dadda_pg_rca32_fa99_or0[0], h_s_dadda_pg_rca32_fa109_xor1, h_s_dadda_pg_rca32_fa109_or0);
  fa fa_h_s_dadda_pg_rca32_fa110_out(h_s_dadda_pg_rca32_fa98_or0[0], h_s_dadda_pg_rca32_fa97_or0[0], h_s_dadda_pg_rca32_fa96_or0[0], h_s_dadda_pg_rca32_fa110_xor1, h_s_dadda_pg_rca32_fa110_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_0(a[20], b[0], h_s_dadda_pg_rca32_and_20_0);
  fa fa_h_s_dadda_pg_rca32_fa111_out(h_s_dadda_pg_rca32_fa95_or0[0], h_s_dadda_pg_rca32_fa94_or0[0], h_s_dadda_pg_rca32_and_20_0[0], h_s_dadda_pg_rca32_fa111_xor1, h_s_dadda_pg_rca32_fa111_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_1(a[19], b[1], h_s_dadda_pg_rca32_and_19_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_2(a[18], b[2], h_s_dadda_pg_rca32_and_18_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_3(a[17], b[3], h_s_dadda_pg_rca32_and_17_3);
  fa fa_h_s_dadda_pg_rca32_fa112_out(h_s_dadda_pg_rca32_and_19_1[0], h_s_dadda_pg_rca32_and_18_2[0], h_s_dadda_pg_rca32_and_17_3[0], h_s_dadda_pg_rca32_fa112_xor1, h_s_dadda_pg_rca32_fa112_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_4(a[16], b[4], h_s_dadda_pg_rca32_and_16_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_5(a[15], b[5], h_s_dadda_pg_rca32_and_15_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_6(a[14], b[6], h_s_dadda_pg_rca32_and_14_6);
  fa fa_h_s_dadda_pg_rca32_fa113_out(h_s_dadda_pg_rca32_and_16_4[0], h_s_dadda_pg_rca32_and_15_5[0], h_s_dadda_pg_rca32_and_14_6[0], h_s_dadda_pg_rca32_fa113_xor1, h_s_dadda_pg_rca32_fa113_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_7(a[13], b[7], h_s_dadda_pg_rca32_and_13_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_8(a[12], b[8], h_s_dadda_pg_rca32_and_12_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_9(a[11], b[9], h_s_dadda_pg_rca32_and_11_9);
  fa fa_h_s_dadda_pg_rca32_fa114_out(h_s_dadda_pg_rca32_and_13_7[0], h_s_dadda_pg_rca32_and_12_8[0], h_s_dadda_pg_rca32_and_11_9[0], h_s_dadda_pg_rca32_fa114_xor1, h_s_dadda_pg_rca32_fa114_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_10(a[10], b[10], h_s_dadda_pg_rca32_and_10_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_11(a[9], b[11], h_s_dadda_pg_rca32_and_9_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_12(a[8], b[12], h_s_dadda_pg_rca32_and_8_12);
  fa fa_h_s_dadda_pg_rca32_fa115_out(h_s_dadda_pg_rca32_and_10_10[0], h_s_dadda_pg_rca32_and_9_11[0], h_s_dadda_pg_rca32_and_8_12[0], h_s_dadda_pg_rca32_fa115_xor1, h_s_dadda_pg_rca32_fa115_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_13(a[7], b[13], h_s_dadda_pg_rca32_and_7_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_14(a[6], b[14], h_s_dadda_pg_rca32_and_6_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_15(a[5], b[15], h_s_dadda_pg_rca32_and_5_15);
  fa fa_h_s_dadda_pg_rca32_fa116_out(h_s_dadda_pg_rca32_and_7_13[0], h_s_dadda_pg_rca32_and_6_14[0], h_s_dadda_pg_rca32_and_5_15[0], h_s_dadda_pg_rca32_fa116_xor1, h_s_dadda_pg_rca32_fa116_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_16(a[4], b[16], h_s_dadda_pg_rca32_and_4_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_17(a[3], b[17], h_s_dadda_pg_rca32_and_3_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_18(a[2], b[18], h_s_dadda_pg_rca32_and_2_18);
  fa fa_h_s_dadda_pg_rca32_fa117_out(h_s_dadda_pg_rca32_and_4_16[0], h_s_dadda_pg_rca32_and_3_17[0], h_s_dadda_pg_rca32_and_2_18[0], h_s_dadda_pg_rca32_fa117_xor1, h_s_dadda_pg_rca32_fa117_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_19(a[1], b[19], h_s_dadda_pg_rca32_and_1_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_20(a[0], b[20], h_s_dadda_pg_rca32_and_0_20);
  fa fa_h_s_dadda_pg_rca32_fa118_out(h_s_dadda_pg_rca32_and_1_19[0], h_s_dadda_pg_rca32_and_0_20[0], h_s_dadda_pg_rca32_fa107_xor1[0], h_s_dadda_pg_rca32_fa118_xor1, h_s_dadda_pg_rca32_fa118_or0);
  fa fa_h_s_dadda_pg_rca32_fa119_out(h_s_dadda_pg_rca32_fa108_xor1[0], h_s_dadda_pg_rca32_fa109_xor1[0], h_s_dadda_pg_rca32_fa110_xor1[0], h_s_dadda_pg_rca32_fa119_xor1, h_s_dadda_pg_rca32_fa119_or0);
  fa fa_h_s_dadda_pg_rca32_fa120_out(h_s_dadda_pg_rca32_fa111_xor1[0], h_s_dadda_pg_rca32_fa112_xor1[0], h_s_dadda_pg_rca32_fa113_xor1[0], h_s_dadda_pg_rca32_fa120_xor1, h_s_dadda_pg_rca32_fa120_or0);
  ha ha_h_s_dadda_pg_rca32_ha18_out(h_s_dadda_pg_rca32_fa114_xor1[0], h_s_dadda_pg_rca32_fa115_xor1[0], h_s_dadda_pg_rca32_ha18_xor0, h_s_dadda_pg_rca32_ha18_and0);
  fa fa_h_s_dadda_pg_rca32_fa121_out(h_s_dadda_pg_rca32_ha18_and0[0], h_s_dadda_pg_rca32_fa120_or0[0], h_s_dadda_pg_rca32_fa119_or0[0], h_s_dadda_pg_rca32_fa121_xor1, h_s_dadda_pg_rca32_fa121_or0);
  fa fa_h_s_dadda_pg_rca32_fa122_out(h_s_dadda_pg_rca32_fa118_or0[0], h_s_dadda_pg_rca32_fa117_or0[0], h_s_dadda_pg_rca32_fa116_or0[0], h_s_dadda_pg_rca32_fa122_xor1, h_s_dadda_pg_rca32_fa122_or0);
  fa fa_h_s_dadda_pg_rca32_fa123_out(h_s_dadda_pg_rca32_fa115_or0[0], h_s_dadda_pg_rca32_fa114_or0[0], h_s_dadda_pg_rca32_fa113_or0[0], h_s_dadda_pg_rca32_fa123_xor1, h_s_dadda_pg_rca32_fa123_or0);
  fa fa_h_s_dadda_pg_rca32_fa124_out(h_s_dadda_pg_rca32_fa112_or0[0], h_s_dadda_pg_rca32_fa111_or0[0], h_s_dadda_pg_rca32_fa110_or0[0], h_s_dadda_pg_rca32_fa124_xor1, h_s_dadda_pg_rca32_fa124_or0);
  fa fa_h_s_dadda_pg_rca32_fa125_out(h_s_dadda_pg_rca32_fa109_or0[0], h_s_dadda_pg_rca32_fa108_or0[0], h_s_dadda_pg_rca32_fa107_or0[0], h_s_dadda_pg_rca32_fa125_xor1, h_s_dadda_pg_rca32_fa125_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_0(a[21], b[0], h_s_dadda_pg_rca32_and_21_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_1(a[20], b[1], h_s_dadda_pg_rca32_and_20_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_2(a[19], b[2], h_s_dadda_pg_rca32_and_19_2);
  fa fa_h_s_dadda_pg_rca32_fa126_out(h_s_dadda_pg_rca32_and_21_0[0], h_s_dadda_pg_rca32_and_20_1[0], h_s_dadda_pg_rca32_and_19_2[0], h_s_dadda_pg_rca32_fa126_xor1, h_s_dadda_pg_rca32_fa126_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_3(a[18], b[3], h_s_dadda_pg_rca32_and_18_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_4(a[17], b[4], h_s_dadda_pg_rca32_and_17_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_5(a[16], b[5], h_s_dadda_pg_rca32_and_16_5);
  fa fa_h_s_dadda_pg_rca32_fa127_out(h_s_dadda_pg_rca32_and_18_3[0], h_s_dadda_pg_rca32_and_17_4[0], h_s_dadda_pg_rca32_and_16_5[0], h_s_dadda_pg_rca32_fa127_xor1, h_s_dadda_pg_rca32_fa127_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_6(a[15], b[6], h_s_dadda_pg_rca32_and_15_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_7(a[14], b[7], h_s_dadda_pg_rca32_and_14_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_8(a[13], b[8], h_s_dadda_pg_rca32_and_13_8);
  fa fa_h_s_dadda_pg_rca32_fa128_out(h_s_dadda_pg_rca32_and_15_6[0], h_s_dadda_pg_rca32_and_14_7[0], h_s_dadda_pg_rca32_and_13_8[0], h_s_dadda_pg_rca32_fa128_xor1, h_s_dadda_pg_rca32_fa128_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_9(a[12], b[9], h_s_dadda_pg_rca32_and_12_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_10(a[11], b[10], h_s_dadda_pg_rca32_and_11_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_11(a[10], b[11], h_s_dadda_pg_rca32_and_10_11);
  fa fa_h_s_dadda_pg_rca32_fa129_out(h_s_dadda_pg_rca32_and_12_9[0], h_s_dadda_pg_rca32_and_11_10[0], h_s_dadda_pg_rca32_and_10_11[0], h_s_dadda_pg_rca32_fa129_xor1, h_s_dadda_pg_rca32_fa129_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_12(a[9], b[12], h_s_dadda_pg_rca32_and_9_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_13(a[8], b[13], h_s_dadda_pg_rca32_and_8_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_14(a[7], b[14], h_s_dadda_pg_rca32_and_7_14);
  fa fa_h_s_dadda_pg_rca32_fa130_out(h_s_dadda_pg_rca32_and_9_12[0], h_s_dadda_pg_rca32_and_8_13[0], h_s_dadda_pg_rca32_and_7_14[0], h_s_dadda_pg_rca32_fa130_xor1, h_s_dadda_pg_rca32_fa130_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_15(a[6], b[15], h_s_dadda_pg_rca32_and_6_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_16(a[5], b[16], h_s_dadda_pg_rca32_and_5_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_17(a[4], b[17], h_s_dadda_pg_rca32_and_4_17);
  fa fa_h_s_dadda_pg_rca32_fa131_out(h_s_dadda_pg_rca32_and_6_15[0], h_s_dadda_pg_rca32_and_5_16[0], h_s_dadda_pg_rca32_and_4_17[0], h_s_dadda_pg_rca32_fa131_xor1, h_s_dadda_pg_rca32_fa131_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_18(a[3], b[18], h_s_dadda_pg_rca32_and_3_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_19(a[2], b[19], h_s_dadda_pg_rca32_and_2_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_20(a[1], b[20], h_s_dadda_pg_rca32_and_1_20);
  fa fa_h_s_dadda_pg_rca32_fa132_out(h_s_dadda_pg_rca32_and_3_18[0], h_s_dadda_pg_rca32_and_2_19[0], h_s_dadda_pg_rca32_and_1_20[0], h_s_dadda_pg_rca32_fa132_xor1, h_s_dadda_pg_rca32_fa132_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_21(a[0], b[21], h_s_dadda_pg_rca32_and_0_21);
  fa fa_h_s_dadda_pg_rca32_fa133_out(h_s_dadda_pg_rca32_and_0_21[0], h_s_dadda_pg_rca32_fa121_xor1[0], h_s_dadda_pg_rca32_fa122_xor1[0], h_s_dadda_pg_rca32_fa133_xor1, h_s_dadda_pg_rca32_fa133_or0);
  fa fa_h_s_dadda_pg_rca32_fa134_out(h_s_dadda_pg_rca32_fa123_xor1[0], h_s_dadda_pg_rca32_fa124_xor1[0], h_s_dadda_pg_rca32_fa125_xor1[0], h_s_dadda_pg_rca32_fa134_xor1, h_s_dadda_pg_rca32_fa134_or0);
  fa fa_h_s_dadda_pg_rca32_fa135_out(h_s_dadda_pg_rca32_fa126_xor1[0], h_s_dadda_pg_rca32_fa127_xor1[0], h_s_dadda_pg_rca32_fa128_xor1[0], h_s_dadda_pg_rca32_fa135_xor1, h_s_dadda_pg_rca32_fa135_or0);
  ha ha_h_s_dadda_pg_rca32_ha19_out(h_s_dadda_pg_rca32_fa129_xor1[0], h_s_dadda_pg_rca32_fa130_xor1[0], h_s_dadda_pg_rca32_ha19_xor0, h_s_dadda_pg_rca32_ha19_and0);
  fa fa_h_s_dadda_pg_rca32_fa136_out(h_s_dadda_pg_rca32_ha19_and0[0], h_s_dadda_pg_rca32_fa135_or0[0], h_s_dadda_pg_rca32_fa134_or0[0], h_s_dadda_pg_rca32_fa136_xor1, h_s_dadda_pg_rca32_fa136_or0);
  fa fa_h_s_dadda_pg_rca32_fa137_out(h_s_dadda_pg_rca32_fa133_or0[0], h_s_dadda_pg_rca32_fa132_or0[0], h_s_dadda_pg_rca32_fa131_or0[0], h_s_dadda_pg_rca32_fa137_xor1, h_s_dadda_pg_rca32_fa137_or0);
  fa fa_h_s_dadda_pg_rca32_fa138_out(h_s_dadda_pg_rca32_fa130_or0[0], h_s_dadda_pg_rca32_fa129_or0[0], h_s_dadda_pg_rca32_fa128_or0[0], h_s_dadda_pg_rca32_fa138_xor1, h_s_dadda_pg_rca32_fa138_or0);
  fa fa_h_s_dadda_pg_rca32_fa139_out(h_s_dadda_pg_rca32_fa127_or0[0], h_s_dadda_pg_rca32_fa126_or0[0], h_s_dadda_pg_rca32_fa125_or0[0], h_s_dadda_pg_rca32_fa139_xor1, h_s_dadda_pg_rca32_fa139_or0);
  fa fa_h_s_dadda_pg_rca32_fa140_out(h_s_dadda_pg_rca32_fa124_or0[0], h_s_dadda_pg_rca32_fa123_or0[0], h_s_dadda_pg_rca32_fa122_or0[0], h_s_dadda_pg_rca32_fa140_xor1, h_s_dadda_pg_rca32_fa140_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_0(a[22], b[0], h_s_dadda_pg_rca32_and_22_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_1(a[21], b[1], h_s_dadda_pg_rca32_and_21_1);
  fa fa_h_s_dadda_pg_rca32_fa141_out(h_s_dadda_pg_rca32_fa121_or0[0], h_s_dadda_pg_rca32_and_22_0[0], h_s_dadda_pg_rca32_and_21_1[0], h_s_dadda_pg_rca32_fa141_xor1, h_s_dadda_pg_rca32_fa141_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_2(a[20], b[2], h_s_dadda_pg_rca32_and_20_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_3(a[19], b[3], h_s_dadda_pg_rca32_and_19_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_4(a[18], b[4], h_s_dadda_pg_rca32_and_18_4);
  fa fa_h_s_dadda_pg_rca32_fa142_out(h_s_dadda_pg_rca32_and_20_2[0], h_s_dadda_pg_rca32_and_19_3[0], h_s_dadda_pg_rca32_and_18_4[0], h_s_dadda_pg_rca32_fa142_xor1, h_s_dadda_pg_rca32_fa142_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_5(a[17], b[5], h_s_dadda_pg_rca32_and_17_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_6(a[16], b[6], h_s_dadda_pg_rca32_and_16_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_7(a[15], b[7], h_s_dadda_pg_rca32_and_15_7);
  fa fa_h_s_dadda_pg_rca32_fa143_out(h_s_dadda_pg_rca32_and_17_5[0], h_s_dadda_pg_rca32_and_16_6[0], h_s_dadda_pg_rca32_and_15_7[0], h_s_dadda_pg_rca32_fa143_xor1, h_s_dadda_pg_rca32_fa143_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_8(a[14], b[8], h_s_dadda_pg_rca32_and_14_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_9(a[13], b[9], h_s_dadda_pg_rca32_and_13_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_10(a[12], b[10], h_s_dadda_pg_rca32_and_12_10);
  fa fa_h_s_dadda_pg_rca32_fa144_out(h_s_dadda_pg_rca32_and_14_8[0], h_s_dadda_pg_rca32_and_13_9[0], h_s_dadda_pg_rca32_and_12_10[0], h_s_dadda_pg_rca32_fa144_xor1, h_s_dadda_pg_rca32_fa144_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_11(a[11], b[11], h_s_dadda_pg_rca32_and_11_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_12(a[10], b[12], h_s_dadda_pg_rca32_and_10_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_13(a[9], b[13], h_s_dadda_pg_rca32_and_9_13);
  fa fa_h_s_dadda_pg_rca32_fa145_out(h_s_dadda_pg_rca32_and_11_11[0], h_s_dadda_pg_rca32_and_10_12[0], h_s_dadda_pg_rca32_and_9_13[0], h_s_dadda_pg_rca32_fa145_xor1, h_s_dadda_pg_rca32_fa145_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_14(a[8], b[14], h_s_dadda_pg_rca32_and_8_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_15(a[7], b[15], h_s_dadda_pg_rca32_and_7_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_16(a[6], b[16], h_s_dadda_pg_rca32_and_6_16);
  fa fa_h_s_dadda_pg_rca32_fa146_out(h_s_dadda_pg_rca32_and_8_14[0], h_s_dadda_pg_rca32_and_7_15[0], h_s_dadda_pg_rca32_and_6_16[0], h_s_dadda_pg_rca32_fa146_xor1, h_s_dadda_pg_rca32_fa146_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_17(a[5], b[17], h_s_dadda_pg_rca32_and_5_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_18(a[4], b[18], h_s_dadda_pg_rca32_and_4_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_19(a[3], b[19], h_s_dadda_pg_rca32_and_3_19);
  fa fa_h_s_dadda_pg_rca32_fa147_out(h_s_dadda_pg_rca32_and_5_17[0], h_s_dadda_pg_rca32_and_4_18[0], h_s_dadda_pg_rca32_and_3_19[0], h_s_dadda_pg_rca32_fa147_xor1, h_s_dadda_pg_rca32_fa147_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_20(a[2], b[20], h_s_dadda_pg_rca32_and_2_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_21(a[1], b[21], h_s_dadda_pg_rca32_and_1_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_22(a[0], b[22], h_s_dadda_pg_rca32_and_0_22);
  fa fa_h_s_dadda_pg_rca32_fa148_out(h_s_dadda_pg_rca32_and_2_20[0], h_s_dadda_pg_rca32_and_1_21[0], h_s_dadda_pg_rca32_and_0_22[0], h_s_dadda_pg_rca32_fa148_xor1, h_s_dadda_pg_rca32_fa148_or0);
  fa fa_h_s_dadda_pg_rca32_fa149_out(h_s_dadda_pg_rca32_fa136_xor1[0], h_s_dadda_pg_rca32_fa137_xor1[0], h_s_dadda_pg_rca32_fa138_xor1[0], h_s_dadda_pg_rca32_fa149_xor1, h_s_dadda_pg_rca32_fa149_or0);
  fa fa_h_s_dadda_pg_rca32_fa150_out(h_s_dadda_pg_rca32_fa139_xor1[0], h_s_dadda_pg_rca32_fa140_xor1[0], h_s_dadda_pg_rca32_fa141_xor1[0], h_s_dadda_pg_rca32_fa150_xor1, h_s_dadda_pg_rca32_fa150_or0);
  fa fa_h_s_dadda_pg_rca32_fa151_out(h_s_dadda_pg_rca32_fa142_xor1[0], h_s_dadda_pg_rca32_fa143_xor1[0], h_s_dadda_pg_rca32_fa144_xor1[0], h_s_dadda_pg_rca32_fa151_xor1, h_s_dadda_pg_rca32_fa151_or0);
  ha ha_h_s_dadda_pg_rca32_ha20_out(h_s_dadda_pg_rca32_fa145_xor1[0], h_s_dadda_pg_rca32_fa146_xor1[0], h_s_dadda_pg_rca32_ha20_xor0, h_s_dadda_pg_rca32_ha20_and0);
  fa fa_h_s_dadda_pg_rca32_fa152_out(h_s_dadda_pg_rca32_ha20_and0[0], h_s_dadda_pg_rca32_fa151_or0[0], h_s_dadda_pg_rca32_fa150_or0[0], h_s_dadda_pg_rca32_fa152_xor1, h_s_dadda_pg_rca32_fa152_or0);
  fa fa_h_s_dadda_pg_rca32_fa153_out(h_s_dadda_pg_rca32_fa149_or0[0], h_s_dadda_pg_rca32_fa148_or0[0], h_s_dadda_pg_rca32_fa147_or0[0], h_s_dadda_pg_rca32_fa153_xor1, h_s_dadda_pg_rca32_fa153_or0);
  fa fa_h_s_dadda_pg_rca32_fa154_out(h_s_dadda_pg_rca32_fa146_or0[0], h_s_dadda_pg_rca32_fa145_or0[0], h_s_dadda_pg_rca32_fa144_or0[0], h_s_dadda_pg_rca32_fa154_xor1, h_s_dadda_pg_rca32_fa154_or0);
  fa fa_h_s_dadda_pg_rca32_fa155_out(h_s_dadda_pg_rca32_fa143_or0[0], h_s_dadda_pg_rca32_fa142_or0[0], h_s_dadda_pg_rca32_fa141_or0[0], h_s_dadda_pg_rca32_fa155_xor1, h_s_dadda_pg_rca32_fa155_or0);
  fa fa_h_s_dadda_pg_rca32_fa156_out(h_s_dadda_pg_rca32_fa140_or0[0], h_s_dadda_pg_rca32_fa139_or0[0], h_s_dadda_pg_rca32_fa138_or0[0], h_s_dadda_pg_rca32_fa156_xor1, h_s_dadda_pg_rca32_fa156_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_0(a[23], b[0], h_s_dadda_pg_rca32_and_23_0);
  fa fa_h_s_dadda_pg_rca32_fa157_out(h_s_dadda_pg_rca32_fa137_or0[0], h_s_dadda_pg_rca32_fa136_or0[0], h_s_dadda_pg_rca32_and_23_0[0], h_s_dadda_pg_rca32_fa157_xor1, h_s_dadda_pg_rca32_fa157_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_1(a[22], b[1], h_s_dadda_pg_rca32_and_22_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_2(a[21], b[2], h_s_dadda_pg_rca32_and_21_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_3(a[20], b[3], h_s_dadda_pg_rca32_and_20_3);
  fa fa_h_s_dadda_pg_rca32_fa158_out(h_s_dadda_pg_rca32_and_22_1[0], h_s_dadda_pg_rca32_and_21_2[0], h_s_dadda_pg_rca32_and_20_3[0], h_s_dadda_pg_rca32_fa158_xor1, h_s_dadda_pg_rca32_fa158_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_4(a[19], b[4], h_s_dadda_pg_rca32_and_19_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_5(a[18], b[5], h_s_dadda_pg_rca32_and_18_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_6(a[17], b[6], h_s_dadda_pg_rca32_and_17_6);
  fa fa_h_s_dadda_pg_rca32_fa159_out(h_s_dadda_pg_rca32_and_19_4[0], h_s_dadda_pg_rca32_and_18_5[0], h_s_dadda_pg_rca32_and_17_6[0], h_s_dadda_pg_rca32_fa159_xor1, h_s_dadda_pg_rca32_fa159_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_7(a[16], b[7], h_s_dadda_pg_rca32_and_16_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_8(a[15], b[8], h_s_dadda_pg_rca32_and_15_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_9(a[14], b[9], h_s_dadda_pg_rca32_and_14_9);
  fa fa_h_s_dadda_pg_rca32_fa160_out(h_s_dadda_pg_rca32_and_16_7[0], h_s_dadda_pg_rca32_and_15_8[0], h_s_dadda_pg_rca32_and_14_9[0], h_s_dadda_pg_rca32_fa160_xor1, h_s_dadda_pg_rca32_fa160_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_10(a[13], b[10], h_s_dadda_pg_rca32_and_13_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_11(a[12], b[11], h_s_dadda_pg_rca32_and_12_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_12(a[11], b[12], h_s_dadda_pg_rca32_and_11_12);
  fa fa_h_s_dadda_pg_rca32_fa161_out(h_s_dadda_pg_rca32_and_13_10[0], h_s_dadda_pg_rca32_and_12_11[0], h_s_dadda_pg_rca32_and_11_12[0], h_s_dadda_pg_rca32_fa161_xor1, h_s_dadda_pg_rca32_fa161_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_13(a[10], b[13], h_s_dadda_pg_rca32_and_10_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_14(a[9], b[14], h_s_dadda_pg_rca32_and_9_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_15(a[8], b[15], h_s_dadda_pg_rca32_and_8_15);
  fa fa_h_s_dadda_pg_rca32_fa162_out(h_s_dadda_pg_rca32_and_10_13[0], h_s_dadda_pg_rca32_and_9_14[0], h_s_dadda_pg_rca32_and_8_15[0], h_s_dadda_pg_rca32_fa162_xor1, h_s_dadda_pg_rca32_fa162_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_16(a[7], b[16], h_s_dadda_pg_rca32_and_7_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_17(a[6], b[17], h_s_dadda_pg_rca32_and_6_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_18(a[5], b[18], h_s_dadda_pg_rca32_and_5_18);
  fa fa_h_s_dadda_pg_rca32_fa163_out(h_s_dadda_pg_rca32_and_7_16[0], h_s_dadda_pg_rca32_and_6_17[0], h_s_dadda_pg_rca32_and_5_18[0], h_s_dadda_pg_rca32_fa163_xor1, h_s_dadda_pg_rca32_fa163_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_19(a[4], b[19], h_s_dadda_pg_rca32_and_4_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_20(a[3], b[20], h_s_dadda_pg_rca32_and_3_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_21(a[2], b[21], h_s_dadda_pg_rca32_and_2_21);
  fa fa_h_s_dadda_pg_rca32_fa164_out(h_s_dadda_pg_rca32_and_4_19[0], h_s_dadda_pg_rca32_and_3_20[0], h_s_dadda_pg_rca32_and_2_21[0], h_s_dadda_pg_rca32_fa164_xor1, h_s_dadda_pg_rca32_fa164_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_22(a[1], b[22], h_s_dadda_pg_rca32_and_1_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_23(a[0], b[23], h_s_dadda_pg_rca32_and_0_23);
  fa fa_h_s_dadda_pg_rca32_fa165_out(h_s_dadda_pg_rca32_and_1_22[0], h_s_dadda_pg_rca32_and_0_23[0], h_s_dadda_pg_rca32_fa152_xor1[0], h_s_dadda_pg_rca32_fa165_xor1, h_s_dadda_pg_rca32_fa165_or0);
  fa fa_h_s_dadda_pg_rca32_fa166_out(h_s_dadda_pg_rca32_fa153_xor1[0], h_s_dadda_pg_rca32_fa154_xor1[0], h_s_dadda_pg_rca32_fa155_xor1[0], h_s_dadda_pg_rca32_fa166_xor1, h_s_dadda_pg_rca32_fa166_or0);
  fa fa_h_s_dadda_pg_rca32_fa167_out(h_s_dadda_pg_rca32_fa156_xor1[0], h_s_dadda_pg_rca32_fa157_xor1[0], h_s_dadda_pg_rca32_fa158_xor1[0], h_s_dadda_pg_rca32_fa167_xor1, h_s_dadda_pg_rca32_fa167_or0);
  fa fa_h_s_dadda_pg_rca32_fa168_out(h_s_dadda_pg_rca32_fa159_xor1[0], h_s_dadda_pg_rca32_fa160_xor1[0], h_s_dadda_pg_rca32_fa161_xor1[0], h_s_dadda_pg_rca32_fa168_xor1, h_s_dadda_pg_rca32_fa168_or0);
  ha ha_h_s_dadda_pg_rca32_ha21_out(h_s_dadda_pg_rca32_fa162_xor1[0], h_s_dadda_pg_rca32_fa163_xor1[0], h_s_dadda_pg_rca32_ha21_xor0, h_s_dadda_pg_rca32_ha21_and0);
  fa fa_h_s_dadda_pg_rca32_fa169_out(h_s_dadda_pg_rca32_ha21_and0[0], h_s_dadda_pg_rca32_fa168_or0[0], h_s_dadda_pg_rca32_fa167_or0[0], h_s_dadda_pg_rca32_fa169_xor1, h_s_dadda_pg_rca32_fa169_or0);
  fa fa_h_s_dadda_pg_rca32_fa170_out(h_s_dadda_pg_rca32_fa166_or0[0], h_s_dadda_pg_rca32_fa165_or0[0], h_s_dadda_pg_rca32_fa164_or0[0], h_s_dadda_pg_rca32_fa170_xor1, h_s_dadda_pg_rca32_fa170_or0);
  fa fa_h_s_dadda_pg_rca32_fa171_out(h_s_dadda_pg_rca32_fa163_or0[0], h_s_dadda_pg_rca32_fa162_or0[0], h_s_dadda_pg_rca32_fa161_or0[0], h_s_dadda_pg_rca32_fa171_xor1, h_s_dadda_pg_rca32_fa171_or0);
  fa fa_h_s_dadda_pg_rca32_fa172_out(h_s_dadda_pg_rca32_fa160_or0[0], h_s_dadda_pg_rca32_fa159_or0[0], h_s_dadda_pg_rca32_fa158_or0[0], h_s_dadda_pg_rca32_fa172_xor1, h_s_dadda_pg_rca32_fa172_or0);
  fa fa_h_s_dadda_pg_rca32_fa173_out(h_s_dadda_pg_rca32_fa157_or0[0], h_s_dadda_pg_rca32_fa156_or0[0], h_s_dadda_pg_rca32_fa155_or0[0], h_s_dadda_pg_rca32_fa173_xor1, h_s_dadda_pg_rca32_fa173_or0);
  fa fa_h_s_dadda_pg_rca32_fa174_out(h_s_dadda_pg_rca32_fa154_or0[0], h_s_dadda_pg_rca32_fa153_or0[0], h_s_dadda_pg_rca32_fa152_or0[0], h_s_dadda_pg_rca32_fa174_xor1, h_s_dadda_pg_rca32_fa174_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_0(a[24], b[0], h_s_dadda_pg_rca32_and_24_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_1(a[23], b[1], h_s_dadda_pg_rca32_and_23_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_2(a[22], b[2], h_s_dadda_pg_rca32_and_22_2);
  fa fa_h_s_dadda_pg_rca32_fa175_out(h_s_dadda_pg_rca32_and_24_0[0], h_s_dadda_pg_rca32_and_23_1[0], h_s_dadda_pg_rca32_and_22_2[0], h_s_dadda_pg_rca32_fa175_xor1, h_s_dadda_pg_rca32_fa175_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_3(a[21], b[3], h_s_dadda_pg_rca32_and_21_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_4(a[20], b[4], h_s_dadda_pg_rca32_and_20_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_5(a[19], b[5], h_s_dadda_pg_rca32_and_19_5);
  fa fa_h_s_dadda_pg_rca32_fa176_out(h_s_dadda_pg_rca32_and_21_3[0], h_s_dadda_pg_rca32_and_20_4[0], h_s_dadda_pg_rca32_and_19_5[0], h_s_dadda_pg_rca32_fa176_xor1, h_s_dadda_pg_rca32_fa176_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_6(a[18], b[6], h_s_dadda_pg_rca32_and_18_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_7(a[17], b[7], h_s_dadda_pg_rca32_and_17_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_8(a[16], b[8], h_s_dadda_pg_rca32_and_16_8);
  fa fa_h_s_dadda_pg_rca32_fa177_out(h_s_dadda_pg_rca32_and_18_6[0], h_s_dadda_pg_rca32_and_17_7[0], h_s_dadda_pg_rca32_and_16_8[0], h_s_dadda_pg_rca32_fa177_xor1, h_s_dadda_pg_rca32_fa177_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_9(a[15], b[9], h_s_dadda_pg_rca32_and_15_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_10(a[14], b[10], h_s_dadda_pg_rca32_and_14_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_11(a[13], b[11], h_s_dadda_pg_rca32_and_13_11);
  fa fa_h_s_dadda_pg_rca32_fa178_out(h_s_dadda_pg_rca32_and_15_9[0], h_s_dadda_pg_rca32_and_14_10[0], h_s_dadda_pg_rca32_and_13_11[0], h_s_dadda_pg_rca32_fa178_xor1, h_s_dadda_pg_rca32_fa178_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_12(a[12], b[12], h_s_dadda_pg_rca32_and_12_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_13(a[11], b[13], h_s_dadda_pg_rca32_and_11_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_14(a[10], b[14], h_s_dadda_pg_rca32_and_10_14);
  fa fa_h_s_dadda_pg_rca32_fa179_out(h_s_dadda_pg_rca32_and_12_12[0], h_s_dadda_pg_rca32_and_11_13[0], h_s_dadda_pg_rca32_and_10_14[0], h_s_dadda_pg_rca32_fa179_xor1, h_s_dadda_pg_rca32_fa179_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_15(a[9], b[15], h_s_dadda_pg_rca32_and_9_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_16(a[8], b[16], h_s_dadda_pg_rca32_and_8_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_17(a[7], b[17], h_s_dadda_pg_rca32_and_7_17);
  fa fa_h_s_dadda_pg_rca32_fa180_out(h_s_dadda_pg_rca32_and_9_15[0], h_s_dadda_pg_rca32_and_8_16[0], h_s_dadda_pg_rca32_and_7_17[0], h_s_dadda_pg_rca32_fa180_xor1, h_s_dadda_pg_rca32_fa180_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_18(a[6], b[18], h_s_dadda_pg_rca32_and_6_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_19(a[5], b[19], h_s_dadda_pg_rca32_and_5_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_20(a[4], b[20], h_s_dadda_pg_rca32_and_4_20);
  fa fa_h_s_dadda_pg_rca32_fa181_out(h_s_dadda_pg_rca32_and_6_18[0], h_s_dadda_pg_rca32_and_5_19[0], h_s_dadda_pg_rca32_and_4_20[0], h_s_dadda_pg_rca32_fa181_xor1, h_s_dadda_pg_rca32_fa181_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_21(a[3], b[21], h_s_dadda_pg_rca32_and_3_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_22(a[2], b[22], h_s_dadda_pg_rca32_and_2_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_23(a[1], b[23], h_s_dadda_pg_rca32_and_1_23);
  fa fa_h_s_dadda_pg_rca32_fa182_out(h_s_dadda_pg_rca32_and_3_21[0], h_s_dadda_pg_rca32_and_2_22[0], h_s_dadda_pg_rca32_and_1_23[0], h_s_dadda_pg_rca32_fa182_xor1, h_s_dadda_pg_rca32_fa182_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_24(a[0], b[24], h_s_dadda_pg_rca32_and_0_24);
  fa fa_h_s_dadda_pg_rca32_fa183_out(h_s_dadda_pg_rca32_and_0_24[0], h_s_dadda_pg_rca32_fa169_xor1[0], h_s_dadda_pg_rca32_fa170_xor1[0], h_s_dadda_pg_rca32_fa183_xor1, h_s_dadda_pg_rca32_fa183_or0);
  fa fa_h_s_dadda_pg_rca32_fa184_out(h_s_dadda_pg_rca32_fa171_xor1[0], h_s_dadda_pg_rca32_fa172_xor1[0], h_s_dadda_pg_rca32_fa173_xor1[0], h_s_dadda_pg_rca32_fa184_xor1, h_s_dadda_pg_rca32_fa184_or0);
  fa fa_h_s_dadda_pg_rca32_fa185_out(h_s_dadda_pg_rca32_fa174_xor1[0], h_s_dadda_pg_rca32_fa175_xor1[0], h_s_dadda_pg_rca32_fa176_xor1[0], h_s_dadda_pg_rca32_fa185_xor1, h_s_dadda_pg_rca32_fa185_or0);
  fa fa_h_s_dadda_pg_rca32_fa186_out(h_s_dadda_pg_rca32_fa177_xor1[0], h_s_dadda_pg_rca32_fa178_xor1[0], h_s_dadda_pg_rca32_fa179_xor1[0], h_s_dadda_pg_rca32_fa186_xor1, h_s_dadda_pg_rca32_fa186_or0);
  ha ha_h_s_dadda_pg_rca32_ha22_out(h_s_dadda_pg_rca32_fa180_xor1[0], h_s_dadda_pg_rca32_fa181_xor1[0], h_s_dadda_pg_rca32_ha22_xor0, h_s_dadda_pg_rca32_ha22_and0);
  fa fa_h_s_dadda_pg_rca32_fa187_out(h_s_dadda_pg_rca32_ha22_and0[0], h_s_dadda_pg_rca32_fa186_or0[0], h_s_dadda_pg_rca32_fa185_or0[0], h_s_dadda_pg_rca32_fa187_xor1, h_s_dadda_pg_rca32_fa187_or0);
  fa fa_h_s_dadda_pg_rca32_fa188_out(h_s_dadda_pg_rca32_fa184_or0[0], h_s_dadda_pg_rca32_fa183_or0[0], h_s_dadda_pg_rca32_fa182_or0[0], h_s_dadda_pg_rca32_fa188_xor1, h_s_dadda_pg_rca32_fa188_or0);
  fa fa_h_s_dadda_pg_rca32_fa189_out(h_s_dadda_pg_rca32_fa181_or0[0], h_s_dadda_pg_rca32_fa180_or0[0], h_s_dadda_pg_rca32_fa179_or0[0], h_s_dadda_pg_rca32_fa189_xor1, h_s_dadda_pg_rca32_fa189_or0);
  fa fa_h_s_dadda_pg_rca32_fa190_out(h_s_dadda_pg_rca32_fa178_or0[0], h_s_dadda_pg_rca32_fa177_or0[0], h_s_dadda_pg_rca32_fa176_or0[0], h_s_dadda_pg_rca32_fa190_xor1, h_s_dadda_pg_rca32_fa190_or0);
  fa fa_h_s_dadda_pg_rca32_fa191_out(h_s_dadda_pg_rca32_fa175_or0[0], h_s_dadda_pg_rca32_fa174_or0[0], h_s_dadda_pg_rca32_fa173_or0[0], h_s_dadda_pg_rca32_fa191_xor1, h_s_dadda_pg_rca32_fa191_or0);
  fa fa_h_s_dadda_pg_rca32_fa192_out(h_s_dadda_pg_rca32_fa172_or0[0], h_s_dadda_pg_rca32_fa171_or0[0], h_s_dadda_pg_rca32_fa170_or0[0], h_s_dadda_pg_rca32_fa192_xor1, h_s_dadda_pg_rca32_fa192_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_0(a[25], b[0], h_s_dadda_pg_rca32_and_25_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_1(a[24], b[1], h_s_dadda_pg_rca32_and_24_1);
  fa fa_h_s_dadda_pg_rca32_fa193_out(h_s_dadda_pg_rca32_fa169_or0[0], h_s_dadda_pg_rca32_and_25_0[0], h_s_dadda_pg_rca32_and_24_1[0], h_s_dadda_pg_rca32_fa193_xor1, h_s_dadda_pg_rca32_fa193_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_2(a[23], b[2], h_s_dadda_pg_rca32_and_23_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_3(a[22], b[3], h_s_dadda_pg_rca32_and_22_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_4(a[21], b[4], h_s_dadda_pg_rca32_and_21_4);
  fa fa_h_s_dadda_pg_rca32_fa194_out(h_s_dadda_pg_rca32_and_23_2[0], h_s_dadda_pg_rca32_and_22_3[0], h_s_dadda_pg_rca32_and_21_4[0], h_s_dadda_pg_rca32_fa194_xor1, h_s_dadda_pg_rca32_fa194_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_5(a[20], b[5], h_s_dadda_pg_rca32_and_20_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_6(a[19], b[6], h_s_dadda_pg_rca32_and_19_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_7(a[18], b[7], h_s_dadda_pg_rca32_and_18_7);
  fa fa_h_s_dadda_pg_rca32_fa195_out(h_s_dadda_pg_rca32_and_20_5[0], h_s_dadda_pg_rca32_and_19_6[0], h_s_dadda_pg_rca32_and_18_7[0], h_s_dadda_pg_rca32_fa195_xor1, h_s_dadda_pg_rca32_fa195_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_8(a[17], b[8], h_s_dadda_pg_rca32_and_17_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_9(a[16], b[9], h_s_dadda_pg_rca32_and_16_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_10(a[15], b[10], h_s_dadda_pg_rca32_and_15_10);
  fa fa_h_s_dadda_pg_rca32_fa196_out(h_s_dadda_pg_rca32_and_17_8[0], h_s_dadda_pg_rca32_and_16_9[0], h_s_dadda_pg_rca32_and_15_10[0], h_s_dadda_pg_rca32_fa196_xor1, h_s_dadda_pg_rca32_fa196_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_11(a[14], b[11], h_s_dadda_pg_rca32_and_14_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_12(a[13], b[12], h_s_dadda_pg_rca32_and_13_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_13(a[12], b[13], h_s_dadda_pg_rca32_and_12_13);
  fa fa_h_s_dadda_pg_rca32_fa197_out(h_s_dadda_pg_rca32_and_14_11[0], h_s_dadda_pg_rca32_and_13_12[0], h_s_dadda_pg_rca32_and_12_13[0], h_s_dadda_pg_rca32_fa197_xor1, h_s_dadda_pg_rca32_fa197_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_14(a[11], b[14], h_s_dadda_pg_rca32_and_11_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_15(a[10], b[15], h_s_dadda_pg_rca32_and_10_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_16(a[9], b[16], h_s_dadda_pg_rca32_and_9_16);
  fa fa_h_s_dadda_pg_rca32_fa198_out(h_s_dadda_pg_rca32_and_11_14[0], h_s_dadda_pg_rca32_and_10_15[0], h_s_dadda_pg_rca32_and_9_16[0], h_s_dadda_pg_rca32_fa198_xor1, h_s_dadda_pg_rca32_fa198_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_17(a[8], b[17], h_s_dadda_pg_rca32_and_8_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_18(a[7], b[18], h_s_dadda_pg_rca32_and_7_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_19(a[6], b[19], h_s_dadda_pg_rca32_and_6_19);
  fa fa_h_s_dadda_pg_rca32_fa199_out(h_s_dadda_pg_rca32_and_8_17[0], h_s_dadda_pg_rca32_and_7_18[0], h_s_dadda_pg_rca32_and_6_19[0], h_s_dadda_pg_rca32_fa199_xor1, h_s_dadda_pg_rca32_fa199_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_20(a[5], b[20], h_s_dadda_pg_rca32_and_5_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_21(a[4], b[21], h_s_dadda_pg_rca32_and_4_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_22(a[3], b[22], h_s_dadda_pg_rca32_and_3_22);
  fa fa_h_s_dadda_pg_rca32_fa200_out(h_s_dadda_pg_rca32_and_5_20[0], h_s_dadda_pg_rca32_and_4_21[0], h_s_dadda_pg_rca32_and_3_22[0], h_s_dadda_pg_rca32_fa200_xor1, h_s_dadda_pg_rca32_fa200_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_23(a[2], b[23], h_s_dadda_pg_rca32_and_2_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_24(a[1], b[24], h_s_dadda_pg_rca32_and_1_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_25(a[0], b[25], h_s_dadda_pg_rca32_and_0_25);
  fa fa_h_s_dadda_pg_rca32_fa201_out(h_s_dadda_pg_rca32_and_2_23[0], h_s_dadda_pg_rca32_and_1_24[0], h_s_dadda_pg_rca32_and_0_25[0], h_s_dadda_pg_rca32_fa201_xor1, h_s_dadda_pg_rca32_fa201_or0);
  fa fa_h_s_dadda_pg_rca32_fa202_out(h_s_dadda_pg_rca32_fa187_xor1[0], h_s_dadda_pg_rca32_fa188_xor1[0], h_s_dadda_pg_rca32_fa189_xor1[0], h_s_dadda_pg_rca32_fa202_xor1, h_s_dadda_pg_rca32_fa202_or0);
  fa fa_h_s_dadda_pg_rca32_fa203_out(h_s_dadda_pg_rca32_fa190_xor1[0], h_s_dadda_pg_rca32_fa191_xor1[0], h_s_dadda_pg_rca32_fa192_xor1[0], h_s_dadda_pg_rca32_fa203_xor1, h_s_dadda_pg_rca32_fa203_or0);
  fa fa_h_s_dadda_pg_rca32_fa204_out(h_s_dadda_pg_rca32_fa193_xor1[0], h_s_dadda_pg_rca32_fa194_xor1[0], h_s_dadda_pg_rca32_fa195_xor1[0], h_s_dadda_pg_rca32_fa204_xor1, h_s_dadda_pg_rca32_fa204_or0);
  fa fa_h_s_dadda_pg_rca32_fa205_out(h_s_dadda_pg_rca32_fa196_xor1[0], h_s_dadda_pg_rca32_fa197_xor1[0], h_s_dadda_pg_rca32_fa198_xor1[0], h_s_dadda_pg_rca32_fa205_xor1, h_s_dadda_pg_rca32_fa205_or0);
  ha ha_h_s_dadda_pg_rca32_ha23_out(h_s_dadda_pg_rca32_fa199_xor1[0], h_s_dadda_pg_rca32_fa200_xor1[0], h_s_dadda_pg_rca32_ha23_xor0, h_s_dadda_pg_rca32_ha23_and0);
  fa fa_h_s_dadda_pg_rca32_fa206_out(h_s_dadda_pg_rca32_ha23_and0[0], h_s_dadda_pg_rca32_fa205_or0[0], h_s_dadda_pg_rca32_fa204_or0[0], h_s_dadda_pg_rca32_fa206_xor1, h_s_dadda_pg_rca32_fa206_or0);
  fa fa_h_s_dadda_pg_rca32_fa207_out(h_s_dadda_pg_rca32_fa203_or0[0], h_s_dadda_pg_rca32_fa202_or0[0], h_s_dadda_pg_rca32_fa201_or0[0], h_s_dadda_pg_rca32_fa207_xor1, h_s_dadda_pg_rca32_fa207_or0);
  fa fa_h_s_dadda_pg_rca32_fa208_out(h_s_dadda_pg_rca32_fa200_or0[0], h_s_dadda_pg_rca32_fa199_or0[0], h_s_dadda_pg_rca32_fa198_or0[0], h_s_dadda_pg_rca32_fa208_xor1, h_s_dadda_pg_rca32_fa208_or0);
  fa fa_h_s_dadda_pg_rca32_fa209_out(h_s_dadda_pg_rca32_fa197_or0[0], h_s_dadda_pg_rca32_fa196_or0[0], h_s_dadda_pg_rca32_fa195_or0[0], h_s_dadda_pg_rca32_fa209_xor1, h_s_dadda_pg_rca32_fa209_or0);
  fa fa_h_s_dadda_pg_rca32_fa210_out(h_s_dadda_pg_rca32_fa194_or0[0], h_s_dadda_pg_rca32_fa193_or0[0], h_s_dadda_pg_rca32_fa192_or0[0], h_s_dadda_pg_rca32_fa210_xor1, h_s_dadda_pg_rca32_fa210_or0);
  fa fa_h_s_dadda_pg_rca32_fa211_out(h_s_dadda_pg_rca32_fa191_or0[0], h_s_dadda_pg_rca32_fa190_or0[0], h_s_dadda_pg_rca32_fa189_or0[0], h_s_dadda_pg_rca32_fa211_xor1, h_s_dadda_pg_rca32_fa211_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_0(a[26], b[0], h_s_dadda_pg_rca32_and_26_0);
  fa fa_h_s_dadda_pg_rca32_fa212_out(h_s_dadda_pg_rca32_fa188_or0[0], h_s_dadda_pg_rca32_fa187_or0[0], h_s_dadda_pg_rca32_and_26_0[0], h_s_dadda_pg_rca32_fa212_xor1, h_s_dadda_pg_rca32_fa212_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_1(a[25], b[1], h_s_dadda_pg_rca32_and_25_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_2(a[24], b[2], h_s_dadda_pg_rca32_and_24_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_3(a[23], b[3], h_s_dadda_pg_rca32_and_23_3);
  fa fa_h_s_dadda_pg_rca32_fa213_out(h_s_dadda_pg_rca32_and_25_1[0], h_s_dadda_pg_rca32_and_24_2[0], h_s_dadda_pg_rca32_and_23_3[0], h_s_dadda_pg_rca32_fa213_xor1, h_s_dadda_pg_rca32_fa213_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_4(a[22], b[4], h_s_dadda_pg_rca32_and_22_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_5(a[21], b[5], h_s_dadda_pg_rca32_and_21_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_6(a[20], b[6], h_s_dadda_pg_rca32_and_20_6);
  fa fa_h_s_dadda_pg_rca32_fa214_out(h_s_dadda_pg_rca32_and_22_4[0], h_s_dadda_pg_rca32_and_21_5[0], h_s_dadda_pg_rca32_and_20_6[0], h_s_dadda_pg_rca32_fa214_xor1, h_s_dadda_pg_rca32_fa214_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_7(a[19], b[7], h_s_dadda_pg_rca32_and_19_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_8(a[18], b[8], h_s_dadda_pg_rca32_and_18_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_9(a[17], b[9], h_s_dadda_pg_rca32_and_17_9);
  fa fa_h_s_dadda_pg_rca32_fa215_out(h_s_dadda_pg_rca32_and_19_7[0], h_s_dadda_pg_rca32_and_18_8[0], h_s_dadda_pg_rca32_and_17_9[0], h_s_dadda_pg_rca32_fa215_xor1, h_s_dadda_pg_rca32_fa215_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_10(a[16], b[10], h_s_dadda_pg_rca32_and_16_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_11(a[15], b[11], h_s_dadda_pg_rca32_and_15_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_12(a[14], b[12], h_s_dadda_pg_rca32_and_14_12);
  fa fa_h_s_dadda_pg_rca32_fa216_out(h_s_dadda_pg_rca32_and_16_10[0], h_s_dadda_pg_rca32_and_15_11[0], h_s_dadda_pg_rca32_and_14_12[0], h_s_dadda_pg_rca32_fa216_xor1, h_s_dadda_pg_rca32_fa216_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_13(a[13], b[13], h_s_dadda_pg_rca32_and_13_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_14(a[12], b[14], h_s_dadda_pg_rca32_and_12_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_15(a[11], b[15], h_s_dadda_pg_rca32_and_11_15);
  fa fa_h_s_dadda_pg_rca32_fa217_out(h_s_dadda_pg_rca32_and_13_13[0], h_s_dadda_pg_rca32_and_12_14[0], h_s_dadda_pg_rca32_and_11_15[0], h_s_dadda_pg_rca32_fa217_xor1, h_s_dadda_pg_rca32_fa217_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_16(a[10], b[16], h_s_dadda_pg_rca32_and_10_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_17(a[9], b[17], h_s_dadda_pg_rca32_and_9_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_18(a[8], b[18], h_s_dadda_pg_rca32_and_8_18);
  fa fa_h_s_dadda_pg_rca32_fa218_out(h_s_dadda_pg_rca32_and_10_16[0], h_s_dadda_pg_rca32_and_9_17[0], h_s_dadda_pg_rca32_and_8_18[0], h_s_dadda_pg_rca32_fa218_xor1, h_s_dadda_pg_rca32_fa218_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_19(a[7], b[19], h_s_dadda_pg_rca32_and_7_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_20(a[6], b[20], h_s_dadda_pg_rca32_and_6_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_21(a[5], b[21], h_s_dadda_pg_rca32_and_5_21);
  fa fa_h_s_dadda_pg_rca32_fa219_out(h_s_dadda_pg_rca32_and_7_19[0], h_s_dadda_pg_rca32_and_6_20[0], h_s_dadda_pg_rca32_and_5_21[0], h_s_dadda_pg_rca32_fa219_xor1, h_s_dadda_pg_rca32_fa219_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_22(a[4], b[22], h_s_dadda_pg_rca32_and_4_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_23(a[3], b[23], h_s_dadda_pg_rca32_and_3_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_24(a[2], b[24], h_s_dadda_pg_rca32_and_2_24);
  fa fa_h_s_dadda_pg_rca32_fa220_out(h_s_dadda_pg_rca32_and_4_22[0], h_s_dadda_pg_rca32_and_3_23[0], h_s_dadda_pg_rca32_and_2_24[0], h_s_dadda_pg_rca32_fa220_xor1, h_s_dadda_pg_rca32_fa220_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_25(a[1], b[25], h_s_dadda_pg_rca32_and_1_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_26(a[0], b[26], h_s_dadda_pg_rca32_and_0_26);
  fa fa_h_s_dadda_pg_rca32_fa221_out(h_s_dadda_pg_rca32_and_1_25[0], h_s_dadda_pg_rca32_and_0_26[0], h_s_dadda_pg_rca32_fa206_xor1[0], h_s_dadda_pg_rca32_fa221_xor1, h_s_dadda_pg_rca32_fa221_or0);
  fa fa_h_s_dadda_pg_rca32_fa222_out(h_s_dadda_pg_rca32_fa207_xor1[0], h_s_dadda_pg_rca32_fa208_xor1[0], h_s_dadda_pg_rca32_fa209_xor1[0], h_s_dadda_pg_rca32_fa222_xor1, h_s_dadda_pg_rca32_fa222_or0);
  fa fa_h_s_dadda_pg_rca32_fa223_out(h_s_dadda_pg_rca32_fa210_xor1[0], h_s_dadda_pg_rca32_fa211_xor1[0], h_s_dadda_pg_rca32_fa212_xor1[0], h_s_dadda_pg_rca32_fa223_xor1, h_s_dadda_pg_rca32_fa223_or0);
  fa fa_h_s_dadda_pg_rca32_fa224_out(h_s_dadda_pg_rca32_fa213_xor1[0], h_s_dadda_pg_rca32_fa214_xor1[0], h_s_dadda_pg_rca32_fa215_xor1[0], h_s_dadda_pg_rca32_fa224_xor1, h_s_dadda_pg_rca32_fa224_or0);
  fa fa_h_s_dadda_pg_rca32_fa225_out(h_s_dadda_pg_rca32_fa216_xor1[0], h_s_dadda_pg_rca32_fa217_xor1[0], h_s_dadda_pg_rca32_fa218_xor1[0], h_s_dadda_pg_rca32_fa225_xor1, h_s_dadda_pg_rca32_fa225_or0);
  ha ha_h_s_dadda_pg_rca32_ha24_out(h_s_dadda_pg_rca32_fa219_xor1[0], h_s_dadda_pg_rca32_fa220_xor1[0], h_s_dadda_pg_rca32_ha24_xor0, h_s_dadda_pg_rca32_ha24_and0);
  fa fa_h_s_dadda_pg_rca32_fa226_out(h_s_dadda_pg_rca32_ha24_and0[0], h_s_dadda_pg_rca32_fa225_or0[0], h_s_dadda_pg_rca32_fa224_or0[0], h_s_dadda_pg_rca32_fa226_xor1, h_s_dadda_pg_rca32_fa226_or0);
  fa fa_h_s_dadda_pg_rca32_fa227_out(h_s_dadda_pg_rca32_fa223_or0[0], h_s_dadda_pg_rca32_fa222_or0[0], h_s_dadda_pg_rca32_fa221_or0[0], h_s_dadda_pg_rca32_fa227_xor1, h_s_dadda_pg_rca32_fa227_or0);
  fa fa_h_s_dadda_pg_rca32_fa228_out(h_s_dadda_pg_rca32_fa220_or0[0], h_s_dadda_pg_rca32_fa219_or0[0], h_s_dadda_pg_rca32_fa218_or0[0], h_s_dadda_pg_rca32_fa228_xor1, h_s_dadda_pg_rca32_fa228_or0);
  fa fa_h_s_dadda_pg_rca32_fa229_out(h_s_dadda_pg_rca32_fa217_or0[0], h_s_dadda_pg_rca32_fa216_or0[0], h_s_dadda_pg_rca32_fa215_or0[0], h_s_dadda_pg_rca32_fa229_xor1, h_s_dadda_pg_rca32_fa229_or0);
  fa fa_h_s_dadda_pg_rca32_fa230_out(h_s_dadda_pg_rca32_fa214_or0[0], h_s_dadda_pg_rca32_fa213_or0[0], h_s_dadda_pg_rca32_fa212_or0[0], h_s_dadda_pg_rca32_fa230_xor1, h_s_dadda_pg_rca32_fa230_or0);
  fa fa_h_s_dadda_pg_rca32_fa231_out(h_s_dadda_pg_rca32_fa211_or0[0], h_s_dadda_pg_rca32_fa210_or0[0], h_s_dadda_pg_rca32_fa209_or0[0], h_s_dadda_pg_rca32_fa231_xor1, h_s_dadda_pg_rca32_fa231_or0);
  fa fa_h_s_dadda_pg_rca32_fa232_out(h_s_dadda_pg_rca32_fa208_or0[0], h_s_dadda_pg_rca32_fa207_or0[0], h_s_dadda_pg_rca32_fa206_or0[0], h_s_dadda_pg_rca32_fa232_xor1, h_s_dadda_pg_rca32_fa232_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_0(a[27], b[0], h_s_dadda_pg_rca32_and_27_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_1(a[26], b[1], h_s_dadda_pg_rca32_and_26_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_2(a[25], b[2], h_s_dadda_pg_rca32_and_25_2);
  fa fa_h_s_dadda_pg_rca32_fa233_out(h_s_dadda_pg_rca32_and_27_0[0], h_s_dadda_pg_rca32_and_26_1[0], h_s_dadda_pg_rca32_and_25_2[0], h_s_dadda_pg_rca32_fa233_xor1, h_s_dadda_pg_rca32_fa233_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_3(a[24], b[3], h_s_dadda_pg_rca32_and_24_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_4(a[23], b[4], h_s_dadda_pg_rca32_and_23_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_5(a[22], b[5], h_s_dadda_pg_rca32_and_22_5);
  fa fa_h_s_dadda_pg_rca32_fa234_out(h_s_dadda_pg_rca32_and_24_3[0], h_s_dadda_pg_rca32_and_23_4[0], h_s_dadda_pg_rca32_and_22_5[0], h_s_dadda_pg_rca32_fa234_xor1, h_s_dadda_pg_rca32_fa234_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_6(a[21], b[6], h_s_dadda_pg_rca32_and_21_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_7(a[20], b[7], h_s_dadda_pg_rca32_and_20_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_8(a[19], b[8], h_s_dadda_pg_rca32_and_19_8);
  fa fa_h_s_dadda_pg_rca32_fa235_out(h_s_dadda_pg_rca32_and_21_6[0], h_s_dadda_pg_rca32_and_20_7[0], h_s_dadda_pg_rca32_and_19_8[0], h_s_dadda_pg_rca32_fa235_xor1, h_s_dadda_pg_rca32_fa235_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_9(a[18], b[9], h_s_dadda_pg_rca32_and_18_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_10(a[17], b[10], h_s_dadda_pg_rca32_and_17_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_11(a[16], b[11], h_s_dadda_pg_rca32_and_16_11);
  fa fa_h_s_dadda_pg_rca32_fa236_out(h_s_dadda_pg_rca32_and_18_9[0], h_s_dadda_pg_rca32_and_17_10[0], h_s_dadda_pg_rca32_and_16_11[0], h_s_dadda_pg_rca32_fa236_xor1, h_s_dadda_pg_rca32_fa236_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_12(a[15], b[12], h_s_dadda_pg_rca32_and_15_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_13(a[14], b[13], h_s_dadda_pg_rca32_and_14_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_14(a[13], b[14], h_s_dadda_pg_rca32_and_13_14);
  fa fa_h_s_dadda_pg_rca32_fa237_out(h_s_dadda_pg_rca32_and_15_12[0], h_s_dadda_pg_rca32_and_14_13[0], h_s_dadda_pg_rca32_and_13_14[0], h_s_dadda_pg_rca32_fa237_xor1, h_s_dadda_pg_rca32_fa237_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_15(a[12], b[15], h_s_dadda_pg_rca32_and_12_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_16(a[11], b[16], h_s_dadda_pg_rca32_and_11_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_17(a[10], b[17], h_s_dadda_pg_rca32_and_10_17);
  fa fa_h_s_dadda_pg_rca32_fa238_out(h_s_dadda_pg_rca32_and_12_15[0], h_s_dadda_pg_rca32_and_11_16[0], h_s_dadda_pg_rca32_and_10_17[0], h_s_dadda_pg_rca32_fa238_xor1, h_s_dadda_pg_rca32_fa238_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_18(a[9], b[18], h_s_dadda_pg_rca32_and_9_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_19(a[8], b[19], h_s_dadda_pg_rca32_and_8_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_20(a[7], b[20], h_s_dadda_pg_rca32_and_7_20);
  fa fa_h_s_dadda_pg_rca32_fa239_out(h_s_dadda_pg_rca32_and_9_18[0], h_s_dadda_pg_rca32_and_8_19[0], h_s_dadda_pg_rca32_and_7_20[0], h_s_dadda_pg_rca32_fa239_xor1, h_s_dadda_pg_rca32_fa239_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_21(a[6], b[21], h_s_dadda_pg_rca32_and_6_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_22(a[5], b[22], h_s_dadda_pg_rca32_and_5_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_23(a[4], b[23], h_s_dadda_pg_rca32_and_4_23);
  fa fa_h_s_dadda_pg_rca32_fa240_out(h_s_dadda_pg_rca32_and_6_21[0], h_s_dadda_pg_rca32_and_5_22[0], h_s_dadda_pg_rca32_and_4_23[0], h_s_dadda_pg_rca32_fa240_xor1, h_s_dadda_pg_rca32_fa240_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_24(a[3], b[24], h_s_dadda_pg_rca32_and_3_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_25(a[2], b[25], h_s_dadda_pg_rca32_and_2_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_26(a[1], b[26], h_s_dadda_pg_rca32_and_1_26);
  fa fa_h_s_dadda_pg_rca32_fa241_out(h_s_dadda_pg_rca32_and_3_24[0], h_s_dadda_pg_rca32_and_2_25[0], h_s_dadda_pg_rca32_and_1_26[0], h_s_dadda_pg_rca32_fa241_xor1, h_s_dadda_pg_rca32_fa241_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_27(a[0], b[27], h_s_dadda_pg_rca32_and_0_27);
  fa fa_h_s_dadda_pg_rca32_fa242_out(h_s_dadda_pg_rca32_and_0_27[0], h_s_dadda_pg_rca32_fa226_xor1[0], h_s_dadda_pg_rca32_fa227_xor1[0], h_s_dadda_pg_rca32_fa242_xor1, h_s_dadda_pg_rca32_fa242_or0);
  fa fa_h_s_dadda_pg_rca32_fa243_out(h_s_dadda_pg_rca32_fa228_xor1[0], h_s_dadda_pg_rca32_fa229_xor1[0], h_s_dadda_pg_rca32_fa230_xor1[0], h_s_dadda_pg_rca32_fa243_xor1, h_s_dadda_pg_rca32_fa243_or0);
  fa fa_h_s_dadda_pg_rca32_fa244_out(h_s_dadda_pg_rca32_fa231_xor1[0], h_s_dadda_pg_rca32_fa232_xor1[0], h_s_dadda_pg_rca32_fa233_xor1[0], h_s_dadda_pg_rca32_fa244_xor1, h_s_dadda_pg_rca32_fa244_or0);
  fa fa_h_s_dadda_pg_rca32_fa245_out(h_s_dadda_pg_rca32_fa234_xor1[0], h_s_dadda_pg_rca32_fa235_xor1[0], h_s_dadda_pg_rca32_fa236_xor1[0], h_s_dadda_pg_rca32_fa245_xor1, h_s_dadda_pg_rca32_fa245_or0);
  fa fa_h_s_dadda_pg_rca32_fa246_out(h_s_dadda_pg_rca32_fa237_xor1[0], h_s_dadda_pg_rca32_fa238_xor1[0], h_s_dadda_pg_rca32_fa239_xor1[0], h_s_dadda_pg_rca32_fa246_xor1, h_s_dadda_pg_rca32_fa246_or0);
  ha ha_h_s_dadda_pg_rca32_ha25_out(h_s_dadda_pg_rca32_fa240_xor1[0], h_s_dadda_pg_rca32_fa241_xor1[0], h_s_dadda_pg_rca32_ha25_xor0, h_s_dadda_pg_rca32_ha25_and0);
  fa fa_h_s_dadda_pg_rca32_fa247_out(h_s_dadda_pg_rca32_ha25_and0[0], h_s_dadda_pg_rca32_fa246_or0[0], h_s_dadda_pg_rca32_fa245_or0[0], h_s_dadda_pg_rca32_fa247_xor1, h_s_dadda_pg_rca32_fa247_or0);
  fa fa_h_s_dadda_pg_rca32_fa248_out(h_s_dadda_pg_rca32_fa244_or0[0], h_s_dadda_pg_rca32_fa243_or0[0], h_s_dadda_pg_rca32_fa242_or0[0], h_s_dadda_pg_rca32_fa248_xor1, h_s_dadda_pg_rca32_fa248_or0);
  fa fa_h_s_dadda_pg_rca32_fa249_out(h_s_dadda_pg_rca32_fa241_or0[0], h_s_dadda_pg_rca32_fa240_or0[0], h_s_dadda_pg_rca32_fa239_or0[0], h_s_dadda_pg_rca32_fa249_xor1, h_s_dadda_pg_rca32_fa249_or0);
  fa fa_h_s_dadda_pg_rca32_fa250_out(h_s_dadda_pg_rca32_fa238_or0[0], h_s_dadda_pg_rca32_fa237_or0[0], h_s_dadda_pg_rca32_fa236_or0[0], h_s_dadda_pg_rca32_fa250_xor1, h_s_dadda_pg_rca32_fa250_or0);
  fa fa_h_s_dadda_pg_rca32_fa251_out(h_s_dadda_pg_rca32_fa235_or0[0], h_s_dadda_pg_rca32_fa234_or0[0], h_s_dadda_pg_rca32_fa233_or0[0], h_s_dadda_pg_rca32_fa251_xor1, h_s_dadda_pg_rca32_fa251_or0);
  fa fa_h_s_dadda_pg_rca32_fa252_out(h_s_dadda_pg_rca32_fa232_or0[0], h_s_dadda_pg_rca32_fa231_or0[0], h_s_dadda_pg_rca32_fa230_or0[0], h_s_dadda_pg_rca32_fa252_xor1, h_s_dadda_pg_rca32_fa252_or0);
  fa fa_h_s_dadda_pg_rca32_fa253_out(h_s_dadda_pg_rca32_fa229_or0[0], h_s_dadda_pg_rca32_fa228_or0[0], h_s_dadda_pg_rca32_fa227_or0[0], h_s_dadda_pg_rca32_fa253_xor1, h_s_dadda_pg_rca32_fa253_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_2(a[26], b[2], h_s_dadda_pg_rca32_and_26_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_3(a[25], b[3], h_s_dadda_pg_rca32_and_25_3);
  fa fa_h_s_dadda_pg_rca32_fa254_out(h_s_dadda_pg_rca32_fa226_or0[0], h_s_dadda_pg_rca32_and_26_2[0], h_s_dadda_pg_rca32_and_25_3[0], h_s_dadda_pg_rca32_fa254_xor1, h_s_dadda_pg_rca32_fa254_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_4(a[24], b[4], h_s_dadda_pg_rca32_and_24_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_5(a[23], b[5], h_s_dadda_pg_rca32_and_23_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_6(a[22], b[6], h_s_dadda_pg_rca32_and_22_6);
  fa fa_h_s_dadda_pg_rca32_fa255_out(h_s_dadda_pg_rca32_and_24_4[0], h_s_dadda_pg_rca32_and_23_5[0], h_s_dadda_pg_rca32_and_22_6[0], h_s_dadda_pg_rca32_fa255_xor1, h_s_dadda_pg_rca32_fa255_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_7(a[21], b[7], h_s_dadda_pg_rca32_and_21_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_8(a[20], b[8], h_s_dadda_pg_rca32_and_20_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_9(a[19], b[9], h_s_dadda_pg_rca32_and_19_9);
  fa fa_h_s_dadda_pg_rca32_fa256_out(h_s_dadda_pg_rca32_and_21_7[0], h_s_dadda_pg_rca32_and_20_8[0], h_s_dadda_pg_rca32_and_19_9[0], h_s_dadda_pg_rca32_fa256_xor1, h_s_dadda_pg_rca32_fa256_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_10(a[18], b[10], h_s_dadda_pg_rca32_and_18_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_11(a[17], b[11], h_s_dadda_pg_rca32_and_17_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_12(a[16], b[12], h_s_dadda_pg_rca32_and_16_12);
  fa fa_h_s_dadda_pg_rca32_fa257_out(h_s_dadda_pg_rca32_and_18_10[0], h_s_dadda_pg_rca32_and_17_11[0], h_s_dadda_pg_rca32_and_16_12[0], h_s_dadda_pg_rca32_fa257_xor1, h_s_dadda_pg_rca32_fa257_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_13(a[15], b[13], h_s_dadda_pg_rca32_and_15_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_14(a[14], b[14], h_s_dadda_pg_rca32_and_14_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_15(a[13], b[15], h_s_dadda_pg_rca32_and_13_15);
  fa fa_h_s_dadda_pg_rca32_fa258_out(h_s_dadda_pg_rca32_and_15_13[0], h_s_dadda_pg_rca32_and_14_14[0], h_s_dadda_pg_rca32_and_13_15[0], h_s_dadda_pg_rca32_fa258_xor1, h_s_dadda_pg_rca32_fa258_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_16(a[12], b[16], h_s_dadda_pg_rca32_and_12_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_17(a[11], b[17], h_s_dadda_pg_rca32_and_11_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_18(a[10], b[18], h_s_dadda_pg_rca32_and_10_18);
  fa fa_h_s_dadda_pg_rca32_fa259_out(h_s_dadda_pg_rca32_and_12_16[0], h_s_dadda_pg_rca32_and_11_17[0], h_s_dadda_pg_rca32_and_10_18[0], h_s_dadda_pg_rca32_fa259_xor1, h_s_dadda_pg_rca32_fa259_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_19(a[9], b[19], h_s_dadda_pg_rca32_and_9_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_20(a[8], b[20], h_s_dadda_pg_rca32_and_8_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_21(a[7], b[21], h_s_dadda_pg_rca32_and_7_21);
  fa fa_h_s_dadda_pg_rca32_fa260_out(h_s_dadda_pg_rca32_and_9_19[0], h_s_dadda_pg_rca32_and_8_20[0], h_s_dadda_pg_rca32_and_7_21[0], h_s_dadda_pg_rca32_fa260_xor1, h_s_dadda_pg_rca32_fa260_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_22(a[6], b[22], h_s_dadda_pg_rca32_and_6_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_23(a[5], b[23], h_s_dadda_pg_rca32_and_5_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_24(a[4], b[24], h_s_dadda_pg_rca32_and_4_24);
  fa fa_h_s_dadda_pg_rca32_fa261_out(h_s_dadda_pg_rca32_and_6_22[0], h_s_dadda_pg_rca32_and_5_23[0], h_s_dadda_pg_rca32_and_4_24[0], h_s_dadda_pg_rca32_fa261_xor1, h_s_dadda_pg_rca32_fa261_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_25(a[3], b[25], h_s_dadda_pg_rca32_and_3_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_26(a[2], b[26], h_s_dadda_pg_rca32_and_2_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_27(a[1], b[27], h_s_dadda_pg_rca32_and_1_27);
  fa fa_h_s_dadda_pg_rca32_fa262_out(h_s_dadda_pg_rca32_and_3_25[0], h_s_dadda_pg_rca32_and_2_26[0], h_s_dadda_pg_rca32_and_1_27[0], h_s_dadda_pg_rca32_fa262_xor1, h_s_dadda_pg_rca32_fa262_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_28(a[0], b[28], h_s_dadda_pg_rca32_and_0_28);
  fa fa_h_s_dadda_pg_rca32_fa263_out(h_s_dadda_pg_rca32_and_0_28[0], h_s_dadda_pg_rca32_ha0_xor0[0], h_s_dadda_pg_rca32_fa247_xor1[0], h_s_dadda_pg_rca32_fa263_xor1, h_s_dadda_pg_rca32_fa263_or0);
  fa fa_h_s_dadda_pg_rca32_fa264_out(h_s_dadda_pg_rca32_fa248_xor1[0], h_s_dadda_pg_rca32_fa249_xor1[0], h_s_dadda_pg_rca32_fa250_xor1[0], h_s_dadda_pg_rca32_fa264_xor1, h_s_dadda_pg_rca32_fa264_or0);
  fa fa_h_s_dadda_pg_rca32_fa265_out(h_s_dadda_pg_rca32_fa251_xor1[0], h_s_dadda_pg_rca32_fa252_xor1[0], h_s_dadda_pg_rca32_fa253_xor1[0], h_s_dadda_pg_rca32_fa265_xor1, h_s_dadda_pg_rca32_fa265_or0);
  fa fa_h_s_dadda_pg_rca32_fa266_out(h_s_dadda_pg_rca32_fa254_xor1[0], h_s_dadda_pg_rca32_fa255_xor1[0], h_s_dadda_pg_rca32_fa256_xor1[0], h_s_dadda_pg_rca32_fa266_xor1, h_s_dadda_pg_rca32_fa266_or0);
  fa fa_h_s_dadda_pg_rca32_fa267_out(h_s_dadda_pg_rca32_fa257_xor1[0], h_s_dadda_pg_rca32_fa258_xor1[0], h_s_dadda_pg_rca32_fa259_xor1[0], h_s_dadda_pg_rca32_fa267_xor1, h_s_dadda_pg_rca32_fa267_or0);
  fa fa_h_s_dadda_pg_rca32_fa268_out(h_s_dadda_pg_rca32_fa260_xor1[0], h_s_dadda_pg_rca32_fa261_xor1[0], h_s_dadda_pg_rca32_fa262_xor1[0], h_s_dadda_pg_rca32_fa268_xor1, h_s_dadda_pg_rca32_fa268_or0);
  fa fa_h_s_dadda_pg_rca32_fa269_out(h_s_dadda_pg_rca32_fa268_or0[0], h_s_dadda_pg_rca32_fa267_or0[0], h_s_dadda_pg_rca32_fa266_or0[0], h_s_dadda_pg_rca32_fa269_xor1, h_s_dadda_pg_rca32_fa269_or0);
  fa fa_h_s_dadda_pg_rca32_fa270_out(h_s_dadda_pg_rca32_fa265_or0[0], h_s_dadda_pg_rca32_fa264_or0[0], h_s_dadda_pg_rca32_fa263_or0[0], h_s_dadda_pg_rca32_fa270_xor1, h_s_dadda_pg_rca32_fa270_or0);
  fa fa_h_s_dadda_pg_rca32_fa271_out(h_s_dadda_pg_rca32_fa262_or0[0], h_s_dadda_pg_rca32_fa261_or0[0], h_s_dadda_pg_rca32_fa260_or0[0], h_s_dadda_pg_rca32_fa271_xor1, h_s_dadda_pg_rca32_fa271_or0);
  fa fa_h_s_dadda_pg_rca32_fa272_out(h_s_dadda_pg_rca32_fa259_or0[0], h_s_dadda_pg_rca32_fa258_or0[0], h_s_dadda_pg_rca32_fa257_or0[0], h_s_dadda_pg_rca32_fa272_xor1, h_s_dadda_pg_rca32_fa272_or0);
  fa fa_h_s_dadda_pg_rca32_fa273_out(h_s_dadda_pg_rca32_fa256_or0[0], h_s_dadda_pg_rca32_fa255_or0[0], h_s_dadda_pg_rca32_fa254_or0[0], h_s_dadda_pg_rca32_fa273_xor1, h_s_dadda_pg_rca32_fa273_or0);
  fa fa_h_s_dadda_pg_rca32_fa274_out(h_s_dadda_pg_rca32_fa253_or0[0], h_s_dadda_pg_rca32_fa252_or0[0], h_s_dadda_pg_rca32_fa251_or0[0], h_s_dadda_pg_rca32_fa274_xor1, h_s_dadda_pg_rca32_fa274_or0);
  fa fa_h_s_dadda_pg_rca32_fa275_out(h_s_dadda_pg_rca32_fa250_or0[0], h_s_dadda_pg_rca32_fa249_or0[0], h_s_dadda_pg_rca32_fa248_or0[0], h_s_dadda_pg_rca32_fa275_xor1, h_s_dadda_pg_rca32_fa275_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_4(a[25], b[4], h_s_dadda_pg_rca32_and_25_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_5(a[24], b[5], h_s_dadda_pg_rca32_and_24_5);
  fa fa_h_s_dadda_pg_rca32_fa276_out(h_s_dadda_pg_rca32_fa247_or0[0], h_s_dadda_pg_rca32_and_25_4[0], h_s_dadda_pg_rca32_and_24_5[0], h_s_dadda_pg_rca32_fa276_xor1, h_s_dadda_pg_rca32_fa276_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_6(a[23], b[6], h_s_dadda_pg_rca32_and_23_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_7(a[22], b[7], h_s_dadda_pg_rca32_and_22_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_8(a[21], b[8], h_s_dadda_pg_rca32_and_21_8);
  fa fa_h_s_dadda_pg_rca32_fa277_out(h_s_dadda_pg_rca32_and_23_6[0], h_s_dadda_pg_rca32_and_22_7[0], h_s_dadda_pg_rca32_and_21_8[0], h_s_dadda_pg_rca32_fa277_xor1, h_s_dadda_pg_rca32_fa277_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_9(a[20], b[9], h_s_dadda_pg_rca32_and_20_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_10(a[19], b[10], h_s_dadda_pg_rca32_and_19_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_11(a[18], b[11], h_s_dadda_pg_rca32_and_18_11);
  fa fa_h_s_dadda_pg_rca32_fa278_out(h_s_dadda_pg_rca32_and_20_9[0], h_s_dadda_pg_rca32_and_19_10[0], h_s_dadda_pg_rca32_and_18_11[0], h_s_dadda_pg_rca32_fa278_xor1, h_s_dadda_pg_rca32_fa278_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_12(a[17], b[12], h_s_dadda_pg_rca32_and_17_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_13(a[16], b[13], h_s_dadda_pg_rca32_and_16_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_14(a[15], b[14], h_s_dadda_pg_rca32_and_15_14);
  fa fa_h_s_dadda_pg_rca32_fa279_out(h_s_dadda_pg_rca32_and_17_12[0], h_s_dadda_pg_rca32_and_16_13[0], h_s_dadda_pg_rca32_and_15_14[0], h_s_dadda_pg_rca32_fa279_xor1, h_s_dadda_pg_rca32_fa279_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_15(a[14], b[15], h_s_dadda_pg_rca32_and_14_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_16(a[13], b[16], h_s_dadda_pg_rca32_and_13_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_17(a[12], b[17], h_s_dadda_pg_rca32_and_12_17);
  fa fa_h_s_dadda_pg_rca32_fa280_out(h_s_dadda_pg_rca32_and_14_15[0], h_s_dadda_pg_rca32_and_13_16[0], h_s_dadda_pg_rca32_and_12_17[0], h_s_dadda_pg_rca32_fa280_xor1, h_s_dadda_pg_rca32_fa280_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_18(a[11], b[18], h_s_dadda_pg_rca32_and_11_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_19(a[10], b[19], h_s_dadda_pg_rca32_and_10_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_20(a[9], b[20], h_s_dadda_pg_rca32_and_9_20);
  fa fa_h_s_dadda_pg_rca32_fa281_out(h_s_dadda_pg_rca32_and_11_18[0], h_s_dadda_pg_rca32_and_10_19[0], h_s_dadda_pg_rca32_and_9_20[0], h_s_dadda_pg_rca32_fa281_xor1, h_s_dadda_pg_rca32_fa281_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_21(a[8], b[21], h_s_dadda_pg_rca32_and_8_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_22(a[7], b[22], h_s_dadda_pg_rca32_and_7_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_23(a[6], b[23], h_s_dadda_pg_rca32_and_6_23);
  fa fa_h_s_dadda_pg_rca32_fa282_out(h_s_dadda_pg_rca32_and_8_21[0], h_s_dadda_pg_rca32_and_7_22[0], h_s_dadda_pg_rca32_and_6_23[0], h_s_dadda_pg_rca32_fa282_xor1, h_s_dadda_pg_rca32_fa282_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_24(a[5], b[24], h_s_dadda_pg_rca32_and_5_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_25(a[4], b[25], h_s_dadda_pg_rca32_and_4_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_26(a[3], b[26], h_s_dadda_pg_rca32_and_3_26);
  fa fa_h_s_dadda_pg_rca32_fa283_out(h_s_dadda_pg_rca32_and_5_24[0], h_s_dadda_pg_rca32_and_4_25[0], h_s_dadda_pg_rca32_and_3_26[0], h_s_dadda_pg_rca32_fa283_xor1, h_s_dadda_pg_rca32_fa283_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_27(a[2], b[27], h_s_dadda_pg_rca32_and_2_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_28(a[1], b[28], h_s_dadda_pg_rca32_and_1_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_29(a[0], b[29], h_s_dadda_pg_rca32_and_0_29);
  fa fa_h_s_dadda_pg_rca32_fa284_out(h_s_dadda_pg_rca32_and_2_27[0], h_s_dadda_pg_rca32_and_1_28[0], h_s_dadda_pg_rca32_and_0_29[0], h_s_dadda_pg_rca32_fa284_xor1, h_s_dadda_pg_rca32_fa284_or0);
  fa fa_h_s_dadda_pg_rca32_fa285_out(h_s_dadda_pg_rca32_fa0_xor1[0], h_s_dadda_pg_rca32_ha1_xor0[0], h_s_dadda_pg_rca32_fa269_xor1[0], h_s_dadda_pg_rca32_fa285_xor1, h_s_dadda_pg_rca32_fa285_or0);
  fa fa_h_s_dadda_pg_rca32_fa286_out(h_s_dadda_pg_rca32_fa270_xor1[0], h_s_dadda_pg_rca32_fa271_xor1[0], h_s_dadda_pg_rca32_fa272_xor1[0], h_s_dadda_pg_rca32_fa286_xor1, h_s_dadda_pg_rca32_fa286_or0);
  fa fa_h_s_dadda_pg_rca32_fa287_out(h_s_dadda_pg_rca32_fa273_xor1[0], h_s_dadda_pg_rca32_fa274_xor1[0], h_s_dadda_pg_rca32_fa275_xor1[0], h_s_dadda_pg_rca32_fa287_xor1, h_s_dadda_pg_rca32_fa287_or0);
  fa fa_h_s_dadda_pg_rca32_fa288_out(h_s_dadda_pg_rca32_fa276_xor1[0], h_s_dadda_pg_rca32_fa277_xor1[0], h_s_dadda_pg_rca32_fa278_xor1[0], h_s_dadda_pg_rca32_fa288_xor1, h_s_dadda_pg_rca32_fa288_or0);
  fa fa_h_s_dadda_pg_rca32_fa289_out(h_s_dadda_pg_rca32_fa279_xor1[0], h_s_dadda_pg_rca32_fa280_xor1[0], h_s_dadda_pg_rca32_fa281_xor1[0], h_s_dadda_pg_rca32_fa289_xor1, h_s_dadda_pg_rca32_fa289_or0);
  fa fa_h_s_dadda_pg_rca32_fa290_out(h_s_dadda_pg_rca32_fa282_xor1[0], h_s_dadda_pg_rca32_fa283_xor1[0], h_s_dadda_pg_rca32_fa284_xor1[0], h_s_dadda_pg_rca32_fa290_xor1, h_s_dadda_pg_rca32_fa290_or0);
  fa fa_h_s_dadda_pg_rca32_fa291_out(h_s_dadda_pg_rca32_fa290_or0[0], h_s_dadda_pg_rca32_fa289_or0[0], h_s_dadda_pg_rca32_fa288_or0[0], h_s_dadda_pg_rca32_fa291_xor1, h_s_dadda_pg_rca32_fa291_or0);
  fa fa_h_s_dadda_pg_rca32_fa292_out(h_s_dadda_pg_rca32_fa287_or0[0], h_s_dadda_pg_rca32_fa286_or0[0], h_s_dadda_pg_rca32_fa285_or0[0], h_s_dadda_pg_rca32_fa292_xor1, h_s_dadda_pg_rca32_fa292_or0);
  fa fa_h_s_dadda_pg_rca32_fa293_out(h_s_dadda_pg_rca32_fa284_or0[0], h_s_dadda_pg_rca32_fa283_or0[0], h_s_dadda_pg_rca32_fa282_or0[0], h_s_dadda_pg_rca32_fa293_xor1, h_s_dadda_pg_rca32_fa293_or0);
  fa fa_h_s_dadda_pg_rca32_fa294_out(h_s_dadda_pg_rca32_fa281_or0[0], h_s_dadda_pg_rca32_fa280_or0[0], h_s_dadda_pg_rca32_fa279_or0[0], h_s_dadda_pg_rca32_fa294_xor1, h_s_dadda_pg_rca32_fa294_or0);
  fa fa_h_s_dadda_pg_rca32_fa295_out(h_s_dadda_pg_rca32_fa278_or0[0], h_s_dadda_pg_rca32_fa277_or0[0], h_s_dadda_pg_rca32_fa276_or0[0], h_s_dadda_pg_rca32_fa295_xor1, h_s_dadda_pg_rca32_fa295_or0);
  fa fa_h_s_dadda_pg_rca32_fa296_out(h_s_dadda_pg_rca32_fa275_or0[0], h_s_dadda_pg_rca32_fa274_or0[0], h_s_dadda_pg_rca32_fa273_or0[0], h_s_dadda_pg_rca32_fa296_xor1, h_s_dadda_pg_rca32_fa296_or0);
  fa fa_h_s_dadda_pg_rca32_fa297_out(h_s_dadda_pg_rca32_fa272_or0[0], h_s_dadda_pg_rca32_fa271_or0[0], h_s_dadda_pg_rca32_fa270_or0[0], h_s_dadda_pg_rca32_fa297_xor1, h_s_dadda_pg_rca32_fa297_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_6(a[24], b[6], h_s_dadda_pg_rca32_and_24_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_7(a[23], b[7], h_s_dadda_pg_rca32_and_23_7);
  fa fa_h_s_dadda_pg_rca32_fa298_out(h_s_dadda_pg_rca32_fa269_or0[0], h_s_dadda_pg_rca32_and_24_6[0], h_s_dadda_pg_rca32_and_23_7[0], h_s_dadda_pg_rca32_fa298_xor1, h_s_dadda_pg_rca32_fa298_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_8(a[22], b[8], h_s_dadda_pg_rca32_and_22_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_9(a[21], b[9], h_s_dadda_pg_rca32_and_21_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_10(a[20], b[10], h_s_dadda_pg_rca32_and_20_10);
  fa fa_h_s_dadda_pg_rca32_fa299_out(h_s_dadda_pg_rca32_and_22_8[0], h_s_dadda_pg_rca32_and_21_9[0], h_s_dadda_pg_rca32_and_20_10[0], h_s_dadda_pg_rca32_fa299_xor1, h_s_dadda_pg_rca32_fa299_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_11(a[19], b[11], h_s_dadda_pg_rca32_and_19_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_12(a[18], b[12], h_s_dadda_pg_rca32_and_18_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_13(a[17], b[13], h_s_dadda_pg_rca32_and_17_13);
  fa fa_h_s_dadda_pg_rca32_fa300_out(h_s_dadda_pg_rca32_and_19_11[0], h_s_dadda_pg_rca32_and_18_12[0], h_s_dadda_pg_rca32_and_17_13[0], h_s_dadda_pg_rca32_fa300_xor1, h_s_dadda_pg_rca32_fa300_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_14(a[16], b[14], h_s_dadda_pg_rca32_and_16_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_15(a[15], b[15], h_s_dadda_pg_rca32_and_15_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_16(a[14], b[16], h_s_dadda_pg_rca32_and_14_16);
  fa fa_h_s_dadda_pg_rca32_fa301_out(h_s_dadda_pg_rca32_and_16_14[0], h_s_dadda_pg_rca32_and_15_15[0], h_s_dadda_pg_rca32_and_14_16[0], h_s_dadda_pg_rca32_fa301_xor1, h_s_dadda_pg_rca32_fa301_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_17(a[13], b[17], h_s_dadda_pg_rca32_and_13_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_18(a[12], b[18], h_s_dadda_pg_rca32_and_12_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_19(a[11], b[19], h_s_dadda_pg_rca32_and_11_19);
  fa fa_h_s_dadda_pg_rca32_fa302_out(h_s_dadda_pg_rca32_and_13_17[0], h_s_dadda_pg_rca32_and_12_18[0], h_s_dadda_pg_rca32_and_11_19[0], h_s_dadda_pg_rca32_fa302_xor1, h_s_dadda_pg_rca32_fa302_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_20(a[10], b[20], h_s_dadda_pg_rca32_and_10_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_21(a[9], b[21], h_s_dadda_pg_rca32_and_9_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_22(a[8], b[22], h_s_dadda_pg_rca32_and_8_22);
  fa fa_h_s_dadda_pg_rca32_fa303_out(h_s_dadda_pg_rca32_and_10_20[0], h_s_dadda_pg_rca32_and_9_21[0], h_s_dadda_pg_rca32_and_8_22[0], h_s_dadda_pg_rca32_fa303_xor1, h_s_dadda_pg_rca32_fa303_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_23(a[7], b[23], h_s_dadda_pg_rca32_and_7_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_24(a[6], b[24], h_s_dadda_pg_rca32_and_6_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_25(a[5], b[25], h_s_dadda_pg_rca32_and_5_25);
  fa fa_h_s_dadda_pg_rca32_fa304_out(h_s_dadda_pg_rca32_and_7_23[0], h_s_dadda_pg_rca32_and_6_24[0], h_s_dadda_pg_rca32_and_5_25[0], h_s_dadda_pg_rca32_fa304_xor1, h_s_dadda_pg_rca32_fa304_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_26(a[4], b[26], h_s_dadda_pg_rca32_and_4_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_27(a[3], b[27], h_s_dadda_pg_rca32_and_3_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_28(a[2], b[28], h_s_dadda_pg_rca32_and_2_28);
  fa fa_h_s_dadda_pg_rca32_fa305_out(h_s_dadda_pg_rca32_and_4_26[0], h_s_dadda_pg_rca32_and_3_27[0], h_s_dadda_pg_rca32_and_2_28[0], h_s_dadda_pg_rca32_fa305_xor1, h_s_dadda_pg_rca32_fa305_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_29(a[1], b[29], h_s_dadda_pg_rca32_and_1_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_30(a[0], b[30], h_s_dadda_pg_rca32_and_0_30);
  fa fa_h_s_dadda_pg_rca32_fa306_out(h_s_dadda_pg_rca32_and_1_29[0], h_s_dadda_pg_rca32_and_0_30[0], h_s_dadda_pg_rca32_fa1_xor1[0], h_s_dadda_pg_rca32_fa306_xor1, h_s_dadda_pg_rca32_fa306_or0);
  fa fa_h_s_dadda_pg_rca32_fa307_out(h_s_dadda_pg_rca32_fa2_xor1[0], h_s_dadda_pg_rca32_ha2_xor0[0], h_s_dadda_pg_rca32_fa291_xor1[0], h_s_dadda_pg_rca32_fa307_xor1, h_s_dadda_pg_rca32_fa307_or0);
  fa fa_h_s_dadda_pg_rca32_fa308_out(h_s_dadda_pg_rca32_fa292_xor1[0], h_s_dadda_pg_rca32_fa293_xor1[0], h_s_dadda_pg_rca32_fa294_xor1[0], h_s_dadda_pg_rca32_fa308_xor1, h_s_dadda_pg_rca32_fa308_or0);
  fa fa_h_s_dadda_pg_rca32_fa309_out(h_s_dadda_pg_rca32_fa295_xor1[0], h_s_dadda_pg_rca32_fa296_xor1[0], h_s_dadda_pg_rca32_fa297_xor1[0], h_s_dadda_pg_rca32_fa309_xor1, h_s_dadda_pg_rca32_fa309_or0);
  fa fa_h_s_dadda_pg_rca32_fa310_out(h_s_dadda_pg_rca32_fa298_xor1[0], h_s_dadda_pg_rca32_fa299_xor1[0], h_s_dadda_pg_rca32_fa300_xor1[0], h_s_dadda_pg_rca32_fa310_xor1, h_s_dadda_pg_rca32_fa310_or0);
  fa fa_h_s_dadda_pg_rca32_fa311_out(h_s_dadda_pg_rca32_fa301_xor1[0], h_s_dadda_pg_rca32_fa302_xor1[0], h_s_dadda_pg_rca32_fa303_xor1[0], h_s_dadda_pg_rca32_fa311_xor1, h_s_dadda_pg_rca32_fa311_or0);
  fa fa_h_s_dadda_pg_rca32_fa312_out(h_s_dadda_pg_rca32_fa304_xor1[0], h_s_dadda_pg_rca32_fa305_xor1[0], h_s_dadda_pg_rca32_fa306_xor1[0], h_s_dadda_pg_rca32_fa312_xor1, h_s_dadda_pg_rca32_fa312_or0);
  fa fa_h_s_dadda_pg_rca32_fa313_out(h_s_dadda_pg_rca32_fa312_or0[0], h_s_dadda_pg_rca32_fa311_or0[0], h_s_dadda_pg_rca32_fa310_or0[0], h_s_dadda_pg_rca32_fa313_xor1, h_s_dadda_pg_rca32_fa313_or0);
  fa fa_h_s_dadda_pg_rca32_fa314_out(h_s_dadda_pg_rca32_fa309_or0[0], h_s_dadda_pg_rca32_fa308_or0[0], h_s_dadda_pg_rca32_fa307_or0[0], h_s_dadda_pg_rca32_fa314_xor1, h_s_dadda_pg_rca32_fa314_or0);
  fa fa_h_s_dadda_pg_rca32_fa315_out(h_s_dadda_pg_rca32_fa306_or0[0], h_s_dadda_pg_rca32_fa305_or0[0], h_s_dadda_pg_rca32_fa304_or0[0], h_s_dadda_pg_rca32_fa315_xor1, h_s_dadda_pg_rca32_fa315_or0);
  fa fa_h_s_dadda_pg_rca32_fa316_out(h_s_dadda_pg_rca32_fa303_or0[0], h_s_dadda_pg_rca32_fa302_or0[0], h_s_dadda_pg_rca32_fa301_or0[0], h_s_dadda_pg_rca32_fa316_xor1, h_s_dadda_pg_rca32_fa316_or0);
  fa fa_h_s_dadda_pg_rca32_fa317_out(h_s_dadda_pg_rca32_fa300_or0[0], h_s_dadda_pg_rca32_fa299_or0[0], h_s_dadda_pg_rca32_fa298_or0[0], h_s_dadda_pg_rca32_fa317_xor1, h_s_dadda_pg_rca32_fa317_or0);
  fa fa_h_s_dadda_pg_rca32_fa318_out(h_s_dadda_pg_rca32_fa297_or0[0], h_s_dadda_pg_rca32_fa296_or0[0], h_s_dadda_pg_rca32_fa295_or0[0], h_s_dadda_pg_rca32_fa318_xor1, h_s_dadda_pg_rca32_fa318_or0);
  fa fa_h_s_dadda_pg_rca32_fa319_out(h_s_dadda_pg_rca32_fa294_or0[0], h_s_dadda_pg_rca32_fa293_or0[0], h_s_dadda_pg_rca32_fa292_or0[0], h_s_dadda_pg_rca32_fa319_xor1, h_s_dadda_pg_rca32_fa319_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_8(a[23], b[8], h_s_dadda_pg_rca32_and_23_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_9(a[22], b[9], h_s_dadda_pg_rca32_and_22_9);
  fa fa_h_s_dadda_pg_rca32_fa320_out(h_s_dadda_pg_rca32_fa291_or0[0], h_s_dadda_pg_rca32_and_23_8[0], h_s_dadda_pg_rca32_and_22_9[0], h_s_dadda_pg_rca32_fa320_xor1, h_s_dadda_pg_rca32_fa320_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_10(a[21], b[10], h_s_dadda_pg_rca32_and_21_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_11(a[20], b[11], h_s_dadda_pg_rca32_and_20_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_12(a[19], b[12], h_s_dadda_pg_rca32_and_19_12);
  fa fa_h_s_dadda_pg_rca32_fa321_out(h_s_dadda_pg_rca32_and_21_10[0], h_s_dadda_pg_rca32_and_20_11[0], h_s_dadda_pg_rca32_and_19_12[0], h_s_dadda_pg_rca32_fa321_xor1, h_s_dadda_pg_rca32_fa321_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_13(a[18], b[13], h_s_dadda_pg_rca32_and_18_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_14(a[17], b[14], h_s_dadda_pg_rca32_and_17_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_15(a[16], b[15], h_s_dadda_pg_rca32_and_16_15);
  fa fa_h_s_dadda_pg_rca32_fa322_out(h_s_dadda_pg_rca32_and_18_13[0], h_s_dadda_pg_rca32_and_17_14[0], h_s_dadda_pg_rca32_and_16_15[0], h_s_dadda_pg_rca32_fa322_xor1, h_s_dadda_pg_rca32_fa322_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_16(a[15], b[16], h_s_dadda_pg_rca32_and_15_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_17(a[14], b[17], h_s_dadda_pg_rca32_and_14_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_18(a[13], b[18], h_s_dadda_pg_rca32_and_13_18);
  fa fa_h_s_dadda_pg_rca32_fa323_out(h_s_dadda_pg_rca32_and_15_16[0], h_s_dadda_pg_rca32_and_14_17[0], h_s_dadda_pg_rca32_and_13_18[0], h_s_dadda_pg_rca32_fa323_xor1, h_s_dadda_pg_rca32_fa323_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_19(a[12], b[19], h_s_dadda_pg_rca32_and_12_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_20(a[11], b[20], h_s_dadda_pg_rca32_and_11_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_21(a[10], b[21], h_s_dadda_pg_rca32_and_10_21);
  fa fa_h_s_dadda_pg_rca32_fa324_out(h_s_dadda_pg_rca32_and_12_19[0], h_s_dadda_pg_rca32_and_11_20[0], h_s_dadda_pg_rca32_and_10_21[0], h_s_dadda_pg_rca32_fa324_xor1, h_s_dadda_pg_rca32_fa324_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_22(a[9], b[22], h_s_dadda_pg_rca32_and_9_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_23(a[8], b[23], h_s_dadda_pg_rca32_and_8_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_24(a[7], b[24], h_s_dadda_pg_rca32_and_7_24);
  fa fa_h_s_dadda_pg_rca32_fa325_out(h_s_dadda_pg_rca32_and_9_22[0], h_s_dadda_pg_rca32_and_8_23[0], h_s_dadda_pg_rca32_and_7_24[0], h_s_dadda_pg_rca32_fa325_xor1, h_s_dadda_pg_rca32_fa325_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_25(a[6], b[25], h_s_dadda_pg_rca32_and_6_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_26(a[5], b[26], h_s_dadda_pg_rca32_and_5_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_27(a[4], b[27], h_s_dadda_pg_rca32_and_4_27);
  fa fa_h_s_dadda_pg_rca32_fa326_out(h_s_dadda_pg_rca32_and_6_25[0], h_s_dadda_pg_rca32_and_5_26[0], h_s_dadda_pg_rca32_and_4_27[0], h_s_dadda_pg_rca32_fa326_xor1, h_s_dadda_pg_rca32_fa326_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_28(a[3], b[28], h_s_dadda_pg_rca32_and_3_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_29(a[2], b[29], h_s_dadda_pg_rca32_and_2_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_30(a[1], b[30], h_s_dadda_pg_rca32_and_1_30);
  fa fa_h_s_dadda_pg_rca32_fa327_out(h_s_dadda_pg_rca32_and_3_28[0], h_s_dadda_pg_rca32_and_2_29[0], h_s_dadda_pg_rca32_and_1_30[0], h_s_dadda_pg_rca32_fa327_xor1, h_s_dadda_pg_rca32_fa327_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_0_31(a[0], b[31], h_s_dadda_pg_rca32_nand_0_31);
  fa fa_h_s_dadda_pg_rca32_fa328_out(h_s_dadda_pg_rca32_nand_0_31[0], h_s_dadda_pg_rca32_fa3_xor1[0], h_s_dadda_pg_rca32_fa4_xor1[0], h_s_dadda_pg_rca32_fa328_xor1, h_s_dadda_pg_rca32_fa328_or0);
  fa fa_h_s_dadda_pg_rca32_fa329_out(h_s_dadda_pg_rca32_fa5_xor1[0], h_s_dadda_pg_rca32_ha3_xor0[0], h_s_dadda_pg_rca32_fa313_xor1[0], h_s_dadda_pg_rca32_fa329_xor1, h_s_dadda_pg_rca32_fa329_or0);
  fa fa_h_s_dadda_pg_rca32_fa330_out(h_s_dadda_pg_rca32_fa314_xor1[0], h_s_dadda_pg_rca32_fa315_xor1[0], h_s_dadda_pg_rca32_fa316_xor1[0], h_s_dadda_pg_rca32_fa330_xor1, h_s_dadda_pg_rca32_fa330_or0);
  fa fa_h_s_dadda_pg_rca32_fa331_out(h_s_dadda_pg_rca32_fa317_xor1[0], h_s_dadda_pg_rca32_fa318_xor1[0], h_s_dadda_pg_rca32_fa319_xor1[0], h_s_dadda_pg_rca32_fa331_xor1, h_s_dadda_pg_rca32_fa331_or0);
  fa fa_h_s_dadda_pg_rca32_fa332_out(h_s_dadda_pg_rca32_fa320_xor1[0], h_s_dadda_pg_rca32_fa321_xor1[0], h_s_dadda_pg_rca32_fa322_xor1[0], h_s_dadda_pg_rca32_fa332_xor1, h_s_dadda_pg_rca32_fa332_or0);
  fa fa_h_s_dadda_pg_rca32_fa333_out(h_s_dadda_pg_rca32_fa323_xor1[0], h_s_dadda_pg_rca32_fa324_xor1[0], h_s_dadda_pg_rca32_fa325_xor1[0], h_s_dadda_pg_rca32_fa333_xor1, h_s_dadda_pg_rca32_fa333_or0);
  fa fa_h_s_dadda_pg_rca32_fa334_out(h_s_dadda_pg_rca32_fa326_xor1[0], h_s_dadda_pg_rca32_fa327_xor1[0], h_s_dadda_pg_rca32_fa328_xor1[0], h_s_dadda_pg_rca32_fa334_xor1, h_s_dadda_pg_rca32_fa334_or0);
  fa fa_h_s_dadda_pg_rca32_fa335_out(h_s_dadda_pg_rca32_fa334_or0[0], h_s_dadda_pg_rca32_fa333_or0[0], h_s_dadda_pg_rca32_fa332_or0[0], h_s_dadda_pg_rca32_fa335_xor1, h_s_dadda_pg_rca32_fa335_or0);
  fa fa_h_s_dadda_pg_rca32_fa336_out(h_s_dadda_pg_rca32_fa331_or0[0], h_s_dadda_pg_rca32_fa330_or0[0], h_s_dadda_pg_rca32_fa329_or0[0], h_s_dadda_pg_rca32_fa336_xor1, h_s_dadda_pg_rca32_fa336_or0);
  fa fa_h_s_dadda_pg_rca32_fa337_out(h_s_dadda_pg_rca32_fa328_or0[0], h_s_dadda_pg_rca32_fa327_or0[0], h_s_dadda_pg_rca32_fa326_or0[0], h_s_dadda_pg_rca32_fa337_xor1, h_s_dadda_pg_rca32_fa337_or0);
  fa fa_h_s_dadda_pg_rca32_fa338_out(h_s_dadda_pg_rca32_fa325_or0[0], h_s_dadda_pg_rca32_fa324_or0[0], h_s_dadda_pg_rca32_fa323_or0[0], h_s_dadda_pg_rca32_fa338_xor1, h_s_dadda_pg_rca32_fa338_or0);
  fa fa_h_s_dadda_pg_rca32_fa339_out(h_s_dadda_pg_rca32_fa322_or0[0], h_s_dadda_pg_rca32_fa321_or0[0], h_s_dadda_pg_rca32_fa320_or0[0], h_s_dadda_pg_rca32_fa339_xor1, h_s_dadda_pg_rca32_fa339_or0);
  fa fa_h_s_dadda_pg_rca32_fa340_out(h_s_dadda_pg_rca32_fa319_or0[0], h_s_dadda_pg_rca32_fa318_or0[0], h_s_dadda_pg_rca32_fa317_or0[0], h_s_dadda_pg_rca32_fa340_xor1, h_s_dadda_pg_rca32_fa340_or0);
  fa fa_h_s_dadda_pg_rca32_fa341_out(h_s_dadda_pg_rca32_fa316_or0[0], h_s_dadda_pg_rca32_fa315_or0[0], h_s_dadda_pg_rca32_fa314_or0[0], h_s_dadda_pg_rca32_fa341_xor1, h_s_dadda_pg_rca32_fa341_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_8(a[24], b[8], h_s_dadda_pg_rca32_and_24_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_9(a[23], b[9], h_s_dadda_pg_rca32_and_23_9);
  fa fa_h_s_dadda_pg_rca32_fa342_out(h_s_dadda_pg_rca32_fa313_or0[0], h_s_dadda_pg_rca32_and_24_8[0], h_s_dadda_pg_rca32_and_23_9[0], h_s_dadda_pg_rca32_fa342_xor1, h_s_dadda_pg_rca32_fa342_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_10(a[22], b[10], h_s_dadda_pg_rca32_and_22_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_11(a[21], b[11], h_s_dadda_pg_rca32_and_21_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_12(a[20], b[12], h_s_dadda_pg_rca32_and_20_12);
  fa fa_h_s_dadda_pg_rca32_fa343_out(h_s_dadda_pg_rca32_and_22_10[0], h_s_dadda_pg_rca32_and_21_11[0], h_s_dadda_pg_rca32_and_20_12[0], h_s_dadda_pg_rca32_fa343_xor1, h_s_dadda_pg_rca32_fa343_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_13(a[19], b[13], h_s_dadda_pg_rca32_and_19_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_14(a[18], b[14], h_s_dadda_pg_rca32_and_18_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_15(a[17], b[15], h_s_dadda_pg_rca32_and_17_15);
  fa fa_h_s_dadda_pg_rca32_fa344_out(h_s_dadda_pg_rca32_and_19_13[0], h_s_dadda_pg_rca32_and_18_14[0], h_s_dadda_pg_rca32_and_17_15[0], h_s_dadda_pg_rca32_fa344_xor1, h_s_dadda_pg_rca32_fa344_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_16(a[16], b[16], h_s_dadda_pg_rca32_and_16_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_17(a[15], b[17], h_s_dadda_pg_rca32_and_15_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_18(a[14], b[18], h_s_dadda_pg_rca32_and_14_18);
  fa fa_h_s_dadda_pg_rca32_fa345_out(h_s_dadda_pg_rca32_and_16_16[0], h_s_dadda_pg_rca32_and_15_17[0], h_s_dadda_pg_rca32_and_14_18[0], h_s_dadda_pg_rca32_fa345_xor1, h_s_dadda_pg_rca32_fa345_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_19(a[13], b[19], h_s_dadda_pg_rca32_and_13_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_20(a[12], b[20], h_s_dadda_pg_rca32_and_12_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_21(a[11], b[21], h_s_dadda_pg_rca32_and_11_21);
  fa fa_h_s_dadda_pg_rca32_fa346_out(h_s_dadda_pg_rca32_and_13_19[0], h_s_dadda_pg_rca32_and_12_20[0], h_s_dadda_pg_rca32_and_11_21[0], h_s_dadda_pg_rca32_fa346_xor1, h_s_dadda_pg_rca32_fa346_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_22(a[10], b[22], h_s_dadda_pg_rca32_and_10_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_23(a[9], b[23], h_s_dadda_pg_rca32_and_9_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_24(a[8], b[24], h_s_dadda_pg_rca32_and_8_24);
  fa fa_h_s_dadda_pg_rca32_fa347_out(h_s_dadda_pg_rca32_and_10_22[0], h_s_dadda_pg_rca32_and_9_23[0], h_s_dadda_pg_rca32_and_8_24[0], h_s_dadda_pg_rca32_fa347_xor1, h_s_dadda_pg_rca32_fa347_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_25(a[7], b[25], h_s_dadda_pg_rca32_and_7_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_26(a[6], b[26], h_s_dadda_pg_rca32_and_6_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_27(a[5], b[27], h_s_dadda_pg_rca32_and_5_27);
  fa fa_h_s_dadda_pg_rca32_fa348_out(h_s_dadda_pg_rca32_and_7_25[0], h_s_dadda_pg_rca32_and_6_26[0], h_s_dadda_pg_rca32_and_5_27[0], h_s_dadda_pg_rca32_fa348_xor1, h_s_dadda_pg_rca32_fa348_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_28(a[4], b[28], h_s_dadda_pg_rca32_and_4_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_29(a[3], b[29], h_s_dadda_pg_rca32_and_3_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_30(a[2], b[30], h_s_dadda_pg_rca32_and_2_30);
  fa fa_h_s_dadda_pg_rca32_fa349_out(h_s_dadda_pg_rca32_and_4_28[0], h_s_dadda_pg_rca32_and_3_29[0], h_s_dadda_pg_rca32_and_2_30[0], h_s_dadda_pg_rca32_fa349_xor1, h_s_dadda_pg_rca32_fa349_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_1_31(a[1], b[31], h_s_dadda_pg_rca32_nand_1_31);
  fa fa_h_s_dadda_pg_rca32_fa350_out(h_s_dadda_pg_rca32_nand_1_31[0], h_s_dadda_pg_rca32_fa6_xor1[0], h_s_dadda_pg_rca32_fa7_xor1[0], h_s_dadda_pg_rca32_fa350_xor1, h_s_dadda_pg_rca32_fa350_or0);
  fa fa_h_s_dadda_pg_rca32_fa351_out(h_s_dadda_pg_rca32_fa8_xor1[0], h_s_dadda_pg_rca32_fa9_xor1[0], h_s_dadda_pg_rca32_fa335_xor1[0], h_s_dadda_pg_rca32_fa351_xor1, h_s_dadda_pg_rca32_fa351_or0);
  fa fa_h_s_dadda_pg_rca32_fa352_out(h_s_dadda_pg_rca32_fa336_xor1[0], h_s_dadda_pg_rca32_fa337_xor1[0], h_s_dadda_pg_rca32_fa338_xor1[0], h_s_dadda_pg_rca32_fa352_xor1, h_s_dadda_pg_rca32_fa352_or0);
  fa fa_h_s_dadda_pg_rca32_fa353_out(h_s_dadda_pg_rca32_fa339_xor1[0], h_s_dadda_pg_rca32_fa340_xor1[0], h_s_dadda_pg_rca32_fa341_xor1[0], h_s_dadda_pg_rca32_fa353_xor1, h_s_dadda_pg_rca32_fa353_or0);
  fa fa_h_s_dadda_pg_rca32_fa354_out(h_s_dadda_pg_rca32_fa342_xor1[0], h_s_dadda_pg_rca32_fa343_xor1[0], h_s_dadda_pg_rca32_fa344_xor1[0], h_s_dadda_pg_rca32_fa354_xor1, h_s_dadda_pg_rca32_fa354_or0);
  fa fa_h_s_dadda_pg_rca32_fa355_out(h_s_dadda_pg_rca32_fa345_xor1[0], h_s_dadda_pg_rca32_fa346_xor1[0], h_s_dadda_pg_rca32_fa347_xor1[0], h_s_dadda_pg_rca32_fa355_xor1, h_s_dadda_pg_rca32_fa355_or0);
  fa fa_h_s_dadda_pg_rca32_fa356_out(h_s_dadda_pg_rca32_fa348_xor1[0], h_s_dadda_pg_rca32_fa349_xor1[0], h_s_dadda_pg_rca32_fa350_xor1[0], h_s_dadda_pg_rca32_fa356_xor1, h_s_dadda_pg_rca32_fa356_or0);
  fa fa_h_s_dadda_pg_rca32_fa357_out(h_s_dadda_pg_rca32_fa356_or0[0], h_s_dadda_pg_rca32_fa355_or0[0], h_s_dadda_pg_rca32_fa354_or0[0], h_s_dadda_pg_rca32_fa357_xor1, h_s_dadda_pg_rca32_fa357_or0);
  fa fa_h_s_dadda_pg_rca32_fa358_out(h_s_dadda_pg_rca32_fa353_or0[0], h_s_dadda_pg_rca32_fa352_or0[0], h_s_dadda_pg_rca32_fa351_or0[0], h_s_dadda_pg_rca32_fa358_xor1, h_s_dadda_pg_rca32_fa358_or0);
  fa fa_h_s_dadda_pg_rca32_fa359_out(h_s_dadda_pg_rca32_fa350_or0[0], h_s_dadda_pg_rca32_fa349_or0[0], h_s_dadda_pg_rca32_fa348_or0[0], h_s_dadda_pg_rca32_fa359_xor1, h_s_dadda_pg_rca32_fa359_or0);
  fa fa_h_s_dadda_pg_rca32_fa360_out(h_s_dadda_pg_rca32_fa347_or0[0], h_s_dadda_pg_rca32_fa346_or0[0], h_s_dadda_pg_rca32_fa345_or0[0], h_s_dadda_pg_rca32_fa360_xor1, h_s_dadda_pg_rca32_fa360_or0);
  fa fa_h_s_dadda_pg_rca32_fa361_out(h_s_dadda_pg_rca32_fa344_or0[0], h_s_dadda_pg_rca32_fa343_or0[0], h_s_dadda_pg_rca32_fa342_or0[0], h_s_dadda_pg_rca32_fa361_xor1, h_s_dadda_pg_rca32_fa361_or0);
  fa fa_h_s_dadda_pg_rca32_fa362_out(h_s_dadda_pg_rca32_fa341_or0[0], h_s_dadda_pg_rca32_fa340_or0[0], h_s_dadda_pg_rca32_fa339_or0[0], h_s_dadda_pg_rca32_fa362_xor1, h_s_dadda_pg_rca32_fa362_or0);
  fa fa_h_s_dadda_pg_rca32_fa363_out(h_s_dadda_pg_rca32_fa338_or0[0], h_s_dadda_pg_rca32_fa337_or0[0], h_s_dadda_pg_rca32_fa336_or0[0], h_s_dadda_pg_rca32_fa363_xor1, h_s_dadda_pg_rca32_fa363_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_7(a[26], b[7], h_s_dadda_pg_rca32_and_26_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_8(a[25], b[8], h_s_dadda_pg_rca32_and_25_8);
  fa fa_h_s_dadda_pg_rca32_fa364_out(h_s_dadda_pg_rca32_fa335_or0[0], h_s_dadda_pg_rca32_and_26_7[0], h_s_dadda_pg_rca32_and_25_8[0], h_s_dadda_pg_rca32_fa364_xor1, h_s_dadda_pg_rca32_fa364_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_9(a[24], b[9], h_s_dadda_pg_rca32_and_24_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_10(a[23], b[10], h_s_dadda_pg_rca32_and_23_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_11(a[22], b[11], h_s_dadda_pg_rca32_and_22_11);
  fa fa_h_s_dadda_pg_rca32_fa365_out(h_s_dadda_pg_rca32_and_24_9[0], h_s_dadda_pg_rca32_and_23_10[0], h_s_dadda_pg_rca32_and_22_11[0], h_s_dadda_pg_rca32_fa365_xor1, h_s_dadda_pg_rca32_fa365_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_12(a[21], b[12], h_s_dadda_pg_rca32_and_21_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_13(a[20], b[13], h_s_dadda_pg_rca32_and_20_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_14(a[19], b[14], h_s_dadda_pg_rca32_and_19_14);
  fa fa_h_s_dadda_pg_rca32_fa366_out(h_s_dadda_pg_rca32_and_21_12[0], h_s_dadda_pg_rca32_and_20_13[0], h_s_dadda_pg_rca32_and_19_14[0], h_s_dadda_pg_rca32_fa366_xor1, h_s_dadda_pg_rca32_fa366_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_15(a[18], b[15], h_s_dadda_pg_rca32_and_18_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_16(a[17], b[16], h_s_dadda_pg_rca32_and_17_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_17(a[16], b[17], h_s_dadda_pg_rca32_and_16_17);
  fa fa_h_s_dadda_pg_rca32_fa367_out(h_s_dadda_pg_rca32_and_18_15[0], h_s_dadda_pg_rca32_and_17_16[0], h_s_dadda_pg_rca32_and_16_17[0], h_s_dadda_pg_rca32_fa367_xor1, h_s_dadda_pg_rca32_fa367_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_18(a[15], b[18], h_s_dadda_pg_rca32_and_15_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_19(a[14], b[19], h_s_dadda_pg_rca32_and_14_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_20(a[13], b[20], h_s_dadda_pg_rca32_and_13_20);
  fa fa_h_s_dadda_pg_rca32_fa368_out(h_s_dadda_pg_rca32_and_15_18[0], h_s_dadda_pg_rca32_and_14_19[0], h_s_dadda_pg_rca32_and_13_20[0], h_s_dadda_pg_rca32_fa368_xor1, h_s_dadda_pg_rca32_fa368_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_21(a[12], b[21], h_s_dadda_pg_rca32_and_12_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_22(a[11], b[22], h_s_dadda_pg_rca32_and_11_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_23(a[10], b[23], h_s_dadda_pg_rca32_and_10_23);
  fa fa_h_s_dadda_pg_rca32_fa369_out(h_s_dadda_pg_rca32_and_12_21[0], h_s_dadda_pg_rca32_and_11_22[0], h_s_dadda_pg_rca32_and_10_23[0], h_s_dadda_pg_rca32_fa369_xor1, h_s_dadda_pg_rca32_fa369_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_24(a[9], b[24], h_s_dadda_pg_rca32_and_9_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_25(a[8], b[25], h_s_dadda_pg_rca32_and_8_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_26(a[7], b[26], h_s_dadda_pg_rca32_and_7_26);
  fa fa_h_s_dadda_pg_rca32_fa370_out(h_s_dadda_pg_rca32_and_9_24[0], h_s_dadda_pg_rca32_and_8_25[0], h_s_dadda_pg_rca32_and_7_26[0], h_s_dadda_pg_rca32_fa370_xor1, h_s_dadda_pg_rca32_fa370_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_27(a[6], b[27], h_s_dadda_pg_rca32_and_6_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_28(a[5], b[28], h_s_dadda_pg_rca32_and_5_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_29(a[4], b[29], h_s_dadda_pg_rca32_and_4_29);
  fa fa_h_s_dadda_pg_rca32_fa371_out(h_s_dadda_pg_rca32_and_6_27[0], h_s_dadda_pg_rca32_and_5_28[0], h_s_dadda_pg_rca32_and_4_29[0], h_s_dadda_pg_rca32_fa371_xor1, h_s_dadda_pg_rca32_fa371_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_30(a[3], b[30], h_s_dadda_pg_rca32_and_3_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_2_31(a[2], b[31], h_s_dadda_pg_rca32_nand_2_31);
  fa fa_h_s_dadda_pg_rca32_fa372_out(h_s_dadda_pg_rca32_and_3_30[0], h_s_dadda_pg_rca32_nand_2_31[0], h_s_dadda_pg_rca32_fa10_xor1[0], h_s_dadda_pg_rca32_fa372_xor1, h_s_dadda_pg_rca32_fa372_or0);
  fa fa_h_s_dadda_pg_rca32_fa373_out(h_s_dadda_pg_rca32_fa11_xor1[0], h_s_dadda_pg_rca32_fa12_xor1[0], h_s_dadda_pg_rca32_fa357_xor1[0], h_s_dadda_pg_rca32_fa373_xor1, h_s_dadda_pg_rca32_fa373_or0);
  fa fa_h_s_dadda_pg_rca32_fa374_out(h_s_dadda_pg_rca32_fa358_xor1[0], h_s_dadda_pg_rca32_fa359_xor1[0], h_s_dadda_pg_rca32_fa360_xor1[0], h_s_dadda_pg_rca32_fa374_xor1, h_s_dadda_pg_rca32_fa374_or0);
  fa fa_h_s_dadda_pg_rca32_fa375_out(h_s_dadda_pg_rca32_fa361_xor1[0], h_s_dadda_pg_rca32_fa362_xor1[0], h_s_dadda_pg_rca32_fa363_xor1[0], h_s_dadda_pg_rca32_fa375_xor1, h_s_dadda_pg_rca32_fa375_or0);
  fa fa_h_s_dadda_pg_rca32_fa376_out(h_s_dadda_pg_rca32_fa364_xor1[0], h_s_dadda_pg_rca32_fa365_xor1[0], h_s_dadda_pg_rca32_fa366_xor1[0], h_s_dadda_pg_rca32_fa376_xor1, h_s_dadda_pg_rca32_fa376_or0);
  fa fa_h_s_dadda_pg_rca32_fa377_out(h_s_dadda_pg_rca32_fa367_xor1[0], h_s_dadda_pg_rca32_fa368_xor1[0], h_s_dadda_pg_rca32_fa369_xor1[0], h_s_dadda_pg_rca32_fa377_xor1, h_s_dadda_pg_rca32_fa377_or0);
  fa fa_h_s_dadda_pg_rca32_fa378_out(h_s_dadda_pg_rca32_fa370_xor1[0], h_s_dadda_pg_rca32_fa371_xor1[0], h_s_dadda_pg_rca32_fa372_xor1[0], h_s_dadda_pg_rca32_fa378_xor1, h_s_dadda_pg_rca32_fa378_or0);
  fa fa_h_s_dadda_pg_rca32_fa379_out(h_s_dadda_pg_rca32_fa378_or0[0], h_s_dadda_pg_rca32_fa377_or0[0], h_s_dadda_pg_rca32_fa376_or0[0], h_s_dadda_pg_rca32_fa379_xor1, h_s_dadda_pg_rca32_fa379_or0);
  fa fa_h_s_dadda_pg_rca32_fa380_out(h_s_dadda_pg_rca32_fa375_or0[0], h_s_dadda_pg_rca32_fa374_or0[0], h_s_dadda_pg_rca32_fa373_or0[0], h_s_dadda_pg_rca32_fa380_xor1, h_s_dadda_pg_rca32_fa380_or0);
  fa fa_h_s_dadda_pg_rca32_fa381_out(h_s_dadda_pg_rca32_fa372_or0[0], h_s_dadda_pg_rca32_fa371_or0[0], h_s_dadda_pg_rca32_fa370_or0[0], h_s_dadda_pg_rca32_fa381_xor1, h_s_dadda_pg_rca32_fa381_or0);
  fa fa_h_s_dadda_pg_rca32_fa382_out(h_s_dadda_pg_rca32_fa369_or0[0], h_s_dadda_pg_rca32_fa368_or0[0], h_s_dadda_pg_rca32_fa367_or0[0], h_s_dadda_pg_rca32_fa382_xor1, h_s_dadda_pg_rca32_fa382_or0);
  fa fa_h_s_dadda_pg_rca32_fa383_out(h_s_dadda_pg_rca32_fa366_or0[0], h_s_dadda_pg_rca32_fa365_or0[0], h_s_dadda_pg_rca32_fa364_or0[0], h_s_dadda_pg_rca32_fa383_xor1, h_s_dadda_pg_rca32_fa383_or0);
  fa fa_h_s_dadda_pg_rca32_fa384_out(h_s_dadda_pg_rca32_fa363_or0[0], h_s_dadda_pg_rca32_fa362_or0[0], h_s_dadda_pg_rca32_fa361_or0[0], h_s_dadda_pg_rca32_fa384_xor1, h_s_dadda_pg_rca32_fa384_or0);
  fa fa_h_s_dadda_pg_rca32_fa385_out(h_s_dadda_pg_rca32_fa360_or0[0], h_s_dadda_pg_rca32_fa359_or0[0], h_s_dadda_pg_rca32_fa358_or0[0], h_s_dadda_pg_rca32_fa385_xor1, h_s_dadda_pg_rca32_fa385_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_6(a[28], b[6], h_s_dadda_pg_rca32_and_28_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_7(a[27], b[7], h_s_dadda_pg_rca32_and_27_7);
  fa fa_h_s_dadda_pg_rca32_fa386_out(h_s_dadda_pg_rca32_fa357_or0[0], h_s_dadda_pg_rca32_and_28_6[0], h_s_dadda_pg_rca32_and_27_7[0], h_s_dadda_pg_rca32_fa386_xor1, h_s_dadda_pg_rca32_fa386_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_8(a[26], b[8], h_s_dadda_pg_rca32_and_26_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_9(a[25], b[9], h_s_dadda_pg_rca32_and_25_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_10(a[24], b[10], h_s_dadda_pg_rca32_and_24_10);
  fa fa_h_s_dadda_pg_rca32_fa387_out(h_s_dadda_pg_rca32_and_26_8[0], h_s_dadda_pg_rca32_and_25_9[0], h_s_dadda_pg_rca32_and_24_10[0], h_s_dadda_pg_rca32_fa387_xor1, h_s_dadda_pg_rca32_fa387_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_11(a[23], b[11], h_s_dadda_pg_rca32_and_23_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_12(a[22], b[12], h_s_dadda_pg_rca32_and_22_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_13(a[21], b[13], h_s_dadda_pg_rca32_and_21_13);
  fa fa_h_s_dadda_pg_rca32_fa388_out(h_s_dadda_pg_rca32_and_23_11[0], h_s_dadda_pg_rca32_and_22_12[0], h_s_dadda_pg_rca32_and_21_13[0], h_s_dadda_pg_rca32_fa388_xor1, h_s_dadda_pg_rca32_fa388_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_14(a[20], b[14], h_s_dadda_pg_rca32_and_20_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_15(a[19], b[15], h_s_dadda_pg_rca32_and_19_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_16(a[18], b[16], h_s_dadda_pg_rca32_and_18_16);
  fa fa_h_s_dadda_pg_rca32_fa389_out(h_s_dadda_pg_rca32_and_20_14[0], h_s_dadda_pg_rca32_and_19_15[0], h_s_dadda_pg_rca32_and_18_16[0], h_s_dadda_pg_rca32_fa389_xor1, h_s_dadda_pg_rca32_fa389_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_17(a[17], b[17], h_s_dadda_pg_rca32_and_17_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_18(a[16], b[18], h_s_dadda_pg_rca32_and_16_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_19(a[15], b[19], h_s_dadda_pg_rca32_and_15_19);
  fa fa_h_s_dadda_pg_rca32_fa390_out(h_s_dadda_pg_rca32_and_17_17[0], h_s_dadda_pg_rca32_and_16_18[0], h_s_dadda_pg_rca32_and_15_19[0], h_s_dadda_pg_rca32_fa390_xor1, h_s_dadda_pg_rca32_fa390_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_20(a[14], b[20], h_s_dadda_pg_rca32_and_14_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_21(a[13], b[21], h_s_dadda_pg_rca32_and_13_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_22(a[12], b[22], h_s_dadda_pg_rca32_and_12_22);
  fa fa_h_s_dadda_pg_rca32_fa391_out(h_s_dadda_pg_rca32_and_14_20[0], h_s_dadda_pg_rca32_and_13_21[0], h_s_dadda_pg_rca32_and_12_22[0], h_s_dadda_pg_rca32_fa391_xor1, h_s_dadda_pg_rca32_fa391_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_23(a[11], b[23], h_s_dadda_pg_rca32_and_11_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_24(a[10], b[24], h_s_dadda_pg_rca32_and_10_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_25(a[9], b[25], h_s_dadda_pg_rca32_and_9_25);
  fa fa_h_s_dadda_pg_rca32_fa392_out(h_s_dadda_pg_rca32_and_11_23[0], h_s_dadda_pg_rca32_and_10_24[0], h_s_dadda_pg_rca32_and_9_25[0], h_s_dadda_pg_rca32_fa392_xor1, h_s_dadda_pg_rca32_fa392_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_26(a[8], b[26], h_s_dadda_pg_rca32_and_8_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_27(a[7], b[27], h_s_dadda_pg_rca32_and_7_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_28(a[6], b[28], h_s_dadda_pg_rca32_and_6_28);
  fa fa_h_s_dadda_pg_rca32_fa393_out(h_s_dadda_pg_rca32_and_8_26[0], h_s_dadda_pg_rca32_and_7_27[0], h_s_dadda_pg_rca32_and_6_28[0], h_s_dadda_pg_rca32_fa393_xor1, h_s_dadda_pg_rca32_fa393_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_29(a[5], b[29], h_s_dadda_pg_rca32_and_5_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_30(a[4], b[30], h_s_dadda_pg_rca32_and_4_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_3_31(a[3], b[31], h_s_dadda_pg_rca32_nand_3_31);
  fa fa_h_s_dadda_pg_rca32_fa394_out(h_s_dadda_pg_rca32_and_5_29[0], h_s_dadda_pg_rca32_and_4_30[0], h_s_dadda_pg_rca32_nand_3_31[0], h_s_dadda_pg_rca32_fa394_xor1, h_s_dadda_pg_rca32_fa394_or0);
  fa fa_h_s_dadda_pg_rca32_fa395_out(h_s_dadda_pg_rca32_fa13_xor1[0], h_s_dadda_pg_rca32_fa14_xor1[0], h_s_dadda_pg_rca32_fa379_xor1[0], h_s_dadda_pg_rca32_fa395_xor1, h_s_dadda_pg_rca32_fa395_or0);
  fa fa_h_s_dadda_pg_rca32_fa396_out(h_s_dadda_pg_rca32_fa380_xor1[0], h_s_dadda_pg_rca32_fa381_xor1[0], h_s_dadda_pg_rca32_fa382_xor1[0], h_s_dadda_pg_rca32_fa396_xor1, h_s_dadda_pg_rca32_fa396_or0);
  fa fa_h_s_dadda_pg_rca32_fa397_out(h_s_dadda_pg_rca32_fa383_xor1[0], h_s_dadda_pg_rca32_fa384_xor1[0], h_s_dadda_pg_rca32_fa385_xor1[0], h_s_dadda_pg_rca32_fa397_xor1, h_s_dadda_pg_rca32_fa397_or0);
  fa fa_h_s_dadda_pg_rca32_fa398_out(h_s_dadda_pg_rca32_fa386_xor1[0], h_s_dadda_pg_rca32_fa387_xor1[0], h_s_dadda_pg_rca32_fa388_xor1[0], h_s_dadda_pg_rca32_fa398_xor1, h_s_dadda_pg_rca32_fa398_or0);
  fa fa_h_s_dadda_pg_rca32_fa399_out(h_s_dadda_pg_rca32_fa389_xor1[0], h_s_dadda_pg_rca32_fa390_xor1[0], h_s_dadda_pg_rca32_fa391_xor1[0], h_s_dadda_pg_rca32_fa399_xor1, h_s_dadda_pg_rca32_fa399_or0);
  fa fa_h_s_dadda_pg_rca32_fa400_out(h_s_dadda_pg_rca32_fa392_xor1[0], h_s_dadda_pg_rca32_fa393_xor1[0], h_s_dadda_pg_rca32_fa394_xor1[0], h_s_dadda_pg_rca32_fa400_xor1, h_s_dadda_pg_rca32_fa400_or0);
  fa fa_h_s_dadda_pg_rca32_fa401_out(h_s_dadda_pg_rca32_fa400_or0[0], h_s_dadda_pg_rca32_fa399_or0[0], h_s_dadda_pg_rca32_fa398_or0[0], h_s_dadda_pg_rca32_fa401_xor1, h_s_dadda_pg_rca32_fa401_or0);
  fa fa_h_s_dadda_pg_rca32_fa402_out(h_s_dadda_pg_rca32_fa397_or0[0], h_s_dadda_pg_rca32_fa396_or0[0], h_s_dadda_pg_rca32_fa395_or0[0], h_s_dadda_pg_rca32_fa402_xor1, h_s_dadda_pg_rca32_fa402_or0);
  fa fa_h_s_dadda_pg_rca32_fa403_out(h_s_dadda_pg_rca32_fa394_or0[0], h_s_dadda_pg_rca32_fa393_or0[0], h_s_dadda_pg_rca32_fa392_or0[0], h_s_dadda_pg_rca32_fa403_xor1, h_s_dadda_pg_rca32_fa403_or0);
  fa fa_h_s_dadda_pg_rca32_fa404_out(h_s_dadda_pg_rca32_fa391_or0[0], h_s_dadda_pg_rca32_fa390_or0[0], h_s_dadda_pg_rca32_fa389_or0[0], h_s_dadda_pg_rca32_fa404_xor1, h_s_dadda_pg_rca32_fa404_or0);
  fa fa_h_s_dadda_pg_rca32_fa405_out(h_s_dadda_pg_rca32_fa388_or0[0], h_s_dadda_pg_rca32_fa387_or0[0], h_s_dadda_pg_rca32_fa386_or0[0], h_s_dadda_pg_rca32_fa405_xor1, h_s_dadda_pg_rca32_fa405_or0);
  fa fa_h_s_dadda_pg_rca32_fa406_out(h_s_dadda_pg_rca32_fa385_or0[0], h_s_dadda_pg_rca32_fa384_or0[0], h_s_dadda_pg_rca32_fa383_or0[0], h_s_dadda_pg_rca32_fa406_xor1, h_s_dadda_pg_rca32_fa406_or0);
  fa fa_h_s_dadda_pg_rca32_fa407_out(h_s_dadda_pg_rca32_fa382_or0[0], h_s_dadda_pg_rca32_fa381_or0[0], h_s_dadda_pg_rca32_fa380_or0[0], h_s_dadda_pg_rca32_fa407_xor1, h_s_dadda_pg_rca32_fa407_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_5(a[30], b[5], h_s_dadda_pg_rca32_and_30_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_6(a[29], b[6], h_s_dadda_pg_rca32_and_29_6);
  fa fa_h_s_dadda_pg_rca32_fa408_out(h_s_dadda_pg_rca32_fa379_or0[0], h_s_dadda_pg_rca32_and_30_5[0], h_s_dadda_pg_rca32_and_29_6[0], h_s_dadda_pg_rca32_fa408_xor1, h_s_dadda_pg_rca32_fa408_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_7(a[28], b[7], h_s_dadda_pg_rca32_and_28_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_8(a[27], b[8], h_s_dadda_pg_rca32_and_27_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_9(a[26], b[9], h_s_dadda_pg_rca32_and_26_9);
  fa fa_h_s_dadda_pg_rca32_fa409_out(h_s_dadda_pg_rca32_and_28_7[0], h_s_dadda_pg_rca32_and_27_8[0], h_s_dadda_pg_rca32_and_26_9[0], h_s_dadda_pg_rca32_fa409_xor1, h_s_dadda_pg_rca32_fa409_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_10(a[25], b[10], h_s_dadda_pg_rca32_and_25_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_11(a[24], b[11], h_s_dadda_pg_rca32_and_24_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_12(a[23], b[12], h_s_dadda_pg_rca32_and_23_12);
  fa fa_h_s_dadda_pg_rca32_fa410_out(h_s_dadda_pg_rca32_and_25_10[0], h_s_dadda_pg_rca32_and_24_11[0], h_s_dadda_pg_rca32_and_23_12[0], h_s_dadda_pg_rca32_fa410_xor1, h_s_dadda_pg_rca32_fa410_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_13(a[22], b[13], h_s_dadda_pg_rca32_and_22_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_14(a[21], b[14], h_s_dadda_pg_rca32_and_21_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_15(a[20], b[15], h_s_dadda_pg_rca32_and_20_15);
  fa fa_h_s_dadda_pg_rca32_fa411_out(h_s_dadda_pg_rca32_and_22_13[0], h_s_dadda_pg_rca32_and_21_14[0], h_s_dadda_pg_rca32_and_20_15[0], h_s_dadda_pg_rca32_fa411_xor1, h_s_dadda_pg_rca32_fa411_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_16(a[19], b[16], h_s_dadda_pg_rca32_and_19_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_17(a[18], b[17], h_s_dadda_pg_rca32_and_18_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_18(a[17], b[18], h_s_dadda_pg_rca32_and_17_18);
  fa fa_h_s_dadda_pg_rca32_fa412_out(h_s_dadda_pg_rca32_and_19_16[0], h_s_dadda_pg_rca32_and_18_17[0], h_s_dadda_pg_rca32_and_17_18[0], h_s_dadda_pg_rca32_fa412_xor1, h_s_dadda_pg_rca32_fa412_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_19(a[16], b[19], h_s_dadda_pg_rca32_and_16_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_20(a[15], b[20], h_s_dadda_pg_rca32_and_15_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_21(a[14], b[21], h_s_dadda_pg_rca32_and_14_21);
  fa fa_h_s_dadda_pg_rca32_fa413_out(h_s_dadda_pg_rca32_and_16_19[0], h_s_dadda_pg_rca32_and_15_20[0], h_s_dadda_pg_rca32_and_14_21[0], h_s_dadda_pg_rca32_fa413_xor1, h_s_dadda_pg_rca32_fa413_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_22(a[13], b[22], h_s_dadda_pg_rca32_and_13_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_23(a[12], b[23], h_s_dadda_pg_rca32_and_12_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_24(a[11], b[24], h_s_dadda_pg_rca32_and_11_24);
  fa fa_h_s_dadda_pg_rca32_fa414_out(h_s_dadda_pg_rca32_and_13_22[0], h_s_dadda_pg_rca32_and_12_23[0], h_s_dadda_pg_rca32_and_11_24[0], h_s_dadda_pg_rca32_fa414_xor1, h_s_dadda_pg_rca32_fa414_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_25(a[10], b[25], h_s_dadda_pg_rca32_and_10_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_26(a[9], b[26], h_s_dadda_pg_rca32_and_9_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_27(a[8], b[27], h_s_dadda_pg_rca32_and_8_27);
  fa fa_h_s_dadda_pg_rca32_fa415_out(h_s_dadda_pg_rca32_and_10_25[0], h_s_dadda_pg_rca32_and_9_26[0], h_s_dadda_pg_rca32_and_8_27[0], h_s_dadda_pg_rca32_fa415_xor1, h_s_dadda_pg_rca32_fa415_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_28(a[7], b[28], h_s_dadda_pg_rca32_and_7_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_29(a[6], b[29], h_s_dadda_pg_rca32_and_6_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_30(a[5], b[30], h_s_dadda_pg_rca32_and_5_30);
  fa fa_h_s_dadda_pg_rca32_fa416_out(h_s_dadda_pg_rca32_and_7_28[0], h_s_dadda_pg_rca32_and_6_29[0], h_s_dadda_pg_rca32_and_5_30[0], h_s_dadda_pg_rca32_fa416_xor1, h_s_dadda_pg_rca32_fa416_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_4_31(a[4], b[31], h_s_dadda_pg_rca32_nand_4_31);
  fa fa_h_s_dadda_pg_rca32_fa417_out(h_s_dadda_pg_rca32_nand_4_31[0], h_s_dadda_pg_rca32_fa15_xor1[0], h_s_dadda_pg_rca32_fa401_xor1[0], h_s_dadda_pg_rca32_fa417_xor1, h_s_dadda_pg_rca32_fa417_or0);
  fa fa_h_s_dadda_pg_rca32_fa418_out(h_s_dadda_pg_rca32_fa402_xor1[0], h_s_dadda_pg_rca32_fa403_xor1[0], h_s_dadda_pg_rca32_fa404_xor1[0], h_s_dadda_pg_rca32_fa418_xor1, h_s_dadda_pg_rca32_fa418_or0);
  fa fa_h_s_dadda_pg_rca32_fa419_out(h_s_dadda_pg_rca32_fa405_xor1[0], h_s_dadda_pg_rca32_fa406_xor1[0], h_s_dadda_pg_rca32_fa407_xor1[0], h_s_dadda_pg_rca32_fa419_xor1, h_s_dadda_pg_rca32_fa419_or0);
  fa fa_h_s_dadda_pg_rca32_fa420_out(h_s_dadda_pg_rca32_fa408_xor1[0], h_s_dadda_pg_rca32_fa409_xor1[0], h_s_dadda_pg_rca32_fa410_xor1[0], h_s_dadda_pg_rca32_fa420_xor1, h_s_dadda_pg_rca32_fa420_or0);
  fa fa_h_s_dadda_pg_rca32_fa421_out(h_s_dadda_pg_rca32_fa411_xor1[0], h_s_dadda_pg_rca32_fa412_xor1[0], h_s_dadda_pg_rca32_fa413_xor1[0], h_s_dadda_pg_rca32_fa421_xor1, h_s_dadda_pg_rca32_fa421_or0);
  fa fa_h_s_dadda_pg_rca32_fa422_out(h_s_dadda_pg_rca32_fa414_xor1[0], h_s_dadda_pg_rca32_fa415_xor1[0], h_s_dadda_pg_rca32_fa416_xor1[0], h_s_dadda_pg_rca32_fa422_xor1, h_s_dadda_pg_rca32_fa422_or0);
  fa fa_h_s_dadda_pg_rca32_fa423_out(h_s_dadda_pg_rca32_fa422_or0[0], h_s_dadda_pg_rca32_fa421_or0[0], h_s_dadda_pg_rca32_fa420_or0[0], h_s_dadda_pg_rca32_fa423_xor1, h_s_dadda_pg_rca32_fa423_or0);
  fa fa_h_s_dadda_pg_rca32_fa424_out(h_s_dadda_pg_rca32_fa419_or0[0], h_s_dadda_pg_rca32_fa418_or0[0], h_s_dadda_pg_rca32_fa417_or0[0], h_s_dadda_pg_rca32_fa424_xor1, h_s_dadda_pg_rca32_fa424_or0);
  fa fa_h_s_dadda_pg_rca32_fa425_out(h_s_dadda_pg_rca32_fa416_or0[0], h_s_dadda_pg_rca32_fa415_or0[0], h_s_dadda_pg_rca32_fa414_or0[0], h_s_dadda_pg_rca32_fa425_xor1, h_s_dadda_pg_rca32_fa425_or0);
  fa fa_h_s_dadda_pg_rca32_fa426_out(h_s_dadda_pg_rca32_fa413_or0[0], h_s_dadda_pg_rca32_fa412_or0[0], h_s_dadda_pg_rca32_fa411_or0[0], h_s_dadda_pg_rca32_fa426_xor1, h_s_dadda_pg_rca32_fa426_or0);
  fa fa_h_s_dadda_pg_rca32_fa427_out(h_s_dadda_pg_rca32_fa410_or0[0], h_s_dadda_pg_rca32_fa409_or0[0], h_s_dadda_pg_rca32_fa408_or0[0], h_s_dadda_pg_rca32_fa427_xor1, h_s_dadda_pg_rca32_fa427_or0);
  fa fa_h_s_dadda_pg_rca32_fa428_out(h_s_dadda_pg_rca32_fa407_or0[0], h_s_dadda_pg_rca32_fa406_or0[0], h_s_dadda_pg_rca32_fa405_or0[0], h_s_dadda_pg_rca32_fa428_xor1, h_s_dadda_pg_rca32_fa428_or0);
  fa fa_h_s_dadda_pg_rca32_fa429_out(h_s_dadda_pg_rca32_fa404_or0[0], h_s_dadda_pg_rca32_fa403_or0[0], h_s_dadda_pg_rca32_fa402_or0[0], h_s_dadda_pg_rca32_fa429_xor1, h_s_dadda_pg_rca32_fa429_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_5(a[31], b[5], h_s_dadda_pg_rca32_nand_31_5);
  fa fa_h_s_dadda_pg_rca32_fa430_out(h_s_dadda_pg_rca32_fa401_or0[0], h_s_dadda_pg_rca32_fa15_or0[0], h_s_dadda_pg_rca32_nand_31_5[0], h_s_dadda_pg_rca32_fa430_xor1, h_s_dadda_pg_rca32_fa430_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_6(a[30], b[6], h_s_dadda_pg_rca32_and_30_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_7(a[29], b[7], h_s_dadda_pg_rca32_and_29_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_8(a[28], b[8], h_s_dadda_pg_rca32_and_28_8);
  fa fa_h_s_dadda_pg_rca32_fa431_out(h_s_dadda_pg_rca32_and_30_6[0], h_s_dadda_pg_rca32_and_29_7[0], h_s_dadda_pg_rca32_and_28_8[0], h_s_dadda_pg_rca32_fa431_xor1, h_s_dadda_pg_rca32_fa431_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_9(a[27], b[9], h_s_dadda_pg_rca32_and_27_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_10(a[26], b[10], h_s_dadda_pg_rca32_and_26_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_11(a[25], b[11], h_s_dadda_pg_rca32_and_25_11);
  fa fa_h_s_dadda_pg_rca32_fa432_out(h_s_dadda_pg_rca32_and_27_9[0], h_s_dadda_pg_rca32_and_26_10[0], h_s_dadda_pg_rca32_and_25_11[0], h_s_dadda_pg_rca32_fa432_xor1, h_s_dadda_pg_rca32_fa432_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_12(a[24], b[12], h_s_dadda_pg_rca32_and_24_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_13(a[23], b[13], h_s_dadda_pg_rca32_and_23_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_14(a[22], b[14], h_s_dadda_pg_rca32_and_22_14);
  fa fa_h_s_dadda_pg_rca32_fa433_out(h_s_dadda_pg_rca32_and_24_12[0], h_s_dadda_pg_rca32_and_23_13[0], h_s_dadda_pg_rca32_and_22_14[0], h_s_dadda_pg_rca32_fa433_xor1, h_s_dadda_pg_rca32_fa433_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_15(a[21], b[15], h_s_dadda_pg_rca32_and_21_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_16(a[20], b[16], h_s_dadda_pg_rca32_and_20_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_17(a[19], b[17], h_s_dadda_pg_rca32_and_19_17);
  fa fa_h_s_dadda_pg_rca32_fa434_out(h_s_dadda_pg_rca32_and_21_15[0], h_s_dadda_pg_rca32_and_20_16[0], h_s_dadda_pg_rca32_and_19_17[0], h_s_dadda_pg_rca32_fa434_xor1, h_s_dadda_pg_rca32_fa434_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_18(a[18], b[18], h_s_dadda_pg_rca32_and_18_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_19(a[17], b[19], h_s_dadda_pg_rca32_and_17_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_20(a[16], b[20], h_s_dadda_pg_rca32_and_16_20);
  fa fa_h_s_dadda_pg_rca32_fa435_out(h_s_dadda_pg_rca32_and_18_18[0], h_s_dadda_pg_rca32_and_17_19[0], h_s_dadda_pg_rca32_and_16_20[0], h_s_dadda_pg_rca32_fa435_xor1, h_s_dadda_pg_rca32_fa435_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_21(a[15], b[21], h_s_dadda_pg_rca32_and_15_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_22(a[14], b[22], h_s_dadda_pg_rca32_and_14_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_23(a[13], b[23], h_s_dadda_pg_rca32_and_13_23);
  fa fa_h_s_dadda_pg_rca32_fa436_out(h_s_dadda_pg_rca32_and_15_21[0], h_s_dadda_pg_rca32_and_14_22[0], h_s_dadda_pg_rca32_and_13_23[0], h_s_dadda_pg_rca32_fa436_xor1, h_s_dadda_pg_rca32_fa436_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_24(a[12], b[24], h_s_dadda_pg_rca32_and_12_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_25(a[11], b[25], h_s_dadda_pg_rca32_and_11_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_26(a[10], b[26], h_s_dadda_pg_rca32_and_10_26);
  fa fa_h_s_dadda_pg_rca32_fa437_out(h_s_dadda_pg_rca32_and_12_24[0], h_s_dadda_pg_rca32_and_11_25[0], h_s_dadda_pg_rca32_and_10_26[0], h_s_dadda_pg_rca32_fa437_xor1, h_s_dadda_pg_rca32_fa437_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_27(a[9], b[27], h_s_dadda_pg_rca32_and_9_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_28(a[8], b[28], h_s_dadda_pg_rca32_and_8_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_29(a[7], b[29], h_s_dadda_pg_rca32_and_7_29);
  fa fa_h_s_dadda_pg_rca32_fa438_out(h_s_dadda_pg_rca32_and_9_27[0], h_s_dadda_pg_rca32_and_8_28[0], h_s_dadda_pg_rca32_and_7_29[0], h_s_dadda_pg_rca32_fa438_xor1, h_s_dadda_pg_rca32_fa438_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_6_30(a[6], b[30], h_s_dadda_pg_rca32_and_6_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_5_31(a[5], b[31], h_s_dadda_pg_rca32_nand_5_31);
  fa fa_h_s_dadda_pg_rca32_fa439_out(h_s_dadda_pg_rca32_and_6_30[0], h_s_dadda_pg_rca32_nand_5_31[0], h_s_dadda_pg_rca32_fa423_xor1[0], h_s_dadda_pg_rca32_fa439_xor1, h_s_dadda_pg_rca32_fa439_or0);
  fa fa_h_s_dadda_pg_rca32_fa440_out(h_s_dadda_pg_rca32_fa424_xor1[0], h_s_dadda_pg_rca32_fa425_xor1[0], h_s_dadda_pg_rca32_fa426_xor1[0], h_s_dadda_pg_rca32_fa440_xor1, h_s_dadda_pg_rca32_fa440_or0);
  fa fa_h_s_dadda_pg_rca32_fa441_out(h_s_dadda_pg_rca32_fa427_xor1[0], h_s_dadda_pg_rca32_fa428_xor1[0], h_s_dadda_pg_rca32_fa429_xor1[0], h_s_dadda_pg_rca32_fa441_xor1, h_s_dadda_pg_rca32_fa441_or0);
  fa fa_h_s_dadda_pg_rca32_fa442_out(h_s_dadda_pg_rca32_fa430_xor1[0], h_s_dadda_pg_rca32_fa431_xor1[0], h_s_dadda_pg_rca32_fa432_xor1[0], h_s_dadda_pg_rca32_fa442_xor1, h_s_dadda_pg_rca32_fa442_or0);
  fa fa_h_s_dadda_pg_rca32_fa443_out(h_s_dadda_pg_rca32_fa433_xor1[0], h_s_dadda_pg_rca32_fa434_xor1[0], h_s_dadda_pg_rca32_fa435_xor1[0], h_s_dadda_pg_rca32_fa443_xor1, h_s_dadda_pg_rca32_fa443_or0);
  fa fa_h_s_dadda_pg_rca32_fa444_out(h_s_dadda_pg_rca32_fa436_xor1[0], h_s_dadda_pg_rca32_fa437_xor1[0], h_s_dadda_pg_rca32_fa438_xor1[0], h_s_dadda_pg_rca32_fa444_xor1, h_s_dadda_pg_rca32_fa444_or0);
  fa fa_h_s_dadda_pg_rca32_fa445_out(h_s_dadda_pg_rca32_fa444_or0[0], h_s_dadda_pg_rca32_fa443_or0[0], h_s_dadda_pg_rca32_fa442_or0[0], h_s_dadda_pg_rca32_fa445_xor1, h_s_dadda_pg_rca32_fa445_or0);
  fa fa_h_s_dadda_pg_rca32_fa446_out(h_s_dadda_pg_rca32_fa441_or0[0], h_s_dadda_pg_rca32_fa440_or0[0], h_s_dadda_pg_rca32_fa439_or0[0], h_s_dadda_pg_rca32_fa446_xor1, h_s_dadda_pg_rca32_fa446_or0);
  fa fa_h_s_dadda_pg_rca32_fa447_out(h_s_dadda_pg_rca32_fa438_or0[0], h_s_dadda_pg_rca32_fa437_or0[0], h_s_dadda_pg_rca32_fa436_or0[0], h_s_dadda_pg_rca32_fa447_xor1, h_s_dadda_pg_rca32_fa447_or0);
  fa fa_h_s_dadda_pg_rca32_fa448_out(h_s_dadda_pg_rca32_fa435_or0[0], h_s_dadda_pg_rca32_fa434_or0[0], h_s_dadda_pg_rca32_fa433_or0[0], h_s_dadda_pg_rca32_fa448_xor1, h_s_dadda_pg_rca32_fa448_or0);
  fa fa_h_s_dadda_pg_rca32_fa449_out(h_s_dadda_pg_rca32_fa432_or0[0], h_s_dadda_pg_rca32_fa431_or0[0], h_s_dadda_pg_rca32_fa430_or0[0], h_s_dadda_pg_rca32_fa449_xor1, h_s_dadda_pg_rca32_fa449_or0);
  fa fa_h_s_dadda_pg_rca32_fa450_out(h_s_dadda_pg_rca32_fa429_or0[0], h_s_dadda_pg_rca32_fa428_or0[0], h_s_dadda_pg_rca32_fa427_or0[0], h_s_dadda_pg_rca32_fa450_xor1, h_s_dadda_pg_rca32_fa450_or0);
  fa fa_h_s_dadda_pg_rca32_fa451_out(h_s_dadda_pg_rca32_fa426_or0[0], h_s_dadda_pg_rca32_fa425_or0[0], h_s_dadda_pg_rca32_fa424_or0[0], h_s_dadda_pg_rca32_fa451_xor1, h_s_dadda_pg_rca32_fa451_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_6(a[31], b[6], h_s_dadda_pg_rca32_nand_31_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_7(a[30], b[7], h_s_dadda_pg_rca32_and_30_7);
  fa fa_h_s_dadda_pg_rca32_fa452_out(h_s_dadda_pg_rca32_fa423_or0[0], h_s_dadda_pg_rca32_nand_31_6[0], h_s_dadda_pg_rca32_and_30_7[0], h_s_dadda_pg_rca32_fa452_xor1, h_s_dadda_pg_rca32_fa452_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_8(a[29], b[8], h_s_dadda_pg_rca32_and_29_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_9(a[28], b[9], h_s_dadda_pg_rca32_and_28_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_10(a[27], b[10], h_s_dadda_pg_rca32_and_27_10);
  fa fa_h_s_dadda_pg_rca32_fa453_out(h_s_dadda_pg_rca32_and_29_8[0], h_s_dadda_pg_rca32_and_28_9[0], h_s_dadda_pg_rca32_and_27_10[0], h_s_dadda_pg_rca32_fa453_xor1, h_s_dadda_pg_rca32_fa453_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_11(a[26], b[11], h_s_dadda_pg_rca32_and_26_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_12(a[25], b[12], h_s_dadda_pg_rca32_and_25_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_13(a[24], b[13], h_s_dadda_pg_rca32_and_24_13);
  fa fa_h_s_dadda_pg_rca32_fa454_out(h_s_dadda_pg_rca32_and_26_11[0], h_s_dadda_pg_rca32_and_25_12[0], h_s_dadda_pg_rca32_and_24_13[0], h_s_dadda_pg_rca32_fa454_xor1, h_s_dadda_pg_rca32_fa454_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_14(a[23], b[14], h_s_dadda_pg_rca32_and_23_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_15(a[22], b[15], h_s_dadda_pg_rca32_and_22_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_16(a[21], b[16], h_s_dadda_pg_rca32_and_21_16);
  fa fa_h_s_dadda_pg_rca32_fa455_out(h_s_dadda_pg_rca32_and_23_14[0], h_s_dadda_pg_rca32_and_22_15[0], h_s_dadda_pg_rca32_and_21_16[0], h_s_dadda_pg_rca32_fa455_xor1, h_s_dadda_pg_rca32_fa455_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_17(a[20], b[17], h_s_dadda_pg_rca32_and_20_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_18(a[19], b[18], h_s_dadda_pg_rca32_and_19_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_19(a[18], b[19], h_s_dadda_pg_rca32_and_18_19);
  fa fa_h_s_dadda_pg_rca32_fa456_out(h_s_dadda_pg_rca32_and_20_17[0], h_s_dadda_pg_rca32_and_19_18[0], h_s_dadda_pg_rca32_and_18_19[0], h_s_dadda_pg_rca32_fa456_xor1, h_s_dadda_pg_rca32_fa456_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_20(a[17], b[20], h_s_dadda_pg_rca32_and_17_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_21(a[16], b[21], h_s_dadda_pg_rca32_and_16_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_22(a[15], b[22], h_s_dadda_pg_rca32_and_15_22);
  fa fa_h_s_dadda_pg_rca32_fa457_out(h_s_dadda_pg_rca32_and_17_20[0], h_s_dadda_pg_rca32_and_16_21[0], h_s_dadda_pg_rca32_and_15_22[0], h_s_dadda_pg_rca32_fa457_xor1, h_s_dadda_pg_rca32_fa457_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_23(a[14], b[23], h_s_dadda_pg_rca32_and_14_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_24(a[13], b[24], h_s_dadda_pg_rca32_and_13_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_25(a[12], b[25], h_s_dadda_pg_rca32_and_12_25);
  fa fa_h_s_dadda_pg_rca32_fa458_out(h_s_dadda_pg_rca32_and_14_23[0], h_s_dadda_pg_rca32_and_13_24[0], h_s_dadda_pg_rca32_and_12_25[0], h_s_dadda_pg_rca32_fa458_xor1, h_s_dadda_pg_rca32_fa458_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_26(a[11], b[26], h_s_dadda_pg_rca32_and_11_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_27(a[10], b[27], h_s_dadda_pg_rca32_and_10_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_28(a[9], b[28], h_s_dadda_pg_rca32_and_9_28);
  fa fa_h_s_dadda_pg_rca32_fa459_out(h_s_dadda_pg_rca32_and_11_26[0], h_s_dadda_pg_rca32_and_10_27[0], h_s_dadda_pg_rca32_and_9_28[0], h_s_dadda_pg_rca32_fa459_xor1, h_s_dadda_pg_rca32_fa459_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_29(a[8], b[29], h_s_dadda_pg_rca32_and_8_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_7_30(a[7], b[30], h_s_dadda_pg_rca32_and_7_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_6_31(a[6], b[31], h_s_dadda_pg_rca32_nand_6_31);
  fa fa_h_s_dadda_pg_rca32_fa460_out(h_s_dadda_pg_rca32_and_8_29[0], h_s_dadda_pg_rca32_and_7_30[0], h_s_dadda_pg_rca32_nand_6_31[0], h_s_dadda_pg_rca32_fa460_xor1, h_s_dadda_pg_rca32_fa460_or0);
  fa fa_h_s_dadda_pg_rca32_fa461_out(h_s_dadda_pg_rca32_fa445_xor1[0], h_s_dadda_pg_rca32_fa446_xor1[0], h_s_dadda_pg_rca32_fa447_xor1[0], h_s_dadda_pg_rca32_fa461_xor1, h_s_dadda_pg_rca32_fa461_or0);
  fa fa_h_s_dadda_pg_rca32_fa462_out(h_s_dadda_pg_rca32_fa448_xor1[0], h_s_dadda_pg_rca32_fa449_xor1[0], h_s_dadda_pg_rca32_fa450_xor1[0], h_s_dadda_pg_rca32_fa462_xor1, h_s_dadda_pg_rca32_fa462_or0);
  fa fa_h_s_dadda_pg_rca32_fa463_out(h_s_dadda_pg_rca32_fa451_xor1[0], h_s_dadda_pg_rca32_fa452_xor1[0], h_s_dadda_pg_rca32_fa453_xor1[0], h_s_dadda_pg_rca32_fa463_xor1, h_s_dadda_pg_rca32_fa463_or0);
  fa fa_h_s_dadda_pg_rca32_fa464_out(h_s_dadda_pg_rca32_fa454_xor1[0], h_s_dadda_pg_rca32_fa455_xor1[0], h_s_dadda_pg_rca32_fa456_xor1[0], h_s_dadda_pg_rca32_fa464_xor1, h_s_dadda_pg_rca32_fa464_or0);
  fa fa_h_s_dadda_pg_rca32_fa465_out(h_s_dadda_pg_rca32_fa457_xor1[0], h_s_dadda_pg_rca32_fa458_xor1[0], h_s_dadda_pg_rca32_fa459_xor1[0], h_s_dadda_pg_rca32_fa465_xor1, h_s_dadda_pg_rca32_fa465_or0);
  fa fa_h_s_dadda_pg_rca32_fa466_out(h_s_dadda_pg_rca32_fa465_or0[0], h_s_dadda_pg_rca32_fa464_or0[0], h_s_dadda_pg_rca32_fa463_or0[0], h_s_dadda_pg_rca32_fa466_xor1, h_s_dadda_pg_rca32_fa466_or0);
  fa fa_h_s_dadda_pg_rca32_fa467_out(h_s_dadda_pg_rca32_fa462_or0[0], h_s_dadda_pg_rca32_fa461_or0[0], h_s_dadda_pg_rca32_fa460_or0[0], h_s_dadda_pg_rca32_fa467_xor1, h_s_dadda_pg_rca32_fa467_or0);
  fa fa_h_s_dadda_pg_rca32_fa468_out(h_s_dadda_pg_rca32_fa459_or0[0], h_s_dadda_pg_rca32_fa458_or0[0], h_s_dadda_pg_rca32_fa457_or0[0], h_s_dadda_pg_rca32_fa468_xor1, h_s_dadda_pg_rca32_fa468_or0);
  fa fa_h_s_dadda_pg_rca32_fa469_out(h_s_dadda_pg_rca32_fa456_or0[0], h_s_dadda_pg_rca32_fa455_or0[0], h_s_dadda_pg_rca32_fa454_or0[0], h_s_dadda_pg_rca32_fa469_xor1, h_s_dadda_pg_rca32_fa469_or0);
  fa fa_h_s_dadda_pg_rca32_fa470_out(h_s_dadda_pg_rca32_fa453_or0[0], h_s_dadda_pg_rca32_fa452_or0[0], h_s_dadda_pg_rca32_fa451_or0[0], h_s_dadda_pg_rca32_fa470_xor1, h_s_dadda_pg_rca32_fa470_or0);
  fa fa_h_s_dadda_pg_rca32_fa471_out(h_s_dadda_pg_rca32_fa450_or0[0], h_s_dadda_pg_rca32_fa449_or0[0], h_s_dadda_pg_rca32_fa448_or0[0], h_s_dadda_pg_rca32_fa471_xor1, h_s_dadda_pg_rca32_fa471_or0);
  fa fa_h_s_dadda_pg_rca32_fa472_out(h_s_dadda_pg_rca32_fa447_or0[0], h_s_dadda_pg_rca32_fa446_or0[0], h_s_dadda_pg_rca32_fa445_or0[0], h_s_dadda_pg_rca32_fa472_xor1, h_s_dadda_pg_rca32_fa472_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_7(a[31], b[7], h_s_dadda_pg_rca32_nand_31_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_8(a[30], b[8], h_s_dadda_pg_rca32_and_30_8);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_9(a[29], b[9], h_s_dadda_pg_rca32_and_29_9);
  fa fa_h_s_dadda_pg_rca32_fa473_out(h_s_dadda_pg_rca32_nand_31_7[0], h_s_dadda_pg_rca32_and_30_8[0], h_s_dadda_pg_rca32_and_29_9[0], h_s_dadda_pg_rca32_fa473_xor1, h_s_dadda_pg_rca32_fa473_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_10(a[28], b[10], h_s_dadda_pg_rca32_and_28_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_11(a[27], b[11], h_s_dadda_pg_rca32_and_27_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_12(a[26], b[12], h_s_dadda_pg_rca32_and_26_12);
  fa fa_h_s_dadda_pg_rca32_fa474_out(h_s_dadda_pg_rca32_and_28_10[0], h_s_dadda_pg_rca32_and_27_11[0], h_s_dadda_pg_rca32_and_26_12[0], h_s_dadda_pg_rca32_fa474_xor1, h_s_dadda_pg_rca32_fa474_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_13(a[25], b[13], h_s_dadda_pg_rca32_and_25_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_14(a[24], b[14], h_s_dadda_pg_rca32_and_24_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_15(a[23], b[15], h_s_dadda_pg_rca32_and_23_15);
  fa fa_h_s_dadda_pg_rca32_fa475_out(h_s_dadda_pg_rca32_and_25_13[0], h_s_dadda_pg_rca32_and_24_14[0], h_s_dadda_pg_rca32_and_23_15[0], h_s_dadda_pg_rca32_fa475_xor1, h_s_dadda_pg_rca32_fa475_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_16(a[22], b[16], h_s_dadda_pg_rca32_and_22_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_17(a[21], b[17], h_s_dadda_pg_rca32_and_21_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_18(a[20], b[18], h_s_dadda_pg_rca32_and_20_18);
  fa fa_h_s_dadda_pg_rca32_fa476_out(h_s_dadda_pg_rca32_and_22_16[0], h_s_dadda_pg_rca32_and_21_17[0], h_s_dadda_pg_rca32_and_20_18[0], h_s_dadda_pg_rca32_fa476_xor1, h_s_dadda_pg_rca32_fa476_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_19(a[19], b[19], h_s_dadda_pg_rca32_and_19_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_20(a[18], b[20], h_s_dadda_pg_rca32_and_18_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_21(a[17], b[21], h_s_dadda_pg_rca32_and_17_21);
  fa fa_h_s_dadda_pg_rca32_fa477_out(h_s_dadda_pg_rca32_and_19_19[0], h_s_dadda_pg_rca32_and_18_20[0], h_s_dadda_pg_rca32_and_17_21[0], h_s_dadda_pg_rca32_fa477_xor1, h_s_dadda_pg_rca32_fa477_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_22(a[16], b[22], h_s_dadda_pg_rca32_and_16_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_23(a[15], b[23], h_s_dadda_pg_rca32_and_15_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_24(a[14], b[24], h_s_dadda_pg_rca32_and_14_24);
  fa fa_h_s_dadda_pg_rca32_fa478_out(h_s_dadda_pg_rca32_and_16_22[0], h_s_dadda_pg_rca32_and_15_23[0], h_s_dadda_pg_rca32_and_14_24[0], h_s_dadda_pg_rca32_fa478_xor1, h_s_dadda_pg_rca32_fa478_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_25(a[13], b[25], h_s_dadda_pg_rca32_and_13_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_26(a[12], b[26], h_s_dadda_pg_rca32_and_12_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_27(a[11], b[27], h_s_dadda_pg_rca32_and_11_27);
  fa fa_h_s_dadda_pg_rca32_fa479_out(h_s_dadda_pg_rca32_and_13_25[0], h_s_dadda_pg_rca32_and_12_26[0], h_s_dadda_pg_rca32_and_11_27[0], h_s_dadda_pg_rca32_fa479_xor1, h_s_dadda_pg_rca32_fa479_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_28(a[10], b[28], h_s_dadda_pg_rca32_and_10_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_29(a[9], b[29], h_s_dadda_pg_rca32_and_9_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_8_30(a[8], b[30], h_s_dadda_pg_rca32_and_8_30);
  fa fa_h_s_dadda_pg_rca32_fa480_out(h_s_dadda_pg_rca32_and_10_28[0], h_s_dadda_pg_rca32_and_9_29[0], h_s_dadda_pg_rca32_and_8_30[0], h_s_dadda_pg_rca32_fa480_xor1, h_s_dadda_pg_rca32_fa480_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_7_31(a[7], b[31], h_s_dadda_pg_rca32_nand_7_31);
  fa fa_h_s_dadda_pg_rca32_fa481_out(h_s_dadda_pg_rca32_nand_7_31[0], h_s_dadda_pg_rca32_fa466_xor1[0], h_s_dadda_pg_rca32_fa467_xor1[0], h_s_dadda_pg_rca32_fa481_xor1, h_s_dadda_pg_rca32_fa481_or0);
  fa fa_h_s_dadda_pg_rca32_fa482_out(h_s_dadda_pg_rca32_fa468_xor1[0], h_s_dadda_pg_rca32_fa469_xor1[0], h_s_dadda_pg_rca32_fa470_xor1[0], h_s_dadda_pg_rca32_fa482_xor1, h_s_dadda_pg_rca32_fa482_or0);
  fa fa_h_s_dadda_pg_rca32_fa483_out(h_s_dadda_pg_rca32_fa471_xor1[0], h_s_dadda_pg_rca32_fa472_xor1[0], h_s_dadda_pg_rca32_fa473_xor1[0], h_s_dadda_pg_rca32_fa483_xor1, h_s_dadda_pg_rca32_fa483_or0);
  fa fa_h_s_dadda_pg_rca32_fa484_out(h_s_dadda_pg_rca32_fa474_xor1[0], h_s_dadda_pg_rca32_fa475_xor1[0], h_s_dadda_pg_rca32_fa476_xor1[0], h_s_dadda_pg_rca32_fa484_xor1, h_s_dadda_pg_rca32_fa484_or0);
  fa fa_h_s_dadda_pg_rca32_fa485_out(h_s_dadda_pg_rca32_fa477_xor1[0], h_s_dadda_pg_rca32_fa478_xor1[0], h_s_dadda_pg_rca32_fa479_xor1[0], h_s_dadda_pg_rca32_fa485_xor1, h_s_dadda_pg_rca32_fa485_or0);
  fa fa_h_s_dadda_pg_rca32_fa486_out(h_s_dadda_pg_rca32_fa485_or0[0], h_s_dadda_pg_rca32_fa484_or0[0], h_s_dadda_pg_rca32_fa483_or0[0], h_s_dadda_pg_rca32_fa486_xor1, h_s_dadda_pg_rca32_fa486_or0);
  fa fa_h_s_dadda_pg_rca32_fa487_out(h_s_dadda_pg_rca32_fa482_or0[0], h_s_dadda_pg_rca32_fa481_or0[0], h_s_dadda_pg_rca32_fa480_or0[0], h_s_dadda_pg_rca32_fa487_xor1, h_s_dadda_pg_rca32_fa487_or0);
  fa fa_h_s_dadda_pg_rca32_fa488_out(h_s_dadda_pg_rca32_fa479_or0[0], h_s_dadda_pg_rca32_fa478_or0[0], h_s_dadda_pg_rca32_fa477_or0[0], h_s_dadda_pg_rca32_fa488_xor1, h_s_dadda_pg_rca32_fa488_or0);
  fa fa_h_s_dadda_pg_rca32_fa489_out(h_s_dadda_pg_rca32_fa476_or0[0], h_s_dadda_pg_rca32_fa475_or0[0], h_s_dadda_pg_rca32_fa474_or0[0], h_s_dadda_pg_rca32_fa489_xor1, h_s_dadda_pg_rca32_fa489_or0);
  fa fa_h_s_dadda_pg_rca32_fa490_out(h_s_dadda_pg_rca32_fa473_or0[0], h_s_dadda_pg_rca32_fa472_or0[0], h_s_dadda_pg_rca32_fa471_or0[0], h_s_dadda_pg_rca32_fa490_xor1, h_s_dadda_pg_rca32_fa490_or0);
  fa fa_h_s_dadda_pg_rca32_fa491_out(h_s_dadda_pg_rca32_fa470_or0[0], h_s_dadda_pg_rca32_fa469_or0[0], h_s_dadda_pg_rca32_fa468_or0[0], h_s_dadda_pg_rca32_fa491_xor1, h_s_dadda_pg_rca32_fa491_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_8(a[31], b[8], h_s_dadda_pg_rca32_nand_31_8);
  fa fa_h_s_dadda_pg_rca32_fa492_out(h_s_dadda_pg_rca32_fa467_or0[0], h_s_dadda_pg_rca32_fa466_or0[0], h_s_dadda_pg_rca32_nand_31_8[0], h_s_dadda_pg_rca32_fa492_xor1, h_s_dadda_pg_rca32_fa492_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_9(a[30], b[9], h_s_dadda_pg_rca32_and_30_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_10(a[29], b[10], h_s_dadda_pg_rca32_and_29_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_11(a[28], b[11], h_s_dadda_pg_rca32_and_28_11);
  fa fa_h_s_dadda_pg_rca32_fa493_out(h_s_dadda_pg_rca32_and_30_9[0], h_s_dadda_pg_rca32_and_29_10[0], h_s_dadda_pg_rca32_and_28_11[0], h_s_dadda_pg_rca32_fa493_xor1, h_s_dadda_pg_rca32_fa493_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_12(a[27], b[12], h_s_dadda_pg_rca32_and_27_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_13(a[26], b[13], h_s_dadda_pg_rca32_and_26_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_14(a[25], b[14], h_s_dadda_pg_rca32_and_25_14);
  fa fa_h_s_dadda_pg_rca32_fa494_out(h_s_dadda_pg_rca32_and_27_12[0], h_s_dadda_pg_rca32_and_26_13[0], h_s_dadda_pg_rca32_and_25_14[0], h_s_dadda_pg_rca32_fa494_xor1, h_s_dadda_pg_rca32_fa494_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_15(a[24], b[15], h_s_dadda_pg_rca32_and_24_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_16(a[23], b[16], h_s_dadda_pg_rca32_and_23_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_17(a[22], b[17], h_s_dadda_pg_rca32_and_22_17);
  fa fa_h_s_dadda_pg_rca32_fa495_out(h_s_dadda_pg_rca32_and_24_15[0], h_s_dadda_pg_rca32_and_23_16[0], h_s_dadda_pg_rca32_and_22_17[0], h_s_dadda_pg_rca32_fa495_xor1, h_s_dadda_pg_rca32_fa495_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_18(a[21], b[18], h_s_dadda_pg_rca32_and_21_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_19(a[20], b[19], h_s_dadda_pg_rca32_and_20_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_20(a[19], b[20], h_s_dadda_pg_rca32_and_19_20);
  fa fa_h_s_dadda_pg_rca32_fa496_out(h_s_dadda_pg_rca32_and_21_18[0], h_s_dadda_pg_rca32_and_20_19[0], h_s_dadda_pg_rca32_and_19_20[0], h_s_dadda_pg_rca32_fa496_xor1, h_s_dadda_pg_rca32_fa496_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_21(a[18], b[21], h_s_dadda_pg_rca32_and_18_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_22(a[17], b[22], h_s_dadda_pg_rca32_and_17_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_23(a[16], b[23], h_s_dadda_pg_rca32_and_16_23);
  fa fa_h_s_dadda_pg_rca32_fa497_out(h_s_dadda_pg_rca32_and_18_21[0], h_s_dadda_pg_rca32_and_17_22[0], h_s_dadda_pg_rca32_and_16_23[0], h_s_dadda_pg_rca32_fa497_xor1, h_s_dadda_pg_rca32_fa497_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_24(a[15], b[24], h_s_dadda_pg_rca32_and_15_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_25(a[14], b[25], h_s_dadda_pg_rca32_and_14_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_26(a[13], b[26], h_s_dadda_pg_rca32_and_13_26);
  fa fa_h_s_dadda_pg_rca32_fa498_out(h_s_dadda_pg_rca32_and_15_24[0], h_s_dadda_pg_rca32_and_14_25[0], h_s_dadda_pg_rca32_and_13_26[0], h_s_dadda_pg_rca32_fa498_xor1, h_s_dadda_pg_rca32_fa498_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_27(a[12], b[27], h_s_dadda_pg_rca32_and_12_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_28(a[11], b[28], h_s_dadda_pg_rca32_and_11_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_29(a[10], b[29], h_s_dadda_pg_rca32_and_10_29);
  fa fa_h_s_dadda_pg_rca32_fa499_out(h_s_dadda_pg_rca32_and_12_27[0], h_s_dadda_pg_rca32_and_11_28[0], h_s_dadda_pg_rca32_and_10_29[0], h_s_dadda_pg_rca32_fa499_xor1, h_s_dadda_pg_rca32_fa499_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_9_30(a[9], b[30], h_s_dadda_pg_rca32_and_9_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_8_31(a[8], b[31], h_s_dadda_pg_rca32_nand_8_31);
  fa fa_h_s_dadda_pg_rca32_fa500_out(h_s_dadda_pg_rca32_and_9_30[0], h_s_dadda_pg_rca32_nand_8_31[0], h_s_dadda_pg_rca32_fa486_xor1[0], h_s_dadda_pg_rca32_fa500_xor1, h_s_dadda_pg_rca32_fa500_or0);
  fa fa_h_s_dadda_pg_rca32_fa501_out(h_s_dadda_pg_rca32_fa487_xor1[0], h_s_dadda_pg_rca32_fa488_xor1[0], h_s_dadda_pg_rca32_fa489_xor1[0], h_s_dadda_pg_rca32_fa501_xor1, h_s_dadda_pg_rca32_fa501_or0);
  fa fa_h_s_dadda_pg_rca32_fa502_out(h_s_dadda_pg_rca32_fa490_xor1[0], h_s_dadda_pg_rca32_fa491_xor1[0], h_s_dadda_pg_rca32_fa492_xor1[0], h_s_dadda_pg_rca32_fa502_xor1, h_s_dadda_pg_rca32_fa502_or0);
  fa fa_h_s_dadda_pg_rca32_fa503_out(h_s_dadda_pg_rca32_fa493_xor1[0], h_s_dadda_pg_rca32_fa494_xor1[0], h_s_dadda_pg_rca32_fa495_xor1[0], h_s_dadda_pg_rca32_fa503_xor1, h_s_dadda_pg_rca32_fa503_or0);
  fa fa_h_s_dadda_pg_rca32_fa504_out(h_s_dadda_pg_rca32_fa496_xor1[0], h_s_dadda_pg_rca32_fa497_xor1[0], h_s_dadda_pg_rca32_fa498_xor1[0], h_s_dadda_pg_rca32_fa504_xor1, h_s_dadda_pg_rca32_fa504_or0);
  fa fa_h_s_dadda_pg_rca32_fa505_out(h_s_dadda_pg_rca32_fa504_or0[0], h_s_dadda_pg_rca32_fa503_or0[0], h_s_dadda_pg_rca32_fa502_or0[0], h_s_dadda_pg_rca32_fa505_xor1, h_s_dadda_pg_rca32_fa505_or0);
  fa fa_h_s_dadda_pg_rca32_fa506_out(h_s_dadda_pg_rca32_fa501_or0[0], h_s_dadda_pg_rca32_fa500_or0[0], h_s_dadda_pg_rca32_fa499_or0[0], h_s_dadda_pg_rca32_fa506_xor1, h_s_dadda_pg_rca32_fa506_or0);
  fa fa_h_s_dadda_pg_rca32_fa507_out(h_s_dadda_pg_rca32_fa498_or0[0], h_s_dadda_pg_rca32_fa497_or0[0], h_s_dadda_pg_rca32_fa496_or0[0], h_s_dadda_pg_rca32_fa507_xor1, h_s_dadda_pg_rca32_fa507_or0);
  fa fa_h_s_dadda_pg_rca32_fa508_out(h_s_dadda_pg_rca32_fa495_or0[0], h_s_dadda_pg_rca32_fa494_or0[0], h_s_dadda_pg_rca32_fa493_or0[0], h_s_dadda_pg_rca32_fa508_xor1, h_s_dadda_pg_rca32_fa508_or0);
  fa fa_h_s_dadda_pg_rca32_fa509_out(h_s_dadda_pg_rca32_fa492_or0[0], h_s_dadda_pg_rca32_fa491_or0[0], h_s_dadda_pg_rca32_fa490_or0[0], h_s_dadda_pg_rca32_fa509_xor1, h_s_dadda_pg_rca32_fa509_or0);
  fa fa_h_s_dadda_pg_rca32_fa510_out(h_s_dadda_pg_rca32_fa489_or0[0], h_s_dadda_pg_rca32_fa488_or0[0], h_s_dadda_pg_rca32_fa487_or0[0], h_s_dadda_pg_rca32_fa510_xor1, h_s_dadda_pg_rca32_fa510_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_9(a[31], b[9], h_s_dadda_pg_rca32_nand_31_9);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_10(a[30], b[10], h_s_dadda_pg_rca32_and_30_10);
  fa fa_h_s_dadda_pg_rca32_fa511_out(h_s_dadda_pg_rca32_fa486_or0[0], h_s_dadda_pg_rca32_nand_31_9[0], h_s_dadda_pg_rca32_and_30_10[0], h_s_dadda_pg_rca32_fa511_xor1, h_s_dadda_pg_rca32_fa511_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_11(a[29], b[11], h_s_dadda_pg_rca32_and_29_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_12(a[28], b[12], h_s_dadda_pg_rca32_and_28_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_13(a[27], b[13], h_s_dadda_pg_rca32_and_27_13);
  fa fa_h_s_dadda_pg_rca32_fa512_out(h_s_dadda_pg_rca32_and_29_11[0], h_s_dadda_pg_rca32_and_28_12[0], h_s_dadda_pg_rca32_and_27_13[0], h_s_dadda_pg_rca32_fa512_xor1, h_s_dadda_pg_rca32_fa512_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_14(a[26], b[14], h_s_dadda_pg_rca32_and_26_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_15(a[25], b[15], h_s_dadda_pg_rca32_and_25_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_16(a[24], b[16], h_s_dadda_pg_rca32_and_24_16);
  fa fa_h_s_dadda_pg_rca32_fa513_out(h_s_dadda_pg_rca32_and_26_14[0], h_s_dadda_pg_rca32_and_25_15[0], h_s_dadda_pg_rca32_and_24_16[0], h_s_dadda_pg_rca32_fa513_xor1, h_s_dadda_pg_rca32_fa513_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_17(a[23], b[17], h_s_dadda_pg_rca32_and_23_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_18(a[22], b[18], h_s_dadda_pg_rca32_and_22_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_19(a[21], b[19], h_s_dadda_pg_rca32_and_21_19);
  fa fa_h_s_dadda_pg_rca32_fa514_out(h_s_dadda_pg_rca32_and_23_17[0], h_s_dadda_pg_rca32_and_22_18[0], h_s_dadda_pg_rca32_and_21_19[0], h_s_dadda_pg_rca32_fa514_xor1, h_s_dadda_pg_rca32_fa514_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_20(a[20], b[20], h_s_dadda_pg_rca32_and_20_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_21(a[19], b[21], h_s_dadda_pg_rca32_and_19_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_22(a[18], b[22], h_s_dadda_pg_rca32_and_18_22);
  fa fa_h_s_dadda_pg_rca32_fa515_out(h_s_dadda_pg_rca32_and_20_20[0], h_s_dadda_pg_rca32_and_19_21[0], h_s_dadda_pg_rca32_and_18_22[0], h_s_dadda_pg_rca32_fa515_xor1, h_s_dadda_pg_rca32_fa515_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_23(a[17], b[23], h_s_dadda_pg_rca32_and_17_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_24(a[16], b[24], h_s_dadda_pg_rca32_and_16_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_25(a[15], b[25], h_s_dadda_pg_rca32_and_15_25);
  fa fa_h_s_dadda_pg_rca32_fa516_out(h_s_dadda_pg_rca32_and_17_23[0], h_s_dadda_pg_rca32_and_16_24[0], h_s_dadda_pg_rca32_and_15_25[0], h_s_dadda_pg_rca32_fa516_xor1, h_s_dadda_pg_rca32_fa516_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_26(a[14], b[26], h_s_dadda_pg_rca32_and_14_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_27(a[13], b[27], h_s_dadda_pg_rca32_and_13_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_28(a[12], b[28], h_s_dadda_pg_rca32_and_12_28);
  fa fa_h_s_dadda_pg_rca32_fa517_out(h_s_dadda_pg_rca32_and_14_26[0], h_s_dadda_pg_rca32_and_13_27[0], h_s_dadda_pg_rca32_and_12_28[0], h_s_dadda_pg_rca32_fa517_xor1, h_s_dadda_pg_rca32_fa517_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_29(a[11], b[29], h_s_dadda_pg_rca32_and_11_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_10_30(a[10], b[30], h_s_dadda_pg_rca32_and_10_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_9_31(a[9], b[31], h_s_dadda_pg_rca32_nand_9_31);
  fa fa_h_s_dadda_pg_rca32_fa518_out(h_s_dadda_pg_rca32_and_11_29[0], h_s_dadda_pg_rca32_and_10_30[0], h_s_dadda_pg_rca32_nand_9_31[0], h_s_dadda_pg_rca32_fa518_xor1, h_s_dadda_pg_rca32_fa518_or0);
  fa fa_h_s_dadda_pg_rca32_fa519_out(h_s_dadda_pg_rca32_fa505_xor1[0], h_s_dadda_pg_rca32_fa506_xor1[0], h_s_dadda_pg_rca32_fa507_xor1[0], h_s_dadda_pg_rca32_fa519_xor1, h_s_dadda_pg_rca32_fa519_or0);
  fa fa_h_s_dadda_pg_rca32_fa520_out(h_s_dadda_pg_rca32_fa508_xor1[0], h_s_dadda_pg_rca32_fa509_xor1[0], h_s_dadda_pg_rca32_fa510_xor1[0], h_s_dadda_pg_rca32_fa520_xor1, h_s_dadda_pg_rca32_fa520_or0);
  fa fa_h_s_dadda_pg_rca32_fa521_out(h_s_dadda_pg_rca32_fa511_xor1[0], h_s_dadda_pg_rca32_fa512_xor1[0], h_s_dadda_pg_rca32_fa513_xor1[0], h_s_dadda_pg_rca32_fa521_xor1, h_s_dadda_pg_rca32_fa521_or0);
  fa fa_h_s_dadda_pg_rca32_fa522_out(h_s_dadda_pg_rca32_fa514_xor1[0], h_s_dadda_pg_rca32_fa515_xor1[0], h_s_dadda_pg_rca32_fa516_xor1[0], h_s_dadda_pg_rca32_fa522_xor1, h_s_dadda_pg_rca32_fa522_or0);
  fa fa_h_s_dadda_pg_rca32_fa523_out(h_s_dadda_pg_rca32_fa522_or0[0], h_s_dadda_pg_rca32_fa521_or0[0], h_s_dadda_pg_rca32_fa520_or0[0], h_s_dadda_pg_rca32_fa523_xor1, h_s_dadda_pg_rca32_fa523_or0);
  fa fa_h_s_dadda_pg_rca32_fa524_out(h_s_dadda_pg_rca32_fa519_or0[0], h_s_dadda_pg_rca32_fa518_or0[0], h_s_dadda_pg_rca32_fa517_or0[0], h_s_dadda_pg_rca32_fa524_xor1, h_s_dadda_pg_rca32_fa524_or0);
  fa fa_h_s_dadda_pg_rca32_fa525_out(h_s_dadda_pg_rca32_fa516_or0[0], h_s_dadda_pg_rca32_fa515_or0[0], h_s_dadda_pg_rca32_fa514_or0[0], h_s_dadda_pg_rca32_fa525_xor1, h_s_dadda_pg_rca32_fa525_or0);
  fa fa_h_s_dadda_pg_rca32_fa526_out(h_s_dadda_pg_rca32_fa513_or0[0], h_s_dadda_pg_rca32_fa512_or0[0], h_s_dadda_pg_rca32_fa511_or0[0], h_s_dadda_pg_rca32_fa526_xor1, h_s_dadda_pg_rca32_fa526_or0);
  fa fa_h_s_dadda_pg_rca32_fa527_out(h_s_dadda_pg_rca32_fa510_or0[0], h_s_dadda_pg_rca32_fa509_or0[0], h_s_dadda_pg_rca32_fa508_or0[0], h_s_dadda_pg_rca32_fa527_xor1, h_s_dadda_pg_rca32_fa527_or0);
  fa fa_h_s_dadda_pg_rca32_fa528_out(h_s_dadda_pg_rca32_fa507_or0[0], h_s_dadda_pg_rca32_fa506_or0[0], h_s_dadda_pg_rca32_fa505_or0[0], h_s_dadda_pg_rca32_fa528_xor1, h_s_dadda_pg_rca32_fa528_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_10(a[31], b[10], h_s_dadda_pg_rca32_nand_31_10);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_11(a[30], b[11], h_s_dadda_pg_rca32_and_30_11);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_12(a[29], b[12], h_s_dadda_pg_rca32_and_29_12);
  fa fa_h_s_dadda_pg_rca32_fa529_out(h_s_dadda_pg_rca32_nand_31_10[0], h_s_dadda_pg_rca32_and_30_11[0], h_s_dadda_pg_rca32_and_29_12[0], h_s_dadda_pg_rca32_fa529_xor1, h_s_dadda_pg_rca32_fa529_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_13(a[28], b[13], h_s_dadda_pg_rca32_and_28_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_14(a[27], b[14], h_s_dadda_pg_rca32_and_27_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_15(a[26], b[15], h_s_dadda_pg_rca32_and_26_15);
  fa fa_h_s_dadda_pg_rca32_fa530_out(h_s_dadda_pg_rca32_and_28_13[0], h_s_dadda_pg_rca32_and_27_14[0], h_s_dadda_pg_rca32_and_26_15[0], h_s_dadda_pg_rca32_fa530_xor1, h_s_dadda_pg_rca32_fa530_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_16(a[25], b[16], h_s_dadda_pg_rca32_and_25_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_17(a[24], b[17], h_s_dadda_pg_rca32_and_24_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_18(a[23], b[18], h_s_dadda_pg_rca32_and_23_18);
  fa fa_h_s_dadda_pg_rca32_fa531_out(h_s_dadda_pg_rca32_and_25_16[0], h_s_dadda_pg_rca32_and_24_17[0], h_s_dadda_pg_rca32_and_23_18[0], h_s_dadda_pg_rca32_fa531_xor1, h_s_dadda_pg_rca32_fa531_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_19(a[22], b[19], h_s_dadda_pg_rca32_and_22_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_20(a[21], b[20], h_s_dadda_pg_rca32_and_21_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_21(a[20], b[21], h_s_dadda_pg_rca32_and_20_21);
  fa fa_h_s_dadda_pg_rca32_fa532_out(h_s_dadda_pg_rca32_and_22_19[0], h_s_dadda_pg_rca32_and_21_20[0], h_s_dadda_pg_rca32_and_20_21[0], h_s_dadda_pg_rca32_fa532_xor1, h_s_dadda_pg_rca32_fa532_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_22(a[19], b[22], h_s_dadda_pg_rca32_and_19_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_23(a[18], b[23], h_s_dadda_pg_rca32_and_18_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_24(a[17], b[24], h_s_dadda_pg_rca32_and_17_24);
  fa fa_h_s_dadda_pg_rca32_fa533_out(h_s_dadda_pg_rca32_and_19_22[0], h_s_dadda_pg_rca32_and_18_23[0], h_s_dadda_pg_rca32_and_17_24[0], h_s_dadda_pg_rca32_fa533_xor1, h_s_dadda_pg_rca32_fa533_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_25(a[16], b[25], h_s_dadda_pg_rca32_and_16_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_26(a[15], b[26], h_s_dadda_pg_rca32_and_15_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_27(a[14], b[27], h_s_dadda_pg_rca32_and_14_27);
  fa fa_h_s_dadda_pg_rca32_fa534_out(h_s_dadda_pg_rca32_and_16_25[0], h_s_dadda_pg_rca32_and_15_26[0], h_s_dadda_pg_rca32_and_14_27[0], h_s_dadda_pg_rca32_fa534_xor1, h_s_dadda_pg_rca32_fa534_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_28(a[13], b[28], h_s_dadda_pg_rca32_and_13_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_29(a[12], b[29], h_s_dadda_pg_rca32_and_12_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_11_30(a[11], b[30], h_s_dadda_pg_rca32_and_11_30);
  fa fa_h_s_dadda_pg_rca32_fa535_out(h_s_dadda_pg_rca32_and_13_28[0], h_s_dadda_pg_rca32_and_12_29[0], h_s_dadda_pg_rca32_and_11_30[0], h_s_dadda_pg_rca32_fa535_xor1, h_s_dadda_pg_rca32_fa535_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_10_31(a[10], b[31], h_s_dadda_pg_rca32_nand_10_31);
  fa fa_h_s_dadda_pg_rca32_fa536_out(h_s_dadda_pg_rca32_nand_10_31[0], h_s_dadda_pg_rca32_fa523_xor1[0], h_s_dadda_pg_rca32_fa524_xor1[0], h_s_dadda_pg_rca32_fa536_xor1, h_s_dadda_pg_rca32_fa536_or0);
  fa fa_h_s_dadda_pg_rca32_fa537_out(h_s_dadda_pg_rca32_fa525_xor1[0], h_s_dadda_pg_rca32_fa526_xor1[0], h_s_dadda_pg_rca32_fa527_xor1[0], h_s_dadda_pg_rca32_fa537_xor1, h_s_dadda_pg_rca32_fa537_or0);
  fa fa_h_s_dadda_pg_rca32_fa538_out(h_s_dadda_pg_rca32_fa528_xor1[0], h_s_dadda_pg_rca32_fa529_xor1[0], h_s_dadda_pg_rca32_fa530_xor1[0], h_s_dadda_pg_rca32_fa538_xor1, h_s_dadda_pg_rca32_fa538_or0);
  fa fa_h_s_dadda_pg_rca32_fa539_out(h_s_dadda_pg_rca32_fa531_xor1[0], h_s_dadda_pg_rca32_fa532_xor1[0], h_s_dadda_pg_rca32_fa533_xor1[0], h_s_dadda_pg_rca32_fa539_xor1, h_s_dadda_pg_rca32_fa539_or0);
  fa fa_h_s_dadda_pg_rca32_fa540_out(h_s_dadda_pg_rca32_fa539_or0[0], h_s_dadda_pg_rca32_fa538_or0[0], h_s_dadda_pg_rca32_fa537_or0[0], h_s_dadda_pg_rca32_fa540_xor1, h_s_dadda_pg_rca32_fa540_or0);
  fa fa_h_s_dadda_pg_rca32_fa541_out(h_s_dadda_pg_rca32_fa536_or0[0], h_s_dadda_pg_rca32_fa535_or0[0], h_s_dadda_pg_rca32_fa534_or0[0], h_s_dadda_pg_rca32_fa541_xor1, h_s_dadda_pg_rca32_fa541_or0);
  fa fa_h_s_dadda_pg_rca32_fa542_out(h_s_dadda_pg_rca32_fa533_or0[0], h_s_dadda_pg_rca32_fa532_or0[0], h_s_dadda_pg_rca32_fa531_or0[0], h_s_dadda_pg_rca32_fa542_xor1, h_s_dadda_pg_rca32_fa542_or0);
  fa fa_h_s_dadda_pg_rca32_fa543_out(h_s_dadda_pg_rca32_fa530_or0[0], h_s_dadda_pg_rca32_fa529_or0[0], h_s_dadda_pg_rca32_fa528_or0[0], h_s_dadda_pg_rca32_fa543_xor1, h_s_dadda_pg_rca32_fa543_or0);
  fa fa_h_s_dadda_pg_rca32_fa544_out(h_s_dadda_pg_rca32_fa527_or0[0], h_s_dadda_pg_rca32_fa526_or0[0], h_s_dadda_pg_rca32_fa525_or0[0], h_s_dadda_pg_rca32_fa544_xor1, h_s_dadda_pg_rca32_fa544_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_11(a[31], b[11], h_s_dadda_pg_rca32_nand_31_11);
  fa fa_h_s_dadda_pg_rca32_fa545_out(h_s_dadda_pg_rca32_fa524_or0[0], h_s_dadda_pg_rca32_fa523_or0[0], h_s_dadda_pg_rca32_nand_31_11[0], h_s_dadda_pg_rca32_fa545_xor1, h_s_dadda_pg_rca32_fa545_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_12(a[30], b[12], h_s_dadda_pg_rca32_and_30_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_13(a[29], b[13], h_s_dadda_pg_rca32_and_29_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_14(a[28], b[14], h_s_dadda_pg_rca32_and_28_14);
  fa fa_h_s_dadda_pg_rca32_fa546_out(h_s_dadda_pg_rca32_and_30_12[0], h_s_dadda_pg_rca32_and_29_13[0], h_s_dadda_pg_rca32_and_28_14[0], h_s_dadda_pg_rca32_fa546_xor1, h_s_dadda_pg_rca32_fa546_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_15(a[27], b[15], h_s_dadda_pg_rca32_and_27_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_16(a[26], b[16], h_s_dadda_pg_rca32_and_26_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_17(a[25], b[17], h_s_dadda_pg_rca32_and_25_17);
  fa fa_h_s_dadda_pg_rca32_fa547_out(h_s_dadda_pg_rca32_and_27_15[0], h_s_dadda_pg_rca32_and_26_16[0], h_s_dadda_pg_rca32_and_25_17[0], h_s_dadda_pg_rca32_fa547_xor1, h_s_dadda_pg_rca32_fa547_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_18(a[24], b[18], h_s_dadda_pg_rca32_and_24_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_19(a[23], b[19], h_s_dadda_pg_rca32_and_23_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_20(a[22], b[20], h_s_dadda_pg_rca32_and_22_20);
  fa fa_h_s_dadda_pg_rca32_fa548_out(h_s_dadda_pg_rca32_and_24_18[0], h_s_dadda_pg_rca32_and_23_19[0], h_s_dadda_pg_rca32_and_22_20[0], h_s_dadda_pg_rca32_fa548_xor1, h_s_dadda_pg_rca32_fa548_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_21(a[21], b[21], h_s_dadda_pg_rca32_and_21_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_22(a[20], b[22], h_s_dadda_pg_rca32_and_20_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_23(a[19], b[23], h_s_dadda_pg_rca32_and_19_23);
  fa fa_h_s_dadda_pg_rca32_fa549_out(h_s_dadda_pg_rca32_and_21_21[0], h_s_dadda_pg_rca32_and_20_22[0], h_s_dadda_pg_rca32_and_19_23[0], h_s_dadda_pg_rca32_fa549_xor1, h_s_dadda_pg_rca32_fa549_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_24(a[18], b[24], h_s_dadda_pg_rca32_and_18_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_25(a[17], b[25], h_s_dadda_pg_rca32_and_17_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_26(a[16], b[26], h_s_dadda_pg_rca32_and_16_26);
  fa fa_h_s_dadda_pg_rca32_fa550_out(h_s_dadda_pg_rca32_and_18_24[0], h_s_dadda_pg_rca32_and_17_25[0], h_s_dadda_pg_rca32_and_16_26[0], h_s_dadda_pg_rca32_fa550_xor1, h_s_dadda_pg_rca32_fa550_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_27(a[15], b[27], h_s_dadda_pg_rca32_and_15_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_28(a[14], b[28], h_s_dadda_pg_rca32_and_14_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_29(a[13], b[29], h_s_dadda_pg_rca32_and_13_29);
  fa fa_h_s_dadda_pg_rca32_fa551_out(h_s_dadda_pg_rca32_and_15_27[0], h_s_dadda_pg_rca32_and_14_28[0], h_s_dadda_pg_rca32_and_13_29[0], h_s_dadda_pg_rca32_fa551_xor1, h_s_dadda_pg_rca32_fa551_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_12_30(a[12], b[30], h_s_dadda_pg_rca32_and_12_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_11_31(a[11], b[31], h_s_dadda_pg_rca32_nand_11_31);
  fa fa_h_s_dadda_pg_rca32_fa552_out(h_s_dadda_pg_rca32_and_12_30[0], h_s_dadda_pg_rca32_nand_11_31[0], h_s_dadda_pg_rca32_fa540_xor1[0], h_s_dadda_pg_rca32_fa552_xor1, h_s_dadda_pg_rca32_fa552_or0);
  fa fa_h_s_dadda_pg_rca32_fa553_out(h_s_dadda_pg_rca32_fa541_xor1[0], h_s_dadda_pg_rca32_fa542_xor1[0], h_s_dadda_pg_rca32_fa543_xor1[0], h_s_dadda_pg_rca32_fa553_xor1, h_s_dadda_pg_rca32_fa553_or0);
  fa fa_h_s_dadda_pg_rca32_fa554_out(h_s_dadda_pg_rca32_fa544_xor1[0], h_s_dadda_pg_rca32_fa545_xor1[0], h_s_dadda_pg_rca32_fa546_xor1[0], h_s_dadda_pg_rca32_fa554_xor1, h_s_dadda_pg_rca32_fa554_or0);
  fa fa_h_s_dadda_pg_rca32_fa555_out(h_s_dadda_pg_rca32_fa547_xor1[0], h_s_dadda_pg_rca32_fa548_xor1[0], h_s_dadda_pg_rca32_fa549_xor1[0], h_s_dadda_pg_rca32_fa555_xor1, h_s_dadda_pg_rca32_fa555_or0);
  fa fa_h_s_dadda_pg_rca32_fa556_out(h_s_dadda_pg_rca32_fa555_or0[0], h_s_dadda_pg_rca32_fa554_or0[0], h_s_dadda_pg_rca32_fa553_or0[0], h_s_dadda_pg_rca32_fa556_xor1, h_s_dadda_pg_rca32_fa556_or0);
  fa fa_h_s_dadda_pg_rca32_fa557_out(h_s_dadda_pg_rca32_fa552_or0[0], h_s_dadda_pg_rca32_fa551_or0[0], h_s_dadda_pg_rca32_fa550_or0[0], h_s_dadda_pg_rca32_fa557_xor1, h_s_dadda_pg_rca32_fa557_or0);
  fa fa_h_s_dadda_pg_rca32_fa558_out(h_s_dadda_pg_rca32_fa549_or0[0], h_s_dadda_pg_rca32_fa548_or0[0], h_s_dadda_pg_rca32_fa547_or0[0], h_s_dadda_pg_rca32_fa558_xor1, h_s_dadda_pg_rca32_fa558_or0);
  fa fa_h_s_dadda_pg_rca32_fa559_out(h_s_dadda_pg_rca32_fa546_or0[0], h_s_dadda_pg_rca32_fa545_or0[0], h_s_dadda_pg_rca32_fa544_or0[0], h_s_dadda_pg_rca32_fa559_xor1, h_s_dadda_pg_rca32_fa559_or0);
  fa fa_h_s_dadda_pg_rca32_fa560_out(h_s_dadda_pg_rca32_fa543_or0[0], h_s_dadda_pg_rca32_fa542_or0[0], h_s_dadda_pg_rca32_fa541_or0[0], h_s_dadda_pg_rca32_fa560_xor1, h_s_dadda_pg_rca32_fa560_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_12(a[31], b[12], h_s_dadda_pg_rca32_nand_31_12);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_13(a[30], b[13], h_s_dadda_pg_rca32_and_30_13);
  fa fa_h_s_dadda_pg_rca32_fa561_out(h_s_dadda_pg_rca32_fa540_or0[0], h_s_dadda_pg_rca32_nand_31_12[0], h_s_dadda_pg_rca32_and_30_13[0], h_s_dadda_pg_rca32_fa561_xor1, h_s_dadda_pg_rca32_fa561_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_14(a[29], b[14], h_s_dadda_pg_rca32_and_29_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_15(a[28], b[15], h_s_dadda_pg_rca32_and_28_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_16(a[27], b[16], h_s_dadda_pg_rca32_and_27_16);
  fa fa_h_s_dadda_pg_rca32_fa562_out(h_s_dadda_pg_rca32_and_29_14[0], h_s_dadda_pg_rca32_and_28_15[0], h_s_dadda_pg_rca32_and_27_16[0], h_s_dadda_pg_rca32_fa562_xor1, h_s_dadda_pg_rca32_fa562_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_17(a[26], b[17], h_s_dadda_pg_rca32_and_26_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_18(a[25], b[18], h_s_dadda_pg_rca32_and_25_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_19(a[24], b[19], h_s_dadda_pg_rca32_and_24_19);
  fa fa_h_s_dadda_pg_rca32_fa563_out(h_s_dadda_pg_rca32_and_26_17[0], h_s_dadda_pg_rca32_and_25_18[0], h_s_dadda_pg_rca32_and_24_19[0], h_s_dadda_pg_rca32_fa563_xor1, h_s_dadda_pg_rca32_fa563_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_20(a[23], b[20], h_s_dadda_pg_rca32_and_23_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_21(a[22], b[21], h_s_dadda_pg_rca32_and_22_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_22(a[21], b[22], h_s_dadda_pg_rca32_and_21_22);
  fa fa_h_s_dadda_pg_rca32_fa564_out(h_s_dadda_pg_rca32_and_23_20[0], h_s_dadda_pg_rca32_and_22_21[0], h_s_dadda_pg_rca32_and_21_22[0], h_s_dadda_pg_rca32_fa564_xor1, h_s_dadda_pg_rca32_fa564_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_23(a[20], b[23], h_s_dadda_pg_rca32_and_20_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_24(a[19], b[24], h_s_dadda_pg_rca32_and_19_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_25(a[18], b[25], h_s_dadda_pg_rca32_and_18_25);
  fa fa_h_s_dadda_pg_rca32_fa565_out(h_s_dadda_pg_rca32_and_20_23[0], h_s_dadda_pg_rca32_and_19_24[0], h_s_dadda_pg_rca32_and_18_25[0], h_s_dadda_pg_rca32_fa565_xor1, h_s_dadda_pg_rca32_fa565_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_26(a[17], b[26], h_s_dadda_pg_rca32_and_17_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_27(a[16], b[27], h_s_dadda_pg_rca32_and_16_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_28(a[15], b[28], h_s_dadda_pg_rca32_and_15_28);
  fa fa_h_s_dadda_pg_rca32_fa566_out(h_s_dadda_pg_rca32_and_17_26[0], h_s_dadda_pg_rca32_and_16_27[0], h_s_dadda_pg_rca32_and_15_28[0], h_s_dadda_pg_rca32_fa566_xor1, h_s_dadda_pg_rca32_fa566_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_29(a[14], b[29], h_s_dadda_pg_rca32_and_14_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_13_30(a[13], b[30], h_s_dadda_pg_rca32_and_13_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_12_31(a[12], b[31], h_s_dadda_pg_rca32_nand_12_31);
  fa fa_h_s_dadda_pg_rca32_fa567_out(h_s_dadda_pg_rca32_and_14_29[0], h_s_dadda_pg_rca32_and_13_30[0], h_s_dadda_pg_rca32_nand_12_31[0], h_s_dadda_pg_rca32_fa567_xor1, h_s_dadda_pg_rca32_fa567_or0);
  fa fa_h_s_dadda_pg_rca32_fa568_out(h_s_dadda_pg_rca32_fa556_xor1[0], h_s_dadda_pg_rca32_fa557_xor1[0], h_s_dadda_pg_rca32_fa558_xor1[0], h_s_dadda_pg_rca32_fa568_xor1, h_s_dadda_pg_rca32_fa568_or0);
  fa fa_h_s_dadda_pg_rca32_fa569_out(h_s_dadda_pg_rca32_fa559_xor1[0], h_s_dadda_pg_rca32_fa560_xor1[0], h_s_dadda_pg_rca32_fa561_xor1[0], h_s_dadda_pg_rca32_fa569_xor1, h_s_dadda_pg_rca32_fa569_or0);
  fa fa_h_s_dadda_pg_rca32_fa570_out(h_s_dadda_pg_rca32_fa562_xor1[0], h_s_dadda_pg_rca32_fa563_xor1[0], h_s_dadda_pg_rca32_fa564_xor1[0], h_s_dadda_pg_rca32_fa570_xor1, h_s_dadda_pg_rca32_fa570_or0);
  fa fa_h_s_dadda_pg_rca32_fa571_out(h_s_dadda_pg_rca32_fa570_or0[0], h_s_dadda_pg_rca32_fa569_or0[0], h_s_dadda_pg_rca32_fa568_or0[0], h_s_dadda_pg_rca32_fa571_xor1, h_s_dadda_pg_rca32_fa571_or0);
  fa fa_h_s_dadda_pg_rca32_fa572_out(h_s_dadda_pg_rca32_fa567_or0[0], h_s_dadda_pg_rca32_fa566_or0[0], h_s_dadda_pg_rca32_fa565_or0[0], h_s_dadda_pg_rca32_fa572_xor1, h_s_dadda_pg_rca32_fa572_or0);
  fa fa_h_s_dadda_pg_rca32_fa573_out(h_s_dadda_pg_rca32_fa564_or0[0], h_s_dadda_pg_rca32_fa563_or0[0], h_s_dadda_pg_rca32_fa562_or0[0], h_s_dadda_pg_rca32_fa573_xor1, h_s_dadda_pg_rca32_fa573_or0);
  fa fa_h_s_dadda_pg_rca32_fa574_out(h_s_dadda_pg_rca32_fa561_or0[0], h_s_dadda_pg_rca32_fa560_or0[0], h_s_dadda_pg_rca32_fa559_or0[0], h_s_dadda_pg_rca32_fa574_xor1, h_s_dadda_pg_rca32_fa574_or0);
  fa fa_h_s_dadda_pg_rca32_fa575_out(h_s_dadda_pg_rca32_fa558_or0[0], h_s_dadda_pg_rca32_fa557_or0[0], h_s_dadda_pg_rca32_fa556_or0[0], h_s_dadda_pg_rca32_fa575_xor1, h_s_dadda_pg_rca32_fa575_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_13(a[31], b[13], h_s_dadda_pg_rca32_nand_31_13);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_14(a[30], b[14], h_s_dadda_pg_rca32_and_30_14);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_15(a[29], b[15], h_s_dadda_pg_rca32_and_29_15);
  fa fa_h_s_dadda_pg_rca32_fa576_out(h_s_dadda_pg_rca32_nand_31_13[0], h_s_dadda_pg_rca32_and_30_14[0], h_s_dadda_pg_rca32_and_29_15[0], h_s_dadda_pg_rca32_fa576_xor1, h_s_dadda_pg_rca32_fa576_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_16(a[28], b[16], h_s_dadda_pg_rca32_and_28_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_17(a[27], b[17], h_s_dadda_pg_rca32_and_27_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_18(a[26], b[18], h_s_dadda_pg_rca32_and_26_18);
  fa fa_h_s_dadda_pg_rca32_fa577_out(h_s_dadda_pg_rca32_and_28_16[0], h_s_dadda_pg_rca32_and_27_17[0], h_s_dadda_pg_rca32_and_26_18[0], h_s_dadda_pg_rca32_fa577_xor1, h_s_dadda_pg_rca32_fa577_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_19(a[25], b[19], h_s_dadda_pg_rca32_and_25_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_20(a[24], b[20], h_s_dadda_pg_rca32_and_24_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_21(a[23], b[21], h_s_dadda_pg_rca32_and_23_21);
  fa fa_h_s_dadda_pg_rca32_fa578_out(h_s_dadda_pg_rca32_and_25_19[0], h_s_dadda_pg_rca32_and_24_20[0], h_s_dadda_pg_rca32_and_23_21[0], h_s_dadda_pg_rca32_fa578_xor1, h_s_dadda_pg_rca32_fa578_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_22(a[22], b[22], h_s_dadda_pg_rca32_and_22_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_23(a[21], b[23], h_s_dadda_pg_rca32_and_21_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_24(a[20], b[24], h_s_dadda_pg_rca32_and_20_24);
  fa fa_h_s_dadda_pg_rca32_fa579_out(h_s_dadda_pg_rca32_and_22_22[0], h_s_dadda_pg_rca32_and_21_23[0], h_s_dadda_pg_rca32_and_20_24[0], h_s_dadda_pg_rca32_fa579_xor1, h_s_dadda_pg_rca32_fa579_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_25(a[19], b[25], h_s_dadda_pg_rca32_and_19_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_26(a[18], b[26], h_s_dadda_pg_rca32_and_18_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_27(a[17], b[27], h_s_dadda_pg_rca32_and_17_27);
  fa fa_h_s_dadda_pg_rca32_fa580_out(h_s_dadda_pg_rca32_and_19_25[0], h_s_dadda_pg_rca32_and_18_26[0], h_s_dadda_pg_rca32_and_17_27[0], h_s_dadda_pg_rca32_fa580_xor1, h_s_dadda_pg_rca32_fa580_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_28(a[16], b[28], h_s_dadda_pg_rca32_and_16_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_29(a[15], b[29], h_s_dadda_pg_rca32_and_15_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_14_30(a[14], b[30], h_s_dadda_pg_rca32_and_14_30);
  fa fa_h_s_dadda_pg_rca32_fa581_out(h_s_dadda_pg_rca32_and_16_28[0], h_s_dadda_pg_rca32_and_15_29[0], h_s_dadda_pg_rca32_and_14_30[0], h_s_dadda_pg_rca32_fa581_xor1, h_s_dadda_pg_rca32_fa581_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_13_31(a[13], b[31], h_s_dadda_pg_rca32_nand_13_31);
  fa fa_h_s_dadda_pg_rca32_fa582_out(h_s_dadda_pg_rca32_nand_13_31[0], h_s_dadda_pg_rca32_fa571_xor1[0], h_s_dadda_pg_rca32_fa572_xor1[0], h_s_dadda_pg_rca32_fa582_xor1, h_s_dadda_pg_rca32_fa582_or0);
  fa fa_h_s_dadda_pg_rca32_fa583_out(h_s_dadda_pg_rca32_fa573_xor1[0], h_s_dadda_pg_rca32_fa574_xor1[0], h_s_dadda_pg_rca32_fa575_xor1[0], h_s_dadda_pg_rca32_fa583_xor1, h_s_dadda_pg_rca32_fa583_or0);
  fa fa_h_s_dadda_pg_rca32_fa584_out(h_s_dadda_pg_rca32_fa576_xor1[0], h_s_dadda_pg_rca32_fa577_xor1[0], h_s_dadda_pg_rca32_fa578_xor1[0], h_s_dadda_pg_rca32_fa584_xor1, h_s_dadda_pg_rca32_fa584_or0);
  fa fa_h_s_dadda_pg_rca32_fa585_out(h_s_dadda_pg_rca32_fa584_or0[0], h_s_dadda_pg_rca32_fa583_or0[0], h_s_dadda_pg_rca32_fa582_or0[0], h_s_dadda_pg_rca32_fa585_xor1, h_s_dadda_pg_rca32_fa585_or0);
  fa fa_h_s_dadda_pg_rca32_fa586_out(h_s_dadda_pg_rca32_fa581_or0[0], h_s_dadda_pg_rca32_fa580_or0[0], h_s_dadda_pg_rca32_fa579_or0[0], h_s_dadda_pg_rca32_fa586_xor1, h_s_dadda_pg_rca32_fa586_or0);
  fa fa_h_s_dadda_pg_rca32_fa587_out(h_s_dadda_pg_rca32_fa578_or0[0], h_s_dadda_pg_rca32_fa577_or0[0], h_s_dadda_pg_rca32_fa576_or0[0], h_s_dadda_pg_rca32_fa587_xor1, h_s_dadda_pg_rca32_fa587_or0);
  fa fa_h_s_dadda_pg_rca32_fa588_out(h_s_dadda_pg_rca32_fa575_or0[0], h_s_dadda_pg_rca32_fa574_or0[0], h_s_dadda_pg_rca32_fa573_or0[0], h_s_dadda_pg_rca32_fa588_xor1, h_s_dadda_pg_rca32_fa588_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_14(a[31], b[14], h_s_dadda_pg_rca32_nand_31_14);
  fa fa_h_s_dadda_pg_rca32_fa589_out(h_s_dadda_pg_rca32_fa572_or0[0], h_s_dadda_pg_rca32_fa571_or0[0], h_s_dadda_pg_rca32_nand_31_14[0], h_s_dadda_pg_rca32_fa589_xor1, h_s_dadda_pg_rca32_fa589_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_15(a[30], b[15], h_s_dadda_pg_rca32_and_30_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_16(a[29], b[16], h_s_dadda_pg_rca32_and_29_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_17(a[28], b[17], h_s_dadda_pg_rca32_and_28_17);
  fa fa_h_s_dadda_pg_rca32_fa590_out(h_s_dadda_pg_rca32_and_30_15[0], h_s_dadda_pg_rca32_and_29_16[0], h_s_dadda_pg_rca32_and_28_17[0], h_s_dadda_pg_rca32_fa590_xor1, h_s_dadda_pg_rca32_fa590_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_18(a[27], b[18], h_s_dadda_pg_rca32_and_27_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_19(a[26], b[19], h_s_dadda_pg_rca32_and_26_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_20(a[25], b[20], h_s_dadda_pg_rca32_and_25_20);
  fa fa_h_s_dadda_pg_rca32_fa591_out(h_s_dadda_pg_rca32_and_27_18[0], h_s_dadda_pg_rca32_and_26_19[0], h_s_dadda_pg_rca32_and_25_20[0], h_s_dadda_pg_rca32_fa591_xor1, h_s_dadda_pg_rca32_fa591_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_21(a[24], b[21], h_s_dadda_pg_rca32_and_24_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_22(a[23], b[22], h_s_dadda_pg_rca32_and_23_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_23(a[22], b[23], h_s_dadda_pg_rca32_and_22_23);
  fa fa_h_s_dadda_pg_rca32_fa592_out(h_s_dadda_pg_rca32_and_24_21[0], h_s_dadda_pg_rca32_and_23_22[0], h_s_dadda_pg_rca32_and_22_23[0], h_s_dadda_pg_rca32_fa592_xor1, h_s_dadda_pg_rca32_fa592_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_24(a[21], b[24], h_s_dadda_pg_rca32_and_21_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_25(a[20], b[25], h_s_dadda_pg_rca32_and_20_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_26(a[19], b[26], h_s_dadda_pg_rca32_and_19_26);
  fa fa_h_s_dadda_pg_rca32_fa593_out(h_s_dadda_pg_rca32_and_21_24[0], h_s_dadda_pg_rca32_and_20_25[0], h_s_dadda_pg_rca32_and_19_26[0], h_s_dadda_pg_rca32_fa593_xor1, h_s_dadda_pg_rca32_fa593_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_27(a[18], b[27], h_s_dadda_pg_rca32_and_18_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_28(a[17], b[28], h_s_dadda_pg_rca32_and_17_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_29(a[16], b[29], h_s_dadda_pg_rca32_and_16_29);
  fa fa_h_s_dadda_pg_rca32_fa594_out(h_s_dadda_pg_rca32_and_18_27[0], h_s_dadda_pg_rca32_and_17_28[0], h_s_dadda_pg_rca32_and_16_29[0], h_s_dadda_pg_rca32_fa594_xor1, h_s_dadda_pg_rca32_fa594_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_15_30(a[15], b[30], h_s_dadda_pg_rca32_and_15_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_14_31(a[14], b[31], h_s_dadda_pg_rca32_nand_14_31);
  fa fa_h_s_dadda_pg_rca32_fa595_out(h_s_dadda_pg_rca32_and_15_30[0], h_s_dadda_pg_rca32_nand_14_31[0], h_s_dadda_pg_rca32_fa585_xor1[0], h_s_dadda_pg_rca32_fa595_xor1, h_s_dadda_pg_rca32_fa595_or0);
  fa fa_h_s_dadda_pg_rca32_fa596_out(h_s_dadda_pg_rca32_fa586_xor1[0], h_s_dadda_pg_rca32_fa587_xor1[0], h_s_dadda_pg_rca32_fa588_xor1[0], h_s_dadda_pg_rca32_fa596_xor1, h_s_dadda_pg_rca32_fa596_or0);
  fa fa_h_s_dadda_pg_rca32_fa597_out(h_s_dadda_pg_rca32_fa589_xor1[0], h_s_dadda_pg_rca32_fa590_xor1[0], h_s_dadda_pg_rca32_fa591_xor1[0], h_s_dadda_pg_rca32_fa597_xor1, h_s_dadda_pg_rca32_fa597_or0);
  fa fa_h_s_dadda_pg_rca32_fa598_out(h_s_dadda_pg_rca32_fa597_or0[0], h_s_dadda_pg_rca32_fa596_or0[0], h_s_dadda_pg_rca32_fa595_or0[0], h_s_dadda_pg_rca32_fa598_xor1, h_s_dadda_pg_rca32_fa598_or0);
  fa fa_h_s_dadda_pg_rca32_fa599_out(h_s_dadda_pg_rca32_fa594_or0[0], h_s_dadda_pg_rca32_fa593_or0[0], h_s_dadda_pg_rca32_fa592_or0[0], h_s_dadda_pg_rca32_fa599_xor1, h_s_dadda_pg_rca32_fa599_or0);
  fa fa_h_s_dadda_pg_rca32_fa600_out(h_s_dadda_pg_rca32_fa591_or0[0], h_s_dadda_pg_rca32_fa590_or0[0], h_s_dadda_pg_rca32_fa589_or0[0], h_s_dadda_pg_rca32_fa600_xor1, h_s_dadda_pg_rca32_fa600_or0);
  fa fa_h_s_dadda_pg_rca32_fa601_out(h_s_dadda_pg_rca32_fa588_or0[0], h_s_dadda_pg_rca32_fa587_or0[0], h_s_dadda_pg_rca32_fa586_or0[0], h_s_dadda_pg_rca32_fa601_xor1, h_s_dadda_pg_rca32_fa601_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_15(a[31], b[15], h_s_dadda_pg_rca32_nand_31_15);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_16(a[30], b[16], h_s_dadda_pg_rca32_and_30_16);
  fa fa_h_s_dadda_pg_rca32_fa602_out(h_s_dadda_pg_rca32_fa585_or0[0], h_s_dadda_pg_rca32_nand_31_15[0], h_s_dadda_pg_rca32_and_30_16[0], h_s_dadda_pg_rca32_fa602_xor1, h_s_dadda_pg_rca32_fa602_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_17(a[29], b[17], h_s_dadda_pg_rca32_and_29_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_18(a[28], b[18], h_s_dadda_pg_rca32_and_28_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_19(a[27], b[19], h_s_dadda_pg_rca32_and_27_19);
  fa fa_h_s_dadda_pg_rca32_fa603_out(h_s_dadda_pg_rca32_and_29_17[0], h_s_dadda_pg_rca32_and_28_18[0], h_s_dadda_pg_rca32_and_27_19[0], h_s_dadda_pg_rca32_fa603_xor1, h_s_dadda_pg_rca32_fa603_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_20(a[26], b[20], h_s_dadda_pg_rca32_and_26_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_21(a[25], b[21], h_s_dadda_pg_rca32_and_25_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_22(a[24], b[22], h_s_dadda_pg_rca32_and_24_22);
  fa fa_h_s_dadda_pg_rca32_fa604_out(h_s_dadda_pg_rca32_and_26_20[0], h_s_dadda_pg_rca32_and_25_21[0], h_s_dadda_pg_rca32_and_24_22[0], h_s_dadda_pg_rca32_fa604_xor1, h_s_dadda_pg_rca32_fa604_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_23(a[23], b[23], h_s_dadda_pg_rca32_and_23_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_24(a[22], b[24], h_s_dadda_pg_rca32_and_22_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_25(a[21], b[25], h_s_dadda_pg_rca32_and_21_25);
  fa fa_h_s_dadda_pg_rca32_fa605_out(h_s_dadda_pg_rca32_and_23_23[0], h_s_dadda_pg_rca32_and_22_24[0], h_s_dadda_pg_rca32_and_21_25[0], h_s_dadda_pg_rca32_fa605_xor1, h_s_dadda_pg_rca32_fa605_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_26(a[20], b[26], h_s_dadda_pg_rca32_and_20_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_27(a[19], b[27], h_s_dadda_pg_rca32_and_19_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_28(a[18], b[28], h_s_dadda_pg_rca32_and_18_28);
  fa fa_h_s_dadda_pg_rca32_fa606_out(h_s_dadda_pg_rca32_and_20_26[0], h_s_dadda_pg_rca32_and_19_27[0], h_s_dadda_pg_rca32_and_18_28[0], h_s_dadda_pg_rca32_fa606_xor1, h_s_dadda_pg_rca32_fa606_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_29(a[17], b[29], h_s_dadda_pg_rca32_and_17_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_16_30(a[16], b[30], h_s_dadda_pg_rca32_and_16_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_15_31(a[15], b[31], h_s_dadda_pg_rca32_nand_15_31);
  fa fa_h_s_dadda_pg_rca32_fa607_out(h_s_dadda_pg_rca32_and_17_29[0], h_s_dadda_pg_rca32_and_16_30[0], h_s_dadda_pg_rca32_nand_15_31[0], h_s_dadda_pg_rca32_fa607_xor1, h_s_dadda_pg_rca32_fa607_or0);
  fa fa_h_s_dadda_pg_rca32_fa608_out(h_s_dadda_pg_rca32_fa598_xor1[0], h_s_dadda_pg_rca32_fa599_xor1[0], h_s_dadda_pg_rca32_fa600_xor1[0], h_s_dadda_pg_rca32_fa608_xor1, h_s_dadda_pg_rca32_fa608_or0);
  fa fa_h_s_dadda_pg_rca32_fa609_out(h_s_dadda_pg_rca32_fa601_xor1[0], h_s_dadda_pg_rca32_fa602_xor1[0], h_s_dadda_pg_rca32_fa603_xor1[0], h_s_dadda_pg_rca32_fa609_xor1, h_s_dadda_pg_rca32_fa609_or0);
  fa fa_h_s_dadda_pg_rca32_fa610_out(h_s_dadda_pg_rca32_fa609_or0[0], h_s_dadda_pg_rca32_fa608_or0[0], h_s_dadda_pg_rca32_fa607_or0[0], h_s_dadda_pg_rca32_fa610_xor1, h_s_dadda_pg_rca32_fa610_or0);
  fa fa_h_s_dadda_pg_rca32_fa611_out(h_s_dadda_pg_rca32_fa606_or0[0], h_s_dadda_pg_rca32_fa605_or0[0], h_s_dadda_pg_rca32_fa604_or0[0], h_s_dadda_pg_rca32_fa611_xor1, h_s_dadda_pg_rca32_fa611_or0);
  fa fa_h_s_dadda_pg_rca32_fa612_out(h_s_dadda_pg_rca32_fa603_or0[0], h_s_dadda_pg_rca32_fa602_or0[0], h_s_dadda_pg_rca32_fa601_or0[0], h_s_dadda_pg_rca32_fa612_xor1, h_s_dadda_pg_rca32_fa612_or0);
  fa fa_h_s_dadda_pg_rca32_fa613_out(h_s_dadda_pg_rca32_fa600_or0[0], h_s_dadda_pg_rca32_fa599_or0[0], h_s_dadda_pg_rca32_fa598_or0[0], h_s_dadda_pg_rca32_fa613_xor1, h_s_dadda_pg_rca32_fa613_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_16(a[31], b[16], h_s_dadda_pg_rca32_nand_31_16);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_17(a[30], b[17], h_s_dadda_pg_rca32_and_30_17);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_18(a[29], b[18], h_s_dadda_pg_rca32_and_29_18);
  fa fa_h_s_dadda_pg_rca32_fa614_out(h_s_dadda_pg_rca32_nand_31_16[0], h_s_dadda_pg_rca32_and_30_17[0], h_s_dadda_pg_rca32_and_29_18[0], h_s_dadda_pg_rca32_fa614_xor1, h_s_dadda_pg_rca32_fa614_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_19(a[28], b[19], h_s_dadda_pg_rca32_and_28_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_20(a[27], b[20], h_s_dadda_pg_rca32_and_27_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_21(a[26], b[21], h_s_dadda_pg_rca32_and_26_21);
  fa fa_h_s_dadda_pg_rca32_fa615_out(h_s_dadda_pg_rca32_and_28_19[0], h_s_dadda_pg_rca32_and_27_20[0], h_s_dadda_pg_rca32_and_26_21[0], h_s_dadda_pg_rca32_fa615_xor1, h_s_dadda_pg_rca32_fa615_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_22(a[25], b[22], h_s_dadda_pg_rca32_and_25_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_23(a[24], b[23], h_s_dadda_pg_rca32_and_24_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_24(a[23], b[24], h_s_dadda_pg_rca32_and_23_24);
  fa fa_h_s_dadda_pg_rca32_fa616_out(h_s_dadda_pg_rca32_and_25_22[0], h_s_dadda_pg_rca32_and_24_23[0], h_s_dadda_pg_rca32_and_23_24[0], h_s_dadda_pg_rca32_fa616_xor1, h_s_dadda_pg_rca32_fa616_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_25(a[22], b[25], h_s_dadda_pg_rca32_and_22_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_26(a[21], b[26], h_s_dadda_pg_rca32_and_21_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_27(a[20], b[27], h_s_dadda_pg_rca32_and_20_27);
  fa fa_h_s_dadda_pg_rca32_fa617_out(h_s_dadda_pg_rca32_and_22_25[0], h_s_dadda_pg_rca32_and_21_26[0], h_s_dadda_pg_rca32_and_20_27[0], h_s_dadda_pg_rca32_fa617_xor1, h_s_dadda_pg_rca32_fa617_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_28(a[19], b[28], h_s_dadda_pg_rca32_and_19_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_29(a[18], b[29], h_s_dadda_pg_rca32_and_18_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_17_30(a[17], b[30], h_s_dadda_pg_rca32_and_17_30);
  fa fa_h_s_dadda_pg_rca32_fa618_out(h_s_dadda_pg_rca32_and_19_28[0], h_s_dadda_pg_rca32_and_18_29[0], h_s_dadda_pg_rca32_and_17_30[0], h_s_dadda_pg_rca32_fa618_xor1, h_s_dadda_pg_rca32_fa618_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_16_31(a[16], b[31], h_s_dadda_pg_rca32_nand_16_31);
  fa fa_h_s_dadda_pg_rca32_fa619_out(h_s_dadda_pg_rca32_nand_16_31[0], h_s_dadda_pg_rca32_fa610_xor1[0], h_s_dadda_pg_rca32_fa611_xor1[0], h_s_dadda_pg_rca32_fa619_xor1, h_s_dadda_pg_rca32_fa619_or0);
  fa fa_h_s_dadda_pg_rca32_fa620_out(h_s_dadda_pg_rca32_fa612_xor1[0], h_s_dadda_pg_rca32_fa613_xor1[0], h_s_dadda_pg_rca32_fa614_xor1[0], h_s_dadda_pg_rca32_fa620_xor1, h_s_dadda_pg_rca32_fa620_or0);
  fa fa_h_s_dadda_pg_rca32_fa621_out(h_s_dadda_pg_rca32_fa620_or0[0], h_s_dadda_pg_rca32_fa619_or0[0], h_s_dadda_pg_rca32_fa618_or0[0], h_s_dadda_pg_rca32_fa621_xor1, h_s_dadda_pg_rca32_fa621_or0);
  fa fa_h_s_dadda_pg_rca32_fa622_out(h_s_dadda_pg_rca32_fa617_or0[0], h_s_dadda_pg_rca32_fa616_or0[0], h_s_dadda_pg_rca32_fa615_or0[0], h_s_dadda_pg_rca32_fa622_xor1, h_s_dadda_pg_rca32_fa622_or0);
  fa fa_h_s_dadda_pg_rca32_fa623_out(h_s_dadda_pg_rca32_fa614_or0[0], h_s_dadda_pg_rca32_fa613_or0[0], h_s_dadda_pg_rca32_fa612_or0[0], h_s_dadda_pg_rca32_fa623_xor1, h_s_dadda_pg_rca32_fa623_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_17(a[31], b[17], h_s_dadda_pg_rca32_nand_31_17);
  fa fa_h_s_dadda_pg_rca32_fa624_out(h_s_dadda_pg_rca32_fa611_or0[0], h_s_dadda_pg_rca32_fa610_or0[0], h_s_dadda_pg_rca32_nand_31_17[0], h_s_dadda_pg_rca32_fa624_xor1, h_s_dadda_pg_rca32_fa624_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_18(a[30], b[18], h_s_dadda_pg_rca32_and_30_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_19(a[29], b[19], h_s_dadda_pg_rca32_and_29_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_20(a[28], b[20], h_s_dadda_pg_rca32_and_28_20);
  fa fa_h_s_dadda_pg_rca32_fa625_out(h_s_dadda_pg_rca32_and_30_18[0], h_s_dadda_pg_rca32_and_29_19[0], h_s_dadda_pg_rca32_and_28_20[0], h_s_dadda_pg_rca32_fa625_xor1, h_s_dadda_pg_rca32_fa625_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_21(a[27], b[21], h_s_dadda_pg_rca32_and_27_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_22(a[26], b[22], h_s_dadda_pg_rca32_and_26_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_23(a[25], b[23], h_s_dadda_pg_rca32_and_25_23);
  fa fa_h_s_dadda_pg_rca32_fa626_out(h_s_dadda_pg_rca32_and_27_21[0], h_s_dadda_pg_rca32_and_26_22[0], h_s_dadda_pg_rca32_and_25_23[0], h_s_dadda_pg_rca32_fa626_xor1, h_s_dadda_pg_rca32_fa626_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_24(a[24], b[24], h_s_dadda_pg_rca32_and_24_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_25(a[23], b[25], h_s_dadda_pg_rca32_and_23_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_26(a[22], b[26], h_s_dadda_pg_rca32_and_22_26);
  fa fa_h_s_dadda_pg_rca32_fa627_out(h_s_dadda_pg_rca32_and_24_24[0], h_s_dadda_pg_rca32_and_23_25[0], h_s_dadda_pg_rca32_and_22_26[0], h_s_dadda_pg_rca32_fa627_xor1, h_s_dadda_pg_rca32_fa627_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_27(a[21], b[27], h_s_dadda_pg_rca32_and_21_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_28(a[20], b[28], h_s_dadda_pg_rca32_and_20_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_29(a[19], b[29], h_s_dadda_pg_rca32_and_19_29);
  fa fa_h_s_dadda_pg_rca32_fa628_out(h_s_dadda_pg_rca32_and_21_27[0], h_s_dadda_pg_rca32_and_20_28[0], h_s_dadda_pg_rca32_and_19_29[0], h_s_dadda_pg_rca32_fa628_xor1, h_s_dadda_pg_rca32_fa628_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_18_30(a[18], b[30], h_s_dadda_pg_rca32_and_18_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_17_31(a[17], b[31], h_s_dadda_pg_rca32_nand_17_31);
  fa fa_h_s_dadda_pg_rca32_fa629_out(h_s_dadda_pg_rca32_and_18_30[0], h_s_dadda_pg_rca32_nand_17_31[0], h_s_dadda_pg_rca32_fa621_xor1[0], h_s_dadda_pg_rca32_fa629_xor1, h_s_dadda_pg_rca32_fa629_or0);
  fa fa_h_s_dadda_pg_rca32_fa630_out(h_s_dadda_pg_rca32_fa622_xor1[0], h_s_dadda_pg_rca32_fa623_xor1[0], h_s_dadda_pg_rca32_fa624_xor1[0], h_s_dadda_pg_rca32_fa630_xor1, h_s_dadda_pg_rca32_fa630_or0);
  fa fa_h_s_dadda_pg_rca32_fa631_out(h_s_dadda_pg_rca32_fa630_or0[0], h_s_dadda_pg_rca32_fa629_or0[0], h_s_dadda_pg_rca32_fa628_or0[0], h_s_dadda_pg_rca32_fa631_xor1, h_s_dadda_pg_rca32_fa631_or0);
  fa fa_h_s_dadda_pg_rca32_fa632_out(h_s_dadda_pg_rca32_fa627_or0[0], h_s_dadda_pg_rca32_fa626_or0[0], h_s_dadda_pg_rca32_fa625_or0[0], h_s_dadda_pg_rca32_fa632_xor1, h_s_dadda_pg_rca32_fa632_or0);
  fa fa_h_s_dadda_pg_rca32_fa633_out(h_s_dadda_pg_rca32_fa624_or0[0], h_s_dadda_pg_rca32_fa623_or0[0], h_s_dadda_pg_rca32_fa622_or0[0], h_s_dadda_pg_rca32_fa633_xor1, h_s_dadda_pg_rca32_fa633_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_18(a[31], b[18], h_s_dadda_pg_rca32_nand_31_18);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_19(a[30], b[19], h_s_dadda_pg_rca32_and_30_19);
  fa fa_h_s_dadda_pg_rca32_fa634_out(h_s_dadda_pg_rca32_fa621_or0[0], h_s_dadda_pg_rca32_nand_31_18[0], h_s_dadda_pg_rca32_and_30_19[0], h_s_dadda_pg_rca32_fa634_xor1, h_s_dadda_pg_rca32_fa634_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_20(a[29], b[20], h_s_dadda_pg_rca32_and_29_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_21(a[28], b[21], h_s_dadda_pg_rca32_and_28_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_22(a[27], b[22], h_s_dadda_pg_rca32_and_27_22);
  fa fa_h_s_dadda_pg_rca32_fa635_out(h_s_dadda_pg_rca32_and_29_20[0], h_s_dadda_pg_rca32_and_28_21[0], h_s_dadda_pg_rca32_and_27_22[0], h_s_dadda_pg_rca32_fa635_xor1, h_s_dadda_pg_rca32_fa635_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_23(a[26], b[23], h_s_dadda_pg_rca32_and_26_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_24(a[25], b[24], h_s_dadda_pg_rca32_and_25_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_25(a[24], b[25], h_s_dadda_pg_rca32_and_24_25);
  fa fa_h_s_dadda_pg_rca32_fa636_out(h_s_dadda_pg_rca32_and_26_23[0], h_s_dadda_pg_rca32_and_25_24[0], h_s_dadda_pg_rca32_and_24_25[0], h_s_dadda_pg_rca32_fa636_xor1, h_s_dadda_pg_rca32_fa636_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_26(a[23], b[26], h_s_dadda_pg_rca32_and_23_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_27(a[22], b[27], h_s_dadda_pg_rca32_and_22_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_28(a[21], b[28], h_s_dadda_pg_rca32_and_21_28);
  fa fa_h_s_dadda_pg_rca32_fa637_out(h_s_dadda_pg_rca32_and_23_26[0], h_s_dadda_pg_rca32_and_22_27[0], h_s_dadda_pg_rca32_and_21_28[0], h_s_dadda_pg_rca32_fa637_xor1, h_s_dadda_pg_rca32_fa637_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_29(a[20], b[29], h_s_dadda_pg_rca32_and_20_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_19_30(a[19], b[30], h_s_dadda_pg_rca32_and_19_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_18_31(a[18], b[31], h_s_dadda_pg_rca32_nand_18_31);
  fa fa_h_s_dadda_pg_rca32_fa638_out(h_s_dadda_pg_rca32_and_20_29[0], h_s_dadda_pg_rca32_and_19_30[0], h_s_dadda_pg_rca32_nand_18_31[0], h_s_dadda_pg_rca32_fa638_xor1, h_s_dadda_pg_rca32_fa638_or0);
  fa fa_h_s_dadda_pg_rca32_fa639_out(h_s_dadda_pg_rca32_fa631_xor1[0], h_s_dadda_pg_rca32_fa632_xor1[0], h_s_dadda_pg_rca32_fa633_xor1[0], h_s_dadda_pg_rca32_fa639_xor1, h_s_dadda_pg_rca32_fa639_or0);
  fa fa_h_s_dadda_pg_rca32_fa640_out(h_s_dadda_pg_rca32_fa639_or0[0], h_s_dadda_pg_rca32_fa638_or0[0], h_s_dadda_pg_rca32_fa637_or0[0], h_s_dadda_pg_rca32_fa640_xor1, h_s_dadda_pg_rca32_fa640_or0);
  fa fa_h_s_dadda_pg_rca32_fa641_out(h_s_dadda_pg_rca32_fa636_or0[0], h_s_dadda_pg_rca32_fa635_or0[0], h_s_dadda_pg_rca32_fa634_or0[0], h_s_dadda_pg_rca32_fa641_xor1, h_s_dadda_pg_rca32_fa641_or0);
  fa fa_h_s_dadda_pg_rca32_fa642_out(h_s_dadda_pg_rca32_fa633_or0[0], h_s_dadda_pg_rca32_fa632_or0[0], h_s_dadda_pg_rca32_fa631_or0[0], h_s_dadda_pg_rca32_fa642_xor1, h_s_dadda_pg_rca32_fa642_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_19(a[31], b[19], h_s_dadda_pg_rca32_nand_31_19);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_20(a[30], b[20], h_s_dadda_pg_rca32_and_30_20);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_21(a[29], b[21], h_s_dadda_pg_rca32_and_29_21);
  fa fa_h_s_dadda_pg_rca32_fa643_out(h_s_dadda_pg_rca32_nand_31_19[0], h_s_dadda_pg_rca32_and_30_20[0], h_s_dadda_pg_rca32_and_29_21[0], h_s_dadda_pg_rca32_fa643_xor1, h_s_dadda_pg_rca32_fa643_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_22(a[28], b[22], h_s_dadda_pg_rca32_and_28_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_23(a[27], b[23], h_s_dadda_pg_rca32_and_27_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_24(a[26], b[24], h_s_dadda_pg_rca32_and_26_24);
  fa fa_h_s_dadda_pg_rca32_fa644_out(h_s_dadda_pg_rca32_and_28_22[0], h_s_dadda_pg_rca32_and_27_23[0], h_s_dadda_pg_rca32_and_26_24[0], h_s_dadda_pg_rca32_fa644_xor1, h_s_dadda_pg_rca32_fa644_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_25(a[25], b[25], h_s_dadda_pg_rca32_and_25_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_26(a[24], b[26], h_s_dadda_pg_rca32_and_24_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_27(a[23], b[27], h_s_dadda_pg_rca32_and_23_27);
  fa fa_h_s_dadda_pg_rca32_fa645_out(h_s_dadda_pg_rca32_and_25_25[0], h_s_dadda_pg_rca32_and_24_26[0], h_s_dadda_pg_rca32_and_23_27[0], h_s_dadda_pg_rca32_fa645_xor1, h_s_dadda_pg_rca32_fa645_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_28(a[22], b[28], h_s_dadda_pg_rca32_and_22_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_29(a[21], b[29], h_s_dadda_pg_rca32_and_21_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_20_30(a[20], b[30], h_s_dadda_pg_rca32_and_20_30);
  fa fa_h_s_dadda_pg_rca32_fa646_out(h_s_dadda_pg_rca32_and_22_28[0], h_s_dadda_pg_rca32_and_21_29[0], h_s_dadda_pg_rca32_and_20_30[0], h_s_dadda_pg_rca32_fa646_xor1, h_s_dadda_pg_rca32_fa646_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_19_31(a[19], b[31], h_s_dadda_pg_rca32_nand_19_31);
  fa fa_h_s_dadda_pg_rca32_fa647_out(h_s_dadda_pg_rca32_nand_19_31[0], h_s_dadda_pg_rca32_fa640_xor1[0], h_s_dadda_pg_rca32_fa641_xor1[0], h_s_dadda_pg_rca32_fa647_xor1, h_s_dadda_pg_rca32_fa647_or0);
  fa fa_h_s_dadda_pg_rca32_fa648_out(h_s_dadda_pg_rca32_fa647_or0[0], h_s_dadda_pg_rca32_fa646_or0[0], h_s_dadda_pg_rca32_fa645_or0[0], h_s_dadda_pg_rca32_fa648_xor1, h_s_dadda_pg_rca32_fa648_or0);
  fa fa_h_s_dadda_pg_rca32_fa649_out(h_s_dadda_pg_rca32_fa644_or0[0], h_s_dadda_pg_rca32_fa643_or0[0], h_s_dadda_pg_rca32_fa642_or0[0], h_s_dadda_pg_rca32_fa649_xor1, h_s_dadda_pg_rca32_fa649_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_20(a[31], b[20], h_s_dadda_pg_rca32_nand_31_20);
  fa fa_h_s_dadda_pg_rca32_fa650_out(h_s_dadda_pg_rca32_fa641_or0[0], h_s_dadda_pg_rca32_fa640_or0[0], h_s_dadda_pg_rca32_nand_31_20[0], h_s_dadda_pg_rca32_fa650_xor1, h_s_dadda_pg_rca32_fa650_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_21(a[30], b[21], h_s_dadda_pg_rca32_and_30_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_22(a[29], b[22], h_s_dadda_pg_rca32_and_29_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_23(a[28], b[23], h_s_dadda_pg_rca32_and_28_23);
  fa fa_h_s_dadda_pg_rca32_fa651_out(h_s_dadda_pg_rca32_and_30_21[0], h_s_dadda_pg_rca32_and_29_22[0], h_s_dadda_pg_rca32_and_28_23[0], h_s_dadda_pg_rca32_fa651_xor1, h_s_dadda_pg_rca32_fa651_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_24(a[27], b[24], h_s_dadda_pg_rca32_and_27_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_25(a[26], b[25], h_s_dadda_pg_rca32_and_26_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_26(a[25], b[26], h_s_dadda_pg_rca32_and_25_26);
  fa fa_h_s_dadda_pg_rca32_fa652_out(h_s_dadda_pg_rca32_and_27_24[0], h_s_dadda_pg_rca32_and_26_25[0], h_s_dadda_pg_rca32_and_25_26[0], h_s_dadda_pg_rca32_fa652_xor1, h_s_dadda_pg_rca32_fa652_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_27(a[24], b[27], h_s_dadda_pg_rca32_and_24_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_28(a[23], b[28], h_s_dadda_pg_rca32_and_23_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_29(a[22], b[29], h_s_dadda_pg_rca32_and_22_29);
  fa fa_h_s_dadda_pg_rca32_fa653_out(h_s_dadda_pg_rca32_and_24_27[0], h_s_dadda_pg_rca32_and_23_28[0], h_s_dadda_pg_rca32_and_22_29[0], h_s_dadda_pg_rca32_fa653_xor1, h_s_dadda_pg_rca32_fa653_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_21_30(a[21], b[30], h_s_dadda_pg_rca32_and_21_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_20_31(a[20], b[31], h_s_dadda_pg_rca32_nand_20_31);
  fa fa_h_s_dadda_pg_rca32_fa654_out(h_s_dadda_pg_rca32_and_21_30[0], h_s_dadda_pg_rca32_nand_20_31[0], h_s_dadda_pg_rca32_fa648_xor1[0], h_s_dadda_pg_rca32_fa654_xor1, h_s_dadda_pg_rca32_fa654_or0);
  fa fa_h_s_dadda_pg_rca32_fa655_out(h_s_dadda_pg_rca32_fa654_or0[0], h_s_dadda_pg_rca32_fa653_or0[0], h_s_dadda_pg_rca32_fa652_or0[0], h_s_dadda_pg_rca32_fa655_xor1, h_s_dadda_pg_rca32_fa655_or0);
  fa fa_h_s_dadda_pg_rca32_fa656_out(h_s_dadda_pg_rca32_fa651_or0[0], h_s_dadda_pg_rca32_fa650_or0[0], h_s_dadda_pg_rca32_fa649_or0[0], h_s_dadda_pg_rca32_fa656_xor1, h_s_dadda_pg_rca32_fa656_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_21(a[31], b[21], h_s_dadda_pg_rca32_nand_31_21);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_22(a[30], b[22], h_s_dadda_pg_rca32_and_30_22);
  fa fa_h_s_dadda_pg_rca32_fa657_out(h_s_dadda_pg_rca32_fa648_or0[0], h_s_dadda_pg_rca32_nand_31_21[0], h_s_dadda_pg_rca32_and_30_22[0], h_s_dadda_pg_rca32_fa657_xor1, h_s_dadda_pg_rca32_fa657_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_23(a[29], b[23], h_s_dadda_pg_rca32_and_29_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_24(a[28], b[24], h_s_dadda_pg_rca32_and_28_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_25(a[27], b[25], h_s_dadda_pg_rca32_and_27_25);
  fa fa_h_s_dadda_pg_rca32_fa658_out(h_s_dadda_pg_rca32_and_29_23[0], h_s_dadda_pg_rca32_and_28_24[0], h_s_dadda_pg_rca32_and_27_25[0], h_s_dadda_pg_rca32_fa658_xor1, h_s_dadda_pg_rca32_fa658_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_26(a[26], b[26], h_s_dadda_pg_rca32_and_26_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_27(a[25], b[27], h_s_dadda_pg_rca32_and_25_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_28(a[24], b[28], h_s_dadda_pg_rca32_and_24_28);
  fa fa_h_s_dadda_pg_rca32_fa659_out(h_s_dadda_pg_rca32_and_26_26[0], h_s_dadda_pg_rca32_and_25_27[0], h_s_dadda_pg_rca32_and_24_28[0], h_s_dadda_pg_rca32_fa659_xor1, h_s_dadda_pg_rca32_fa659_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_29(a[23], b[29], h_s_dadda_pg_rca32_and_23_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_22_30(a[22], b[30], h_s_dadda_pg_rca32_and_22_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_21_31(a[21], b[31], h_s_dadda_pg_rca32_nand_21_31);
  fa fa_h_s_dadda_pg_rca32_fa660_out(h_s_dadda_pg_rca32_and_23_29[0], h_s_dadda_pg_rca32_and_22_30[0], h_s_dadda_pg_rca32_nand_21_31[0], h_s_dadda_pg_rca32_fa660_xor1, h_s_dadda_pg_rca32_fa660_or0);
  fa fa_h_s_dadda_pg_rca32_fa661_out(h_s_dadda_pg_rca32_fa660_or0[0], h_s_dadda_pg_rca32_fa659_or0[0], h_s_dadda_pg_rca32_fa658_or0[0], h_s_dadda_pg_rca32_fa661_xor1, h_s_dadda_pg_rca32_fa661_or0);
  fa fa_h_s_dadda_pg_rca32_fa662_out(h_s_dadda_pg_rca32_fa657_or0[0], h_s_dadda_pg_rca32_fa656_or0[0], h_s_dadda_pg_rca32_fa655_or0[0], h_s_dadda_pg_rca32_fa662_xor1, h_s_dadda_pg_rca32_fa662_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_22(a[31], b[22], h_s_dadda_pg_rca32_nand_31_22);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_23(a[30], b[23], h_s_dadda_pg_rca32_and_30_23);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_24(a[29], b[24], h_s_dadda_pg_rca32_and_29_24);
  fa fa_h_s_dadda_pg_rca32_fa663_out(h_s_dadda_pg_rca32_nand_31_22[0], h_s_dadda_pg_rca32_and_30_23[0], h_s_dadda_pg_rca32_and_29_24[0], h_s_dadda_pg_rca32_fa663_xor1, h_s_dadda_pg_rca32_fa663_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_25(a[28], b[25], h_s_dadda_pg_rca32_and_28_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_26(a[27], b[26], h_s_dadda_pg_rca32_and_27_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_27(a[26], b[27], h_s_dadda_pg_rca32_and_26_27);
  fa fa_h_s_dadda_pg_rca32_fa664_out(h_s_dadda_pg_rca32_and_28_25[0], h_s_dadda_pg_rca32_and_27_26[0], h_s_dadda_pg_rca32_and_26_27[0], h_s_dadda_pg_rca32_fa664_xor1, h_s_dadda_pg_rca32_fa664_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_28(a[25], b[28], h_s_dadda_pg_rca32_and_25_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_29(a[24], b[29], h_s_dadda_pg_rca32_and_24_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_23_30(a[23], b[30], h_s_dadda_pg_rca32_and_23_30);
  fa fa_h_s_dadda_pg_rca32_fa665_out(h_s_dadda_pg_rca32_and_25_28[0], h_s_dadda_pg_rca32_and_24_29[0], h_s_dadda_pg_rca32_and_23_30[0], h_s_dadda_pg_rca32_fa665_xor1, h_s_dadda_pg_rca32_fa665_or0);
  fa fa_h_s_dadda_pg_rca32_fa666_out(h_s_dadda_pg_rca32_fa665_or0[0], h_s_dadda_pg_rca32_fa664_or0[0], h_s_dadda_pg_rca32_fa663_or0[0], h_s_dadda_pg_rca32_fa666_xor1, h_s_dadda_pg_rca32_fa666_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_23(a[31], b[23], h_s_dadda_pg_rca32_nand_31_23);
  fa fa_h_s_dadda_pg_rca32_fa667_out(h_s_dadda_pg_rca32_fa662_or0[0], h_s_dadda_pg_rca32_fa661_or0[0], h_s_dadda_pg_rca32_nand_31_23[0], h_s_dadda_pg_rca32_fa667_xor1, h_s_dadda_pg_rca32_fa667_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_24(a[30], b[24], h_s_dadda_pg_rca32_and_30_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_25(a[29], b[25], h_s_dadda_pg_rca32_and_29_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_26(a[28], b[26], h_s_dadda_pg_rca32_and_28_26);
  fa fa_h_s_dadda_pg_rca32_fa668_out(h_s_dadda_pg_rca32_and_30_24[0], h_s_dadda_pg_rca32_and_29_25[0], h_s_dadda_pg_rca32_and_28_26[0], h_s_dadda_pg_rca32_fa668_xor1, h_s_dadda_pg_rca32_fa668_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_27(a[27], b[27], h_s_dadda_pg_rca32_and_27_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_28(a[26], b[28], h_s_dadda_pg_rca32_and_26_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_29(a[25], b[29], h_s_dadda_pg_rca32_and_25_29);
  fa fa_h_s_dadda_pg_rca32_fa669_out(h_s_dadda_pg_rca32_and_27_27[0], h_s_dadda_pg_rca32_and_26_28[0], h_s_dadda_pg_rca32_and_25_29[0], h_s_dadda_pg_rca32_fa669_xor1, h_s_dadda_pg_rca32_fa669_or0);
  fa fa_h_s_dadda_pg_rca32_fa670_out(h_s_dadda_pg_rca32_fa669_or0[0], h_s_dadda_pg_rca32_fa668_or0[0], h_s_dadda_pg_rca32_fa667_or0[0], h_s_dadda_pg_rca32_fa670_xor1, h_s_dadda_pg_rca32_fa670_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_24(a[31], b[24], h_s_dadda_pg_rca32_nand_31_24);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_25(a[30], b[25], h_s_dadda_pg_rca32_and_30_25);
  fa fa_h_s_dadda_pg_rca32_fa671_out(h_s_dadda_pg_rca32_fa666_or0[0], h_s_dadda_pg_rca32_nand_31_24[0], h_s_dadda_pg_rca32_and_30_25[0], h_s_dadda_pg_rca32_fa671_xor1, h_s_dadda_pg_rca32_fa671_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_26(a[29], b[26], h_s_dadda_pg_rca32_and_29_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_27(a[28], b[27], h_s_dadda_pg_rca32_and_28_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_28(a[27], b[28], h_s_dadda_pg_rca32_and_27_28);
  fa fa_h_s_dadda_pg_rca32_fa672_out(h_s_dadda_pg_rca32_and_29_26[0], h_s_dadda_pg_rca32_and_28_27[0], h_s_dadda_pg_rca32_and_27_28[0], h_s_dadda_pg_rca32_fa672_xor1, h_s_dadda_pg_rca32_fa672_or0);
  fa fa_h_s_dadda_pg_rca32_fa673_out(h_s_dadda_pg_rca32_fa672_or0[0], h_s_dadda_pg_rca32_fa671_or0[0], h_s_dadda_pg_rca32_fa670_or0[0], h_s_dadda_pg_rca32_fa673_xor1, h_s_dadda_pg_rca32_fa673_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_25(a[31], b[25], h_s_dadda_pg_rca32_nand_31_25);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_26(a[30], b[26], h_s_dadda_pg_rca32_and_30_26);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_27(a[29], b[27], h_s_dadda_pg_rca32_and_29_27);
  fa fa_h_s_dadda_pg_rca32_fa674_out(h_s_dadda_pg_rca32_nand_31_25[0], h_s_dadda_pg_rca32_and_30_26[0], h_s_dadda_pg_rca32_and_29_27[0], h_s_dadda_pg_rca32_fa674_xor1, h_s_dadda_pg_rca32_fa674_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_26(a[31], b[26], h_s_dadda_pg_rca32_nand_31_26);
  fa fa_h_s_dadda_pg_rca32_fa675_out(h_s_dadda_pg_rca32_fa674_or0[0], h_s_dadda_pg_rca32_fa673_or0[0], h_s_dadda_pg_rca32_nand_31_26[0], h_s_dadda_pg_rca32_fa675_xor1, h_s_dadda_pg_rca32_fa675_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_0(a[4], b[0], h_s_dadda_pg_rca32_and_4_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_1(a[3], b[1], h_s_dadda_pg_rca32_and_3_1);
  ha ha_h_s_dadda_pg_rca32_ha26_out(h_s_dadda_pg_rca32_and_4_0[0], h_s_dadda_pg_rca32_and_3_1[0], h_s_dadda_pg_rca32_ha26_xor0, h_s_dadda_pg_rca32_ha26_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_5_0(a[5], b[0], h_s_dadda_pg_rca32_and_5_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_1(a[4], b[1], h_s_dadda_pg_rca32_and_4_1);
  fa fa_h_s_dadda_pg_rca32_fa676_out(h_s_dadda_pg_rca32_ha26_and0[0], h_s_dadda_pg_rca32_and_5_0[0], h_s_dadda_pg_rca32_and_4_1[0], h_s_dadda_pg_rca32_fa676_xor1, h_s_dadda_pg_rca32_fa676_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_2(a[3], b[2], h_s_dadda_pg_rca32_and_3_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_3(a[2], b[3], h_s_dadda_pg_rca32_and_2_3);
  ha ha_h_s_dadda_pg_rca32_ha27_out(h_s_dadda_pg_rca32_and_3_2[0], h_s_dadda_pg_rca32_and_2_3[0], h_s_dadda_pg_rca32_ha27_xor0, h_s_dadda_pg_rca32_ha27_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_4_2(a[4], b[2], h_s_dadda_pg_rca32_and_4_2);
  fa fa_h_s_dadda_pg_rca32_fa677_out(h_s_dadda_pg_rca32_ha27_and0[0], h_s_dadda_pg_rca32_fa676_or0[0], h_s_dadda_pg_rca32_and_4_2[0], h_s_dadda_pg_rca32_fa677_xor1, h_s_dadda_pg_rca32_fa677_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_3(a[3], b[3], h_s_dadda_pg_rca32_and_3_3);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_4(a[2], b[4], h_s_dadda_pg_rca32_and_2_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_5(a[1], b[5], h_s_dadda_pg_rca32_and_1_5);
  fa fa_h_s_dadda_pg_rca32_fa678_out(h_s_dadda_pg_rca32_and_3_3[0], h_s_dadda_pg_rca32_and_2_4[0], h_s_dadda_pg_rca32_and_1_5[0], h_s_dadda_pg_rca32_fa678_xor1, h_s_dadda_pg_rca32_fa678_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_4(a[3], b[4], h_s_dadda_pg_rca32_and_3_4);
  fa fa_h_s_dadda_pg_rca32_fa679_out(h_s_dadda_pg_rca32_fa678_or0[0], h_s_dadda_pg_rca32_fa677_or0[0], h_s_dadda_pg_rca32_and_3_4[0], h_s_dadda_pg_rca32_fa679_xor1, h_s_dadda_pg_rca32_fa679_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_5(a[2], b[5], h_s_dadda_pg_rca32_and_2_5);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_6(a[1], b[6], h_s_dadda_pg_rca32_and_1_6);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_7(a[0], b[7], h_s_dadda_pg_rca32_and_0_7);
  fa fa_h_s_dadda_pg_rca32_fa680_out(h_s_dadda_pg_rca32_and_2_5[0], h_s_dadda_pg_rca32_and_1_6[0], h_s_dadda_pg_rca32_and_0_7[0], h_s_dadda_pg_rca32_fa680_xor1, h_s_dadda_pg_rca32_fa680_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_6(a[2], b[6], h_s_dadda_pg_rca32_and_2_6);
  fa fa_h_s_dadda_pg_rca32_fa681_out(h_s_dadda_pg_rca32_fa680_or0[0], h_s_dadda_pg_rca32_fa679_or0[0], h_s_dadda_pg_rca32_and_2_6[0], h_s_dadda_pg_rca32_fa681_xor1, h_s_dadda_pg_rca32_fa681_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_7(a[1], b[7], h_s_dadda_pg_rca32_and_1_7);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_8(a[0], b[8], h_s_dadda_pg_rca32_and_0_8);
  fa fa_h_s_dadda_pg_rca32_fa682_out(h_s_dadda_pg_rca32_and_1_7[0], h_s_dadda_pg_rca32_and_0_8[0], h_s_dadda_pg_rca32_fa17_xor1[0], h_s_dadda_pg_rca32_fa682_xor1, h_s_dadda_pg_rca32_fa682_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_8(a[1], b[8], h_s_dadda_pg_rca32_and_1_8);
  fa fa_h_s_dadda_pg_rca32_fa683_out(h_s_dadda_pg_rca32_fa682_or0[0], h_s_dadda_pg_rca32_fa681_or0[0], h_s_dadda_pg_rca32_and_1_8[0], h_s_dadda_pg_rca32_fa683_xor1, h_s_dadda_pg_rca32_fa683_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_9(a[0], b[9], h_s_dadda_pg_rca32_and_0_9);
  fa fa_h_s_dadda_pg_rca32_fa684_out(h_s_dadda_pg_rca32_and_0_9[0], h_s_dadda_pg_rca32_fa19_xor1[0], h_s_dadda_pg_rca32_fa20_xor1[0], h_s_dadda_pg_rca32_fa684_xor1, h_s_dadda_pg_rca32_fa684_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_10(a[0], b[10], h_s_dadda_pg_rca32_and_0_10);
  fa fa_h_s_dadda_pg_rca32_fa685_out(h_s_dadda_pg_rca32_fa684_or0[0], h_s_dadda_pg_rca32_fa683_or0[0], h_s_dadda_pg_rca32_and_0_10[0], h_s_dadda_pg_rca32_fa685_xor1, h_s_dadda_pg_rca32_fa685_or0);
  fa fa_h_s_dadda_pg_rca32_fa686_out(h_s_dadda_pg_rca32_fa22_xor1[0], h_s_dadda_pg_rca32_fa23_xor1[0], h_s_dadda_pg_rca32_fa24_xor1[0], h_s_dadda_pg_rca32_fa686_xor1, h_s_dadda_pg_rca32_fa686_or0);
  fa fa_h_s_dadda_pg_rca32_fa687_out(h_s_dadda_pg_rca32_fa686_or0[0], h_s_dadda_pg_rca32_fa685_or0[0], h_s_dadda_pg_rca32_fa26_xor1[0], h_s_dadda_pg_rca32_fa687_xor1, h_s_dadda_pg_rca32_fa687_or0);
  fa fa_h_s_dadda_pg_rca32_fa688_out(h_s_dadda_pg_rca32_fa27_xor1[0], h_s_dadda_pg_rca32_fa28_xor1[0], h_s_dadda_pg_rca32_fa29_xor1[0], h_s_dadda_pg_rca32_fa688_xor1, h_s_dadda_pg_rca32_fa688_or0);
  fa fa_h_s_dadda_pg_rca32_fa689_out(h_s_dadda_pg_rca32_fa688_or0[0], h_s_dadda_pg_rca32_fa687_or0[0], h_s_dadda_pg_rca32_fa32_xor1[0], h_s_dadda_pg_rca32_fa689_xor1, h_s_dadda_pg_rca32_fa689_or0);
  fa fa_h_s_dadda_pg_rca32_fa690_out(h_s_dadda_pg_rca32_fa33_xor1[0], h_s_dadda_pg_rca32_fa34_xor1[0], h_s_dadda_pg_rca32_fa35_xor1[0], h_s_dadda_pg_rca32_fa690_xor1, h_s_dadda_pg_rca32_fa690_or0);
  fa fa_h_s_dadda_pg_rca32_fa691_out(h_s_dadda_pg_rca32_fa690_or0[0], h_s_dadda_pg_rca32_fa689_or0[0], h_s_dadda_pg_rca32_fa39_xor1[0], h_s_dadda_pg_rca32_fa691_xor1, h_s_dadda_pg_rca32_fa691_or0);
  fa fa_h_s_dadda_pg_rca32_fa692_out(h_s_dadda_pg_rca32_fa40_xor1[0], h_s_dadda_pg_rca32_fa41_xor1[0], h_s_dadda_pg_rca32_fa42_xor1[0], h_s_dadda_pg_rca32_fa692_xor1, h_s_dadda_pg_rca32_fa692_or0);
  fa fa_h_s_dadda_pg_rca32_fa693_out(h_s_dadda_pg_rca32_fa692_or0[0], h_s_dadda_pg_rca32_fa691_or0[0], h_s_dadda_pg_rca32_fa47_xor1[0], h_s_dadda_pg_rca32_fa693_xor1, h_s_dadda_pg_rca32_fa693_or0);
  fa fa_h_s_dadda_pg_rca32_fa694_out(h_s_dadda_pg_rca32_fa48_xor1[0], h_s_dadda_pg_rca32_fa49_xor1[0], h_s_dadda_pg_rca32_fa50_xor1[0], h_s_dadda_pg_rca32_fa694_xor1, h_s_dadda_pg_rca32_fa694_or0);
  fa fa_h_s_dadda_pg_rca32_fa695_out(h_s_dadda_pg_rca32_fa694_or0[0], h_s_dadda_pg_rca32_fa693_or0[0], h_s_dadda_pg_rca32_fa56_xor1[0], h_s_dadda_pg_rca32_fa695_xor1, h_s_dadda_pg_rca32_fa695_or0);
  fa fa_h_s_dadda_pg_rca32_fa696_out(h_s_dadda_pg_rca32_fa57_xor1[0], h_s_dadda_pg_rca32_fa58_xor1[0], h_s_dadda_pg_rca32_fa59_xor1[0], h_s_dadda_pg_rca32_fa696_xor1, h_s_dadda_pg_rca32_fa696_or0);
  fa fa_h_s_dadda_pg_rca32_fa697_out(h_s_dadda_pg_rca32_fa696_or0[0], h_s_dadda_pg_rca32_fa695_or0[0], h_s_dadda_pg_rca32_fa66_xor1[0], h_s_dadda_pg_rca32_fa697_xor1, h_s_dadda_pg_rca32_fa697_or0);
  fa fa_h_s_dadda_pg_rca32_fa698_out(h_s_dadda_pg_rca32_fa67_xor1[0], h_s_dadda_pg_rca32_fa68_xor1[0], h_s_dadda_pg_rca32_fa69_xor1[0], h_s_dadda_pg_rca32_fa698_xor1, h_s_dadda_pg_rca32_fa698_or0);
  fa fa_h_s_dadda_pg_rca32_fa699_out(h_s_dadda_pg_rca32_fa698_or0[0], h_s_dadda_pg_rca32_fa697_or0[0], h_s_dadda_pg_rca32_fa77_xor1[0], h_s_dadda_pg_rca32_fa699_xor1, h_s_dadda_pg_rca32_fa699_or0);
  fa fa_h_s_dadda_pg_rca32_fa700_out(h_s_dadda_pg_rca32_fa78_xor1[0], h_s_dadda_pg_rca32_fa79_xor1[0], h_s_dadda_pg_rca32_fa80_xor1[0], h_s_dadda_pg_rca32_fa700_xor1, h_s_dadda_pg_rca32_fa700_or0);
  fa fa_h_s_dadda_pg_rca32_fa701_out(h_s_dadda_pg_rca32_fa700_or0[0], h_s_dadda_pg_rca32_fa699_or0[0], h_s_dadda_pg_rca32_fa89_xor1[0], h_s_dadda_pg_rca32_fa701_xor1, h_s_dadda_pg_rca32_fa701_or0);
  fa fa_h_s_dadda_pg_rca32_fa702_out(h_s_dadda_pg_rca32_fa90_xor1[0], h_s_dadda_pg_rca32_fa91_xor1[0], h_s_dadda_pg_rca32_fa92_xor1[0], h_s_dadda_pg_rca32_fa702_xor1, h_s_dadda_pg_rca32_fa702_or0);
  fa fa_h_s_dadda_pg_rca32_fa703_out(h_s_dadda_pg_rca32_fa702_or0[0], h_s_dadda_pg_rca32_fa701_or0[0], h_s_dadda_pg_rca32_fa102_xor1[0], h_s_dadda_pg_rca32_fa703_xor1, h_s_dadda_pg_rca32_fa703_or0);
  fa fa_h_s_dadda_pg_rca32_fa704_out(h_s_dadda_pg_rca32_fa103_xor1[0], h_s_dadda_pg_rca32_fa104_xor1[0], h_s_dadda_pg_rca32_fa105_xor1[0], h_s_dadda_pg_rca32_fa704_xor1, h_s_dadda_pg_rca32_fa704_or0);
  fa fa_h_s_dadda_pg_rca32_fa705_out(h_s_dadda_pg_rca32_fa704_or0[0], h_s_dadda_pg_rca32_fa703_or0[0], h_s_dadda_pg_rca32_fa116_xor1[0], h_s_dadda_pg_rca32_fa705_xor1, h_s_dadda_pg_rca32_fa705_or0);
  fa fa_h_s_dadda_pg_rca32_fa706_out(h_s_dadda_pg_rca32_fa117_xor1[0], h_s_dadda_pg_rca32_fa118_xor1[0], h_s_dadda_pg_rca32_fa119_xor1[0], h_s_dadda_pg_rca32_fa706_xor1, h_s_dadda_pg_rca32_fa706_or0);
  fa fa_h_s_dadda_pg_rca32_fa707_out(h_s_dadda_pg_rca32_fa706_or0[0], h_s_dadda_pg_rca32_fa705_or0[0], h_s_dadda_pg_rca32_fa131_xor1[0], h_s_dadda_pg_rca32_fa707_xor1, h_s_dadda_pg_rca32_fa707_or0);
  fa fa_h_s_dadda_pg_rca32_fa708_out(h_s_dadda_pg_rca32_fa132_xor1[0], h_s_dadda_pg_rca32_fa133_xor1[0], h_s_dadda_pg_rca32_fa134_xor1[0], h_s_dadda_pg_rca32_fa708_xor1, h_s_dadda_pg_rca32_fa708_or0);
  fa fa_h_s_dadda_pg_rca32_fa709_out(h_s_dadda_pg_rca32_fa708_or0[0], h_s_dadda_pg_rca32_fa707_or0[0], h_s_dadda_pg_rca32_fa147_xor1[0], h_s_dadda_pg_rca32_fa709_xor1, h_s_dadda_pg_rca32_fa709_or0);
  fa fa_h_s_dadda_pg_rca32_fa710_out(h_s_dadda_pg_rca32_fa148_xor1[0], h_s_dadda_pg_rca32_fa149_xor1[0], h_s_dadda_pg_rca32_fa150_xor1[0], h_s_dadda_pg_rca32_fa710_xor1, h_s_dadda_pg_rca32_fa710_or0);
  fa fa_h_s_dadda_pg_rca32_fa711_out(h_s_dadda_pg_rca32_fa710_or0[0], h_s_dadda_pg_rca32_fa709_or0[0], h_s_dadda_pg_rca32_fa164_xor1[0], h_s_dadda_pg_rca32_fa711_xor1, h_s_dadda_pg_rca32_fa711_or0);
  fa fa_h_s_dadda_pg_rca32_fa712_out(h_s_dadda_pg_rca32_fa165_xor1[0], h_s_dadda_pg_rca32_fa166_xor1[0], h_s_dadda_pg_rca32_fa167_xor1[0], h_s_dadda_pg_rca32_fa712_xor1, h_s_dadda_pg_rca32_fa712_or0);
  fa fa_h_s_dadda_pg_rca32_fa713_out(h_s_dadda_pg_rca32_fa712_or0[0], h_s_dadda_pg_rca32_fa711_or0[0], h_s_dadda_pg_rca32_fa182_xor1[0], h_s_dadda_pg_rca32_fa713_xor1, h_s_dadda_pg_rca32_fa713_or0);
  fa fa_h_s_dadda_pg_rca32_fa714_out(h_s_dadda_pg_rca32_fa183_xor1[0], h_s_dadda_pg_rca32_fa184_xor1[0], h_s_dadda_pg_rca32_fa185_xor1[0], h_s_dadda_pg_rca32_fa714_xor1, h_s_dadda_pg_rca32_fa714_or0);
  fa fa_h_s_dadda_pg_rca32_fa715_out(h_s_dadda_pg_rca32_fa714_or0[0], h_s_dadda_pg_rca32_fa713_or0[0], h_s_dadda_pg_rca32_fa201_xor1[0], h_s_dadda_pg_rca32_fa715_xor1, h_s_dadda_pg_rca32_fa715_or0);
  fa fa_h_s_dadda_pg_rca32_fa716_out(h_s_dadda_pg_rca32_fa202_xor1[0], h_s_dadda_pg_rca32_fa203_xor1[0], h_s_dadda_pg_rca32_fa204_xor1[0], h_s_dadda_pg_rca32_fa716_xor1, h_s_dadda_pg_rca32_fa716_or0);
  fa fa_h_s_dadda_pg_rca32_fa717_out(h_s_dadda_pg_rca32_fa716_or0[0], h_s_dadda_pg_rca32_fa715_or0[0], h_s_dadda_pg_rca32_fa221_xor1[0], h_s_dadda_pg_rca32_fa717_xor1, h_s_dadda_pg_rca32_fa717_or0);
  fa fa_h_s_dadda_pg_rca32_fa718_out(h_s_dadda_pg_rca32_fa222_xor1[0], h_s_dadda_pg_rca32_fa223_xor1[0], h_s_dadda_pg_rca32_fa224_xor1[0], h_s_dadda_pg_rca32_fa718_xor1, h_s_dadda_pg_rca32_fa718_or0);
  fa fa_h_s_dadda_pg_rca32_fa719_out(h_s_dadda_pg_rca32_fa718_or0[0], h_s_dadda_pg_rca32_fa717_or0[0], h_s_dadda_pg_rca32_fa242_xor1[0], h_s_dadda_pg_rca32_fa719_xor1, h_s_dadda_pg_rca32_fa719_or0);
  fa fa_h_s_dadda_pg_rca32_fa720_out(h_s_dadda_pg_rca32_fa243_xor1[0], h_s_dadda_pg_rca32_fa244_xor1[0], h_s_dadda_pg_rca32_fa245_xor1[0], h_s_dadda_pg_rca32_fa720_xor1, h_s_dadda_pg_rca32_fa720_or0);
  fa fa_h_s_dadda_pg_rca32_fa721_out(h_s_dadda_pg_rca32_fa720_or0[0], h_s_dadda_pg_rca32_fa719_or0[0], h_s_dadda_pg_rca32_fa263_xor1[0], h_s_dadda_pg_rca32_fa721_xor1, h_s_dadda_pg_rca32_fa721_or0);
  fa fa_h_s_dadda_pg_rca32_fa722_out(h_s_dadda_pg_rca32_fa264_xor1[0], h_s_dadda_pg_rca32_fa265_xor1[0], h_s_dadda_pg_rca32_fa266_xor1[0], h_s_dadda_pg_rca32_fa722_xor1, h_s_dadda_pg_rca32_fa722_or0);
  fa fa_h_s_dadda_pg_rca32_fa723_out(h_s_dadda_pg_rca32_fa722_or0[0], h_s_dadda_pg_rca32_fa721_or0[0], h_s_dadda_pg_rca32_fa285_xor1[0], h_s_dadda_pg_rca32_fa723_xor1, h_s_dadda_pg_rca32_fa723_or0);
  fa fa_h_s_dadda_pg_rca32_fa724_out(h_s_dadda_pg_rca32_fa286_xor1[0], h_s_dadda_pg_rca32_fa287_xor1[0], h_s_dadda_pg_rca32_fa288_xor1[0], h_s_dadda_pg_rca32_fa724_xor1, h_s_dadda_pg_rca32_fa724_or0);
  fa fa_h_s_dadda_pg_rca32_fa725_out(h_s_dadda_pg_rca32_fa724_or0[0], h_s_dadda_pg_rca32_fa723_or0[0], h_s_dadda_pg_rca32_fa307_xor1[0], h_s_dadda_pg_rca32_fa725_xor1, h_s_dadda_pg_rca32_fa725_or0);
  fa fa_h_s_dadda_pg_rca32_fa726_out(h_s_dadda_pg_rca32_fa308_xor1[0], h_s_dadda_pg_rca32_fa309_xor1[0], h_s_dadda_pg_rca32_fa310_xor1[0], h_s_dadda_pg_rca32_fa726_xor1, h_s_dadda_pg_rca32_fa726_or0);
  fa fa_h_s_dadda_pg_rca32_fa727_out(h_s_dadda_pg_rca32_fa726_or0[0], h_s_dadda_pg_rca32_fa725_or0[0], h_s_dadda_pg_rca32_fa329_xor1[0], h_s_dadda_pg_rca32_fa727_xor1, h_s_dadda_pg_rca32_fa727_or0);
  fa fa_h_s_dadda_pg_rca32_fa728_out(h_s_dadda_pg_rca32_fa330_xor1[0], h_s_dadda_pg_rca32_fa331_xor1[0], h_s_dadda_pg_rca32_fa332_xor1[0], h_s_dadda_pg_rca32_fa728_xor1, h_s_dadda_pg_rca32_fa728_or0);
  fa fa_h_s_dadda_pg_rca32_fa729_out(h_s_dadda_pg_rca32_fa728_or0[0], h_s_dadda_pg_rca32_fa727_or0[0], h_s_dadda_pg_rca32_fa351_xor1[0], h_s_dadda_pg_rca32_fa729_xor1, h_s_dadda_pg_rca32_fa729_or0);
  fa fa_h_s_dadda_pg_rca32_fa730_out(h_s_dadda_pg_rca32_fa352_xor1[0], h_s_dadda_pg_rca32_fa353_xor1[0], h_s_dadda_pg_rca32_fa354_xor1[0], h_s_dadda_pg_rca32_fa730_xor1, h_s_dadda_pg_rca32_fa730_or0);
  fa fa_h_s_dadda_pg_rca32_fa731_out(h_s_dadda_pg_rca32_fa730_or0[0], h_s_dadda_pg_rca32_fa729_or0[0], h_s_dadda_pg_rca32_fa373_xor1[0], h_s_dadda_pg_rca32_fa731_xor1, h_s_dadda_pg_rca32_fa731_or0);
  fa fa_h_s_dadda_pg_rca32_fa732_out(h_s_dadda_pg_rca32_fa374_xor1[0], h_s_dadda_pg_rca32_fa375_xor1[0], h_s_dadda_pg_rca32_fa376_xor1[0], h_s_dadda_pg_rca32_fa732_xor1, h_s_dadda_pg_rca32_fa732_or0);
  fa fa_h_s_dadda_pg_rca32_fa733_out(h_s_dadda_pg_rca32_fa732_or0[0], h_s_dadda_pg_rca32_fa731_or0[0], h_s_dadda_pg_rca32_fa395_xor1[0], h_s_dadda_pg_rca32_fa733_xor1, h_s_dadda_pg_rca32_fa733_or0);
  fa fa_h_s_dadda_pg_rca32_fa734_out(h_s_dadda_pg_rca32_fa396_xor1[0], h_s_dadda_pg_rca32_fa397_xor1[0], h_s_dadda_pg_rca32_fa398_xor1[0], h_s_dadda_pg_rca32_fa734_xor1, h_s_dadda_pg_rca32_fa734_or0);
  fa fa_h_s_dadda_pg_rca32_fa735_out(h_s_dadda_pg_rca32_fa734_or0[0], h_s_dadda_pg_rca32_fa733_or0[0], h_s_dadda_pg_rca32_fa417_xor1[0], h_s_dadda_pg_rca32_fa735_xor1, h_s_dadda_pg_rca32_fa735_or0);
  fa fa_h_s_dadda_pg_rca32_fa736_out(h_s_dadda_pg_rca32_fa418_xor1[0], h_s_dadda_pg_rca32_fa419_xor1[0], h_s_dadda_pg_rca32_fa420_xor1[0], h_s_dadda_pg_rca32_fa736_xor1, h_s_dadda_pg_rca32_fa736_or0);
  fa fa_h_s_dadda_pg_rca32_fa737_out(h_s_dadda_pg_rca32_fa736_or0[0], h_s_dadda_pg_rca32_fa735_or0[0], h_s_dadda_pg_rca32_fa439_xor1[0], h_s_dadda_pg_rca32_fa737_xor1, h_s_dadda_pg_rca32_fa737_or0);
  fa fa_h_s_dadda_pg_rca32_fa738_out(h_s_dadda_pg_rca32_fa440_xor1[0], h_s_dadda_pg_rca32_fa441_xor1[0], h_s_dadda_pg_rca32_fa442_xor1[0], h_s_dadda_pg_rca32_fa738_xor1, h_s_dadda_pg_rca32_fa738_or0);
  fa fa_h_s_dadda_pg_rca32_fa739_out(h_s_dadda_pg_rca32_fa738_or0[0], h_s_dadda_pg_rca32_fa737_or0[0], h_s_dadda_pg_rca32_fa460_xor1[0], h_s_dadda_pg_rca32_fa739_xor1, h_s_dadda_pg_rca32_fa739_or0);
  fa fa_h_s_dadda_pg_rca32_fa740_out(h_s_dadda_pg_rca32_fa461_xor1[0], h_s_dadda_pg_rca32_fa462_xor1[0], h_s_dadda_pg_rca32_fa463_xor1[0], h_s_dadda_pg_rca32_fa740_xor1, h_s_dadda_pg_rca32_fa740_or0);
  fa fa_h_s_dadda_pg_rca32_fa741_out(h_s_dadda_pg_rca32_fa740_or0[0], h_s_dadda_pg_rca32_fa739_or0[0], h_s_dadda_pg_rca32_fa480_xor1[0], h_s_dadda_pg_rca32_fa741_xor1, h_s_dadda_pg_rca32_fa741_or0);
  fa fa_h_s_dadda_pg_rca32_fa742_out(h_s_dadda_pg_rca32_fa481_xor1[0], h_s_dadda_pg_rca32_fa482_xor1[0], h_s_dadda_pg_rca32_fa483_xor1[0], h_s_dadda_pg_rca32_fa742_xor1, h_s_dadda_pg_rca32_fa742_or0);
  fa fa_h_s_dadda_pg_rca32_fa743_out(h_s_dadda_pg_rca32_fa742_or0[0], h_s_dadda_pg_rca32_fa741_or0[0], h_s_dadda_pg_rca32_fa499_xor1[0], h_s_dadda_pg_rca32_fa743_xor1, h_s_dadda_pg_rca32_fa743_or0);
  fa fa_h_s_dadda_pg_rca32_fa744_out(h_s_dadda_pg_rca32_fa500_xor1[0], h_s_dadda_pg_rca32_fa501_xor1[0], h_s_dadda_pg_rca32_fa502_xor1[0], h_s_dadda_pg_rca32_fa744_xor1, h_s_dadda_pg_rca32_fa744_or0);
  fa fa_h_s_dadda_pg_rca32_fa745_out(h_s_dadda_pg_rca32_fa744_or0[0], h_s_dadda_pg_rca32_fa743_or0[0], h_s_dadda_pg_rca32_fa517_xor1[0], h_s_dadda_pg_rca32_fa745_xor1, h_s_dadda_pg_rca32_fa745_or0);
  fa fa_h_s_dadda_pg_rca32_fa746_out(h_s_dadda_pg_rca32_fa518_xor1[0], h_s_dadda_pg_rca32_fa519_xor1[0], h_s_dadda_pg_rca32_fa520_xor1[0], h_s_dadda_pg_rca32_fa746_xor1, h_s_dadda_pg_rca32_fa746_or0);
  fa fa_h_s_dadda_pg_rca32_fa747_out(h_s_dadda_pg_rca32_fa746_or0[0], h_s_dadda_pg_rca32_fa745_or0[0], h_s_dadda_pg_rca32_fa534_xor1[0], h_s_dadda_pg_rca32_fa747_xor1, h_s_dadda_pg_rca32_fa747_or0);
  fa fa_h_s_dadda_pg_rca32_fa748_out(h_s_dadda_pg_rca32_fa535_xor1[0], h_s_dadda_pg_rca32_fa536_xor1[0], h_s_dadda_pg_rca32_fa537_xor1[0], h_s_dadda_pg_rca32_fa748_xor1, h_s_dadda_pg_rca32_fa748_or0);
  fa fa_h_s_dadda_pg_rca32_fa749_out(h_s_dadda_pg_rca32_fa748_or0[0], h_s_dadda_pg_rca32_fa747_or0[0], h_s_dadda_pg_rca32_fa550_xor1[0], h_s_dadda_pg_rca32_fa749_xor1, h_s_dadda_pg_rca32_fa749_or0);
  fa fa_h_s_dadda_pg_rca32_fa750_out(h_s_dadda_pg_rca32_fa551_xor1[0], h_s_dadda_pg_rca32_fa552_xor1[0], h_s_dadda_pg_rca32_fa553_xor1[0], h_s_dadda_pg_rca32_fa750_xor1, h_s_dadda_pg_rca32_fa750_or0);
  fa fa_h_s_dadda_pg_rca32_fa751_out(h_s_dadda_pg_rca32_fa750_or0[0], h_s_dadda_pg_rca32_fa749_or0[0], h_s_dadda_pg_rca32_fa565_xor1[0], h_s_dadda_pg_rca32_fa751_xor1, h_s_dadda_pg_rca32_fa751_or0);
  fa fa_h_s_dadda_pg_rca32_fa752_out(h_s_dadda_pg_rca32_fa566_xor1[0], h_s_dadda_pg_rca32_fa567_xor1[0], h_s_dadda_pg_rca32_fa568_xor1[0], h_s_dadda_pg_rca32_fa752_xor1, h_s_dadda_pg_rca32_fa752_or0);
  fa fa_h_s_dadda_pg_rca32_fa753_out(h_s_dadda_pg_rca32_fa752_or0[0], h_s_dadda_pg_rca32_fa751_or0[0], h_s_dadda_pg_rca32_fa579_xor1[0], h_s_dadda_pg_rca32_fa753_xor1, h_s_dadda_pg_rca32_fa753_or0);
  fa fa_h_s_dadda_pg_rca32_fa754_out(h_s_dadda_pg_rca32_fa580_xor1[0], h_s_dadda_pg_rca32_fa581_xor1[0], h_s_dadda_pg_rca32_fa582_xor1[0], h_s_dadda_pg_rca32_fa754_xor1, h_s_dadda_pg_rca32_fa754_or0);
  fa fa_h_s_dadda_pg_rca32_fa755_out(h_s_dadda_pg_rca32_fa754_or0[0], h_s_dadda_pg_rca32_fa753_or0[0], h_s_dadda_pg_rca32_fa592_xor1[0], h_s_dadda_pg_rca32_fa755_xor1, h_s_dadda_pg_rca32_fa755_or0);
  fa fa_h_s_dadda_pg_rca32_fa756_out(h_s_dadda_pg_rca32_fa593_xor1[0], h_s_dadda_pg_rca32_fa594_xor1[0], h_s_dadda_pg_rca32_fa595_xor1[0], h_s_dadda_pg_rca32_fa756_xor1, h_s_dadda_pg_rca32_fa756_or0);
  fa fa_h_s_dadda_pg_rca32_fa757_out(h_s_dadda_pg_rca32_fa756_or0[0], h_s_dadda_pg_rca32_fa755_or0[0], h_s_dadda_pg_rca32_fa604_xor1[0], h_s_dadda_pg_rca32_fa757_xor1, h_s_dadda_pg_rca32_fa757_or0);
  fa fa_h_s_dadda_pg_rca32_fa758_out(h_s_dadda_pg_rca32_fa605_xor1[0], h_s_dadda_pg_rca32_fa606_xor1[0], h_s_dadda_pg_rca32_fa607_xor1[0], h_s_dadda_pg_rca32_fa758_xor1, h_s_dadda_pg_rca32_fa758_or0);
  fa fa_h_s_dadda_pg_rca32_fa759_out(h_s_dadda_pg_rca32_fa758_or0[0], h_s_dadda_pg_rca32_fa757_or0[0], h_s_dadda_pg_rca32_fa615_xor1[0], h_s_dadda_pg_rca32_fa759_xor1, h_s_dadda_pg_rca32_fa759_or0);
  fa fa_h_s_dadda_pg_rca32_fa760_out(h_s_dadda_pg_rca32_fa616_xor1[0], h_s_dadda_pg_rca32_fa617_xor1[0], h_s_dadda_pg_rca32_fa618_xor1[0], h_s_dadda_pg_rca32_fa760_xor1, h_s_dadda_pg_rca32_fa760_or0);
  fa fa_h_s_dadda_pg_rca32_fa761_out(h_s_dadda_pg_rca32_fa760_or0[0], h_s_dadda_pg_rca32_fa759_or0[0], h_s_dadda_pg_rca32_fa625_xor1[0], h_s_dadda_pg_rca32_fa761_xor1, h_s_dadda_pg_rca32_fa761_or0);
  fa fa_h_s_dadda_pg_rca32_fa762_out(h_s_dadda_pg_rca32_fa626_xor1[0], h_s_dadda_pg_rca32_fa627_xor1[0], h_s_dadda_pg_rca32_fa628_xor1[0], h_s_dadda_pg_rca32_fa762_xor1, h_s_dadda_pg_rca32_fa762_or0);
  fa fa_h_s_dadda_pg_rca32_fa763_out(h_s_dadda_pg_rca32_fa762_or0[0], h_s_dadda_pg_rca32_fa761_or0[0], h_s_dadda_pg_rca32_fa634_xor1[0], h_s_dadda_pg_rca32_fa763_xor1, h_s_dadda_pg_rca32_fa763_or0);
  fa fa_h_s_dadda_pg_rca32_fa764_out(h_s_dadda_pg_rca32_fa635_xor1[0], h_s_dadda_pg_rca32_fa636_xor1[0], h_s_dadda_pg_rca32_fa637_xor1[0], h_s_dadda_pg_rca32_fa764_xor1, h_s_dadda_pg_rca32_fa764_or0);
  fa fa_h_s_dadda_pg_rca32_fa765_out(h_s_dadda_pg_rca32_fa764_or0[0], h_s_dadda_pg_rca32_fa763_or0[0], h_s_dadda_pg_rca32_fa642_xor1[0], h_s_dadda_pg_rca32_fa765_xor1, h_s_dadda_pg_rca32_fa765_or0);
  fa fa_h_s_dadda_pg_rca32_fa766_out(h_s_dadda_pg_rca32_fa643_xor1[0], h_s_dadda_pg_rca32_fa644_xor1[0], h_s_dadda_pg_rca32_fa645_xor1[0], h_s_dadda_pg_rca32_fa766_xor1, h_s_dadda_pg_rca32_fa766_or0);
  fa fa_h_s_dadda_pg_rca32_fa767_out(h_s_dadda_pg_rca32_fa766_or0[0], h_s_dadda_pg_rca32_fa765_or0[0], h_s_dadda_pg_rca32_fa649_xor1[0], h_s_dadda_pg_rca32_fa767_xor1, h_s_dadda_pg_rca32_fa767_or0);
  fa fa_h_s_dadda_pg_rca32_fa768_out(h_s_dadda_pg_rca32_fa650_xor1[0], h_s_dadda_pg_rca32_fa651_xor1[0], h_s_dadda_pg_rca32_fa652_xor1[0], h_s_dadda_pg_rca32_fa768_xor1, h_s_dadda_pg_rca32_fa768_or0);
  fa fa_h_s_dadda_pg_rca32_fa769_out(h_s_dadda_pg_rca32_fa768_or0[0], h_s_dadda_pg_rca32_fa767_or0[0], h_s_dadda_pg_rca32_fa655_xor1[0], h_s_dadda_pg_rca32_fa769_xor1, h_s_dadda_pg_rca32_fa769_or0);
  fa fa_h_s_dadda_pg_rca32_fa770_out(h_s_dadda_pg_rca32_fa656_xor1[0], h_s_dadda_pg_rca32_fa657_xor1[0], h_s_dadda_pg_rca32_fa658_xor1[0], h_s_dadda_pg_rca32_fa770_xor1, h_s_dadda_pg_rca32_fa770_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_22_31(a[22], b[31], h_s_dadda_pg_rca32_nand_22_31);
  fa fa_h_s_dadda_pg_rca32_fa771_out(h_s_dadda_pg_rca32_fa770_or0[0], h_s_dadda_pg_rca32_fa769_or0[0], h_s_dadda_pg_rca32_nand_22_31[0], h_s_dadda_pg_rca32_fa771_xor1, h_s_dadda_pg_rca32_fa771_or0);
  fa fa_h_s_dadda_pg_rca32_fa772_out(h_s_dadda_pg_rca32_fa661_xor1[0], h_s_dadda_pg_rca32_fa662_xor1[0], h_s_dadda_pg_rca32_fa663_xor1[0], h_s_dadda_pg_rca32_fa772_xor1, h_s_dadda_pg_rca32_fa772_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_24_30(a[24], b[30], h_s_dadda_pg_rca32_and_24_30);
  fa fa_h_s_dadda_pg_rca32_fa773_out(h_s_dadda_pg_rca32_fa772_or0[0], h_s_dadda_pg_rca32_fa771_or0[0], h_s_dadda_pg_rca32_and_24_30[0], h_s_dadda_pg_rca32_fa773_xor1, h_s_dadda_pg_rca32_fa773_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_23_31(a[23], b[31], h_s_dadda_pg_rca32_nand_23_31);
  fa fa_h_s_dadda_pg_rca32_fa774_out(h_s_dadda_pg_rca32_nand_23_31[0], h_s_dadda_pg_rca32_fa666_xor1[0], h_s_dadda_pg_rca32_fa667_xor1[0], h_s_dadda_pg_rca32_fa774_xor1, h_s_dadda_pg_rca32_fa774_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_29(a[26], b[29], h_s_dadda_pg_rca32_and_26_29);
  fa fa_h_s_dadda_pg_rca32_fa775_out(h_s_dadda_pg_rca32_fa774_or0[0], h_s_dadda_pg_rca32_fa773_or0[0], h_s_dadda_pg_rca32_and_26_29[0], h_s_dadda_pg_rca32_fa775_xor1, h_s_dadda_pg_rca32_fa775_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_25_30(a[25], b[30], h_s_dadda_pg_rca32_and_25_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_24_31(a[24], b[31], h_s_dadda_pg_rca32_nand_24_31);
  fa fa_h_s_dadda_pg_rca32_fa776_out(h_s_dadda_pg_rca32_and_25_30[0], h_s_dadda_pg_rca32_nand_24_31[0], h_s_dadda_pg_rca32_fa670_xor1[0], h_s_dadda_pg_rca32_fa776_xor1, h_s_dadda_pg_rca32_fa776_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_28(a[28], b[28], h_s_dadda_pg_rca32_and_28_28);
  fa fa_h_s_dadda_pg_rca32_fa777_out(h_s_dadda_pg_rca32_fa776_or0[0], h_s_dadda_pg_rca32_fa775_or0[0], h_s_dadda_pg_rca32_and_28_28[0], h_s_dadda_pg_rca32_fa777_xor1, h_s_dadda_pg_rca32_fa777_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_29(a[27], b[29], h_s_dadda_pg_rca32_and_27_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_26_30(a[26], b[30], h_s_dadda_pg_rca32_and_26_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_25_31(a[25], b[31], h_s_dadda_pg_rca32_nand_25_31);
  fa fa_h_s_dadda_pg_rca32_fa778_out(h_s_dadda_pg_rca32_and_27_29[0], h_s_dadda_pg_rca32_and_26_30[0], h_s_dadda_pg_rca32_nand_25_31[0], h_s_dadda_pg_rca32_fa778_xor1, h_s_dadda_pg_rca32_fa778_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_27(a[30], b[27], h_s_dadda_pg_rca32_and_30_27);
  fa fa_h_s_dadda_pg_rca32_fa779_out(h_s_dadda_pg_rca32_fa778_or0[0], h_s_dadda_pg_rca32_fa777_or0[0], h_s_dadda_pg_rca32_and_30_27[0], h_s_dadda_pg_rca32_fa779_xor1, h_s_dadda_pg_rca32_fa779_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_28(a[29], b[28], h_s_dadda_pg_rca32_and_29_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_29(a[28], b[29], h_s_dadda_pg_rca32_and_28_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_27_30(a[27], b[30], h_s_dadda_pg_rca32_and_27_30);
  fa fa_h_s_dadda_pg_rca32_fa780_out(h_s_dadda_pg_rca32_and_29_28[0], h_s_dadda_pg_rca32_and_28_29[0], h_s_dadda_pg_rca32_and_27_30[0], h_s_dadda_pg_rca32_fa780_xor1, h_s_dadda_pg_rca32_fa780_or0);
  fa fa_h_s_dadda_pg_rca32_fa781_out(h_s_dadda_pg_rca32_fa780_or0[0], h_s_dadda_pg_rca32_fa779_or0[0], h_s_dadda_pg_rca32_fa675_or0[0], h_s_dadda_pg_rca32_fa781_xor1, h_s_dadda_pg_rca32_fa781_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_27(a[31], b[27], h_s_dadda_pg_rca32_nand_31_27);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_28(a[30], b[28], h_s_dadda_pg_rca32_and_30_28);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_29(a[29], b[29], h_s_dadda_pg_rca32_and_29_29);
  fa fa_h_s_dadda_pg_rca32_fa782_out(h_s_dadda_pg_rca32_nand_31_27[0], h_s_dadda_pg_rca32_and_30_28[0], h_s_dadda_pg_rca32_and_29_29[0], h_s_dadda_pg_rca32_fa782_xor1, h_s_dadda_pg_rca32_fa782_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_28(a[31], b[28], h_s_dadda_pg_rca32_nand_31_28);
  fa fa_h_s_dadda_pg_rca32_fa783_out(h_s_dadda_pg_rca32_fa782_or0[0], h_s_dadda_pg_rca32_fa781_or0[0], h_s_dadda_pg_rca32_nand_31_28[0], h_s_dadda_pg_rca32_fa783_xor1, h_s_dadda_pg_rca32_fa783_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_3_0(a[3], b[0], h_s_dadda_pg_rca32_and_3_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_1(a[2], b[1], h_s_dadda_pg_rca32_and_2_1);
  ha ha_h_s_dadda_pg_rca32_ha28_out(h_s_dadda_pg_rca32_and_3_0[0], h_s_dadda_pg_rca32_and_2_1[0], h_s_dadda_pg_rca32_ha28_xor0, h_s_dadda_pg_rca32_ha28_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_2(a[2], b[2], h_s_dadda_pg_rca32_and_2_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_3(a[1], b[3], h_s_dadda_pg_rca32_and_1_3);
  fa fa_h_s_dadda_pg_rca32_fa784_out(h_s_dadda_pg_rca32_ha28_and0[0], h_s_dadda_pg_rca32_and_2_2[0], h_s_dadda_pg_rca32_and_1_3[0], h_s_dadda_pg_rca32_fa784_xor1, h_s_dadda_pg_rca32_fa784_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_4(a[1], b[4], h_s_dadda_pg_rca32_and_1_4);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_5(a[0], b[5], h_s_dadda_pg_rca32_and_0_5);
  fa fa_h_s_dadda_pg_rca32_fa785_out(h_s_dadda_pg_rca32_fa784_or0[0], h_s_dadda_pg_rca32_and_1_4[0], h_s_dadda_pg_rca32_and_0_5[0], h_s_dadda_pg_rca32_fa785_xor1, h_s_dadda_pg_rca32_fa785_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_6(a[0], b[6], h_s_dadda_pg_rca32_and_0_6);
  fa fa_h_s_dadda_pg_rca32_fa786_out(h_s_dadda_pg_rca32_fa785_or0[0], h_s_dadda_pg_rca32_and_0_6[0], h_s_dadda_pg_rca32_ha4_xor0[0], h_s_dadda_pg_rca32_fa786_xor1, h_s_dadda_pg_rca32_fa786_or0);
  fa fa_h_s_dadda_pg_rca32_fa787_out(h_s_dadda_pg_rca32_fa786_or0[0], h_s_dadda_pg_rca32_fa16_xor1[0], h_s_dadda_pg_rca32_ha5_xor0[0], h_s_dadda_pg_rca32_fa787_xor1, h_s_dadda_pg_rca32_fa787_or0);
  fa fa_h_s_dadda_pg_rca32_fa788_out(h_s_dadda_pg_rca32_fa787_or0[0], h_s_dadda_pg_rca32_fa18_xor1[0], h_s_dadda_pg_rca32_ha6_xor0[0], h_s_dadda_pg_rca32_fa788_xor1, h_s_dadda_pg_rca32_fa788_or0);
  fa fa_h_s_dadda_pg_rca32_fa789_out(h_s_dadda_pg_rca32_fa788_or0[0], h_s_dadda_pg_rca32_fa21_xor1[0], h_s_dadda_pg_rca32_ha7_xor0[0], h_s_dadda_pg_rca32_fa789_xor1, h_s_dadda_pg_rca32_fa789_or0);
  fa fa_h_s_dadda_pg_rca32_fa790_out(h_s_dadda_pg_rca32_fa789_or0[0], h_s_dadda_pg_rca32_fa25_xor1[0], h_s_dadda_pg_rca32_ha8_xor0[0], h_s_dadda_pg_rca32_fa790_xor1, h_s_dadda_pg_rca32_fa790_or0);
  fa fa_h_s_dadda_pg_rca32_fa791_out(h_s_dadda_pg_rca32_fa790_or0[0], h_s_dadda_pg_rca32_fa30_xor1[0], h_s_dadda_pg_rca32_ha9_xor0[0], h_s_dadda_pg_rca32_fa791_xor1, h_s_dadda_pg_rca32_fa791_or0);
  fa fa_h_s_dadda_pg_rca32_fa792_out(h_s_dadda_pg_rca32_fa791_or0[0], h_s_dadda_pg_rca32_fa36_xor1[0], h_s_dadda_pg_rca32_ha10_xor0[0], h_s_dadda_pg_rca32_fa792_xor1, h_s_dadda_pg_rca32_fa792_or0);
  fa fa_h_s_dadda_pg_rca32_fa793_out(h_s_dadda_pg_rca32_fa792_or0[0], h_s_dadda_pg_rca32_fa43_xor1[0], h_s_dadda_pg_rca32_ha11_xor0[0], h_s_dadda_pg_rca32_fa793_xor1, h_s_dadda_pg_rca32_fa793_or0);
  fa fa_h_s_dadda_pg_rca32_fa794_out(h_s_dadda_pg_rca32_fa793_or0[0], h_s_dadda_pg_rca32_fa51_xor1[0], h_s_dadda_pg_rca32_ha12_xor0[0], h_s_dadda_pg_rca32_fa794_xor1, h_s_dadda_pg_rca32_fa794_or0);
  fa fa_h_s_dadda_pg_rca32_fa795_out(h_s_dadda_pg_rca32_fa794_or0[0], h_s_dadda_pg_rca32_fa60_xor1[0], h_s_dadda_pg_rca32_ha13_xor0[0], h_s_dadda_pg_rca32_fa795_xor1, h_s_dadda_pg_rca32_fa795_or0);
  fa fa_h_s_dadda_pg_rca32_fa796_out(h_s_dadda_pg_rca32_fa795_or0[0], h_s_dadda_pg_rca32_fa70_xor1[0], h_s_dadda_pg_rca32_ha14_xor0[0], h_s_dadda_pg_rca32_fa796_xor1, h_s_dadda_pg_rca32_fa796_or0);
  fa fa_h_s_dadda_pg_rca32_fa797_out(h_s_dadda_pg_rca32_fa796_or0[0], h_s_dadda_pg_rca32_fa81_xor1[0], h_s_dadda_pg_rca32_ha15_xor0[0], h_s_dadda_pg_rca32_fa797_xor1, h_s_dadda_pg_rca32_fa797_or0);
  fa fa_h_s_dadda_pg_rca32_fa798_out(h_s_dadda_pg_rca32_fa797_or0[0], h_s_dadda_pg_rca32_fa93_xor1[0], h_s_dadda_pg_rca32_ha16_xor0[0], h_s_dadda_pg_rca32_fa798_xor1, h_s_dadda_pg_rca32_fa798_or0);
  fa fa_h_s_dadda_pg_rca32_fa799_out(h_s_dadda_pg_rca32_fa798_or0[0], h_s_dadda_pg_rca32_fa106_xor1[0], h_s_dadda_pg_rca32_ha17_xor0[0], h_s_dadda_pg_rca32_fa799_xor1, h_s_dadda_pg_rca32_fa799_or0);
  fa fa_h_s_dadda_pg_rca32_fa800_out(h_s_dadda_pg_rca32_fa799_or0[0], h_s_dadda_pg_rca32_fa120_xor1[0], h_s_dadda_pg_rca32_ha18_xor0[0], h_s_dadda_pg_rca32_fa800_xor1, h_s_dadda_pg_rca32_fa800_or0);
  fa fa_h_s_dadda_pg_rca32_fa801_out(h_s_dadda_pg_rca32_fa800_or0[0], h_s_dadda_pg_rca32_fa135_xor1[0], h_s_dadda_pg_rca32_ha19_xor0[0], h_s_dadda_pg_rca32_fa801_xor1, h_s_dadda_pg_rca32_fa801_or0);
  fa fa_h_s_dadda_pg_rca32_fa802_out(h_s_dadda_pg_rca32_fa801_or0[0], h_s_dadda_pg_rca32_fa151_xor1[0], h_s_dadda_pg_rca32_ha20_xor0[0], h_s_dadda_pg_rca32_fa802_xor1, h_s_dadda_pg_rca32_fa802_or0);
  fa fa_h_s_dadda_pg_rca32_fa803_out(h_s_dadda_pg_rca32_fa802_or0[0], h_s_dadda_pg_rca32_fa168_xor1[0], h_s_dadda_pg_rca32_ha21_xor0[0], h_s_dadda_pg_rca32_fa803_xor1, h_s_dadda_pg_rca32_fa803_or0);
  fa fa_h_s_dadda_pg_rca32_fa804_out(h_s_dadda_pg_rca32_fa803_or0[0], h_s_dadda_pg_rca32_fa186_xor1[0], h_s_dadda_pg_rca32_ha22_xor0[0], h_s_dadda_pg_rca32_fa804_xor1, h_s_dadda_pg_rca32_fa804_or0);
  fa fa_h_s_dadda_pg_rca32_fa805_out(h_s_dadda_pg_rca32_fa804_or0[0], h_s_dadda_pg_rca32_fa205_xor1[0], h_s_dadda_pg_rca32_ha23_xor0[0], h_s_dadda_pg_rca32_fa805_xor1, h_s_dadda_pg_rca32_fa805_or0);
  fa fa_h_s_dadda_pg_rca32_fa806_out(h_s_dadda_pg_rca32_fa805_or0[0], h_s_dadda_pg_rca32_fa225_xor1[0], h_s_dadda_pg_rca32_ha24_xor0[0], h_s_dadda_pg_rca32_fa806_xor1, h_s_dadda_pg_rca32_fa806_or0);
  fa fa_h_s_dadda_pg_rca32_fa807_out(h_s_dadda_pg_rca32_fa806_or0[0], h_s_dadda_pg_rca32_fa246_xor1[0], h_s_dadda_pg_rca32_ha25_xor0[0], h_s_dadda_pg_rca32_fa807_xor1, h_s_dadda_pg_rca32_fa807_or0);
  fa fa_h_s_dadda_pg_rca32_fa808_out(h_s_dadda_pg_rca32_fa807_or0[0], h_s_dadda_pg_rca32_fa267_xor1[0], h_s_dadda_pg_rca32_fa268_xor1[0], h_s_dadda_pg_rca32_fa808_xor1, h_s_dadda_pg_rca32_fa808_or0);
  fa fa_h_s_dadda_pg_rca32_fa809_out(h_s_dadda_pg_rca32_fa808_or0[0], h_s_dadda_pg_rca32_fa289_xor1[0], h_s_dadda_pg_rca32_fa290_xor1[0], h_s_dadda_pg_rca32_fa809_xor1, h_s_dadda_pg_rca32_fa809_or0);
  fa fa_h_s_dadda_pg_rca32_fa810_out(h_s_dadda_pg_rca32_fa809_or0[0], h_s_dadda_pg_rca32_fa311_xor1[0], h_s_dadda_pg_rca32_fa312_xor1[0], h_s_dadda_pg_rca32_fa810_xor1, h_s_dadda_pg_rca32_fa810_or0);
  fa fa_h_s_dadda_pg_rca32_fa811_out(h_s_dadda_pg_rca32_fa810_or0[0], h_s_dadda_pg_rca32_fa333_xor1[0], h_s_dadda_pg_rca32_fa334_xor1[0], h_s_dadda_pg_rca32_fa811_xor1, h_s_dadda_pg_rca32_fa811_or0);
  fa fa_h_s_dadda_pg_rca32_fa812_out(h_s_dadda_pg_rca32_fa811_or0[0], h_s_dadda_pg_rca32_fa355_xor1[0], h_s_dadda_pg_rca32_fa356_xor1[0], h_s_dadda_pg_rca32_fa812_xor1, h_s_dadda_pg_rca32_fa812_or0);
  fa fa_h_s_dadda_pg_rca32_fa813_out(h_s_dadda_pg_rca32_fa812_or0[0], h_s_dadda_pg_rca32_fa377_xor1[0], h_s_dadda_pg_rca32_fa378_xor1[0], h_s_dadda_pg_rca32_fa813_xor1, h_s_dadda_pg_rca32_fa813_or0);
  fa fa_h_s_dadda_pg_rca32_fa814_out(h_s_dadda_pg_rca32_fa813_or0[0], h_s_dadda_pg_rca32_fa399_xor1[0], h_s_dadda_pg_rca32_fa400_xor1[0], h_s_dadda_pg_rca32_fa814_xor1, h_s_dadda_pg_rca32_fa814_or0);
  fa fa_h_s_dadda_pg_rca32_fa815_out(h_s_dadda_pg_rca32_fa814_or0[0], h_s_dadda_pg_rca32_fa421_xor1[0], h_s_dadda_pg_rca32_fa422_xor1[0], h_s_dadda_pg_rca32_fa815_xor1, h_s_dadda_pg_rca32_fa815_or0);
  fa fa_h_s_dadda_pg_rca32_fa816_out(h_s_dadda_pg_rca32_fa815_or0[0], h_s_dadda_pg_rca32_fa443_xor1[0], h_s_dadda_pg_rca32_fa444_xor1[0], h_s_dadda_pg_rca32_fa816_xor1, h_s_dadda_pg_rca32_fa816_or0);
  fa fa_h_s_dadda_pg_rca32_fa817_out(h_s_dadda_pg_rca32_fa816_or0[0], h_s_dadda_pg_rca32_fa464_xor1[0], h_s_dadda_pg_rca32_fa465_xor1[0], h_s_dadda_pg_rca32_fa817_xor1, h_s_dadda_pg_rca32_fa817_or0);
  fa fa_h_s_dadda_pg_rca32_fa818_out(h_s_dadda_pg_rca32_fa817_or0[0], h_s_dadda_pg_rca32_fa484_xor1[0], h_s_dadda_pg_rca32_fa485_xor1[0], h_s_dadda_pg_rca32_fa818_xor1, h_s_dadda_pg_rca32_fa818_or0);
  fa fa_h_s_dadda_pg_rca32_fa819_out(h_s_dadda_pg_rca32_fa818_or0[0], h_s_dadda_pg_rca32_fa503_xor1[0], h_s_dadda_pg_rca32_fa504_xor1[0], h_s_dadda_pg_rca32_fa819_xor1, h_s_dadda_pg_rca32_fa819_or0);
  fa fa_h_s_dadda_pg_rca32_fa820_out(h_s_dadda_pg_rca32_fa819_or0[0], h_s_dadda_pg_rca32_fa521_xor1[0], h_s_dadda_pg_rca32_fa522_xor1[0], h_s_dadda_pg_rca32_fa820_xor1, h_s_dadda_pg_rca32_fa820_or0);
  fa fa_h_s_dadda_pg_rca32_fa821_out(h_s_dadda_pg_rca32_fa820_or0[0], h_s_dadda_pg_rca32_fa538_xor1[0], h_s_dadda_pg_rca32_fa539_xor1[0], h_s_dadda_pg_rca32_fa821_xor1, h_s_dadda_pg_rca32_fa821_or0);
  fa fa_h_s_dadda_pg_rca32_fa822_out(h_s_dadda_pg_rca32_fa821_or0[0], h_s_dadda_pg_rca32_fa554_xor1[0], h_s_dadda_pg_rca32_fa555_xor1[0], h_s_dadda_pg_rca32_fa822_xor1, h_s_dadda_pg_rca32_fa822_or0);
  fa fa_h_s_dadda_pg_rca32_fa823_out(h_s_dadda_pg_rca32_fa822_or0[0], h_s_dadda_pg_rca32_fa569_xor1[0], h_s_dadda_pg_rca32_fa570_xor1[0], h_s_dadda_pg_rca32_fa823_xor1, h_s_dadda_pg_rca32_fa823_or0);
  fa fa_h_s_dadda_pg_rca32_fa824_out(h_s_dadda_pg_rca32_fa823_or0[0], h_s_dadda_pg_rca32_fa583_xor1[0], h_s_dadda_pg_rca32_fa584_xor1[0], h_s_dadda_pg_rca32_fa824_xor1, h_s_dadda_pg_rca32_fa824_or0);
  fa fa_h_s_dadda_pg_rca32_fa825_out(h_s_dadda_pg_rca32_fa824_or0[0], h_s_dadda_pg_rca32_fa596_xor1[0], h_s_dadda_pg_rca32_fa597_xor1[0], h_s_dadda_pg_rca32_fa825_xor1, h_s_dadda_pg_rca32_fa825_or0);
  fa fa_h_s_dadda_pg_rca32_fa826_out(h_s_dadda_pg_rca32_fa825_or0[0], h_s_dadda_pg_rca32_fa608_xor1[0], h_s_dadda_pg_rca32_fa609_xor1[0], h_s_dadda_pg_rca32_fa826_xor1, h_s_dadda_pg_rca32_fa826_or0);
  fa fa_h_s_dadda_pg_rca32_fa827_out(h_s_dadda_pg_rca32_fa826_or0[0], h_s_dadda_pg_rca32_fa619_xor1[0], h_s_dadda_pg_rca32_fa620_xor1[0], h_s_dadda_pg_rca32_fa827_xor1, h_s_dadda_pg_rca32_fa827_or0);
  fa fa_h_s_dadda_pg_rca32_fa828_out(h_s_dadda_pg_rca32_fa827_or0[0], h_s_dadda_pg_rca32_fa629_xor1[0], h_s_dadda_pg_rca32_fa630_xor1[0], h_s_dadda_pg_rca32_fa828_xor1, h_s_dadda_pg_rca32_fa828_or0);
  fa fa_h_s_dadda_pg_rca32_fa829_out(h_s_dadda_pg_rca32_fa828_or0[0], h_s_dadda_pg_rca32_fa638_xor1[0], h_s_dadda_pg_rca32_fa639_xor1[0], h_s_dadda_pg_rca32_fa829_xor1, h_s_dadda_pg_rca32_fa829_or0);
  fa fa_h_s_dadda_pg_rca32_fa830_out(h_s_dadda_pg_rca32_fa829_or0[0], h_s_dadda_pg_rca32_fa646_xor1[0], h_s_dadda_pg_rca32_fa647_xor1[0], h_s_dadda_pg_rca32_fa830_xor1, h_s_dadda_pg_rca32_fa830_or0);
  fa fa_h_s_dadda_pg_rca32_fa831_out(h_s_dadda_pg_rca32_fa830_or0[0], h_s_dadda_pg_rca32_fa653_xor1[0], h_s_dadda_pg_rca32_fa654_xor1[0], h_s_dadda_pg_rca32_fa831_xor1, h_s_dadda_pg_rca32_fa831_or0);
  fa fa_h_s_dadda_pg_rca32_fa832_out(h_s_dadda_pg_rca32_fa831_or0[0], h_s_dadda_pg_rca32_fa659_xor1[0], h_s_dadda_pg_rca32_fa660_xor1[0], h_s_dadda_pg_rca32_fa832_xor1, h_s_dadda_pg_rca32_fa832_or0);
  fa fa_h_s_dadda_pg_rca32_fa833_out(h_s_dadda_pg_rca32_fa832_or0[0], h_s_dadda_pg_rca32_fa664_xor1[0], h_s_dadda_pg_rca32_fa665_xor1[0], h_s_dadda_pg_rca32_fa833_xor1, h_s_dadda_pg_rca32_fa833_or0);
  fa fa_h_s_dadda_pg_rca32_fa834_out(h_s_dadda_pg_rca32_fa833_or0[0], h_s_dadda_pg_rca32_fa668_xor1[0], h_s_dadda_pg_rca32_fa669_xor1[0], h_s_dadda_pg_rca32_fa834_xor1, h_s_dadda_pg_rca32_fa834_or0);
  fa fa_h_s_dadda_pg_rca32_fa835_out(h_s_dadda_pg_rca32_fa834_or0[0], h_s_dadda_pg_rca32_fa671_xor1[0], h_s_dadda_pg_rca32_fa672_xor1[0], h_s_dadda_pg_rca32_fa835_xor1, h_s_dadda_pg_rca32_fa835_or0);
  fa fa_h_s_dadda_pg_rca32_fa836_out(h_s_dadda_pg_rca32_fa835_or0[0], h_s_dadda_pg_rca32_fa673_xor1[0], h_s_dadda_pg_rca32_fa674_xor1[0], h_s_dadda_pg_rca32_fa836_xor1, h_s_dadda_pg_rca32_fa836_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_26_31(a[26], b[31], h_s_dadda_pg_rca32_nand_26_31);
  fa fa_h_s_dadda_pg_rca32_fa837_out(h_s_dadda_pg_rca32_fa836_or0[0], h_s_dadda_pg_rca32_nand_26_31[0], h_s_dadda_pg_rca32_fa675_xor1[0], h_s_dadda_pg_rca32_fa837_xor1, h_s_dadda_pg_rca32_fa837_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_28_30(a[28], b[30], h_s_dadda_pg_rca32_and_28_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_27_31(a[27], b[31], h_s_dadda_pg_rca32_nand_27_31);
  fa fa_h_s_dadda_pg_rca32_fa838_out(h_s_dadda_pg_rca32_fa837_or0[0], h_s_dadda_pg_rca32_and_28_30[0], h_s_dadda_pg_rca32_nand_27_31[0], h_s_dadda_pg_rca32_fa838_xor1, h_s_dadda_pg_rca32_fa838_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_29(a[30], b[29], h_s_dadda_pg_rca32_and_30_29);
  and_gate and_gate_h_s_dadda_pg_rca32_and_29_30(a[29], b[30], h_s_dadda_pg_rca32_and_29_30);
  fa fa_h_s_dadda_pg_rca32_fa839_out(h_s_dadda_pg_rca32_fa838_or0[0], h_s_dadda_pg_rca32_and_30_29[0], h_s_dadda_pg_rca32_and_29_30[0], h_s_dadda_pg_rca32_fa839_xor1, h_s_dadda_pg_rca32_fa839_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_29(a[31], b[29], h_s_dadda_pg_rca32_nand_31_29);
  fa fa_h_s_dadda_pg_rca32_fa840_out(h_s_dadda_pg_rca32_fa839_or0[0], h_s_dadda_pg_rca32_fa783_or0[0], h_s_dadda_pg_rca32_nand_31_29[0], h_s_dadda_pg_rca32_fa840_xor1, h_s_dadda_pg_rca32_fa840_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_2_0(a[2], b[0], h_s_dadda_pg_rca32_and_2_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_1(a[1], b[1], h_s_dadda_pg_rca32_and_1_1);
  ha ha_h_s_dadda_pg_rca32_ha29_out(h_s_dadda_pg_rca32_and_2_0[0], h_s_dadda_pg_rca32_and_1_1[0], h_s_dadda_pg_rca32_ha29_xor0, h_s_dadda_pg_rca32_ha29_and0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_2(a[1], b[2], h_s_dadda_pg_rca32_and_1_2);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_3(a[0], b[3], h_s_dadda_pg_rca32_and_0_3);
  fa fa_h_s_dadda_pg_rca32_fa841_out(h_s_dadda_pg_rca32_ha29_and0[0], h_s_dadda_pg_rca32_and_1_2[0], h_s_dadda_pg_rca32_and_0_3[0], h_s_dadda_pg_rca32_fa841_xor1, h_s_dadda_pg_rca32_fa841_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_4(a[0], b[4], h_s_dadda_pg_rca32_and_0_4);
  fa fa_h_s_dadda_pg_rca32_fa842_out(h_s_dadda_pg_rca32_fa841_or0[0], h_s_dadda_pg_rca32_and_0_4[0], h_s_dadda_pg_rca32_ha26_xor0[0], h_s_dadda_pg_rca32_fa842_xor1, h_s_dadda_pg_rca32_fa842_or0);
  fa fa_h_s_dadda_pg_rca32_fa843_out(h_s_dadda_pg_rca32_fa842_or0[0], h_s_dadda_pg_rca32_fa676_xor1[0], h_s_dadda_pg_rca32_ha27_xor0[0], h_s_dadda_pg_rca32_fa843_xor1, h_s_dadda_pg_rca32_fa843_or0);
  fa fa_h_s_dadda_pg_rca32_fa844_out(h_s_dadda_pg_rca32_fa843_or0[0], h_s_dadda_pg_rca32_fa677_xor1[0], h_s_dadda_pg_rca32_fa678_xor1[0], h_s_dadda_pg_rca32_fa844_xor1, h_s_dadda_pg_rca32_fa844_or0);
  fa fa_h_s_dadda_pg_rca32_fa845_out(h_s_dadda_pg_rca32_fa844_or0[0], h_s_dadda_pg_rca32_fa679_xor1[0], h_s_dadda_pg_rca32_fa680_xor1[0], h_s_dadda_pg_rca32_fa845_xor1, h_s_dadda_pg_rca32_fa845_or0);
  fa fa_h_s_dadda_pg_rca32_fa846_out(h_s_dadda_pg_rca32_fa845_or0[0], h_s_dadda_pg_rca32_fa681_xor1[0], h_s_dadda_pg_rca32_fa682_xor1[0], h_s_dadda_pg_rca32_fa846_xor1, h_s_dadda_pg_rca32_fa846_or0);
  fa fa_h_s_dadda_pg_rca32_fa847_out(h_s_dadda_pg_rca32_fa846_or0[0], h_s_dadda_pg_rca32_fa683_xor1[0], h_s_dadda_pg_rca32_fa684_xor1[0], h_s_dadda_pg_rca32_fa847_xor1, h_s_dadda_pg_rca32_fa847_or0);
  fa fa_h_s_dadda_pg_rca32_fa848_out(h_s_dadda_pg_rca32_fa847_or0[0], h_s_dadda_pg_rca32_fa685_xor1[0], h_s_dadda_pg_rca32_fa686_xor1[0], h_s_dadda_pg_rca32_fa848_xor1, h_s_dadda_pg_rca32_fa848_or0);
  fa fa_h_s_dadda_pg_rca32_fa849_out(h_s_dadda_pg_rca32_fa848_or0[0], h_s_dadda_pg_rca32_fa687_xor1[0], h_s_dadda_pg_rca32_fa688_xor1[0], h_s_dadda_pg_rca32_fa849_xor1, h_s_dadda_pg_rca32_fa849_or0);
  fa fa_h_s_dadda_pg_rca32_fa850_out(h_s_dadda_pg_rca32_fa849_or0[0], h_s_dadda_pg_rca32_fa689_xor1[0], h_s_dadda_pg_rca32_fa690_xor1[0], h_s_dadda_pg_rca32_fa850_xor1, h_s_dadda_pg_rca32_fa850_or0);
  fa fa_h_s_dadda_pg_rca32_fa851_out(h_s_dadda_pg_rca32_fa850_or0[0], h_s_dadda_pg_rca32_fa691_xor1[0], h_s_dadda_pg_rca32_fa692_xor1[0], h_s_dadda_pg_rca32_fa851_xor1, h_s_dadda_pg_rca32_fa851_or0);
  fa fa_h_s_dadda_pg_rca32_fa852_out(h_s_dadda_pg_rca32_fa851_or0[0], h_s_dadda_pg_rca32_fa693_xor1[0], h_s_dadda_pg_rca32_fa694_xor1[0], h_s_dadda_pg_rca32_fa852_xor1, h_s_dadda_pg_rca32_fa852_or0);
  fa fa_h_s_dadda_pg_rca32_fa853_out(h_s_dadda_pg_rca32_fa852_or0[0], h_s_dadda_pg_rca32_fa695_xor1[0], h_s_dadda_pg_rca32_fa696_xor1[0], h_s_dadda_pg_rca32_fa853_xor1, h_s_dadda_pg_rca32_fa853_or0);
  fa fa_h_s_dadda_pg_rca32_fa854_out(h_s_dadda_pg_rca32_fa853_or0[0], h_s_dadda_pg_rca32_fa697_xor1[0], h_s_dadda_pg_rca32_fa698_xor1[0], h_s_dadda_pg_rca32_fa854_xor1, h_s_dadda_pg_rca32_fa854_or0);
  fa fa_h_s_dadda_pg_rca32_fa855_out(h_s_dadda_pg_rca32_fa854_or0[0], h_s_dadda_pg_rca32_fa699_xor1[0], h_s_dadda_pg_rca32_fa700_xor1[0], h_s_dadda_pg_rca32_fa855_xor1, h_s_dadda_pg_rca32_fa855_or0);
  fa fa_h_s_dadda_pg_rca32_fa856_out(h_s_dadda_pg_rca32_fa855_or0[0], h_s_dadda_pg_rca32_fa701_xor1[0], h_s_dadda_pg_rca32_fa702_xor1[0], h_s_dadda_pg_rca32_fa856_xor1, h_s_dadda_pg_rca32_fa856_or0);
  fa fa_h_s_dadda_pg_rca32_fa857_out(h_s_dadda_pg_rca32_fa856_or0[0], h_s_dadda_pg_rca32_fa703_xor1[0], h_s_dadda_pg_rca32_fa704_xor1[0], h_s_dadda_pg_rca32_fa857_xor1, h_s_dadda_pg_rca32_fa857_or0);
  fa fa_h_s_dadda_pg_rca32_fa858_out(h_s_dadda_pg_rca32_fa857_or0[0], h_s_dadda_pg_rca32_fa705_xor1[0], h_s_dadda_pg_rca32_fa706_xor1[0], h_s_dadda_pg_rca32_fa858_xor1, h_s_dadda_pg_rca32_fa858_or0);
  fa fa_h_s_dadda_pg_rca32_fa859_out(h_s_dadda_pg_rca32_fa858_or0[0], h_s_dadda_pg_rca32_fa707_xor1[0], h_s_dadda_pg_rca32_fa708_xor1[0], h_s_dadda_pg_rca32_fa859_xor1, h_s_dadda_pg_rca32_fa859_or0);
  fa fa_h_s_dadda_pg_rca32_fa860_out(h_s_dadda_pg_rca32_fa859_or0[0], h_s_dadda_pg_rca32_fa709_xor1[0], h_s_dadda_pg_rca32_fa710_xor1[0], h_s_dadda_pg_rca32_fa860_xor1, h_s_dadda_pg_rca32_fa860_or0);
  fa fa_h_s_dadda_pg_rca32_fa861_out(h_s_dadda_pg_rca32_fa860_or0[0], h_s_dadda_pg_rca32_fa711_xor1[0], h_s_dadda_pg_rca32_fa712_xor1[0], h_s_dadda_pg_rca32_fa861_xor1, h_s_dadda_pg_rca32_fa861_or0);
  fa fa_h_s_dadda_pg_rca32_fa862_out(h_s_dadda_pg_rca32_fa861_or0[0], h_s_dadda_pg_rca32_fa713_xor1[0], h_s_dadda_pg_rca32_fa714_xor1[0], h_s_dadda_pg_rca32_fa862_xor1, h_s_dadda_pg_rca32_fa862_or0);
  fa fa_h_s_dadda_pg_rca32_fa863_out(h_s_dadda_pg_rca32_fa862_or0[0], h_s_dadda_pg_rca32_fa715_xor1[0], h_s_dadda_pg_rca32_fa716_xor1[0], h_s_dadda_pg_rca32_fa863_xor1, h_s_dadda_pg_rca32_fa863_or0);
  fa fa_h_s_dadda_pg_rca32_fa864_out(h_s_dadda_pg_rca32_fa863_or0[0], h_s_dadda_pg_rca32_fa717_xor1[0], h_s_dadda_pg_rca32_fa718_xor1[0], h_s_dadda_pg_rca32_fa864_xor1, h_s_dadda_pg_rca32_fa864_or0);
  fa fa_h_s_dadda_pg_rca32_fa865_out(h_s_dadda_pg_rca32_fa864_or0[0], h_s_dadda_pg_rca32_fa719_xor1[0], h_s_dadda_pg_rca32_fa720_xor1[0], h_s_dadda_pg_rca32_fa865_xor1, h_s_dadda_pg_rca32_fa865_or0);
  fa fa_h_s_dadda_pg_rca32_fa866_out(h_s_dadda_pg_rca32_fa865_or0[0], h_s_dadda_pg_rca32_fa721_xor1[0], h_s_dadda_pg_rca32_fa722_xor1[0], h_s_dadda_pg_rca32_fa866_xor1, h_s_dadda_pg_rca32_fa866_or0);
  fa fa_h_s_dadda_pg_rca32_fa867_out(h_s_dadda_pg_rca32_fa866_or0[0], h_s_dadda_pg_rca32_fa723_xor1[0], h_s_dadda_pg_rca32_fa724_xor1[0], h_s_dadda_pg_rca32_fa867_xor1, h_s_dadda_pg_rca32_fa867_or0);
  fa fa_h_s_dadda_pg_rca32_fa868_out(h_s_dadda_pg_rca32_fa867_or0[0], h_s_dadda_pg_rca32_fa725_xor1[0], h_s_dadda_pg_rca32_fa726_xor1[0], h_s_dadda_pg_rca32_fa868_xor1, h_s_dadda_pg_rca32_fa868_or0);
  fa fa_h_s_dadda_pg_rca32_fa869_out(h_s_dadda_pg_rca32_fa868_or0[0], h_s_dadda_pg_rca32_fa727_xor1[0], h_s_dadda_pg_rca32_fa728_xor1[0], h_s_dadda_pg_rca32_fa869_xor1, h_s_dadda_pg_rca32_fa869_or0);
  fa fa_h_s_dadda_pg_rca32_fa870_out(h_s_dadda_pg_rca32_fa869_or0[0], h_s_dadda_pg_rca32_fa729_xor1[0], h_s_dadda_pg_rca32_fa730_xor1[0], h_s_dadda_pg_rca32_fa870_xor1, h_s_dadda_pg_rca32_fa870_or0);
  fa fa_h_s_dadda_pg_rca32_fa871_out(h_s_dadda_pg_rca32_fa870_or0[0], h_s_dadda_pg_rca32_fa731_xor1[0], h_s_dadda_pg_rca32_fa732_xor1[0], h_s_dadda_pg_rca32_fa871_xor1, h_s_dadda_pg_rca32_fa871_or0);
  fa fa_h_s_dadda_pg_rca32_fa872_out(h_s_dadda_pg_rca32_fa871_or0[0], h_s_dadda_pg_rca32_fa733_xor1[0], h_s_dadda_pg_rca32_fa734_xor1[0], h_s_dadda_pg_rca32_fa872_xor1, h_s_dadda_pg_rca32_fa872_or0);
  fa fa_h_s_dadda_pg_rca32_fa873_out(h_s_dadda_pg_rca32_fa872_or0[0], h_s_dadda_pg_rca32_fa735_xor1[0], h_s_dadda_pg_rca32_fa736_xor1[0], h_s_dadda_pg_rca32_fa873_xor1, h_s_dadda_pg_rca32_fa873_or0);
  fa fa_h_s_dadda_pg_rca32_fa874_out(h_s_dadda_pg_rca32_fa873_or0[0], h_s_dadda_pg_rca32_fa737_xor1[0], h_s_dadda_pg_rca32_fa738_xor1[0], h_s_dadda_pg_rca32_fa874_xor1, h_s_dadda_pg_rca32_fa874_or0);
  fa fa_h_s_dadda_pg_rca32_fa875_out(h_s_dadda_pg_rca32_fa874_or0[0], h_s_dadda_pg_rca32_fa739_xor1[0], h_s_dadda_pg_rca32_fa740_xor1[0], h_s_dadda_pg_rca32_fa875_xor1, h_s_dadda_pg_rca32_fa875_or0);
  fa fa_h_s_dadda_pg_rca32_fa876_out(h_s_dadda_pg_rca32_fa875_or0[0], h_s_dadda_pg_rca32_fa741_xor1[0], h_s_dadda_pg_rca32_fa742_xor1[0], h_s_dadda_pg_rca32_fa876_xor1, h_s_dadda_pg_rca32_fa876_or0);
  fa fa_h_s_dadda_pg_rca32_fa877_out(h_s_dadda_pg_rca32_fa876_or0[0], h_s_dadda_pg_rca32_fa743_xor1[0], h_s_dadda_pg_rca32_fa744_xor1[0], h_s_dadda_pg_rca32_fa877_xor1, h_s_dadda_pg_rca32_fa877_or0);
  fa fa_h_s_dadda_pg_rca32_fa878_out(h_s_dadda_pg_rca32_fa877_or0[0], h_s_dadda_pg_rca32_fa745_xor1[0], h_s_dadda_pg_rca32_fa746_xor1[0], h_s_dadda_pg_rca32_fa878_xor1, h_s_dadda_pg_rca32_fa878_or0);
  fa fa_h_s_dadda_pg_rca32_fa879_out(h_s_dadda_pg_rca32_fa878_or0[0], h_s_dadda_pg_rca32_fa747_xor1[0], h_s_dadda_pg_rca32_fa748_xor1[0], h_s_dadda_pg_rca32_fa879_xor1, h_s_dadda_pg_rca32_fa879_or0);
  fa fa_h_s_dadda_pg_rca32_fa880_out(h_s_dadda_pg_rca32_fa879_or0[0], h_s_dadda_pg_rca32_fa749_xor1[0], h_s_dadda_pg_rca32_fa750_xor1[0], h_s_dadda_pg_rca32_fa880_xor1, h_s_dadda_pg_rca32_fa880_or0);
  fa fa_h_s_dadda_pg_rca32_fa881_out(h_s_dadda_pg_rca32_fa880_or0[0], h_s_dadda_pg_rca32_fa751_xor1[0], h_s_dadda_pg_rca32_fa752_xor1[0], h_s_dadda_pg_rca32_fa881_xor1, h_s_dadda_pg_rca32_fa881_or0);
  fa fa_h_s_dadda_pg_rca32_fa882_out(h_s_dadda_pg_rca32_fa881_or0[0], h_s_dadda_pg_rca32_fa753_xor1[0], h_s_dadda_pg_rca32_fa754_xor1[0], h_s_dadda_pg_rca32_fa882_xor1, h_s_dadda_pg_rca32_fa882_or0);
  fa fa_h_s_dadda_pg_rca32_fa883_out(h_s_dadda_pg_rca32_fa882_or0[0], h_s_dadda_pg_rca32_fa755_xor1[0], h_s_dadda_pg_rca32_fa756_xor1[0], h_s_dadda_pg_rca32_fa883_xor1, h_s_dadda_pg_rca32_fa883_or0);
  fa fa_h_s_dadda_pg_rca32_fa884_out(h_s_dadda_pg_rca32_fa883_or0[0], h_s_dadda_pg_rca32_fa757_xor1[0], h_s_dadda_pg_rca32_fa758_xor1[0], h_s_dadda_pg_rca32_fa884_xor1, h_s_dadda_pg_rca32_fa884_or0);
  fa fa_h_s_dadda_pg_rca32_fa885_out(h_s_dadda_pg_rca32_fa884_or0[0], h_s_dadda_pg_rca32_fa759_xor1[0], h_s_dadda_pg_rca32_fa760_xor1[0], h_s_dadda_pg_rca32_fa885_xor1, h_s_dadda_pg_rca32_fa885_or0);
  fa fa_h_s_dadda_pg_rca32_fa886_out(h_s_dadda_pg_rca32_fa885_or0[0], h_s_dadda_pg_rca32_fa761_xor1[0], h_s_dadda_pg_rca32_fa762_xor1[0], h_s_dadda_pg_rca32_fa886_xor1, h_s_dadda_pg_rca32_fa886_or0);
  fa fa_h_s_dadda_pg_rca32_fa887_out(h_s_dadda_pg_rca32_fa886_or0[0], h_s_dadda_pg_rca32_fa763_xor1[0], h_s_dadda_pg_rca32_fa764_xor1[0], h_s_dadda_pg_rca32_fa887_xor1, h_s_dadda_pg_rca32_fa887_or0);
  fa fa_h_s_dadda_pg_rca32_fa888_out(h_s_dadda_pg_rca32_fa887_or0[0], h_s_dadda_pg_rca32_fa765_xor1[0], h_s_dadda_pg_rca32_fa766_xor1[0], h_s_dadda_pg_rca32_fa888_xor1, h_s_dadda_pg_rca32_fa888_or0);
  fa fa_h_s_dadda_pg_rca32_fa889_out(h_s_dadda_pg_rca32_fa888_or0[0], h_s_dadda_pg_rca32_fa767_xor1[0], h_s_dadda_pg_rca32_fa768_xor1[0], h_s_dadda_pg_rca32_fa889_xor1, h_s_dadda_pg_rca32_fa889_or0);
  fa fa_h_s_dadda_pg_rca32_fa890_out(h_s_dadda_pg_rca32_fa889_or0[0], h_s_dadda_pg_rca32_fa769_xor1[0], h_s_dadda_pg_rca32_fa770_xor1[0], h_s_dadda_pg_rca32_fa890_xor1, h_s_dadda_pg_rca32_fa890_or0);
  fa fa_h_s_dadda_pg_rca32_fa891_out(h_s_dadda_pg_rca32_fa890_or0[0], h_s_dadda_pg_rca32_fa771_xor1[0], h_s_dadda_pg_rca32_fa772_xor1[0], h_s_dadda_pg_rca32_fa891_xor1, h_s_dadda_pg_rca32_fa891_or0);
  fa fa_h_s_dadda_pg_rca32_fa892_out(h_s_dadda_pg_rca32_fa891_or0[0], h_s_dadda_pg_rca32_fa773_xor1[0], h_s_dadda_pg_rca32_fa774_xor1[0], h_s_dadda_pg_rca32_fa892_xor1, h_s_dadda_pg_rca32_fa892_or0);
  fa fa_h_s_dadda_pg_rca32_fa893_out(h_s_dadda_pg_rca32_fa892_or0[0], h_s_dadda_pg_rca32_fa775_xor1[0], h_s_dadda_pg_rca32_fa776_xor1[0], h_s_dadda_pg_rca32_fa893_xor1, h_s_dadda_pg_rca32_fa893_or0);
  fa fa_h_s_dadda_pg_rca32_fa894_out(h_s_dadda_pg_rca32_fa893_or0[0], h_s_dadda_pg_rca32_fa777_xor1[0], h_s_dadda_pg_rca32_fa778_xor1[0], h_s_dadda_pg_rca32_fa894_xor1, h_s_dadda_pg_rca32_fa894_or0);
  fa fa_h_s_dadda_pg_rca32_fa895_out(h_s_dadda_pg_rca32_fa894_or0[0], h_s_dadda_pg_rca32_fa779_xor1[0], h_s_dadda_pg_rca32_fa780_xor1[0], h_s_dadda_pg_rca32_fa895_xor1, h_s_dadda_pg_rca32_fa895_or0);
  fa fa_h_s_dadda_pg_rca32_fa896_out(h_s_dadda_pg_rca32_fa895_or0[0], h_s_dadda_pg_rca32_fa781_xor1[0], h_s_dadda_pg_rca32_fa782_xor1[0], h_s_dadda_pg_rca32_fa896_xor1, h_s_dadda_pg_rca32_fa896_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_28_31(a[28], b[31], h_s_dadda_pg_rca32_nand_28_31);
  fa fa_h_s_dadda_pg_rca32_fa897_out(h_s_dadda_pg_rca32_fa896_or0[0], h_s_dadda_pg_rca32_nand_28_31[0], h_s_dadda_pg_rca32_fa783_xor1[0], h_s_dadda_pg_rca32_fa897_xor1, h_s_dadda_pg_rca32_fa897_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_30_30(a[30], b[30], h_s_dadda_pg_rca32_and_30_30);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_29_31(a[29], b[31], h_s_dadda_pg_rca32_nand_29_31);
  fa fa_h_s_dadda_pg_rca32_fa898_out(h_s_dadda_pg_rca32_fa897_or0[0], h_s_dadda_pg_rca32_and_30_30[0], h_s_dadda_pg_rca32_nand_29_31[0], h_s_dadda_pg_rca32_fa898_xor1, h_s_dadda_pg_rca32_fa898_or0);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_31_30(a[31], b[30], h_s_dadda_pg_rca32_nand_31_30);
  fa fa_h_s_dadda_pg_rca32_fa899_out(h_s_dadda_pg_rca32_fa898_or0[0], h_s_dadda_pg_rca32_fa840_or0[0], h_s_dadda_pg_rca32_nand_31_30[0], h_s_dadda_pg_rca32_fa899_xor1, h_s_dadda_pg_rca32_fa899_or0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_0(a[0], b[0], h_s_dadda_pg_rca32_and_0_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_1_0(a[1], b[0], h_s_dadda_pg_rca32_and_1_0);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_2(a[0], b[2], h_s_dadda_pg_rca32_and_0_2);
  nand_gate nand_gate_h_s_dadda_pg_rca32_nand_30_31(a[30], b[31], h_s_dadda_pg_rca32_nand_30_31);
  and_gate and_gate_h_s_dadda_pg_rca32_and_0_1(a[0], b[1], h_s_dadda_pg_rca32_and_0_1);
  and_gate and_gate_h_s_dadda_pg_rca32_and_31_31(a[31], b[31], h_s_dadda_pg_rca32_and_31_31);
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[0] = h_s_dadda_pg_rca32_and_1_0[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[1] = h_s_dadda_pg_rca32_and_0_2[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[2] = h_s_dadda_pg_rca32_ha28_xor0[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[3] = h_s_dadda_pg_rca32_fa784_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[4] = h_s_dadda_pg_rca32_fa785_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[5] = h_s_dadda_pg_rca32_fa786_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[6] = h_s_dadda_pg_rca32_fa787_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[7] = h_s_dadda_pg_rca32_fa788_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[8] = h_s_dadda_pg_rca32_fa789_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[9] = h_s_dadda_pg_rca32_fa790_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[10] = h_s_dadda_pg_rca32_fa791_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[11] = h_s_dadda_pg_rca32_fa792_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[12] = h_s_dadda_pg_rca32_fa793_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[13] = h_s_dadda_pg_rca32_fa794_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[14] = h_s_dadda_pg_rca32_fa795_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[15] = h_s_dadda_pg_rca32_fa796_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[16] = h_s_dadda_pg_rca32_fa797_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[17] = h_s_dadda_pg_rca32_fa798_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[18] = h_s_dadda_pg_rca32_fa799_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[19] = h_s_dadda_pg_rca32_fa800_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[20] = h_s_dadda_pg_rca32_fa801_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[21] = h_s_dadda_pg_rca32_fa802_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[22] = h_s_dadda_pg_rca32_fa803_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[23] = h_s_dadda_pg_rca32_fa804_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[24] = h_s_dadda_pg_rca32_fa805_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[25] = h_s_dadda_pg_rca32_fa806_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[26] = h_s_dadda_pg_rca32_fa807_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[27] = h_s_dadda_pg_rca32_fa808_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[28] = h_s_dadda_pg_rca32_fa809_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[29] = h_s_dadda_pg_rca32_fa810_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[30] = h_s_dadda_pg_rca32_fa811_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[31] = h_s_dadda_pg_rca32_fa812_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[32] = h_s_dadda_pg_rca32_fa813_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[33] = h_s_dadda_pg_rca32_fa814_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[34] = h_s_dadda_pg_rca32_fa815_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[35] = h_s_dadda_pg_rca32_fa816_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[36] = h_s_dadda_pg_rca32_fa817_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[37] = h_s_dadda_pg_rca32_fa818_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[38] = h_s_dadda_pg_rca32_fa819_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[39] = h_s_dadda_pg_rca32_fa820_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[40] = h_s_dadda_pg_rca32_fa821_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[41] = h_s_dadda_pg_rca32_fa822_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[42] = h_s_dadda_pg_rca32_fa823_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[43] = h_s_dadda_pg_rca32_fa824_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[44] = h_s_dadda_pg_rca32_fa825_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[45] = h_s_dadda_pg_rca32_fa826_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[46] = h_s_dadda_pg_rca32_fa827_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[47] = h_s_dadda_pg_rca32_fa828_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[48] = h_s_dadda_pg_rca32_fa829_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[49] = h_s_dadda_pg_rca32_fa830_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[50] = h_s_dadda_pg_rca32_fa831_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[51] = h_s_dadda_pg_rca32_fa832_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[52] = h_s_dadda_pg_rca32_fa833_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[53] = h_s_dadda_pg_rca32_fa834_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[54] = h_s_dadda_pg_rca32_fa835_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[55] = h_s_dadda_pg_rca32_fa836_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[56] = h_s_dadda_pg_rca32_fa837_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[57] = h_s_dadda_pg_rca32_fa838_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[58] = h_s_dadda_pg_rca32_fa839_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[59] = h_s_dadda_pg_rca32_fa840_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[60] = h_s_dadda_pg_rca32_nand_30_31[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_a[61] = h_s_dadda_pg_rca32_fa899_or0[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[0] = h_s_dadda_pg_rca32_and_0_1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[1] = h_s_dadda_pg_rca32_ha29_xor0[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[2] = h_s_dadda_pg_rca32_fa841_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[3] = h_s_dadda_pg_rca32_fa842_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[4] = h_s_dadda_pg_rca32_fa843_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[5] = h_s_dadda_pg_rca32_fa844_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[6] = h_s_dadda_pg_rca32_fa845_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[7] = h_s_dadda_pg_rca32_fa846_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[8] = h_s_dadda_pg_rca32_fa847_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[9] = h_s_dadda_pg_rca32_fa848_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[10] = h_s_dadda_pg_rca32_fa849_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[11] = h_s_dadda_pg_rca32_fa850_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[12] = h_s_dadda_pg_rca32_fa851_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[13] = h_s_dadda_pg_rca32_fa852_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[14] = h_s_dadda_pg_rca32_fa853_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[15] = h_s_dadda_pg_rca32_fa854_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[16] = h_s_dadda_pg_rca32_fa855_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[17] = h_s_dadda_pg_rca32_fa856_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[18] = h_s_dadda_pg_rca32_fa857_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[19] = h_s_dadda_pg_rca32_fa858_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[20] = h_s_dadda_pg_rca32_fa859_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[21] = h_s_dadda_pg_rca32_fa860_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[22] = h_s_dadda_pg_rca32_fa861_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[23] = h_s_dadda_pg_rca32_fa862_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[24] = h_s_dadda_pg_rca32_fa863_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[25] = h_s_dadda_pg_rca32_fa864_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[26] = h_s_dadda_pg_rca32_fa865_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[27] = h_s_dadda_pg_rca32_fa866_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[28] = h_s_dadda_pg_rca32_fa867_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[29] = h_s_dadda_pg_rca32_fa868_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[30] = h_s_dadda_pg_rca32_fa869_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[31] = h_s_dadda_pg_rca32_fa870_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[32] = h_s_dadda_pg_rca32_fa871_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[33] = h_s_dadda_pg_rca32_fa872_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[34] = h_s_dadda_pg_rca32_fa873_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[35] = h_s_dadda_pg_rca32_fa874_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[36] = h_s_dadda_pg_rca32_fa875_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[37] = h_s_dadda_pg_rca32_fa876_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[38] = h_s_dadda_pg_rca32_fa877_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[39] = h_s_dadda_pg_rca32_fa878_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[40] = h_s_dadda_pg_rca32_fa879_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[41] = h_s_dadda_pg_rca32_fa880_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[42] = h_s_dadda_pg_rca32_fa881_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[43] = h_s_dadda_pg_rca32_fa882_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[44] = h_s_dadda_pg_rca32_fa883_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[45] = h_s_dadda_pg_rca32_fa884_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[46] = h_s_dadda_pg_rca32_fa885_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[47] = h_s_dadda_pg_rca32_fa886_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[48] = h_s_dadda_pg_rca32_fa887_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[49] = h_s_dadda_pg_rca32_fa888_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[50] = h_s_dadda_pg_rca32_fa889_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[51] = h_s_dadda_pg_rca32_fa890_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[52] = h_s_dadda_pg_rca32_fa891_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[53] = h_s_dadda_pg_rca32_fa892_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[54] = h_s_dadda_pg_rca32_fa893_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[55] = h_s_dadda_pg_rca32_fa894_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[56] = h_s_dadda_pg_rca32_fa895_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[57] = h_s_dadda_pg_rca32_fa896_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[58] = h_s_dadda_pg_rca32_fa897_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[59] = h_s_dadda_pg_rca32_fa898_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[60] = h_s_dadda_pg_rca32_fa899_xor1[0];
  assign h_s_dadda_pg_rca32_u_pg_rca62_b[61] = h_s_dadda_pg_rca32_and_31_31[0];
  u_pg_rca62 u_pg_rca62_h_s_dadda_pg_rca32_u_pg_rca62_out(h_s_dadda_pg_rca32_u_pg_rca62_a, h_s_dadda_pg_rca32_u_pg_rca62_b, h_s_dadda_pg_rca32_u_pg_rca62_out);
  not_gate not_gate_h_s_dadda_pg_rca32_xor0(h_s_dadda_pg_rca32_u_pg_rca62_out[62], h_s_dadda_pg_rca32_xor0);

  assign h_s_dadda_pg_rca32_out[0] = h_s_dadda_pg_rca32_and_0_0[0];
  assign h_s_dadda_pg_rca32_out[1] = h_s_dadda_pg_rca32_u_pg_rca62_out[0];
  assign h_s_dadda_pg_rca32_out[2] = h_s_dadda_pg_rca32_u_pg_rca62_out[1];
  assign h_s_dadda_pg_rca32_out[3] = h_s_dadda_pg_rca32_u_pg_rca62_out[2];
  assign h_s_dadda_pg_rca32_out[4] = h_s_dadda_pg_rca32_u_pg_rca62_out[3];
  assign h_s_dadda_pg_rca32_out[5] = h_s_dadda_pg_rca32_u_pg_rca62_out[4];
  assign h_s_dadda_pg_rca32_out[6] = h_s_dadda_pg_rca32_u_pg_rca62_out[5];
  assign h_s_dadda_pg_rca32_out[7] = h_s_dadda_pg_rca32_u_pg_rca62_out[6];
  assign h_s_dadda_pg_rca32_out[8] = h_s_dadda_pg_rca32_u_pg_rca62_out[7];
  assign h_s_dadda_pg_rca32_out[9] = h_s_dadda_pg_rca32_u_pg_rca62_out[8];
  assign h_s_dadda_pg_rca32_out[10] = h_s_dadda_pg_rca32_u_pg_rca62_out[9];
  assign h_s_dadda_pg_rca32_out[11] = h_s_dadda_pg_rca32_u_pg_rca62_out[10];
  assign h_s_dadda_pg_rca32_out[12] = h_s_dadda_pg_rca32_u_pg_rca62_out[11];
  assign h_s_dadda_pg_rca32_out[13] = h_s_dadda_pg_rca32_u_pg_rca62_out[12];
  assign h_s_dadda_pg_rca32_out[14] = h_s_dadda_pg_rca32_u_pg_rca62_out[13];
  assign h_s_dadda_pg_rca32_out[15] = h_s_dadda_pg_rca32_u_pg_rca62_out[14];
  assign h_s_dadda_pg_rca32_out[16] = h_s_dadda_pg_rca32_u_pg_rca62_out[15];
  assign h_s_dadda_pg_rca32_out[17] = h_s_dadda_pg_rca32_u_pg_rca62_out[16];
  assign h_s_dadda_pg_rca32_out[18] = h_s_dadda_pg_rca32_u_pg_rca62_out[17];
  assign h_s_dadda_pg_rca32_out[19] = h_s_dadda_pg_rca32_u_pg_rca62_out[18];
  assign h_s_dadda_pg_rca32_out[20] = h_s_dadda_pg_rca32_u_pg_rca62_out[19];
  assign h_s_dadda_pg_rca32_out[21] = h_s_dadda_pg_rca32_u_pg_rca62_out[20];
  assign h_s_dadda_pg_rca32_out[22] = h_s_dadda_pg_rca32_u_pg_rca62_out[21];
  assign h_s_dadda_pg_rca32_out[23] = h_s_dadda_pg_rca32_u_pg_rca62_out[22];
  assign h_s_dadda_pg_rca32_out[24] = h_s_dadda_pg_rca32_u_pg_rca62_out[23];
  assign h_s_dadda_pg_rca32_out[25] = h_s_dadda_pg_rca32_u_pg_rca62_out[24];
  assign h_s_dadda_pg_rca32_out[26] = h_s_dadda_pg_rca32_u_pg_rca62_out[25];
  assign h_s_dadda_pg_rca32_out[27] = h_s_dadda_pg_rca32_u_pg_rca62_out[26];
  assign h_s_dadda_pg_rca32_out[28] = h_s_dadda_pg_rca32_u_pg_rca62_out[27];
  assign h_s_dadda_pg_rca32_out[29] = h_s_dadda_pg_rca32_u_pg_rca62_out[28];
  assign h_s_dadda_pg_rca32_out[30] = h_s_dadda_pg_rca32_u_pg_rca62_out[29];
  assign h_s_dadda_pg_rca32_out[31] = h_s_dadda_pg_rca32_u_pg_rca62_out[30];
  assign h_s_dadda_pg_rca32_out[32] = h_s_dadda_pg_rca32_u_pg_rca62_out[31];
  assign h_s_dadda_pg_rca32_out[33] = h_s_dadda_pg_rca32_u_pg_rca62_out[32];
  assign h_s_dadda_pg_rca32_out[34] = h_s_dadda_pg_rca32_u_pg_rca62_out[33];
  assign h_s_dadda_pg_rca32_out[35] = h_s_dadda_pg_rca32_u_pg_rca62_out[34];
  assign h_s_dadda_pg_rca32_out[36] = h_s_dadda_pg_rca32_u_pg_rca62_out[35];
  assign h_s_dadda_pg_rca32_out[37] = h_s_dadda_pg_rca32_u_pg_rca62_out[36];
  assign h_s_dadda_pg_rca32_out[38] = h_s_dadda_pg_rca32_u_pg_rca62_out[37];
  assign h_s_dadda_pg_rca32_out[39] = h_s_dadda_pg_rca32_u_pg_rca62_out[38];
  assign h_s_dadda_pg_rca32_out[40] = h_s_dadda_pg_rca32_u_pg_rca62_out[39];
  assign h_s_dadda_pg_rca32_out[41] = h_s_dadda_pg_rca32_u_pg_rca62_out[40];
  assign h_s_dadda_pg_rca32_out[42] = h_s_dadda_pg_rca32_u_pg_rca62_out[41];
  assign h_s_dadda_pg_rca32_out[43] = h_s_dadda_pg_rca32_u_pg_rca62_out[42];
  assign h_s_dadda_pg_rca32_out[44] = h_s_dadda_pg_rca32_u_pg_rca62_out[43];
  assign h_s_dadda_pg_rca32_out[45] = h_s_dadda_pg_rca32_u_pg_rca62_out[44];
  assign h_s_dadda_pg_rca32_out[46] = h_s_dadda_pg_rca32_u_pg_rca62_out[45];
  assign h_s_dadda_pg_rca32_out[47] = h_s_dadda_pg_rca32_u_pg_rca62_out[46];
  assign h_s_dadda_pg_rca32_out[48] = h_s_dadda_pg_rca32_u_pg_rca62_out[47];
  assign h_s_dadda_pg_rca32_out[49] = h_s_dadda_pg_rca32_u_pg_rca62_out[48];
  assign h_s_dadda_pg_rca32_out[50] = h_s_dadda_pg_rca32_u_pg_rca62_out[49];
  assign h_s_dadda_pg_rca32_out[51] = h_s_dadda_pg_rca32_u_pg_rca62_out[50];
  assign h_s_dadda_pg_rca32_out[52] = h_s_dadda_pg_rca32_u_pg_rca62_out[51];
  assign h_s_dadda_pg_rca32_out[53] = h_s_dadda_pg_rca32_u_pg_rca62_out[52];
  assign h_s_dadda_pg_rca32_out[54] = h_s_dadda_pg_rca32_u_pg_rca62_out[53];
  assign h_s_dadda_pg_rca32_out[55] = h_s_dadda_pg_rca32_u_pg_rca62_out[54];
  assign h_s_dadda_pg_rca32_out[56] = h_s_dadda_pg_rca32_u_pg_rca62_out[55];
  assign h_s_dadda_pg_rca32_out[57] = h_s_dadda_pg_rca32_u_pg_rca62_out[56];
  assign h_s_dadda_pg_rca32_out[58] = h_s_dadda_pg_rca32_u_pg_rca62_out[57];
  assign h_s_dadda_pg_rca32_out[59] = h_s_dadda_pg_rca32_u_pg_rca62_out[58];
  assign h_s_dadda_pg_rca32_out[60] = h_s_dadda_pg_rca32_u_pg_rca62_out[59];
  assign h_s_dadda_pg_rca32_out[61] = h_s_dadda_pg_rca32_u_pg_rca62_out[60];
  assign h_s_dadda_pg_rca32_out[62] = h_s_dadda_pg_rca32_u_pg_rca62_out[61];
  assign h_s_dadda_pg_rca32_out[63] = h_s_dadda_pg_rca32_xor0[0];
endmodule