module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;
  wire constant_wire_value_1_y0;
  wire constant_wire_value_1_y1;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_y0;
  wire fa_y1;
  wire fa_cin;
  wire fa_y3;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module u_rca62(input [61:0] a, input [61:0] b, output [62:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire a_30;
  wire a_31;
  wire a_32;
  wire a_33;
  wire a_34;
  wire a_35;
  wire a_36;
  wire a_37;
  wire a_38;
  wire a_39;
  wire a_40;
  wire a_41;
  wire a_42;
  wire a_43;
  wire a_44;
  wire a_45;
  wire a_46;
  wire a_47;
  wire a_48;
  wire a_49;
  wire a_50;
  wire a_51;
  wire a_52;
  wire a_53;
  wire a_54;
  wire a_55;
  wire a_56;
  wire a_57;
  wire a_58;
  wire a_59;
  wire a_60;
  wire a_61;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire b_30;
  wire b_31;
  wire b_32;
  wire b_33;
  wire b_34;
  wire b_35;
  wire b_36;
  wire b_37;
  wire b_38;
  wire b_39;
  wire b_40;
  wire b_41;
  wire b_42;
  wire b_43;
  wire b_44;
  wire b_45;
  wire b_46;
  wire b_47;
  wire b_48;
  wire b_49;
  wire b_50;
  wire b_51;
  wire b_52;
  wire b_53;
  wire b_54;
  wire b_55;
  wire b_56;
  wire b_57;
  wire b_58;
  wire b_59;
  wire b_60;
  wire b_61;
  wire u_rca62_ha_y0;
  wire u_rca62_ha_y1;
  wire u_rca62_fa1_y2;
  wire u_rca62_fa1_y4;
  wire u_rca62_fa2_y2;
  wire u_rca62_fa2_y4;
  wire u_rca62_fa3_y2;
  wire u_rca62_fa3_y4;
  wire u_rca62_fa4_y2;
  wire u_rca62_fa4_y4;
  wire u_rca62_fa5_y2;
  wire u_rca62_fa5_y4;
  wire u_rca62_fa6_y2;
  wire u_rca62_fa6_y4;
  wire u_rca62_fa7_y2;
  wire u_rca62_fa7_y4;
  wire u_rca62_fa8_y2;
  wire u_rca62_fa8_y4;
  wire u_rca62_fa9_y2;
  wire u_rca62_fa9_y4;
  wire u_rca62_fa10_y2;
  wire u_rca62_fa10_y4;
  wire u_rca62_fa11_y2;
  wire u_rca62_fa11_y4;
  wire u_rca62_fa12_y2;
  wire u_rca62_fa12_y4;
  wire u_rca62_fa13_y2;
  wire u_rca62_fa13_y4;
  wire u_rca62_fa14_y2;
  wire u_rca62_fa14_y4;
  wire u_rca62_fa15_y2;
  wire u_rca62_fa15_y4;
  wire u_rca62_fa16_y2;
  wire u_rca62_fa16_y4;
  wire u_rca62_fa17_y2;
  wire u_rca62_fa17_y4;
  wire u_rca62_fa18_y2;
  wire u_rca62_fa18_y4;
  wire u_rca62_fa19_y2;
  wire u_rca62_fa19_y4;
  wire u_rca62_fa20_y2;
  wire u_rca62_fa20_y4;
  wire u_rca62_fa21_y2;
  wire u_rca62_fa21_y4;
  wire u_rca62_fa22_y2;
  wire u_rca62_fa22_y4;
  wire u_rca62_fa23_y2;
  wire u_rca62_fa23_y4;
  wire u_rca62_fa24_y2;
  wire u_rca62_fa24_y4;
  wire u_rca62_fa25_y2;
  wire u_rca62_fa25_y4;
  wire u_rca62_fa26_y2;
  wire u_rca62_fa26_y4;
  wire u_rca62_fa27_y2;
  wire u_rca62_fa27_y4;
  wire u_rca62_fa28_y2;
  wire u_rca62_fa28_y4;
  wire u_rca62_fa29_y2;
  wire u_rca62_fa29_y4;
  wire u_rca62_fa30_y2;
  wire u_rca62_fa30_y4;
  wire u_rca62_fa31_y2;
  wire u_rca62_fa31_y4;
  wire u_rca62_fa32_y2;
  wire u_rca62_fa32_y4;
  wire u_rca62_fa33_y2;
  wire u_rca62_fa33_y4;
  wire u_rca62_fa34_y2;
  wire u_rca62_fa34_y4;
  wire u_rca62_fa35_y2;
  wire u_rca62_fa35_y4;
  wire u_rca62_fa36_y2;
  wire u_rca62_fa36_y4;
  wire u_rca62_fa37_y2;
  wire u_rca62_fa37_y4;
  wire u_rca62_fa38_y2;
  wire u_rca62_fa38_y4;
  wire u_rca62_fa39_y2;
  wire u_rca62_fa39_y4;
  wire u_rca62_fa40_y2;
  wire u_rca62_fa40_y4;
  wire u_rca62_fa41_y2;
  wire u_rca62_fa41_y4;
  wire u_rca62_fa42_y2;
  wire u_rca62_fa42_y4;
  wire u_rca62_fa43_y2;
  wire u_rca62_fa43_y4;
  wire u_rca62_fa44_y2;
  wire u_rca62_fa44_y4;
  wire u_rca62_fa45_y2;
  wire u_rca62_fa45_y4;
  wire u_rca62_fa46_y2;
  wire u_rca62_fa46_y4;
  wire u_rca62_fa47_y2;
  wire u_rca62_fa47_y4;
  wire u_rca62_fa48_y2;
  wire u_rca62_fa48_y4;
  wire u_rca62_fa49_y2;
  wire u_rca62_fa49_y4;
  wire u_rca62_fa50_y2;
  wire u_rca62_fa50_y4;
  wire u_rca62_fa51_y2;
  wire u_rca62_fa51_y4;
  wire u_rca62_fa52_y2;
  wire u_rca62_fa52_y4;
  wire u_rca62_fa53_y2;
  wire u_rca62_fa53_y4;
  wire u_rca62_fa54_y2;
  wire u_rca62_fa54_y4;
  wire u_rca62_fa55_y2;
  wire u_rca62_fa55_y4;
  wire u_rca62_fa56_y2;
  wire u_rca62_fa56_y4;
  wire u_rca62_fa57_y2;
  wire u_rca62_fa57_y4;
  wire u_rca62_fa58_y2;
  wire u_rca62_fa58_y4;
  wire u_rca62_fa59_y2;
  wire u_rca62_fa59_y4;
  wire u_rca62_fa60_y2;
  wire u_rca62_fa60_y4;
  wire u_rca62_fa61_y2;
  wire u_rca62_fa61_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign a_30 = a[30];
  assign a_31 = a[31];
  assign a_32 = a[32];
  assign a_33 = a[33];
  assign a_34 = a[34];
  assign a_35 = a[35];
  assign a_36 = a[36];
  assign a_37 = a[37];
  assign a_38 = a[38];
  assign a_39 = a[39];
  assign a_40 = a[40];
  assign a_41 = a[41];
  assign a_42 = a[42];
  assign a_43 = a[43];
  assign a_44 = a[44];
  assign a_45 = a[45];
  assign a_46 = a[46];
  assign a_47 = a[47];
  assign a_48 = a[48];
  assign a_49 = a[49];
  assign a_50 = a[50];
  assign a_51 = a[51];
  assign a_52 = a[52];
  assign a_53 = a[53];
  assign a_54 = a[54];
  assign a_55 = a[55];
  assign a_56 = a[56];
  assign a_57 = a[57];
  assign a_58 = a[58];
  assign a_59 = a[59];
  assign a_60 = a[60];
  assign a_61 = a[61];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  assign b_30 = b[30];
  assign b_31 = b[31];
  assign b_32 = b[32];
  assign b_33 = b[33];
  assign b_34 = b[34];
  assign b_35 = b[35];
  assign b_36 = b[36];
  assign b_37 = b[37];
  assign b_38 = b[38];
  assign b_39 = b[39];
  assign b_40 = b[40];
  assign b_41 = b[41];
  assign b_42 = b[42];
  assign b_43 = b[43];
  assign b_44 = b[44];
  assign b_45 = b[45];
  assign b_46 = b[46];
  assign b_47 = b[47];
  assign b_48 = b[48];
  assign b_49 = b[49];
  assign b_50 = b[50];
  assign b_51 = b[51];
  assign b_52 = b[52];
  assign b_53 = b[53];
  assign b_54 = b[54];
  assign b_55 = b[55];
  assign b_56 = b[56];
  assign b_57 = b[57];
  assign b_58 = b[58];
  assign b_59 = b[59];
  assign b_60 = b[60];
  assign b_61 = b[61];
  ha ha_u_rca62_ha_y0(a_0, b_0, u_rca62_ha_y0, u_rca62_ha_y1);
  fa fa_u_rca62_fa1_y2(a_1, b_1, u_rca62_ha_y1, u_rca62_fa1_y2, u_rca62_fa1_y4);
  fa fa_u_rca62_fa2_y2(a_2, b_2, u_rca62_fa1_y4, u_rca62_fa2_y2, u_rca62_fa2_y4);
  fa fa_u_rca62_fa3_y2(a_3, b_3, u_rca62_fa2_y4, u_rca62_fa3_y2, u_rca62_fa3_y4);
  fa fa_u_rca62_fa4_y2(a_4, b_4, u_rca62_fa3_y4, u_rca62_fa4_y2, u_rca62_fa4_y4);
  fa fa_u_rca62_fa5_y2(a_5, b_5, u_rca62_fa4_y4, u_rca62_fa5_y2, u_rca62_fa5_y4);
  fa fa_u_rca62_fa6_y2(a_6, b_6, u_rca62_fa5_y4, u_rca62_fa6_y2, u_rca62_fa6_y4);
  fa fa_u_rca62_fa7_y2(a_7, b_7, u_rca62_fa6_y4, u_rca62_fa7_y2, u_rca62_fa7_y4);
  fa fa_u_rca62_fa8_y2(a_8, b_8, u_rca62_fa7_y4, u_rca62_fa8_y2, u_rca62_fa8_y4);
  fa fa_u_rca62_fa9_y2(a_9, b_9, u_rca62_fa8_y4, u_rca62_fa9_y2, u_rca62_fa9_y4);
  fa fa_u_rca62_fa10_y2(a_10, b_10, u_rca62_fa9_y4, u_rca62_fa10_y2, u_rca62_fa10_y4);
  fa fa_u_rca62_fa11_y2(a_11, b_11, u_rca62_fa10_y4, u_rca62_fa11_y2, u_rca62_fa11_y4);
  fa fa_u_rca62_fa12_y2(a_12, b_12, u_rca62_fa11_y4, u_rca62_fa12_y2, u_rca62_fa12_y4);
  fa fa_u_rca62_fa13_y2(a_13, b_13, u_rca62_fa12_y4, u_rca62_fa13_y2, u_rca62_fa13_y4);
  fa fa_u_rca62_fa14_y2(a_14, b_14, u_rca62_fa13_y4, u_rca62_fa14_y2, u_rca62_fa14_y4);
  fa fa_u_rca62_fa15_y2(a_15, b_15, u_rca62_fa14_y4, u_rca62_fa15_y2, u_rca62_fa15_y4);
  fa fa_u_rca62_fa16_y2(a_16, b_16, u_rca62_fa15_y4, u_rca62_fa16_y2, u_rca62_fa16_y4);
  fa fa_u_rca62_fa17_y2(a_17, b_17, u_rca62_fa16_y4, u_rca62_fa17_y2, u_rca62_fa17_y4);
  fa fa_u_rca62_fa18_y2(a_18, b_18, u_rca62_fa17_y4, u_rca62_fa18_y2, u_rca62_fa18_y4);
  fa fa_u_rca62_fa19_y2(a_19, b_19, u_rca62_fa18_y4, u_rca62_fa19_y2, u_rca62_fa19_y4);
  fa fa_u_rca62_fa20_y2(a_20, b_20, u_rca62_fa19_y4, u_rca62_fa20_y2, u_rca62_fa20_y4);
  fa fa_u_rca62_fa21_y2(a_21, b_21, u_rca62_fa20_y4, u_rca62_fa21_y2, u_rca62_fa21_y4);
  fa fa_u_rca62_fa22_y2(a_22, b_22, u_rca62_fa21_y4, u_rca62_fa22_y2, u_rca62_fa22_y4);
  fa fa_u_rca62_fa23_y2(a_23, b_23, u_rca62_fa22_y4, u_rca62_fa23_y2, u_rca62_fa23_y4);
  fa fa_u_rca62_fa24_y2(a_24, b_24, u_rca62_fa23_y4, u_rca62_fa24_y2, u_rca62_fa24_y4);
  fa fa_u_rca62_fa25_y2(a_25, b_25, u_rca62_fa24_y4, u_rca62_fa25_y2, u_rca62_fa25_y4);
  fa fa_u_rca62_fa26_y2(a_26, b_26, u_rca62_fa25_y4, u_rca62_fa26_y2, u_rca62_fa26_y4);
  fa fa_u_rca62_fa27_y2(a_27, b_27, u_rca62_fa26_y4, u_rca62_fa27_y2, u_rca62_fa27_y4);
  fa fa_u_rca62_fa28_y2(a_28, b_28, u_rca62_fa27_y4, u_rca62_fa28_y2, u_rca62_fa28_y4);
  fa fa_u_rca62_fa29_y2(a_29, b_29, u_rca62_fa28_y4, u_rca62_fa29_y2, u_rca62_fa29_y4);
  fa fa_u_rca62_fa30_y2(a_30, b_30, u_rca62_fa29_y4, u_rca62_fa30_y2, u_rca62_fa30_y4);
  fa fa_u_rca62_fa31_y2(a_31, b_31, u_rca62_fa30_y4, u_rca62_fa31_y2, u_rca62_fa31_y4);
  fa fa_u_rca62_fa32_y2(a_32, b_32, u_rca62_fa31_y4, u_rca62_fa32_y2, u_rca62_fa32_y4);
  fa fa_u_rca62_fa33_y2(a_33, b_33, u_rca62_fa32_y4, u_rca62_fa33_y2, u_rca62_fa33_y4);
  fa fa_u_rca62_fa34_y2(a_34, b_34, u_rca62_fa33_y4, u_rca62_fa34_y2, u_rca62_fa34_y4);
  fa fa_u_rca62_fa35_y2(a_35, b_35, u_rca62_fa34_y4, u_rca62_fa35_y2, u_rca62_fa35_y4);
  fa fa_u_rca62_fa36_y2(a_36, b_36, u_rca62_fa35_y4, u_rca62_fa36_y2, u_rca62_fa36_y4);
  fa fa_u_rca62_fa37_y2(a_37, b_37, u_rca62_fa36_y4, u_rca62_fa37_y2, u_rca62_fa37_y4);
  fa fa_u_rca62_fa38_y2(a_38, b_38, u_rca62_fa37_y4, u_rca62_fa38_y2, u_rca62_fa38_y4);
  fa fa_u_rca62_fa39_y2(a_39, b_39, u_rca62_fa38_y4, u_rca62_fa39_y2, u_rca62_fa39_y4);
  fa fa_u_rca62_fa40_y2(a_40, b_40, u_rca62_fa39_y4, u_rca62_fa40_y2, u_rca62_fa40_y4);
  fa fa_u_rca62_fa41_y2(a_41, b_41, u_rca62_fa40_y4, u_rca62_fa41_y2, u_rca62_fa41_y4);
  fa fa_u_rca62_fa42_y2(a_42, b_42, u_rca62_fa41_y4, u_rca62_fa42_y2, u_rca62_fa42_y4);
  fa fa_u_rca62_fa43_y2(a_43, b_43, u_rca62_fa42_y4, u_rca62_fa43_y2, u_rca62_fa43_y4);
  fa fa_u_rca62_fa44_y2(a_44, b_44, u_rca62_fa43_y4, u_rca62_fa44_y2, u_rca62_fa44_y4);
  fa fa_u_rca62_fa45_y2(a_45, b_45, u_rca62_fa44_y4, u_rca62_fa45_y2, u_rca62_fa45_y4);
  fa fa_u_rca62_fa46_y2(a_46, b_46, u_rca62_fa45_y4, u_rca62_fa46_y2, u_rca62_fa46_y4);
  fa fa_u_rca62_fa47_y2(a_47, b_47, u_rca62_fa46_y4, u_rca62_fa47_y2, u_rca62_fa47_y4);
  fa fa_u_rca62_fa48_y2(a_48, b_48, u_rca62_fa47_y4, u_rca62_fa48_y2, u_rca62_fa48_y4);
  fa fa_u_rca62_fa49_y2(a_49, b_49, u_rca62_fa48_y4, u_rca62_fa49_y2, u_rca62_fa49_y4);
  fa fa_u_rca62_fa50_y2(a_50, b_50, u_rca62_fa49_y4, u_rca62_fa50_y2, u_rca62_fa50_y4);
  fa fa_u_rca62_fa51_y2(a_51, b_51, u_rca62_fa50_y4, u_rca62_fa51_y2, u_rca62_fa51_y4);
  fa fa_u_rca62_fa52_y2(a_52, b_52, u_rca62_fa51_y4, u_rca62_fa52_y2, u_rca62_fa52_y4);
  fa fa_u_rca62_fa53_y2(a_53, b_53, u_rca62_fa52_y4, u_rca62_fa53_y2, u_rca62_fa53_y4);
  fa fa_u_rca62_fa54_y2(a_54, b_54, u_rca62_fa53_y4, u_rca62_fa54_y2, u_rca62_fa54_y4);
  fa fa_u_rca62_fa55_y2(a_55, b_55, u_rca62_fa54_y4, u_rca62_fa55_y2, u_rca62_fa55_y4);
  fa fa_u_rca62_fa56_y2(a_56, b_56, u_rca62_fa55_y4, u_rca62_fa56_y2, u_rca62_fa56_y4);
  fa fa_u_rca62_fa57_y2(a_57, b_57, u_rca62_fa56_y4, u_rca62_fa57_y2, u_rca62_fa57_y4);
  fa fa_u_rca62_fa58_y2(a_58, b_58, u_rca62_fa57_y4, u_rca62_fa58_y2, u_rca62_fa58_y4);
  fa fa_u_rca62_fa59_y2(a_59, b_59, u_rca62_fa58_y4, u_rca62_fa59_y2, u_rca62_fa59_y4);
  fa fa_u_rca62_fa60_y2(a_60, b_60, u_rca62_fa59_y4, u_rca62_fa60_y2, u_rca62_fa60_y4);
  fa fa_u_rca62_fa61_y2(a_61, b_61, u_rca62_fa60_y4, u_rca62_fa61_y2, u_rca62_fa61_y4);

  assign out[0] = u_rca62_ha_y0;
  assign out[1] = u_rca62_fa1_y2;
  assign out[2] = u_rca62_fa2_y2;
  assign out[3] = u_rca62_fa3_y2;
  assign out[4] = u_rca62_fa4_y2;
  assign out[5] = u_rca62_fa5_y2;
  assign out[6] = u_rca62_fa6_y2;
  assign out[7] = u_rca62_fa7_y2;
  assign out[8] = u_rca62_fa8_y2;
  assign out[9] = u_rca62_fa9_y2;
  assign out[10] = u_rca62_fa10_y2;
  assign out[11] = u_rca62_fa11_y2;
  assign out[12] = u_rca62_fa12_y2;
  assign out[13] = u_rca62_fa13_y2;
  assign out[14] = u_rca62_fa14_y2;
  assign out[15] = u_rca62_fa15_y2;
  assign out[16] = u_rca62_fa16_y2;
  assign out[17] = u_rca62_fa17_y2;
  assign out[18] = u_rca62_fa18_y2;
  assign out[19] = u_rca62_fa19_y2;
  assign out[20] = u_rca62_fa20_y2;
  assign out[21] = u_rca62_fa21_y2;
  assign out[22] = u_rca62_fa22_y2;
  assign out[23] = u_rca62_fa23_y2;
  assign out[24] = u_rca62_fa24_y2;
  assign out[25] = u_rca62_fa25_y2;
  assign out[26] = u_rca62_fa26_y2;
  assign out[27] = u_rca62_fa27_y2;
  assign out[28] = u_rca62_fa28_y2;
  assign out[29] = u_rca62_fa29_y2;
  assign out[30] = u_rca62_fa30_y2;
  assign out[31] = u_rca62_fa31_y2;
  assign out[32] = u_rca62_fa32_y2;
  assign out[33] = u_rca62_fa33_y2;
  assign out[34] = u_rca62_fa34_y2;
  assign out[35] = u_rca62_fa35_y2;
  assign out[36] = u_rca62_fa36_y2;
  assign out[37] = u_rca62_fa37_y2;
  assign out[38] = u_rca62_fa38_y2;
  assign out[39] = u_rca62_fa39_y2;
  assign out[40] = u_rca62_fa40_y2;
  assign out[41] = u_rca62_fa41_y2;
  assign out[42] = u_rca62_fa42_y2;
  assign out[43] = u_rca62_fa43_y2;
  assign out[44] = u_rca62_fa44_y2;
  assign out[45] = u_rca62_fa45_y2;
  assign out[46] = u_rca62_fa46_y2;
  assign out[47] = u_rca62_fa47_y2;
  assign out[48] = u_rca62_fa48_y2;
  assign out[49] = u_rca62_fa49_y2;
  assign out[50] = u_rca62_fa50_y2;
  assign out[51] = u_rca62_fa51_y2;
  assign out[52] = u_rca62_fa52_y2;
  assign out[53] = u_rca62_fa53_y2;
  assign out[54] = u_rca62_fa54_y2;
  assign out[55] = u_rca62_fa55_y2;
  assign out[56] = u_rca62_fa56_y2;
  assign out[57] = u_rca62_fa57_y2;
  assign out[58] = u_rca62_fa58_y2;
  assign out[59] = u_rca62_fa59_y2;
  assign out[60] = u_rca62_fa60_y2;
  assign out[61] = u_rca62_fa61_y2;
  assign out[62] = u_rca62_fa61_y4;
endmodule

module h_s_dadda_rca32(input [31:0] a, input [31:0] b, output [63:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire a_30;
  wire a_31;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire b_30;
  wire b_31;
  wire constant_wire_1;
  wire h_s_dadda_rca32_and_28_0_y0;
  wire h_s_dadda_rca32_and_27_1_y0;
  wire h_s_dadda_rca32_ha0_y0;
  wire h_s_dadda_rca32_ha0_y1;
  wire h_s_dadda_rca32_and_29_0_y0;
  wire h_s_dadda_rca32_and_28_1_y0;
  wire h_s_dadda_rca32_fa0_y2;
  wire h_s_dadda_rca32_fa0_y4;
  wire h_s_dadda_rca32_and_27_2_y0;
  wire h_s_dadda_rca32_and_26_3_y0;
  wire h_s_dadda_rca32_ha1_y0;
  wire h_s_dadda_rca32_ha1_y1;
  wire h_s_dadda_rca32_and_30_0_y0;
  wire h_s_dadda_rca32_fa1_y2;
  wire h_s_dadda_rca32_fa1_y4;
  wire h_s_dadda_rca32_and_29_1_y0;
  wire h_s_dadda_rca32_and_28_2_y0;
  wire h_s_dadda_rca32_and_27_3_y0;
  wire h_s_dadda_rca32_fa2_y2;
  wire h_s_dadda_rca32_fa2_y4;
  wire h_s_dadda_rca32_and_26_4_y0;
  wire h_s_dadda_rca32_and_25_5_y0;
  wire h_s_dadda_rca32_ha2_y0;
  wire h_s_dadda_rca32_ha2_y1;
  wire h_s_dadda_rca32_fa3_y2;
  wire h_s_dadda_rca32_fa3_y4;
  wire h_s_dadda_rca32_nand_31_0_y0;
  wire h_s_dadda_rca32_and_30_1_y0;
  wire h_s_dadda_rca32_and_29_2_y0;
  wire h_s_dadda_rca32_fa4_y2;
  wire h_s_dadda_rca32_fa4_y4;
  wire h_s_dadda_rca32_and_28_3_y0;
  wire h_s_dadda_rca32_and_27_4_y0;
  wire h_s_dadda_rca32_and_26_5_y0;
  wire h_s_dadda_rca32_fa5_y2;
  wire h_s_dadda_rca32_fa5_y4;
  wire h_s_dadda_rca32_and_25_6_y0;
  wire h_s_dadda_rca32_and_24_7_y0;
  wire h_s_dadda_rca32_ha3_y0;
  wire h_s_dadda_rca32_ha3_y1;
  wire h_s_dadda_rca32_fa6_y2;
  wire h_s_dadda_rca32_fa6_y4;
  wire h_s_dadda_rca32_nand_31_1_y0;
  wire h_s_dadda_rca32_fa7_y2;
  wire h_s_dadda_rca32_fa7_y4;
  wire h_s_dadda_rca32_and_30_2_y0;
  wire h_s_dadda_rca32_and_29_3_y0;
  wire h_s_dadda_rca32_and_28_4_y0;
  wire h_s_dadda_rca32_fa8_y2;
  wire h_s_dadda_rca32_fa8_y4;
  wire h_s_dadda_rca32_and_27_5_y0;
  wire h_s_dadda_rca32_and_26_6_y0;
  wire h_s_dadda_rca32_and_25_7_y0;
  wire h_s_dadda_rca32_fa9_y2;
  wire h_s_dadda_rca32_fa9_y4;
  wire h_s_dadda_rca32_fa10_y2;
  wire h_s_dadda_rca32_fa10_y4;
  wire h_s_dadda_rca32_nand_31_2_y0;
  wire h_s_dadda_rca32_and_30_3_y0;
  wire h_s_dadda_rca32_fa11_y2;
  wire h_s_dadda_rca32_fa11_y4;
  wire h_s_dadda_rca32_and_29_4_y0;
  wire h_s_dadda_rca32_and_28_5_y0;
  wire h_s_dadda_rca32_and_27_6_y0;
  wire h_s_dadda_rca32_fa12_y2;
  wire h_s_dadda_rca32_fa12_y4;
  wire h_s_dadda_rca32_fa13_y2;
  wire h_s_dadda_rca32_fa13_y4;
  wire h_s_dadda_rca32_nand_31_3_y0;
  wire h_s_dadda_rca32_and_30_4_y0;
  wire h_s_dadda_rca32_and_29_5_y0;
  wire h_s_dadda_rca32_fa14_y2;
  wire h_s_dadda_rca32_fa14_y4;
  wire h_s_dadda_rca32_nand_31_4_y0;
  wire h_s_dadda_rca32_fa15_y2;
  wire h_s_dadda_rca32_fa15_y4;
  wire h_s_dadda_rca32_and_6_0_y0;
  wire h_s_dadda_rca32_and_5_1_y0;
  wire h_s_dadda_rca32_ha4_y0;
  wire h_s_dadda_rca32_ha4_y1;
  wire h_s_dadda_rca32_and_7_0_y0;
  wire h_s_dadda_rca32_and_6_1_y0;
  wire h_s_dadda_rca32_fa16_y2;
  wire h_s_dadda_rca32_fa16_y4;
  wire h_s_dadda_rca32_and_5_2_y0;
  wire h_s_dadda_rca32_and_4_3_y0;
  wire h_s_dadda_rca32_ha5_y0;
  wire h_s_dadda_rca32_ha5_y1;
  wire h_s_dadda_rca32_and_8_0_y0;
  wire h_s_dadda_rca32_fa17_y2;
  wire h_s_dadda_rca32_fa17_y4;
  wire h_s_dadda_rca32_and_7_1_y0;
  wire h_s_dadda_rca32_and_6_2_y0;
  wire h_s_dadda_rca32_and_5_3_y0;
  wire h_s_dadda_rca32_fa18_y2;
  wire h_s_dadda_rca32_fa18_y4;
  wire h_s_dadda_rca32_and_4_4_y0;
  wire h_s_dadda_rca32_and_3_5_y0;
  wire h_s_dadda_rca32_ha6_y0;
  wire h_s_dadda_rca32_ha6_y1;
  wire h_s_dadda_rca32_fa19_y2;
  wire h_s_dadda_rca32_fa19_y4;
  wire h_s_dadda_rca32_and_9_0_y0;
  wire h_s_dadda_rca32_and_8_1_y0;
  wire h_s_dadda_rca32_and_7_2_y0;
  wire h_s_dadda_rca32_fa20_y2;
  wire h_s_dadda_rca32_fa20_y4;
  wire h_s_dadda_rca32_and_6_3_y0;
  wire h_s_dadda_rca32_and_5_4_y0;
  wire h_s_dadda_rca32_and_4_5_y0;
  wire h_s_dadda_rca32_fa21_y2;
  wire h_s_dadda_rca32_fa21_y4;
  wire h_s_dadda_rca32_and_3_6_y0;
  wire h_s_dadda_rca32_and_2_7_y0;
  wire h_s_dadda_rca32_ha7_y0;
  wire h_s_dadda_rca32_ha7_y1;
  wire h_s_dadda_rca32_fa22_y2;
  wire h_s_dadda_rca32_fa22_y4;
  wire h_s_dadda_rca32_and_10_0_y0;
  wire h_s_dadda_rca32_and_9_1_y0;
  wire h_s_dadda_rca32_fa23_y2;
  wire h_s_dadda_rca32_fa23_y4;
  wire h_s_dadda_rca32_and_8_2_y0;
  wire h_s_dadda_rca32_and_7_3_y0;
  wire h_s_dadda_rca32_and_6_4_y0;
  wire h_s_dadda_rca32_fa24_y2;
  wire h_s_dadda_rca32_fa24_y4;
  wire h_s_dadda_rca32_and_5_5_y0;
  wire h_s_dadda_rca32_and_4_6_y0;
  wire h_s_dadda_rca32_and_3_7_y0;
  wire h_s_dadda_rca32_fa25_y2;
  wire h_s_dadda_rca32_fa25_y4;
  wire h_s_dadda_rca32_and_2_8_y0;
  wire h_s_dadda_rca32_and_1_9_y0;
  wire h_s_dadda_rca32_ha8_y0;
  wire h_s_dadda_rca32_ha8_y1;
  wire h_s_dadda_rca32_fa26_y2;
  wire h_s_dadda_rca32_fa26_y4;
  wire h_s_dadda_rca32_and_11_0_y0;
  wire h_s_dadda_rca32_fa27_y2;
  wire h_s_dadda_rca32_fa27_y4;
  wire h_s_dadda_rca32_and_10_1_y0;
  wire h_s_dadda_rca32_and_9_2_y0;
  wire h_s_dadda_rca32_and_8_3_y0;
  wire h_s_dadda_rca32_fa28_y2;
  wire h_s_dadda_rca32_fa28_y4;
  wire h_s_dadda_rca32_and_7_4_y0;
  wire h_s_dadda_rca32_and_6_5_y0;
  wire h_s_dadda_rca32_and_5_6_y0;
  wire h_s_dadda_rca32_fa29_y2;
  wire h_s_dadda_rca32_fa29_y4;
  wire h_s_dadda_rca32_and_4_7_y0;
  wire h_s_dadda_rca32_and_3_8_y0;
  wire h_s_dadda_rca32_and_2_9_y0;
  wire h_s_dadda_rca32_fa30_y2;
  wire h_s_dadda_rca32_fa30_y4;
  wire h_s_dadda_rca32_and_1_10_y0;
  wire h_s_dadda_rca32_and_0_11_y0;
  wire h_s_dadda_rca32_ha9_y0;
  wire h_s_dadda_rca32_ha9_y1;
  wire h_s_dadda_rca32_fa31_y2;
  wire h_s_dadda_rca32_fa31_y4;
  wire h_s_dadda_rca32_fa32_y2;
  wire h_s_dadda_rca32_fa32_y4;
  wire h_s_dadda_rca32_and_12_0_y0;
  wire h_s_dadda_rca32_and_11_1_y0;
  wire h_s_dadda_rca32_and_10_2_y0;
  wire h_s_dadda_rca32_fa33_y2;
  wire h_s_dadda_rca32_fa33_y4;
  wire h_s_dadda_rca32_and_9_3_y0;
  wire h_s_dadda_rca32_and_8_4_y0;
  wire h_s_dadda_rca32_and_7_5_y0;
  wire h_s_dadda_rca32_fa34_y2;
  wire h_s_dadda_rca32_fa34_y4;
  wire h_s_dadda_rca32_and_6_6_y0;
  wire h_s_dadda_rca32_and_5_7_y0;
  wire h_s_dadda_rca32_and_4_8_y0;
  wire h_s_dadda_rca32_fa35_y2;
  wire h_s_dadda_rca32_fa35_y4;
  wire h_s_dadda_rca32_and_3_9_y0;
  wire h_s_dadda_rca32_and_2_10_y0;
  wire h_s_dadda_rca32_and_1_11_y0;
  wire h_s_dadda_rca32_fa36_y2;
  wire h_s_dadda_rca32_fa36_y4;
  wire h_s_dadda_rca32_and_0_12_y0;
  wire h_s_dadda_rca32_ha10_y0;
  wire h_s_dadda_rca32_ha10_y1;
  wire h_s_dadda_rca32_fa37_y2;
  wire h_s_dadda_rca32_fa37_y4;
  wire h_s_dadda_rca32_fa38_y2;
  wire h_s_dadda_rca32_fa38_y4;
  wire h_s_dadda_rca32_and_13_0_y0;
  wire h_s_dadda_rca32_and_12_1_y0;
  wire h_s_dadda_rca32_fa39_y2;
  wire h_s_dadda_rca32_fa39_y4;
  wire h_s_dadda_rca32_and_11_2_y0;
  wire h_s_dadda_rca32_and_10_3_y0;
  wire h_s_dadda_rca32_and_9_4_y0;
  wire h_s_dadda_rca32_fa40_y2;
  wire h_s_dadda_rca32_fa40_y4;
  wire h_s_dadda_rca32_and_8_5_y0;
  wire h_s_dadda_rca32_and_7_6_y0;
  wire h_s_dadda_rca32_and_6_7_y0;
  wire h_s_dadda_rca32_fa41_y2;
  wire h_s_dadda_rca32_fa41_y4;
  wire h_s_dadda_rca32_and_5_8_y0;
  wire h_s_dadda_rca32_and_4_9_y0;
  wire h_s_dadda_rca32_and_3_10_y0;
  wire h_s_dadda_rca32_fa42_y2;
  wire h_s_dadda_rca32_fa42_y4;
  wire h_s_dadda_rca32_and_2_11_y0;
  wire h_s_dadda_rca32_and_1_12_y0;
  wire h_s_dadda_rca32_and_0_13_y0;
  wire h_s_dadda_rca32_fa43_y2;
  wire h_s_dadda_rca32_fa43_y4;
  wire h_s_dadda_rca32_ha11_y0;
  wire h_s_dadda_rca32_ha11_y1;
  wire h_s_dadda_rca32_fa44_y2;
  wire h_s_dadda_rca32_fa44_y4;
  wire h_s_dadda_rca32_fa45_y2;
  wire h_s_dadda_rca32_fa45_y4;
  wire h_s_dadda_rca32_and_14_0_y0;
  wire h_s_dadda_rca32_fa46_y2;
  wire h_s_dadda_rca32_fa46_y4;
  wire h_s_dadda_rca32_and_13_1_y0;
  wire h_s_dadda_rca32_and_12_2_y0;
  wire h_s_dadda_rca32_and_11_3_y0;
  wire h_s_dadda_rca32_fa47_y2;
  wire h_s_dadda_rca32_fa47_y4;
  wire h_s_dadda_rca32_and_10_4_y0;
  wire h_s_dadda_rca32_and_9_5_y0;
  wire h_s_dadda_rca32_and_8_6_y0;
  wire h_s_dadda_rca32_fa48_y2;
  wire h_s_dadda_rca32_fa48_y4;
  wire h_s_dadda_rca32_and_7_7_y0;
  wire h_s_dadda_rca32_and_6_8_y0;
  wire h_s_dadda_rca32_and_5_9_y0;
  wire h_s_dadda_rca32_fa49_y2;
  wire h_s_dadda_rca32_fa49_y4;
  wire h_s_dadda_rca32_and_4_10_y0;
  wire h_s_dadda_rca32_and_3_11_y0;
  wire h_s_dadda_rca32_and_2_12_y0;
  wire h_s_dadda_rca32_fa50_y2;
  wire h_s_dadda_rca32_fa50_y4;
  wire h_s_dadda_rca32_and_1_13_y0;
  wire h_s_dadda_rca32_and_0_14_y0;
  wire h_s_dadda_rca32_fa51_y2;
  wire h_s_dadda_rca32_fa51_y4;
  wire h_s_dadda_rca32_ha12_y0;
  wire h_s_dadda_rca32_ha12_y1;
  wire h_s_dadda_rca32_fa52_y2;
  wire h_s_dadda_rca32_fa52_y4;
  wire h_s_dadda_rca32_fa53_y2;
  wire h_s_dadda_rca32_fa53_y4;
  wire h_s_dadda_rca32_fa54_y2;
  wire h_s_dadda_rca32_fa54_y4;
  wire h_s_dadda_rca32_and_15_0_y0;
  wire h_s_dadda_rca32_and_14_1_y0;
  wire h_s_dadda_rca32_and_13_2_y0;
  wire h_s_dadda_rca32_fa55_y2;
  wire h_s_dadda_rca32_fa55_y4;
  wire h_s_dadda_rca32_and_12_3_y0;
  wire h_s_dadda_rca32_and_11_4_y0;
  wire h_s_dadda_rca32_and_10_5_y0;
  wire h_s_dadda_rca32_fa56_y2;
  wire h_s_dadda_rca32_fa56_y4;
  wire h_s_dadda_rca32_and_9_6_y0;
  wire h_s_dadda_rca32_and_8_7_y0;
  wire h_s_dadda_rca32_and_7_8_y0;
  wire h_s_dadda_rca32_fa57_y2;
  wire h_s_dadda_rca32_fa57_y4;
  wire h_s_dadda_rca32_and_6_9_y0;
  wire h_s_dadda_rca32_and_5_10_y0;
  wire h_s_dadda_rca32_and_4_11_y0;
  wire h_s_dadda_rca32_fa58_y2;
  wire h_s_dadda_rca32_fa58_y4;
  wire h_s_dadda_rca32_and_3_12_y0;
  wire h_s_dadda_rca32_and_2_13_y0;
  wire h_s_dadda_rca32_and_1_14_y0;
  wire h_s_dadda_rca32_fa59_y2;
  wire h_s_dadda_rca32_fa59_y4;
  wire h_s_dadda_rca32_and_0_15_y0;
  wire h_s_dadda_rca32_fa60_y2;
  wire h_s_dadda_rca32_fa60_y4;
  wire h_s_dadda_rca32_ha13_y0;
  wire h_s_dadda_rca32_ha13_y1;
  wire h_s_dadda_rca32_fa61_y2;
  wire h_s_dadda_rca32_fa61_y4;
  wire h_s_dadda_rca32_fa62_y2;
  wire h_s_dadda_rca32_fa62_y4;
  wire h_s_dadda_rca32_fa63_y2;
  wire h_s_dadda_rca32_fa63_y4;
  wire h_s_dadda_rca32_and_16_0_y0;
  wire h_s_dadda_rca32_and_15_1_y0;
  wire h_s_dadda_rca32_fa64_y2;
  wire h_s_dadda_rca32_fa64_y4;
  wire h_s_dadda_rca32_and_14_2_y0;
  wire h_s_dadda_rca32_and_13_3_y0;
  wire h_s_dadda_rca32_and_12_4_y0;
  wire h_s_dadda_rca32_fa65_y2;
  wire h_s_dadda_rca32_fa65_y4;
  wire h_s_dadda_rca32_and_11_5_y0;
  wire h_s_dadda_rca32_and_10_6_y0;
  wire h_s_dadda_rca32_and_9_7_y0;
  wire h_s_dadda_rca32_fa66_y2;
  wire h_s_dadda_rca32_fa66_y4;
  wire h_s_dadda_rca32_and_8_8_y0;
  wire h_s_dadda_rca32_and_7_9_y0;
  wire h_s_dadda_rca32_and_6_10_y0;
  wire h_s_dadda_rca32_fa67_y2;
  wire h_s_dadda_rca32_fa67_y4;
  wire h_s_dadda_rca32_and_5_11_y0;
  wire h_s_dadda_rca32_and_4_12_y0;
  wire h_s_dadda_rca32_and_3_13_y0;
  wire h_s_dadda_rca32_fa68_y2;
  wire h_s_dadda_rca32_fa68_y4;
  wire h_s_dadda_rca32_and_2_14_y0;
  wire h_s_dadda_rca32_and_1_15_y0;
  wire h_s_dadda_rca32_and_0_16_y0;
  wire h_s_dadda_rca32_fa69_y2;
  wire h_s_dadda_rca32_fa69_y4;
  wire h_s_dadda_rca32_fa70_y2;
  wire h_s_dadda_rca32_fa70_y4;
  wire h_s_dadda_rca32_ha14_y0;
  wire h_s_dadda_rca32_ha14_y1;
  wire h_s_dadda_rca32_fa71_y2;
  wire h_s_dadda_rca32_fa71_y4;
  wire h_s_dadda_rca32_fa72_y2;
  wire h_s_dadda_rca32_fa72_y4;
  wire h_s_dadda_rca32_fa73_y2;
  wire h_s_dadda_rca32_fa73_y4;
  wire h_s_dadda_rca32_and_17_0_y0;
  wire h_s_dadda_rca32_fa74_y2;
  wire h_s_dadda_rca32_fa74_y4;
  wire h_s_dadda_rca32_and_16_1_y0;
  wire h_s_dadda_rca32_and_15_2_y0;
  wire h_s_dadda_rca32_and_14_3_y0;
  wire h_s_dadda_rca32_fa75_y2;
  wire h_s_dadda_rca32_fa75_y4;
  wire h_s_dadda_rca32_and_13_4_y0;
  wire h_s_dadda_rca32_and_12_5_y0;
  wire h_s_dadda_rca32_and_11_6_y0;
  wire h_s_dadda_rca32_fa76_y2;
  wire h_s_dadda_rca32_fa76_y4;
  wire h_s_dadda_rca32_and_10_7_y0;
  wire h_s_dadda_rca32_and_9_8_y0;
  wire h_s_dadda_rca32_and_8_9_y0;
  wire h_s_dadda_rca32_fa77_y2;
  wire h_s_dadda_rca32_fa77_y4;
  wire h_s_dadda_rca32_and_7_10_y0;
  wire h_s_dadda_rca32_and_6_11_y0;
  wire h_s_dadda_rca32_and_5_12_y0;
  wire h_s_dadda_rca32_fa78_y2;
  wire h_s_dadda_rca32_fa78_y4;
  wire h_s_dadda_rca32_and_4_13_y0;
  wire h_s_dadda_rca32_and_3_14_y0;
  wire h_s_dadda_rca32_and_2_15_y0;
  wire h_s_dadda_rca32_fa79_y2;
  wire h_s_dadda_rca32_fa79_y4;
  wire h_s_dadda_rca32_and_1_16_y0;
  wire h_s_dadda_rca32_and_0_17_y0;
  wire h_s_dadda_rca32_fa80_y2;
  wire h_s_dadda_rca32_fa80_y4;
  wire h_s_dadda_rca32_fa81_y2;
  wire h_s_dadda_rca32_fa81_y4;
  wire h_s_dadda_rca32_ha15_y0;
  wire h_s_dadda_rca32_ha15_y1;
  wire h_s_dadda_rca32_fa82_y2;
  wire h_s_dadda_rca32_fa82_y4;
  wire h_s_dadda_rca32_fa83_y2;
  wire h_s_dadda_rca32_fa83_y4;
  wire h_s_dadda_rca32_fa84_y2;
  wire h_s_dadda_rca32_fa84_y4;
  wire h_s_dadda_rca32_fa85_y2;
  wire h_s_dadda_rca32_fa85_y4;
  wire h_s_dadda_rca32_and_18_0_y0;
  wire h_s_dadda_rca32_and_17_1_y0;
  wire h_s_dadda_rca32_and_16_2_y0;
  wire h_s_dadda_rca32_fa86_y2;
  wire h_s_dadda_rca32_fa86_y4;
  wire h_s_dadda_rca32_and_15_3_y0;
  wire h_s_dadda_rca32_and_14_4_y0;
  wire h_s_dadda_rca32_and_13_5_y0;
  wire h_s_dadda_rca32_fa87_y2;
  wire h_s_dadda_rca32_fa87_y4;
  wire h_s_dadda_rca32_and_12_6_y0;
  wire h_s_dadda_rca32_and_11_7_y0;
  wire h_s_dadda_rca32_and_10_8_y0;
  wire h_s_dadda_rca32_fa88_y2;
  wire h_s_dadda_rca32_fa88_y4;
  wire h_s_dadda_rca32_and_9_9_y0;
  wire h_s_dadda_rca32_and_8_10_y0;
  wire h_s_dadda_rca32_and_7_11_y0;
  wire h_s_dadda_rca32_fa89_y2;
  wire h_s_dadda_rca32_fa89_y4;
  wire h_s_dadda_rca32_and_6_12_y0;
  wire h_s_dadda_rca32_and_5_13_y0;
  wire h_s_dadda_rca32_and_4_14_y0;
  wire h_s_dadda_rca32_fa90_y2;
  wire h_s_dadda_rca32_fa90_y4;
  wire h_s_dadda_rca32_and_3_15_y0;
  wire h_s_dadda_rca32_and_2_16_y0;
  wire h_s_dadda_rca32_and_1_17_y0;
  wire h_s_dadda_rca32_fa91_y2;
  wire h_s_dadda_rca32_fa91_y4;
  wire h_s_dadda_rca32_and_0_18_y0;
  wire h_s_dadda_rca32_fa92_y2;
  wire h_s_dadda_rca32_fa92_y4;
  wire h_s_dadda_rca32_fa93_y2;
  wire h_s_dadda_rca32_fa93_y4;
  wire h_s_dadda_rca32_ha16_y0;
  wire h_s_dadda_rca32_ha16_y1;
  wire h_s_dadda_rca32_fa94_y2;
  wire h_s_dadda_rca32_fa94_y4;
  wire h_s_dadda_rca32_fa95_y2;
  wire h_s_dadda_rca32_fa95_y4;
  wire h_s_dadda_rca32_fa96_y2;
  wire h_s_dadda_rca32_fa96_y4;
  wire h_s_dadda_rca32_fa97_y2;
  wire h_s_dadda_rca32_fa97_y4;
  wire h_s_dadda_rca32_and_19_0_y0;
  wire h_s_dadda_rca32_and_18_1_y0;
  wire h_s_dadda_rca32_fa98_y2;
  wire h_s_dadda_rca32_fa98_y4;
  wire h_s_dadda_rca32_and_17_2_y0;
  wire h_s_dadda_rca32_and_16_3_y0;
  wire h_s_dadda_rca32_and_15_4_y0;
  wire h_s_dadda_rca32_fa99_y2;
  wire h_s_dadda_rca32_fa99_y4;
  wire h_s_dadda_rca32_and_14_5_y0;
  wire h_s_dadda_rca32_and_13_6_y0;
  wire h_s_dadda_rca32_and_12_7_y0;
  wire h_s_dadda_rca32_fa100_y2;
  wire h_s_dadda_rca32_fa100_y4;
  wire h_s_dadda_rca32_and_11_8_y0;
  wire h_s_dadda_rca32_and_10_9_y0;
  wire h_s_dadda_rca32_and_9_10_y0;
  wire h_s_dadda_rca32_fa101_y2;
  wire h_s_dadda_rca32_fa101_y4;
  wire h_s_dadda_rca32_and_8_11_y0;
  wire h_s_dadda_rca32_and_7_12_y0;
  wire h_s_dadda_rca32_and_6_13_y0;
  wire h_s_dadda_rca32_fa102_y2;
  wire h_s_dadda_rca32_fa102_y4;
  wire h_s_dadda_rca32_and_5_14_y0;
  wire h_s_dadda_rca32_and_4_15_y0;
  wire h_s_dadda_rca32_and_3_16_y0;
  wire h_s_dadda_rca32_fa103_y2;
  wire h_s_dadda_rca32_fa103_y4;
  wire h_s_dadda_rca32_and_2_17_y0;
  wire h_s_dadda_rca32_and_1_18_y0;
  wire h_s_dadda_rca32_and_0_19_y0;
  wire h_s_dadda_rca32_fa104_y2;
  wire h_s_dadda_rca32_fa104_y4;
  wire h_s_dadda_rca32_fa105_y2;
  wire h_s_dadda_rca32_fa105_y4;
  wire h_s_dadda_rca32_fa106_y2;
  wire h_s_dadda_rca32_fa106_y4;
  wire h_s_dadda_rca32_ha17_y0;
  wire h_s_dadda_rca32_ha17_y1;
  wire h_s_dadda_rca32_fa107_y2;
  wire h_s_dadda_rca32_fa107_y4;
  wire h_s_dadda_rca32_fa108_y2;
  wire h_s_dadda_rca32_fa108_y4;
  wire h_s_dadda_rca32_fa109_y2;
  wire h_s_dadda_rca32_fa109_y4;
  wire h_s_dadda_rca32_fa110_y2;
  wire h_s_dadda_rca32_fa110_y4;
  wire h_s_dadda_rca32_and_20_0_y0;
  wire h_s_dadda_rca32_fa111_y2;
  wire h_s_dadda_rca32_fa111_y4;
  wire h_s_dadda_rca32_and_19_1_y0;
  wire h_s_dadda_rca32_and_18_2_y0;
  wire h_s_dadda_rca32_and_17_3_y0;
  wire h_s_dadda_rca32_fa112_y2;
  wire h_s_dadda_rca32_fa112_y4;
  wire h_s_dadda_rca32_and_16_4_y0;
  wire h_s_dadda_rca32_and_15_5_y0;
  wire h_s_dadda_rca32_and_14_6_y0;
  wire h_s_dadda_rca32_fa113_y2;
  wire h_s_dadda_rca32_fa113_y4;
  wire h_s_dadda_rca32_and_13_7_y0;
  wire h_s_dadda_rca32_and_12_8_y0;
  wire h_s_dadda_rca32_and_11_9_y0;
  wire h_s_dadda_rca32_fa114_y2;
  wire h_s_dadda_rca32_fa114_y4;
  wire h_s_dadda_rca32_and_10_10_y0;
  wire h_s_dadda_rca32_and_9_11_y0;
  wire h_s_dadda_rca32_and_8_12_y0;
  wire h_s_dadda_rca32_fa115_y2;
  wire h_s_dadda_rca32_fa115_y4;
  wire h_s_dadda_rca32_and_7_13_y0;
  wire h_s_dadda_rca32_and_6_14_y0;
  wire h_s_dadda_rca32_and_5_15_y0;
  wire h_s_dadda_rca32_fa116_y2;
  wire h_s_dadda_rca32_fa116_y4;
  wire h_s_dadda_rca32_and_4_16_y0;
  wire h_s_dadda_rca32_and_3_17_y0;
  wire h_s_dadda_rca32_and_2_18_y0;
  wire h_s_dadda_rca32_fa117_y2;
  wire h_s_dadda_rca32_fa117_y4;
  wire h_s_dadda_rca32_and_1_19_y0;
  wire h_s_dadda_rca32_and_0_20_y0;
  wire h_s_dadda_rca32_fa118_y2;
  wire h_s_dadda_rca32_fa118_y4;
  wire h_s_dadda_rca32_fa119_y2;
  wire h_s_dadda_rca32_fa119_y4;
  wire h_s_dadda_rca32_fa120_y2;
  wire h_s_dadda_rca32_fa120_y4;
  wire h_s_dadda_rca32_ha18_y0;
  wire h_s_dadda_rca32_ha18_y1;
  wire h_s_dadda_rca32_fa121_y2;
  wire h_s_dadda_rca32_fa121_y4;
  wire h_s_dadda_rca32_fa122_y2;
  wire h_s_dadda_rca32_fa122_y4;
  wire h_s_dadda_rca32_fa123_y2;
  wire h_s_dadda_rca32_fa123_y4;
  wire h_s_dadda_rca32_fa124_y2;
  wire h_s_dadda_rca32_fa124_y4;
  wire h_s_dadda_rca32_fa125_y2;
  wire h_s_dadda_rca32_fa125_y4;
  wire h_s_dadda_rca32_and_21_0_y0;
  wire h_s_dadda_rca32_and_20_1_y0;
  wire h_s_dadda_rca32_and_19_2_y0;
  wire h_s_dadda_rca32_fa126_y2;
  wire h_s_dadda_rca32_fa126_y4;
  wire h_s_dadda_rca32_and_18_3_y0;
  wire h_s_dadda_rca32_and_17_4_y0;
  wire h_s_dadda_rca32_and_16_5_y0;
  wire h_s_dadda_rca32_fa127_y2;
  wire h_s_dadda_rca32_fa127_y4;
  wire h_s_dadda_rca32_and_15_6_y0;
  wire h_s_dadda_rca32_and_14_7_y0;
  wire h_s_dadda_rca32_and_13_8_y0;
  wire h_s_dadda_rca32_fa128_y2;
  wire h_s_dadda_rca32_fa128_y4;
  wire h_s_dadda_rca32_and_12_9_y0;
  wire h_s_dadda_rca32_and_11_10_y0;
  wire h_s_dadda_rca32_and_10_11_y0;
  wire h_s_dadda_rca32_fa129_y2;
  wire h_s_dadda_rca32_fa129_y4;
  wire h_s_dadda_rca32_and_9_12_y0;
  wire h_s_dadda_rca32_and_8_13_y0;
  wire h_s_dadda_rca32_and_7_14_y0;
  wire h_s_dadda_rca32_fa130_y2;
  wire h_s_dadda_rca32_fa130_y4;
  wire h_s_dadda_rca32_and_6_15_y0;
  wire h_s_dadda_rca32_and_5_16_y0;
  wire h_s_dadda_rca32_and_4_17_y0;
  wire h_s_dadda_rca32_fa131_y2;
  wire h_s_dadda_rca32_fa131_y4;
  wire h_s_dadda_rca32_and_3_18_y0;
  wire h_s_dadda_rca32_and_2_19_y0;
  wire h_s_dadda_rca32_and_1_20_y0;
  wire h_s_dadda_rca32_fa132_y2;
  wire h_s_dadda_rca32_fa132_y4;
  wire h_s_dadda_rca32_and_0_21_y0;
  wire h_s_dadda_rca32_fa133_y2;
  wire h_s_dadda_rca32_fa133_y4;
  wire h_s_dadda_rca32_fa134_y2;
  wire h_s_dadda_rca32_fa134_y4;
  wire h_s_dadda_rca32_fa135_y2;
  wire h_s_dadda_rca32_fa135_y4;
  wire h_s_dadda_rca32_ha19_y0;
  wire h_s_dadda_rca32_ha19_y1;
  wire h_s_dadda_rca32_fa136_y2;
  wire h_s_dadda_rca32_fa136_y4;
  wire h_s_dadda_rca32_fa137_y2;
  wire h_s_dadda_rca32_fa137_y4;
  wire h_s_dadda_rca32_fa138_y2;
  wire h_s_dadda_rca32_fa138_y4;
  wire h_s_dadda_rca32_fa139_y2;
  wire h_s_dadda_rca32_fa139_y4;
  wire h_s_dadda_rca32_fa140_y2;
  wire h_s_dadda_rca32_fa140_y4;
  wire h_s_dadda_rca32_and_22_0_y0;
  wire h_s_dadda_rca32_and_21_1_y0;
  wire h_s_dadda_rca32_fa141_y2;
  wire h_s_dadda_rca32_fa141_y4;
  wire h_s_dadda_rca32_and_20_2_y0;
  wire h_s_dadda_rca32_and_19_3_y0;
  wire h_s_dadda_rca32_and_18_4_y0;
  wire h_s_dadda_rca32_fa142_y2;
  wire h_s_dadda_rca32_fa142_y4;
  wire h_s_dadda_rca32_and_17_5_y0;
  wire h_s_dadda_rca32_and_16_6_y0;
  wire h_s_dadda_rca32_and_15_7_y0;
  wire h_s_dadda_rca32_fa143_y2;
  wire h_s_dadda_rca32_fa143_y4;
  wire h_s_dadda_rca32_and_14_8_y0;
  wire h_s_dadda_rca32_and_13_9_y0;
  wire h_s_dadda_rca32_and_12_10_y0;
  wire h_s_dadda_rca32_fa144_y2;
  wire h_s_dadda_rca32_fa144_y4;
  wire h_s_dadda_rca32_and_11_11_y0;
  wire h_s_dadda_rca32_and_10_12_y0;
  wire h_s_dadda_rca32_and_9_13_y0;
  wire h_s_dadda_rca32_fa145_y2;
  wire h_s_dadda_rca32_fa145_y4;
  wire h_s_dadda_rca32_and_8_14_y0;
  wire h_s_dadda_rca32_and_7_15_y0;
  wire h_s_dadda_rca32_and_6_16_y0;
  wire h_s_dadda_rca32_fa146_y2;
  wire h_s_dadda_rca32_fa146_y4;
  wire h_s_dadda_rca32_and_5_17_y0;
  wire h_s_dadda_rca32_and_4_18_y0;
  wire h_s_dadda_rca32_and_3_19_y0;
  wire h_s_dadda_rca32_fa147_y2;
  wire h_s_dadda_rca32_fa147_y4;
  wire h_s_dadda_rca32_and_2_20_y0;
  wire h_s_dadda_rca32_and_1_21_y0;
  wire h_s_dadda_rca32_and_0_22_y0;
  wire h_s_dadda_rca32_fa148_y2;
  wire h_s_dadda_rca32_fa148_y4;
  wire h_s_dadda_rca32_fa149_y2;
  wire h_s_dadda_rca32_fa149_y4;
  wire h_s_dadda_rca32_fa150_y2;
  wire h_s_dadda_rca32_fa150_y4;
  wire h_s_dadda_rca32_fa151_y2;
  wire h_s_dadda_rca32_fa151_y4;
  wire h_s_dadda_rca32_ha20_y0;
  wire h_s_dadda_rca32_ha20_y1;
  wire h_s_dadda_rca32_fa152_y2;
  wire h_s_dadda_rca32_fa152_y4;
  wire h_s_dadda_rca32_fa153_y2;
  wire h_s_dadda_rca32_fa153_y4;
  wire h_s_dadda_rca32_fa154_y2;
  wire h_s_dadda_rca32_fa154_y4;
  wire h_s_dadda_rca32_fa155_y2;
  wire h_s_dadda_rca32_fa155_y4;
  wire h_s_dadda_rca32_fa156_y2;
  wire h_s_dadda_rca32_fa156_y4;
  wire h_s_dadda_rca32_and_23_0_y0;
  wire h_s_dadda_rca32_fa157_y2;
  wire h_s_dadda_rca32_fa157_y4;
  wire h_s_dadda_rca32_and_22_1_y0;
  wire h_s_dadda_rca32_and_21_2_y0;
  wire h_s_dadda_rca32_and_20_3_y0;
  wire h_s_dadda_rca32_fa158_y2;
  wire h_s_dadda_rca32_fa158_y4;
  wire h_s_dadda_rca32_and_19_4_y0;
  wire h_s_dadda_rca32_and_18_5_y0;
  wire h_s_dadda_rca32_and_17_6_y0;
  wire h_s_dadda_rca32_fa159_y2;
  wire h_s_dadda_rca32_fa159_y4;
  wire h_s_dadda_rca32_and_16_7_y0;
  wire h_s_dadda_rca32_and_15_8_y0;
  wire h_s_dadda_rca32_and_14_9_y0;
  wire h_s_dadda_rca32_fa160_y2;
  wire h_s_dadda_rca32_fa160_y4;
  wire h_s_dadda_rca32_and_13_10_y0;
  wire h_s_dadda_rca32_and_12_11_y0;
  wire h_s_dadda_rca32_and_11_12_y0;
  wire h_s_dadda_rca32_fa161_y2;
  wire h_s_dadda_rca32_fa161_y4;
  wire h_s_dadda_rca32_and_10_13_y0;
  wire h_s_dadda_rca32_and_9_14_y0;
  wire h_s_dadda_rca32_and_8_15_y0;
  wire h_s_dadda_rca32_fa162_y2;
  wire h_s_dadda_rca32_fa162_y4;
  wire h_s_dadda_rca32_and_7_16_y0;
  wire h_s_dadda_rca32_and_6_17_y0;
  wire h_s_dadda_rca32_and_5_18_y0;
  wire h_s_dadda_rca32_fa163_y2;
  wire h_s_dadda_rca32_fa163_y4;
  wire h_s_dadda_rca32_and_4_19_y0;
  wire h_s_dadda_rca32_and_3_20_y0;
  wire h_s_dadda_rca32_and_2_21_y0;
  wire h_s_dadda_rca32_fa164_y2;
  wire h_s_dadda_rca32_fa164_y4;
  wire h_s_dadda_rca32_and_1_22_y0;
  wire h_s_dadda_rca32_and_0_23_y0;
  wire h_s_dadda_rca32_fa165_y2;
  wire h_s_dadda_rca32_fa165_y4;
  wire h_s_dadda_rca32_fa166_y2;
  wire h_s_dadda_rca32_fa166_y4;
  wire h_s_dadda_rca32_fa167_y2;
  wire h_s_dadda_rca32_fa167_y4;
  wire h_s_dadda_rca32_fa168_y2;
  wire h_s_dadda_rca32_fa168_y4;
  wire h_s_dadda_rca32_ha21_y0;
  wire h_s_dadda_rca32_ha21_y1;
  wire h_s_dadda_rca32_fa169_y2;
  wire h_s_dadda_rca32_fa169_y4;
  wire h_s_dadda_rca32_fa170_y2;
  wire h_s_dadda_rca32_fa170_y4;
  wire h_s_dadda_rca32_fa171_y2;
  wire h_s_dadda_rca32_fa171_y4;
  wire h_s_dadda_rca32_fa172_y2;
  wire h_s_dadda_rca32_fa172_y4;
  wire h_s_dadda_rca32_fa173_y2;
  wire h_s_dadda_rca32_fa173_y4;
  wire h_s_dadda_rca32_fa174_y2;
  wire h_s_dadda_rca32_fa174_y4;
  wire h_s_dadda_rca32_and_24_0_y0;
  wire h_s_dadda_rca32_and_23_1_y0;
  wire h_s_dadda_rca32_and_22_2_y0;
  wire h_s_dadda_rca32_fa175_y2;
  wire h_s_dadda_rca32_fa175_y4;
  wire h_s_dadda_rca32_and_21_3_y0;
  wire h_s_dadda_rca32_and_20_4_y0;
  wire h_s_dadda_rca32_and_19_5_y0;
  wire h_s_dadda_rca32_fa176_y2;
  wire h_s_dadda_rca32_fa176_y4;
  wire h_s_dadda_rca32_and_18_6_y0;
  wire h_s_dadda_rca32_and_17_7_y0;
  wire h_s_dadda_rca32_and_16_8_y0;
  wire h_s_dadda_rca32_fa177_y2;
  wire h_s_dadda_rca32_fa177_y4;
  wire h_s_dadda_rca32_and_15_9_y0;
  wire h_s_dadda_rca32_and_14_10_y0;
  wire h_s_dadda_rca32_and_13_11_y0;
  wire h_s_dadda_rca32_fa178_y2;
  wire h_s_dadda_rca32_fa178_y4;
  wire h_s_dadda_rca32_and_12_12_y0;
  wire h_s_dadda_rca32_and_11_13_y0;
  wire h_s_dadda_rca32_and_10_14_y0;
  wire h_s_dadda_rca32_fa179_y2;
  wire h_s_dadda_rca32_fa179_y4;
  wire h_s_dadda_rca32_and_9_15_y0;
  wire h_s_dadda_rca32_and_8_16_y0;
  wire h_s_dadda_rca32_and_7_17_y0;
  wire h_s_dadda_rca32_fa180_y2;
  wire h_s_dadda_rca32_fa180_y4;
  wire h_s_dadda_rca32_and_6_18_y0;
  wire h_s_dadda_rca32_and_5_19_y0;
  wire h_s_dadda_rca32_and_4_20_y0;
  wire h_s_dadda_rca32_fa181_y2;
  wire h_s_dadda_rca32_fa181_y4;
  wire h_s_dadda_rca32_and_3_21_y0;
  wire h_s_dadda_rca32_and_2_22_y0;
  wire h_s_dadda_rca32_and_1_23_y0;
  wire h_s_dadda_rca32_fa182_y2;
  wire h_s_dadda_rca32_fa182_y4;
  wire h_s_dadda_rca32_and_0_24_y0;
  wire h_s_dadda_rca32_fa183_y2;
  wire h_s_dadda_rca32_fa183_y4;
  wire h_s_dadda_rca32_fa184_y2;
  wire h_s_dadda_rca32_fa184_y4;
  wire h_s_dadda_rca32_fa185_y2;
  wire h_s_dadda_rca32_fa185_y4;
  wire h_s_dadda_rca32_fa186_y2;
  wire h_s_dadda_rca32_fa186_y4;
  wire h_s_dadda_rca32_ha22_y0;
  wire h_s_dadda_rca32_ha22_y1;
  wire h_s_dadda_rca32_fa187_y2;
  wire h_s_dadda_rca32_fa187_y4;
  wire h_s_dadda_rca32_fa188_y2;
  wire h_s_dadda_rca32_fa188_y4;
  wire h_s_dadda_rca32_fa189_y2;
  wire h_s_dadda_rca32_fa189_y4;
  wire h_s_dadda_rca32_fa190_y2;
  wire h_s_dadda_rca32_fa190_y4;
  wire h_s_dadda_rca32_fa191_y2;
  wire h_s_dadda_rca32_fa191_y4;
  wire h_s_dadda_rca32_fa192_y2;
  wire h_s_dadda_rca32_fa192_y4;
  wire h_s_dadda_rca32_and_25_0_y0;
  wire h_s_dadda_rca32_and_24_1_y0;
  wire h_s_dadda_rca32_fa193_y2;
  wire h_s_dadda_rca32_fa193_y4;
  wire h_s_dadda_rca32_and_23_2_y0;
  wire h_s_dadda_rca32_and_22_3_y0;
  wire h_s_dadda_rca32_and_21_4_y0;
  wire h_s_dadda_rca32_fa194_y2;
  wire h_s_dadda_rca32_fa194_y4;
  wire h_s_dadda_rca32_and_20_5_y0;
  wire h_s_dadda_rca32_and_19_6_y0;
  wire h_s_dadda_rca32_and_18_7_y0;
  wire h_s_dadda_rca32_fa195_y2;
  wire h_s_dadda_rca32_fa195_y4;
  wire h_s_dadda_rca32_and_17_8_y0;
  wire h_s_dadda_rca32_and_16_9_y0;
  wire h_s_dadda_rca32_and_15_10_y0;
  wire h_s_dadda_rca32_fa196_y2;
  wire h_s_dadda_rca32_fa196_y4;
  wire h_s_dadda_rca32_and_14_11_y0;
  wire h_s_dadda_rca32_and_13_12_y0;
  wire h_s_dadda_rca32_and_12_13_y0;
  wire h_s_dadda_rca32_fa197_y2;
  wire h_s_dadda_rca32_fa197_y4;
  wire h_s_dadda_rca32_and_11_14_y0;
  wire h_s_dadda_rca32_and_10_15_y0;
  wire h_s_dadda_rca32_and_9_16_y0;
  wire h_s_dadda_rca32_fa198_y2;
  wire h_s_dadda_rca32_fa198_y4;
  wire h_s_dadda_rca32_and_8_17_y0;
  wire h_s_dadda_rca32_and_7_18_y0;
  wire h_s_dadda_rca32_and_6_19_y0;
  wire h_s_dadda_rca32_fa199_y2;
  wire h_s_dadda_rca32_fa199_y4;
  wire h_s_dadda_rca32_and_5_20_y0;
  wire h_s_dadda_rca32_and_4_21_y0;
  wire h_s_dadda_rca32_and_3_22_y0;
  wire h_s_dadda_rca32_fa200_y2;
  wire h_s_dadda_rca32_fa200_y4;
  wire h_s_dadda_rca32_and_2_23_y0;
  wire h_s_dadda_rca32_and_1_24_y0;
  wire h_s_dadda_rca32_and_0_25_y0;
  wire h_s_dadda_rca32_fa201_y2;
  wire h_s_dadda_rca32_fa201_y4;
  wire h_s_dadda_rca32_fa202_y2;
  wire h_s_dadda_rca32_fa202_y4;
  wire h_s_dadda_rca32_fa203_y2;
  wire h_s_dadda_rca32_fa203_y4;
  wire h_s_dadda_rca32_fa204_y2;
  wire h_s_dadda_rca32_fa204_y4;
  wire h_s_dadda_rca32_fa205_y2;
  wire h_s_dadda_rca32_fa205_y4;
  wire h_s_dadda_rca32_ha23_y0;
  wire h_s_dadda_rca32_ha23_y1;
  wire h_s_dadda_rca32_fa206_y2;
  wire h_s_dadda_rca32_fa206_y4;
  wire h_s_dadda_rca32_fa207_y2;
  wire h_s_dadda_rca32_fa207_y4;
  wire h_s_dadda_rca32_fa208_y2;
  wire h_s_dadda_rca32_fa208_y4;
  wire h_s_dadda_rca32_fa209_y2;
  wire h_s_dadda_rca32_fa209_y4;
  wire h_s_dadda_rca32_fa210_y2;
  wire h_s_dadda_rca32_fa210_y4;
  wire h_s_dadda_rca32_fa211_y2;
  wire h_s_dadda_rca32_fa211_y4;
  wire h_s_dadda_rca32_and_26_0_y0;
  wire h_s_dadda_rca32_fa212_y2;
  wire h_s_dadda_rca32_fa212_y4;
  wire h_s_dadda_rca32_and_25_1_y0;
  wire h_s_dadda_rca32_and_24_2_y0;
  wire h_s_dadda_rca32_and_23_3_y0;
  wire h_s_dadda_rca32_fa213_y2;
  wire h_s_dadda_rca32_fa213_y4;
  wire h_s_dadda_rca32_and_22_4_y0;
  wire h_s_dadda_rca32_and_21_5_y0;
  wire h_s_dadda_rca32_and_20_6_y0;
  wire h_s_dadda_rca32_fa214_y2;
  wire h_s_dadda_rca32_fa214_y4;
  wire h_s_dadda_rca32_and_19_7_y0;
  wire h_s_dadda_rca32_and_18_8_y0;
  wire h_s_dadda_rca32_and_17_9_y0;
  wire h_s_dadda_rca32_fa215_y2;
  wire h_s_dadda_rca32_fa215_y4;
  wire h_s_dadda_rca32_and_16_10_y0;
  wire h_s_dadda_rca32_and_15_11_y0;
  wire h_s_dadda_rca32_and_14_12_y0;
  wire h_s_dadda_rca32_fa216_y2;
  wire h_s_dadda_rca32_fa216_y4;
  wire h_s_dadda_rca32_and_13_13_y0;
  wire h_s_dadda_rca32_and_12_14_y0;
  wire h_s_dadda_rca32_and_11_15_y0;
  wire h_s_dadda_rca32_fa217_y2;
  wire h_s_dadda_rca32_fa217_y4;
  wire h_s_dadda_rca32_and_10_16_y0;
  wire h_s_dadda_rca32_and_9_17_y0;
  wire h_s_dadda_rca32_and_8_18_y0;
  wire h_s_dadda_rca32_fa218_y2;
  wire h_s_dadda_rca32_fa218_y4;
  wire h_s_dadda_rca32_and_7_19_y0;
  wire h_s_dadda_rca32_and_6_20_y0;
  wire h_s_dadda_rca32_and_5_21_y0;
  wire h_s_dadda_rca32_fa219_y2;
  wire h_s_dadda_rca32_fa219_y4;
  wire h_s_dadda_rca32_and_4_22_y0;
  wire h_s_dadda_rca32_and_3_23_y0;
  wire h_s_dadda_rca32_and_2_24_y0;
  wire h_s_dadda_rca32_fa220_y2;
  wire h_s_dadda_rca32_fa220_y4;
  wire h_s_dadda_rca32_and_1_25_y0;
  wire h_s_dadda_rca32_and_0_26_y0;
  wire h_s_dadda_rca32_fa221_y2;
  wire h_s_dadda_rca32_fa221_y4;
  wire h_s_dadda_rca32_fa222_y2;
  wire h_s_dadda_rca32_fa222_y4;
  wire h_s_dadda_rca32_fa223_y2;
  wire h_s_dadda_rca32_fa223_y4;
  wire h_s_dadda_rca32_fa224_y2;
  wire h_s_dadda_rca32_fa224_y4;
  wire h_s_dadda_rca32_fa225_y2;
  wire h_s_dadda_rca32_fa225_y4;
  wire h_s_dadda_rca32_ha24_y0;
  wire h_s_dadda_rca32_ha24_y1;
  wire h_s_dadda_rca32_fa226_y2;
  wire h_s_dadda_rca32_fa226_y4;
  wire h_s_dadda_rca32_fa227_y2;
  wire h_s_dadda_rca32_fa227_y4;
  wire h_s_dadda_rca32_fa228_y2;
  wire h_s_dadda_rca32_fa228_y4;
  wire h_s_dadda_rca32_fa229_y2;
  wire h_s_dadda_rca32_fa229_y4;
  wire h_s_dadda_rca32_fa230_y2;
  wire h_s_dadda_rca32_fa230_y4;
  wire h_s_dadda_rca32_fa231_y2;
  wire h_s_dadda_rca32_fa231_y4;
  wire h_s_dadda_rca32_fa232_y2;
  wire h_s_dadda_rca32_fa232_y4;
  wire h_s_dadda_rca32_and_27_0_y0;
  wire h_s_dadda_rca32_and_26_1_y0;
  wire h_s_dadda_rca32_and_25_2_y0;
  wire h_s_dadda_rca32_fa233_y2;
  wire h_s_dadda_rca32_fa233_y4;
  wire h_s_dadda_rca32_and_24_3_y0;
  wire h_s_dadda_rca32_and_23_4_y0;
  wire h_s_dadda_rca32_and_22_5_y0;
  wire h_s_dadda_rca32_fa234_y2;
  wire h_s_dadda_rca32_fa234_y4;
  wire h_s_dadda_rca32_and_21_6_y0;
  wire h_s_dadda_rca32_and_20_7_y0;
  wire h_s_dadda_rca32_and_19_8_y0;
  wire h_s_dadda_rca32_fa235_y2;
  wire h_s_dadda_rca32_fa235_y4;
  wire h_s_dadda_rca32_and_18_9_y0;
  wire h_s_dadda_rca32_and_17_10_y0;
  wire h_s_dadda_rca32_and_16_11_y0;
  wire h_s_dadda_rca32_fa236_y2;
  wire h_s_dadda_rca32_fa236_y4;
  wire h_s_dadda_rca32_and_15_12_y0;
  wire h_s_dadda_rca32_and_14_13_y0;
  wire h_s_dadda_rca32_and_13_14_y0;
  wire h_s_dadda_rca32_fa237_y2;
  wire h_s_dadda_rca32_fa237_y4;
  wire h_s_dadda_rca32_and_12_15_y0;
  wire h_s_dadda_rca32_and_11_16_y0;
  wire h_s_dadda_rca32_and_10_17_y0;
  wire h_s_dadda_rca32_fa238_y2;
  wire h_s_dadda_rca32_fa238_y4;
  wire h_s_dadda_rca32_and_9_18_y0;
  wire h_s_dadda_rca32_and_8_19_y0;
  wire h_s_dadda_rca32_and_7_20_y0;
  wire h_s_dadda_rca32_fa239_y2;
  wire h_s_dadda_rca32_fa239_y4;
  wire h_s_dadda_rca32_and_6_21_y0;
  wire h_s_dadda_rca32_and_5_22_y0;
  wire h_s_dadda_rca32_and_4_23_y0;
  wire h_s_dadda_rca32_fa240_y2;
  wire h_s_dadda_rca32_fa240_y4;
  wire h_s_dadda_rca32_and_3_24_y0;
  wire h_s_dadda_rca32_and_2_25_y0;
  wire h_s_dadda_rca32_and_1_26_y0;
  wire h_s_dadda_rca32_fa241_y2;
  wire h_s_dadda_rca32_fa241_y4;
  wire h_s_dadda_rca32_and_0_27_y0;
  wire h_s_dadda_rca32_fa242_y2;
  wire h_s_dadda_rca32_fa242_y4;
  wire h_s_dadda_rca32_fa243_y2;
  wire h_s_dadda_rca32_fa243_y4;
  wire h_s_dadda_rca32_fa244_y2;
  wire h_s_dadda_rca32_fa244_y4;
  wire h_s_dadda_rca32_fa245_y2;
  wire h_s_dadda_rca32_fa245_y4;
  wire h_s_dadda_rca32_fa246_y2;
  wire h_s_dadda_rca32_fa246_y4;
  wire h_s_dadda_rca32_ha25_y0;
  wire h_s_dadda_rca32_ha25_y1;
  wire h_s_dadda_rca32_fa247_y2;
  wire h_s_dadda_rca32_fa247_y4;
  wire h_s_dadda_rca32_fa248_y2;
  wire h_s_dadda_rca32_fa248_y4;
  wire h_s_dadda_rca32_fa249_y2;
  wire h_s_dadda_rca32_fa249_y4;
  wire h_s_dadda_rca32_fa250_y2;
  wire h_s_dadda_rca32_fa250_y4;
  wire h_s_dadda_rca32_fa251_y2;
  wire h_s_dadda_rca32_fa251_y4;
  wire h_s_dadda_rca32_fa252_y2;
  wire h_s_dadda_rca32_fa252_y4;
  wire h_s_dadda_rca32_fa253_y2;
  wire h_s_dadda_rca32_fa253_y4;
  wire h_s_dadda_rca32_and_26_2_y0;
  wire h_s_dadda_rca32_and_25_3_y0;
  wire h_s_dadda_rca32_fa254_y2;
  wire h_s_dadda_rca32_fa254_y4;
  wire h_s_dadda_rca32_and_24_4_y0;
  wire h_s_dadda_rca32_and_23_5_y0;
  wire h_s_dadda_rca32_and_22_6_y0;
  wire h_s_dadda_rca32_fa255_y2;
  wire h_s_dadda_rca32_fa255_y4;
  wire h_s_dadda_rca32_and_21_7_y0;
  wire h_s_dadda_rca32_and_20_8_y0;
  wire h_s_dadda_rca32_and_19_9_y0;
  wire h_s_dadda_rca32_fa256_y2;
  wire h_s_dadda_rca32_fa256_y4;
  wire h_s_dadda_rca32_and_18_10_y0;
  wire h_s_dadda_rca32_and_17_11_y0;
  wire h_s_dadda_rca32_and_16_12_y0;
  wire h_s_dadda_rca32_fa257_y2;
  wire h_s_dadda_rca32_fa257_y4;
  wire h_s_dadda_rca32_and_15_13_y0;
  wire h_s_dadda_rca32_and_14_14_y0;
  wire h_s_dadda_rca32_and_13_15_y0;
  wire h_s_dadda_rca32_fa258_y2;
  wire h_s_dadda_rca32_fa258_y4;
  wire h_s_dadda_rca32_and_12_16_y0;
  wire h_s_dadda_rca32_and_11_17_y0;
  wire h_s_dadda_rca32_and_10_18_y0;
  wire h_s_dadda_rca32_fa259_y2;
  wire h_s_dadda_rca32_fa259_y4;
  wire h_s_dadda_rca32_and_9_19_y0;
  wire h_s_dadda_rca32_and_8_20_y0;
  wire h_s_dadda_rca32_and_7_21_y0;
  wire h_s_dadda_rca32_fa260_y2;
  wire h_s_dadda_rca32_fa260_y4;
  wire h_s_dadda_rca32_and_6_22_y0;
  wire h_s_dadda_rca32_and_5_23_y0;
  wire h_s_dadda_rca32_and_4_24_y0;
  wire h_s_dadda_rca32_fa261_y2;
  wire h_s_dadda_rca32_fa261_y4;
  wire h_s_dadda_rca32_and_3_25_y0;
  wire h_s_dadda_rca32_and_2_26_y0;
  wire h_s_dadda_rca32_and_1_27_y0;
  wire h_s_dadda_rca32_fa262_y2;
  wire h_s_dadda_rca32_fa262_y4;
  wire h_s_dadda_rca32_and_0_28_y0;
  wire h_s_dadda_rca32_fa263_y2;
  wire h_s_dadda_rca32_fa263_y4;
  wire h_s_dadda_rca32_fa264_y2;
  wire h_s_dadda_rca32_fa264_y4;
  wire h_s_dadda_rca32_fa265_y2;
  wire h_s_dadda_rca32_fa265_y4;
  wire h_s_dadda_rca32_fa266_y2;
  wire h_s_dadda_rca32_fa266_y4;
  wire h_s_dadda_rca32_fa267_y2;
  wire h_s_dadda_rca32_fa267_y4;
  wire h_s_dadda_rca32_fa268_y2;
  wire h_s_dadda_rca32_fa268_y4;
  wire h_s_dadda_rca32_fa269_y2;
  wire h_s_dadda_rca32_fa269_y4;
  wire h_s_dadda_rca32_fa270_y2;
  wire h_s_dadda_rca32_fa270_y4;
  wire h_s_dadda_rca32_fa271_y2;
  wire h_s_dadda_rca32_fa271_y4;
  wire h_s_dadda_rca32_fa272_y2;
  wire h_s_dadda_rca32_fa272_y4;
  wire h_s_dadda_rca32_fa273_y2;
  wire h_s_dadda_rca32_fa273_y4;
  wire h_s_dadda_rca32_fa274_y2;
  wire h_s_dadda_rca32_fa274_y4;
  wire h_s_dadda_rca32_fa275_y2;
  wire h_s_dadda_rca32_fa275_y4;
  wire h_s_dadda_rca32_and_25_4_y0;
  wire h_s_dadda_rca32_and_24_5_y0;
  wire h_s_dadda_rca32_fa276_y2;
  wire h_s_dadda_rca32_fa276_y4;
  wire h_s_dadda_rca32_and_23_6_y0;
  wire h_s_dadda_rca32_and_22_7_y0;
  wire h_s_dadda_rca32_and_21_8_y0;
  wire h_s_dadda_rca32_fa277_y2;
  wire h_s_dadda_rca32_fa277_y4;
  wire h_s_dadda_rca32_and_20_9_y0;
  wire h_s_dadda_rca32_and_19_10_y0;
  wire h_s_dadda_rca32_and_18_11_y0;
  wire h_s_dadda_rca32_fa278_y2;
  wire h_s_dadda_rca32_fa278_y4;
  wire h_s_dadda_rca32_and_17_12_y0;
  wire h_s_dadda_rca32_and_16_13_y0;
  wire h_s_dadda_rca32_and_15_14_y0;
  wire h_s_dadda_rca32_fa279_y2;
  wire h_s_dadda_rca32_fa279_y4;
  wire h_s_dadda_rca32_and_14_15_y0;
  wire h_s_dadda_rca32_and_13_16_y0;
  wire h_s_dadda_rca32_and_12_17_y0;
  wire h_s_dadda_rca32_fa280_y2;
  wire h_s_dadda_rca32_fa280_y4;
  wire h_s_dadda_rca32_and_11_18_y0;
  wire h_s_dadda_rca32_and_10_19_y0;
  wire h_s_dadda_rca32_and_9_20_y0;
  wire h_s_dadda_rca32_fa281_y2;
  wire h_s_dadda_rca32_fa281_y4;
  wire h_s_dadda_rca32_and_8_21_y0;
  wire h_s_dadda_rca32_and_7_22_y0;
  wire h_s_dadda_rca32_and_6_23_y0;
  wire h_s_dadda_rca32_fa282_y2;
  wire h_s_dadda_rca32_fa282_y4;
  wire h_s_dadda_rca32_and_5_24_y0;
  wire h_s_dadda_rca32_and_4_25_y0;
  wire h_s_dadda_rca32_and_3_26_y0;
  wire h_s_dadda_rca32_fa283_y2;
  wire h_s_dadda_rca32_fa283_y4;
  wire h_s_dadda_rca32_and_2_27_y0;
  wire h_s_dadda_rca32_and_1_28_y0;
  wire h_s_dadda_rca32_and_0_29_y0;
  wire h_s_dadda_rca32_fa284_y2;
  wire h_s_dadda_rca32_fa284_y4;
  wire h_s_dadda_rca32_fa285_y2;
  wire h_s_dadda_rca32_fa285_y4;
  wire h_s_dadda_rca32_fa286_y2;
  wire h_s_dadda_rca32_fa286_y4;
  wire h_s_dadda_rca32_fa287_y2;
  wire h_s_dadda_rca32_fa287_y4;
  wire h_s_dadda_rca32_fa288_y2;
  wire h_s_dadda_rca32_fa288_y4;
  wire h_s_dadda_rca32_fa289_y2;
  wire h_s_dadda_rca32_fa289_y4;
  wire h_s_dadda_rca32_fa290_y2;
  wire h_s_dadda_rca32_fa290_y4;
  wire h_s_dadda_rca32_fa291_y2;
  wire h_s_dadda_rca32_fa291_y4;
  wire h_s_dadda_rca32_fa292_y2;
  wire h_s_dadda_rca32_fa292_y4;
  wire h_s_dadda_rca32_fa293_y2;
  wire h_s_dadda_rca32_fa293_y4;
  wire h_s_dadda_rca32_fa294_y2;
  wire h_s_dadda_rca32_fa294_y4;
  wire h_s_dadda_rca32_fa295_y2;
  wire h_s_dadda_rca32_fa295_y4;
  wire h_s_dadda_rca32_fa296_y2;
  wire h_s_dadda_rca32_fa296_y4;
  wire h_s_dadda_rca32_fa297_y2;
  wire h_s_dadda_rca32_fa297_y4;
  wire h_s_dadda_rca32_and_24_6_y0;
  wire h_s_dadda_rca32_and_23_7_y0;
  wire h_s_dadda_rca32_fa298_y2;
  wire h_s_dadda_rca32_fa298_y4;
  wire h_s_dadda_rca32_and_22_8_y0;
  wire h_s_dadda_rca32_and_21_9_y0;
  wire h_s_dadda_rca32_and_20_10_y0;
  wire h_s_dadda_rca32_fa299_y2;
  wire h_s_dadda_rca32_fa299_y4;
  wire h_s_dadda_rca32_and_19_11_y0;
  wire h_s_dadda_rca32_and_18_12_y0;
  wire h_s_dadda_rca32_and_17_13_y0;
  wire h_s_dadda_rca32_fa300_y2;
  wire h_s_dadda_rca32_fa300_y4;
  wire h_s_dadda_rca32_and_16_14_y0;
  wire h_s_dadda_rca32_and_15_15_y0;
  wire h_s_dadda_rca32_and_14_16_y0;
  wire h_s_dadda_rca32_fa301_y2;
  wire h_s_dadda_rca32_fa301_y4;
  wire h_s_dadda_rca32_and_13_17_y0;
  wire h_s_dadda_rca32_and_12_18_y0;
  wire h_s_dadda_rca32_and_11_19_y0;
  wire h_s_dadda_rca32_fa302_y2;
  wire h_s_dadda_rca32_fa302_y4;
  wire h_s_dadda_rca32_and_10_20_y0;
  wire h_s_dadda_rca32_and_9_21_y0;
  wire h_s_dadda_rca32_and_8_22_y0;
  wire h_s_dadda_rca32_fa303_y2;
  wire h_s_dadda_rca32_fa303_y4;
  wire h_s_dadda_rca32_and_7_23_y0;
  wire h_s_dadda_rca32_and_6_24_y0;
  wire h_s_dadda_rca32_and_5_25_y0;
  wire h_s_dadda_rca32_fa304_y2;
  wire h_s_dadda_rca32_fa304_y4;
  wire h_s_dadda_rca32_and_4_26_y0;
  wire h_s_dadda_rca32_and_3_27_y0;
  wire h_s_dadda_rca32_and_2_28_y0;
  wire h_s_dadda_rca32_fa305_y2;
  wire h_s_dadda_rca32_fa305_y4;
  wire h_s_dadda_rca32_and_1_29_y0;
  wire h_s_dadda_rca32_and_0_30_y0;
  wire h_s_dadda_rca32_fa306_y2;
  wire h_s_dadda_rca32_fa306_y4;
  wire h_s_dadda_rca32_fa307_y2;
  wire h_s_dadda_rca32_fa307_y4;
  wire h_s_dadda_rca32_fa308_y2;
  wire h_s_dadda_rca32_fa308_y4;
  wire h_s_dadda_rca32_fa309_y2;
  wire h_s_dadda_rca32_fa309_y4;
  wire h_s_dadda_rca32_fa310_y2;
  wire h_s_dadda_rca32_fa310_y4;
  wire h_s_dadda_rca32_fa311_y2;
  wire h_s_dadda_rca32_fa311_y4;
  wire h_s_dadda_rca32_fa312_y2;
  wire h_s_dadda_rca32_fa312_y4;
  wire h_s_dadda_rca32_fa313_y2;
  wire h_s_dadda_rca32_fa313_y4;
  wire h_s_dadda_rca32_fa314_y2;
  wire h_s_dadda_rca32_fa314_y4;
  wire h_s_dadda_rca32_fa315_y2;
  wire h_s_dadda_rca32_fa315_y4;
  wire h_s_dadda_rca32_fa316_y2;
  wire h_s_dadda_rca32_fa316_y4;
  wire h_s_dadda_rca32_fa317_y2;
  wire h_s_dadda_rca32_fa317_y4;
  wire h_s_dadda_rca32_fa318_y2;
  wire h_s_dadda_rca32_fa318_y4;
  wire h_s_dadda_rca32_fa319_y2;
  wire h_s_dadda_rca32_fa319_y4;
  wire h_s_dadda_rca32_and_23_8_y0;
  wire h_s_dadda_rca32_and_22_9_y0;
  wire h_s_dadda_rca32_fa320_y2;
  wire h_s_dadda_rca32_fa320_y4;
  wire h_s_dadda_rca32_and_21_10_y0;
  wire h_s_dadda_rca32_and_20_11_y0;
  wire h_s_dadda_rca32_and_19_12_y0;
  wire h_s_dadda_rca32_fa321_y2;
  wire h_s_dadda_rca32_fa321_y4;
  wire h_s_dadda_rca32_and_18_13_y0;
  wire h_s_dadda_rca32_and_17_14_y0;
  wire h_s_dadda_rca32_and_16_15_y0;
  wire h_s_dadda_rca32_fa322_y2;
  wire h_s_dadda_rca32_fa322_y4;
  wire h_s_dadda_rca32_and_15_16_y0;
  wire h_s_dadda_rca32_and_14_17_y0;
  wire h_s_dadda_rca32_and_13_18_y0;
  wire h_s_dadda_rca32_fa323_y2;
  wire h_s_dadda_rca32_fa323_y4;
  wire h_s_dadda_rca32_and_12_19_y0;
  wire h_s_dadda_rca32_and_11_20_y0;
  wire h_s_dadda_rca32_and_10_21_y0;
  wire h_s_dadda_rca32_fa324_y2;
  wire h_s_dadda_rca32_fa324_y4;
  wire h_s_dadda_rca32_and_9_22_y0;
  wire h_s_dadda_rca32_and_8_23_y0;
  wire h_s_dadda_rca32_and_7_24_y0;
  wire h_s_dadda_rca32_fa325_y2;
  wire h_s_dadda_rca32_fa325_y4;
  wire h_s_dadda_rca32_and_6_25_y0;
  wire h_s_dadda_rca32_and_5_26_y0;
  wire h_s_dadda_rca32_and_4_27_y0;
  wire h_s_dadda_rca32_fa326_y2;
  wire h_s_dadda_rca32_fa326_y4;
  wire h_s_dadda_rca32_and_3_28_y0;
  wire h_s_dadda_rca32_and_2_29_y0;
  wire h_s_dadda_rca32_and_1_30_y0;
  wire h_s_dadda_rca32_fa327_y2;
  wire h_s_dadda_rca32_fa327_y4;
  wire h_s_dadda_rca32_nand_0_31_y0;
  wire h_s_dadda_rca32_fa328_y2;
  wire h_s_dadda_rca32_fa328_y4;
  wire h_s_dadda_rca32_fa329_y2;
  wire h_s_dadda_rca32_fa329_y4;
  wire h_s_dadda_rca32_fa330_y2;
  wire h_s_dadda_rca32_fa330_y4;
  wire h_s_dadda_rca32_fa331_y2;
  wire h_s_dadda_rca32_fa331_y4;
  wire h_s_dadda_rca32_fa332_y2;
  wire h_s_dadda_rca32_fa332_y4;
  wire h_s_dadda_rca32_fa333_y2;
  wire h_s_dadda_rca32_fa333_y4;
  wire h_s_dadda_rca32_fa334_y2;
  wire h_s_dadda_rca32_fa334_y4;
  wire h_s_dadda_rca32_fa335_y2;
  wire h_s_dadda_rca32_fa335_y4;
  wire h_s_dadda_rca32_fa336_y2;
  wire h_s_dadda_rca32_fa336_y4;
  wire h_s_dadda_rca32_fa337_y2;
  wire h_s_dadda_rca32_fa337_y4;
  wire h_s_dadda_rca32_fa338_y2;
  wire h_s_dadda_rca32_fa338_y4;
  wire h_s_dadda_rca32_fa339_y2;
  wire h_s_dadda_rca32_fa339_y4;
  wire h_s_dadda_rca32_fa340_y2;
  wire h_s_dadda_rca32_fa340_y4;
  wire h_s_dadda_rca32_fa341_y2;
  wire h_s_dadda_rca32_fa341_y4;
  wire h_s_dadda_rca32_and_24_8_y0;
  wire h_s_dadda_rca32_and_23_9_y0;
  wire h_s_dadda_rca32_fa342_y2;
  wire h_s_dadda_rca32_fa342_y4;
  wire h_s_dadda_rca32_and_22_10_y0;
  wire h_s_dadda_rca32_and_21_11_y0;
  wire h_s_dadda_rca32_and_20_12_y0;
  wire h_s_dadda_rca32_fa343_y2;
  wire h_s_dadda_rca32_fa343_y4;
  wire h_s_dadda_rca32_and_19_13_y0;
  wire h_s_dadda_rca32_and_18_14_y0;
  wire h_s_dadda_rca32_and_17_15_y0;
  wire h_s_dadda_rca32_fa344_y2;
  wire h_s_dadda_rca32_fa344_y4;
  wire h_s_dadda_rca32_and_16_16_y0;
  wire h_s_dadda_rca32_and_15_17_y0;
  wire h_s_dadda_rca32_and_14_18_y0;
  wire h_s_dadda_rca32_fa345_y2;
  wire h_s_dadda_rca32_fa345_y4;
  wire h_s_dadda_rca32_and_13_19_y0;
  wire h_s_dadda_rca32_and_12_20_y0;
  wire h_s_dadda_rca32_and_11_21_y0;
  wire h_s_dadda_rca32_fa346_y2;
  wire h_s_dadda_rca32_fa346_y4;
  wire h_s_dadda_rca32_and_10_22_y0;
  wire h_s_dadda_rca32_and_9_23_y0;
  wire h_s_dadda_rca32_and_8_24_y0;
  wire h_s_dadda_rca32_fa347_y2;
  wire h_s_dadda_rca32_fa347_y4;
  wire h_s_dadda_rca32_and_7_25_y0;
  wire h_s_dadda_rca32_and_6_26_y0;
  wire h_s_dadda_rca32_and_5_27_y0;
  wire h_s_dadda_rca32_fa348_y2;
  wire h_s_dadda_rca32_fa348_y4;
  wire h_s_dadda_rca32_and_4_28_y0;
  wire h_s_dadda_rca32_and_3_29_y0;
  wire h_s_dadda_rca32_and_2_30_y0;
  wire h_s_dadda_rca32_fa349_y2;
  wire h_s_dadda_rca32_fa349_y4;
  wire h_s_dadda_rca32_nand_1_31_y0;
  wire h_s_dadda_rca32_fa350_y2;
  wire h_s_dadda_rca32_fa350_y4;
  wire h_s_dadda_rca32_fa351_y2;
  wire h_s_dadda_rca32_fa351_y4;
  wire h_s_dadda_rca32_fa352_y2;
  wire h_s_dadda_rca32_fa352_y4;
  wire h_s_dadda_rca32_fa353_y2;
  wire h_s_dadda_rca32_fa353_y4;
  wire h_s_dadda_rca32_fa354_y2;
  wire h_s_dadda_rca32_fa354_y4;
  wire h_s_dadda_rca32_fa355_y2;
  wire h_s_dadda_rca32_fa355_y4;
  wire h_s_dadda_rca32_fa356_y2;
  wire h_s_dadda_rca32_fa356_y4;
  wire h_s_dadda_rca32_fa357_y2;
  wire h_s_dadda_rca32_fa357_y4;
  wire h_s_dadda_rca32_fa358_y2;
  wire h_s_dadda_rca32_fa358_y4;
  wire h_s_dadda_rca32_fa359_y2;
  wire h_s_dadda_rca32_fa359_y4;
  wire h_s_dadda_rca32_fa360_y2;
  wire h_s_dadda_rca32_fa360_y4;
  wire h_s_dadda_rca32_fa361_y2;
  wire h_s_dadda_rca32_fa361_y4;
  wire h_s_dadda_rca32_fa362_y2;
  wire h_s_dadda_rca32_fa362_y4;
  wire h_s_dadda_rca32_fa363_y2;
  wire h_s_dadda_rca32_fa363_y4;
  wire h_s_dadda_rca32_and_26_7_y0;
  wire h_s_dadda_rca32_and_25_8_y0;
  wire h_s_dadda_rca32_fa364_y2;
  wire h_s_dadda_rca32_fa364_y4;
  wire h_s_dadda_rca32_and_24_9_y0;
  wire h_s_dadda_rca32_and_23_10_y0;
  wire h_s_dadda_rca32_and_22_11_y0;
  wire h_s_dadda_rca32_fa365_y2;
  wire h_s_dadda_rca32_fa365_y4;
  wire h_s_dadda_rca32_and_21_12_y0;
  wire h_s_dadda_rca32_and_20_13_y0;
  wire h_s_dadda_rca32_and_19_14_y0;
  wire h_s_dadda_rca32_fa366_y2;
  wire h_s_dadda_rca32_fa366_y4;
  wire h_s_dadda_rca32_and_18_15_y0;
  wire h_s_dadda_rca32_and_17_16_y0;
  wire h_s_dadda_rca32_and_16_17_y0;
  wire h_s_dadda_rca32_fa367_y2;
  wire h_s_dadda_rca32_fa367_y4;
  wire h_s_dadda_rca32_and_15_18_y0;
  wire h_s_dadda_rca32_and_14_19_y0;
  wire h_s_dadda_rca32_and_13_20_y0;
  wire h_s_dadda_rca32_fa368_y2;
  wire h_s_dadda_rca32_fa368_y4;
  wire h_s_dadda_rca32_and_12_21_y0;
  wire h_s_dadda_rca32_and_11_22_y0;
  wire h_s_dadda_rca32_and_10_23_y0;
  wire h_s_dadda_rca32_fa369_y2;
  wire h_s_dadda_rca32_fa369_y4;
  wire h_s_dadda_rca32_and_9_24_y0;
  wire h_s_dadda_rca32_and_8_25_y0;
  wire h_s_dadda_rca32_and_7_26_y0;
  wire h_s_dadda_rca32_fa370_y2;
  wire h_s_dadda_rca32_fa370_y4;
  wire h_s_dadda_rca32_and_6_27_y0;
  wire h_s_dadda_rca32_and_5_28_y0;
  wire h_s_dadda_rca32_and_4_29_y0;
  wire h_s_dadda_rca32_fa371_y2;
  wire h_s_dadda_rca32_fa371_y4;
  wire h_s_dadda_rca32_and_3_30_y0;
  wire h_s_dadda_rca32_nand_2_31_y0;
  wire h_s_dadda_rca32_fa372_y2;
  wire h_s_dadda_rca32_fa372_y4;
  wire h_s_dadda_rca32_fa373_y2;
  wire h_s_dadda_rca32_fa373_y4;
  wire h_s_dadda_rca32_fa374_y2;
  wire h_s_dadda_rca32_fa374_y4;
  wire h_s_dadda_rca32_fa375_y2;
  wire h_s_dadda_rca32_fa375_y4;
  wire h_s_dadda_rca32_fa376_y2;
  wire h_s_dadda_rca32_fa376_y4;
  wire h_s_dadda_rca32_fa377_y2;
  wire h_s_dadda_rca32_fa377_y4;
  wire h_s_dadda_rca32_fa378_y2;
  wire h_s_dadda_rca32_fa378_y4;
  wire h_s_dadda_rca32_fa379_y2;
  wire h_s_dadda_rca32_fa379_y4;
  wire h_s_dadda_rca32_fa380_y2;
  wire h_s_dadda_rca32_fa380_y4;
  wire h_s_dadda_rca32_fa381_y2;
  wire h_s_dadda_rca32_fa381_y4;
  wire h_s_dadda_rca32_fa382_y2;
  wire h_s_dadda_rca32_fa382_y4;
  wire h_s_dadda_rca32_fa383_y2;
  wire h_s_dadda_rca32_fa383_y4;
  wire h_s_dadda_rca32_fa384_y2;
  wire h_s_dadda_rca32_fa384_y4;
  wire h_s_dadda_rca32_fa385_y2;
  wire h_s_dadda_rca32_fa385_y4;
  wire h_s_dadda_rca32_and_28_6_y0;
  wire h_s_dadda_rca32_and_27_7_y0;
  wire h_s_dadda_rca32_fa386_y2;
  wire h_s_dadda_rca32_fa386_y4;
  wire h_s_dadda_rca32_and_26_8_y0;
  wire h_s_dadda_rca32_and_25_9_y0;
  wire h_s_dadda_rca32_and_24_10_y0;
  wire h_s_dadda_rca32_fa387_y2;
  wire h_s_dadda_rca32_fa387_y4;
  wire h_s_dadda_rca32_and_23_11_y0;
  wire h_s_dadda_rca32_and_22_12_y0;
  wire h_s_dadda_rca32_and_21_13_y0;
  wire h_s_dadda_rca32_fa388_y2;
  wire h_s_dadda_rca32_fa388_y4;
  wire h_s_dadda_rca32_and_20_14_y0;
  wire h_s_dadda_rca32_and_19_15_y0;
  wire h_s_dadda_rca32_and_18_16_y0;
  wire h_s_dadda_rca32_fa389_y2;
  wire h_s_dadda_rca32_fa389_y4;
  wire h_s_dadda_rca32_and_17_17_y0;
  wire h_s_dadda_rca32_and_16_18_y0;
  wire h_s_dadda_rca32_and_15_19_y0;
  wire h_s_dadda_rca32_fa390_y2;
  wire h_s_dadda_rca32_fa390_y4;
  wire h_s_dadda_rca32_and_14_20_y0;
  wire h_s_dadda_rca32_and_13_21_y0;
  wire h_s_dadda_rca32_and_12_22_y0;
  wire h_s_dadda_rca32_fa391_y2;
  wire h_s_dadda_rca32_fa391_y4;
  wire h_s_dadda_rca32_and_11_23_y0;
  wire h_s_dadda_rca32_and_10_24_y0;
  wire h_s_dadda_rca32_and_9_25_y0;
  wire h_s_dadda_rca32_fa392_y2;
  wire h_s_dadda_rca32_fa392_y4;
  wire h_s_dadda_rca32_and_8_26_y0;
  wire h_s_dadda_rca32_and_7_27_y0;
  wire h_s_dadda_rca32_and_6_28_y0;
  wire h_s_dadda_rca32_fa393_y2;
  wire h_s_dadda_rca32_fa393_y4;
  wire h_s_dadda_rca32_and_5_29_y0;
  wire h_s_dadda_rca32_and_4_30_y0;
  wire h_s_dadda_rca32_nand_3_31_y0;
  wire h_s_dadda_rca32_fa394_y2;
  wire h_s_dadda_rca32_fa394_y4;
  wire h_s_dadda_rca32_fa395_y2;
  wire h_s_dadda_rca32_fa395_y4;
  wire h_s_dadda_rca32_fa396_y2;
  wire h_s_dadda_rca32_fa396_y4;
  wire h_s_dadda_rca32_fa397_y2;
  wire h_s_dadda_rca32_fa397_y4;
  wire h_s_dadda_rca32_fa398_y2;
  wire h_s_dadda_rca32_fa398_y4;
  wire h_s_dadda_rca32_fa399_y2;
  wire h_s_dadda_rca32_fa399_y4;
  wire h_s_dadda_rca32_fa400_y2;
  wire h_s_dadda_rca32_fa400_y4;
  wire h_s_dadda_rca32_fa401_y2;
  wire h_s_dadda_rca32_fa401_y4;
  wire h_s_dadda_rca32_fa402_y2;
  wire h_s_dadda_rca32_fa402_y4;
  wire h_s_dadda_rca32_fa403_y2;
  wire h_s_dadda_rca32_fa403_y4;
  wire h_s_dadda_rca32_fa404_y2;
  wire h_s_dadda_rca32_fa404_y4;
  wire h_s_dadda_rca32_fa405_y2;
  wire h_s_dadda_rca32_fa405_y4;
  wire h_s_dadda_rca32_fa406_y2;
  wire h_s_dadda_rca32_fa406_y4;
  wire h_s_dadda_rca32_fa407_y2;
  wire h_s_dadda_rca32_fa407_y4;
  wire h_s_dadda_rca32_and_30_5_y0;
  wire h_s_dadda_rca32_and_29_6_y0;
  wire h_s_dadda_rca32_fa408_y2;
  wire h_s_dadda_rca32_fa408_y4;
  wire h_s_dadda_rca32_and_28_7_y0;
  wire h_s_dadda_rca32_and_27_8_y0;
  wire h_s_dadda_rca32_and_26_9_y0;
  wire h_s_dadda_rca32_fa409_y2;
  wire h_s_dadda_rca32_fa409_y4;
  wire h_s_dadda_rca32_and_25_10_y0;
  wire h_s_dadda_rca32_and_24_11_y0;
  wire h_s_dadda_rca32_and_23_12_y0;
  wire h_s_dadda_rca32_fa410_y2;
  wire h_s_dadda_rca32_fa410_y4;
  wire h_s_dadda_rca32_and_22_13_y0;
  wire h_s_dadda_rca32_and_21_14_y0;
  wire h_s_dadda_rca32_and_20_15_y0;
  wire h_s_dadda_rca32_fa411_y2;
  wire h_s_dadda_rca32_fa411_y4;
  wire h_s_dadda_rca32_and_19_16_y0;
  wire h_s_dadda_rca32_and_18_17_y0;
  wire h_s_dadda_rca32_and_17_18_y0;
  wire h_s_dadda_rca32_fa412_y2;
  wire h_s_dadda_rca32_fa412_y4;
  wire h_s_dadda_rca32_and_16_19_y0;
  wire h_s_dadda_rca32_and_15_20_y0;
  wire h_s_dadda_rca32_and_14_21_y0;
  wire h_s_dadda_rca32_fa413_y2;
  wire h_s_dadda_rca32_fa413_y4;
  wire h_s_dadda_rca32_and_13_22_y0;
  wire h_s_dadda_rca32_and_12_23_y0;
  wire h_s_dadda_rca32_and_11_24_y0;
  wire h_s_dadda_rca32_fa414_y2;
  wire h_s_dadda_rca32_fa414_y4;
  wire h_s_dadda_rca32_and_10_25_y0;
  wire h_s_dadda_rca32_and_9_26_y0;
  wire h_s_dadda_rca32_and_8_27_y0;
  wire h_s_dadda_rca32_fa415_y2;
  wire h_s_dadda_rca32_fa415_y4;
  wire h_s_dadda_rca32_and_7_28_y0;
  wire h_s_dadda_rca32_and_6_29_y0;
  wire h_s_dadda_rca32_and_5_30_y0;
  wire h_s_dadda_rca32_fa416_y2;
  wire h_s_dadda_rca32_fa416_y4;
  wire h_s_dadda_rca32_nand_4_31_y0;
  wire h_s_dadda_rca32_fa417_y2;
  wire h_s_dadda_rca32_fa417_y4;
  wire h_s_dadda_rca32_fa418_y2;
  wire h_s_dadda_rca32_fa418_y4;
  wire h_s_dadda_rca32_fa419_y2;
  wire h_s_dadda_rca32_fa419_y4;
  wire h_s_dadda_rca32_fa420_y2;
  wire h_s_dadda_rca32_fa420_y4;
  wire h_s_dadda_rca32_fa421_y2;
  wire h_s_dadda_rca32_fa421_y4;
  wire h_s_dadda_rca32_fa422_y2;
  wire h_s_dadda_rca32_fa422_y4;
  wire h_s_dadda_rca32_fa423_y2;
  wire h_s_dadda_rca32_fa423_y4;
  wire h_s_dadda_rca32_fa424_y2;
  wire h_s_dadda_rca32_fa424_y4;
  wire h_s_dadda_rca32_fa425_y2;
  wire h_s_dadda_rca32_fa425_y4;
  wire h_s_dadda_rca32_fa426_y2;
  wire h_s_dadda_rca32_fa426_y4;
  wire h_s_dadda_rca32_fa427_y2;
  wire h_s_dadda_rca32_fa427_y4;
  wire h_s_dadda_rca32_fa428_y2;
  wire h_s_dadda_rca32_fa428_y4;
  wire h_s_dadda_rca32_fa429_y2;
  wire h_s_dadda_rca32_fa429_y4;
  wire h_s_dadda_rca32_nand_31_5_y0;
  wire h_s_dadda_rca32_fa430_y2;
  wire h_s_dadda_rca32_fa430_y4;
  wire h_s_dadda_rca32_and_30_6_y0;
  wire h_s_dadda_rca32_and_29_7_y0;
  wire h_s_dadda_rca32_and_28_8_y0;
  wire h_s_dadda_rca32_fa431_y2;
  wire h_s_dadda_rca32_fa431_y4;
  wire h_s_dadda_rca32_and_27_9_y0;
  wire h_s_dadda_rca32_and_26_10_y0;
  wire h_s_dadda_rca32_and_25_11_y0;
  wire h_s_dadda_rca32_fa432_y2;
  wire h_s_dadda_rca32_fa432_y4;
  wire h_s_dadda_rca32_and_24_12_y0;
  wire h_s_dadda_rca32_and_23_13_y0;
  wire h_s_dadda_rca32_and_22_14_y0;
  wire h_s_dadda_rca32_fa433_y2;
  wire h_s_dadda_rca32_fa433_y4;
  wire h_s_dadda_rca32_and_21_15_y0;
  wire h_s_dadda_rca32_and_20_16_y0;
  wire h_s_dadda_rca32_and_19_17_y0;
  wire h_s_dadda_rca32_fa434_y2;
  wire h_s_dadda_rca32_fa434_y4;
  wire h_s_dadda_rca32_and_18_18_y0;
  wire h_s_dadda_rca32_and_17_19_y0;
  wire h_s_dadda_rca32_and_16_20_y0;
  wire h_s_dadda_rca32_fa435_y2;
  wire h_s_dadda_rca32_fa435_y4;
  wire h_s_dadda_rca32_and_15_21_y0;
  wire h_s_dadda_rca32_and_14_22_y0;
  wire h_s_dadda_rca32_and_13_23_y0;
  wire h_s_dadda_rca32_fa436_y2;
  wire h_s_dadda_rca32_fa436_y4;
  wire h_s_dadda_rca32_and_12_24_y0;
  wire h_s_dadda_rca32_and_11_25_y0;
  wire h_s_dadda_rca32_and_10_26_y0;
  wire h_s_dadda_rca32_fa437_y2;
  wire h_s_dadda_rca32_fa437_y4;
  wire h_s_dadda_rca32_and_9_27_y0;
  wire h_s_dadda_rca32_and_8_28_y0;
  wire h_s_dadda_rca32_and_7_29_y0;
  wire h_s_dadda_rca32_fa438_y2;
  wire h_s_dadda_rca32_fa438_y4;
  wire h_s_dadda_rca32_and_6_30_y0;
  wire h_s_dadda_rca32_nand_5_31_y0;
  wire h_s_dadda_rca32_fa439_y2;
  wire h_s_dadda_rca32_fa439_y4;
  wire h_s_dadda_rca32_fa440_y2;
  wire h_s_dadda_rca32_fa440_y4;
  wire h_s_dadda_rca32_fa441_y2;
  wire h_s_dadda_rca32_fa441_y4;
  wire h_s_dadda_rca32_fa442_y2;
  wire h_s_dadda_rca32_fa442_y4;
  wire h_s_dadda_rca32_fa443_y2;
  wire h_s_dadda_rca32_fa443_y4;
  wire h_s_dadda_rca32_fa444_y2;
  wire h_s_dadda_rca32_fa444_y4;
  wire h_s_dadda_rca32_fa445_y2;
  wire h_s_dadda_rca32_fa445_y4;
  wire h_s_dadda_rca32_fa446_y2;
  wire h_s_dadda_rca32_fa446_y4;
  wire h_s_dadda_rca32_fa447_y2;
  wire h_s_dadda_rca32_fa447_y4;
  wire h_s_dadda_rca32_fa448_y2;
  wire h_s_dadda_rca32_fa448_y4;
  wire h_s_dadda_rca32_fa449_y2;
  wire h_s_dadda_rca32_fa449_y4;
  wire h_s_dadda_rca32_fa450_y2;
  wire h_s_dadda_rca32_fa450_y4;
  wire h_s_dadda_rca32_fa451_y2;
  wire h_s_dadda_rca32_fa451_y4;
  wire h_s_dadda_rca32_nand_31_6_y0;
  wire h_s_dadda_rca32_and_30_7_y0;
  wire h_s_dadda_rca32_fa452_y2;
  wire h_s_dadda_rca32_fa452_y4;
  wire h_s_dadda_rca32_and_29_8_y0;
  wire h_s_dadda_rca32_and_28_9_y0;
  wire h_s_dadda_rca32_and_27_10_y0;
  wire h_s_dadda_rca32_fa453_y2;
  wire h_s_dadda_rca32_fa453_y4;
  wire h_s_dadda_rca32_and_26_11_y0;
  wire h_s_dadda_rca32_and_25_12_y0;
  wire h_s_dadda_rca32_and_24_13_y0;
  wire h_s_dadda_rca32_fa454_y2;
  wire h_s_dadda_rca32_fa454_y4;
  wire h_s_dadda_rca32_and_23_14_y0;
  wire h_s_dadda_rca32_and_22_15_y0;
  wire h_s_dadda_rca32_and_21_16_y0;
  wire h_s_dadda_rca32_fa455_y2;
  wire h_s_dadda_rca32_fa455_y4;
  wire h_s_dadda_rca32_and_20_17_y0;
  wire h_s_dadda_rca32_and_19_18_y0;
  wire h_s_dadda_rca32_and_18_19_y0;
  wire h_s_dadda_rca32_fa456_y2;
  wire h_s_dadda_rca32_fa456_y4;
  wire h_s_dadda_rca32_and_17_20_y0;
  wire h_s_dadda_rca32_and_16_21_y0;
  wire h_s_dadda_rca32_and_15_22_y0;
  wire h_s_dadda_rca32_fa457_y2;
  wire h_s_dadda_rca32_fa457_y4;
  wire h_s_dadda_rca32_and_14_23_y0;
  wire h_s_dadda_rca32_and_13_24_y0;
  wire h_s_dadda_rca32_and_12_25_y0;
  wire h_s_dadda_rca32_fa458_y2;
  wire h_s_dadda_rca32_fa458_y4;
  wire h_s_dadda_rca32_and_11_26_y0;
  wire h_s_dadda_rca32_and_10_27_y0;
  wire h_s_dadda_rca32_and_9_28_y0;
  wire h_s_dadda_rca32_fa459_y2;
  wire h_s_dadda_rca32_fa459_y4;
  wire h_s_dadda_rca32_and_8_29_y0;
  wire h_s_dadda_rca32_and_7_30_y0;
  wire h_s_dadda_rca32_nand_6_31_y0;
  wire h_s_dadda_rca32_fa460_y2;
  wire h_s_dadda_rca32_fa460_y4;
  wire h_s_dadda_rca32_fa461_y2;
  wire h_s_dadda_rca32_fa461_y4;
  wire h_s_dadda_rca32_fa462_y2;
  wire h_s_dadda_rca32_fa462_y4;
  wire h_s_dadda_rca32_fa463_y2;
  wire h_s_dadda_rca32_fa463_y4;
  wire h_s_dadda_rca32_fa464_y2;
  wire h_s_dadda_rca32_fa464_y4;
  wire h_s_dadda_rca32_fa465_y2;
  wire h_s_dadda_rca32_fa465_y4;
  wire h_s_dadda_rca32_fa466_y2;
  wire h_s_dadda_rca32_fa466_y4;
  wire h_s_dadda_rca32_fa467_y2;
  wire h_s_dadda_rca32_fa467_y4;
  wire h_s_dadda_rca32_fa468_y2;
  wire h_s_dadda_rca32_fa468_y4;
  wire h_s_dadda_rca32_fa469_y2;
  wire h_s_dadda_rca32_fa469_y4;
  wire h_s_dadda_rca32_fa470_y2;
  wire h_s_dadda_rca32_fa470_y4;
  wire h_s_dadda_rca32_fa471_y2;
  wire h_s_dadda_rca32_fa471_y4;
  wire h_s_dadda_rca32_fa472_y2;
  wire h_s_dadda_rca32_fa472_y4;
  wire h_s_dadda_rca32_nand_31_7_y0;
  wire h_s_dadda_rca32_and_30_8_y0;
  wire h_s_dadda_rca32_and_29_9_y0;
  wire h_s_dadda_rca32_fa473_y2;
  wire h_s_dadda_rca32_fa473_y4;
  wire h_s_dadda_rca32_and_28_10_y0;
  wire h_s_dadda_rca32_and_27_11_y0;
  wire h_s_dadda_rca32_and_26_12_y0;
  wire h_s_dadda_rca32_fa474_y2;
  wire h_s_dadda_rca32_fa474_y4;
  wire h_s_dadda_rca32_and_25_13_y0;
  wire h_s_dadda_rca32_and_24_14_y0;
  wire h_s_dadda_rca32_and_23_15_y0;
  wire h_s_dadda_rca32_fa475_y2;
  wire h_s_dadda_rca32_fa475_y4;
  wire h_s_dadda_rca32_and_22_16_y0;
  wire h_s_dadda_rca32_and_21_17_y0;
  wire h_s_dadda_rca32_and_20_18_y0;
  wire h_s_dadda_rca32_fa476_y2;
  wire h_s_dadda_rca32_fa476_y4;
  wire h_s_dadda_rca32_and_19_19_y0;
  wire h_s_dadda_rca32_and_18_20_y0;
  wire h_s_dadda_rca32_and_17_21_y0;
  wire h_s_dadda_rca32_fa477_y2;
  wire h_s_dadda_rca32_fa477_y4;
  wire h_s_dadda_rca32_and_16_22_y0;
  wire h_s_dadda_rca32_and_15_23_y0;
  wire h_s_dadda_rca32_and_14_24_y0;
  wire h_s_dadda_rca32_fa478_y2;
  wire h_s_dadda_rca32_fa478_y4;
  wire h_s_dadda_rca32_and_13_25_y0;
  wire h_s_dadda_rca32_and_12_26_y0;
  wire h_s_dadda_rca32_and_11_27_y0;
  wire h_s_dadda_rca32_fa479_y2;
  wire h_s_dadda_rca32_fa479_y4;
  wire h_s_dadda_rca32_and_10_28_y0;
  wire h_s_dadda_rca32_and_9_29_y0;
  wire h_s_dadda_rca32_and_8_30_y0;
  wire h_s_dadda_rca32_fa480_y2;
  wire h_s_dadda_rca32_fa480_y4;
  wire h_s_dadda_rca32_nand_7_31_y0;
  wire h_s_dadda_rca32_fa481_y2;
  wire h_s_dadda_rca32_fa481_y4;
  wire h_s_dadda_rca32_fa482_y2;
  wire h_s_dadda_rca32_fa482_y4;
  wire h_s_dadda_rca32_fa483_y2;
  wire h_s_dadda_rca32_fa483_y4;
  wire h_s_dadda_rca32_fa484_y2;
  wire h_s_dadda_rca32_fa484_y4;
  wire h_s_dadda_rca32_fa485_y2;
  wire h_s_dadda_rca32_fa485_y4;
  wire h_s_dadda_rca32_fa486_y2;
  wire h_s_dadda_rca32_fa486_y4;
  wire h_s_dadda_rca32_fa487_y2;
  wire h_s_dadda_rca32_fa487_y4;
  wire h_s_dadda_rca32_fa488_y2;
  wire h_s_dadda_rca32_fa488_y4;
  wire h_s_dadda_rca32_fa489_y2;
  wire h_s_dadda_rca32_fa489_y4;
  wire h_s_dadda_rca32_fa490_y2;
  wire h_s_dadda_rca32_fa490_y4;
  wire h_s_dadda_rca32_fa491_y2;
  wire h_s_dadda_rca32_fa491_y4;
  wire h_s_dadda_rca32_nand_31_8_y0;
  wire h_s_dadda_rca32_fa492_y2;
  wire h_s_dadda_rca32_fa492_y4;
  wire h_s_dadda_rca32_and_30_9_y0;
  wire h_s_dadda_rca32_and_29_10_y0;
  wire h_s_dadda_rca32_and_28_11_y0;
  wire h_s_dadda_rca32_fa493_y2;
  wire h_s_dadda_rca32_fa493_y4;
  wire h_s_dadda_rca32_and_27_12_y0;
  wire h_s_dadda_rca32_and_26_13_y0;
  wire h_s_dadda_rca32_and_25_14_y0;
  wire h_s_dadda_rca32_fa494_y2;
  wire h_s_dadda_rca32_fa494_y4;
  wire h_s_dadda_rca32_and_24_15_y0;
  wire h_s_dadda_rca32_and_23_16_y0;
  wire h_s_dadda_rca32_and_22_17_y0;
  wire h_s_dadda_rca32_fa495_y2;
  wire h_s_dadda_rca32_fa495_y4;
  wire h_s_dadda_rca32_and_21_18_y0;
  wire h_s_dadda_rca32_and_20_19_y0;
  wire h_s_dadda_rca32_and_19_20_y0;
  wire h_s_dadda_rca32_fa496_y2;
  wire h_s_dadda_rca32_fa496_y4;
  wire h_s_dadda_rca32_and_18_21_y0;
  wire h_s_dadda_rca32_and_17_22_y0;
  wire h_s_dadda_rca32_and_16_23_y0;
  wire h_s_dadda_rca32_fa497_y2;
  wire h_s_dadda_rca32_fa497_y4;
  wire h_s_dadda_rca32_and_15_24_y0;
  wire h_s_dadda_rca32_and_14_25_y0;
  wire h_s_dadda_rca32_and_13_26_y0;
  wire h_s_dadda_rca32_fa498_y2;
  wire h_s_dadda_rca32_fa498_y4;
  wire h_s_dadda_rca32_and_12_27_y0;
  wire h_s_dadda_rca32_and_11_28_y0;
  wire h_s_dadda_rca32_and_10_29_y0;
  wire h_s_dadda_rca32_fa499_y2;
  wire h_s_dadda_rca32_fa499_y4;
  wire h_s_dadda_rca32_and_9_30_y0;
  wire h_s_dadda_rca32_nand_8_31_y0;
  wire h_s_dadda_rca32_fa500_y2;
  wire h_s_dadda_rca32_fa500_y4;
  wire h_s_dadda_rca32_fa501_y2;
  wire h_s_dadda_rca32_fa501_y4;
  wire h_s_dadda_rca32_fa502_y2;
  wire h_s_dadda_rca32_fa502_y4;
  wire h_s_dadda_rca32_fa503_y2;
  wire h_s_dadda_rca32_fa503_y4;
  wire h_s_dadda_rca32_fa504_y2;
  wire h_s_dadda_rca32_fa504_y4;
  wire h_s_dadda_rca32_fa505_y2;
  wire h_s_dadda_rca32_fa505_y4;
  wire h_s_dadda_rca32_fa506_y2;
  wire h_s_dadda_rca32_fa506_y4;
  wire h_s_dadda_rca32_fa507_y2;
  wire h_s_dadda_rca32_fa507_y4;
  wire h_s_dadda_rca32_fa508_y2;
  wire h_s_dadda_rca32_fa508_y4;
  wire h_s_dadda_rca32_fa509_y2;
  wire h_s_dadda_rca32_fa509_y4;
  wire h_s_dadda_rca32_fa510_y2;
  wire h_s_dadda_rca32_fa510_y4;
  wire h_s_dadda_rca32_nand_31_9_y0;
  wire h_s_dadda_rca32_and_30_10_y0;
  wire h_s_dadda_rca32_fa511_y2;
  wire h_s_dadda_rca32_fa511_y4;
  wire h_s_dadda_rca32_and_29_11_y0;
  wire h_s_dadda_rca32_and_28_12_y0;
  wire h_s_dadda_rca32_and_27_13_y0;
  wire h_s_dadda_rca32_fa512_y2;
  wire h_s_dadda_rca32_fa512_y4;
  wire h_s_dadda_rca32_and_26_14_y0;
  wire h_s_dadda_rca32_and_25_15_y0;
  wire h_s_dadda_rca32_and_24_16_y0;
  wire h_s_dadda_rca32_fa513_y2;
  wire h_s_dadda_rca32_fa513_y4;
  wire h_s_dadda_rca32_and_23_17_y0;
  wire h_s_dadda_rca32_and_22_18_y0;
  wire h_s_dadda_rca32_and_21_19_y0;
  wire h_s_dadda_rca32_fa514_y2;
  wire h_s_dadda_rca32_fa514_y4;
  wire h_s_dadda_rca32_and_20_20_y0;
  wire h_s_dadda_rca32_and_19_21_y0;
  wire h_s_dadda_rca32_and_18_22_y0;
  wire h_s_dadda_rca32_fa515_y2;
  wire h_s_dadda_rca32_fa515_y4;
  wire h_s_dadda_rca32_and_17_23_y0;
  wire h_s_dadda_rca32_and_16_24_y0;
  wire h_s_dadda_rca32_and_15_25_y0;
  wire h_s_dadda_rca32_fa516_y2;
  wire h_s_dadda_rca32_fa516_y4;
  wire h_s_dadda_rca32_and_14_26_y0;
  wire h_s_dadda_rca32_and_13_27_y0;
  wire h_s_dadda_rca32_and_12_28_y0;
  wire h_s_dadda_rca32_fa517_y2;
  wire h_s_dadda_rca32_fa517_y4;
  wire h_s_dadda_rca32_and_11_29_y0;
  wire h_s_dadda_rca32_and_10_30_y0;
  wire h_s_dadda_rca32_nand_9_31_y0;
  wire h_s_dadda_rca32_fa518_y2;
  wire h_s_dadda_rca32_fa518_y4;
  wire h_s_dadda_rca32_fa519_y2;
  wire h_s_dadda_rca32_fa519_y4;
  wire h_s_dadda_rca32_fa520_y2;
  wire h_s_dadda_rca32_fa520_y4;
  wire h_s_dadda_rca32_fa521_y2;
  wire h_s_dadda_rca32_fa521_y4;
  wire h_s_dadda_rca32_fa522_y2;
  wire h_s_dadda_rca32_fa522_y4;
  wire h_s_dadda_rca32_fa523_y2;
  wire h_s_dadda_rca32_fa523_y4;
  wire h_s_dadda_rca32_fa524_y2;
  wire h_s_dadda_rca32_fa524_y4;
  wire h_s_dadda_rca32_fa525_y2;
  wire h_s_dadda_rca32_fa525_y4;
  wire h_s_dadda_rca32_fa526_y2;
  wire h_s_dadda_rca32_fa526_y4;
  wire h_s_dadda_rca32_fa527_y2;
  wire h_s_dadda_rca32_fa527_y4;
  wire h_s_dadda_rca32_fa528_y2;
  wire h_s_dadda_rca32_fa528_y4;
  wire h_s_dadda_rca32_nand_31_10_y0;
  wire h_s_dadda_rca32_and_30_11_y0;
  wire h_s_dadda_rca32_and_29_12_y0;
  wire h_s_dadda_rca32_fa529_y2;
  wire h_s_dadda_rca32_fa529_y4;
  wire h_s_dadda_rca32_and_28_13_y0;
  wire h_s_dadda_rca32_and_27_14_y0;
  wire h_s_dadda_rca32_and_26_15_y0;
  wire h_s_dadda_rca32_fa530_y2;
  wire h_s_dadda_rca32_fa530_y4;
  wire h_s_dadda_rca32_and_25_16_y0;
  wire h_s_dadda_rca32_and_24_17_y0;
  wire h_s_dadda_rca32_and_23_18_y0;
  wire h_s_dadda_rca32_fa531_y2;
  wire h_s_dadda_rca32_fa531_y4;
  wire h_s_dadda_rca32_and_22_19_y0;
  wire h_s_dadda_rca32_and_21_20_y0;
  wire h_s_dadda_rca32_and_20_21_y0;
  wire h_s_dadda_rca32_fa532_y2;
  wire h_s_dadda_rca32_fa532_y4;
  wire h_s_dadda_rca32_and_19_22_y0;
  wire h_s_dadda_rca32_and_18_23_y0;
  wire h_s_dadda_rca32_and_17_24_y0;
  wire h_s_dadda_rca32_fa533_y2;
  wire h_s_dadda_rca32_fa533_y4;
  wire h_s_dadda_rca32_and_16_25_y0;
  wire h_s_dadda_rca32_and_15_26_y0;
  wire h_s_dadda_rca32_and_14_27_y0;
  wire h_s_dadda_rca32_fa534_y2;
  wire h_s_dadda_rca32_fa534_y4;
  wire h_s_dadda_rca32_and_13_28_y0;
  wire h_s_dadda_rca32_and_12_29_y0;
  wire h_s_dadda_rca32_and_11_30_y0;
  wire h_s_dadda_rca32_fa535_y2;
  wire h_s_dadda_rca32_fa535_y4;
  wire h_s_dadda_rca32_nand_10_31_y0;
  wire h_s_dadda_rca32_fa536_y2;
  wire h_s_dadda_rca32_fa536_y4;
  wire h_s_dadda_rca32_fa537_y2;
  wire h_s_dadda_rca32_fa537_y4;
  wire h_s_dadda_rca32_fa538_y2;
  wire h_s_dadda_rca32_fa538_y4;
  wire h_s_dadda_rca32_fa539_y2;
  wire h_s_dadda_rca32_fa539_y4;
  wire h_s_dadda_rca32_fa540_y2;
  wire h_s_dadda_rca32_fa540_y4;
  wire h_s_dadda_rca32_fa541_y2;
  wire h_s_dadda_rca32_fa541_y4;
  wire h_s_dadda_rca32_fa542_y2;
  wire h_s_dadda_rca32_fa542_y4;
  wire h_s_dadda_rca32_fa543_y2;
  wire h_s_dadda_rca32_fa543_y4;
  wire h_s_dadda_rca32_fa544_y2;
  wire h_s_dadda_rca32_fa544_y4;
  wire h_s_dadda_rca32_nand_31_11_y0;
  wire h_s_dadda_rca32_fa545_y2;
  wire h_s_dadda_rca32_fa545_y4;
  wire h_s_dadda_rca32_and_30_12_y0;
  wire h_s_dadda_rca32_and_29_13_y0;
  wire h_s_dadda_rca32_and_28_14_y0;
  wire h_s_dadda_rca32_fa546_y2;
  wire h_s_dadda_rca32_fa546_y4;
  wire h_s_dadda_rca32_and_27_15_y0;
  wire h_s_dadda_rca32_and_26_16_y0;
  wire h_s_dadda_rca32_and_25_17_y0;
  wire h_s_dadda_rca32_fa547_y2;
  wire h_s_dadda_rca32_fa547_y4;
  wire h_s_dadda_rca32_and_24_18_y0;
  wire h_s_dadda_rca32_and_23_19_y0;
  wire h_s_dadda_rca32_and_22_20_y0;
  wire h_s_dadda_rca32_fa548_y2;
  wire h_s_dadda_rca32_fa548_y4;
  wire h_s_dadda_rca32_and_21_21_y0;
  wire h_s_dadda_rca32_and_20_22_y0;
  wire h_s_dadda_rca32_and_19_23_y0;
  wire h_s_dadda_rca32_fa549_y2;
  wire h_s_dadda_rca32_fa549_y4;
  wire h_s_dadda_rca32_and_18_24_y0;
  wire h_s_dadda_rca32_and_17_25_y0;
  wire h_s_dadda_rca32_and_16_26_y0;
  wire h_s_dadda_rca32_fa550_y2;
  wire h_s_dadda_rca32_fa550_y4;
  wire h_s_dadda_rca32_and_15_27_y0;
  wire h_s_dadda_rca32_and_14_28_y0;
  wire h_s_dadda_rca32_and_13_29_y0;
  wire h_s_dadda_rca32_fa551_y2;
  wire h_s_dadda_rca32_fa551_y4;
  wire h_s_dadda_rca32_and_12_30_y0;
  wire h_s_dadda_rca32_nand_11_31_y0;
  wire h_s_dadda_rca32_fa552_y2;
  wire h_s_dadda_rca32_fa552_y4;
  wire h_s_dadda_rca32_fa553_y2;
  wire h_s_dadda_rca32_fa553_y4;
  wire h_s_dadda_rca32_fa554_y2;
  wire h_s_dadda_rca32_fa554_y4;
  wire h_s_dadda_rca32_fa555_y2;
  wire h_s_dadda_rca32_fa555_y4;
  wire h_s_dadda_rca32_fa556_y2;
  wire h_s_dadda_rca32_fa556_y4;
  wire h_s_dadda_rca32_fa557_y2;
  wire h_s_dadda_rca32_fa557_y4;
  wire h_s_dadda_rca32_fa558_y2;
  wire h_s_dadda_rca32_fa558_y4;
  wire h_s_dadda_rca32_fa559_y2;
  wire h_s_dadda_rca32_fa559_y4;
  wire h_s_dadda_rca32_fa560_y2;
  wire h_s_dadda_rca32_fa560_y4;
  wire h_s_dadda_rca32_nand_31_12_y0;
  wire h_s_dadda_rca32_and_30_13_y0;
  wire h_s_dadda_rca32_fa561_y2;
  wire h_s_dadda_rca32_fa561_y4;
  wire h_s_dadda_rca32_and_29_14_y0;
  wire h_s_dadda_rca32_and_28_15_y0;
  wire h_s_dadda_rca32_and_27_16_y0;
  wire h_s_dadda_rca32_fa562_y2;
  wire h_s_dadda_rca32_fa562_y4;
  wire h_s_dadda_rca32_and_26_17_y0;
  wire h_s_dadda_rca32_and_25_18_y0;
  wire h_s_dadda_rca32_and_24_19_y0;
  wire h_s_dadda_rca32_fa563_y2;
  wire h_s_dadda_rca32_fa563_y4;
  wire h_s_dadda_rca32_and_23_20_y0;
  wire h_s_dadda_rca32_and_22_21_y0;
  wire h_s_dadda_rca32_and_21_22_y0;
  wire h_s_dadda_rca32_fa564_y2;
  wire h_s_dadda_rca32_fa564_y4;
  wire h_s_dadda_rca32_and_20_23_y0;
  wire h_s_dadda_rca32_and_19_24_y0;
  wire h_s_dadda_rca32_and_18_25_y0;
  wire h_s_dadda_rca32_fa565_y2;
  wire h_s_dadda_rca32_fa565_y4;
  wire h_s_dadda_rca32_and_17_26_y0;
  wire h_s_dadda_rca32_and_16_27_y0;
  wire h_s_dadda_rca32_and_15_28_y0;
  wire h_s_dadda_rca32_fa566_y2;
  wire h_s_dadda_rca32_fa566_y4;
  wire h_s_dadda_rca32_and_14_29_y0;
  wire h_s_dadda_rca32_and_13_30_y0;
  wire h_s_dadda_rca32_nand_12_31_y0;
  wire h_s_dadda_rca32_fa567_y2;
  wire h_s_dadda_rca32_fa567_y4;
  wire h_s_dadda_rca32_fa568_y2;
  wire h_s_dadda_rca32_fa568_y4;
  wire h_s_dadda_rca32_fa569_y2;
  wire h_s_dadda_rca32_fa569_y4;
  wire h_s_dadda_rca32_fa570_y2;
  wire h_s_dadda_rca32_fa570_y4;
  wire h_s_dadda_rca32_fa571_y2;
  wire h_s_dadda_rca32_fa571_y4;
  wire h_s_dadda_rca32_fa572_y2;
  wire h_s_dadda_rca32_fa572_y4;
  wire h_s_dadda_rca32_fa573_y2;
  wire h_s_dadda_rca32_fa573_y4;
  wire h_s_dadda_rca32_fa574_y2;
  wire h_s_dadda_rca32_fa574_y4;
  wire h_s_dadda_rca32_fa575_y2;
  wire h_s_dadda_rca32_fa575_y4;
  wire h_s_dadda_rca32_nand_31_13_y0;
  wire h_s_dadda_rca32_and_30_14_y0;
  wire h_s_dadda_rca32_and_29_15_y0;
  wire h_s_dadda_rca32_fa576_y2;
  wire h_s_dadda_rca32_fa576_y4;
  wire h_s_dadda_rca32_and_28_16_y0;
  wire h_s_dadda_rca32_and_27_17_y0;
  wire h_s_dadda_rca32_and_26_18_y0;
  wire h_s_dadda_rca32_fa577_y2;
  wire h_s_dadda_rca32_fa577_y4;
  wire h_s_dadda_rca32_and_25_19_y0;
  wire h_s_dadda_rca32_and_24_20_y0;
  wire h_s_dadda_rca32_and_23_21_y0;
  wire h_s_dadda_rca32_fa578_y2;
  wire h_s_dadda_rca32_fa578_y4;
  wire h_s_dadda_rca32_and_22_22_y0;
  wire h_s_dadda_rca32_and_21_23_y0;
  wire h_s_dadda_rca32_and_20_24_y0;
  wire h_s_dadda_rca32_fa579_y2;
  wire h_s_dadda_rca32_fa579_y4;
  wire h_s_dadda_rca32_and_19_25_y0;
  wire h_s_dadda_rca32_and_18_26_y0;
  wire h_s_dadda_rca32_and_17_27_y0;
  wire h_s_dadda_rca32_fa580_y2;
  wire h_s_dadda_rca32_fa580_y4;
  wire h_s_dadda_rca32_and_16_28_y0;
  wire h_s_dadda_rca32_and_15_29_y0;
  wire h_s_dadda_rca32_and_14_30_y0;
  wire h_s_dadda_rca32_fa581_y2;
  wire h_s_dadda_rca32_fa581_y4;
  wire h_s_dadda_rca32_nand_13_31_y0;
  wire h_s_dadda_rca32_fa582_y2;
  wire h_s_dadda_rca32_fa582_y4;
  wire h_s_dadda_rca32_fa583_y2;
  wire h_s_dadda_rca32_fa583_y4;
  wire h_s_dadda_rca32_fa584_y2;
  wire h_s_dadda_rca32_fa584_y4;
  wire h_s_dadda_rca32_fa585_y2;
  wire h_s_dadda_rca32_fa585_y4;
  wire h_s_dadda_rca32_fa586_y2;
  wire h_s_dadda_rca32_fa586_y4;
  wire h_s_dadda_rca32_fa587_y2;
  wire h_s_dadda_rca32_fa587_y4;
  wire h_s_dadda_rca32_fa588_y2;
  wire h_s_dadda_rca32_fa588_y4;
  wire h_s_dadda_rca32_nand_31_14_y0;
  wire h_s_dadda_rca32_fa589_y2;
  wire h_s_dadda_rca32_fa589_y4;
  wire h_s_dadda_rca32_and_30_15_y0;
  wire h_s_dadda_rca32_and_29_16_y0;
  wire h_s_dadda_rca32_and_28_17_y0;
  wire h_s_dadda_rca32_fa590_y2;
  wire h_s_dadda_rca32_fa590_y4;
  wire h_s_dadda_rca32_and_27_18_y0;
  wire h_s_dadda_rca32_and_26_19_y0;
  wire h_s_dadda_rca32_and_25_20_y0;
  wire h_s_dadda_rca32_fa591_y2;
  wire h_s_dadda_rca32_fa591_y4;
  wire h_s_dadda_rca32_and_24_21_y0;
  wire h_s_dadda_rca32_and_23_22_y0;
  wire h_s_dadda_rca32_and_22_23_y0;
  wire h_s_dadda_rca32_fa592_y2;
  wire h_s_dadda_rca32_fa592_y4;
  wire h_s_dadda_rca32_and_21_24_y0;
  wire h_s_dadda_rca32_and_20_25_y0;
  wire h_s_dadda_rca32_and_19_26_y0;
  wire h_s_dadda_rca32_fa593_y2;
  wire h_s_dadda_rca32_fa593_y4;
  wire h_s_dadda_rca32_and_18_27_y0;
  wire h_s_dadda_rca32_and_17_28_y0;
  wire h_s_dadda_rca32_and_16_29_y0;
  wire h_s_dadda_rca32_fa594_y2;
  wire h_s_dadda_rca32_fa594_y4;
  wire h_s_dadda_rca32_and_15_30_y0;
  wire h_s_dadda_rca32_nand_14_31_y0;
  wire h_s_dadda_rca32_fa595_y2;
  wire h_s_dadda_rca32_fa595_y4;
  wire h_s_dadda_rca32_fa596_y2;
  wire h_s_dadda_rca32_fa596_y4;
  wire h_s_dadda_rca32_fa597_y2;
  wire h_s_dadda_rca32_fa597_y4;
  wire h_s_dadda_rca32_fa598_y2;
  wire h_s_dadda_rca32_fa598_y4;
  wire h_s_dadda_rca32_fa599_y2;
  wire h_s_dadda_rca32_fa599_y4;
  wire h_s_dadda_rca32_fa600_y2;
  wire h_s_dadda_rca32_fa600_y4;
  wire h_s_dadda_rca32_fa601_y2;
  wire h_s_dadda_rca32_fa601_y4;
  wire h_s_dadda_rca32_nand_31_15_y0;
  wire h_s_dadda_rca32_and_30_16_y0;
  wire h_s_dadda_rca32_fa602_y2;
  wire h_s_dadda_rca32_fa602_y4;
  wire h_s_dadda_rca32_and_29_17_y0;
  wire h_s_dadda_rca32_and_28_18_y0;
  wire h_s_dadda_rca32_and_27_19_y0;
  wire h_s_dadda_rca32_fa603_y2;
  wire h_s_dadda_rca32_fa603_y4;
  wire h_s_dadda_rca32_and_26_20_y0;
  wire h_s_dadda_rca32_and_25_21_y0;
  wire h_s_dadda_rca32_and_24_22_y0;
  wire h_s_dadda_rca32_fa604_y2;
  wire h_s_dadda_rca32_fa604_y4;
  wire h_s_dadda_rca32_and_23_23_y0;
  wire h_s_dadda_rca32_and_22_24_y0;
  wire h_s_dadda_rca32_and_21_25_y0;
  wire h_s_dadda_rca32_fa605_y2;
  wire h_s_dadda_rca32_fa605_y4;
  wire h_s_dadda_rca32_and_20_26_y0;
  wire h_s_dadda_rca32_and_19_27_y0;
  wire h_s_dadda_rca32_and_18_28_y0;
  wire h_s_dadda_rca32_fa606_y2;
  wire h_s_dadda_rca32_fa606_y4;
  wire h_s_dadda_rca32_and_17_29_y0;
  wire h_s_dadda_rca32_and_16_30_y0;
  wire h_s_dadda_rca32_nand_15_31_y0;
  wire h_s_dadda_rca32_fa607_y2;
  wire h_s_dadda_rca32_fa607_y4;
  wire h_s_dadda_rca32_fa608_y2;
  wire h_s_dadda_rca32_fa608_y4;
  wire h_s_dadda_rca32_fa609_y2;
  wire h_s_dadda_rca32_fa609_y4;
  wire h_s_dadda_rca32_fa610_y2;
  wire h_s_dadda_rca32_fa610_y4;
  wire h_s_dadda_rca32_fa611_y2;
  wire h_s_dadda_rca32_fa611_y4;
  wire h_s_dadda_rca32_fa612_y2;
  wire h_s_dadda_rca32_fa612_y4;
  wire h_s_dadda_rca32_fa613_y2;
  wire h_s_dadda_rca32_fa613_y4;
  wire h_s_dadda_rca32_nand_31_16_y0;
  wire h_s_dadda_rca32_and_30_17_y0;
  wire h_s_dadda_rca32_and_29_18_y0;
  wire h_s_dadda_rca32_fa614_y2;
  wire h_s_dadda_rca32_fa614_y4;
  wire h_s_dadda_rca32_and_28_19_y0;
  wire h_s_dadda_rca32_and_27_20_y0;
  wire h_s_dadda_rca32_and_26_21_y0;
  wire h_s_dadda_rca32_fa615_y2;
  wire h_s_dadda_rca32_fa615_y4;
  wire h_s_dadda_rca32_and_25_22_y0;
  wire h_s_dadda_rca32_and_24_23_y0;
  wire h_s_dadda_rca32_and_23_24_y0;
  wire h_s_dadda_rca32_fa616_y2;
  wire h_s_dadda_rca32_fa616_y4;
  wire h_s_dadda_rca32_and_22_25_y0;
  wire h_s_dadda_rca32_and_21_26_y0;
  wire h_s_dadda_rca32_and_20_27_y0;
  wire h_s_dadda_rca32_fa617_y2;
  wire h_s_dadda_rca32_fa617_y4;
  wire h_s_dadda_rca32_and_19_28_y0;
  wire h_s_dadda_rca32_and_18_29_y0;
  wire h_s_dadda_rca32_and_17_30_y0;
  wire h_s_dadda_rca32_fa618_y2;
  wire h_s_dadda_rca32_fa618_y4;
  wire h_s_dadda_rca32_nand_16_31_y0;
  wire h_s_dadda_rca32_fa619_y2;
  wire h_s_dadda_rca32_fa619_y4;
  wire h_s_dadda_rca32_fa620_y2;
  wire h_s_dadda_rca32_fa620_y4;
  wire h_s_dadda_rca32_fa621_y2;
  wire h_s_dadda_rca32_fa621_y4;
  wire h_s_dadda_rca32_fa622_y2;
  wire h_s_dadda_rca32_fa622_y4;
  wire h_s_dadda_rca32_fa623_y2;
  wire h_s_dadda_rca32_fa623_y4;
  wire h_s_dadda_rca32_nand_31_17_y0;
  wire h_s_dadda_rca32_fa624_y2;
  wire h_s_dadda_rca32_fa624_y4;
  wire h_s_dadda_rca32_and_30_18_y0;
  wire h_s_dadda_rca32_and_29_19_y0;
  wire h_s_dadda_rca32_and_28_20_y0;
  wire h_s_dadda_rca32_fa625_y2;
  wire h_s_dadda_rca32_fa625_y4;
  wire h_s_dadda_rca32_and_27_21_y0;
  wire h_s_dadda_rca32_and_26_22_y0;
  wire h_s_dadda_rca32_and_25_23_y0;
  wire h_s_dadda_rca32_fa626_y2;
  wire h_s_dadda_rca32_fa626_y4;
  wire h_s_dadda_rca32_and_24_24_y0;
  wire h_s_dadda_rca32_and_23_25_y0;
  wire h_s_dadda_rca32_and_22_26_y0;
  wire h_s_dadda_rca32_fa627_y2;
  wire h_s_dadda_rca32_fa627_y4;
  wire h_s_dadda_rca32_and_21_27_y0;
  wire h_s_dadda_rca32_and_20_28_y0;
  wire h_s_dadda_rca32_and_19_29_y0;
  wire h_s_dadda_rca32_fa628_y2;
  wire h_s_dadda_rca32_fa628_y4;
  wire h_s_dadda_rca32_and_18_30_y0;
  wire h_s_dadda_rca32_nand_17_31_y0;
  wire h_s_dadda_rca32_fa629_y2;
  wire h_s_dadda_rca32_fa629_y4;
  wire h_s_dadda_rca32_fa630_y2;
  wire h_s_dadda_rca32_fa630_y4;
  wire h_s_dadda_rca32_fa631_y2;
  wire h_s_dadda_rca32_fa631_y4;
  wire h_s_dadda_rca32_fa632_y2;
  wire h_s_dadda_rca32_fa632_y4;
  wire h_s_dadda_rca32_fa633_y2;
  wire h_s_dadda_rca32_fa633_y4;
  wire h_s_dadda_rca32_nand_31_18_y0;
  wire h_s_dadda_rca32_and_30_19_y0;
  wire h_s_dadda_rca32_fa634_y2;
  wire h_s_dadda_rca32_fa634_y4;
  wire h_s_dadda_rca32_and_29_20_y0;
  wire h_s_dadda_rca32_and_28_21_y0;
  wire h_s_dadda_rca32_and_27_22_y0;
  wire h_s_dadda_rca32_fa635_y2;
  wire h_s_dadda_rca32_fa635_y4;
  wire h_s_dadda_rca32_and_26_23_y0;
  wire h_s_dadda_rca32_and_25_24_y0;
  wire h_s_dadda_rca32_and_24_25_y0;
  wire h_s_dadda_rca32_fa636_y2;
  wire h_s_dadda_rca32_fa636_y4;
  wire h_s_dadda_rca32_and_23_26_y0;
  wire h_s_dadda_rca32_and_22_27_y0;
  wire h_s_dadda_rca32_and_21_28_y0;
  wire h_s_dadda_rca32_fa637_y2;
  wire h_s_dadda_rca32_fa637_y4;
  wire h_s_dadda_rca32_and_20_29_y0;
  wire h_s_dadda_rca32_and_19_30_y0;
  wire h_s_dadda_rca32_nand_18_31_y0;
  wire h_s_dadda_rca32_fa638_y2;
  wire h_s_dadda_rca32_fa638_y4;
  wire h_s_dadda_rca32_fa639_y2;
  wire h_s_dadda_rca32_fa639_y4;
  wire h_s_dadda_rca32_fa640_y2;
  wire h_s_dadda_rca32_fa640_y4;
  wire h_s_dadda_rca32_fa641_y2;
  wire h_s_dadda_rca32_fa641_y4;
  wire h_s_dadda_rca32_fa642_y2;
  wire h_s_dadda_rca32_fa642_y4;
  wire h_s_dadda_rca32_nand_31_19_y0;
  wire h_s_dadda_rca32_and_30_20_y0;
  wire h_s_dadda_rca32_and_29_21_y0;
  wire h_s_dadda_rca32_fa643_y2;
  wire h_s_dadda_rca32_fa643_y4;
  wire h_s_dadda_rca32_and_28_22_y0;
  wire h_s_dadda_rca32_and_27_23_y0;
  wire h_s_dadda_rca32_and_26_24_y0;
  wire h_s_dadda_rca32_fa644_y2;
  wire h_s_dadda_rca32_fa644_y4;
  wire h_s_dadda_rca32_and_25_25_y0;
  wire h_s_dadda_rca32_and_24_26_y0;
  wire h_s_dadda_rca32_and_23_27_y0;
  wire h_s_dadda_rca32_fa645_y2;
  wire h_s_dadda_rca32_fa645_y4;
  wire h_s_dadda_rca32_and_22_28_y0;
  wire h_s_dadda_rca32_and_21_29_y0;
  wire h_s_dadda_rca32_and_20_30_y0;
  wire h_s_dadda_rca32_fa646_y2;
  wire h_s_dadda_rca32_fa646_y4;
  wire h_s_dadda_rca32_nand_19_31_y0;
  wire h_s_dadda_rca32_fa647_y2;
  wire h_s_dadda_rca32_fa647_y4;
  wire h_s_dadda_rca32_fa648_y2;
  wire h_s_dadda_rca32_fa648_y4;
  wire h_s_dadda_rca32_fa649_y2;
  wire h_s_dadda_rca32_fa649_y4;
  wire h_s_dadda_rca32_nand_31_20_y0;
  wire h_s_dadda_rca32_fa650_y2;
  wire h_s_dadda_rca32_fa650_y4;
  wire h_s_dadda_rca32_and_30_21_y0;
  wire h_s_dadda_rca32_and_29_22_y0;
  wire h_s_dadda_rca32_and_28_23_y0;
  wire h_s_dadda_rca32_fa651_y2;
  wire h_s_dadda_rca32_fa651_y4;
  wire h_s_dadda_rca32_and_27_24_y0;
  wire h_s_dadda_rca32_and_26_25_y0;
  wire h_s_dadda_rca32_and_25_26_y0;
  wire h_s_dadda_rca32_fa652_y2;
  wire h_s_dadda_rca32_fa652_y4;
  wire h_s_dadda_rca32_and_24_27_y0;
  wire h_s_dadda_rca32_and_23_28_y0;
  wire h_s_dadda_rca32_and_22_29_y0;
  wire h_s_dadda_rca32_fa653_y2;
  wire h_s_dadda_rca32_fa653_y4;
  wire h_s_dadda_rca32_and_21_30_y0;
  wire h_s_dadda_rca32_nand_20_31_y0;
  wire h_s_dadda_rca32_fa654_y2;
  wire h_s_dadda_rca32_fa654_y4;
  wire h_s_dadda_rca32_fa655_y2;
  wire h_s_dadda_rca32_fa655_y4;
  wire h_s_dadda_rca32_fa656_y2;
  wire h_s_dadda_rca32_fa656_y4;
  wire h_s_dadda_rca32_nand_31_21_y0;
  wire h_s_dadda_rca32_and_30_22_y0;
  wire h_s_dadda_rca32_fa657_y2;
  wire h_s_dadda_rca32_fa657_y4;
  wire h_s_dadda_rca32_and_29_23_y0;
  wire h_s_dadda_rca32_and_28_24_y0;
  wire h_s_dadda_rca32_and_27_25_y0;
  wire h_s_dadda_rca32_fa658_y2;
  wire h_s_dadda_rca32_fa658_y4;
  wire h_s_dadda_rca32_and_26_26_y0;
  wire h_s_dadda_rca32_and_25_27_y0;
  wire h_s_dadda_rca32_and_24_28_y0;
  wire h_s_dadda_rca32_fa659_y2;
  wire h_s_dadda_rca32_fa659_y4;
  wire h_s_dadda_rca32_and_23_29_y0;
  wire h_s_dadda_rca32_and_22_30_y0;
  wire h_s_dadda_rca32_nand_21_31_y0;
  wire h_s_dadda_rca32_fa660_y2;
  wire h_s_dadda_rca32_fa660_y4;
  wire h_s_dadda_rca32_fa661_y2;
  wire h_s_dadda_rca32_fa661_y4;
  wire h_s_dadda_rca32_fa662_y2;
  wire h_s_dadda_rca32_fa662_y4;
  wire h_s_dadda_rca32_nand_31_22_y0;
  wire h_s_dadda_rca32_and_30_23_y0;
  wire h_s_dadda_rca32_and_29_24_y0;
  wire h_s_dadda_rca32_fa663_y2;
  wire h_s_dadda_rca32_fa663_y4;
  wire h_s_dadda_rca32_and_28_25_y0;
  wire h_s_dadda_rca32_and_27_26_y0;
  wire h_s_dadda_rca32_and_26_27_y0;
  wire h_s_dadda_rca32_fa664_y2;
  wire h_s_dadda_rca32_fa664_y4;
  wire h_s_dadda_rca32_and_25_28_y0;
  wire h_s_dadda_rca32_and_24_29_y0;
  wire h_s_dadda_rca32_and_23_30_y0;
  wire h_s_dadda_rca32_fa665_y2;
  wire h_s_dadda_rca32_fa665_y4;
  wire h_s_dadda_rca32_fa666_y2;
  wire h_s_dadda_rca32_fa666_y4;
  wire h_s_dadda_rca32_nand_31_23_y0;
  wire h_s_dadda_rca32_fa667_y2;
  wire h_s_dadda_rca32_fa667_y4;
  wire h_s_dadda_rca32_and_30_24_y0;
  wire h_s_dadda_rca32_and_29_25_y0;
  wire h_s_dadda_rca32_and_28_26_y0;
  wire h_s_dadda_rca32_fa668_y2;
  wire h_s_dadda_rca32_fa668_y4;
  wire h_s_dadda_rca32_and_27_27_y0;
  wire h_s_dadda_rca32_and_26_28_y0;
  wire h_s_dadda_rca32_and_25_29_y0;
  wire h_s_dadda_rca32_fa669_y2;
  wire h_s_dadda_rca32_fa669_y4;
  wire h_s_dadda_rca32_fa670_y2;
  wire h_s_dadda_rca32_fa670_y4;
  wire h_s_dadda_rca32_nand_31_24_y0;
  wire h_s_dadda_rca32_and_30_25_y0;
  wire h_s_dadda_rca32_fa671_y2;
  wire h_s_dadda_rca32_fa671_y4;
  wire h_s_dadda_rca32_and_29_26_y0;
  wire h_s_dadda_rca32_and_28_27_y0;
  wire h_s_dadda_rca32_and_27_28_y0;
  wire h_s_dadda_rca32_fa672_y2;
  wire h_s_dadda_rca32_fa672_y4;
  wire h_s_dadda_rca32_fa673_y2;
  wire h_s_dadda_rca32_fa673_y4;
  wire h_s_dadda_rca32_nand_31_25_y0;
  wire h_s_dadda_rca32_and_30_26_y0;
  wire h_s_dadda_rca32_and_29_27_y0;
  wire h_s_dadda_rca32_fa674_y2;
  wire h_s_dadda_rca32_fa674_y4;
  wire h_s_dadda_rca32_nand_31_26_y0;
  wire h_s_dadda_rca32_fa675_y2;
  wire h_s_dadda_rca32_fa675_y4;
  wire h_s_dadda_rca32_and_4_0_y0;
  wire h_s_dadda_rca32_and_3_1_y0;
  wire h_s_dadda_rca32_ha26_y0;
  wire h_s_dadda_rca32_ha26_y1;
  wire h_s_dadda_rca32_and_5_0_y0;
  wire h_s_dadda_rca32_and_4_1_y0;
  wire h_s_dadda_rca32_fa676_y2;
  wire h_s_dadda_rca32_fa676_y4;
  wire h_s_dadda_rca32_and_3_2_y0;
  wire h_s_dadda_rca32_and_2_3_y0;
  wire h_s_dadda_rca32_ha27_y0;
  wire h_s_dadda_rca32_ha27_y1;
  wire h_s_dadda_rca32_and_4_2_y0;
  wire h_s_dadda_rca32_fa677_y2;
  wire h_s_dadda_rca32_fa677_y4;
  wire h_s_dadda_rca32_and_3_3_y0;
  wire h_s_dadda_rca32_and_2_4_y0;
  wire h_s_dadda_rca32_and_1_5_y0;
  wire h_s_dadda_rca32_fa678_y2;
  wire h_s_dadda_rca32_fa678_y4;
  wire h_s_dadda_rca32_and_3_4_y0;
  wire h_s_dadda_rca32_fa679_y2;
  wire h_s_dadda_rca32_fa679_y4;
  wire h_s_dadda_rca32_and_2_5_y0;
  wire h_s_dadda_rca32_and_1_6_y0;
  wire h_s_dadda_rca32_and_0_7_y0;
  wire h_s_dadda_rca32_fa680_y2;
  wire h_s_dadda_rca32_fa680_y4;
  wire h_s_dadda_rca32_and_2_6_y0;
  wire h_s_dadda_rca32_fa681_y2;
  wire h_s_dadda_rca32_fa681_y4;
  wire h_s_dadda_rca32_and_1_7_y0;
  wire h_s_dadda_rca32_and_0_8_y0;
  wire h_s_dadda_rca32_fa682_y2;
  wire h_s_dadda_rca32_fa682_y4;
  wire h_s_dadda_rca32_and_1_8_y0;
  wire h_s_dadda_rca32_fa683_y2;
  wire h_s_dadda_rca32_fa683_y4;
  wire h_s_dadda_rca32_and_0_9_y0;
  wire h_s_dadda_rca32_fa684_y2;
  wire h_s_dadda_rca32_fa684_y4;
  wire h_s_dadda_rca32_and_0_10_y0;
  wire h_s_dadda_rca32_fa685_y2;
  wire h_s_dadda_rca32_fa685_y4;
  wire h_s_dadda_rca32_fa686_y2;
  wire h_s_dadda_rca32_fa686_y4;
  wire h_s_dadda_rca32_fa687_y2;
  wire h_s_dadda_rca32_fa687_y4;
  wire h_s_dadda_rca32_fa688_y2;
  wire h_s_dadda_rca32_fa688_y4;
  wire h_s_dadda_rca32_fa689_y2;
  wire h_s_dadda_rca32_fa689_y4;
  wire h_s_dadda_rca32_fa690_y2;
  wire h_s_dadda_rca32_fa690_y4;
  wire h_s_dadda_rca32_fa691_y2;
  wire h_s_dadda_rca32_fa691_y4;
  wire h_s_dadda_rca32_fa692_y2;
  wire h_s_dadda_rca32_fa692_y4;
  wire h_s_dadda_rca32_fa693_y2;
  wire h_s_dadda_rca32_fa693_y4;
  wire h_s_dadda_rca32_fa694_y2;
  wire h_s_dadda_rca32_fa694_y4;
  wire h_s_dadda_rca32_fa695_y2;
  wire h_s_dadda_rca32_fa695_y4;
  wire h_s_dadda_rca32_fa696_y2;
  wire h_s_dadda_rca32_fa696_y4;
  wire h_s_dadda_rca32_fa697_y2;
  wire h_s_dadda_rca32_fa697_y4;
  wire h_s_dadda_rca32_fa698_y2;
  wire h_s_dadda_rca32_fa698_y4;
  wire h_s_dadda_rca32_fa699_y2;
  wire h_s_dadda_rca32_fa699_y4;
  wire h_s_dadda_rca32_fa700_y2;
  wire h_s_dadda_rca32_fa700_y4;
  wire h_s_dadda_rca32_fa701_y2;
  wire h_s_dadda_rca32_fa701_y4;
  wire h_s_dadda_rca32_fa702_y2;
  wire h_s_dadda_rca32_fa702_y4;
  wire h_s_dadda_rca32_fa703_y2;
  wire h_s_dadda_rca32_fa703_y4;
  wire h_s_dadda_rca32_fa704_y2;
  wire h_s_dadda_rca32_fa704_y4;
  wire h_s_dadda_rca32_fa705_y2;
  wire h_s_dadda_rca32_fa705_y4;
  wire h_s_dadda_rca32_fa706_y2;
  wire h_s_dadda_rca32_fa706_y4;
  wire h_s_dadda_rca32_fa707_y2;
  wire h_s_dadda_rca32_fa707_y4;
  wire h_s_dadda_rca32_fa708_y2;
  wire h_s_dadda_rca32_fa708_y4;
  wire h_s_dadda_rca32_fa709_y2;
  wire h_s_dadda_rca32_fa709_y4;
  wire h_s_dadda_rca32_fa710_y2;
  wire h_s_dadda_rca32_fa710_y4;
  wire h_s_dadda_rca32_fa711_y2;
  wire h_s_dadda_rca32_fa711_y4;
  wire h_s_dadda_rca32_fa712_y2;
  wire h_s_dadda_rca32_fa712_y4;
  wire h_s_dadda_rca32_fa713_y2;
  wire h_s_dadda_rca32_fa713_y4;
  wire h_s_dadda_rca32_fa714_y2;
  wire h_s_dadda_rca32_fa714_y4;
  wire h_s_dadda_rca32_fa715_y2;
  wire h_s_dadda_rca32_fa715_y4;
  wire h_s_dadda_rca32_fa716_y2;
  wire h_s_dadda_rca32_fa716_y4;
  wire h_s_dadda_rca32_fa717_y2;
  wire h_s_dadda_rca32_fa717_y4;
  wire h_s_dadda_rca32_fa718_y2;
  wire h_s_dadda_rca32_fa718_y4;
  wire h_s_dadda_rca32_fa719_y2;
  wire h_s_dadda_rca32_fa719_y4;
  wire h_s_dadda_rca32_fa720_y2;
  wire h_s_dadda_rca32_fa720_y4;
  wire h_s_dadda_rca32_fa721_y2;
  wire h_s_dadda_rca32_fa721_y4;
  wire h_s_dadda_rca32_fa722_y2;
  wire h_s_dadda_rca32_fa722_y4;
  wire h_s_dadda_rca32_fa723_y2;
  wire h_s_dadda_rca32_fa723_y4;
  wire h_s_dadda_rca32_fa724_y2;
  wire h_s_dadda_rca32_fa724_y4;
  wire h_s_dadda_rca32_fa725_y2;
  wire h_s_dadda_rca32_fa725_y4;
  wire h_s_dadda_rca32_fa726_y2;
  wire h_s_dadda_rca32_fa726_y4;
  wire h_s_dadda_rca32_fa727_y2;
  wire h_s_dadda_rca32_fa727_y4;
  wire h_s_dadda_rca32_fa728_y2;
  wire h_s_dadda_rca32_fa728_y4;
  wire h_s_dadda_rca32_fa729_y2;
  wire h_s_dadda_rca32_fa729_y4;
  wire h_s_dadda_rca32_fa730_y2;
  wire h_s_dadda_rca32_fa730_y4;
  wire h_s_dadda_rca32_fa731_y2;
  wire h_s_dadda_rca32_fa731_y4;
  wire h_s_dadda_rca32_fa732_y2;
  wire h_s_dadda_rca32_fa732_y4;
  wire h_s_dadda_rca32_fa733_y2;
  wire h_s_dadda_rca32_fa733_y4;
  wire h_s_dadda_rca32_fa734_y2;
  wire h_s_dadda_rca32_fa734_y4;
  wire h_s_dadda_rca32_fa735_y2;
  wire h_s_dadda_rca32_fa735_y4;
  wire h_s_dadda_rca32_fa736_y2;
  wire h_s_dadda_rca32_fa736_y4;
  wire h_s_dadda_rca32_fa737_y2;
  wire h_s_dadda_rca32_fa737_y4;
  wire h_s_dadda_rca32_fa738_y2;
  wire h_s_dadda_rca32_fa738_y4;
  wire h_s_dadda_rca32_fa739_y2;
  wire h_s_dadda_rca32_fa739_y4;
  wire h_s_dadda_rca32_fa740_y2;
  wire h_s_dadda_rca32_fa740_y4;
  wire h_s_dadda_rca32_fa741_y2;
  wire h_s_dadda_rca32_fa741_y4;
  wire h_s_dadda_rca32_fa742_y2;
  wire h_s_dadda_rca32_fa742_y4;
  wire h_s_dadda_rca32_fa743_y2;
  wire h_s_dadda_rca32_fa743_y4;
  wire h_s_dadda_rca32_fa744_y2;
  wire h_s_dadda_rca32_fa744_y4;
  wire h_s_dadda_rca32_fa745_y2;
  wire h_s_dadda_rca32_fa745_y4;
  wire h_s_dadda_rca32_fa746_y2;
  wire h_s_dadda_rca32_fa746_y4;
  wire h_s_dadda_rca32_fa747_y2;
  wire h_s_dadda_rca32_fa747_y4;
  wire h_s_dadda_rca32_fa748_y2;
  wire h_s_dadda_rca32_fa748_y4;
  wire h_s_dadda_rca32_fa749_y2;
  wire h_s_dadda_rca32_fa749_y4;
  wire h_s_dadda_rca32_fa750_y2;
  wire h_s_dadda_rca32_fa750_y4;
  wire h_s_dadda_rca32_fa751_y2;
  wire h_s_dadda_rca32_fa751_y4;
  wire h_s_dadda_rca32_fa752_y2;
  wire h_s_dadda_rca32_fa752_y4;
  wire h_s_dadda_rca32_fa753_y2;
  wire h_s_dadda_rca32_fa753_y4;
  wire h_s_dadda_rca32_fa754_y2;
  wire h_s_dadda_rca32_fa754_y4;
  wire h_s_dadda_rca32_fa755_y2;
  wire h_s_dadda_rca32_fa755_y4;
  wire h_s_dadda_rca32_fa756_y2;
  wire h_s_dadda_rca32_fa756_y4;
  wire h_s_dadda_rca32_fa757_y2;
  wire h_s_dadda_rca32_fa757_y4;
  wire h_s_dadda_rca32_fa758_y2;
  wire h_s_dadda_rca32_fa758_y4;
  wire h_s_dadda_rca32_fa759_y2;
  wire h_s_dadda_rca32_fa759_y4;
  wire h_s_dadda_rca32_fa760_y2;
  wire h_s_dadda_rca32_fa760_y4;
  wire h_s_dadda_rca32_fa761_y2;
  wire h_s_dadda_rca32_fa761_y4;
  wire h_s_dadda_rca32_fa762_y2;
  wire h_s_dadda_rca32_fa762_y4;
  wire h_s_dadda_rca32_fa763_y2;
  wire h_s_dadda_rca32_fa763_y4;
  wire h_s_dadda_rca32_fa764_y2;
  wire h_s_dadda_rca32_fa764_y4;
  wire h_s_dadda_rca32_fa765_y2;
  wire h_s_dadda_rca32_fa765_y4;
  wire h_s_dadda_rca32_fa766_y2;
  wire h_s_dadda_rca32_fa766_y4;
  wire h_s_dadda_rca32_fa767_y2;
  wire h_s_dadda_rca32_fa767_y4;
  wire h_s_dadda_rca32_fa768_y2;
  wire h_s_dadda_rca32_fa768_y4;
  wire h_s_dadda_rca32_fa769_y2;
  wire h_s_dadda_rca32_fa769_y4;
  wire h_s_dadda_rca32_fa770_y2;
  wire h_s_dadda_rca32_fa770_y4;
  wire h_s_dadda_rca32_nand_22_31_y0;
  wire h_s_dadda_rca32_fa771_y2;
  wire h_s_dadda_rca32_fa771_y4;
  wire h_s_dadda_rca32_fa772_y2;
  wire h_s_dadda_rca32_fa772_y4;
  wire h_s_dadda_rca32_and_24_30_y0;
  wire h_s_dadda_rca32_fa773_y2;
  wire h_s_dadda_rca32_fa773_y4;
  wire h_s_dadda_rca32_nand_23_31_y0;
  wire h_s_dadda_rca32_fa774_y2;
  wire h_s_dadda_rca32_fa774_y4;
  wire h_s_dadda_rca32_and_26_29_y0;
  wire h_s_dadda_rca32_fa775_y2;
  wire h_s_dadda_rca32_fa775_y4;
  wire h_s_dadda_rca32_and_25_30_y0;
  wire h_s_dadda_rca32_nand_24_31_y0;
  wire h_s_dadda_rca32_fa776_y2;
  wire h_s_dadda_rca32_fa776_y4;
  wire h_s_dadda_rca32_and_28_28_y0;
  wire h_s_dadda_rca32_fa777_y2;
  wire h_s_dadda_rca32_fa777_y4;
  wire h_s_dadda_rca32_and_27_29_y0;
  wire h_s_dadda_rca32_and_26_30_y0;
  wire h_s_dadda_rca32_nand_25_31_y0;
  wire h_s_dadda_rca32_fa778_y2;
  wire h_s_dadda_rca32_fa778_y4;
  wire h_s_dadda_rca32_and_30_27_y0;
  wire h_s_dadda_rca32_fa779_y2;
  wire h_s_dadda_rca32_fa779_y4;
  wire h_s_dadda_rca32_and_29_28_y0;
  wire h_s_dadda_rca32_and_28_29_y0;
  wire h_s_dadda_rca32_and_27_30_y0;
  wire h_s_dadda_rca32_fa780_y2;
  wire h_s_dadda_rca32_fa780_y4;
  wire h_s_dadda_rca32_fa781_y2;
  wire h_s_dadda_rca32_fa781_y4;
  wire h_s_dadda_rca32_nand_31_27_y0;
  wire h_s_dadda_rca32_and_30_28_y0;
  wire h_s_dadda_rca32_and_29_29_y0;
  wire h_s_dadda_rca32_fa782_y2;
  wire h_s_dadda_rca32_fa782_y4;
  wire h_s_dadda_rca32_nand_31_28_y0;
  wire h_s_dadda_rca32_fa783_y2;
  wire h_s_dadda_rca32_fa783_y4;
  wire h_s_dadda_rca32_and_3_0_y0;
  wire h_s_dadda_rca32_and_2_1_y0;
  wire h_s_dadda_rca32_ha28_y0;
  wire h_s_dadda_rca32_ha28_y1;
  wire h_s_dadda_rca32_and_2_2_y0;
  wire h_s_dadda_rca32_and_1_3_y0;
  wire h_s_dadda_rca32_fa784_y2;
  wire h_s_dadda_rca32_fa784_y4;
  wire h_s_dadda_rca32_and_1_4_y0;
  wire h_s_dadda_rca32_and_0_5_y0;
  wire h_s_dadda_rca32_fa785_y2;
  wire h_s_dadda_rca32_fa785_y4;
  wire h_s_dadda_rca32_and_0_6_y0;
  wire h_s_dadda_rca32_fa786_y2;
  wire h_s_dadda_rca32_fa786_y4;
  wire h_s_dadda_rca32_fa787_y2;
  wire h_s_dadda_rca32_fa787_y4;
  wire h_s_dadda_rca32_fa788_y2;
  wire h_s_dadda_rca32_fa788_y4;
  wire h_s_dadda_rca32_fa789_y2;
  wire h_s_dadda_rca32_fa789_y4;
  wire h_s_dadda_rca32_fa790_y2;
  wire h_s_dadda_rca32_fa790_y4;
  wire h_s_dadda_rca32_fa791_y2;
  wire h_s_dadda_rca32_fa791_y4;
  wire h_s_dadda_rca32_fa792_y2;
  wire h_s_dadda_rca32_fa792_y4;
  wire h_s_dadda_rca32_fa793_y2;
  wire h_s_dadda_rca32_fa793_y4;
  wire h_s_dadda_rca32_fa794_y2;
  wire h_s_dadda_rca32_fa794_y4;
  wire h_s_dadda_rca32_fa795_y2;
  wire h_s_dadda_rca32_fa795_y4;
  wire h_s_dadda_rca32_fa796_y2;
  wire h_s_dadda_rca32_fa796_y4;
  wire h_s_dadda_rca32_fa797_y2;
  wire h_s_dadda_rca32_fa797_y4;
  wire h_s_dadda_rca32_fa798_y2;
  wire h_s_dadda_rca32_fa798_y4;
  wire h_s_dadda_rca32_fa799_y2;
  wire h_s_dadda_rca32_fa799_y4;
  wire h_s_dadda_rca32_fa800_y2;
  wire h_s_dadda_rca32_fa800_y4;
  wire h_s_dadda_rca32_fa801_y2;
  wire h_s_dadda_rca32_fa801_y4;
  wire h_s_dadda_rca32_fa802_y2;
  wire h_s_dadda_rca32_fa802_y4;
  wire h_s_dadda_rca32_fa803_y2;
  wire h_s_dadda_rca32_fa803_y4;
  wire h_s_dadda_rca32_fa804_y2;
  wire h_s_dadda_rca32_fa804_y4;
  wire h_s_dadda_rca32_fa805_y2;
  wire h_s_dadda_rca32_fa805_y4;
  wire h_s_dadda_rca32_fa806_y2;
  wire h_s_dadda_rca32_fa806_y4;
  wire h_s_dadda_rca32_fa807_y2;
  wire h_s_dadda_rca32_fa807_y4;
  wire h_s_dadda_rca32_fa808_y2;
  wire h_s_dadda_rca32_fa808_y4;
  wire h_s_dadda_rca32_fa809_y2;
  wire h_s_dadda_rca32_fa809_y4;
  wire h_s_dadda_rca32_fa810_y2;
  wire h_s_dadda_rca32_fa810_y4;
  wire h_s_dadda_rca32_fa811_y2;
  wire h_s_dadda_rca32_fa811_y4;
  wire h_s_dadda_rca32_fa812_y2;
  wire h_s_dadda_rca32_fa812_y4;
  wire h_s_dadda_rca32_fa813_y2;
  wire h_s_dadda_rca32_fa813_y4;
  wire h_s_dadda_rca32_fa814_y2;
  wire h_s_dadda_rca32_fa814_y4;
  wire h_s_dadda_rca32_fa815_y2;
  wire h_s_dadda_rca32_fa815_y4;
  wire h_s_dadda_rca32_fa816_y2;
  wire h_s_dadda_rca32_fa816_y4;
  wire h_s_dadda_rca32_fa817_y2;
  wire h_s_dadda_rca32_fa817_y4;
  wire h_s_dadda_rca32_fa818_y2;
  wire h_s_dadda_rca32_fa818_y4;
  wire h_s_dadda_rca32_fa819_y2;
  wire h_s_dadda_rca32_fa819_y4;
  wire h_s_dadda_rca32_fa820_y2;
  wire h_s_dadda_rca32_fa820_y4;
  wire h_s_dadda_rca32_fa821_y2;
  wire h_s_dadda_rca32_fa821_y4;
  wire h_s_dadda_rca32_fa822_y2;
  wire h_s_dadda_rca32_fa822_y4;
  wire h_s_dadda_rca32_fa823_y2;
  wire h_s_dadda_rca32_fa823_y4;
  wire h_s_dadda_rca32_fa824_y2;
  wire h_s_dadda_rca32_fa824_y4;
  wire h_s_dadda_rca32_fa825_y2;
  wire h_s_dadda_rca32_fa825_y4;
  wire h_s_dadda_rca32_fa826_y2;
  wire h_s_dadda_rca32_fa826_y4;
  wire h_s_dadda_rca32_fa827_y2;
  wire h_s_dadda_rca32_fa827_y4;
  wire h_s_dadda_rca32_fa828_y2;
  wire h_s_dadda_rca32_fa828_y4;
  wire h_s_dadda_rca32_fa829_y2;
  wire h_s_dadda_rca32_fa829_y4;
  wire h_s_dadda_rca32_fa830_y2;
  wire h_s_dadda_rca32_fa830_y4;
  wire h_s_dadda_rca32_fa831_y2;
  wire h_s_dadda_rca32_fa831_y4;
  wire h_s_dadda_rca32_fa832_y2;
  wire h_s_dadda_rca32_fa832_y4;
  wire h_s_dadda_rca32_fa833_y2;
  wire h_s_dadda_rca32_fa833_y4;
  wire h_s_dadda_rca32_fa834_y2;
  wire h_s_dadda_rca32_fa834_y4;
  wire h_s_dadda_rca32_fa835_y2;
  wire h_s_dadda_rca32_fa835_y4;
  wire h_s_dadda_rca32_fa836_y2;
  wire h_s_dadda_rca32_fa836_y4;
  wire h_s_dadda_rca32_nand_26_31_y0;
  wire h_s_dadda_rca32_fa837_y2;
  wire h_s_dadda_rca32_fa837_y4;
  wire h_s_dadda_rca32_and_28_30_y0;
  wire h_s_dadda_rca32_nand_27_31_y0;
  wire h_s_dadda_rca32_fa838_y2;
  wire h_s_dadda_rca32_fa838_y4;
  wire h_s_dadda_rca32_and_30_29_y0;
  wire h_s_dadda_rca32_and_29_30_y0;
  wire h_s_dadda_rca32_fa839_y2;
  wire h_s_dadda_rca32_fa839_y4;
  wire h_s_dadda_rca32_nand_31_29_y0;
  wire h_s_dadda_rca32_fa840_y2;
  wire h_s_dadda_rca32_fa840_y4;
  wire h_s_dadda_rca32_and_2_0_y0;
  wire h_s_dadda_rca32_and_1_1_y0;
  wire h_s_dadda_rca32_ha29_y0;
  wire h_s_dadda_rca32_ha29_y1;
  wire h_s_dadda_rca32_and_1_2_y0;
  wire h_s_dadda_rca32_and_0_3_y0;
  wire h_s_dadda_rca32_fa841_y2;
  wire h_s_dadda_rca32_fa841_y4;
  wire h_s_dadda_rca32_and_0_4_y0;
  wire h_s_dadda_rca32_fa842_y2;
  wire h_s_dadda_rca32_fa842_y4;
  wire h_s_dadda_rca32_fa843_y2;
  wire h_s_dadda_rca32_fa843_y4;
  wire h_s_dadda_rca32_fa844_y2;
  wire h_s_dadda_rca32_fa844_y4;
  wire h_s_dadda_rca32_fa845_y2;
  wire h_s_dadda_rca32_fa845_y4;
  wire h_s_dadda_rca32_fa846_y2;
  wire h_s_dadda_rca32_fa846_y4;
  wire h_s_dadda_rca32_fa847_y2;
  wire h_s_dadda_rca32_fa847_y4;
  wire h_s_dadda_rca32_fa848_y2;
  wire h_s_dadda_rca32_fa848_y4;
  wire h_s_dadda_rca32_fa849_y2;
  wire h_s_dadda_rca32_fa849_y4;
  wire h_s_dadda_rca32_fa850_y2;
  wire h_s_dadda_rca32_fa850_y4;
  wire h_s_dadda_rca32_fa851_y2;
  wire h_s_dadda_rca32_fa851_y4;
  wire h_s_dadda_rca32_fa852_y2;
  wire h_s_dadda_rca32_fa852_y4;
  wire h_s_dadda_rca32_fa853_y2;
  wire h_s_dadda_rca32_fa853_y4;
  wire h_s_dadda_rca32_fa854_y2;
  wire h_s_dadda_rca32_fa854_y4;
  wire h_s_dadda_rca32_fa855_y2;
  wire h_s_dadda_rca32_fa855_y4;
  wire h_s_dadda_rca32_fa856_y2;
  wire h_s_dadda_rca32_fa856_y4;
  wire h_s_dadda_rca32_fa857_y2;
  wire h_s_dadda_rca32_fa857_y4;
  wire h_s_dadda_rca32_fa858_y2;
  wire h_s_dadda_rca32_fa858_y4;
  wire h_s_dadda_rca32_fa859_y2;
  wire h_s_dadda_rca32_fa859_y4;
  wire h_s_dadda_rca32_fa860_y2;
  wire h_s_dadda_rca32_fa860_y4;
  wire h_s_dadda_rca32_fa861_y2;
  wire h_s_dadda_rca32_fa861_y4;
  wire h_s_dadda_rca32_fa862_y2;
  wire h_s_dadda_rca32_fa862_y4;
  wire h_s_dadda_rca32_fa863_y2;
  wire h_s_dadda_rca32_fa863_y4;
  wire h_s_dadda_rca32_fa864_y2;
  wire h_s_dadda_rca32_fa864_y4;
  wire h_s_dadda_rca32_fa865_y2;
  wire h_s_dadda_rca32_fa865_y4;
  wire h_s_dadda_rca32_fa866_y2;
  wire h_s_dadda_rca32_fa866_y4;
  wire h_s_dadda_rca32_fa867_y2;
  wire h_s_dadda_rca32_fa867_y4;
  wire h_s_dadda_rca32_fa868_y2;
  wire h_s_dadda_rca32_fa868_y4;
  wire h_s_dadda_rca32_fa869_y2;
  wire h_s_dadda_rca32_fa869_y4;
  wire h_s_dadda_rca32_fa870_y2;
  wire h_s_dadda_rca32_fa870_y4;
  wire h_s_dadda_rca32_fa871_y2;
  wire h_s_dadda_rca32_fa871_y4;
  wire h_s_dadda_rca32_fa872_y2;
  wire h_s_dadda_rca32_fa872_y4;
  wire h_s_dadda_rca32_fa873_y2;
  wire h_s_dadda_rca32_fa873_y4;
  wire h_s_dadda_rca32_fa874_y2;
  wire h_s_dadda_rca32_fa874_y4;
  wire h_s_dadda_rca32_fa875_y2;
  wire h_s_dadda_rca32_fa875_y4;
  wire h_s_dadda_rca32_fa876_y2;
  wire h_s_dadda_rca32_fa876_y4;
  wire h_s_dadda_rca32_fa877_y2;
  wire h_s_dadda_rca32_fa877_y4;
  wire h_s_dadda_rca32_fa878_y2;
  wire h_s_dadda_rca32_fa878_y4;
  wire h_s_dadda_rca32_fa879_y2;
  wire h_s_dadda_rca32_fa879_y4;
  wire h_s_dadda_rca32_fa880_y2;
  wire h_s_dadda_rca32_fa880_y4;
  wire h_s_dadda_rca32_fa881_y2;
  wire h_s_dadda_rca32_fa881_y4;
  wire h_s_dadda_rca32_fa882_y2;
  wire h_s_dadda_rca32_fa882_y4;
  wire h_s_dadda_rca32_fa883_y2;
  wire h_s_dadda_rca32_fa883_y4;
  wire h_s_dadda_rca32_fa884_y2;
  wire h_s_dadda_rca32_fa884_y4;
  wire h_s_dadda_rca32_fa885_y2;
  wire h_s_dadda_rca32_fa885_y4;
  wire h_s_dadda_rca32_fa886_y2;
  wire h_s_dadda_rca32_fa886_y4;
  wire h_s_dadda_rca32_fa887_y2;
  wire h_s_dadda_rca32_fa887_y4;
  wire h_s_dadda_rca32_fa888_y2;
  wire h_s_dadda_rca32_fa888_y4;
  wire h_s_dadda_rca32_fa889_y2;
  wire h_s_dadda_rca32_fa889_y4;
  wire h_s_dadda_rca32_fa890_y2;
  wire h_s_dadda_rca32_fa890_y4;
  wire h_s_dadda_rca32_fa891_y2;
  wire h_s_dadda_rca32_fa891_y4;
  wire h_s_dadda_rca32_fa892_y2;
  wire h_s_dadda_rca32_fa892_y4;
  wire h_s_dadda_rca32_fa893_y2;
  wire h_s_dadda_rca32_fa893_y4;
  wire h_s_dadda_rca32_fa894_y2;
  wire h_s_dadda_rca32_fa894_y4;
  wire h_s_dadda_rca32_fa895_y2;
  wire h_s_dadda_rca32_fa895_y4;
  wire h_s_dadda_rca32_fa896_y2;
  wire h_s_dadda_rca32_fa896_y4;
  wire h_s_dadda_rca32_nand_28_31_y0;
  wire h_s_dadda_rca32_fa897_y2;
  wire h_s_dadda_rca32_fa897_y4;
  wire h_s_dadda_rca32_and_30_30_y0;
  wire h_s_dadda_rca32_nand_29_31_y0;
  wire h_s_dadda_rca32_fa898_y2;
  wire h_s_dadda_rca32_fa898_y4;
  wire h_s_dadda_rca32_nand_31_30_y0;
  wire h_s_dadda_rca32_fa899_y2;
  wire h_s_dadda_rca32_fa899_y4;
  wire h_s_dadda_rca32_and_0_0_y0;
  wire h_s_dadda_rca32_and_1_0_y0;
  wire h_s_dadda_rca32_and_0_2_y0;
  wire h_s_dadda_rca32_nand_30_31_y0;
  wire h_s_dadda_rca32_and_0_1_y0;
  wire h_s_dadda_rca32_and_31_31_y0;
  wire [61:0] h_s_dadda_rca32_u_rca62_u_rca62_a;
  wire [61:0] h_s_dadda_rca32_u_rca62_u_rca62_b;
  wire [62:0] h_s_dadda_rca32_u_rca62_out;
  wire h_s_dadda_rca32_u_rca62_ha_y0;
  wire h_s_dadda_rca32_u_rca62_fa1_y2;
  wire h_s_dadda_rca32_u_rca62_fa2_y2;
  wire h_s_dadda_rca32_u_rca62_fa3_y2;
  wire h_s_dadda_rca32_u_rca62_fa4_y2;
  wire h_s_dadda_rca32_u_rca62_fa5_y2;
  wire h_s_dadda_rca32_u_rca62_fa6_y2;
  wire h_s_dadda_rca32_u_rca62_fa7_y2;
  wire h_s_dadda_rca32_u_rca62_fa8_y2;
  wire h_s_dadda_rca32_u_rca62_fa9_y2;
  wire h_s_dadda_rca32_u_rca62_fa10_y2;
  wire h_s_dadda_rca32_u_rca62_fa11_y2;
  wire h_s_dadda_rca32_u_rca62_fa12_y2;
  wire h_s_dadda_rca32_u_rca62_fa13_y2;
  wire h_s_dadda_rca32_u_rca62_fa14_y2;
  wire h_s_dadda_rca32_u_rca62_fa15_y2;
  wire h_s_dadda_rca32_u_rca62_fa16_y2;
  wire h_s_dadda_rca32_u_rca62_fa17_y2;
  wire h_s_dadda_rca32_u_rca62_fa18_y2;
  wire h_s_dadda_rca32_u_rca62_fa19_y2;
  wire h_s_dadda_rca32_u_rca62_fa20_y2;
  wire h_s_dadda_rca32_u_rca62_fa21_y2;
  wire h_s_dadda_rca32_u_rca62_fa22_y2;
  wire h_s_dadda_rca32_u_rca62_fa23_y2;
  wire h_s_dadda_rca32_u_rca62_fa24_y2;
  wire h_s_dadda_rca32_u_rca62_fa25_y2;
  wire h_s_dadda_rca32_u_rca62_fa26_y2;
  wire h_s_dadda_rca32_u_rca62_fa27_y2;
  wire h_s_dadda_rca32_u_rca62_fa28_y2;
  wire h_s_dadda_rca32_u_rca62_fa29_y2;
  wire h_s_dadda_rca32_u_rca62_fa30_y2;
  wire h_s_dadda_rca32_u_rca62_fa31_y2;
  wire h_s_dadda_rca32_u_rca62_fa32_y2;
  wire h_s_dadda_rca32_u_rca62_fa33_y2;
  wire h_s_dadda_rca32_u_rca62_fa34_y2;
  wire h_s_dadda_rca32_u_rca62_fa35_y2;
  wire h_s_dadda_rca32_u_rca62_fa36_y2;
  wire h_s_dadda_rca32_u_rca62_fa37_y2;
  wire h_s_dadda_rca32_u_rca62_fa38_y2;
  wire h_s_dadda_rca32_u_rca62_fa39_y2;
  wire h_s_dadda_rca32_u_rca62_fa40_y2;
  wire h_s_dadda_rca32_u_rca62_fa41_y2;
  wire h_s_dadda_rca32_u_rca62_fa42_y2;
  wire h_s_dadda_rca32_u_rca62_fa43_y2;
  wire h_s_dadda_rca32_u_rca62_fa44_y2;
  wire h_s_dadda_rca32_u_rca62_fa45_y2;
  wire h_s_dadda_rca32_u_rca62_fa46_y2;
  wire h_s_dadda_rca32_u_rca62_fa47_y2;
  wire h_s_dadda_rca32_u_rca62_fa48_y2;
  wire h_s_dadda_rca32_u_rca62_fa49_y2;
  wire h_s_dadda_rca32_u_rca62_fa50_y2;
  wire h_s_dadda_rca32_u_rca62_fa51_y2;
  wire h_s_dadda_rca32_u_rca62_fa52_y2;
  wire h_s_dadda_rca32_u_rca62_fa53_y2;
  wire h_s_dadda_rca32_u_rca62_fa54_y2;
  wire h_s_dadda_rca32_u_rca62_fa55_y2;
  wire h_s_dadda_rca32_u_rca62_fa56_y2;
  wire h_s_dadda_rca32_u_rca62_fa57_y2;
  wire h_s_dadda_rca32_u_rca62_fa58_y2;
  wire h_s_dadda_rca32_u_rca62_fa59_y2;
  wire h_s_dadda_rca32_u_rca62_fa60_y2;
  wire h_s_dadda_rca32_u_rca62_fa61_y2;
  wire h_s_dadda_rca32_u_rca62_fa61_y4;
  wire h_s_dadda_rca32_xor0_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign a_30 = a[30];
  assign a_31 = a[31];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  assign b_30 = b[30];
  assign b_31 = b[31];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_dadda_rca32_and_28_0_y0(a_28, b_0, h_s_dadda_rca32_and_28_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_1_y0(a_27, b_1, h_s_dadda_rca32_and_27_1_y0);
  ha ha_h_s_dadda_rca32_ha0_y0(h_s_dadda_rca32_and_28_0_y0, h_s_dadda_rca32_and_27_1_y0, h_s_dadda_rca32_ha0_y0, h_s_dadda_rca32_ha0_y1);
  and_gate and_gate_h_s_dadda_rca32_and_29_0_y0(a_29, b_0, h_s_dadda_rca32_and_29_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_1_y0(a_28, b_1, h_s_dadda_rca32_and_28_1_y0);
  fa fa_h_s_dadda_rca32_fa0_y2(h_s_dadda_rca32_ha0_y1, h_s_dadda_rca32_and_29_0_y0, h_s_dadda_rca32_and_28_1_y0, h_s_dadda_rca32_fa0_y2, h_s_dadda_rca32_fa0_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_2_y0(a_27, b_2, h_s_dadda_rca32_and_27_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_3_y0(a_26, b_3, h_s_dadda_rca32_and_26_3_y0);
  ha ha_h_s_dadda_rca32_ha1_y0(h_s_dadda_rca32_and_27_2_y0, h_s_dadda_rca32_and_26_3_y0, h_s_dadda_rca32_ha1_y0, h_s_dadda_rca32_ha1_y1);
  and_gate and_gate_h_s_dadda_rca32_and_30_0_y0(a_30, b_0, h_s_dadda_rca32_and_30_0_y0);
  fa fa_h_s_dadda_rca32_fa1_y2(h_s_dadda_rca32_ha1_y1, h_s_dadda_rca32_fa0_y4, h_s_dadda_rca32_and_30_0_y0, h_s_dadda_rca32_fa1_y2, h_s_dadda_rca32_fa1_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_1_y0(a_29, b_1, h_s_dadda_rca32_and_29_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_2_y0(a_28, b_2, h_s_dadda_rca32_and_28_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_3_y0(a_27, b_3, h_s_dadda_rca32_and_27_3_y0);
  fa fa_h_s_dadda_rca32_fa2_y2(h_s_dadda_rca32_and_29_1_y0, h_s_dadda_rca32_and_28_2_y0, h_s_dadda_rca32_and_27_3_y0, h_s_dadda_rca32_fa2_y2, h_s_dadda_rca32_fa2_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_4_y0(a_26, b_4, h_s_dadda_rca32_and_26_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_5_y0(a_25, b_5, h_s_dadda_rca32_and_25_5_y0);
  ha ha_h_s_dadda_rca32_ha2_y0(h_s_dadda_rca32_and_26_4_y0, h_s_dadda_rca32_and_25_5_y0, h_s_dadda_rca32_ha2_y0, h_s_dadda_rca32_ha2_y1);
  fa fa_h_s_dadda_rca32_fa3_y2(h_s_dadda_rca32_ha2_y1, h_s_dadda_rca32_fa2_y4, h_s_dadda_rca32_fa1_y4, h_s_dadda_rca32_fa3_y2, h_s_dadda_rca32_fa3_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_0_y0(a_31, b_0, h_s_dadda_rca32_nand_31_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_1_y0(a_30, b_1, h_s_dadda_rca32_and_30_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_2_y0(a_29, b_2, h_s_dadda_rca32_and_29_2_y0);
  fa fa_h_s_dadda_rca32_fa4_y2(h_s_dadda_rca32_nand_31_0_y0, h_s_dadda_rca32_and_30_1_y0, h_s_dadda_rca32_and_29_2_y0, h_s_dadda_rca32_fa4_y2, h_s_dadda_rca32_fa4_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_3_y0(a_28, b_3, h_s_dadda_rca32_and_28_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_4_y0(a_27, b_4, h_s_dadda_rca32_and_27_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_5_y0(a_26, b_5, h_s_dadda_rca32_and_26_5_y0);
  fa fa_h_s_dadda_rca32_fa5_y2(h_s_dadda_rca32_and_28_3_y0, h_s_dadda_rca32_and_27_4_y0, h_s_dadda_rca32_and_26_5_y0, h_s_dadda_rca32_fa5_y2, h_s_dadda_rca32_fa5_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_6_y0(a_25, b_6, h_s_dadda_rca32_and_25_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_7_y0(a_24, b_7, h_s_dadda_rca32_and_24_7_y0);
  ha ha_h_s_dadda_rca32_ha3_y0(h_s_dadda_rca32_and_25_6_y0, h_s_dadda_rca32_and_24_7_y0, h_s_dadda_rca32_ha3_y0, h_s_dadda_rca32_ha3_y1);
  fa fa_h_s_dadda_rca32_fa6_y2(h_s_dadda_rca32_ha3_y1, h_s_dadda_rca32_fa5_y4, h_s_dadda_rca32_fa4_y4, h_s_dadda_rca32_fa6_y2, h_s_dadda_rca32_fa6_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_1_y0(a_31, b_1, h_s_dadda_rca32_nand_31_1_y0);
  fa fa_h_s_dadda_rca32_fa7_y2(h_s_dadda_rca32_fa3_y4, constant_wire_1, h_s_dadda_rca32_nand_31_1_y0, h_s_dadda_rca32_fa7_y2, h_s_dadda_rca32_fa7_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_2_y0(a_30, b_2, h_s_dadda_rca32_and_30_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_3_y0(a_29, b_3, h_s_dadda_rca32_and_29_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_4_y0(a_28, b_4, h_s_dadda_rca32_and_28_4_y0);
  fa fa_h_s_dadda_rca32_fa8_y2(h_s_dadda_rca32_and_30_2_y0, h_s_dadda_rca32_and_29_3_y0, h_s_dadda_rca32_and_28_4_y0, h_s_dadda_rca32_fa8_y2, h_s_dadda_rca32_fa8_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_5_y0(a_27, b_5, h_s_dadda_rca32_and_27_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_6_y0(a_26, b_6, h_s_dadda_rca32_and_26_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_7_y0(a_25, b_7, h_s_dadda_rca32_and_25_7_y0);
  fa fa_h_s_dadda_rca32_fa9_y2(h_s_dadda_rca32_and_27_5_y0, h_s_dadda_rca32_and_26_6_y0, h_s_dadda_rca32_and_25_7_y0, h_s_dadda_rca32_fa9_y2, h_s_dadda_rca32_fa9_y4);
  fa fa_h_s_dadda_rca32_fa10_y2(h_s_dadda_rca32_fa9_y4, h_s_dadda_rca32_fa8_y4, h_s_dadda_rca32_fa7_y4, h_s_dadda_rca32_fa10_y2, h_s_dadda_rca32_fa10_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_2_y0(a_31, b_2, h_s_dadda_rca32_nand_31_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_3_y0(a_30, b_3, h_s_dadda_rca32_and_30_3_y0);
  fa fa_h_s_dadda_rca32_fa11_y2(h_s_dadda_rca32_fa6_y4, h_s_dadda_rca32_nand_31_2_y0, h_s_dadda_rca32_and_30_3_y0, h_s_dadda_rca32_fa11_y2, h_s_dadda_rca32_fa11_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_4_y0(a_29, b_4, h_s_dadda_rca32_and_29_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_5_y0(a_28, b_5, h_s_dadda_rca32_and_28_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_6_y0(a_27, b_6, h_s_dadda_rca32_and_27_6_y0);
  fa fa_h_s_dadda_rca32_fa12_y2(h_s_dadda_rca32_and_29_4_y0, h_s_dadda_rca32_and_28_5_y0, h_s_dadda_rca32_and_27_6_y0, h_s_dadda_rca32_fa12_y2, h_s_dadda_rca32_fa12_y4);
  fa fa_h_s_dadda_rca32_fa13_y2(h_s_dadda_rca32_fa12_y4, h_s_dadda_rca32_fa11_y4, h_s_dadda_rca32_fa10_y4, h_s_dadda_rca32_fa13_y2, h_s_dadda_rca32_fa13_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_3_y0(a_31, b_3, h_s_dadda_rca32_nand_31_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_4_y0(a_30, b_4, h_s_dadda_rca32_and_30_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_5_y0(a_29, b_5, h_s_dadda_rca32_and_29_5_y0);
  fa fa_h_s_dadda_rca32_fa14_y2(h_s_dadda_rca32_nand_31_3_y0, h_s_dadda_rca32_and_30_4_y0, h_s_dadda_rca32_and_29_5_y0, h_s_dadda_rca32_fa14_y2, h_s_dadda_rca32_fa14_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_4_y0(a_31, b_4, h_s_dadda_rca32_nand_31_4_y0);
  fa fa_h_s_dadda_rca32_fa15_y2(h_s_dadda_rca32_fa14_y4, h_s_dadda_rca32_fa13_y4, h_s_dadda_rca32_nand_31_4_y0, h_s_dadda_rca32_fa15_y2, h_s_dadda_rca32_fa15_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_0_y0(a_6, b_0, h_s_dadda_rca32_and_6_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_1_y0(a_5, b_1, h_s_dadda_rca32_and_5_1_y0);
  ha ha_h_s_dadda_rca32_ha4_y0(h_s_dadda_rca32_and_6_0_y0, h_s_dadda_rca32_and_5_1_y0, h_s_dadda_rca32_ha4_y0, h_s_dadda_rca32_ha4_y1);
  and_gate and_gate_h_s_dadda_rca32_and_7_0_y0(a_7, b_0, h_s_dadda_rca32_and_7_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_1_y0(a_6, b_1, h_s_dadda_rca32_and_6_1_y0);
  fa fa_h_s_dadda_rca32_fa16_y2(h_s_dadda_rca32_ha4_y1, h_s_dadda_rca32_and_7_0_y0, h_s_dadda_rca32_and_6_1_y0, h_s_dadda_rca32_fa16_y2, h_s_dadda_rca32_fa16_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_2_y0(a_5, b_2, h_s_dadda_rca32_and_5_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_3_y0(a_4, b_3, h_s_dadda_rca32_and_4_3_y0);
  ha ha_h_s_dadda_rca32_ha5_y0(h_s_dadda_rca32_and_5_2_y0, h_s_dadda_rca32_and_4_3_y0, h_s_dadda_rca32_ha5_y0, h_s_dadda_rca32_ha5_y1);
  and_gate and_gate_h_s_dadda_rca32_and_8_0_y0(a_8, b_0, h_s_dadda_rca32_and_8_0_y0);
  fa fa_h_s_dadda_rca32_fa17_y2(h_s_dadda_rca32_ha5_y1, h_s_dadda_rca32_fa16_y4, h_s_dadda_rca32_and_8_0_y0, h_s_dadda_rca32_fa17_y2, h_s_dadda_rca32_fa17_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_1_y0(a_7, b_1, h_s_dadda_rca32_and_7_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_2_y0(a_6, b_2, h_s_dadda_rca32_and_6_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_3_y0(a_5, b_3, h_s_dadda_rca32_and_5_3_y0);
  fa fa_h_s_dadda_rca32_fa18_y2(h_s_dadda_rca32_and_7_1_y0, h_s_dadda_rca32_and_6_2_y0, h_s_dadda_rca32_and_5_3_y0, h_s_dadda_rca32_fa18_y2, h_s_dadda_rca32_fa18_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_4_y0(a_4, b_4, h_s_dadda_rca32_and_4_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_5_y0(a_3, b_5, h_s_dadda_rca32_and_3_5_y0);
  ha ha_h_s_dadda_rca32_ha6_y0(h_s_dadda_rca32_and_4_4_y0, h_s_dadda_rca32_and_3_5_y0, h_s_dadda_rca32_ha6_y0, h_s_dadda_rca32_ha6_y1);
  fa fa_h_s_dadda_rca32_fa19_y2(h_s_dadda_rca32_ha6_y1, h_s_dadda_rca32_fa18_y4, h_s_dadda_rca32_fa17_y4, h_s_dadda_rca32_fa19_y2, h_s_dadda_rca32_fa19_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_0_y0(a_9, b_0, h_s_dadda_rca32_and_9_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_1_y0(a_8, b_1, h_s_dadda_rca32_and_8_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_2_y0(a_7, b_2, h_s_dadda_rca32_and_7_2_y0);
  fa fa_h_s_dadda_rca32_fa20_y2(h_s_dadda_rca32_and_9_0_y0, h_s_dadda_rca32_and_8_1_y0, h_s_dadda_rca32_and_7_2_y0, h_s_dadda_rca32_fa20_y2, h_s_dadda_rca32_fa20_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_3_y0(a_6, b_3, h_s_dadda_rca32_and_6_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_4_y0(a_5, b_4, h_s_dadda_rca32_and_5_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_5_y0(a_4, b_5, h_s_dadda_rca32_and_4_5_y0);
  fa fa_h_s_dadda_rca32_fa21_y2(h_s_dadda_rca32_and_6_3_y0, h_s_dadda_rca32_and_5_4_y0, h_s_dadda_rca32_and_4_5_y0, h_s_dadda_rca32_fa21_y2, h_s_dadda_rca32_fa21_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_6_y0(a_3, b_6, h_s_dadda_rca32_and_3_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_7_y0(a_2, b_7, h_s_dadda_rca32_and_2_7_y0);
  ha ha_h_s_dadda_rca32_ha7_y0(h_s_dadda_rca32_and_3_6_y0, h_s_dadda_rca32_and_2_7_y0, h_s_dadda_rca32_ha7_y0, h_s_dadda_rca32_ha7_y1);
  fa fa_h_s_dadda_rca32_fa22_y2(h_s_dadda_rca32_ha7_y1, h_s_dadda_rca32_fa21_y4, h_s_dadda_rca32_fa20_y4, h_s_dadda_rca32_fa22_y2, h_s_dadda_rca32_fa22_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_0_y0(a_10, b_0, h_s_dadda_rca32_and_10_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_1_y0(a_9, b_1, h_s_dadda_rca32_and_9_1_y0);
  fa fa_h_s_dadda_rca32_fa23_y2(h_s_dadda_rca32_fa19_y4, h_s_dadda_rca32_and_10_0_y0, h_s_dadda_rca32_and_9_1_y0, h_s_dadda_rca32_fa23_y2, h_s_dadda_rca32_fa23_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_2_y0(a_8, b_2, h_s_dadda_rca32_and_8_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_3_y0(a_7, b_3, h_s_dadda_rca32_and_7_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_4_y0(a_6, b_4, h_s_dadda_rca32_and_6_4_y0);
  fa fa_h_s_dadda_rca32_fa24_y2(h_s_dadda_rca32_and_8_2_y0, h_s_dadda_rca32_and_7_3_y0, h_s_dadda_rca32_and_6_4_y0, h_s_dadda_rca32_fa24_y2, h_s_dadda_rca32_fa24_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_5_y0(a_5, b_5, h_s_dadda_rca32_and_5_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_6_y0(a_4, b_6, h_s_dadda_rca32_and_4_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_7_y0(a_3, b_7, h_s_dadda_rca32_and_3_7_y0);
  fa fa_h_s_dadda_rca32_fa25_y2(h_s_dadda_rca32_and_5_5_y0, h_s_dadda_rca32_and_4_6_y0, h_s_dadda_rca32_and_3_7_y0, h_s_dadda_rca32_fa25_y2, h_s_dadda_rca32_fa25_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_8_y0(a_2, b_8, h_s_dadda_rca32_and_2_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_9_y0(a_1, b_9, h_s_dadda_rca32_and_1_9_y0);
  ha ha_h_s_dadda_rca32_ha8_y0(h_s_dadda_rca32_and_2_8_y0, h_s_dadda_rca32_and_1_9_y0, h_s_dadda_rca32_ha8_y0, h_s_dadda_rca32_ha8_y1);
  fa fa_h_s_dadda_rca32_fa26_y2(h_s_dadda_rca32_ha8_y1, h_s_dadda_rca32_fa25_y4, h_s_dadda_rca32_fa24_y4, h_s_dadda_rca32_fa26_y2, h_s_dadda_rca32_fa26_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_0_y0(a_11, b_0, h_s_dadda_rca32_and_11_0_y0);
  fa fa_h_s_dadda_rca32_fa27_y2(h_s_dadda_rca32_fa23_y4, h_s_dadda_rca32_fa22_y4, h_s_dadda_rca32_and_11_0_y0, h_s_dadda_rca32_fa27_y2, h_s_dadda_rca32_fa27_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_1_y0(a_10, b_1, h_s_dadda_rca32_and_10_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_2_y0(a_9, b_2, h_s_dadda_rca32_and_9_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_3_y0(a_8, b_3, h_s_dadda_rca32_and_8_3_y0);
  fa fa_h_s_dadda_rca32_fa28_y2(h_s_dadda_rca32_and_10_1_y0, h_s_dadda_rca32_and_9_2_y0, h_s_dadda_rca32_and_8_3_y0, h_s_dadda_rca32_fa28_y2, h_s_dadda_rca32_fa28_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_4_y0(a_7, b_4, h_s_dadda_rca32_and_7_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_5_y0(a_6, b_5, h_s_dadda_rca32_and_6_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_6_y0(a_5, b_6, h_s_dadda_rca32_and_5_6_y0);
  fa fa_h_s_dadda_rca32_fa29_y2(h_s_dadda_rca32_and_7_4_y0, h_s_dadda_rca32_and_6_5_y0, h_s_dadda_rca32_and_5_6_y0, h_s_dadda_rca32_fa29_y2, h_s_dadda_rca32_fa29_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_7_y0(a_4, b_7, h_s_dadda_rca32_and_4_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_8_y0(a_3, b_8, h_s_dadda_rca32_and_3_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_9_y0(a_2, b_9, h_s_dadda_rca32_and_2_9_y0);
  fa fa_h_s_dadda_rca32_fa30_y2(h_s_dadda_rca32_and_4_7_y0, h_s_dadda_rca32_and_3_8_y0, h_s_dadda_rca32_and_2_9_y0, h_s_dadda_rca32_fa30_y2, h_s_dadda_rca32_fa30_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_10_y0(a_1, b_10, h_s_dadda_rca32_and_1_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_11_y0(a_0, b_11, h_s_dadda_rca32_and_0_11_y0);
  ha ha_h_s_dadda_rca32_ha9_y0(h_s_dadda_rca32_and_1_10_y0, h_s_dadda_rca32_and_0_11_y0, h_s_dadda_rca32_ha9_y0, h_s_dadda_rca32_ha9_y1);
  fa fa_h_s_dadda_rca32_fa31_y2(h_s_dadda_rca32_ha9_y1, h_s_dadda_rca32_fa30_y4, h_s_dadda_rca32_fa29_y4, h_s_dadda_rca32_fa31_y2, h_s_dadda_rca32_fa31_y4);
  fa fa_h_s_dadda_rca32_fa32_y2(h_s_dadda_rca32_fa28_y4, h_s_dadda_rca32_fa27_y4, h_s_dadda_rca32_fa26_y4, h_s_dadda_rca32_fa32_y2, h_s_dadda_rca32_fa32_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_0_y0(a_12, b_0, h_s_dadda_rca32_and_12_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_1_y0(a_11, b_1, h_s_dadda_rca32_and_11_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_2_y0(a_10, b_2, h_s_dadda_rca32_and_10_2_y0);
  fa fa_h_s_dadda_rca32_fa33_y2(h_s_dadda_rca32_and_12_0_y0, h_s_dadda_rca32_and_11_1_y0, h_s_dadda_rca32_and_10_2_y0, h_s_dadda_rca32_fa33_y2, h_s_dadda_rca32_fa33_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_3_y0(a_9, b_3, h_s_dadda_rca32_and_9_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_4_y0(a_8, b_4, h_s_dadda_rca32_and_8_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_5_y0(a_7, b_5, h_s_dadda_rca32_and_7_5_y0);
  fa fa_h_s_dadda_rca32_fa34_y2(h_s_dadda_rca32_and_9_3_y0, h_s_dadda_rca32_and_8_4_y0, h_s_dadda_rca32_and_7_5_y0, h_s_dadda_rca32_fa34_y2, h_s_dadda_rca32_fa34_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_6_y0(a_6, b_6, h_s_dadda_rca32_and_6_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_7_y0(a_5, b_7, h_s_dadda_rca32_and_5_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_8_y0(a_4, b_8, h_s_dadda_rca32_and_4_8_y0);
  fa fa_h_s_dadda_rca32_fa35_y2(h_s_dadda_rca32_and_6_6_y0, h_s_dadda_rca32_and_5_7_y0, h_s_dadda_rca32_and_4_8_y0, h_s_dadda_rca32_fa35_y2, h_s_dadda_rca32_fa35_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_9_y0(a_3, b_9, h_s_dadda_rca32_and_3_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_10_y0(a_2, b_10, h_s_dadda_rca32_and_2_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_11_y0(a_1, b_11, h_s_dadda_rca32_and_1_11_y0);
  fa fa_h_s_dadda_rca32_fa36_y2(h_s_dadda_rca32_and_3_9_y0, h_s_dadda_rca32_and_2_10_y0, h_s_dadda_rca32_and_1_11_y0, h_s_dadda_rca32_fa36_y2, h_s_dadda_rca32_fa36_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_12_y0(a_0, b_12, h_s_dadda_rca32_and_0_12_y0);
  ha ha_h_s_dadda_rca32_ha10_y0(h_s_dadda_rca32_and_0_12_y0, h_s_dadda_rca32_fa31_y2, h_s_dadda_rca32_ha10_y0, h_s_dadda_rca32_ha10_y1);
  fa fa_h_s_dadda_rca32_fa37_y2(h_s_dadda_rca32_ha10_y1, h_s_dadda_rca32_fa36_y4, h_s_dadda_rca32_fa35_y4, h_s_dadda_rca32_fa37_y2, h_s_dadda_rca32_fa37_y4);
  fa fa_h_s_dadda_rca32_fa38_y2(h_s_dadda_rca32_fa34_y4, h_s_dadda_rca32_fa33_y4, h_s_dadda_rca32_fa32_y4, h_s_dadda_rca32_fa38_y2, h_s_dadda_rca32_fa38_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_0_y0(a_13, b_0, h_s_dadda_rca32_and_13_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_1_y0(a_12, b_1, h_s_dadda_rca32_and_12_1_y0);
  fa fa_h_s_dadda_rca32_fa39_y2(h_s_dadda_rca32_fa31_y4, h_s_dadda_rca32_and_13_0_y0, h_s_dadda_rca32_and_12_1_y0, h_s_dadda_rca32_fa39_y2, h_s_dadda_rca32_fa39_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_2_y0(a_11, b_2, h_s_dadda_rca32_and_11_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_3_y0(a_10, b_3, h_s_dadda_rca32_and_10_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_4_y0(a_9, b_4, h_s_dadda_rca32_and_9_4_y0);
  fa fa_h_s_dadda_rca32_fa40_y2(h_s_dadda_rca32_and_11_2_y0, h_s_dadda_rca32_and_10_3_y0, h_s_dadda_rca32_and_9_4_y0, h_s_dadda_rca32_fa40_y2, h_s_dadda_rca32_fa40_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_5_y0(a_8, b_5, h_s_dadda_rca32_and_8_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_6_y0(a_7, b_6, h_s_dadda_rca32_and_7_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_7_y0(a_6, b_7, h_s_dadda_rca32_and_6_7_y0);
  fa fa_h_s_dadda_rca32_fa41_y2(h_s_dadda_rca32_and_8_5_y0, h_s_dadda_rca32_and_7_6_y0, h_s_dadda_rca32_and_6_7_y0, h_s_dadda_rca32_fa41_y2, h_s_dadda_rca32_fa41_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_8_y0(a_5, b_8, h_s_dadda_rca32_and_5_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_9_y0(a_4, b_9, h_s_dadda_rca32_and_4_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_10_y0(a_3, b_10, h_s_dadda_rca32_and_3_10_y0);
  fa fa_h_s_dadda_rca32_fa42_y2(h_s_dadda_rca32_and_5_8_y0, h_s_dadda_rca32_and_4_9_y0, h_s_dadda_rca32_and_3_10_y0, h_s_dadda_rca32_fa42_y2, h_s_dadda_rca32_fa42_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_11_y0(a_2, b_11, h_s_dadda_rca32_and_2_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_12_y0(a_1, b_12, h_s_dadda_rca32_and_1_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_13_y0(a_0, b_13, h_s_dadda_rca32_and_0_13_y0);
  fa fa_h_s_dadda_rca32_fa43_y2(h_s_dadda_rca32_and_2_11_y0, h_s_dadda_rca32_and_1_12_y0, h_s_dadda_rca32_and_0_13_y0, h_s_dadda_rca32_fa43_y2, h_s_dadda_rca32_fa43_y4);
  ha ha_h_s_dadda_rca32_ha11_y0(h_s_dadda_rca32_fa37_y2, h_s_dadda_rca32_fa38_y2, h_s_dadda_rca32_ha11_y0, h_s_dadda_rca32_ha11_y1);
  fa fa_h_s_dadda_rca32_fa44_y2(h_s_dadda_rca32_ha11_y1, h_s_dadda_rca32_fa43_y4, h_s_dadda_rca32_fa42_y4, h_s_dadda_rca32_fa44_y2, h_s_dadda_rca32_fa44_y4);
  fa fa_h_s_dadda_rca32_fa45_y2(h_s_dadda_rca32_fa41_y4, h_s_dadda_rca32_fa40_y4, h_s_dadda_rca32_fa39_y4, h_s_dadda_rca32_fa45_y2, h_s_dadda_rca32_fa45_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_0_y0(a_14, b_0, h_s_dadda_rca32_and_14_0_y0);
  fa fa_h_s_dadda_rca32_fa46_y2(h_s_dadda_rca32_fa38_y4, h_s_dadda_rca32_fa37_y4, h_s_dadda_rca32_and_14_0_y0, h_s_dadda_rca32_fa46_y2, h_s_dadda_rca32_fa46_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_1_y0(a_13, b_1, h_s_dadda_rca32_and_13_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_2_y0(a_12, b_2, h_s_dadda_rca32_and_12_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_3_y0(a_11, b_3, h_s_dadda_rca32_and_11_3_y0);
  fa fa_h_s_dadda_rca32_fa47_y2(h_s_dadda_rca32_and_13_1_y0, h_s_dadda_rca32_and_12_2_y0, h_s_dadda_rca32_and_11_3_y0, h_s_dadda_rca32_fa47_y2, h_s_dadda_rca32_fa47_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_4_y0(a_10, b_4, h_s_dadda_rca32_and_10_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_5_y0(a_9, b_5, h_s_dadda_rca32_and_9_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_6_y0(a_8, b_6, h_s_dadda_rca32_and_8_6_y0);
  fa fa_h_s_dadda_rca32_fa48_y2(h_s_dadda_rca32_and_10_4_y0, h_s_dadda_rca32_and_9_5_y0, h_s_dadda_rca32_and_8_6_y0, h_s_dadda_rca32_fa48_y2, h_s_dadda_rca32_fa48_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_7_y0(a_7, b_7, h_s_dadda_rca32_and_7_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_8_y0(a_6, b_8, h_s_dadda_rca32_and_6_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_9_y0(a_5, b_9, h_s_dadda_rca32_and_5_9_y0);
  fa fa_h_s_dadda_rca32_fa49_y2(h_s_dadda_rca32_and_7_7_y0, h_s_dadda_rca32_and_6_8_y0, h_s_dadda_rca32_and_5_9_y0, h_s_dadda_rca32_fa49_y2, h_s_dadda_rca32_fa49_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_10_y0(a_4, b_10, h_s_dadda_rca32_and_4_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_11_y0(a_3, b_11, h_s_dadda_rca32_and_3_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_12_y0(a_2, b_12, h_s_dadda_rca32_and_2_12_y0);
  fa fa_h_s_dadda_rca32_fa50_y2(h_s_dadda_rca32_and_4_10_y0, h_s_dadda_rca32_and_3_11_y0, h_s_dadda_rca32_and_2_12_y0, h_s_dadda_rca32_fa50_y2, h_s_dadda_rca32_fa50_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_13_y0(a_1, b_13, h_s_dadda_rca32_and_1_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_14_y0(a_0, b_14, h_s_dadda_rca32_and_0_14_y0);
  fa fa_h_s_dadda_rca32_fa51_y2(h_s_dadda_rca32_and_1_13_y0, h_s_dadda_rca32_and_0_14_y0, h_s_dadda_rca32_fa44_y2, h_s_dadda_rca32_fa51_y2, h_s_dadda_rca32_fa51_y4);
  ha ha_h_s_dadda_rca32_ha12_y0(h_s_dadda_rca32_fa45_y2, h_s_dadda_rca32_fa46_y2, h_s_dadda_rca32_ha12_y0, h_s_dadda_rca32_ha12_y1);
  fa fa_h_s_dadda_rca32_fa52_y2(h_s_dadda_rca32_ha12_y1, h_s_dadda_rca32_fa51_y4, h_s_dadda_rca32_fa50_y4, h_s_dadda_rca32_fa52_y2, h_s_dadda_rca32_fa52_y4);
  fa fa_h_s_dadda_rca32_fa53_y2(h_s_dadda_rca32_fa49_y4, h_s_dadda_rca32_fa48_y4, h_s_dadda_rca32_fa47_y4, h_s_dadda_rca32_fa53_y2, h_s_dadda_rca32_fa53_y4);
  fa fa_h_s_dadda_rca32_fa54_y2(h_s_dadda_rca32_fa46_y4, h_s_dadda_rca32_fa45_y4, h_s_dadda_rca32_fa44_y4, h_s_dadda_rca32_fa54_y2, h_s_dadda_rca32_fa54_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_0_y0(a_15, b_0, h_s_dadda_rca32_and_15_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_1_y0(a_14, b_1, h_s_dadda_rca32_and_14_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_2_y0(a_13, b_2, h_s_dadda_rca32_and_13_2_y0);
  fa fa_h_s_dadda_rca32_fa55_y2(h_s_dadda_rca32_and_15_0_y0, h_s_dadda_rca32_and_14_1_y0, h_s_dadda_rca32_and_13_2_y0, h_s_dadda_rca32_fa55_y2, h_s_dadda_rca32_fa55_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_3_y0(a_12, b_3, h_s_dadda_rca32_and_12_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_4_y0(a_11, b_4, h_s_dadda_rca32_and_11_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_5_y0(a_10, b_5, h_s_dadda_rca32_and_10_5_y0);
  fa fa_h_s_dadda_rca32_fa56_y2(h_s_dadda_rca32_and_12_3_y0, h_s_dadda_rca32_and_11_4_y0, h_s_dadda_rca32_and_10_5_y0, h_s_dadda_rca32_fa56_y2, h_s_dadda_rca32_fa56_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_6_y0(a_9, b_6, h_s_dadda_rca32_and_9_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_7_y0(a_8, b_7, h_s_dadda_rca32_and_8_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_8_y0(a_7, b_8, h_s_dadda_rca32_and_7_8_y0);
  fa fa_h_s_dadda_rca32_fa57_y2(h_s_dadda_rca32_and_9_6_y0, h_s_dadda_rca32_and_8_7_y0, h_s_dadda_rca32_and_7_8_y0, h_s_dadda_rca32_fa57_y2, h_s_dadda_rca32_fa57_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_9_y0(a_6, b_9, h_s_dadda_rca32_and_6_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_10_y0(a_5, b_10, h_s_dadda_rca32_and_5_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_11_y0(a_4, b_11, h_s_dadda_rca32_and_4_11_y0);
  fa fa_h_s_dadda_rca32_fa58_y2(h_s_dadda_rca32_and_6_9_y0, h_s_dadda_rca32_and_5_10_y0, h_s_dadda_rca32_and_4_11_y0, h_s_dadda_rca32_fa58_y2, h_s_dadda_rca32_fa58_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_12_y0(a_3, b_12, h_s_dadda_rca32_and_3_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_13_y0(a_2, b_13, h_s_dadda_rca32_and_2_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_14_y0(a_1, b_14, h_s_dadda_rca32_and_1_14_y0);
  fa fa_h_s_dadda_rca32_fa59_y2(h_s_dadda_rca32_and_3_12_y0, h_s_dadda_rca32_and_2_13_y0, h_s_dadda_rca32_and_1_14_y0, h_s_dadda_rca32_fa59_y2, h_s_dadda_rca32_fa59_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_15_y0(a_0, b_15, h_s_dadda_rca32_and_0_15_y0);
  fa fa_h_s_dadda_rca32_fa60_y2(h_s_dadda_rca32_and_0_15_y0, h_s_dadda_rca32_fa52_y2, h_s_dadda_rca32_fa53_y2, h_s_dadda_rca32_fa60_y2, h_s_dadda_rca32_fa60_y4);
  ha ha_h_s_dadda_rca32_ha13_y0(h_s_dadda_rca32_fa54_y2, h_s_dadda_rca32_fa55_y2, h_s_dadda_rca32_ha13_y0, h_s_dadda_rca32_ha13_y1);
  fa fa_h_s_dadda_rca32_fa61_y2(h_s_dadda_rca32_ha13_y1, h_s_dadda_rca32_fa60_y4, h_s_dadda_rca32_fa59_y4, h_s_dadda_rca32_fa61_y2, h_s_dadda_rca32_fa61_y4);
  fa fa_h_s_dadda_rca32_fa62_y2(h_s_dadda_rca32_fa58_y4, h_s_dadda_rca32_fa57_y4, h_s_dadda_rca32_fa56_y4, h_s_dadda_rca32_fa62_y2, h_s_dadda_rca32_fa62_y4);
  fa fa_h_s_dadda_rca32_fa63_y2(h_s_dadda_rca32_fa55_y4, h_s_dadda_rca32_fa54_y4, h_s_dadda_rca32_fa53_y4, h_s_dadda_rca32_fa63_y2, h_s_dadda_rca32_fa63_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_0_y0(a_16, b_0, h_s_dadda_rca32_and_16_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_1_y0(a_15, b_1, h_s_dadda_rca32_and_15_1_y0);
  fa fa_h_s_dadda_rca32_fa64_y2(h_s_dadda_rca32_fa52_y4, h_s_dadda_rca32_and_16_0_y0, h_s_dadda_rca32_and_15_1_y0, h_s_dadda_rca32_fa64_y2, h_s_dadda_rca32_fa64_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_2_y0(a_14, b_2, h_s_dadda_rca32_and_14_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_3_y0(a_13, b_3, h_s_dadda_rca32_and_13_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_4_y0(a_12, b_4, h_s_dadda_rca32_and_12_4_y0);
  fa fa_h_s_dadda_rca32_fa65_y2(h_s_dadda_rca32_and_14_2_y0, h_s_dadda_rca32_and_13_3_y0, h_s_dadda_rca32_and_12_4_y0, h_s_dadda_rca32_fa65_y2, h_s_dadda_rca32_fa65_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_5_y0(a_11, b_5, h_s_dadda_rca32_and_11_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_6_y0(a_10, b_6, h_s_dadda_rca32_and_10_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_7_y0(a_9, b_7, h_s_dadda_rca32_and_9_7_y0);
  fa fa_h_s_dadda_rca32_fa66_y2(h_s_dadda_rca32_and_11_5_y0, h_s_dadda_rca32_and_10_6_y0, h_s_dadda_rca32_and_9_7_y0, h_s_dadda_rca32_fa66_y2, h_s_dadda_rca32_fa66_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_8_y0(a_8, b_8, h_s_dadda_rca32_and_8_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_9_y0(a_7, b_9, h_s_dadda_rca32_and_7_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_10_y0(a_6, b_10, h_s_dadda_rca32_and_6_10_y0);
  fa fa_h_s_dadda_rca32_fa67_y2(h_s_dadda_rca32_and_8_8_y0, h_s_dadda_rca32_and_7_9_y0, h_s_dadda_rca32_and_6_10_y0, h_s_dadda_rca32_fa67_y2, h_s_dadda_rca32_fa67_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_11_y0(a_5, b_11, h_s_dadda_rca32_and_5_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_12_y0(a_4, b_12, h_s_dadda_rca32_and_4_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_13_y0(a_3, b_13, h_s_dadda_rca32_and_3_13_y0);
  fa fa_h_s_dadda_rca32_fa68_y2(h_s_dadda_rca32_and_5_11_y0, h_s_dadda_rca32_and_4_12_y0, h_s_dadda_rca32_and_3_13_y0, h_s_dadda_rca32_fa68_y2, h_s_dadda_rca32_fa68_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_14_y0(a_2, b_14, h_s_dadda_rca32_and_2_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_15_y0(a_1, b_15, h_s_dadda_rca32_and_1_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_16_y0(a_0, b_16, h_s_dadda_rca32_and_0_16_y0);
  fa fa_h_s_dadda_rca32_fa69_y2(h_s_dadda_rca32_and_2_14_y0, h_s_dadda_rca32_and_1_15_y0, h_s_dadda_rca32_and_0_16_y0, h_s_dadda_rca32_fa69_y2, h_s_dadda_rca32_fa69_y4);
  fa fa_h_s_dadda_rca32_fa70_y2(h_s_dadda_rca32_fa61_y2, h_s_dadda_rca32_fa62_y2, h_s_dadda_rca32_fa63_y2, h_s_dadda_rca32_fa70_y2, h_s_dadda_rca32_fa70_y4);
  ha ha_h_s_dadda_rca32_ha14_y0(h_s_dadda_rca32_fa64_y2, h_s_dadda_rca32_fa65_y2, h_s_dadda_rca32_ha14_y0, h_s_dadda_rca32_ha14_y1);
  fa fa_h_s_dadda_rca32_fa71_y2(h_s_dadda_rca32_ha14_y1, h_s_dadda_rca32_fa70_y4, h_s_dadda_rca32_fa69_y4, h_s_dadda_rca32_fa71_y2, h_s_dadda_rca32_fa71_y4);
  fa fa_h_s_dadda_rca32_fa72_y2(h_s_dadda_rca32_fa68_y4, h_s_dadda_rca32_fa67_y4, h_s_dadda_rca32_fa66_y4, h_s_dadda_rca32_fa72_y2, h_s_dadda_rca32_fa72_y4);
  fa fa_h_s_dadda_rca32_fa73_y2(h_s_dadda_rca32_fa65_y4, h_s_dadda_rca32_fa64_y4, h_s_dadda_rca32_fa63_y4, h_s_dadda_rca32_fa73_y2, h_s_dadda_rca32_fa73_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_0_y0(a_17, b_0, h_s_dadda_rca32_and_17_0_y0);
  fa fa_h_s_dadda_rca32_fa74_y2(h_s_dadda_rca32_fa62_y4, h_s_dadda_rca32_fa61_y4, h_s_dadda_rca32_and_17_0_y0, h_s_dadda_rca32_fa74_y2, h_s_dadda_rca32_fa74_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_1_y0(a_16, b_1, h_s_dadda_rca32_and_16_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_2_y0(a_15, b_2, h_s_dadda_rca32_and_15_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_3_y0(a_14, b_3, h_s_dadda_rca32_and_14_3_y0);
  fa fa_h_s_dadda_rca32_fa75_y2(h_s_dadda_rca32_and_16_1_y0, h_s_dadda_rca32_and_15_2_y0, h_s_dadda_rca32_and_14_3_y0, h_s_dadda_rca32_fa75_y2, h_s_dadda_rca32_fa75_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_4_y0(a_13, b_4, h_s_dadda_rca32_and_13_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_5_y0(a_12, b_5, h_s_dadda_rca32_and_12_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_6_y0(a_11, b_6, h_s_dadda_rca32_and_11_6_y0);
  fa fa_h_s_dadda_rca32_fa76_y2(h_s_dadda_rca32_and_13_4_y0, h_s_dadda_rca32_and_12_5_y0, h_s_dadda_rca32_and_11_6_y0, h_s_dadda_rca32_fa76_y2, h_s_dadda_rca32_fa76_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_7_y0(a_10, b_7, h_s_dadda_rca32_and_10_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_8_y0(a_9, b_8, h_s_dadda_rca32_and_9_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_9_y0(a_8, b_9, h_s_dadda_rca32_and_8_9_y0);
  fa fa_h_s_dadda_rca32_fa77_y2(h_s_dadda_rca32_and_10_7_y0, h_s_dadda_rca32_and_9_8_y0, h_s_dadda_rca32_and_8_9_y0, h_s_dadda_rca32_fa77_y2, h_s_dadda_rca32_fa77_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_10_y0(a_7, b_10, h_s_dadda_rca32_and_7_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_11_y0(a_6, b_11, h_s_dadda_rca32_and_6_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_12_y0(a_5, b_12, h_s_dadda_rca32_and_5_12_y0);
  fa fa_h_s_dadda_rca32_fa78_y2(h_s_dadda_rca32_and_7_10_y0, h_s_dadda_rca32_and_6_11_y0, h_s_dadda_rca32_and_5_12_y0, h_s_dadda_rca32_fa78_y2, h_s_dadda_rca32_fa78_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_13_y0(a_4, b_13, h_s_dadda_rca32_and_4_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_14_y0(a_3, b_14, h_s_dadda_rca32_and_3_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_15_y0(a_2, b_15, h_s_dadda_rca32_and_2_15_y0);
  fa fa_h_s_dadda_rca32_fa79_y2(h_s_dadda_rca32_and_4_13_y0, h_s_dadda_rca32_and_3_14_y0, h_s_dadda_rca32_and_2_15_y0, h_s_dadda_rca32_fa79_y2, h_s_dadda_rca32_fa79_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_16_y0(a_1, b_16, h_s_dadda_rca32_and_1_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_17_y0(a_0, b_17, h_s_dadda_rca32_and_0_17_y0);
  fa fa_h_s_dadda_rca32_fa80_y2(h_s_dadda_rca32_and_1_16_y0, h_s_dadda_rca32_and_0_17_y0, h_s_dadda_rca32_fa71_y2, h_s_dadda_rca32_fa80_y2, h_s_dadda_rca32_fa80_y4);
  fa fa_h_s_dadda_rca32_fa81_y2(h_s_dadda_rca32_fa72_y2, h_s_dadda_rca32_fa73_y2, h_s_dadda_rca32_fa74_y2, h_s_dadda_rca32_fa81_y2, h_s_dadda_rca32_fa81_y4);
  ha ha_h_s_dadda_rca32_ha15_y0(h_s_dadda_rca32_fa75_y2, h_s_dadda_rca32_fa76_y2, h_s_dadda_rca32_ha15_y0, h_s_dadda_rca32_ha15_y1);
  fa fa_h_s_dadda_rca32_fa82_y2(h_s_dadda_rca32_ha15_y1, h_s_dadda_rca32_fa81_y4, h_s_dadda_rca32_fa80_y4, h_s_dadda_rca32_fa82_y2, h_s_dadda_rca32_fa82_y4);
  fa fa_h_s_dadda_rca32_fa83_y2(h_s_dadda_rca32_fa79_y4, h_s_dadda_rca32_fa78_y4, h_s_dadda_rca32_fa77_y4, h_s_dadda_rca32_fa83_y2, h_s_dadda_rca32_fa83_y4);
  fa fa_h_s_dadda_rca32_fa84_y2(h_s_dadda_rca32_fa76_y4, h_s_dadda_rca32_fa75_y4, h_s_dadda_rca32_fa74_y4, h_s_dadda_rca32_fa84_y2, h_s_dadda_rca32_fa84_y4);
  fa fa_h_s_dadda_rca32_fa85_y2(h_s_dadda_rca32_fa73_y4, h_s_dadda_rca32_fa72_y4, h_s_dadda_rca32_fa71_y4, h_s_dadda_rca32_fa85_y2, h_s_dadda_rca32_fa85_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_0_y0(a_18, b_0, h_s_dadda_rca32_and_18_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_1_y0(a_17, b_1, h_s_dadda_rca32_and_17_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_2_y0(a_16, b_2, h_s_dadda_rca32_and_16_2_y0);
  fa fa_h_s_dadda_rca32_fa86_y2(h_s_dadda_rca32_and_18_0_y0, h_s_dadda_rca32_and_17_1_y0, h_s_dadda_rca32_and_16_2_y0, h_s_dadda_rca32_fa86_y2, h_s_dadda_rca32_fa86_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_3_y0(a_15, b_3, h_s_dadda_rca32_and_15_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_4_y0(a_14, b_4, h_s_dadda_rca32_and_14_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_5_y0(a_13, b_5, h_s_dadda_rca32_and_13_5_y0);
  fa fa_h_s_dadda_rca32_fa87_y2(h_s_dadda_rca32_and_15_3_y0, h_s_dadda_rca32_and_14_4_y0, h_s_dadda_rca32_and_13_5_y0, h_s_dadda_rca32_fa87_y2, h_s_dadda_rca32_fa87_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_6_y0(a_12, b_6, h_s_dadda_rca32_and_12_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_7_y0(a_11, b_7, h_s_dadda_rca32_and_11_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_8_y0(a_10, b_8, h_s_dadda_rca32_and_10_8_y0);
  fa fa_h_s_dadda_rca32_fa88_y2(h_s_dadda_rca32_and_12_6_y0, h_s_dadda_rca32_and_11_7_y0, h_s_dadda_rca32_and_10_8_y0, h_s_dadda_rca32_fa88_y2, h_s_dadda_rca32_fa88_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_9_y0(a_9, b_9, h_s_dadda_rca32_and_9_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_10_y0(a_8, b_10, h_s_dadda_rca32_and_8_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_11_y0(a_7, b_11, h_s_dadda_rca32_and_7_11_y0);
  fa fa_h_s_dadda_rca32_fa89_y2(h_s_dadda_rca32_and_9_9_y0, h_s_dadda_rca32_and_8_10_y0, h_s_dadda_rca32_and_7_11_y0, h_s_dadda_rca32_fa89_y2, h_s_dadda_rca32_fa89_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_12_y0(a_6, b_12, h_s_dadda_rca32_and_6_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_13_y0(a_5, b_13, h_s_dadda_rca32_and_5_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_14_y0(a_4, b_14, h_s_dadda_rca32_and_4_14_y0);
  fa fa_h_s_dadda_rca32_fa90_y2(h_s_dadda_rca32_and_6_12_y0, h_s_dadda_rca32_and_5_13_y0, h_s_dadda_rca32_and_4_14_y0, h_s_dadda_rca32_fa90_y2, h_s_dadda_rca32_fa90_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_15_y0(a_3, b_15, h_s_dadda_rca32_and_3_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_16_y0(a_2, b_16, h_s_dadda_rca32_and_2_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_17_y0(a_1, b_17, h_s_dadda_rca32_and_1_17_y0);
  fa fa_h_s_dadda_rca32_fa91_y2(h_s_dadda_rca32_and_3_15_y0, h_s_dadda_rca32_and_2_16_y0, h_s_dadda_rca32_and_1_17_y0, h_s_dadda_rca32_fa91_y2, h_s_dadda_rca32_fa91_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_18_y0(a_0, b_18, h_s_dadda_rca32_and_0_18_y0);
  fa fa_h_s_dadda_rca32_fa92_y2(h_s_dadda_rca32_and_0_18_y0, h_s_dadda_rca32_fa82_y2, h_s_dadda_rca32_fa83_y2, h_s_dadda_rca32_fa92_y2, h_s_dadda_rca32_fa92_y4);
  fa fa_h_s_dadda_rca32_fa93_y2(h_s_dadda_rca32_fa84_y2, h_s_dadda_rca32_fa85_y2, h_s_dadda_rca32_fa86_y2, h_s_dadda_rca32_fa93_y2, h_s_dadda_rca32_fa93_y4);
  ha ha_h_s_dadda_rca32_ha16_y0(h_s_dadda_rca32_fa87_y2, h_s_dadda_rca32_fa88_y2, h_s_dadda_rca32_ha16_y0, h_s_dadda_rca32_ha16_y1);
  fa fa_h_s_dadda_rca32_fa94_y2(h_s_dadda_rca32_ha16_y1, h_s_dadda_rca32_fa93_y4, h_s_dadda_rca32_fa92_y4, h_s_dadda_rca32_fa94_y2, h_s_dadda_rca32_fa94_y4);
  fa fa_h_s_dadda_rca32_fa95_y2(h_s_dadda_rca32_fa91_y4, h_s_dadda_rca32_fa90_y4, h_s_dadda_rca32_fa89_y4, h_s_dadda_rca32_fa95_y2, h_s_dadda_rca32_fa95_y4);
  fa fa_h_s_dadda_rca32_fa96_y2(h_s_dadda_rca32_fa88_y4, h_s_dadda_rca32_fa87_y4, h_s_dadda_rca32_fa86_y4, h_s_dadda_rca32_fa96_y2, h_s_dadda_rca32_fa96_y4);
  fa fa_h_s_dadda_rca32_fa97_y2(h_s_dadda_rca32_fa85_y4, h_s_dadda_rca32_fa84_y4, h_s_dadda_rca32_fa83_y4, h_s_dadda_rca32_fa97_y2, h_s_dadda_rca32_fa97_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_0_y0(a_19, b_0, h_s_dadda_rca32_and_19_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_1_y0(a_18, b_1, h_s_dadda_rca32_and_18_1_y0);
  fa fa_h_s_dadda_rca32_fa98_y2(h_s_dadda_rca32_fa82_y4, h_s_dadda_rca32_and_19_0_y0, h_s_dadda_rca32_and_18_1_y0, h_s_dadda_rca32_fa98_y2, h_s_dadda_rca32_fa98_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_2_y0(a_17, b_2, h_s_dadda_rca32_and_17_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_3_y0(a_16, b_3, h_s_dadda_rca32_and_16_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_4_y0(a_15, b_4, h_s_dadda_rca32_and_15_4_y0);
  fa fa_h_s_dadda_rca32_fa99_y2(h_s_dadda_rca32_and_17_2_y0, h_s_dadda_rca32_and_16_3_y0, h_s_dadda_rca32_and_15_4_y0, h_s_dadda_rca32_fa99_y2, h_s_dadda_rca32_fa99_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_5_y0(a_14, b_5, h_s_dadda_rca32_and_14_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_6_y0(a_13, b_6, h_s_dadda_rca32_and_13_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_7_y0(a_12, b_7, h_s_dadda_rca32_and_12_7_y0);
  fa fa_h_s_dadda_rca32_fa100_y2(h_s_dadda_rca32_and_14_5_y0, h_s_dadda_rca32_and_13_6_y0, h_s_dadda_rca32_and_12_7_y0, h_s_dadda_rca32_fa100_y2, h_s_dadda_rca32_fa100_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_8_y0(a_11, b_8, h_s_dadda_rca32_and_11_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_9_y0(a_10, b_9, h_s_dadda_rca32_and_10_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_10_y0(a_9, b_10, h_s_dadda_rca32_and_9_10_y0);
  fa fa_h_s_dadda_rca32_fa101_y2(h_s_dadda_rca32_and_11_8_y0, h_s_dadda_rca32_and_10_9_y0, h_s_dadda_rca32_and_9_10_y0, h_s_dadda_rca32_fa101_y2, h_s_dadda_rca32_fa101_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_11_y0(a_8, b_11, h_s_dadda_rca32_and_8_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_12_y0(a_7, b_12, h_s_dadda_rca32_and_7_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_13_y0(a_6, b_13, h_s_dadda_rca32_and_6_13_y0);
  fa fa_h_s_dadda_rca32_fa102_y2(h_s_dadda_rca32_and_8_11_y0, h_s_dadda_rca32_and_7_12_y0, h_s_dadda_rca32_and_6_13_y0, h_s_dadda_rca32_fa102_y2, h_s_dadda_rca32_fa102_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_14_y0(a_5, b_14, h_s_dadda_rca32_and_5_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_15_y0(a_4, b_15, h_s_dadda_rca32_and_4_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_16_y0(a_3, b_16, h_s_dadda_rca32_and_3_16_y0);
  fa fa_h_s_dadda_rca32_fa103_y2(h_s_dadda_rca32_and_5_14_y0, h_s_dadda_rca32_and_4_15_y0, h_s_dadda_rca32_and_3_16_y0, h_s_dadda_rca32_fa103_y2, h_s_dadda_rca32_fa103_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_17_y0(a_2, b_17, h_s_dadda_rca32_and_2_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_18_y0(a_1, b_18, h_s_dadda_rca32_and_1_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_19_y0(a_0, b_19, h_s_dadda_rca32_and_0_19_y0);
  fa fa_h_s_dadda_rca32_fa104_y2(h_s_dadda_rca32_and_2_17_y0, h_s_dadda_rca32_and_1_18_y0, h_s_dadda_rca32_and_0_19_y0, h_s_dadda_rca32_fa104_y2, h_s_dadda_rca32_fa104_y4);
  fa fa_h_s_dadda_rca32_fa105_y2(h_s_dadda_rca32_fa94_y2, h_s_dadda_rca32_fa95_y2, h_s_dadda_rca32_fa96_y2, h_s_dadda_rca32_fa105_y2, h_s_dadda_rca32_fa105_y4);
  fa fa_h_s_dadda_rca32_fa106_y2(h_s_dadda_rca32_fa97_y2, h_s_dadda_rca32_fa98_y2, h_s_dadda_rca32_fa99_y2, h_s_dadda_rca32_fa106_y2, h_s_dadda_rca32_fa106_y4);
  ha ha_h_s_dadda_rca32_ha17_y0(h_s_dadda_rca32_fa100_y2, h_s_dadda_rca32_fa101_y2, h_s_dadda_rca32_ha17_y0, h_s_dadda_rca32_ha17_y1);
  fa fa_h_s_dadda_rca32_fa107_y2(h_s_dadda_rca32_ha17_y1, h_s_dadda_rca32_fa106_y4, h_s_dadda_rca32_fa105_y4, h_s_dadda_rca32_fa107_y2, h_s_dadda_rca32_fa107_y4);
  fa fa_h_s_dadda_rca32_fa108_y2(h_s_dadda_rca32_fa104_y4, h_s_dadda_rca32_fa103_y4, h_s_dadda_rca32_fa102_y4, h_s_dadda_rca32_fa108_y2, h_s_dadda_rca32_fa108_y4);
  fa fa_h_s_dadda_rca32_fa109_y2(h_s_dadda_rca32_fa101_y4, h_s_dadda_rca32_fa100_y4, h_s_dadda_rca32_fa99_y4, h_s_dadda_rca32_fa109_y2, h_s_dadda_rca32_fa109_y4);
  fa fa_h_s_dadda_rca32_fa110_y2(h_s_dadda_rca32_fa98_y4, h_s_dadda_rca32_fa97_y4, h_s_dadda_rca32_fa96_y4, h_s_dadda_rca32_fa110_y2, h_s_dadda_rca32_fa110_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_0_y0(a_20, b_0, h_s_dadda_rca32_and_20_0_y0);
  fa fa_h_s_dadda_rca32_fa111_y2(h_s_dadda_rca32_fa95_y4, h_s_dadda_rca32_fa94_y4, h_s_dadda_rca32_and_20_0_y0, h_s_dadda_rca32_fa111_y2, h_s_dadda_rca32_fa111_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_1_y0(a_19, b_1, h_s_dadda_rca32_and_19_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_2_y0(a_18, b_2, h_s_dadda_rca32_and_18_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_3_y0(a_17, b_3, h_s_dadda_rca32_and_17_3_y0);
  fa fa_h_s_dadda_rca32_fa112_y2(h_s_dadda_rca32_and_19_1_y0, h_s_dadda_rca32_and_18_2_y0, h_s_dadda_rca32_and_17_3_y0, h_s_dadda_rca32_fa112_y2, h_s_dadda_rca32_fa112_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_4_y0(a_16, b_4, h_s_dadda_rca32_and_16_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_5_y0(a_15, b_5, h_s_dadda_rca32_and_15_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_6_y0(a_14, b_6, h_s_dadda_rca32_and_14_6_y0);
  fa fa_h_s_dadda_rca32_fa113_y2(h_s_dadda_rca32_and_16_4_y0, h_s_dadda_rca32_and_15_5_y0, h_s_dadda_rca32_and_14_6_y0, h_s_dadda_rca32_fa113_y2, h_s_dadda_rca32_fa113_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_7_y0(a_13, b_7, h_s_dadda_rca32_and_13_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_8_y0(a_12, b_8, h_s_dadda_rca32_and_12_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_9_y0(a_11, b_9, h_s_dadda_rca32_and_11_9_y0);
  fa fa_h_s_dadda_rca32_fa114_y2(h_s_dadda_rca32_and_13_7_y0, h_s_dadda_rca32_and_12_8_y0, h_s_dadda_rca32_and_11_9_y0, h_s_dadda_rca32_fa114_y2, h_s_dadda_rca32_fa114_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_10_y0(a_10, b_10, h_s_dadda_rca32_and_10_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_11_y0(a_9, b_11, h_s_dadda_rca32_and_9_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_12_y0(a_8, b_12, h_s_dadda_rca32_and_8_12_y0);
  fa fa_h_s_dadda_rca32_fa115_y2(h_s_dadda_rca32_and_10_10_y0, h_s_dadda_rca32_and_9_11_y0, h_s_dadda_rca32_and_8_12_y0, h_s_dadda_rca32_fa115_y2, h_s_dadda_rca32_fa115_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_13_y0(a_7, b_13, h_s_dadda_rca32_and_7_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_14_y0(a_6, b_14, h_s_dadda_rca32_and_6_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_15_y0(a_5, b_15, h_s_dadda_rca32_and_5_15_y0);
  fa fa_h_s_dadda_rca32_fa116_y2(h_s_dadda_rca32_and_7_13_y0, h_s_dadda_rca32_and_6_14_y0, h_s_dadda_rca32_and_5_15_y0, h_s_dadda_rca32_fa116_y2, h_s_dadda_rca32_fa116_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_16_y0(a_4, b_16, h_s_dadda_rca32_and_4_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_17_y0(a_3, b_17, h_s_dadda_rca32_and_3_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_18_y0(a_2, b_18, h_s_dadda_rca32_and_2_18_y0);
  fa fa_h_s_dadda_rca32_fa117_y2(h_s_dadda_rca32_and_4_16_y0, h_s_dadda_rca32_and_3_17_y0, h_s_dadda_rca32_and_2_18_y0, h_s_dadda_rca32_fa117_y2, h_s_dadda_rca32_fa117_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_19_y0(a_1, b_19, h_s_dadda_rca32_and_1_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_20_y0(a_0, b_20, h_s_dadda_rca32_and_0_20_y0);
  fa fa_h_s_dadda_rca32_fa118_y2(h_s_dadda_rca32_and_1_19_y0, h_s_dadda_rca32_and_0_20_y0, h_s_dadda_rca32_fa107_y2, h_s_dadda_rca32_fa118_y2, h_s_dadda_rca32_fa118_y4);
  fa fa_h_s_dadda_rca32_fa119_y2(h_s_dadda_rca32_fa108_y2, h_s_dadda_rca32_fa109_y2, h_s_dadda_rca32_fa110_y2, h_s_dadda_rca32_fa119_y2, h_s_dadda_rca32_fa119_y4);
  fa fa_h_s_dadda_rca32_fa120_y2(h_s_dadda_rca32_fa111_y2, h_s_dadda_rca32_fa112_y2, h_s_dadda_rca32_fa113_y2, h_s_dadda_rca32_fa120_y2, h_s_dadda_rca32_fa120_y4);
  ha ha_h_s_dadda_rca32_ha18_y0(h_s_dadda_rca32_fa114_y2, h_s_dadda_rca32_fa115_y2, h_s_dadda_rca32_ha18_y0, h_s_dadda_rca32_ha18_y1);
  fa fa_h_s_dadda_rca32_fa121_y2(h_s_dadda_rca32_ha18_y1, h_s_dadda_rca32_fa120_y4, h_s_dadda_rca32_fa119_y4, h_s_dadda_rca32_fa121_y2, h_s_dadda_rca32_fa121_y4);
  fa fa_h_s_dadda_rca32_fa122_y2(h_s_dadda_rca32_fa118_y4, h_s_dadda_rca32_fa117_y4, h_s_dadda_rca32_fa116_y4, h_s_dadda_rca32_fa122_y2, h_s_dadda_rca32_fa122_y4);
  fa fa_h_s_dadda_rca32_fa123_y2(h_s_dadda_rca32_fa115_y4, h_s_dadda_rca32_fa114_y4, h_s_dadda_rca32_fa113_y4, h_s_dadda_rca32_fa123_y2, h_s_dadda_rca32_fa123_y4);
  fa fa_h_s_dadda_rca32_fa124_y2(h_s_dadda_rca32_fa112_y4, h_s_dadda_rca32_fa111_y4, h_s_dadda_rca32_fa110_y4, h_s_dadda_rca32_fa124_y2, h_s_dadda_rca32_fa124_y4);
  fa fa_h_s_dadda_rca32_fa125_y2(h_s_dadda_rca32_fa109_y4, h_s_dadda_rca32_fa108_y4, h_s_dadda_rca32_fa107_y4, h_s_dadda_rca32_fa125_y2, h_s_dadda_rca32_fa125_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_0_y0(a_21, b_0, h_s_dadda_rca32_and_21_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_1_y0(a_20, b_1, h_s_dadda_rca32_and_20_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_2_y0(a_19, b_2, h_s_dadda_rca32_and_19_2_y0);
  fa fa_h_s_dadda_rca32_fa126_y2(h_s_dadda_rca32_and_21_0_y0, h_s_dadda_rca32_and_20_1_y0, h_s_dadda_rca32_and_19_2_y0, h_s_dadda_rca32_fa126_y2, h_s_dadda_rca32_fa126_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_3_y0(a_18, b_3, h_s_dadda_rca32_and_18_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_4_y0(a_17, b_4, h_s_dadda_rca32_and_17_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_5_y0(a_16, b_5, h_s_dadda_rca32_and_16_5_y0);
  fa fa_h_s_dadda_rca32_fa127_y2(h_s_dadda_rca32_and_18_3_y0, h_s_dadda_rca32_and_17_4_y0, h_s_dadda_rca32_and_16_5_y0, h_s_dadda_rca32_fa127_y2, h_s_dadda_rca32_fa127_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_6_y0(a_15, b_6, h_s_dadda_rca32_and_15_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_7_y0(a_14, b_7, h_s_dadda_rca32_and_14_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_8_y0(a_13, b_8, h_s_dadda_rca32_and_13_8_y0);
  fa fa_h_s_dadda_rca32_fa128_y2(h_s_dadda_rca32_and_15_6_y0, h_s_dadda_rca32_and_14_7_y0, h_s_dadda_rca32_and_13_8_y0, h_s_dadda_rca32_fa128_y2, h_s_dadda_rca32_fa128_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_9_y0(a_12, b_9, h_s_dadda_rca32_and_12_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_10_y0(a_11, b_10, h_s_dadda_rca32_and_11_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_11_y0(a_10, b_11, h_s_dadda_rca32_and_10_11_y0);
  fa fa_h_s_dadda_rca32_fa129_y2(h_s_dadda_rca32_and_12_9_y0, h_s_dadda_rca32_and_11_10_y0, h_s_dadda_rca32_and_10_11_y0, h_s_dadda_rca32_fa129_y2, h_s_dadda_rca32_fa129_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_12_y0(a_9, b_12, h_s_dadda_rca32_and_9_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_13_y0(a_8, b_13, h_s_dadda_rca32_and_8_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_14_y0(a_7, b_14, h_s_dadda_rca32_and_7_14_y0);
  fa fa_h_s_dadda_rca32_fa130_y2(h_s_dadda_rca32_and_9_12_y0, h_s_dadda_rca32_and_8_13_y0, h_s_dadda_rca32_and_7_14_y0, h_s_dadda_rca32_fa130_y2, h_s_dadda_rca32_fa130_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_15_y0(a_6, b_15, h_s_dadda_rca32_and_6_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_16_y0(a_5, b_16, h_s_dadda_rca32_and_5_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_17_y0(a_4, b_17, h_s_dadda_rca32_and_4_17_y0);
  fa fa_h_s_dadda_rca32_fa131_y2(h_s_dadda_rca32_and_6_15_y0, h_s_dadda_rca32_and_5_16_y0, h_s_dadda_rca32_and_4_17_y0, h_s_dadda_rca32_fa131_y2, h_s_dadda_rca32_fa131_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_18_y0(a_3, b_18, h_s_dadda_rca32_and_3_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_19_y0(a_2, b_19, h_s_dadda_rca32_and_2_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_20_y0(a_1, b_20, h_s_dadda_rca32_and_1_20_y0);
  fa fa_h_s_dadda_rca32_fa132_y2(h_s_dadda_rca32_and_3_18_y0, h_s_dadda_rca32_and_2_19_y0, h_s_dadda_rca32_and_1_20_y0, h_s_dadda_rca32_fa132_y2, h_s_dadda_rca32_fa132_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_21_y0(a_0, b_21, h_s_dadda_rca32_and_0_21_y0);
  fa fa_h_s_dadda_rca32_fa133_y2(h_s_dadda_rca32_and_0_21_y0, h_s_dadda_rca32_fa121_y2, h_s_dadda_rca32_fa122_y2, h_s_dadda_rca32_fa133_y2, h_s_dadda_rca32_fa133_y4);
  fa fa_h_s_dadda_rca32_fa134_y2(h_s_dadda_rca32_fa123_y2, h_s_dadda_rca32_fa124_y2, h_s_dadda_rca32_fa125_y2, h_s_dadda_rca32_fa134_y2, h_s_dadda_rca32_fa134_y4);
  fa fa_h_s_dadda_rca32_fa135_y2(h_s_dadda_rca32_fa126_y2, h_s_dadda_rca32_fa127_y2, h_s_dadda_rca32_fa128_y2, h_s_dadda_rca32_fa135_y2, h_s_dadda_rca32_fa135_y4);
  ha ha_h_s_dadda_rca32_ha19_y0(h_s_dadda_rca32_fa129_y2, h_s_dadda_rca32_fa130_y2, h_s_dadda_rca32_ha19_y0, h_s_dadda_rca32_ha19_y1);
  fa fa_h_s_dadda_rca32_fa136_y2(h_s_dadda_rca32_ha19_y1, h_s_dadda_rca32_fa135_y4, h_s_dadda_rca32_fa134_y4, h_s_dadda_rca32_fa136_y2, h_s_dadda_rca32_fa136_y4);
  fa fa_h_s_dadda_rca32_fa137_y2(h_s_dadda_rca32_fa133_y4, h_s_dadda_rca32_fa132_y4, h_s_dadda_rca32_fa131_y4, h_s_dadda_rca32_fa137_y2, h_s_dadda_rca32_fa137_y4);
  fa fa_h_s_dadda_rca32_fa138_y2(h_s_dadda_rca32_fa130_y4, h_s_dadda_rca32_fa129_y4, h_s_dadda_rca32_fa128_y4, h_s_dadda_rca32_fa138_y2, h_s_dadda_rca32_fa138_y4);
  fa fa_h_s_dadda_rca32_fa139_y2(h_s_dadda_rca32_fa127_y4, h_s_dadda_rca32_fa126_y4, h_s_dadda_rca32_fa125_y4, h_s_dadda_rca32_fa139_y2, h_s_dadda_rca32_fa139_y4);
  fa fa_h_s_dadda_rca32_fa140_y2(h_s_dadda_rca32_fa124_y4, h_s_dadda_rca32_fa123_y4, h_s_dadda_rca32_fa122_y4, h_s_dadda_rca32_fa140_y2, h_s_dadda_rca32_fa140_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_0_y0(a_22, b_0, h_s_dadda_rca32_and_22_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_1_y0(a_21, b_1, h_s_dadda_rca32_and_21_1_y0);
  fa fa_h_s_dadda_rca32_fa141_y2(h_s_dadda_rca32_fa121_y4, h_s_dadda_rca32_and_22_0_y0, h_s_dadda_rca32_and_21_1_y0, h_s_dadda_rca32_fa141_y2, h_s_dadda_rca32_fa141_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_2_y0(a_20, b_2, h_s_dadda_rca32_and_20_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_3_y0(a_19, b_3, h_s_dadda_rca32_and_19_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_4_y0(a_18, b_4, h_s_dadda_rca32_and_18_4_y0);
  fa fa_h_s_dadda_rca32_fa142_y2(h_s_dadda_rca32_and_20_2_y0, h_s_dadda_rca32_and_19_3_y0, h_s_dadda_rca32_and_18_4_y0, h_s_dadda_rca32_fa142_y2, h_s_dadda_rca32_fa142_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_5_y0(a_17, b_5, h_s_dadda_rca32_and_17_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_6_y0(a_16, b_6, h_s_dadda_rca32_and_16_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_7_y0(a_15, b_7, h_s_dadda_rca32_and_15_7_y0);
  fa fa_h_s_dadda_rca32_fa143_y2(h_s_dadda_rca32_and_17_5_y0, h_s_dadda_rca32_and_16_6_y0, h_s_dadda_rca32_and_15_7_y0, h_s_dadda_rca32_fa143_y2, h_s_dadda_rca32_fa143_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_8_y0(a_14, b_8, h_s_dadda_rca32_and_14_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_9_y0(a_13, b_9, h_s_dadda_rca32_and_13_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_10_y0(a_12, b_10, h_s_dadda_rca32_and_12_10_y0);
  fa fa_h_s_dadda_rca32_fa144_y2(h_s_dadda_rca32_and_14_8_y0, h_s_dadda_rca32_and_13_9_y0, h_s_dadda_rca32_and_12_10_y0, h_s_dadda_rca32_fa144_y2, h_s_dadda_rca32_fa144_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_11_y0(a_11, b_11, h_s_dadda_rca32_and_11_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_12_y0(a_10, b_12, h_s_dadda_rca32_and_10_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_13_y0(a_9, b_13, h_s_dadda_rca32_and_9_13_y0);
  fa fa_h_s_dadda_rca32_fa145_y2(h_s_dadda_rca32_and_11_11_y0, h_s_dadda_rca32_and_10_12_y0, h_s_dadda_rca32_and_9_13_y0, h_s_dadda_rca32_fa145_y2, h_s_dadda_rca32_fa145_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_14_y0(a_8, b_14, h_s_dadda_rca32_and_8_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_15_y0(a_7, b_15, h_s_dadda_rca32_and_7_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_16_y0(a_6, b_16, h_s_dadda_rca32_and_6_16_y0);
  fa fa_h_s_dadda_rca32_fa146_y2(h_s_dadda_rca32_and_8_14_y0, h_s_dadda_rca32_and_7_15_y0, h_s_dadda_rca32_and_6_16_y0, h_s_dadda_rca32_fa146_y2, h_s_dadda_rca32_fa146_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_17_y0(a_5, b_17, h_s_dadda_rca32_and_5_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_18_y0(a_4, b_18, h_s_dadda_rca32_and_4_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_19_y0(a_3, b_19, h_s_dadda_rca32_and_3_19_y0);
  fa fa_h_s_dadda_rca32_fa147_y2(h_s_dadda_rca32_and_5_17_y0, h_s_dadda_rca32_and_4_18_y0, h_s_dadda_rca32_and_3_19_y0, h_s_dadda_rca32_fa147_y2, h_s_dadda_rca32_fa147_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_20_y0(a_2, b_20, h_s_dadda_rca32_and_2_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_21_y0(a_1, b_21, h_s_dadda_rca32_and_1_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_22_y0(a_0, b_22, h_s_dadda_rca32_and_0_22_y0);
  fa fa_h_s_dadda_rca32_fa148_y2(h_s_dadda_rca32_and_2_20_y0, h_s_dadda_rca32_and_1_21_y0, h_s_dadda_rca32_and_0_22_y0, h_s_dadda_rca32_fa148_y2, h_s_dadda_rca32_fa148_y4);
  fa fa_h_s_dadda_rca32_fa149_y2(h_s_dadda_rca32_fa136_y2, h_s_dadda_rca32_fa137_y2, h_s_dadda_rca32_fa138_y2, h_s_dadda_rca32_fa149_y2, h_s_dadda_rca32_fa149_y4);
  fa fa_h_s_dadda_rca32_fa150_y2(h_s_dadda_rca32_fa139_y2, h_s_dadda_rca32_fa140_y2, h_s_dadda_rca32_fa141_y2, h_s_dadda_rca32_fa150_y2, h_s_dadda_rca32_fa150_y4);
  fa fa_h_s_dadda_rca32_fa151_y2(h_s_dadda_rca32_fa142_y2, h_s_dadda_rca32_fa143_y2, h_s_dadda_rca32_fa144_y2, h_s_dadda_rca32_fa151_y2, h_s_dadda_rca32_fa151_y4);
  ha ha_h_s_dadda_rca32_ha20_y0(h_s_dadda_rca32_fa145_y2, h_s_dadda_rca32_fa146_y2, h_s_dadda_rca32_ha20_y0, h_s_dadda_rca32_ha20_y1);
  fa fa_h_s_dadda_rca32_fa152_y2(h_s_dadda_rca32_ha20_y1, h_s_dadda_rca32_fa151_y4, h_s_dadda_rca32_fa150_y4, h_s_dadda_rca32_fa152_y2, h_s_dadda_rca32_fa152_y4);
  fa fa_h_s_dadda_rca32_fa153_y2(h_s_dadda_rca32_fa149_y4, h_s_dadda_rca32_fa148_y4, h_s_dadda_rca32_fa147_y4, h_s_dadda_rca32_fa153_y2, h_s_dadda_rca32_fa153_y4);
  fa fa_h_s_dadda_rca32_fa154_y2(h_s_dadda_rca32_fa146_y4, h_s_dadda_rca32_fa145_y4, h_s_dadda_rca32_fa144_y4, h_s_dadda_rca32_fa154_y2, h_s_dadda_rca32_fa154_y4);
  fa fa_h_s_dadda_rca32_fa155_y2(h_s_dadda_rca32_fa143_y4, h_s_dadda_rca32_fa142_y4, h_s_dadda_rca32_fa141_y4, h_s_dadda_rca32_fa155_y2, h_s_dadda_rca32_fa155_y4);
  fa fa_h_s_dadda_rca32_fa156_y2(h_s_dadda_rca32_fa140_y4, h_s_dadda_rca32_fa139_y4, h_s_dadda_rca32_fa138_y4, h_s_dadda_rca32_fa156_y2, h_s_dadda_rca32_fa156_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_0_y0(a_23, b_0, h_s_dadda_rca32_and_23_0_y0);
  fa fa_h_s_dadda_rca32_fa157_y2(h_s_dadda_rca32_fa137_y4, h_s_dadda_rca32_fa136_y4, h_s_dadda_rca32_and_23_0_y0, h_s_dadda_rca32_fa157_y2, h_s_dadda_rca32_fa157_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_1_y0(a_22, b_1, h_s_dadda_rca32_and_22_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_2_y0(a_21, b_2, h_s_dadda_rca32_and_21_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_3_y0(a_20, b_3, h_s_dadda_rca32_and_20_3_y0);
  fa fa_h_s_dadda_rca32_fa158_y2(h_s_dadda_rca32_and_22_1_y0, h_s_dadda_rca32_and_21_2_y0, h_s_dadda_rca32_and_20_3_y0, h_s_dadda_rca32_fa158_y2, h_s_dadda_rca32_fa158_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_4_y0(a_19, b_4, h_s_dadda_rca32_and_19_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_5_y0(a_18, b_5, h_s_dadda_rca32_and_18_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_6_y0(a_17, b_6, h_s_dadda_rca32_and_17_6_y0);
  fa fa_h_s_dadda_rca32_fa159_y2(h_s_dadda_rca32_and_19_4_y0, h_s_dadda_rca32_and_18_5_y0, h_s_dadda_rca32_and_17_6_y0, h_s_dadda_rca32_fa159_y2, h_s_dadda_rca32_fa159_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_7_y0(a_16, b_7, h_s_dadda_rca32_and_16_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_8_y0(a_15, b_8, h_s_dadda_rca32_and_15_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_9_y0(a_14, b_9, h_s_dadda_rca32_and_14_9_y0);
  fa fa_h_s_dadda_rca32_fa160_y2(h_s_dadda_rca32_and_16_7_y0, h_s_dadda_rca32_and_15_8_y0, h_s_dadda_rca32_and_14_9_y0, h_s_dadda_rca32_fa160_y2, h_s_dadda_rca32_fa160_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_10_y0(a_13, b_10, h_s_dadda_rca32_and_13_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_11_y0(a_12, b_11, h_s_dadda_rca32_and_12_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_12_y0(a_11, b_12, h_s_dadda_rca32_and_11_12_y0);
  fa fa_h_s_dadda_rca32_fa161_y2(h_s_dadda_rca32_and_13_10_y0, h_s_dadda_rca32_and_12_11_y0, h_s_dadda_rca32_and_11_12_y0, h_s_dadda_rca32_fa161_y2, h_s_dadda_rca32_fa161_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_13_y0(a_10, b_13, h_s_dadda_rca32_and_10_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_14_y0(a_9, b_14, h_s_dadda_rca32_and_9_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_15_y0(a_8, b_15, h_s_dadda_rca32_and_8_15_y0);
  fa fa_h_s_dadda_rca32_fa162_y2(h_s_dadda_rca32_and_10_13_y0, h_s_dadda_rca32_and_9_14_y0, h_s_dadda_rca32_and_8_15_y0, h_s_dadda_rca32_fa162_y2, h_s_dadda_rca32_fa162_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_16_y0(a_7, b_16, h_s_dadda_rca32_and_7_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_17_y0(a_6, b_17, h_s_dadda_rca32_and_6_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_18_y0(a_5, b_18, h_s_dadda_rca32_and_5_18_y0);
  fa fa_h_s_dadda_rca32_fa163_y2(h_s_dadda_rca32_and_7_16_y0, h_s_dadda_rca32_and_6_17_y0, h_s_dadda_rca32_and_5_18_y0, h_s_dadda_rca32_fa163_y2, h_s_dadda_rca32_fa163_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_19_y0(a_4, b_19, h_s_dadda_rca32_and_4_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_20_y0(a_3, b_20, h_s_dadda_rca32_and_3_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_21_y0(a_2, b_21, h_s_dadda_rca32_and_2_21_y0);
  fa fa_h_s_dadda_rca32_fa164_y2(h_s_dadda_rca32_and_4_19_y0, h_s_dadda_rca32_and_3_20_y0, h_s_dadda_rca32_and_2_21_y0, h_s_dadda_rca32_fa164_y2, h_s_dadda_rca32_fa164_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_22_y0(a_1, b_22, h_s_dadda_rca32_and_1_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_23_y0(a_0, b_23, h_s_dadda_rca32_and_0_23_y0);
  fa fa_h_s_dadda_rca32_fa165_y2(h_s_dadda_rca32_and_1_22_y0, h_s_dadda_rca32_and_0_23_y0, h_s_dadda_rca32_fa152_y2, h_s_dadda_rca32_fa165_y2, h_s_dadda_rca32_fa165_y4);
  fa fa_h_s_dadda_rca32_fa166_y2(h_s_dadda_rca32_fa153_y2, h_s_dadda_rca32_fa154_y2, h_s_dadda_rca32_fa155_y2, h_s_dadda_rca32_fa166_y2, h_s_dadda_rca32_fa166_y4);
  fa fa_h_s_dadda_rca32_fa167_y2(h_s_dadda_rca32_fa156_y2, h_s_dadda_rca32_fa157_y2, h_s_dadda_rca32_fa158_y2, h_s_dadda_rca32_fa167_y2, h_s_dadda_rca32_fa167_y4);
  fa fa_h_s_dadda_rca32_fa168_y2(h_s_dadda_rca32_fa159_y2, h_s_dadda_rca32_fa160_y2, h_s_dadda_rca32_fa161_y2, h_s_dadda_rca32_fa168_y2, h_s_dadda_rca32_fa168_y4);
  ha ha_h_s_dadda_rca32_ha21_y0(h_s_dadda_rca32_fa162_y2, h_s_dadda_rca32_fa163_y2, h_s_dadda_rca32_ha21_y0, h_s_dadda_rca32_ha21_y1);
  fa fa_h_s_dadda_rca32_fa169_y2(h_s_dadda_rca32_ha21_y1, h_s_dadda_rca32_fa168_y4, h_s_dadda_rca32_fa167_y4, h_s_dadda_rca32_fa169_y2, h_s_dadda_rca32_fa169_y4);
  fa fa_h_s_dadda_rca32_fa170_y2(h_s_dadda_rca32_fa166_y4, h_s_dadda_rca32_fa165_y4, h_s_dadda_rca32_fa164_y4, h_s_dadda_rca32_fa170_y2, h_s_dadda_rca32_fa170_y4);
  fa fa_h_s_dadda_rca32_fa171_y2(h_s_dadda_rca32_fa163_y4, h_s_dadda_rca32_fa162_y4, h_s_dadda_rca32_fa161_y4, h_s_dadda_rca32_fa171_y2, h_s_dadda_rca32_fa171_y4);
  fa fa_h_s_dadda_rca32_fa172_y2(h_s_dadda_rca32_fa160_y4, h_s_dadda_rca32_fa159_y4, h_s_dadda_rca32_fa158_y4, h_s_dadda_rca32_fa172_y2, h_s_dadda_rca32_fa172_y4);
  fa fa_h_s_dadda_rca32_fa173_y2(h_s_dadda_rca32_fa157_y4, h_s_dadda_rca32_fa156_y4, h_s_dadda_rca32_fa155_y4, h_s_dadda_rca32_fa173_y2, h_s_dadda_rca32_fa173_y4);
  fa fa_h_s_dadda_rca32_fa174_y2(h_s_dadda_rca32_fa154_y4, h_s_dadda_rca32_fa153_y4, h_s_dadda_rca32_fa152_y4, h_s_dadda_rca32_fa174_y2, h_s_dadda_rca32_fa174_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_0_y0(a_24, b_0, h_s_dadda_rca32_and_24_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_1_y0(a_23, b_1, h_s_dadda_rca32_and_23_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_2_y0(a_22, b_2, h_s_dadda_rca32_and_22_2_y0);
  fa fa_h_s_dadda_rca32_fa175_y2(h_s_dadda_rca32_and_24_0_y0, h_s_dadda_rca32_and_23_1_y0, h_s_dadda_rca32_and_22_2_y0, h_s_dadda_rca32_fa175_y2, h_s_dadda_rca32_fa175_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_3_y0(a_21, b_3, h_s_dadda_rca32_and_21_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_4_y0(a_20, b_4, h_s_dadda_rca32_and_20_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_5_y0(a_19, b_5, h_s_dadda_rca32_and_19_5_y0);
  fa fa_h_s_dadda_rca32_fa176_y2(h_s_dadda_rca32_and_21_3_y0, h_s_dadda_rca32_and_20_4_y0, h_s_dadda_rca32_and_19_5_y0, h_s_dadda_rca32_fa176_y2, h_s_dadda_rca32_fa176_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_6_y0(a_18, b_6, h_s_dadda_rca32_and_18_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_7_y0(a_17, b_7, h_s_dadda_rca32_and_17_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_8_y0(a_16, b_8, h_s_dadda_rca32_and_16_8_y0);
  fa fa_h_s_dadda_rca32_fa177_y2(h_s_dadda_rca32_and_18_6_y0, h_s_dadda_rca32_and_17_7_y0, h_s_dadda_rca32_and_16_8_y0, h_s_dadda_rca32_fa177_y2, h_s_dadda_rca32_fa177_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_9_y0(a_15, b_9, h_s_dadda_rca32_and_15_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_10_y0(a_14, b_10, h_s_dadda_rca32_and_14_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_11_y0(a_13, b_11, h_s_dadda_rca32_and_13_11_y0);
  fa fa_h_s_dadda_rca32_fa178_y2(h_s_dadda_rca32_and_15_9_y0, h_s_dadda_rca32_and_14_10_y0, h_s_dadda_rca32_and_13_11_y0, h_s_dadda_rca32_fa178_y2, h_s_dadda_rca32_fa178_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_12_y0(a_12, b_12, h_s_dadda_rca32_and_12_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_13_y0(a_11, b_13, h_s_dadda_rca32_and_11_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_14_y0(a_10, b_14, h_s_dadda_rca32_and_10_14_y0);
  fa fa_h_s_dadda_rca32_fa179_y2(h_s_dadda_rca32_and_12_12_y0, h_s_dadda_rca32_and_11_13_y0, h_s_dadda_rca32_and_10_14_y0, h_s_dadda_rca32_fa179_y2, h_s_dadda_rca32_fa179_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_15_y0(a_9, b_15, h_s_dadda_rca32_and_9_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_16_y0(a_8, b_16, h_s_dadda_rca32_and_8_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_17_y0(a_7, b_17, h_s_dadda_rca32_and_7_17_y0);
  fa fa_h_s_dadda_rca32_fa180_y2(h_s_dadda_rca32_and_9_15_y0, h_s_dadda_rca32_and_8_16_y0, h_s_dadda_rca32_and_7_17_y0, h_s_dadda_rca32_fa180_y2, h_s_dadda_rca32_fa180_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_18_y0(a_6, b_18, h_s_dadda_rca32_and_6_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_19_y0(a_5, b_19, h_s_dadda_rca32_and_5_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_20_y0(a_4, b_20, h_s_dadda_rca32_and_4_20_y0);
  fa fa_h_s_dadda_rca32_fa181_y2(h_s_dadda_rca32_and_6_18_y0, h_s_dadda_rca32_and_5_19_y0, h_s_dadda_rca32_and_4_20_y0, h_s_dadda_rca32_fa181_y2, h_s_dadda_rca32_fa181_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_21_y0(a_3, b_21, h_s_dadda_rca32_and_3_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_22_y0(a_2, b_22, h_s_dadda_rca32_and_2_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_23_y0(a_1, b_23, h_s_dadda_rca32_and_1_23_y0);
  fa fa_h_s_dadda_rca32_fa182_y2(h_s_dadda_rca32_and_3_21_y0, h_s_dadda_rca32_and_2_22_y0, h_s_dadda_rca32_and_1_23_y0, h_s_dadda_rca32_fa182_y2, h_s_dadda_rca32_fa182_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_24_y0(a_0, b_24, h_s_dadda_rca32_and_0_24_y0);
  fa fa_h_s_dadda_rca32_fa183_y2(h_s_dadda_rca32_and_0_24_y0, h_s_dadda_rca32_fa169_y2, h_s_dadda_rca32_fa170_y2, h_s_dadda_rca32_fa183_y2, h_s_dadda_rca32_fa183_y4);
  fa fa_h_s_dadda_rca32_fa184_y2(h_s_dadda_rca32_fa171_y2, h_s_dadda_rca32_fa172_y2, h_s_dadda_rca32_fa173_y2, h_s_dadda_rca32_fa184_y2, h_s_dadda_rca32_fa184_y4);
  fa fa_h_s_dadda_rca32_fa185_y2(h_s_dadda_rca32_fa174_y2, h_s_dadda_rca32_fa175_y2, h_s_dadda_rca32_fa176_y2, h_s_dadda_rca32_fa185_y2, h_s_dadda_rca32_fa185_y4);
  fa fa_h_s_dadda_rca32_fa186_y2(h_s_dadda_rca32_fa177_y2, h_s_dadda_rca32_fa178_y2, h_s_dadda_rca32_fa179_y2, h_s_dadda_rca32_fa186_y2, h_s_dadda_rca32_fa186_y4);
  ha ha_h_s_dadda_rca32_ha22_y0(h_s_dadda_rca32_fa180_y2, h_s_dadda_rca32_fa181_y2, h_s_dadda_rca32_ha22_y0, h_s_dadda_rca32_ha22_y1);
  fa fa_h_s_dadda_rca32_fa187_y2(h_s_dadda_rca32_ha22_y1, h_s_dadda_rca32_fa186_y4, h_s_dadda_rca32_fa185_y4, h_s_dadda_rca32_fa187_y2, h_s_dadda_rca32_fa187_y4);
  fa fa_h_s_dadda_rca32_fa188_y2(h_s_dadda_rca32_fa184_y4, h_s_dadda_rca32_fa183_y4, h_s_dadda_rca32_fa182_y4, h_s_dadda_rca32_fa188_y2, h_s_dadda_rca32_fa188_y4);
  fa fa_h_s_dadda_rca32_fa189_y2(h_s_dadda_rca32_fa181_y4, h_s_dadda_rca32_fa180_y4, h_s_dadda_rca32_fa179_y4, h_s_dadda_rca32_fa189_y2, h_s_dadda_rca32_fa189_y4);
  fa fa_h_s_dadda_rca32_fa190_y2(h_s_dadda_rca32_fa178_y4, h_s_dadda_rca32_fa177_y4, h_s_dadda_rca32_fa176_y4, h_s_dadda_rca32_fa190_y2, h_s_dadda_rca32_fa190_y4);
  fa fa_h_s_dadda_rca32_fa191_y2(h_s_dadda_rca32_fa175_y4, h_s_dadda_rca32_fa174_y4, h_s_dadda_rca32_fa173_y4, h_s_dadda_rca32_fa191_y2, h_s_dadda_rca32_fa191_y4);
  fa fa_h_s_dadda_rca32_fa192_y2(h_s_dadda_rca32_fa172_y4, h_s_dadda_rca32_fa171_y4, h_s_dadda_rca32_fa170_y4, h_s_dadda_rca32_fa192_y2, h_s_dadda_rca32_fa192_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_0_y0(a_25, b_0, h_s_dadda_rca32_and_25_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_1_y0(a_24, b_1, h_s_dadda_rca32_and_24_1_y0);
  fa fa_h_s_dadda_rca32_fa193_y2(h_s_dadda_rca32_fa169_y4, h_s_dadda_rca32_and_25_0_y0, h_s_dadda_rca32_and_24_1_y0, h_s_dadda_rca32_fa193_y2, h_s_dadda_rca32_fa193_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_2_y0(a_23, b_2, h_s_dadda_rca32_and_23_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_3_y0(a_22, b_3, h_s_dadda_rca32_and_22_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_4_y0(a_21, b_4, h_s_dadda_rca32_and_21_4_y0);
  fa fa_h_s_dadda_rca32_fa194_y2(h_s_dadda_rca32_and_23_2_y0, h_s_dadda_rca32_and_22_3_y0, h_s_dadda_rca32_and_21_4_y0, h_s_dadda_rca32_fa194_y2, h_s_dadda_rca32_fa194_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_5_y0(a_20, b_5, h_s_dadda_rca32_and_20_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_6_y0(a_19, b_6, h_s_dadda_rca32_and_19_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_7_y0(a_18, b_7, h_s_dadda_rca32_and_18_7_y0);
  fa fa_h_s_dadda_rca32_fa195_y2(h_s_dadda_rca32_and_20_5_y0, h_s_dadda_rca32_and_19_6_y0, h_s_dadda_rca32_and_18_7_y0, h_s_dadda_rca32_fa195_y2, h_s_dadda_rca32_fa195_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_8_y0(a_17, b_8, h_s_dadda_rca32_and_17_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_9_y0(a_16, b_9, h_s_dadda_rca32_and_16_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_10_y0(a_15, b_10, h_s_dadda_rca32_and_15_10_y0);
  fa fa_h_s_dadda_rca32_fa196_y2(h_s_dadda_rca32_and_17_8_y0, h_s_dadda_rca32_and_16_9_y0, h_s_dadda_rca32_and_15_10_y0, h_s_dadda_rca32_fa196_y2, h_s_dadda_rca32_fa196_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_11_y0(a_14, b_11, h_s_dadda_rca32_and_14_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_12_y0(a_13, b_12, h_s_dadda_rca32_and_13_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_13_y0(a_12, b_13, h_s_dadda_rca32_and_12_13_y0);
  fa fa_h_s_dadda_rca32_fa197_y2(h_s_dadda_rca32_and_14_11_y0, h_s_dadda_rca32_and_13_12_y0, h_s_dadda_rca32_and_12_13_y0, h_s_dadda_rca32_fa197_y2, h_s_dadda_rca32_fa197_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_14_y0(a_11, b_14, h_s_dadda_rca32_and_11_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_15_y0(a_10, b_15, h_s_dadda_rca32_and_10_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_16_y0(a_9, b_16, h_s_dadda_rca32_and_9_16_y0);
  fa fa_h_s_dadda_rca32_fa198_y2(h_s_dadda_rca32_and_11_14_y0, h_s_dadda_rca32_and_10_15_y0, h_s_dadda_rca32_and_9_16_y0, h_s_dadda_rca32_fa198_y2, h_s_dadda_rca32_fa198_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_17_y0(a_8, b_17, h_s_dadda_rca32_and_8_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_18_y0(a_7, b_18, h_s_dadda_rca32_and_7_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_19_y0(a_6, b_19, h_s_dadda_rca32_and_6_19_y0);
  fa fa_h_s_dadda_rca32_fa199_y2(h_s_dadda_rca32_and_8_17_y0, h_s_dadda_rca32_and_7_18_y0, h_s_dadda_rca32_and_6_19_y0, h_s_dadda_rca32_fa199_y2, h_s_dadda_rca32_fa199_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_20_y0(a_5, b_20, h_s_dadda_rca32_and_5_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_21_y0(a_4, b_21, h_s_dadda_rca32_and_4_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_22_y0(a_3, b_22, h_s_dadda_rca32_and_3_22_y0);
  fa fa_h_s_dadda_rca32_fa200_y2(h_s_dadda_rca32_and_5_20_y0, h_s_dadda_rca32_and_4_21_y0, h_s_dadda_rca32_and_3_22_y0, h_s_dadda_rca32_fa200_y2, h_s_dadda_rca32_fa200_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_23_y0(a_2, b_23, h_s_dadda_rca32_and_2_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_24_y0(a_1, b_24, h_s_dadda_rca32_and_1_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_25_y0(a_0, b_25, h_s_dadda_rca32_and_0_25_y0);
  fa fa_h_s_dadda_rca32_fa201_y2(h_s_dadda_rca32_and_2_23_y0, h_s_dadda_rca32_and_1_24_y0, h_s_dadda_rca32_and_0_25_y0, h_s_dadda_rca32_fa201_y2, h_s_dadda_rca32_fa201_y4);
  fa fa_h_s_dadda_rca32_fa202_y2(h_s_dadda_rca32_fa187_y2, h_s_dadda_rca32_fa188_y2, h_s_dadda_rca32_fa189_y2, h_s_dadda_rca32_fa202_y2, h_s_dadda_rca32_fa202_y4);
  fa fa_h_s_dadda_rca32_fa203_y2(h_s_dadda_rca32_fa190_y2, h_s_dadda_rca32_fa191_y2, h_s_dadda_rca32_fa192_y2, h_s_dadda_rca32_fa203_y2, h_s_dadda_rca32_fa203_y4);
  fa fa_h_s_dadda_rca32_fa204_y2(h_s_dadda_rca32_fa193_y2, h_s_dadda_rca32_fa194_y2, h_s_dadda_rca32_fa195_y2, h_s_dadda_rca32_fa204_y2, h_s_dadda_rca32_fa204_y4);
  fa fa_h_s_dadda_rca32_fa205_y2(h_s_dadda_rca32_fa196_y2, h_s_dadda_rca32_fa197_y2, h_s_dadda_rca32_fa198_y2, h_s_dadda_rca32_fa205_y2, h_s_dadda_rca32_fa205_y4);
  ha ha_h_s_dadda_rca32_ha23_y0(h_s_dadda_rca32_fa199_y2, h_s_dadda_rca32_fa200_y2, h_s_dadda_rca32_ha23_y0, h_s_dadda_rca32_ha23_y1);
  fa fa_h_s_dadda_rca32_fa206_y2(h_s_dadda_rca32_ha23_y1, h_s_dadda_rca32_fa205_y4, h_s_dadda_rca32_fa204_y4, h_s_dadda_rca32_fa206_y2, h_s_dadda_rca32_fa206_y4);
  fa fa_h_s_dadda_rca32_fa207_y2(h_s_dadda_rca32_fa203_y4, h_s_dadda_rca32_fa202_y4, h_s_dadda_rca32_fa201_y4, h_s_dadda_rca32_fa207_y2, h_s_dadda_rca32_fa207_y4);
  fa fa_h_s_dadda_rca32_fa208_y2(h_s_dadda_rca32_fa200_y4, h_s_dadda_rca32_fa199_y4, h_s_dadda_rca32_fa198_y4, h_s_dadda_rca32_fa208_y2, h_s_dadda_rca32_fa208_y4);
  fa fa_h_s_dadda_rca32_fa209_y2(h_s_dadda_rca32_fa197_y4, h_s_dadda_rca32_fa196_y4, h_s_dadda_rca32_fa195_y4, h_s_dadda_rca32_fa209_y2, h_s_dadda_rca32_fa209_y4);
  fa fa_h_s_dadda_rca32_fa210_y2(h_s_dadda_rca32_fa194_y4, h_s_dadda_rca32_fa193_y4, h_s_dadda_rca32_fa192_y4, h_s_dadda_rca32_fa210_y2, h_s_dadda_rca32_fa210_y4);
  fa fa_h_s_dadda_rca32_fa211_y2(h_s_dadda_rca32_fa191_y4, h_s_dadda_rca32_fa190_y4, h_s_dadda_rca32_fa189_y4, h_s_dadda_rca32_fa211_y2, h_s_dadda_rca32_fa211_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_0_y0(a_26, b_0, h_s_dadda_rca32_and_26_0_y0);
  fa fa_h_s_dadda_rca32_fa212_y2(h_s_dadda_rca32_fa188_y4, h_s_dadda_rca32_fa187_y4, h_s_dadda_rca32_and_26_0_y0, h_s_dadda_rca32_fa212_y2, h_s_dadda_rca32_fa212_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_1_y0(a_25, b_1, h_s_dadda_rca32_and_25_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_2_y0(a_24, b_2, h_s_dadda_rca32_and_24_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_3_y0(a_23, b_3, h_s_dadda_rca32_and_23_3_y0);
  fa fa_h_s_dadda_rca32_fa213_y2(h_s_dadda_rca32_and_25_1_y0, h_s_dadda_rca32_and_24_2_y0, h_s_dadda_rca32_and_23_3_y0, h_s_dadda_rca32_fa213_y2, h_s_dadda_rca32_fa213_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_4_y0(a_22, b_4, h_s_dadda_rca32_and_22_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_5_y0(a_21, b_5, h_s_dadda_rca32_and_21_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_6_y0(a_20, b_6, h_s_dadda_rca32_and_20_6_y0);
  fa fa_h_s_dadda_rca32_fa214_y2(h_s_dadda_rca32_and_22_4_y0, h_s_dadda_rca32_and_21_5_y0, h_s_dadda_rca32_and_20_6_y0, h_s_dadda_rca32_fa214_y2, h_s_dadda_rca32_fa214_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_7_y0(a_19, b_7, h_s_dadda_rca32_and_19_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_8_y0(a_18, b_8, h_s_dadda_rca32_and_18_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_9_y0(a_17, b_9, h_s_dadda_rca32_and_17_9_y0);
  fa fa_h_s_dadda_rca32_fa215_y2(h_s_dadda_rca32_and_19_7_y0, h_s_dadda_rca32_and_18_8_y0, h_s_dadda_rca32_and_17_9_y0, h_s_dadda_rca32_fa215_y2, h_s_dadda_rca32_fa215_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_10_y0(a_16, b_10, h_s_dadda_rca32_and_16_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_11_y0(a_15, b_11, h_s_dadda_rca32_and_15_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_12_y0(a_14, b_12, h_s_dadda_rca32_and_14_12_y0);
  fa fa_h_s_dadda_rca32_fa216_y2(h_s_dadda_rca32_and_16_10_y0, h_s_dadda_rca32_and_15_11_y0, h_s_dadda_rca32_and_14_12_y0, h_s_dadda_rca32_fa216_y2, h_s_dadda_rca32_fa216_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_13_y0(a_13, b_13, h_s_dadda_rca32_and_13_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_14_y0(a_12, b_14, h_s_dadda_rca32_and_12_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_15_y0(a_11, b_15, h_s_dadda_rca32_and_11_15_y0);
  fa fa_h_s_dadda_rca32_fa217_y2(h_s_dadda_rca32_and_13_13_y0, h_s_dadda_rca32_and_12_14_y0, h_s_dadda_rca32_and_11_15_y0, h_s_dadda_rca32_fa217_y2, h_s_dadda_rca32_fa217_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_16_y0(a_10, b_16, h_s_dadda_rca32_and_10_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_17_y0(a_9, b_17, h_s_dadda_rca32_and_9_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_18_y0(a_8, b_18, h_s_dadda_rca32_and_8_18_y0);
  fa fa_h_s_dadda_rca32_fa218_y2(h_s_dadda_rca32_and_10_16_y0, h_s_dadda_rca32_and_9_17_y0, h_s_dadda_rca32_and_8_18_y0, h_s_dadda_rca32_fa218_y2, h_s_dadda_rca32_fa218_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_19_y0(a_7, b_19, h_s_dadda_rca32_and_7_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_20_y0(a_6, b_20, h_s_dadda_rca32_and_6_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_21_y0(a_5, b_21, h_s_dadda_rca32_and_5_21_y0);
  fa fa_h_s_dadda_rca32_fa219_y2(h_s_dadda_rca32_and_7_19_y0, h_s_dadda_rca32_and_6_20_y0, h_s_dadda_rca32_and_5_21_y0, h_s_dadda_rca32_fa219_y2, h_s_dadda_rca32_fa219_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_22_y0(a_4, b_22, h_s_dadda_rca32_and_4_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_23_y0(a_3, b_23, h_s_dadda_rca32_and_3_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_24_y0(a_2, b_24, h_s_dadda_rca32_and_2_24_y0);
  fa fa_h_s_dadda_rca32_fa220_y2(h_s_dadda_rca32_and_4_22_y0, h_s_dadda_rca32_and_3_23_y0, h_s_dadda_rca32_and_2_24_y0, h_s_dadda_rca32_fa220_y2, h_s_dadda_rca32_fa220_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_25_y0(a_1, b_25, h_s_dadda_rca32_and_1_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_26_y0(a_0, b_26, h_s_dadda_rca32_and_0_26_y0);
  fa fa_h_s_dadda_rca32_fa221_y2(h_s_dadda_rca32_and_1_25_y0, h_s_dadda_rca32_and_0_26_y0, h_s_dadda_rca32_fa206_y2, h_s_dadda_rca32_fa221_y2, h_s_dadda_rca32_fa221_y4);
  fa fa_h_s_dadda_rca32_fa222_y2(h_s_dadda_rca32_fa207_y2, h_s_dadda_rca32_fa208_y2, h_s_dadda_rca32_fa209_y2, h_s_dadda_rca32_fa222_y2, h_s_dadda_rca32_fa222_y4);
  fa fa_h_s_dadda_rca32_fa223_y2(h_s_dadda_rca32_fa210_y2, h_s_dadda_rca32_fa211_y2, h_s_dadda_rca32_fa212_y2, h_s_dadda_rca32_fa223_y2, h_s_dadda_rca32_fa223_y4);
  fa fa_h_s_dadda_rca32_fa224_y2(h_s_dadda_rca32_fa213_y2, h_s_dadda_rca32_fa214_y2, h_s_dadda_rca32_fa215_y2, h_s_dadda_rca32_fa224_y2, h_s_dadda_rca32_fa224_y4);
  fa fa_h_s_dadda_rca32_fa225_y2(h_s_dadda_rca32_fa216_y2, h_s_dadda_rca32_fa217_y2, h_s_dadda_rca32_fa218_y2, h_s_dadda_rca32_fa225_y2, h_s_dadda_rca32_fa225_y4);
  ha ha_h_s_dadda_rca32_ha24_y0(h_s_dadda_rca32_fa219_y2, h_s_dadda_rca32_fa220_y2, h_s_dadda_rca32_ha24_y0, h_s_dadda_rca32_ha24_y1);
  fa fa_h_s_dadda_rca32_fa226_y2(h_s_dadda_rca32_ha24_y1, h_s_dadda_rca32_fa225_y4, h_s_dadda_rca32_fa224_y4, h_s_dadda_rca32_fa226_y2, h_s_dadda_rca32_fa226_y4);
  fa fa_h_s_dadda_rca32_fa227_y2(h_s_dadda_rca32_fa223_y4, h_s_dadda_rca32_fa222_y4, h_s_dadda_rca32_fa221_y4, h_s_dadda_rca32_fa227_y2, h_s_dadda_rca32_fa227_y4);
  fa fa_h_s_dadda_rca32_fa228_y2(h_s_dadda_rca32_fa220_y4, h_s_dadda_rca32_fa219_y4, h_s_dadda_rca32_fa218_y4, h_s_dadda_rca32_fa228_y2, h_s_dadda_rca32_fa228_y4);
  fa fa_h_s_dadda_rca32_fa229_y2(h_s_dadda_rca32_fa217_y4, h_s_dadda_rca32_fa216_y4, h_s_dadda_rca32_fa215_y4, h_s_dadda_rca32_fa229_y2, h_s_dadda_rca32_fa229_y4);
  fa fa_h_s_dadda_rca32_fa230_y2(h_s_dadda_rca32_fa214_y4, h_s_dadda_rca32_fa213_y4, h_s_dadda_rca32_fa212_y4, h_s_dadda_rca32_fa230_y2, h_s_dadda_rca32_fa230_y4);
  fa fa_h_s_dadda_rca32_fa231_y2(h_s_dadda_rca32_fa211_y4, h_s_dadda_rca32_fa210_y4, h_s_dadda_rca32_fa209_y4, h_s_dadda_rca32_fa231_y2, h_s_dadda_rca32_fa231_y4);
  fa fa_h_s_dadda_rca32_fa232_y2(h_s_dadda_rca32_fa208_y4, h_s_dadda_rca32_fa207_y4, h_s_dadda_rca32_fa206_y4, h_s_dadda_rca32_fa232_y2, h_s_dadda_rca32_fa232_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_0_y0(a_27, b_0, h_s_dadda_rca32_and_27_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_1_y0(a_26, b_1, h_s_dadda_rca32_and_26_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_2_y0(a_25, b_2, h_s_dadda_rca32_and_25_2_y0);
  fa fa_h_s_dadda_rca32_fa233_y2(h_s_dadda_rca32_and_27_0_y0, h_s_dadda_rca32_and_26_1_y0, h_s_dadda_rca32_and_25_2_y0, h_s_dadda_rca32_fa233_y2, h_s_dadda_rca32_fa233_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_3_y0(a_24, b_3, h_s_dadda_rca32_and_24_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_4_y0(a_23, b_4, h_s_dadda_rca32_and_23_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_5_y0(a_22, b_5, h_s_dadda_rca32_and_22_5_y0);
  fa fa_h_s_dadda_rca32_fa234_y2(h_s_dadda_rca32_and_24_3_y0, h_s_dadda_rca32_and_23_4_y0, h_s_dadda_rca32_and_22_5_y0, h_s_dadda_rca32_fa234_y2, h_s_dadda_rca32_fa234_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_6_y0(a_21, b_6, h_s_dadda_rca32_and_21_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_7_y0(a_20, b_7, h_s_dadda_rca32_and_20_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_8_y0(a_19, b_8, h_s_dadda_rca32_and_19_8_y0);
  fa fa_h_s_dadda_rca32_fa235_y2(h_s_dadda_rca32_and_21_6_y0, h_s_dadda_rca32_and_20_7_y0, h_s_dadda_rca32_and_19_8_y0, h_s_dadda_rca32_fa235_y2, h_s_dadda_rca32_fa235_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_9_y0(a_18, b_9, h_s_dadda_rca32_and_18_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_10_y0(a_17, b_10, h_s_dadda_rca32_and_17_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_11_y0(a_16, b_11, h_s_dadda_rca32_and_16_11_y0);
  fa fa_h_s_dadda_rca32_fa236_y2(h_s_dadda_rca32_and_18_9_y0, h_s_dadda_rca32_and_17_10_y0, h_s_dadda_rca32_and_16_11_y0, h_s_dadda_rca32_fa236_y2, h_s_dadda_rca32_fa236_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_12_y0(a_15, b_12, h_s_dadda_rca32_and_15_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_13_y0(a_14, b_13, h_s_dadda_rca32_and_14_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_14_y0(a_13, b_14, h_s_dadda_rca32_and_13_14_y0);
  fa fa_h_s_dadda_rca32_fa237_y2(h_s_dadda_rca32_and_15_12_y0, h_s_dadda_rca32_and_14_13_y0, h_s_dadda_rca32_and_13_14_y0, h_s_dadda_rca32_fa237_y2, h_s_dadda_rca32_fa237_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_15_y0(a_12, b_15, h_s_dadda_rca32_and_12_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_16_y0(a_11, b_16, h_s_dadda_rca32_and_11_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_17_y0(a_10, b_17, h_s_dadda_rca32_and_10_17_y0);
  fa fa_h_s_dadda_rca32_fa238_y2(h_s_dadda_rca32_and_12_15_y0, h_s_dadda_rca32_and_11_16_y0, h_s_dadda_rca32_and_10_17_y0, h_s_dadda_rca32_fa238_y2, h_s_dadda_rca32_fa238_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_18_y0(a_9, b_18, h_s_dadda_rca32_and_9_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_19_y0(a_8, b_19, h_s_dadda_rca32_and_8_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_20_y0(a_7, b_20, h_s_dadda_rca32_and_7_20_y0);
  fa fa_h_s_dadda_rca32_fa239_y2(h_s_dadda_rca32_and_9_18_y0, h_s_dadda_rca32_and_8_19_y0, h_s_dadda_rca32_and_7_20_y0, h_s_dadda_rca32_fa239_y2, h_s_dadda_rca32_fa239_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_21_y0(a_6, b_21, h_s_dadda_rca32_and_6_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_22_y0(a_5, b_22, h_s_dadda_rca32_and_5_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_23_y0(a_4, b_23, h_s_dadda_rca32_and_4_23_y0);
  fa fa_h_s_dadda_rca32_fa240_y2(h_s_dadda_rca32_and_6_21_y0, h_s_dadda_rca32_and_5_22_y0, h_s_dadda_rca32_and_4_23_y0, h_s_dadda_rca32_fa240_y2, h_s_dadda_rca32_fa240_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_24_y0(a_3, b_24, h_s_dadda_rca32_and_3_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_25_y0(a_2, b_25, h_s_dadda_rca32_and_2_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_26_y0(a_1, b_26, h_s_dadda_rca32_and_1_26_y0);
  fa fa_h_s_dadda_rca32_fa241_y2(h_s_dadda_rca32_and_3_24_y0, h_s_dadda_rca32_and_2_25_y0, h_s_dadda_rca32_and_1_26_y0, h_s_dadda_rca32_fa241_y2, h_s_dadda_rca32_fa241_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_27_y0(a_0, b_27, h_s_dadda_rca32_and_0_27_y0);
  fa fa_h_s_dadda_rca32_fa242_y2(h_s_dadda_rca32_and_0_27_y0, h_s_dadda_rca32_fa226_y2, h_s_dadda_rca32_fa227_y2, h_s_dadda_rca32_fa242_y2, h_s_dadda_rca32_fa242_y4);
  fa fa_h_s_dadda_rca32_fa243_y2(h_s_dadda_rca32_fa228_y2, h_s_dadda_rca32_fa229_y2, h_s_dadda_rca32_fa230_y2, h_s_dadda_rca32_fa243_y2, h_s_dadda_rca32_fa243_y4);
  fa fa_h_s_dadda_rca32_fa244_y2(h_s_dadda_rca32_fa231_y2, h_s_dadda_rca32_fa232_y2, h_s_dadda_rca32_fa233_y2, h_s_dadda_rca32_fa244_y2, h_s_dadda_rca32_fa244_y4);
  fa fa_h_s_dadda_rca32_fa245_y2(h_s_dadda_rca32_fa234_y2, h_s_dadda_rca32_fa235_y2, h_s_dadda_rca32_fa236_y2, h_s_dadda_rca32_fa245_y2, h_s_dadda_rca32_fa245_y4);
  fa fa_h_s_dadda_rca32_fa246_y2(h_s_dadda_rca32_fa237_y2, h_s_dadda_rca32_fa238_y2, h_s_dadda_rca32_fa239_y2, h_s_dadda_rca32_fa246_y2, h_s_dadda_rca32_fa246_y4);
  ha ha_h_s_dadda_rca32_ha25_y0(h_s_dadda_rca32_fa240_y2, h_s_dadda_rca32_fa241_y2, h_s_dadda_rca32_ha25_y0, h_s_dadda_rca32_ha25_y1);
  fa fa_h_s_dadda_rca32_fa247_y2(h_s_dadda_rca32_ha25_y1, h_s_dadda_rca32_fa246_y4, h_s_dadda_rca32_fa245_y4, h_s_dadda_rca32_fa247_y2, h_s_dadda_rca32_fa247_y4);
  fa fa_h_s_dadda_rca32_fa248_y2(h_s_dadda_rca32_fa244_y4, h_s_dadda_rca32_fa243_y4, h_s_dadda_rca32_fa242_y4, h_s_dadda_rca32_fa248_y2, h_s_dadda_rca32_fa248_y4);
  fa fa_h_s_dadda_rca32_fa249_y2(h_s_dadda_rca32_fa241_y4, h_s_dadda_rca32_fa240_y4, h_s_dadda_rca32_fa239_y4, h_s_dadda_rca32_fa249_y2, h_s_dadda_rca32_fa249_y4);
  fa fa_h_s_dadda_rca32_fa250_y2(h_s_dadda_rca32_fa238_y4, h_s_dadda_rca32_fa237_y4, h_s_dadda_rca32_fa236_y4, h_s_dadda_rca32_fa250_y2, h_s_dadda_rca32_fa250_y4);
  fa fa_h_s_dadda_rca32_fa251_y2(h_s_dadda_rca32_fa235_y4, h_s_dadda_rca32_fa234_y4, h_s_dadda_rca32_fa233_y4, h_s_dadda_rca32_fa251_y2, h_s_dadda_rca32_fa251_y4);
  fa fa_h_s_dadda_rca32_fa252_y2(h_s_dadda_rca32_fa232_y4, h_s_dadda_rca32_fa231_y4, h_s_dadda_rca32_fa230_y4, h_s_dadda_rca32_fa252_y2, h_s_dadda_rca32_fa252_y4);
  fa fa_h_s_dadda_rca32_fa253_y2(h_s_dadda_rca32_fa229_y4, h_s_dadda_rca32_fa228_y4, h_s_dadda_rca32_fa227_y4, h_s_dadda_rca32_fa253_y2, h_s_dadda_rca32_fa253_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_2_y0(a_26, b_2, h_s_dadda_rca32_and_26_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_3_y0(a_25, b_3, h_s_dadda_rca32_and_25_3_y0);
  fa fa_h_s_dadda_rca32_fa254_y2(h_s_dadda_rca32_fa226_y4, h_s_dadda_rca32_and_26_2_y0, h_s_dadda_rca32_and_25_3_y0, h_s_dadda_rca32_fa254_y2, h_s_dadda_rca32_fa254_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_4_y0(a_24, b_4, h_s_dadda_rca32_and_24_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_5_y0(a_23, b_5, h_s_dadda_rca32_and_23_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_6_y0(a_22, b_6, h_s_dadda_rca32_and_22_6_y0);
  fa fa_h_s_dadda_rca32_fa255_y2(h_s_dadda_rca32_and_24_4_y0, h_s_dadda_rca32_and_23_5_y0, h_s_dadda_rca32_and_22_6_y0, h_s_dadda_rca32_fa255_y2, h_s_dadda_rca32_fa255_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_7_y0(a_21, b_7, h_s_dadda_rca32_and_21_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_8_y0(a_20, b_8, h_s_dadda_rca32_and_20_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_9_y0(a_19, b_9, h_s_dadda_rca32_and_19_9_y0);
  fa fa_h_s_dadda_rca32_fa256_y2(h_s_dadda_rca32_and_21_7_y0, h_s_dadda_rca32_and_20_8_y0, h_s_dadda_rca32_and_19_9_y0, h_s_dadda_rca32_fa256_y2, h_s_dadda_rca32_fa256_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_10_y0(a_18, b_10, h_s_dadda_rca32_and_18_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_11_y0(a_17, b_11, h_s_dadda_rca32_and_17_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_12_y0(a_16, b_12, h_s_dadda_rca32_and_16_12_y0);
  fa fa_h_s_dadda_rca32_fa257_y2(h_s_dadda_rca32_and_18_10_y0, h_s_dadda_rca32_and_17_11_y0, h_s_dadda_rca32_and_16_12_y0, h_s_dadda_rca32_fa257_y2, h_s_dadda_rca32_fa257_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_13_y0(a_15, b_13, h_s_dadda_rca32_and_15_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_14_y0(a_14, b_14, h_s_dadda_rca32_and_14_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_15_y0(a_13, b_15, h_s_dadda_rca32_and_13_15_y0);
  fa fa_h_s_dadda_rca32_fa258_y2(h_s_dadda_rca32_and_15_13_y0, h_s_dadda_rca32_and_14_14_y0, h_s_dadda_rca32_and_13_15_y0, h_s_dadda_rca32_fa258_y2, h_s_dadda_rca32_fa258_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_16_y0(a_12, b_16, h_s_dadda_rca32_and_12_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_17_y0(a_11, b_17, h_s_dadda_rca32_and_11_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_18_y0(a_10, b_18, h_s_dadda_rca32_and_10_18_y0);
  fa fa_h_s_dadda_rca32_fa259_y2(h_s_dadda_rca32_and_12_16_y0, h_s_dadda_rca32_and_11_17_y0, h_s_dadda_rca32_and_10_18_y0, h_s_dadda_rca32_fa259_y2, h_s_dadda_rca32_fa259_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_19_y0(a_9, b_19, h_s_dadda_rca32_and_9_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_20_y0(a_8, b_20, h_s_dadda_rca32_and_8_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_21_y0(a_7, b_21, h_s_dadda_rca32_and_7_21_y0);
  fa fa_h_s_dadda_rca32_fa260_y2(h_s_dadda_rca32_and_9_19_y0, h_s_dadda_rca32_and_8_20_y0, h_s_dadda_rca32_and_7_21_y0, h_s_dadda_rca32_fa260_y2, h_s_dadda_rca32_fa260_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_22_y0(a_6, b_22, h_s_dadda_rca32_and_6_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_23_y0(a_5, b_23, h_s_dadda_rca32_and_5_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_24_y0(a_4, b_24, h_s_dadda_rca32_and_4_24_y0);
  fa fa_h_s_dadda_rca32_fa261_y2(h_s_dadda_rca32_and_6_22_y0, h_s_dadda_rca32_and_5_23_y0, h_s_dadda_rca32_and_4_24_y0, h_s_dadda_rca32_fa261_y2, h_s_dadda_rca32_fa261_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_25_y0(a_3, b_25, h_s_dadda_rca32_and_3_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_26_y0(a_2, b_26, h_s_dadda_rca32_and_2_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_27_y0(a_1, b_27, h_s_dadda_rca32_and_1_27_y0);
  fa fa_h_s_dadda_rca32_fa262_y2(h_s_dadda_rca32_and_3_25_y0, h_s_dadda_rca32_and_2_26_y0, h_s_dadda_rca32_and_1_27_y0, h_s_dadda_rca32_fa262_y2, h_s_dadda_rca32_fa262_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_28_y0(a_0, b_28, h_s_dadda_rca32_and_0_28_y0);
  fa fa_h_s_dadda_rca32_fa263_y2(h_s_dadda_rca32_and_0_28_y0, h_s_dadda_rca32_ha0_y0, h_s_dadda_rca32_fa247_y2, h_s_dadda_rca32_fa263_y2, h_s_dadda_rca32_fa263_y4);
  fa fa_h_s_dadda_rca32_fa264_y2(h_s_dadda_rca32_fa248_y2, h_s_dadda_rca32_fa249_y2, h_s_dadda_rca32_fa250_y2, h_s_dadda_rca32_fa264_y2, h_s_dadda_rca32_fa264_y4);
  fa fa_h_s_dadda_rca32_fa265_y2(h_s_dadda_rca32_fa251_y2, h_s_dadda_rca32_fa252_y2, h_s_dadda_rca32_fa253_y2, h_s_dadda_rca32_fa265_y2, h_s_dadda_rca32_fa265_y4);
  fa fa_h_s_dadda_rca32_fa266_y2(h_s_dadda_rca32_fa254_y2, h_s_dadda_rca32_fa255_y2, h_s_dadda_rca32_fa256_y2, h_s_dadda_rca32_fa266_y2, h_s_dadda_rca32_fa266_y4);
  fa fa_h_s_dadda_rca32_fa267_y2(h_s_dadda_rca32_fa257_y2, h_s_dadda_rca32_fa258_y2, h_s_dadda_rca32_fa259_y2, h_s_dadda_rca32_fa267_y2, h_s_dadda_rca32_fa267_y4);
  fa fa_h_s_dadda_rca32_fa268_y2(h_s_dadda_rca32_fa260_y2, h_s_dadda_rca32_fa261_y2, h_s_dadda_rca32_fa262_y2, h_s_dadda_rca32_fa268_y2, h_s_dadda_rca32_fa268_y4);
  fa fa_h_s_dadda_rca32_fa269_y2(h_s_dadda_rca32_fa268_y4, h_s_dadda_rca32_fa267_y4, h_s_dadda_rca32_fa266_y4, h_s_dadda_rca32_fa269_y2, h_s_dadda_rca32_fa269_y4);
  fa fa_h_s_dadda_rca32_fa270_y2(h_s_dadda_rca32_fa265_y4, h_s_dadda_rca32_fa264_y4, h_s_dadda_rca32_fa263_y4, h_s_dadda_rca32_fa270_y2, h_s_dadda_rca32_fa270_y4);
  fa fa_h_s_dadda_rca32_fa271_y2(h_s_dadda_rca32_fa262_y4, h_s_dadda_rca32_fa261_y4, h_s_dadda_rca32_fa260_y4, h_s_dadda_rca32_fa271_y2, h_s_dadda_rca32_fa271_y4);
  fa fa_h_s_dadda_rca32_fa272_y2(h_s_dadda_rca32_fa259_y4, h_s_dadda_rca32_fa258_y4, h_s_dadda_rca32_fa257_y4, h_s_dadda_rca32_fa272_y2, h_s_dadda_rca32_fa272_y4);
  fa fa_h_s_dadda_rca32_fa273_y2(h_s_dadda_rca32_fa256_y4, h_s_dadda_rca32_fa255_y4, h_s_dadda_rca32_fa254_y4, h_s_dadda_rca32_fa273_y2, h_s_dadda_rca32_fa273_y4);
  fa fa_h_s_dadda_rca32_fa274_y2(h_s_dadda_rca32_fa253_y4, h_s_dadda_rca32_fa252_y4, h_s_dadda_rca32_fa251_y4, h_s_dadda_rca32_fa274_y2, h_s_dadda_rca32_fa274_y4);
  fa fa_h_s_dadda_rca32_fa275_y2(h_s_dadda_rca32_fa250_y4, h_s_dadda_rca32_fa249_y4, h_s_dadda_rca32_fa248_y4, h_s_dadda_rca32_fa275_y2, h_s_dadda_rca32_fa275_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_4_y0(a_25, b_4, h_s_dadda_rca32_and_25_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_5_y0(a_24, b_5, h_s_dadda_rca32_and_24_5_y0);
  fa fa_h_s_dadda_rca32_fa276_y2(h_s_dadda_rca32_fa247_y4, h_s_dadda_rca32_and_25_4_y0, h_s_dadda_rca32_and_24_5_y0, h_s_dadda_rca32_fa276_y2, h_s_dadda_rca32_fa276_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_6_y0(a_23, b_6, h_s_dadda_rca32_and_23_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_7_y0(a_22, b_7, h_s_dadda_rca32_and_22_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_8_y0(a_21, b_8, h_s_dadda_rca32_and_21_8_y0);
  fa fa_h_s_dadda_rca32_fa277_y2(h_s_dadda_rca32_and_23_6_y0, h_s_dadda_rca32_and_22_7_y0, h_s_dadda_rca32_and_21_8_y0, h_s_dadda_rca32_fa277_y2, h_s_dadda_rca32_fa277_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_9_y0(a_20, b_9, h_s_dadda_rca32_and_20_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_10_y0(a_19, b_10, h_s_dadda_rca32_and_19_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_11_y0(a_18, b_11, h_s_dadda_rca32_and_18_11_y0);
  fa fa_h_s_dadda_rca32_fa278_y2(h_s_dadda_rca32_and_20_9_y0, h_s_dadda_rca32_and_19_10_y0, h_s_dadda_rca32_and_18_11_y0, h_s_dadda_rca32_fa278_y2, h_s_dadda_rca32_fa278_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_12_y0(a_17, b_12, h_s_dadda_rca32_and_17_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_13_y0(a_16, b_13, h_s_dadda_rca32_and_16_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_14_y0(a_15, b_14, h_s_dadda_rca32_and_15_14_y0);
  fa fa_h_s_dadda_rca32_fa279_y2(h_s_dadda_rca32_and_17_12_y0, h_s_dadda_rca32_and_16_13_y0, h_s_dadda_rca32_and_15_14_y0, h_s_dadda_rca32_fa279_y2, h_s_dadda_rca32_fa279_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_15_y0(a_14, b_15, h_s_dadda_rca32_and_14_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_16_y0(a_13, b_16, h_s_dadda_rca32_and_13_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_17_y0(a_12, b_17, h_s_dadda_rca32_and_12_17_y0);
  fa fa_h_s_dadda_rca32_fa280_y2(h_s_dadda_rca32_and_14_15_y0, h_s_dadda_rca32_and_13_16_y0, h_s_dadda_rca32_and_12_17_y0, h_s_dadda_rca32_fa280_y2, h_s_dadda_rca32_fa280_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_18_y0(a_11, b_18, h_s_dadda_rca32_and_11_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_19_y0(a_10, b_19, h_s_dadda_rca32_and_10_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_20_y0(a_9, b_20, h_s_dadda_rca32_and_9_20_y0);
  fa fa_h_s_dadda_rca32_fa281_y2(h_s_dadda_rca32_and_11_18_y0, h_s_dadda_rca32_and_10_19_y0, h_s_dadda_rca32_and_9_20_y0, h_s_dadda_rca32_fa281_y2, h_s_dadda_rca32_fa281_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_21_y0(a_8, b_21, h_s_dadda_rca32_and_8_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_22_y0(a_7, b_22, h_s_dadda_rca32_and_7_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_23_y0(a_6, b_23, h_s_dadda_rca32_and_6_23_y0);
  fa fa_h_s_dadda_rca32_fa282_y2(h_s_dadda_rca32_and_8_21_y0, h_s_dadda_rca32_and_7_22_y0, h_s_dadda_rca32_and_6_23_y0, h_s_dadda_rca32_fa282_y2, h_s_dadda_rca32_fa282_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_24_y0(a_5, b_24, h_s_dadda_rca32_and_5_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_25_y0(a_4, b_25, h_s_dadda_rca32_and_4_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_26_y0(a_3, b_26, h_s_dadda_rca32_and_3_26_y0);
  fa fa_h_s_dadda_rca32_fa283_y2(h_s_dadda_rca32_and_5_24_y0, h_s_dadda_rca32_and_4_25_y0, h_s_dadda_rca32_and_3_26_y0, h_s_dadda_rca32_fa283_y2, h_s_dadda_rca32_fa283_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_27_y0(a_2, b_27, h_s_dadda_rca32_and_2_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_28_y0(a_1, b_28, h_s_dadda_rca32_and_1_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_29_y0(a_0, b_29, h_s_dadda_rca32_and_0_29_y0);
  fa fa_h_s_dadda_rca32_fa284_y2(h_s_dadda_rca32_and_2_27_y0, h_s_dadda_rca32_and_1_28_y0, h_s_dadda_rca32_and_0_29_y0, h_s_dadda_rca32_fa284_y2, h_s_dadda_rca32_fa284_y4);
  fa fa_h_s_dadda_rca32_fa285_y2(h_s_dadda_rca32_fa0_y2, h_s_dadda_rca32_ha1_y0, h_s_dadda_rca32_fa269_y2, h_s_dadda_rca32_fa285_y2, h_s_dadda_rca32_fa285_y4);
  fa fa_h_s_dadda_rca32_fa286_y2(h_s_dadda_rca32_fa270_y2, h_s_dadda_rca32_fa271_y2, h_s_dadda_rca32_fa272_y2, h_s_dadda_rca32_fa286_y2, h_s_dadda_rca32_fa286_y4);
  fa fa_h_s_dadda_rca32_fa287_y2(h_s_dadda_rca32_fa273_y2, h_s_dadda_rca32_fa274_y2, h_s_dadda_rca32_fa275_y2, h_s_dadda_rca32_fa287_y2, h_s_dadda_rca32_fa287_y4);
  fa fa_h_s_dadda_rca32_fa288_y2(h_s_dadda_rca32_fa276_y2, h_s_dadda_rca32_fa277_y2, h_s_dadda_rca32_fa278_y2, h_s_dadda_rca32_fa288_y2, h_s_dadda_rca32_fa288_y4);
  fa fa_h_s_dadda_rca32_fa289_y2(h_s_dadda_rca32_fa279_y2, h_s_dadda_rca32_fa280_y2, h_s_dadda_rca32_fa281_y2, h_s_dadda_rca32_fa289_y2, h_s_dadda_rca32_fa289_y4);
  fa fa_h_s_dadda_rca32_fa290_y2(h_s_dadda_rca32_fa282_y2, h_s_dadda_rca32_fa283_y2, h_s_dadda_rca32_fa284_y2, h_s_dadda_rca32_fa290_y2, h_s_dadda_rca32_fa290_y4);
  fa fa_h_s_dadda_rca32_fa291_y2(h_s_dadda_rca32_fa290_y4, h_s_dadda_rca32_fa289_y4, h_s_dadda_rca32_fa288_y4, h_s_dadda_rca32_fa291_y2, h_s_dadda_rca32_fa291_y4);
  fa fa_h_s_dadda_rca32_fa292_y2(h_s_dadda_rca32_fa287_y4, h_s_dadda_rca32_fa286_y4, h_s_dadda_rca32_fa285_y4, h_s_dadda_rca32_fa292_y2, h_s_dadda_rca32_fa292_y4);
  fa fa_h_s_dadda_rca32_fa293_y2(h_s_dadda_rca32_fa284_y4, h_s_dadda_rca32_fa283_y4, h_s_dadda_rca32_fa282_y4, h_s_dadda_rca32_fa293_y2, h_s_dadda_rca32_fa293_y4);
  fa fa_h_s_dadda_rca32_fa294_y2(h_s_dadda_rca32_fa281_y4, h_s_dadda_rca32_fa280_y4, h_s_dadda_rca32_fa279_y4, h_s_dadda_rca32_fa294_y2, h_s_dadda_rca32_fa294_y4);
  fa fa_h_s_dadda_rca32_fa295_y2(h_s_dadda_rca32_fa278_y4, h_s_dadda_rca32_fa277_y4, h_s_dadda_rca32_fa276_y4, h_s_dadda_rca32_fa295_y2, h_s_dadda_rca32_fa295_y4);
  fa fa_h_s_dadda_rca32_fa296_y2(h_s_dadda_rca32_fa275_y4, h_s_dadda_rca32_fa274_y4, h_s_dadda_rca32_fa273_y4, h_s_dadda_rca32_fa296_y2, h_s_dadda_rca32_fa296_y4);
  fa fa_h_s_dadda_rca32_fa297_y2(h_s_dadda_rca32_fa272_y4, h_s_dadda_rca32_fa271_y4, h_s_dadda_rca32_fa270_y4, h_s_dadda_rca32_fa297_y2, h_s_dadda_rca32_fa297_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_6_y0(a_24, b_6, h_s_dadda_rca32_and_24_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_7_y0(a_23, b_7, h_s_dadda_rca32_and_23_7_y0);
  fa fa_h_s_dadda_rca32_fa298_y2(h_s_dadda_rca32_fa269_y4, h_s_dadda_rca32_and_24_6_y0, h_s_dadda_rca32_and_23_7_y0, h_s_dadda_rca32_fa298_y2, h_s_dadda_rca32_fa298_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_8_y0(a_22, b_8, h_s_dadda_rca32_and_22_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_9_y0(a_21, b_9, h_s_dadda_rca32_and_21_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_10_y0(a_20, b_10, h_s_dadda_rca32_and_20_10_y0);
  fa fa_h_s_dadda_rca32_fa299_y2(h_s_dadda_rca32_and_22_8_y0, h_s_dadda_rca32_and_21_9_y0, h_s_dadda_rca32_and_20_10_y0, h_s_dadda_rca32_fa299_y2, h_s_dadda_rca32_fa299_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_11_y0(a_19, b_11, h_s_dadda_rca32_and_19_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_12_y0(a_18, b_12, h_s_dadda_rca32_and_18_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_13_y0(a_17, b_13, h_s_dadda_rca32_and_17_13_y0);
  fa fa_h_s_dadda_rca32_fa300_y2(h_s_dadda_rca32_and_19_11_y0, h_s_dadda_rca32_and_18_12_y0, h_s_dadda_rca32_and_17_13_y0, h_s_dadda_rca32_fa300_y2, h_s_dadda_rca32_fa300_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_14_y0(a_16, b_14, h_s_dadda_rca32_and_16_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_15_y0(a_15, b_15, h_s_dadda_rca32_and_15_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_16_y0(a_14, b_16, h_s_dadda_rca32_and_14_16_y0);
  fa fa_h_s_dadda_rca32_fa301_y2(h_s_dadda_rca32_and_16_14_y0, h_s_dadda_rca32_and_15_15_y0, h_s_dadda_rca32_and_14_16_y0, h_s_dadda_rca32_fa301_y2, h_s_dadda_rca32_fa301_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_17_y0(a_13, b_17, h_s_dadda_rca32_and_13_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_18_y0(a_12, b_18, h_s_dadda_rca32_and_12_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_19_y0(a_11, b_19, h_s_dadda_rca32_and_11_19_y0);
  fa fa_h_s_dadda_rca32_fa302_y2(h_s_dadda_rca32_and_13_17_y0, h_s_dadda_rca32_and_12_18_y0, h_s_dadda_rca32_and_11_19_y0, h_s_dadda_rca32_fa302_y2, h_s_dadda_rca32_fa302_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_20_y0(a_10, b_20, h_s_dadda_rca32_and_10_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_21_y0(a_9, b_21, h_s_dadda_rca32_and_9_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_22_y0(a_8, b_22, h_s_dadda_rca32_and_8_22_y0);
  fa fa_h_s_dadda_rca32_fa303_y2(h_s_dadda_rca32_and_10_20_y0, h_s_dadda_rca32_and_9_21_y0, h_s_dadda_rca32_and_8_22_y0, h_s_dadda_rca32_fa303_y2, h_s_dadda_rca32_fa303_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_23_y0(a_7, b_23, h_s_dadda_rca32_and_7_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_24_y0(a_6, b_24, h_s_dadda_rca32_and_6_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_25_y0(a_5, b_25, h_s_dadda_rca32_and_5_25_y0);
  fa fa_h_s_dadda_rca32_fa304_y2(h_s_dadda_rca32_and_7_23_y0, h_s_dadda_rca32_and_6_24_y0, h_s_dadda_rca32_and_5_25_y0, h_s_dadda_rca32_fa304_y2, h_s_dadda_rca32_fa304_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_26_y0(a_4, b_26, h_s_dadda_rca32_and_4_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_27_y0(a_3, b_27, h_s_dadda_rca32_and_3_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_28_y0(a_2, b_28, h_s_dadda_rca32_and_2_28_y0);
  fa fa_h_s_dadda_rca32_fa305_y2(h_s_dadda_rca32_and_4_26_y0, h_s_dadda_rca32_and_3_27_y0, h_s_dadda_rca32_and_2_28_y0, h_s_dadda_rca32_fa305_y2, h_s_dadda_rca32_fa305_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_29_y0(a_1, b_29, h_s_dadda_rca32_and_1_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_30_y0(a_0, b_30, h_s_dadda_rca32_and_0_30_y0);
  fa fa_h_s_dadda_rca32_fa306_y2(h_s_dadda_rca32_and_1_29_y0, h_s_dadda_rca32_and_0_30_y0, h_s_dadda_rca32_fa1_y2, h_s_dadda_rca32_fa306_y2, h_s_dadda_rca32_fa306_y4);
  fa fa_h_s_dadda_rca32_fa307_y2(h_s_dadda_rca32_fa2_y2, h_s_dadda_rca32_ha2_y0, h_s_dadda_rca32_fa291_y2, h_s_dadda_rca32_fa307_y2, h_s_dadda_rca32_fa307_y4);
  fa fa_h_s_dadda_rca32_fa308_y2(h_s_dadda_rca32_fa292_y2, h_s_dadda_rca32_fa293_y2, h_s_dadda_rca32_fa294_y2, h_s_dadda_rca32_fa308_y2, h_s_dadda_rca32_fa308_y4);
  fa fa_h_s_dadda_rca32_fa309_y2(h_s_dadda_rca32_fa295_y2, h_s_dadda_rca32_fa296_y2, h_s_dadda_rca32_fa297_y2, h_s_dadda_rca32_fa309_y2, h_s_dadda_rca32_fa309_y4);
  fa fa_h_s_dadda_rca32_fa310_y2(h_s_dadda_rca32_fa298_y2, h_s_dadda_rca32_fa299_y2, h_s_dadda_rca32_fa300_y2, h_s_dadda_rca32_fa310_y2, h_s_dadda_rca32_fa310_y4);
  fa fa_h_s_dadda_rca32_fa311_y2(h_s_dadda_rca32_fa301_y2, h_s_dadda_rca32_fa302_y2, h_s_dadda_rca32_fa303_y2, h_s_dadda_rca32_fa311_y2, h_s_dadda_rca32_fa311_y4);
  fa fa_h_s_dadda_rca32_fa312_y2(h_s_dadda_rca32_fa304_y2, h_s_dadda_rca32_fa305_y2, h_s_dadda_rca32_fa306_y2, h_s_dadda_rca32_fa312_y2, h_s_dadda_rca32_fa312_y4);
  fa fa_h_s_dadda_rca32_fa313_y2(h_s_dadda_rca32_fa312_y4, h_s_dadda_rca32_fa311_y4, h_s_dadda_rca32_fa310_y4, h_s_dadda_rca32_fa313_y2, h_s_dadda_rca32_fa313_y4);
  fa fa_h_s_dadda_rca32_fa314_y2(h_s_dadda_rca32_fa309_y4, h_s_dadda_rca32_fa308_y4, h_s_dadda_rca32_fa307_y4, h_s_dadda_rca32_fa314_y2, h_s_dadda_rca32_fa314_y4);
  fa fa_h_s_dadda_rca32_fa315_y2(h_s_dadda_rca32_fa306_y4, h_s_dadda_rca32_fa305_y4, h_s_dadda_rca32_fa304_y4, h_s_dadda_rca32_fa315_y2, h_s_dadda_rca32_fa315_y4);
  fa fa_h_s_dadda_rca32_fa316_y2(h_s_dadda_rca32_fa303_y4, h_s_dadda_rca32_fa302_y4, h_s_dadda_rca32_fa301_y4, h_s_dadda_rca32_fa316_y2, h_s_dadda_rca32_fa316_y4);
  fa fa_h_s_dadda_rca32_fa317_y2(h_s_dadda_rca32_fa300_y4, h_s_dadda_rca32_fa299_y4, h_s_dadda_rca32_fa298_y4, h_s_dadda_rca32_fa317_y2, h_s_dadda_rca32_fa317_y4);
  fa fa_h_s_dadda_rca32_fa318_y2(h_s_dadda_rca32_fa297_y4, h_s_dadda_rca32_fa296_y4, h_s_dadda_rca32_fa295_y4, h_s_dadda_rca32_fa318_y2, h_s_dadda_rca32_fa318_y4);
  fa fa_h_s_dadda_rca32_fa319_y2(h_s_dadda_rca32_fa294_y4, h_s_dadda_rca32_fa293_y4, h_s_dadda_rca32_fa292_y4, h_s_dadda_rca32_fa319_y2, h_s_dadda_rca32_fa319_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_8_y0(a_23, b_8, h_s_dadda_rca32_and_23_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_9_y0(a_22, b_9, h_s_dadda_rca32_and_22_9_y0);
  fa fa_h_s_dadda_rca32_fa320_y2(h_s_dadda_rca32_fa291_y4, h_s_dadda_rca32_and_23_8_y0, h_s_dadda_rca32_and_22_9_y0, h_s_dadda_rca32_fa320_y2, h_s_dadda_rca32_fa320_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_10_y0(a_21, b_10, h_s_dadda_rca32_and_21_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_11_y0(a_20, b_11, h_s_dadda_rca32_and_20_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_12_y0(a_19, b_12, h_s_dadda_rca32_and_19_12_y0);
  fa fa_h_s_dadda_rca32_fa321_y2(h_s_dadda_rca32_and_21_10_y0, h_s_dadda_rca32_and_20_11_y0, h_s_dadda_rca32_and_19_12_y0, h_s_dadda_rca32_fa321_y2, h_s_dadda_rca32_fa321_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_13_y0(a_18, b_13, h_s_dadda_rca32_and_18_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_14_y0(a_17, b_14, h_s_dadda_rca32_and_17_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_15_y0(a_16, b_15, h_s_dadda_rca32_and_16_15_y0);
  fa fa_h_s_dadda_rca32_fa322_y2(h_s_dadda_rca32_and_18_13_y0, h_s_dadda_rca32_and_17_14_y0, h_s_dadda_rca32_and_16_15_y0, h_s_dadda_rca32_fa322_y2, h_s_dadda_rca32_fa322_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_16_y0(a_15, b_16, h_s_dadda_rca32_and_15_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_17_y0(a_14, b_17, h_s_dadda_rca32_and_14_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_18_y0(a_13, b_18, h_s_dadda_rca32_and_13_18_y0);
  fa fa_h_s_dadda_rca32_fa323_y2(h_s_dadda_rca32_and_15_16_y0, h_s_dadda_rca32_and_14_17_y0, h_s_dadda_rca32_and_13_18_y0, h_s_dadda_rca32_fa323_y2, h_s_dadda_rca32_fa323_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_19_y0(a_12, b_19, h_s_dadda_rca32_and_12_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_20_y0(a_11, b_20, h_s_dadda_rca32_and_11_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_21_y0(a_10, b_21, h_s_dadda_rca32_and_10_21_y0);
  fa fa_h_s_dadda_rca32_fa324_y2(h_s_dadda_rca32_and_12_19_y0, h_s_dadda_rca32_and_11_20_y0, h_s_dadda_rca32_and_10_21_y0, h_s_dadda_rca32_fa324_y2, h_s_dadda_rca32_fa324_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_22_y0(a_9, b_22, h_s_dadda_rca32_and_9_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_23_y0(a_8, b_23, h_s_dadda_rca32_and_8_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_24_y0(a_7, b_24, h_s_dadda_rca32_and_7_24_y0);
  fa fa_h_s_dadda_rca32_fa325_y2(h_s_dadda_rca32_and_9_22_y0, h_s_dadda_rca32_and_8_23_y0, h_s_dadda_rca32_and_7_24_y0, h_s_dadda_rca32_fa325_y2, h_s_dadda_rca32_fa325_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_25_y0(a_6, b_25, h_s_dadda_rca32_and_6_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_26_y0(a_5, b_26, h_s_dadda_rca32_and_5_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_27_y0(a_4, b_27, h_s_dadda_rca32_and_4_27_y0);
  fa fa_h_s_dadda_rca32_fa326_y2(h_s_dadda_rca32_and_6_25_y0, h_s_dadda_rca32_and_5_26_y0, h_s_dadda_rca32_and_4_27_y0, h_s_dadda_rca32_fa326_y2, h_s_dadda_rca32_fa326_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_28_y0(a_3, b_28, h_s_dadda_rca32_and_3_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_29_y0(a_2, b_29, h_s_dadda_rca32_and_2_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_30_y0(a_1, b_30, h_s_dadda_rca32_and_1_30_y0);
  fa fa_h_s_dadda_rca32_fa327_y2(h_s_dadda_rca32_and_3_28_y0, h_s_dadda_rca32_and_2_29_y0, h_s_dadda_rca32_and_1_30_y0, h_s_dadda_rca32_fa327_y2, h_s_dadda_rca32_fa327_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_0_31_y0(a_0, b_31, h_s_dadda_rca32_nand_0_31_y0);
  fa fa_h_s_dadda_rca32_fa328_y2(h_s_dadda_rca32_nand_0_31_y0, h_s_dadda_rca32_fa3_y2, h_s_dadda_rca32_fa4_y2, h_s_dadda_rca32_fa328_y2, h_s_dadda_rca32_fa328_y4);
  fa fa_h_s_dadda_rca32_fa329_y2(h_s_dadda_rca32_fa5_y2, h_s_dadda_rca32_ha3_y0, h_s_dadda_rca32_fa313_y2, h_s_dadda_rca32_fa329_y2, h_s_dadda_rca32_fa329_y4);
  fa fa_h_s_dadda_rca32_fa330_y2(h_s_dadda_rca32_fa314_y2, h_s_dadda_rca32_fa315_y2, h_s_dadda_rca32_fa316_y2, h_s_dadda_rca32_fa330_y2, h_s_dadda_rca32_fa330_y4);
  fa fa_h_s_dadda_rca32_fa331_y2(h_s_dadda_rca32_fa317_y2, h_s_dadda_rca32_fa318_y2, h_s_dadda_rca32_fa319_y2, h_s_dadda_rca32_fa331_y2, h_s_dadda_rca32_fa331_y4);
  fa fa_h_s_dadda_rca32_fa332_y2(h_s_dadda_rca32_fa320_y2, h_s_dadda_rca32_fa321_y2, h_s_dadda_rca32_fa322_y2, h_s_dadda_rca32_fa332_y2, h_s_dadda_rca32_fa332_y4);
  fa fa_h_s_dadda_rca32_fa333_y2(h_s_dadda_rca32_fa323_y2, h_s_dadda_rca32_fa324_y2, h_s_dadda_rca32_fa325_y2, h_s_dadda_rca32_fa333_y2, h_s_dadda_rca32_fa333_y4);
  fa fa_h_s_dadda_rca32_fa334_y2(h_s_dadda_rca32_fa326_y2, h_s_dadda_rca32_fa327_y2, h_s_dadda_rca32_fa328_y2, h_s_dadda_rca32_fa334_y2, h_s_dadda_rca32_fa334_y4);
  fa fa_h_s_dadda_rca32_fa335_y2(h_s_dadda_rca32_fa334_y4, h_s_dadda_rca32_fa333_y4, h_s_dadda_rca32_fa332_y4, h_s_dadda_rca32_fa335_y2, h_s_dadda_rca32_fa335_y4);
  fa fa_h_s_dadda_rca32_fa336_y2(h_s_dadda_rca32_fa331_y4, h_s_dadda_rca32_fa330_y4, h_s_dadda_rca32_fa329_y4, h_s_dadda_rca32_fa336_y2, h_s_dadda_rca32_fa336_y4);
  fa fa_h_s_dadda_rca32_fa337_y2(h_s_dadda_rca32_fa328_y4, h_s_dadda_rca32_fa327_y4, h_s_dadda_rca32_fa326_y4, h_s_dadda_rca32_fa337_y2, h_s_dadda_rca32_fa337_y4);
  fa fa_h_s_dadda_rca32_fa338_y2(h_s_dadda_rca32_fa325_y4, h_s_dadda_rca32_fa324_y4, h_s_dadda_rca32_fa323_y4, h_s_dadda_rca32_fa338_y2, h_s_dadda_rca32_fa338_y4);
  fa fa_h_s_dadda_rca32_fa339_y2(h_s_dadda_rca32_fa322_y4, h_s_dadda_rca32_fa321_y4, h_s_dadda_rca32_fa320_y4, h_s_dadda_rca32_fa339_y2, h_s_dadda_rca32_fa339_y4);
  fa fa_h_s_dadda_rca32_fa340_y2(h_s_dadda_rca32_fa319_y4, h_s_dadda_rca32_fa318_y4, h_s_dadda_rca32_fa317_y4, h_s_dadda_rca32_fa340_y2, h_s_dadda_rca32_fa340_y4);
  fa fa_h_s_dadda_rca32_fa341_y2(h_s_dadda_rca32_fa316_y4, h_s_dadda_rca32_fa315_y4, h_s_dadda_rca32_fa314_y4, h_s_dadda_rca32_fa341_y2, h_s_dadda_rca32_fa341_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_8_y0(a_24, b_8, h_s_dadda_rca32_and_24_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_9_y0(a_23, b_9, h_s_dadda_rca32_and_23_9_y0);
  fa fa_h_s_dadda_rca32_fa342_y2(h_s_dadda_rca32_fa313_y4, h_s_dadda_rca32_and_24_8_y0, h_s_dadda_rca32_and_23_9_y0, h_s_dadda_rca32_fa342_y2, h_s_dadda_rca32_fa342_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_10_y0(a_22, b_10, h_s_dadda_rca32_and_22_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_11_y0(a_21, b_11, h_s_dadda_rca32_and_21_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_12_y0(a_20, b_12, h_s_dadda_rca32_and_20_12_y0);
  fa fa_h_s_dadda_rca32_fa343_y2(h_s_dadda_rca32_and_22_10_y0, h_s_dadda_rca32_and_21_11_y0, h_s_dadda_rca32_and_20_12_y0, h_s_dadda_rca32_fa343_y2, h_s_dadda_rca32_fa343_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_13_y0(a_19, b_13, h_s_dadda_rca32_and_19_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_14_y0(a_18, b_14, h_s_dadda_rca32_and_18_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_15_y0(a_17, b_15, h_s_dadda_rca32_and_17_15_y0);
  fa fa_h_s_dadda_rca32_fa344_y2(h_s_dadda_rca32_and_19_13_y0, h_s_dadda_rca32_and_18_14_y0, h_s_dadda_rca32_and_17_15_y0, h_s_dadda_rca32_fa344_y2, h_s_dadda_rca32_fa344_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_16_y0(a_16, b_16, h_s_dadda_rca32_and_16_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_17_y0(a_15, b_17, h_s_dadda_rca32_and_15_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_18_y0(a_14, b_18, h_s_dadda_rca32_and_14_18_y0);
  fa fa_h_s_dadda_rca32_fa345_y2(h_s_dadda_rca32_and_16_16_y0, h_s_dadda_rca32_and_15_17_y0, h_s_dadda_rca32_and_14_18_y0, h_s_dadda_rca32_fa345_y2, h_s_dadda_rca32_fa345_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_19_y0(a_13, b_19, h_s_dadda_rca32_and_13_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_20_y0(a_12, b_20, h_s_dadda_rca32_and_12_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_21_y0(a_11, b_21, h_s_dadda_rca32_and_11_21_y0);
  fa fa_h_s_dadda_rca32_fa346_y2(h_s_dadda_rca32_and_13_19_y0, h_s_dadda_rca32_and_12_20_y0, h_s_dadda_rca32_and_11_21_y0, h_s_dadda_rca32_fa346_y2, h_s_dadda_rca32_fa346_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_22_y0(a_10, b_22, h_s_dadda_rca32_and_10_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_23_y0(a_9, b_23, h_s_dadda_rca32_and_9_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_24_y0(a_8, b_24, h_s_dadda_rca32_and_8_24_y0);
  fa fa_h_s_dadda_rca32_fa347_y2(h_s_dadda_rca32_and_10_22_y0, h_s_dadda_rca32_and_9_23_y0, h_s_dadda_rca32_and_8_24_y0, h_s_dadda_rca32_fa347_y2, h_s_dadda_rca32_fa347_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_25_y0(a_7, b_25, h_s_dadda_rca32_and_7_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_26_y0(a_6, b_26, h_s_dadda_rca32_and_6_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_27_y0(a_5, b_27, h_s_dadda_rca32_and_5_27_y0);
  fa fa_h_s_dadda_rca32_fa348_y2(h_s_dadda_rca32_and_7_25_y0, h_s_dadda_rca32_and_6_26_y0, h_s_dadda_rca32_and_5_27_y0, h_s_dadda_rca32_fa348_y2, h_s_dadda_rca32_fa348_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_28_y0(a_4, b_28, h_s_dadda_rca32_and_4_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_29_y0(a_3, b_29, h_s_dadda_rca32_and_3_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_30_y0(a_2, b_30, h_s_dadda_rca32_and_2_30_y0);
  fa fa_h_s_dadda_rca32_fa349_y2(h_s_dadda_rca32_and_4_28_y0, h_s_dadda_rca32_and_3_29_y0, h_s_dadda_rca32_and_2_30_y0, h_s_dadda_rca32_fa349_y2, h_s_dadda_rca32_fa349_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_1_31_y0(a_1, b_31, h_s_dadda_rca32_nand_1_31_y0);
  fa fa_h_s_dadda_rca32_fa350_y2(h_s_dadda_rca32_nand_1_31_y0, h_s_dadda_rca32_fa6_y2, h_s_dadda_rca32_fa7_y2, h_s_dadda_rca32_fa350_y2, h_s_dadda_rca32_fa350_y4);
  fa fa_h_s_dadda_rca32_fa351_y2(h_s_dadda_rca32_fa8_y2, h_s_dadda_rca32_fa9_y2, h_s_dadda_rca32_fa335_y2, h_s_dadda_rca32_fa351_y2, h_s_dadda_rca32_fa351_y4);
  fa fa_h_s_dadda_rca32_fa352_y2(h_s_dadda_rca32_fa336_y2, h_s_dadda_rca32_fa337_y2, h_s_dadda_rca32_fa338_y2, h_s_dadda_rca32_fa352_y2, h_s_dadda_rca32_fa352_y4);
  fa fa_h_s_dadda_rca32_fa353_y2(h_s_dadda_rca32_fa339_y2, h_s_dadda_rca32_fa340_y2, h_s_dadda_rca32_fa341_y2, h_s_dadda_rca32_fa353_y2, h_s_dadda_rca32_fa353_y4);
  fa fa_h_s_dadda_rca32_fa354_y2(h_s_dadda_rca32_fa342_y2, h_s_dadda_rca32_fa343_y2, h_s_dadda_rca32_fa344_y2, h_s_dadda_rca32_fa354_y2, h_s_dadda_rca32_fa354_y4);
  fa fa_h_s_dadda_rca32_fa355_y2(h_s_dadda_rca32_fa345_y2, h_s_dadda_rca32_fa346_y2, h_s_dadda_rca32_fa347_y2, h_s_dadda_rca32_fa355_y2, h_s_dadda_rca32_fa355_y4);
  fa fa_h_s_dadda_rca32_fa356_y2(h_s_dadda_rca32_fa348_y2, h_s_dadda_rca32_fa349_y2, h_s_dadda_rca32_fa350_y2, h_s_dadda_rca32_fa356_y2, h_s_dadda_rca32_fa356_y4);
  fa fa_h_s_dadda_rca32_fa357_y2(h_s_dadda_rca32_fa356_y4, h_s_dadda_rca32_fa355_y4, h_s_dadda_rca32_fa354_y4, h_s_dadda_rca32_fa357_y2, h_s_dadda_rca32_fa357_y4);
  fa fa_h_s_dadda_rca32_fa358_y2(h_s_dadda_rca32_fa353_y4, h_s_dadda_rca32_fa352_y4, h_s_dadda_rca32_fa351_y4, h_s_dadda_rca32_fa358_y2, h_s_dadda_rca32_fa358_y4);
  fa fa_h_s_dadda_rca32_fa359_y2(h_s_dadda_rca32_fa350_y4, h_s_dadda_rca32_fa349_y4, h_s_dadda_rca32_fa348_y4, h_s_dadda_rca32_fa359_y2, h_s_dadda_rca32_fa359_y4);
  fa fa_h_s_dadda_rca32_fa360_y2(h_s_dadda_rca32_fa347_y4, h_s_dadda_rca32_fa346_y4, h_s_dadda_rca32_fa345_y4, h_s_dadda_rca32_fa360_y2, h_s_dadda_rca32_fa360_y4);
  fa fa_h_s_dadda_rca32_fa361_y2(h_s_dadda_rca32_fa344_y4, h_s_dadda_rca32_fa343_y4, h_s_dadda_rca32_fa342_y4, h_s_dadda_rca32_fa361_y2, h_s_dadda_rca32_fa361_y4);
  fa fa_h_s_dadda_rca32_fa362_y2(h_s_dadda_rca32_fa341_y4, h_s_dadda_rca32_fa340_y4, h_s_dadda_rca32_fa339_y4, h_s_dadda_rca32_fa362_y2, h_s_dadda_rca32_fa362_y4);
  fa fa_h_s_dadda_rca32_fa363_y2(h_s_dadda_rca32_fa338_y4, h_s_dadda_rca32_fa337_y4, h_s_dadda_rca32_fa336_y4, h_s_dadda_rca32_fa363_y2, h_s_dadda_rca32_fa363_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_7_y0(a_26, b_7, h_s_dadda_rca32_and_26_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_8_y0(a_25, b_8, h_s_dadda_rca32_and_25_8_y0);
  fa fa_h_s_dadda_rca32_fa364_y2(h_s_dadda_rca32_fa335_y4, h_s_dadda_rca32_and_26_7_y0, h_s_dadda_rca32_and_25_8_y0, h_s_dadda_rca32_fa364_y2, h_s_dadda_rca32_fa364_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_9_y0(a_24, b_9, h_s_dadda_rca32_and_24_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_10_y0(a_23, b_10, h_s_dadda_rca32_and_23_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_11_y0(a_22, b_11, h_s_dadda_rca32_and_22_11_y0);
  fa fa_h_s_dadda_rca32_fa365_y2(h_s_dadda_rca32_and_24_9_y0, h_s_dadda_rca32_and_23_10_y0, h_s_dadda_rca32_and_22_11_y0, h_s_dadda_rca32_fa365_y2, h_s_dadda_rca32_fa365_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_12_y0(a_21, b_12, h_s_dadda_rca32_and_21_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_13_y0(a_20, b_13, h_s_dadda_rca32_and_20_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_14_y0(a_19, b_14, h_s_dadda_rca32_and_19_14_y0);
  fa fa_h_s_dadda_rca32_fa366_y2(h_s_dadda_rca32_and_21_12_y0, h_s_dadda_rca32_and_20_13_y0, h_s_dadda_rca32_and_19_14_y0, h_s_dadda_rca32_fa366_y2, h_s_dadda_rca32_fa366_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_15_y0(a_18, b_15, h_s_dadda_rca32_and_18_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_16_y0(a_17, b_16, h_s_dadda_rca32_and_17_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_17_y0(a_16, b_17, h_s_dadda_rca32_and_16_17_y0);
  fa fa_h_s_dadda_rca32_fa367_y2(h_s_dadda_rca32_and_18_15_y0, h_s_dadda_rca32_and_17_16_y0, h_s_dadda_rca32_and_16_17_y0, h_s_dadda_rca32_fa367_y2, h_s_dadda_rca32_fa367_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_18_y0(a_15, b_18, h_s_dadda_rca32_and_15_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_19_y0(a_14, b_19, h_s_dadda_rca32_and_14_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_20_y0(a_13, b_20, h_s_dadda_rca32_and_13_20_y0);
  fa fa_h_s_dadda_rca32_fa368_y2(h_s_dadda_rca32_and_15_18_y0, h_s_dadda_rca32_and_14_19_y0, h_s_dadda_rca32_and_13_20_y0, h_s_dadda_rca32_fa368_y2, h_s_dadda_rca32_fa368_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_21_y0(a_12, b_21, h_s_dadda_rca32_and_12_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_22_y0(a_11, b_22, h_s_dadda_rca32_and_11_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_23_y0(a_10, b_23, h_s_dadda_rca32_and_10_23_y0);
  fa fa_h_s_dadda_rca32_fa369_y2(h_s_dadda_rca32_and_12_21_y0, h_s_dadda_rca32_and_11_22_y0, h_s_dadda_rca32_and_10_23_y0, h_s_dadda_rca32_fa369_y2, h_s_dadda_rca32_fa369_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_24_y0(a_9, b_24, h_s_dadda_rca32_and_9_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_25_y0(a_8, b_25, h_s_dadda_rca32_and_8_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_26_y0(a_7, b_26, h_s_dadda_rca32_and_7_26_y0);
  fa fa_h_s_dadda_rca32_fa370_y2(h_s_dadda_rca32_and_9_24_y0, h_s_dadda_rca32_and_8_25_y0, h_s_dadda_rca32_and_7_26_y0, h_s_dadda_rca32_fa370_y2, h_s_dadda_rca32_fa370_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_27_y0(a_6, b_27, h_s_dadda_rca32_and_6_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_28_y0(a_5, b_28, h_s_dadda_rca32_and_5_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_29_y0(a_4, b_29, h_s_dadda_rca32_and_4_29_y0);
  fa fa_h_s_dadda_rca32_fa371_y2(h_s_dadda_rca32_and_6_27_y0, h_s_dadda_rca32_and_5_28_y0, h_s_dadda_rca32_and_4_29_y0, h_s_dadda_rca32_fa371_y2, h_s_dadda_rca32_fa371_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_30_y0(a_3, b_30, h_s_dadda_rca32_and_3_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_2_31_y0(a_2, b_31, h_s_dadda_rca32_nand_2_31_y0);
  fa fa_h_s_dadda_rca32_fa372_y2(h_s_dadda_rca32_and_3_30_y0, h_s_dadda_rca32_nand_2_31_y0, h_s_dadda_rca32_fa10_y2, h_s_dadda_rca32_fa372_y2, h_s_dadda_rca32_fa372_y4);
  fa fa_h_s_dadda_rca32_fa373_y2(h_s_dadda_rca32_fa11_y2, h_s_dadda_rca32_fa12_y2, h_s_dadda_rca32_fa357_y2, h_s_dadda_rca32_fa373_y2, h_s_dadda_rca32_fa373_y4);
  fa fa_h_s_dadda_rca32_fa374_y2(h_s_dadda_rca32_fa358_y2, h_s_dadda_rca32_fa359_y2, h_s_dadda_rca32_fa360_y2, h_s_dadda_rca32_fa374_y2, h_s_dadda_rca32_fa374_y4);
  fa fa_h_s_dadda_rca32_fa375_y2(h_s_dadda_rca32_fa361_y2, h_s_dadda_rca32_fa362_y2, h_s_dadda_rca32_fa363_y2, h_s_dadda_rca32_fa375_y2, h_s_dadda_rca32_fa375_y4);
  fa fa_h_s_dadda_rca32_fa376_y2(h_s_dadda_rca32_fa364_y2, h_s_dadda_rca32_fa365_y2, h_s_dadda_rca32_fa366_y2, h_s_dadda_rca32_fa376_y2, h_s_dadda_rca32_fa376_y4);
  fa fa_h_s_dadda_rca32_fa377_y2(h_s_dadda_rca32_fa367_y2, h_s_dadda_rca32_fa368_y2, h_s_dadda_rca32_fa369_y2, h_s_dadda_rca32_fa377_y2, h_s_dadda_rca32_fa377_y4);
  fa fa_h_s_dadda_rca32_fa378_y2(h_s_dadda_rca32_fa370_y2, h_s_dadda_rca32_fa371_y2, h_s_dadda_rca32_fa372_y2, h_s_dadda_rca32_fa378_y2, h_s_dadda_rca32_fa378_y4);
  fa fa_h_s_dadda_rca32_fa379_y2(h_s_dadda_rca32_fa378_y4, h_s_dadda_rca32_fa377_y4, h_s_dadda_rca32_fa376_y4, h_s_dadda_rca32_fa379_y2, h_s_dadda_rca32_fa379_y4);
  fa fa_h_s_dadda_rca32_fa380_y2(h_s_dadda_rca32_fa375_y4, h_s_dadda_rca32_fa374_y4, h_s_dadda_rca32_fa373_y4, h_s_dadda_rca32_fa380_y2, h_s_dadda_rca32_fa380_y4);
  fa fa_h_s_dadda_rca32_fa381_y2(h_s_dadda_rca32_fa372_y4, h_s_dadda_rca32_fa371_y4, h_s_dadda_rca32_fa370_y4, h_s_dadda_rca32_fa381_y2, h_s_dadda_rca32_fa381_y4);
  fa fa_h_s_dadda_rca32_fa382_y2(h_s_dadda_rca32_fa369_y4, h_s_dadda_rca32_fa368_y4, h_s_dadda_rca32_fa367_y4, h_s_dadda_rca32_fa382_y2, h_s_dadda_rca32_fa382_y4);
  fa fa_h_s_dadda_rca32_fa383_y2(h_s_dadda_rca32_fa366_y4, h_s_dadda_rca32_fa365_y4, h_s_dadda_rca32_fa364_y4, h_s_dadda_rca32_fa383_y2, h_s_dadda_rca32_fa383_y4);
  fa fa_h_s_dadda_rca32_fa384_y2(h_s_dadda_rca32_fa363_y4, h_s_dadda_rca32_fa362_y4, h_s_dadda_rca32_fa361_y4, h_s_dadda_rca32_fa384_y2, h_s_dadda_rca32_fa384_y4);
  fa fa_h_s_dadda_rca32_fa385_y2(h_s_dadda_rca32_fa360_y4, h_s_dadda_rca32_fa359_y4, h_s_dadda_rca32_fa358_y4, h_s_dadda_rca32_fa385_y2, h_s_dadda_rca32_fa385_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_6_y0(a_28, b_6, h_s_dadda_rca32_and_28_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_7_y0(a_27, b_7, h_s_dadda_rca32_and_27_7_y0);
  fa fa_h_s_dadda_rca32_fa386_y2(h_s_dadda_rca32_fa357_y4, h_s_dadda_rca32_and_28_6_y0, h_s_dadda_rca32_and_27_7_y0, h_s_dadda_rca32_fa386_y2, h_s_dadda_rca32_fa386_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_8_y0(a_26, b_8, h_s_dadda_rca32_and_26_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_9_y0(a_25, b_9, h_s_dadda_rca32_and_25_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_10_y0(a_24, b_10, h_s_dadda_rca32_and_24_10_y0);
  fa fa_h_s_dadda_rca32_fa387_y2(h_s_dadda_rca32_and_26_8_y0, h_s_dadda_rca32_and_25_9_y0, h_s_dadda_rca32_and_24_10_y0, h_s_dadda_rca32_fa387_y2, h_s_dadda_rca32_fa387_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_11_y0(a_23, b_11, h_s_dadda_rca32_and_23_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_12_y0(a_22, b_12, h_s_dadda_rca32_and_22_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_13_y0(a_21, b_13, h_s_dadda_rca32_and_21_13_y0);
  fa fa_h_s_dadda_rca32_fa388_y2(h_s_dadda_rca32_and_23_11_y0, h_s_dadda_rca32_and_22_12_y0, h_s_dadda_rca32_and_21_13_y0, h_s_dadda_rca32_fa388_y2, h_s_dadda_rca32_fa388_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_14_y0(a_20, b_14, h_s_dadda_rca32_and_20_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_15_y0(a_19, b_15, h_s_dadda_rca32_and_19_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_16_y0(a_18, b_16, h_s_dadda_rca32_and_18_16_y0);
  fa fa_h_s_dadda_rca32_fa389_y2(h_s_dadda_rca32_and_20_14_y0, h_s_dadda_rca32_and_19_15_y0, h_s_dadda_rca32_and_18_16_y0, h_s_dadda_rca32_fa389_y2, h_s_dadda_rca32_fa389_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_17_y0(a_17, b_17, h_s_dadda_rca32_and_17_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_18_y0(a_16, b_18, h_s_dadda_rca32_and_16_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_19_y0(a_15, b_19, h_s_dadda_rca32_and_15_19_y0);
  fa fa_h_s_dadda_rca32_fa390_y2(h_s_dadda_rca32_and_17_17_y0, h_s_dadda_rca32_and_16_18_y0, h_s_dadda_rca32_and_15_19_y0, h_s_dadda_rca32_fa390_y2, h_s_dadda_rca32_fa390_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_20_y0(a_14, b_20, h_s_dadda_rca32_and_14_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_21_y0(a_13, b_21, h_s_dadda_rca32_and_13_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_22_y0(a_12, b_22, h_s_dadda_rca32_and_12_22_y0);
  fa fa_h_s_dadda_rca32_fa391_y2(h_s_dadda_rca32_and_14_20_y0, h_s_dadda_rca32_and_13_21_y0, h_s_dadda_rca32_and_12_22_y0, h_s_dadda_rca32_fa391_y2, h_s_dadda_rca32_fa391_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_23_y0(a_11, b_23, h_s_dadda_rca32_and_11_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_24_y0(a_10, b_24, h_s_dadda_rca32_and_10_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_25_y0(a_9, b_25, h_s_dadda_rca32_and_9_25_y0);
  fa fa_h_s_dadda_rca32_fa392_y2(h_s_dadda_rca32_and_11_23_y0, h_s_dadda_rca32_and_10_24_y0, h_s_dadda_rca32_and_9_25_y0, h_s_dadda_rca32_fa392_y2, h_s_dadda_rca32_fa392_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_26_y0(a_8, b_26, h_s_dadda_rca32_and_8_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_27_y0(a_7, b_27, h_s_dadda_rca32_and_7_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_28_y0(a_6, b_28, h_s_dadda_rca32_and_6_28_y0);
  fa fa_h_s_dadda_rca32_fa393_y2(h_s_dadda_rca32_and_8_26_y0, h_s_dadda_rca32_and_7_27_y0, h_s_dadda_rca32_and_6_28_y0, h_s_dadda_rca32_fa393_y2, h_s_dadda_rca32_fa393_y4);
  and_gate and_gate_h_s_dadda_rca32_and_5_29_y0(a_5, b_29, h_s_dadda_rca32_and_5_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_30_y0(a_4, b_30, h_s_dadda_rca32_and_4_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_3_31_y0(a_3, b_31, h_s_dadda_rca32_nand_3_31_y0);
  fa fa_h_s_dadda_rca32_fa394_y2(h_s_dadda_rca32_and_5_29_y0, h_s_dadda_rca32_and_4_30_y0, h_s_dadda_rca32_nand_3_31_y0, h_s_dadda_rca32_fa394_y2, h_s_dadda_rca32_fa394_y4);
  fa fa_h_s_dadda_rca32_fa395_y2(h_s_dadda_rca32_fa13_y2, h_s_dadda_rca32_fa14_y2, h_s_dadda_rca32_fa379_y2, h_s_dadda_rca32_fa395_y2, h_s_dadda_rca32_fa395_y4);
  fa fa_h_s_dadda_rca32_fa396_y2(h_s_dadda_rca32_fa380_y2, h_s_dadda_rca32_fa381_y2, h_s_dadda_rca32_fa382_y2, h_s_dadda_rca32_fa396_y2, h_s_dadda_rca32_fa396_y4);
  fa fa_h_s_dadda_rca32_fa397_y2(h_s_dadda_rca32_fa383_y2, h_s_dadda_rca32_fa384_y2, h_s_dadda_rca32_fa385_y2, h_s_dadda_rca32_fa397_y2, h_s_dadda_rca32_fa397_y4);
  fa fa_h_s_dadda_rca32_fa398_y2(h_s_dadda_rca32_fa386_y2, h_s_dadda_rca32_fa387_y2, h_s_dadda_rca32_fa388_y2, h_s_dadda_rca32_fa398_y2, h_s_dadda_rca32_fa398_y4);
  fa fa_h_s_dadda_rca32_fa399_y2(h_s_dadda_rca32_fa389_y2, h_s_dadda_rca32_fa390_y2, h_s_dadda_rca32_fa391_y2, h_s_dadda_rca32_fa399_y2, h_s_dadda_rca32_fa399_y4);
  fa fa_h_s_dadda_rca32_fa400_y2(h_s_dadda_rca32_fa392_y2, h_s_dadda_rca32_fa393_y2, h_s_dadda_rca32_fa394_y2, h_s_dadda_rca32_fa400_y2, h_s_dadda_rca32_fa400_y4);
  fa fa_h_s_dadda_rca32_fa401_y2(h_s_dadda_rca32_fa400_y4, h_s_dadda_rca32_fa399_y4, h_s_dadda_rca32_fa398_y4, h_s_dadda_rca32_fa401_y2, h_s_dadda_rca32_fa401_y4);
  fa fa_h_s_dadda_rca32_fa402_y2(h_s_dadda_rca32_fa397_y4, h_s_dadda_rca32_fa396_y4, h_s_dadda_rca32_fa395_y4, h_s_dadda_rca32_fa402_y2, h_s_dadda_rca32_fa402_y4);
  fa fa_h_s_dadda_rca32_fa403_y2(h_s_dadda_rca32_fa394_y4, h_s_dadda_rca32_fa393_y4, h_s_dadda_rca32_fa392_y4, h_s_dadda_rca32_fa403_y2, h_s_dadda_rca32_fa403_y4);
  fa fa_h_s_dadda_rca32_fa404_y2(h_s_dadda_rca32_fa391_y4, h_s_dadda_rca32_fa390_y4, h_s_dadda_rca32_fa389_y4, h_s_dadda_rca32_fa404_y2, h_s_dadda_rca32_fa404_y4);
  fa fa_h_s_dadda_rca32_fa405_y2(h_s_dadda_rca32_fa388_y4, h_s_dadda_rca32_fa387_y4, h_s_dadda_rca32_fa386_y4, h_s_dadda_rca32_fa405_y2, h_s_dadda_rca32_fa405_y4);
  fa fa_h_s_dadda_rca32_fa406_y2(h_s_dadda_rca32_fa385_y4, h_s_dadda_rca32_fa384_y4, h_s_dadda_rca32_fa383_y4, h_s_dadda_rca32_fa406_y2, h_s_dadda_rca32_fa406_y4);
  fa fa_h_s_dadda_rca32_fa407_y2(h_s_dadda_rca32_fa382_y4, h_s_dadda_rca32_fa381_y4, h_s_dadda_rca32_fa380_y4, h_s_dadda_rca32_fa407_y2, h_s_dadda_rca32_fa407_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_5_y0(a_30, b_5, h_s_dadda_rca32_and_30_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_6_y0(a_29, b_6, h_s_dadda_rca32_and_29_6_y0);
  fa fa_h_s_dadda_rca32_fa408_y2(h_s_dadda_rca32_fa379_y4, h_s_dadda_rca32_and_30_5_y0, h_s_dadda_rca32_and_29_6_y0, h_s_dadda_rca32_fa408_y2, h_s_dadda_rca32_fa408_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_7_y0(a_28, b_7, h_s_dadda_rca32_and_28_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_8_y0(a_27, b_8, h_s_dadda_rca32_and_27_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_9_y0(a_26, b_9, h_s_dadda_rca32_and_26_9_y0);
  fa fa_h_s_dadda_rca32_fa409_y2(h_s_dadda_rca32_and_28_7_y0, h_s_dadda_rca32_and_27_8_y0, h_s_dadda_rca32_and_26_9_y0, h_s_dadda_rca32_fa409_y2, h_s_dadda_rca32_fa409_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_10_y0(a_25, b_10, h_s_dadda_rca32_and_25_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_11_y0(a_24, b_11, h_s_dadda_rca32_and_24_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_12_y0(a_23, b_12, h_s_dadda_rca32_and_23_12_y0);
  fa fa_h_s_dadda_rca32_fa410_y2(h_s_dadda_rca32_and_25_10_y0, h_s_dadda_rca32_and_24_11_y0, h_s_dadda_rca32_and_23_12_y0, h_s_dadda_rca32_fa410_y2, h_s_dadda_rca32_fa410_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_13_y0(a_22, b_13, h_s_dadda_rca32_and_22_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_14_y0(a_21, b_14, h_s_dadda_rca32_and_21_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_15_y0(a_20, b_15, h_s_dadda_rca32_and_20_15_y0);
  fa fa_h_s_dadda_rca32_fa411_y2(h_s_dadda_rca32_and_22_13_y0, h_s_dadda_rca32_and_21_14_y0, h_s_dadda_rca32_and_20_15_y0, h_s_dadda_rca32_fa411_y2, h_s_dadda_rca32_fa411_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_16_y0(a_19, b_16, h_s_dadda_rca32_and_19_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_17_y0(a_18, b_17, h_s_dadda_rca32_and_18_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_18_y0(a_17, b_18, h_s_dadda_rca32_and_17_18_y0);
  fa fa_h_s_dadda_rca32_fa412_y2(h_s_dadda_rca32_and_19_16_y0, h_s_dadda_rca32_and_18_17_y0, h_s_dadda_rca32_and_17_18_y0, h_s_dadda_rca32_fa412_y2, h_s_dadda_rca32_fa412_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_19_y0(a_16, b_19, h_s_dadda_rca32_and_16_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_20_y0(a_15, b_20, h_s_dadda_rca32_and_15_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_21_y0(a_14, b_21, h_s_dadda_rca32_and_14_21_y0);
  fa fa_h_s_dadda_rca32_fa413_y2(h_s_dadda_rca32_and_16_19_y0, h_s_dadda_rca32_and_15_20_y0, h_s_dadda_rca32_and_14_21_y0, h_s_dadda_rca32_fa413_y2, h_s_dadda_rca32_fa413_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_22_y0(a_13, b_22, h_s_dadda_rca32_and_13_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_23_y0(a_12, b_23, h_s_dadda_rca32_and_12_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_24_y0(a_11, b_24, h_s_dadda_rca32_and_11_24_y0);
  fa fa_h_s_dadda_rca32_fa414_y2(h_s_dadda_rca32_and_13_22_y0, h_s_dadda_rca32_and_12_23_y0, h_s_dadda_rca32_and_11_24_y0, h_s_dadda_rca32_fa414_y2, h_s_dadda_rca32_fa414_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_25_y0(a_10, b_25, h_s_dadda_rca32_and_10_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_26_y0(a_9, b_26, h_s_dadda_rca32_and_9_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_27_y0(a_8, b_27, h_s_dadda_rca32_and_8_27_y0);
  fa fa_h_s_dadda_rca32_fa415_y2(h_s_dadda_rca32_and_10_25_y0, h_s_dadda_rca32_and_9_26_y0, h_s_dadda_rca32_and_8_27_y0, h_s_dadda_rca32_fa415_y2, h_s_dadda_rca32_fa415_y4);
  and_gate and_gate_h_s_dadda_rca32_and_7_28_y0(a_7, b_28, h_s_dadda_rca32_and_7_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_6_29_y0(a_6, b_29, h_s_dadda_rca32_and_6_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_5_30_y0(a_5, b_30, h_s_dadda_rca32_and_5_30_y0);
  fa fa_h_s_dadda_rca32_fa416_y2(h_s_dadda_rca32_and_7_28_y0, h_s_dadda_rca32_and_6_29_y0, h_s_dadda_rca32_and_5_30_y0, h_s_dadda_rca32_fa416_y2, h_s_dadda_rca32_fa416_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_4_31_y0(a_4, b_31, h_s_dadda_rca32_nand_4_31_y0);
  fa fa_h_s_dadda_rca32_fa417_y2(h_s_dadda_rca32_nand_4_31_y0, h_s_dadda_rca32_fa15_y2, h_s_dadda_rca32_fa401_y2, h_s_dadda_rca32_fa417_y2, h_s_dadda_rca32_fa417_y4);
  fa fa_h_s_dadda_rca32_fa418_y2(h_s_dadda_rca32_fa402_y2, h_s_dadda_rca32_fa403_y2, h_s_dadda_rca32_fa404_y2, h_s_dadda_rca32_fa418_y2, h_s_dadda_rca32_fa418_y4);
  fa fa_h_s_dadda_rca32_fa419_y2(h_s_dadda_rca32_fa405_y2, h_s_dadda_rca32_fa406_y2, h_s_dadda_rca32_fa407_y2, h_s_dadda_rca32_fa419_y2, h_s_dadda_rca32_fa419_y4);
  fa fa_h_s_dadda_rca32_fa420_y2(h_s_dadda_rca32_fa408_y2, h_s_dadda_rca32_fa409_y2, h_s_dadda_rca32_fa410_y2, h_s_dadda_rca32_fa420_y2, h_s_dadda_rca32_fa420_y4);
  fa fa_h_s_dadda_rca32_fa421_y2(h_s_dadda_rca32_fa411_y2, h_s_dadda_rca32_fa412_y2, h_s_dadda_rca32_fa413_y2, h_s_dadda_rca32_fa421_y2, h_s_dadda_rca32_fa421_y4);
  fa fa_h_s_dadda_rca32_fa422_y2(h_s_dadda_rca32_fa414_y2, h_s_dadda_rca32_fa415_y2, h_s_dadda_rca32_fa416_y2, h_s_dadda_rca32_fa422_y2, h_s_dadda_rca32_fa422_y4);
  fa fa_h_s_dadda_rca32_fa423_y2(h_s_dadda_rca32_fa422_y4, h_s_dadda_rca32_fa421_y4, h_s_dadda_rca32_fa420_y4, h_s_dadda_rca32_fa423_y2, h_s_dadda_rca32_fa423_y4);
  fa fa_h_s_dadda_rca32_fa424_y2(h_s_dadda_rca32_fa419_y4, h_s_dadda_rca32_fa418_y4, h_s_dadda_rca32_fa417_y4, h_s_dadda_rca32_fa424_y2, h_s_dadda_rca32_fa424_y4);
  fa fa_h_s_dadda_rca32_fa425_y2(h_s_dadda_rca32_fa416_y4, h_s_dadda_rca32_fa415_y4, h_s_dadda_rca32_fa414_y4, h_s_dadda_rca32_fa425_y2, h_s_dadda_rca32_fa425_y4);
  fa fa_h_s_dadda_rca32_fa426_y2(h_s_dadda_rca32_fa413_y4, h_s_dadda_rca32_fa412_y4, h_s_dadda_rca32_fa411_y4, h_s_dadda_rca32_fa426_y2, h_s_dadda_rca32_fa426_y4);
  fa fa_h_s_dadda_rca32_fa427_y2(h_s_dadda_rca32_fa410_y4, h_s_dadda_rca32_fa409_y4, h_s_dadda_rca32_fa408_y4, h_s_dadda_rca32_fa427_y2, h_s_dadda_rca32_fa427_y4);
  fa fa_h_s_dadda_rca32_fa428_y2(h_s_dadda_rca32_fa407_y4, h_s_dadda_rca32_fa406_y4, h_s_dadda_rca32_fa405_y4, h_s_dadda_rca32_fa428_y2, h_s_dadda_rca32_fa428_y4);
  fa fa_h_s_dadda_rca32_fa429_y2(h_s_dadda_rca32_fa404_y4, h_s_dadda_rca32_fa403_y4, h_s_dadda_rca32_fa402_y4, h_s_dadda_rca32_fa429_y2, h_s_dadda_rca32_fa429_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_5_y0(a_31, b_5, h_s_dadda_rca32_nand_31_5_y0);
  fa fa_h_s_dadda_rca32_fa430_y2(h_s_dadda_rca32_fa401_y4, h_s_dadda_rca32_fa15_y4, h_s_dadda_rca32_nand_31_5_y0, h_s_dadda_rca32_fa430_y2, h_s_dadda_rca32_fa430_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_6_y0(a_30, b_6, h_s_dadda_rca32_and_30_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_7_y0(a_29, b_7, h_s_dadda_rca32_and_29_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_8_y0(a_28, b_8, h_s_dadda_rca32_and_28_8_y0);
  fa fa_h_s_dadda_rca32_fa431_y2(h_s_dadda_rca32_and_30_6_y0, h_s_dadda_rca32_and_29_7_y0, h_s_dadda_rca32_and_28_8_y0, h_s_dadda_rca32_fa431_y2, h_s_dadda_rca32_fa431_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_9_y0(a_27, b_9, h_s_dadda_rca32_and_27_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_10_y0(a_26, b_10, h_s_dadda_rca32_and_26_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_11_y0(a_25, b_11, h_s_dadda_rca32_and_25_11_y0);
  fa fa_h_s_dadda_rca32_fa432_y2(h_s_dadda_rca32_and_27_9_y0, h_s_dadda_rca32_and_26_10_y0, h_s_dadda_rca32_and_25_11_y0, h_s_dadda_rca32_fa432_y2, h_s_dadda_rca32_fa432_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_12_y0(a_24, b_12, h_s_dadda_rca32_and_24_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_13_y0(a_23, b_13, h_s_dadda_rca32_and_23_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_14_y0(a_22, b_14, h_s_dadda_rca32_and_22_14_y0);
  fa fa_h_s_dadda_rca32_fa433_y2(h_s_dadda_rca32_and_24_12_y0, h_s_dadda_rca32_and_23_13_y0, h_s_dadda_rca32_and_22_14_y0, h_s_dadda_rca32_fa433_y2, h_s_dadda_rca32_fa433_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_15_y0(a_21, b_15, h_s_dadda_rca32_and_21_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_16_y0(a_20, b_16, h_s_dadda_rca32_and_20_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_17_y0(a_19, b_17, h_s_dadda_rca32_and_19_17_y0);
  fa fa_h_s_dadda_rca32_fa434_y2(h_s_dadda_rca32_and_21_15_y0, h_s_dadda_rca32_and_20_16_y0, h_s_dadda_rca32_and_19_17_y0, h_s_dadda_rca32_fa434_y2, h_s_dadda_rca32_fa434_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_18_y0(a_18, b_18, h_s_dadda_rca32_and_18_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_19_y0(a_17, b_19, h_s_dadda_rca32_and_17_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_20_y0(a_16, b_20, h_s_dadda_rca32_and_16_20_y0);
  fa fa_h_s_dadda_rca32_fa435_y2(h_s_dadda_rca32_and_18_18_y0, h_s_dadda_rca32_and_17_19_y0, h_s_dadda_rca32_and_16_20_y0, h_s_dadda_rca32_fa435_y2, h_s_dadda_rca32_fa435_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_21_y0(a_15, b_21, h_s_dadda_rca32_and_15_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_22_y0(a_14, b_22, h_s_dadda_rca32_and_14_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_23_y0(a_13, b_23, h_s_dadda_rca32_and_13_23_y0);
  fa fa_h_s_dadda_rca32_fa436_y2(h_s_dadda_rca32_and_15_21_y0, h_s_dadda_rca32_and_14_22_y0, h_s_dadda_rca32_and_13_23_y0, h_s_dadda_rca32_fa436_y2, h_s_dadda_rca32_fa436_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_24_y0(a_12, b_24, h_s_dadda_rca32_and_12_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_25_y0(a_11, b_25, h_s_dadda_rca32_and_11_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_26_y0(a_10, b_26, h_s_dadda_rca32_and_10_26_y0);
  fa fa_h_s_dadda_rca32_fa437_y2(h_s_dadda_rca32_and_12_24_y0, h_s_dadda_rca32_and_11_25_y0, h_s_dadda_rca32_and_10_26_y0, h_s_dadda_rca32_fa437_y2, h_s_dadda_rca32_fa437_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_27_y0(a_9, b_27, h_s_dadda_rca32_and_9_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_28_y0(a_8, b_28, h_s_dadda_rca32_and_8_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_29_y0(a_7, b_29, h_s_dadda_rca32_and_7_29_y0);
  fa fa_h_s_dadda_rca32_fa438_y2(h_s_dadda_rca32_and_9_27_y0, h_s_dadda_rca32_and_8_28_y0, h_s_dadda_rca32_and_7_29_y0, h_s_dadda_rca32_fa438_y2, h_s_dadda_rca32_fa438_y4);
  and_gate and_gate_h_s_dadda_rca32_and_6_30_y0(a_6, b_30, h_s_dadda_rca32_and_6_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_5_31_y0(a_5, b_31, h_s_dadda_rca32_nand_5_31_y0);
  fa fa_h_s_dadda_rca32_fa439_y2(h_s_dadda_rca32_and_6_30_y0, h_s_dadda_rca32_nand_5_31_y0, h_s_dadda_rca32_fa423_y2, h_s_dadda_rca32_fa439_y2, h_s_dadda_rca32_fa439_y4);
  fa fa_h_s_dadda_rca32_fa440_y2(h_s_dadda_rca32_fa424_y2, h_s_dadda_rca32_fa425_y2, h_s_dadda_rca32_fa426_y2, h_s_dadda_rca32_fa440_y2, h_s_dadda_rca32_fa440_y4);
  fa fa_h_s_dadda_rca32_fa441_y2(h_s_dadda_rca32_fa427_y2, h_s_dadda_rca32_fa428_y2, h_s_dadda_rca32_fa429_y2, h_s_dadda_rca32_fa441_y2, h_s_dadda_rca32_fa441_y4);
  fa fa_h_s_dadda_rca32_fa442_y2(h_s_dadda_rca32_fa430_y2, h_s_dadda_rca32_fa431_y2, h_s_dadda_rca32_fa432_y2, h_s_dadda_rca32_fa442_y2, h_s_dadda_rca32_fa442_y4);
  fa fa_h_s_dadda_rca32_fa443_y2(h_s_dadda_rca32_fa433_y2, h_s_dadda_rca32_fa434_y2, h_s_dadda_rca32_fa435_y2, h_s_dadda_rca32_fa443_y2, h_s_dadda_rca32_fa443_y4);
  fa fa_h_s_dadda_rca32_fa444_y2(h_s_dadda_rca32_fa436_y2, h_s_dadda_rca32_fa437_y2, h_s_dadda_rca32_fa438_y2, h_s_dadda_rca32_fa444_y2, h_s_dadda_rca32_fa444_y4);
  fa fa_h_s_dadda_rca32_fa445_y2(h_s_dadda_rca32_fa444_y4, h_s_dadda_rca32_fa443_y4, h_s_dadda_rca32_fa442_y4, h_s_dadda_rca32_fa445_y2, h_s_dadda_rca32_fa445_y4);
  fa fa_h_s_dadda_rca32_fa446_y2(h_s_dadda_rca32_fa441_y4, h_s_dadda_rca32_fa440_y4, h_s_dadda_rca32_fa439_y4, h_s_dadda_rca32_fa446_y2, h_s_dadda_rca32_fa446_y4);
  fa fa_h_s_dadda_rca32_fa447_y2(h_s_dadda_rca32_fa438_y4, h_s_dadda_rca32_fa437_y4, h_s_dadda_rca32_fa436_y4, h_s_dadda_rca32_fa447_y2, h_s_dadda_rca32_fa447_y4);
  fa fa_h_s_dadda_rca32_fa448_y2(h_s_dadda_rca32_fa435_y4, h_s_dadda_rca32_fa434_y4, h_s_dadda_rca32_fa433_y4, h_s_dadda_rca32_fa448_y2, h_s_dadda_rca32_fa448_y4);
  fa fa_h_s_dadda_rca32_fa449_y2(h_s_dadda_rca32_fa432_y4, h_s_dadda_rca32_fa431_y4, h_s_dadda_rca32_fa430_y4, h_s_dadda_rca32_fa449_y2, h_s_dadda_rca32_fa449_y4);
  fa fa_h_s_dadda_rca32_fa450_y2(h_s_dadda_rca32_fa429_y4, h_s_dadda_rca32_fa428_y4, h_s_dadda_rca32_fa427_y4, h_s_dadda_rca32_fa450_y2, h_s_dadda_rca32_fa450_y4);
  fa fa_h_s_dadda_rca32_fa451_y2(h_s_dadda_rca32_fa426_y4, h_s_dadda_rca32_fa425_y4, h_s_dadda_rca32_fa424_y4, h_s_dadda_rca32_fa451_y2, h_s_dadda_rca32_fa451_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_6_y0(a_31, b_6, h_s_dadda_rca32_nand_31_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_7_y0(a_30, b_7, h_s_dadda_rca32_and_30_7_y0);
  fa fa_h_s_dadda_rca32_fa452_y2(h_s_dadda_rca32_fa423_y4, h_s_dadda_rca32_nand_31_6_y0, h_s_dadda_rca32_and_30_7_y0, h_s_dadda_rca32_fa452_y2, h_s_dadda_rca32_fa452_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_8_y0(a_29, b_8, h_s_dadda_rca32_and_29_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_9_y0(a_28, b_9, h_s_dadda_rca32_and_28_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_10_y0(a_27, b_10, h_s_dadda_rca32_and_27_10_y0);
  fa fa_h_s_dadda_rca32_fa453_y2(h_s_dadda_rca32_and_29_8_y0, h_s_dadda_rca32_and_28_9_y0, h_s_dadda_rca32_and_27_10_y0, h_s_dadda_rca32_fa453_y2, h_s_dadda_rca32_fa453_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_11_y0(a_26, b_11, h_s_dadda_rca32_and_26_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_12_y0(a_25, b_12, h_s_dadda_rca32_and_25_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_13_y0(a_24, b_13, h_s_dadda_rca32_and_24_13_y0);
  fa fa_h_s_dadda_rca32_fa454_y2(h_s_dadda_rca32_and_26_11_y0, h_s_dadda_rca32_and_25_12_y0, h_s_dadda_rca32_and_24_13_y0, h_s_dadda_rca32_fa454_y2, h_s_dadda_rca32_fa454_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_14_y0(a_23, b_14, h_s_dadda_rca32_and_23_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_15_y0(a_22, b_15, h_s_dadda_rca32_and_22_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_16_y0(a_21, b_16, h_s_dadda_rca32_and_21_16_y0);
  fa fa_h_s_dadda_rca32_fa455_y2(h_s_dadda_rca32_and_23_14_y0, h_s_dadda_rca32_and_22_15_y0, h_s_dadda_rca32_and_21_16_y0, h_s_dadda_rca32_fa455_y2, h_s_dadda_rca32_fa455_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_17_y0(a_20, b_17, h_s_dadda_rca32_and_20_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_18_y0(a_19, b_18, h_s_dadda_rca32_and_19_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_19_y0(a_18, b_19, h_s_dadda_rca32_and_18_19_y0);
  fa fa_h_s_dadda_rca32_fa456_y2(h_s_dadda_rca32_and_20_17_y0, h_s_dadda_rca32_and_19_18_y0, h_s_dadda_rca32_and_18_19_y0, h_s_dadda_rca32_fa456_y2, h_s_dadda_rca32_fa456_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_20_y0(a_17, b_20, h_s_dadda_rca32_and_17_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_21_y0(a_16, b_21, h_s_dadda_rca32_and_16_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_22_y0(a_15, b_22, h_s_dadda_rca32_and_15_22_y0);
  fa fa_h_s_dadda_rca32_fa457_y2(h_s_dadda_rca32_and_17_20_y0, h_s_dadda_rca32_and_16_21_y0, h_s_dadda_rca32_and_15_22_y0, h_s_dadda_rca32_fa457_y2, h_s_dadda_rca32_fa457_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_23_y0(a_14, b_23, h_s_dadda_rca32_and_14_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_24_y0(a_13, b_24, h_s_dadda_rca32_and_13_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_25_y0(a_12, b_25, h_s_dadda_rca32_and_12_25_y0);
  fa fa_h_s_dadda_rca32_fa458_y2(h_s_dadda_rca32_and_14_23_y0, h_s_dadda_rca32_and_13_24_y0, h_s_dadda_rca32_and_12_25_y0, h_s_dadda_rca32_fa458_y2, h_s_dadda_rca32_fa458_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_26_y0(a_11, b_26, h_s_dadda_rca32_and_11_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_27_y0(a_10, b_27, h_s_dadda_rca32_and_10_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_28_y0(a_9, b_28, h_s_dadda_rca32_and_9_28_y0);
  fa fa_h_s_dadda_rca32_fa459_y2(h_s_dadda_rca32_and_11_26_y0, h_s_dadda_rca32_and_10_27_y0, h_s_dadda_rca32_and_9_28_y0, h_s_dadda_rca32_fa459_y2, h_s_dadda_rca32_fa459_y4);
  and_gate and_gate_h_s_dadda_rca32_and_8_29_y0(a_8, b_29, h_s_dadda_rca32_and_8_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_7_30_y0(a_7, b_30, h_s_dadda_rca32_and_7_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_6_31_y0(a_6, b_31, h_s_dadda_rca32_nand_6_31_y0);
  fa fa_h_s_dadda_rca32_fa460_y2(h_s_dadda_rca32_and_8_29_y0, h_s_dadda_rca32_and_7_30_y0, h_s_dadda_rca32_nand_6_31_y0, h_s_dadda_rca32_fa460_y2, h_s_dadda_rca32_fa460_y4);
  fa fa_h_s_dadda_rca32_fa461_y2(h_s_dadda_rca32_fa445_y2, h_s_dadda_rca32_fa446_y2, h_s_dadda_rca32_fa447_y2, h_s_dadda_rca32_fa461_y2, h_s_dadda_rca32_fa461_y4);
  fa fa_h_s_dadda_rca32_fa462_y2(h_s_dadda_rca32_fa448_y2, h_s_dadda_rca32_fa449_y2, h_s_dadda_rca32_fa450_y2, h_s_dadda_rca32_fa462_y2, h_s_dadda_rca32_fa462_y4);
  fa fa_h_s_dadda_rca32_fa463_y2(h_s_dadda_rca32_fa451_y2, h_s_dadda_rca32_fa452_y2, h_s_dadda_rca32_fa453_y2, h_s_dadda_rca32_fa463_y2, h_s_dadda_rca32_fa463_y4);
  fa fa_h_s_dadda_rca32_fa464_y2(h_s_dadda_rca32_fa454_y2, h_s_dadda_rca32_fa455_y2, h_s_dadda_rca32_fa456_y2, h_s_dadda_rca32_fa464_y2, h_s_dadda_rca32_fa464_y4);
  fa fa_h_s_dadda_rca32_fa465_y2(h_s_dadda_rca32_fa457_y2, h_s_dadda_rca32_fa458_y2, h_s_dadda_rca32_fa459_y2, h_s_dadda_rca32_fa465_y2, h_s_dadda_rca32_fa465_y4);
  fa fa_h_s_dadda_rca32_fa466_y2(h_s_dadda_rca32_fa465_y4, h_s_dadda_rca32_fa464_y4, h_s_dadda_rca32_fa463_y4, h_s_dadda_rca32_fa466_y2, h_s_dadda_rca32_fa466_y4);
  fa fa_h_s_dadda_rca32_fa467_y2(h_s_dadda_rca32_fa462_y4, h_s_dadda_rca32_fa461_y4, h_s_dadda_rca32_fa460_y4, h_s_dadda_rca32_fa467_y2, h_s_dadda_rca32_fa467_y4);
  fa fa_h_s_dadda_rca32_fa468_y2(h_s_dadda_rca32_fa459_y4, h_s_dadda_rca32_fa458_y4, h_s_dadda_rca32_fa457_y4, h_s_dadda_rca32_fa468_y2, h_s_dadda_rca32_fa468_y4);
  fa fa_h_s_dadda_rca32_fa469_y2(h_s_dadda_rca32_fa456_y4, h_s_dadda_rca32_fa455_y4, h_s_dadda_rca32_fa454_y4, h_s_dadda_rca32_fa469_y2, h_s_dadda_rca32_fa469_y4);
  fa fa_h_s_dadda_rca32_fa470_y2(h_s_dadda_rca32_fa453_y4, h_s_dadda_rca32_fa452_y4, h_s_dadda_rca32_fa451_y4, h_s_dadda_rca32_fa470_y2, h_s_dadda_rca32_fa470_y4);
  fa fa_h_s_dadda_rca32_fa471_y2(h_s_dadda_rca32_fa450_y4, h_s_dadda_rca32_fa449_y4, h_s_dadda_rca32_fa448_y4, h_s_dadda_rca32_fa471_y2, h_s_dadda_rca32_fa471_y4);
  fa fa_h_s_dadda_rca32_fa472_y2(h_s_dadda_rca32_fa447_y4, h_s_dadda_rca32_fa446_y4, h_s_dadda_rca32_fa445_y4, h_s_dadda_rca32_fa472_y2, h_s_dadda_rca32_fa472_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_7_y0(a_31, b_7, h_s_dadda_rca32_nand_31_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_8_y0(a_30, b_8, h_s_dadda_rca32_and_30_8_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_9_y0(a_29, b_9, h_s_dadda_rca32_and_29_9_y0);
  fa fa_h_s_dadda_rca32_fa473_y2(h_s_dadda_rca32_nand_31_7_y0, h_s_dadda_rca32_and_30_8_y0, h_s_dadda_rca32_and_29_9_y0, h_s_dadda_rca32_fa473_y2, h_s_dadda_rca32_fa473_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_10_y0(a_28, b_10, h_s_dadda_rca32_and_28_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_11_y0(a_27, b_11, h_s_dadda_rca32_and_27_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_12_y0(a_26, b_12, h_s_dadda_rca32_and_26_12_y0);
  fa fa_h_s_dadda_rca32_fa474_y2(h_s_dadda_rca32_and_28_10_y0, h_s_dadda_rca32_and_27_11_y0, h_s_dadda_rca32_and_26_12_y0, h_s_dadda_rca32_fa474_y2, h_s_dadda_rca32_fa474_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_13_y0(a_25, b_13, h_s_dadda_rca32_and_25_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_14_y0(a_24, b_14, h_s_dadda_rca32_and_24_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_15_y0(a_23, b_15, h_s_dadda_rca32_and_23_15_y0);
  fa fa_h_s_dadda_rca32_fa475_y2(h_s_dadda_rca32_and_25_13_y0, h_s_dadda_rca32_and_24_14_y0, h_s_dadda_rca32_and_23_15_y0, h_s_dadda_rca32_fa475_y2, h_s_dadda_rca32_fa475_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_16_y0(a_22, b_16, h_s_dadda_rca32_and_22_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_17_y0(a_21, b_17, h_s_dadda_rca32_and_21_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_18_y0(a_20, b_18, h_s_dadda_rca32_and_20_18_y0);
  fa fa_h_s_dadda_rca32_fa476_y2(h_s_dadda_rca32_and_22_16_y0, h_s_dadda_rca32_and_21_17_y0, h_s_dadda_rca32_and_20_18_y0, h_s_dadda_rca32_fa476_y2, h_s_dadda_rca32_fa476_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_19_y0(a_19, b_19, h_s_dadda_rca32_and_19_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_20_y0(a_18, b_20, h_s_dadda_rca32_and_18_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_21_y0(a_17, b_21, h_s_dadda_rca32_and_17_21_y0);
  fa fa_h_s_dadda_rca32_fa477_y2(h_s_dadda_rca32_and_19_19_y0, h_s_dadda_rca32_and_18_20_y0, h_s_dadda_rca32_and_17_21_y0, h_s_dadda_rca32_fa477_y2, h_s_dadda_rca32_fa477_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_22_y0(a_16, b_22, h_s_dadda_rca32_and_16_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_23_y0(a_15, b_23, h_s_dadda_rca32_and_15_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_24_y0(a_14, b_24, h_s_dadda_rca32_and_14_24_y0);
  fa fa_h_s_dadda_rca32_fa478_y2(h_s_dadda_rca32_and_16_22_y0, h_s_dadda_rca32_and_15_23_y0, h_s_dadda_rca32_and_14_24_y0, h_s_dadda_rca32_fa478_y2, h_s_dadda_rca32_fa478_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_25_y0(a_13, b_25, h_s_dadda_rca32_and_13_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_26_y0(a_12, b_26, h_s_dadda_rca32_and_12_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_27_y0(a_11, b_27, h_s_dadda_rca32_and_11_27_y0);
  fa fa_h_s_dadda_rca32_fa479_y2(h_s_dadda_rca32_and_13_25_y0, h_s_dadda_rca32_and_12_26_y0, h_s_dadda_rca32_and_11_27_y0, h_s_dadda_rca32_fa479_y2, h_s_dadda_rca32_fa479_y4);
  and_gate and_gate_h_s_dadda_rca32_and_10_28_y0(a_10, b_28, h_s_dadda_rca32_and_10_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_9_29_y0(a_9, b_29, h_s_dadda_rca32_and_9_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_8_30_y0(a_8, b_30, h_s_dadda_rca32_and_8_30_y0);
  fa fa_h_s_dadda_rca32_fa480_y2(h_s_dadda_rca32_and_10_28_y0, h_s_dadda_rca32_and_9_29_y0, h_s_dadda_rca32_and_8_30_y0, h_s_dadda_rca32_fa480_y2, h_s_dadda_rca32_fa480_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_7_31_y0(a_7, b_31, h_s_dadda_rca32_nand_7_31_y0);
  fa fa_h_s_dadda_rca32_fa481_y2(h_s_dadda_rca32_nand_7_31_y0, h_s_dadda_rca32_fa466_y2, h_s_dadda_rca32_fa467_y2, h_s_dadda_rca32_fa481_y2, h_s_dadda_rca32_fa481_y4);
  fa fa_h_s_dadda_rca32_fa482_y2(h_s_dadda_rca32_fa468_y2, h_s_dadda_rca32_fa469_y2, h_s_dadda_rca32_fa470_y2, h_s_dadda_rca32_fa482_y2, h_s_dadda_rca32_fa482_y4);
  fa fa_h_s_dadda_rca32_fa483_y2(h_s_dadda_rca32_fa471_y2, h_s_dadda_rca32_fa472_y2, h_s_dadda_rca32_fa473_y2, h_s_dadda_rca32_fa483_y2, h_s_dadda_rca32_fa483_y4);
  fa fa_h_s_dadda_rca32_fa484_y2(h_s_dadda_rca32_fa474_y2, h_s_dadda_rca32_fa475_y2, h_s_dadda_rca32_fa476_y2, h_s_dadda_rca32_fa484_y2, h_s_dadda_rca32_fa484_y4);
  fa fa_h_s_dadda_rca32_fa485_y2(h_s_dadda_rca32_fa477_y2, h_s_dadda_rca32_fa478_y2, h_s_dadda_rca32_fa479_y2, h_s_dadda_rca32_fa485_y2, h_s_dadda_rca32_fa485_y4);
  fa fa_h_s_dadda_rca32_fa486_y2(h_s_dadda_rca32_fa485_y4, h_s_dadda_rca32_fa484_y4, h_s_dadda_rca32_fa483_y4, h_s_dadda_rca32_fa486_y2, h_s_dadda_rca32_fa486_y4);
  fa fa_h_s_dadda_rca32_fa487_y2(h_s_dadda_rca32_fa482_y4, h_s_dadda_rca32_fa481_y4, h_s_dadda_rca32_fa480_y4, h_s_dadda_rca32_fa487_y2, h_s_dadda_rca32_fa487_y4);
  fa fa_h_s_dadda_rca32_fa488_y2(h_s_dadda_rca32_fa479_y4, h_s_dadda_rca32_fa478_y4, h_s_dadda_rca32_fa477_y4, h_s_dadda_rca32_fa488_y2, h_s_dadda_rca32_fa488_y4);
  fa fa_h_s_dadda_rca32_fa489_y2(h_s_dadda_rca32_fa476_y4, h_s_dadda_rca32_fa475_y4, h_s_dadda_rca32_fa474_y4, h_s_dadda_rca32_fa489_y2, h_s_dadda_rca32_fa489_y4);
  fa fa_h_s_dadda_rca32_fa490_y2(h_s_dadda_rca32_fa473_y4, h_s_dadda_rca32_fa472_y4, h_s_dadda_rca32_fa471_y4, h_s_dadda_rca32_fa490_y2, h_s_dadda_rca32_fa490_y4);
  fa fa_h_s_dadda_rca32_fa491_y2(h_s_dadda_rca32_fa470_y4, h_s_dadda_rca32_fa469_y4, h_s_dadda_rca32_fa468_y4, h_s_dadda_rca32_fa491_y2, h_s_dadda_rca32_fa491_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_8_y0(a_31, b_8, h_s_dadda_rca32_nand_31_8_y0);
  fa fa_h_s_dadda_rca32_fa492_y2(h_s_dadda_rca32_fa467_y4, h_s_dadda_rca32_fa466_y4, h_s_dadda_rca32_nand_31_8_y0, h_s_dadda_rca32_fa492_y2, h_s_dadda_rca32_fa492_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_9_y0(a_30, b_9, h_s_dadda_rca32_and_30_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_10_y0(a_29, b_10, h_s_dadda_rca32_and_29_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_11_y0(a_28, b_11, h_s_dadda_rca32_and_28_11_y0);
  fa fa_h_s_dadda_rca32_fa493_y2(h_s_dadda_rca32_and_30_9_y0, h_s_dadda_rca32_and_29_10_y0, h_s_dadda_rca32_and_28_11_y0, h_s_dadda_rca32_fa493_y2, h_s_dadda_rca32_fa493_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_12_y0(a_27, b_12, h_s_dadda_rca32_and_27_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_13_y0(a_26, b_13, h_s_dadda_rca32_and_26_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_14_y0(a_25, b_14, h_s_dadda_rca32_and_25_14_y0);
  fa fa_h_s_dadda_rca32_fa494_y2(h_s_dadda_rca32_and_27_12_y0, h_s_dadda_rca32_and_26_13_y0, h_s_dadda_rca32_and_25_14_y0, h_s_dadda_rca32_fa494_y2, h_s_dadda_rca32_fa494_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_15_y0(a_24, b_15, h_s_dadda_rca32_and_24_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_16_y0(a_23, b_16, h_s_dadda_rca32_and_23_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_17_y0(a_22, b_17, h_s_dadda_rca32_and_22_17_y0);
  fa fa_h_s_dadda_rca32_fa495_y2(h_s_dadda_rca32_and_24_15_y0, h_s_dadda_rca32_and_23_16_y0, h_s_dadda_rca32_and_22_17_y0, h_s_dadda_rca32_fa495_y2, h_s_dadda_rca32_fa495_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_18_y0(a_21, b_18, h_s_dadda_rca32_and_21_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_19_y0(a_20, b_19, h_s_dadda_rca32_and_20_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_20_y0(a_19, b_20, h_s_dadda_rca32_and_19_20_y0);
  fa fa_h_s_dadda_rca32_fa496_y2(h_s_dadda_rca32_and_21_18_y0, h_s_dadda_rca32_and_20_19_y0, h_s_dadda_rca32_and_19_20_y0, h_s_dadda_rca32_fa496_y2, h_s_dadda_rca32_fa496_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_21_y0(a_18, b_21, h_s_dadda_rca32_and_18_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_22_y0(a_17, b_22, h_s_dadda_rca32_and_17_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_23_y0(a_16, b_23, h_s_dadda_rca32_and_16_23_y0);
  fa fa_h_s_dadda_rca32_fa497_y2(h_s_dadda_rca32_and_18_21_y0, h_s_dadda_rca32_and_17_22_y0, h_s_dadda_rca32_and_16_23_y0, h_s_dadda_rca32_fa497_y2, h_s_dadda_rca32_fa497_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_24_y0(a_15, b_24, h_s_dadda_rca32_and_15_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_25_y0(a_14, b_25, h_s_dadda_rca32_and_14_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_26_y0(a_13, b_26, h_s_dadda_rca32_and_13_26_y0);
  fa fa_h_s_dadda_rca32_fa498_y2(h_s_dadda_rca32_and_15_24_y0, h_s_dadda_rca32_and_14_25_y0, h_s_dadda_rca32_and_13_26_y0, h_s_dadda_rca32_fa498_y2, h_s_dadda_rca32_fa498_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_27_y0(a_12, b_27, h_s_dadda_rca32_and_12_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_28_y0(a_11, b_28, h_s_dadda_rca32_and_11_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_29_y0(a_10, b_29, h_s_dadda_rca32_and_10_29_y0);
  fa fa_h_s_dadda_rca32_fa499_y2(h_s_dadda_rca32_and_12_27_y0, h_s_dadda_rca32_and_11_28_y0, h_s_dadda_rca32_and_10_29_y0, h_s_dadda_rca32_fa499_y2, h_s_dadda_rca32_fa499_y4);
  and_gate and_gate_h_s_dadda_rca32_and_9_30_y0(a_9, b_30, h_s_dadda_rca32_and_9_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_8_31_y0(a_8, b_31, h_s_dadda_rca32_nand_8_31_y0);
  fa fa_h_s_dadda_rca32_fa500_y2(h_s_dadda_rca32_and_9_30_y0, h_s_dadda_rca32_nand_8_31_y0, h_s_dadda_rca32_fa486_y2, h_s_dadda_rca32_fa500_y2, h_s_dadda_rca32_fa500_y4);
  fa fa_h_s_dadda_rca32_fa501_y2(h_s_dadda_rca32_fa487_y2, h_s_dadda_rca32_fa488_y2, h_s_dadda_rca32_fa489_y2, h_s_dadda_rca32_fa501_y2, h_s_dadda_rca32_fa501_y4);
  fa fa_h_s_dadda_rca32_fa502_y2(h_s_dadda_rca32_fa490_y2, h_s_dadda_rca32_fa491_y2, h_s_dadda_rca32_fa492_y2, h_s_dadda_rca32_fa502_y2, h_s_dadda_rca32_fa502_y4);
  fa fa_h_s_dadda_rca32_fa503_y2(h_s_dadda_rca32_fa493_y2, h_s_dadda_rca32_fa494_y2, h_s_dadda_rca32_fa495_y2, h_s_dadda_rca32_fa503_y2, h_s_dadda_rca32_fa503_y4);
  fa fa_h_s_dadda_rca32_fa504_y2(h_s_dadda_rca32_fa496_y2, h_s_dadda_rca32_fa497_y2, h_s_dadda_rca32_fa498_y2, h_s_dadda_rca32_fa504_y2, h_s_dadda_rca32_fa504_y4);
  fa fa_h_s_dadda_rca32_fa505_y2(h_s_dadda_rca32_fa504_y4, h_s_dadda_rca32_fa503_y4, h_s_dadda_rca32_fa502_y4, h_s_dadda_rca32_fa505_y2, h_s_dadda_rca32_fa505_y4);
  fa fa_h_s_dadda_rca32_fa506_y2(h_s_dadda_rca32_fa501_y4, h_s_dadda_rca32_fa500_y4, h_s_dadda_rca32_fa499_y4, h_s_dadda_rca32_fa506_y2, h_s_dadda_rca32_fa506_y4);
  fa fa_h_s_dadda_rca32_fa507_y2(h_s_dadda_rca32_fa498_y4, h_s_dadda_rca32_fa497_y4, h_s_dadda_rca32_fa496_y4, h_s_dadda_rca32_fa507_y2, h_s_dadda_rca32_fa507_y4);
  fa fa_h_s_dadda_rca32_fa508_y2(h_s_dadda_rca32_fa495_y4, h_s_dadda_rca32_fa494_y4, h_s_dadda_rca32_fa493_y4, h_s_dadda_rca32_fa508_y2, h_s_dadda_rca32_fa508_y4);
  fa fa_h_s_dadda_rca32_fa509_y2(h_s_dadda_rca32_fa492_y4, h_s_dadda_rca32_fa491_y4, h_s_dadda_rca32_fa490_y4, h_s_dadda_rca32_fa509_y2, h_s_dadda_rca32_fa509_y4);
  fa fa_h_s_dadda_rca32_fa510_y2(h_s_dadda_rca32_fa489_y4, h_s_dadda_rca32_fa488_y4, h_s_dadda_rca32_fa487_y4, h_s_dadda_rca32_fa510_y2, h_s_dadda_rca32_fa510_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_9_y0(a_31, b_9, h_s_dadda_rca32_nand_31_9_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_10_y0(a_30, b_10, h_s_dadda_rca32_and_30_10_y0);
  fa fa_h_s_dadda_rca32_fa511_y2(h_s_dadda_rca32_fa486_y4, h_s_dadda_rca32_nand_31_9_y0, h_s_dadda_rca32_and_30_10_y0, h_s_dadda_rca32_fa511_y2, h_s_dadda_rca32_fa511_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_11_y0(a_29, b_11, h_s_dadda_rca32_and_29_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_12_y0(a_28, b_12, h_s_dadda_rca32_and_28_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_13_y0(a_27, b_13, h_s_dadda_rca32_and_27_13_y0);
  fa fa_h_s_dadda_rca32_fa512_y2(h_s_dadda_rca32_and_29_11_y0, h_s_dadda_rca32_and_28_12_y0, h_s_dadda_rca32_and_27_13_y0, h_s_dadda_rca32_fa512_y2, h_s_dadda_rca32_fa512_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_14_y0(a_26, b_14, h_s_dadda_rca32_and_26_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_15_y0(a_25, b_15, h_s_dadda_rca32_and_25_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_16_y0(a_24, b_16, h_s_dadda_rca32_and_24_16_y0);
  fa fa_h_s_dadda_rca32_fa513_y2(h_s_dadda_rca32_and_26_14_y0, h_s_dadda_rca32_and_25_15_y0, h_s_dadda_rca32_and_24_16_y0, h_s_dadda_rca32_fa513_y2, h_s_dadda_rca32_fa513_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_17_y0(a_23, b_17, h_s_dadda_rca32_and_23_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_18_y0(a_22, b_18, h_s_dadda_rca32_and_22_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_19_y0(a_21, b_19, h_s_dadda_rca32_and_21_19_y0);
  fa fa_h_s_dadda_rca32_fa514_y2(h_s_dadda_rca32_and_23_17_y0, h_s_dadda_rca32_and_22_18_y0, h_s_dadda_rca32_and_21_19_y0, h_s_dadda_rca32_fa514_y2, h_s_dadda_rca32_fa514_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_20_y0(a_20, b_20, h_s_dadda_rca32_and_20_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_21_y0(a_19, b_21, h_s_dadda_rca32_and_19_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_22_y0(a_18, b_22, h_s_dadda_rca32_and_18_22_y0);
  fa fa_h_s_dadda_rca32_fa515_y2(h_s_dadda_rca32_and_20_20_y0, h_s_dadda_rca32_and_19_21_y0, h_s_dadda_rca32_and_18_22_y0, h_s_dadda_rca32_fa515_y2, h_s_dadda_rca32_fa515_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_23_y0(a_17, b_23, h_s_dadda_rca32_and_17_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_24_y0(a_16, b_24, h_s_dadda_rca32_and_16_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_25_y0(a_15, b_25, h_s_dadda_rca32_and_15_25_y0);
  fa fa_h_s_dadda_rca32_fa516_y2(h_s_dadda_rca32_and_17_23_y0, h_s_dadda_rca32_and_16_24_y0, h_s_dadda_rca32_and_15_25_y0, h_s_dadda_rca32_fa516_y2, h_s_dadda_rca32_fa516_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_26_y0(a_14, b_26, h_s_dadda_rca32_and_14_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_27_y0(a_13, b_27, h_s_dadda_rca32_and_13_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_28_y0(a_12, b_28, h_s_dadda_rca32_and_12_28_y0);
  fa fa_h_s_dadda_rca32_fa517_y2(h_s_dadda_rca32_and_14_26_y0, h_s_dadda_rca32_and_13_27_y0, h_s_dadda_rca32_and_12_28_y0, h_s_dadda_rca32_fa517_y2, h_s_dadda_rca32_fa517_y4);
  and_gate and_gate_h_s_dadda_rca32_and_11_29_y0(a_11, b_29, h_s_dadda_rca32_and_11_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_10_30_y0(a_10, b_30, h_s_dadda_rca32_and_10_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_9_31_y0(a_9, b_31, h_s_dadda_rca32_nand_9_31_y0);
  fa fa_h_s_dadda_rca32_fa518_y2(h_s_dadda_rca32_and_11_29_y0, h_s_dadda_rca32_and_10_30_y0, h_s_dadda_rca32_nand_9_31_y0, h_s_dadda_rca32_fa518_y2, h_s_dadda_rca32_fa518_y4);
  fa fa_h_s_dadda_rca32_fa519_y2(h_s_dadda_rca32_fa505_y2, h_s_dadda_rca32_fa506_y2, h_s_dadda_rca32_fa507_y2, h_s_dadda_rca32_fa519_y2, h_s_dadda_rca32_fa519_y4);
  fa fa_h_s_dadda_rca32_fa520_y2(h_s_dadda_rca32_fa508_y2, h_s_dadda_rca32_fa509_y2, h_s_dadda_rca32_fa510_y2, h_s_dadda_rca32_fa520_y2, h_s_dadda_rca32_fa520_y4);
  fa fa_h_s_dadda_rca32_fa521_y2(h_s_dadda_rca32_fa511_y2, h_s_dadda_rca32_fa512_y2, h_s_dadda_rca32_fa513_y2, h_s_dadda_rca32_fa521_y2, h_s_dadda_rca32_fa521_y4);
  fa fa_h_s_dadda_rca32_fa522_y2(h_s_dadda_rca32_fa514_y2, h_s_dadda_rca32_fa515_y2, h_s_dadda_rca32_fa516_y2, h_s_dadda_rca32_fa522_y2, h_s_dadda_rca32_fa522_y4);
  fa fa_h_s_dadda_rca32_fa523_y2(h_s_dadda_rca32_fa522_y4, h_s_dadda_rca32_fa521_y4, h_s_dadda_rca32_fa520_y4, h_s_dadda_rca32_fa523_y2, h_s_dadda_rca32_fa523_y4);
  fa fa_h_s_dadda_rca32_fa524_y2(h_s_dadda_rca32_fa519_y4, h_s_dadda_rca32_fa518_y4, h_s_dadda_rca32_fa517_y4, h_s_dadda_rca32_fa524_y2, h_s_dadda_rca32_fa524_y4);
  fa fa_h_s_dadda_rca32_fa525_y2(h_s_dadda_rca32_fa516_y4, h_s_dadda_rca32_fa515_y4, h_s_dadda_rca32_fa514_y4, h_s_dadda_rca32_fa525_y2, h_s_dadda_rca32_fa525_y4);
  fa fa_h_s_dadda_rca32_fa526_y2(h_s_dadda_rca32_fa513_y4, h_s_dadda_rca32_fa512_y4, h_s_dadda_rca32_fa511_y4, h_s_dadda_rca32_fa526_y2, h_s_dadda_rca32_fa526_y4);
  fa fa_h_s_dadda_rca32_fa527_y2(h_s_dadda_rca32_fa510_y4, h_s_dadda_rca32_fa509_y4, h_s_dadda_rca32_fa508_y4, h_s_dadda_rca32_fa527_y2, h_s_dadda_rca32_fa527_y4);
  fa fa_h_s_dadda_rca32_fa528_y2(h_s_dadda_rca32_fa507_y4, h_s_dadda_rca32_fa506_y4, h_s_dadda_rca32_fa505_y4, h_s_dadda_rca32_fa528_y2, h_s_dadda_rca32_fa528_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_10_y0(a_31, b_10, h_s_dadda_rca32_nand_31_10_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_11_y0(a_30, b_11, h_s_dadda_rca32_and_30_11_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_12_y0(a_29, b_12, h_s_dadda_rca32_and_29_12_y0);
  fa fa_h_s_dadda_rca32_fa529_y2(h_s_dadda_rca32_nand_31_10_y0, h_s_dadda_rca32_and_30_11_y0, h_s_dadda_rca32_and_29_12_y0, h_s_dadda_rca32_fa529_y2, h_s_dadda_rca32_fa529_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_13_y0(a_28, b_13, h_s_dadda_rca32_and_28_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_14_y0(a_27, b_14, h_s_dadda_rca32_and_27_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_15_y0(a_26, b_15, h_s_dadda_rca32_and_26_15_y0);
  fa fa_h_s_dadda_rca32_fa530_y2(h_s_dadda_rca32_and_28_13_y0, h_s_dadda_rca32_and_27_14_y0, h_s_dadda_rca32_and_26_15_y0, h_s_dadda_rca32_fa530_y2, h_s_dadda_rca32_fa530_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_16_y0(a_25, b_16, h_s_dadda_rca32_and_25_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_17_y0(a_24, b_17, h_s_dadda_rca32_and_24_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_18_y0(a_23, b_18, h_s_dadda_rca32_and_23_18_y0);
  fa fa_h_s_dadda_rca32_fa531_y2(h_s_dadda_rca32_and_25_16_y0, h_s_dadda_rca32_and_24_17_y0, h_s_dadda_rca32_and_23_18_y0, h_s_dadda_rca32_fa531_y2, h_s_dadda_rca32_fa531_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_19_y0(a_22, b_19, h_s_dadda_rca32_and_22_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_20_y0(a_21, b_20, h_s_dadda_rca32_and_21_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_21_y0(a_20, b_21, h_s_dadda_rca32_and_20_21_y0);
  fa fa_h_s_dadda_rca32_fa532_y2(h_s_dadda_rca32_and_22_19_y0, h_s_dadda_rca32_and_21_20_y0, h_s_dadda_rca32_and_20_21_y0, h_s_dadda_rca32_fa532_y2, h_s_dadda_rca32_fa532_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_22_y0(a_19, b_22, h_s_dadda_rca32_and_19_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_23_y0(a_18, b_23, h_s_dadda_rca32_and_18_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_24_y0(a_17, b_24, h_s_dadda_rca32_and_17_24_y0);
  fa fa_h_s_dadda_rca32_fa533_y2(h_s_dadda_rca32_and_19_22_y0, h_s_dadda_rca32_and_18_23_y0, h_s_dadda_rca32_and_17_24_y0, h_s_dadda_rca32_fa533_y2, h_s_dadda_rca32_fa533_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_25_y0(a_16, b_25, h_s_dadda_rca32_and_16_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_26_y0(a_15, b_26, h_s_dadda_rca32_and_15_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_27_y0(a_14, b_27, h_s_dadda_rca32_and_14_27_y0);
  fa fa_h_s_dadda_rca32_fa534_y2(h_s_dadda_rca32_and_16_25_y0, h_s_dadda_rca32_and_15_26_y0, h_s_dadda_rca32_and_14_27_y0, h_s_dadda_rca32_fa534_y2, h_s_dadda_rca32_fa534_y4);
  and_gate and_gate_h_s_dadda_rca32_and_13_28_y0(a_13, b_28, h_s_dadda_rca32_and_13_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_12_29_y0(a_12, b_29, h_s_dadda_rca32_and_12_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_11_30_y0(a_11, b_30, h_s_dadda_rca32_and_11_30_y0);
  fa fa_h_s_dadda_rca32_fa535_y2(h_s_dadda_rca32_and_13_28_y0, h_s_dadda_rca32_and_12_29_y0, h_s_dadda_rca32_and_11_30_y0, h_s_dadda_rca32_fa535_y2, h_s_dadda_rca32_fa535_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_10_31_y0(a_10, b_31, h_s_dadda_rca32_nand_10_31_y0);
  fa fa_h_s_dadda_rca32_fa536_y2(h_s_dadda_rca32_nand_10_31_y0, h_s_dadda_rca32_fa523_y2, h_s_dadda_rca32_fa524_y2, h_s_dadda_rca32_fa536_y2, h_s_dadda_rca32_fa536_y4);
  fa fa_h_s_dadda_rca32_fa537_y2(h_s_dadda_rca32_fa525_y2, h_s_dadda_rca32_fa526_y2, h_s_dadda_rca32_fa527_y2, h_s_dadda_rca32_fa537_y2, h_s_dadda_rca32_fa537_y4);
  fa fa_h_s_dadda_rca32_fa538_y2(h_s_dadda_rca32_fa528_y2, h_s_dadda_rca32_fa529_y2, h_s_dadda_rca32_fa530_y2, h_s_dadda_rca32_fa538_y2, h_s_dadda_rca32_fa538_y4);
  fa fa_h_s_dadda_rca32_fa539_y2(h_s_dadda_rca32_fa531_y2, h_s_dadda_rca32_fa532_y2, h_s_dadda_rca32_fa533_y2, h_s_dadda_rca32_fa539_y2, h_s_dadda_rca32_fa539_y4);
  fa fa_h_s_dadda_rca32_fa540_y2(h_s_dadda_rca32_fa539_y4, h_s_dadda_rca32_fa538_y4, h_s_dadda_rca32_fa537_y4, h_s_dadda_rca32_fa540_y2, h_s_dadda_rca32_fa540_y4);
  fa fa_h_s_dadda_rca32_fa541_y2(h_s_dadda_rca32_fa536_y4, h_s_dadda_rca32_fa535_y4, h_s_dadda_rca32_fa534_y4, h_s_dadda_rca32_fa541_y2, h_s_dadda_rca32_fa541_y4);
  fa fa_h_s_dadda_rca32_fa542_y2(h_s_dadda_rca32_fa533_y4, h_s_dadda_rca32_fa532_y4, h_s_dadda_rca32_fa531_y4, h_s_dadda_rca32_fa542_y2, h_s_dadda_rca32_fa542_y4);
  fa fa_h_s_dadda_rca32_fa543_y2(h_s_dadda_rca32_fa530_y4, h_s_dadda_rca32_fa529_y4, h_s_dadda_rca32_fa528_y4, h_s_dadda_rca32_fa543_y2, h_s_dadda_rca32_fa543_y4);
  fa fa_h_s_dadda_rca32_fa544_y2(h_s_dadda_rca32_fa527_y4, h_s_dadda_rca32_fa526_y4, h_s_dadda_rca32_fa525_y4, h_s_dadda_rca32_fa544_y2, h_s_dadda_rca32_fa544_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_11_y0(a_31, b_11, h_s_dadda_rca32_nand_31_11_y0);
  fa fa_h_s_dadda_rca32_fa545_y2(h_s_dadda_rca32_fa524_y4, h_s_dadda_rca32_fa523_y4, h_s_dadda_rca32_nand_31_11_y0, h_s_dadda_rca32_fa545_y2, h_s_dadda_rca32_fa545_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_12_y0(a_30, b_12, h_s_dadda_rca32_and_30_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_13_y0(a_29, b_13, h_s_dadda_rca32_and_29_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_14_y0(a_28, b_14, h_s_dadda_rca32_and_28_14_y0);
  fa fa_h_s_dadda_rca32_fa546_y2(h_s_dadda_rca32_and_30_12_y0, h_s_dadda_rca32_and_29_13_y0, h_s_dadda_rca32_and_28_14_y0, h_s_dadda_rca32_fa546_y2, h_s_dadda_rca32_fa546_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_15_y0(a_27, b_15, h_s_dadda_rca32_and_27_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_16_y0(a_26, b_16, h_s_dadda_rca32_and_26_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_17_y0(a_25, b_17, h_s_dadda_rca32_and_25_17_y0);
  fa fa_h_s_dadda_rca32_fa547_y2(h_s_dadda_rca32_and_27_15_y0, h_s_dadda_rca32_and_26_16_y0, h_s_dadda_rca32_and_25_17_y0, h_s_dadda_rca32_fa547_y2, h_s_dadda_rca32_fa547_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_18_y0(a_24, b_18, h_s_dadda_rca32_and_24_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_19_y0(a_23, b_19, h_s_dadda_rca32_and_23_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_20_y0(a_22, b_20, h_s_dadda_rca32_and_22_20_y0);
  fa fa_h_s_dadda_rca32_fa548_y2(h_s_dadda_rca32_and_24_18_y0, h_s_dadda_rca32_and_23_19_y0, h_s_dadda_rca32_and_22_20_y0, h_s_dadda_rca32_fa548_y2, h_s_dadda_rca32_fa548_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_21_y0(a_21, b_21, h_s_dadda_rca32_and_21_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_22_y0(a_20, b_22, h_s_dadda_rca32_and_20_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_23_y0(a_19, b_23, h_s_dadda_rca32_and_19_23_y0);
  fa fa_h_s_dadda_rca32_fa549_y2(h_s_dadda_rca32_and_21_21_y0, h_s_dadda_rca32_and_20_22_y0, h_s_dadda_rca32_and_19_23_y0, h_s_dadda_rca32_fa549_y2, h_s_dadda_rca32_fa549_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_24_y0(a_18, b_24, h_s_dadda_rca32_and_18_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_25_y0(a_17, b_25, h_s_dadda_rca32_and_17_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_26_y0(a_16, b_26, h_s_dadda_rca32_and_16_26_y0);
  fa fa_h_s_dadda_rca32_fa550_y2(h_s_dadda_rca32_and_18_24_y0, h_s_dadda_rca32_and_17_25_y0, h_s_dadda_rca32_and_16_26_y0, h_s_dadda_rca32_fa550_y2, h_s_dadda_rca32_fa550_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_27_y0(a_15, b_27, h_s_dadda_rca32_and_15_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_28_y0(a_14, b_28, h_s_dadda_rca32_and_14_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_29_y0(a_13, b_29, h_s_dadda_rca32_and_13_29_y0);
  fa fa_h_s_dadda_rca32_fa551_y2(h_s_dadda_rca32_and_15_27_y0, h_s_dadda_rca32_and_14_28_y0, h_s_dadda_rca32_and_13_29_y0, h_s_dadda_rca32_fa551_y2, h_s_dadda_rca32_fa551_y4);
  and_gate and_gate_h_s_dadda_rca32_and_12_30_y0(a_12, b_30, h_s_dadda_rca32_and_12_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_11_31_y0(a_11, b_31, h_s_dadda_rca32_nand_11_31_y0);
  fa fa_h_s_dadda_rca32_fa552_y2(h_s_dadda_rca32_and_12_30_y0, h_s_dadda_rca32_nand_11_31_y0, h_s_dadda_rca32_fa540_y2, h_s_dadda_rca32_fa552_y2, h_s_dadda_rca32_fa552_y4);
  fa fa_h_s_dadda_rca32_fa553_y2(h_s_dadda_rca32_fa541_y2, h_s_dadda_rca32_fa542_y2, h_s_dadda_rca32_fa543_y2, h_s_dadda_rca32_fa553_y2, h_s_dadda_rca32_fa553_y4);
  fa fa_h_s_dadda_rca32_fa554_y2(h_s_dadda_rca32_fa544_y2, h_s_dadda_rca32_fa545_y2, h_s_dadda_rca32_fa546_y2, h_s_dadda_rca32_fa554_y2, h_s_dadda_rca32_fa554_y4);
  fa fa_h_s_dadda_rca32_fa555_y2(h_s_dadda_rca32_fa547_y2, h_s_dadda_rca32_fa548_y2, h_s_dadda_rca32_fa549_y2, h_s_dadda_rca32_fa555_y2, h_s_dadda_rca32_fa555_y4);
  fa fa_h_s_dadda_rca32_fa556_y2(h_s_dadda_rca32_fa555_y4, h_s_dadda_rca32_fa554_y4, h_s_dadda_rca32_fa553_y4, h_s_dadda_rca32_fa556_y2, h_s_dadda_rca32_fa556_y4);
  fa fa_h_s_dadda_rca32_fa557_y2(h_s_dadda_rca32_fa552_y4, h_s_dadda_rca32_fa551_y4, h_s_dadda_rca32_fa550_y4, h_s_dadda_rca32_fa557_y2, h_s_dadda_rca32_fa557_y4);
  fa fa_h_s_dadda_rca32_fa558_y2(h_s_dadda_rca32_fa549_y4, h_s_dadda_rca32_fa548_y4, h_s_dadda_rca32_fa547_y4, h_s_dadda_rca32_fa558_y2, h_s_dadda_rca32_fa558_y4);
  fa fa_h_s_dadda_rca32_fa559_y2(h_s_dadda_rca32_fa546_y4, h_s_dadda_rca32_fa545_y4, h_s_dadda_rca32_fa544_y4, h_s_dadda_rca32_fa559_y2, h_s_dadda_rca32_fa559_y4);
  fa fa_h_s_dadda_rca32_fa560_y2(h_s_dadda_rca32_fa543_y4, h_s_dadda_rca32_fa542_y4, h_s_dadda_rca32_fa541_y4, h_s_dadda_rca32_fa560_y2, h_s_dadda_rca32_fa560_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_12_y0(a_31, b_12, h_s_dadda_rca32_nand_31_12_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_13_y0(a_30, b_13, h_s_dadda_rca32_and_30_13_y0);
  fa fa_h_s_dadda_rca32_fa561_y2(h_s_dadda_rca32_fa540_y4, h_s_dadda_rca32_nand_31_12_y0, h_s_dadda_rca32_and_30_13_y0, h_s_dadda_rca32_fa561_y2, h_s_dadda_rca32_fa561_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_14_y0(a_29, b_14, h_s_dadda_rca32_and_29_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_15_y0(a_28, b_15, h_s_dadda_rca32_and_28_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_16_y0(a_27, b_16, h_s_dadda_rca32_and_27_16_y0);
  fa fa_h_s_dadda_rca32_fa562_y2(h_s_dadda_rca32_and_29_14_y0, h_s_dadda_rca32_and_28_15_y0, h_s_dadda_rca32_and_27_16_y0, h_s_dadda_rca32_fa562_y2, h_s_dadda_rca32_fa562_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_17_y0(a_26, b_17, h_s_dadda_rca32_and_26_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_18_y0(a_25, b_18, h_s_dadda_rca32_and_25_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_19_y0(a_24, b_19, h_s_dadda_rca32_and_24_19_y0);
  fa fa_h_s_dadda_rca32_fa563_y2(h_s_dadda_rca32_and_26_17_y0, h_s_dadda_rca32_and_25_18_y0, h_s_dadda_rca32_and_24_19_y0, h_s_dadda_rca32_fa563_y2, h_s_dadda_rca32_fa563_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_20_y0(a_23, b_20, h_s_dadda_rca32_and_23_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_21_y0(a_22, b_21, h_s_dadda_rca32_and_22_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_22_y0(a_21, b_22, h_s_dadda_rca32_and_21_22_y0);
  fa fa_h_s_dadda_rca32_fa564_y2(h_s_dadda_rca32_and_23_20_y0, h_s_dadda_rca32_and_22_21_y0, h_s_dadda_rca32_and_21_22_y0, h_s_dadda_rca32_fa564_y2, h_s_dadda_rca32_fa564_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_23_y0(a_20, b_23, h_s_dadda_rca32_and_20_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_24_y0(a_19, b_24, h_s_dadda_rca32_and_19_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_25_y0(a_18, b_25, h_s_dadda_rca32_and_18_25_y0);
  fa fa_h_s_dadda_rca32_fa565_y2(h_s_dadda_rca32_and_20_23_y0, h_s_dadda_rca32_and_19_24_y0, h_s_dadda_rca32_and_18_25_y0, h_s_dadda_rca32_fa565_y2, h_s_dadda_rca32_fa565_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_26_y0(a_17, b_26, h_s_dadda_rca32_and_17_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_27_y0(a_16, b_27, h_s_dadda_rca32_and_16_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_28_y0(a_15, b_28, h_s_dadda_rca32_and_15_28_y0);
  fa fa_h_s_dadda_rca32_fa566_y2(h_s_dadda_rca32_and_17_26_y0, h_s_dadda_rca32_and_16_27_y0, h_s_dadda_rca32_and_15_28_y0, h_s_dadda_rca32_fa566_y2, h_s_dadda_rca32_fa566_y4);
  and_gate and_gate_h_s_dadda_rca32_and_14_29_y0(a_14, b_29, h_s_dadda_rca32_and_14_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_13_30_y0(a_13, b_30, h_s_dadda_rca32_and_13_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_12_31_y0(a_12, b_31, h_s_dadda_rca32_nand_12_31_y0);
  fa fa_h_s_dadda_rca32_fa567_y2(h_s_dadda_rca32_and_14_29_y0, h_s_dadda_rca32_and_13_30_y0, h_s_dadda_rca32_nand_12_31_y0, h_s_dadda_rca32_fa567_y2, h_s_dadda_rca32_fa567_y4);
  fa fa_h_s_dadda_rca32_fa568_y2(h_s_dadda_rca32_fa556_y2, h_s_dadda_rca32_fa557_y2, h_s_dadda_rca32_fa558_y2, h_s_dadda_rca32_fa568_y2, h_s_dadda_rca32_fa568_y4);
  fa fa_h_s_dadda_rca32_fa569_y2(h_s_dadda_rca32_fa559_y2, h_s_dadda_rca32_fa560_y2, h_s_dadda_rca32_fa561_y2, h_s_dadda_rca32_fa569_y2, h_s_dadda_rca32_fa569_y4);
  fa fa_h_s_dadda_rca32_fa570_y2(h_s_dadda_rca32_fa562_y2, h_s_dadda_rca32_fa563_y2, h_s_dadda_rca32_fa564_y2, h_s_dadda_rca32_fa570_y2, h_s_dadda_rca32_fa570_y4);
  fa fa_h_s_dadda_rca32_fa571_y2(h_s_dadda_rca32_fa570_y4, h_s_dadda_rca32_fa569_y4, h_s_dadda_rca32_fa568_y4, h_s_dadda_rca32_fa571_y2, h_s_dadda_rca32_fa571_y4);
  fa fa_h_s_dadda_rca32_fa572_y2(h_s_dadda_rca32_fa567_y4, h_s_dadda_rca32_fa566_y4, h_s_dadda_rca32_fa565_y4, h_s_dadda_rca32_fa572_y2, h_s_dadda_rca32_fa572_y4);
  fa fa_h_s_dadda_rca32_fa573_y2(h_s_dadda_rca32_fa564_y4, h_s_dadda_rca32_fa563_y4, h_s_dadda_rca32_fa562_y4, h_s_dadda_rca32_fa573_y2, h_s_dadda_rca32_fa573_y4);
  fa fa_h_s_dadda_rca32_fa574_y2(h_s_dadda_rca32_fa561_y4, h_s_dadda_rca32_fa560_y4, h_s_dadda_rca32_fa559_y4, h_s_dadda_rca32_fa574_y2, h_s_dadda_rca32_fa574_y4);
  fa fa_h_s_dadda_rca32_fa575_y2(h_s_dadda_rca32_fa558_y4, h_s_dadda_rca32_fa557_y4, h_s_dadda_rca32_fa556_y4, h_s_dadda_rca32_fa575_y2, h_s_dadda_rca32_fa575_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_13_y0(a_31, b_13, h_s_dadda_rca32_nand_31_13_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_14_y0(a_30, b_14, h_s_dadda_rca32_and_30_14_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_15_y0(a_29, b_15, h_s_dadda_rca32_and_29_15_y0);
  fa fa_h_s_dadda_rca32_fa576_y2(h_s_dadda_rca32_nand_31_13_y0, h_s_dadda_rca32_and_30_14_y0, h_s_dadda_rca32_and_29_15_y0, h_s_dadda_rca32_fa576_y2, h_s_dadda_rca32_fa576_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_16_y0(a_28, b_16, h_s_dadda_rca32_and_28_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_17_y0(a_27, b_17, h_s_dadda_rca32_and_27_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_18_y0(a_26, b_18, h_s_dadda_rca32_and_26_18_y0);
  fa fa_h_s_dadda_rca32_fa577_y2(h_s_dadda_rca32_and_28_16_y0, h_s_dadda_rca32_and_27_17_y0, h_s_dadda_rca32_and_26_18_y0, h_s_dadda_rca32_fa577_y2, h_s_dadda_rca32_fa577_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_19_y0(a_25, b_19, h_s_dadda_rca32_and_25_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_20_y0(a_24, b_20, h_s_dadda_rca32_and_24_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_21_y0(a_23, b_21, h_s_dadda_rca32_and_23_21_y0);
  fa fa_h_s_dadda_rca32_fa578_y2(h_s_dadda_rca32_and_25_19_y0, h_s_dadda_rca32_and_24_20_y0, h_s_dadda_rca32_and_23_21_y0, h_s_dadda_rca32_fa578_y2, h_s_dadda_rca32_fa578_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_22_y0(a_22, b_22, h_s_dadda_rca32_and_22_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_23_y0(a_21, b_23, h_s_dadda_rca32_and_21_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_24_y0(a_20, b_24, h_s_dadda_rca32_and_20_24_y0);
  fa fa_h_s_dadda_rca32_fa579_y2(h_s_dadda_rca32_and_22_22_y0, h_s_dadda_rca32_and_21_23_y0, h_s_dadda_rca32_and_20_24_y0, h_s_dadda_rca32_fa579_y2, h_s_dadda_rca32_fa579_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_25_y0(a_19, b_25, h_s_dadda_rca32_and_19_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_26_y0(a_18, b_26, h_s_dadda_rca32_and_18_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_27_y0(a_17, b_27, h_s_dadda_rca32_and_17_27_y0);
  fa fa_h_s_dadda_rca32_fa580_y2(h_s_dadda_rca32_and_19_25_y0, h_s_dadda_rca32_and_18_26_y0, h_s_dadda_rca32_and_17_27_y0, h_s_dadda_rca32_fa580_y2, h_s_dadda_rca32_fa580_y4);
  and_gate and_gate_h_s_dadda_rca32_and_16_28_y0(a_16, b_28, h_s_dadda_rca32_and_16_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_15_29_y0(a_15, b_29, h_s_dadda_rca32_and_15_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_14_30_y0(a_14, b_30, h_s_dadda_rca32_and_14_30_y0);
  fa fa_h_s_dadda_rca32_fa581_y2(h_s_dadda_rca32_and_16_28_y0, h_s_dadda_rca32_and_15_29_y0, h_s_dadda_rca32_and_14_30_y0, h_s_dadda_rca32_fa581_y2, h_s_dadda_rca32_fa581_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_13_31_y0(a_13, b_31, h_s_dadda_rca32_nand_13_31_y0);
  fa fa_h_s_dadda_rca32_fa582_y2(h_s_dadda_rca32_nand_13_31_y0, h_s_dadda_rca32_fa571_y2, h_s_dadda_rca32_fa572_y2, h_s_dadda_rca32_fa582_y2, h_s_dadda_rca32_fa582_y4);
  fa fa_h_s_dadda_rca32_fa583_y2(h_s_dadda_rca32_fa573_y2, h_s_dadda_rca32_fa574_y2, h_s_dadda_rca32_fa575_y2, h_s_dadda_rca32_fa583_y2, h_s_dadda_rca32_fa583_y4);
  fa fa_h_s_dadda_rca32_fa584_y2(h_s_dadda_rca32_fa576_y2, h_s_dadda_rca32_fa577_y2, h_s_dadda_rca32_fa578_y2, h_s_dadda_rca32_fa584_y2, h_s_dadda_rca32_fa584_y4);
  fa fa_h_s_dadda_rca32_fa585_y2(h_s_dadda_rca32_fa584_y4, h_s_dadda_rca32_fa583_y4, h_s_dadda_rca32_fa582_y4, h_s_dadda_rca32_fa585_y2, h_s_dadda_rca32_fa585_y4);
  fa fa_h_s_dadda_rca32_fa586_y2(h_s_dadda_rca32_fa581_y4, h_s_dadda_rca32_fa580_y4, h_s_dadda_rca32_fa579_y4, h_s_dadda_rca32_fa586_y2, h_s_dadda_rca32_fa586_y4);
  fa fa_h_s_dadda_rca32_fa587_y2(h_s_dadda_rca32_fa578_y4, h_s_dadda_rca32_fa577_y4, h_s_dadda_rca32_fa576_y4, h_s_dadda_rca32_fa587_y2, h_s_dadda_rca32_fa587_y4);
  fa fa_h_s_dadda_rca32_fa588_y2(h_s_dadda_rca32_fa575_y4, h_s_dadda_rca32_fa574_y4, h_s_dadda_rca32_fa573_y4, h_s_dadda_rca32_fa588_y2, h_s_dadda_rca32_fa588_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_14_y0(a_31, b_14, h_s_dadda_rca32_nand_31_14_y0);
  fa fa_h_s_dadda_rca32_fa589_y2(h_s_dadda_rca32_fa572_y4, h_s_dadda_rca32_fa571_y4, h_s_dadda_rca32_nand_31_14_y0, h_s_dadda_rca32_fa589_y2, h_s_dadda_rca32_fa589_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_15_y0(a_30, b_15, h_s_dadda_rca32_and_30_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_16_y0(a_29, b_16, h_s_dadda_rca32_and_29_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_17_y0(a_28, b_17, h_s_dadda_rca32_and_28_17_y0);
  fa fa_h_s_dadda_rca32_fa590_y2(h_s_dadda_rca32_and_30_15_y0, h_s_dadda_rca32_and_29_16_y0, h_s_dadda_rca32_and_28_17_y0, h_s_dadda_rca32_fa590_y2, h_s_dadda_rca32_fa590_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_18_y0(a_27, b_18, h_s_dadda_rca32_and_27_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_19_y0(a_26, b_19, h_s_dadda_rca32_and_26_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_20_y0(a_25, b_20, h_s_dadda_rca32_and_25_20_y0);
  fa fa_h_s_dadda_rca32_fa591_y2(h_s_dadda_rca32_and_27_18_y0, h_s_dadda_rca32_and_26_19_y0, h_s_dadda_rca32_and_25_20_y0, h_s_dadda_rca32_fa591_y2, h_s_dadda_rca32_fa591_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_21_y0(a_24, b_21, h_s_dadda_rca32_and_24_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_22_y0(a_23, b_22, h_s_dadda_rca32_and_23_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_23_y0(a_22, b_23, h_s_dadda_rca32_and_22_23_y0);
  fa fa_h_s_dadda_rca32_fa592_y2(h_s_dadda_rca32_and_24_21_y0, h_s_dadda_rca32_and_23_22_y0, h_s_dadda_rca32_and_22_23_y0, h_s_dadda_rca32_fa592_y2, h_s_dadda_rca32_fa592_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_24_y0(a_21, b_24, h_s_dadda_rca32_and_21_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_25_y0(a_20, b_25, h_s_dadda_rca32_and_20_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_26_y0(a_19, b_26, h_s_dadda_rca32_and_19_26_y0);
  fa fa_h_s_dadda_rca32_fa593_y2(h_s_dadda_rca32_and_21_24_y0, h_s_dadda_rca32_and_20_25_y0, h_s_dadda_rca32_and_19_26_y0, h_s_dadda_rca32_fa593_y2, h_s_dadda_rca32_fa593_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_27_y0(a_18, b_27, h_s_dadda_rca32_and_18_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_28_y0(a_17, b_28, h_s_dadda_rca32_and_17_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_29_y0(a_16, b_29, h_s_dadda_rca32_and_16_29_y0);
  fa fa_h_s_dadda_rca32_fa594_y2(h_s_dadda_rca32_and_18_27_y0, h_s_dadda_rca32_and_17_28_y0, h_s_dadda_rca32_and_16_29_y0, h_s_dadda_rca32_fa594_y2, h_s_dadda_rca32_fa594_y4);
  and_gate and_gate_h_s_dadda_rca32_and_15_30_y0(a_15, b_30, h_s_dadda_rca32_and_15_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_14_31_y0(a_14, b_31, h_s_dadda_rca32_nand_14_31_y0);
  fa fa_h_s_dadda_rca32_fa595_y2(h_s_dadda_rca32_and_15_30_y0, h_s_dadda_rca32_nand_14_31_y0, h_s_dadda_rca32_fa585_y2, h_s_dadda_rca32_fa595_y2, h_s_dadda_rca32_fa595_y4);
  fa fa_h_s_dadda_rca32_fa596_y2(h_s_dadda_rca32_fa586_y2, h_s_dadda_rca32_fa587_y2, h_s_dadda_rca32_fa588_y2, h_s_dadda_rca32_fa596_y2, h_s_dadda_rca32_fa596_y4);
  fa fa_h_s_dadda_rca32_fa597_y2(h_s_dadda_rca32_fa589_y2, h_s_dadda_rca32_fa590_y2, h_s_dadda_rca32_fa591_y2, h_s_dadda_rca32_fa597_y2, h_s_dadda_rca32_fa597_y4);
  fa fa_h_s_dadda_rca32_fa598_y2(h_s_dadda_rca32_fa597_y4, h_s_dadda_rca32_fa596_y4, h_s_dadda_rca32_fa595_y4, h_s_dadda_rca32_fa598_y2, h_s_dadda_rca32_fa598_y4);
  fa fa_h_s_dadda_rca32_fa599_y2(h_s_dadda_rca32_fa594_y4, h_s_dadda_rca32_fa593_y4, h_s_dadda_rca32_fa592_y4, h_s_dadda_rca32_fa599_y2, h_s_dadda_rca32_fa599_y4);
  fa fa_h_s_dadda_rca32_fa600_y2(h_s_dadda_rca32_fa591_y4, h_s_dadda_rca32_fa590_y4, h_s_dadda_rca32_fa589_y4, h_s_dadda_rca32_fa600_y2, h_s_dadda_rca32_fa600_y4);
  fa fa_h_s_dadda_rca32_fa601_y2(h_s_dadda_rca32_fa588_y4, h_s_dadda_rca32_fa587_y4, h_s_dadda_rca32_fa586_y4, h_s_dadda_rca32_fa601_y2, h_s_dadda_rca32_fa601_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_15_y0(a_31, b_15, h_s_dadda_rca32_nand_31_15_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_16_y0(a_30, b_16, h_s_dadda_rca32_and_30_16_y0);
  fa fa_h_s_dadda_rca32_fa602_y2(h_s_dadda_rca32_fa585_y4, h_s_dadda_rca32_nand_31_15_y0, h_s_dadda_rca32_and_30_16_y0, h_s_dadda_rca32_fa602_y2, h_s_dadda_rca32_fa602_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_17_y0(a_29, b_17, h_s_dadda_rca32_and_29_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_18_y0(a_28, b_18, h_s_dadda_rca32_and_28_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_19_y0(a_27, b_19, h_s_dadda_rca32_and_27_19_y0);
  fa fa_h_s_dadda_rca32_fa603_y2(h_s_dadda_rca32_and_29_17_y0, h_s_dadda_rca32_and_28_18_y0, h_s_dadda_rca32_and_27_19_y0, h_s_dadda_rca32_fa603_y2, h_s_dadda_rca32_fa603_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_20_y0(a_26, b_20, h_s_dadda_rca32_and_26_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_21_y0(a_25, b_21, h_s_dadda_rca32_and_25_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_22_y0(a_24, b_22, h_s_dadda_rca32_and_24_22_y0);
  fa fa_h_s_dadda_rca32_fa604_y2(h_s_dadda_rca32_and_26_20_y0, h_s_dadda_rca32_and_25_21_y0, h_s_dadda_rca32_and_24_22_y0, h_s_dadda_rca32_fa604_y2, h_s_dadda_rca32_fa604_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_23_y0(a_23, b_23, h_s_dadda_rca32_and_23_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_24_y0(a_22, b_24, h_s_dadda_rca32_and_22_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_25_y0(a_21, b_25, h_s_dadda_rca32_and_21_25_y0);
  fa fa_h_s_dadda_rca32_fa605_y2(h_s_dadda_rca32_and_23_23_y0, h_s_dadda_rca32_and_22_24_y0, h_s_dadda_rca32_and_21_25_y0, h_s_dadda_rca32_fa605_y2, h_s_dadda_rca32_fa605_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_26_y0(a_20, b_26, h_s_dadda_rca32_and_20_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_27_y0(a_19, b_27, h_s_dadda_rca32_and_19_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_28_y0(a_18, b_28, h_s_dadda_rca32_and_18_28_y0);
  fa fa_h_s_dadda_rca32_fa606_y2(h_s_dadda_rca32_and_20_26_y0, h_s_dadda_rca32_and_19_27_y0, h_s_dadda_rca32_and_18_28_y0, h_s_dadda_rca32_fa606_y2, h_s_dadda_rca32_fa606_y4);
  and_gate and_gate_h_s_dadda_rca32_and_17_29_y0(a_17, b_29, h_s_dadda_rca32_and_17_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_16_30_y0(a_16, b_30, h_s_dadda_rca32_and_16_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_15_31_y0(a_15, b_31, h_s_dadda_rca32_nand_15_31_y0);
  fa fa_h_s_dadda_rca32_fa607_y2(h_s_dadda_rca32_and_17_29_y0, h_s_dadda_rca32_and_16_30_y0, h_s_dadda_rca32_nand_15_31_y0, h_s_dadda_rca32_fa607_y2, h_s_dadda_rca32_fa607_y4);
  fa fa_h_s_dadda_rca32_fa608_y2(h_s_dadda_rca32_fa598_y2, h_s_dadda_rca32_fa599_y2, h_s_dadda_rca32_fa600_y2, h_s_dadda_rca32_fa608_y2, h_s_dadda_rca32_fa608_y4);
  fa fa_h_s_dadda_rca32_fa609_y2(h_s_dadda_rca32_fa601_y2, h_s_dadda_rca32_fa602_y2, h_s_dadda_rca32_fa603_y2, h_s_dadda_rca32_fa609_y2, h_s_dadda_rca32_fa609_y4);
  fa fa_h_s_dadda_rca32_fa610_y2(h_s_dadda_rca32_fa609_y4, h_s_dadda_rca32_fa608_y4, h_s_dadda_rca32_fa607_y4, h_s_dadda_rca32_fa610_y2, h_s_dadda_rca32_fa610_y4);
  fa fa_h_s_dadda_rca32_fa611_y2(h_s_dadda_rca32_fa606_y4, h_s_dadda_rca32_fa605_y4, h_s_dadda_rca32_fa604_y4, h_s_dadda_rca32_fa611_y2, h_s_dadda_rca32_fa611_y4);
  fa fa_h_s_dadda_rca32_fa612_y2(h_s_dadda_rca32_fa603_y4, h_s_dadda_rca32_fa602_y4, h_s_dadda_rca32_fa601_y4, h_s_dadda_rca32_fa612_y2, h_s_dadda_rca32_fa612_y4);
  fa fa_h_s_dadda_rca32_fa613_y2(h_s_dadda_rca32_fa600_y4, h_s_dadda_rca32_fa599_y4, h_s_dadda_rca32_fa598_y4, h_s_dadda_rca32_fa613_y2, h_s_dadda_rca32_fa613_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_16_y0(a_31, b_16, h_s_dadda_rca32_nand_31_16_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_17_y0(a_30, b_17, h_s_dadda_rca32_and_30_17_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_18_y0(a_29, b_18, h_s_dadda_rca32_and_29_18_y0);
  fa fa_h_s_dadda_rca32_fa614_y2(h_s_dadda_rca32_nand_31_16_y0, h_s_dadda_rca32_and_30_17_y0, h_s_dadda_rca32_and_29_18_y0, h_s_dadda_rca32_fa614_y2, h_s_dadda_rca32_fa614_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_19_y0(a_28, b_19, h_s_dadda_rca32_and_28_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_20_y0(a_27, b_20, h_s_dadda_rca32_and_27_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_21_y0(a_26, b_21, h_s_dadda_rca32_and_26_21_y0);
  fa fa_h_s_dadda_rca32_fa615_y2(h_s_dadda_rca32_and_28_19_y0, h_s_dadda_rca32_and_27_20_y0, h_s_dadda_rca32_and_26_21_y0, h_s_dadda_rca32_fa615_y2, h_s_dadda_rca32_fa615_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_22_y0(a_25, b_22, h_s_dadda_rca32_and_25_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_23_y0(a_24, b_23, h_s_dadda_rca32_and_24_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_24_y0(a_23, b_24, h_s_dadda_rca32_and_23_24_y0);
  fa fa_h_s_dadda_rca32_fa616_y2(h_s_dadda_rca32_and_25_22_y0, h_s_dadda_rca32_and_24_23_y0, h_s_dadda_rca32_and_23_24_y0, h_s_dadda_rca32_fa616_y2, h_s_dadda_rca32_fa616_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_25_y0(a_22, b_25, h_s_dadda_rca32_and_22_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_26_y0(a_21, b_26, h_s_dadda_rca32_and_21_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_27_y0(a_20, b_27, h_s_dadda_rca32_and_20_27_y0);
  fa fa_h_s_dadda_rca32_fa617_y2(h_s_dadda_rca32_and_22_25_y0, h_s_dadda_rca32_and_21_26_y0, h_s_dadda_rca32_and_20_27_y0, h_s_dadda_rca32_fa617_y2, h_s_dadda_rca32_fa617_y4);
  and_gate and_gate_h_s_dadda_rca32_and_19_28_y0(a_19, b_28, h_s_dadda_rca32_and_19_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_18_29_y0(a_18, b_29, h_s_dadda_rca32_and_18_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_17_30_y0(a_17, b_30, h_s_dadda_rca32_and_17_30_y0);
  fa fa_h_s_dadda_rca32_fa618_y2(h_s_dadda_rca32_and_19_28_y0, h_s_dadda_rca32_and_18_29_y0, h_s_dadda_rca32_and_17_30_y0, h_s_dadda_rca32_fa618_y2, h_s_dadda_rca32_fa618_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_16_31_y0(a_16, b_31, h_s_dadda_rca32_nand_16_31_y0);
  fa fa_h_s_dadda_rca32_fa619_y2(h_s_dadda_rca32_nand_16_31_y0, h_s_dadda_rca32_fa610_y2, h_s_dadda_rca32_fa611_y2, h_s_dadda_rca32_fa619_y2, h_s_dadda_rca32_fa619_y4);
  fa fa_h_s_dadda_rca32_fa620_y2(h_s_dadda_rca32_fa612_y2, h_s_dadda_rca32_fa613_y2, h_s_dadda_rca32_fa614_y2, h_s_dadda_rca32_fa620_y2, h_s_dadda_rca32_fa620_y4);
  fa fa_h_s_dadda_rca32_fa621_y2(h_s_dadda_rca32_fa620_y4, h_s_dadda_rca32_fa619_y4, h_s_dadda_rca32_fa618_y4, h_s_dadda_rca32_fa621_y2, h_s_dadda_rca32_fa621_y4);
  fa fa_h_s_dadda_rca32_fa622_y2(h_s_dadda_rca32_fa617_y4, h_s_dadda_rca32_fa616_y4, h_s_dadda_rca32_fa615_y4, h_s_dadda_rca32_fa622_y2, h_s_dadda_rca32_fa622_y4);
  fa fa_h_s_dadda_rca32_fa623_y2(h_s_dadda_rca32_fa614_y4, h_s_dadda_rca32_fa613_y4, h_s_dadda_rca32_fa612_y4, h_s_dadda_rca32_fa623_y2, h_s_dadda_rca32_fa623_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_17_y0(a_31, b_17, h_s_dadda_rca32_nand_31_17_y0);
  fa fa_h_s_dadda_rca32_fa624_y2(h_s_dadda_rca32_fa611_y4, h_s_dadda_rca32_fa610_y4, h_s_dadda_rca32_nand_31_17_y0, h_s_dadda_rca32_fa624_y2, h_s_dadda_rca32_fa624_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_18_y0(a_30, b_18, h_s_dadda_rca32_and_30_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_19_y0(a_29, b_19, h_s_dadda_rca32_and_29_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_20_y0(a_28, b_20, h_s_dadda_rca32_and_28_20_y0);
  fa fa_h_s_dadda_rca32_fa625_y2(h_s_dadda_rca32_and_30_18_y0, h_s_dadda_rca32_and_29_19_y0, h_s_dadda_rca32_and_28_20_y0, h_s_dadda_rca32_fa625_y2, h_s_dadda_rca32_fa625_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_21_y0(a_27, b_21, h_s_dadda_rca32_and_27_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_22_y0(a_26, b_22, h_s_dadda_rca32_and_26_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_23_y0(a_25, b_23, h_s_dadda_rca32_and_25_23_y0);
  fa fa_h_s_dadda_rca32_fa626_y2(h_s_dadda_rca32_and_27_21_y0, h_s_dadda_rca32_and_26_22_y0, h_s_dadda_rca32_and_25_23_y0, h_s_dadda_rca32_fa626_y2, h_s_dadda_rca32_fa626_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_24_y0(a_24, b_24, h_s_dadda_rca32_and_24_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_25_y0(a_23, b_25, h_s_dadda_rca32_and_23_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_26_y0(a_22, b_26, h_s_dadda_rca32_and_22_26_y0);
  fa fa_h_s_dadda_rca32_fa627_y2(h_s_dadda_rca32_and_24_24_y0, h_s_dadda_rca32_and_23_25_y0, h_s_dadda_rca32_and_22_26_y0, h_s_dadda_rca32_fa627_y2, h_s_dadda_rca32_fa627_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_27_y0(a_21, b_27, h_s_dadda_rca32_and_21_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_28_y0(a_20, b_28, h_s_dadda_rca32_and_20_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_29_y0(a_19, b_29, h_s_dadda_rca32_and_19_29_y0);
  fa fa_h_s_dadda_rca32_fa628_y2(h_s_dadda_rca32_and_21_27_y0, h_s_dadda_rca32_and_20_28_y0, h_s_dadda_rca32_and_19_29_y0, h_s_dadda_rca32_fa628_y2, h_s_dadda_rca32_fa628_y4);
  and_gate and_gate_h_s_dadda_rca32_and_18_30_y0(a_18, b_30, h_s_dadda_rca32_and_18_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_17_31_y0(a_17, b_31, h_s_dadda_rca32_nand_17_31_y0);
  fa fa_h_s_dadda_rca32_fa629_y2(h_s_dadda_rca32_and_18_30_y0, h_s_dadda_rca32_nand_17_31_y0, h_s_dadda_rca32_fa621_y2, h_s_dadda_rca32_fa629_y2, h_s_dadda_rca32_fa629_y4);
  fa fa_h_s_dadda_rca32_fa630_y2(h_s_dadda_rca32_fa622_y2, h_s_dadda_rca32_fa623_y2, h_s_dadda_rca32_fa624_y2, h_s_dadda_rca32_fa630_y2, h_s_dadda_rca32_fa630_y4);
  fa fa_h_s_dadda_rca32_fa631_y2(h_s_dadda_rca32_fa630_y4, h_s_dadda_rca32_fa629_y4, h_s_dadda_rca32_fa628_y4, h_s_dadda_rca32_fa631_y2, h_s_dadda_rca32_fa631_y4);
  fa fa_h_s_dadda_rca32_fa632_y2(h_s_dadda_rca32_fa627_y4, h_s_dadda_rca32_fa626_y4, h_s_dadda_rca32_fa625_y4, h_s_dadda_rca32_fa632_y2, h_s_dadda_rca32_fa632_y4);
  fa fa_h_s_dadda_rca32_fa633_y2(h_s_dadda_rca32_fa624_y4, h_s_dadda_rca32_fa623_y4, h_s_dadda_rca32_fa622_y4, h_s_dadda_rca32_fa633_y2, h_s_dadda_rca32_fa633_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_18_y0(a_31, b_18, h_s_dadda_rca32_nand_31_18_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_19_y0(a_30, b_19, h_s_dadda_rca32_and_30_19_y0);
  fa fa_h_s_dadda_rca32_fa634_y2(h_s_dadda_rca32_fa621_y4, h_s_dadda_rca32_nand_31_18_y0, h_s_dadda_rca32_and_30_19_y0, h_s_dadda_rca32_fa634_y2, h_s_dadda_rca32_fa634_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_20_y0(a_29, b_20, h_s_dadda_rca32_and_29_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_21_y0(a_28, b_21, h_s_dadda_rca32_and_28_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_22_y0(a_27, b_22, h_s_dadda_rca32_and_27_22_y0);
  fa fa_h_s_dadda_rca32_fa635_y2(h_s_dadda_rca32_and_29_20_y0, h_s_dadda_rca32_and_28_21_y0, h_s_dadda_rca32_and_27_22_y0, h_s_dadda_rca32_fa635_y2, h_s_dadda_rca32_fa635_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_23_y0(a_26, b_23, h_s_dadda_rca32_and_26_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_24_y0(a_25, b_24, h_s_dadda_rca32_and_25_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_25_y0(a_24, b_25, h_s_dadda_rca32_and_24_25_y0);
  fa fa_h_s_dadda_rca32_fa636_y2(h_s_dadda_rca32_and_26_23_y0, h_s_dadda_rca32_and_25_24_y0, h_s_dadda_rca32_and_24_25_y0, h_s_dadda_rca32_fa636_y2, h_s_dadda_rca32_fa636_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_26_y0(a_23, b_26, h_s_dadda_rca32_and_23_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_27_y0(a_22, b_27, h_s_dadda_rca32_and_22_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_28_y0(a_21, b_28, h_s_dadda_rca32_and_21_28_y0);
  fa fa_h_s_dadda_rca32_fa637_y2(h_s_dadda_rca32_and_23_26_y0, h_s_dadda_rca32_and_22_27_y0, h_s_dadda_rca32_and_21_28_y0, h_s_dadda_rca32_fa637_y2, h_s_dadda_rca32_fa637_y4);
  and_gate and_gate_h_s_dadda_rca32_and_20_29_y0(a_20, b_29, h_s_dadda_rca32_and_20_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_19_30_y0(a_19, b_30, h_s_dadda_rca32_and_19_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_18_31_y0(a_18, b_31, h_s_dadda_rca32_nand_18_31_y0);
  fa fa_h_s_dadda_rca32_fa638_y2(h_s_dadda_rca32_and_20_29_y0, h_s_dadda_rca32_and_19_30_y0, h_s_dadda_rca32_nand_18_31_y0, h_s_dadda_rca32_fa638_y2, h_s_dadda_rca32_fa638_y4);
  fa fa_h_s_dadda_rca32_fa639_y2(h_s_dadda_rca32_fa631_y2, h_s_dadda_rca32_fa632_y2, h_s_dadda_rca32_fa633_y2, h_s_dadda_rca32_fa639_y2, h_s_dadda_rca32_fa639_y4);
  fa fa_h_s_dadda_rca32_fa640_y2(h_s_dadda_rca32_fa639_y4, h_s_dadda_rca32_fa638_y4, h_s_dadda_rca32_fa637_y4, h_s_dadda_rca32_fa640_y2, h_s_dadda_rca32_fa640_y4);
  fa fa_h_s_dadda_rca32_fa641_y2(h_s_dadda_rca32_fa636_y4, h_s_dadda_rca32_fa635_y4, h_s_dadda_rca32_fa634_y4, h_s_dadda_rca32_fa641_y2, h_s_dadda_rca32_fa641_y4);
  fa fa_h_s_dadda_rca32_fa642_y2(h_s_dadda_rca32_fa633_y4, h_s_dadda_rca32_fa632_y4, h_s_dadda_rca32_fa631_y4, h_s_dadda_rca32_fa642_y2, h_s_dadda_rca32_fa642_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_19_y0(a_31, b_19, h_s_dadda_rca32_nand_31_19_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_20_y0(a_30, b_20, h_s_dadda_rca32_and_30_20_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_21_y0(a_29, b_21, h_s_dadda_rca32_and_29_21_y0);
  fa fa_h_s_dadda_rca32_fa643_y2(h_s_dadda_rca32_nand_31_19_y0, h_s_dadda_rca32_and_30_20_y0, h_s_dadda_rca32_and_29_21_y0, h_s_dadda_rca32_fa643_y2, h_s_dadda_rca32_fa643_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_22_y0(a_28, b_22, h_s_dadda_rca32_and_28_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_23_y0(a_27, b_23, h_s_dadda_rca32_and_27_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_24_y0(a_26, b_24, h_s_dadda_rca32_and_26_24_y0);
  fa fa_h_s_dadda_rca32_fa644_y2(h_s_dadda_rca32_and_28_22_y0, h_s_dadda_rca32_and_27_23_y0, h_s_dadda_rca32_and_26_24_y0, h_s_dadda_rca32_fa644_y2, h_s_dadda_rca32_fa644_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_25_y0(a_25, b_25, h_s_dadda_rca32_and_25_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_26_y0(a_24, b_26, h_s_dadda_rca32_and_24_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_27_y0(a_23, b_27, h_s_dadda_rca32_and_23_27_y0);
  fa fa_h_s_dadda_rca32_fa645_y2(h_s_dadda_rca32_and_25_25_y0, h_s_dadda_rca32_and_24_26_y0, h_s_dadda_rca32_and_23_27_y0, h_s_dadda_rca32_fa645_y2, h_s_dadda_rca32_fa645_y4);
  and_gate and_gate_h_s_dadda_rca32_and_22_28_y0(a_22, b_28, h_s_dadda_rca32_and_22_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_21_29_y0(a_21, b_29, h_s_dadda_rca32_and_21_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_20_30_y0(a_20, b_30, h_s_dadda_rca32_and_20_30_y0);
  fa fa_h_s_dadda_rca32_fa646_y2(h_s_dadda_rca32_and_22_28_y0, h_s_dadda_rca32_and_21_29_y0, h_s_dadda_rca32_and_20_30_y0, h_s_dadda_rca32_fa646_y2, h_s_dadda_rca32_fa646_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_19_31_y0(a_19, b_31, h_s_dadda_rca32_nand_19_31_y0);
  fa fa_h_s_dadda_rca32_fa647_y2(h_s_dadda_rca32_nand_19_31_y0, h_s_dadda_rca32_fa640_y2, h_s_dadda_rca32_fa641_y2, h_s_dadda_rca32_fa647_y2, h_s_dadda_rca32_fa647_y4);
  fa fa_h_s_dadda_rca32_fa648_y2(h_s_dadda_rca32_fa647_y4, h_s_dadda_rca32_fa646_y4, h_s_dadda_rca32_fa645_y4, h_s_dadda_rca32_fa648_y2, h_s_dadda_rca32_fa648_y4);
  fa fa_h_s_dadda_rca32_fa649_y2(h_s_dadda_rca32_fa644_y4, h_s_dadda_rca32_fa643_y4, h_s_dadda_rca32_fa642_y4, h_s_dadda_rca32_fa649_y2, h_s_dadda_rca32_fa649_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_20_y0(a_31, b_20, h_s_dadda_rca32_nand_31_20_y0);
  fa fa_h_s_dadda_rca32_fa650_y2(h_s_dadda_rca32_fa641_y4, h_s_dadda_rca32_fa640_y4, h_s_dadda_rca32_nand_31_20_y0, h_s_dadda_rca32_fa650_y2, h_s_dadda_rca32_fa650_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_21_y0(a_30, b_21, h_s_dadda_rca32_and_30_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_22_y0(a_29, b_22, h_s_dadda_rca32_and_29_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_23_y0(a_28, b_23, h_s_dadda_rca32_and_28_23_y0);
  fa fa_h_s_dadda_rca32_fa651_y2(h_s_dadda_rca32_and_30_21_y0, h_s_dadda_rca32_and_29_22_y0, h_s_dadda_rca32_and_28_23_y0, h_s_dadda_rca32_fa651_y2, h_s_dadda_rca32_fa651_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_24_y0(a_27, b_24, h_s_dadda_rca32_and_27_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_25_y0(a_26, b_25, h_s_dadda_rca32_and_26_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_26_y0(a_25, b_26, h_s_dadda_rca32_and_25_26_y0);
  fa fa_h_s_dadda_rca32_fa652_y2(h_s_dadda_rca32_and_27_24_y0, h_s_dadda_rca32_and_26_25_y0, h_s_dadda_rca32_and_25_26_y0, h_s_dadda_rca32_fa652_y2, h_s_dadda_rca32_fa652_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_27_y0(a_24, b_27, h_s_dadda_rca32_and_24_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_28_y0(a_23, b_28, h_s_dadda_rca32_and_23_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_29_y0(a_22, b_29, h_s_dadda_rca32_and_22_29_y0);
  fa fa_h_s_dadda_rca32_fa653_y2(h_s_dadda_rca32_and_24_27_y0, h_s_dadda_rca32_and_23_28_y0, h_s_dadda_rca32_and_22_29_y0, h_s_dadda_rca32_fa653_y2, h_s_dadda_rca32_fa653_y4);
  and_gate and_gate_h_s_dadda_rca32_and_21_30_y0(a_21, b_30, h_s_dadda_rca32_and_21_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_20_31_y0(a_20, b_31, h_s_dadda_rca32_nand_20_31_y0);
  fa fa_h_s_dadda_rca32_fa654_y2(h_s_dadda_rca32_and_21_30_y0, h_s_dadda_rca32_nand_20_31_y0, h_s_dadda_rca32_fa648_y2, h_s_dadda_rca32_fa654_y2, h_s_dadda_rca32_fa654_y4);
  fa fa_h_s_dadda_rca32_fa655_y2(h_s_dadda_rca32_fa654_y4, h_s_dadda_rca32_fa653_y4, h_s_dadda_rca32_fa652_y4, h_s_dadda_rca32_fa655_y2, h_s_dadda_rca32_fa655_y4);
  fa fa_h_s_dadda_rca32_fa656_y2(h_s_dadda_rca32_fa651_y4, h_s_dadda_rca32_fa650_y4, h_s_dadda_rca32_fa649_y4, h_s_dadda_rca32_fa656_y2, h_s_dadda_rca32_fa656_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_21_y0(a_31, b_21, h_s_dadda_rca32_nand_31_21_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_22_y0(a_30, b_22, h_s_dadda_rca32_and_30_22_y0);
  fa fa_h_s_dadda_rca32_fa657_y2(h_s_dadda_rca32_fa648_y4, h_s_dadda_rca32_nand_31_21_y0, h_s_dadda_rca32_and_30_22_y0, h_s_dadda_rca32_fa657_y2, h_s_dadda_rca32_fa657_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_23_y0(a_29, b_23, h_s_dadda_rca32_and_29_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_24_y0(a_28, b_24, h_s_dadda_rca32_and_28_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_25_y0(a_27, b_25, h_s_dadda_rca32_and_27_25_y0);
  fa fa_h_s_dadda_rca32_fa658_y2(h_s_dadda_rca32_and_29_23_y0, h_s_dadda_rca32_and_28_24_y0, h_s_dadda_rca32_and_27_25_y0, h_s_dadda_rca32_fa658_y2, h_s_dadda_rca32_fa658_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_26_y0(a_26, b_26, h_s_dadda_rca32_and_26_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_27_y0(a_25, b_27, h_s_dadda_rca32_and_25_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_28_y0(a_24, b_28, h_s_dadda_rca32_and_24_28_y0);
  fa fa_h_s_dadda_rca32_fa659_y2(h_s_dadda_rca32_and_26_26_y0, h_s_dadda_rca32_and_25_27_y0, h_s_dadda_rca32_and_24_28_y0, h_s_dadda_rca32_fa659_y2, h_s_dadda_rca32_fa659_y4);
  and_gate and_gate_h_s_dadda_rca32_and_23_29_y0(a_23, b_29, h_s_dadda_rca32_and_23_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_22_30_y0(a_22, b_30, h_s_dadda_rca32_and_22_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_21_31_y0(a_21, b_31, h_s_dadda_rca32_nand_21_31_y0);
  fa fa_h_s_dadda_rca32_fa660_y2(h_s_dadda_rca32_and_23_29_y0, h_s_dadda_rca32_and_22_30_y0, h_s_dadda_rca32_nand_21_31_y0, h_s_dadda_rca32_fa660_y2, h_s_dadda_rca32_fa660_y4);
  fa fa_h_s_dadda_rca32_fa661_y2(h_s_dadda_rca32_fa660_y4, h_s_dadda_rca32_fa659_y4, h_s_dadda_rca32_fa658_y4, h_s_dadda_rca32_fa661_y2, h_s_dadda_rca32_fa661_y4);
  fa fa_h_s_dadda_rca32_fa662_y2(h_s_dadda_rca32_fa657_y4, h_s_dadda_rca32_fa656_y4, h_s_dadda_rca32_fa655_y4, h_s_dadda_rca32_fa662_y2, h_s_dadda_rca32_fa662_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_22_y0(a_31, b_22, h_s_dadda_rca32_nand_31_22_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_23_y0(a_30, b_23, h_s_dadda_rca32_and_30_23_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_24_y0(a_29, b_24, h_s_dadda_rca32_and_29_24_y0);
  fa fa_h_s_dadda_rca32_fa663_y2(h_s_dadda_rca32_nand_31_22_y0, h_s_dadda_rca32_and_30_23_y0, h_s_dadda_rca32_and_29_24_y0, h_s_dadda_rca32_fa663_y2, h_s_dadda_rca32_fa663_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_25_y0(a_28, b_25, h_s_dadda_rca32_and_28_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_26_y0(a_27, b_26, h_s_dadda_rca32_and_27_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_27_y0(a_26, b_27, h_s_dadda_rca32_and_26_27_y0);
  fa fa_h_s_dadda_rca32_fa664_y2(h_s_dadda_rca32_and_28_25_y0, h_s_dadda_rca32_and_27_26_y0, h_s_dadda_rca32_and_26_27_y0, h_s_dadda_rca32_fa664_y2, h_s_dadda_rca32_fa664_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_28_y0(a_25, b_28, h_s_dadda_rca32_and_25_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_24_29_y0(a_24, b_29, h_s_dadda_rca32_and_24_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_23_30_y0(a_23, b_30, h_s_dadda_rca32_and_23_30_y0);
  fa fa_h_s_dadda_rca32_fa665_y2(h_s_dadda_rca32_and_25_28_y0, h_s_dadda_rca32_and_24_29_y0, h_s_dadda_rca32_and_23_30_y0, h_s_dadda_rca32_fa665_y2, h_s_dadda_rca32_fa665_y4);
  fa fa_h_s_dadda_rca32_fa666_y2(h_s_dadda_rca32_fa665_y4, h_s_dadda_rca32_fa664_y4, h_s_dadda_rca32_fa663_y4, h_s_dadda_rca32_fa666_y2, h_s_dadda_rca32_fa666_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_23_y0(a_31, b_23, h_s_dadda_rca32_nand_31_23_y0);
  fa fa_h_s_dadda_rca32_fa667_y2(h_s_dadda_rca32_fa662_y4, h_s_dadda_rca32_fa661_y4, h_s_dadda_rca32_nand_31_23_y0, h_s_dadda_rca32_fa667_y2, h_s_dadda_rca32_fa667_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_24_y0(a_30, b_24, h_s_dadda_rca32_and_30_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_25_y0(a_29, b_25, h_s_dadda_rca32_and_29_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_26_y0(a_28, b_26, h_s_dadda_rca32_and_28_26_y0);
  fa fa_h_s_dadda_rca32_fa668_y2(h_s_dadda_rca32_and_30_24_y0, h_s_dadda_rca32_and_29_25_y0, h_s_dadda_rca32_and_28_26_y0, h_s_dadda_rca32_fa668_y2, h_s_dadda_rca32_fa668_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_27_y0(a_27, b_27, h_s_dadda_rca32_and_27_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_28_y0(a_26, b_28, h_s_dadda_rca32_and_26_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_25_29_y0(a_25, b_29, h_s_dadda_rca32_and_25_29_y0);
  fa fa_h_s_dadda_rca32_fa669_y2(h_s_dadda_rca32_and_27_27_y0, h_s_dadda_rca32_and_26_28_y0, h_s_dadda_rca32_and_25_29_y0, h_s_dadda_rca32_fa669_y2, h_s_dadda_rca32_fa669_y4);
  fa fa_h_s_dadda_rca32_fa670_y2(h_s_dadda_rca32_fa669_y4, h_s_dadda_rca32_fa668_y4, h_s_dadda_rca32_fa667_y4, h_s_dadda_rca32_fa670_y2, h_s_dadda_rca32_fa670_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_24_y0(a_31, b_24, h_s_dadda_rca32_nand_31_24_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_25_y0(a_30, b_25, h_s_dadda_rca32_and_30_25_y0);
  fa fa_h_s_dadda_rca32_fa671_y2(h_s_dadda_rca32_fa666_y4, h_s_dadda_rca32_nand_31_24_y0, h_s_dadda_rca32_and_30_25_y0, h_s_dadda_rca32_fa671_y2, h_s_dadda_rca32_fa671_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_26_y0(a_29, b_26, h_s_dadda_rca32_and_29_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_27_y0(a_28, b_27, h_s_dadda_rca32_and_28_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_28_y0(a_27, b_28, h_s_dadda_rca32_and_27_28_y0);
  fa fa_h_s_dadda_rca32_fa672_y2(h_s_dadda_rca32_and_29_26_y0, h_s_dadda_rca32_and_28_27_y0, h_s_dadda_rca32_and_27_28_y0, h_s_dadda_rca32_fa672_y2, h_s_dadda_rca32_fa672_y4);
  fa fa_h_s_dadda_rca32_fa673_y2(h_s_dadda_rca32_fa672_y4, h_s_dadda_rca32_fa671_y4, h_s_dadda_rca32_fa670_y4, h_s_dadda_rca32_fa673_y2, h_s_dadda_rca32_fa673_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_25_y0(a_31, b_25, h_s_dadda_rca32_nand_31_25_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_26_y0(a_30, b_26, h_s_dadda_rca32_and_30_26_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_27_y0(a_29, b_27, h_s_dadda_rca32_and_29_27_y0);
  fa fa_h_s_dadda_rca32_fa674_y2(h_s_dadda_rca32_nand_31_25_y0, h_s_dadda_rca32_and_30_26_y0, h_s_dadda_rca32_and_29_27_y0, h_s_dadda_rca32_fa674_y2, h_s_dadda_rca32_fa674_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_26_y0(a_31, b_26, h_s_dadda_rca32_nand_31_26_y0);
  fa fa_h_s_dadda_rca32_fa675_y2(h_s_dadda_rca32_fa674_y4, h_s_dadda_rca32_fa673_y4, h_s_dadda_rca32_nand_31_26_y0, h_s_dadda_rca32_fa675_y2, h_s_dadda_rca32_fa675_y4);
  and_gate and_gate_h_s_dadda_rca32_and_4_0_y0(a_4, b_0, h_s_dadda_rca32_and_4_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_3_1_y0(a_3, b_1, h_s_dadda_rca32_and_3_1_y0);
  ha ha_h_s_dadda_rca32_ha26_y0(h_s_dadda_rca32_and_4_0_y0, h_s_dadda_rca32_and_3_1_y0, h_s_dadda_rca32_ha26_y0, h_s_dadda_rca32_ha26_y1);
  and_gate and_gate_h_s_dadda_rca32_and_5_0_y0(a_5, b_0, h_s_dadda_rca32_and_5_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_4_1_y0(a_4, b_1, h_s_dadda_rca32_and_4_1_y0);
  fa fa_h_s_dadda_rca32_fa676_y2(h_s_dadda_rca32_ha26_y1, h_s_dadda_rca32_and_5_0_y0, h_s_dadda_rca32_and_4_1_y0, h_s_dadda_rca32_fa676_y2, h_s_dadda_rca32_fa676_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_2_y0(a_3, b_2, h_s_dadda_rca32_and_3_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_3_y0(a_2, b_3, h_s_dadda_rca32_and_2_3_y0);
  ha ha_h_s_dadda_rca32_ha27_y0(h_s_dadda_rca32_and_3_2_y0, h_s_dadda_rca32_and_2_3_y0, h_s_dadda_rca32_ha27_y0, h_s_dadda_rca32_ha27_y1);
  and_gate and_gate_h_s_dadda_rca32_and_4_2_y0(a_4, b_2, h_s_dadda_rca32_and_4_2_y0);
  fa fa_h_s_dadda_rca32_fa677_y2(h_s_dadda_rca32_ha27_y1, h_s_dadda_rca32_fa676_y4, h_s_dadda_rca32_and_4_2_y0, h_s_dadda_rca32_fa677_y2, h_s_dadda_rca32_fa677_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_3_y0(a_3, b_3, h_s_dadda_rca32_and_3_3_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_4_y0(a_2, b_4, h_s_dadda_rca32_and_2_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_5_y0(a_1, b_5, h_s_dadda_rca32_and_1_5_y0);
  fa fa_h_s_dadda_rca32_fa678_y2(h_s_dadda_rca32_and_3_3_y0, h_s_dadda_rca32_and_2_4_y0, h_s_dadda_rca32_and_1_5_y0, h_s_dadda_rca32_fa678_y2, h_s_dadda_rca32_fa678_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_4_y0(a_3, b_4, h_s_dadda_rca32_and_3_4_y0);
  fa fa_h_s_dadda_rca32_fa679_y2(h_s_dadda_rca32_fa678_y4, h_s_dadda_rca32_fa677_y4, h_s_dadda_rca32_and_3_4_y0, h_s_dadda_rca32_fa679_y2, h_s_dadda_rca32_fa679_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_5_y0(a_2, b_5, h_s_dadda_rca32_and_2_5_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_6_y0(a_1, b_6, h_s_dadda_rca32_and_1_6_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_7_y0(a_0, b_7, h_s_dadda_rca32_and_0_7_y0);
  fa fa_h_s_dadda_rca32_fa680_y2(h_s_dadda_rca32_and_2_5_y0, h_s_dadda_rca32_and_1_6_y0, h_s_dadda_rca32_and_0_7_y0, h_s_dadda_rca32_fa680_y2, h_s_dadda_rca32_fa680_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_6_y0(a_2, b_6, h_s_dadda_rca32_and_2_6_y0);
  fa fa_h_s_dadda_rca32_fa681_y2(h_s_dadda_rca32_fa680_y4, h_s_dadda_rca32_fa679_y4, h_s_dadda_rca32_and_2_6_y0, h_s_dadda_rca32_fa681_y2, h_s_dadda_rca32_fa681_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_7_y0(a_1, b_7, h_s_dadda_rca32_and_1_7_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_8_y0(a_0, b_8, h_s_dadda_rca32_and_0_8_y0);
  fa fa_h_s_dadda_rca32_fa682_y2(h_s_dadda_rca32_and_1_7_y0, h_s_dadda_rca32_and_0_8_y0, h_s_dadda_rca32_fa17_y2, h_s_dadda_rca32_fa682_y2, h_s_dadda_rca32_fa682_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_8_y0(a_1, b_8, h_s_dadda_rca32_and_1_8_y0);
  fa fa_h_s_dadda_rca32_fa683_y2(h_s_dadda_rca32_fa682_y4, h_s_dadda_rca32_fa681_y4, h_s_dadda_rca32_and_1_8_y0, h_s_dadda_rca32_fa683_y2, h_s_dadda_rca32_fa683_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_9_y0(a_0, b_9, h_s_dadda_rca32_and_0_9_y0);
  fa fa_h_s_dadda_rca32_fa684_y2(h_s_dadda_rca32_and_0_9_y0, h_s_dadda_rca32_fa19_y2, h_s_dadda_rca32_fa20_y2, h_s_dadda_rca32_fa684_y2, h_s_dadda_rca32_fa684_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_10_y0(a_0, b_10, h_s_dadda_rca32_and_0_10_y0);
  fa fa_h_s_dadda_rca32_fa685_y2(h_s_dadda_rca32_fa684_y4, h_s_dadda_rca32_fa683_y4, h_s_dadda_rca32_and_0_10_y0, h_s_dadda_rca32_fa685_y2, h_s_dadda_rca32_fa685_y4);
  fa fa_h_s_dadda_rca32_fa686_y2(h_s_dadda_rca32_fa22_y2, h_s_dadda_rca32_fa23_y2, h_s_dadda_rca32_fa24_y2, h_s_dadda_rca32_fa686_y2, h_s_dadda_rca32_fa686_y4);
  fa fa_h_s_dadda_rca32_fa687_y2(h_s_dadda_rca32_fa686_y4, h_s_dadda_rca32_fa685_y4, h_s_dadda_rca32_fa26_y2, h_s_dadda_rca32_fa687_y2, h_s_dadda_rca32_fa687_y4);
  fa fa_h_s_dadda_rca32_fa688_y2(h_s_dadda_rca32_fa27_y2, h_s_dadda_rca32_fa28_y2, h_s_dadda_rca32_fa29_y2, h_s_dadda_rca32_fa688_y2, h_s_dadda_rca32_fa688_y4);
  fa fa_h_s_dadda_rca32_fa689_y2(h_s_dadda_rca32_fa688_y4, h_s_dadda_rca32_fa687_y4, h_s_dadda_rca32_fa32_y2, h_s_dadda_rca32_fa689_y2, h_s_dadda_rca32_fa689_y4);
  fa fa_h_s_dadda_rca32_fa690_y2(h_s_dadda_rca32_fa33_y2, h_s_dadda_rca32_fa34_y2, h_s_dadda_rca32_fa35_y2, h_s_dadda_rca32_fa690_y2, h_s_dadda_rca32_fa690_y4);
  fa fa_h_s_dadda_rca32_fa691_y2(h_s_dadda_rca32_fa690_y4, h_s_dadda_rca32_fa689_y4, h_s_dadda_rca32_fa39_y2, h_s_dadda_rca32_fa691_y2, h_s_dadda_rca32_fa691_y4);
  fa fa_h_s_dadda_rca32_fa692_y2(h_s_dadda_rca32_fa40_y2, h_s_dadda_rca32_fa41_y2, h_s_dadda_rca32_fa42_y2, h_s_dadda_rca32_fa692_y2, h_s_dadda_rca32_fa692_y4);
  fa fa_h_s_dadda_rca32_fa693_y2(h_s_dadda_rca32_fa692_y4, h_s_dadda_rca32_fa691_y4, h_s_dadda_rca32_fa47_y2, h_s_dadda_rca32_fa693_y2, h_s_dadda_rca32_fa693_y4);
  fa fa_h_s_dadda_rca32_fa694_y2(h_s_dadda_rca32_fa48_y2, h_s_dadda_rca32_fa49_y2, h_s_dadda_rca32_fa50_y2, h_s_dadda_rca32_fa694_y2, h_s_dadda_rca32_fa694_y4);
  fa fa_h_s_dadda_rca32_fa695_y2(h_s_dadda_rca32_fa694_y4, h_s_dadda_rca32_fa693_y4, h_s_dadda_rca32_fa56_y2, h_s_dadda_rca32_fa695_y2, h_s_dadda_rca32_fa695_y4);
  fa fa_h_s_dadda_rca32_fa696_y2(h_s_dadda_rca32_fa57_y2, h_s_dadda_rca32_fa58_y2, h_s_dadda_rca32_fa59_y2, h_s_dadda_rca32_fa696_y2, h_s_dadda_rca32_fa696_y4);
  fa fa_h_s_dadda_rca32_fa697_y2(h_s_dadda_rca32_fa696_y4, h_s_dadda_rca32_fa695_y4, h_s_dadda_rca32_fa66_y2, h_s_dadda_rca32_fa697_y2, h_s_dadda_rca32_fa697_y4);
  fa fa_h_s_dadda_rca32_fa698_y2(h_s_dadda_rca32_fa67_y2, h_s_dadda_rca32_fa68_y2, h_s_dadda_rca32_fa69_y2, h_s_dadda_rca32_fa698_y2, h_s_dadda_rca32_fa698_y4);
  fa fa_h_s_dadda_rca32_fa699_y2(h_s_dadda_rca32_fa698_y4, h_s_dadda_rca32_fa697_y4, h_s_dadda_rca32_fa77_y2, h_s_dadda_rca32_fa699_y2, h_s_dadda_rca32_fa699_y4);
  fa fa_h_s_dadda_rca32_fa700_y2(h_s_dadda_rca32_fa78_y2, h_s_dadda_rca32_fa79_y2, h_s_dadda_rca32_fa80_y2, h_s_dadda_rca32_fa700_y2, h_s_dadda_rca32_fa700_y4);
  fa fa_h_s_dadda_rca32_fa701_y2(h_s_dadda_rca32_fa700_y4, h_s_dadda_rca32_fa699_y4, h_s_dadda_rca32_fa89_y2, h_s_dadda_rca32_fa701_y2, h_s_dadda_rca32_fa701_y4);
  fa fa_h_s_dadda_rca32_fa702_y2(h_s_dadda_rca32_fa90_y2, h_s_dadda_rca32_fa91_y2, h_s_dadda_rca32_fa92_y2, h_s_dadda_rca32_fa702_y2, h_s_dadda_rca32_fa702_y4);
  fa fa_h_s_dadda_rca32_fa703_y2(h_s_dadda_rca32_fa702_y4, h_s_dadda_rca32_fa701_y4, h_s_dadda_rca32_fa102_y2, h_s_dadda_rca32_fa703_y2, h_s_dadda_rca32_fa703_y4);
  fa fa_h_s_dadda_rca32_fa704_y2(h_s_dadda_rca32_fa103_y2, h_s_dadda_rca32_fa104_y2, h_s_dadda_rca32_fa105_y2, h_s_dadda_rca32_fa704_y2, h_s_dadda_rca32_fa704_y4);
  fa fa_h_s_dadda_rca32_fa705_y2(h_s_dadda_rca32_fa704_y4, h_s_dadda_rca32_fa703_y4, h_s_dadda_rca32_fa116_y2, h_s_dadda_rca32_fa705_y2, h_s_dadda_rca32_fa705_y4);
  fa fa_h_s_dadda_rca32_fa706_y2(h_s_dadda_rca32_fa117_y2, h_s_dadda_rca32_fa118_y2, h_s_dadda_rca32_fa119_y2, h_s_dadda_rca32_fa706_y2, h_s_dadda_rca32_fa706_y4);
  fa fa_h_s_dadda_rca32_fa707_y2(h_s_dadda_rca32_fa706_y4, h_s_dadda_rca32_fa705_y4, h_s_dadda_rca32_fa131_y2, h_s_dadda_rca32_fa707_y2, h_s_dadda_rca32_fa707_y4);
  fa fa_h_s_dadda_rca32_fa708_y2(h_s_dadda_rca32_fa132_y2, h_s_dadda_rca32_fa133_y2, h_s_dadda_rca32_fa134_y2, h_s_dadda_rca32_fa708_y2, h_s_dadda_rca32_fa708_y4);
  fa fa_h_s_dadda_rca32_fa709_y2(h_s_dadda_rca32_fa708_y4, h_s_dadda_rca32_fa707_y4, h_s_dadda_rca32_fa147_y2, h_s_dadda_rca32_fa709_y2, h_s_dadda_rca32_fa709_y4);
  fa fa_h_s_dadda_rca32_fa710_y2(h_s_dadda_rca32_fa148_y2, h_s_dadda_rca32_fa149_y2, h_s_dadda_rca32_fa150_y2, h_s_dadda_rca32_fa710_y2, h_s_dadda_rca32_fa710_y4);
  fa fa_h_s_dadda_rca32_fa711_y2(h_s_dadda_rca32_fa710_y4, h_s_dadda_rca32_fa709_y4, h_s_dadda_rca32_fa164_y2, h_s_dadda_rca32_fa711_y2, h_s_dadda_rca32_fa711_y4);
  fa fa_h_s_dadda_rca32_fa712_y2(h_s_dadda_rca32_fa165_y2, h_s_dadda_rca32_fa166_y2, h_s_dadda_rca32_fa167_y2, h_s_dadda_rca32_fa712_y2, h_s_dadda_rca32_fa712_y4);
  fa fa_h_s_dadda_rca32_fa713_y2(h_s_dadda_rca32_fa712_y4, h_s_dadda_rca32_fa711_y4, h_s_dadda_rca32_fa182_y2, h_s_dadda_rca32_fa713_y2, h_s_dadda_rca32_fa713_y4);
  fa fa_h_s_dadda_rca32_fa714_y2(h_s_dadda_rca32_fa183_y2, h_s_dadda_rca32_fa184_y2, h_s_dadda_rca32_fa185_y2, h_s_dadda_rca32_fa714_y2, h_s_dadda_rca32_fa714_y4);
  fa fa_h_s_dadda_rca32_fa715_y2(h_s_dadda_rca32_fa714_y4, h_s_dadda_rca32_fa713_y4, h_s_dadda_rca32_fa201_y2, h_s_dadda_rca32_fa715_y2, h_s_dadda_rca32_fa715_y4);
  fa fa_h_s_dadda_rca32_fa716_y2(h_s_dadda_rca32_fa202_y2, h_s_dadda_rca32_fa203_y2, h_s_dadda_rca32_fa204_y2, h_s_dadda_rca32_fa716_y2, h_s_dadda_rca32_fa716_y4);
  fa fa_h_s_dadda_rca32_fa717_y2(h_s_dadda_rca32_fa716_y4, h_s_dadda_rca32_fa715_y4, h_s_dadda_rca32_fa221_y2, h_s_dadda_rca32_fa717_y2, h_s_dadda_rca32_fa717_y4);
  fa fa_h_s_dadda_rca32_fa718_y2(h_s_dadda_rca32_fa222_y2, h_s_dadda_rca32_fa223_y2, h_s_dadda_rca32_fa224_y2, h_s_dadda_rca32_fa718_y2, h_s_dadda_rca32_fa718_y4);
  fa fa_h_s_dadda_rca32_fa719_y2(h_s_dadda_rca32_fa718_y4, h_s_dadda_rca32_fa717_y4, h_s_dadda_rca32_fa242_y2, h_s_dadda_rca32_fa719_y2, h_s_dadda_rca32_fa719_y4);
  fa fa_h_s_dadda_rca32_fa720_y2(h_s_dadda_rca32_fa243_y2, h_s_dadda_rca32_fa244_y2, h_s_dadda_rca32_fa245_y2, h_s_dadda_rca32_fa720_y2, h_s_dadda_rca32_fa720_y4);
  fa fa_h_s_dadda_rca32_fa721_y2(h_s_dadda_rca32_fa720_y4, h_s_dadda_rca32_fa719_y4, h_s_dadda_rca32_fa263_y2, h_s_dadda_rca32_fa721_y2, h_s_dadda_rca32_fa721_y4);
  fa fa_h_s_dadda_rca32_fa722_y2(h_s_dadda_rca32_fa264_y2, h_s_dadda_rca32_fa265_y2, h_s_dadda_rca32_fa266_y2, h_s_dadda_rca32_fa722_y2, h_s_dadda_rca32_fa722_y4);
  fa fa_h_s_dadda_rca32_fa723_y2(h_s_dadda_rca32_fa722_y4, h_s_dadda_rca32_fa721_y4, h_s_dadda_rca32_fa285_y2, h_s_dadda_rca32_fa723_y2, h_s_dadda_rca32_fa723_y4);
  fa fa_h_s_dadda_rca32_fa724_y2(h_s_dadda_rca32_fa286_y2, h_s_dadda_rca32_fa287_y2, h_s_dadda_rca32_fa288_y2, h_s_dadda_rca32_fa724_y2, h_s_dadda_rca32_fa724_y4);
  fa fa_h_s_dadda_rca32_fa725_y2(h_s_dadda_rca32_fa724_y4, h_s_dadda_rca32_fa723_y4, h_s_dadda_rca32_fa307_y2, h_s_dadda_rca32_fa725_y2, h_s_dadda_rca32_fa725_y4);
  fa fa_h_s_dadda_rca32_fa726_y2(h_s_dadda_rca32_fa308_y2, h_s_dadda_rca32_fa309_y2, h_s_dadda_rca32_fa310_y2, h_s_dadda_rca32_fa726_y2, h_s_dadda_rca32_fa726_y4);
  fa fa_h_s_dadda_rca32_fa727_y2(h_s_dadda_rca32_fa726_y4, h_s_dadda_rca32_fa725_y4, h_s_dadda_rca32_fa329_y2, h_s_dadda_rca32_fa727_y2, h_s_dadda_rca32_fa727_y4);
  fa fa_h_s_dadda_rca32_fa728_y2(h_s_dadda_rca32_fa330_y2, h_s_dadda_rca32_fa331_y2, h_s_dadda_rca32_fa332_y2, h_s_dadda_rca32_fa728_y2, h_s_dadda_rca32_fa728_y4);
  fa fa_h_s_dadda_rca32_fa729_y2(h_s_dadda_rca32_fa728_y4, h_s_dadda_rca32_fa727_y4, h_s_dadda_rca32_fa351_y2, h_s_dadda_rca32_fa729_y2, h_s_dadda_rca32_fa729_y4);
  fa fa_h_s_dadda_rca32_fa730_y2(h_s_dadda_rca32_fa352_y2, h_s_dadda_rca32_fa353_y2, h_s_dadda_rca32_fa354_y2, h_s_dadda_rca32_fa730_y2, h_s_dadda_rca32_fa730_y4);
  fa fa_h_s_dadda_rca32_fa731_y2(h_s_dadda_rca32_fa730_y4, h_s_dadda_rca32_fa729_y4, h_s_dadda_rca32_fa373_y2, h_s_dadda_rca32_fa731_y2, h_s_dadda_rca32_fa731_y4);
  fa fa_h_s_dadda_rca32_fa732_y2(h_s_dadda_rca32_fa374_y2, h_s_dadda_rca32_fa375_y2, h_s_dadda_rca32_fa376_y2, h_s_dadda_rca32_fa732_y2, h_s_dadda_rca32_fa732_y4);
  fa fa_h_s_dadda_rca32_fa733_y2(h_s_dadda_rca32_fa732_y4, h_s_dadda_rca32_fa731_y4, h_s_dadda_rca32_fa395_y2, h_s_dadda_rca32_fa733_y2, h_s_dadda_rca32_fa733_y4);
  fa fa_h_s_dadda_rca32_fa734_y2(h_s_dadda_rca32_fa396_y2, h_s_dadda_rca32_fa397_y2, h_s_dadda_rca32_fa398_y2, h_s_dadda_rca32_fa734_y2, h_s_dadda_rca32_fa734_y4);
  fa fa_h_s_dadda_rca32_fa735_y2(h_s_dadda_rca32_fa734_y4, h_s_dadda_rca32_fa733_y4, h_s_dadda_rca32_fa417_y2, h_s_dadda_rca32_fa735_y2, h_s_dadda_rca32_fa735_y4);
  fa fa_h_s_dadda_rca32_fa736_y2(h_s_dadda_rca32_fa418_y2, h_s_dadda_rca32_fa419_y2, h_s_dadda_rca32_fa420_y2, h_s_dadda_rca32_fa736_y2, h_s_dadda_rca32_fa736_y4);
  fa fa_h_s_dadda_rca32_fa737_y2(h_s_dadda_rca32_fa736_y4, h_s_dadda_rca32_fa735_y4, h_s_dadda_rca32_fa439_y2, h_s_dadda_rca32_fa737_y2, h_s_dadda_rca32_fa737_y4);
  fa fa_h_s_dadda_rca32_fa738_y2(h_s_dadda_rca32_fa440_y2, h_s_dadda_rca32_fa441_y2, h_s_dadda_rca32_fa442_y2, h_s_dadda_rca32_fa738_y2, h_s_dadda_rca32_fa738_y4);
  fa fa_h_s_dadda_rca32_fa739_y2(h_s_dadda_rca32_fa738_y4, h_s_dadda_rca32_fa737_y4, h_s_dadda_rca32_fa460_y2, h_s_dadda_rca32_fa739_y2, h_s_dadda_rca32_fa739_y4);
  fa fa_h_s_dadda_rca32_fa740_y2(h_s_dadda_rca32_fa461_y2, h_s_dadda_rca32_fa462_y2, h_s_dadda_rca32_fa463_y2, h_s_dadda_rca32_fa740_y2, h_s_dadda_rca32_fa740_y4);
  fa fa_h_s_dadda_rca32_fa741_y2(h_s_dadda_rca32_fa740_y4, h_s_dadda_rca32_fa739_y4, h_s_dadda_rca32_fa480_y2, h_s_dadda_rca32_fa741_y2, h_s_dadda_rca32_fa741_y4);
  fa fa_h_s_dadda_rca32_fa742_y2(h_s_dadda_rca32_fa481_y2, h_s_dadda_rca32_fa482_y2, h_s_dadda_rca32_fa483_y2, h_s_dadda_rca32_fa742_y2, h_s_dadda_rca32_fa742_y4);
  fa fa_h_s_dadda_rca32_fa743_y2(h_s_dadda_rca32_fa742_y4, h_s_dadda_rca32_fa741_y4, h_s_dadda_rca32_fa499_y2, h_s_dadda_rca32_fa743_y2, h_s_dadda_rca32_fa743_y4);
  fa fa_h_s_dadda_rca32_fa744_y2(h_s_dadda_rca32_fa500_y2, h_s_dadda_rca32_fa501_y2, h_s_dadda_rca32_fa502_y2, h_s_dadda_rca32_fa744_y2, h_s_dadda_rca32_fa744_y4);
  fa fa_h_s_dadda_rca32_fa745_y2(h_s_dadda_rca32_fa744_y4, h_s_dadda_rca32_fa743_y4, h_s_dadda_rca32_fa517_y2, h_s_dadda_rca32_fa745_y2, h_s_dadda_rca32_fa745_y4);
  fa fa_h_s_dadda_rca32_fa746_y2(h_s_dadda_rca32_fa518_y2, h_s_dadda_rca32_fa519_y2, h_s_dadda_rca32_fa520_y2, h_s_dadda_rca32_fa746_y2, h_s_dadda_rca32_fa746_y4);
  fa fa_h_s_dadda_rca32_fa747_y2(h_s_dadda_rca32_fa746_y4, h_s_dadda_rca32_fa745_y4, h_s_dadda_rca32_fa534_y2, h_s_dadda_rca32_fa747_y2, h_s_dadda_rca32_fa747_y4);
  fa fa_h_s_dadda_rca32_fa748_y2(h_s_dadda_rca32_fa535_y2, h_s_dadda_rca32_fa536_y2, h_s_dadda_rca32_fa537_y2, h_s_dadda_rca32_fa748_y2, h_s_dadda_rca32_fa748_y4);
  fa fa_h_s_dadda_rca32_fa749_y2(h_s_dadda_rca32_fa748_y4, h_s_dadda_rca32_fa747_y4, h_s_dadda_rca32_fa550_y2, h_s_dadda_rca32_fa749_y2, h_s_dadda_rca32_fa749_y4);
  fa fa_h_s_dadda_rca32_fa750_y2(h_s_dadda_rca32_fa551_y2, h_s_dadda_rca32_fa552_y2, h_s_dadda_rca32_fa553_y2, h_s_dadda_rca32_fa750_y2, h_s_dadda_rca32_fa750_y4);
  fa fa_h_s_dadda_rca32_fa751_y2(h_s_dadda_rca32_fa750_y4, h_s_dadda_rca32_fa749_y4, h_s_dadda_rca32_fa565_y2, h_s_dadda_rca32_fa751_y2, h_s_dadda_rca32_fa751_y4);
  fa fa_h_s_dadda_rca32_fa752_y2(h_s_dadda_rca32_fa566_y2, h_s_dadda_rca32_fa567_y2, h_s_dadda_rca32_fa568_y2, h_s_dadda_rca32_fa752_y2, h_s_dadda_rca32_fa752_y4);
  fa fa_h_s_dadda_rca32_fa753_y2(h_s_dadda_rca32_fa752_y4, h_s_dadda_rca32_fa751_y4, h_s_dadda_rca32_fa579_y2, h_s_dadda_rca32_fa753_y2, h_s_dadda_rca32_fa753_y4);
  fa fa_h_s_dadda_rca32_fa754_y2(h_s_dadda_rca32_fa580_y2, h_s_dadda_rca32_fa581_y2, h_s_dadda_rca32_fa582_y2, h_s_dadda_rca32_fa754_y2, h_s_dadda_rca32_fa754_y4);
  fa fa_h_s_dadda_rca32_fa755_y2(h_s_dadda_rca32_fa754_y4, h_s_dadda_rca32_fa753_y4, h_s_dadda_rca32_fa592_y2, h_s_dadda_rca32_fa755_y2, h_s_dadda_rca32_fa755_y4);
  fa fa_h_s_dadda_rca32_fa756_y2(h_s_dadda_rca32_fa593_y2, h_s_dadda_rca32_fa594_y2, h_s_dadda_rca32_fa595_y2, h_s_dadda_rca32_fa756_y2, h_s_dadda_rca32_fa756_y4);
  fa fa_h_s_dadda_rca32_fa757_y2(h_s_dadda_rca32_fa756_y4, h_s_dadda_rca32_fa755_y4, h_s_dadda_rca32_fa604_y2, h_s_dadda_rca32_fa757_y2, h_s_dadda_rca32_fa757_y4);
  fa fa_h_s_dadda_rca32_fa758_y2(h_s_dadda_rca32_fa605_y2, h_s_dadda_rca32_fa606_y2, h_s_dadda_rca32_fa607_y2, h_s_dadda_rca32_fa758_y2, h_s_dadda_rca32_fa758_y4);
  fa fa_h_s_dadda_rca32_fa759_y2(h_s_dadda_rca32_fa758_y4, h_s_dadda_rca32_fa757_y4, h_s_dadda_rca32_fa615_y2, h_s_dadda_rca32_fa759_y2, h_s_dadda_rca32_fa759_y4);
  fa fa_h_s_dadda_rca32_fa760_y2(h_s_dadda_rca32_fa616_y2, h_s_dadda_rca32_fa617_y2, h_s_dadda_rca32_fa618_y2, h_s_dadda_rca32_fa760_y2, h_s_dadda_rca32_fa760_y4);
  fa fa_h_s_dadda_rca32_fa761_y2(h_s_dadda_rca32_fa760_y4, h_s_dadda_rca32_fa759_y4, h_s_dadda_rca32_fa625_y2, h_s_dadda_rca32_fa761_y2, h_s_dadda_rca32_fa761_y4);
  fa fa_h_s_dadda_rca32_fa762_y2(h_s_dadda_rca32_fa626_y2, h_s_dadda_rca32_fa627_y2, h_s_dadda_rca32_fa628_y2, h_s_dadda_rca32_fa762_y2, h_s_dadda_rca32_fa762_y4);
  fa fa_h_s_dadda_rca32_fa763_y2(h_s_dadda_rca32_fa762_y4, h_s_dadda_rca32_fa761_y4, h_s_dadda_rca32_fa634_y2, h_s_dadda_rca32_fa763_y2, h_s_dadda_rca32_fa763_y4);
  fa fa_h_s_dadda_rca32_fa764_y2(h_s_dadda_rca32_fa635_y2, h_s_dadda_rca32_fa636_y2, h_s_dadda_rca32_fa637_y2, h_s_dadda_rca32_fa764_y2, h_s_dadda_rca32_fa764_y4);
  fa fa_h_s_dadda_rca32_fa765_y2(h_s_dadda_rca32_fa764_y4, h_s_dadda_rca32_fa763_y4, h_s_dadda_rca32_fa642_y2, h_s_dadda_rca32_fa765_y2, h_s_dadda_rca32_fa765_y4);
  fa fa_h_s_dadda_rca32_fa766_y2(h_s_dadda_rca32_fa643_y2, h_s_dadda_rca32_fa644_y2, h_s_dadda_rca32_fa645_y2, h_s_dadda_rca32_fa766_y2, h_s_dadda_rca32_fa766_y4);
  fa fa_h_s_dadda_rca32_fa767_y2(h_s_dadda_rca32_fa766_y4, h_s_dadda_rca32_fa765_y4, h_s_dadda_rca32_fa649_y2, h_s_dadda_rca32_fa767_y2, h_s_dadda_rca32_fa767_y4);
  fa fa_h_s_dadda_rca32_fa768_y2(h_s_dadda_rca32_fa650_y2, h_s_dadda_rca32_fa651_y2, h_s_dadda_rca32_fa652_y2, h_s_dadda_rca32_fa768_y2, h_s_dadda_rca32_fa768_y4);
  fa fa_h_s_dadda_rca32_fa769_y2(h_s_dadda_rca32_fa768_y4, h_s_dadda_rca32_fa767_y4, h_s_dadda_rca32_fa655_y2, h_s_dadda_rca32_fa769_y2, h_s_dadda_rca32_fa769_y4);
  fa fa_h_s_dadda_rca32_fa770_y2(h_s_dadda_rca32_fa656_y2, h_s_dadda_rca32_fa657_y2, h_s_dadda_rca32_fa658_y2, h_s_dadda_rca32_fa770_y2, h_s_dadda_rca32_fa770_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_22_31_y0(a_22, b_31, h_s_dadda_rca32_nand_22_31_y0);
  fa fa_h_s_dadda_rca32_fa771_y2(h_s_dadda_rca32_fa770_y4, h_s_dadda_rca32_fa769_y4, h_s_dadda_rca32_nand_22_31_y0, h_s_dadda_rca32_fa771_y2, h_s_dadda_rca32_fa771_y4);
  fa fa_h_s_dadda_rca32_fa772_y2(h_s_dadda_rca32_fa661_y2, h_s_dadda_rca32_fa662_y2, h_s_dadda_rca32_fa663_y2, h_s_dadda_rca32_fa772_y2, h_s_dadda_rca32_fa772_y4);
  and_gate and_gate_h_s_dadda_rca32_and_24_30_y0(a_24, b_30, h_s_dadda_rca32_and_24_30_y0);
  fa fa_h_s_dadda_rca32_fa773_y2(h_s_dadda_rca32_fa772_y4, h_s_dadda_rca32_fa771_y4, h_s_dadda_rca32_and_24_30_y0, h_s_dadda_rca32_fa773_y2, h_s_dadda_rca32_fa773_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_23_31_y0(a_23, b_31, h_s_dadda_rca32_nand_23_31_y0);
  fa fa_h_s_dadda_rca32_fa774_y2(h_s_dadda_rca32_nand_23_31_y0, h_s_dadda_rca32_fa666_y2, h_s_dadda_rca32_fa667_y2, h_s_dadda_rca32_fa774_y2, h_s_dadda_rca32_fa774_y4);
  and_gate and_gate_h_s_dadda_rca32_and_26_29_y0(a_26, b_29, h_s_dadda_rca32_and_26_29_y0);
  fa fa_h_s_dadda_rca32_fa775_y2(h_s_dadda_rca32_fa774_y4, h_s_dadda_rca32_fa773_y4, h_s_dadda_rca32_and_26_29_y0, h_s_dadda_rca32_fa775_y2, h_s_dadda_rca32_fa775_y4);
  and_gate and_gate_h_s_dadda_rca32_and_25_30_y0(a_25, b_30, h_s_dadda_rca32_and_25_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_24_31_y0(a_24, b_31, h_s_dadda_rca32_nand_24_31_y0);
  fa fa_h_s_dadda_rca32_fa776_y2(h_s_dadda_rca32_and_25_30_y0, h_s_dadda_rca32_nand_24_31_y0, h_s_dadda_rca32_fa670_y2, h_s_dadda_rca32_fa776_y2, h_s_dadda_rca32_fa776_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_28_y0(a_28, b_28, h_s_dadda_rca32_and_28_28_y0);
  fa fa_h_s_dadda_rca32_fa777_y2(h_s_dadda_rca32_fa776_y4, h_s_dadda_rca32_fa775_y4, h_s_dadda_rca32_and_28_28_y0, h_s_dadda_rca32_fa777_y2, h_s_dadda_rca32_fa777_y4);
  and_gate and_gate_h_s_dadda_rca32_and_27_29_y0(a_27, b_29, h_s_dadda_rca32_and_27_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_26_30_y0(a_26, b_30, h_s_dadda_rca32_and_26_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_25_31_y0(a_25, b_31, h_s_dadda_rca32_nand_25_31_y0);
  fa fa_h_s_dadda_rca32_fa778_y2(h_s_dadda_rca32_and_27_29_y0, h_s_dadda_rca32_and_26_30_y0, h_s_dadda_rca32_nand_25_31_y0, h_s_dadda_rca32_fa778_y2, h_s_dadda_rca32_fa778_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_27_y0(a_30, b_27, h_s_dadda_rca32_and_30_27_y0);
  fa fa_h_s_dadda_rca32_fa779_y2(h_s_dadda_rca32_fa778_y4, h_s_dadda_rca32_fa777_y4, h_s_dadda_rca32_and_30_27_y0, h_s_dadda_rca32_fa779_y2, h_s_dadda_rca32_fa779_y4);
  and_gate and_gate_h_s_dadda_rca32_and_29_28_y0(a_29, b_28, h_s_dadda_rca32_and_29_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_28_29_y0(a_28, b_29, h_s_dadda_rca32_and_28_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_27_30_y0(a_27, b_30, h_s_dadda_rca32_and_27_30_y0);
  fa fa_h_s_dadda_rca32_fa780_y2(h_s_dadda_rca32_and_29_28_y0, h_s_dadda_rca32_and_28_29_y0, h_s_dadda_rca32_and_27_30_y0, h_s_dadda_rca32_fa780_y2, h_s_dadda_rca32_fa780_y4);
  fa fa_h_s_dadda_rca32_fa781_y2(h_s_dadda_rca32_fa780_y4, h_s_dadda_rca32_fa779_y4, h_s_dadda_rca32_fa675_y4, h_s_dadda_rca32_fa781_y2, h_s_dadda_rca32_fa781_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_27_y0(a_31, b_27, h_s_dadda_rca32_nand_31_27_y0);
  and_gate and_gate_h_s_dadda_rca32_and_30_28_y0(a_30, b_28, h_s_dadda_rca32_and_30_28_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_29_y0(a_29, b_29, h_s_dadda_rca32_and_29_29_y0);
  fa fa_h_s_dadda_rca32_fa782_y2(h_s_dadda_rca32_nand_31_27_y0, h_s_dadda_rca32_and_30_28_y0, h_s_dadda_rca32_and_29_29_y0, h_s_dadda_rca32_fa782_y2, h_s_dadda_rca32_fa782_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_28_y0(a_31, b_28, h_s_dadda_rca32_nand_31_28_y0);
  fa fa_h_s_dadda_rca32_fa783_y2(h_s_dadda_rca32_fa782_y4, h_s_dadda_rca32_fa781_y4, h_s_dadda_rca32_nand_31_28_y0, h_s_dadda_rca32_fa783_y2, h_s_dadda_rca32_fa783_y4);
  and_gate and_gate_h_s_dadda_rca32_and_3_0_y0(a_3, b_0, h_s_dadda_rca32_and_3_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_2_1_y0(a_2, b_1, h_s_dadda_rca32_and_2_1_y0);
  ha ha_h_s_dadda_rca32_ha28_y0(h_s_dadda_rca32_and_3_0_y0, h_s_dadda_rca32_and_2_1_y0, h_s_dadda_rca32_ha28_y0, h_s_dadda_rca32_ha28_y1);
  and_gate and_gate_h_s_dadda_rca32_and_2_2_y0(a_2, b_2, h_s_dadda_rca32_and_2_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_3_y0(a_1, b_3, h_s_dadda_rca32_and_1_3_y0);
  fa fa_h_s_dadda_rca32_fa784_y2(h_s_dadda_rca32_ha28_y1, h_s_dadda_rca32_and_2_2_y0, h_s_dadda_rca32_and_1_3_y0, h_s_dadda_rca32_fa784_y2, h_s_dadda_rca32_fa784_y4);
  and_gate and_gate_h_s_dadda_rca32_and_1_4_y0(a_1, b_4, h_s_dadda_rca32_and_1_4_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_5_y0(a_0, b_5, h_s_dadda_rca32_and_0_5_y0);
  fa fa_h_s_dadda_rca32_fa785_y2(h_s_dadda_rca32_fa784_y4, h_s_dadda_rca32_and_1_4_y0, h_s_dadda_rca32_and_0_5_y0, h_s_dadda_rca32_fa785_y2, h_s_dadda_rca32_fa785_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_6_y0(a_0, b_6, h_s_dadda_rca32_and_0_6_y0);
  fa fa_h_s_dadda_rca32_fa786_y2(h_s_dadda_rca32_fa785_y4, h_s_dadda_rca32_and_0_6_y0, h_s_dadda_rca32_ha4_y0, h_s_dadda_rca32_fa786_y2, h_s_dadda_rca32_fa786_y4);
  fa fa_h_s_dadda_rca32_fa787_y2(h_s_dadda_rca32_fa786_y4, h_s_dadda_rca32_fa16_y2, h_s_dadda_rca32_ha5_y0, h_s_dadda_rca32_fa787_y2, h_s_dadda_rca32_fa787_y4);
  fa fa_h_s_dadda_rca32_fa788_y2(h_s_dadda_rca32_fa787_y4, h_s_dadda_rca32_fa18_y2, h_s_dadda_rca32_ha6_y0, h_s_dadda_rca32_fa788_y2, h_s_dadda_rca32_fa788_y4);
  fa fa_h_s_dadda_rca32_fa789_y2(h_s_dadda_rca32_fa788_y4, h_s_dadda_rca32_fa21_y2, h_s_dadda_rca32_ha7_y0, h_s_dadda_rca32_fa789_y2, h_s_dadda_rca32_fa789_y4);
  fa fa_h_s_dadda_rca32_fa790_y2(h_s_dadda_rca32_fa789_y4, h_s_dadda_rca32_fa25_y2, h_s_dadda_rca32_ha8_y0, h_s_dadda_rca32_fa790_y2, h_s_dadda_rca32_fa790_y4);
  fa fa_h_s_dadda_rca32_fa791_y2(h_s_dadda_rca32_fa790_y4, h_s_dadda_rca32_fa30_y2, h_s_dadda_rca32_ha9_y0, h_s_dadda_rca32_fa791_y2, h_s_dadda_rca32_fa791_y4);
  fa fa_h_s_dadda_rca32_fa792_y2(h_s_dadda_rca32_fa791_y4, h_s_dadda_rca32_fa36_y2, h_s_dadda_rca32_ha10_y0, h_s_dadda_rca32_fa792_y2, h_s_dadda_rca32_fa792_y4);
  fa fa_h_s_dadda_rca32_fa793_y2(h_s_dadda_rca32_fa792_y4, h_s_dadda_rca32_fa43_y2, h_s_dadda_rca32_ha11_y0, h_s_dadda_rca32_fa793_y2, h_s_dadda_rca32_fa793_y4);
  fa fa_h_s_dadda_rca32_fa794_y2(h_s_dadda_rca32_fa793_y4, h_s_dadda_rca32_fa51_y2, h_s_dadda_rca32_ha12_y0, h_s_dadda_rca32_fa794_y2, h_s_dadda_rca32_fa794_y4);
  fa fa_h_s_dadda_rca32_fa795_y2(h_s_dadda_rca32_fa794_y4, h_s_dadda_rca32_fa60_y2, h_s_dadda_rca32_ha13_y0, h_s_dadda_rca32_fa795_y2, h_s_dadda_rca32_fa795_y4);
  fa fa_h_s_dadda_rca32_fa796_y2(h_s_dadda_rca32_fa795_y4, h_s_dadda_rca32_fa70_y2, h_s_dadda_rca32_ha14_y0, h_s_dadda_rca32_fa796_y2, h_s_dadda_rca32_fa796_y4);
  fa fa_h_s_dadda_rca32_fa797_y2(h_s_dadda_rca32_fa796_y4, h_s_dadda_rca32_fa81_y2, h_s_dadda_rca32_ha15_y0, h_s_dadda_rca32_fa797_y2, h_s_dadda_rca32_fa797_y4);
  fa fa_h_s_dadda_rca32_fa798_y2(h_s_dadda_rca32_fa797_y4, h_s_dadda_rca32_fa93_y2, h_s_dadda_rca32_ha16_y0, h_s_dadda_rca32_fa798_y2, h_s_dadda_rca32_fa798_y4);
  fa fa_h_s_dadda_rca32_fa799_y2(h_s_dadda_rca32_fa798_y4, h_s_dadda_rca32_fa106_y2, h_s_dadda_rca32_ha17_y0, h_s_dadda_rca32_fa799_y2, h_s_dadda_rca32_fa799_y4);
  fa fa_h_s_dadda_rca32_fa800_y2(h_s_dadda_rca32_fa799_y4, h_s_dadda_rca32_fa120_y2, h_s_dadda_rca32_ha18_y0, h_s_dadda_rca32_fa800_y2, h_s_dadda_rca32_fa800_y4);
  fa fa_h_s_dadda_rca32_fa801_y2(h_s_dadda_rca32_fa800_y4, h_s_dadda_rca32_fa135_y2, h_s_dadda_rca32_ha19_y0, h_s_dadda_rca32_fa801_y2, h_s_dadda_rca32_fa801_y4);
  fa fa_h_s_dadda_rca32_fa802_y2(h_s_dadda_rca32_fa801_y4, h_s_dadda_rca32_fa151_y2, h_s_dadda_rca32_ha20_y0, h_s_dadda_rca32_fa802_y2, h_s_dadda_rca32_fa802_y4);
  fa fa_h_s_dadda_rca32_fa803_y2(h_s_dadda_rca32_fa802_y4, h_s_dadda_rca32_fa168_y2, h_s_dadda_rca32_ha21_y0, h_s_dadda_rca32_fa803_y2, h_s_dadda_rca32_fa803_y4);
  fa fa_h_s_dadda_rca32_fa804_y2(h_s_dadda_rca32_fa803_y4, h_s_dadda_rca32_fa186_y2, h_s_dadda_rca32_ha22_y0, h_s_dadda_rca32_fa804_y2, h_s_dadda_rca32_fa804_y4);
  fa fa_h_s_dadda_rca32_fa805_y2(h_s_dadda_rca32_fa804_y4, h_s_dadda_rca32_fa205_y2, h_s_dadda_rca32_ha23_y0, h_s_dadda_rca32_fa805_y2, h_s_dadda_rca32_fa805_y4);
  fa fa_h_s_dadda_rca32_fa806_y2(h_s_dadda_rca32_fa805_y4, h_s_dadda_rca32_fa225_y2, h_s_dadda_rca32_ha24_y0, h_s_dadda_rca32_fa806_y2, h_s_dadda_rca32_fa806_y4);
  fa fa_h_s_dadda_rca32_fa807_y2(h_s_dadda_rca32_fa806_y4, h_s_dadda_rca32_fa246_y2, h_s_dadda_rca32_ha25_y0, h_s_dadda_rca32_fa807_y2, h_s_dadda_rca32_fa807_y4);
  fa fa_h_s_dadda_rca32_fa808_y2(h_s_dadda_rca32_fa807_y4, h_s_dadda_rca32_fa267_y2, h_s_dadda_rca32_fa268_y2, h_s_dadda_rca32_fa808_y2, h_s_dadda_rca32_fa808_y4);
  fa fa_h_s_dadda_rca32_fa809_y2(h_s_dadda_rca32_fa808_y4, h_s_dadda_rca32_fa289_y2, h_s_dadda_rca32_fa290_y2, h_s_dadda_rca32_fa809_y2, h_s_dadda_rca32_fa809_y4);
  fa fa_h_s_dadda_rca32_fa810_y2(h_s_dadda_rca32_fa809_y4, h_s_dadda_rca32_fa311_y2, h_s_dadda_rca32_fa312_y2, h_s_dadda_rca32_fa810_y2, h_s_dadda_rca32_fa810_y4);
  fa fa_h_s_dadda_rca32_fa811_y2(h_s_dadda_rca32_fa810_y4, h_s_dadda_rca32_fa333_y2, h_s_dadda_rca32_fa334_y2, h_s_dadda_rca32_fa811_y2, h_s_dadda_rca32_fa811_y4);
  fa fa_h_s_dadda_rca32_fa812_y2(h_s_dadda_rca32_fa811_y4, h_s_dadda_rca32_fa355_y2, h_s_dadda_rca32_fa356_y2, h_s_dadda_rca32_fa812_y2, h_s_dadda_rca32_fa812_y4);
  fa fa_h_s_dadda_rca32_fa813_y2(h_s_dadda_rca32_fa812_y4, h_s_dadda_rca32_fa377_y2, h_s_dadda_rca32_fa378_y2, h_s_dadda_rca32_fa813_y2, h_s_dadda_rca32_fa813_y4);
  fa fa_h_s_dadda_rca32_fa814_y2(h_s_dadda_rca32_fa813_y4, h_s_dadda_rca32_fa399_y2, h_s_dadda_rca32_fa400_y2, h_s_dadda_rca32_fa814_y2, h_s_dadda_rca32_fa814_y4);
  fa fa_h_s_dadda_rca32_fa815_y2(h_s_dadda_rca32_fa814_y4, h_s_dadda_rca32_fa421_y2, h_s_dadda_rca32_fa422_y2, h_s_dadda_rca32_fa815_y2, h_s_dadda_rca32_fa815_y4);
  fa fa_h_s_dadda_rca32_fa816_y2(h_s_dadda_rca32_fa815_y4, h_s_dadda_rca32_fa443_y2, h_s_dadda_rca32_fa444_y2, h_s_dadda_rca32_fa816_y2, h_s_dadda_rca32_fa816_y4);
  fa fa_h_s_dadda_rca32_fa817_y2(h_s_dadda_rca32_fa816_y4, h_s_dadda_rca32_fa464_y2, h_s_dadda_rca32_fa465_y2, h_s_dadda_rca32_fa817_y2, h_s_dadda_rca32_fa817_y4);
  fa fa_h_s_dadda_rca32_fa818_y2(h_s_dadda_rca32_fa817_y4, h_s_dadda_rca32_fa484_y2, h_s_dadda_rca32_fa485_y2, h_s_dadda_rca32_fa818_y2, h_s_dadda_rca32_fa818_y4);
  fa fa_h_s_dadda_rca32_fa819_y2(h_s_dadda_rca32_fa818_y4, h_s_dadda_rca32_fa503_y2, h_s_dadda_rca32_fa504_y2, h_s_dadda_rca32_fa819_y2, h_s_dadda_rca32_fa819_y4);
  fa fa_h_s_dadda_rca32_fa820_y2(h_s_dadda_rca32_fa819_y4, h_s_dadda_rca32_fa521_y2, h_s_dadda_rca32_fa522_y2, h_s_dadda_rca32_fa820_y2, h_s_dadda_rca32_fa820_y4);
  fa fa_h_s_dadda_rca32_fa821_y2(h_s_dadda_rca32_fa820_y4, h_s_dadda_rca32_fa538_y2, h_s_dadda_rca32_fa539_y2, h_s_dadda_rca32_fa821_y2, h_s_dadda_rca32_fa821_y4);
  fa fa_h_s_dadda_rca32_fa822_y2(h_s_dadda_rca32_fa821_y4, h_s_dadda_rca32_fa554_y2, h_s_dadda_rca32_fa555_y2, h_s_dadda_rca32_fa822_y2, h_s_dadda_rca32_fa822_y4);
  fa fa_h_s_dadda_rca32_fa823_y2(h_s_dadda_rca32_fa822_y4, h_s_dadda_rca32_fa569_y2, h_s_dadda_rca32_fa570_y2, h_s_dadda_rca32_fa823_y2, h_s_dadda_rca32_fa823_y4);
  fa fa_h_s_dadda_rca32_fa824_y2(h_s_dadda_rca32_fa823_y4, h_s_dadda_rca32_fa583_y2, h_s_dadda_rca32_fa584_y2, h_s_dadda_rca32_fa824_y2, h_s_dadda_rca32_fa824_y4);
  fa fa_h_s_dadda_rca32_fa825_y2(h_s_dadda_rca32_fa824_y4, h_s_dadda_rca32_fa596_y2, h_s_dadda_rca32_fa597_y2, h_s_dadda_rca32_fa825_y2, h_s_dadda_rca32_fa825_y4);
  fa fa_h_s_dadda_rca32_fa826_y2(h_s_dadda_rca32_fa825_y4, h_s_dadda_rca32_fa608_y2, h_s_dadda_rca32_fa609_y2, h_s_dadda_rca32_fa826_y2, h_s_dadda_rca32_fa826_y4);
  fa fa_h_s_dadda_rca32_fa827_y2(h_s_dadda_rca32_fa826_y4, h_s_dadda_rca32_fa619_y2, h_s_dadda_rca32_fa620_y2, h_s_dadda_rca32_fa827_y2, h_s_dadda_rca32_fa827_y4);
  fa fa_h_s_dadda_rca32_fa828_y2(h_s_dadda_rca32_fa827_y4, h_s_dadda_rca32_fa629_y2, h_s_dadda_rca32_fa630_y2, h_s_dadda_rca32_fa828_y2, h_s_dadda_rca32_fa828_y4);
  fa fa_h_s_dadda_rca32_fa829_y2(h_s_dadda_rca32_fa828_y4, h_s_dadda_rca32_fa638_y2, h_s_dadda_rca32_fa639_y2, h_s_dadda_rca32_fa829_y2, h_s_dadda_rca32_fa829_y4);
  fa fa_h_s_dadda_rca32_fa830_y2(h_s_dadda_rca32_fa829_y4, h_s_dadda_rca32_fa646_y2, h_s_dadda_rca32_fa647_y2, h_s_dadda_rca32_fa830_y2, h_s_dadda_rca32_fa830_y4);
  fa fa_h_s_dadda_rca32_fa831_y2(h_s_dadda_rca32_fa830_y4, h_s_dadda_rca32_fa653_y2, h_s_dadda_rca32_fa654_y2, h_s_dadda_rca32_fa831_y2, h_s_dadda_rca32_fa831_y4);
  fa fa_h_s_dadda_rca32_fa832_y2(h_s_dadda_rca32_fa831_y4, h_s_dadda_rca32_fa659_y2, h_s_dadda_rca32_fa660_y2, h_s_dadda_rca32_fa832_y2, h_s_dadda_rca32_fa832_y4);
  fa fa_h_s_dadda_rca32_fa833_y2(h_s_dadda_rca32_fa832_y4, h_s_dadda_rca32_fa664_y2, h_s_dadda_rca32_fa665_y2, h_s_dadda_rca32_fa833_y2, h_s_dadda_rca32_fa833_y4);
  fa fa_h_s_dadda_rca32_fa834_y2(h_s_dadda_rca32_fa833_y4, h_s_dadda_rca32_fa668_y2, h_s_dadda_rca32_fa669_y2, h_s_dadda_rca32_fa834_y2, h_s_dadda_rca32_fa834_y4);
  fa fa_h_s_dadda_rca32_fa835_y2(h_s_dadda_rca32_fa834_y4, h_s_dadda_rca32_fa671_y2, h_s_dadda_rca32_fa672_y2, h_s_dadda_rca32_fa835_y2, h_s_dadda_rca32_fa835_y4);
  fa fa_h_s_dadda_rca32_fa836_y2(h_s_dadda_rca32_fa835_y4, h_s_dadda_rca32_fa673_y2, h_s_dadda_rca32_fa674_y2, h_s_dadda_rca32_fa836_y2, h_s_dadda_rca32_fa836_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_26_31_y0(a_26, b_31, h_s_dadda_rca32_nand_26_31_y0);
  fa fa_h_s_dadda_rca32_fa837_y2(h_s_dadda_rca32_fa836_y4, h_s_dadda_rca32_nand_26_31_y0, h_s_dadda_rca32_fa675_y2, h_s_dadda_rca32_fa837_y2, h_s_dadda_rca32_fa837_y4);
  and_gate and_gate_h_s_dadda_rca32_and_28_30_y0(a_28, b_30, h_s_dadda_rca32_and_28_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_27_31_y0(a_27, b_31, h_s_dadda_rca32_nand_27_31_y0);
  fa fa_h_s_dadda_rca32_fa838_y2(h_s_dadda_rca32_fa837_y4, h_s_dadda_rca32_and_28_30_y0, h_s_dadda_rca32_nand_27_31_y0, h_s_dadda_rca32_fa838_y2, h_s_dadda_rca32_fa838_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_29_y0(a_30, b_29, h_s_dadda_rca32_and_30_29_y0);
  and_gate and_gate_h_s_dadda_rca32_and_29_30_y0(a_29, b_30, h_s_dadda_rca32_and_29_30_y0);
  fa fa_h_s_dadda_rca32_fa839_y2(h_s_dadda_rca32_fa838_y4, h_s_dadda_rca32_and_30_29_y0, h_s_dadda_rca32_and_29_30_y0, h_s_dadda_rca32_fa839_y2, h_s_dadda_rca32_fa839_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_29_y0(a_31, b_29, h_s_dadda_rca32_nand_31_29_y0);
  fa fa_h_s_dadda_rca32_fa840_y2(h_s_dadda_rca32_fa839_y4, h_s_dadda_rca32_fa783_y4, h_s_dadda_rca32_nand_31_29_y0, h_s_dadda_rca32_fa840_y2, h_s_dadda_rca32_fa840_y4);
  and_gate and_gate_h_s_dadda_rca32_and_2_0_y0(a_2, b_0, h_s_dadda_rca32_and_2_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_1_y0(a_1, b_1, h_s_dadda_rca32_and_1_1_y0);
  ha ha_h_s_dadda_rca32_ha29_y0(h_s_dadda_rca32_and_2_0_y0, h_s_dadda_rca32_and_1_1_y0, h_s_dadda_rca32_ha29_y0, h_s_dadda_rca32_ha29_y1);
  and_gate and_gate_h_s_dadda_rca32_and_1_2_y0(a_1, b_2, h_s_dadda_rca32_and_1_2_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_3_y0(a_0, b_3, h_s_dadda_rca32_and_0_3_y0);
  fa fa_h_s_dadda_rca32_fa841_y2(h_s_dadda_rca32_ha29_y1, h_s_dadda_rca32_and_1_2_y0, h_s_dadda_rca32_and_0_3_y0, h_s_dadda_rca32_fa841_y2, h_s_dadda_rca32_fa841_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_4_y0(a_0, b_4, h_s_dadda_rca32_and_0_4_y0);
  fa fa_h_s_dadda_rca32_fa842_y2(h_s_dadda_rca32_fa841_y4, h_s_dadda_rca32_and_0_4_y0, h_s_dadda_rca32_ha26_y0, h_s_dadda_rca32_fa842_y2, h_s_dadda_rca32_fa842_y4);
  fa fa_h_s_dadda_rca32_fa843_y2(h_s_dadda_rca32_fa842_y4, h_s_dadda_rca32_fa676_y2, h_s_dadda_rca32_ha27_y0, h_s_dadda_rca32_fa843_y2, h_s_dadda_rca32_fa843_y4);
  fa fa_h_s_dadda_rca32_fa844_y2(h_s_dadda_rca32_fa843_y4, h_s_dadda_rca32_fa677_y2, h_s_dadda_rca32_fa678_y2, h_s_dadda_rca32_fa844_y2, h_s_dadda_rca32_fa844_y4);
  fa fa_h_s_dadda_rca32_fa845_y2(h_s_dadda_rca32_fa844_y4, h_s_dadda_rca32_fa679_y2, h_s_dadda_rca32_fa680_y2, h_s_dadda_rca32_fa845_y2, h_s_dadda_rca32_fa845_y4);
  fa fa_h_s_dadda_rca32_fa846_y2(h_s_dadda_rca32_fa845_y4, h_s_dadda_rca32_fa681_y2, h_s_dadda_rca32_fa682_y2, h_s_dadda_rca32_fa846_y2, h_s_dadda_rca32_fa846_y4);
  fa fa_h_s_dadda_rca32_fa847_y2(h_s_dadda_rca32_fa846_y4, h_s_dadda_rca32_fa683_y2, h_s_dadda_rca32_fa684_y2, h_s_dadda_rca32_fa847_y2, h_s_dadda_rca32_fa847_y4);
  fa fa_h_s_dadda_rca32_fa848_y2(h_s_dadda_rca32_fa847_y4, h_s_dadda_rca32_fa685_y2, h_s_dadda_rca32_fa686_y2, h_s_dadda_rca32_fa848_y2, h_s_dadda_rca32_fa848_y4);
  fa fa_h_s_dadda_rca32_fa849_y2(h_s_dadda_rca32_fa848_y4, h_s_dadda_rca32_fa687_y2, h_s_dadda_rca32_fa688_y2, h_s_dadda_rca32_fa849_y2, h_s_dadda_rca32_fa849_y4);
  fa fa_h_s_dadda_rca32_fa850_y2(h_s_dadda_rca32_fa849_y4, h_s_dadda_rca32_fa689_y2, h_s_dadda_rca32_fa690_y2, h_s_dadda_rca32_fa850_y2, h_s_dadda_rca32_fa850_y4);
  fa fa_h_s_dadda_rca32_fa851_y2(h_s_dadda_rca32_fa850_y4, h_s_dadda_rca32_fa691_y2, h_s_dadda_rca32_fa692_y2, h_s_dadda_rca32_fa851_y2, h_s_dadda_rca32_fa851_y4);
  fa fa_h_s_dadda_rca32_fa852_y2(h_s_dadda_rca32_fa851_y4, h_s_dadda_rca32_fa693_y2, h_s_dadda_rca32_fa694_y2, h_s_dadda_rca32_fa852_y2, h_s_dadda_rca32_fa852_y4);
  fa fa_h_s_dadda_rca32_fa853_y2(h_s_dadda_rca32_fa852_y4, h_s_dadda_rca32_fa695_y2, h_s_dadda_rca32_fa696_y2, h_s_dadda_rca32_fa853_y2, h_s_dadda_rca32_fa853_y4);
  fa fa_h_s_dadda_rca32_fa854_y2(h_s_dadda_rca32_fa853_y4, h_s_dadda_rca32_fa697_y2, h_s_dadda_rca32_fa698_y2, h_s_dadda_rca32_fa854_y2, h_s_dadda_rca32_fa854_y4);
  fa fa_h_s_dadda_rca32_fa855_y2(h_s_dadda_rca32_fa854_y4, h_s_dadda_rca32_fa699_y2, h_s_dadda_rca32_fa700_y2, h_s_dadda_rca32_fa855_y2, h_s_dadda_rca32_fa855_y4);
  fa fa_h_s_dadda_rca32_fa856_y2(h_s_dadda_rca32_fa855_y4, h_s_dadda_rca32_fa701_y2, h_s_dadda_rca32_fa702_y2, h_s_dadda_rca32_fa856_y2, h_s_dadda_rca32_fa856_y4);
  fa fa_h_s_dadda_rca32_fa857_y2(h_s_dadda_rca32_fa856_y4, h_s_dadda_rca32_fa703_y2, h_s_dadda_rca32_fa704_y2, h_s_dadda_rca32_fa857_y2, h_s_dadda_rca32_fa857_y4);
  fa fa_h_s_dadda_rca32_fa858_y2(h_s_dadda_rca32_fa857_y4, h_s_dadda_rca32_fa705_y2, h_s_dadda_rca32_fa706_y2, h_s_dadda_rca32_fa858_y2, h_s_dadda_rca32_fa858_y4);
  fa fa_h_s_dadda_rca32_fa859_y2(h_s_dadda_rca32_fa858_y4, h_s_dadda_rca32_fa707_y2, h_s_dadda_rca32_fa708_y2, h_s_dadda_rca32_fa859_y2, h_s_dadda_rca32_fa859_y4);
  fa fa_h_s_dadda_rca32_fa860_y2(h_s_dadda_rca32_fa859_y4, h_s_dadda_rca32_fa709_y2, h_s_dadda_rca32_fa710_y2, h_s_dadda_rca32_fa860_y2, h_s_dadda_rca32_fa860_y4);
  fa fa_h_s_dadda_rca32_fa861_y2(h_s_dadda_rca32_fa860_y4, h_s_dadda_rca32_fa711_y2, h_s_dadda_rca32_fa712_y2, h_s_dadda_rca32_fa861_y2, h_s_dadda_rca32_fa861_y4);
  fa fa_h_s_dadda_rca32_fa862_y2(h_s_dadda_rca32_fa861_y4, h_s_dadda_rca32_fa713_y2, h_s_dadda_rca32_fa714_y2, h_s_dadda_rca32_fa862_y2, h_s_dadda_rca32_fa862_y4);
  fa fa_h_s_dadda_rca32_fa863_y2(h_s_dadda_rca32_fa862_y4, h_s_dadda_rca32_fa715_y2, h_s_dadda_rca32_fa716_y2, h_s_dadda_rca32_fa863_y2, h_s_dadda_rca32_fa863_y4);
  fa fa_h_s_dadda_rca32_fa864_y2(h_s_dadda_rca32_fa863_y4, h_s_dadda_rca32_fa717_y2, h_s_dadda_rca32_fa718_y2, h_s_dadda_rca32_fa864_y2, h_s_dadda_rca32_fa864_y4);
  fa fa_h_s_dadda_rca32_fa865_y2(h_s_dadda_rca32_fa864_y4, h_s_dadda_rca32_fa719_y2, h_s_dadda_rca32_fa720_y2, h_s_dadda_rca32_fa865_y2, h_s_dadda_rca32_fa865_y4);
  fa fa_h_s_dadda_rca32_fa866_y2(h_s_dadda_rca32_fa865_y4, h_s_dadda_rca32_fa721_y2, h_s_dadda_rca32_fa722_y2, h_s_dadda_rca32_fa866_y2, h_s_dadda_rca32_fa866_y4);
  fa fa_h_s_dadda_rca32_fa867_y2(h_s_dadda_rca32_fa866_y4, h_s_dadda_rca32_fa723_y2, h_s_dadda_rca32_fa724_y2, h_s_dadda_rca32_fa867_y2, h_s_dadda_rca32_fa867_y4);
  fa fa_h_s_dadda_rca32_fa868_y2(h_s_dadda_rca32_fa867_y4, h_s_dadda_rca32_fa725_y2, h_s_dadda_rca32_fa726_y2, h_s_dadda_rca32_fa868_y2, h_s_dadda_rca32_fa868_y4);
  fa fa_h_s_dadda_rca32_fa869_y2(h_s_dadda_rca32_fa868_y4, h_s_dadda_rca32_fa727_y2, h_s_dadda_rca32_fa728_y2, h_s_dadda_rca32_fa869_y2, h_s_dadda_rca32_fa869_y4);
  fa fa_h_s_dadda_rca32_fa870_y2(h_s_dadda_rca32_fa869_y4, h_s_dadda_rca32_fa729_y2, h_s_dadda_rca32_fa730_y2, h_s_dadda_rca32_fa870_y2, h_s_dadda_rca32_fa870_y4);
  fa fa_h_s_dadda_rca32_fa871_y2(h_s_dadda_rca32_fa870_y4, h_s_dadda_rca32_fa731_y2, h_s_dadda_rca32_fa732_y2, h_s_dadda_rca32_fa871_y2, h_s_dadda_rca32_fa871_y4);
  fa fa_h_s_dadda_rca32_fa872_y2(h_s_dadda_rca32_fa871_y4, h_s_dadda_rca32_fa733_y2, h_s_dadda_rca32_fa734_y2, h_s_dadda_rca32_fa872_y2, h_s_dadda_rca32_fa872_y4);
  fa fa_h_s_dadda_rca32_fa873_y2(h_s_dadda_rca32_fa872_y4, h_s_dadda_rca32_fa735_y2, h_s_dadda_rca32_fa736_y2, h_s_dadda_rca32_fa873_y2, h_s_dadda_rca32_fa873_y4);
  fa fa_h_s_dadda_rca32_fa874_y2(h_s_dadda_rca32_fa873_y4, h_s_dadda_rca32_fa737_y2, h_s_dadda_rca32_fa738_y2, h_s_dadda_rca32_fa874_y2, h_s_dadda_rca32_fa874_y4);
  fa fa_h_s_dadda_rca32_fa875_y2(h_s_dadda_rca32_fa874_y4, h_s_dadda_rca32_fa739_y2, h_s_dadda_rca32_fa740_y2, h_s_dadda_rca32_fa875_y2, h_s_dadda_rca32_fa875_y4);
  fa fa_h_s_dadda_rca32_fa876_y2(h_s_dadda_rca32_fa875_y4, h_s_dadda_rca32_fa741_y2, h_s_dadda_rca32_fa742_y2, h_s_dadda_rca32_fa876_y2, h_s_dadda_rca32_fa876_y4);
  fa fa_h_s_dadda_rca32_fa877_y2(h_s_dadda_rca32_fa876_y4, h_s_dadda_rca32_fa743_y2, h_s_dadda_rca32_fa744_y2, h_s_dadda_rca32_fa877_y2, h_s_dadda_rca32_fa877_y4);
  fa fa_h_s_dadda_rca32_fa878_y2(h_s_dadda_rca32_fa877_y4, h_s_dadda_rca32_fa745_y2, h_s_dadda_rca32_fa746_y2, h_s_dadda_rca32_fa878_y2, h_s_dadda_rca32_fa878_y4);
  fa fa_h_s_dadda_rca32_fa879_y2(h_s_dadda_rca32_fa878_y4, h_s_dadda_rca32_fa747_y2, h_s_dadda_rca32_fa748_y2, h_s_dadda_rca32_fa879_y2, h_s_dadda_rca32_fa879_y4);
  fa fa_h_s_dadda_rca32_fa880_y2(h_s_dadda_rca32_fa879_y4, h_s_dadda_rca32_fa749_y2, h_s_dadda_rca32_fa750_y2, h_s_dadda_rca32_fa880_y2, h_s_dadda_rca32_fa880_y4);
  fa fa_h_s_dadda_rca32_fa881_y2(h_s_dadda_rca32_fa880_y4, h_s_dadda_rca32_fa751_y2, h_s_dadda_rca32_fa752_y2, h_s_dadda_rca32_fa881_y2, h_s_dadda_rca32_fa881_y4);
  fa fa_h_s_dadda_rca32_fa882_y2(h_s_dadda_rca32_fa881_y4, h_s_dadda_rca32_fa753_y2, h_s_dadda_rca32_fa754_y2, h_s_dadda_rca32_fa882_y2, h_s_dadda_rca32_fa882_y4);
  fa fa_h_s_dadda_rca32_fa883_y2(h_s_dadda_rca32_fa882_y4, h_s_dadda_rca32_fa755_y2, h_s_dadda_rca32_fa756_y2, h_s_dadda_rca32_fa883_y2, h_s_dadda_rca32_fa883_y4);
  fa fa_h_s_dadda_rca32_fa884_y2(h_s_dadda_rca32_fa883_y4, h_s_dadda_rca32_fa757_y2, h_s_dadda_rca32_fa758_y2, h_s_dadda_rca32_fa884_y2, h_s_dadda_rca32_fa884_y4);
  fa fa_h_s_dadda_rca32_fa885_y2(h_s_dadda_rca32_fa884_y4, h_s_dadda_rca32_fa759_y2, h_s_dadda_rca32_fa760_y2, h_s_dadda_rca32_fa885_y2, h_s_dadda_rca32_fa885_y4);
  fa fa_h_s_dadda_rca32_fa886_y2(h_s_dadda_rca32_fa885_y4, h_s_dadda_rca32_fa761_y2, h_s_dadda_rca32_fa762_y2, h_s_dadda_rca32_fa886_y2, h_s_dadda_rca32_fa886_y4);
  fa fa_h_s_dadda_rca32_fa887_y2(h_s_dadda_rca32_fa886_y4, h_s_dadda_rca32_fa763_y2, h_s_dadda_rca32_fa764_y2, h_s_dadda_rca32_fa887_y2, h_s_dadda_rca32_fa887_y4);
  fa fa_h_s_dadda_rca32_fa888_y2(h_s_dadda_rca32_fa887_y4, h_s_dadda_rca32_fa765_y2, h_s_dadda_rca32_fa766_y2, h_s_dadda_rca32_fa888_y2, h_s_dadda_rca32_fa888_y4);
  fa fa_h_s_dadda_rca32_fa889_y2(h_s_dadda_rca32_fa888_y4, h_s_dadda_rca32_fa767_y2, h_s_dadda_rca32_fa768_y2, h_s_dadda_rca32_fa889_y2, h_s_dadda_rca32_fa889_y4);
  fa fa_h_s_dadda_rca32_fa890_y2(h_s_dadda_rca32_fa889_y4, h_s_dadda_rca32_fa769_y2, h_s_dadda_rca32_fa770_y2, h_s_dadda_rca32_fa890_y2, h_s_dadda_rca32_fa890_y4);
  fa fa_h_s_dadda_rca32_fa891_y2(h_s_dadda_rca32_fa890_y4, h_s_dadda_rca32_fa771_y2, h_s_dadda_rca32_fa772_y2, h_s_dadda_rca32_fa891_y2, h_s_dadda_rca32_fa891_y4);
  fa fa_h_s_dadda_rca32_fa892_y2(h_s_dadda_rca32_fa891_y4, h_s_dadda_rca32_fa773_y2, h_s_dadda_rca32_fa774_y2, h_s_dadda_rca32_fa892_y2, h_s_dadda_rca32_fa892_y4);
  fa fa_h_s_dadda_rca32_fa893_y2(h_s_dadda_rca32_fa892_y4, h_s_dadda_rca32_fa775_y2, h_s_dadda_rca32_fa776_y2, h_s_dadda_rca32_fa893_y2, h_s_dadda_rca32_fa893_y4);
  fa fa_h_s_dadda_rca32_fa894_y2(h_s_dadda_rca32_fa893_y4, h_s_dadda_rca32_fa777_y2, h_s_dadda_rca32_fa778_y2, h_s_dadda_rca32_fa894_y2, h_s_dadda_rca32_fa894_y4);
  fa fa_h_s_dadda_rca32_fa895_y2(h_s_dadda_rca32_fa894_y4, h_s_dadda_rca32_fa779_y2, h_s_dadda_rca32_fa780_y2, h_s_dadda_rca32_fa895_y2, h_s_dadda_rca32_fa895_y4);
  fa fa_h_s_dadda_rca32_fa896_y2(h_s_dadda_rca32_fa895_y4, h_s_dadda_rca32_fa781_y2, h_s_dadda_rca32_fa782_y2, h_s_dadda_rca32_fa896_y2, h_s_dadda_rca32_fa896_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_28_31_y0(a_28, b_31, h_s_dadda_rca32_nand_28_31_y0);
  fa fa_h_s_dadda_rca32_fa897_y2(h_s_dadda_rca32_fa896_y4, h_s_dadda_rca32_nand_28_31_y0, h_s_dadda_rca32_fa783_y2, h_s_dadda_rca32_fa897_y2, h_s_dadda_rca32_fa897_y4);
  and_gate and_gate_h_s_dadda_rca32_and_30_30_y0(a_30, b_30, h_s_dadda_rca32_and_30_30_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_29_31_y0(a_29, b_31, h_s_dadda_rca32_nand_29_31_y0);
  fa fa_h_s_dadda_rca32_fa898_y2(h_s_dadda_rca32_fa897_y4, h_s_dadda_rca32_and_30_30_y0, h_s_dadda_rca32_nand_29_31_y0, h_s_dadda_rca32_fa898_y2, h_s_dadda_rca32_fa898_y4);
  nand_gate nand_gate_h_s_dadda_rca32_nand_31_30_y0(a_31, b_30, h_s_dadda_rca32_nand_31_30_y0);
  fa fa_h_s_dadda_rca32_fa899_y2(h_s_dadda_rca32_fa898_y4, h_s_dadda_rca32_fa840_y4, h_s_dadda_rca32_nand_31_30_y0, h_s_dadda_rca32_fa899_y2, h_s_dadda_rca32_fa899_y4);
  and_gate and_gate_h_s_dadda_rca32_and_0_0_y0(a_0, b_0, h_s_dadda_rca32_and_0_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_1_0_y0(a_1, b_0, h_s_dadda_rca32_and_1_0_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_2_y0(a_0, b_2, h_s_dadda_rca32_and_0_2_y0);
  nand_gate nand_gate_h_s_dadda_rca32_nand_30_31_y0(a_30, b_31, h_s_dadda_rca32_nand_30_31_y0);
  and_gate and_gate_h_s_dadda_rca32_and_0_1_y0(a_0, b_1, h_s_dadda_rca32_and_0_1_y0);
  and_gate and_gate_h_s_dadda_rca32_and_31_31_y0(a_31, b_31, h_s_dadda_rca32_and_31_31_y0);
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[0] = h_s_dadda_rca32_and_1_0_y0;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[1] = h_s_dadda_rca32_and_0_2_y0;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[2] = h_s_dadda_rca32_ha28_y0;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[3] = h_s_dadda_rca32_fa784_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[4] = h_s_dadda_rca32_fa785_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[5] = h_s_dadda_rca32_fa786_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[6] = h_s_dadda_rca32_fa787_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[7] = h_s_dadda_rca32_fa788_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[8] = h_s_dadda_rca32_fa789_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[9] = h_s_dadda_rca32_fa790_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[10] = h_s_dadda_rca32_fa791_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[11] = h_s_dadda_rca32_fa792_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[12] = h_s_dadda_rca32_fa793_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[13] = h_s_dadda_rca32_fa794_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[14] = h_s_dadda_rca32_fa795_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[15] = h_s_dadda_rca32_fa796_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[16] = h_s_dadda_rca32_fa797_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[17] = h_s_dadda_rca32_fa798_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[18] = h_s_dadda_rca32_fa799_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[19] = h_s_dadda_rca32_fa800_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[20] = h_s_dadda_rca32_fa801_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[21] = h_s_dadda_rca32_fa802_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[22] = h_s_dadda_rca32_fa803_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[23] = h_s_dadda_rca32_fa804_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[24] = h_s_dadda_rca32_fa805_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[25] = h_s_dadda_rca32_fa806_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[26] = h_s_dadda_rca32_fa807_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[27] = h_s_dadda_rca32_fa808_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[28] = h_s_dadda_rca32_fa809_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[29] = h_s_dadda_rca32_fa810_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[30] = h_s_dadda_rca32_fa811_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[31] = h_s_dadda_rca32_fa812_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[32] = h_s_dadda_rca32_fa813_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[33] = h_s_dadda_rca32_fa814_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[34] = h_s_dadda_rca32_fa815_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[35] = h_s_dadda_rca32_fa816_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[36] = h_s_dadda_rca32_fa817_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[37] = h_s_dadda_rca32_fa818_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[38] = h_s_dadda_rca32_fa819_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[39] = h_s_dadda_rca32_fa820_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[40] = h_s_dadda_rca32_fa821_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[41] = h_s_dadda_rca32_fa822_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[42] = h_s_dadda_rca32_fa823_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[43] = h_s_dadda_rca32_fa824_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[44] = h_s_dadda_rca32_fa825_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[45] = h_s_dadda_rca32_fa826_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[46] = h_s_dadda_rca32_fa827_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[47] = h_s_dadda_rca32_fa828_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[48] = h_s_dadda_rca32_fa829_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[49] = h_s_dadda_rca32_fa830_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[50] = h_s_dadda_rca32_fa831_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[51] = h_s_dadda_rca32_fa832_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[52] = h_s_dadda_rca32_fa833_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[53] = h_s_dadda_rca32_fa834_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[54] = h_s_dadda_rca32_fa835_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[55] = h_s_dadda_rca32_fa836_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[56] = h_s_dadda_rca32_fa837_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[57] = h_s_dadda_rca32_fa838_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[58] = h_s_dadda_rca32_fa839_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[59] = h_s_dadda_rca32_fa840_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[60] = h_s_dadda_rca32_nand_30_31_y0;
  assign h_s_dadda_rca32_u_rca62_u_rca62_a[61] = h_s_dadda_rca32_fa899_y4;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[0] = h_s_dadda_rca32_and_0_1_y0;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[1] = h_s_dadda_rca32_ha29_y0;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[2] = h_s_dadda_rca32_fa841_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[3] = h_s_dadda_rca32_fa842_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[4] = h_s_dadda_rca32_fa843_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[5] = h_s_dadda_rca32_fa844_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[6] = h_s_dadda_rca32_fa845_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[7] = h_s_dadda_rca32_fa846_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[8] = h_s_dadda_rca32_fa847_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[9] = h_s_dadda_rca32_fa848_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[10] = h_s_dadda_rca32_fa849_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[11] = h_s_dadda_rca32_fa850_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[12] = h_s_dadda_rca32_fa851_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[13] = h_s_dadda_rca32_fa852_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[14] = h_s_dadda_rca32_fa853_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[15] = h_s_dadda_rca32_fa854_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[16] = h_s_dadda_rca32_fa855_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[17] = h_s_dadda_rca32_fa856_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[18] = h_s_dadda_rca32_fa857_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[19] = h_s_dadda_rca32_fa858_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[20] = h_s_dadda_rca32_fa859_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[21] = h_s_dadda_rca32_fa860_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[22] = h_s_dadda_rca32_fa861_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[23] = h_s_dadda_rca32_fa862_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[24] = h_s_dadda_rca32_fa863_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[25] = h_s_dadda_rca32_fa864_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[26] = h_s_dadda_rca32_fa865_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[27] = h_s_dadda_rca32_fa866_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[28] = h_s_dadda_rca32_fa867_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[29] = h_s_dadda_rca32_fa868_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[30] = h_s_dadda_rca32_fa869_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[31] = h_s_dadda_rca32_fa870_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[32] = h_s_dadda_rca32_fa871_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[33] = h_s_dadda_rca32_fa872_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[34] = h_s_dadda_rca32_fa873_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[35] = h_s_dadda_rca32_fa874_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[36] = h_s_dadda_rca32_fa875_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[37] = h_s_dadda_rca32_fa876_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[38] = h_s_dadda_rca32_fa877_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[39] = h_s_dadda_rca32_fa878_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[40] = h_s_dadda_rca32_fa879_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[41] = h_s_dadda_rca32_fa880_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[42] = h_s_dadda_rca32_fa881_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[43] = h_s_dadda_rca32_fa882_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[44] = h_s_dadda_rca32_fa883_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[45] = h_s_dadda_rca32_fa884_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[46] = h_s_dadda_rca32_fa885_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[47] = h_s_dadda_rca32_fa886_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[48] = h_s_dadda_rca32_fa887_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[49] = h_s_dadda_rca32_fa888_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[50] = h_s_dadda_rca32_fa889_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[51] = h_s_dadda_rca32_fa890_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[52] = h_s_dadda_rca32_fa891_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[53] = h_s_dadda_rca32_fa892_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[54] = h_s_dadda_rca32_fa893_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[55] = h_s_dadda_rca32_fa894_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[56] = h_s_dadda_rca32_fa895_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[57] = h_s_dadda_rca32_fa896_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[58] = h_s_dadda_rca32_fa897_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[59] = h_s_dadda_rca32_fa898_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[60] = h_s_dadda_rca32_fa899_y2;
  assign h_s_dadda_rca32_u_rca62_u_rca62_b[61] = h_s_dadda_rca32_and_31_31_y0;
  u_rca62 u_rca62_out(h_s_dadda_rca32_u_rca62_u_rca62_a, h_s_dadda_rca32_u_rca62_u_rca62_b, h_s_dadda_rca32_u_rca62_out);
  assign h_s_dadda_rca32_u_rca62_ha_y0 = h_s_dadda_rca32_u_rca62_out[0];
  assign h_s_dadda_rca32_u_rca62_fa1_y2 = h_s_dadda_rca32_u_rca62_out[1];
  assign h_s_dadda_rca32_u_rca62_fa2_y2 = h_s_dadda_rca32_u_rca62_out[2];
  assign h_s_dadda_rca32_u_rca62_fa3_y2 = h_s_dadda_rca32_u_rca62_out[3];
  assign h_s_dadda_rca32_u_rca62_fa4_y2 = h_s_dadda_rca32_u_rca62_out[4];
  assign h_s_dadda_rca32_u_rca62_fa5_y2 = h_s_dadda_rca32_u_rca62_out[5];
  assign h_s_dadda_rca32_u_rca62_fa6_y2 = h_s_dadda_rca32_u_rca62_out[6];
  assign h_s_dadda_rca32_u_rca62_fa7_y2 = h_s_dadda_rca32_u_rca62_out[7];
  assign h_s_dadda_rca32_u_rca62_fa8_y2 = h_s_dadda_rca32_u_rca62_out[8];
  assign h_s_dadda_rca32_u_rca62_fa9_y2 = h_s_dadda_rca32_u_rca62_out[9];
  assign h_s_dadda_rca32_u_rca62_fa10_y2 = h_s_dadda_rca32_u_rca62_out[10];
  assign h_s_dadda_rca32_u_rca62_fa11_y2 = h_s_dadda_rca32_u_rca62_out[11];
  assign h_s_dadda_rca32_u_rca62_fa12_y2 = h_s_dadda_rca32_u_rca62_out[12];
  assign h_s_dadda_rca32_u_rca62_fa13_y2 = h_s_dadda_rca32_u_rca62_out[13];
  assign h_s_dadda_rca32_u_rca62_fa14_y2 = h_s_dadda_rca32_u_rca62_out[14];
  assign h_s_dadda_rca32_u_rca62_fa15_y2 = h_s_dadda_rca32_u_rca62_out[15];
  assign h_s_dadda_rca32_u_rca62_fa16_y2 = h_s_dadda_rca32_u_rca62_out[16];
  assign h_s_dadda_rca32_u_rca62_fa17_y2 = h_s_dadda_rca32_u_rca62_out[17];
  assign h_s_dadda_rca32_u_rca62_fa18_y2 = h_s_dadda_rca32_u_rca62_out[18];
  assign h_s_dadda_rca32_u_rca62_fa19_y2 = h_s_dadda_rca32_u_rca62_out[19];
  assign h_s_dadda_rca32_u_rca62_fa20_y2 = h_s_dadda_rca32_u_rca62_out[20];
  assign h_s_dadda_rca32_u_rca62_fa21_y2 = h_s_dadda_rca32_u_rca62_out[21];
  assign h_s_dadda_rca32_u_rca62_fa22_y2 = h_s_dadda_rca32_u_rca62_out[22];
  assign h_s_dadda_rca32_u_rca62_fa23_y2 = h_s_dadda_rca32_u_rca62_out[23];
  assign h_s_dadda_rca32_u_rca62_fa24_y2 = h_s_dadda_rca32_u_rca62_out[24];
  assign h_s_dadda_rca32_u_rca62_fa25_y2 = h_s_dadda_rca32_u_rca62_out[25];
  assign h_s_dadda_rca32_u_rca62_fa26_y2 = h_s_dadda_rca32_u_rca62_out[26];
  assign h_s_dadda_rca32_u_rca62_fa27_y2 = h_s_dadda_rca32_u_rca62_out[27];
  assign h_s_dadda_rca32_u_rca62_fa28_y2 = h_s_dadda_rca32_u_rca62_out[28];
  assign h_s_dadda_rca32_u_rca62_fa29_y2 = h_s_dadda_rca32_u_rca62_out[29];
  assign h_s_dadda_rca32_u_rca62_fa30_y2 = h_s_dadda_rca32_u_rca62_out[30];
  assign h_s_dadda_rca32_u_rca62_fa31_y2 = h_s_dadda_rca32_u_rca62_out[31];
  assign h_s_dadda_rca32_u_rca62_fa32_y2 = h_s_dadda_rca32_u_rca62_out[32];
  assign h_s_dadda_rca32_u_rca62_fa33_y2 = h_s_dadda_rca32_u_rca62_out[33];
  assign h_s_dadda_rca32_u_rca62_fa34_y2 = h_s_dadda_rca32_u_rca62_out[34];
  assign h_s_dadda_rca32_u_rca62_fa35_y2 = h_s_dadda_rca32_u_rca62_out[35];
  assign h_s_dadda_rca32_u_rca62_fa36_y2 = h_s_dadda_rca32_u_rca62_out[36];
  assign h_s_dadda_rca32_u_rca62_fa37_y2 = h_s_dadda_rca32_u_rca62_out[37];
  assign h_s_dadda_rca32_u_rca62_fa38_y2 = h_s_dadda_rca32_u_rca62_out[38];
  assign h_s_dadda_rca32_u_rca62_fa39_y2 = h_s_dadda_rca32_u_rca62_out[39];
  assign h_s_dadda_rca32_u_rca62_fa40_y2 = h_s_dadda_rca32_u_rca62_out[40];
  assign h_s_dadda_rca32_u_rca62_fa41_y2 = h_s_dadda_rca32_u_rca62_out[41];
  assign h_s_dadda_rca32_u_rca62_fa42_y2 = h_s_dadda_rca32_u_rca62_out[42];
  assign h_s_dadda_rca32_u_rca62_fa43_y2 = h_s_dadda_rca32_u_rca62_out[43];
  assign h_s_dadda_rca32_u_rca62_fa44_y2 = h_s_dadda_rca32_u_rca62_out[44];
  assign h_s_dadda_rca32_u_rca62_fa45_y2 = h_s_dadda_rca32_u_rca62_out[45];
  assign h_s_dadda_rca32_u_rca62_fa46_y2 = h_s_dadda_rca32_u_rca62_out[46];
  assign h_s_dadda_rca32_u_rca62_fa47_y2 = h_s_dadda_rca32_u_rca62_out[47];
  assign h_s_dadda_rca32_u_rca62_fa48_y2 = h_s_dadda_rca32_u_rca62_out[48];
  assign h_s_dadda_rca32_u_rca62_fa49_y2 = h_s_dadda_rca32_u_rca62_out[49];
  assign h_s_dadda_rca32_u_rca62_fa50_y2 = h_s_dadda_rca32_u_rca62_out[50];
  assign h_s_dadda_rca32_u_rca62_fa51_y2 = h_s_dadda_rca32_u_rca62_out[51];
  assign h_s_dadda_rca32_u_rca62_fa52_y2 = h_s_dadda_rca32_u_rca62_out[52];
  assign h_s_dadda_rca32_u_rca62_fa53_y2 = h_s_dadda_rca32_u_rca62_out[53];
  assign h_s_dadda_rca32_u_rca62_fa54_y2 = h_s_dadda_rca32_u_rca62_out[54];
  assign h_s_dadda_rca32_u_rca62_fa55_y2 = h_s_dadda_rca32_u_rca62_out[55];
  assign h_s_dadda_rca32_u_rca62_fa56_y2 = h_s_dadda_rca32_u_rca62_out[56];
  assign h_s_dadda_rca32_u_rca62_fa57_y2 = h_s_dadda_rca32_u_rca62_out[57];
  assign h_s_dadda_rca32_u_rca62_fa58_y2 = h_s_dadda_rca32_u_rca62_out[58];
  assign h_s_dadda_rca32_u_rca62_fa59_y2 = h_s_dadda_rca32_u_rca62_out[59];
  assign h_s_dadda_rca32_u_rca62_fa60_y2 = h_s_dadda_rca32_u_rca62_out[60];
  assign h_s_dadda_rca32_u_rca62_fa61_y2 = h_s_dadda_rca32_u_rca62_out[61];
  assign h_s_dadda_rca32_u_rca62_fa61_y4 = h_s_dadda_rca32_u_rca62_out[62];
  xor_gate xor_gate_h_s_dadda_rca32_xor0_y0(constant_wire_1, h_s_dadda_rca32_u_rca62_fa61_y4, h_s_dadda_rca32_xor0_y0);

  assign out[0] = h_s_dadda_rca32_and_0_0_y0;
  assign out[1] = h_s_dadda_rca32_u_rca62_ha_y0;
  assign out[2] = h_s_dadda_rca32_u_rca62_fa1_y2;
  assign out[3] = h_s_dadda_rca32_u_rca62_fa2_y2;
  assign out[4] = h_s_dadda_rca32_u_rca62_fa3_y2;
  assign out[5] = h_s_dadda_rca32_u_rca62_fa4_y2;
  assign out[6] = h_s_dadda_rca32_u_rca62_fa5_y2;
  assign out[7] = h_s_dadda_rca32_u_rca62_fa6_y2;
  assign out[8] = h_s_dadda_rca32_u_rca62_fa7_y2;
  assign out[9] = h_s_dadda_rca32_u_rca62_fa8_y2;
  assign out[10] = h_s_dadda_rca32_u_rca62_fa9_y2;
  assign out[11] = h_s_dadda_rca32_u_rca62_fa10_y2;
  assign out[12] = h_s_dadda_rca32_u_rca62_fa11_y2;
  assign out[13] = h_s_dadda_rca32_u_rca62_fa12_y2;
  assign out[14] = h_s_dadda_rca32_u_rca62_fa13_y2;
  assign out[15] = h_s_dadda_rca32_u_rca62_fa14_y2;
  assign out[16] = h_s_dadda_rca32_u_rca62_fa15_y2;
  assign out[17] = h_s_dadda_rca32_u_rca62_fa16_y2;
  assign out[18] = h_s_dadda_rca32_u_rca62_fa17_y2;
  assign out[19] = h_s_dadda_rca32_u_rca62_fa18_y2;
  assign out[20] = h_s_dadda_rca32_u_rca62_fa19_y2;
  assign out[21] = h_s_dadda_rca32_u_rca62_fa20_y2;
  assign out[22] = h_s_dadda_rca32_u_rca62_fa21_y2;
  assign out[23] = h_s_dadda_rca32_u_rca62_fa22_y2;
  assign out[24] = h_s_dadda_rca32_u_rca62_fa23_y2;
  assign out[25] = h_s_dadda_rca32_u_rca62_fa24_y2;
  assign out[26] = h_s_dadda_rca32_u_rca62_fa25_y2;
  assign out[27] = h_s_dadda_rca32_u_rca62_fa26_y2;
  assign out[28] = h_s_dadda_rca32_u_rca62_fa27_y2;
  assign out[29] = h_s_dadda_rca32_u_rca62_fa28_y2;
  assign out[30] = h_s_dadda_rca32_u_rca62_fa29_y2;
  assign out[31] = h_s_dadda_rca32_u_rca62_fa30_y2;
  assign out[32] = h_s_dadda_rca32_u_rca62_fa31_y2;
  assign out[33] = h_s_dadda_rca32_u_rca62_fa32_y2;
  assign out[34] = h_s_dadda_rca32_u_rca62_fa33_y2;
  assign out[35] = h_s_dadda_rca32_u_rca62_fa34_y2;
  assign out[36] = h_s_dadda_rca32_u_rca62_fa35_y2;
  assign out[37] = h_s_dadda_rca32_u_rca62_fa36_y2;
  assign out[38] = h_s_dadda_rca32_u_rca62_fa37_y2;
  assign out[39] = h_s_dadda_rca32_u_rca62_fa38_y2;
  assign out[40] = h_s_dadda_rca32_u_rca62_fa39_y2;
  assign out[41] = h_s_dadda_rca32_u_rca62_fa40_y2;
  assign out[42] = h_s_dadda_rca32_u_rca62_fa41_y2;
  assign out[43] = h_s_dadda_rca32_u_rca62_fa42_y2;
  assign out[44] = h_s_dadda_rca32_u_rca62_fa43_y2;
  assign out[45] = h_s_dadda_rca32_u_rca62_fa44_y2;
  assign out[46] = h_s_dadda_rca32_u_rca62_fa45_y2;
  assign out[47] = h_s_dadda_rca32_u_rca62_fa46_y2;
  assign out[48] = h_s_dadda_rca32_u_rca62_fa47_y2;
  assign out[49] = h_s_dadda_rca32_u_rca62_fa48_y2;
  assign out[50] = h_s_dadda_rca32_u_rca62_fa49_y2;
  assign out[51] = h_s_dadda_rca32_u_rca62_fa50_y2;
  assign out[52] = h_s_dadda_rca32_u_rca62_fa51_y2;
  assign out[53] = h_s_dadda_rca32_u_rca62_fa52_y2;
  assign out[54] = h_s_dadda_rca32_u_rca62_fa53_y2;
  assign out[55] = h_s_dadda_rca32_u_rca62_fa54_y2;
  assign out[56] = h_s_dadda_rca32_u_rca62_fa55_y2;
  assign out[57] = h_s_dadda_rca32_u_rca62_fa56_y2;
  assign out[58] = h_s_dadda_rca32_u_rca62_fa57_y2;
  assign out[59] = h_s_dadda_rca32_u_rca62_fa58_y2;
  assign out[60] = h_s_dadda_rca32_u_rca62_fa59_y2;
  assign out[61] = h_s_dadda_rca32_u_rca62_fa60_y2;
  assign out[62] = h_s_dadda_rca32_u_rca62_fa61_y2;
  assign out[63] = h_s_dadda_rca32_xor0_y0;
endmodule