module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module u_rca46(input [45:0] a, input [45:0] b, output [46:0] u_rca46_out);
  wire [0:0] u_rca46_ha_xor0;
  wire [0:0] u_rca46_ha_and0;
  wire [0:0] u_rca46_fa1_xor1;
  wire [0:0] u_rca46_fa1_or0;
  wire [0:0] u_rca46_fa2_xor1;
  wire [0:0] u_rca46_fa2_or0;
  wire [0:0] u_rca46_fa3_xor1;
  wire [0:0] u_rca46_fa3_or0;
  wire [0:0] u_rca46_fa4_xor1;
  wire [0:0] u_rca46_fa4_or0;
  wire [0:0] u_rca46_fa5_xor1;
  wire [0:0] u_rca46_fa5_or0;
  wire [0:0] u_rca46_fa6_xor1;
  wire [0:0] u_rca46_fa6_or0;
  wire [0:0] u_rca46_fa7_xor1;
  wire [0:0] u_rca46_fa7_or0;
  wire [0:0] u_rca46_fa8_xor1;
  wire [0:0] u_rca46_fa8_or0;
  wire [0:0] u_rca46_fa9_xor1;
  wire [0:0] u_rca46_fa9_or0;
  wire [0:0] u_rca46_fa10_xor1;
  wire [0:0] u_rca46_fa10_or0;
  wire [0:0] u_rca46_fa11_xor1;
  wire [0:0] u_rca46_fa11_or0;
  wire [0:0] u_rca46_fa12_xor1;
  wire [0:0] u_rca46_fa12_or0;
  wire [0:0] u_rca46_fa13_xor1;
  wire [0:0] u_rca46_fa13_or0;
  wire [0:0] u_rca46_fa14_xor1;
  wire [0:0] u_rca46_fa14_or0;
  wire [0:0] u_rca46_fa15_xor1;
  wire [0:0] u_rca46_fa15_or0;
  wire [0:0] u_rca46_fa16_xor1;
  wire [0:0] u_rca46_fa16_or0;
  wire [0:0] u_rca46_fa17_xor1;
  wire [0:0] u_rca46_fa17_or0;
  wire [0:0] u_rca46_fa18_xor1;
  wire [0:0] u_rca46_fa18_or0;
  wire [0:0] u_rca46_fa19_xor1;
  wire [0:0] u_rca46_fa19_or0;
  wire [0:0] u_rca46_fa20_xor1;
  wire [0:0] u_rca46_fa20_or0;
  wire [0:0] u_rca46_fa21_xor1;
  wire [0:0] u_rca46_fa21_or0;
  wire [0:0] u_rca46_fa22_xor1;
  wire [0:0] u_rca46_fa22_or0;
  wire [0:0] u_rca46_fa23_xor1;
  wire [0:0] u_rca46_fa23_or0;
  wire [0:0] u_rca46_fa24_xor1;
  wire [0:0] u_rca46_fa24_or0;
  wire [0:0] u_rca46_fa25_xor1;
  wire [0:0] u_rca46_fa25_or0;
  wire [0:0] u_rca46_fa26_xor1;
  wire [0:0] u_rca46_fa26_or0;
  wire [0:0] u_rca46_fa27_xor1;
  wire [0:0] u_rca46_fa27_or0;
  wire [0:0] u_rca46_fa28_xor1;
  wire [0:0] u_rca46_fa28_or0;
  wire [0:0] u_rca46_fa29_xor1;
  wire [0:0] u_rca46_fa29_or0;
  wire [0:0] u_rca46_fa30_xor1;
  wire [0:0] u_rca46_fa30_or0;
  wire [0:0] u_rca46_fa31_xor1;
  wire [0:0] u_rca46_fa31_or0;
  wire [0:0] u_rca46_fa32_xor1;
  wire [0:0] u_rca46_fa32_or0;
  wire [0:0] u_rca46_fa33_xor1;
  wire [0:0] u_rca46_fa33_or0;
  wire [0:0] u_rca46_fa34_xor1;
  wire [0:0] u_rca46_fa34_or0;
  wire [0:0] u_rca46_fa35_xor1;
  wire [0:0] u_rca46_fa35_or0;
  wire [0:0] u_rca46_fa36_xor1;
  wire [0:0] u_rca46_fa36_or0;
  wire [0:0] u_rca46_fa37_xor1;
  wire [0:0] u_rca46_fa37_or0;
  wire [0:0] u_rca46_fa38_xor1;
  wire [0:0] u_rca46_fa38_or0;
  wire [0:0] u_rca46_fa39_xor1;
  wire [0:0] u_rca46_fa39_or0;
  wire [0:0] u_rca46_fa40_xor1;
  wire [0:0] u_rca46_fa40_or0;
  wire [0:0] u_rca46_fa41_xor1;
  wire [0:0] u_rca46_fa41_or0;
  wire [0:0] u_rca46_fa42_xor1;
  wire [0:0] u_rca46_fa42_or0;
  wire [0:0] u_rca46_fa43_xor1;
  wire [0:0] u_rca46_fa43_or0;
  wire [0:0] u_rca46_fa44_xor1;
  wire [0:0] u_rca46_fa44_or0;
  wire [0:0] u_rca46_fa45_xor1;
  wire [0:0] u_rca46_fa45_or0;

  ha ha_u_rca46_ha_out(.a(a[0]), .b(b[0]), .ha_xor0(u_rca46_ha_xor0), .ha_and0(u_rca46_ha_and0));
  fa fa_u_rca46_fa1_out(.a(a[1]), .b(b[1]), .cin(u_rca46_ha_and0[0]), .fa_xor1(u_rca46_fa1_xor1), .fa_or0(u_rca46_fa1_or0));
  fa fa_u_rca46_fa2_out(.a(a[2]), .b(b[2]), .cin(u_rca46_fa1_or0[0]), .fa_xor1(u_rca46_fa2_xor1), .fa_or0(u_rca46_fa2_or0));
  fa fa_u_rca46_fa3_out(.a(a[3]), .b(b[3]), .cin(u_rca46_fa2_or0[0]), .fa_xor1(u_rca46_fa3_xor1), .fa_or0(u_rca46_fa3_or0));
  fa fa_u_rca46_fa4_out(.a(a[4]), .b(b[4]), .cin(u_rca46_fa3_or0[0]), .fa_xor1(u_rca46_fa4_xor1), .fa_or0(u_rca46_fa4_or0));
  fa fa_u_rca46_fa5_out(.a(a[5]), .b(b[5]), .cin(u_rca46_fa4_or0[0]), .fa_xor1(u_rca46_fa5_xor1), .fa_or0(u_rca46_fa5_or0));
  fa fa_u_rca46_fa6_out(.a(a[6]), .b(b[6]), .cin(u_rca46_fa5_or0[0]), .fa_xor1(u_rca46_fa6_xor1), .fa_or0(u_rca46_fa6_or0));
  fa fa_u_rca46_fa7_out(.a(a[7]), .b(b[7]), .cin(u_rca46_fa6_or0[0]), .fa_xor1(u_rca46_fa7_xor1), .fa_or0(u_rca46_fa7_or0));
  fa fa_u_rca46_fa8_out(.a(a[8]), .b(b[8]), .cin(u_rca46_fa7_or0[0]), .fa_xor1(u_rca46_fa8_xor1), .fa_or0(u_rca46_fa8_or0));
  fa fa_u_rca46_fa9_out(.a(a[9]), .b(b[9]), .cin(u_rca46_fa8_or0[0]), .fa_xor1(u_rca46_fa9_xor1), .fa_or0(u_rca46_fa9_or0));
  fa fa_u_rca46_fa10_out(.a(a[10]), .b(b[10]), .cin(u_rca46_fa9_or0[0]), .fa_xor1(u_rca46_fa10_xor1), .fa_or0(u_rca46_fa10_or0));
  fa fa_u_rca46_fa11_out(.a(a[11]), .b(b[11]), .cin(u_rca46_fa10_or0[0]), .fa_xor1(u_rca46_fa11_xor1), .fa_or0(u_rca46_fa11_or0));
  fa fa_u_rca46_fa12_out(.a(a[12]), .b(b[12]), .cin(u_rca46_fa11_or0[0]), .fa_xor1(u_rca46_fa12_xor1), .fa_or0(u_rca46_fa12_or0));
  fa fa_u_rca46_fa13_out(.a(a[13]), .b(b[13]), .cin(u_rca46_fa12_or0[0]), .fa_xor1(u_rca46_fa13_xor1), .fa_or0(u_rca46_fa13_or0));
  fa fa_u_rca46_fa14_out(.a(a[14]), .b(b[14]), .cin(u_rca46_fa13_or0[0]), .fa_xor1(u_rca46_fa14_xor1), .fa_or0(u_rca46_fa14_or0));
  fa fa_u_rca46_fa15_out(.a(a[15]), .b(b[15]), .cin(u_rca46_fa14_or0[0]), .fa_xor1(u_rca46_fa15_xor1), .fa_or0(u_rca46_fa15_or0));
  fa fa_u_rca46_fa16_out(.a(a[16]), .b(b[16]), .cin(u_rca46_fa15_or0[0]), .fa_xor1(u_rca46_fa16_xor1), .fa_or0(u_rca46_fa16_or0));
  fa fa_u_rca46_fa17_out(.a(a[17]), .b(b[17]), .cin(u_rca46_fa16_or0[0]), .fa_xor1(u_rca46_fa17_xor1), .fa_or0(u_rca46_fa17_or0));
  fa fa_u_rca46_fa18_out(.a(a[18]), .b(b[18]), .cin(u_rca46_fa17_or0[0]), .fa_xor1(u_rca46_fa18_xor1), .fa_or0(u_rca46_fa18_or0));
  fa fa_u_rca46_fa19_out(.a(a[19]), .b(b[19]), .cin(u_rca46_fa18_or0[0]), .fa_xor1(u_rca46_fa19_xor1), .fa_or0(u_rca46_fa19_or0));
  fa fa_u_rca46_fa20_out(.a(a[20]), .b(b[20]), .cin(u_rca46_fa19_or0[0]), .fa_xor1(u_rca46_fa20_xor1), .fa_or0(u_rca46_fa20_or0));
  fa fa_u_rca46_fa21_out(.a(a[21]), .b(b[21]), .cin(u_rca46_fa20_or0[0]), .fa_xor1(u_rca46_fa21_xor1), .fa_or0(u_rca46_fa21_or0));
  fa fa_u_rca46_fa22_out(.a(a[22]), .b(b[22]), .cin(u_rca46_fa21_or0[0]), .fa_xor1(u_rca46_fa22_xor1), .fa_or0(u_rca46_fa22_or0));
  fa fa_u_rca46_fa23_out(.a(a[23]), .b(b[23]), .cin(u_rca46_fa22_or0[0]), .fa_xor1(u_rca46_fa23_xor1), .fa_or0(u_rca46_fa23_or0));
  fa fa_u_rca46_fa24_out(.a(a[24]), .b(b[24]), .cin(u_rca46_fa23_or0[0]), .fa_xor1(u_rca46_fa24_xor1), .fa_or0(u_rca46_fa24_or0));
  fa fa_u_rca46_fa25_out(.a(a[25]), .b(b[25]), .cin(u_rca46_fa24_or0[0]), .fa_xor1(u_rca46_fa25_xor1), .fa_or0(u_rca46_fa25_or0));
  fa fa_u_rca46_fa26_out(.a(a[26]), .b(b[26]), .cin(u_rca46_fa25_or0[0]), .fa_xor1(u_rca46_fa26_xor1), .fa_or0(u_rca46_fa26_or0));
  fa fa_u_rca46_fa27_out(.a(a[27]), .b(b[27]), .cin(u_rca46_fa26_or0[0]), .fa_xor1(u_rca46_fa27_xor1), .fa_or0(u_rca46_fa27_or0));
  fa fa_u_rca46_fa28_out(.a(a[28]), .b(b[28]), .cin(u_rca46_fa27_or0[0]), .fa_xor1(u_rca46_fa28_xor1), .fa_or0(u_rca46_fa28_or0));
  fa fa_u_rca46_fa29_out(.a(a[29]), .b(b[29]), .cin(u_rca46_fa28_or0[0]), .fa_xor1(u_rca46_fa29_xor1), .fa_or0(u_rca46_fa29_or0));
  fa fa_u_rca46_fa30_out(.a(a[30]), .b(b[30]), .cin(u_rca46_fa29_or0[0]), .fa_xor1(u_rca46_fa30_xor1), .fa_or0(u_rca46_fa30_or0));
  fa fa_u_rca46_fa31_out(.a(a[31]), .b(b[31]), .cin(u_rca46_fa30_or0[0]), .fa_xor1(u_rca46_fa31_xor1), .fa_or0(u_rca46_fa31_or0));
  fa fa_u_rca46_fa32_out(.a(a[32]), .b(b[32]), .cin(u_rca46_fa31_or0[0]), .fa_xor1(u_rca46_fa32_xor1), .fa_or0(u_rca46_fa32_or0));
  fa fa_u_rca46_fa33_out(.a(a[33]), .b(b[33]), .cin(u_rca46_fa32_or0[0]), .fa_xor1(u_rca46_fa33_xor1), .fa_or0(u_rca46_fa33_or0));
  fa fa_u_rca46_fa34_out(.a(a[34]), .b(b[34]), .cin(u_rca46_fa33_or0[0]), .fa_xor1(u_rca46_fa34_xor1), .fa_or0(u_rca46_fa34_or0));
  fa fa_u_rca46_fa35_out(.a(a[35]), .b(b[35]), .cin(u_rca46_fa34_or0[0]), .fa_xor1(u_rca46_fa35_xor1), .fa_or0(u_rca46_fa35_or0));
  fa fa_u_rca46_fa36_out(.a(a[36]), .b(b[36]), .cin(u_rca46_fa35_or0[0]), .fa_xor1(u_rca46_fa36_xor1), .fa_or0(u_rca46_fa36_or0));
  fa fa_u_rca46_fa37_out(.a(a[37]), .b(b[37]), .cin(u_rca46_fa36_or0[0]), .fa_xor1(u_rca46_fa37_xor1), .fa_or0(u_rca46_fa37_or0));
  fa fa_u_rca46_fa38_out(.a(a[38]), .b(b[38]), .cin(u_rca46_fa37_or0[0]), .fa_xor1(u_rca46_fa38_xor1), .fa_or0(u_rca46_fa38_or0));
  fa fa_u_rca46_fa39_out(.a(a[39]), .b(b[39]), .cin(u_rca46_fa38_or0[0]), .fa_xor1(u_rca46_fa39_xor1), .fa_or0(u_rca46_fa39_or0));
  fa fa_u_rca46_fa40_out(.a(a[40]), .b(b[40]), .cin(u_rca46_fa39_or0[0]), .fa_xor1(u_rca46_fa40_xor1), .fa_or0(u_rca46_fa40_or0));
  fa fa_u_rca46_fa41_out(.a(a[41]), .b(b[41]), .cin(u_rca46_fa40_or0[0]), .fa_xor1(u_rca46_fa41_xor1), .fa_or0(u_rca46_fa41_or0));
  fa fa_u_rca46_fa42_out(.a(a[42]), .b(b[42]), .cin(u_rca46_fa41_or0[0]), .fa_xor1(u_rca46_fa42_xor1), .fa_or0(u_rca46_fa42_or0));
  fa fa_u_rca46_fa43_out(.a(a[43]), .b(b[43]), .cin(u_rca46_fa42_or0[0]), .fa_xor1(u_rca46_fa43_xor1), .fa_or0(u_rca46_fa43_or0));
  fa fa_u_rca46_fa44_out(.a(a[44]), .b(b[44]), .cin(u_rca46_fa43_or0[0]), .fa_xor1(u_rca46_fa44_xor1), .fa_or0(u_rca46_fa44_or0));
  fa fa_u_rca46_fa45_out(.a(a[45]), .b(b[45]), .cin(u_rca46_fa44_or0[0]), .fa_xor1(u_rca46_fa45_xor1), .fa_or0(u_rca46_fa45_or0));

  assign u_rca46_out[0] = u_rca46_ha_xor0[0];
  assign u_rca46_out[1] = u_rca46_fa1_xor1[0];
  assign u_rca46_out[2] = u_rca46_fa2_xor1[0];
  assign u_rca46_out[3] = u_rca46_fa3_xor1[0];
  assign u_rca46_out[4] = u_rca46_fa4_xor1[0];
  assign u_rca46_out[5] = u_rca46_fa5_xor1[0];
  assign u_rca46_out[6] = u_rca46_fa6_xor1[0];
  assign u_rca46_out[7] = u_rca46_fa7_xor1[0];
  assign u_rca46_out[8] = u_rca46_fa8_xor1[0];
  assign u_rca46_out[9] = u_rca46_fa9_xor1[0];
  assign u_rca46_out[10] = u_rca46_fa10_xor1[0];
  assign u_rca46_out[11] = u_rca46_fa11_xor1[0];
  assign u_rca46_out[12] = u_rca46_fa12_xor1[0];
  assign u_rca46_out[13] = u_rca46_fa13_xor1[0];
  assign u_rca46_out[14] = u_rca46_fa14_xor1[0];
  assign u_rca46_out[15] = u_rca46_fa15_xor1[0];
  assign u_rca46_out[16] = u_rca46_fa16_xor1[0];
  assign u_rca46_out[17] = u_rca46_fa17_xor1[0];
  assign u_rca46_out[18] = u_rca46_fa18_xor1[0];
  assign u_rca46_out[19] = u_rca46_fa19_xor1[0];
  assign u_rca46_out[20] = u_rca46_fa20_xor1[0];
  assign u_rca46_out[21] = u_rca46_fa21_xor1[0];
  assign u_rca46_out[22] = u_rca46_fa22_xor1[0];
  assign u_rca46_out[23] = u_rca46_fa23_xor1[0];
  assign u_rca46_out[24] = u_rca46_fa24_xor1[0];
  assign u_rca46_out[25] = u_rca46_fa25_xor1[0];
  assign u_rca46_out[26] = u_rca46_fa26_xor1[0];
  assign u_rca46_out[27] = u_rca46_fa27_xor1[0];
  assign u_rca46_out[28] = u_rca46_fa28_xor1[0];
  assign u_rca46_out[29] = u_rca46_fa29_xor1[0];
  assign u_rca46_out[30] = u_rca46_fa30_xor1[0];
  assign u_rca46_out[31] = u_rca46_fa31_xor1[0];
  assign u_rca46_out[32] = u_rca46_fa32_xor1[0];
  assign u_rca46_out[33] = u_rca46_fa33_xor1[0];
  assign u_rca46_out[34] = u_rca46_fa34_xor1[0];
  assign u_rca46_out[35] = u_rca46_fa35_xor1[0];
  assign u_rca46_out[36] = u_rca46_fa36_xor1[0];
  assign u_rca46_out[37] = u_rca46_fa37_xor1[0];
  assign u_rca46_out[38] = u_rca46_fa38_xor1[0];
  assign u_rca46_out[39] = u_rca46_fa39_xor1[0];
  assign u_rca46_out[40] = u_rca46_fa40_xor1[0];
  assign u_rca46_out[41] = u_rca46_fa41_xor1[0];
  assign u_rca46_out[42] = u_rca46_fa42_xor1[0];
  assign u_rca46_out[43] = u_rca46_fa43_xor1[0];
  assign u_rca46_out[44] = u_rca46_fa44_xor1[0];
  assign u_rca46_out[45] = u_rca46_fa45_xor1[0];
  assign u_rca46_out[46] = u_rca46_fa45_or0[0];
endmodule

module s_wallace_rca24(input [23:0] a, input [23:0] b, output [47:0] s_wallace_rca24_out);
  wire [0:0] s_wallace_rca24_and_2_0;
  wire [0:0] s_wallace_rca24_and_1_1;
  wire [0:0] s_wallace_rca24_ha0_xor0;
  wire [0:0] s_wallace_rca24_ha0_and0;
  wire [0:0] s_wallace_rca24_and_3_0;
  wire [0:0] s_wallace_rca24_and_2_1;
  wire [0:0] s_wallace_rca24_fa0_xor1;
  wire [0:0] s_wallace_rca24_fa0_or0;
  wire [0:0] s_wallace_rca24_and_4_0;
  wire [0:0] s_wallace_rca24_and_3_1;
  wire [0:0] s_wallace_rca24_fa1_xor1;
  wire [0:0] s_wallace_rca24_fa1_or0;
  wire [0:0] s_wallace_rca24_and_5_0;
  wire [0:0] s_wallace_rca24_and_4_1;
  wire [0:0] s_wallace_rca24_fa2_xor1;
  wire [0:0] s_wallace_rca24_fa2_or0;
  wire [0:0] s_wallace_rca24_and_6_0;
  wire [0:0] s_wallace_rca24_and_5_1;
  wire [0:0] s_wallace_rca24_fa3_xor1;
  wire [0:0] s_wallace_rca24_fa3_or0;
  wire [0:0] s_wallace_rca24_and_7_0;
  wire [0:0] s_wallace_rca24_and_6_1;
  wire [0:0] s_wallace_rca24_fa4_xor1;
  wire [0:0] s_wallace_rca24_fa4_or0;
  wire [0:0] s_wallace_rca24_and_8_0;
  wire [0:0] s_wallace_rca24_and_7_1;
  wire [0:0] s_wallace_rca24_fa5_xor1;
  wire [0:0] s_wallace_rca24_fa5_or0;
  wire [0:0] s_wallace_rca24_and_9_0;
  wire [0:0] s_wallace_rca24_and_8_1;
  wire [0:0] s_wallace_rca24_fa6_xor1;
  wire [0:0] s_wallace_rca24_fa6_or0;
  wire [0:0] s_wallace_rca24_and_10_0;
  wire [0:0] s_wallace_rca24_and_9_1;
  wire [0:0] s_wallace_rca24_fa7_xor1;
  wire [0:0] s_wallace_rca24_fa7_or0;
  wire [0:0] s_wallace_rca24_and_11_0;
  wire [0:0] s_wallace_rca24_and_10_1;
  wire [0:0] s_wallace_rca24_fa8_xor1;
  wire [0:0] s_wallace_rca24_fa8_or0;
  wire [0:0] s_wallace_rca24_and_12_0;
  wire [0:0] s_wallace_rca24_and_11_1;
  wire [0:0] s_wallace_rca24_fa9_xor1;
  wire [0:0] s_wallace_rca24_fa9_or0;
  wire [0:0] s_wallace_rca24_and_13_0;
  wire [0:0] s_wallace_rca24_and_12_1;
  wire [0:0] s_wallace_rca24_fa10_xor1;
  wire [0:0] s_wallace_rca24_fa10_or0;
  wire [0:0] s_wallace_rca24_and_14_0;
  wire [0:0] s_wallace_rca24_and_13_1;
  wire [0:0] s_wallace_rca24_fa11_xor1;
  wire [0:0] s_wallace_rca24_fa11_or0;
  wire [0:0] s_wallace_rca24_and_15_0;
  wire [0:0] s_wallace_rca24_and_14_1;
  wire [0:0] s_wallace_rca24_fa12_xor1;
  wire [0:0] s_wallace_rca24_fa12_or0;
  wire [0:0] s_wallace_rca24_and_16_0;
  wire [0:0] s_wallace_rca24_and_15_1;
  wire [0:0] s_wallace_rca24_fa13_xor1;
  wire [0:0] s_wallace_rca24_fa13_or0;
  wire [0:0] s_wallace_rca24_and_17_0;
  wire [0:0] s_wallace_rca24_and_16_1;
  wire [0:0] s_wallace_rca24_fa14_xor1;
  wire [0:0] s_wallace_rca24_fa14_or0;
  wire [0:0] s_wallace_rca24_and_18_0;
  wire [0:0] s_wallace_rca24_and_17_1;
  wire [0:0] s_wallace_rca24_fa15_xor1;
  wire [0:0] s_wallace_rca24_fa15_or0;
  wire [0:0] s_wallace_rca24_and_19_0;
  wire [0:0] s_wallace_rca24_and_18_1;
  wire [0:0] s_wallace_rca24_fa16_xor1;
  wire [0:0] s_wallace_rca24_fa16_or0;
  wire [0:0] s_wallace_rca24_and_20_0;
  wire [0:0] s_wallace_rca24_and_19_1;
  wire [0:0] s_wallace_rca24_fa17_xor1;
  wire [0:0] s_wallace_rca24_fa17_or0;
  wire [0:0] s_wallace_rca24_and_21_0;
  wire [0:0] s_wallace_rca24_and_20_1;
  wire [0:0] s_wallace_rca24_fa18_xor1;
  wire [0:0] s_wallace_rca24_fa18_or0;
  wire [0:0] s_wallace_rca24_and_22_0;
  wire [0:0] s_wallace_rca24_and_21_1;
  wire [0:0] s_wallace_rca24_fa19_xor1;
  wire [0:0] s_wallace_rca24_fa19_or0;
  wire [0:0] s_wallace_rca24_nand_23_0;
  wire [0:0] s_wallace_rca24_and_22_1;
  wire [0:0] s_wallace_rca24_fa20_xor1;
  wire [0:0] s_wallace_rca24_fa20_or0;
  wire [0:0] s_wallace_rca24_nand_23_1;
  wire [0:0] s_wallace_rca24_fa21_xor1;
  wire [0:0] s_wallace_rca24_fa21_or0;
  wire [0:0] s_wallace_rca24_nand_23_2;
  wire [0:0] s_wallace_rca24_and_22_3;
  wire [0:0] s_wallace_rca24_fa22_xor1;
  wire [0:0] s_wallace_rca24_fa22_or0;
  wire [0:0] s_wallace_rca24_nand_23_3;
  wire [0:0] s_wallace_rca24_and_22_4;
  wire [0:0] s_wallace_rca24_fa23_xor1;
  wire [0:0] s_wallace_rca24_fa23_or0;
  wire [0:0] s_wallace_rca24_nand_23_4;
  wire [0:0] s_wallace_rca24_and_22_5;
  wire [0:0] s_wallace_rca24_fa24_xor1;
  wire [0:0] s_wallace_rca24_fa24_or0;
  wire [0:0] s_wallace_rca24_nand_23_5;
  wire [0:0] s_wallace_rca24_and_22_6;
  wire [0:0] s_wallace_rca24_fa25_xor1;
  wire [0:0] s_wallace_rca24_fa25_or0;
  wire [0:0] s_wallace_rca24_nand_23_6;
  wire [0:0] s_wallace_rca24_and_22_7;
  wire [0:0] s_wallace_rca24_fa26_xor1;
  wire [0:0] s_wallace_rca24_fa26_or0;
  wire [0:0] s_wallace_rca24_nand_23_7;
  wire [0:0] s_wallace_rca24_and_22_8;
  wire [0:0] s_wallace_rca24_fa27_xor1;
  wire [0:0] s_wallace_rca24_fa27_or0;
  wire [0:0] s_wallace_rca24_nand_23_8;
  wire [0:0] s_wallace_rca24_and_22_9;
  wire [0:0] s_wallace_rca24_fa28_xor1;
  wire [0:0] s_wallace_rca24_fa28_or0;
  wire [0:0] s_wallace_rca24_nand_23_9;
  wire [0:0] s_wallace_rca24_and_22_10;
  wire [0:0] s_wallace_rca24_fa29_xor1;
  wire [0:0] s_wallace_rca24_fa29_or0;
  wire [0:0] s_wallace_rca24_nand_23_10;
  wire [0:0] s_wallace_rca24_and_22_11;
  wire [0:0] s_wallace_rca24_fa30_xor1;
  wire [0:0] s_wallace_rca24_fa30_or0;
  wire [0:0] s_wallace_rca24_nand_23_11;
  wire [0:0] s_wallace_rca24_and_22_12;
  wire [0:0] s_wallace_rca24_fa31_xor1;
  wire [0:0] s_wallace_rca24_fa31_or0;
  wire [0:0] s_wallace_rca24_nand_23_12;
  wire [0:0] s_wallace_rca24_and_22_13;
  wire [0:0] s_wallace_rca24_fa32_xor1;
  wire [0:0] s_wallace_rca24_fa32_or0;
  wire [0:0] s_wallace_rca24_nand_23_13;
  wire [0:0] s_wallace_rca24_and_22_14;
  wire [0:0] s_wallace_rca24_fa33_xor1;
  wire [0:0] s_wallace_rca24_fa33_or0;
  wire [0:0] s_wallace_rca24_nand_23_14;
  wire [0:0] s_wallace_rca24_and_22_15;
  wire [0:0] s_wallace_rca24_fa34_xor1;
  wire [0:0] s_wallace_rca24_fa34_or0;
  wire [0:0] s_wallace_rca24_nand_23_15;
  wire [0:0] s_wallace_rca24_and_22_16;
  wire [0:0] s_wallace_rca24_fa35_xor1;
  wire [0:0] s_wallace_rca24_fa35_or0;
  wire [0:0] s_wallace_rca24_nand_23_16;
  wire [0:0] s_wallace_rca24_and_22_17;
  wire [0:0] s_wallace_rca24_fa36_xor1;
  wire [0:0] s_wallace_rca24_fa36_or0;
  wire [0:0] s_wallace_rca24_nand_23_17;
  wire [0:0] s_wallace_rca24_and_22_18;
  wire [0:0] s_wallace_rca24_fa37_xor1;
  wire [0:0] s_wallace_rca24_fa37_or0;
  wire [0:0] s_wallace_rca24_nand_23_18;
  wire [0:0] s_wallace_rca24_and_22_19;
  wire [0:0] s_wallace_rca24_fa38_xor1;
  wire [0:0] s_wallace_rca24_fa38_or0;
  wire [0:0] s_wallace_rca24_nand_23_19;
  wire [0:0] s_wallace_rca24_and_22_20;
  wire [0:0] s_wallace_rca24_fa39_xor1;
  wire [0:0] s_wallace_rca24_fa39_or0;
  wire [0:0] s_wallace_rca24_nand_23_20;
  wire [0:0] s_wallace_rca24_and_22_21;
  wire [0:0] s_wallace_rca24_fa40_xor1;
  wire [0:0] s_wallace_rca24_fa40_or0;
  wire [0:0] s_wallace_rca24_nand_23_21;
  wire [0:0] s_wallace_rca24_and_22_22;
  wire [0:0] s_wallace_rca24_fa41_xor1;
  wire [0:0] s_wallace_rca24_fa41_or0;
  wire [0:0] s_wallace_rca24_and_1_2;
  wire [0:0] s_wallace_rca24_and_0_3;
  wire [0:0] s_wallace_rca24_ha1_xor0;
  wire [0:0] s_wallace_rca24_ha1_and0;
  wire [0:0] s_wallace_rca24_and_2_2;
  wire [0:0] s_wallace_rca24_and_1_3;
  wire [0:0] s_wallace_rca24_fa42_xor1;
  wire [0:0] s_wallace_rca24_fa42_or0;
  wire [0:0] s_wallace_rca24_and_3_2;
  wire [0:0] s_wallace_rca24_and_2_3;
  wire [0:0] s_wallace_rca24_fa43_xor1;
  wire [0:0] s_wallace_rca24_fa43_or0;
  wire [0:0] s_wallace_rca24_and_4_2;
  wire [0:0] s_wallace_rca24_and_3_3;
  wire [0:0] s_wallace_rca24_fa44_xor1;
  wire [0:0] s_wallace_rca24_fa44_or0;
  wire [0:0] s_wallace_rca24_and_5_2;
  wire [0:0] s_wallace_rca24_and_4_3;
  wire [0:0] s_wallace_rca24_fa45_xor1;
  wire [0:0] s_wallace_rca24_fa45_or0;
  wire [0:0] s_wallace_rca24_and_6_2;
  wire [0:0] s_wallace_rca24_and_5_3;
  wire [0:0] s_wallace_rca24_fa46_xor1;
  wire [0:0] s_wallace_rca24_fa46_or0;
  wire [0:0] s_wallace_rca24_and_7_2;
  wire [0:0] s_wallace_rca24_and_6_3;
  wire [0:0] s_wallace_rca24_fa47_xor1;
  wire [0:0] s_wallace_rca24_fa47_or0;
  wire [0:0] s_wallace_rca24_and_8_2;
  wire [0:0] s_wallace_rca24_and_7_3;
  wire [0:0] s_wallace_rca24_fa48_xor1;
  wire [0:0] s_wallace_rca24_fa48_or0;
  wire [0:0] s_wallace_rca24_and_9_2;
  wire [0:0] s_wallace_rca24_and_8_3;
  wire [0:0] s_wallace_rca24_fa49_xor1;
  wire [0:0] s_wallace_rca24_fa49_or0;
  wire [0:0] s_wallace_rca24_and_10_2;
  wire [0:0] s_wallace_rca24_and_9_3;
  wire [0:0] s_wallace_rca24_fa50_xor1;
  wire [0:0] s_wallace_rca24_fa50_or0;
  wire [0:0] s_wallace_rca24_and_11_2;
  wire [0:0] s_wallace_rca24_and_10_3;
  wire [0:0] s_wallace_rca24_fa51_xor1;
  wire [0:0] s_wallace_rca24_fa51_or0;
  wire [0:0] s_wallace_rca24_and_12_2;
  wire [0:0] s_wallace_rca24_and_11_3;
  wire [0:0] s_wallace_rca24_fa52_xor1;
  wire [0:0] s_wallace_rca24_fa52_or0;
  wire [0:0] s_wallace_rca24_and_13_2;
  wire [0:0] s_wallace_rca24_and_12_3;
  wire [0:0] s_wallace_rca24_fa53_xor1;
  wire [0:0] s_wallace_rca24_fa53_or0;
  wire [0:0] s_wallace_rca24_and_14_2;
  wire [0:0] s_wallace_rca24_and_13_3;
  wire [0:0] s_wallace_rca24_fa54_xor1;
  wire [0:0] s_wallace_rca24_fa54_or0;
  wire [0:0] s_wallace_rca24_and_15_2;
  wire [0:0] s_wallace_rca24_and_14_3;
  wire [0:0] s_wallace_rca24_fa55_xor1;
  wire [0:0] s_wallace_rca24_fa55_or0;
  wire [0:0] s_wallace_rca24_and_16_2;
  wire [0:0] s_wallace_rca24_and_15_3;
  wire [0:0] s_wallace_rca24_fa56_xor1;
  wire [0:0] s_wallace_rca24_fa56_or0;
  wire [0:0] s_wallace_rca24_and_17_2;
  wire [0:0] s_wallace_rca24_and_16_3;
  wire [0:0] s_wallace_rca24_fa57_xor1;
  wire [0:0] s_wallace_rca24_fa57_or0;
  wire [0:0] s_wallace_rca24_and_18_2;
  wire [0:0] s_wallace_rca24_and_17_3;
  wire [0:0] s_wallace_rca24_fa58_xor1;
  wire [0:0] s_wallace_rca24_fa58_or0;
  wire [0:0] s_wallace_rca24_and_19_2;
  wire [0:0] s_wallace_rca24_and_18_3;
  wire [0:0] s_wallace_rca24_fa59_xor1;
  wire [0:0] s_wallace_rca24_fa59_or0;
  wire [0:0] s_wallace_rca24_and_20_2;
  wire [0:0] s_wallace_rca24_and_19_3;
  wire [0:0] s_wallace_rca24_fa60_xor1;
  wire [0:0] s_wallace_rca24_fa60_or0;
  wire [0:0] s_wallace_rca24_and_21_2;
  wire [0:0] s_wallace_rca24_and_20_3;
  wire [0:0] s_wallace_rca24_fa61_xor1;
  wire [0:0] s_wallace_rca24_fa61_or0;
  wire [0:0] s_wallace_rca24_and_22_2;
  wire [0:0] s_wallace_rca24_and_21_3;
  wire [0:0] s_wallace_rca24_fa62_xor1;
  wire [0:0] s_wallace_rca24_fa62_or0;
  wire [0:0] s_wallace_rca24_and_21_4;
  wire [0:0] s_wallace_rca24_and_20_5;
  wire [0:0] s_wallace_rca24_fa63_xor1;
  wire [0:0] s_wallace_rca24_fa63_or0;
  wire [0:0] s_wallace_rca24_and_21_5;
  wire [0:0] s_wallace_rca24_and_20_6;
  wire [0:0] s_wallace_rca24_fa64_xor1;
  wire [0:0] s_wallace_rca24_fa64_or0;
  wire [0:0] s_wallace_rca24_and_21_6;
  wire [0:0] s_wallace_rca24_and_20_7;
  wire [0:0] s_wallace_rca24_fa65_xor1;
  wire [0:0] s_wallace_rca24_fa65_or0;
  wire [0:0] s_wallace_rca24_and_21_7;
  wire [0:0] s_wallace_rca24_and_20_8;
  wire [0:0] s_wallace_rca24_fa66_xor1;
  wire [0:0] s_wallace_rca24_fa66_or0;
  wire [0:0] s_wallace_rca24_and_21_8;
  wire [0:0] s_wallace_rca24_and_20_9;
  wire [0:0] s_wallace_rca24_fa67_xor1;
  wire [0:0] s_wallace_rca24_fa67_or0;
  wire [0:0] s_wallace_rca24_and_21_9;
  wire [0:0] s_wallace_rca24_and_20_10;
  wire [0:0] s_wallace_rca24_fa68_xor1;
  wire [0:0] s_wallace_rca24_fa68_or0;
  wire [0:0] s_wallace_rca24_and_21_10;
  wire [0:0] s_wallace_rca24_and_20_11;
  wire [0:0] s_wallace_rca24_fa69_xor1;
  wire [0:0] s_wallace_rca24_fa69_or0;
  wire [0:0] s_wallace_rca24_and_21_11;
  wire [0:0] s_wallace_rca24_and_20_12;
  wire [0:0] s_wallace_rca24_fa70_xor1;
  wire [0:0] s_wallace_rca24_fa70_or0;
  wire [0:0] s_wallace_rca24_and_21_12;
  wire [0:0] s_wallace_rca24_and_20_13;
  wire [0:0] s_wallace_rca24_fa71_xor1;
  wire [0:0] s_wallace_rca24_fa71_or0;
  wire [0:0] s_wallace_rca24_and_21_13;
  wire [0:0] s_wallace_rca24_and_20_14;
  wire [0:0] s_wallace_rca24_fa72_xor1;
  wire [0:0] s_wallace_rca24_fa72_or0;
  wire [0:0] s_wallace_rca24_and_21_14;
  wire [0:0] s_wallace_rca24_and_20_15;
  wire [0:0] s_wallace_rca24_fa73_xor1;
  wire [0:0] s_wallace_rca24_fa73_or0;
  wire [0:0] s_wallace_rca24_and_21_15;
  wire [0:0] s_wallace_rca24_and_20_16;
  wire [0:0] s_wallace_rca24_fa74_xor1;
  wire [0:0] s_wallace_rca24_fa74_or0;
  wire [0:0] s_wallace_rca24_and_21_16;
  wire [0:0] s_wallace_rca24_and_20_17;
  wire [0:0] s_wallace_rca24_fa75_xor1;
  wire [0:0] s_wallace_rca24_fa75_or0;
  wire [0:0] s_wallace_rca24_and_21_17;
  wire [0:0] s_wallace_rca24_and_20_18;
  wire [0:0] s_wallace_rca24_fa76_xor1;
  wire [0:0] s_wallace_rca24_fa76_or0;
  wire [0:0] s_wallace_rca24_and_21_18;
  wire [0:0] s_wallace_rca24_and_20_19;
  wire [0:0] s_wallace_rca24_fa77_xor1;
  wire [0:0] s_wallace_rca24_fa77_or0;
  wire [0:0] s_wallace_rca24_and_21_19;
  wire [0:0] s_wallace_rca24_and_20_20;
  wire [0:0] s_wallace_rca24_fa78_xor1;
  wire [0:0] s_wallace_rca24_fa78_or0;
  wire [0:0] s_wallace_rca24_and_21_20;
  wire [0:0] s_wallace_rca24_and_20_21;
  wire [0:0] s_wallace_rca24_fa79_xor1;
  wire [0:0] s_wallace_rca24_fa79_or0;
  wire [0:0] s_wallace_rca24_and_21_21;
  wire [0:0] s_wallace_rca24_and_20_22;
  wire [0:0] s_wallace_rca24_fa80_xor1;
  wire [0:0] s_wallace_rca24_fa80_or0;
  wire [0:0] s_wallace_rca24_and_21_22;
  wire [0:0] s_wallace_rca24_nand_20_23;
  wire [0:0] s_wallace_rca24_fa81_xor1;
  wire [0:0] s_wallace_rca24_fa81_or0;
  wire [0:0] s_wallace_rca24_and_0_4;
  wire [0:0] s_wallace_rca24_ha2_xor0;
  wire [0:0] s_wallace_rca24_ha2_and0;
  wire [0:0] s_wallace_rca24_and_1_4;
  wire [0:0] s_wallace_rca24_and_0_5;
  wire [0:0] s_wallace_rca24_fa82_xor1;
  wire [0:0] s_wallace_rca24_fa82_or0;
  wire [0:0] s_wallace_rca24_and_2_4;
  wire [0:0] s_wallace_rca24_and_1_5;
  wire [0:0] s_wallace_rca24_fa83_xor1;
  wire [0:0] s_wallace_rca24_fa83_or0;
  wire [0:0] s_wallace_rca24_and_3_4;
  wire [0:0] s_wallace_rca24_and_2_5;
  wire [0:0] s_wallace_rca24_fa84_xor1;
  wire [0:0] s_wallace_rca24_fa84_or0;
  wire [0:0] s_wallace_rca24_and_4_4;
  wire [0:0] s_wallace_rca24_and_3_5;
  wire [0:0] s_wallace_rca24_fa85_xor1;
  wire [0:0] s_wallace_rca24_fa85_or0;
  wire [0:0] s_wallace_rca24_and_5_4;
  wire [0:0] s_wallace_rca24_and_4_5;
  wire [0:0] s_wallace_rca24_fa86_xor1;
  wire [0:0] s_wallace_rca24_fa86_or0;
  wire [0:0] s_wallace_rca24_and_6_4;
  wire [0:0] s_wallace_rca24_and_5_5;
  wire [0:0] s_wallace_rca24_fa87_xor1;
  wire [0:0] s_wallace_rca24_fa87_or0;
  wire [0:0] s_wallace_rca24_and_7_4;
  wire [0:0] s_wallace_rca24_and_6_5;
  wire [0:0] s_wallace_rca24_fa88_xor1;
  wire [0:0] s_wallace_rca24_fa88_or0;
  wire [0:0] s_wallace_rca24_and_8_4;
  wire [0:0] s_wallace_rca24_and_7_5;
  wire [0:0] s_wallace_rca24_fa89_xor1;
  wire [0:0] s_wallace_rca24_fa89_or0;
  wire [0:0] s_wallace_rca24_and_9_4;
  wire [0:0] s_wallace_rca24_and_8_5;
  wire [0:0] s_wallace_rca24_fa90_xor1;
  wire [0:0] s_wallace_rca24_fa90_or0;
  wire [0:0] s_wallace_rca24_and_10_4;
  wire [0:0] s_wallace_rca24_and_9_5;
  wire [0:0] s_wallace_rca24_fa91_xor1;
  wire [0:0] s_wallace_rca24_fa91_or0;
  wire [0:0] s_wallace_rca24_and_11_4;
  wire [0:0] s_wallace_rca24_and_10_5;
  wire [0:0] s_wallace_rca24_fa92_xor1;
  wire [0:0] s_wallace_rca24_fa92_or0;
  wire [0:0] s_wallace_rca24_and_12_4;
  wire [0:0] s_wallace_rca24_and_11_5;
  wire [0:0] s_wallace_rca24_fa93_xor1;
  wire [0:0] s_wallace_rca24_fa93_or0;
  wire [0:0] s_wallace_rca24_and_13_4;
  wire [0:0] s_wallace_rca24_and_12_5;
  wire [0:0] s_wallace_rca24_fa94_xor1;
  wire [0:0] s_wallace_rca24_fa94_or0;
  wire [0:0] s_wallace_rca24_and_14_4;
  wire [0:0] s_wallace_rca24_and_13_5;
  wire [0:0] s_wallace_rca24_fa95_xor1;
  wire [0:0] s_wallace_rca24_fa95_or0;
  wire [0:0] s_wallace_rca24_and_15_4;
  wire [0:0] s_wallace_rca24_and_14_5;
  wire [0:0] s_wallace_rca24_fa96_xor1;
  wire [0:0] s_wallace_rca24_fa96_or0;
  wire [0:0] s_wallace_rca24_and_16_4;
  wire [0:0] s_wallace_rca24_and_15_5;
  wire [0:0] s_wallace_rca24_fa97_xor1;
  wire [0:0] s_wallace_rca24_fa97_or0;
  wire [0:0] s_wallace_rca24_and_17_4;
  wire [0:0] s_wallace_rca24_and_16_5;
  wire [0:0] s_wallace_rca24_fa98_xor1;
  wire [0:0] s_wallace_rca24_fa98_or0;
  wire [0:0] s_wallace_rca24_and_18_4;
  wire [0:0] s_wallace_rca24_and_17_5;
  wire [0:0] s_wallace_rca24_fa99_xor1;
  wire [0:0] s_wallace_rca24_fa99_or0;
  wire [0:0] s_wallace_rca24_and_19_4;
  wire [0:0] s_wallace_rca24_and_18_5;
  wire [0:0] s_wallace_rca24_fa100_xor1;
  wire [0:0] s_wallace_rca24_fa100_or0;
  wire [0:0] s_wallace_rca24_and_20_4;
  wire [0:0] s_wallace_rca24_and_19_5;
  wire [0:0] s_wallace_rca24_fa101_xor1;
  wire [0:0] s_wallace_rca24_fa101_or0;
  wire [0:0] s_wallace_rca24_and_19_6;
  wire [0:0] s_wallace_rca24_and_18_7;
  wire [0:0] s_wallace_rca24_fa102_xor1;
  wire [0:0] s_wallace_rca24_fa102_or0;
  wire [0:0] s_wallace_rca24_and_19_7;
  wire [0:0] s_wallace_rca24_and_18_8;
  wire [0:0] s_wallace_rca24_fa103_xor1;
  wire [0:0] s_wallace_rca24_fa103_or0;
  wire [0:0] s_wallace_rca24_and_19_8;
  wire [0:0] s_wallace_rca24_and_18_9;
  wire [0:0] s_wallace_rca24_fa104_xor1;
  wire [0:0] s_wallace_rca24_fa104_or0;
  wire [0:0] s_wallace_rca24_and_19_9;
  wire [0:0] s_wallace_rca24_and_18_10;
  wire [0:0] s_wallace_rca24_fa105_xor1;
  wire [0:0] s_wallace_rca24_fa105_or0;
  wire [0:0] s_wallace_rca24_and_19_10;
  wire [0:0] s_wallace_rca24_and_18_11;
  wire [0:0] s_wallace_rca24_fa106_xor1;
  wire [0:0] s_wallace_rca24_fa106_or0;
  wire [0:0] s_wallace_rca24_and_19_11;
  wire [0:0] s_wallace_rca24_and_18_12;
  wire [0:0] s_wallace_rca24_fa107_xor1;
  wire [0:0] s_wallace_rca24_fa107_or0;
  wire [0:0] s_wallace_rca24_and_19_12;
  wire [0:0] s_wallace_rca24_and_18_13;
  wire [0:0] s_wallace_rca24_fa108_xor1;
  wire [0:0] s_wallace_rca24_fa108_or0;
  wire [0:0] s_wallace_rca24_and_19_13;
  wire [0:0] s_wallace_rca24_and_18_14;
  wire [0:0] s_wallace_rca24_fa109_xor1;
  wire [0:0] s_wallace_rca24_fa109_or0;
  wire [0:0] s_wallace_rca24_and_19_14;
  wire [0:0] s_wallace_rca24_and_18_15;
  wire [0:0] s_wallace_rca24_fa110_xor1;
  wire [0:0] s_wallace_rca24_fa110_or0;
  wire [0:0] s_wallace_rca24_and_19_15;
  wire [0:0] s_wallace_rca24_and_18_16;
  wire [0:0] s_wallace_rca24_fa111_xor1;
  wire [0:0] s_wallace_rca24_fa111_or0;
  wire [0:0] s_wallace_rca24_and_19_16;
  wire [0:0] s_wallace_rca24_and_18_17;
  wire [0:0] s_wallace_rca24_fa112_xor1;
  wire [0:0] s_wallace_rca24_fa112_or0;
  wire [0:0] s_wallace_rca24_and_19_17;
  wire [0:0] s_wallace_rca24_and_18_18;
  wire [0:0] s_wallace_rca24_fa113_xor1;
  wire [0:0] s_wallace_rca24_fa113_or0;
  wire [0:0] s_wallace_rca24_and_19_18;
  wire [0:0] s_wallace_rca24_and_18_19;
  wire [0:0] s_wallace_rca24_fa114_xor1;
  wire [0:0] s_wallace_rca24_fa114_or0;
  wire [0:0] s_wallace_rca24_and_19_19;
  wire [0:0] s_wallace_rca24_and_18_20;
  wire [0:0] s_wallace_rca24_fa115_xor1;
  wire [0:0] s_wallace_rca24_fa115_or0;
  wire [0:0] s_wallace_rca24_and_19_20;
  wire [0:0] s_wallace_rca24_and_18_21;
  wire [0:0] s_wallace_rca24_fa116_xor1;
  wire [0:0] s_wallace_rca24_fa116_or0;
  wire [0:0] s_wallace_rca24_and_19_21;
  wire [0:0] s_wallace_rca24_and_18_22;
  wire [0:0] s_wallace_rca24_fa117_xor1;
  wire [0:0] s_wallace_rca24_fa117_or0;
  wire [0:0] s_wallace_rca24_and_19_22;
  wire [0:0] s_wallace_rca24_nand_18_23;
  wire [0:0] s_wallace_rca24_fa118_xor1;
  wire [0:0] s_wallace_rca24_fa118_or0;
  wire [0:0] s_wallace_rca24_nand_19_23;
  wire [0:0] s_wallace_rca24_fa119_xor1;
  wire [0:0] s_wallace_rca24_fa119_or0;
  wire [0:0] s_wallace_rca24_ha3_xor0;
  wire [0:0] s_wallace_rca24_ha3_and0;
  wire [0:0] s_wallace_rca24_and_0_6;
  wire [0:0] s_wallace_rca24_fa120_xor1;
  wire [0:0] s_wallace_rca24_fa120_or0;
  wire [0:0] s_wallace_rca24_and_1_6;
  wire [0:0] s_wallace_rca24_and_0_7;
  wire [0:0] s_wallace_rca24_fa121_xor1;
  wire [0:0] s_wallace_rca24_fa121_or0;
  wire [0:0] s_wallace_rca24_and_2_6;
  wire [0:0] s_wallace_rca24_and_1_7;
  wire [0:0] s_wallace_rca24_fa122_xor1;
  wire [0:0] s_wallace_rca24_fa122_or0;
  wire [0:0] s_wallace_rca24_and_3_6;
  wire [0:0] s_wallace_rca24_and_2_7;
  wire [0:0] s_wallace_rca24_fa123_xor1;
  wire [0:0] s_wallace_rca24_fa123_or0;
  wire [0:0] s_wallace_rca24_and_4_6;
  wire [0:0] s_wallace_rca24_and_3_7;
  wire [0:0] s_wallace_rca24_fa124_xor1;
  wire [0:0] s_wallace_rca24_fa124_or0;
  wire [0:0] s_wallace_rca24_and_5_6;
  wire [0:0] s_wallace_rca24_and_4_7;
  wire [0:0] s_wallace_rca24_fa125_xor1;
  wire [0:0] s_wallace_rca24_fa125_or0;
  wire [0:0] s_wallace_rca24_and_6_6;
  wire [0:0] s_wallace_rca24_and_5_7;
  wire [0:0] s_wallace_rca24_fa126_xor1;
  wire [0:0] s_wallace_rca24_fa126_or0;
  wire [0:0] s_wallace_rca24_and_7_6;
  wire [0:0] s_wallace_rca24_and_6_7;
  wire [0:0] s_wallace_rca24_fa127_xor1;
  wire [0:0] s_wallace_rca24_fa127_or0;
  wire [0:0] s_wallace_rca24_and_8_6;
  wire [0:0] s_wallace_rca24_and_7_7;
  wire [0:0] s_wallace_rca24_fa128_xor1;
  wire [0:0] s_wallace_rca24_fa128_or0;
  wire [0:0] s_wallace_rca24_and_9_6;
  wire [0:0] s_wallace_rca24_and_8_7;
  wire [0:0] s_wallace_rca24_fa129_xor1;
  wire [0:0] s_wallace_rca24_fa129_or0;
  wire [0:0] s_wallace_rca24_and_10_6;
  wire [0:0] s_wallace_rca24_and_9_7;
  wire [0:0] s_wallace_rca24_fa130_xor1;
  wire [0:0] s_wallace_rca24_fa130_or0;
  wire [0:0] s_wallace_rca24_and_11_6;
  wire [0:0] s_wallace_rca24_and_10_7;
  wire [0:0] s_wallace_rca24_fa131_xor1;
  wire [0:0] s_wallace_rca24_fa131_or0;
  wire [0:0] s_wallace_rca24_and_12_6;
  wire [0:0] s_wallace_rca24_and_11_7;
  wire [0:0] s_wallace_rca24_fa132_xor1;
  wire [0:0] s_wallace_rca24_fa132_or0;
  wire [0:0] s_wallace_rca24_and_13_6;
  wire [0:0] s_wallace_rca24_and_12_7;
  wire [0:0] s_wallace_rca24_fa133_xor1;
  wire [0:0] s_wallace_rca24_fa133_or0;
  wire [0:0] s_wallace_rca24_and_14_6;
  wire [0:0] s_wallace_rca24_and_13_7;
  wire [0:0] s_wallace_rca24_fa134_xor1;
  wire [0:0] s_wallace_rca24_fa134_or0;
  wire [0:0] s_wallace_rca24_and_15_6;
  wire [0:0] s_wallace_rca24_and_14_7;
  wire [0:0] s_wallace_rca24_fa135_xor1;
  wire [0:0] s_wallace_rca24_fa135_or0;
  wire [0:0] s_wallace_rca24_and_16_6;
  wire [0:0] s_wallace_rca24_and_15_7;
  wire [0:0] s_wallace_rca24_fa136_xor1;
  wire [0:0] s_wallace_rca24_fa136_or0;
  wire [0:0] s_wallace_rca24_and_17_6;
  wire [0:0] s_wallace_rca24_and_16_7;
  wire [0:0] s_wallace_rca24_fa137_xor1;
  wire [0:0] s_wallace_rca24_fa137_or0;
  wire [0:0] s_wallace_rca24_and_18_6;
  wire [0:0] s_wallace_rca24_and_17_7;
  wire [0:0] s_wallace_rca24_fa138_xor1;
  wire [0:0] s_wallace_rca24_fa138_or0;
  wire [0:0] s_wallace_rca24_and_17_8;
  wire [0:0] s_wallace_rca24_and_16_9;
  wire [0:0] s_wallace_rca24_fa139_xor1;
  wire [0:0] s_wallace_rca24_fa139_or0;
  wire [0:0] s_wallace_rca24_and_17_9;
  wire [0:0] s_wallace_rca24_and_16_10;
  wire [0:0] s_wallace_rca24_fa140_xor1;
  wire [0:0] s_wallace_rca24_fa140_or0;
  wire [0:0] s_wallace_rca24_and_17_10;
  wire [0:0] s_wallace_rca24_and_16_11;
  wire [0:0] s_wallace_rca24_fa141_xor1;
  wire [0:0] s_wallace_rca24_fa141_or0;
  wire [0:0] s_wallace_rca24_and_17_11;
  wire [0:0] s_wallace_rca24_and_16_12;
  wire [0:0] s_wallace_rca24_fa142_xor1;
  wire [0:0] s_wallace_rca24_fa142_or0;
  wire [0:0] s_wallace_rca24_and_17_12;
  wire [0:0] s_wallace_rca24_and_16_13;
  wire [0:0] s_wallace_rca24_fa143_xor1;
  wire [0:0] s_wallace_rca24_fa143_or0;
  wire [0:0] s_wallace_rca24_and_17_13;
  wire [0:0] s_wallace_rca24_and_16_14;
  wire [0:0] s_wallace_rca24_fa144_xor1;
  wire [0:0] s_wallace_rca24_fa144_or0;
  wire [0:0] s_wallace_rca24_and_17_14;
  wire [0:0] s_wallace_rca24_and_16_15;
  wire [0:0] s_wallace_rca24_fa145_xor1;
  wire [0:0] s_wallace_rca24_fa145_or0;
  wire [0:0] s_wallace_rca24_and_17_15;
  wire [0:0] s_wallace_rca24_and_16_16;
  wire [0:0] s_wallace_rca24_fa146_xor1;
  wire [0:0] s_wallace_rca24_fa146_or0;
  wire [0:0] s_wallace_rca24_and_17_16;
  wire [0:0] s_wallace_rca24_and_16_17;
  wire [0:0] s_wallace_rca24_fa147_xor1;
  wire [0:0] s_wallace_rca24_fa147_or0;
  wire [0:0] s_wallace_rca24_and_17_17;
  wire [0:0] s_wallace_rca24_and_16_18;
  wire [0:0] s_wallace_rca24_fa148_xor1;
  wire [0:0] s_wallace_rca24_fa148_or0;
  wire [0:0] s_wallace_rca24_and_17_18;
  wire [0:0] s_wallace_rca24_and_16_19;
  wire [0:0] s_wallace_rca24_fa149_xor1;
  wire [0:0] s_wallace_rca24_fa149_or0;
  wire [0:0] s_wallace_rca24_and_17_19;
  wire [0:0] s_wallace_rca24_and_16_20;
  wire [0:0] s_wallace_rca24_fa150_xor1;
  wire [0:0] s_wallace_rca24_fa150_or0;
  wire [0:0] s_wallace_rca24_and_17_20;
  wire [0:0] s_wallace_rca24_and_16_21;
  wire [0:0] s_wallace_rca24_fa151_xor1;
  wire [0:0] s_wallace_rca24_fa151_or0;
  wire [0:0] s_wallace_rca24_and_17_21;
  wire [0:0] s_wallace_rca24_and_16_22;
  wire [0:0] s_wallace_rca24_fa152_xor1;
  wire [0:0] s_wallace_rca24_fa152_or0;
  wire [0:0] s_wallace_rca24_and_17_22;
  wire [0:0] s_wallace_rca24_nand_16_23;
  wire [0:0] s_wallace_rca24_fa153_xor1;
  wire [0:0] s_wallace_rca24_fa153_or0;
  wire [0:0] s_wallace_rca24_nand_17_23;
  wire [0:0] s_wallace_rca24_fa154_xor1;
  wire [0:0] s_wallace_rca24_fa154_or0;
  wire [0:0] s_wallace_rca24_fa155_xor1;
  wire [0:0] s_wallace_rca24_fa155_or0;
  wire [0:0] s_wallace_rca24_ha4_xor0;
  wire [0:0] s_wallace_rca24_ha4_and0;
  wire [0:0] s_wallace_rca24_fa156_xor1;
  wire [0:0] s_wallace_rca24_fa156_or0;
  wire [0:0] s_wallace_rca24_and_0_8;
  wire [0:0] s_wallace_rca24_fa157_xor1;
  wire [0:0] s_wallace_rca24_fa157_or0;
  wire [0:0] s_wallace_rca24_and_1_8;
  wire [0:0] s_wallace_rca24_and_0_9;
  wire [0:0] s_wallace_rca24_fa158_xor1;
  wire [0:0] s_wallace_rca24_fa158_or0;
  wire [0:0] s_wallace_rca24_and_2_8;
  wire [0:0] s_wallace_rca24_and_1_9;
  wire [0:0] s_wallace_rca24_fa159_xor1;
  wire [0:0] s_wallace_rca24_fa159_or0;
  wire [0:0] s_wallace_rca24_and_3_8;
  wire [0:0] s_wallace_rca24_and_2_9;
  wire [0:0] s_wallace_rca24_fa160_xor1;
  wire [0:0] s_wallace_rca24_fa160_or0;
  wire [0:0] s_wallace_rca24_and_4_8;
  wire [0:0] s_wallace_rca24_and_3_9;
  wire [0:0] s_wallace_rca24_fa161_xor1;
  wire [0:0] s_wallace_rca24_fa161_or0;
  wire [0:0] s_wallace_rca24_and_5_8;
  wire [0:0] s_wallace_rca24_and_4_9;
  wire [0:0] s_wallace_rca24_fa162_xor1;
  wire [0:0] s_wallace_rca24_fa162_or0;
  wire [0:0] s_wallace_rca24_and_6_8;
  wire [0:0] s_wallace_rca24_and_5_9;
  wire [0:0] s_wallace_rca24_fa163_xor1;
  wire [0:0] s_wallace_rca24_fa163_or0;
  wire [0:0] s_wallace_rca24_and_7_8;
  wire [0:0] s_wallace_rca24_and_6_9;
  wire [0:0] s_wallace_rca24_fa164_xor1;
  wire [0:0] s_wallace_rca24_fa164_or0;
  wire [0:0] s_wallace_rca24_and_8_8;
  wire [0:0] s_wallace_rca24_and_7_9;
  wire [0:0] s_wallace_rca24_fa165_xor1;
  wire [0:0] s_wallace_rca24_fa165_or0;
  wire [0:0] s_wallace_rca24_and_9_8;
  wire [0:0] s_wallace_rca24_and_8_9;
  wire [0:0] s_wallace_rca24_fa166_xor1;
  wire [0:0] s_wallace_rca24_fa166_or0;
  wire [0:0] s_wallace_rca24_and_10_8;
  wire [0:0] s_wallace_rca24_and_9_9;
  wire [0:0] s_wallace_rca24_fa167_xor1;
  wire [0:0] s_wallace_rca24_fa167_or0;
  wire [0:0] s_wallace_rca24_and_11_8;
  wire [0:0] s_wallace_rca24_and_10_9;
  wire [0:0] s_wallace_rca24_fa168_xor1;
  wire [0:0] s_wallace_rca24_fa168_or0;
  wire [0:0] s_wallace_rca24_and_12_8;
  wire [0:0] s_wallace_rca24_and_11_9;
  wire [0:0] s_wallace_rca24_fa169_xor1;
  wire [0:0] s_wallace_rca24_fa169_or0;
  wire [0:0] s_wallace_rca24_and_13_8;
  wire [0:0] s_wallace_rca24_and_12_9;
  wire [0:0] s_wallace_rca24_fa170_xor1;
  wire [0:0] s_wallace_rca24_fa170_or0;
  wire [0:0] s_wallace_rca24_and_14_8;
  wire [0:0] s_wallace_rca24_and_13_9;
  wire [0:0] s_wallace_rca24_fa171_xor1;
  wire [0:0] s_wallace_rca24_fa171_or0;
  wire [0:0] s_wallace_rca24_and_15_8;
  wire [0:0] s_wallace_rca24_and_14_9;
  wire [0:0] s_wallace_rca24_fa172_xor1;
  wire [0:0] s_wallace_rca24_fa172_or0;
  wire [0:0] s_wallace_rca24_and_16_8;
  wire [0:0] s_wallace_rca24_and_15_9;
  wire [0:0] s_wallace_rca24_fa173_xor1;
  wire [0:0] s_wallace_rca24_fa173_or0;
  wire [0:0] s_wallace_rca24_and_15_10;
  wire [0:0] s_wallace_rca24_and_14_11;
  wire [0:0] s_wallace_rca24_fa174_xor1;
  wire [0:0] s_wallace_rca24_fa174_or0;
  wire [0:0] s_wallace_rca24_and_15_11;
  wire [0:0] s_wallace_rca24_and_14_12;
  wire [0:0] s_wallace_rca24_fa175_xor1;
  wire [0:0] s_wallace_rca24_fa175_or0;
  wire [0:0] s_wallace_rca24_and_15_12;
  wire [0:0] s_wallace_rca24_and_14_13;
  wire [0:0] s_wallace_rca24_fa176_xor1;
  wire [0:0] s_wallace_rca24_fa176_or0;
  wire [0:0] s_wallace_rca24_and_15_13;
  wire [0:0] s_wallace_rca24_and_14_14;
  wire [0:0] s_wallace_rca24_fa177_xor1;
  wire [0:0] s_wallace_rca24_fa177_or0;
  wire [0:0] s_wallace_rca24_and_15_14;
  wire [0:0] s_wallace_rca24_and_14_15;
  wire [0:0] s_wallace_rca24_fa178_xor1;
  wire [0:0] s_wallace_rca24_fa178_or0;
  wire [0:0] s_wallace_rca24_and_15_15;
  wire [0:0] s_wallace_rca24_and_14_16;
  wire [0:0] s_wallace_rca24_fa179_xor1;
  wire [0:0] s_wallace_rca24_fa179_or0;
  wire [0:0] s_wallace_rca24_and_15_16;
  wire [0:0] s_wallace_rca24_and_14_17;
  wire [0:0] s_wallace_rca24_fa180_xor1;
  wire [0:0] s_wallace_rca24_fa180_or0;
  wire [0:0] s_wallace_rca24_and_15_17;
  wire [0:0] s_wallace_rca24_and_14_18;
  wire [0:0] s_wallace_rca24_fa181_xor1;
  wire [0:0] s_wallace_rca24_fa181_or0;
  wire [0:0] s_wallace_rca24_and_15_18;
  wire [0:0] s_wallace_rca24_and_14_19;
  wire [0:0] s_wallace_rca24_fa182_xor1;
  wire [0:0] s_wallace_rca24_fa182_or0;
  wire [0:0] s_wallace_rca24_and_15_19;
  wire [0:0] s_wallace_rca24_and_14_20;
  wire [0:0] s_wallace_rca24_fa183_xor1;
  wire [0:0] s_wallace_rca24_fa183_or0;
  wire [0:0] s_wallace_rca24_and_15_20;
  wire [0:0] s_wallace_rca24_and_14_21;
  wire [0:0] s_wallace_rca24_fa184_xor1;
  wire [0:0] s_wallace_rca24_fa184_or0;
  wire [0:0] s_wallace_rca24_and_15_21;
  wire [0:0] s_wallace_rca24_and_14_22;
  wire [0:0] s_wallace_rca24_fa185_xor1;
  wire [0:0] s_wallace_rca24_fa185_or0;
  wire [0:0] s_wallace_rca24_and_15_22;
  wire [0:0] s_wallace_rca24_nand_14_23;
  wire [0:0] s_wallace_rca24_fa186_xor1;
  wire [0:0] s_wallace_rca24_fa186_or0;
  wire [0:0] s_wallace_rca24_nand_15_23;
  wire [0:0] s_wallace_rca24_fa187_xor1;
  wire [0:0] s_wallace_rca24_fa187_or0;
  wire [0:0] s_wallace_rca24_fa188_xor1;
  wire [0:0] s_wallace_rca24_fa188_or0;
  wire [0:0] s_wallace_rca24_fa189_xor1;
  wire [0:0] s_wallace_rca24_fa189_or0;
  wire [0:0] s_wallace_rca24_ha5_xor0;
  wire [0:0] s_wallace_rca24_ha5_and0;
  wire [0:0] s_wallace_rca24_fa190_xor1;
  wire [0:0] s_wallace_rca24_fa190_or0;
  wire [0:0] s_wallace_rca24_fa191_xor1;
  wire [0:0] s_wallace_rca24_fa191_or0;
  wire [0:0] s_wallace_rca24_and_0_10;
  wire [0:0] s_wallace_rca24_fa192_xor1;
  wire [0:0] s_wallace_rca24_fa192_or0;
  wire [0:0] s_wallace_rca24_and_1_10;
  wire [0:0] s_wallace_rca24_and_0_11;
  wire [0:0] s_wallace_rca24_fa193_xor1;
  wire [0:0] s_wallace_rca24_fa193_or0;
  wire [0:0] s_wallace_rca24_and_2_10;
  wire [0:0] s_wallace_rca24_and_1_11;
  wire [0:0] s_wallace_rca24_fa194_xor1;
  wire [0:0] s_wallace_rca24_fa194_or0;
  wire [0:0] s_wallace_rca24_and_3_10;
  wire [0:0] s_wallace_rca24_and_2_11;
  wire [0:0] s_wallace_rca24_fa195_xor1;
  wire [0:0] s_wallace_rca24_fa195_or0;
  wire [0:0] s_wallace_rca24_and_4_10;
  wire [0:0] s_wallace_rca24_and_3_11;
  wire [0:0] s_wallace_rca24_fa196_xor1;
  wire [0:0] s_wallace_rca24_fa196_or0;
  wire [0:0] s_wallace_rca24_and_5_10;
  wire [0:0] s_wallace_rca24_and_4_11;
  wire [0:0] s_wallace_rca24_fa197_xor1;
  wire [0:0] s_wallace_rca24_fa197_or0;
  wire [0:0] s_wallace_rca24_and_6_10;
  wire [0:0] s_wallace_rca24_and_5_11;
  wire [0:0] s_wallace_rca24_fa198_xor1;
  wire [0:0] s_wallace_rca24_fa198_or0;
  wire [0:0] s_wallace_rca24_and_7_10;
  wire [0:0] s_wallace_rca24_and_6_11;
  wire [0:0] s_wallace_rca24_fa199_xor1;
  wire [0:0] s_wallace_rca24_fa199_or0;
  wire [0:0] s_wallace_rca24_and_8_10;
  wire [0:0] s_wallace_rca24_and_7_11;
  wire [0:0] s_wallace_rca24_fa200_xor1;
  wire [0:0] s_wallace_rca24_fa200_or0;
  wire [0:0] s_wallace_rca24_and_9_10;
  wire [0:0] s_wallace_rca24_and_8_11;
  wire [0:0] s_wallace_rca24_fa201_xor1;
  wire [0:0] s_wallace_rca24_fa201_or0;
  wire [0:0] s_wallace_rca24_and_10_10;
  wire [0:0] s_wallace_rca24_and_9_11;
  wire [0:0] s_wallace_rca24_fa202_xor1;
  wire [0:0] s_wallace_rca24_fa202_or0;
  wire [0:0] s_wallace_rca24_and_11_10;
  wire [0:0] s_wallace_rca24_and_10_11;
  wire [0:0] s_wallace_rca24_fa203_xor1;
  wire [0:0] s_wallace_rca24_fa203_or0;
  wire [0:0] s_wallace_rca24_and_12_10;
  wire [0:0] s_wallace_rca24_and_11_11;
  wire [0:0] s_wallace_rca24_fa204_xor1;
  wire [0:0] s_wallace_rca24_fa204_or0;
  wire [0:0] s_wallace_rca24_and_13_10;
  wire [0:0] s_wallace_rca24_and_12_11;
  wire [0:0] s_wallace_rca24_fa205_xor1;
  wire [0:0] s_wallace_rca24_fa205_or0;
  wire [0:0] s_wallace_rca24_and_14_10;
  wire [0:0] s_wallace_rca24_and_13_11;
  wire [0:0] s_wallace_rca24_fa206_xor1;
  wire [0:0] s_wallace_rca24_fa206_or0;
  wire [0:0] s_wallace_rca24_and_13_12;
  wire [0:0] s_wallace_rca24_and_12_13;
  wire [0:0] s_wallace_rca24_fa207_xor1;
  wire [0:0] s_wallace_rca24_fa207_or0;
  wire [0:0] s_wallace_rca24_and_13_13;
  wire [0:0] s_wallace_rca24_and_12_14;
  wire [0:0] s_wallace_rca24_fa208_xor1;
  wire [0:0] s_wallace_rca24_fa208_or0;
  wire [0:0] s_wallace_rca24_and_13_14;
  wire [0:0] s_wallace_rca24_and_12_15;
  wire [0:0] s_wallace_rca24_fa209_xor1;
  wire [0:0] s_wallace_rca24_fa209_or0;
  wire [0:0] s_wallace_rca24_and_13_15;
  wire [0:0] s_wallace_rca24_and_12_16;
  wire [0:0] s_wallace_rca24_fa210_xor1;
  wire [0:0] s_wallace_rca24_fa210_or0;
  wire [0:0] s_wallace_rca24_and_13_16;
  wire [0:0] s_wallace_rca24_and_12_17;
  wire [0:0] s_wallace_rca24_fa211_xor1;
  wire [0:0] s_wallace_rca24_fa211_or0;
  wire [0:0] s_wallace_rca24_and_13_17;
  wire [0:0] s_wallace_rca24_and_12_18;
  wire [0:0] s_wallace_rca24_fa212_xor1;
  wire [0:0] s_wallace_rca24_fa212_or0;
  wire [0:0] s_wallace_rca24_and_13_18;
  wire [0:0] s_wallace_rca24_and_12_19;
  wire [0:0] s_wallace_rca24_fa213_xor1;
  wire [0:0] s_wallace_rca24_fa213_or0;
  wire [0:0] s_wallace_rca24_and_13_19;
  wire [0:0] s_wallace_rca24_and_12_20;
  wire [0:0] s_wallace_rca24_fa214_xor1;
  wire [0:0] s_wallace_rca24_fa214_or0;
  wire [0:0] s_wallace_rca24_and_13_20;
  wire [0:0] s_wallace_rca24_and_12_21;
  wire [0:0] s_wallace_rca24_fa215_xor1;
  wire [0:0] s_wallace_rca24_fa215_or0;
  wire [0:0] s_wallace_rca24_and_13_21;
  wire [0:0] s_wallace_rca24_and_12_22;
  wire [0:0] s_wallace_rca24_fa216_xor1;
  wire [0:0] s_wallace_rca24_fa216_or0;
  wire [0:0] s_wallace_rca24_and_13_22;
  wire [0:0] s_wallace_rca24_nand_12_23;
  wire [0:0] s_wallace_rca24_fa217_xor1;
  wire [0:0] s_wallace_rca24_fa217_or0;
  wire [0:0] s_wallace_rca24_nand_13_23;
  wire [0:0] s_wallace_rca24_fa218_xor1;
  wire [0:0] s_wallace_rca24_fa218_or0;
  wire [0:0] s_wallace_rca24_fa219_xor1;
  wire [0:0] s_wallace_rca24_fa219_or0;
  wire [0:0] s_wallace_rca24_fa220_xor1;
  wire [0:0] s_wallace_rca24_fa220_or0;
  wire [0:0] s_wallace_rca24_fa221_xor1;
  wire [0:0] s_wallace_rca24_fa221_or0;
  wire [0:0] s_wallace_rca24_ha6_xor0;
  wire [0:0] s_wallace_rca24_ha6_and0;
  wire [0:0] s_wallace_rca24_fa222_xor1;
  wire [0:0] s_wallace_rca24_fa222_or0;
  wire [0:0] s_wallace_rca24_fa223_xor1;
  wire [0:0] s_wallace_rca24_fa223_or0;
  wire [0:0] s_wallace_rca24_fa224_xor1;
  wire [0:0] s_wallace_rca24_fa224_or0;
  wire [0:0] s_wallace_rca24_and_0_12;
  wire [0:0] s_wallace_rca24_fa225_xor1;
  wire [0:0] s_wallace_rca24_fa225_or0;
  wire [0:0] s_wallace_rca24_and_1_12;
  wire [0:0] s_wallace_rca24_and_0_13;
  wire [0:0] s_wallace_rca24_fa226_xor1;
  wire [0:0] s_wallace_rca24_fa226_or0;
  wire [0:0] s_wallace_rca24_and_2_12;
  wire [0:0] s_wallace_rca24_and_1_13;
  wire [0:0] s_wallace_rca24_fa227_xor1;
  wire [0:0] s_wallace_rca24_fa227_or0;
  wire [0:0] s_wallace_rca24_and_3_12;
  wire [0:0] s_wallace_rca24_and_2_13;
  wire [0:0] s_wallace_rca24_fa228_xor1;
  wire [0:0] s_wallace_rca24_fa228_or0;
  wire [0:0] s_wallace_rca24_and_4_12;
  wire [0:0] s_wallace_rca24_and_3_13;
  wire [0:0] s_wallace_rca24_fa229_xor1;
  wire [0:0] s_wallace_rca24_fa229_or0;
  wire [0:0] s_wallace_rca24_and_5_12;
  wire [0:0] s_wallace_rca24_and_4_13;
  wire [0:0] s_wallace_rca24_fa230_xor1;
  wire [0:0] s_wallace_rca24_fa230_or0;
  wire [0:0] s_wallace_rca24_and_6_12;
  wire [0:0] s_wallace_rca24_and_5_13;
  wire [0:0] s_wallace_rca24_fa231_xor1;
  wire [0:0] s_wallace_rca24_fa231_or0;
  wire [0:0] s_wallace_rca24_and_7_12;
  wire [0:0] s_wallace_rca24_and_6_13;
  wire [0:0] s_wallace_rca24_fa232_xor1;
  wire [0:0] s_wallace_rca24_fa232_or0;
  wire [0:0] s_wallace_rca24_and_8_12;
  wire [0:0] s_wallace_rca24_and_7_13;
  wire [0:0] s_wallace_rca24_fa233_xor1;
  wire [0:0] s_wallace_rca24_fa233_or0;
  wire [0:0] s_wallace_rca24_and_9_12;
  wire [0:0] s_wallace_rca24_and_8_13;
  wire [0:0] s_wallace_rca24_fa234_xor1;
  wire [0:0] s_wallace_rca24_fa234_or0;
  wire [0:0] s_wallace_rca24_and_10_12;
  wire [0:0] s_wallace_rca24_and_9_13;
  wire [0:0] s_wallace_rca24_fa235_xor1;
  wire [0:0] s_wallace_rca24_fa235_or0;
  wire [0:0] s_wallace_rca24_and_11_12;
  wire [0:0] s_wallace_rca24_and_10_13;
  wire [0:0] s_wallace_rca24_fa236_xor1;
  wire [0:0] s_wallace_rca24_fa236_or0;
  wire [0:0] s_wallace_rca24_and_12_12;
  wire [0:0] s_wallace_rca24_and_11_13;
  wire [0:0] s_wallace_rca24_fa237_xor1;
  wire [0:0] s_wallace_rca24_fa237_or0;
  wire [0:0] s_wallace_rca24_and_11_14;
  wire [0:0] s_wallace_rca24_and_10_15;
  wire [0:0] s_wallace_rca24_fa238_xor1;
  wire [0:0] s_wallace_rca24_fa238_or0;
  wire [0:0] s_wallace_rca24_and_11_15;
  wire [0:0] s_wallace_rca24_and_10_16;
  wire [0:0] s_wallace_rca24_fa239_xor1;
  wire [0:0] s_wallace_rca24_fa239_or0;
  wire [0:0] s_wallace_rca24_and_11_16;
  wire [0:0] s_wallace_rca24_and_10_17;
  wire [0:0] s_wallace_rca24_fa240_xor1;
  wire [0:0] s_wallace_rca24_fa240_or0;
  wire [0:0] s_wallace_rca24_and_11_17;
  wire [0:0] s_wallace_rca24_and_10_18;
  wire [0:0] s_wallace_rca24_fa241_xor1;
  wire [0:0] s_wallace_rca24_fa241_or0;
  wire [0:0] s_wallace_rca24_and_11_18;
  wire [0:0] s_wallace_rca24_and_10_19;
  wire [0:0] s_wallace_rca24_fa242_xor1;
  wire [0:0] s_wallace_rca24_fa242_or0;
  wire [0:0] s_wallace_rca24_and_11_19;
  wire [0:0] s_wallace_rca24_and_10_20;
  wire [0:0] s_wallace_rca24_fa243_xor1;
  wire [0:0] s_wallace_rca24_fa243_or0;
  wire [0:0] s_wallace_rca24_and_11_20;
  wire [0:0] s_wallace_rca24_and_10_21;
  wire [0:0] s_wallace_rca24_fa244_xor1;
  wire [0:0] s_wallace_rca24_fa244_or0;
  wire [0:0] s_wallace_rca24_and_11_21;
  wire [0:0] s_wallace_rca24_and_10_22;
  wire [0:0] s_wallace_rca24_fa245_xor1;
  wire [0:0] s_wallace_rca24_fa245_or0;
  wire [0:0] s_wallace_rca24_and_11_22;
  wire [0:0] s_wallace_rca24_nand_10_23;
  wire [0:0] s_wallace_rca24_fa246_xor1;
  wire [0:0] s_wallace_rca24_fa246_or0;
  wire [0:0] s_wallace_rca24_nand_11_23;
  wire [0:0] s_wallace_rca24_fa247_xor1;
  wire [0:0] s_wallace_rca24_fa247_or0;
  wire [0:0] s_wallace_rca24_fa248_xor1;
  wire [0:0] s_wallace_rca24_fa248_or0;
  wire [0:0] s_wallace_rca24_fa249_xor1;
  wire [0:0] s_wallace_rca24_fa249_or0;
  wire [0:0] s_wallace_rca24_fa250_xor1;
  wire [0:0] s_wallace_rca24_fa250_or0;
  wire [0:0] s_wallace_rca24_fa251_xor1;
  wire [0:0] s_wallace_rca24_fa251_or0;
  wire [0:0] s_wallace_rca24_ha7_xor0;
  wire [0:0] s_wallace_rca24_ha7_and0;
  wire [0:0] s_wallace_rca24_fa252_xor1;
  wire [0:0] s_wallace_rca24_fa252_or0;
  wire [0:0] s_wallace_rca24_fa253_xor1;
  wire [0:0] s_wallace_rca24_fa253_or0;
  wire [0:0] s_wallace_rca24_fa254_xor1;
  wire [0:0] s_wallace_rca24_fa254_or0;
  wire [0:0] s_wallace_rca24_fa255_xor1;
  wire [0:0] s_wallace_rca24_fa255_or0;
  wire [0:0] s_wallace_rca24_and_0_14;
  wire [0:0] s_wallace_rca24_fa256_xor1;
  wire [0:0] s_wallace_rca24_fa256_or0;
  wire [0:0] s_wallace_rca24_and_1_14;
  wire [0:0] s_wallace_rca24_and_0_15;
  wire [0:0] s_wallace_rca24_fa257_xor1;
  wire [0:0] s_wallace_rca24_fa257_or0;
  wire [0:0] s_wallace_rca24_and_2_14;
  wire [0:0] s_wallace_rca24_and_1_15;
  wire [0:0] s_wallace_rca24_fa258_xor1;
  wire [0:0] s_wallace_rca24_fa258_or0;
  wire [0:0] s_wallace_rca24_and_3_14;
  wire [0:0] s_wallace_rca24_and_2_15;
  wire [0:0] s_wallace_rca24_fa259_xor1;
  wire [0:0] s_wallace_rca24_fa259_or0;
  wire [0:0] s_wallace_rca24_and_4_14;
  wire [0:0] s_wallace_rca24_and_3_15;
  wire [0:0] s_wallace_rca24_fa260_xor1;
  wire [0:0] s_wallace_rca24_fa260_or0;
  wire [0:0] s_wallace_rca24_and_5_14;
  wire [0:0] s_wallace_rca24_and_4_15;
  wire [0:0] s_wallace_rca24_fa261_xor1;
  wire [0:0] s_wallace_rca24_fa261_or0;
  wire [0:0] s_wallace_rca24_and_6_14;
  wire [0:0] s_wallace_rca24_and_5_15;
  wire [0:0] s_wallace_rca24_fa262_xor1;
  wire [0:0] s_wallace_rca24_fa262_or0;
  wire [0:0] s_wallace_rca24_and_7_14;
  wire [0:0] s_wallace_rca24_and_6_15;
  wire [0:0] s_wallace_rca24_fa263_xor1;
  wire [0:0] s_wallace_rca24_fa263_or0;
  wire [0:0] s_wallace_rca24_and_8_14;
  wire [0:0] s_wallace_rca24_and_7_15;
  wire [0:0] s_wallace_rca24_fa264_xor1;
  wire [0:0] s_wallace_rca24_fa264_or0;
  wire [0:0] s_wallace_rca24_and_9_14;
  wire [0:0] s_wallace_rca24_and_8_15;
  wire [0:0] s_wallace_rca24_fa265_xor1;
  wire [0:0] s_wallace_rca24_fa265_or0;
  wire [0:0] s_wallace_rca24_and_10_14;
  wire [0:0] s_wallace_rca24_and_9_15;
  wire [0:0] s_wallace_rca24_fa266_xor1;
  wire [0:0] s_wallace_rca24_fa266_or0;
  wire [0:0] s_wallace_rca24_and_9_16;
  wire [0:0] s_wallace_rca24_and_8_17;
  wire [0:0] s_wallace_rca24_fa267_xor1;
  wire [0:0] s_wallace_rca24_fa267_or0;
  wire [0:0] s_wallace_rca24_and_9_17;
  wire [0:0] s_wallace_rca24_and_8_18;
  wire [0:0] s_wallace_rca24_fa268_xor1;
  wire [0:0] s_wallace_rca24_fa268_or0;
  wire [0:0] s_wallace_rca24_and_9_18;
  wire [0:0] s_wallace_rca24_and_8_19;
  wire [0:0] s_wallace_rca24_fa269_xor1;
  wire [0:0] s_wallace_rca24_fa269_or0;
  wire [0:0] s_wallace_rca24_and_9_19;
  wire [0:0] s_wallace_rca24_and_8_20;
  wire [0:0] s_wallace_rca24_fa270_xor1;
  wire [0:0] s_wallace_rca24_fa270_or0;
  wire [0:0] s_wallace_rca24_and_9_20;
  wire [0:0] s_wallace_rca24_and_8_21;
  wire [0:0] s_wallace_rca24_fa271_xor1;
  wire [0:0] s_wallace_rca24_fa271_or0;
  wire [0:0] s_wallace_rca24_and_9_21;
  wire [0:0] s_wallace_rca24_and_8_22;
  wire [0:0] s_wallace_rca24_fa272_xor1;
  wire [0:0] s_wallace_rca24_fa272_or0;
  wire [0:0] s_wallace_rca24_and_9_22;
  wire [0:0] s_wallace_rca24_nand_8_23;
  wire [0:0] s_wallace_rca24_fa273_xor1;
  wire [0:0] s_wallace_rca24_fa273_or0;
  wire [0:0] s_wallace_rca24_nand_9_23;
  wire [0:0] s_wallace_rca24_fa274_xor1;
  wire [0:0] s_wallace_rca24_fa274_or0;
  wire [0:0] s_wallace_rca24_fa275_xor1;
  wire [0:0] s_wallace_rca24_fa275_or0;
  wire [0:0] s_wallace_rca24_fa276_xor1;
  wire [0:0] s_wallace_rca24_fa276_or0;
  wire [0:0] s_wallace_rca24_fa277_xor1;
  wire [0:0] s_wallace_rca24_fa277_or0;
  wire [0:0] s_wallace_rca24_fa278_xor1;
  wire [0:0] s_wallace_rca24_fa278_or0;
  wire [0:0] s_wallace_rca24_fa279_xor1;
  wire [0:0] s_wallace_rca24_fa279_or0;
  wire [0:0] s_wallace_rca24_ha8_xor0;
  wire [0:0] s_wallace_rca24_ha8_and0;
  wire [0:0] s_wallace_rca24_fa280_xor1;
  wire [0:0] s_wallace_rca24_fa280_or0;
  wire [0:0] s_wallace_rca24_fa281_xor1;
  wire [0:0] s_wallace_rca24_fa281_or0;
  wire [0:0] s_wallace_rca24_fa282_xor1;
  wire [0:0] s_wallace_rca24_fa282_or0;
  wire [0:0] s_wallace_rca24_fa283_xor1;
  wire [0:0] s_wallace_rca24_fa283_or0;
  wire [0:0] s_wallace_rca24_fa284_xor1;
  wire [0:0] s_wallace_rca24_fa284_or0;
  wire [0:0] s_wallace_rca24_and_0_16;
  wire [0:0] s_wallace_rca24_fa285_xor1;
  wire [0:0] s_wallace_rca24_fa285_or0;
  wire [0:0] s_wallace_rca24_and_1_16;
  wire [0:0] s_wallace_rca24_and_0_17;
  wire [0:0] s_wallace_rca24_fa286_xor1;
  wire [0:0] s_wallace_rca24_fa286_or0;
  wire [0:0] s_wallace_rca24_and_2_16;
  wire [0:0] s_wallace_rca24_and_1_17;
  wire [0:0] s_wallace_rca24_fa287_xor1;
  wire [0:0] s_wallace_rca24_fa287_or0;
  wire [0:0] s_wallace_rca24_and_3_16;
  wire [0:0] s_wallace_rca24_and_2_17;
  wire [0:0] s_wallace_rca24_fa288_xor1;
  wire [0:0] s_wallace_rca24_fa288_or0;
  wire [0:0] s_wallace_rca24_and_4_16;
  wire [0:0] s_wallace_rca24_and_3_17;
  wire [0:0] s_wallace_rca24_fa289_xor1;
  wire [0:0] s_wallace_rca24_fa289_or0;
  wire [0:0] s_wallace_rca24_and_5_16;
  wire [0:0] s_wallace_rca24_and_4_17;
  wire [0:0] s_wallace_rca24_fa290_xor1;
  wire [0:0] s_wallace_rca24_fa290_or0;
  wire [0:0] s_wallace_rca24_and_6_16;
  wire [0:0] s_wallace_rca24_and_5_17;
  wire [0:0] s_wallace_rca24_fa291_xor1;
  wire [0:0] s_wallace_rca24_fa291_or0;
  wire [0:0] s_wallace_rca24_and_7_16;
  wire [0:0] s_wallace_rca24_and_6_17;
  wire [0:0] s_wallace_rca24_fa292_xor1;
  wire [0:0] s_wallace_rca24_fa292_or0;
  wire [0:0] s_wallace_rca24_and_8_16;
  wire [0:0] s_wallace_rca24_and_7_17;
  wire [0:0] s_wallace_rca24_fa293_xor1;
  wire [0:0] s_wallace_rca24_fa293_or0;
  wire [0:0] s_wallace_rca24_and_7_18;
  wire [0:0] s_wallace_rca24_and_6_19;
  wire [0:0] s_wallace_rca24_fa294_xor1;
  wire [0:0] s_wallace_rca24_fa294_or0;
  wire [0:0] s_wallace_rca24_and_7_19;
  wire [0:0] s_wallace_rca24_and_6_20;
  wire [0:0] s_wallace_rca24_fa295_xor1;
  wire [0:0] s_wallace_rca24_fa295_or0;
  wire [0:0] s_wallace_rca24_and_7_20;
  wire [0:0] s_wallace_rca24_and_6_21;
  wire [0:0] s_wallace_rca24_fa296_xor1;
  wire [0:0] s_wallace_rca24_fa296_or0;
  wire [0:0] s_wallace_rca24_and_7_21;
  wire [0:0] s_wallace_rca24_and_6_22;
  wire [0:0] s_wallace_rca24_fa297_xor1;
  wire [0:0] s_wallace_rca24_fa297_or0;
  wire [0:0] s_wallace_rca24_and_7_22;
  wire [0:0] s_wallace_rca24_nand_6_23;
  wire [0:0] s_wallace_rca24_fa298_xor1;
  wire [0:0] s_wallace_rca24_fa298_or0;
  wire [0:0] s_wallace_rca24_nand_7_23;
  wire [0:0] s_wallace_rca24_fa299_xor1;
  wire [0:0] s_wallace_rca24_fa299_or0;
  wire [0:0] s_wallace_rca24_fa300_xor1;
  wire [0:0] s_wallace_rca24_fa300_or0;
  wire [0:0] s_wallace_rca24_fa301_xor1;
  wire [0:0] s_wallace_rca24_fa301_or0;
  wire [0:0] s_wallace_rca24_fa302_xor1;
  wire [0:0] s_wallace_rca24_fa302_or0;
  wire [0:0] s_wallace_rca24_fa303_xor1;
  wire [0:0] s_wallace_rca24_fa303_or0;
  wire [0:0] s_wallace_rca24_fa304_xor1;
  wire [0:0] s_wallace_rca24_fa304_or0;
  wire [0:0] s_wallace_rca24_fa305_xor1;
  wire [0:0] s_wallace_rca24_fa305_or0;
  wire [0:0] s_wallace_rca24_ha9_xor0;
  wire [0:0] s_wallace_rca24_ha9_and0;
  wire [0:0] s_wallace_rca24_fa306_xor1;
  wire [0:0] s_wallace_rca24_fa306_or0;
  wire [0:0] s_wallace_rca24_fa307_xor1;
  wire [0:0] s_wallace_rca24_fa307_or0;
  wire [0:0] s_wallace_rca24_fa308_xor1;
  wire [0:0] s_wallace_rca24_fa308_or0;
  wire [0:0] s_wallace_rca24_fa309_xor1;
  wire [0:0] s_wallace_rca24_fa309_or0;
  wire [0:0] s_wallace_rca24_fa310_xor1;
  wire [0:0] s_wallace_rca24_fa310_or0;
  wire [0:0] s_wallace_rca24_fa311_xor1;
  wire [0:0] s_wallace_rca24_fa311_or0;
  wire [0:0] s_wallace_rca24_and_0_18;
  wire [0:0] s_wallace_rca24_fa312_xor1;
  wire [0:0] s_wallace_rca24_fa312_or0;
  wire [0:0] s_wallace_rca24_and_1_18;
  wire [0:0] s_wallace_rca24_and_0_19;
  wire [0:0] s_wallace_rca24_fa313_xor1;
  wire [0:0] s_wallace_rca24_fa313_or0;
  wire [0:0] s_wallace_rca24_and_2_18;
  wire [0:0] s_wallace_rca24_and_1_19;
  wire [0:0] s_wallace_rca24_fa314_xor1;
  wire [0:0] s_wallace_rca24_fa314_or0;
  wire [0:0] s_wallace_rca24_and_3_18;
  wire [0:0] s_wallace_rca24_and_2_19;
  wire [0:0] s_wallace_rca24_fa315_xor1;
  wire [0:0] s_wallace_rca24_fa315_or0;
  wire [0:0] s_wallace_rca24_and_4_18;
  wire [0:0] s_wallace_rca24_and_3_19;
  wire [0:0] s_wallace_rca24_fa316_xor1;
  wire [0:0] s_wallace_rca24_fa316_or0;
  wire [0:0] s_wallace_rca24_and_5_18;
  wire [0:0] s_wallace_rca24_and_4_19;
  wire [0:0] s_wallace_rca24_fa317_xor1;
  wire [0:0] s_wallace_rca24_fa317_or0;
  wire [0:0] s_wallace_rca24_and_6_18;
  wire [0:0] s_wallace_rca24_and_5_19;
  wire [0:0] s_wallace_rca24_fa318_xor1;
  wire [0:0] s_wallace_rca24_fa318_or0;
  wire [0:0] s_wallace_rca24_and_5_20;
  wire [0:0] s_wallace_rca24_and_4_21;
  wire [0:0] s_wallace_rca24_fa319_xor1;
  wire [0:0] s_wallace_rca24_fa319_or0;
  wire [0:0] s_wallace_rca24_and_5_21;
  wire [0:0] s_wallace_rca24_and_4_22;
  wire [0:0] s_wallace_rca24_fa320_xor1;
  wire [0:0] s_wallace_rca24_fa320_or0;
  wire [0:0] s_wallace_rca24_and_5_22;
  wire [0:0] s_wallace_rca24_nand_4_23;
  wire [0:0] s_wallace_rca24_fa321_xor1;
  wire [0:0] s_wallace_rca24_fa321_or0;
  wire [0:0] s_wallace_rca24_nand_5_23;
  wire [0:0] s_wallace_rca24_fa322_xor1;
  wire [0:0] s_wallace_rca24_fa322_or0;
  wire [0:0] s_wallace_rca24_fa323_xor1;
  wire [0:0] s_wallace_rca24_fa323_or0;
  wire [0:0] s_wallace_rca24_fa324_xor1;
  wire [0:0] s_wallace_rca24_fa324_or0;
  wire [0:0] s_wallace_rca24_fa325_xor1;
  wire [0:0] s_wallace_rca24_fa325_or0;
  wire [0:0] s_wallace_rca24_fa326_xor1;
  wire [0:0] s_wallace_rca24_fa326_or0;
  wire [0:0] s_wallace_rca24_fa327_xor1;
  wire [0:0] s_wallace_rca24_fa327_or0;
  wire [0:0] s_wallace_rca24_fa328_xor1;
  wire [0:0] s_wallace_rca24_fa328_or0;
  wire [0:0] s_wallace_rca24_fa329_xor1;
  wire [0:0] s_wallace_rca24_fa329_or0;
  wire [0:0] s_wallace_rca24_ha10_xor0;
  wire [0:0] s_wallace_rca24_ha10_and0;
  wire [0:0] s_wallace_rca24_fa330_xor1;
  wire [0:0] s_wallace_rca24_fa330_or0;
  wire [0:0] s_wallace_rca24_fa331_xor1;
  wire [0:0] s_wallace_rca24_fa331_or0;
  wire [0:0] s_wallace_rca24_fa332_xor1;
  wire [0:0] s_wallace_rca24_fa332_or0;
  wire [0:0] s_wallace_rca24_fa333_xor1;
  wire [0:0] s_wallace_rca24_fa333_or0;
  wire [0:0] s_wallace_rca24_fa334_xor1;
  wire [0:0] s_wallace_rca24_fa334_or0;
  wire [0:0] s_wallace_rca24_fa335_xor1;
  wire [0:0] s_wallace_rca24_fa335_or0;
  wire [0:0] s_wallace_rca24_fa336_xor1;
  wire [0:0] s_wallace_rca24_fa336_or0;
  wire [0:0] s_wallace_rca24_and_0_20;
  wire [0:0] s_wallace_rca24_fa337_xor1;
  wire [0:0] s_wallace_rca24_fa337_or0;
  wire [0:0] s_wallace_rca24_and_1_20;
  wire [0:0] s_wallace_rca24_and_0_21;
  wire [0:0] s_wallace_rca24_fa338_xor1;
  wire [0:0] s_wallace_rca24_fa338_or0;
  wire [0:0] s_wallace_rca24_and_2_20;
  wire [0:0] s_wallace_rca24_and_1_21;
  wire [0:0] s_wallace_rca24_fa339_xor1;
  wire [0:0] s_wallace_rca24_fa339_or0;
  wire [0:0] s_wallace_rca24_and_3_20;
  wire [0:0] s_wallace_rca24_and_2_21;
  wire [0:0] s_wallace_rca24_fa340_xor1;
  wire [0:0] s_wallace_rca24_fa340_or0;
  wire [0:0] s_wallace_rca24_and_4_20;
  wire [0:0] s_wallace_rca24_and_3_21;
  wire [0:0] s_wallace_rca24_fa341_xor1;
  wire [0:0] s_wallace_rca24_fa341_or0;
  wire [0:0] s_wallace_rca24_and_3_22;
  wire [0:0] s_wallace_rca24_nand_2_23;
  wire [0:0] s_wallace_rca24_fa342_xor1;
  wire [0:0] s_wallace_rca24_fa342_or0;
  wire [0:0] s_wallace_rca24_nand_3_23;
  wire [0:0] s_wallace_rca24_fa343_xor1;
  wire [0:0] s_wallace_rca24_fa343_or0;
  wire [0:0] s_wallace_rca24_fa344_xor1;
  wire [0:0] s_wallace_rca24_fa344_or0;
  wire [0:0] s_wallace_rca24_fa345_xor1;
  wire [0:0] s_wallace_rca24_fa345_or0;
  wire [0:0] s_wallace_rca24_fa346_xor1;
  wire [0:0] s_wallace_rca24_fa346_or0;
  wire [0:0] s_wallace_rca24_fa347_xor1;
  wire [0:0] s_wallace_rca24_fa347_or0;
  wire [0:0] s_wallace_rca24_fa348_xor1;
  wire [0:0] s_wallace_rca24_fa348_or0;
  wire [0:0] s_wallace_rca24_fa349_xor1;
  wire [0:0] s_wallace_rca24_fa349_or0;
  wire [0:0] s_wallace_rca24_fa350_xor1;
  wire [0:0] s_wallace_rca24_fa350_or0;
  wire [0:0] s_wallace_rca24_fa351_xor1;
  wire [0:0] s_wallace_rca24_fa351_or0;
  wire [0:0] s_wallace_rca24_ha11_xor0;
  wire [0:0] s_wallace_rca24_ha11_and0;
  wire [0:0] s_wallace_rca24_fa352_xor1;
  wire [0:0] s_wallace_rca24_fa352_or0;
  wire [0:0] s_wallace_rca24_fa353_xor1;
  wire [0:0] s_wallace_rca24_fa353_or0;
  wire [0:0] s_wallace_rca24_fa354_xor1;
  wire [0:0] s_wallace_rca24_fa354_or0;
  wire [0:0] s_wallace_rca24_fa355_xor1;
  wire [0:0] s_wallace_rca24_fa355_or0;
  wire [0:0] s_wallace_rca24_fa356_xor1;
  wire [0:0] s_wallace_rca24_fa356_or0;
  wire [0:0] s_wallace_rca24_fa357_xor1;
  wire [0:0] s_wallace_rca24_fa357_or0;
  wire [0:0] s_wallace_rca24_fa358_xor1;
  wire [0:0] s_wallace_rca24_fa358_or0;
  wire [0:0] s_wallace_rca24_fa359_xor1;
  wire [0:0] s_wallace_rca24_fa359_or0;
  wire [0:0] s_wallace_rca24_and_0_22;
  wire [0:0] s_wallace_rca24_fa360_xor1;
  wire [0:0] s_wallace_rca24_fa360_or0;
  wire [0:0] s_wallace_rca24_and_1_22;
  wire [0:0] s_wallace_rca24_nand_0_23;
  wire [0:0] s_wallace_rca24_fa361_xor1;
  wire [0:0] s_wallace_rca24_fa361_or0;
  wire [0:0] s_wallace_rca24_and_2_22;
  wire [0:0] s_wallace_rca24_nand_1_23;
  wire [0:0] s_wallace_rca24_fa362_xor1;
  wire [0:0] s_wallace_rca24_fa362_or0;
  wire [0:0] s_wallace_rca24_fa363_xor1;
  wire [0:0] s_wallace_rca24_fa363_or0;
  wire [0:0] s_wallace_rca24_fa364_xor1;
  wire [0:0] s_wallace_rca24_fa364_or0;
  wire [0:0] s_wallace_rca24_fa365_xor1;
  wire [0:0] s_wallace_rca24_fa365_or0;
  wire [0:0] s_wallace_rca24_fa366_xor1;
  wire [0:0] s_wallace_rca24_fa366_or0;
  wire [0:0] s_wallace_rca24_fa367_xor1;
  wire [0:0] s_wallace_rca24_fa367_or0;
  wire [0:0] s_wallace_rca24_fa368_xor1;
  wire [0:0] s_wallace_rca24_fa368_or0;
  wire [0:0] s_wallace_rca24_fa369_xor1;
  wire [0:0] s_wallace_rca24_fa369_or0;
  wire [0:0] s_wallace_rca24_fa370_xor1;
  wire [0:0] s_wallace_rca24_fa370_or0;
  wire [0:0] s_wallace_rca24_fa371_xor1;
  wire [0:0] s_wallace_rca24_fa371_or0;
  wire [0:0] s_wallace_rca24_ha12_xor0;
  wire [0:0] s_wallace_rca24_ha12_and0;
  wire [0:0] s_wallace_rca24_fa372_xor1;
  wire [0:0] s_wallace_rca24_fa372_or0;
  wire [0:0] s_wallace_rca24_fa373_xor1;
  wire [0:0] s_wallace_rca24_fa373_or0;
  wire [0:0] s_wallace_rca24_fa374_xor1;
  wire [0:0] s_wallace_rca24_fa374_or0;
  wire [0:0] s_wallace_rca24_fa375_xor1;
  wire [0:0] s_wallace_rca24_fa375_or0;
  wire [0:0] s_wallace_rca24_fa376_xor1;
  wire [0:0] s_wallace_rca24_fa376_or0;
  wire [0:0] s_wallace_rca24_fa377_xor1;
  wire [0:0] s_wallace_rca24_fa377_or0;
  wire [0:0] s_wallace_rca24_fa378_xor1;
  wire [0:0] s_wallace_rca24_fa378_or0;
  wire [0:0] s_wallace_rca24_fa379_xor1;
  wire [0:0] s_wallace_rca24_fa379_or0;
  wire [0:0] s_wallace_rca24_fa380_xor1;
  wire [0:0] s_wallace_rca24_fa380_or0;
  wire [0:0] s_wallace_rca24_fa381_xor1;
  wire [0:0] s_wallace_rca24_fa381_or0;
  wire [0:0] s_wallace_rca24_fa382_xor1;
  wire [0:0] s_wallace_rca24_fa382_or0;
  wire [0:0] s_wallace_rca24_fa383_xor1;
  wire [0:0] s_wallace_rca24_fa383_or0;
  wire [0:0] s_wallace_rca24_fa384_xor1;
  wire [0:0] s_wallace_rca24_fa384_or0;
  wire [0:0] s_wallace_rca24_fa385_xor1;
  wire [0:0] s_wallace_rca24_fa385_or0;
  wire [0:0] s_wallace_rca24_fa386_xor1;
  wire [0:0] s_wallace_rca24_fa386_or0;
  wire [0:0] s_wallace_rca24_fa387_xor1;
  wire [0:0] s_wallace_rca24_fa387_or0;
  wire [0:0] s_wallace_rca24_fa388_xor1;
  wire [0:0] s_wallace_rca24_fa388_or0;
  wire [0:0] s_wallace_rca24_fa389_xor1;
  wire [0:0] s_wallace_rca24_fa389_or0;
  wire [0:0] s_wallace_rca24_ha13_xor0;
  wire [0:0] s_wallace_rca24_ha13_and0;
  wire [0:0] s_wallace_rca24_fa390_xor1;
  wire [0:0] s_wallace_rca24_fa390_or0;
  wire [0:0] s_wallace_rca24_fa391_xor1;
  wire [0:0] s_wallace_rca24_fa391_or0;
  wire [0:0] s_wallace_rca24_fa392_xor1;
  wire [0:0] s_wallace_rca24_fa392_or0;
  wire [0:0] s_wallace_rca24_fa393_xor1;
  wire [0:0] s_wallace_rca24_fa393_or0;
  wire [0:0] s_wallace_rca24_fa394_xor1;
  wire [0:0] s_wallace_rca24_fa394_or0;
  wire [0:0] s_wallace_rca24_fa395_xor1;
  wire [0:0] s_wallace_rca24_fa395_or0;
  wire [0:0] s_wallace_rca24_fa396_xor1;
  wire [0:0] s_wallace_rca24_fa396_or0;
  wire [0:0] s_wallace_rca24_fa397_xor1;
  wire [0:0] s_wallace_rca24_fa397_or0;
  wire [0:0] s_wallace_rca24_fa398_xor1;
  wire [0:0] s_wallace_rca24_fa398_or0;
  wire [0:0] s_wallace_rca24_fa399_xor1;
  wire [0:0] s_wallace_rca24_fa399_or0;
  wire [0:0] s_wallace_rca24_fa400_xor1;
  wire [0:0] s_wallace_rca24_fa400_or0;
  wire [0:0] s_wallace_rca24_fa401_xor1;
  wire [0:0] s_wallace_rca24_fa401_or0;
  wire [0:0] s_wallace_rca24_fa402_xor1;
  wire [0:0] s_wallace_rca24_fa402_or0;
  wire [0:0] s_wallace_rca24_fa403_xor1;
  wire [0:0] s_wallace_rca24_fa403_or0;
  wire [0:0] s_wallace_rca24_fa404_xor1;
  wire [0:0] s_wallace_rca24_fa404_or0;
  wire [0:0] s_wallace_rca24_fa405_xor1;
  wire [0:0] s_wallace_rca24_fa405_or0;
  wire [0:0] s_wallace_rca24_ha14_xor0;
  wire [0:0] s_wallace_rca24_ha14_and0;
  wire [0:0] s_wallace_rca24_fa406_xor1;
  wire [0:0] s_wallace_rca24_fa406_or0;
  wire [0:0] s_wallace_rca24_fa407_xor1;
  wire [0:0] s_wallace_rca24_fa407_or0;
  wire [0:0] s_wallace_rca24_fa408_xor1;
  wire [0:0] s_wallace_rca24_fa408_or0;
  wire [0:0] s_wallace_rca24_fa409_xor1;
  wire [0:0] s_wallace_rca24_fa409_or0;
  wire [0:0] s_wallace_rca24_fa410_xor1;
  wire [0:0] s_wallace_rca24_fa410_or0;
  wire [0:0] s_wallace_rca24_fa411_xor1;
  wire [0:0] s_wallace_rca24_fa411_or0;
  wire [0:0] s_wallace_rca24_fa412_xor1;
  wire [0:0] s_wallace_rca24_fa412_or0;
  wire [0:0] s_wallace_rca24_fa413_xor1;
  wire [0:0] s_wallace_rca24_fa413_or0;
  wire [0:0] s_wallace_rca24_fa414_xor1;
  wire [0:0] s_wallace_rca24_fa414_or0;
  wire [0:0] s_wallace_rca24_fa415_xor1;
  wire [0:0] s_wallace_rca24_fa415_or0;
  wire [0:0] s_wallace_rca24_fa416_xor1;
  wire [0:0] s_wallace_rca24_fa416_or0;
  wire [0:0] s_wallace_rca24_fa417_xor1;
  wire [0:0] s_wallace_rca24_fa417_or0;
  wire [0:0] s_wallace_rca24_fa418_xor1;
  wire [0:0] s_wallace_rca24_fa418_or0;
  wire [0:0] s_wallace_rca24_fa419_xor1;
  wire [0:0] s_wallace_rca24_fa419_or0;
  wire [0:0] s_wallace_rca24_ha15_xor0;
  wire [0:0] s_wallace_rca24_ha15_and0;
  wire [0:0] s_wallace_rca24_fa420_xor1;
  wire [0:0] s_wallace_rca24_fa420_or0;
  wire [0:0] s_wallace_rca24_fa421_xor1;
  wire [0:0] s_wallace_rca24_fa421_or0;
  wire [0:0] s_wallace_rca24_fa422_xor1;
  wire [0:0] s_wallace_rca24_fa422_or0;
  wire [0:0] s_wallace_rca24_fa423_xor1;
  wire [0:0] s_wallace_rca24_fa423_or0;
  wire [0:0] s_wallace_rca24_fa424_xor1;
  wire [0:0] s_wallace_rca24_fa424_or0;
  wire [0:0] s_wallace_rca24_fa425_xor1;
  wire [0:0] s_wallace_rca24_fa425_or0;
  wire [0:0] s_wallace_rca24_fa426_xor1;
  wire [0:0] s_wallace_rca24_fa426_or0;
  wire [0:0] s_wallace_rca24_fa427_xor1;
  wire [0:0] s_wallace_rca24_fa427_or0;
  wire [0:0] s_wallace_rca24_fa428_xor1;
  wire [0:0] s_wallace_rca24_fa428_or0;
  wire [0:0] s_wallace_rca24_fa429_xor1;
  wire [0:0] s_wallace_rca24_fa429_or0;
  wire [0:0] s_wallace_rca24_fa430_xor1;
  wire [0:0] s_wallace_rca24_fa430_or0;
  wire [0:0] s_wallace_rca24_fa431_xor1;
  wire [0:0] s_wallace_rca24_fa431_or0;
  wire [0:0] s_wallace_rca24_ha16_xor0;
  wire [0:0] s_wallace_rca24_ha16_and0;
  wire [0:0] s_wallace_rca24_fa432_xor1;
  wire [0:0] s_wallace_rca24_fa432_or0;
  wire [0:0] s_wallace_rca24_fa433_xor1;
  wire [0:0] s_wallace_rca24_fa433_or0;
  wire [0:0] s_wallace_rca24_fa434_xor1;
  wire [0:0] s_wallace_rca24_fa434_or0;
  wire [0:0] s_wallace_rca24_fa435_xor1;
  wire [0:0] s_wallace_rca24_fa435_or0;
  wire [0:0] s_wallace_rca24_fa436_xor1;
  wire [0:0] s_wallace_rca24_fa436_or0;
  wire [0:0] s_wallace_rca24_fa437_xor1;
  wire [0:0] s_wallace_rca24_fa437_or0;
  wire [0:0] s_wallace_rca24_fa438_xor1;
  wire [0:0] s_wallace_rca24_fa438_or0;
  wire [0:0] s_wallace_rca24_fa439_xor1;
  wire [0:0] s_wallace_rca24_fa439_or0;
  wire [0:0] s_wallace_rca24_fa440_xor1;
  wire [0:0] s_wallace_rca24_fa440_or0;
  wire [0:0] s_wallace_rca24_fa441_xor1;
  wire [0:0] s_wallace_rca24_fa441_or0;
  wire [0:0] s_wallace_rca24_ha17_xor0;
  wire [0:0] s_wallace_rca24_ha17_and0;
  wire [0:0] s_wallace_rca24_fa442_xor1;
  wire [0:0] s_wallace_rca24_fa442_or0;
  wire [0:0] s_wallace_rca24_fa443_xor1;
  wire [0:0] s_wallace_rca24_fa443_or0;
  wire [0:0] s_wallace_rca24_fa444_xor1;
  wire [0:0] s_wallace_rca24_fa444_or0;
  wire [0:0] s_wallace_rca24_fa445_xor1;
  wire [0:0] s_wallace_rca24_fa445_or0;
  wire [0:0] s_wallace_rca24_fa446_xor1;
  wire [0:0] s_wallace_rca24_fa446_or0;
  wire [0:0] s_wallace_rca24_fa447_xor1;
  wire [0:0] s_wallace_rca24_fa447_or0;
  wire [0:0] s_wallace_rca24_fa448_xor1;
  wire [0:0] s_wallace_rca24_fa448_or0;
  wire [0:0] s_wallace_rca24_fa449_xor1;
  wire [0:0] s_wallace_rca24_fa449_or0;
  wire [0:0] s_wallace_rca24_ha18_xor0;
  wire [0:0] s_wallace_rca24_ha18_and0;
  wire [0:0] s_wallace_rca24_fa450_xor1;
  wire [0:0] s_wallace_rca24_fa450_or0;
  wire [0:0] s_wallace_rca24_fa451_xor1;
  wire [0:0] s_wallace_rca24_fa451_or0;
  wire [0:0] s_wallace_rca24_fa452_xor1;
  wire [0:0] s_wallace_rca24_fa452_or0;
  wire [0:0] s_wallace_rca24_fa453_xor1;
  wire [0:0] s_wallace_rca24_fa453_or0;
  wire [0:0] s_wallace_rca24_fa454_xor1;
  wire [0:0] s_wallace_rca24_fa454_or0;
  wire [0:0] s_wallace_rca24_fa455_xor1;
  wire [0:0] s_wallace_rca24_fa455_or0;
  wire [0:0] s_wallace_rca24_ha19_xor0;
  wire [0:0] s_wallace_rca24_ha19_and0;
  wire [0:0] s_wallace_rca24_fa456_xor1;
  wire [0:0] s_wallace_rca24_fa456_or0;
  wire [0:0] s_wallace_rca24_fa457_xor1;
  wire [0:0] s_wallace_rca24_fa457_or0;
  wire [0:0] s_wallace_rca24_fa458_xor1;
  wire [0:0] s_wallace_rca24_fa458_or0;
  wire [0:0] s_wallace_rca24_fa459_xor1;
  wire [0:0] s_wallace_rca24_fa459_or0;
  wire [0:0] s_wallace_rca24_ha20_xor0;
  wire [0:0] s_wallace_rca24_ha20_and0;
  wire [0:0] s_wallace_rca24_fa460_xor1;
  wire [0:0] s_wallace_rca24_fa460_or0;
  wire [0:0] s_wallace_rca24_fa461_xor1;
  wire [0:0] s_wallace_rca24_fa461_or0;
  wire [0:0] s_wallace_rca24_ha21_xor0;
  wire [0:0] s_wallace_rca24_ha21_and0;
  wire [0:0] s_wallace_rca24_fa462_xor1;
  wire [0:0] s_wallace_rca24_fa462_or0;
  wire [0:0] s_wallace_rca24_fa463_xor1;
  wire [0:0] s_wallace_rca24_fa463_or0;
  wire [0:0] s_wallace_rca24_fa464_xor1;
  wire [0:0] s_wallace_rca24_fa464_or0;
  wire [0:0] s_wallace_rca24_fa465_xor1;
  wire [0:0] s_wallace_rca24_fa465_or0;
  wire [0:0] s_wallace_rca24_fa466_xor1;
  wire [0:0] s_wallace_rca24_fa466_or0;
  wire [0:0] s_wallace_rca24_fa467_xor1;
  wire [0:0] s_wallace_rca24_fa467_or0;
  wire [0:0] s_wallace_rca24_fa468_xor1;
  wire [0:0] s_wallace_rca24_fa468_or0;
  wire [0:0] s_wallace_rca24_fa469_xor1;
  wire [0:0] s_wallace_rca24_fa469_or0;
  wire [0:0] s_wallace_rca24_fa470_xor1;
  wire [0:0] s_wallace_rca24_fa470_or0;
  wire [0:0] s_wallace_rca24_fa471_xor1;
  wire [0:0] s_wallace_rca24_fa471_or0;
  wire [0:0] s_wallace_rca24_fa472_xor1;
  wire [0:0] s_wallace_rca24_fa472_or0;
  wire [0:0] s_wallace_rca24_fa473_xor1;
  wire [0:0] s_wallace_rca24_fa473_or0;
  wire [0:0] s_wallace_rca24_fa474_xor1;
  wire [0:0] s_wallace_rca24_fa474_or0;
  wire [0:0] s_wallace_rca24_fa475_xor1;
  wire [0:0] s_wallace_rca24_fa475_or0;
  wire [0:0] s_wallace_rca24_fa476_xor1;
  wire [0:0] s_wallace_rca24_fa476_or0;
  wire [0:0] s_wallace_rca24_fa477_xor1;
  wire [0:0] s_wallace_rca24_fa477_or0;
  wire [0:0] s_wallace_rca24_fa478_xor1;
  wire [0:0] s_wallace_rca24_fa478_or0;
  wire [0:0] s_wallace_rca24_fa479_xor1;
  wire [0:0] s_wallace_rca24_fa479_or0;
  wire [0:0] s_wallace_rca24_fa480_xor1;
  wire [0:0] s_wallace_rca24_fa480_or0;
  wire [0:0] s_wallace_rca24_fa481_xor1;
  wire [0:0] s_wallace_rca24_fa481_or0;
  wire [0:0] s_wallace_rca24_nand_21_23;
  wire [0:0] s_wallace_rca24_fa482_xor1;
  wire [0:0] s_wallace_rca24_fa482_or0;
  wire [0:0] s_wallace_rca24_nand_23_22;
  wire [0:0] s_wallace_rca24_fa483_xor1;
  wire [0:0] s_wallace_rca24_fa483_or0;
  wire [0:0] s_wallace_rca24_and_0_0;
  wire [0:0] s_wallace_rca24_and_1_0;
  wire [0:0] s_wallace_rca24_and_0_2;
  wire [0:0] s_wallace_rca24_nand_22_23;
  wire [0:0] s_wallace_rca24_and_0_1;
  wire [0:0] s_wallace_rca24_and_23_23;
  wire [45:0] s_wallace_rca24_u_rca46_a;
  wire [45:0] s_wallace_rca24_u_rca46_b;
  wire [46:0] s_wallace_rca24_u_rca46_out;
  wire [0:0] s_wallace_rca24_xor0;

  and_gate and_gate_s_wallace_rca24_and_2_0(.a(a[2]), .b(b[0]), .out(s_wallace_rca24_and_2_0));
  and_gate and_gate_s_wallace_rca24_and_1_1(.a(a[1]), .b(b[1]), .out(s_wallace_rca24_and_1_1));
  ha ha_s_wallace_rca24_ha0_out(.a(s_wallace_rca24_and_2_0[0]), .b(s_wallace_rca24_and_1_1[0]), .ha_xor0(s_wallace_rca24_ha0_xor0), .ha_and0(s_wallace_rca24_ha0_and0));
  and_gate and_gate_s_wallace_rca24_and_3_0(.a(a[3]), .b(b[0]), .out(s_wallace_rca24_and_3_0));
  and_gate and_gate_s_wallace_rca24_and_2_1(.a(a[2]), .b(b[1]), .out(s_wallace_rca24_and_2_1));
  fa fa_s_wallace_rca24_fa0_out(.a(s_wallace_rca24_ha0_and0[0]), .b(s_wallace_rca24_and_3_0[0]), .cin(s_wallace_rca24_and_2_1[0]), .fa_xor1(s_wallace_rca24_fa0_xor1), .fa_or0(s_wallace_rca24_fa0_or0));
  and_gate and_gate_s_wallace_rca24_and_4_0(.a(a[4]), .b(b[0]), .out(s_wallace_rca24_and_4_0));
  and_gate and_gate_s_wallace_rca24_and_3_1(.a(a[3]), .b(b[1]), .out(s_wallace_rca24_and_3_1));
  fa fa_s_wallace_rca24_fa1_out(.a(s_wallace_rca24_fa0_or0[0]), .b(s_wallace_rca24_and_4_0[0]), .cin(s_wallace_rca24_and_3_1[0]), .fa_xor1(s_wallace_rca24_fa1_xor1), .fa_or0(s_wallace_rca24_fa1_or0));
  and_gate and_gate_s_wallace_rca24_and_5_0(.a(a[5]), .b(b[0]), .out(s_wallace_rca24_and_5_0));
  and_gate and_gate_s_wallace_rca24_and_4_1(.a(a[4]), .b(b[1]), .out(s_wallace_rca24_and_4_1));
  fa fa_s_wallace_rca24_fa2_out(.a(s_wallace_rca24_fa1_or0[0]), .b(s_wallace_rca24_and_5_0[0]), .cin(s_wallace_rca24_and_4_1[0]), .fa_xor1(s_wallace_rca24_fa2_xor1), .fa_or0(s_wallace_rca24_fa2_or0));
  and_gate and_gate_s_wallace_rca24_and_6_0(.a(a[6]), .b(b[0]), .out(s_wallace_rca24_and_6_0));
  and_gate and_gate_s_wallace_rca24_and_5_1(.a(a[5]), .b(b[1]), .out(s_wallace_rca24_and_5_1));
  fa fa_s_wallace_rca24_fa3_out(.a(s_wallace_rca24_fa2_or0[0]), .b(s_wallace_rca24_and_6_0[0]), .cin(s_wallace_rca24_and_5_1[0]), .fa_xor1(s_wallace_rca24_fa3_xor1), .fa_or0(s_wallace_rca24_fa3_or0));
  and_gate and_gate_s_wallace_rca24_and_7_0(.a(a[7]), .b(b[0]), .out(s_wallace_rca24_and_7_0));
  and_gate and_gate_s_wallace_rca24_and_6_1(.a(a[6]), .b(b[1]), .out(s_wallace_rca24_and_6_1));
  fa fa_s_wallace_rca24_fa4_out(.a(s_wallace_rca24_fa3_or0[0]), .b(s_wallace_rca24_and_7_0[0]), .cin(s_wallace_rca24_and_6_1[0]), .fa_xor1(s_wallace_rca24_fa4_xor1), .fa_or0(s_wallace_rca24_fa4_or0));
  and_gate and_gate_s_wallace_rca24_and_8_0(.a(a[8]), .b(b[0]), .out(s_wallace_rca24_and_8_0));
  and_gate and_gate_s_wallace_rca24_and_7_1(.a(a[7]), .b(b[1]), .out(s_wallace_rca24_and_7_1));
  fa fa_s_wallace_rca24_fa5_out(.a(s_wallace_rca24_fa4_or0[0]), .b(s_wallace_rca24_and_8_0[0]), .cin(s_wallace_rca24_and_7_1[0]), .fa_xor1(s_wallace_rca24_fa5_xor1), .fa_or0(s_wallace_rca24_fa5_or0));
  and_gate and_gate_s_wallace_rca24_and_9_0(.a(a[9]), .b(b[0]), .out(s_wallace_rca24_and_9_0));
  and_gate and_gate_s_wallace_rca24_and_8_1(.a(a[8]), .b(b[1]), .out(s_wallace_rca24_and_8_1));
  fa fa_s_wallace_rca24_fa6_out(.a(s_wallace_rca24_fa5_or0[0]), .b(s_wallace_rca24_and_9_0[0]), .cin(s_wallace_rca24_and_8_1[0]), .fa_xor1(s_wallace_rca24_fa6_xor1), .fa_or0(s_wallace_rca24_fa6_or0));
  and_gate and_gate_s_wallace_rca24_and_10_0(.a(a[10]), .b(b[0]), .out(s_wallace_rca24_and_10_0));
  and_gate and_gate_s_wallace_rca24_and_9_1(.a(a[9]), .b(b[1]), .out(s_wallace_rca24_and_9_1));
  fa fa_s_wallace_rca24_fa7_out(.a(s_wallace_rca24_fa6_or0[0]), .b(s_wallace_rca24_and_10_0[0]), .cin(s_wallace_rca24_and_9_1[0]), .fa_xor1(s_wallace_rca24_fa7_xor1), .fa_or0(s_wallace_rca24_fa7_or0));
  and_gate and_gate_s_wallace_rca24_and_11_0(.a(a[11]), .b(b[0]), .out(s_wallace_rca24_and_11_0));
  and_gate and_gate_s_wallace_rca24_and_10_1(.a(a[10]), .b(b[1]), .out(s_wallace_rca24_and_10_1));
  fa fa_s_wallace_rca24_fa8_out(.a(s_wallace_rca24_fa7_or0[0]), .b(s_wallace_rca24_and_11_0[0]), .cin(s_wallace_rca24_and_10_1[0]), .fa_xor1(s_wallace_rca24_fa8_xor1), .fa_or0(s_wallace_rca24_fa8_or0));
  and_gate and_gate_s_wallace_rca24_and_12_0(.a(a[12]), .b(b[0]), .out(s_wallace_rca24_and_12_0));
  and_gate and_gate_s_wallace_rca24_and_11_1(.a(a[11]), .b(b[1]), .out(s_wallace_rca24_and_11_1));
  fa fa_s_wallace_rca24_fa9_out(.a(s_wallace_rca24_fa8_or0[0]), .b(s_wallace_rca24_and_12_0[0]), .cin(s_wallace_rca24_and_11_1[0]), .fa_xor1(s_wallace_rca24_fa9_xor1), .fa_or0(s_wallace_rca24_fa9_or0));
  and_gate and_gate_s_wallace_rca24_and_13_0(.a(a[13]), .b(b[0]), .out(s_wallace_rca24_and_13_0));
  and_gate and_gate_s_wallace_rca24_and_12_1(.a(a[12]), .b(b[1]), .out(s_wallace_rca24_and_12_1));
  fa fa_s_wallace_rca24_fa10_out(.a(s_wallace_rca24_fa9_or0[0]), .b(s_wallace_rca24_and_13_0[0]), .cin(s_wallace_rca24_and_12_1[0]), .fa_xor1(s_wallace_rca24_fa10_xor1), .fa_or0(s_wallace_rca24_fa10_or0));
  and_gate and_gate_s_wallace_rca24_and_14_0(.a(a[14]), .b(b[0]), .out(s_wallace_rca24_and_14_0));
  and_gate and_gate_s_wallace_rca24_and_13_1(.a(a[13]), .b(b[1]), .out(s_wallace_rca24_and_13_1));
  fa fa_s_wallace_rca24_fa11_out(.a(s_wallace_rca24_fa10_or0[0]), .b(s_wallace_rca24_and_14_0[0]), .cin(s_wallace_rca24_and_13_1[0]), .fa_xor1(s_wallace_rca24_fa11_xor1), .fa_or0(s_wallace_rca24_fa11_or0));
  and_gate and_gate_s_wallace_rca24_and_15_0(.a(a[15]), .b(b[0]), .out(s_wallace_rca24_and_15_0));
  and_gate and_gate_s_wallace_rca24_and_14_1(.a(a[14]), .b(b[1]), .out(s_wallace_rca24_and_14_1));
  fa fa_s_wallace_rca24_fa12_out(.a(s_wallace_rca24_fa11_or0[0]), .b(s_wallace_rca24_and_15_0[0]), .cin(s_wallace_rca24_and_14_1[0]), .fa_xor1(s_wallace_rca24_fa12_xor1), .fa_or0(s_wallace_rca24_fa12_or0));
  and_gate and_gate_s_wallace_rca24_and_16_0(.a(a[16]), .b(b[0]), .out(s_wallace_rca24_and_16_0));
  and_gate and_gate_s_wallace_rca24_and_15_1(.a(a[15]), .b(b[1]), .out(s_wallace_rca24_and_15_1));
  fa fa_s_wallace_rca24_fa13_out(.a(s_wallace_rca24_fa12_or0[0]), .b(s_wallace_rca24_and_16_0[0]), .cin(s_wallace_rca24_and_15_1[0]), .fa_xor1(s_wallace_rca24_fa13_xor1), .fa_or0(s_wallace_rca24_fa13_or0));
  and_gate and_gate_s_wallace_rca24_and_17_0(.a(a[17]), .b(b[0]), .out(s_wallace_rca24_and_17_0));
  and_gate and_gate_s_wallace_rca24_and_16_1(.a(a[16]), .b(b[1]), .out(s_wallace_rca24_and_16_1));
  fa fa_s_wallace_rca24_fa14_out(.a(s_wallace_rca24_fa13_or0[0]), .b(s_wallace_rca24_and_17_0[0]), .cin(s_wallace_rca24_and_16_1[0]), .fa_xor1(s_wallace_rca24_fa14_xor1), .fa_or0(s_wallace_rca24_fa14_or0));
  and_gate and_gate_s_wallace_rca24_and_18_0(.a(a[18]), .b(b[0]), .out(s_wallace_rca24_and_18_0));
  and_gate and_gate_s_wallace_rca24_and_17_1(.a(a[17]), .b(b[1]), .out(s_wallace_rca24_and_17_1));
  fa fa_s_wallace_rca24_fa15_out(.a(s_wallace_rca24_fa14_or0[0]), .b(s_wallace_rca24_and_18_0[0]), .cin(s_wallace_rca24_and_17_1[0]), .fa_xor1(s_wallace_rca24_fa15_xor1), .fa_or0(s_wallace_rca24_fa15_or0));
  and_gate and_gate_s_wallace_rca24_and_19_0(.a(a[19]), .b(b[0]), .out(s_wallace_rca24_and_19_0));
  and_gate and_gate_s_wallace_rca24_and_18_1(.a(a[18]), .b(b[1]), .out(s_wallace_rca24_and_18_1));
  fa fa_s_wallace_rca24_fa16_out(.a(s_wallace_rca24_fa15_or0[0]), .b(s_wallace_rca24_and_19_0[0]), .cin(s_wallace_rca24_and_18_1[0]), .fa_xor1(s_wallace_rca24_fa16_xor1), .fa_or0(s_wallace_rca24_fa16_or0));
  and_gate and_gate_s_wallace_rca24_and_20_0(.a(a[20]), .b(b[0]), .out(s_wallace_rca24_and_20_0));
  and_gate and_gate_s_wallace_rca24_and_19_1(.a(a[19]), .b(b[1]), .out(s_wallace_rca24_and_19_1));
  fa fa_s_wallace_rca24_fa17_out(.a(s_wallace_rca24_fa16_or0[0]), .b(s_wallace_rca24_and_20_0[0]), .cin(s_wallace_rca24_and_19_1[0]), .fa_xor1(s_wallace_rca24_fa17_xor1), .fa_or0(s_wallace_rca24_fa17_or0));
  and_gate and_gate_s_wallace_rca24_and_21_0(.a(a[21]), .b(b[0]), .out(s_wallace_rca24_and_21_0));
  and_gate and_gate_s_wallace_rca24_and_20_1(.a(a[20]), .b(b[1]), .out(s_wallace_rca24_and_20_1));
  fa fa_s_wallace_rca24_fa18_out(.a(s_wallace_rca24_fa17_or0[0]), .b(s_wallace_rca24_and_21_0[0]), .cin(s_wallace_rca24_and_20_1[0]), .fa_xor1(s_wallace_rca24_fa18_xor1), .fa_or0(s_wallace_rca24_fa18_or0));
  and_gate and_gate_s_wallace_rca24_and_22_0(.a(a[22]), .b(b[0]), .out(s_wallace_rca24_and_22_0));
  and_gate and_gate_s_wallace_rca24_and_21_1(.a(a[21]), .b(b[1]), .out(s_wallace_rca24_and_21_1));
  fa fa_s_wallace_rca24_fa19_out(.a(s_wallace_rca24_fa18_or0[0]), .b(s_wallace_rca24_and_22_0[0]), .cin(s_wallace_rca24_and_21_1[0]), .fa_xor1(s_wallace_rca24_fa19_xor1), .fa_or0(s_wallace_rca24_fa19_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_0(.a(a[23]), .b(b[0]), .out(s_wallace_rca24_nand_23_0));
  and_gate and_gate_s_wallace_rca24_and_22_1(.a(a[22]), .b(b[1]), .out(s_wallace_rca24_and_22_1));
  fa fa_s_wallace_rca24_fa20_out(.a(s_wallace_rca24_fa19_or0[0]), .b(s_wallace_rca24_nand_23_0[0]), .cin(s_wallace_rca24_and_22_1[0]), .fa_xor1(s_wallace_rca24_fa20_xor1), .fa_or0(s_wallace_rca24_fa20_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_1(.a(a[23]), .b(b[1]), .out(s_wallace_rca24_nand_23_1));
  fa fa_s_wallace_rca24_fa21_out(.a(s_wallace_rca24_fa20_or0[0]), .b(1'b1), .cin(s_wallace_rca24_nand_23_1[0]), .fa_xor1(s_wallace_rca24_fa21_xor1), .fa_or0(s_wallace_rca24_fa21_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_2(.a(a[23]), .b(b[2]), .out(s_wallace_rca24_nand_23_2));
  and_gate and_gate_s_wallace_rca24_and_22_3(.a(a[22]), .b(b[3]), .out(s_wallace_rca24_and_22_3));
  fa fa_s_wallace_rca24_fa22_out(.a(s_wallace_rca24_fa21_or0[0]), .b(s_wallace_rca24_nand_23_2[0]), .cin(s_wallace_rca24_and_22_3[0]), .fa_xor1(s_wallace_rca24_fa22_xor1), .fa_or0(s_wallace_rca24_fa22_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_3(.a(a[23]), .b(b[3]), .out(s_wallace_rca24_nand_23_3));
  and_gate and_gate_s_wallace_rca24_and_22_4(.a(a[22]), .b(b[4]), .out(s_wallace_rca24_and_22_4));
  fa fa_s_wallace_rca24_fa23_out(.a(s_wallace_rca24_fa22_or0[0]), .b(s_wallace_rca24_nand_23_3[0]), .cin(s_wallace_rca24_and_22_4[0]), .fa_xor1(s_wallace_rca24_fa23_xor1), .fa_or0(s_wallace_rca24_fa23_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_4(.a(a[23]), .b(b[4]), .out(s_wallace_rca24_nand_23_4));
  and_gate and_gate_s_wallace_rca24_and_22_5(.a(a[22]), .b(b[5]), .out(s_wallace_rca24_and_22_5));
  fa fa_s_wallace_rca24_fa24_out(.a(s_wallace_rca24_fa23_or0[0]), .b(s_wallace_rca24_nand_23_4[0]), .cin(s_wallace_rca24_and_22_5[0]), .fa_xor1(s_wallace_rca24_fa24_xor1), .fa_or0(s_wallace_rca24_fa24_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_5(.a(a[23]), .b(b[5]), .out(s_wallace_rca24_nand_23_5));
  and_gate and_gate_s_wallace_rca24_and_22_6(.a(a[22]), .b(b[6]), .out(s_wallace_rca24_and_22_6));
  fa fa_s_wallace_rca24_fa25_out(.a(s_wallace_rca24_fa24_or0[0]), .b(s_wallace_rca24_nand_23_5[0]), .cin(s_wallace_rca24_and_22_6[0]), .fa_xor1(s_wallace_rca24_fa25_xor1), .fa_or0(s_wallace_rca24_fa25_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_6(.a(a[23]), .b(b[6]), .out(s_wallace_rca24_nand_23_6));
  and_gate and_gate_s_wallace_rca24_and_22_7(.a(a[22]), .b(b[7]), .out(s_wallace_rca24_and_22_7));
  fa fa_s_wallace_rca24_fa26_out(.a(s_wallace_rca24_fa25_or0[0]), .b(s_wallace_rca24_nand_23_6[0]), .cin(s_wallace_rca24_and_22_7[0]), .fa_xor1(s_wallace_rca24_fa26_xor1), .fa_or0(s_wallace_rca24_fa26_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_7(.a(a[23]), .b(b[7]), .out(s_wallace_rca24_nand_23_7));
  and_gate and_gate_s_wallace_rca24_and_22_8(.a(a[22]), .b(b[8]), .out(s_wallace_rca24_and_22_8));
  fa fa_s_wallace_rca24_fa27_out(.a(s_wallace_rca24_fa26_or0[0]), .b(s_wallace_rca24_nand_23_7[0]), .cin(s_wallace_rca24_and_22_8[0]), .fa_xor1(s_wallace_rca24_fa27_xor1), .fa_or0(s_wallace_rca24_fa27_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_8(.a(a[23]), .b(b[8]), .out(s_wallace_rca24_nand_23_8));
  and_gate and_gate_s_wallace_rca24_and_22_9(.a(a[22]), .b(b[9]), .out(s_wallace_rca24_and_22_9));
  fa fa_s_wallace_rca24_fa28_out(.a(s_wallace_rca24_fa27_or0[0]), .b(s_wallace_rca24_nand_23_8[0]), .cin(s_wallace_rca24_and_22_9[0]), .fa_xor1(s_wallace_rca24_fa28_xor1), .fa_or0(s_wallace_rca24_fa28_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_9(.a(a[23]), .b(b[9]), .out(s_wallace_rca24_nand_23_9));
  and_gate and_gate_s_wallace_rca24_and_22_10(.a(a[22]), .b(b[10]), .out(s_wallace_rca24_and_22_10));
  fa fa_s_wallace_rca24_fa29_out(.a(s_wallace_rca24_fa28_or0[0]), .b(s_wallace_rca24_nand_23_9[0]), .cin(s_wallace_rca24_and_22_10[0]), .fa_xor1(s_wallace_rca24_fa29_xor1), .fa_or0(s_wallace_rca24_fa29_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_10(.a(a[23]), .b(b[10]), .out(s_wallace_rca24_nand_23_10));
  and_gate and_gate_s_wallace_rca24_and_22_11(.a(a[22]), .b(b[11]), .out(s_wallace_rca24_and_22_11));
  fa fa_s_wallace_rca24_fa30_out(.a(s_wallace_rca24_fa29_or0[0]), .b(s_wallace_rca24_nand_23_10[0]), .cin(s_wallace_rca24_and_22_11[0]), .fa_xor1(s_wallace_rca24_fa30_xor1), .fa_or0(s_wallace_rca24_fa30_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_11(.a(a[23]), .b(b[11]), .out(s_wallace_rca24_nand_23_11));
  and_gate and_gate_s_wallace_rca24_and_22_12(.a(a[22]), .b(b[12]), .out(s_wallace_rca24_and_22_12));
  fa fa_s_wallace_rca24_fa31_out(.a(s_wallace_rca24_fa30_or0[0]), .b(s_wallace_rca24_nand_23_11[0]), .cin(s_wallace_rca24_and_22_12[0]), .fa_xor1(s_wallace_rca24_fa31_xor1), .fa_or0(s_wallace_rca24_fa31_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_12(.a(a[23]), .b(b[12]), .out(s_wallace_rca24_nand_23_12));
  and_gate and_gate_s_wallace_rca24_and_22_13(.a(a[22]), .b(b[13]), .out(s_wallace_rca24_and_22_13));
  fa fa_s_wallace_rca24_fa32_out(.a(s_wallace_rca24_fa31_or0[0]), .b(s_wallace_rca24_nand_23_12[0]), .cin(s_wallace_rca24_and_22_13[0]), .fa_xor1(s_wallace_rca24_fa32_xor1), .fa_or0(s_wallace_rca24_fa32_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_13(.a(a[23]), .b(b[13]), .out(s_wallace_rca24_nand_23_13));
  and_gate and_gate_s_wallace_rca24_and_22_14(.a(a[22]), .b(b[14]), .out(s_wallace_rca24_and_22_14));
  fa fa_s_wallace_rca24_fa33_out(.a(s_wallace_rca24_fa32_or0[0]), .b(s_wallace_rca24_nand_23_13[0]), .cin(s_wallace_rca24_and_22_14[0]), .fa_xor1(s_wallace_rca24_fa33_xor1), .fa_or0(s_wallace_rca24_fa33_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_14(.a(a[23]), .b(b[14]), .out(s_wallace_rca24_nand_23_14));
  and_gate and_gate_s_wallace_rca24_and_22_15(.a(a[22]), .b(b[15]), .out(s_wallace_rca24_and_22_15));
  fa fa_s_wallace_rca24_fa34_out(.a(s_wallace_rca24_fa33_or0[0]), .b(s_wallace_rca24_nand_23_14[0]), .cin(s_wallace_rca24_and_22_15[0]), .fa_xor1(s_wallace_rca24_fa34_xor1), .fa_or0(s_wallace_rca24_fa34_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_15(.a(a[23]), .b(b[15]), .out(s_wallace_rca24_nand_23_15));
  and_gate and_gate_s_wallace_rca24_and_22_16(.a(a[22]), .b(b[16]), .out(s_wallace_rca24_and_22_16));
  fa fa_s_wallace_rca24_fa35_out(.a(s_wallace_rca24_fa34_or0[0]), .b(s_wallace_rca24_nand_23_15[0]), .cin(s_wallace_rca24_and_22_16[0]), .fa_xor1(s_wallace_rca24_fa35_xor1), .fa_or0(s_wallace_rca24_fa35_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_16(.a(a[23]), .b(b[16]), .out(s_wallace_rca24_nand_23_16));
  and_gate and_gate_s_wallace_rca24_and_22_17(.a(a[22]), .b(b[17]), .out(s_wallace_rca24_and_22_17));
  fa fa_s_wallace_rca24_fa36_out(.a(s_wallace_rca24_fa35_or0[0]), .b(s_wallace_rca24_nand_23_16[0]), .cin(s_wallace_rca24_and_22_17[0]), .fa_xor1(s_wallace_rca24_fa36_xor1), .fa_or0(s_wallace_rca24_fa36_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_17(.a(a[23]), .b(b[17]), .out(s_wallace_rca24_nand_23_17));
  and_gate and_gate_s_wallace_rca24_and_22_18(.a(a[22]), .b(b[18]), .out(s_wallace_rca24_and_22_18));
  fa fa_s_wallace_rca24_fa37_out(.a(s_wallace_rca24_fa36_or0[0]), .b(s_wallace_rca24_nand_23_17[0]), .cin(s_wallace_rca24_and_22_18[0]), .fa_xor1(s_wallace_rca24_fa37_xor1), .fa_or0(s_wallace_rca24_fa37_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_18(.a(a[23]), .b(b[18]), .out(s_wallace_rca24_nand_23_18));
  and_gate and_gate_s_wallace_rca24_and_22_19(.a(a[22]), .b(b[19]), .out(s_wallace_rca24_and_22_19));
  fa fa_s_wallace_rca24_fa38_out(.a(s_wallace_rca24_fa37_or0[0]), .b(s_wallace_rca24_nand_23_18[0]), .cin(s_wallace_rca24_and_22_19[0]), .fa_xor1(s_wallace_rca24_fa38_xor1), .fa_or0(s_wallace_rca24_fa38_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_19(.a(a[23]), .b(b[19]), .out(s_wallace_rca24_nand_23_19));
  and_gate and_gate_s_wallace_rca24_and_22_20(.a(a[22]), .b(b[20]), .out(s_wallace_rca24_and_22_20));
  fa fa_s_wallace_rca24_fa39_out(.a(s_wallace_rca24_fa38_or0[0]), .b(s_wallace_rca24_nand_23_19[0]), .cin(s_wallace_rca24_and_22_20[0]), .fa_xor1(s_wallace_rca24_fa39_xor1), .fa_or0(s_wallace_rca24_fa39_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_20(.a(a[23]), .b(b[20]), .out(s_wallace_rca24_nand_23_20));
  and_gate and_gate_s_wallace_rca24_and_22_21(.a(a[22]), .b(b[21]), .out(s_wallace_rca24_and_22_21));
  fa fa_s_wallace_rca24_fa40_out(.a(s_wallace_rca24_fa39_or0[0]), .b(s_wallace_rca24_nand_23_20[0]), .cin(s_wallace_rca24_and_22_21[0]), .fa_xor1(s_wallace_rca24_fa40_xor1), .fa_or0(s_wallace_rca24_fa40_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_21(.a(a[23]), .b(b[21]), .out(s_wallace_rca24_nand_23_21));
  and_gate and_gate_s_wallace_rca24_and_22_22(.a(a[22]), .b(b[22]), .out(s_wallace_rca24_and_22_22));
  fa fa_s_wallace_rca24_fa41_out(.a(s_wallace_rca24_fa40_or0[0]), .b(s_wallace_rca24_nand_23_21[0]), .cin(s_wallace_rca24_and_22_22[0]), .fa_xor1(s_wallace_rca24_fa41_xor1), .fa_or0(s_wallace_rca24_fa41_or0));
  and_gate and_gate_s_wallace_rca24_and_1_2(.a(a[1]), .b(b[2]), .out(s_wallace_rca24_and_1_2));
  and_gate and_gate_s_wallace_rca24_and_0_3(.a(a[0]), .b(b[3]), .out(s_wallace_rca24_and_0_3));
  ha ha_s_wallace_rca24_ha1_out(.a(s_wallace_rca24_and_1_2[0]), .b(s_wallace_rca24_and_0_3[0]), .ha_xor0(s_wallace_rca24_ha1_xor0), .ha_and0(s_wallace_rca24_ha1_and0));
  and_gate and_gate_s_wallace_rca24_and_2_2(.a(a[2]), .b(b[2]), .out(s_wallace_rca24_and_2_2));
  and_gate and_gate_s_wallace_rca24_and_1_3(.a(a[1]), .b(b[3]), .out(s_wallace_rca24_and_1_3));
  fa fa_s_wallace_rca24_fa42_out(.a(s_wallace_rca24_ha1_and0[0]), .b(s_wallace_rca24_and_2_2[0]), .cin(s_wallace_rca24_and_1_3[0]), .fa_xor1(s_wallace_rca24_fa42_xor1), .fa_or0(s_wallace_rca24_fa42_or0));
  and_gate and_gate_s_wallace_rca24_and_3_2(.a(a[3]), .b(b[2]), .out(s_wallace_rca24_and_3_2));
  and_gate and_gate_s_wallace_rca24_and_2_3(.a(a[2]), .b(b[3]), .out(s_wallace_rca24_and_2_3));
  fa fa_s_wallace_rca24_fa43_out(.a(s_wallace_rca24_fa42_or0[0]), .b(s_wallace_rca24_and_3_2[0]), .cin(s_wallace_rca24_and_2_3[0]), .fa_xor1(s_wallace_rca24_fa43_xor1), .fa_or0(s_wallace_rca24_fa43_or0));
  and_gate and_gate_s_wallace_rca24_and_4_2(.a(a[4]), .b(b[2]), .out(s_wallace_rca24_and_4_2));
  and_gate and_gate_s_wallace_rca24_and_3_3(.a(a[3]), .b(b[3]), .out(s_wallace_rca24_and_3_3));
  fa fa_s_wallace_rca24_fa44_out(.a(s_wallace_rca24_fa43_or0[0]), .b(s_wallace_rca24_and_4_2[0]), .cin(s_wallace_rca24_and_3_3[0]), .fa_xor1(s_wallace_rca24_fa44_xor1), .fa_or0(s_wallace_rca24_fa44_or0));
  and_gate and_gate_s_wallace_rca24_and_5_2(.a(a[5]), .b(b[2]), .out(s_wallace_rca24_and_5_2));
  and_gate and_gate_s_wallace_rca24_and_4_3(.a(a[4]), .b(b[3]), .out(s_wallace_rca24_and_4_3));
  fa fa_s_wallace_rca24_fa45_out(.a(s_wallace_rca24_fa44_or0[0]), .b(s_wallace_rca24_and_5_2[0]), .cin(s_wallace_rca24_and_4_3[0]), .fa_xor1(s_wallace_rca24_fa45_xor1), .fa_or0(s_wallace_rca24_fa45_or0));
  and_gate and_gate_s_wallace_rca24_and_6_2(.a(a[6]), .b(b[2]), .out(s_wallace_rca24_and_6_2));
  and_gate and_gate_s_wallace_rca24_and_5_3(.a(a[5]), .b(b[3]), .out(s_wallace_rca24_and_5_3));
  fa fa_s_wallace_rca24_fa46_out(.a(s_wallace_rca24_fa45_or0[0]), .b(s_wallace_rca24_and_6_2[0]), .cin(s_wallace_rca24_and_5_3[0]), .fa_xor1(s_wallace_rca24_fa46_xor1), .fa_or0(s_wallace_rca24_fa46_or0));
  and_gate and_gate_s_wallace_rca24_and_7_2(.a(a[7]), .b(b[2]), .out(s_wallace_rca24_and_7_2));
  and_gate and_gate_s_wallace_rca24_and_6_3(.a(a[6]), .b(b[3]), .out(s_wallace_rca24_and_6_3));
  fa fa_s_wallace_rca24_fa47_out(.a(s_wallace_rca24_fa46_or0[0]), .b(s_wallace_rca24_and_7_2[0]), .cin(s_wallace_rca24_and_6_3[0]), .fa_xor1(s_wallace_rca24_fa47_xor1), .fa_or0(s_wallace_rca24_fa47_or0));
  and_gate and_gate_s_wallace_rca24_and_8_2(.a(a[8]), .b(b[2]), .out(s_wallace_rca24_and_8_2));
  and_gate and_gate_s_wallace_rca24_and_7_3(.a(a[7]), .b(b[3]), .out(s_wallace_rca24_and_7_3));
  fa fa_s_wallace_rca24_fa48_out(.a(s_wallace_rca24_fa47_or0[0]), .b(s_wallace_rca24_and_8_2[0]), .cin(s_wallace_rca24_and_7_3[0]), .fa_xor1(s_wallace_rca24_fa48_xor1), .fa_or0(s_wallace_rca24_fa48_or0));
  and_gate and_gate_s_wallace_rca24_and_9_2(.a(a[9]), .b(b[2]), .out(s_wallace_rca24_and_9_2));
  and_gate and_gate_s_wallace_rca24_and_8_3(.a(a[8]), .b(b[3]), .out(s_wallace_rca24_and_8_3));
  fa fa_s_wallace_rca24_fa49_out(.a(s_wallace_rca24_fa48_or0[0]), .b(s_wallace_rca24_and_9_2[0]), .cin(s_wallace_rca24_and_8_3[0]), .fa_xor1(s_wallace_rca24_fa49_xor1), .fa_or0(s_wallace_rca24_fa49_or0));
  and_gate and_gate_s_wallace_rca24_and_10_2(.a(a[10]), .b(b[2]), .out(s_wallace_rca24_and_10_2));
  and_gate and_gate_s_wallace_rca24_and_9_3(.a(a[9]), .b(b[3]), .out(s_wallace_rca24_and_9_3));
  fa fa_s_wallace_rca24_fa50_out(.a(s_wallace_rca24_fa49_or0[0]), .b(s_wallace_rca24_and_10_2[0]), .cin(s_wallace_rca24_and_9_3[0]), .fa_xor1(s_wallace_rca24_fa50_xor1), .fa_or0(s_wallace_rca24_fa50_or0));
  and_gate and_gate_s_wallace_rca24_and_11_2(.a(a[11]), .b(b[2]), .out(s_wallace_rca24_and_11_2));
  and_gate and_gate_s_wallace_rca24_and_10_3(.a(a[10]), .b(b[3]), .out(s_wallace_rca24_and_10_3));
  fa fa_s_wallace_rca24_fa51_out(.a(s_wallace_rca24_fa50_or0[0]), .b(s_wallace_rca24_and_11_2[0]), .cin(s_wallace_rca24_and_10_3[0]), .fa_xor1(s_wallace_rca24_fa51_xor1), .fa_or0(s_wallace_rca24_fa51_or0));
  and_gate and_gate_s_wallace_rca24_and_12_2(.a(a[12]), .b(b[2]), .out(s_wallace_rca24_and_12_2));
  and_gate and_gate_s_wallace_rca24_and_11_3(.a(a[11]), .b(b[3]), .out(s_wallace_rca24_and_11_3));
  fa fa_s_wallace_rca24_fa52_out(.a(s_wallace_rca24_fa51_or0[0]), .b(s_wallace_rca24_and_12_2[0]), .cin(s_wallace_rca24_and_11_3[0]), .fa_xor1(s_wallace_rca24_fa52_xor1), .fa_or0(s_wallace_rca24_fa52_or0));
  and_gate and_gate_s_wallace_rca24_and_13_2(.a(a[13]), .b(b[2]), .out(s_wallace_rca24_and_13_2));
  and_gate and_gate_s_wallace_rca24_and_12_3(.a(a[12]), .b(b[3]), .out(s_wallace_rca24_and_12_3));
  fa fa_s_wallace_rca24_fa53_out(.a(s_wallace_rca24_fa52_or0[0]), .b(s_wallace_rca24_and_13_2[0]), .cin(s_wallace_rca24_and_12_3[0]), .fa_xor1(s_wallace_rca24_fa53_xor1), .fa_or0(s_wallace_rca24_fa53_or0));
  and_gate and_gate_s_wallace_rca24_and_14_2(.a(a[14]), .b(b[2]), .out(s_wallace_rca24_and_14_2));
  and_gate and_gate_s_wallace_rca24_and_13_3(.a(a[13]), .b(b[3]), .out(s_wallace_rca24_and_13_3));
  fa fa_s_wallace_rca24_fa54_out(.a(s_wallace_rca24_fa53_or0[0]), .b(s_wallace_rca24_and_14_2[0]), .cin(s_wallace_rca24_and_13_3[0]), .fa_xor1(s_wallace_rca24_fa54_xor1), .fa_or0(s_wallace_rca24_fa54_or0));
  and_gate and_gate_s_wallace_rca24_and_15_2(.a(a[15]), .b(b[2]), .out(s_wallace_rca24_and_15_2));
  and_gate and_gate_s_wallace_rca24_and_14_3(.a(a[14]), .b(b[3]), .out(s_wallace_rca24_and_14_3));
  fa fa_s_wallace_rca24_fa55_out(.a(s_wallace_rca24_fa54_or0[0]), .b(s_wallace_rca24_and_15_2[0]), .cin(s_wallace_rca24_and_14_3[0]), .fa_xor1(s_wallace_rca24_fa55_xor1), .fa_or0(s_wallace_rca24_fa55_or0));
  and_gate and_gate_s_wallace_rca24_and_16_2(.a(a[16]), .b(b[2]), .out(s_wallace_rca24_and_16_2));
  and_gate and_gate_s_wallace_rca24_and_15_3(.a(a[15]), .b(b[3]), .out(s_wallace_rca24_and_15_3));
  fa fa_s_wallace_rca24_fa56_out(.a(s_wallace_rca24_fa55_or0[0]), .b(s_wallace_rca24_and_16_2[0]), .cin(s_wallace_rca24_and_15_3[0]), .fa_xor1(s_wallace_rca24_fa56_xor1), .fa_or0(s_wallace_rca24_fa56_or0));
  and_gate and_gate_s_wallace_rca24_and_17_2(.a(a[17]), .b(b[2]), .out(s_wallace_rca24_and_17_2));
  and_gate and_gate_s_wallace_rca24_and_16_3(.a(a[16]), .b(b[3]), .out(s_wallace_rca24_and_16_3));
  fa fa_s_wallace_rca24_fa57_out(.a(s_wallace_rca24_fa56_or0[0]), .b(s_wallace_rca24_and_17_2[0]), .cin(s_wallace_rca24_and_16_3[0]), .fa_xor1(s_wallace_rca24_fa57_xor1), .fa_or0(s_wallace_rca24_fa57_or0));
  and_gate and_gate_s_wallace_rca24_and_18_2(.a(a[18]), .b(b[2]), .out(s_wallace_rca24_and_18_2));
  and_gate and_gate_s_wallace_rca24_and_17_3(.a(a[17]), .b(b[3]), .out(s_wallace_rca24_and_17_3));
  fa fa_s_wallace_rca24_fa58_out(.a(s_wallace_rca24_fa57_or0[0]), .b(s_wallace_rca24_and_18_2[0]), .cin(s_wallace_rca24_and_17_3[0]), .fa_xor1(s_wallace_rca24_fa58_xor1), .fa_or0(s_wallace_rca24_fa58_or0));
  and_gate and_gate_s_wallace_rca24_and_19_2(.a(a[19]), .b(b[2]), .out(s_wallace_rca24_and_19_2));
  and_gate and_gate_s_wallace_rca24_and_18_3(.a(a[18]), .b(b[3]), .out(s_wallace_rca24_and_18_3));
  fa fa_s_wallace_rca24_fa59_out(.a(s_wallace_rca24_fa58_or0[0]), .b(s_wallace_rca24_and_19_2[0]), .cin(s_wallace_rca24_and_18_3[0]), .fa_xor1(s_wallace_rca24_fa59_xor1), .fa_or0(s_wallace_rca24_fa59_or0));
  and_gate and_gate_s_wallace_rca24_and_20_2(.a(a[20]), .b(b[2]), .out(s_wallace_rca24_and_20_2));
  and_gate and_gate_s_wallace_rca24_and_19_3(.a(a[19]), .b(b[3]), .out(s_wallace_rca24_and_19_3));
  fa fa_s_wallace_rca24_fa60_out(.a(s_wallace_rca24_fa59_or0[0]), .b(s_wallace_rca24_and_20_2[0]), .cin(s_wallace_rca24_and_19_3[0]), .fa_xor1(s_wallace_rca24_fa60_xor1), .fa_or0(s_wallace_rca24_fa60_or0));
  and_gate and_gate_s_wallace_rca24_and_21_2(.a(a[21]), .b(b[2]), .out(s_wallace_rca24_and_21_2));
  and_gate and_gate_s_wallace_rca24_and_20_3(.a(a[20]), .b(b[3]), .out(s_wallace_rca24_and_20_3));
  fa fa_s_wallace_rca24_fa61_out(.a(s_wallace_rca24_fa60_or0[0]), .b(s_wallace_rca24_and_21_2[0]), .cin(s_wallace_rca24_and_20_3[0]), .fa_xor1(s_wallace_rca24_fa61_xor1), .fa_or0(s_wallace_rca24_fa61_or0));
  and_gate and_gate_s_wallace_rca24_and_22_2(.a(a[22]), .b(b[2]), .out(s_wallace_rca24_and_22_2));
  and_gate and_gate_s_wallace_rca24_and_21_3(.a(a[21]), .b(b[3]), .out(s_wallace_rca24_and_21_3));
  fa fa_s_wallace_rca24_fa62_out(.a(s_wallace_rca24_fa61_or0[0]), .b(s_wallace_rca24_and_22_2[0]), .cin(s_wallace_rca24_and_21_3[0]), .fa_xor1(s_wallace_rca24_fa62_xor1), .fa_or0(s_wallace_rca24_fa62_or0));
  and_gate and_gate_s_wallace_rca24_and_21_4(.a(a[21]), .b(b[4]), .out(s_wallace_rca24_and_21_4));
  and_gate and_gate_s_wallace_rca24_and_20_5(.a(a[20]), .b(b[5]), .out(s_wallace_rca24_and_20_5));
  fa fa_s_wallace_rca24_fa63_out(.a(s_wallace_rca24_fa62_or0[0]), .b(s_wallace_rca24_and_21_4[0]), .cin(s_wallace_rca24_and_20_5[0]), .fa_xor1(s_wallace_rca24_fa63_xor1), .fa_or0(s_wallace_rca24_fa63_or0));
  and_gate and_gate_s_wallace_rca24_and_21_5(.a(a[21]), .b(b[5]), .out(s_wallace_rca24_and_21_5));
  and_gate and_gate_s_wallace_rca24_and_20_6(.a(a[20]), .b(b[6]), .out(s_wallace_rca24_and_20_6));
  fa fa_s_wallace_rca24_fa64_out(.a(s_wallace_rca24_fa63_or0[0]), .b(s_wallace_rca24_and_21_5[0]), .cin(s_wallace_rca24_and_20_6[0]), .fa_xor1(s_wallace_rca24_fa64_xor1), .fa_or0(s_wallace_rca24_fa64_or0));
  and_gate and_gate_s_wallace_rca24_and_21_6(.a(a[21]), .b(b[6]), .out(s_wallace_rca24_and_21_6));
  and_gate and_gate_s_wallace_rca24_and_20_7(.a(a[20]), .b(b[7]), .out(s_wallace_rca24_and_20_7));
  fa fa_s_wallace_rca24_fa65_out(.a(s_wallace_rca24_fa64_or0[0]), .b(s_wallace_rca24_and_21_6[0]), .cin(s_wallace_rca24_and_20_7[0]), .fa_xor1(s_wallace_rca24_fa65_xor1), .fa_or0(s_wallace_rca24_fa65_or0));
  and_gate and_gate_s_wallace_rca24_and_21_7(.a(a[21]), .b(b[7]), .out(s_wallace_rca24_and_21_7));
  and_gate and_gate_s_wallace_rca24_and_20_8(.a(a[20]), .b(b[8]), .out(s_wallace_rca24_and_20_8));
  fa fa_s_wallace_rca24_fa66_out(.a(s_wallace_rca24_fa65_or0[0]), .b(s_wallace_rca24_and_21_7[0]), .cin(s_wallace_rca24_and_20_8[0]), .fa_xor1(s_wallace_rca24_fa66_xor1), .fa_or0(s_wallace_rca24_fa66_or0));
  and_gate and_gate_s_wallace_rca24_and_21_8(.a(a[21]), .b(b[8]), .out(s_wallace_rca24_and_21_8));
  and_gate and_gate_s_wallace_rca24_and_20_9(.a(a[20]), .b(b[9]), .out(s_wallace_rca24_and_20_9));
  fa fa_s_wallace_rca24_fa67_out(.a(s_wallace_rca24_fa66_or0[0]), .b(s_wallace_rca24_and_21_8[0]), .cin(s_wallace_rca24_and_20_9[0]), .fa_xor1(s_wallace_rca24_fa67_xor1), .fa_or0(s_wallace_rca24_fa67_or0));
  and_gate and_gate_s_wallace_rca24_and_21_9(.a(a[21]), .b(b[9]), .out(s_wallace_rca24_and_21_9));
  and_gate and_gate_s_wallace_rca24_and_20_10(.a(a[20]), .b(b[10]), .out(s_wallace_rca24_and_20_10));
  fa fa_s_wallace_rca24_fa68_out(.a(s_wallace_rca24_fa67_or0[0]), .b(s_wallace_rca24_and_21_9[0]), .cin(s_wallace_rca24_and_20_10[0]), .fa_xor1(s_wallace_rca24_fa68_xor1), .fa_or0(s_wallace_rca24_fa68_or0));
  and_gate and_gate_s_wallace_rca24_and_21_10(.a(a[21]), .b(b[10]), .out(s_wallace_rca24_and_21_10));
  and_gate and_gate_s_wallace_rca24_and_20_11(.a(a[20]), .b(b[11]), .out(s_wallace_rca24_and_20_11));
  fa fa_s_wallace_rca24_fa69_out(.a(s_wallace_rca24_fa68_or0[0]), .b(s_wallace_rca24_and_21_10[0]), .cin(s_wallace_rca24_and_20_11[0]), .fa_xor1(s_wallace_rca24_fa69_xor1), .fa_or0(s_wallace_rca24_fa69_or0));
  and_gate and_gate_s_wallace_rca24_and_21_11(.a(a[21]), .b(b[11]), .out(s_wallace_rca24_and_21_11));
  and_gate and_gate_s_wallace_rca24_and_20_12(.a(a[20]), .b(b[12]), .out(s_wallace_rca24_and_20_12));
  fa fa_s_wallace_rca24_fa70_out(.a(s_wallace_rca24_fa69_or0[0]), .b(s_wallace_rca24_and_21_11[0]), .cin(s_wallace_rca24_and_20_12[0]), .fa_xor1(s_wallace_rca24_fa70_xor1), .fa_or0(s_wallace_rca24_fa70_or0));
  and_gate and_gate_s_wallace_rca24_and_21_12(.a(a[21]), .b(b[12]), .out(s_wallace_rca24_and_21_12));
  and_gate and_gate_s_wallace_rca24_and_20_13(.a(a[20]), .b(b[13]), .out(s_wallace_rca24_and_20_13));
  fa fa_s_wallace_rca24_fa71_out(.a(s_wallace_rca24_fa70_or0[0]), .b(s_wallace_rca24_and_21_12[0]), .cin(s_wallace_rca24_and_20_13[0]), .fa_xor1(s_wallace_rca24_fa71_xor1), .fa_or0(s_wallace_rca24_fa71_or0));
  and_gate and_gate_s_wallace_rca24_and_21_13(.a(a[21]), .b(b[13]), .out(s_wallace_rca24_and_21_13));
  and_gate and_gate_s_wallace_rca24_and_20_14(.a(a[20]), .b(b[14]), .out(s_wallace_rca24_and_20_14));
  fa fa_s_wallace_rca24_fa72_out(.a(s_wallace_rca24_fa71_or0[0]), .b(s_wallace_rca24_and_21_13[0]), .cin(s_wallace_rca24_and_20_14[0]), .fa_xor1(s_wallace_rca24_fa72_xor1), .fa_or0(s_wallace_rca24_fa72_or0));
  and_gate and_gate_s_wallace_rca24_and_21_14(.a(a[21]), .b(b[14]), .out(s_wallace_rca24_and_21_14));
  and_gate and_gate_s_wallace_rca24_and_20_15(.a(a[20]), .b(b[15]), .out(s_wallace_rca24_and_20_15));
  fa fa_s_wallace_rca24_fa73_out(.a(s_wallace_rca24_fa72_or0[0]), .b(s_wallace_rca24_and_21_14[0]), .cin(s_wallace_rca24_and_20_15[0]), .fa_xor1(s_wallace_rca24_fa73_xor1), .fa_or0(s_wallace_rca24_fa73_or0));
  and_gate and_gate_s_wallace_rca24_and_21_15(.a(a[21]), .b(b[15]), .out(s_wallace_rca24_and_21_15));
  and_gate and_gate_s_wallace_rca24_and_20_16(.a(a[20]), .b(b[16]), .out(s_wallace_rca24_and_20_16));
  fa fa_s_wallace_rca24_fa74_out(.a(s_wallace_rca24_fa73_or0[0]), .b(s_wallace_rca24_and_21_15[0]), .cin(s_wallace_rca24_and_20_16[0]), .fa_xor1(s_wallace_rca24_fa74_xor1), .fa_or0(s_wallace_rca24_fa74_or0));
  and_gate and_gate_s_wallace_rca24_and_21_16(.a(a[21]), .b(b[16]), .out(s_wallace_rca24_and_21_16));
  and_gate and_gate_s_wallace_rca24_and_20_17(.a(a[20]), .b(b[17]), .out(s_wallace_rca24_and_20_17));
  fa fa_s_wallace_rca24_fa75_out(.a(s_wallace_rca24_fa74_or0[0]), .b(s_wallace_rca24_and_21_16[0]), .cin(s_wallace_rca24_and_20_17[0]), .fa_xor1(s_wallace_rca24_fa75_xor1), .fa_or0(s_wallace_rca24_fa75_or0));
  and_gate and_gate_s_wallace_rca24_and_21_17(.a(a[21]), .b(b[17]), .out(s_wallace_rca24_and_21_17));
  and_gate and_gate_s_wallace_rca24_and_20_18(.a(a[20]), .b(b[18]), .out(s_wallace_rca24_and_20_18));
  fa fa_s_wallace_rca24_fa76_out(.a(s_wallace_rca24_fa75_or0[0]), .b(s_wallace_rca24_and_21_17[0]), .cin(s_wallace_rca24_and_20_18[0]), .fa_xor1(s_wallace_rca24_fa76_xor1), .fa_or0(s_wallace_rca24_fa76_or0));
  and_gate and_gate_s_wallace_rca24_and_21_18(.a(a[21]), .b(b[18]), .out(s_wallace_rca24_and_21_18));
  and_gate and_gate_s_wallace_rca24_and_20_19(.a(a[20]), .b(b[19]), .out(s_wallace_rca24_and_20_19));
  fa fa_s_wallace_rca24_fa77_out(.a(s_wallace_rca24_fa76_or0[0]), .b(s_wallace_rca24_and_21_18[0]), .cin(s_wallace_rca24_and_20_19[0]), .fa_xor1(s_wallace_rca24_fa77_xor1), .fa_or0(s_wallace_rca24_fa77_or0));
  and_gate and_gate_s_wallace_rca24_and_21_19(.a(a[21]), .b(b[19]), .out(s_wallace_rca24_and_21_19));
  and_gate and_gate_s_wallace_rca24_and_20_20(.a(a[20]), .b(b[20]), .out(s_wallace_rca24_and_20_20));
  fa fa_s_wallace_rca24_fa78_out(.a(s_wallace_rca24_fa77_or0[0]), .b(s_wallace_rca24_and_21_19[0]), .cin(s_wallace_rca24_and_20_20[0]), .fa_xor1(s_wallace_rca24_fa78_xor1), .fa_or0(s_wallace_rca24_fa78_or0));
  and_gate and_gate_s_wallace_rca24_and_21_20(.a(a[21]), .b(b[20]), .out(s_wallace_rca24_and_21_20));
  and_gate and_gate_s_wallace_rca24_and_20_21(.a(a[20]), .b(b[21]), .out(s_wallace_rca24_and_20_21));
  fa fa_s_wallace_rca24_fa79_out(.a(s_wallace_rca24_fa78_or0[0]), .b(s_wallace_rca24_and_21_20[0]), .cin(s_wallace_rca24_and_20_21[0]), .fa_xor1(s_wallace_rca24_fa79_xor1), .fa_or0(s_wallace_rca24_fa79_or0));
  and_gate and_gate_s_wallace_rca24_and_21_21(.a(a[21]), .b(b[21]), .out(s_wallace_rca24_and_21_21));
  and_gate and_gate_s_wallace_rca24_and_20_22(.a(a[20]), .b(b[22]), .out(s_wallace_rca24_and_20_22));
  fa fa_s_wallace_rca24_fa80_out(.a(s_wallace_rca24_fa79_or0[0]), .b(s_wallace_rca24_and_21_21[0]), .cin(s_wallace_rca24_and_20_22[0]), .fa_xor1(s_wallace_rca24_fa80_xor1), .fa_or0(s_wallace_rca24_fa80_or0));
  and_gate and_gate_s_wallace_rca24_and_21_22(.a(a[21]), .b(b[22]), .out(s_wallace_rca24_and_21_22));
  nand_gate nand_gate_s_wallace_rca24_nand_20_23(.a(a[20]), .b(b[23]), .out(s_wallace_rca24_nand_20_23));
  fa fa_s_wallace_rca24_fa81_out(.a(s_wallace_rca24_fa80_or0[0]), .b(s_wallace_rca24_and_21_22[0]), .cin(s_wallace_rca24_nand_20_23[0]), .fa_xor1(s_wallace_rca24_fa81_xor1), .fa_or0(s_wallace_rca24_fa81_or0));
  and_gate and_gate_s_wallace_rca24_and_0_4(.a(a[0]), .b(b[4]), .out(s_wallace_rca24_and_0_4));
  ha ha_s_wallace_rca24_ha2_out(.a(s_wallace_rca24_and_0_4[0]), .b(s_wallace_rca24_fa1_xor1[0]), .ha_xor0(s_wallace_rca24_ha2_xor0), .ha_and0(s_wallace_rca24_ha2_and0));
  and_gate and_gate_s_wallace_rca24_and_1_4(.a(a[1]), .b(b[4]), .out(s_wallace_rca24_and_1_4));
  and_gate and_gate_s_wallace_rca24_and_0_5(.a(a[0]), .b(b[5]), .out(s_wallace_rca24_and_0_5));
  fa fa_s_wallace_rca24_fa82_out(.a(s_wallace_rca24_ha2_and0[0]), .b(s_wallace_rca24_and_1_4[0]), .cin(s_wallace_rca24_and_0_5[0]), .fa_xor1(s_wallace_rca24_fa82_xor1), .fa_or0(s_wallace_rca24_fa82_or0));
  and_gate and_gate_s_wallace_rca24_and_2_4(.a(a[2]), .b(b[4]), .out(s_wallace_rca24_and_2_4));
  and_gate and_gate_s_wallace_rca24_and_1_5(.a(a[1]), .b(b[5]), .out(s_wallace_rca24_and_1_5));
  fa fa_s_wallace_rca24_fa83_out(.a(s_wallace_rca24_fa82_or0[0]), .b(s_wallace_rca24_and_2_4[0]), .cin(s_wallace_rca24_and_1_5[0]), .fa_xor1(s_wallace_rca24_fa83_xor1), .fa_or0(s_wallace_rca24_fa83_or0));
  and_gate and_gate_s_wallace_rca24_and_3_4(.a(a[3]), .b(b[4]), .out(s_wallace_rca24_and_3_4));
  and_gate and_gate_s_wallace_rca24_and_2_5(.a(a[2]), .b(b[5]), .out(s_wallace_rca24_and_2_5));
  fa fa_s_wallace_rca24_fa84_out(.a(s_wallace_rca24_fa83_or0[0]), .b(s_wallace_rca24_and_3_4[0]), .cin(s_wallace_rca24_and_2_5[0]), .fa_xor1(s_wallace_rca24_fa84_xor1), .fa_or0(s_wallace_rca24_fa84_or0));
  and_gate and_gate_s_wallace_rca24_and_4_4(.a(a[4]), .b(b[4]), .out(s_wallace_rca24_and_4_4));
  and_gate and_gate_s_wallace_rca24_and_3_5(.a(a[3]), .b(b[5]), .out(s_wallace_rca24_and_3_5));
  fa fa_s_wallace_rca24_fa85_out(.a(s_wallace_rca24_fa84_or0[0]), .b(s_wallace_rca24_and_4_4[0]), .cin(s_wallace_rca24_and_3_5[0]), .fa_xor1(s_wallace_rca24_fa85_xor1), .fa_or0(s_wallace_rca24_fa85_or0));
  and_gate and_gate_s_wallace_rca24_and_5_4(.a(a[5]), .b(b[4]), .out(s_wallace_rca24_and_5_4));
  and_gate and_gate_s_wallace_rca24_and_4_5(.a(a[4]), .b(b[5]), .out(s_wallace_rca24_and_4_5));
  fa fa_s_wallace_rca24_fa86_out(.a(s_wallace_rca24_fa85_or0[0]), .b(s_wallace_rca24_and_5_4[0]), .cin(s_wallace_rca24_and_4_5[0]), .fa_xor1(s_wallace_rca24_fa86_xor1), .fa_or0(s_wallace_rca24_fa86_or0));
  and_gate and_gate_s_wallace_rca24_and_6_4(.a(a[6]), .b(b[4]), .out(s_wallace_rca24_and_6_4));
  and_gate and_gate_s_wallace_rca24_and_5_5(.a(a[5]), .b(b[5]), .out(s_wallace_rca24_and_5_5));
  fa fa_s_wallace_rca24_fa87_out(.a(s_wallace_rca24_fa86_or0[0]), .b(s_wallace_rca24_and_6_4[0]), .cin(s_wallace_rca24_and_5_5[0]), .fa_xor1(s_wallace_rca24_fa87_xor1), .fa_or0(s_wallace_rca24_fa87_or0));
  and_gate and_gate_s_wallace_rca24_and_7_4(.a(a[7]), .b(b[4]), .out(s_wallace_rca24_and_7_4));
  and_gate and_gate_s_wallace_rca24_and_6_5(.a(a[6]), .b(b[5]), .out(s_wallace_rca24_and_6_5));
  fa fa_s_wallace_rca24_fa88_out(.a(s_wallace_rca24_fa87_or0[0]), .b(s_wallace_rca24_and_7_4[0]), .cin(s_wallace_rca24_and_6_5[0]), .fa_xor1(s_wallace_rca24_fa88_xor1), .fa_or0(s_wallace_rca24_fa88_or0));
  and_gate and_gate_s_wallace_rca24_and_8_4(.a(a[8]), .b(b[4]), .out(s_wallace_rca24_and_8_4));
  and_gate and_gate_s_wallace_rca24_and_7_5(.a(a[7]), .b(b[5]), .out(s_wallace_rca24_and_7_5));
  fa fa_s_wallace_rca24_fa89_out(.a(s_wallace_rca24_fa88_or0[0]), .b(s_wallace_rca24_and_8_4[0]), .cin(s_wallace_rca24_and_7_5[0]), .fa_xor1(s_wallace_rca24_fa89_xor1), .fa_or0(s_wallace_rca24_fa89_or0));
  and_gate and_gate_s_wallace_rca24_and_9_4(.a(a[9]), .b(b[4]), .out(s_wallace_rca24_and_9_4));
  and_gate and_gate_s_wallace_rca24_and_8_5(.a(a[8]), .b(b[5]), .out(s_wallace_rca24_and_8_5));
  fa fa_s_wallace_rca24_fa90_out(.a(s_wallace_rca24_fa89_or0[0]), .b(s_wallace_rca24_and_9_4[0]), .cin(s_wallace_rca24_and_8_5[0]), .fa_xor1(s_wallace_rca24_fa90_xor1), .fa_or0(s_wallace_rca24_fa90_or0));
  and_gate and_gate_s_wallace_rca24_and_10_4(.a(a[10]), .b(b[4]), .out(s_wallace_rca24_and_10_4));
  and_gate and_gate_s_wallace_rca24_and_9_5(.a(a[9]), .b(b[5]), .out(s_wallace_rca24_and_9_5));
  fa fa_s_wallace_rca24_fa91_out(.a(s_wallace_rca24_fa90_or0[0]), .b(s_wallace_rca24_and_10_4[0]), .cin(s_wallace_rca24_and_9_5[0]), .fa_xor1(s_wallace_rca24_fa91_xor1), .fa_or0(s_wallace_rca24_fa91_or0));
  and_gate and_gate_s_wallace_rca24_and_11_4(.a(a[11]), .b(b[4]), .out(s_wallace_rca24_and_11_4));
  and_gate and_gate_s_wallace_rca24_and_10_5(.a(a[10]), .b(b[5]), .out(s_wallace_rca24_and_10_5));
  fa fa_s_wallace_rca24_fa92_out(.a(s_wallace_rca24_fa91_or0[0]), .b(s_wallace_rca24_and_11_4[0]), .cin(s_wallace_rca24_and_10_5[0]), .fa_xor1(s_wallace_rca24_fa92_xor1), .fa_or0(s_wallace_rca24_fa92_or0));
  and_gate and_gate_s_wallace_rca24_and_12_4(.a(a[12]), .b(b[4]), .out(s_wallace_rca24_and_12_4));
  and_gate and_gate_s_wallace_rca24_and_11_5(.a(a[11]), .b(b[5]), .out(s_wallace_rca24_and_11_5));
  fa fa_s_wallace_rca24_fa93_out(.a(s_wallace_rca24_fa92_or0[0]), .b(s_wallace_rca24_and_12_4[0]), .cin(s_wallace_rca24_and_11_5[0]), .fa_xor1(s_wallace_rca24_fa93_xor1), .fa_or0(s_wallace_rca24_fa93_or0));
  and_gate and_gate_s_wallace_rca24_and_13_4(.a(a[13]), .b(b[4]), .out(s_wallace_rca24_and_13_4));
  and_gate and_gate_s_wallace_rca24_and_12_5(.a(a[12]), .b(b[5]), .out(s_wallace_rca24_and_12_5));
  fa fa_s_wallace_rca24_fa94_out(.a(s_wallace_rca24_fa93_or0[0]), .b(s_wallace_rca24_and_13_4[0]), .cin(s_wallace_rca24_and_12_5[0]), .fa_xor1(s_wallace_rca24_fa94_xor1), .fa_or0(s_wallace_rca24_fa94_or0));
  and_gate and_gate_s_wallace_rca24_and_14_4(.a(a[14]), .b(b[4]), .out(s_wallace_rca24_and_14_4));
  and_gate and_gate_s_wallace_rca24_and_13_5(.a(a[13]), .b(b[5]), .out(s_wallace_rca24_and_13_5));
  fa fa_s_wallace_rca24_fa95_out(.a(s_wallace_rca24_fa94_or0[0]), .b(s_wallace_rca24_and_14_4[0]), .cin(s_wallace_rca24_and_13_5[0]), .fa_xor1(s_wallace_rca24_fa95_xor1), .fa_or0(s_wallace_rca24_fa95_or0));
  and_gate and_gate_s_wallace_rca24_and_15_4(.a(a[15]), .b(b[4]), .out(s_wallace_rca24_and_15_4));
  and_gate and_gate_s_wallace_rca24_and_14_5(.a(a[14]), .b(b[5]), .out(s_wallace_rca24_and_14_5));
  fa fa_s_wallace_rca24_fa96_out(.a(s_wallace_rca24_fa95_or0[0]), .b(s_wallace_rca24_and_15_4[0]), .cin(s_wallace_rca24_and_14_5[0]), .fa_xor1(s_wallace_rca24_fa96_xor1), .fa_or0(s_wallace_rca24_fa96_or0));
  and_gate and_gate_s_wallace_rca24_and_16_4(.a(a[16]), .b(b[4]), .out(s_wallace_rca24_and_16_4));
  and_gate and_gate_s_wallace_rca24_and_15_5(.a(a[15]), .b(b[5]), .out(s_wallace_rca24_and_15_5));
  fa fa_s_wallace_rca24_fa97_out(.a(s_wallace_rca24_fa96_or0[0]), .b(s_wallace_rca24_and_16_4[0]), .cin(s_wallace_rca24_and_15_5[0]), .fa_xor1(s_wallace_rca24_fa97_xor1), .fa_or0(s_wallace_rca24_fa97_or0));
  and_gate and_gate_s_wallace_rca24_and_17_4(.a(a[17]), .b(b[4]), .out(s_wallace_rca24_and_17_4));
  and_gate and_gate_s_wallace_rca24_and_16_5(.a(a[16]), .b(b[5]), .out(s_wallace_rca24_and_16_5));
  fa fa_s_wallace_rca24_fa98_out(.a(s_wallace_rca24_fa97_or0[0]), .b(s_wallace_rca24_and_17_4[0]), .cin(s_wallace_rca24_and_16_5[0]), .fa_xor1(s_wallace_rca24_fa98_xor1), .fa_or0(s_wallace_rca24_fa98_or0));
  and_gate and_gate_s_wallace_rca24_and_18_4(.a(a[18]), .b(b[4]), .out(s_wallace_rca24_and_18_4));
  and_gate and_gate_s_wallace_rca24_and_17_5(.a(a[17]), .b(b[5]), .out(s_wallace_rca24_and_17_5));
  fa fa_s_wallace_rca24_fa99_out(.a(s_wallace_rca24_fa98_or0[0]), .b(s_wallace_rca24_and_18_4[0]), .cin(s_wallace_rca24_and_17_5[0]), .fa_xor1(s_wallace_rca24_fa99_xor1), .fa_or0(s_wallace_rca24_fa99_or0));
  and_gate and_gate_s_wallace_rca24_and_19_4(.a(a[19]), .b(b[4]), .out(s_wallace_rca24_and_19_4));
  and_gate and_gate_s_wallace_rca24_and_18_5(.a(a[18]), .b(b[5]), .out(s_wallace_rca24_and_18_5));
  fa fa_s_wallace_rca24_fa100_out(.a(s_wallace_rca24_fa99_or0[0]), .b(s_wallace_rca24_and_19_4[0]), .cin(s_wallace_rca24_and_18_5[0]), .fa_xor1(s_wallace_rca24_fa100_xor1), .fa_or0(s_wallace_rca24_fa100_or0));
  and_gate and_gate_s_wallace_rca24_and_20_4(.a(a[20]), .b(b[4]), .out(s_wallace_rca24_and_20_4));
  and_gate and_gate_s_wallace_rca24_and_19_5(.a(a[19]), .b(b[5]), .out(s_wallace_rca24_and_19_5));
  fa fa_s_wallace_rca24_fa101_out(.a(s_wallace_rca24_fa100_or0[0]), .b(s_wallace_rca24_and_20_4[0]), .cin(s_wallace_rca24_and_19_5[0]), .fa_xor1(s_wallace_rca24_fa101_xor1), .fa_or0(s_wallace_rca24_fa101_or0));
  and_gate and_gate_s_wallace_rca24_and_19_6(.a(a[19]), .b(b[6]), .out(s_wallace_rca24_and_19_6));
  and_gate and_gate_s_wallace_rca24_and_18_7(.a(a[18]), .b(b[7]), .out(s_wallace_rca24_and_18_7));
  fa fa_s_wallace_rca24_fa102_out(.a(s_wallace_rca24_fa101_or0[0]), .b(s_wallace_rca24_and_19_6[0]), .cin(s_wallace_rca24_and_18_7[0]), .fa_xor1(s_wallace_rca24_fa102_xor1), .fa_or0(s_wallace_rca24_fa102_or0));
  and_gate and_gate_s_wallace_rca24_and_19_7(.a(a[19]), .b(b[7]), .out(s_wallace_rca24_and_19_7));
  and_gate and_gate_s_wallace_rca24_and_18_8(.a(a[18]), .b(b[8]), .out(s_wallace_rca24_and_18_8));
  fa fa_s_wallace_rca24_fa103_out(.a(s_wallace_rca24_fa102_or0[0]), .b(s_wallace_rca24_and_19_7[0]), .cin(s_wallace_rca24_and_18_8[0]), .fa_xor1(s_wallace_rca24_fa103_xor1), .fa_or0(s_wallace_rca24_fa103_or0));
  and_gate and_gate_s_wallace_rca24_and_19_8(.a(a[19]), .b(b[8]), .out(s_wallace_rca24_and_19_8));
  and_gate and_gate_s_wallace_rca24_and_18_9(.a(a[18]), .b(b[9]), .out(s_wallace_rca24_and_18_9));
  fa fa_s_wallace_rca24_fa104_out(.a(s_wallace_rca24_fa103_or0[0]), .b(s_wallace_rca24_and_19_8[0]), .cin(s_wallace_rca24_and_18_9[0]), .fa_xor1(s_wallace_rca24_fa104_xor1), .fa_or0(s_wallace_rca24_fa104_or0));
  and_gate and_gate_s_wallace_rca24_and_19_9(.a(a[19]), .b(b[9]), .out(s_wallace_rca24_and_19_9));
  and_gate and_gate_s_wallace_rca24_and_18_10(.a(a[18]), .b(b[10]), .out(s_wallace_rca24_and_18_10));
  fa fa_s_wallace_rca24_fa105_out(.a(s_wallace_rca24_fa104_or0[0]), .b(s_wallace_rca24_and_19_9[0]), .cin(s_wallace_rca24_and_18_10[0]), .fa_xor1(s_wallace_rca24_fa105_xor1), .fa_or0(s_wallace_rca24_fa105_or0));
  and_gate and_gate_s_wallace_rca24_and_19_10(.a(a[19]), .b(b[10]), .out(s_wallace_rca24_and_19_10));
  and_gate and_gate_s_wallace_rca24_and_18_11(.a(a[18]), .b(b[11]), .out(s_wallace_rca24_and_18_11));
  fa fa_s_wallace_rca24_fa106_out(.a(s_wallace_rca24_fa105_or0[0]), .b(s_wallace_rca24_and_19_10[0]), .cin(s_wallace_rca24_and_18_11[0]), .fa_xor1(s_wallace_rca24_fa106_xor1), .fa_or0(s_wallace_rca24_fa106_or0));
  and_gate and_gate_s_wallace_rca24_and_19_11(.a(a[19]), .b(b[11]), .out(s_wallace_rca24_and_19_11));
  and_gate and_gate_s_wallace_rca24_and_18_12(.a(a[18]), .b(b[12]), .out(s_wallace_rca24_and_18_12));
  fa fa_s_wallace_rca24_fa107_out(.a(s_wallace_rca24_fa106_or0[0]), .b(s_wallace_rca24_and_19_11[0]), .cin(s_wallace_rca24_and_18_12[0]), .fa_xor1(s_wallace_rca24_fa107_xor1), .fa_or0(s_wallace_rca24_fa107_or0));
  and_gate and_gate_s_wallace_rca24_and_19_12(.a(a[19]), .b(b[12]), .out(s_wallace_rca24_and_19_12));
  and_gate and_gate_s_wallace_rca24_and_18_13(.a(a[18]), .b(b[13]), .out(s_wallace_rca24_and_18_13));
  fa fa_s_wallace_rca24_fa108_out(.a(s_wallace_rca24_fa107_or0[0]), .b(s_wallace_rca24_and_19_12[0]), .cin(s_wallace_rca24_and_18_13[0]), .fa_xor1(s_wallace_rca24_fa108_xor1), .fa_or0(s_wallace_rca24_fa108_or0));
  and_gate and_gate_s_wallace_rca24_and_19_13(.a(a[19]), .b(b[13]), .out(s_wallace_rca24_and_19_13));
  and_gate and_gate_s_wallace_rca24_and_18_14(.a(a[18]), .b(b[14]), .out(s_wallace_rca24_and_18_14));
  fa fa_s_wallace_rca24_fa109_out(.a(s_wallace_rca24_fa108_or0[0]), .b(s_wallace_rca24_and_19_13[0]), .cin(s_wallace_rca24_and_18_14[0]), .fa_xor1(s_wallace_rca24_fa109_xor1), .fa_or0(s_wallace_rca24_fa109_or0));
  and_gate and_gate_s_wallace_rca24_and_19_14(.a(a[19]), .b(b[14]), .out(s_wallace_rca24_and_19_14));
  and_gate and_gate_s_wallace_rca24_and_18_15(.a(a[18]), .b(b[15]), .out(s_wallace_rca24_and_18_15));
  fa fa_s_wallace_rca24_fa110_out(.a(s_wallace_rca24_fa109_or0[0]), .b(s_wallace_rca24_and_19_14[0]), .cin(s_wallace_rca24_and_18_15[0]), .fa_xor1(s_wallace_rca24_fa110_xor1), .fa_or0(s_wallace_rca24_fa110_or0));
  and_gate and_gate_s_wallace_rca24_and_19_15(.a(a[19]), .b(b[15]), .out(s_wallace_rca24_and_19_15));
  and_gate and_gate_s_wallace_rca24_and_18_16(.a(a[18]), .b(b[16]), .out(s_wallace_rca24_and_18_16));
  fa fa_s_wallace_rca24_fa111_out(.a(s_wallace_rca24_fa110_or0[0]), .b(s_wallace_rca24_and_19_15[0]), .cin(s_wallace_rca24_and_18_16[0]), .fa_xor1(s_wallace_rca24_fa111_xor1), .fa_or0(s_wallace_rca24_fa111_or0));
  and_gate and_gate_s_wallace_rca24_and_19_16(.a(a[19]), .b(b[16]), .out(s_wallace_rca24_and_19_16));
  and_gate and_gate_s_wallace_rca24_and_18_17(.a(a[18]), .b(b[17]), .out(s_wallace_rca24_and_18_17));
  fa fa_s_wallace_rca24_fa112_out(.a(s_wallace_rca24_fa111_or0[0]), .b(s_wallace_rca24_and_19_16[0]), .cin(s_wallace_rca24_and_18_17[0]), .fa_xor1(s_wallace_rca24_fa112_xor1), .fa_or0(s_wallace_rca24_fa112_or0));
  and_gate and_gate_s_wallace_rca24_and_19_17(.a(a[19]), .b(b[17]), .out(s_wallace_rca24_and_19_17));
  and_gate and_gate_s_wallace_rca24_and_18_18(.a(a[18]), .b(b[18]), .out(s_wallace_rca24_and_18_18));
  fa fa_s_wallace_rca24_fa113_out(.a(s_wallace_rca24_fa112_or0[0]), .b(s_wallace_rca24_and_19_17[0]), .cin(s_wallace_rca24_and_18_18[0]), .fa_xor1(s_wallace_rca24_fa113_xor1), .fa_or0(s_wallace_rca24_fa113_or0));
  and_gate and_gate_s_wallace_rca24_and_19_18(.a(a[19]), .b(b[18]), .out(s_wallace_rca24_and_19_18));
  and_gate and_gate_s_wallace_rca24_and_18_19(.a(a[18]), .b(b[19]), .out(s_wallace_rca24_and_18_19));
  fa fa_s_wallace_rca24_fa114_out(.a(s_wallace_rca24_fa113_or0[0]), .b(s_wallace_rca24_and_19_18[0]), .cin(s_wallace_rca24_and_18_19[0]), .fa_xor1(s_wallace_rca24_fa114_xor1), .fa_or0(s_wallace_rca24_fa114_or0));
  and_gate and_gate_s_wallace_rca24_and_19_19(.a(a[19]), .b(b[19]), .out(s_wallace_rca24_and_19_19));
  and_gate and_gate_s_wallace_rca24_and_18_20(.a(a[18]), .b(b[20]), .out(s_wallace_rca24_and_18_20));
  fa fa_s_wallace_rca24_fa115_out(.a(s_wallace_rca24_fa114_or0[0]), .b(s_wallace_rca24_and_19_19[0]), .cin(s_wallace_rca24_and_18_20[0]), .fa_xor1(s_wallace_rca24_fa115_xor1), .fa_or0(s_wallace_rca24_fa115_or0));
  and_gate and_gate_s_wallace_rca24_and_19_20(.a(a[19]), .b(b[20]), .out(s_wallace_rca24_and_19_20));
  and_gate and_gate_s_wallace_rca24_and_18_21(.a(a[18]), .b(b[21]), .out(s_wallace_rca24_and_18_21));
  fa fa_s_wallace_rca24_fa116_out(.a(s_wallace_rca24_fa115_or0[0]), .b(s_wallace_rca24_and_19_20[0]), .cin(s_wallace_rca24_and_18_21[0]), .fa_xor1(s_wallace_rca24_fa116_xor1), .fa_or0(s_wallace_rca24_fa116_or0));
  and_gate and_gate_s_wallace_rca24_and_19_21(.a(a[19]), .b(b[21]), .out(s_wallace_rca24_and_19_21));
  and_gate and_gate_s_wallace_rca24_and_18_22(.a(a[18]), .b(b[22]), .out(s_wallace_rca24_and_18_22));
  fa fa_s_wallace_rca24_fa117_out(.a(s_wallace_rca24_fa116_or0[0]), .b(s_wallace_rca24_and_19_21[0]), .cin(s_wallace_rca24_and_18_22[0]), .fa_xor1(s_wallace_rca24_fa117_xor1), .fa_or0(s_wallace_rca24_fa117_or0));
  and_gate and_gate_s_wallace_rca24_and_19_22(.a(a[19]), .b(b[22]), .out(s_wallace_rca24_and_19_22));
  nand_gate nand_gate_s_wallace_rca24_nand_18_23(.a(a[18]), .b(b[23]), .out(s_wallace_rca24_nand_18_23));
  fa fa_s_wallace_rca24_fa118_out(.a(s_wallace_rca24_fa117_or0[0]), .b(s_wallace_rca24_and_19_22[0]), .cin(s_wallace_rca24_nand_18_23[0]), .fa_xor1(s_wallace_rca24_fa118_xor1), .fa_or0(s_wallace_rca24_fa118_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_19_23(.a(a[19]), .b(b[23]), .out(s_wallace_rca24_nand_19_23));
  fa fa_s_wallace_rca24_fa119_out(.a(s_wallace_rca24_fa118_or0[0]), .b(s_wallace_rca24_nand_19_23[0]), .cin(s_wallace_rca24_fa39_xor1[0]), .fa_xor1(s_wallace_rca24_fa119_xor1), .fa_or0(s_wallace_rca24_fa119_or0));
  ha ha_s_wallace_rca24_ha3_out(.a(s_wallace_rca24_fa2_xor1[0]), .b(s_wallace_rca24_fa43_xor1[0]), .ha_xor0(s_wallace_rca24_ha3_xor0), .ha_and0(s_wallace_rca24_ha3_and0));
  and_gate and_gate_s_wallace_rca24_and_0_6(.a(a[0]), .b(b[6]), .out(s_wallace_rca24_and_0_6));
  fa fa_s_wallace_rca24_fa120_out(.a(s_wallace_rca24_ha3_and0[0]), .b(s_wallace_rca24_and_0_6[0]), .cin(s_wallace_rca24_fa3_xor1[0]), .fa_xor1(s_wallace_rca24_fa120_xor1), .fa_or0(s_wallace_rca24_fa120_or0));
  and_gate and_gate_s_wallace_rca24_and_1_6(.a(a[1]), .b(b[6]), .out(s_wallace_rca24_and_1_6));
  and_gate and_gate_s_wallace_rca24_and_0_7(.a(a[0]), .b(b[7]), .out(s_wallace_rca24_and_0_7));
  fa fa_s_wallace_rca24_fa121_out(.a(s_wallace_rca24_fa120_or0[0]), .b(s_wallace_rca24_and_1_6[0]), .cin(s_wallace_rca24_and_0_7[0]), .fa_xor1(s_wallace_rca24_fa121_xor1), .fa_or0(s_wallace_rca24_fa121_or0));
  and_gate and_gate_s_wallace_rca24_and_2_6(.a(a[2]), .b(b[6]), .out(s_wallace_rca24_and_2_6));
  and_gate and_gate_s_wallace_rca24_and_1_7(.a(a[1]), .b(b[7]), .out(s_wallace_rca24_and_1_7));
  fa fa_s_wallace_rca24_fa122_out(.a(s_wallace_rca24_fa121_or0[0]), .b(s_wallace_rca24_and_2_6[0]), .cin(s_wallace_rca24_and_1_7[0]), .fa_xor1(s_wallace_rca24_fa122_xor1), .fa_or0(s_wallace_rca24_fa122_or0));
  and_gate and_gate_s_wallace_rca24_and_3_6(.a(a[3]), .b(b[6]), .out(s_wallace_rca24_and_3_6));
  and_gate and_gate_s_wallace_rca24_and_2_7(.a(a[2]), .b(b[7]), .out(s_wallace_rca24_and_2_7));
  fa fa_s_wallace_rca24_fa123_out(.a(s_wallace_rca24_fa122_or0[0]), .b(s_wallace_rca24_and_3_6[0]), .cin(s_wallace_rca24_and_2_7[0]), .fa_xor1(s_wallace_rca24_fa123_xor1), .fa_or0(s_wallace_rca24_fa123_or0));
  and_gate and_gate_s_wallace_rca24_and_4_6(.a(a[4]), .b(b[6]), .out(s_wallace_rca24_and_4_6));
  and_gate and_gate_s_wallace_rca24_and_3_7(.a(a[3]), .b(b[7]), .out(s_wallace_rca24_and_3_7));
  fa fa_s_wallace_rca24_fa124_out(.a(s_wallace_rca24_fa123_or0[0]), .b(s_wallace_rca24_and_4_6[0]), .cin(s_wallace_rca24_and_3_7[0]), .fa_xor1(s_wallace_rca24_fa124_xor1), .fa_or0(s_wallace_rca24_fa124_or0));
  and_gate and_gate_s_wallace_rca24_and_5_6(.a(a[5]), .b(b[6]), .out(s_wallace_rca24_and_5_6));
  and_gate and_gate_s_wallace_rca24_and_4_7(.a(a[4]), .b(b[7]), .out(s_wallace_rca24_and_4_7));
  fa fa_s_wallace_rca24_fa125_out(.a(s_wallace_rca24_fa124_or0[0]), .b(s_wallace_rca24_and_5_6[0]), .cin(s_wallace_rca24_and_4_7[0]), .fa_xor1(s_wallace_rca24_fa125_xor1), .fa_or0(s_wallace_rca24_fa125_or0));
  and_gate and_gate_s_wallace_rca24_and_6_6(.a(a[6]), .b(b[6]), .out(s_wallace_rca24_and_6_6));
  and_gate and_gate_s_wallace_rca24_and_5_7(.a(a[5]), .b(b[7]), .out(s_wallace_rca24_and_5_7));
  fa fa_s_wallace_rca24_fa126_out(.a(s_wallace_rca24_fa125_or0[0]), .b(s_wallace_rca24_and_6_6[0]), .cin(s_wallace_rca24_and_5_7[0]), .fa_xor1(s_wallace_rca24_fa126_xor1), .fa_or0(s_wallace_rca24_fa126_or0));
  and_gate and_gate_s_wallace_rca24_and_7_6(.a(a[7]), .b(b[6]), .out(s_wallace_rca24_and_7_6));
  and_gate and_gate_s_wallace_rca24_and_6_7(.a(a[6]), .b(b[7]), .out(s_wallace_rca24_and_6_7));
  fa fa_s_wallace_rca24_fa127_out(.a(s_wallace_rca24_fa126_or0[0]), .b(s_wallace_rca24_and_7_6[0]), .cin(s_wallace_rca24_and_6_7[0]), .fa_xor1(s_wallace_rca24_fa127_xor1), .fa_or0(s_wallace_rca24_fa127_or0));
  and_gate and_gate_s_wallace_rca24_and_8_6(.a(a[8]), .b(b[6]), .out(s_wallace_rca24_and_8_6));
  and_gate and_gate_s_wallace_rca24_and_7_7(.a(a[7]), .b(b[7]), .out(s_wallace_rca24_and_7_7));
  fa fa_s_wallace_rca24_fa128_out(.a(s_wallace_rca24_fa127_or0[0]), .b(s_wallace_rca24_and_8_6[0]), .cin(s_wallace_rca24_and_7_7[0]), .fa_xor1(s_wallace_rca24_fa128_xor1), .fa_or0(s_wallace_rca24_fa128_or0));
  and_gate and_gate_s_wallace_rca24_and_9_6(.a(a[9]), .b(b[6]), .out(s_wallace_rca24_and_9_6));
  and_gate and_gate_s_wallace_rca24_and_8_7(.a(a[8]), .b(b[7]), .out(s_wallace_rca24_and_8_7));
  fa fa_s_wallace_rca24_fa129_out(.a(s_wallace_rca24_fa128_or0[0]), .b(s_wallace_rca24_and_9_6[0]), .cin(s_wallace_rca24_and_8_7[0]), .fa_xor1(s_wallace_rca24_fa129_xor1), .fa_or0(s_wallace_rca24_fa129_or0));
  and_gate and_gate_s_wallace_rca24_and_10_6(.a(a[10]), .b(b[6]), .out(s_wallace_rca24_and_10_6));
  and_gate and_gate_s_wallace_rca24_and_9_7(.a(a[9]), .b(b[7]), .out(s_wallace_rca24_and_9_7));
  fa fa_s_wallace_rca24_fa130_out(.a(s_wallace_rca24_fa129_or0[0]), .b(s_wallace_rca24_and_10_6[0]), .cin(s_wallace_rca24_and_9_7[0]), .fa_xor1(s_wallace_rca24_fa130_xor1), .fa_or0(s_wallace_rca24_fa130_or0));
  and_gate and_gate_s_wallace_rca24_and_11_6(.a(a[11]), .b(b[6]), .out(s_wallace_rca24_and_11_6));
  and_gate and_gate_s_wallace_rca24_and_10_7(.a(a[10]), .b(b[7]), .out(s_wallace_rca24_and_10_7));
  fa fa_s_wallace_rca24_fa131_out(.a(s_wallace_rca24_fa130_or0[0]), .b(s_wallace_rca24_and_11_6[0]), .cin(s_wallace_rca24_and_10_7[0]), .fa_xor1(s_wallace_rca24_fa131_xor1), .fa_or0(s_wallace_rca24_fa131_or0));
  and_gate and_gate_s_wallace_rca24_and_12_6(.a(a[12]), .b(b[6]), .out(s_wallace_rca24_and_12_6));
  and_gate and_gate_s_wallace_rca24_and_11_7(.a(a[11]), .b(b[7]), .out(s_wallace_rca24_and_11_7));
  fa fa_s_wallace_rca24_fa132_out(.a(s_wallace_rca24_fa131_or0[0]), .b(s_wallace_rca24_and_12_6[0]), .cin(s_wallace_rca24_and_11_7[0]), .fa_xor1(s_wallace_rca24_fa132_xor1), .fa_or0(s_wallace_rca24_fa132_or0));
  and_gate and_gate_s_wallace_rca24_and_13_6(.a(a[13]), .b(b[6]), .out(s_wallace_rca24_and_13_6));
  and_gate and_gate_s_wallace_rca24_and_12_7(.a(a[12]), .b(b[7]), .out(s_wallace_rca24_and_12_7));
  fa fa_s_wallace_rca24_fa133_out(.a(s_wallace_rca24_fa132_or0[0]), .b(s_wallace_rca24_and_13_6[0]), .cin(s_wallace_rca24_and_12_7[0]), .fa_xor1(s_wallace_rca24_fa133_xor1), .fa_or0(s_wallace_rca24_fa133_or0));
  and_gate and_gate_s_wallace_rca24_and_14_6(.a(a[14]), .b(b[6]), .out(s_wallace_rca24_and_14_6));
  and_gate and_gate_s_wallace_rca24_and_13_7(.a(a[13]), .b(b[7]), .out(s_wallace_rca24_and_13_7));
  fa fa_s_wallace_rca24_fa134_out(.a(s_wallace_rca24_fa133_or0[0]), .b(s_wallace_rca24_and_14_6[0]), .cin(s_wallace_rca24_and_13_7[0]), .fa_xor1(s_wallace_rca24_fa134_xor1), .fa_or0(s_wallace_rca24_fa134_or0));
  and_gate and_gate_s_wallace_rca24_and_15_6(.a(a[15]), .b(b[6]), .out(s_wallace_rca24_and_15_6));
  and_gate and_gate_s_wallace_rca24_and_14_7(.a(a[14]), .b(b[7]), .out(s_wallace_rca24_and_14_7));
  fa fa_s_wallace_rca24_fa135_out(.a(s_wallace_rca24_fa134_or0[0]), .b(s_wallace_rca24_and_15_6[0]), .cin(s_wallace_rca24_and_14_7[0]), .fa_xor1(s_wallace_rca24_fa135_xor1), .fa_or0(s_wallace_rca24_fa135_or0));
  and_gate and_gate_s_wallace_rca24_and_16_6(.a(a[16]), .b(b[6]), .out(s_wallace_rca24_and_16_6));
  and_gate and_gate_s_wallace_rca24_and_15_7(.a(a[15]), .b(b[7]), .out(s_wallace_rca24_and_15_7));
  fa fa_s_wallace_rca24_fa136_out(.a(s_wallace_rca24_fa135_or0[0]), .b(s_wallace_rca24_and_16_6[0]), .cin(s_wallace_rca24_and_15_7[0]), .fa_xor1(s_wallace_rca24_fa136_xor1), .fa_or0(s_wallace_rca24_fa136_or0));
  and_gate and_gate_s_wallace_rca24_and_17_6(.a(a[17]), .b(b[6]), .out(s_wallace_rca24_and_17_6));
  and_gate and_gate_s_wallace_rca24_and_16_7(.a(a[16]), .b(b[7]), .out(s_wallace_rca24_and_16_7));
  fa fa_s_wallace_rca24_fa137_out(.a(s_wallace_rca24_fa136_or0[0]), .b(s_wallace_rca24_and_17_6[0]), .cin(s_wallace_rca24_and_16_7[0]), .fa_xor1(s_wallace_rca24_fa137_xor1), .fa_or0(s_wallace_rca24_fa137_or0));
  and_gate and_gate_s_wallace_rca24_and_18_6(.a(a[18]), .b(b[6]), .out(s_wallace_rca24_and_18_6));
  and_gate and_gate_s_wallace_rca24_and_17_7(.a(a[17]), .b(b[7]), .out(s_wallace_rca24_and_17_7));
  fa fa_s_wallace_rca24_fa138_out(.a(s_wallace_rca24_fa137_or0[0]), .b(s_wallace_rca24_and_18_6[0]), .cin(s_wallace_rca24_and_17_7[0]), .fa_xor1(s_wallace_rca24_fa138_xor1), .fa_or0(s_wallace_rca24_fa138_or0));
  and_gate and_gate_s_wallace_rca24_and_17_8(.a(a[17]), .b(b[8]), .out(s_wallace_rca24_and_17_8));
  and_gate and_gate_s_wallace_rca24_and_16_9(.a(a[16]), .b(b[9]), .out(s_wallace_rca24_and_16_9));
  fa fa_s_wallace_rca24_fa139_out(.a(s_wallace_rca24_fa138_or0[0]), .b(s_wallace_rca24_and_17_8[0]), .cin(s_wallace_rca24_and_16_9[0]), .fa_xor1(s_wallace_rca24_fa139_xor1), .fa_or0(s_wallace_rca24_fa139_or0));
  and_gate and_gate_s_wallace_rca24_and_17_9(.a(a[17]), .b(b[9]), .out(s_wallace_rca24_and_17_9));
  and_gate and_gate_s_wallace_rca24_and_16_10(.a(a[16]), .b(b[10]), .out(s_wallace_rca24_and_16_10));
  fa fa_s_wallace_rca24_fa140_out(.a(s_wallace_rca24_fa139_or0[0]), .b(s_wallace_rca24_and_17_9[0]), .cin(s_wallace_rca24_and_16_10[0]), .fa_xor1(s_wallace_rca24_fa140_xor1), .fa_or0(s_wallace_rca24_fa140_or0));
  and_gate and_gate_s_wallace_rca24_and_17_10(.a(a[17]), .b(b[10]), .out(s_wallace_rca24_and_17_10));
  and_gate and_gate_s_wallace_rca24_and_16_11(.a(a[16]), .b(b[11]), .out(s_wallace_rca24_and_16_11));
  fa fa_s_wallace_rca24_fa141_out(.a(s_wallace_rca24_fa140_or0[0]), .b(s_wallace_rca24_and_17_10[0]), .cin(s_wallace_rca24_and_16_11[0]), .fa_xor1(s_wallace_rca24_fa141_xor1), .fa_or0(s_wallace_rca24_fa141_or0));
  and_gate and_gate_s_wallace_rca24_and_17_11(.a(a[17]), .b(b[11]), .out(s_wallace_rca24_and_17_11));
  and_gate and_gate_s_wallace_rca24_and_16_12(.a(a[16]), .b(b[12]), .out(s_wallace_rca24_and_16_12));
  fa fa_s_wallace_rca24_fa142_out(.a(s_wallace_rca24_fa141_or0[0]), .b(s_wallace_rca24_and_17_11[0]), .cin(s_wallace_rca24_and_16_12[0]), .fa_xor1(s_wallace_rca24_fa142_xor1), .fa_or0(s_wallace_rca24_fa142_or0));
  and_gate and_gate_s_wallace_rca24_and_17_12(.a(a[17]), .b(b[12]), .out(s_wallace_rca24_and_17_12));
  and_gate and_gate_s_wallace_rca24_and_16_13(.a(a[16]), .b(b[13]), .out(s_wallace_rca24_and_16_13));
  fa fa_s_wallace_rca24_fa143_out(.a(s_wallace_rca24_fa142_or0[0]), .b(s_wallace_rca24_and_17_12[0]), .cin(s_wallace_rca24_and_16_13[0]), .fa_xor1(s_wallace_rca24_fa143_xor1), .fa_or0(s_wallace_rca24_fa143_or0));
  and_gate and_gate_s_wallace_rca24_and_17_13(.a(a[17]), .b(b[13]), .out(s_wallace_rca24_and_17_13));
  and_gate and_gate_s_wallace_rca24_and_16_14(.a(a[16]), .b(b[14]), .out(s_wallace_rca24_and_16_14));
  fa fa_s_wallace_rca24_fa144_out(.a(s_wallace_rca24_fa143_or0[0]), .b(s_wallace_rca24_and_17_13[0]), .cin(s_wallace_rca24_and_16_14[0]), .fa_xor1(s_wallace_rca24_fa144_xor1), .fa_or0(s_wallace_rca24_fa144_or0));
  and_gate and_gate_s_wallace_rca24_and_17_14(.a(a[17]), .b(b[14]), .out(s_wallace_rca24_and_17_14));
  and_gate and_gate_s_wallace_rca24_and_16_15(.a(a[16]), .b(b[15]), .out(s_wallace_rca24_and_16_15));
  fa fa_s_wallace_rca24_fa145_out(.a(s_wallace_rca24_fa144_or0[0]), .b(s_wallace_rca24_and_17_14[0]), .cin(s_wallace_rca24_and_16_15[0]), .fa_xor1(s_wallace_rca24_fa145_xor1), .fa_or0(s_wallace_rca24_fa145_or0));
  and_gate and_gate_s_wallace_rca24_and_17_15(.a(a[17]), .b(b[15]), .out(s_wallace_rca24_and_17_15));
  and_gate and_gate_s_wallace_rca24_and_16_16(.a(a[16]), .b(b[16]), .out(s_wallace_rca24_and_16_16));
  fa fa_s_wallace_rca24_fa146_out(.a(s_wallace_rca24_fa145_or0[0]), .b(s_wallace_rca24_and_17_15[0]), .cin(s_wallace_rca24_and_16_16[0]), .fa_xor1(s_wallace_rca24_fa146_xor1), .fa_or0(s_wallace_rca24_fa146_or0));
  and_gate and_gate_s_wallace_rca24_and_17_16(.a(a[17]), .b(b[16]), .out(s_wallace_rca24_and_17_16));
  and_gate and_gate_s_wallace_rca24_and_16_17(.a(a[16]), .b(b[17]), .out(s_wallace_rca24_and_16_17));
  fa fa_s_wallace_rca24_fa147_out(.a(s_wallace_rca24_fa146_or0[0]), .b(s_wallace_rca24_and_17_16[0]), .cin(s_wallace_rca24_and_16_17[0]), .fa_xor1(s_wallace_rca24_fa147_xor1), .fa_or0(s_wallace_rca24_fa147_or0));
  and_gate and_gate_s_wallace_rca24_and_17_17(.a(a[17]), .b(b[17]), .out(s_wallace_rca24_and_17_17));
  and_gate and_gate_s_wallace_rca24_and_16_18(.a(a[16]), .b(b[18]), .out(s_wallace_rca24_and_16_18));
  fa fa_s_wallace_rca24_fa148_out(.a(s_wallace_rca24_fa147_or0[0]), .b(s_wallace_rca24_and_17_17[0]), .cin(s_wallace_rca24_and_16_18[0]), .fa_xor1(s_wallace_rca24_fa148_xor1), .fa_or0(s_wallace_rca24_fa148_or0));
  and_gate and_gate_s_wallace_rca24_and_17_18(.a(a[17]), .b(b[18]), .out(s_wallace_rca24_and_17_18));
  and_gate and_gate_s_wallace_rca24_and_16_19(.a(a[16]), .b(b[19]), .out(s_wallace_rca24_and_16_19));
  fa fa_s_wallace_rca24_fa149_out(.a(s_wallace_rca24_fa148_or0[0]), .b(s_wallace_rca24_and_17_18[0]), .cin(s_wallace_rca24_and_16_19[0]), .fa_xor1(s_wallace_rca24_fa149_xor1), .fa_or0(s_wallace_rca24_fa149_or0));
  and_gate and_gate_s_wallace_rca24_and_17_19(.a(a[17]), .b(b[19]), .out(s_wallace_rca24_and_17_19));
  and_gate and_gate_s_wallace_rca24_and_16_20(.a(a[16]), .b(b[20]), .out(s_wallace_rca24_and_16_20));
  fa fa_s_wallace_rca24_fa150_out(.a(s_wallace_rca24_fa149_or0[0]), .b(s_wallace_rca24_and_17_19[0]), .cin(s_wallace_rca24_and_16_20[0]), .fa_xor1(s_wallace_rca24_fa150_xor1), .fa_or0(s_wallace_rca24_fa150_or0));
  and_gate and_gate_s_wallace_rca24_and_17_20(.a(a[17]), .b(b[20]), .out(s_wallace_rca24_and_17_20));
  and_gate and_gate_s_wallace_rca24_and_16_21(.a(a[16]), .b(b[21]), .out(s_wallace_rca24_and_16_21));
  fa fa_s_wallace_rca24_fa151_out(.a(s_wallace_rca24_fa150_or0[0]), .b(s_wallace_rca24_and_17_20[0]), .cin(s_wallace_rca24_and_16_21[0]), .fa_xor1(s_wallace_rca24_fa151_xor1), .fa_or0(s_wallace_rca24_fa151_or0));
  and_gate and_gate_s_wallace_rca24_and_17_21(.a(a[17]), .b(b[21]), .out(s_wallace_rca24_and_17_21));
  and_gate and_gate_s_wallace_rca24_and_16_22(.a(a[16]), .b(b[22]), .out(s_wallace_rca24_and_16_22));
  fa fa_s_wallace_rca24_fa152_out(.a(s_wallace_rca24_fa151_or0[0]), .b(s_wallace_rca24_and_17_21[0]), .cin(s_wallace_rca24_and_16_22[0]), .fa_xor1(s_wallace_rca24_fa152_xor1), .fa_or0(s_wallace_rca24_fa152_or0));
  and_gate and_gate_s_wallace_rca24_and_17_22(.a(a[17]), .b(b[22]), .out(s_wallace_rca24_and_17_22));
  nand_gate nand_gate_s_wallace_rca24_nand_16_23(.a(a[16]), .b(b[23]), .out(s_wallace_rca24_nand_16_23));
  fa fa_s_wallace_rca24_fa153_out(.a(s_wallace_rca24_fa152_or0[0]), .b(s_wallace_rca24_and_17_22[0]), .cin(s_wallace_rca24_nand_16_23[0]), .fa_xor1(s_wallace_rca24_fa153_xor1), .fa_or0(s_wallace_rca24_fa153_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_17_23(.a(a[17]), .b(b[23]), .out(s_wallace_rca24_nand_17_23));
  fa fa_s_wallace_rca24_fa154_out(.a(s_wallace_rca24_fa153_or0[0]), .b(s_wallace_rca24_nand_17_23[0]), .cin(s_wallace_rca24_fa37_xor1[0]), .fa_xor1(s_wallace_rca24_fa154_xor1), .fa_or0(s_wallace_rca24_fa154_or0));
  fa fa_s_wallace_rca24_fa155_out(.a(s_wallace_rca24_fa154_or0[0]), .b(s_wallace_rca24_fa38_xor1[0]), .cin(s_wallace_rca24_fa79_xor1[0]), .fa_xor1(s_wallace_rca24_fa155_xor1), .fa_or0(s_wallace_rca24_fa155_or0));
  ha ha_s_wallace_rca24_ha4_out(.a(s_wallace_rca24_fa44_xor1[0]), .b(s_wallace_rca24_fa83_xor1[0]), .ha_xor0(s_wallace_rca24_ha4_xor0), .ha_and0(s_wallace_rca24_ha4_and0));
  fa fa_s_wallace_rca24_fa156_out(.a(s_wallace_rca24_ha4_and0[0]), .b(s_wallace_rca24_fa4_xor1[0]), .cin(s_wallace_rca24_fa45_xor1[0]), .fa_xor1(s_wallace_rca24_fa156_xor1), .fa_or0(s_wallace_rca24_fa156_or0));
  and_gate and_gate_s_wallace_rca24_and_0_8(.a(a[0]), .b(b[8]), .out(s_wallace_rca24_and_0_8));
  fa fa_s_wallace_rca24_fa157_out(.a(s_wallace_rca24_fa156_or0[0]), .b(s_wallace_rca24_and_0_8[0]), .cin(s_wallace_rca24_fa5_xor1[0]), .fa_xor1(s_wallace_rca24_fa157_xor1), .fa_or0(s_wallace_rca24_fa157_or0));
  and_gate and_gate_s_wallace_rca24_and_1_8(.a(a[1]), .b(b[8]), .out(s_wallace_rca24_and_1_8));
  and_gate and_gate_s_wallace_rca24_and_0_9(.a(a[0]), .b(b[9]), .out(s_wallace_rca24_and_0_9));
  fa fa_s_wallace_rca24_fa158_out(.a(s_wallace_rca24_fa157_or0[0]), .b(s_wallace_rca24_and_1_8[0]), .cin(s_wallace_rca24_and_0_9[0]), .fa_xor1(s_wallace_rca24_fa158_xor1), .fa_or0(s_wallace_rca24_fa158_or0));
  and_gate and_gate_s_wallace_rca24_and_2_8(.a(a[2]), .b(b[8]), .out(s_wallace_rca24_and_2_8));
  and_gate and_gate_s_wallace_rca24_and_1_9(.a(a[1]), .b(b[9]), .out(s_wallace_rca24_and_1_9));
  fa fa_s_wallace_rca24_fa159_out(.a(s_wallace_rca24_fa158_or0[0]), .b(s_wallace_rca24_and_2_8[0]), .cin(s_wallace_rca24_and_1_9[0]), .fa_xor1(s_wallace_rca24_fa159_xor1), .fa_or0(s_wallace_rca24_fa159_or0));
  and_gate and_gate_s_wallace_rca24_and_3_8(.a(a[3]), .b(b[8]), .out(s_wallace_rca24_and_3_8));
  and_gate and_gate_s_wallace_rca24_and_2_9(.a(a[2]), .b(b[9]), .out(s_wallace_rca24_and_2_9));
  fa fa_s_wallace_rca24_fa160_out(.a(s_wallace_rca24_fa159_or0[0]), .b(s_wallace_rca24_and_3_8[0]), .cin(s_wallace_rca24_and_2_9[0]), .fa_xor1(s_wallace_rca24_fa160_xor1), .fa_or0(s_wallace_rca24_fa160_or0));
  and_gate and_gate_s_wallace_rca24_and_4_8(.a(a[4]), .b(b[8]), .out(s_wallace_rca24_and_4_8));
  and_gate and_gate_s_wallace_rca24_and_3_9(.a(a[3]), .b(b[9]), .out(s_wallace_rca24_and_3_9));
  fa fa_s_wallace_rca24_fa161_out(.a(s_wallace_rca24_fa160_or0[0]), .b(s_wallace_rca24_and_4_8[0]), .cin(s_wallace_rca24_and_3_9[0]), .fa_xor1(s_wallace_rca24_fa161_xor1), .fa_or0(s_wallace_rca24_fa161_or0));
  and_gate and_gate_s_wallace_rca24_and_5_8(.a(a[5]), .b(b[8]), .out(s_wallace_rca24_and_5_8));
  and_gate and_gate_s_wallace_rca24_and_4_9(.a(a[4]), .b(b[9]), .out(s_wallace_rca24_and_4_9));
  fa fa_s_wallace_rca24_fa162_out(.a(s_wallace_rca24_fa161_or0[0]), .b(s_wallace_rca24_and_5_8[0]), .cin(s_wallace_rca24_and_4_9[0]), .fa_xor1(s_wallace_rca24_fa162_xor1), .fa_or0(s_wallace_rca24_fa162_or0));
  and_gate and_gate_s_wallace_rca24_and_6_8(.a(a[6]), .b(b[8]), .out(s_wallace_rca24_and_6_8));
  and_gate and_gate_s_wallace_rca24_and_5_9(.a(a[5]), .b(b[9]), .out(s_wallace_rca24_and_5_9));
  fa fa_s_wallace_rca24_fa163_out(.a(s_wallace_rca24_fa162_or0[0]), .b(s_wallace_rca24_and_6_8[0]), .cin(s_wallace_rca24_and_5_9[0]), .fa_xor1(s_wallace_rca24_fa163_xor1), .fa_or0(s_wallace_rca24_fa163_or0));
  and_gate and_gate_s_wallace_rca24_and_7_8(.a(a[7]), .b(b[8]), .out(s_wallace_rca24_and_7_8));
  and_gate and_gate_s_wallace_rca24_and_6_9(.a(a[6]), .b(b[9]), .out(s_wallace_rca24_and_6_9));
  fa fa_s_wallace_rca24_fa164_out(.a(s_wallace_rca24_fa163_or0[0]), .b(s_wallace_rca24_and_7_8[0]), .cin(s_wallace_rca24_and_6_9[0]), .fa_xor1(s_wallace_rca24_fa164_xor1), .fa_or0(s_wallace_rca24_fa164_or0));
  and_gate and_gate_s_wallace_rca24_and_8_8(.a(a[8]), .b(b[8]), .out(s_wallace_rca24_and_8_8));
  and_gate and_gate_s_wallace_rca24_and_7_9(.a(a[7]), .b(b[9]), .out(s_wallace_rca24_and_7_9));
  fa fa_s_wallace_rca24_fa165_out(.a(s_wallace_rca24_fa164_or0[0]), .b(s_wallace_rca24_and_8_8[0]), .cin(s_wallace_rca24_and_7_9[0]), .fa_xor1(s_wallace_rca24_fa165_xor1), .fa_or0(s_wallace_rca24_fa165_or0));
  and_gate and_gate_s_wallace_rca24_and_9_8(.a(a[9]), .b(b[8]), .out(s_wallace_rca24_and_9_8));
  and_gate and_gate_s_wallace_rca24_and_8_9(.a(a[8]), .b(b[9]), .out(s_wallace_rca24_and_8_9));
  fa fa_s_wallace_rca24_fa166_out(.a(s_wallace_rca24_fa165_or0[0]), .b(s_wallace_rca24_and_9_8[0]), .cin(s_wallace_rca24_and_8_9[0]), .fa_xor1(s_wallace_rca24_fa166_xor1), .fa_or0(s_wallace_rca24_fa166_or0));
  and_gate and_gate_s_wallace_rca24_and_10_8(.a(a[10]), .b(b[8]), .out(s_wallace_rca24_and_10_8));
  and_gate and_gate_s_wallace_rca24_and_9_9(.a(a[9]), .b(b[9]), .out(s_wallace_rca24_and_9_9));
  fa fa_s_wallace_rca24_fa167_out(.a(s_wallace_rca24_fa166_or0[0]), .b(s_wallace_rca24_and_10_8[0]), .cin(s_wallace_rca24_and_9_9[0]), .fa_xor1(s_wallace_rca24_fa167_xor1), .fa_or0(s_wallace_rca24_fa167_or0));
  and_gate and_gate_s_wallace_rca24_and_11_8(.a(a[11]), .b(b[8]), .out(s_wallace_rca24_and_11_8));
  and_gate and_gate_s_wallace_rca24_and_10_9(.a(a[10]), .b(b[9]), .out(s_wallace_rca24_and_10_9));
  fa fa_s_wallace_rca24_fa168_out(.a(s_wallace_rca24_fa167_or0[0]), .b(s_wallace_rca24_and_11_8[0]), .cin(s_wallace_rca24_and_10_9[0]), .fa_xor1(s_wallace_rca24_fa168_xor1), .fa_or0(s_wallace_rca24_fa168_or0));
  and_gate and_gate_s_wallace_rca24_and_12_8(.a(a[12]), .b(b[8]), .out(s_wallace_rca24_and_12_8));
  and_gate and_gate_s_wallace_rca24_and_11_9(.a(a[11]), .b(b[9]), .out(s_wallace_rca24_and_11_9));
  fa fa_s_wallace_rca24_fa169_out(.a(s_wallace_rca24_fa168_or0[0]), .b(s_wallace_rca24_and_12_8[0]), .cin(s_wallace_rca24_and_11_9[0]), .fa_xor1(s_wallace_rca24_fa169_xor1), .fa_or0(s_wallace_rca24_fa169_or0));
  and_gate and_gate_s_wallace_rca24_and_13_8(.a(a[13]), .b(b[8]), .out(s_wallace_rca24_and_13_8));
  and_gate and_gate_s_wallace_rca24_and_12_9(.a(a[12]), .b(b[9]), .out(s_wallace_rca24_and_12_9));
  fa fa_s_wallace_rca24_fa170_out(.a(s_wallace_rca24_fa169_or0[0]), .b(s_wallace_rca24_and_13_8[0]), .cin(s_wallace_rca24_and_12_9[0]), .fa_xor1(s_wallace_rca24_fa170_xor1), .fa_or0(s_wallace_rca24_fa170_or0));
  and_gate and_gate_s_wallace_rca24_and_14_8(.a(a[14]), .b(b[8]), .out(s_wallace_rca24_and_14_8));
  and_gate and_gate_s_wallace_rca24_and_13_9(.a(a[13]), .b(b[9]), .out(s_wallace_rca24_and_13_9));
  fa fa_s_wallace_rca24_fa171_out(.a(s_wallace_rca24_fa170_or0[0]), .b(s_wallace_rca24_and_14_8[0]), .cin(s_wallace_rca24_and_13_9[0]), .fa_xor1(s_wallace_rca24_fa171_xor1), .fa_or0(s_wallace_rca24_fa171_or0));
  and_gate and_gate_s_wallace_rca24_and_15_8(.a(a[15]), .b(b[8]), .out(s_wallace_rca24_and_15_8));
  and_gate and_gate_s_wallace_rca24_and_14_9(.a(a[14]), .b(b[9]), .out(s_wallace_rca24_and_14_9));
  fa fa_s_wallace_rca24_fa172_out(.a(s_wallace_rca24_fa171_or0[0]), .b(s_wallace_rca24_and_15_8[0]), .cin(s_wallace_rca24_and_14_9[0]), .fa_xor1(s_wallace_rca24_fa172_xor1), .fa_or0(s_wallace_rca24_fa172_or0));
  and_gate and_gate_s_wallace_rca24_and_16_8(.a(a[16]), .b(b[8]), .out(s_wallace_rca24_and_16_8));
  and_gate and_gate_s_wallace_rca24_and_15_9(.a(a[15]), .b(b[9]), .out(s_wallace_rca24_and_15_9));
  fa fa_s_wallace_rca24_fa173_out(.a(s_wallace_rca24_fa172_or0[0]), .b(s_wallace_rca24_and_16_8[0]), .cin(s_wallace_rca24_and_15_9[0]), .fa_xor1(s_wallace_rca24_fa173_xor1), .fa_or0(s_wallace_rca24_fa173_or0));
  and_gate and_gate_s_wallace_rca24_and_15_10(.a(a[15]), .b(b[10]), .out(s_wallace_rca24_and_15_10));
  and_gate and_gate_s_wallace_rca24_and_14_11(.a(a[14]), .b(b[11]), .out(s_wallace_rca24_and_14_11));
  fa fa_s_wallace_rca24_fa174_out(.a(s_wallace_rca24_fa173_or0[0]), .b(s_wallace_rca24_and_15_10[0]), .cin(s_wallace_rca24_and_14_11[0]), .fa_xor1(s_wallace_rca24_fa174_xor1), .fa_or0(s_wallace_rca24_fa174_or0));
  and_gate and_gate_s_wallace_rca24_and_15_11(.a(a[15]), .b(b[11]), .out(s_wallace_rca24_and_15_11));
  and_gate and_gate_s_wallace_rca24_and_14_12(.a(a[14]), .b(b[12]), .out(s_wallace_rca24_and_14_12));
  fa fa_s_wallace_rca24_fa175_out(.a(s_wallace_rca24_fa174_or0[0]), .b(s_wallace_rca24_and_15_11[0]), .cin(s_wallace_rca24_and_14_12[0]), .fa_xor1(s_wallace_rca24_fa175_xor1), .fa_or0(s_wallace_rca24_fa175_or0));
  and_gate and_gate_s_wallace_rca24_and_15_12(.a(a[15]), .b(b[12]), .out(s_wallace_rca24_and_15_12));
  and_gate and_gate_s_wallace_rca24_and_14_13(.a(a[14]), .b(b[13]), .out(s_wallace_rca24_and_14_13));
  fa fa_s_wallace_rca24_fa176_out(.a(s_wallace_rca24_fa175_or0[0]), .b(s_wallace_rca24_and_15_12[0]), .cin(s_wallace_rca24_and_14_13[0]), .fa_xor1(s_wallace_rca24_fa176_xor1), .fa_or0(s_wallace_rca24_fa176_or0));
  and_gate and_gate_s_wallace_rca24_and_15_13(.a(a[15]), .b(b[13]), .out(s_wallace_rca24_and_15_13));
  and_gate and_gate_s_wallace_rca24_and_14_14(.a(a[14]), .b(b[14]), .out(s_wallace_rca24_and_14_14));
  fa fa_s_wallace_rca24_fa177_out(.a(s_wallace_rca24_fa176_or0[0]), .b(s_wallace_rca24_and_15_13[0]), .cin(s_wallace_rca24_and_14_14[0]), .fa_xor1(s_wallace_rca24_fa177_xor1), .fa_or0(s_wallace_rca24_fa177_or0));
  and_gate and_gate_s_wallace_rca24_and_15_14(.a(a[15]), .b(b[14]), .out(s_wallace_rca24_and_15_14));
  and_gate and_gate_s_wallace_rca24_and_14_15(.a(a[14]), .b(b[15]), .out(s_wallace_rca24_and_14_15));
  fa fa_s_wallace_rca24_fa178_out(.a(s_wallace_rca24_fa177_or0[0]), .b(s_wallace_rca24_and_15_14[0]), .cin(s_wallace_rca24_and_14_15[0]), .fa_xor1(s_wallace_rca24_fa178_xor1), .fa_or0(s_wallace_rca24_fa178_or0));
  and_gate and_gate_s_wallace_rca24_and_15_15(.a(a[15]), .b(b[15]), .out(s_wallace_rca24_and_15_15));
  and_gate and_gate_s_wallace_rca24_and_14_16(.a(a[14]), .b(b[16]), .out(s_wallace_rca24_and_14_16));
  fa fa_s_wallace_rca24_fa179_out(.a(s_wallace_rca24_fa178_or0[0]), .b(s_wallace_rca24_and_15_15[0]), .cin(s_wallace_rca24_and_14_16[0]), .fa_xor1(s_wallace_rca24_fa179_xor1), .fa_or0(s_wallace_rca24_fa179_or0));
  and_gate and_gate_s_wallace_rca24_and_15_16(.a(a[15]), .b(b[16]), .out(s_wallace_rca24_and_15_16));
  and_gate and_gate_s_wallace_rca24_and_14_17(.a(a[14]), .b(b[17]), .out(s_wallace_rca24_and_14_17));
  fa fa_s_wallace_rca24_fa180_out(.a(s_wallace_rca24_fa179_or0[0]), .b(s_wallace_rca24_and_15_16[0]), .cin(s_wallace_rca24_and_14_17[0]), .fa_xor1(s_wallace_rca24_fa180_xor1), .fa_or0(s_wallace_rca24_fa180_or0));
  and_gate and_gate_s_wallace_rca24_and_15_17(.a(a[15]), .b(b[17]), .out(s_wallace_rca24_and_15_17));
  and_gate and_gate_s_wallace_rca24_and_14_18(.a(a[14]), .b(b[18]), .out(s_wallace_rca24_and_14_18));
  fa fa_s_wallace_rca24_fa181_out(.a(s_wallace_rca24_fa180_or0[0]), .b(s_wallace_rca24_and_15_17[0]), .cin(s_wallace_rca24_and_14_18[0]), .fa_xor1(s_wallace_rca24_fa181_xor1), .fa_or0(s_wallace_rca24_fa181_or0));
  and_gate and_gate_s_wallace_rca24_and_15_18(.a(a[15]), .b(b[18]), .out(s_wallace_rca24_and_15_18));
  and_gate and_gate_s_wallace_rca24_and_14_19(.a(a[14]), .b(b[19]), .out(s_wallace_rca24_and_14_19));
  fa fa_s_wallace_rca24_fa182_out(.a(s_wallace_rca24_fa181_or0[0]), .b(s_wallace_rca24_and_15_18[0]), .cin(s_wallace_rca24_and_14_19[0]), .fa_xor1(s_wallace_rca24_fa182_xor1), .fa_or0(s_wallace_rca24_fa182_or0));
  and_gate and_gate_s_wallace_rca24_and_15_19(.a(a[15]), .b(b[19]), .out(s_wallace_rca24_and_15_19));
  and_gate and_gate_s_wallace_rca24_and_14_20(.a(a[14]), .b(b[20]), .out(s_wallace_rca24_and_14_20));
  fa fa_s_wallace_rca24_fa183_out(.a(s_wallace_rca24_fa182_or0[0]), .b(s_wallace_rca24_and_15_19[0]), .cin(s_wallace_rca24_and_14_20[0]), .fa_xor1(s_wallace_rca24_fa183_xor1), .fa_or0(s_wallace_rca24_fa183_or0));
  and_gate and_gate_s_wallace_rca24_and_15_20(.a(a[15]), .b(b[20]), .out(s_wallace_rca24_and_15_20));
  and_gate and_gate_s_wallace_rca24_and_14_21(.a(a[14]), .b(b[21]), .out(s_wallace_rca24_and_14_21));
  fa fa_s_wallace_rca24_fa184_out(.a(s_wallace_rca24_fa183_or0[0]), .b(s_wallace_rca24_and_15_20[0]), .cin(s_wallace_rca24_and_14_21[0]), .fa_xor1(s_wallace_rca24_fa184_xor1), .fa_or0(s_wallace_rca24_fa184_or0));
  and_gate and_gate_s_wallace_rca24_and_15_21(.a(a[15]), .b(b[21]), .out(s_wallace_rca24_and_15_21));
  and_gate and_gate_s_wallace_rca24_and_14_22(.a(a[14]), .b(b[22]), .out(s_wallace_rca24_and_14_22));
  fa fa_s_wallace_rca24_fa185_out(.a(s_wallace_rca24_fa184_or0[0]), .b(s_wallace_rca24_and_15_21[0]), .cin(s_wallace_rca24_and_14_22[0]), .fa_xor1(s_wallace_rca24_fa185_xor1), .fa_or0(s_wallace_rca24_fa185_or0));
  and_gate and_gate_s_wallace_rca24_and_15_22(.a(a[15]), .b(b[22]), .out(s_wallace_rca24_and_15_22));
  nand_gate nand_gate_s_wallace_rca24_nand_14_23(.a(a[14]), .b(b[23]), .out(s_wallace_rca24_nand_14_23));
  fa fa_s_wallace_rca24_fa186_out(.a(s_wallace_rca24_fa185_or0[0]), .b(s_wallace_rca24_and_15_22[0]), .cin(s_wallace_rca24_nand_14_23[0]), .fa_xor1(s_wallace_rca24_fa186_xor1), .fa_or0(s_wallace_rca24_fa186_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_15_23(.a(a[15]), .b(b[23]), .out(s_wallace_rca24_nand_15_23));
  fa fa_s_wallace_rca24_fa187_out(.a(s_wallace_rca24_fa186_or0[0]), .b(s_wallace_rca24_nand_15_23[0]), .cin(s_wallace_rca24_fa35_xor1[0]), .fa_xor1(s_wallace_rca24_fa187_xor1), .fa_or0(s_wallace_rca24_fa187_or0));
  fa fa_s_wallace_rca24_fa188_out(.a(s_wallace_rca24_fa187_or0[0]), .b(s_wallace_rca24_fa36_xor1[0]), .cin(s_wallace_rca24_fa77_xor1[0]), .fa_xor1(s_wallace_rca24_fa188_xor1), .fa_or0(s_wallace_rca24_fa188_or0));
  fa fa_s_wallace_rca24_fa189_out(.a(s_wallace_rca24_fa188_or0[0]), .b(s_wallace_rca24_fa78_xor1[0]), .cin(s_wallace_rca24_fa117_xor1[0]), .fa_xor1(s_wallace_rca24_fa189_xor1), .fa_or0(s_wallace_rca24_fa189_or0));
  ha ha_s_wallace_rca24_ha5_out(.a(s_wallace_rca24_fa84_xor1[0]), .b(s_wallace_rca24_fa121_xor1[0]), .ha_xor0(s_wallace_rca24_ha5_xor0), .ha_and0(s_wallace_rca24_ha5_and0));
  fa fa_s_wallace_rca24_fa190_out(.a(s_wallace_rca24_ha5_and0[0]), .b(s_wallace_rca24_fa46_xor1[0]), .cin(s_wallace_rca24_fa85_xor1[0]), .fa_xor1(s_wallace_rca24_fa190_xor1), .fa_or0(s_wallace_rca24_fa190_or0));
  fa fa_s_wallace_rca24_fa191_out(.a(s_wallace_rca24_fa190_or0[0]), .b(s_wallace_rca24_fa6_xor1[0]), .cin(s_wallace_rca24_fa47_xor1[0]), .fa_xor1(s_wallace_rca24_fa191_xor1), .fa_or0(s_wallace_rca24_fa191_or0));
  and_gate and_gate_s_wallace_rca24_and_0_10(.a(a[0]), .b(b[10]), .out(s_wallace_rca24_and_0_10));
  fa fa_s_wallace_rca24_fa192_out(.a(s_wallace_rca24_fa191_or0[0]), .b(s_wallace_rca24_and_0_10[0]), .cin(s_wallace_rca24_fa7_xor1[0]), .fa_xor1(s_wallace_rca24_fa192_xor1), .fa_or0(s_wallace_rca24_fa192_or0));
  and_gate and_gate_s_wallace_rca24_and_1_10(.a(a[1]), .b(b[10]), .out(s_wallace_rca24_and_1_10));
  and_gate and_gate_s_wallace_rca24_and_0_11(.a(a[0]), .b(b[11]), .out(s_wallace_rca24_and_0_11));
  fa fa_s_wallace_rca24_fa193_out(.a(s_wallace_rca24_fa192_or0[0]), .b(s_wallace_rca24_and_1_10[0]), .cin(s_wallace_rca24_and_0_11[0]), .fa_xor1(s_wallace_rca24_fa193_xor1), .fa_or0(s_wallace_rca24_fa193_or0));
  and_gate and_gate_s_wallace_rca24_and_2_10(.a(a[2]), .b(b[10]), .out(s_wallace_rca24_and_2_10));
  and_gate and_gate_s_wallace_rca24_and_1_11(.a(a[1]), .b(b[11]), .out(s_wallace_rca24_and_1_11));
  fa fa_s_wallace_rca24_fa194_out(.a(s_wallace_rca24_fa193_or0[0]), .b(s_wallace_rca24_and_2_10[0]), .cin(s_wallace_rca24_and_1_11[0]), .fa_xor1(s_wallace_rca24_fa194_xor1), .fa_or0(s_wallace_rca24_fa194_or0));
  and_gate and_gate_s_wallace_rca24_and_3_10(.a(a[3]), .b(b[10]), .out(s_wallace_rca24_and_3_10));
  and_gate and_gate_s_wallace_rca24_and_2_11(.a(a[2]), .b(b[11]), .out(s_wallace_rca24_and_2_11));
  fa fa_s_wallace_rca24_fa195_out(.a(s_wallace_rca24_fa194_or0[0]), .b(s_wallace_rca24_and_3_10[0]), .cin(s_wallace_rca24_and_2_11[0]), .fa_xor1(s_wallace_rca24_fa195_xor1), .fa_or0(s_wallace_rca24_fa195_or0));
  and_gate and_gate_s_wallace_rca24_and_4_10(.a(a[4]), .b(b[10]), .out(s_wallace_rca24_and_4_10));
  and_gate and_gate_s_wallace_rca24_and_3_11(.a(a[3]), .b(b[11]), .out(s_wallace_rca24_and_3_11));
  fa fa_s_wallace_rca24_fa196_out(.a(s_wallace_rca24_fa195_or0[0]), .b(s_wallace_rca24_and_4_10[0]), .cin(s_wallace_rca24_and_3_11[0]), .fa_xor1(s_wallace_rca24_fa196_xor1), .fa_or0(s_wallace_rca24_fa196_or0));
  and_gate and_gate_s_wallace_rca24_and_5_10(.a(a[5]), .b(b[10]), .out(s_wallace_rca24_and_5_10));
  and_gate and_gate_s_wallace_rca24_and_4_11(.a(a[4]), .b(b[11]), .out(s_wallace_rca24_and_4_11));
  fa fa_s_wallace_rca24_fa197_out(.a(s_wallace_rca24_fa196_or0[0]), .b(s_wallace_rca24_and_5_10[0]), .cin(s_wallace_rca24_and_4_11[0]), .fa_xor1(s_wallace_rca24_fa197_xor1), .fa_or0(s_wallace_rca24_fa197_or0));
  and_gate and_gate_s_wallace_rca24_and_6_10(.a(a[6]), .b(b[10]), .out(s_wallace_rca24_and_6_10));
  and_gate and_gate_s_wallace_rca24_and_5_11(.a(a[5]), .b(b[11]), .out(s_wallace_rca24_and_5_11));
  fa fa_s_wallace_rca24_fa198_out(.a(s_wallace_rca24_fa197_or0[0]), .b(s_wallace_rca24_and_6_10[0]), .cin(s_wallace_rca24_and_5_11[0]), .fa_xor1(s_wallace_rca24_fa198_xor1), .fa_or0(s_wallace_rca24_fa198_or0));
  and_gate and_gate_s_wallace_rca24_and_7_10(.a(a[7]), .b(b[10]), .out(s_wallace_rca24_and_7_10));
  and_gate and_gate_s_wallace_rca24_and_6_11(.a(a[6]), .b(b[11]), .out(s_wallace_rca24_and_6_11));
  fa fa_s_wallace_rca24_fa199_out(.a(s_wallace_rca24_fa198_or0[0]), .b(s_wallace_rca24_and_7_10[0]), .cin(s_wallace_rca24_and_6_11[0]), .fa_xor1(s_wallace_rca24_fa199_xor1), .fa_or0(s_wallace_rca24_fa199_or0));
  and_gate and_gate_s_wallace_rca24_and_8_10(.a(a[8]), .b(b[10]), .out(s_wallace_rca24_and_8_10));
  and_gate and_gate_s_wallace_rca24_and_7_11(.a(a[7]), .b(b[11]), .out(s_wallace_rca24_and_7_11));
  fa fa_s_wallace_rca24_fa200_out(.a(s_wallace_rca24_fa199_or0[0]), .b(s_wallace_rca24_and_8_10[0]), .cin(s_wallace_rca24_and_7_11[0]), .fa_xor1(s_wallace_rca24_fa200_xor1), .fa_or0(s_wallace_rca24_fa200_or0));
  and_gate and_gate_s_wallace_rca24_and_9_10(.a(a[9]), .b(b[10]), .out(s_wallace_rca24_and_9_10));
  and_gate and_gate_s_wallace_rca24_and_8_11(.a(a[8]), .b(b[11]), .out(s_wallace_rca24_and_8_11));
  fa fa_s_wallace_rca24_fa201_out(.a(s_wallace_rca24_fa200_or0[0]), .b(s_wallace_rca24_and_9_10[0]), .cin(s_wallace_rca24_and_8_11[0]), .fa_xor1(s_wallace_rca24_fa201_xor1), .fa_or0(s_wallace_rca24_fa201_or0));
  and_gate and_gate_s_wallace_rca24_and_10_10(.a(a[10]), .b(b[10]), .out(s_wallace_rca24_and_10_10));
  and_gate and_gate_s_wallace_rca24_and_9_11(.a(a[9]), .b(b[11]), .out(s_wallace_rca24_and_9_11));
  fa fa_s_wallace_rca24_fa202_out(.a(s_wallace_rca24_fa201_or0[0]), .b(s_wallace_rca24_and_10_10[0]), .cin(s_wallace_rca24_and_9_11[0]), .fa_xor1(s_wallace_rca24_fa202_xor1), .fa_or0(s_wallace_rca24_fa202_or0));
  and_gate and_gate_s_wallace_rca24_and_11_10(.a(a[11]), .b(b[10]), .out(s_wallace_rca24_and_11_10));
  and_gate and_gate_s_wallace_rca24_and_10_11(.a(a[10]), .b(b[11]), .out(s_wallace_rca24_and_10_11));
  fa fa_s_wallace_rca24_fa203_out(.a(s_wallace_rca24_fa202_or0[0]), .b(s_wallace_rca24_and_11_10[0]), .cin(s_wallace_rca24_and_10_11[0]), .fa_xor1(s_wallace_rca24_fa203_xor1), .fa_or0(s_wallace_rca24_fa203_or0));
  and_gate and_gate_s_wallace_rca24_and_12_10(.a(a[12]), .b(b[10]), .out(s_wallace_rca24_and_12_10));
  and_gate and_gate_s_wallace_rca24_and_11_11(.a(a[11]), .b(b[11]), .out(s_wallace_rca24_and_11_11));
  fa fa_s_wallace_rca24_fa204_out(.a(s_wallace_rca24_fa203_or0[0]), .b(s_wallace_rca24_and_12_10[0]), .cin(s_wallace_rca24_and_11_11[0]), .fa_xor1(s_wallace_rca24_fa204_xor1), .fa_or0(s_wallace_rca24_fa204_or0));
  and_gate and_gate_s_wallace_rca24_and_13_10(.a(a[13]), .b(b[10]), .out(s_wallace_rca24_and_13_10));
  and_gate and_gate_s_wallace_rca24_and_12_11(.a(a[12]), .b(b[11]), .out(s_wallace_rca24_and_12_11));
  fa fa_s_wallace_rca24_fa205_out(.a(s_wallace_rca24_fa204_or0[0]), .b(s_wallace_rca24_and_13_10[0]), .cin(s_wallace_rca24_and_12_11[0]), .fa_xor1(s_wallace_rca24_fa205_xor1), .fa_or0(s_wallace_rca24_fa205_or0));
  and_gate and_gate_s_wallace_rca24_and_14_10(.a(a[14]), .b(b[10]), .out(s_wallace_rca24_and_14_10));
  and_gate and_gate_s_wallace_rca24_and_13_11(.a(a[13]), .b(b[11]), .out(s_wallace_rca24_and_13_11));
  fa fa_s_wallace_rca24_fa206_out(.a(s_wallace_rca24_fa205_or0[0]), .b(s_wallace_rca24_and_14_10[0]), .cin(s_wallace_rca24_and_13_11[0]), .fa_xor1(s_wallace_rca24_fa206_xor1), .fa_or0(s_wallace_rca24_fa206_or0));
  and_gate and_gate_s_wallace_rca24_and_13_12(.a(a[13]), .b(b[12]), .out(s_wallace_rca24_and_13_12));
  and_gate and_gate_s_wallace_rca24_and_12_13(.a(a[12]), .b(b[13]), .out(s_wallace_rca24_and_12_13));
  fa fa_s_wallace_rca24_fa207_out(.a(s_wallace_rca24_fa206_or0[0]), .b(s_wallace_rca24_and_13_12[0]), .cin(s_wallace_rca24_and_12_13[0]), .fa_xor1(s_wallace_rca24_fa207_xor1), .fa_or0(s_wallace_rca24_fa207_or0));
  and_gate and_gate_s_wallace_rca24_and_13_13(.a(a[13]), .b(b[13]), .out(s_wallace_rca24_and_13_13));
  and_gate and_gate_s_wallace_rca24_and_12_14(.a(a[12]), .b(b[14]), .out(s_wallace_rca24_and_12_14));
  fa fa_s_wallace_rca24_fa208_out(.a(s_wallace_rca24_fa207_or0[0]), .b(s_wallace_rca24_and_13_13[0]), .cin(s_wallace_rca24_and_12_14[0]), .fa_xor1(s_wallace_rca24_fa208_xor1), .fa_or0(s_wallace_rca24_fa208_or0));
  and_gate and_gate_s_wallace_rca24_and_13_14(.a(a[13]), .b(b[14]), .out(s_wallace_rca24_and_13_14));
  and_gate and_gate_s_wallace_rca24_and_12_15(.a(a[12]), .b(b[15]), .out(s_wallace_rca24_and_12_15));
  fa fa_s_wallace_rca24_fa209_out(.a(s_wallace_rca24_fa208_or0[0]), .b(s_wallace_rca24_and_13_14[0]), .cin(s_wallace_rca24_and_12_15[0]), .fa_xor1(s_wallace_rca24_fa209_xor1), .fa_or0(s_wallace_rca24_fa209_or0));
  and_gate and_gate_s_wallace_rca24_and_13_15(.a(a[13]), .b(b[15]), .out(s_wallace_rca24_and_13_15));
  and_gate and_gate_s_wallace_rca24_and_12_16(.a(a[12]), .b(b[16]), .out(s_wallace_rca24_and_12_16));
  fa fa_s_wallace_rca24_fa210_out(.a(s_wallace_rca24_fa209_or0[0]), .b(s_wallace_rca24_and_13_15[0]), .cin(s_wallace_rca24_and_12_16[0]), .fa_xor1(s_wallace_rca24_fa210_xor1), .fa_or0(s_wallace_rca24_fa210_or0));
  and_gate and_gate_s_wallace_rca24_and_13_16(.a(a[13]), .b(b[16]), .out(s_wallace_rca24_and_13_16));
  and_gate and_gate_s_wallace_rca24_and_12_17(.a(a[12]), .b(b[17]), .out(s_wallace_rca24_and_12_17));
  fa fa_s_wallace_rca24_fa211_out(.a(s_wallace_rca24_fa210_or0[0]), .b(s_wallace_rca24_and_13_16[0]), .cin(s_wallace_rca24_and_12_17[0]), .fa_xor1(s_wallace_rca24_fa211_xor1), .fa_or0(s_wallace_rca24_fa211_or0));
  and_gate and_gate_s_wallace_rca24_and_13_17(.a(a[13]), .b(b[17]), .out(s_wallace_rca24_and_13_17));
  and_gate and_gate_s_wallace_rca24_and_12_18(.a(a[12]), .b(b[18]), .out(s_wallace_rca24_and_12_18));
  fa fa_s_wallace_rca24_fa212_out(.a(s_wallace_rca24_fa211_or0[0]), .b(s_wallace_rca24_and_13_17[0]), .cin(s_wallace_rca24_and_12_18[0]), .fa_xor1(s_wallace_rca24_fa212_xor1), .fa_or0(s_wallace_rca24_fa212_or0));
  and_gate and_gate_s_wallace_rca24_and_13_18(.a(a[13]), .b(b[18]), .out(s_wallace_rca24_and_13_18));
  and_gate and_gate_s_wallace_rca24_and_12_19(.a(a[12]), .b(b[19]), .out(s_wallace_rca24_and_12_19));
  fa fa_s_wallace_rca24_fa213_out(.a(s_wallace_rca24_fa212_or0[0]), .b(s_wallace_rca24_and_13_18[0]), .cin(s_wallace_rca24_and_12_19[0]), .fa_xor1(s_wallace_rca24_fa213_xor1), .fa_or0(s_wallace_rca24_fa213_or0));
  and_gate and_gate_s_wallace_rca24_and_13_19(.a(a[13]), .b(b[19]), .out(s_wallace_rca24_and_13_19));
  and_gate and_gate_s_wallace_rca24_and_12_20(.a(a[12]), .b(b[20]), .out(s_wallace_rca24_and_12_20));
  fa fa_s_wallace_rca24_fa214_out(.a(s_wallace_rca24_fa213_or0[0]), .b(s_wallace_rca24_and_13_19[0]), .cin(s_wallace_rca24_and_12_20[0]), .fa_xor1(s_wallace_rca24_fa214_xor1), .fa_or0(s_wallace_rca24_fa214_or0));
  and_gate and_gate_s_wallace_rca24_and_13_20(.a(a[13]), .b(b[20]), .out(s_wallace_rca24_and_13_20));
  and_gate and_gate_s_wallace_rca24_and_12_21(.a(a[12]), .b(b[21]), .out(s_wallace_rca24_and_12_21));
  fa fa_s_wallace_rca24_fa215_out(.a(s_wallace_rca24_fa214_or0[0]), .b(s_wallace_rca24_and_13_20[0]), .cin(s_wallace_rca24_and_12_21[0]), .fa_xor1(s_wallace_rca24_fa215_xor1), .fa_or0(s_wallace_rca24_fa215_or0));
  and_gate and_gate_s_wallace_rca24_and_13_21(.a(a[13]), .b(b[21]), .out(s_wallace_rca24_and_13_21));
  and_gate and_gate_s_wallace_rca24_and_12_22(.a(a[12]), .b(b[22]), .out(s_wallace_rca24_and_12_22));
  fa fa_s_wallace_rca24_fa216_out(.a(s_wallace_rca24_fa215_or0[0]), .b(s_wallace_rca24_and_13_21[0]), .cin(s_wallace_rca24_and_12_22[0]), .fa_xor1(s_wallace_rca24_fa216_xor1), .fa_or0(s_wallace_rca24_fa216_or0));
  and_gate and_gate_s_wallace_rca24_and_13_22(.a(a[13]), .b(b[22]), .out(s_wallace_rca24_and_13_22));
  nand_gate nand_gate_s_wallace_rca24_nand_12_23(.a(a[12]), .b(b[23]), .out(s_wallace_rca24_nand_12_23));
  fa fa_s_wallace_rca24_fa217_out(.a(s_wallace_rca24_fa216_or0[0]), .b(s_wallace_rca24_and_13_22[0]), .cin(s_wallace_rca24_nand_12_23[0]), .fa_xor1(s_wallace_rca24_fa217_xor1), .fa_or0(s_wallace_rca24_fa217_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_13_23(.a(a[13]), .b(b[23]), .out(s_wallace_rca24_nand_13_23));
  fa fa_s_wallace_rca24_fa218_out(.a(s_wallace_rca24_fa217_or0[0]), .b(s_wallace_rca24_nand_13_23[0]), .cin(s_wallace_rca24_fa33_xor1[0]), .fa_xor1(s_wallace_rca24_fa218_xor1), .fa_or0(s_wallace_rca24_fa218_or0));
  fa fa_s_wallace_rca24_fa219_out(.a(s_wallace_rca24_fa218_or0[0]), .b(s_wallace_rca24_fa34_xor1[0]), .cin(s_wallace_rca24_fa75_xor1[0]), .fa_xor1(s_wallace_rca24_fa219_xor1), .fa_or0(s_wallace_rca24_fa219_or0));
  fa fa_s_wallace_rca24_fa220_out(.a(s_wallace_rca24_fa219_or0[0]), .b(s_wallace_rca24_fa76_xor1[0]), .cin(s_wallace_rca24_fa115_xor1[0]), .fa_xor1(s_wallace_rca24_fa220_xor1), .fa_or0(s_wallace_rca24_fa220_or0));
  fa fa_s_wallace_rca24_fa221_out(.a(s_wallace_rca24_fa220_or0[0]), .b(s_wallace_rca24_fa116_xor1[0]), .cin(s_wallace_rca24_fa153_xor1[0]), .fa_xor1(s_wallace_rca24_fa221_xor1), .fa_or0(s_wallace_rca24_fa221_or0));
  ha ha_s_wallace_rca24_ha6_out(.a(s_wallace_rca24_fa122_xor1[0]), .b(s_wallace_rca24_fa157_xor1[0]), .ha_xor0(s_wallace_rca24_ha6_xor0), .ha_and0(s_wallace_rca24_ha6_and0));
  fa fa_s_wallace_rca24_fa222_out(.a(s_wallace_rca24_ha6_and0[0]), .b(s_wallace_rca24_fa86_xor1[0]), .cin(s_wallace_rca24_fa123_xor1[0]), .fa_xor1(s_wallace_rca24_fa222_xor1), .fa_or0(s_wallace_rca24_fa222_or0));
  fa fa_s_wallace_rca24_fa223_out(.a(s_wallace_rca24_fa222_or0[0]), .b(s_wallace_rca24_fa48_xor1[0]), .cin(s_wallace_rca24_fa87_xor1[0]), .fa_xor1(s_wallace_rca24_fa223_xor1), .fa_or0(s_wallace_rca24_fa223_or0));
  fa fa_s_wallace_rca24_fa224_out(.a(s_wallace_rca24_fa223_or0[0]), .b(s_wallace_rca24_fa8_xor1[0]), .cin(s_wallace_rca24_fa49_xor1[0]), .fa_xor1(s_wallace_rca24_fa224_xor1), .fa_or0(s_wallace_rca24_fa224_or0));
  and_gate and_gate_s_wallace_rca24_and_0_12(.a(a[0]), .b(b[12]), .out(s_wallace_rca24_and_0_12));
  fa fa_s_wallace_rca24_fa225_out(.a(s_wallace_rca24_fa224_or0[0]), .b(s_wallace_rca24_and_0_12[0]), .cin(s_wallace_rca24_fa9_xor1[0]), .fa_xor1(s_wallace_rca24_fa225_xor1), .fa_or0(s_wallace_rca24_fa225_or0));
  and_gate and_gate_s_wallace_rca24_and_1_12(.a(a[1]), .b(b[12]), .out(s_wallace_rca24_and_1_12));
  and_gate and_gate_s_wallace_rca24_and_0_13(.a(a[0]), .b(b[13]), .out(s_wallace_rca24_and_0_13));
  fa fa_s_wallace_rca24_fa226_out(.a(s_wallace_rca24_fa225_or0[0]), .b(s_wallace_rca24_and_1_12[0]), .cin(s_wallace_rca24_and_0_13[0]), .fa_xor1(s_wallace_rca24_fa226_xor1), .fa_or0(s_wallace_rca24_fa226_or0));
  and_gate and_gate_s_wallace_rca24_and_2_12(.a(a[2]), .b(b[12]), .out(s_wallace_rca24_and_2_12));
  and_gate and_gate_s_wallace_rca24_and_1_13(.a(a[1]), .b(b[13]), .out(s_wallace_rca24_and_1_13));
  fa fa_s_wallace_rca24_fa227_out(.a(s_wallace_rca24_fa226_or0[0]), .b(s_wallace_rca24_and_2_12[0]), .cin(s_wallace_rca24_and_1_13[0]), .fa_xor1(s_wallace_rca24_fa227_xor1), .fa_or0(s_wallace_rca24_fa227_or0));
  and_gate and_gate_s_wallace_rca24_and_3_12(.a(a[3]), .b(b[12]), .out(s_wallace_rca24_and_3_12));
  and_gate and_gate_s_wallace_rca24_and_2_13(.a(a[2]), .b(b[13]), .out(s_wallace_rca24_and_2_13));
  fa fa_s_wallace_rca24_fa228_out(.a(s_wallace_rca24_fa227_or0[0]), .b(s_wallace_rca24_and_3_12[0]), .cin(s_wallace_rca24_and_2_13[0]), .fa_xor1(s_wallace_rca24_fa228_xor1), .fa_or0(s_wallace_rca24_fa228_or0));
  and_gate and_gate_s_wallace_rca24_and_4_12(.a(a[4]), .b(b[12]), .out(s_wallace_rca24_and_4_12));
  and_gate and_gate_s_wallace_rca24_and_3_13(.a(a[3]), .b(b[13]), .out(s_wallace_rca24_and_3_13));
  fa fa_s_wallace_rca24_fa229_out(.a(s_wallace_rca24_fa228_or0[0]), .b(s_wallace_rca24_and_4_12[0]), .cin(s_wallace_rca24_and_3_13[0]), .fa_xor1(s_wallace_rca24_fa229_xor1), .fa_or0(s_wallace_rca24_fa229_or0));
  and_gate and_gate_s_wallace_rca24_and_5_12(.a(a[5]), .b(b[12]), .out(s_wallace_rca24_and_5_12));
  and_gate and_gate_s_wallace_rca24_and_4_13(.a(a[4]), .b(b[13]), .out(s_wallace_rca24_and_4_13));
  fa fa_s_wallace_rca24_fa230_out(.a(s_wallace_rca24_fa229_or0[0]), .b(s_wallace_rca24_and_5_12[0]), .cin(s_wallace_rca24_and_4_13[0]), .fa_xor1(s_wallace_rca24_fa230_xor1), .fa_or0(s_wallace_rca24_fa230_or0));
  and_gate and_gate_s_wallace_rca24_and_6_12(.a(a[6]), .b(b[12]), .out(s_wallace_rca24_and_6_12));
  and_gate and_gate_s_wallace_rca24_and_5_13(.a(a[5]), .b(b[13]), .out(s_wallace_rca24_and_5_13));
  fa fa_s_wallace_rca24_fa231_out(.a(s_wallace_rca24_fa230_or0[0]), .b(s_wallace_rca24_and_6_12[0]), .cin(s_wallace_rca24_and_5_13[0]), .fa_xor1(s_wallace_rca24_fa231_xor1), .fa_or0(s_wallace_rca24_fa231_or0));
  and_gate and_gate_s_wallace_rca24_and_7_12(.a(a[7]), .b(b[12]), .out(s_wallace_rca24_and_7_12));
  and_gate and_gate_s_wallace_rca24_and_6_13(.a(a[6]), .b(b[13]), .out(s_wallace_rca24_and_6_13));
  fa fa_s_wallace_rca24_fa232_out(.a(s_wallace_rca24_fa231_or0[0]), .b(s_wallace_rca24_and_7_12[0]), .cin(s_wallace_rca24_and_6_13[0]), .fa_xor1(s_wallace_rca24_fa232_xor1), .fa_or0(s_wallace_rca24_fa232_or0));
  and_gate and_gate_s_wallace_rca24_and_8_12(.a(a[8]), .b(b[12]), .out(s_wallace_rca24_and_8_12));
  and_gate and_gate_s_wallace_rca24_and_7_13(.a(a[7]), .b(b[13]), .out(s_wallace_rca24_and_7_13));
  fa fa_s_wallace_rca24_fa233_out(.a(s_wallace_rca24_fa232_or0[0]), .b(s_wallace_rca24_and_8_12[0]), .cin(s_wallace_rca24_and_7_13[0]), .fa_xor1(s_wallace_rca24_fa233_xor1), .fa_or0(s_wallace_rca24_fa233_or0));
  and_gate and_gate_s_wallace_rca24_and_9_12(.a(a[9]), .b(b[12]), .out(s_wallace_rca24_and_9_12));
  and_gate and_gate_s_wallace_rca24_and_8_13(.a(a[8]), .b(b[13]), .out(s_wallace_rca24_and_8_13));
  fa fa_s_wallace_rca24_fa234_out(.a(s_wallace_rca24_fa233_or0[0]), .b(s_wallace_rca24_and_9_12[0]), .cin(s_wallace_rca24_and_8_13[0]), .fa_xor1(s_wallace_rca24_fa234_xor1), .fa_or0(s_wallace_rca24_fa234_or0));
  and_gate and_gate_s_wallace_rca24_and_10_12(.a(a[10]), .b(b[12]), .out(s_wallace_rca24_and_10_12));
  and_gate and_gate_s_wallace_rca24_and_9_13(.a(a[9]), .b(b[13]), .out(s_wallace_rca24_and_9_13));
  fa fa_s_wallace_rca24_fa235_out(.a(s_wallace_rca24_fa234_or0[0]), .b(s_wallace_rca24_and_10_12[0]), .cin(s_wallace_rca24_and_9_13[0]), .fa_xor1(s_wallace_rca24_fa235_xor1), .fa_or0(s_wallace_rca24_fa235_or0));
  and_gate and_gate_s_wallace_rca24_and_11_12(.a(a[11]), .b(b[12]), .out(s_wallace_rca24_and_11_12));
  and_gate and_gate_s_wallace_rca24_and_10_13(.a(a[10]), .b(b[13]), .out(s_wallace_rca24_and_10_13));
  fa fa_s_wallace_rca24_fa236_out(.a(s_wallace_rca24_fa235_or0[0]), .b(s_wallace_rca24_and_11_12[0]), .cin(s_wallace_rca24_and_10_13[0]), .fa_xor1(s_wallace_rca24_fa236_xor1), .fa_or0(s_wallace_rca24_fa236_or0));
  and_gate and_gate_s_wallace_rca24_and_12_12(.a(a[12]), .b(b[12]), .out(s_wallace_rca24_and_12_12));
  and_gate and_gate_s_wallace_rca24_and_11_13(.a(a[11]), .b(b[13]), .out(s_wallace_rca24_and_11_13));
  fa fa_s_wallace_rca24_fa237_out(.a(s_wallace_rca24_fa236_or0[0]), .b(s_wallace_rca24_and_12_12[0]), .cin(s_wallace_rca24_and_11_13[0]), .fa_xor1(s_wallace_rca24_fa237_xor1), .fa_or0(s_wallace_rca24_fa237_or0));
  and_gate and_gate_s_wallace_rca24_and_11_14(.a(a[11]), .b(b[14]), .out(s_wallace_rca24_and_11_14));
  and_gate and_gate_s_wallace_rca24_and_10_15(.a(a[10]), .b(b[15]), .out(s_wallace_rca24_and_10_15));
  fa fa_s_wallace_rca24_fa238_out(.a(s_wallace_rca24_fa237_or0[0]), .b(s_wallace_rca24_and_11_14[0]), .cin(s_wallace_rca24_and_10_15[0]), .fa_xor1(s_wallace_rca24_fa238_xor1), .fa_or0(s_wallace_rca24_fa238_or0));
  and_gate and_gate_s_wallace_rca24_and_11_15(.a(a[11]), .b(b[15]), .out(s_wallace_rca24_and_11_15));
  and_gate and_gate_s_wallace_rca24_and_10_16(.a(a[10]), .b(b[16]), .out(s_wallace_rca24_and_10_16));
  fa fa_s_wallace_rca24_fa239_out(.a(s_wallace_rca24_fa238_or0[0]), .b(s_wallace_rca24_and_11_15[0]), .cin(s_wallace_rca24_and_10_16[0]), .fa_xor1(s_wallace_rca24_fa239_xor1), .fa_or0(s_wallace_rca24_fa239_or0));
  and_gate and_gate_s_wallace_rca24_and_11_16(.a(a[11]), .b(b[16]), .out(s_wallace_rca24_and_11_16));
  and_gate and_gate_s_wallace_rca24_and_10_17(.a(a[10]), .b(b[17]), .out(s_wallace_rca24_and_10_17));
  fa fa_s_wallace_rca24_fa240_out(.a(s_wallace_rca24_fa239_or0[0]), .b(s_wallace_rca24_and_11_16[0]), .cin(s_wallace_rca24_and_10_17[0]), .fa_xor1(s_wallace_rca24_fa240_xor1), .fa_or0(s_wallace_rca24_fa240_or0));
  and_gate and_gate_s_wallace_rca24_and_11_17(.a(a[11]), .b(b[17]), .out(s_wallace_rca24_and_11_17));
  and_gate and_gate_s_wallace_rca24_and_10_18(.a(a[10]), .b(b[18]), .out(s_wallace_rca24_and_10_18));
  fa fa_s_wallace_rca24_fa241_out(.a(s_wallace_rca24_fa240_or0[0]), .b(s_wallace_rca24_and_11_17[0]), .cin(s_wallace_rca24_and_10_18[0]), .fa_xor1(s_wallace_rca24_fa241_xor1), .fa_or0(s_wallace_rca24_fa241_or0));
  and_gate and_gate_s_wallace_rca24_and_11_18(.a(a[11]), .b(b[18]), .out(s_wallace_rca24_and_11_18));
  and_gate and_gate_s_wallace_rca24_and_10_19(.a(a[10]), .b(b[19]), .out(s_wallace_rca24_and_10_19));
  fa fa_s_wallace_rca24_fa242_out(.a(s_wallace_rca24_fa241_or0[0]), .b(s_wallace_rca24_and_11_18[0]), .cin(s_wallace_rca24_and_10_19[0]), .fa_xor1(s_wallace_rca24_fa242_xor1), .fa_or0(s_wallace_rca24_fa242_or0));
  and_gate and_gate_s_wallace_rca24_and_11_19(.a(a[11]), .b(b[19]), .out(s_wallace_rca24_and_11_19));
  and_gate and_gate_s_wallace_rca24_and_10_20(.a(a[10]), .b(b[20]), .out(s_wallace_rca24_and_10_20));
  fa fa_s_wallace_rca24_fa243_out(.a(s_wallace_rca24_fa242_or0[0]), .b(s_wallace_rca24_and_11_19[0]), .cin(s_wallace_rca24_and_10_20[0]), .fa_xor1(s_wallace_rca24_fa243_xor1), .fa_or0(s_wallace_rca24_fa243_or0));
  and_gate and_gate_s_wallace_rca24_and_11_20(.a(a[11]), .b(b[20]), .out(s_wallace_rca24_and_11_20));
  and_gate and_gate_s_wallace_rca24_and_10_21(.a(a[10]), .b(b[21]), .out(s_wallace_rca24_and_10_21));
  fa fa_s_wallace_rca24_fa244_out(.a(s_wallace_rca24_fa243_or0[0]), .b(s_wallace_rca24_and_11_20[0]), .cin(s_wallace_rca24_and_10_21[0]), .fa_xor1(s_wallace_rca24_fa244_xor1), .fa_or0(s_wallace_rca24_fa244_or0));
  and_gate and_gate_s_wallace_rca24_and_11_21(.a(a[11]), .b(b[21]), .out(s_wallace_rca24_and_11_21));
  and_gate and_gate_s_wallace_rca24_and_10_22(.a(a[10]), .b(b[22]), .out(s_wallace_rca24_and_10_22));
  fa fa_s_wallace_rca24_fa245_out(.a(s_wallace_rca24_fa244_or0[0]), .b(s_wallace_rca24_and_11_21[0]), .cin(s_wallace_rca24_and_10_22[0]), .fa_xor1(s_wallace_rca24_fa245_xor1), .fa_or0(s_wallace_rca24_fa245_or0));
  and_gate and_gate_s_wallace_rca24_and_11_22(.a(a[11]), .b(b[22]), .out(s_wallace_rca24_and_11_22));
  nand_gate nand_gate_s_wallace_rca24_nand_10_23(.a(a[10]), .b(b[23]), .out(s_wallace_rca24_nand_10_23));
  fa fa_s_wallace_rca24_fa246_out(.a(s_wallace_rca24_fa245_or0[0]), .b(s_wallace_rca24_and_11_22[0]), .cin(s_wallace_rca24_nand_10_23[0]), .fa_xor1(s_wallace_rca24_fa246_xor1), .fa_or0(s_wallace_rca24_fa246_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_11_23(.a(a[11]), .b(b[23]), .out(s_wallace_rca24_nand_11_23));
  fa fa_s_wallace_rca24_fa247_out(.a(s_wallace_rca24_fa246_or0[0]), .b(s_wallace_rca24_nand_11_23[0]), .cin(s_wallace_rca24_fa31_xor1[0]), .fa_xor1(s_wallace_rca24_fa247_xor1), .fa_or0(s_wallace_rca24_fa247_or0));
  fa fa_s_wallace_rca24_fa248_out(.a(s_wallace_rca24_fa247_or0[0]), .b(s_wallace_rca24_fa32_xor1[0]), .cin(s_wallace_rca24_fa73_xor1[0]), .fa_xor1(s_wallace_rca24_fa248_xor1), .fa_or0(s_wallace_rca24_fa248_or0));
  fa fa_s_wallace_rca24_fa249_out(.a(s_wallace_rca24_fa248_or0[0]), .b(s_wallace_rca24_fa74_xor1[0]), .cin(s_wallace_rca24_fa113_xor1[0]), .fa_xor1(s_wallace_rca24_fa249_xor1), .fa_or0(s_wallace_rca24_fa249_or0));
  fa fa_s_wallace_rca24_fa250_out(.a(s_wallace_rca24_fa249_or0[0]), .b(s_wallace_rca24_fa114_xor1[0]), .cin(s_wallace_rca24_fa151_xor1[0]), .fa_xor1(s_wallace_rca24_fa250_xor1), .fa_or0(s_wallace_rca24_fa250_or0));
  fa fa_s_wallace_rca24_fa251_out(.a(s_wallace_rca24_fa250_or0[0]), .b(s_wallace_rca24_fa152_xor1[0]), .cin(s_wallace_rca24_fa187_xor1[0]), .fa_xor1(s_wallace_rca24_fa251_xor1), .fa_or0(s_wallace_rca24_fa251_or0));
  ha ha_s_wallace_rca24_ha7_out(.a(s_wallace_rca24_fa158_xor1[0]), .b(s_wallace_rca24_fa191_xor1[0]), .ha_xor0(s_wallace_rca24_ha7_xor0), .ha_and0(s_wallace_rca24_ha7_and0));
  fa fa_s_wallace_rca24_fa252_out(.a(s_wallace_rca24_ha7_and0[0]), .b(s_wallace_rca24_fa124_xor1[0]), .cin(s_wallace_rca24_fa159_xor1[0]), .fa_xor1(s_wallace_rca24_fa252_xor1), .fa_or0(s_wallace_rca24_fa252_or0));
  fa fa_s_wallace_rca24_fa253_out(.a(s_wallace_rca24_fa252_or0[0]), .b(s_wallace_rca24_fa88_xor1[0]), .cin(s_wallace_rca24_fa125_xor1[0]), .fa_xor1(s_wallace_rca24_fa253_xor1), .fa_or0(s_wallace_rca24_fa253_or0));
  fa fa_s_wallace_rca24_fa254_out(.a(s_wallace_rca24_fa253_or0[0]), .b(s_wallace_rca24_fa50_xor1[0]), .cin(s_wallace_rca24_fa89_xor1[0]), .fa_xor1(s_wallace_rca24_fa254_xor1), .fa_or0(s_wallace_rca24_fa254_or0));
  fa fa_s_wallace_rca24_fa255_out(.a(s_wallace_rca24_fa254_or0[0]), .b(s_wallace_rca24_fa10_xor1[0]), .cin(s_wallace_rca24_fa51_xor1[0]), .fa_xor1(s_wallace_rca24_fa255_xor1), .fa_or0(s_wallace_rca24_fa255_or0));
  and_gate and_gate_s_wallace_rca24_and_0_14(.a(a[0]), .b(b[14]), .out(s_wallace_rca24_and_0_14));
  fa fa_s_wallace_rca24_fa256_out(.a(s_wallace_rca24_fa255_or0[0]), .b(s_wallace_rca24_and_0_14[0]), .cin(s_wallace_rca24_fa11_xor1[0]), .fa_xor1(s_wallace_rca24_fa256_xor1), .fa_or0(s_wallace_rca24_fa256_or0));
  and_gate and_gate_s_wallace_rca24_and_1_14(.a(a[1]), .b(b[14]), .out(s_wallace_rca24_and_1_14));
  and_gate and_gate_s_wallace_rca24_and_0_15(.a(a[0]), .b(b[15]), .out(s_wallace_rca24_and_0_15));
  fa fa_s_wallace_rca24_fa257_out(.a(s_wallace_rca24_fa256_or0[0]), .b(s_wallace_rca24_and_1_14[0]), .cin(s_wallace_rca24_and_0_15[0]), .fa_xor1(s_wallace_rca24_fa257_xor1), .fa_or0(s_wallace_rca24_fa257_or0));
  and_gate and_gate_s_wallace_rca24_and_2_14(.a(a[2]), .b(b[14]), .out(s_wallace_rca24_and_2_14));
  and_gate and_gate_s_wallace_rca24_and_1_15(.a(a[1]), .b(b[15]), .out(s_wallace_rca24_and_1_15));
  fa fa_s_wallace_rca24_fa258_out(.a(s_wallace_rca24_fa257_or0[0]), .b(s_wallace_rca24_and_2_14[0]), .cin(s_wallace_rca24_and_1_15[0]), .fa_xor1(s_wallace_rca24_fa258_xor1), .fa_or0(s_wallace_rca24_fa258_or0));
  and_gate and_gate_s_wallace_rca24_and_3_14(.a(a[3]), .b(b[14]), .out(s_wallace_rca24_and_3_14));
  and_gate and_gate_s_wallace_rca24_and_2_15(.a(a[2]), .b(b[15]), .out(s_wallace_rca24_and_2_15));
  fa fa_s_wallace_rca24_fa259_out(.a(s_wallace_rca24_fa258_or0[0]), .b(s_wallace_rca24_and_3_14[0]), .cin(s_wallace_rca24_and_2_15[0]), .fa_xor1(s_wallace_rca24_fa259_xor1), .fa_or0(s_wallace_rca24_fa259_or0));
  and_gate and_gate_s_wallace_rca24_and_4_14(.a(a[4]), .b(b[14]), .out(s_wallace_rca24_and_4_14));
  and_gate and_gate_s_wallace_rca24_and_3_15(.a(a[3]), .b(b[15]), .out(s_wallace_rca24_and_3_15));
  fa fa_s_wallace_rca24_fa260_out(.a(s_wallace_rca24_fa259_or0[0]), .b(s_wallace_rca24_and_4_14[0]), .cin(s_wallace_rca24_and_3_15[0]), .fa_xor1(s_wallace_rca24_fa260_xor1), .fa_or0(s_wallace_rca24_fa260_or0));
  and_gate and_gate_s_wallace_rca24_and_5_14(.a(a[5]), .b(b[14]), .out(s_wallace_rca24_and_5_14));
  and_gate and_gate_s_wallace_rca24_and_4_15(.a(a[4]), .b(b[15]), .out(s_wallace_rca24_and_4_15));
  fa fa_s_wallace_rca24_fa261_out(.a(s_wallace_rca24_fa260_or0[0]), .b(s_wallace_rca24_and_5_14[0]), .cin(s_wallace_rca24_and_4_15[0]), .fa_xor1(s_wallace_rca24_fa261_xor1), .fa_or0(s_wallace_rca24_fa261_or0));
  and_gate and_gate_s_wallace_rca24_and_6_14(.a(a[6]), .b(b[14]), .out(s_wallace_rca24_and_6_14));
  and_gate and_gate_s_wallace_rca24_and_5_15(.a(a[5]), .b(b[15]), .out(s_wallace_rca24_and_5_15));
  fa fa_s_wallace_rca24_fa262_out(.a(s_wallace_rca24_fa261_or0[0]), .b(s_wallace_rca24_and_6_14[0]), .cin(s_wallace_rca24_and_5_15[0]), .fa_xor1(s_wallace_rca24_fa262_xor1), .fa_or0(s_wallace_rca24_fa262_or0));
  and_gate and_gate_s_wallace_rca24_and_7_14(.a(a[7]), .b(b[14]), .out(s_wallace_rca24_and_7_14));
  and_gate and_gate_s_wallace_rca24_and_6_15(.a(a[6]), .b(b[15]), .out(s_wallace_rca24_and_6_15));
  fa fa_s_wallace_rca24_fa263_out(.a(s_wallace_rca24_fa262_or0[0]), .b(s_wallace_rca24_and_7_14[0]), .cin(s_wallace_rca24_and_6_15[0]), .fa_xor1(s_wallace_rca24_fa263_xor1), .fa_or0(s_wallace_rca24_fa263_or0));
  and_gate and_gate_s_wallace_rca24_and_8_14(.a(a[8]), .b(b[14]), .out(s_wallace_rca24_and_8_14));
  and_gate and_gate_s_wallace_rca24_and_7_15(.a(a[7]), .b(b[15]), .out(s_wallace_rca24_and_7_15));
  fa fa_s_wallace_rca24_fa264_out(.a(s_wallace_rca24_fa263_or0[0]), .b(s_wallace_rca24_and_8_14[0]), .cin(s_wallace_rca24_and_7_15[0]), .fa_xor1(s_wallace_rca24_fa264_xor1), .fa_or0(s_wallace_rca24_fa264_or0));
  and_gate and_gate_s_wallace_rca24_and_9_14(.a(a[9]), .b(b[14]), .out(s_wallace_rca24_and_9_14));
  and_gate and_gate_s_wallace_rca24_and_8_15(.a(a[8]), .b(b[15]), .out(s_wallace_rca24_and_8_15));
  fa fa_s_wallace_rca24_fa265_out(.a(s_wallace_rca24_fa264_or0[0]), .b(s_wallace_rca24_and_9_14[0]), .cin(s_wallace_rca24_and_8_15[0]), .fa_xor1(s_wallace_rca24_fa265_xor1), .fa_or0(s_wallace_rca24_fa265_or0));
  and_gate and_gate_s_wallace_rca24_and_10_14(.a(a[10]), .b(b[14]), .out(s_wallace_rca24_and_10_14));
  and_gate and_gate_s_wallace_rca24_and_9_15(.a(a[9]), .b(b[15]), .out(s_wallace_rca24_and_9_15));
  fa fa_s_wallace_rca24_fa266_out(.a(s_wallace_rca24_fa265_or0[0]), .b(s_wallace_rca24_and_10_14[0]), .cin(s_wallace_rca24_and_9_15[0]), .fa_xor1(s_wallace_rca24_fa266_xor1), .fa_or0(s_wallace_rca24_fa266_or0));
  and_gate and_gate_s_wallace_rca24_and_9_16(.a(a[9]), .b(b[16]), .out(s_wallace_rca24_and_9_16));
  and_gate and_gate_s_wallace_rca24_and_8_17(.a(a[8]), .b(b[17]), .out(s_wallace_rca24_and_8_17));
  fa fa_s_wallace_rca24_fa267_out(.a(s_wallace_rca24_fa266_or0[0]), .b(s_wallace_rca24_and_9_16[0]), .cin(s_wallace_rca24_and_8_17[0]), .fa_xor1(s_wallace_rca24_fa267_xor1), .fa_or0(s_wallace_rca24_fa267_or0));
  and_gate and_gate_s_wallace_rca24_and_9_17(.a(a[9]), .b(b[17]), .out(s_wallace_rca24_and_9_17));
  and_gate and_gate_s_wallace_rca24_and_8_18(.a(a[8]), .b(b[18]), .out(s_wallace_rca24_and_8_18));
  fa fa_s_wallace_rca24_fa268_out(.a(s_wallace_rca24_fa267_or0[0]), .b(s_wallace_rca24_and_9_17[0]), .cin(s_wallace_rca24_and_8_18[0]), .fa_xor1(s_wallace_rca24_fa268_xor1), .fa_or0(s_wallace_rca24_fa268_or0));
  and_gate and_gate_s_wallace_rca24_and_9_18(.a(a[9]), .b(b[18]), .out(s_wallace_rca24_and_9_18));
  and_gate and_gate_s_wallace_rca24_and_8_19(.a(a[8]), .b(b[19]), .out(s_wallace_rca24_and_8_19));
  fa fa_s_wallace_rca24_fa269_out(.a(s_wallace_rca24_fa268_or0[0]), .b(s_wallace_rca24_and_9_18[0]), .cin(s_wallace_rca24_and_8_19[0]), .fa_xor1(s_wallace_rca24_fa269_xor1), .fa_or0(s_wallace_rca24_fa269_or0));
  and_gate and_gate_s_wallace_rca24_and_9_19(.a(a[9]), .b(b[19]), .out(s_wallace_rca24_and_9_19));
  and_gate and_gate_s_wallace_rca24_and_8_20(.a(a[8]), .b(b[20]), .out(s_wallace_rca24_and_8_20));
  fa fa_s_wallace_rca24_fa270_out(.a(s_wallace_rca24_fa269_or0[0]), .b(s_wallace_rca24_and_9_19[0]), .cin(s_wallace_rca24_and_8_20[0]), .fa_xor1(s_wallace_rca24_fa270_xor1), .fa_or0(s_wallace_rca24_fa270_or0));
  and_gate and_gate_s_wallace_rca24_and_9_20(.a(a[9]), .b(b[20]), .out(s_wallace_rca24_and_9_20));
  and_gate and_gate_s_wallace_rca24_and_8_21(.a(a[8]), .b(b[21]), .out(s_wallace_rca24_and_8_21));
  fa fa_s_wallace_rca24_fa271_out(.a(s_wallace_rca24_fa270_or0[0]), .b(s_wallace_rca24_and_9_20[0]), .cin(s_wallace_rca24_and_8_21[0]), .fa_xor1(s_wallace_rca24_fa271_xor1), .fa_or0(s_wallace_rca24_fa271_or0));
  and_gate and_gate_s_wallace_rca24_and_9_21(.a(a[9]), .b(b[21]), .out(s_wallace_rca24_and_9_21));
  and_gate and_gate_s_wallace_rca24_and_8_22(.a(a[8]), .b(b[22]), .out(s_wallace_rca24_and_8_22));
  fa fa_s_wallace_rca24_fa272_out(.a(s_wallace_rca24_fa271_or0[0]), .b(s_wallace_rca24_and_9_21[0]), .cin(s_wallace_rca24_and_8_22[0]), .fa_xor1(s_wallace_rca24_fa272_xor1), .fa_or0(s_wallace_rca24_fa272_or0));
  and_gate and_gate_s_wallace_rca24_and_9_22(.a(a[9]), .b(b[22]), .out(s_wallace_rca24_and_9_22));
  nand_gate nand_gate_s_wallace_rca24_nand_8_23(.a(a[8]), .b(b[23]), .out(s_wallace_rca24_nand_8_23));
  fa fa_s_wallace_rca24_fa273_out(.a(s_wallace_rca24_fa272_or0[0]), .b(s_wallace_rca24_and_9_22[0]), .cin(s_wallace_rca24_nand_8_23[0]), .fa_xor1(s_wallace_rca24_fa273_xor1), .fa_or0(s_wallace_rca24_fa273_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_9_23(.a(a[9]), .b(b[23]), .out(s_wallace_rca24_nand_9_23));
  fa fa_s_wallace_rca24_fa274_out(.a(s_wallace_rca24_fa273_or0[0]), .b(s_wallace_rca24_nand_9_23[0]), .cin(s_wallace_rca24_fa29_xor1[0]), .fa_xor1(s_wallace_rca24_fa274_xor1), .fa_or0(s_wallace_rca24_fa274_or0));
  fa fa_s_wallace_rca24_fa275_out(.a(s_wallace_rca24_fa274_or0[0]), .b(s_wallace_rca24_fa30_xor1[0]), .cin(s_wallace_rca24_fa71_xor1[0]), .fa_xor1(s_wallace_rca24_fa275_xor1), .fa_or0(s_wallace_rca24_fa275_or0));
  fa fa_s_wallace_rca24_fa276_out(.a(s_wallace_rca24_fa275_or0[0]), .b(s_wallace_rca24_fa72_xor1[0]), .cin(s_wallace_rca24_fa111_xor1[0]), .fa_xor1(s_wallace_rca24_fa276_xor1), .fa_or0(s_wallace_rca24_fa276_or0));
  fa fa_s_wallace_rca24_fa277_out(.a(s_wallace_rca24_fa276_or0[0]), .b(s_wallace_rca24_fa112_xor1[0]), .cin(s_wallace_rca24_fa149_xor1[0]), .fa_xor1(s_wallace_rca24_fa277_xor1), .fa_or0(s_wallace_rca24_fa277_or0));
  fa fa_s_wallace_rca24_fa278_out(.a(s_wallace_rca24_fa277_or0[0]), .b(s_wallace_rca24_fa150_xor1[0]), .cin(s_wallace_rca24_fa185_xor1[0]), .fa_xor1(s_wallace_rca24_fa278_xor1), .fa_or0(s_wallace_rca24_fa278_or0));
  fa fa_s_wallace_rca24_fa279_out(.a(s_wallace_rca24_fa278_or0[0]), .b(s_wallace_rca24_fa186_xor1[0]), .cin(s_wallace_rca24_fa219_xor1[0]), .fa_xor1(s_wallace_rca24_fa279_xor1), .fa_or0(s_wallace_rca24_fa279_or0));
  ha ha_s_wallace_rca24_ha8_out(.a(s_wallace_rca24_fa192_xor1[0]), .b(s_wallace_rca24_fa223_xor1[0]), .ha_xor0(s_wallace_rca24_ha8_xor0), .ha_and0(s_wallace_rca24_ha8_and0));
  fa fa_s_wallace_rca24_fa280_out(.a(s_wallace_rca24_ha8_and0[0]), .b(s_wallace_rca24_fa160_xor1[0]), .cin(s_wallace_rca24_fa193_xor1[0]), .fa_xor1(s_wallace_rca24_fa280_xor1), .fa_or0(s_wallace_rca24_fa280_or0));
  fa fa_s_wallace_rca24_fa281_out(.a(s_wallace_rca24_fa280_or0[0]), .b(s_wallace_rca24_fa126_xor1[0]), .cin(s_wallace_rca24_fa161_xor1[0]), .fa_xor1(s_wallace_rca24_fa281_xor1), .fa_or0(s_wallace_rca24_fa281_or0));
  fa fa_s_wallace_rca24_fa282_out(.a(s_wallace_rca24_fa281_or0[0]), .b(s_wallace_rca24_fa90_xor1[0]), .cin(s_wallace_rca24_fa127_xor1[0]), .fa_xor1(s_wallace_rca24_fa282_xor1), .fa_or0(s_wallace_rca24_fa282_or0));
  fa fa_s_wallace_rca24_fa283_out(.a(s_wallace_rca24_fa282_or0[0]), .b(s_wallace_rca24_fa52_xor1[0]), .cin(s_wallace_rca24_fa91_xor1[0]), .fa_xor1(s_wallace_rca24_fa283_xor1), .fa_or0(s_wallace_rca24_fa283_or0));
  fa fa_s_wallace_rca24_fa284_out(.a(s_wallace_rca24_fa283_or0[0]), .b(s_wallace_rca24_fa12_xor1[0]), .cin(s_wallace_rca24_fa53_xor1[0]), .fa_xor1(s_wallace_rca24_fa284_xor1), .fa_or0(s_wallace_rca24_fa284_or0));
  and_gate and_gate_s_wallace_rca24_and_0_16(.a(a[0]), .b(b[16]), .out(s_wallace_rca24_and_0_16));
  fa fa_s_wallace_rca24_fa285_out(.a(s_wallace_rca24_fa284_or0[0]), .b(s_wallace_rca24_and_0_16[0]), .cin(s_wallace_rca24_fa13_xor1[0]), .fa_xor1(s_wallace_rca24_fa285_xor1), .fa_or0(s_wallace_rca24_fa285_or0));
  and_gate and_gate_s_wallace_rca24_and_1_16(.a(a[1]), .b(b[16]), .out(s_wallace_rca24_and_1_16));
  and_gate and_gate_s_wallace_rca24_and_0_17(.a(a[0]), .b(b[17]), .out(s_wallace_rca24_and_0_17));
  fa fa_s_wallace_rca24_fa286_out(.a(s_wallace_rca24_fa285_or0[0]), .b(s_wallace_rca24_and_1_16[0]), .cin(s_wallace_rca24_and_0_17[0]), .fa_xor1(s_wallace_rca24_fa286_xor1), .fa_or0(s_wallace_rca24_fa286_or0));
  and_gate and_gate_s_wallace_rca24_and_2_16(.a(a[2]), .b(b[16]), .out(s_wallace_rca24_and_2_16));
  and_gate and_gate_s_wallace_rca24_and_1_17(.a(a[1]), .b(b[17]), .out(s_wallace_rca24_and_1_17));
  fa fa_s_wallace_rca24_fa287_out(.a(s_wallace_rca24_fa286_or0[0]), .b(s_wallace_rca24_and_2_16[0]), .cin(s_wallace_rca24_and_1_17[0]), .fa_xor1(s_wallace_rca24_fa287_xor1), .fa_or0(s_wallace_rca24_fa287_or0));
  and_gate and_gate_s_wallace_rca24_and_3_16(.a(a[3]), .b(b[16]), .out(s_wallace_rca24_and_3_16));
  and_gate and_gate_s_wallace_rca24_and_2_17(.a(a[2]), .b(b[17]), .out(s_wallace_rca24_and_2_17));
  fa fa_s_wallace_rca24_fa288_out(.a(s_wallace_rca24_fa287_or0[0]), .b(s_wallace_rca24_and_3_16[0]), .cin(s_wallace_rca24_and_2_17[0]), .fa_xor1(s_wallace_rca24_fa288_xor1), .fa_or0(s_wallace_rca24_fa288_or0));
  and_gate and_gate_s_wallace_rca24_and_4_16(.a(a[4]), .b(b[16]), .out(s_wallace_rca24_and_4_16));
  and_gate and_gate_s_wallace_rca24_and_3_17(.a(a[3]), .b(b[17]), .out(s_wallace_rca24_and_3_17));
  fa fa_s_wallace_rca24_fa289_out(.a(s_wallace_rca24_fa288_or0[0]), .b(s_wallace_rca24_and_4_16[0]), .cin(s_wallace_rca24_and_3_17[0]), .fa_xor1(s_wallace_rca24_fa289_xor1), .fa_or0(s_wallace_rca24_fa289_or0));
  and_gate and_gate_s_wallace_rca24_and_5_16(.a(a[5]), .b(b[16]), .out(s_wallace_rca24_and_5_16));
  and_gate and_gate_s_wallace_rca24_and_4_17(.a(a[4]), .b(b[17]), .out(s_wallace_rca24_and_4_17));
  fa fa_s_wallace_rca24_fa290_out(.a(s_wallace_rca24_fa289_or0[0]), .b(s_wallace_rca24_and_5_16[0]), .cin(s_wallace_rca24_and_4_17[0]), .fa_xor1(s_wallace_rca24_fa290_xor1), .fa_or0(s_wallace_rca24_fa290_or0));
  and_gate and_gate_s_wallace_rca24_and_6_16(.a(a[6]), .b(b[16]), .out(s_wallace_rca24_and_6_16));
  and_gate and_gate_s_wallace_rca24_and_5_17(.a(a[5]), .b(b[17]), .out(s_wallace_rca24_and_5_17));
  fa fa_s_wallace_rca24_fa291_out(.a(s_wallace_rca24_fa290_or0[0]), .b(s_wallace_rca24_and_6_16[0]), .cin(s_wallace_rca24_and_5_17[0]), .fa_xor1(s_wallace_rca24_fa291_xor1), .fa_or0(s_wallace_rca24_fa291_or0));
  and_gate and_gate_s_wallace_rca24_and_7_16(.a(a[7]), .b(b[16]), .out(s_wallace_rca24_and_7_16));
  and_gate and_gate_s_wallace_rca24_and_6_17(.a(a[6]), .b(b[17]), .out(s_wallace_rca24_and_6_17));
  fa fa_s_wallace_rca24_fa292_out(.a(s_wallace_rca24_fa291_or0[0]), .b(s_wallace_rca24_and_7_16[0]), .cin(s_wallace_rca24_and_6_17[0]), .fa_xor1(s_wallace_rca24_fa292_xor1), .fa_or0(s_wallace_rca24_fa292_or0));
  and_gate and_gate_s_wallace_rca24_and_8_16(.a(a[8]), .b(b[16]), .out(s_wallace_rca24_and_8_16));
  and_gate and_gate_s_wallace_rca24_and_7_17(.a(a[7]), .b(b[17]), .out(s_wallace_rca24_and_7_17));
  fa fa_s_wallace_rca24_fa293_out(.a(s_wallace_rca24_fa292_or0[0]), .b(s_wallace_rca24_and_8_16[0]), .cin(s_wallace_rca24_and_7_17[0]), .fa_xor1(s_wallace_rca24_fa293_xor1), .fa_or0(s_wallace_rca24_fa293_or0));
  and_gate and_gate_s_wallace_rca24_and_7_18(.a(a[7]), .b(b[18]), .out(s_wallace_rca24_and_7_18));
  and_gate and_gate_s_wallace_rca24_and_6_19(.a(a[6]), .b(b[19]), .out(s_wallace_rca24_and_6_19));
  fa fa_s_wallace_rca24_fa294_out(.a(s_wallace_rca24_fa293_or0[0]), .b(s_wallace_rca24_and_7_18[0]), .cin(s_wallace_rca24_and_6_19[0]), .fa_xor1(s_wallace_rca24_fa294_xor1), .fa_or0(s_wallace_rca24_fa294_or0));
  and_gate and_gate_s_wallace_rca24_and_7_19(.a(a[7]), .b(b[19]), .out(s_wallace_rca24_and_7_19));
  and_gate and_gate_s_wallace_rca24_and_6_20(.a(a[6]), .b(b[20]), .out(s_wallace_rca24_and_6_20));
  fa fa_s_wallace_rca24_fa295_out(.a(s_wallace_rca24_fa294_or0[0]), .b(s_wallace_rca24_and_7_19[0]), .cin(s_wallace_rca24_and_6_20[0]), .fa_xor1(s_wallace_rca24_fa295_xor1), .fa_or0(s_wallace_rca24_fa295_or0));
  and_gate and_gate_s_wallace_rca24_and_7_20(.a(a[7]), .b(b[20]), .out(s_wallace_rca24_and_7_20));
  and_gate and_gate_s_wallace_rca24_and_6_21(.a(a[6]), .b(b[21]), .out(s_wallace_rca24_and_6_21));
  fa fa_s_wallace_rca24_fa296_out(.a(s_wallace_rca24_fa295_or0[0]), .b(s_wallace_rca24_and_7_20[0]), .cin(s_wallace_rca24_and_6_21[0]), .fa_xor1(s_wallace_rca24_fa296_xor1), .fa_or0(s_wallace_rca24_fa296_or0));
  and_gate and_gate_s_wallace_rca24_and_7_21(.a(a[7]), .b(b[21]), .out(s_wallace_rca24_and_7_21));
  and_gate and_gate_s_wallace_rca24_and_6_22(.a(a[6]), .b(b[22]), .out(s_wallace_rca24_and_6_22));
  fa fa_s_wallace_rca24_fa297_out(.a(s_wallace_rca24_fa296_or0[0]), .b(s_wallace_rca24_and_7_21[0]), .cin(s_wallace_rca24_and_6_22[0]), .fa_xor1(s_wallace_rca24_fa297_xor1), .fa_or0(s_wallace_rca24_fa297_or0));
  and_gate and_gate_s_wallace_rca24_and_7_22(.a(a[7]), .b(b[22]), .out(s_wallace_rca24_and_7_22));
  nand_gate nand_gate_s_wallace_rca24_nand_6_23(.a(a[6]), .b(b[23]), .out(s_wallace_rca24_nand_6_23));
  fa fa_s_wallace_rca24_fa298_out(.a(s_wallace_rca24_fa297_or0[0]), .b(s_wallace_rca24_and_7_22[0]), .cin(s_wallace_rca24_nand_6_23[0]), .fa_xor1(s_wallace_rca24_fa298_xor1), .fa_or0(s_wallace_rca24_fa298_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_7_23(.a(a[7]), .b(b[23]), .out(s_wallace_rca24_nand_7_23));
  fa fa_s_wallace_rca24_fa299_out(.a(s_wallace_rca24_fa298_or0[0]), .b(s_wallace_rca24_nand_7_23[0]), .cin(s_wallace_rca24_fa27_xor1[0]), .fa_xor1(s_wallace_rca24_fa299_xor1), .fa_or0(s_wallace_rca24_fa299_or0));
  fa fa_s_wallace_rca24_fa300_out(.a(s_wallace_rca24_fa299_or0[0]), .b(s_wallace_rca24_fa28_xor1[0]), .cin(s_wallace_rca24_fa69_xor1[0]), .fa_xor1(s_wallace_rca24_fa300_xor1), .fa_or0(s_wallace_rca24_fa300_or0));
  fa fa_s_wallace_rca24_fa301_out(.a(s_wallace_rca24_fa300_or0[0]), .b(s_wallace_rca24_fa70_xor1[0]), .cin(s_wallace_rca24_fa109_xor1[0]), .fa_xor1(s_wallace_rca24_fa301_xor1), .fa_or0(s_wallace_rca24_fa301_or0));
  fa fa_s_wallace_rca24_fa302_out(.a(s_wallace_rca24_fa301_or0[0]), .b(s_wallace_rca24_fa110_xor1[0]), .cin(s_wallace_rca24_fa147_xor1[0]), .fa_xor1(s_wallace_rca24_fa302_xor1), .fa_or0(s_wallace_rca24_fa302_or0));
  fa fa_s_wallace_rca24_fa303_out(.a(s_wallace_rca24_fa302_or0[0]), .b(s_wallace_rca24_fa148_xor1[0]), .cin(s_wallace_rca24_fa183_xor1[0]), .fa_xor1(s_wallace_rca24_fa303_xor1), .fa_or0(s_wallace_rca24_fa303_or0));
  fa fa_s_wallace_rca24_fa304_out(.a(s_wallace_rca24_fa303_or0[0]), .b(s_wallace_rca24_fa184_xor1[0]), .cin(s_wallace_rca24_fa217_xor1[0]), .fa_xor1(s_wallace_rca24_fa304_xor1), .fa_or0(s_wallace_rca24_fa304_or0));
  fa fa_s_wallace_rca24_fa305_out(.a(s_wallace_rca24_fa304_or0[0]), .b(s_wallace_rca24_fa218_xor1[0]), .cin(s_wallace_rca24_fa249_xor1[0]), .fa_xor1(s_wallace_rca24_fa305_xor1), .fa_or0(s_wallace_rca24_fa305_or0));
  ha ha_s_wallace_rca24_ha9_out(.a(s_wallace_rca24_fa224_xor1[0]), .b(s_wallace_rca24_fa253_xor1[0]), .ha_xor0(s_wallace_rca24_ha9_xor0), .ha_and0(s_wallace_rca24_ha9_and0));
  fa fa_s_wallace_rca24_fa306_out(.a(s_wallace_rca24_ha9_and0[0]), .b(s_wallace_rca24_fa194_xor1[0]), .cin(s_wallace_rca24_fa225_xor1[0]), .fa_xor1(s_wallace_rca24_fa306_xor1), .fa_or0(s_wallace_rca24_fa306_or0));
  fa fa_s_wallace_rca24_fa307_out(.a(s_wallace_rca24_fa306_or0[0]), .b(s_wallace_rca24_fa162_xor1[0]), .cin(s_wallace_rca24_fa195_xor1[0]), .fa_xor1(s_wallace_rca24_fa307_xor1), .fa_or0(s_wallace_rca24_fa307_or0));
  fa fa_s_wallace_rca24_fa308_out(.a(s_wallace_rca24_fa307_or0[0]), .b(s_wallace_rca24_fa128_xor1[0]), .cin(s_wallace_rca24_fa163_xor1[0]), .fa_xor1(s_wallace_rca24_fa308_xor1), .fa_or0(s_wallace_rca24_fa308_or0));
  fa fa_s_wallace_rca24_fa309_out(.a(s_wallace_rca24_fa308_or0[0]), .b(s_wallace_rca24_fa92_xor1[0]), .cin(s_wallace_rca24_fa129_xor1[0]), .fa_xor1(s_wallace_rca24_fa309_xor1), .fa_or0(s_wallace_rca24_fa309_or0));
  fa fa_s_wallace_rca24_fa310_out(.a(s_wallace_rca24_fa309_or0[0]), .b(s_wallace_rca24_fa54_xor1[0]), .cin(s_wallace_rca24_fa93_xor1[0]), .fa_xor1(s_wallace_rca24_fa310_xor1), .fa_or0(s_wallace_rca24_fa310_or0));
  fa fa_s_wallace_rca24_fa311_out(.a(s_wallace_rca24_fa310_or0[0]), .b(s_wallace_rca24_fa14_xor1[0]), .cin(s_wallace_rca24_fa55_xor1[0]), .fa_xor1(s_wallace_rca24_fa311_xor1), .fa_or0(s_wallace_rca24_fa311_or0));
  and_gate and_gate_s_wallace_rca24_and_0_18(.a(a[0]), .b(b[18]), .out(s_wallace_rca24_and_0_18));
  fa fa_s_wallace_rca24_fa312_out(.a(s_wallace_rca24_fa311_or0[0]), .b(s_wallace_rca24_and_0_18[0]), .cin(s_wallace_rca24_fa15_xor1[0]), .fa_xor1(s_wallace_rca24_fa312_xor1), .fa_or0(s_wallace_rca24_fa312_or0));
  and_gate and_gate_s_wallace_rca24_and_1_18(.a(a[1]), .b(b[18]), .out(s_wallace_rca24_and_1_18));
  and_gate and_gate_s_wallace_rca24_and_0_19(.a(a[0]), .b(b[19]), .out(s_wallace_rca24_and_0_19));
  fa fa_s_wallace_rca24_fa313_out(.a(s_wallace_rca24_fa312_or0[0]), .b(s_wallace_rca24_and_1_18[0]), .cin(s_wallace_rca24_and_0_19[0]), .fa_xor1(s_wallace_rca24_fa313_xor1), .fa_or0(s_wallace_rca24_fa313_or0));
  and_gate and_gate_s_wallace_rca24_and_2_18(.a(a[2]), .b(b[18]), .out(s_wallace_rca24_and_2_18));
  and_gate and_gate_s_wallace_rca24_and_1_19(.a(a[1]), .b(b[19]), .out(s_wallace_rca24_and_1_19));
  fa fa_s_wallace_rca24_fa314_out(.a(s_wallace_rca24_fa313_or0[0]), .b(s_wallace_rca24_and_2_18[0]), .cin(s_wallace_rca24_and_1_19[0]), .fa_xor1(s_wallace_rca24_fa314_xor1), .fa_or0(s_wallace_rca24_fa314_or0));
  and_gate and_gate_s_wallace_rca24_and_3_18(.a(a[3]), .b(b[18]), .out(s_wallace_rca24_and_3_18));
  and_gate and_gate_s_wallace_rca24_and_2_19(.a(a[2]), .b(b[19]), .out(s_wallace_rca24_and_2_19));
  fa fa_s_wallace_rca24_fa315_out(.a(s_wallace_rca24_fa314_or0[0]), .b(s_wallace_rca24_and_3_18[0]), .cin(s_wallace_rca24_and_2_19[0]), .fa_xor1(s_wallace_rca24_fa315_xor1), .fa_or0(s_wallace_rca24_fa315_or0));
  and_gate and_gate_s_wallace_rca24_and_4_18(.a(a[4]), .b(b[18]), .out(s_wallace_rca24_and_4_18));
  and_gate and_gate_s_wallace_rca24_and_3_19(.a(a[3]), .b(b[19]), .out(s_wallace_rca24_and_3_19));
  fa fa_s_wallace_rca24_fa316_out(.a(s_wallace_rca24_fa315_or0[0]), .b(s_wallace_rca24_and_4_18[0]), .cin(s_wallace_rca24_and_3_19[0]), .fa_xor1(s_wallace_rca24_fa316_xor1), .fa_or0(s_wallace_rca24_fa316_or0));
  and_gate and_gate_s_wallace_rca24_and_5_18(.a(a[5]), .b(b[18]), .out(s_wallace_rca24_and_5_18));
  and_gate and_gate_s_wallace_rca24_and_4_19(.a(a[4]), .b(b[19]), .out(s_wallace_rca24_and_4_19));
  fa fa_s_wallace_rca24_fa317_out(.a(s_wallace_rca24_fa316_or0[0]), .b(s_wallace_rca24_and_5_18[0]), .cin(s_wallace_rca24_and_4_19[0]), .fa_xor1(s_wallace_rca24_fa317_xor1), .fa_or0(s_wallace_rca24_fa317_or0));
  and_gate and_gate_s_wallace_rca24_and_6_18(.a(a[6]), .b(b[18]), .out(s_wallace_rca24_and_6_18));
  and_gate and_gate_s_wallace_rca24_and_5_19(.a(a[5]), .b(b[19]), .out(s_wallace_rca24_and_5_19));
  fa fa_s_wallace_rca24_fa318_out(.a(s_wallace_rca24_fa317_or0[0]), .b(s_wallace_rca24_and_6_18[0]), .cin(s_wallace_rca24_and_5_19[0]), .fa_xor1(s_wallace_rca24_fa318_xor1), .fa_or0(s_wallace_rca24_fa318_or0));
  and_gate and_gate_s_wallace_rca24_and_5_20(.a(a[5]), .b(b[20]), .out(s_wallace_rca24_and_5_20));
  and_gate and_gate_s_wallace_rca24_and_4_21(.a(a[4]), .b(b[21]), .out(s_wallace_rca24_and_4_21));
  fa fa_s_wallace_rca24_fa319_out(.a(s_wallace_rca24_fa318_or0[0]), .b(s_wallace_rca24_and_5_20[0]), .cin(s_wallace_rca24_and_4_21[0]), .fa_xor1(s_wallace_rca24_fa319_xor1), .fa_or0(s_wallace_rca24_fa319_or0));
  and_gate and_gate_s_wallace_rca24_and_5_21(.a(a[5]), .b(b[21]), .out(s_wallace_rca24_and_5_21));
  and_gate and_gate_s_wallace_rca24_and_4_22(.a(a[4]), .b(b[22]), .out(s_wallace_rca24_and_4_22));
  fa fa_s_wallace_rca24_fa320_out(.a(s_wallace_rca24_fa319_or0[0]), .b(s_wallace_rca24_and_5_21[0]), .cin(s_wallace_rca24_and_4_22[0]), .fa_xor1(s_wallace_rca24_fa320_xor1), .fa_or0(s_wallace_rca24_fa320_or0));
  and_gate and_gate_s_wallace_rca24_and_5_22(.a(a[5]), .b(b[22]), .out(s_wallace_rca24_and_5_22));
  nand_gate nand_gate_s_wallace_rca24_nand_4_23(.a(a[4]), .b(b[23]), .out(s_wallace_rca24_nand_4_23));
  fa fa_s_wallace_rca24_fa321_out(.a(s_wallace_rca24_fa320_or0[0]), .b(s_wallace_rca24_and_5_22[0]), .cin(s_wallace_rca24_nand_4_23[0]), .fa_xor1(s_wallace_rca24_fa321_xor1), .fa_or0(s_wallace_rca24_fa321_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_5_23(.a(a[5]), .b(b[23]), .out(s_wallace_rca24_nand_5_23));
  fa fa_s_wallace_rca24_fa322_out(.a(s_wallace_rca24_fa321_or0[0]), .b(s_wallace_rca24_nand_5_23[0]), .cin(s_wallace_rca24_fa25_xor1[0]), .fa_xor1(s_wallace_rca24_fa322_xor1), .fa_or0(s_wallace_rca24_fa322_or0));
  fa fa_s_wallace_rca24_fa323_out(.a(s_wallace_rca24_fa322_or0[0]), .b(s_wallace_rca24_fa26_xor1[0]), .cin(s_wallace_rca24_fa67_xor1[0]), .fa_xor1(s_wallace_rca24_fa323_xor1), .fa_or0(s_wallace_rca24_fa323_or0));
  fa fa_s_wallace_rca24_fa324_out(.a(s_wallace_rca24_fa323_or0[0]), .b(s_wallace_rca24_fa68_xor1[0]), .cin(s_wallace_rca24_fa107_xor1[0]), .fa_xor1(s_wallace_rca24_fa324_xor1), .fa_or0(s_wallace_rca24_fa324_or0));
  fa fa_s_wallace_rca24_fa325_out(.a(s_wallace_rca24_fa324_or0[0]), .b(s_wallace_rca24_fa108_xor1[0]), .cin(s_wallace_rca24_fa145_xor1[0]), .fa_xor1(s_wallace_rca24_fa325_xor1), .fa_or0(s_wallace_rca24_fa325_or0));
  fa fa_s_wallace_rca24_fa326_out(.a(s_wallace_rca24_fa325_or0[0]), .b(s_wallace_rca24_fa146_xor1[0]), .cin(s_wallace_rca24_fa181_xor1[0]), .fa_xor1(s_wallace_rca24_fa326_xor1), .fa_or0(s_wallace_rca24_fa326_or0));
  fa fa_s_wallace_rca24_fa327_out(.a(s_wallace_rca24_fa326_or0[0]), .b(s_wallace_rca24_fa182_xor1[0]), .cin(s_wallace_rca24_fa215_xor1[0]), .fa_xor1(s_wallace_rca24_fa327_xor1), .fa_or0(s_wallace_rca24_fa327_or0));
  fa fa_s_wallace_rca24_fa328_out(.a(s_wallace_rca24_fa327_or0[0]), .b(s_wallace_rca24_fa216_xor1[0]), .cin(s_wallace_rca24_fa247_xor1[0]), .fa_xor1(s_wallace_rca24_fa328_xor1), .fa_or0(s_wallace_rca24_fa328_or0));
  fa fa_s_wallace_rca24_fa329_out(.a(s_wallace_rca24_fa328_or0[0]), .b(s_wallace_rca24_fa248_xor1[0]), .cin(s_wallace_rca24_fa277_xor1[0]), .fa_xor1(s_wallace_rca24_fa329_xor1), .fa_or0(s_wallace_rca24_fa329_or0));
  ha ha_s_wallace_rca24_ha10_out(.a(s_wallace_rca24_fa254_xor1[0]), .b(s_wallace_rca24_fa281_xor1[0]), .ha_xor0(s_wallace_rca24_ha10_xor0), .ha_and0(s_wallace_rca24_ha10_and0));
  fa fa_s_wallace_rca24_fa330_out(.a(s_wallace_rca24_ha10_and0[0]), .b(s_wallace_rca24_fa226_xor1[0]), .cin(s_wallace_rca24_fa255_xor1[0]), .fa_xor1(s_wallace_rca24_fa330_xor1), .fa_or0(s_wallace_rca24_fa330_or0));
  fa fa_s_wallace_rca24_fa331_out(.a(s_wallace_rca24_fa330_or0[0]), .b(s_wallace_rca24_fa196_xor1[0]), .cin(s_wallace_rca24_fa227_xor1[0]), .fa_xor1(s_wallace_rca24_fa331_xor1), .fa_or0(s_wallace_rca24_fa331_or0));
  fa fa_s_wallace_rca24_fa332_out(.a(s_wallace_rca24_fa331_or0[0]), .b(s_wallace_rca24_fa164_xor1[0]), .cin(s_wallace_rca24_fa197_xor1[0]), .fa_xor1(s_wallace_rca24_fa332_xor1), .fa_or0(s_wallace_rca24_fa332_or0));
  fa fa_s_wallace_rca24_fa333_out(.a(s_wallace_rca24_fa332_or0[0]), .b(s_wallace_rca24_fa130_xor1[0]), .cin(s_wallace_rca24_fa165_xor1[0]), .fa_xor1(s_wallace_rca24_fa333_xor1), .fa_or0(s_wallace_rca24_fa333_or0));
  fa fa_s_wallace_rca24_fa334_out(.a(s_wallace_rca24_fa333_or0[0]), .b(s_wallace_rca24_fa94_xor1[0]), .cin(s_wallace_rca24_fa131_xor1[0]), .fa_xor1(s_wallace_rca24_fa334_xor1), .fa_or0(s_wallace_rca24_fa334_or0));
  fa fa_s_wallace_rca24_fa335_out(.a(s_wallace_rca24_fa334_or0[0]), .b(s_wallace_rca24_fa56_xor1[0]), .cin(s_wallace_rca24_fa95_xor1[0]), .fa_xor1(s_wallace_rca24_fa335_xor1), .fa_or0(s_wallace_rca24_fa335_or0));
  fa fa_s_wallace_rca24_fa336_out(.a(s_wallace_rca24_fa335_or0[0]), .b(s_wallace_rca24_fa16_xor1[0]), .cin(s_wallace_rca24_fa57_xor1[0]), .fa_xor1(s_wallace_rca24_fa336_xor1), .fa_or0(s_wallace_rca24_fa336_or0));
  and_gate and_gate_s_wallace_rca24_and_0_20(.a(a[0]), .b(b[20]), .out(s_wallace_rca24_and_0_20));
  fa fa_s_wallace_rca24_fa337_out(.a(s_wallace_rca24_fa336_or0[0]), .b(s_wallace_rca24_and_0_20[0]), .cin(s_wallace_rca24_fa17_xor1[0]), .fa_xor1(s_wallace_rca24_fa337_xor1), .fa_or0(s_wallace_rca24_fa337_or0));
  and_gate and_gate_s_wallace_rca24_and_1_20(.a(a[1]), .b(b[20]), .out(s_wallace_rca24_and_1_20));
  and_gate and_gate_s_wallace_rca24_and_0_21(.a(a[0]), .b(b[21]), .out(s_wallace_rca24_and_0_21));
  fa fa_s_wallace_rca24_fa338_out(.a(s_wallace_rca24_fa337_or0[0]), .b(s_wallace_rca24_and_1_20[0]), .cin(s_wallace_rca24_and_0_21[0]), .fa_xor1(s_wallace_rca24_fa338_xor1), .fa_or0(s_wallace_rca24_fa338_or0));
  and_gate and_gate_s_wallace_rca24_and_2_20(.a(a[2]), .b(b[20]), .out(s_wallace_rca24_and_2_20));
  and_gate and_gate_s_wallace_rca24_and_1_21(.a(a[1]), .b(b[21]), .out(s_wallace_rca24_and_1_21));
  fa fa_s_wallace_rca24_fa339_out(.a(s_wallace_rca24_fa338_or0[0]), .b(s_wallace_rca24_and_2_20[0]), .cin(s_wallace_rca24_and_1_21[0]), .fa_xor1(s_wallace_rca24_fa339_xor1), .fa_or0(s_wallace_rca24_fa339_or0));
  and_gate and_gate_s_wallace_rca24_and_3_20(.a(a[3]), .b(b[20]), .out(s_wallace_rca24_and_3_20));
  and_gate and_gate_s_wallace_rca24_and_2_21(.a(a[2]), .b(b[21]), .out(s_wallace_rca24_and_2_21));
  fa fa_s_wallace_rca24_fa340_out(.a(s_wallace_rca24_fa339_or0[0]), .b(s_wallace_rca24_and_3_20[0]), .cin(s_wallace_rca24_and_2_21[0]), .fa_xor1(s_wallace_rca24_fa340_xor1), .fa_or0(s_wallace_rca24_fa340_or0));
  and_gate and_gate_s_wallace_rca24_and_4_20(.a(a[4]), .b(b[20]), .out(s_wallace_rca24_and_4_20));
  and_gate and_gate_s_wallace_rca24_and_3_21(.a(a[3]), .b(b[21]), .out(s_wallace_rca24_and_3_21));
  fa fa_s_wallace_rca24_fa341_out(.a(s_wallace_rca24_fa340_or0[0]), .b(s_wallace_rca24_and_4_20[0]), .cin(s_wallace_rca24_and_3_21[0]), .fa_xor1(s_wallace_rca24_fa341_xor1), .fa_or0(s_wallace_rca24_fa341_or0));
  and_gate and_gate_s_wallace_rca24_and_3_22(.a(a[3]), .b(b[22]), .out(s_wallace_rca24_and_3_22));
  nand_gate nand_gate_s_wallace_rca24_nand_2_23(.a(a[2]), .b(b[23]), .out(s_wallace_rca24_nand_2_23));
  fa fa_s_wallace_rca24_fa342_out(.a(s_wallace_rca24_fa341_or0[0]), .b(s_wallace_rca24_and_3_22[0]), .cin(s_wallace_rca24_nand_2_23[0]), .fa_xor1(s_wallace_rca24_fa342_xor1), .fa_or0(s_wallace_rca24_fa342_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_3_23(.a(a[3]), .b(b[23]), .out(s_wallace_rca24_nand_3_23));
  fa fa_s_wallace_rca24_fa343_out(.a(s_wallace_rca24_fa342_or0[0]), .b(s_wallace_rca24_nand_3_23[0]), .cin(s_wallace_rca24_fa23_xor1[0]), .fa_xor1(s_wallace_rca24_fa343_xor1), .fa_or0(s_wallace_rca24_fa343_or0));
  fa fa_s_wallace_rca24_fa344_out(.a(s_wallace_rca24_fa343_or0[0]), .b(s_wallace_rca24_fa24_xor1[0]), .cin(s_wallace_rca24_fa65_xor1[0]), .fa_xor1(s_wallace_rca24_fa344_xor1), .fa_or0(s_wallace_rca24_fa344_or0));
  fa fa_s_wallace_rca24_fa345_out(.a(s_wallace_rca24_fa344_or0[0]), .b(s_wallace_rca24_fa66_xor1[0]), .cin(s_wallace_rca24_fa105_xor1[0]), .fa_xor1(s_wallace_rca24_fa345_xor1), .fa_or0(s_wallace_rca24_fa345_or0));
  fa fa_s_wallace_rca24_fa346_out(.a(s_wallace_rca24_fa345_or0[0]), .b(s_wallace_rca24_fa106_xor1[0]), .cin(s_wallace_rca24_fa143_xor1[0]), .fa_xor1(s_wallace_rca24_fa346_xor1), .fa_or0(s_wallace_rca24_fa346_or0));
  fa fa_s_wallace_rca24_fa347_out(.a(s_wallace_rca24_fa346_or0[0]), .b(s_wallace_rca24_fa144_xor1[0]), .cin(s_wallace_rca24_fa179_xor1[0]), .fa_xor1(s_wallace_rca24_fa347_xor1), .fa_or0(s_wallace_rca24_fa347_or0));
  fa fa_s_wallace_rca24_fa348_out(.a(s_wallace_rca24_fa347_or0[0]), .b(s_wallace_rca24_fa180_xor1[0]), .cin(s_wallace_rca24_fa213_xor1[0]), .fa_xor1(s_wallace_rca24_fa348_xor1), .fa_or0(s_wallace_rca24_fa348_or0));
  fa fa_s_wallace_rca24_fa349_out(.a(s_wallace_rca24_fa348_or0[0]), .b(s_wallace_rca24_fa214_xor1[0]), .cin(s_wallace_rca24_fa245_xor1[0]), .fa_xor1(s_wallace_rca24_fa349_xor1), .fa_or0(s_wallace_rca24_fa349_or0));
  fa fa_s_wallace_rca24_fa350_out(.a(s_wallace_rca24_fa349_or0[0]), .b(s_wallace_rca24_fa246_xor1[0]), .cin(s_wallace_rca24_fa275_xor1[0]), .fa_xor1(s_wallace_rca24_fa350_xor1), .fa_or0(s_wallace_rca24_fa350_or0));
  fa fa_s_wallace_rca24_fa351_out(.a(s_wallace_rca24_fa350_or0[0]), .b(s_wallace_rca24_fa276_xor1[0]), .cin(s_wallace_rca24_fa303_xor1[0]), .fa_xor1(s_wallace_rca24_fa351_xor1), .fa_or0(s_wallace_rca24_fa351_or0));
  ha ha_s_wallace_rca24_ha11_out(.a(s_wallace_rca24_fa282_xor1[0]), .b(s_wallace_rca24_fa307_xor1[0]), .ha_xor0(s_wallace_rca24_ha11_xor0), .ha_and0(s_wallace_rca24_ha11_and0));
  fa fa_s_wallace_rca24_fa352_out(.a(s_wallace_rca24_ha11_and0[0]), .b(s_wallace_rca24_fa256_xor1[0]), .cin(s_wallace_rca24_fa283_xor1[0]), .fa_xor1(s_wallace_rca24_fa352_xor1), .fa_or0(s_wallace_rca24_fa352_or0));
  fa fa_s_wallace_rca24_fa353_out(.a(s_wallace_rca24_fa352_or0[0]), .b(s_wallace_rca24_fa228_xor1[0]), .cin(s_wallace_rca24_fa257_xor1[0]), .fa_xor1(s_wallace_rca24_fa353_xor1), .fa_or0(s_wallace_rca24_fa353_or0));
  fa fa_s_wallace_rca24_fa354_out(.a(s_wallace_rca24_fa353_or0[0]), .b(s_wallace_rca24_fa198_xor1[0]), .cin(s_wallace_rca24_fa229_xor1[0]), .fa_xor1(s_wallace_rca24_fa354_xor1), .fa_or0(s_wallace_rca24_fa354_or0));
  fa fa_s_wallace_rca24_fa355_out(.a(s_wallace_rca24_fa354_or0[0]), .b(s_wallace_rca24_fa166_xor1[0]), .cin(s_wallace_rca24_fa199_xor1[0]), .fa_xor1(s_wallace_rca24_fa355_xor1), .fa_or0(s_wallace_rca24_fa355_or0));
  fa fa_s_wallace_rca24_fa356_out(.a(s_wallace_rca24_fa355_or0[0]), .b(s_wallace_rca24_fa132_xor1[0]), .cin(s_wallace_rca24_fa167_xor1[0]), .fa_xor1(s_wallace_rca24_fa356_xor1), .fa_or0(s_wallace_rca24_fa356_or0));
  fa fa_s_wallace_rca24_fa357_out(.a(s_wallace_rca24_fa356_or0[0]), .b(s_wallace_rca24_fa96_xor1[0]), .cin(s_wallace_rca24_fa133_xor1[0]), .fa_xor1(s_wallace_rca24_fa357_xor1), .fa_or0(s_wallace_rca24_fa357_or0));
  fa fa_s_wallace_rca24_fa358_out(.a(s_wallace_rca24_fa357_or0[0]), .b(s_wallace_rca24_fa58_xor1[0]), .cin(s_wallace_rca24_fa97_xor1[0]), .fa_xor1(s_wallace_rca24_fa358_xor1), .fa_or0(s_wallace_rca24_fa358_or0));
  fa fa_s_wallace_rca24_fa359_out(.a(s_wallace_rca24_fa358_or0[0]), .b(s_wallace_rca24_fa18_xor1[0]), .cin(s_wallace_rca24_fa59_xor1[0]), .fa_xor1(s_wallace_rca24_fa359_xor1), .fa_or0(s_wallace_rca24_fa359_or0));
  and_gate and_gate_s_wallace_rca24_and_0_22(.a(a[0]), .b(b[22]), .out(s_wallace_rca24_and_0_22));
  fa fa_s_wallace_rca24_fa360_out(.a(s_wallace_rca24_fa359_or0[0]), .b(s_wallace_rca24_and_0_22[0]), .cin(s_wallace_rca24_fa19_xor1[0]), .fa_xor1(s_wallace_rca24_fa360_xor1), .fa_or0(s_wallace_rca24_fa360_or0));
  and_gate and_gate_s_wallace_rca24_and_1_22(.a(a[1]), .b(b[22]), .out(s_wallace_rca24_and_1_22));
  nand_gate nand_gate_s_wallace_rca24_nand_0_23(.a(a[0]), .b(b[23]), .out(s_wallace_rca24_nand_0_23));
  fa fa_s_wallace_rca24_fa361_out(.a(s_wallace_rca24_fa360_or0[0]), .b(s_wallace_rca24_and_1_22[0]), .cin(s_wallace_rca24_nand_0_23[0]), .fa_xor1(s_wallace_rca24_fa361_xor1), .fa_or0(s_wallace_rca24_fa361_or0));
  and_gate and_gate_s_wallace_rca24_and_2_22(.a(a[2]), .b(b[22]), .out(s_wallace_rca24_and_2_22));
  nand_gate nand_gate_s_wallace_rca24_nand_1_23(.a(a[1]), .b(b[23]), .out(s_wallace_rca24_nand_1_23));
  fa fa_s_wallace_rca24_fa362_out(.a(s_wallace_rca24_fa361_or0[0]), .b(s_wallace_rca24_and_2_22[0]), .cin(s_wallace_rca24_nand_1_23[0]), .fa_xor1(s_wallace_rca24_fa362_xor1), .fa_or0(s_wallace_rca24_fa362_or0));
  fa fa_s_wallace_rca24_fa363_out(.a(s_wallace_rca24_fa362_or0[0]), .b(s_wallace_rca24_fa22_xor1[0]), .cin(s_wallace_rca24_fa63_xor1[0]), .fa_xor1(s_wallace_rca24_fa363_xor1), .fa_or0(s_wallace_rca24_fa363_or0));
  fa fa_s_wallace_rca24_fa364_out(.a(s_wallace_rca24_fa363_or0[0]), .b(s_wallace_rca24_fa64_xor1[0]), .cin(s_wallace_rca24_fa103_xor1[0]), .fa_xor1(s_wallace_rca24_fa364_xor1), .fa_or0(s_wallace_rca24_fa364_or0));
  fa fa_s_wallace_rca24_fa365_out(.a(s_wallace_rca24_fa364_or0[0]), .b(s_wallace_rca24_fa104_xor1[0]), .cin(s_wallace_rca24_fa141_xor1[0]), .fa_xor1(s_wallace_rca24_fa365_xor1), .fa_or0(s_wallace_rca24_fa365_or0));
  fa fa_s_wallace_rca24_fa366_out(.a(s_wallace_rca24_fa365_or0[0]), .b(s_wallace_rca24_fa142_xor1[0]), .cin(s_wallace_rca24_fa177_xor1[0]), .fa_xor1(s_wallace_rca24_fa366_xor1), .fa_or0(s_wallace_rca24_fa366_or0));
  fa fa_s_wallace_rca24_fa367_out(.a(s_wallace_rca24_fa366_or0[0]), .b(s_wallace_rca24_fa178_xor1[0]), .cin(s_wallace_rca24_fa211_xor1[0]), .fa_xor1(s_wallace_rca24_fa367_xor1), .fa_or0(s_wallace_rca24_fa367_or0));
  fa fa_s_wallace_rca24_fa368_out(.a(s_wallace_rca24_fa367_or0[0]), .b(s_wallace_rca24_fa212_xor1[0]), .cin(s_wallace_rca24_fa243_xor1[0]), .fa_xor1(s_wallace_rca24_fa368_xor1), .fa_or0(s_wallace_rca24_fa368_or0));
  fa fa_s_wallace_rca24_fa369_out(.a(s_wallace_rca24_fa368_or0[0]), .b(s_wallace_rca24_fa244_xor1[0]), .cin(s_wallace_rca24_fa273_xor1[0]), .fa_xor1(s_wallace_rca24_fa369_xor1), .fa_or0(s_wallace_rca24_fa369_or0));
  fa fa_s_wallace_rca24_fa370_out(.a(s_wallace_rca24_fa369_or0[0]), .b(s_wallace_rca24_fa274_xor1[0]), .cin(s_wallace_rca24_fa301_xor1[0]), .fa_xor1(s_wallace_rca24_fa370_xor1), .fa_or0(s_wallace_rca24_fa370_or0));
  fa fa_s_wallace_rca24_fa371_out(.a(s_wallace_rca24_fa370_or0[0]), .b(s_wallace_rca24_fa302_xor1[0]), .cin(s_wallace_rca24_fa327_xor1[0]), .fa_xor1(s_wallace_rca24_fa371_xor1), .fa_or0(s_wallace_rca24_fa371_or0));
  ha ha_s_wallace_rca24_ha12_out(.a(s_wallace_rca24_fa308_xor1[0]), .b(s_wallace_rca24_fa331_xor1[0]), .ha_xor0(s_wallace_rca24_ha12_xor0), .ha_and0(s_wallace_rca24_ha12_and0));
  fa fa_s_wallace_rca24_fa372_out(.a(s_wallace_rca24_ha12_and0[0]), .b(s_wallace_rca24_fa284_xor1[0]), .cin(s_wallace_rca24_fa309_xor1[0]), .fa_xor1(s_wallace_rca24_fa372_xor1), .fa_or0(s_wallace_rca24_fa372_or0));
  fa fa_s_wallace_rca24_fa373_out(.a(s_wallace_rca24_fa372_or0[0]), .b(s_wallace_rca24_fa258_xor1[0]), .cin(s_wallace_rca24_fa285_xor1[0]), .fa_xor1(s_wallace_rca24_fa373_xor1), .fa_or0(s_wallace_rca24_fa373_or0));
  fa fa_s_wallace_rca24_fa374_out(.a(s_wallace_rca24_fa373_or0[0]), .b(s_wallace_rca24_fa230_xor1[0]), .cin(s_wallace_rca24_fa259_xor1[0]), .fa_xor1(s_wallace_rca24_fa374_xor1), .fa_or0(s_wallace_rca24_fa374_or0));
  fa fa_s_wallace_rca24_fa375_out(.a(s_wallace_rca24_fa374_or0[0]), .b(s_wallace_rca24_fa200_xor1[0]), .cin(s_wallace_rca24_fa231_xor1[0]), .fa_xor1(s_wallace_rca24_fa375_xor1), .fa_or0(s_wallace_rca24_fa375_or0));
  fa fa_s_wallace_rca24_fa376_out(.a(s_wallace_rca24_fa375_or0[0]), .b(s_wallace_rca24_fa168_xor1[0]), .cin(s_wallace_rca24_fa201_xor1[0]), .fa_xor1(s_wallace_rca24_fa376_xor1), .fa_or0(s_wallace_rca24_fa376_or0));
  fa fa_s_wallace_rca24_fa377_out(.a(s_wallace_rca24_fa376_or0[0]), .b(s_wallace_rca24_fa134_xor1[0]), .cin(s_wallace_rca24_fa169_xor1[0]), .fa_xor1(s_wallace_rca24_fa377_xor1), .fa_or0(s_wallace_rca24_fa377_or0));
  fa fa_s_wallace_rca24_fa378_out(.a(s_wallace_rca24_fa377_or0[0]), .b(s_wallace_rca24_fa98_xor1[0]), .cin(s_wallace_rca24_fa135_xor1[0]), .fa_xor1(s_wallace_rca24_fa378_xor1), .fa_or0(s_wallace_rca24_fa378_or0));
  fa fa_s_wallace_rca24_fa379_out(.a(s_wallace_rca24_fa378_or0[0]), .b(s_wallace_rca24_fa60_xor1[0]), .cin(s_wallace_rca24_fa99_xor1[0]), .fa_xor1(s_wallace_rca24_fa379_xor1), .fa_or0(s_wallace_rca24_fa379_or0));
  fa fa_s_wallace_rca24_fa380_out(.a(s_wallace_rca24_fa379_or0[0]), .b(s_wallace_rca24_fa20_xor1[0]), .cin(s_wallace_rca24_fa61_xor1[0]), .fa_xor1(s_wallace_rca24_fa380_xor1), .fa_or0(s_wallace_rca24_fa380_or0));
  fa fa_s_wallace_rca24_fa381_out(.a(s_wallace_rca24_fa380_or0[0]), .b(s_wallace_rca24_fa21_xor1[0]), .cin(s_wallace_rca24_fa62_xor1[0]), .fa_xor1(s_wallace_rca24_fa381_xor1), .fa_or0(s_wallace_rca24_fa381_or0));
  fa fa_s_wallace_rca24_fa382_out(.a(s_wallace_rca24_fa381_or0[0]), .b(s_wallace_rca24_fa102_xor1[0]), .cin(s_wallace_rca24_fa139_xor1[0]), .fa_xor1(s_wallace_rca24_fa382_xor1), .fa_or0(s_wallace_rca24_fa382_or0));
  fa fa_s_wallace_rca24_fa383_out(.a(s_wallace_rca24_fa382_or0[0]), .b(s_wallace_rca24_fa140_xor1[0]), .cin(s_wallace_rca24_fa175_xor1[0]), .fa_xor1(s_wallace_rca24_fa383_xor1), .fa_or0(s_wallace_rca24_fa383_or0));
  fa fa_s_wallace_rca24_fa384_out(.a(s_wallace_rca24_fa383_or0[0]), .b(s_wallace_rca24_fa176_xor1[0]), .cin(s_wallace_rca24_fa209_xor1[0]), .fa_xor1(s_wallace_rca24_fa384_xor1), .fa_or0(s_wallace_rca24_fa384_or0));
  fa fa_s_wallace_rca24_fa385_out(.a(s_wallace_rca24_fa384_or0[0]), .b(s_wallace_rca24_fa210_xor1[0]), .cin(s_wallace_rca24_fa241_xor1[0]), .fa_xor1(s_wallace_rca24_fa385_xor1), .fa_or0(s_wallace_rca24_fa385_or0));
  fa fa_s_wallace_rca24_fa386_out(.a(s_wallace_rca24_fa385_or0[0]), .b(s_wallace_rca24_fa242_xor1[0]), .cin(s_wallace_rca24_fa271_xor1[0]), .fa_xor1(s_wallace_rca24_fa386_xor1), .fa_or0(s_wallace_rca24_fa386_or0));
  fa fa_s_wallace_rca24_fa387_out(.a(s_wallace_rca24_fa386_or0[0]), .b(s_wallace_rca24_fa272_xor1[0]), .cin(s_wallace_rca24_fa299_xor1[0]), .fa_xor1(s_wallace_rca24_fa387_xor1), .fa_or0(s_wallace_rca24_fa387_or0));
  fa fa_s_wallace_rca24_fa388_out(.a(s_wallace_rca24_fa387_or0[0]), .b(s_wallace_rca24_fa300_xor1[0]), .cin(s_wallace_rca24_fa325_xor1[0]), .fa_xor1(s_wallace_rca24_fa388_xor1), .fa_or0(s_wallace_rca24_fa388_or0));
  fa fa_s_wallace_rca24_fa389_out(.a(s_wallace_rca24_fa388_or0[0]), .b(s_wallace_rca24_fa326_xor1[0]), .cin(s_wallace_rca24_fa349_xor1[0]), .fa_xor1(s_wallace_rca24_fa389_xor1), .fa_or0(s_wallace_rca24_fa389_or0));
  ha ha_s_wallace_rca24_ha13_out(.a(s_wallace_rca24_fa332_xor1[0]), .b(s_wallace_rca24_fa353_xor1[0]), .ha_xor0(s_wallace_rca24_ha13_xor0), .ha_and0(s_wallace_rca24_ha13_and0));
  fa fa_s_wallace_rca24_fa390_out(.a(s_wallace_rca24_ha13_and0[0]), .b(s_wallace_rca24_fa310_xor1[0]), .cin(s_wallace_rca24_fa333_xor1[0]), .fa_xor1(s_wallace_rca24_fa390_xor1), .fa_or0(s_wallace_rca24_fa390_or0));
  fa fa_s_wallace_rca24_fa391_out(.a(s_wallace_rca24_fa390_or0[0]), .b(s_wallace_rca24_fa286_xor1[0]), .cin(s_wallace_rca24_fa311_xor1[0]), .fa_xor1(s_wallace_rca24_fa391_xor1), .fa_or0(s_wallace_rca24_fa391_or0));
  fa fa_s_wallace_rca24_fa392_out(.a(s_wallace_rca24_fa391_or0[0]), .b(s_wallace_rca24_fa260_xor1[0]), .cin(s_wallace_rca24_fa287_xor1[0]), .fa_xor1(s_wallace_rca24_fa392_xor1), .fa_or0(s_wallace_rca24_fa392_or0));
  fa fa_s_wallace_rca24_fa393_out(.a(s_wallace_rca24_fa392_or0[0]), .b(s_wallace_rca24_fa232_xor1[0]), .cin(s_wallace_rca24_fa261_xor1[0]), .fa_xor1(s_wallace_rca24_fa393_xor1), .fa_or0(s_wallace_rca24_fa393_or0));
  fa fa_s_wallace_rca24_fa394_out(.a(s_wallace_rca24_fa393_or0[0]), .b(s_wallace_rca24_fa202_xor1[0]), .cin(s_wallace_rca24_fa233_xor1[0]), .fa_xor1(s_wallace_rca24_fa394_xor1), .fa_or0(s_wallace_rca24_fa394_or0));
  fa fa_s_wallace_rca24_fa395_out(.a(s_wallace_rca24_fa394_or0[0]), .b(s_wallace_rca24_fa170_xor1[0]), .cin(s_wallace_rca24_fa203_xor1[0]), .fa_xor1(s_wallace_rca24_fa395_xor1), .fa_or0(s_wallace_rca24_fa395_or0));
  fa fa_s_wallace_rca24_fa396_out(.a(s_wallace_rca24_fa395_or0[0]), .b(s_wallace_rca24_fa136_xor1[0]), .cin(s_wallace_rca24_fa171_xor1[0]), .fa_xor1(s_wallace_rca24_fa396_xor1), .fa_or0(s_wallace_rca24_fa396_or0));
  fa fa_s_wallace_rca24_fa397_out(.a(s_wallace_rca24_fa396_or0[0]), .b(s_wallace_rca24_fa100_xor1[0]), .cin(s_wallace_rca24_fa137_xor1[0]), .fa_xor1(s_wallace_rca24_fa397_xor1), .fa_or0(s_wallace_rca24_fa397_or0));
  fa fa_s_wallace_rca24_fa398_out(.a(s_wallace_rca24_fa397_or0[0]), .b(s_wallace_rca24_fa101_xor1[0]), .cin(s_wallace_rca24_fa138_xor1[0]), .fa_xor1(s_wallace_rca24_fa398_xor1), .fa_or0(s_wallace_rca24_fa398_or0));
  fa fa_s_wallace_rca24_fa399_out(.a(s_wallace_rca24_fa398_or0[0]), .b(s_wallace_rca24_fa174_xor1[0]), .cin(s_wallace_rca24_fa207_xor1[0]), .fa_xor1(s_wallace_rca24_fa399_xor1), .fa_or0(s_wallace_rca24_fa399_or0));
  fa fa_s_wallace_rca24_fa400_out(.a(s_wallace_rca24_fa399_or0[0]), .b(s_wallace_rca24_fa208_xor1[0]), .cin(s_wallace_rca24_fa239_xor1[0]), .fa_xor1(s_wallace_rca24_fa400_xor1), .fa_or0(s_wallace_rca24_fa400_or0));
  fa fa_s_wallace_rca24_fa401_out(.a(s_wallace_rca24_fa400_or0[0]), .b(s_wallace_rca24_fa240_xor1[0]), .cin(s_wallace_rca24_fa269_xor1[0]), .fa_xor1(s_wallace_rca24_fa401_xor1), .fa_or0(s_wallace_rca24_fa401_or0));
  fa fa_s_wallace_rca24_fa402_out(.a(s_wallace_rca24_fa401_or0[0]), .b(s_wallace_rca24_fa270_xor1[0]), .cin(s_wallace_rca24_fa297_xor1[0]), .fa_xor1(s_wallace_rca24_fa402_xor1), .fa_or0(s_wallace_rca24_fa402_or0));
  fa fa_s_wallace_rca24_fa403_out(.a(s_wallace_rca24_fa402_or0[0]), .b(s_wallace_rca24_fa298_xor1[0]), .cin(s_wallace_rca24_fa323_xor1[0]), .fa_xor1(s_wallace_rca24_fa403_xor1), .fa_or0(s_wallace_rca24_fa403_or0));
  fa fa_s_wallace_rca24_fa404_out(.a(s_wallace_rca24_fa403_or0[0]), .b(s_wallace_rca24_fa324_xor1[0]), .cin(s_wallace_rca24_fa347_xor1[0]), .fa_xor1(s_wallace_rca24_fa404_xor1), .fa_or0(s_wallace_rca24_fa404_or0));
  fa fa_s_wallace_rca24_fa405_out(.a(s_wallace_rca24_fa404_or0[0]), .b(s_wallace_rca24_fa348_xor1[0]), .cin(s_wallace_rca24_fa369_xor1[0]), .fa_xor1(s_wallace_rca24_fa405_xor1), .fa_or0(s_wallace_rca24_fa405_or0));
  ha ha_s_wallace_rca24_ha14_out(.a(s_wallace_rca24_fa354_xor1[0]), .b(s_wallace_rca24_fa373_xor1[0]), .ha_xor0(s_wallace_rca24_ha14_xor0), .ha_and0(s_wallace_rca24_ha14_and0));
  fa fa_s_wallace_rca24_fa406_out(.a(s_wallace_rca24_ha14_and0[0]), .b(s_wallace_rca24_fa334_xor1[0]), .cin(s_wallace_rca24_fa355_xor1[0]), .fa_xor1(s_wallace_rca24_fa406_xor1), .fa_or0(s_wallace_rca24_fa406_or0));
  fa fa_s_wallace_rca24_fa407_out(.a(s_wallace_rca24_fa406_or0[0]), .b(s_wallace_rca24_fa312_xor1[0]), .cin(s_wallace_rca24_fa335_xor1[0]), .fa_xor1(s_wallace_rca24_fa407_xor1), .fa_or0(s_wallace_rca24_fa407_or0));
  fa fa_s_wallace_rca24_fa408_out(.a(s_wallace_rca24_fa407_or0[0]), .b(s_wallace_rca24_fa288_xor1[0]), .cin(s_wallace_rca24_fa313_xor1[0]), .fa_xor1(s_wallace_rca24_fa408_xor1), .fa_or0(s_wallace_rca24_fa408_or0));
  fa fa_s_wallace_rca24_fa409_out(.a(s_wallace_rca24_fa408_or0[0]), .b(s_wallace_rca24_fa262_xor1[0]), .cin(s_wallace_rca24_fa289_xor1[0]), .fa_xor1(s_wallace_rca24_fa409_xor1), .fa_or0(s_wallace_rca24_fa409_or0));
  fa fa_s_wallace_rca24_fa410_out(.a(s_wallace_rca24_fa409_or0[0]), .b(s_wallace_rca24_fa234_xor1[0]), .cin(s_wallace_rca24_fa263_xor1[0]), .fa_xor1(s_wallace_rca24_fa410_xor1), .fa_or0(s_wallace_rca24_fa410_or0));
  fa fa_s_wallace_rca24_fa411_out(.a(s_wallace_rca24_fa410_or0[0]), .b(s_wallace_rca24_fa204_xor1[0]), .cin(s_wallace_rca24_fa235_xor1[0]), .fa_xor1(s_wallace_rca24_fa411_xor1), .fa_or0(s_wallace_rca24_fa411_or0));
  fa fa_s_wallace_rca24_fa412_out(.a(s_wallace_rca24_fa411_or0[0]), .b(s_wallace_rca24_fa172_xor1[0]), .cin(s_wallace_rca24_fa205_xor1[0]), .fa_xor1(s_wallace_rca24_fa412_xor1), .fa_or0(s_wallace_rca24_fa412_or0));
  fa fa_s_wallace_rca24_fa413_out(.a(s_wallace_rca24_fa412_or0[0]), .b(s_wallace_rca24_fa173_xor1[0]), .cin(s_wallace_rca24_fa206_xor1[0]), .fa_xor1(s_wallace_rca24_fa413_xor1), .fa_or0(s_wallace_rca24_fa413_or0));
  fa fa_s_wallace_rca24_fa414_out(.a(s_wallace_rca24_fa413_or0[0]), .b(s_wallace_rca24_fa238_xor1[0]), .cin(s_wallace_rca24_fa267_xor1[0]), .fa_xor1(s_wallace_rca24_fa414_xor1), .fa_or0(s_wallace_rca24_fa414_or0));
  fa fa_s_wallace_rca24_fa415_out(.a(s_wallace_rca24_fa414_or0[0]), .b(s_wallace_rca24_fa268_xor1[0]), .cin(s_wallace_rca24_fa295_xor1[0]), .fa_xor1(s_wallace_rca24_fa415_xor1), .fa_or0(s_wallace_rca24_fa415_or0));
  fa fa_s_wallace_rca24_fa416_out(.a(s_wallace_rca24_fa415_or0[0]), .b(s_wallace_rca24_fa296_xor1[0]), .cin(s_wallace_rca24_fa321_xor1[0]), .fa_xor1(s_wallace_rca24_fa416_xor1), .fa_or0(s_wallace_rca24_fa416_or0));
  fa fa_s_wallace_rca24_fa417_out(.a(s_wallace_rca24_fa416_or0[0]), .b(s_wallace_rca24_fa322_xor1[0]), .cin(s_wallace_rca24_fa345_xor1[0]), .fa_xor1(s_wallace_rca24_fa417_xor1), .fa_or0(s_wallace_rca24_fa417_or0));
  fa fa_s_wallace_rca24_fa418_out(.a(s_wallace_rca24_fa417_or0[0]), .b(s_wallace_rca24_fa346_xor1[0]), .cin(s_wallace_rca24_fa367_xor1[0]), .fa_xor1(s_wallace_rca24_fa418_xor1), .fa_or0(s_wallace_rca24_fa418_or0));
  fa fa_s_wallace_rca24_fa419_out(.a(s_wallace_rca24_fa418_or0[0]), .b(s_wallace_rca24_fa368_xor1[0]), .cin(s_wallace_rca24_fa387_xor1[0]), .fa_xor1(s_wallace_rca24_fa419_xor1), .fa_or0(s_wallace_rca24_fa419_or0));
  ha ha_s_wallace_rca24_ha15_out(.a(s_wallace_rca24_fa374_xor1[0]), .b(s_wallace_rca24_fa391_xor1[0]), .ha_xor0(s_wallace_rca24_ha15_xor0), .ha_and0(s_wallace_rca24_ha15_and0));
  fa fa_s_wallace_rca24_fa420_out(.a(s_wallace_rca24_ha15_and0[0]), .b(s_wallace_rca24_fa356_xor1[0]), .cin(s_wallace_rca24_fa375_xor1[0]), .fa_xor1(s_wallace_rca24_fa420_xor1), .fa_or0(s_wallace_rca24_fa420_or0));
  fa fa_s_wallace_rca24_fa421_out(.a(s_wallace_rca24_fa420_or0[0]), .b(s_wallace_rca24_fa336_xor1[0]), .cin(s_wallace_rca24_fa357_xor1[0]), .fa_xor1(s_wallace_rca24_fa421_xor1), .fa_or0(s_wallace_rca24_fa421_or0));
  fa fa_s_wallace_rca24_fa422_out(.a(s_wallace_rca24_fa421_or0[0]), .b(s_wallace_rca24_fa314_xor1[0]), .cin(s_wallace_rca24_fa337_xor1[0]), .fa_xor1(s_wallace_rca24_fa422_xor1), .fa_or0(s_wallace_rca24_fa422_or0));
  fa fa_s_wallace_rca24_fa423_out(.a(s_wallace_rca24_fa422_or0[0]), .b(s_wallace_rca24_fa290_xor1[0]), .cin(s_wallace_rca24_fa315_xor1[0]), .fa_xor1(s_wallace_rca24_fa423_xor1), .fa_or0(s_wallace_rca24_fa423_or0));
  fa fa_s_wallace_rca24_fa424_out(.a(s_wallace_rca24_fa423_or0[0]), .b(s_wallace_rca24_fa264_xor1[0]), .cin(s_wallace_rca24_fa291_xor1[0]), .fa_xor1(s_wallace_rca24_fa424_xor1), .fa_or0(s_wallace_rca24_fa424_or0));
  fa fa_s_wallace_rca24_fa425_out(.a(s_wallace_rca24_fa424_or0[0]), .b(s_wallace_rca24_fa236_xor1[0]), .cin(s_wallace_rca24_fa265_xor1[0]), .fa_xor1(s_wallace_rca24_fa425_xor1), .fa_or0(s_wallace_rca24_fa425_or0));
  fa fa_s_wallace_rca24_fa426_out(.a(s_wallace_rca24_fa425_or0[0]), .b(s_wallace_rca24_fa237_xor1[0]), .cin(s_wallace_rca24_fa266_xor1[0]), .fa_xor1(s_wallace_rca24_fa426_xor1), .fa_or0(s_wallace_rca24_fa426_or0));
  fa fa_s_wallace_rca24_fa427_out(.a(s_wallace_rca24_fa426_or0[0]), .b(s_wallace_rca24_fa294_xor1[0]), .cin(s_wallace_rca24_fa319_xor1[0]), .fa_xor1(s_wallace_rca24_fa427_xor1), .fa_or0(s_wallace_rca24_fa427_or0));
  fa fa_s_wallace_rca24_fa428_out(.a(s_wallace_rca24_fa427_or0[0]), .b(s_wallace_rca24_fa320_xor1[0]), .cin(s_wallace_rca24_fa343_xor1[0]), .fa_xor1(s_wallace_rca24_fa428_xor1), .fa_or0(s_wallace_rca24_fa428_or0));
  fa fa_s_wallace_rca24_fa429_out(.a(s_wallace_rca24_fa428_or0[0]), .b(s_wallace_rca24_fa344_xor1[0]), .cin(s_wallace_rca24_fa365_xor1[0]), .fa_xor1(s_wallace_rca24_fa429_xor1), .fa_or0(s_wallace_rca24_fa429_or0));
  fa fa_s_wallace_rca24_fa430_out(.a(s_wallace_rca24_fa429_or0[0]), .b(s_wallace_rca24_fa366_xor1[0]), .cin(s_wallace_rca24_fa385_xor1[0]), .fa_xor1(s_wallace_rca24_fa430_xor1), .fa_or0(s_wallace_rca24_fa430_or0));
  fa fa_s_wallace_rca24_fa431_out(.a(s_wallace_rca24_fa430_or0[0]), .b(s_wallace_rca24_fa386_xor1[0]), .cin(s_wallace_rca24_fa403_xor1[0]), .fa_xor1(s_wallace_rca24_fa431_xor1), .fa_or0(s_wallace_rca24_fa431_or0));
  ha ha_s_wallace_rca24_ha16_out(.a(s_wallace_rca24_fa392_xor1[0]), .b(s_wallace_rca24_fa407_xor1[0]), .ha_xor0(s_wallace_rca24_ha16_xor0), .ha_and0(s_wallace_rca24_ha16_and0));
  fa fa_s_wallace_rca24_fa432_out(.a(s_wallace_rca24_ha16_and0[0]), .b(s_wallace_rca24_fa376_xor1[0]), .cin(s_wallace_rca24_fa393_xor1[0]), .fa_xor1(s_wallace_rca24_fa432_xor1), .fa_or0(s_wallace_rca24_fa432_or0));
  fa fa_s_wallace_rca24_fa433_out(.a(s_wallace_rca24_fa432_or0[0]), .b(s_wallace_rca24_fa358_xor1[0]), .cin(s_wallace_rca24_fa377_xor1[0]), .fa_xor1(s_wallace_rca24_fa433_xor1), .fa_or0(s_wallace_rca24_fa433_or0));
  fa fa_s_wallace_rca24_fa434_out(.a(s_wallace_rca24_fa433_or0[0]), .b(s_wallace_rca24_fa338_xor1[0]), .cin(s_wallace_rca24_fa359_xor1[0]), .fa_xor1(s_wallace_rca24_fa434_xor1), .fa_or0(s_wallace_rca24_fa434_or0));
  fa fa_s_wallace_rca24_fa435_out(.a(s_wallace_rca24_fa434_or0[0]), .b(s_wallace_rca24_fa316_xor1[0]), .cin(s_wallace_rca24_fa339_xor1[0]), .fa_xor1(s_wallace_rca24_fa435_xor1), .fa_or0(s_wallace_rca24_fa435_or0));
  fa fa_s_wallace_rca24_fa436_out(.a(s_wallace_rca24_fa435_or0[0]), .b(s_wallace_rca24_fa292_xor1[0]), .cin(s_wallace_rca24_fa317_xor1[0]), .fa_xor1(s_wallace_rca24_fa436_xor1), .fa_or0(s_wallace_rca24_fa436_or0));
  fa fa_s_wallace_rca24_fa437_out(.a(s_wallace_rca24_fa436_or0[0]), .b(s_wallace_rca24_fa293_xor1[0]), .cin(s_wallace_rca24_fa318_xor1[0]), .fa_xor1(s_wallace_rca24_fa437_xor1), .fa_or0(s_wallace_rca24_fa437_or0));
  fa fa_s_wallace_rca24_fa438_out(.a(s_wallace_rca24_fa437_or0[0]), .b(s_wallace_rca24_fa342_xor1[0]), .cin(s_wallace_rca24_fa363_xor1[0]), .fa_xor1(s_wallace_rca24_fa438_xor1), .fa_or0(s_wallace_rca24_fa438_or0));
  fa fa_s_wallace_rca24_fa439_out(.a(s_wallace_rca24_fa438_or0[0]), .b(s_wallace_rca24_fa364_xor1[0]), .cin(s_wallace_rca24_fa383_xor1[0]), .fa_xor1(s_wallace_rca24_fa439_xor1), .fa_or0(s_wallace_rca24_fa439_or0));
  fa fa_s_wallace_rca24_fa440_out(.a(s_wallace_rca24_fa439_or0[0]), .b(s_wallace_rca24_fa384_xor1[0]), .cin(s_wallace_rca24_fa401_xor1[0]), .fa_xor1(s_wallace_rca24_fa440_xor1), .fa_or0(s_wallace_rca24_fa440_or0));
  fa fa_s_wallace_rca24_fa441_out(.a(s_wallace_rca24_fa440_or0[0]), .b(s_wallace_rca24_fa402_xor1[0]), .cin(s_wallace_rca24_fa417_xor1[0]), .fa_xor1(s_wallace_rca24_fa441_xor1), .fa_or0(s_wallace_rca24_fa441_or0));
  ha ha_s_wallace_rca24_ha17_out(.a(s_wallace_rca24_fa408_xor1[0]), .b(s_wallace_rca24_fa421_xor1[0]), .ha_xor0(s_wallace_rca24_ha17_xor0), .ha_and0(s_wallace_rca24_ha17_and0));
  fa fa_s_wallace_rca24_fa442_out(.a(s_wallace_rca24_ha17_and0[0]), .b(s_wallace_rca24_fa394_xor1[0]), .cin(s_wallace_rca24_fa409_xor1[0]), .fa_xor1(s_wallace_rca24_fa442_xor1), .fa_or0(s_wallace_rca24_fa442_or0));
  fa fa_s_wallace_rca24_fa443_out(.a(s_wallace_rca24_fa442_or0[0]), .b(s_wallace_rca24_fa378_xor1[0]), .cin(s_wallace_rca24_fa395_xor1[0]), .fa_xor1(s_wallace_rca24_fa443_xor1), .fa_or0(s_wallace_rca24_fa443_or0));
  fa fa_s_wallace_rca24_fa444_out(.a(s_wallace_rca24_fa443_or0[0]), .b(s_wallace_rca24_fa360_xor1[0]), .cin(s_wallace_rca24_fa379_xor1[0]), .fa_xor1(s_wallace_rca24_fa444_xor1), .fa_or0(s_wallace_rca24_fa444_or0));
  fa fa_s_wallace_rca24_fa445_out(.a(s_wallace_rca24_fa444_or0[0]), .b(s_wallace_rca24_fa340_xor1[0]), .cin(s_wallace_rca24_fa361_xor1[0]), .fa_xor1(s_wallace_rca24_fa445_xor1), .fa_or0(s_wallace_rca24_fa445_or0));
  fa fa_s_wallace_rca24_fa446_out(.a(s_wallace_rca24_fa445_or0[0]), .b(s_wallace_rca24_fa341_xor1[0]), .cin(s_wallace_rca24_fa362_xor1[0]), .fa_xor1(s_wallace_rca24_fa446_xor1), .fa_or0(s_wallace_rca24_fa446_or0));
  fa fa_s_wallace_rca24_fa447_out(.a(s_wallace_rca24_fa446_or0[0]), .b(s_wallace_rca24_fa382_xor1[0]), .cin(s_wallace_rca24_fa399_xor1[0]), .fa_xor1(s_wallace_rca24_fa447_xor1), .fa_or0(s_wallace_rca24_fa447_or0));
  fa fa_s_wallace_rca24_fa448_out(.a(s_wallace_rca24_fa447_or0[0]), .b(s_wallace_rca24_fa400_xor1[0]), .cin(s_wallace_rca24_fa415_xor1[0]), .fa_xor1(s_wallace_rca24_fa448_xor1), .fa_or0(s_wallace_rca24_fa448_or0));
  fa fa_s_wallace_rca24_fa449_out(.a(s_wallace_rca24_fa448_or0[0]), .b(s_wallace_rca24_fa416_xor1[0]), .cin(s_wallace_rca24_fa429_xor1[0]), .fa_xor1(s_wallace_rca24_fa449_xor1), .fa_or0(s_wallace_rca24_fa449_or0));
  ha ha_s_wallace_rca24_ha18_out(.a(s_wallace_rca24_fa422_xor1[0]), .b(s_wallace_rca24_fa433_xor1[0]), .ha_xor0(s_wallace_rca24_ha18_xor0), .ha_and0(s_wallace_rca24_ha18_and0));
  fa fa_s_wallace_rca24_fa450_out(.a(s_wallace_rca24_ha18_and0[0]), .b(s_wallace_rca24_fa410_xor1[0]), .cin(s_wallace_rca24_fa423_xor1[0]), .fa_xor1(s_wallace_rca24_fa450_xor1), .fa_or0(s_wallace_rca24_fa450_or0));
  fa fa_s_wallace_rca24_fa451_out(.a(s_wallace_rca24_fa450_or0[0]), .b(s_wallace_rca24_fa396_xor1[0]), .cin(s_wallace_rca24_fa411_xor1[0]), .fa_xor1(s_wallace_rca24_fa451_xor1), .fa_or0(s_wallace_rca24_fa451_or0));
  fa fa_s_wallace_rca24_fa452_out(.a(s_wallace_rca24_fa451_or0[0]), .b(s_wallace_rca24_fa380_xor1[0]), .cin(s_wallace_rca24_fa397_xor1[0]), .fa_xor1(s_wallace_rca24_fa452_xor1), .fa_or0(s_wallace_rca24_fa452_or0));
  fa fa_s_wallace_rca24_fa453_out(.a(s_wallace_rca24_fa452_or0[0]), .b(s_wallace_rca24_fa381_xor1[0]), .cin(s_wallace_rca24_fa398_xor1[0]), .fa_xor1(s_wallace_rca24_fa453_xor1), .fa_or0(s_wallace_rca24_fa453_or0));
  fa fa_s_wallace_rca24_fa454_out(.a(s_wallace_rca24_fa453_or0[0]), .b(s_wallace_rca24_fa414_xor1[0]), .cin(s_wallace_rca24_fa427_xor1[0]), .fa_xor1(s_wallace_rca24_fa454_xor1), .fa_or0(s_wallace_rca24_fa454_or0));
  fa fa_s_wallace_rca24_fa455_out(.a(s_wallace_rca24_fa454_or0[0]), .b(s_wallace_rca24_fa428_xor1[0]), .cin(s_wallace_rca24_fa439_xor1[0]), .fa_xor1(s_wallace_rca24_fa455_xor1), .fa_or0(s_wallace_rca24_fa455_or0));
  ha ha_s_wallace_rca24_ha19_out(.a(s_wallace_rca24_fa434_xor1[0]), .b(s_wallace_rca24_fa443_xor1[0]), .ha_xor0(s_wallace_rca24_ha19_xor0), .ha_and0(s_wallace_rca24_ha19_and0));
  fa fa_s_wallace_rca24_fa456_out(.a(s_wallace_rca24_ha19_and0[0]), .b(s_wallace_rca24_fa424_xor1[0]), .cin(s_wallace_rca24_fa435_xor1[0]), .fa_xor1(s_wallace_rca24_fa456_xor1), .fa_or0(s_wallace_rca24_fa456_or0));
  fa fa_s_wallace_rca24_fa457_out(.a(s_wallace_rca24_fa456_or0[0]), .b(s_wallace_rca24_fa412_xor1[0]), .cin(s_wallace_rca24_fa425_xor1[0]), .fa_xor1(s_wallace_rca24_fa457_xor1), .fa_or0(s_wallace_rca24_fa457_or0));
  fa fa_s_wallace_rca24_fa458_out(.a(s_wallace_rca24_fa457_or0[0]), .b(s_wallace_rca24_fa413_xor1[0]), .cin(s_wallace_rca24_fa426_xor1[0]), .fa_xor1(s_wallace_rca24_fa458_xor1), .fa_or0(s_wallace_rca24_fa458_or0));
  fa fa_s_wallace_rca24_fa459_out(.a(s_wallace_rca24_fa458_or0[0]), .b(s_wallace_rca24_fa438_xor1[0]), .cin(s_wallace_rca24_fa447_xor1[0]), .fa_xor1(s_wallace_rca24_fa459_xor1), .fa_or0(s_wallace_rca24_fa459_or0));
  ha ha_s_wallace_rca24_ha20_out(.a(s_wallace_rca24_fa444_xor1[0]), .b(s_wallace_rca24_fa451_xor1[0]), .ha_xor0(s_wallace_rca24_ha20_xor0), .ha_and0(s_wallace_rca24_ha20_and0));
  fa fa_s_wallace_rca24_fa460_out(.a(s_wallace_rca24_ha20_and0[0]), .b(s_wallace_rca24_fa436_xor1[0]), .cin(s_wallace_rca24_fa445_xor1[0]), .fa_xor1(s_wallace_rca24_fa460_xor1), .fa_or0(s_wallace_rca24_fa460_or0));
  fa fa_s_wallace_rca24_fa461_out(.a(s_wallace_rca24_fa460_or0[0]), .b(s_wallace_rca24_fa437_xor1[0]), .cin(s_wallace_rca24_fa446_xor1[0]), .fa_xor1(s_wallace_rca24_fa461_xor1), .fa_or0(s_wallace_rca24_fa461_or0));
  ha ha_s_wallace_rca24_ha21_out(.a(s_wallace_rca24_fa452_xor1[0]), .b(s_wallace_rca24_fa457_xor1[0]), .ha_xor0(s_wallace_rca24_ha21_xor0), .ha_and0(s_wallace_rca24_ha21_and0));
  fa fa_s_wallace_rca24_fa462_out(.a(s_wallace_rca24_ha21_and0[0]), .b(s_wallace_rca24_fa453_xor1[0]), .cin(s_wallace_rca24_fa458_xor1[0]), .fa_xor1(s_wallace_rca24_fa462_xor1), .fa_or0(s_wallace_rca24_fa462_or0));
  fa fa_s_wallace_rca24_fa463_out(.a(s_wallace_rca24_fa462_or0[0]), .b(s_wallace_rca24_fa461_or0[0]), .cin(s_wallace_rca24_fa454_xor1[0]), .fa_xor1(s_wallace_rca24_fa463_xor1), .fa_or0(s_wallace_rca24_fa463_or0));
  fa fa_s_wallace_rca24_fa464_out(.a(s_wallace_rca24_fa463_or0[0]), .b(s_wallace_rca24_fa459_or0[0]), .cin(s_wallace_rca24_fa448_xor1[0]), .fa_xor1(s_wallace_rca24_fa464_xor1), .fa_or0(s_wallace_rca24_fa464_or0));
  fa fa_s_wallace_rca24_fa465_out(.a(s_wallace_rca24_fa464_or0[0]), .b(s_wallace_rca24_fa455_or0[0]), .cin(s_wallace_rca24_fa440_xor1[0]), .fa_xor1(s_wallace_rca24_fa465_xor1), .fa_or0(s_wallace_rca24_fa465_or0));
  fa fa_s_wallace_rca24_fa466_out(.a(s_wallace_rca24_fa465_or0[0]), .b(s_wallace_rca24_fa449_or0[0]), .cin(s_wallace_rca24_fa430_xor1[0]), .fa_xor1(s_wallace_rca24_fa466_xor1), .fa_or0(s_wallace_rca24_fa466_or0));
  fa fa_s_wallace_rca24_fa467_out(.a(s_wallace_rca24_fa466_or0[0]), .b(s_wallace_rca24_fa441_or0[0]), .cin(s_wallace_rca24_fa418_xor1[0]), .fa_xor1(s_wallace_rca24_fa467_xor1), .fa_or0(s_wallace_rca24_fa467_or0));
  fa fa_s_wallace_rca24_fa468_out(.a(s_wallace_rca24_fa467_or0[0]), .b(s_wallace_rca24_fa431_or0[0]), .cin(s_wallace_rca24_fa404_xor1[0]), .fa_xor1(s_wallace_rca24_fa468_xor1), .fa_or0(s_wallace_rca24_fa468_or0));
  fa fa_s_wallace_rca24_fa469_out(.a(s_wallace_rca24_fa468_or0[0]), .b(s_wallace_rca24_fa419_or0[0]), .cin(s_wallace_rca24_fa388_xor1[0]), .fa_xor1(s_wallace_rca24_fa469_xor1), .fa_or0(s_wallace_rca24_fa469_or0));
  fa fa_s_wallace_rca24_fa470_out(.a(s_wallace_rca24_fa469_or0[0]), .b(s_wallace_rca24_fa405_or0[0]), .cin(s_wallace_rca24_fa370_xor1[0]), .fa_xor1(s_wallace_rca24_fa470_xor1), .fa_or0(s_wallace_rca24_fa470_or0));
  fa fa_s_wallace_rca24_fa471_out(.a(s_wallace_rca24_fa470_or0[0]), .b(s_wallace_rca24_fa389_or0[0]), .cin(s_wallace_rca24_fa350_xor1[0]), .fa_xor1(s_wallace_rca24_fa471_xor1), .fa_or0(s_wallace_rca24_fa471_or0));
  fa fa_s_wallace_rca24_fa472_out(.a(s_wallace_rca24_fa471_or0[0]), .b(s_wallace_rca24_fa371_or0[0]), .cin(s_wallace_rca24_fa328_xor1[0]), .fa_xor1(s_wallace_rca24_fa472_xor1), .fa_or0(s_wallace_rca24_fa472_or0));
  fa fa_s_wallace_rca24_fa473_out(.a(s_wallace_rca24_fa472_or0[0]), .b(s_wallace_rca24_fa351_or0[0]), .cin(s_wallace_rca24_fa304_xor1[0]), .fa_xor1(s_wallace_rca24_fa473_xor1), .fa_or0(s_wallace_rca24_fa473_or0));
  fa fa_s_wallace_rca24_fa474_out(.a(s_wallace_rca24_fa473_or0[0]), .b(s_wallace_rca24_fa329_or0[0]), .cin(s_wallace_rca24_fa278_xor1[0]), .fa_xor1(s_wallace_rca24_fa474_xor1), .fa_or0(s_wallace_rca24_fa474_or0));
  fa fa_s_wallace_rca24_fa475_out(.a(s_wallace_rca24_fa474_or0[0]), .b(s_wallace_rca24_fa305_or0[0]), .cin(s_wallace_rca24_fa250_xor1[0]), .fa_xor1(s_wallace_rca24_fa475_xor1), .fa_or0(s_wallace_rca24_fa475_or0));
  fa fa_s_wallace_rca24_fa476_out(.a(s_wallace_rca24_fa475_or0[0]), .b(s_wallace_rca24_fa279_or0[0]), .cin(s_wallace_rca24_fa220_xor1[0]), .fa_xor1(s_wallace_rca24_fa476_xor1), .fa_or0(s_wallace_rca24_fa476_or0));
  fa fa_s_wallace_rca24_fa477_out(.a(s_wallace_rca24_fa476_or0[0]), .b(s_wallace_rca24_fa251_or0[0]), .cin(s_wallace_rca24_fa188_xor1[0]), .fa_xor1(s_wallace_rca24_fa477_xor1), .fa_or0(s_wallace_rca24_fa477_or0));
  fa fa_s_wallace_rca24_fa478_out(.a(s_wallace_rca24_fa477_or0[0]), .b(s_wallace_rca24_fa221_or0[0]), .cin(s_wallace_rca24_fa154_xor1[0]), .fa_xor1(s_wallace_rca24_fa478_xor1), .fa_or0(s_wallace_rca24_fa478_or0));
  fa fa_s_wallace_rca24_fa479_out(.a(s_wallace_rca24_fa478_or0[0]), .b(s_wallace_rca24_fa189_or0[0]), .cin(s_wallace_rca24_fa118_xor1[0]), .fa_xor1(s_wallace_rca24_fa479_xor1), .fa_or0(s_wallace_rca24_fa479_or0));
  fa fa_s_wallace_rca24_fa480_out(.a(s_wallace_rca24_fa479_or0[0]), .b(s_wallace_rca24_fa155_or0[0]), .cin(s_wallace_rca24_fa80_xor1[0]), .fa_xor1(s_wallace_rca24_fa480_xor1), .fa_or0(s_wallace_rca24_fa480_or0));
  fa fa_s_wallace_rca24_fa481_out(.a(s_wallace_rca24_fa480_or0[0]), .b(s_wallace_rca24_fa119_or0[0]), .cin(s_wallace_rca24_fa40_xor1[0]), .fa_xor1(s_wallace_rca24_fa481_xor1), .fa_or0(s_wallace_rca24_fa481_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_21_23(.a(a[21]), .b(b[23]), .out(s_wallace_rca24_nand_21_23));
  fa fa_s_wallace_rca24_fa482_out(.a(s_wallace_rca24_fa481_or0[0]), .b(s_wallace_rca24_fa81_or0[0]), .cin(s_wallace_rca24_nand_21_23[0]), .fa_xor1(s_wallace_rca24_fa482_xor1), .fa_or0(s_wallace_rca24_fa482_or0));
  nand_gate nand_gate_s_wallace_rca24_nand_23_22(.a(a[23]), .b(b[22]), .out(s_wallace_rca24_nand_23_22));
  fa fa_s_wallace_rca24_fa483_out(.a(s_wallace_rca24_fa482_or0[0]), .b(s_wallace_rca24_fa41_or0[0]), .cin(s_wallace_rca24_nand_23_22[0]), .fa_xor1(s_wallace_rca24_fa483_xor1), .fa_or0(s_wallace_rca24_fa483_or0));
  and_gate and_gate_s_wallace_rca24_and_0_0(.a(a[0]), .b(b[0]), .out(s_wallace_rca24_and_0_0));
  and_gate and_gate_s_wallace_rca24_and_1_0(.a(a[1]), .b(b[0]), .out(s_wallace_rca24_and_1_0));
  and_gate and_gate_s_wallace_rca24_and_0_2(.a(a[0]), .b(b[2]), .out(s_wallace_rca24_and_0_2));
  nand_gate nand_gate_s_wallace_rca24_nand_22_23(.a(a[22]), .b(b[23]), .out(s_wallace_rca24_nand_22_23));
  and_gate and_gate_s_wallace_rca24_and_0_1(.a(a[0]), .b(b[1]), .out(s_wallace_rca24_and_0_1));
  and_gate and_gate_s_wallace_rca24_and_23_23(.a(a[23]), .b(b[23]), .out(s_wallace_rca24_and_23_23));
  assign s_wallace_rca24_u_rca46_a[0] = s_wallace_rca24_and_1_0[0];
  assign s_wallace_rca24_u_rca46_a[1] = s_wallace_rca24_and_0_2[0];
  assign s_wallace_rca24_u_rca46_a[2] = s_wallace_rca24_fa0_xor1[0];
  assign s_wallace_rca24_u_rca46_a[3] = s_wallace_rca24_fa42_xor1[0];
  assign s_wallace_rca24_u_rca46_a[4] = s_wallace_rca24_fa82_xor1[0];
  assign s_wallace_rca24_u_rca46_a[5] = s_wallace_rca24_fa120_xor1[0];
  assign s_wallace_rca24_u_rca46_a[6] = s_wallace_rca24_fa156_xor1[0];
  assign s_wallace_rca24_u_rca46_a[7] = s_wallace_rca24_fa190_xor1[0];
  assign s_wallace_rca24_u_rca46_a[8] = s_wallace_rca24_fa222_xor1[0];
  assign s_wallace_rca24_u_rca46_a[9] = s_wallace_rca24_fa252_xor1[0];
  assign s_wallace_rca24_u_rca46_a[10] = s_wallace_rca24_fa280_xor1[0];
  assign s_wallace_rca24_u_rca46_a[11] = s_wallace_rca24_fa306_xor1[0];
  assign s_wallace_rca24_u_rca46_a[12] = s_wallace_rca24_fa330_xor1[0];
  assign s_wallace_rca24_u_rca46_a[13] = s_wallace_rca24_fa352_xor1[0];
  assign s_wallace_rca24_u_rca46_a[14] = s_wallace_rca24_fa372_xor1[0];
  assign s_wallace_rca24_u_rca46_a[15] = s_wallace_rca24_fa390_xor1[0];
  assign s_wallace_rca24_u_rca46_a[16] = s_wallace_rca24_fa406_xor1[0];
  assign s_wallace_rca24_u_rca46_a[17] = s_wallace_rca24_fa420_xor1[0];
  assign s_wallace_rca24_u_rca46_a[18] = s_wallace_rca24_fa432_xor1[0];
  assign s_wallace_rca24_u_rca46_a[19] = s_wallace_rca24_fa442_xor1[0];
  assign s_wallace_rca24_u_rca46_a[20] = s_wallace_rca24_fa450_xor1[0];
  assign s_wallace_rca24_u_rca46_a[21] = s_wallace_rca24_fa456_xor1[0];
  assign s_wallace_rca24_u_rca46_a[22] = s_wallace_rca24_fa460_xor1[0];
  assign s_wallace_rca24_u_rca46_a[23] = s_wallace_rca24_fa461_xor1[0];
  assign s_wallace_rca24_u_rca46_a[24] = s_wallace_rca24_fa459_xor1[0];
  assign s_wallace_rca24_u_rca46_a[25] = s_wallace_rca24_fa455_xor1[0];
  assign s_wallace_rca24_u_rca46_a[26] = s_wallace_rca24_fa449_xor1[0];
  assign s_wallace_rca24_u_rca46_a[27] = s_wallace_rca24_fa441_xor1[0];
  assign s_wallace_rca24_u_rca46_a[28] = s_wallace_rca24_fa431_xor1[0];
  assign s_wallace_rca24_u_rca46_a[29] = s_wallace_rca24_fa419_xor1[0];
  assign s_wallace_rca24_u_rca46_a[30] = s_wallace_rca24_fa405_xor1[0];
  assign s_wallace_rca24_u_rca46_a[31] = s_wallace_rca24_fa389_xor1[0];
  assign s_wallace_rca24_u_rca46_a[32] = s_wallace_rca24_fa371_xor1[0];
  assign s_wallace_rca24_u_rca46_a[33] = s_wallace_rca24_fa351_xor1[0];
  assign s_wallace_rca24_u_rca46_a[34] = s_wallace_rca24_fa329_xor1[0];
  assign s_wallace_rca24_u_rca46_a[35] = s_wallace_rca24_fa305_xor1[0];
  assign s_wallace_rca24_u_rca46_a[36] = s_wallace_rca24_fa279_xor1[0];
  assign s_wallace_rca24_u_rca46_a[37] = s_wallace_rca24_fa251_xor1[0];
  assign s_wallace_rca24_u_rca46_a[38] = s_wallace_rca24_fa221_xor1[0];
  assign s_wallace_rca24_u_rca46_a[39] = s_wallace_rca24_fa189_xor1[0];
  assign s_wallace_rca24_u_rca46_a[40] = s_wallace_rca24_fa155_xor1[0];
  assign s_wallace_rca24_u_rca46_a[41] = s_wallace_rca24_fa119_xor1[0];
  assign s_wallace_rca24_u_rca46_a[42] = s_wallace_rca24_fa81_xor1[0];
  assign s_wallace_rca24_u_rca46_a[43] = s_wallace_rca24_fa41_xor1[0];
  assign s_wallace_rca24_u_rca46_a[44] = s_wallace_rca24_nand_22_23[0];
  assign s_wallace_rca24_u_rca46_a[45] = s_wallace_rca24_fa483_or0[0];
  assign s_wallace_rca24_u_rca46_b[0] = s_wallace_rca24_and_0_1[0];
  assign s_wallace_rca24_u_rca46_b[1] = s_wallace_rca24_ha0_xor0[0];
  assign s_wallace_rca24_u_rca46_b[2] = s_wallace_rca24_ha1_xor0[0];
  assign s_wallace_rca24_u_rca46_b[3] = s_wallace_rca24_ha2_xor0[0];
  assign s_wallace_rca24_u_rca46_b[4] = s_wallace_rca24_ha3_xor0[0];
  assign s_wallace_rca24_u_rca46_b[5] = s_wallace_rca24_ha4_xor0[0];
  assign s_wallace_rca24_u_rca46_b[6] = s_wallace_rca24_ha5_xor0[0];
  assign s_wallace_rca24_u_rca46_b[7] = s_wallace_rca24_ha6_xor0[0];
  assign s_wallace_rca24_u_rca46_b[8] = s_wallace_rca24_ha7_xor0[0];
  assign s_wallace_rca24_u_rca46_b[9] = s_wallace_rca24_ha8_xor0[0];
  assign s_wallace_rca24_u_rca46_b[10] = s_wallace_rca24_ha9_xor0[0];
  assign s_wallace_rca24_u_rca46_b[11] = s_wallace_rca24_ha10_xor0[0];
  assign s_wallace_rca24_u_rca46_b[12] = s_wallace_rca24_ha11_xor0[0];
  assign s_wallace_rca24_u_rca46_b[13] = s_wallace_rca24_ha12_xor0[0];
  assign s_wallace_rca24_u_rca46_b[14] = s_wallace_rca24_ha13_xor0[0];
  assign s_wallace_rca24_u_rca46_b[15] = s_wallace_rca24_ha14_xor0[0];
  assign s_wallace_rca24_u_rca46_b[16] = s_wallace_rca24_ha15_xor0[0];
  assign s_wallace_rca24_u_rca46_b[17] = s_wallace_rca24_ha16_xor0[0];
  assign s_wallace_rca24_u_rca46_b[18] = s_wallace_rca24_ha17_xor0[0];
  assign s_wallace_rca24_u_rca46_b[19] = s_wallace_rca24_ha18_xor0[0];
  assign s_wallace_rca24_u_rca46_b[20] = s_wallace_rca24_ha19_xor0[0];
  assign s_wallace_rca24_u_rca46_b[21] = s_wallace_rca24_ha20_xor0[0];
  assign s_wallace_rca24_u_rca46_b[22] = s_wallace_rca24_ha21_xor0[0];
  assign s_wallace_rca24_u_rca46_b[23] = s_wallace_rca24_fa462_xor1[0];
  assign s_wallace_rca24_u_rca46_b[24] = s_wallace_rca24_fa463_xor1[0];
  assign s_wallace_rca24_u_rca46_b[25] = s_wallace_rca24_fa464_xor1[0];
  assign s_wallace_rca24_u_rca46_b[26] = s_wallace_rca24_fa465_xor1[0];
  assign s_wallace_rca24_u_rca46_b[27] = s_wallace_rca24_fa466_xor1[0];
  assign s_wallace_rca24_u_rca46_b[28] = s_wallace_rca24_fa467_xor1[0];
  assign s_wallace_rca24_u_rca46_b[29] = s_wallace_rca24_fa468_xor1[0];
  assign s_wallace_rca24_u_rca46_b[30] = s_wallace_rca24_fa469_xor1[0];
  assign s_wallace_rca24_u_rca46_b[31] = s_wallace_rca24_fa470_xor1[0];
  assign s_wallace_rca24_u_rca46_b[32] = s_wallace_rca24_fa471_xor1[0];
  assign s_wallace_rca24_u_rca46_b[33] = s_wallace_rca24_fa472_xor1[0];
  assign s_wallace_rca24_u_rca46_b[34] = s_wallace_rca24_fa473_xor1[0];
  assign s_wallace_rca24_u_rca46_b[35] = s_wallace_rca24_fa474_xor1[0];
  assign s_wallace_rca24_u_rca46_b[36] = s_wallace_rca24_fa475_xor1[0];
  assign s_wallace_rca24_u_rca46_b[37] = s_wallace_rca24_fa476_xor1[0];
  assign s_wallace_rca24_u_rca46_b[38] = s_wallace_rca24_fa477_xor1[0];
  assign s_wallace_rca24_u_rca46_b[39] = s_wallace_rca24_fa478_xor1[0];
  assign s_wallace_rca24_u_rca46_b[40] = s_wallace_rca24_fa479_xor1[0];
  assign s_wallace_rca24_u_rca46_b[41] = s_wallace_rca24_fa480_xor1[0];
  assign s_wallace_rca24_u_rca46_b[42] = s_wallace_rca24_fa481_xor1[0];
  assign s_wallace_rca24_u_rca46_b[43] = s_wallace_rca24_fa482_xor1[0];
  assign s_wallace_rca24_u_rca46_b[44] = s_wallace_rca24_fa483_xor1[0];
  assign s_wallace_rca24_u_rca46_b[45] = s_wallace_rca24_and_23_23[0];
  u_rca46 u_rca46_s_wallace_rca24_u_rca46_out(.a(s_wallace_rca24_u_rca46_a), .b(s_wallace_rca24_u_rca46_b), .u_rca46_out(s_wallace_rca24_u_rca46_out));
  not_gate not_gate_s_wallace_rca24_xor0(.a(s_wallace_rca24_u_rca46_out[46]), .out(s_wallace_rca24_xor0));

  assign s_wallace_rca24_out[0] = s_wallace_rca24_and_0_0[0];
  assign s_wallace_rca24_out[1] = s_wallace_rca24_u_rca46_out[0];
  assign s_wallace_rca24_out[2] = s_wallace_rca24_u_rca46_out[1];
  assign s_wallace_rca24_out[3] = s_wallace_rca24_u_rca46_out[2];
  assign s_wallace_rca24_out[4] = s_wallace_rca24_u_rca46_out[3];
  assign s_wallace_rca24_out[5] = s_wallace_rca24_u_rca46_out[4];
  assign s_wallace_rca24_out[6] = s_wallace_rca24_u_rca46_out[5];
  assign s_wallace_rca24_out[7] = s_wallace_rca24_u_rca46_out[6];
  assign s_wallace_rca24_out[8] = s_wallace_rca24_u_rca46_out[7];
  assign s_wallace_rca24_out[9] = s_wallace_rca24_u_rca46_out[8];
  assign s_wallace_rca24_out[10] = s_wallace_rca24_u_rca46_out[9];
  assign s_wallace_rca24_out[11] = s_wallace_rca24_u_rca46_out[10];
  assign s_wallace_rca24_out[12] = s_wallace_rca24_u_rca46_out[11];
  assign s_wallace_rca24_out[13] = s_wallace_rca24_u_rca46_out[12];
  assign s_wallace_rca24_out[14] = s_wallace_rca24_u_rca46_out[13];
  assign s_wallace_rca24_out[15] = s_wallace_rca24_u_rca46_out[14];
  assign s_wallace_rca24_out[16] = s_wallace_rca24_u_rca46_out[15];
  assign s_wallace_rca24_out[17] = s_wallace_rca24_u_rca46_out[16];
  assign s_wallace_rca24_out[18] = s_wallace_rca24_u_rca46_out[17];
  assign s_wallace_rca24_out[19] = s_wallace_rca24_u_rca46_out[18];
  assign s_wallace_rca24_out[20] = s_wallace_rca24_u_rca46_out[19];
  assign s_wallace_rca24_out[21] = s_wallace_rca24_u_rca46_out[20];
  assign s_wallace_rca24_out[22] = s_wallace_rca24_u_rca46_out[21];
  assign s_wallace_rca24_out[23] = s_wallace_rca24_u_rca46_out[22];
  assign s_wallace_rca24_out[24] = s_wallace_rca24_u_rca46_out[23];
  assign s_wallace_rca24_out[25] = s_wallace_rca24_u_rca46_out[24];
  assign s_wallace_rca24_out[26] = s_wallace_rca24_u_rca46_out[25];
  assign s_wallace_rca24_out[27] = s_wallace_rca24_u_rca46_out[26];
  assign s_wallace_rca24_out[28] = s_wallace_rca24_u_rca46_out[27];
  assign s_wallace_rca24_out[29] = s_wallace_rca24_u_rca46_out[28];
  assign s_wallace_rca24_out[30] = s_wallace_rca24_u_rca46_out[29];
  assign s_wallace_rca24_out[31] = s_wallace_rca24_u_rca46_out[30];
  assign s_wallace_rca24_out[32] = s_wallace_rca24_u_rca46_out[31];
  assign s_wallace_rca24_out[33] = s_wallace_rca24_u_rca46_out[32];
  assign s_wallace_rca24_out[34] = s_wallace_rca24_u_rca46_out[33];
  assign s_wallace_rca24_out[35] = s_wallace_rca24_u_rca46_out[34];
  assign s_wallace_rca24_out[36] = s_wallace_rca24_u_rca46_out[35];
  assign s_wallace_rca24_out[37] = s_wallace_rca24_u_rca46_out[36];
  assign s_wallace_rca24_out[38] = s_wallace_rca24_u_rca46_out[37];
  assign s_wallace_rca24_out[39] = s_wallace_rca24_u_rca46_out[38];
  assign s_wallace_rca24_out[40] = s_wallace_rca24_u_rca46_out[39];
  assign s_wallace_rca24_out[41] = s_wallace_rca24_u_rca46_out[40];
  assign s_wallace_rca24_out[42] = s_wallace_rca24_u_rca46_out[41];
  assign s_wallace_rca24_out[43] = s_wallace_rca24_u_rca46_out[42];
  assign s_wallace_rca24_out[44] = s_wallace_rca24_u_rca46_out[43];
  assign s_wallace_rca24_out[45] = s_wallace_rca24_u_rca46_out[44];
  assign s_wallace_rca24_out[46] = s_wallace_rca24_u_rca46_out[45];
  assign s_wallace_rca24_out[47] = s_wallace_rca24_xor0[0];
endmodule