module u_csamul_pg_rca8(input [7:0] a, input [7:0] b, output [15:0] u_csamul_pg_rca8_out);
  wire u_csamul_pg_rca8_and0_0;
  wire u_csamul_pg_rca8_and1_0;
  wire u_csamul_pg_rca8_and2_0;
  wire u_csamul_pg_rca8_and3_0;
  wire u_csamul_pg_rca8_and4_0;
  wire u_csamul_pg_rca8_and5_0;
  wire u_csamul_pg_rca8_and6_0;
  wire u_csamul_pg_rca8_and7_0;
  wire u_csamul_pg_rca8_and0_1;
  wire u_csamul_pg_rca8_ha0_1_xor0;
  wire u_csamul_pg_rca8_ha0_1_and0;
  wire u_csamul_pg_rca8_and1_1;
  wire u_csamul_pg_rca8_ha1_1_xor0;
  wire u_csamul_pg_rca8_ha1_1_and0;
  wire u_csamul_pg_rca8_and2_1;
  wire u_csamul_pg_rca8_ha2_1_xor0;
  wire u_csamul_pg_rca8_ha2_1_and0;
  wire u_csamul_pg_rca8_and3_1;
  wire u_csamul_pg_rca8_ha3_1_xor0;
  wire u_csamul_pg_rca8_ha3_1_and0;
  wire u_csamul_pg_rca8_and4_1;
  wire u_csamul_pg_rca8_ha4_1_xor0;
  wire u_csamul_pg_rca8_ha4_1_and0;
  wire u_csamul_pg_rca8_and5_1;
  wire u_csamul_pg_rca8_ha5_1_xor0;
  wire u_csamul_pg_rca8_ha5_1_and0;
  wire u_csamul_pg_rca8_and6_1;
  wire u_csamul_pg_rca8_ha6_1_xor0;
  wire u_csamul_pg_rca8_ha6_1_and0;
  wire u_csamul_pg_rca8_and7_1;
  wire u_csamul_pg_rca8_and0_2;
  wire u_csamul_pg_rca8_fa0_2_xor0;
  wire u_csamul_pg_rca8_fa0_2_and0;
  wire u_csamul_pg_rca8_fa0_2_xor1;
  wire u_csamul_pg_rca8_fa0_2_and1;
  wire u_csamul_pg_rca8_fa0_2_or0;
  wire u_csamul_pg_rca8_and1_2;
  wire u_csamul_pg_rca8_fa1_2_xor0;
  wire u_csamul_pg_rca8_fa1_2_and0;
  wire u_csamul_pg_rca8_fa1_2_xor1;
  wire u_csamul_pg_rca8_fa1_2_and1;
  wire u_csamul_pg_rca8_fa1_2_or0;
  wire u_csamul_pg_rca8_and2_2;
  wire u_csamul_pg_rca8_fa2_2_xor0;
  wire u_csamul_pg_rca8_fa2_2_and0;
  wire u_csamul_pg_rca8_fa2_2_xor1;
  wire u_csamul_pg_rca8_fa2_2_and1;
  wire u_csamul_pg_rca8_fa2_2_or0;
  wire u_csamul_pg_rca8_and3_2;
  wire u_csamul_pg_rca8_fa3_2_xor0;
  wire u_csamul_pg_rca8_fa3_2_and0;
  wire u_csamul_pg_rca8_fa3_2_xor1;
  wire u_csamul_pg_rca8_fa3_2_and1;
  wire u_csamul_pg_rca8_fa3_2_or0;
  wire u_csamul_pg_rca8_and4_2;
  wire u_csamul_pg_rca8_fa4_2_xor0;
  wire u_csamul_pg_rca8_fa4_2_and0;
  wire u_csamul_pg_rca8_fa4_2_xor1;
  wire u_csamul_pg_rca8_fa4_2_and1;
  wire u_csamul_pg_rca8_fa4_2_or0;
  wire u_csamul_pg_rca8_and5_2;
  wire u_csamul_pg_rca8_fa5_2_xor0;
  wire u_csamul_pg_rca8_fa5_2_and0;
  wire u_csamul_pg_rca8_fa5_2_xor1;
  wire u_csamul_pg_rca8_fa5_2_and1;
  wire u_csamul_pg_rca8_fa5_2_or0;
  wire u_csamul_pg_rca8_and6_2;
  wire u_csamul_pg_rca8_fa6_2_xor0;
  wire u_csamul_pg_rca8_fa6_2_and0;
  wire u_csamul_pg_rca8_fa6_2_xor1;
  wire u_csamul_pg_rca8_fa6_2_and1;
  wire u_csamul_pg_rca8_fa6_2_or0;
  wire u_csamul_pg_rca8_and7_2;
  wire u_csamul_pg_rca8_and0_3;
  wire u_csamul_pg_rca8_fa0_3_xor0;
  wire u_csamul_pg_rca8_fa0_3_and0;
  wire u_csamul_pg_rca8_fa0_3_xor1;
  wire u_csamul_pg_rca8_fa0_3_and1;
  wire u_csamul_pg_rca8_fa0_3_or0;
  wire u_csamul_pg_rca8_and1_3;
  wire u_csamul_pg_rca8_fa1_3_xor0;
  wire u_csamul_pg_rca8_fa1_3_and0;
  wire u_csamul_pg_rca8_fa1_3_xor1;
  wire u_csamul_pg_rca8_fa1_3_and1;
  wire u_csamul_pg_rca8_fa1_3_or0;
  wire u_csamul_pg_rca8_and2_3;
  wire u_csamul_pg_rca8_fa2_3_xor0;
  wire u_csamul_pg_rca8_fa2_3_and0;
  wire u_csamul_pg_rca8_fa2_3_xor1;
  wire u_csamul_pg_rca8_fa2_3_and1;
  wire u_csamul_pg_rca8_fa2_3_or0;
  wire u_csamul_pg_rca8_and3_3;
  wire u_csamul_pg_rca8_fa3_3_xor0;
  wire u_csamul_pg_rca8_fa3_3_and0;
  wire u_csamul_pg_rca8_fa3_3_xor1;
  wire u_csamul_pg_rca8_fa3_3_and1;
  wire u_csamul_pg_rca8_fa3_3_or0;
  wire u_csamul_pg_rca8_and4_3;
  wire u_csamul_pg_rca8_fa4_3_xor0;
  wire u_csamul_pg_rca8_fa4_3_and0;
  wire u_csamul_pg_rca8_fa4_3_xor1;
  wire u_csamul_pg_rca8_fa4_3_and1;
  wire u_csamul_pg_rca8_fa4_3_or0;
  wire u_csamul_pg_rca8_and5_3;
  wire u_csamul_pg_rca8_fa5_3_xor0;
  wire u_csamul_pg_rca8_fa5_3_and0;
  wire u_csamul_pg_rca8_fa5_3_xor1;
  wire u_csamul_pg_rca8_fa5_3_and1;
  wire u_csamul_pg_rca8_fa5_3_or0;
  wire u_csamul_pg_rca8_and6_3;
  wire u_csamul_pg_rca8_fa6_3_xor0;
  wire u_csamul_pg_rca8_fa6_3_and0;
  wire u_csamul_pg_rca8_fa6_3_xor1;
  wire u_csamul_pg_rca8_fa6_3_and1;
  wire u_csamul_pg_rca8_fa6_3_or0;
  wire u_csamul_pg_rca8_and7_3;
  wire u_csamul_pg_rca8_and0_4;
  wire u_csamul_pg_rca8_fa0_4_xor0;
  wire u_csamul_pg_rca8_fa0_4_and0;
  wire u_csamul_pg_rca8_fa0_4_xor1;
  wire u_csamul_pg_rca8_fa0_4_and1;
  wire u_csamul_pg_rca8_fa0_4_or0;
  wire u_csamul_pg_rca8_and1_4;
  wire u_csamul_pg_rca8_fa1_4_xor0;
  wire u_csamul_pg_rca8_fa1_4_and0;
  wire u_csamul_pg_rca8_fa1_4_xor1;
  wire u_csamul_pg_rca8_fa1_4_and1;
  wire u_csamul_pg_rca8_fa1_4_or0;
  wire u_csamul_pg_rca8_and2_4;
  wire u_csamul_pg_rca8_fa2_4_xor0;
  wire u_csamul_pg_rca8_fa2_4_and0;
  wire u_csamul_pg_rca8_fa2_4_xor1;
  wire u_csamul_pg_rca8_fa2_4_and1;
  wire u_csamul_pg_rca8_fa2_4_or0;
  wire u_csamul_pg_rca8_and3_4;
  wire u_csamul_pg_rca8_fa3_4_xor0;
  wire u_csamul_pg_rca8_fa3_4_and0;
  wire u_csamul_pg_rca8_fa3_4_xor1;
  wire u_csamul_pg_rca8_fa3_4_and1;
  wire u_csamul_pg_rca8_fa3_4_or0;
  wire u_csamul_pg_rca8_and4_4;
  wire u_csamul_pg_rca8_fa4_4_xor0;
  wire u_csamul_pg_rca8_fa4_4_and0;
  wire u_csamul_pg_rca8_fa4_4_xor1;
  wire u_csamul_pg_rca8_fa4_4_and1;
  wire u_csamul_pg_rca8_fa4_4_or0;
  wire u_csamul_pg_rca8_and5_4;
  wire u_csamul_pg_rca8_fa5_4_xor0;
  wire u_csamul_pg_rca8_fa5_4_and0;
  wire u_csamul_pg_rca8_fa5_4_xor1;
  wire u_csamul_pg_rca8_fa5_4_and1;
  wire u_csamul_pg_rca8_fa5_4_or0;
  wire u_csamul_pg_rca8_and6_4;
  wire u_csamul_pg_rca8_fa6_4_xor0;
  wire u_csamul_pg_rca8_fa6_4_and0;
  wire u_csamul_pg_rca8_fa6_4_xor1;
  wire u_csamul_pg_rca8_fa6_4_and1;
  wire u_csamul_pg_rca8_fa6_4_or0;
  wire u_csamul_pg_rca8_and7_4;
  wire u_csamul_pg_rca8_and0_5;
  wire u_csamul_pg_rca8_fa0_5_xor0;
  wire u_csamul_pg_rca8_fa0_5_and0;
  wire u_csamul_pg_rca8_fa0_5_xor1;
  wire u_csamul_pg_rca8_fa0_5_and1;
  wire u_csamul_pg_rca8_fa0_5_or0;
  wire u_csamul_pg_rca8_and1_5;
  wire u_csamul_pg_rca8_fa1_5_xor0;
  wire u_csamul_pg_rca8_fa1_5_and0;
  wire u_csamul_pg_rca8_fa1_5_xor1;
  wire u_csamul_pg_rca8_fa1_5_and1;
  wire u_csamul_pg_rca8_fa1_5_or0;
  wire u_csamul_pg_rca8_and2_5;
  wire u_csamul_pg_rca8_fa2_5_xor0;
  wire u_csamul_pg_rca8_fa2_5_and0;
  wire u_csamul_pg_rca8_fa2_5_xor1;
  wire u_csamul_pg_rca8_fa2_5_and1;
  wire u_csamul_pg_rca8_fa2_5_or0;
  wire u_csamul_pg_rca8_and3_5;
  wire u_csamul_pg_rca8_fa3_5_xor0;
  wire u_csamul_pg_rca8_fa3_5_and0;
  wire u_csamul_pg_rca8_fa3_5_xor1;
  wire u_csamul_pg_rca8_fa3_5_and1;
  wire u_csamul_pg_rca8_fa3_5_or0;
  wire u_csamul_pg_rca8_and4_5;
  wire u_csamul_pg_rca8_fa4_5_xor0;
  wire u_csamul_pg_rca8_fa4_5_and0;
  wire u_csamul_pg_rca8_fa4_5_xor1;
  wire u_csamul_pg_rca8_fa4_5_and1;
  wire u_csamul_pg_rca8_fa4_5_or0;
  wire u_csamul_pg_rca8_and5_5;
  wire u_csamul_pg_rca8_fa5_5_xor0;
  wire u_csamul_pg_rca8_fa5_5_and0;
  wire u_csamul_pg_rca8_fa5_5_xor1;
  wire u_csamul_pg_rca8_fa5_5_and1;
  wire u_csamul_pg_rca8_fa5_5_or0;
  wire u_csamul_pg_rca8_and6_5;
  wire u_csamul_pg_rca8_fa6_5_xor0;
  wire u_csamul_pg_rca8_fa6_5_and0;
  wire u_csamul_pg_rca8_fa6_5_xor1;
  wire u_csamul_pg_rca8_fa6_5_and1;
  wire u_csamul_pg_rca8_fa6_5_or0;
  wire u_csamul_pg_rca8_and7_5;
  wire u_csamul_pg_rca8_and0_6;
  wire u_csamul_pg_rca8_fa0_6_xor0;
  wire u_csamul_pg_rca8_fa0_6_and0;
  wire u_csamul_pg_rca8_fa0_6_xor1;
  wire u_csamul_pg_rca8_fa0_6_and1;
  wire u_csamul_pg_rca8_fa0_6_or0;
  wire u_csamul_pg_rca8_and1_6;
  wire u_csamul_pg_rca8_fa1_6_xor0;
  wire u_csamul_pg_rca8_fa1_6_and0;
  wire u_csamul_pg_rca8_fa1_6_xor1;
  wire u_csamul_pg_rca8_fa1_6_and1;
  wire u_csamul_pg_rca8_fa1_6_or0;
  wire u_csamul_pg_rca8_and2_6;
  wire u_csamul_pg_rca8_fa2_6_xor0;
  wire u_csamul_pg_rca8_fa2_6_and0;
  wire u_csamul_pg_rca8_fa2_6_xor1;
  wire u_csamul_pg_rca8_fa2_6_and1;
  wire u_csamul_pg_rca8_fa2_6_or0;
  wire u_csamul_pg_rca8_and3_6;
  wire u_csamul_pg_rca8_fa3_6_xor0;
  wire u_csamul_pg_rca8_fa3_6_and0;
  wire u_csamul_pg_rca8_fa3_6_xor1;
  wire u_csamul_pg_rca8_fa3_6_and1;
  wire u_csamul_pg_rca8_fa3_6_or0;
  wire u_csamul_pg_rca8_and4_6;
  wire u_csamul_pg_rca8_fa4_6_xor0;
  wire u_csamul_pg_rca8_fa4_6_and0;
  wire u_csamul_pg_rca8_fa4_6_xor1;
  wire u_csamul_pg_rca8_fa4_6_and1;
  wire u_csamul_pg_rca8_fa4_6_or0;
  wire u_csamul_pg_rca8_and5_6;
  wire u_csamul_pg_rca8_fa5_6_xor0;
  wire u_csamul_pg_rca8_fa5_6_and0;
  wire u_csamul_pg_rca8_fa5_6_xor1;
  wire u_csamul_pg_rca8_fa5_6_and1;
  wire u_csamul_pg_rca8_fa5_6_or0;
  wire u_csamul_pg_rca8_and6_6;
  wire u_csamul_pg_rca8_fa6_6_xor0;
  wire u_csamul_pg_rca8_fa6_6_and0;
  wire u_csamul_pg_rca8_fa6_6_xor1;
  wire u_csamul_pg_rca8_fa6_6_and1;
  wire u_csamul_pg_rca8_fa6_6_or0;
  wire u_csamul_pg_rca8_and7_6;
  wire u_csamul_pg_rca8_and0_7;
  wire u_csamul_pg_rca8_fa0_7_xor0;
  wire u_csamul_pg_rca8_fa0_7_and0;
  wire u_csamul_pg_rca8_fa0_7_xor1;
  wire u_csamul_pg_rca8_fa0_7_and1;
  wire u_csamul_pg_rca8_fa0_7_or0;
  wire u_csamul_pg_rca8_and1_7;
  wire u_csamul_pg_rca8_fa1_7_xor0;
  wire u_csamul_pg_rca8_fa1_7_and0;
  wire u_csamul_pg_rca8_fa1_7_xor1;
  wire u_csamul_pg_rca8_fa1_7_and1;
  wire u_csamul_pg_rca8_fa1_7_or0;
  wire u_csamul_pg_rca8_and2_7;
  wire u_csamul_pg_rca8_fa2_7_xor0;
  wire u_csamul_pg_rca8_fa2_7_and0;
  wire u_csamul_pg_rca8_fa2_7_xor1;
  wire u_csamul_pg_rca8_fa2_7_and1;
  wire u_csamul_pg_rca8_fa2_7_or0;
  wire u_csamul_pg_rca8_and3_7;
  wire u_csamul_pg_rca8_fa3_7_xor0;
  wire u_csamul_pg_rca8_fa3_7_and0;
  wire u_csamul_pg_rca8_fa3_7_xor1;
  wire u_csamul_pg_rca8_fa3_7_and1;
  wire u_csamul_pg_rca8_fa3_7_or0;
  wire u_csamul_pg_rca8_and4_7;
  wire u_csamul_pg_rca8_fa4_7_xor0;
  wire u_csamul_pg_rca8_fa4_7_and0;
  wire u_csamul_pg_rca8_fa4_7_xor1;
  wire u_csamul_pg_rca8_fa4_7_and1;
  wire u_csamul_pg_rca8_fa4_7_or0;
  wire u_csamul_pg_rca8_and5_7;
  wire u_csamul_pg_rca8_fa5_7_xor0;
  wire u_csamul_pg_rca8_fa5_7_and0;
  wire u_csamul_pg_rca8_fa5_7_xor1;
  wire u_csamul_pg_rca8_fa5_7_and1;
  wire u_csamul_pg_rca8_fa5_7_or0;
  wire u_csamul_pg_rca8_and6_7;
  wire u_csamul_pg_rca8_fa6_7_xor0;
  wire u_csamul_pg_rca8_fa6_7_and0;
  wire u_csamul_pg_rca8_fa6_7_xor1;
  wire u_csamul_pg_rca8_fa6_7_and1;
  wire u_csamul_pg_rca8_fa6_7_or0;
  wire u_csamul_pg_rca8_and7_7;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa0_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa0_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa1_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor1;
  wire u_csamul_pg_rca8_u_pg_rca8_and1;
  wire u_csamul_pg_rca8_u_pg_rca8_or1;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa2_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor1;
  wire u_csamul_pg_rca8_u_pg_rca8_and2;
  wire u_csamul_pg_rca8_u_pg_rca8_or2;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa3_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor1;
  wire u_csamul_pg_rca8_u_pg_rca8_and3;
  wire u_csamul_pg_rca8_u_pg_rca8_or3;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa4_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor1;
  wire u_csamul_pg_rca8_u_pg_rca8_and4;
  wire u_csamul_pg_rca8_u_pg_rca8_or4;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa5_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor1;
  wire u_csamul_pg_rca8_u_pg_rca8_and5;
  wire u_csamul_pg_rca8_u_pg_rca8_or5;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa6_and0;
  wire u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor1;
  wire u_csamul_pg_rca8_u_pg_rca8_and6;
  wire u_csamul_pg_rca8_u_pg_rca8_or6;

  assign u_csamul_pg_rca8_and0_0 = a[0] & b[0];
  assign u_csamul_pg_rca8_and1_0 = a[1] & b[0];
  assign u_csamul_pg_rca8_and2_0 = a[2] & b[0];
  assign u_csamul_pg_rca8_and3_0 = a[3] & b[0];
  assign u_csamul_pg_rca8_and4_0 = a[4] & b[0];
  assign u_csamul_pg_rca8_and5_0 = a[5] & b[0];
  assign u_csamul_pg_rca8_and6_0 = a[6] & b[0];
  assign u_csamul_pg_rca8_and7_0 = a[7] & b[0];
  assign u_csamul_pg_rca8_and0_1 = a[0] & b[1];
  assign u_csamul_pg_rca8_ha0_1_xor0 = u_csamul_pg_rca8_and0_1 ^ u_csamul_pg_rca8_and1_0;
  assign u_csamul_pg_rca8_ha0_1_and0 = u_csamul_pg_rca8_and0_1 & u_csamul_pg_rca8_and1_0;
  assign u_csamul_pg_rca8_and1_1 = a[1] & b[1];
  assign u_csamul_pg_rca8_ha1_1_xor0 = u_csamul_pg_rca8_and1_1 ^ u_csamul_pg_rca8_and2_0;
  assign u_csamul_pg_rca8_ha1_1_and0 = u_csamul_pg_rca8_and1_1 & u_csamul_pg_rca8_and2_0;
  assign u_csamul_pg_rca8_and2_1 = a[2] & b[1];
  assign u_csamul_pg_rca8_ha2_1_xor0 = u_csamul_pg_rca8_and2_1 ^ u_csamul_pg_rca8_and3_0;
  assign u_csamul_pg_rca8_ha2_1_and0 = u_csamul_pg_rca8_and2_1 & u_csamul_pg_rca8_and3_0;
  assign u_csamul_pg_rca8_and3_1 = a[3] & b[1];
  assign u_csamul_pg_rca8_ha3_1_xor0 = u_csamul_pg_rca8_and3_1 ^ u_csamul_pg_rca8_and4_0;
  assign u_csamul_pg_rca8_ha3_1_and0 = u_csamul_pg_rca8_and3_1 & u_csamul_pg_rca8_and4_0;
  assign u_csamul_pg_rca8_and4_1 = a[4] & b[1];
  assign u_csamul_pg_rca8_ha4_1_xor0 = u_csamul_pg_rca8_and4_1 ^ u_csamul_pg_rca8_and5_0;
  assign u_csamul_pg_rca8_ha4_1_and0 = u_csamul_pg_rca8_and4_1 & u_csamul_pg_rca8_and5_0;
  assign u_csamul_pg_rca8_and5_1 = a[5] & b[1];
  assign u_csamul_pg_rca8_ha5_1_xor0 = u_csamul_pg_rca8_and5_1 ^ u_csamul_pg_rca8_and6_0;
  assign u_csamul_pg_rca8_ha5_1_and0 = u_csamul_pg_rca8_and5_1 & u_csamul_pg_rca8_and6_0;
  assign u_csamul_pg_rca8_and6_1 = a[6] & b[1];
  assign u_csamul_pg_rca8_ha6_1_xor0 = u_csamul_pg_rca8_and6_1 ^ u_csamul_pg_rca8_and7_0;
  assign u_csamul_pg_rca8_ha6_1_and0 = u_csamul_pg_rca8_and6_1 & u_csamul_pg_rca8_and7_0;
  assign u_csamul_pg_rca8_and7_1 = a[7] & b[1];
  assign u_csamul_pg_rca8_and0_2 = a[0] & b[2];
  assign u_csamul_pg_rca8_fa0_2_xor0 = u_csamul_pg_rca8_and0_2 ^ u_csamul_pg_rca8_ha1_1_xor0;
  assign u_csamul_pg_rca8_fa0_2_and0 = u_csamul_pg_rca8_and0_2 & u_csamul_pg_rca8_ha1_1_xor0;
  assign u_csamul_pg_rca8_fa0_2_xor1 = u_csamul_pg_rca8_fa0_2_xor0 ^ u_csamul_pg_rca8_ha0_1_and0;
  assign u_csamul_pg_rca8_fa0_2_and1 = u_csamul_pg_rca8_fa0_2_xor0 & u_csamul_pg_rca8_ha0_1_and0;
  assign u_csamul_pg_rca8_fa0_2_or0 = u_csamul_pg_rca8_fa0_2_and0 | u_csamul_pg_rca8_fa0_2_and1;
  assign u_csamul_pg_rca8_and1_2 = a[1] & b[2];
  assign u_csamul_pg_rca8_fa1_2_xor0 = u_csamul_pg_rca8_and1_2 ^ u_csamul_pg_rca8_ha2_1_xor0;
  assign u_csamul_pg_rca8_fa1_2_and0 = u_csamul_pg_rca8_and1_2 & u_csamul_pg_rca8_ha2_1_xor0;
  assign u_csamul_pg_rca8_fa1_2_xor1 = u_csamul_pg_rca8_fa1_2_xor0 ^ u_csamul_pg_rca8_ha1_1_and0;
  assign u_csamul_pg_rca8_fa1_2_and1 = u_csamul_pg_rca8_fa1_2_xor0 & u_csamul_pg_rca8_ha1_1_and0;
  assign u_csamul_pg_rca8_fa1_2_or0 = u_csamul_pg_rca8_fa1_2_and0 | u_csamul_pg_rca8_fa1_2_and1;
  assign u_csamul_pg_rca8_and2_2 = a[2] & b[2];
  assign u_csamul_pg_rca8_fa2_2_xor0 = u_csamul_pg_rca8_and2_2 ^ u_csamul_pg_rca8_ha3_1_xor0;
  assign u_csamul_pg_rca8_fa2_2_and0 = u_csamul_pg_rca8_and2_2 & u_csamul_pg_rca8_ha3_1_xor0;
  assign u_csamul_pg_rca8_fa2_2_xor1 = u_csamul_pg_rca8_fa2_2_xor0 ^ u_csamul_pg_rca8_ha2_1_and0;
  assign u_csamul_pg_rca8_fa2_2_and1 = u_csamul_pg_rca8_fa2_2_xor0 & u_csamul_pg_rca8_ha2_1_and0;
  assign u_csamul_pg_rca8_fa2_2_or0 = u_csamul_pg_rca8_fa2_2_and0 | u_csamul_pg_rca8_fa2_2_and1;
  assign u_csamul_pg_rca8_and3_2 = a[3] & b[2];
  assign u_csamul_pg_rca8_fa3_2_xor0 = u_csamul_pg_rca8_and3_2 ^ u_csamul_pg_rca8_ha4_1_xor0;
  assign u_csamul_pg_rca8_fa3_2_and0 = u_csamul_pg_rca8_and3_2 & u_csamul_pg_rca8_ha4_1_xor0;
  assign u_csamul_pg_rca8_fa3_2_xor1 = u_csamul_pg_rca8_fa3_2_xor0 ^ u_csamul_pg_rca8_ha3_1_and0;
  assign u_csamul_pg_rca8_fa3_2_and1 = u_csamul_pg_rca8_fa3_2_xor0 & u_csamul_pg_rca8_ha3_1_and0;
  assign u_csamul_pg_rca8_fa3_2_or0 = u_csamul_pg_rca8_fa3_2_and0 | u_csamul_pg_rca8_fa3_2_and1;
  assign u_csamul_pg_rca8_and4_2 = a[4] & b[2];
  assign u_csamul_pg_rca8_fa4_2_xor0 = u_csamul_pg_rca8_and4_2 ^ u_csamul_pg_rca8_ha5_1_xor0;
  assign u_csamul_pg_rca8_fa4_2_and0 = u_csamul_pg_rca8_and4_2 & u_csamul_pg_rca8_ha5_1_xor0;
  assign u_csamul_pg_rca8_fa4_2_xor1 = u_csamul_pg_rca8_fa4_2_xor0 ^ u_csamul_pg_rca8_ha4_1_and0;
  assign u_csamul_pg_rca8_fa4_2_and1 = u_csamul_pg_rca8_fa4_2_xor0 & u_csamul_pg_rca8_ha4_1_and0;
  assign u_csamul_pg_rca8_fa4_2_or0 = u_csamul_pg_rca8_fa4_2_and0 | u_csamul_pg_rca8_fa4_2_and1;
  assign u_csamul_pg_rca8_and5_2 = a[5] & b[2];
  assign u_csamul_pg_rca8_fa5_2_xor0 = u_csamul_pg_rca8_and5_2 ^ u_csamul_pg_rca8_ha6_1_xor0;
  assign u_csamul_pg_rca8_fa5_2_and0 = u_csamul_pg_rca8_and5_2 & u_csamul_pg_rca8_ha6_1_xor0;
  assign u_csamul_pg_rca8_fa5_2_xor1 = u_csamul_pg_rca8_fa5_2_xor0 ^ u_csamul_pg_rca8_ha5_1_and0;
  assign u_csamul_pg_rca8_fa5_2_and1 = u_csamul_pg_rca8_fa5_2_xor0 & u_csamul_pg_rca8_ha5_1_and0;
  assign u_csamul_pg_rca8_fa5_2_or0 = u_csamul_pg_rca8_fa5_2_and0 | u_csamul_pg_rca8_fa5_2_and1;
  assign u_csamul_pg_rca8_and6_2 = a[6] & b[2];
  assign u_csamul_pg_rca8_fa6_2_xor0 = u_csamul_pg_rca8_and6_2 ^ u_csamul_pg_rca8_and7_1;
  assign u_csamul_pg_rca8_fa6_2_and0 = u_csamul_pg_rca8_and6_2 & u_csamul_pg_rca8_and7_1;
  assign u_csamul_pg_rca8_fa6_2_xor1 = u_csamul_pg_rca8_fa6_2_xor0 ^ u_csamul_pg_rca8_ha6_1_and0;
  assign u_csamul_pg_rca8_fa6_2_and1 = u_csamul_pg_rca8_fa6_2_xor0 & u_csamul_pg_rca8_ha6_1_and0;
  assign u_csamul_pg_rca8_fa6_2_or0 = u_csamul_pg_rca8_fa6_2_and0 | u_csamul_pg_rca8_fa6_2_and1;
  assign u_csamul_pg_rca8_and7_2 = a[7] & b[2];
  assign u_csamul_pg_rca8_and0_3 = a[0] & b[3];
  assign u_csamul_pg_rca8_fa0_3_xor0 = u_csamul_pg_rca8_and0_3 ^ u_csamul_pg_rca8_fa1_2_xor1;
  assign u_csamul_pg_rca8_fa0_3_and0 = u_csamul_pg_rca8_and0_3 & u_csamul_pg_rca8_fa1_2_xor1;
  assign u_csamul_pg_rca8_fa0_3_xor1 = u_csamul_pg_rca8_fa0_3_xor0 ^ u_csamul_pg_rca8_fa0_2_or0;
  assign u_csamul_pg_rca8_fa0_3_and1 = u_csamul_pg_rca8_fa0_3_xor0 & u_csamul_pg_rca8_fa0_2_or0;
  assign u_csamul_pg_rca8_fa0_3_or0 = u_csamul_pg_rca8_fa0_3_and0 | u_csamul_pg_rca8_fa0_3_and1;
  assign u_csamul_pg_rca8_and1_3 = a[1] & b[3];
  assign u_csamul_pg_rca8_fa1_3_xor0 = u_csamul_pg_rca8_and1_3 ^ u_csamul_pg_rca8_fa2_2_xor1;
  assign u_csamul_pg_rca8_fa1_3_and0 = u_csamul_pg_rca8_and1_3 & u_csamul_pg_rca8_fa2_2_xor1;
  assign u_csamul_pg_rca8_fa1_3_xor1 = u_csamul_pg_rca8_fa1_3_xor0 ^ u_csamul_pg_rca8_fa1_2_or0;
  assign u_csamul_pg_rca8_fa1_3_and1 = u_csamul_pg_rca8_fa1_3_xor0 & u_csamul_pg_rca8_fa1_2_or0;
  assign u_csamul_pg_rca8_fa1_3_or0 = u_csamul_pg_rca8_fa1_3_and0 | u_csamul_pg_rca8_fa1_3_and1;
  assign u_csamul_pg_rca8_and2_3 = a[2] & b[3];
  assign u_csamul_pg_rca8_fa2_3_xor0 = u_csamul_pg_rca8_and2_3 ^ u_csamul_pg_rca8_fa3_2_xor1;
  assign u_csamul_pg_rca8_fa2_3_and0 = u_csamul_pg_rca8_and2_3 & u_csamul_pg_rca8_fa3_2_xor1;
  assign u_csamul_pg_rca8_fa2_3_xor1 = u_csamul_pg_rca8_fa2_3_xor0 ^ u_csamul_pg_rca8_fa2_2_or0;
  assign u_csamul_pg_rca8_fa2_3_and1 = u_csamul_pg_rca8_fa2_3_xor0 & u_csamul_pg_rca8_fa2_2_or0;
  assign u_csamul_pg_rca8_fa2_3_or0 = u_csamul_pg_rca8_fa2_3_and0 | u_csamul_pg_rca8_fa2_3_and1;
  assign u_csamul_pg_rca8_and3_3 = a[3] & b[3];
  assign u_csamul_pg_rca8_fa3_3_xor0 = u_csamul_pg_rca8_and3_3 ^ u_csamul_pg_rca8_fa4_2_xor1;
  assign u_csamul_pg_rca8_fa3_3_and0 = u_csamul_pg_rca8_and3_3 & u_csamul_pg_rca8_fa4_2_xor1;
  assign u_csamul_pg_rca8_fa3_3_xor1 = u_csamul_pg_rca8_fa3_3_xor0 ^ u_csamul_pg_rca8_fa3_2_or0;
  assign u_csamul_pg_rca8_fa3_3_and1 = u_csamul_pg_rca8_fa3_3_xor0 & u_csamul_pg_rca8_fa3_2_or0;
  assign u_csamul_pg_rca8_fa3_3_or0 = u_csamul_pg_rca8_fa3_3_and0 | u_csamul_pg_rca8_fa3_3_and1;
  assign u_csamul_pg_rca8_and4_3 = a[4] & b[3];
  assign u_csamul_pg_rca8_fa4_3_xor0 = u_csamul_pg_rca8_and4_3 ^ u_csamul_pg_rca8_fa5_2_xor1;
  assign u_csamul_pg_rca8_fa4_3_and0 = u_csamul_pg_rca8_and4_3 & u_csamul_pg_rca8_fa5_2_xor1;
  assign u_csamul_pg_rca8_fa4_3_xor1 = u_csamul_pg_rca8_fa4_3_xor0 ^ u_csamul_pg_rca8_fa4_2_or0;
  assign u_csamul_pg_rca8_fa4_3_and1 = u_csamul_pg_rca8_fa4_3_xor0 & u_csamul_pg_rca8_fa4_2_or0;
  assign u_csamul_pg_rca8_fa4_3_or0 = u_csamul_pg_rca8_fa4_3_and0 | u_csamul_pg_rca8_fa4_3_and1;
  assign u_csamul_pg_rca8_and5_3 = a[5] & b[3];
  assign u_csamul_pg_rca8_fa5_3_xor0 = u_csamul_pg_rca8_and5_3 ^ u_csamul_pg_rca8_fa6_2_xor1;
  assign u_csamul_pg_rca8_fa5_3_and0 = u_csamul_pg_rca8_and5_3 & u_csamul_pg_rca8_fa6_2_xor1;
  assign u_csamul_pg_rca8_fa5_3_xor1 = u_csamul_pg_rca8_fa5_3_xor0 ^ u_csamul_pg_rca8_fa5_2_or0;
  assign u_csamul_pg_rca8_fa5_3_and1 = u_csamul_pg_rca8_fa5_3_xor0 & u_csamul_pg_rca8_fa5_2_or0;
  assign u_csamul_pg_rca8_fa5_3_or0 = u_csamul_pg_rca8_fa5_3_and0 | u_csamul_pg_rca8_fa5_3_and1;
  assign u_csamul_pg_rca8_and6_3 = a[6] & b[3];
  assign u_csamul_pg_rca8_fa6_3_xor0 = u_csamul_pg_rca8_and6_3 ^ u_csamul_pg_rca8_and7_2;
  assign u_csamul_pg_rca8_fa6_3_and0 = u_csamul_pg_rca8_and6_3 & u_csamul_pg_rca8_and7_2;
  assign u_csamul_pg_rca8_fa6_3_xor1 = u_csamul_pg_rca8_fa6_3_xor0 ^ u_csamul_pg_rca8_fa6_2_or0;
  assign u_csamul_pg_rca8_fa6_3_and1 = u_csamul_pg_rca8_fa6_3_xor0 & u_csamul_pg_rca8_fa6_2_or0;
  assign u_csamul_pg_rca8_fa6_3_or0 = u_csamul_pg_rca8_fa6_3_and0 | u_csamul_pg_rca8_fa6_3_and1;
  assign u_csamul_pg_rca8_and7_3 = a[7] & b[3];
  assign u_csamul_pg_rca8_and0_4 = a[0] & b[4];
  assign u_csamul_pg_rca8_fa0_4_xor0 = u_csamul_pg_rca8_and0_4 ^ u_csamul_pg_rca8_fa1_3_xor1;
  assign u_csamul_pg_rca8_fa0_4_and0 = u_csamul_pg_rca8_and0_4 & u_csamul_pg_rca8_fa1_3_xor1;
  assign u_csamul_pg_rca8_fa0_4_xor1 = u_csamul_pg_rca8_fa0_4_xor0 ^ u_csamul_pg_rca8_fa0_3_or0;
  assign u_csamul_pg_rca8_fa0_4_and1 = u_csamul_pg_rca8_fa0_4_xor0 & u_csamul_pg_rca8_fa0_3_or0;
  assign u_csamul_pg_rca8_fa0_4_or0 = u_csamul_pg_rca8_fa0_4_and0 | u_csamul_pg_rca8_fa0_4_and1;
  assign u_csamul_pg_rca8_and1_4 = a[1] & b[4];
  assign u_csamul_pg_rca8_fa1_4_xor0 = u_csamul_pg_rca8_and1_4 ^ u_csamul_pg_rca8_fa2_3_xor1;
  assign u_csamul_pg_rca8_fa1_4_and0 = u_csamul_pg_rca8_and1_4 & u_csamul_pg_rca8_fa2_3_xor1;
  assign u_csamul_pg_rca8_fa1_4_xor1 = u_csamul_pg_rca8_fa1_4_xor0 ^ u_csamul_pg_rca8_fa1_3_or0;
  assign u_csamul_pg_rca8_fa1_4_and1 = u_csamul_pg_rca8_fa1_4_xor0 & u_csamul_pg_rca8_fa1_3_or0;
  assign u_csamul_pg_rca8_fa1_4_or0 = u_csamul_pg_rca8_fa1_4_and0 | u_csamul_pg_rca8_fa1_4_and1;
  assign u_csamul_pg_rca8_and2_4 = a[2] & b[4];
  assign u_csamul_pg_rca8_fa2_4_xor0 = u_csamul_pg_rca8_and2_4 ^ u_csamul_pg_rca8_fa3_3_xor1;
  assign u_csamul_pg_rca8_fa2_4_and0 = u_csamul_pg_rca8_and2_4 & u_csamul_pg_rca8_fa3_3_xor1;
  assign u_csamul_pg_rca8_fa2_4_xor1 = u_csamul_pg_rca8_fa2_4_xor0 ^ u_csamul_pg_rca8_fa2_3_or0;
  assign u_csamul_pg_rca8_fa2_4_and1 = u_csamul_pg_rca8_fa2_4_xor0 & u_csamul_pg_rca8_fa2_3_or0;
  assign u_csamul_pg_rca8_fa2_4_or0 = u_csamul_pg_rca8_fa2_4_and0 | u_csamul_pg_rca8_fa2_4_and1;
  assign u_csamul_pg_rca8_and3_4 = a[3] & b[4];
  assign u_csamul_pg_rca8_fa3_4_xor0 = u_csamul_pg_rca8_and3_4 ^ u_csamul_pg_rca8_fa4_3_xor1;
  assign u_csamul_pg_rca8_fa3_4_and0 = u_csamul_pg_rca8_and3_4 & u_csamul_pg_rca8_fa4_3_xor1;
  assign u_csamul_pg_rca8_fa3_4_xor1 = u_csamul_pg_rca8_fa3_4_xor0 ^ u_csamul_pg_rca8_fa3_3_or0;
  assign u_csamul_pg_rca8_fa3_4_and1 = u_csamul_pg_rca8_fa3_4_xor0 & u_csamul_pg_rca8_fa3_3_or0;
  assign u_csamul_pg_rca8_fa3_4_or0 = u_csamul_pg_rca8_fa3_4_and0 | u_csamul_pg_rca8_fa3_4_and1;
  assign u_csamul_pg_rca8_and4_4 = a[4] & b[4];
  assign u_csamul_pg_rca8_fa4_4_xor0 = u_csamul_pg_rca8_and4_4 ^ u_csamul_pg_rca8_fa5_3_xor1;
  assign u_csamul_pg_rca8_fa4_4_and0 = u_csamul_pg_rca8_and4_4 & u_csamul_pg_rca8_fa5_3_xor1;
  assign u_csamul_pg_rca8_fa4_4_xor1 = u_csamul_pg_rca8_fa4_4_xor0 ^ u_csamul_pg_rca8_fa4_3_or0;
  assign u_csamul_pg_rca8_fa4_4_and1 = u_csamul_pg_rca8_fa4_4_xor0 & u_csamul_pg_rca8_fa4_3_or0;
  assign u_csamul_pg_rca8_fa4_4_or0 = u_csamul_pg_rca8_fa4_4_and0 | u_csamul_pg_rca8_fa4_4_and1;
  assign u_csamul_pg_rca8_and5_4 = a[5] & b[4];
  assign u_csamul_pg_rca8_fa5_4_xor0 = u_csamul_pg_rca8_and5_4 ^ u_csamul_pg_rca8_fa6_3_xor1;
  assign u_csamul_pg_rca8_fa5_4_and0 = u_csamul_pg_rca8_and5_4 & u_csamul_pg_rca8_fa6_3_xor1;
  assign u_csamul_pg_rca8_fa5_4_xor1 = u_csamul_pg_rca8_fa5_4_xor0 ^ u_csamul_pg_rca8_fa5_3_or0;
  assign u_csamul_pg_rca8_fa5_4_and1 = u_csamul_pg_rca8_fa5_4_xor0 & u_csamul_pg_rca8_fa5_3_or0;
  assign u_csamul_pg_rca8_fa5_4_or0 = u_csamul_pg_rca8_fa5_4_and0 | u_csamul_pg_rca8_fa5_4_and1;
  assign u_csamul_pg_rca8_and6_4 = a[6] & b[4];
  assign u_csamul_pg_rca8_fa6_4_xor0 = u_csamul_pg_rca8_and6_4 ^ u_csamul_pg_rca8_and7_3;
  assign u_csamul_pg_rca8_fa6_4_and0 = u_csamul_pg_rca8_and6_4 & u_csamul_pg_rca8_and7_3;
  assign u_csamul_pg_rca8_fa6_4_xor1 = u_csamul_pg_rca8_fa6_4_xor0 ^ u_csamul_pg_rca8_fa6_3_or0;
  assign u_csamul_pg_rca8_fa6_4_and1 = u_csamul_pg_rca8_fa6_4_xor0 & u_csamul_pg_rca8_fa6_3_or0;
  assign u_csamul_pg_rca8_fa6_4_or0 = u_csamul_pg_rca8_fa6_4_and0 | u_csamul_pg_rca8_fa6_4_and1;
  assign u_csamul_pg_rca8_and7_4 = a[7] & b[4];
  assign u_csamul_pg_rca8_and0_5 = a[0] & b[5];
  assign u_csamul_pg_rca8_fa0_5_xor0 = u_csamul_pg_rca8_and0_5 ^ u_csamul_pg_rca8_fa1_4_xor1;
  assign u_csamul_pg_rca8_fa0_5_and0 = u_csamul_pg_rca8_and0_5 & u_csamul_pg_rca8_fa1_4_xor1;
  assign u_csamul_pg_rca8_fa0_5_xor1 = u_csamul_pg_rca8_fa0_5_xor0 ^ u_csamul_pg_rca8_fa0_4_or0;
  assign u_csamul_pg_rca8_fa0_5_and1 = u_csamul_pg_rca8_fa0_5_xor0 & u_csamul_pg_rca8_fa0_4_or0;
  assign u_csamul_pg_rca8_fa0_5_or0 = u_csamul_pg_rca8_fa0_5_and0 | u_csamul_pg_rca8_fa0_5_and1;
  assign u_csamul_pg_rca8_and1_5 = a[1] & b[5];
  assign u_csamul_pg_rca8_fa1_5_xor0 = u_csamul_pg_rca8_and1_5 ^ u_csamul_pg_rca8_fa2_4_xor1;
  assign u_csamul_pg_rca8_fa1_5_and0 = u_csamul_pg_rca8_and1_5 & u_csamul_pg_rca8_fa2_4_xor1;
  assign u_csamul_pg_rca8_fa1_5_xor1 = u_csamul_pg_rca8_fa1_5_xor0 ^ u_csamul_pg_rca8_fa1_4_or0;
  assign u_csamul_pg_rca8_fa1_5_and1 = u_csamul_pg_rca8_fa1_5_xor0 & u_csamul_pg_rca8_fa1_4_or0;
  assign u_csamul_pg_rca8_fa1_5_or0 = u_csamul_pg_rca8_fa1_5_and0 | u_csamul_pg_rca8_fa1_5_and1;
  assign u_csamul_pg_rca8_and2_5 = a[2] & b[5];
  assign u_csamul_pg_rca8_fa2_5_xor0 = u_csamul_pg_rca8_and2_5 ^ u_csamul_pg_rca8_fa3_4_xor1;
  assign u_csamul_pg_rca8_fa2_5_and0 = u_csamul_pg_rca8_and2_5 & u_csamul_pg_rca8_fa3_4_xor1;
  assign u_csamul_pg_rca8_fa2_5_xor1 = u_csamul_pg_rca8_fa2_5_xor0 ^ u_csamul_pg_rca8_fa2_4_or0;
  assign u_csamul_pg_rca8_fa2_5_and1 = u_csamul_pg_rca8_fa2_5_xor0 & u_csamul_pg_rca8_fa2_4_or0;
  assign u_csamul_pg_rca8_fa2_5_or0 = u_csamul_pg_rca8_fa2_5_and0 | u_csamul_pg_rca8_fa2_5_and1;
  assign u_csamul_pg_rca8_and3_5 = a[3] & b[5];
  assign u_csamul_pg_rca8_fa3_5_xor0 = u_csamul_pg_rca8_and3_5 ^ u_csamul_pg_rca8_fa4_4_xor1;
  assign u_csamul_pg_rca8_fa3_5_and0 = u_csamul_pg_rca8_and3_5 & u_csamul_pg_rca8_fa4_4_xor1;
  assign u_csamul_pg_rca8_fa3_5_xor1 = u_csamul_pg_rca8_fa3_5_xor0 ^ u_csamul_pg_rca8_fa3_4_or0;
  assign u_csamul_pg_rca8_fa3_5_and1 = u_csamul_pg_rca8_fa3_5_xor0 & u_csamul_pg_rca8_fa3_4_or0;
  assign u_csamul_pg_rca8_fa3_5_or0 = u_csamul_pg_rca8_fa3_5_and0 | u_csamul_pg_rca8_fa3_5_and1;
  assign u_csamul_pg_rca8_and4_5 = a[4] & b[5];
  assign u_csamul_pg_rca8_fa4_5_xor0 = u_csamul_pg_rca8_and4_5 ^ u_csamul_pg_rca8_fa5_4_xor1;
  assign u_csamul_pg_rca8_fa4_5_and0 = u_csamul_pg_rca8_and4_5 & u_csamul_pg_rca8_fa5_4_xor1;
  assign u_csamul_pg_rca8_fa4_5_xor1 = u_csamul_pg_rca8_fa4_5_xor0 ^ u_csamul_pg_rca8_fa4_4_or0;
  assign u_csamul_pg_rca8_fa4_5_and1 = u_csamul_pg_rca8_fa4_5_xor0 & u_csamul_pg_rca8_fa4_4_or0;
  assign u_csamul_pg_rca8_fa4_5_or0 = u_csamul_pg_rca8_fa4_5_and0 | u_csamul_pg_rca8_fa4_5_and1;
  assign u_csamul_pg_rca8_and5_5 = a[5] & b[5];
  assign u_csamul_pg_rca8_fa5_5_xor0 = u_csamul_pg_rca8_and5_5 ^ u_csamul_pg_rca8_fa6_4_xor1;
  assign u_csamul_pg_rca8_fa5_5_and0 = u_csamul_pg_rca8_and5_5 & u_csamul_pg_rca8_fa6_4_xor1;
  assign u_csamul_pg_rca8_fa5_5_xor1 = u_csamul_pg_rca8_fa5_5_xor0 ^ u_csamul_pg_rca8_fa5_4_or0;
  assign u_csamul_pg_rca8_fa5_5_and1 = u_csamul_pg_rca8_fa5_5_xor0 & u_csamul_pg_rca8_fa5_4_or0;
  assign u_csamul_pg_rca8_fa5_5_or0 = u_csamul_pg_rca8_fa5_5_and0 | u_csamul_pg_rca8_fa5_5_and1;
  assign u_csamul_pg_rca8_and6_5 = a[6] & b[5];
  assign u_csamul_pg_rca8_fa6_5_xor0 = u_csamul_pg_rca8_and6_5 ^ u_csamul_pg_rca8_and7_4;
  assign u_csamul_pg_rca8_fa6_5_and0 = u_csamul_pg_rca8_and6_5 & u_csamul_pg_rca8_and7_4;
  assign u_csamul_pg_rca8_fa6_5_xor1 = u_csamul_pg_rca8_fa6_5_xor0 ^ u_csamul_pg_rca8_fa6_4_or0;
  assign u_csamul_pg_rca8_fa6_5_and1 = u_csamul_pg_rca8_fa6_5_xor0 & u_csamul_pg_rca8_fa6_4_or0;
  assign u_csamul_pg_rca8_fa6_5_or0 = u_csamul_pg_rca8_fa6_5_and0 | u_csamul_pg_rca8_fa6_5_and1;
  assign u_csamul_pg_rca8_and7_5 = a[7] & b[5];
  assign u_csamul_pg_rca8_and0_6 = a[0] & b[6];
  assign u_csamul_pg_rca8_fa0_6_xor0 = u_csamul_pg_rca8_and0_6 ^ u_csamul_pg_rca8_fa1_5_xor1;
  assign u_csamul_pg_rca8_fa0_6_and0 = u_csamul_pg_rca8_and0_6 & u_csamul_pg_rca8_fa1_5_xor1;
  assign u_csamul_pg_rca8_fa0_6_xor1 = u_csamul_pg_rca8_fa0_6_xor0 ^ u_csamul_pg_rca8_fa0_5_or0;
  assign u_csamul_pg_rca8_fa0_6_and1 = u_csamul_pg_rca8_fa0_6_xor0 & u_csamul_pg_rca8_fa0_5_or0;
  assign u_csamul_pg_rca8_fa0_6_or0 = u_csamul_pg_rca8_fa0_6_and0 | u_csamul_pg_rca8_fa0_6_and1;
  assign u_csamul_pg_rca8_and1_6 = a[1] & b[6];
  assign u_csamul_pg_rca8_fa1_6_xor0 = u_csamul_pg_rca8_and1_6 ^ u_csamul_pg_rca8_fa2_5_xor1;
  assign u_csamul_pg_rca8_fa1_6_and0 = u_csamul_pg_rca8_and1_6 & u_csamul_pg_rca8_fa2_5_xor1;
  assign u_csamul_pg_rca8_fa1_6_xor1 = u_csamul_pg_rca8_fa1_6_xor0 ^ u_csamul_pg_rca8_fa1_5_or0;
  assign u_csamul_pg_rca8_fa1_6_and1 = u_csamul_pg_rca8_fa1_6_xor0 & u_csamul_pg_rca8_fa1_5_or0;
  assign u_csamul_pg_rca8_fa1_6_or0 = u_csamul_pg_rca8_fa1_6_and0 | u_csamul_pg_rca8_fa1_6_and1;
  assign u_csamul_pg_rca8_and2_6 = a[2] & b[6];
  assign u_csamul_pg_rca8_fa2_6_xor0 = u_csamul_pg_rca8_and2_6 ^ u_csamul_pg_rca8_fa3_5_xor1;
  assign u_csamul_pg_rca8_fa2_6_and0 = u_csamul_pg_rca8_and2_6 & u_csamul_pg_rca8_fa3_5_xor1;
  assign u_csamul_pg_rca8_fa2_6_xor1 = u_csamul_pg_rca8_fa2_6_xor0 ^ u_csamul_pg_rca8_fa2_5_or0;
  assign u_csamul_pg_rca8_fa2_6_and1 = u_csamul_pg_rca8_fa2_6_xor0 & u_csamul_pg_rca8_fa2_5_or0;
  assign u_csamul_pg_rca8_fa2_6_or0 = u_csamul_pg_rca8_fa2_6_and0 | u_csamul_pg_rca8_fa2_6_and1;
  assign u_csamul_pg_rca8_and3_6 = a[3] & b[6];
  assign u_csamul_pg_rca8_fa3_6_xor0 = u_csamul_pg_rca8_and3_6 ^ u_csamul_pg_rca8_fa4_5_xor1;
  assign u_csamul_pg_rca8_fa3_6_and0 = u_csamul_pg_rca8_and3_6 & u_csamul_pg_rca8_fa4_5_xor1;
  assign u_csamul_pg_rca8_fa3_6_xor1 = u_csamul_pg_rca8_fa3_6_xor0 ^ u_csamul_pg_rca8_fa3_5_or0;
  assign u_csamul_pg_rca8_fa3_6_and1 = u_csamul_pg_rca8_fa3_6_xor0 & u_csamul_pg_rca8_fa3_5_or0;
  assign u_csamul_pg_rca8_fa3_6_or0 = u_csamul_pg_rca8_fa3_6_and0 | u_csamul_pg_rca8_fa3_6_and1;
  assign u_csamul_pg_rca8_and4_6 = a[4] & b[6];
  assign u_csamul_pg_rca8_fa4_6_xor0 = u_csamul_pg_rca8_and4_6 ^ u_csamul_pg_rca8_fa5_5_xor1;
  assign u_csamul_pg_rca8_fa4_6_and0 = u_csamul_pg_rca8_and4_6 & u_csamul_pg_rca8_fa5_5_xor1;
  assign u_csamul_pg_rca8_fa4_6_xor1 = u_csamul_pg_rca8_fa4_6_xor0 ^ u_csamul_pg_rca8_fa4_5_or0;
  assign u_csamul_pg_rca8_fa4_6_and1 = u_csamul_pg_rca8_fa4_6_xor0 & u_csamul_pg_rca8_fa4_5_or0;
  assign u_csamul_pg_rca8_fa4_6_or0 = u_csamul_pg_rca8_fa4_6_and0 | u_csamul_pg_rca8_fa4_6_and1;
  assign u_csamul_pg_rca8_and5_6 = a[5] & b[6];
  assign u_csamul_pg_rca8_fa5_6_xor0 = u_csamul_pg_rca8_and5_6 ^ u_csamul_pg_rca8_fa6_5_xor1;
  assign u_csamul_pg_rca8_fa5_6_and0 = u_csamul_pg_rca8_and5_6 & u_csamul_pg_rca8_fa6_5_xor1;
  assign u_csamul_pg_rca8_fa5_6_xor1 = u_csamul_pg_rca8_fa5_6_xor0 ^ u_csamul_pg_rca8_fa5_5_or0;
  assign u_csamul_pg_rca8_fa5_6_and1 = u_csamul_pg_rca8_fa5_6_xor0 & u_csamul_pg_rca8_fa5_5_or0;
  assign u_csamul_pg_rca8_fa5_6_or0 = u_csamul_pg_rca8_fa5_6_and0 | u_csamul_pg_rca8_fa5_6_and1;
  assign u_csamul_pg_rca8_and6_6 = a[6] & b[6];
  assign u_csamul_pg_rca8_fa6_6_xor0 = u_csamul_pg_rca8_and6_6 ^ u_csamul_pg_rca8_and7_5;
  assign u_csamul_pg_rca8_fa6_6_and0 = u_csamul_pg_rca8_and6_6 & u_csamul_pg_rca8_and7_5;
  assign u_csamul_pg_rca8_fa6_6_xor1 = u_csamul_pg_rca8_fa6_6_xor0 ^ u_csamul_pg_rca8_fa6_5_or0;
  assign u_csamul_pg_rca8_fa6_6_and1 = u_csamul_pg_rca8_fa6_6_xor0 & u_csamul_pg_rca8_fa6_5_or0;
  assign u_csamul_pg_rca8_fa6_6_or0 = u_csamul_pg_rca8_fa6_6_and0 | u_csamul_pg_rca8_fa6_6_and1;
  assign u_csamul_pg_rca8_and7_6 = a[7] & b[6];
  assign u_csamul_pg_rca8_and0_7 = a[0] & b[7];
  assign u_csamul_pg_rca8_fa0_7_xor0 = u_csamul_pg_rca8_and0_7 ^ u_csamul_pg_rca8_fa1_6_xor1;
  assign u_csamul_pg_rca8_fa0_7_and0 = u_csamul_pg_rca8_and0_7 & u_csamul_pg_rca8_fa1_6_xor1;
  assign u_csamul_pg_rca8_fa0_7_xor1 = u_csamul_pg_rca8_fa0_7_xor0 ^ u_csamul_pg_rca8_fa0_6_or0;
  assign u_csamul_pg_rca8_fa0_7_and1 = u_csamul_pg_rca8_fa0_7_xor0 & u_csamul_pg_rca8_fa0_6_or0;
  assign u_csamul_pg_rca8_fa0_7_or0 = u_csamul_pg_rca8_fa0_7_and0 | u_csamul_pg_rca8_fa0_7_and1;
  assign u_csamul_pg_rca8_and1_7 = a[1] & b[7];
  assign u_csamul_pg_rca8_fa1_7_xor0 = u_csamul_pg_rca8_and1_7 ^ u_csamul_pg_rca8_fa2_6_xor1;
  assign u_csamul_pg_rca8_fa1_7_and0 = u_csamul_pg_rca8_and1_7 & u_csamul_pg_rca8_fa2_6_xor1;
  assign u_csamul_pg_rca8_fa1_7_xor1 = u_csamul_pg_rca8_fa1_7_xor0 ^ u_csamul_pg_rca8_fa1_6_or0;
  assign u_csamul_pg_rca8_fa1_7_and1 = u_csamul_pg_rca8_fa1_7_xor0 & u_csamul_pg_rca8_fa1_6_or0;
  assign u_csamul_pg_rca8_fa1_7_or0 = u_csamul_pg_rca8_fa1_7_and0 | u_csamul_pg_rca8_fa1_7_and1;
  assign u_csamul_pg_rca8_and2_7 = a[2] & b[7];
  assign u_csamul_pg_rca8_fa2_7_xor0 = u_csamul_pg_rca8_and2_7 ^ u_csamul_pg_rca8_fa3_6_xor1;
  assign u_csamul_pg_rca8_fa2_7_and0 = u_csamul_pg_rca8_and2_7 & u_csamul_pg_rca8_fa3_6_xor1;
  assign u_csamul_pg_rca8_fa2_7_xor1 = u_csamul_pg_rca8_fa2_7_xor0 ^ u_csamul_pg_rca8_fa2_6_or0;
  assign u_csamul_pg_rca8_fa2_7_and1 = u_csamul_pg_rca8_fa2_7_xor0 & u_csamul_pg_rca8_fa2_6_or0;
  assign u_csamul_pg_rca8_fa2_7_or0 = u_csamul_pg_rca8_fa2_7_and0 | u_csamul_pg_rca8_fa2_7_and1;
  assign u_csamul_pg_rca8_and3_7 = a[3] & b[7];
  assign u_csamul_pg_rca8_fa3_7_xor0 = u_csamul_pg_rca8_and3_7 ^ u_csamul_pg_rca8_fa4_6_xor1;
  assign u_csamul_pg_rca8_fa3_7_and0 = u_csamul_pg_rca8_and3_7 & u_csamul_pg_rca8_fa4_6_xor1;
  assign u_csamul_pg_rca8_fa3_7_xor1 = u_csamul_pg_rca8_fa3_7_xor0 ^ u_csamul_pg_rca8_fa3_6_or0;
  assign u_csamul_pg_rca8_fa3_7_and1 = u_csamul_pg_rca8_fa3_7_xor0 & u_csamul_pg_rca8_fa3_6_or0;
  assign u_csamul_pg_rca8_fa3_7_or0 = u_csamul_pg_rca8_fa3_7_and0 | u_csamul_pg_rca8_fa3_7_and1;
  assign u_csamul_pg_rca8_and4_7 = a[4] & b[7];
  assign u_csamul_pg_rca8_fa4_7_xor0 = u_csamul_pg_rca8_and4_7 ^ u_csamul_pg_rca8_fa5_6_xor1;
  assign u_csamul_pg_rca8_fa4_7_and0 = u_csamul_pg_rca8_and4_7 & u_csamul_pg_rca8_fa5_6_xor1;
  assign u_csamul_pg_rca8_fa4_7_xor1 = u_csamul_pg_rca8_fa4_7_xor0 ^ u_csamul_pg_rca8_fa4_6_or0;
  assign u_csamul_pg_rca8_fa4_7_and1 = u_csamul_pg_rca8_fa4_7_xor0 & u_csamul_pg_rca8_fa4_6_or0;
  assign u_csamul_pg_rca8_fa4_7_or0 = u_csamul_pg_rca8_fa4_7_and0 | u_csamul_pg_rca8_fa4_7_and1;
  assign u_csamul_pg_rca8_and5_7 = a[5] & b[7];
  assign u_csamul_pg_rca8_fa5_7_xor0 = u_csamul_pg_rca8_and5_7 ^ u_csamul_pg_rca8_fa6_6_xor1;
  assign u_csamul_pg_rca8_fa5_7_and0 = u_csamul_pg_rca8_and5_7 & u_csamul_pg_rca8_fa6_6_xor1;
  assign u_csamul_pg_rca8_fa5_7_xor1 = u_csamul_pg_rca8_fa5_7_xor0 ^ u_csamul_pg_rca8_fa5_6_or0;
  assign u_csamul_pg_rca8_fa5_7_and1 = u_csamul_pg_rca8_fa5_7_xor0 & u_csamul_pg_rca8_fa5_6_or0;
  assign u_csamul_pg_rca8_fa5_7_or0 = u_csamul_pg_rca8_fa5_7_and0 | u_csamul_pg_rca8_fa5_7_and1;
  assign u_csamul_pg_rca8_and6_7 = a[6] & b[7];
  assign u_csamul_pg_rca8_fa6_7_xor0 = u_csamul_pg_rca8_and6_7 ^ u_csamul_pg_rca8_and7_6;
  assign u_csamul_pg_rca8_fa6_7_and0 = u_csamul_pg_rca8_and6_7 & u_csamul_pg_rca8_and7_6;
  assign u_csamul_pg_rca8_fa6_7_xor1 = u_csamul_pg_rca8_fa6_7_xor0 ^ u_csamul_pg_rca8_fa6_6_or0;
  assign u_csamul_pg_rca8_fa6_7_and1 = u_csamul_pg_rca8_fa6_7_xor0 & u_csamul_pg_rca8_fa6_6_or0;
  assign u_csamul_pg_rca8_fa6_7_or0 = u_csamul_pg_rca8_fa6_7_and0 | u_csamul_pg_rca8_fa6_7_and1;
  assign u_csamul_pg_rca8_and7_7 = a[7] & b[7];
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa0_xor0 = u_csamul_pg_rca8_fa1_7_xor1 ^ u_csamul_pg_rca8_fa0_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa0_and0 = u_csamul_pg_rca8_fa1_7_xor1 & u_csamul_pg_rca8_fa0_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor0 = u_csamul_pg_rca8_fa2_7_xor1 ^ u_csamul_pg_rca8_fa1_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa1_and0 = u_csamul_pg_rca8_fa2_7_xor1 & u_csamul_pg_rca8_fa1_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor0 ^ u_csamul_pg_rca8_u_pg_rca8_pg_fa0_and0;
  assign u_csamul_pg_rca8_u_pg_rca8_and1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa0_and0 & u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor0;
  assign u_csamul_pg_rca8_u_pg_rca8_or1 = u_csamul_pg_rca8_u_pg_rca8_and1 | u_csamul_pg_rca8_u_pg_rca8_pg_fa1_and0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor0 = u_csamul_pg_rca8_fa3_7_xor1 ^ u_csamul_pg_rca8_fa2_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa2_and0 = u_csamul_pg_rca8_fa3_7_xor1 & u_csamul_pg_rca8_fa2_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor0 ^ u_csamul_pg_rca8_u_pg_rca8_or1;
  assign u_csamul_pg_rca8_u_pg_rca8_and2 = u_csamul_pg_rca8_u_pg_rca8_or1 & u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor0;
  assign u_csamul_pg_rca8_u_pg_rca8_or2 = u_csamul_pg_rca8_u_pg_rca8_and2 | u_csamul_pg_rca8_u_pg_rca8_pg_fa2_and0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor0 = u_csamul_pg_rca8_fa4_7_xor1 ^ u_csamul_pg_rca8_fa3_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa3_and0 = u_csamul_pg_rca8_fa4_7_xor1 & u_csamul_pg_rca8_fa3_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor0 ^ u_csamul_pg_rca8_u_pg_rca8_or2;
  assign u_csamul_pg_rca8_u_pg_rca8_and3 = u_csamul_pg_rca8_u_pg_rca8_or2 & u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor0;
  assign u_csamul_pg_rca8_u_pg_rca8_or3 = u_csamul_pg_rca8_u_pg_rca8_and3 | u_csamul_pg_rca8_u_pg_rca8_pg_fa3_and0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor0 = u_csamul_pg_rca8_fa5_7_xor1 ^ u_csamul_pg_rca8_fa4_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa4_and0 = u_csamul_pg_rca8_fa5_7_xor1 & u_csamul_pg_rca8_fa4_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor0 ^ u_csamul_pg_rca8_u_pg_rca8_or3;
  assign u_csamul_pg_rca8_u_pg_rca8_and4 = u_csamul_pg_rca8_u_pg_rca8_or3 & u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor0;
  assign u_csamul_pg_rca8_u_pg_rca8_or4 = u_csamul_pg_rca8_u_pg_rca8_and4 | u_csamul_pg_rca8_u_pg_rca8_pg_fa4_and0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor0 = u_csamul_pg_rca8_fa6_7_xor1 ^ u_csamul_pg_rca8_fa5_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa5_and0 = u_csamul_pg_rca8_fa6_7_xor1 & u_csamul_pg_rca8_fa5_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor0 ^ u_csamul_pg_rca8_u_pg_rca8_or4;
  assign u_csamul_pg_rca8_u_pg_rca8_and5 = u_csamul_pg_rca8_u_pg_rca8_or4 & u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor0;
  assign u_csamul_pg_rca8_u_pg_rca8_or5 = u_csamul_pg_rca8_u_pg_rca8_and5 | u_csamul_pg_rca8_u_pg_rca8_pg_fa5_and0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor0 = u_csamul_pg_rca8_and7_7 ^ u_csamul_pg_rca8_fa6_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa6_and0 = u_csamul_pg_rca8_and7_7 & u_csamul_pg_rca8_fa6_7_or0;
  assign u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor1 = u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor0 ^ u_csamul_pg_rca8_u_pg_rca8_or5;
  assign u_csamul_pg_rca8_u_pg_rca8_and6 = u_csamul_pg_rca8_u_pg_rca8_or5 & u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor0;
  assign u_csamul_pg_rca8_u_pg_rca8_or6 = u_csamul_pg_rca8_u_pg_rca8_and6 | u_csamul_pg_rca8_u_pg_rca8_pg_fa6_and0;

  assign u_csamul_pg_rca8_out[0] = u_csamul_pg_rca8_and0_0;
  assign u_csamul_pg_rca8_out[1] = u_csamul_pg_rca8_ha0_1_xor0;
  assign u_csamul_pg_rca8_out[2] = u_csamul_pg_rca8_fa0_2_xor1;
  assign u_csamul_pg_rca8_out[3] = u_csamul_pg_rca8_fa0_3_xor1;
  assign u_csamul_pg_rca8_out[4] = u_csamul_pg_rca8_fa0_4_xor1;
  assign u_csamul_pg_rca8_out[5] = u_csamul_pg_rca8_fa0_5_xor1;
  assign u_csamul_pg_rca8_out[6] = u_csamul_pg_rca8_fa0_6_xor1;
  assign u_csamul_pg_rca8_out[7] = u_csamul_pg_rca8_fa0_7_xor1;
  assign u_csamul_pg_rca8_out[8] = u_csamul_pg_rca8_u_pg_rca8_pg_fa0_xor0;
  assign u_csamul_pg_rca8_out[9] = u_csamul_pg_rca8_u_pg_rca8_pg_fa1_xor1;
  assign u_csamul_pg_rca8_out[10] = u_csamul_pg_rca8_u_pg_rca8_pg_fa2_xor1;
  assign u_csamul_pg_rca8_out[11] = u_csamul_pg_rca8_u_pg_rca8_pg_fa3_xor1;
  assign u_csamul_pg_rca8_out[12] = u_csamul_pg_rca8_u_pg_rca8_pg_fa4_xor1;
  assign u_csamul_pg_rca8_out[13] = u_csamul_pg_rca8_u_pg_rca8_pg_fa5_xor1;
  assign u_csamul_pg_rca8_out[14] = u_csamul_pg_rca8_u_pg_rca8_pg_fa6_xor1;
  assign u_csamul_pg_rca8_out[15] = u_csamul_pg_rca8_u_pg_rca8_or6;
endmodule