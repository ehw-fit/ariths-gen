module f_arrdiv16(input [15:0] a, input [15:0] b, output [15:0] f_arrdiv16_out);
  wire f_arrdiv16_fs0_xor0;
  wire f_arrdiv16_fs0_not0;
  wire f_arrdiv16_fs0_and0;
  wire f_arrdiv16_fs0_not1;
  wire f_arrdiv16_fs1_xor1;
  wire f_arrdiv16_fs1_not1;
  wire f_arrdiv16_fs1_and1;
  wire f_arrdiv16_fs1_or0;
  wire f_arrdiv16_fs2_xor1;
  wire f_arrdiv16_fs2_not1;
  wire f_arrdiv16_fs2_and1;
  wire f_arrdiv16_fs2_or0;
  wire f_arrdiv16_fs3_xor1;
  wire f_arrdiv16_fs3_not1;
  wire f_arrdiv16_fs3_and1;
  wire f_arrdiv16_fs3_or0;
  wire f_arrdiv16_fs4_xor1;
  wire f_arrdiv16_fs4_not1;
  wire f_arrdiv16_fs4_and1;
  wire f_arrdiv16_fs4_or0;
  wire f_arrdiv16_fs5_xor1;
  wire f_arrdiv16_fs5_not1;
  wire f_arrdiv16_fs5_and1;
  wire f_arrdiv16_fs5_or0;
  wire f_arrdiv16_fs6_xor1;
  wire f_arrdiv16_fs6_not1;
  wire f_arrdiv16_fs6_and1;
  wire f_arrdiv16_fs6_or0;
  wire f_arrdiv16_fs7_xor1;
  wire f_arrdiv16_fs7_not1;
  wire f_arrdiv16_fs7_and1;
  wire f_arrdiv16_fs7_or0;
  wire f_arrdiv16_fs8_xor1;
  wire f_arrdiv16_fs8_not1;
  wire f_arrdiv16_fs8_and1;
  wire f_arrdiv16_fs8_or0;
  wire f_arrdiv16_fs9_xor1;
  wire f_arrdiv16_fs9_not1;
  wire f_arrdiv16_fs9_and1;
  wire f_arrdiv16_fs9_or0;
  wire f_arrdiv16_fs10_xor1;
  wire f_arrdiv16_fs10_not1;
  wire f_arrdiv16_fs10_and1;
  wire f_arrdiv16_fs10_or0;
  wire f_arrdiv16_fs11_xor1;
  wire f_arrdiv16_fs11_not1;
  wire f_arrdiv16_fs11_and1;
  wire f_arrdiv16_fs11_or0;
  wire f_arrdiv16_fs12_xor1;
  wire f_arrdiv16_fs12_not1;
  wire f_arrdiv16_fs12_and1;
  wire f_arrdiv16_fs12_or0;
  wire f_arrdiv16_fs13_xor1;
  wire f_arrdiv16_fs13_not1;
  wire f_arrdiv16_fs13_and1;
  wire f_arrdiv16_fs13_or0;
  wire f_arrdiv16_fs14_xor1;
  wire f_arrdiv16_fs14_not1;
  wire f_arrdiv16_fs14_and1;
  wire f_arrdiv16_fs14_or0;
  wire f_arrdiv16_fs15_xor1;
  wire f_arrdiv16_fs15_not1;
  wire f_arrdiv16_fs15_and1;
  wire f_arrdiv16_fs15_or0;
  wire f_arrdiv16_mux2to10_and0;
  wire f_arrdiv16_mux2to10_not0;
  wire f_arrdiv16_mux2to10_and1;
  wire f_arrdiv16_mux2to10_xor0;
  wire f_arrdiv16_mux2to11_not0;
  wire f_arrdiv16_mux2to11_and1;
  wire f_arrdiv16_mux2to12_not0;
  wire f_arrdiv16_mux2to12_and1;
  wire f_arrdiv16_mux2to13_not0;
  wire f_arrdiv16_mux2to13_and1;
  wire f_arrdiv16_mux2to14_not0;
  wire f_arrdiv16_mux2to14_and1;
  wire f_arrdiv16_mux2to15_not0;
  wire f_arrdiv16_mux2to15_and1;
  wire f_arrdiv16_mux2to16_not0;
  wire f_arrdiv16_mux2to16_and1;
  wire f_arrdiv16_mux2to17_not0;
  wire f_arrdiv16_mux2to17_and1;
  wire f_arrdiv16_mux2to18_not0;
  wire f_arrdiv16_mux2to18_and1;
  wire f_arrdiv16_mux2to19_not0;
  wire f_arrdiv16_mux2to19_and1;
  wire f_arrdiv16_mux2to110_not0;
  wire f_arrdiv16_mux2to110_and1;
  wire f_arrdiv16_mux2to111_not0;
  wire f_arrdiv16_mux2to111_and1;
  wire f_arrdiv16_mux2to112_not0;
  wire f_arrdiv16_mux2to112_and1;
  wire f_arrdiv16_mux2to113_not0;
  wire f_arrdiv16_mux2to113_and1;
  wire f_arrdiv16_mux2to114_not0;
  wire f_arrdiv16_mux2to114_and1;
  wire f_arrdiv16_not0;
  wire f_arrdiv16_fs16_xor0;
  wire f_arrdiv16_fs16_not0;
  wire f_arrdiv16_fs16_and0;
  wire f_arrdiv16_fs16_not1;
  wire f_arrdiv16_fs17_xor0;
  wire f_arrdiv16_fs17_not0;
  wire f_arrdiv16_fs17_and0;
  wire f_arrdiv16_fs17_xor1;
  wire f_arrdiv16_fs17_not1;
  wire f_arrdiv16_fs17_and1;
  wire f_arrdiv16_fs17_or0;
  wire f_arrdiv16_fs18_xor0;
  wire f_arrdiv16_fs18_not0;
  wire f_arrdiv16_fs18_and0;
  wire f_arrdiv16_fs18_xor1;
  wire f_arrdiv16_fs18_not1;
  wire f_arrdiv16_fs18_and1;
  wire f_arrdiv16_fs18_or0;
  wire f_arrdiv16_fs19_xor0;
  wire f_arrdiv16_fs19_not0;
  wire f_arrdiv16_fs19_and0;
  wire f_arrdiv16_fs19_xor1;
  wire f_arrdiv16_fs19_not1;
  wire f_arrdiv16_fs19_and1;
  wire f_arrdiv16_fs19_or0;
  wire f_arrdiv16_fs20_xor0;
  wire f_arrdiv16_fs20_not0;
  wire f_arrdiv16_fs20_and0;
  wire f_arrdiv16_fs20_xor1;
  wire f_arrdiv16_fs20_not1;
  wire f_arrdiv16_fs20_and1;
  wire f_arrdiv16_fs20_or0;
  wire f_arrdiv16_fs21_xor0;
  wire f_arrdiv16_fs21_not0;
  wire f_arrdiv16_fs21_and0;
  wire f_arrdiv16_fs21_xor1;
  wire f_arrdiv16_fs21_not1;
  wire f_arrdiv16_fs21_and1;
  wire f_arrdiv16_fs21_or0;
  wire f_arrdiv16_fs22_xor0;
  wire f_arrdiv16_fs22_not0;
  wire f_arrdiv16_fs22_and0;
  wire f_arrdiv16_fs22_xor1;
  wire f_arrdiv16_fs22_not1;
  wire f_arrdiv16_fs22_and1;
  wire f_arrdiv16_fs22_or0;
  wire f_arrdiv16_fs23_xor0;
  wire f_arrdiv16_fs23_not0;
  wire f_arrdiv16_fs23_and0;
  wire f_arrdiv16_fs23_xor1;
  wire f_arrdiv16_fs23_not1;
  wire f_arrdiv16_fs23_and1;
  wire f_arrdiv16_fs23_or0;
  wire f_arrdiv16_fs24_xor0;
  wire f_arrdiv16_fs24_not0;
  wire f_arrdiv16_fs24_and0;
  wire f_arrdiv16_fs24_xor1;
  wire f_arrdiv16_fs24_not1;
  wire f_arrdiv16_fs24_and1;
  wire f_arrdiv16_fs24_or0;
  wire f_arrdiv16_fs25_xor0;
  wire f_arrdiv16_fs25_not0;
  wire f_arrdiv16_fs25_and0;
  wire f_arrdiv16_fs25_xor1;
  wire f_arrdiv16_fs25_not1;
  wire f_arrdiv16_fs25_and1;
  wire f_arrdiv16_fs25_or0;
  wire f_arrdiv16_fs26_xor0;
  wire f_arrdiv16_fs26_not0;
  wire f_arrdiv16_fs26_and0;
  wire f_arrdiv16_fs26_xor1;
  wire f_arrdiv16_fs26_not1;
  wire f_arrdiv16_fs26_and1;
  wire f_arrdiv16_fs26_or0;
  wire f_arrdiv16_fs27_xor0;
  wire f_arrdiv16_fs27_not0;
  wire f_arrdiv16_fs27_and0;
  wire f_arrdiv16_fs27_xor1;
  wire f_arrdiv16_fs27_not1;
  wire f_arrdiv16_fs27_and1;
  wire f_arrdiv16_fs27_or0;
  wire f_arrdiv16_fs28_xor0;
  wire f_arrdiv16_fs28_not0;
  wire f_arrdiv16_fs28_and0;
  wire f_arrdiv16_fs28_xor1;
  wire f_arrdiv16_fs28_not1;
  wire f_arrdiv16_fs28_and1;
  wire f_arrdiv16_fs28_or0;
  wire f_arrdiv16_fs29_xor0;
  wire f_arrdiv16_fs29_not0;
  wire f_arrdiv16_fs29_and0;
  wire f_arrdiv16_fs29_xor1;
  wire f_arrdiv16_fs29_not1;
  wire f_arrdiv16_fs29_and1;
  wire f_arrdiv16_fs29_or0;
  wire f_arrdiv16_fs30_xor0;
  wire f_arrdiv16_fs30_not0;
  wire f_arrdiv16_fs30_and0;
  wire f_arrdiv16_fs30_xor1;
  wire f_arrdiv16_fs30_not1;
  wire f_arrdiv16_fs30_and1;
  wire f_arrdiv16_fs30_or0;
  wire f_arrdiv16_fs31_xor0;
  wire f_arrdiv16_fs31_not0;
  wire f_arrdiv16_fs31_and0;
  wire f_arrdiv16_fs31_xor1;
  wire f_arrdiv16_fs31_not1;
  wire f_arrdiv16_fs31_and1;
  wire f_arrdiv16_fs31_or0;
  wire f_arrdiv16_mux2to115_and0;
  wire f_arrdiv16_mux2to115_not0;
  wire f_arrdiv16_mux2to115_and1;
  wire f_arrdiv16_mux2to115_xor0;
  wire f_arrdiv16_mux2to116_and0;
  wire f_arrdiv16_mux2to116_not0;
  wire f_arrdiv16_mux2to116_and1;
  wire f_arrdiv16_mux2to116_xor0;
  wire f_arrdiv16_mux2to117_and0;
  wire f_arrdiv16_mux2to117_not0;
  wire f_arrdiv16_mux2to117_and1;
  wire f_arrdiv16_mux2to117_xor0;
  wire f_arrdiv16_mux2to118_and0;
  wire f_arrdiv16_mux2to118_not0;
  wire f_arrdiv16_mux2to118_and1;
  wire f_arrdiv16_mux2to118_xor0;
  wire f_arrdiv16_mux2to119_and0;
  wire f_arrdiv16_mux2to119_not0;
  wire f_arrdiv16_mux2to119_and1;
  wire f_arrdiv16_mux2to119_xor0;
  wire f_arrdiv16_mux2to120_and0;
  wire f_arrdiv16_mux2to120_not0;
  wire f_arrdiv16_mux2to120_and1;
  wire f_arrdiv16_mux2to120_xor0;
  wire f_arrdiv16_mux2to121_and0;
  wire f_arrdiv16_mux2to121_not0;
  wire f_arrdiv16_mux2to121_and1;
  wire f_arrdiv16_mux2to121_xor0;
  wire f_arrdiv16_mux2to122_and0;
  wire f_arrdiv16_mux2to122_not0;
  wire f_arrdiv16_mux2to122_and1;
  wire f_arrdiv16_mux2to122_xor0;
  wire f_arrdiv16_mux2to123_and0;
  wire f_arrdiv16_mux2to123_not0;
  wire f_arrdiv16_mux2to123_and1;
  wire f_arrdiv16_mux2to123_xor0;
  wire f_arrdiv16_mux2to124_and0;
  wire f_arrdiv16_mux2to124_not0;
  wire f_arrdiv16_mux2to124_and1;
  wire f_arrdiv16_mux2to124_xor0;
  wire f_arrdiv16_mux2to125_and0;
  wire f_arrdiv16_mux2to125_not0;
  wire f_arrdiv16_mux2to125_and1;
  wire f_arrdiv16_mux2to125_xor0;
  wire f_arrdiv16_mux2to126_and0;
  wire f_arrdiv16_mux2to126_not0;
  wire f_arrdiv16_mux2to126_and1;
  wire f_arrdiv16_mux2to126_xor0;
  wire f_arrdiv16_mux2to127_and0;
  wire f_arrdiv16_mux2to127_not0;
  wire f_arrdiv16_mux2to127_and1;
  wire f_arrdiv16_mux2to127_xor0;
  wire f_arrdiv16_mux2to128_and0;
  wire f_arrdiv16_mux2to128_not0;
  wire f_arrdiv16_mux2to128_and1;
  wire f_arrdiv16_mux2to128_xor0;
  wire f_arrdiv16_mux2to129_and0;
  wire f_arrdiv16_mux2to129_not0;
  wire f_arrdiv16_mux2to129_and1;
  wire f_arrdiv16_mux2to129_xor0;
  wire f_arrdiv16_not1;
  wire f_arrdiv16_fs32_xor0;
  wire f_arrdiv16_fs32_not0;
  wire f_arrdiv16_fs32_and0;
  wire f_arrdiv16_fs32_not1;
  wire f_arrdiv16_fs33_xor0;
  wire f_arrdiv16_fs33_not0;
  wire f_arrdiv16_fs33_and0;
  wire f_arrdiv16_fs33_xor1;
  wire f_arrdiv16_fs33_not1;
  wire f_arrdiv16_fs33_and1;
  wire f_arrdiv16_fs33_or0;
  wire f_arrdiv16_fs34_xor0;
  wire f_arrdiv16_fs34_not0;
  wire f_arrdiv16_fs34_and0;
  wire f_arrdiv16_fs34_xor1;
  wire f_arrdiv16_fs34_not1;
  wire f_arrdiv16_fs34_and1;
  wire f_arrdiv16_fs34_or0;
  wire f_arrdiv16_fs35_xor0;
  wire f_arrdiv16_fs35_not0;
  wire f_arrdiv16_fs35_and0;
  wire f_arrdiv16_fs35_xor1;
  wire f_arrdiv16_fs35_not1;
  wire f_arrdiv16_fs35_and1;
  wire f_arrdiv16_fs35_or0;
  wire f_arrdiv16_fs36_xor0;
  wire f_arrdiv16_fs36_not0;
  wire f_arrdiv16_fs36_and0;
  wire f_arrdiv16_fs36_xor1;
  wire f_arrdiv16_fs36_not1;
  wire f_arrdiv16_fs36_and1;
  wire f_arrdiv16_fs36_or0;
  wire f_arrdiv16_fs37_xor0;
  wire f_arrdiv16_fs37_not0;
  wire f_arrdiv16_fs37_and0;
  wire f_arrdiv16_fs37_xor1;
  wire f_arrdiv16_fs37_not1;
  wire f_arrdiv16_fs37_and1;
  wire f_arrdiv16_fs37_or0;
  wire f_arrdiv16_fs38_xor0;
  wire f_arrdiv16_fs38_not0;
  wire f_arrdiv16_fs38_and0;
  wire f_arrdiv16_fs38_xor1;
  wire f_arrdiv16_fs38_not1;
  wire f_arrdiv16_fs38_and1;
  wire f_arrdiv16_fs38_or0;
  wire f_arrdiv16_fs39_xor0;
  wire f_arrdiv16_fs39_not0;
  wire f_arrdiv16_fs39_and0;
  wire f_arrdiv16_fs39_xor1;
  wire f_arrdiv16_fs39_not1;
  wire f_arrdiv16_fs39_and1;
  wire f_arrdiv16_fs39_or0;
  wire f_arrdiv16_fs40_xor0;
  wire f_arrdiv16_fs40_not0;
  wire f_arrdiv16_fs40_and0;
  wire f_arrdiv16_fs40_xor1;
  wire f_arrdiv16_fs40_not1;
  wire f_arrdiv16_fs40_and1;
  wire f_arrdiv16_fs40_or0;
  wire f_arrdiv16_fs41_xor0;
  wire f_arrdiv16_fs41_not0;
  wire f_arrdiv16_fs41_and0;
  wire f_arrdiv16_fs41_xor1;
  wire f_arrdiv16_fs41_not1;
  wire f_arrdiv16_fs41_and1;
  wire f_arrdiv16_fs41_or0;
  wire f_arrdiv16_fs42_xor0;
  wire f_arrdiv16_fs42_not0;
  wire f_arrdiv16_fs42_and0;
  wire f_arrdiv16_fs42_xor1;
  wire f_arrdiv16_fs42_not1;
  wire f_arrdiv16_fs42_and1;
  wire f_arrdiv16_fs42_or0;
  wire f_arrdiv16_fs43_xor0;
  wire f_arrdiv16_fs43_not0;
  wire f_arrdiv16_fs43_and0;
  wire f_arrdiv16_fs43_xor1;
  wire f_arrdiv16_fs43_not1;
  wire f_arrdiv16_fs43_and1;
  wire f_arrdiv16_fs43_or0;
  wire f_arrdiv16_fs44_xor0;
  wire f_arrdiv16_fs44_not0;
  wire f_arrdiv16_fs44_and0;
  wire f_arrdiv16_fs44_xor1;
  wire f_arrdiv16_fs44_not1;
  wire f_arrdiv16_fs44_and1;
  wire f_arrdiv16_fs44_or0;
  wire f_arrdiv16_fs45_xor0;
  wire f_arrdiv16_fs45_not0;
  wire f_arrdiv16_fs45_and0;
  wire f_arrdiv16_fs45_xor1;
  wire f_arrdiv16_fs45_not1;
  wire f_arrdiv16_fs45_and1;
  wire f_arrdiv16_fs45_or0;
  wire f_arrdiv16_fs46_xor0;
  wire f_arrdiv16_fs46_not0;
  wire f_arrdiv16_fs46_and0;
  wire f_arrdiv16_fs46_xor1;
  wire f_arrdiv16_fs46_not1;
  wire f_arrdiv16_fs46_and1;
  wire f_arrdiv16_fs46_or0;
  wire f_arrdiv16_fs47_xor0;
  wire f_arrdiv16_fs47_not0;
  wire f_arrdiv16_fs47_and0;
  wire f_arrdiv16_fs47_xor1;
  wire f_arrdiv16_fs47_not1;
  wire f_arrdiv16_fs47_and1;
  wire f_arrdiv16_fs47_or0;
  wire f_arrdiv16_mux2to130_and0;
  wire f_arrdiv16_mux2to130_not0;
  wire f_arrdiv16_mux2to130_and1;
  wire f_arrdiv16_mux2to130_xor0;
  wire f_arrdiv16_mux2to131_and0;
  wire f_arrdiv16_mux2to131_not0;
  wire f_arrdiv16_mux2to131_and1;
  wire f_arrdiv16_mux2to131_xor0;
  wire f_arrdiv16_mux2to132_and0;
  wire f_arrdiv16_mux2to132_not0;
  wire f_arrdiv16_mux2to132_and1;
  wire f_arrdiv16_mux2to132_xor0;
  wire f_arrdiv16_mux2to133_and0;
  wire f_arrdiv16_mux2to133_not0;
  wire f_arrdiv16_mux2to133_and1;
  wire f_arrdiv16_mux2to133_xor0;
  wire f_arrdiv16_mux2to134_and0;
  wire f_arrdiv16_mux2to134_not0;
  wire f_arrdiv16_mux2to134_and1;
  wire f_arrdiv16_mux2to134_xor0;
  wire f_arrdiv16_mux2to135_and0;
  wire f_arrdiv16_mux2to135_not0;
  wire f_arrdiv16_mux2to135_and1;
  wire f_arrdiv16_mux2to135_xor0;
  wire f_arrdiv16_mux2to136_and0;
  wire f_arrdiv16_mux2to136_not0;
  wire f_arrdiv16_mux2to136_and1;
  wire f_arrdiv16_mux2to136_xor0;
  wire f_arrdiv16_mux2to137_and0;
  wire f_arrdiv16_mux2to137_not0;
  wire f_arrdiv16_mux2to137_and1;
  wire f_arrdiv16_mux2to137_xor0;
  wire f_arrdiv16_mux2to138_and0;
  wire f_arrdiv16_mux2to138_not0;
  wire f_arrdiv16_mux2to138_and1;
  wire f_arrdiv16_mux2to138_xor0;
  wire f_arrdiv16_mux2to139_and0;
  wire f_arrdiv16_mux2to139_not0;
  wire f_arrdiv16_mux2to139_and1;
  wire f_arrdiv16_mux2to139_xor0;
  wire f_arrdiv16_mux2to140_and0;
  wire f_arrdiv16_mux2to140_not0;
  wire f_arrdiv16_mux2to140_and1;
  wire f_arrdiv16_mux2to140_xor0;
  wire f_arrdiv16_mux2to141_and0;
  wire f_arrdiv16_mux2to141_not0;
  wire f_arrdiv16_mux2to141_and1;
  wire f_arrdiv16_mux2to141_xor0;
  wire f_arrdiv16_mux2to142_and0;
  wire f_arrdiv16_mux2to142_not0;
  wire f_arrdiv16_mux2to142_and1;
  wire f_arrdiv16_mux2to142_xor0;
  wire f_arrdiv16_mux2to143_and0;
  wire f_arrdiv16_mux2to143_not0;
  wire f_arrdiv16_mux2to143_and1;
  wire f_arrdiv16_mux2to143_xor0;
  wire f_arrdiv16_mux2to144_and0;
  wire f_arrdiv16_mux2to144_not0;
  wire f_arrdiv16_mux2to144_and1;
  wire f_arrdiv16_mux2to144_xor0;
  wire f_arrdiv16_not2;
  wire f_arrdiv16_fs48_xor0;
  wire f_arrdiv16_fs48_not0;
  wire f_arrdiv16_fs48_and0;
  wire f_arrdiv16_fs48_not1;
  wire f_arrdiv16_fs49_xor0;
  wire f_arrdiv16_fs49_not0;
  wire f_arrdiv16_fs49_and0;
  wire f_arrdiv16_fs49_xor1;
  wire f_arrdiv16_fs49_not1;
  wire f_arrdiv16_fs49_and1;
  wire f_arrdiv16_fs49_or0;
  wire f_arrdiv16_fs50_xor0;
  wire f_arrdiv16_fs50_not0;
  wire f_arrdiv16_fs50_and0;
  wire f_arrdiv16_fs50_xor1;
  wire f_arrdiv16_fs50_not1;
  wire f_arrdiv16_fs50_and1;
  wire f_arrdiv16_fs50_or0;
  wire f_arrdiv16_fs51_xor0;
  wire f_arrdiv16_fs51_not0;
  wire f_arrdiv16_fs51_and0;
  wire f_arrdiv16_fs51_xor1;
  wire f_arrdiv16_fs51_not1;
  wire f_arrdiv16_fs51_and1;
  wire f_arrdiv16_fs51_or0;
  wire f_arrdiv16_fs52_xor0;
  wire f_arrdiv16_fs52_not0;
  wire f_arrdiv16_fs52_and0;
  wire f_arrdiv16_fs52_xor1;
  wire f_arrdiv16_fs52_not1;
  wire f_arrdiv16_fs52_and1;
  wire f_arrdiv16_fs52_or0;
  wire f_arrdiv16_fs53_xor0;
  wire f_arrdiv16_fs53_not0;
  wire f_arrdiv16_fs53_and0;
  wire f_arrdiv16_fs53_xor1;
  wire f_arrdiv16_fs53_not1;
  wire f_arrdiv16_fs53_and1;
  wire f_arrdiv16_fs53_or0;
  wire f_arrdiv16_fs54_xor0;
  wire f_arrdiv16_fs54_not0;
  wire f_arrdiv16_fs54_and0;
  wire f_arrdiv16_fs54_xor1;
  wire f_arrdiv16_fs54_not1;
  wire f_arrdiv16_fs54_and1;
  wire f_arrdiv16_fs54_or0;
  wire f_arrdiv16_fs55_xor0;
  wire f_arrdiv16_fs55_not0;
  wire f_arrdiv16_fs55_and0;
  wire f_arrdiv16_fs55_xor1;
  wire f_arrdiv16_fs55_not1;
  wire f_arrdiv16_fs55_and1;
  wire f_arrdiv16_fs55_or0;
  wire f_arrdiv16_fs56_xor0;
  wire f_arrdiv16_fs56_not0;
  wire f_arrdiv16_fs56_and0;
  wire f_arrdiv16_fs56_xor1;
  wire f_arrdiv16_fs56_not1;
  wire f_arrdiv16_fs56_and1;
  wire f_arrdiv16_fs56_or0;
  wire f_arrdiv16_fs57_xor0;
  wire f_arrdiv16_fs57_not0;
  wire f_arrdiv16_fs57_and0;
  wire f_arrdiv16_fs57_xor1;
  wire f_arrdiv16_fs57_not1;
  wire f_arrdiv16_fs57_and1;
  wire f_arrdiv16_fs57_or0;
  wire f_arrdiv16_fs58_xor0;
  wire f_arrdiv16_fs58_not0;
  wire f_arrdiv16_fs58_and0;
  wire f_arrdiv16_fs58_xor1;
  wire f_arrdiv16_fs58_not1;
  wire f_arrdiv16_fs58_and1;
  wire f_arrdiv16_fs58_or0;
  wire f_arrdiv16_fs59_xor0;
  wire f_arrdiv16_fs59_not0;
  wire f_arrdiv16_fs59_and0;
  wire f_arrdiv16_fs59_xor1;
  wire f_arrdiv16_fs59_not1;
  wire f_arrdiv16_fs59_and1;
  wire f_arrdiv16_fs59_or0;
  wire f_arrdiv16_fs60_xor0;
  wire f_arrdiv16_fs60_not0;
  wire f_arrdiv16_fs60_and0;
  wire f_arrdiv16_fs60_xor1;
  wire f_arrdiv16_fs60_not1;
  wire f_arrdiv16_fs60_and1;
  wire f_arrdiv16_fs60_or0;
  wire f_arrdiv16_fs61_xor0;
  wire f_arrdiv16_fs61_not0;
  wire f_arrdiv16_fs61_and0;
  wire f_arrdiv16_fs61_xor1;
  wire f_arrdiv16_fs61_not1;
  wire f_arrdiv16_fs61_and1;
  wire f_arrdiv16_fs61_or0;
  wire f_arrdiv16_fs62_xor0;
  wire f_arrdiv16_fs62_not0;
  wire f_arrdiv16_fs62_and0;
  wire f_arrdiv16_fs62_xor1;
  wire f_arrdiv16_fs62_not1;
  wire f_arrdiv16_fs62_and1;
  wire f_arrdiv16_fs62_or0;
  wire f_arrdiv16_fs63_xor0;
  wire f_arrdiv16_fs63_not0;
  wire f_arrdiv16_fs63_and0;
  wire f_arrdiv16_fs63_xor1;
  wire f_arrdiv16_fs63_not1;
  wire f_arrdiv16_fs63_and1;
  wire f_arrdiv16_fs63_or0;
  wire f_arrdiv16_mux2to145_and0;
  wire f_arrdiv16_mux2to145_not0;
  wire f_arrdiv16_mux2to145_and1;
  wire f_arrdiv16_mux2to145_xor0;
  wire f_arrdiv16_mux2to146_and0;
  wire f_arrdiv16_mux2to146_not0;
  wire f_arrdiv16_mux2to146_and1;
  wire f_arrdiv16_mux2to146_xor0;
  wire f_arrdiv16_mux2to147_and0;
  wire f_arrdiv16_mux2to147_not0;
  wire f_arrdiv16_mux2to147_and1;
  wire f_arrdiv16_mux2to147_xor0;
  wire f_arrdiv16_mux2to148_and0;
  wire f_arrdiv16_mux2to148_not0;
  wire f_arrdiv16_mux2to148_and1;
  wire f_arrdiv16_mux2to148_xor0;
  wire f_arrdiv16_mux2to149_and0;
  wire f_arrdiv16_mux2to149_not0;
  wire f_arrdiv16_mux2to149_and1;
  wire f_arrdiv16_mux2to149_xor0;
  wire f_arrdiv16_mux2to150_and0;
  wire f_arrdiv16_mux2to150_not0;
  wire f_arrdiv16_mux2to150_and1;
  wire f_arrdiv16_mux2to150_xor0;
  wire f_arrdiv16_mux2to151_and0;
  wire f_arrdiv16_mux2to151_not0;
  wire f_arrdiv16_mux2to151_and1;
  wire f_arrdiv16_mux2to151_xor0;
  wire f_arrdiv16_mux2to152_and0;
  wire f_arrdiv16_mux2to152_not0;
  wire f_arrdiv16_mux2to152_and1;
  wire f_arrdiv16_mux2to152_xor0;
  wire f_arrdiv16_mux2to153_and0;
  wire f_arrdiv16_mux2to153_not0;
  wire f_arrdiv16_mux2to153_and1;
  wire f_arrdiv16_mux2to153_xor0;
  wire f_arrdiv16_mux2to154_and0;
  wire f_arrdiv16_mux2to154_not0;
  wire f_arrdiv16_mux2to154_and1;
  wire f_arrdiv16_mux2to154_xor0;
  wire f_arrdiv16_mux2to155_and0;
  wire f_arrdiv16_mux2to155_not0;
  wire f_arrdiv16_mux2to155_and1;
  wire f_arrdiv16_mux2to155_xor0;
  wire f_arrdiv16_mux2to156_and0;
  wire f_arrdiv16_mux2to156_not0;
  wire f_arrdiv16_mux2to156_and1;
  wire f_arrdiv16_mux2to156_xor0;
  wire f_arrdiv16_mux2to157_and0;
  wire f_arrdiv16_mux2to157_not0;
  wire f_arrdiv16_mux2to157_and1;
  wire f_arrdiv16_mux2to157_xor0;
  wire f_arrdiv16_mux2to158_and0;
  wire f_arrdiv16_mux2to158_not0;
  wire f_arrdiv16_mux2to158_and1;
  wire f_arrdiv16_mux2to158_xor0;
  wire f_arrdiv16_mux2to159_and0;
  wire f_arrdiv16_mux2to159_not0;
  wire f_arrdiv16_mux2to159_and1;
  wire f_arrdiv16_mux2to159_xor0;
  wire f_arrdiv16_not3;
  wire f_arrdiv16_fs64_xor0;
  wire f_arrdiv16_fs64_not0;
  wire f_arrdiv16_fs64_and0;
  wire f_arrdiv16_fs64_not1;
  wire f_arrdiv16_fs65_xor0;
  wire f_arrdiv16_fs65_not0;
  wire f_arrdiv16_fs65_and0;
  wire f_arrdiv16_fs65_xor1;
  wire f_arrdiv16_fs65_not1;
  wire f_arrdiv16_fs65_and1;
  wire f_arrdiv16_fs65_or0;
  wire f_arrdiv16_fs66_xor0;
  wire f_arrdiv16_fs66_not0;
  wire f_arrdiv16_fs66_and0;
  wire f_arrdiv16_fs66_xor1;
  wire f_arrdiv16_fs66_not1;
  wire f_arrdiv16_fs66_and1;
  wire f_arrdiv16_fs66_or0;
  wire f_arrdiv16_fs67_xor0;
  wire f_arrdiv16_fs67_not0;
  wire f_arrdiv16_fs67_and0;
  wire f_arrdiv16_fs67_xor1;
  wire f_arrdiv16_fs67_not1;
  wire f_arrdiv16_fs67_and1;
  wire f_arrdiv16_fs67_or0;
  wire f_arrdiv16_fs68_xor0;
  wire f_arrdiv16_fs68_not0;
  wire f_arrdiv16_fs68_and0;
  wire f_arrdiv16_fs68_xor1;
  wire f_arrdiv16_fs68_not1;
  wire f_arrdiv16_fs68_and1;
  wire f_arrdiv16_fs68_or0;
  wire f_arrdiv16_fs69_xor0;
  wire f_arrdiv16_fs69_not0;
  wire f_arrdiv16_fs69_and0;
  wire f_arrdiv16_fs69_xor1;
  wire f_arrdiv16_fs69_not1;
  wire f_arrdiv16_fs69_and1;
  wire f_arrdiv16_fs69_or0;
  wire f_arrdiv16_fs70_xor0;
  wire f_arrdiv16_fs70_not0;
  wire f_arrdiv16_fs70_and0;
  wire f_arrdiv16_fs70_xor1;
  wire f_arrdiv16_fs70_not1;
  wire f_arrdiv16_fs70_and1;
  wire f_arrdiv16_fs70_or0;
  wire f_arrdiv16_fs71_xor0;
  wire f_arrdiv16_fs71_not0;
  wire f_arrdiv16_fs71_and0;
  wire f_arrdiv16_fs71_xor1;
  wire f_arrdiv16_fs71_not1;
  wire f_arrdiv16_fs71_and1;
  wire f_arrdiv16_fs71_or0;
  wire f_arrdiv16_fs72_xor0;
  wire f_arrdiv16_fs72_not0;
  wire f_arrdiv16_fs72_and0;
  wire f_arrdiv16_fs72_xor1;
  wire f_arrdiv16_fs72_not1;
  wire f_arrdiv16_fs72_and1;
  wire f_arrdiv16_fs72_or0;
  wire f_arrdiv16_fs73_xor0;
  wire f_arrdiv16_fs73_not0;
  wire f_arrdiv16_fs73_and0;
  wire f_arrdiv16_fs73_xor1;
  wire f_arrdiv16_fs73_not1;
  wire f_arrdiv16_fs73_and1;
  wire f_arrdiv16_fs73_or0;
  wire f_arrdiv16_fs74_xor0;
  wire f_arrdiv16_fs74_not0;
  wire f_arrdiv16_fs74_and0;
  wire f_arrdiv16_fs74_xor1;
  wire f_arrdiv16_fs74_not1;
  wire f_arrdiv16_fs74_and1;
  wire f_arrdiv16_fs74_or0;
  wire f_arrdiv16_fs75_xor0;
  wire f_arrdiv16_fs75_not0;
  wire f_arrdiv16_fs75_and0;
  wire f_arrdiv16_fs75_xor1;
  wire f_arrdiv16_fs75_not1;
  wire f_arrdiv16_fs75_and1;
  wire f_arrdiv16_fs75_or0;
  wire f_arrdiv16_fs76_xor0;
  wire f_arrdiv16_fs76_not0;
  wire f_arrdiv16_fs76_and0;
  wire f_arrdiv16_fs76_xor1;
  wire f_arrdiv16_fs76_not1;
  wire f_arrdiv16_fs76_and1;
  wire f_arrdiv16_fs76_or0;
  wire f_arrdiv16_fs77_xor0;
  wire f_arrdiv16_fs77_not0;
  wire f_arrdiv16_fs77_and0;
  wire f_arrdiv16_fs77_xor1;
  wire f_arrdiv16_fs77_not1;
  wire f_arrdiv16_fs77_and1;
  wire f_arrdiv16_fs77_or0;
  wire f_arrdiv16_fs78_xor0;
  wire f_arrdiv16_fs78_not0;
  wire f_arrdiv16_fs78_and0;
  wire f_arrdiv16_fs78_xor1;
  wire f_arrdiv16_fs78_not1;
  wire f_arrdiv16_fs78_and1;
  wire f_arrdiv16_fs78_or0;
  wire f_arrdiv16_fs79_xor0;
  wire f_arrdiv16_fs79_not0;
  wire f_arrdiv16_fs79_and0;
  wire f_arrdiv16_fs79_xor1;
  wire f_arrdiv16_fs79_not1;
  wire f_arrdiv16_fs79_and1;
  wire f_arrdiv16_fs79_or0;
  wire f_arrdiv16_mux2to160_and0;
  wire f_arrdiv16_mux2to160_not0;
  wire f_arrdiv16_mux2to160_and1;
  wire f_arrdiv16_mux2to160_xor0;
  wire f_arrdiv16_mux2to161_and0;
  wire f_arrdiv16_mux2to161_not0;
  wire f_arrdiv16_mux2to161_and1;
  wire f_arrdiv16_mux2to161_xor0;
  wire f_arrdiv16_mux2to162_and0;
  wire f_arrdiv16_mux2to162_not0;
  wire f_arrdiv16_mux2to162_and1;
  wire f_arrdiv16_mux2to162_xor0;
  wire f_arrdiv16_mux2to163_and0;
  wire f_arrdiv16_mux2to163_not0;
  wire f_arrdiv16_mux2to163_and1;
  wire f_arrdiv16_mux2to163_xor0;
  wire f_arrdiv16_mux2to164_and0;
  wire f_arrdiv16_mux2to164_not0;
  wire f_arrdiv16_mux2to164_and1;
  wire f_arrdiv16_mux2to164_xor0;
  wire f_arrdiv16_mux2to165_and0;
  wire f_arrdiv16_mux2to165_not0;
  wire f_arrdiv16_mux2to165_and1;
  wire f_arrdiv16_mux2to165_xor0;
  wire f_arrdiv16_mux2to166_and0;
  wire f_arrdiv16_mux2to166_not0;
  wire f_arrdiv16_mux2to166_and1;
  wire f_arrdiv16_mux2to166_xor0;
  wire f_arrdiv16_mux2to167_and0;
  wire f_arrdiv16_mux2to167_not0;
  wire f_arrdiv16_mux2to167_and1;
  wire f_arrdiv16_mux2to167_xor0;
  wire f_arrdiv16_mux2to168_and0;
  wire f_arrdiv16_mux2to168_not0;
  wire f_arrdiv16_mux2to168_and1;
  wire f_arrdiv16_mux2to168_xor0;
  wire f_arrdiv16_mux2to169_and0;
  wire f_arrdiv16_mux2to169_not0;
  wire f_arrdiv16_mux2to169_and1;
  wire f_arrdiv16_mux2to169_xor0;
  wire f_arrdiv16_mux2to170_and0;
  wire f_arrdiv16_mux2to170_not0;
  wire f_arrdiv16_mux2to170_and1;
  wire f_arrdiv16_mux2to170_xor0;
  wire f_arrdiv16_mux2to171_and0;
  wire f_arrdiv16_mux2to171_not0;
  wire f_arrdiv16_mux2to171_and1;
  wire f_arrdiv16_mux2to171_xor0;
  wire f_arrdiv16_mux2to172_and0;
  wire f_arrdiv16_mux2to172_not0;
  wire f_arrdiv16_mux2to172_and1;
  wire f_arrdiv16_mux2to172_xor0;
  wire f_arrdiv16_mux2to173_and0;
  wire f_arrdiv16_mux2to173_not0;
  wire f_arrdiv16_mux2to173_and1;
  wire f_arrdiv16_mux2to173_xor0;
  wire f_arrdiv16_mux2to174_and0;
  wire f_arrdiv16_mux2to174_not0;
  wire f_arrdiv16_mux2to174_and1;
  wire f_arrdiv16_mux2to174_xor0;
  wire f_arrdiv16_not4;
  wire f_arrdiv16_fs80_xor0;
  wire f_arrdiv16_fs80_not0;
  wire f_arrdiv16_fs80_and0;
  wire f_arrdiv16_fs80_not1;
  wire f_arrdiv16_fs81_xor0;
  wire f_arrdiv16_fs81_not0;
  wire f_arrdiv16_fs81_and0;
  wire f_arrdiv16_fs81_xor1;
  wire f_arrdiv16_fs81_not1;
  wire f_arrdiv16_fs81_and1;
  wire f_arrdiv16_fs81_or0;
  wire f_arrdiv16_fs82_xor0;
  wire f_arrdiv16_fs82_not0;
  wire f_arrdiv16_fs82_and0;
  wire f_arrdiv16_fs82_xor1;
  wire f_arrdiv16_fs82_not1;
  wire f_arrdiv16_fs82_and1;
  wire f_arrdiv16_fs82_or0;
  wire f_arrdiv16_fs83_xor0;
  wire f_arrdiv16_fs83_not0;
  wire f_arrdiv16_fs83_and0;
  wire f_arrdiv16_fs83_xor1;
  wire f_arrdiv16_fs83_not1;
  wire f_arrdiv16_fs83_and1;
  wire f_arrdiv16_fs83_or0;
  wire f_arrdiv16_fs84_xor0;
  wire f_arrdiv16_fs84_not0;
  wire f_arrdiv16_fs84_and0;
  wire f_arrdiv16_fs84_xor1;
  wire f_arrdiv16_fs84_not1;
  wire f_arrdiv16_fs84_and1;
  wire f_arrdiv16_fs84_or0;
  wire f_arrdiv16_fs85_xor0;
  wire f_arrdiv16_fs85_not0;
  wire f_arrdiv16_fs85_and0;
  wire f_arrdiv16_fs85_xor1;
  wire f_arrdiv16_fs85_not1;
  wire f_arrdiv16_fs85_and1;
  wire f_arrdiv16_fs85_or0;
  wire f_arrdiv16_fs86_xor0;
  wire f_arrdiv16_fs86_not0;
  wire f_arrdiv16_fs86_and0;
  wire f_arrdiv16_fs86_xor1;
  wire f_arrdiv16_fs86_not1;
  wire f_arrdiv16_fs86_and1;
  wire f_arrdiv16_fs86_or0;
  wire f_arrdiv16_fs87_xor0;
  wire f_arrdiv16_fs87_not0;
  wire f_arrdiv16_fs87_and0;
  wire f_arrdiv16_fs87_xor1;
  wire f_arrdiv16_fs87_not1;
  wire f_arrdiv16_fs87_and1;
  wire f_arrdiv16_fs87_or0;
  wire f_arrdiv16_fs88_xor0;
  wire f_arrdiv16_fs88_not0;
  wire f_arrdiv16_fs88_and0;
  wire f_arrdiv16_fs88_xor1;
  wire f_arrdiv16_fs88_not1;
  wire f_arrdiv16_fs88_and1;
  wire f_arrdiv16_fs88_or0;
  wire f_arrdiv16_fs89_xor0;
  wire f_arrdiv16_fs89_not0;
  wire f_arrdiv16_fs89_and0;
  wire f_arrdiv16_fs89_xor1;
  wire f_arrdiv16_fs89_not1;
  wire f_arrdiv16_fs89_and1;
  wire f_arrdiv16_fs89_or0;
  wire f_arrdiv16_fs90_xor0;
  wire f_arrdiv16_fs90_not0;
  wire f_arrdiv16_fs90_and0;
  wire f_arrdiv16_fs90_xor1;
  wire f_arrdiv16_fs90_not1;
  wire f_arrdiv16_fs90_and1;
  wire f_arrdiv16_fs90_or0;
  wire f_arrdiv16_fs91_xor0;
  wire f_arrdiv16_fs91_not0;
  wire f_arrdiv16_fs91_and0;
  wire f_arrdiv16_fs91_xor1;
  wire f_arrdiv16_fs91_not1;
  wire f_arrdiv16_fs91_and1;
  wire f_arrdiv16_fs91_or0;
  wire f_arrdiv16_fs92_xor0;
  wire f_arrdiv16_fs92_not0;
  wire f_arrdiv16_fs92_and0;
  wire f_arrdiv16_fs92_xor1;
  wire f_arrdiv16_fs92_not1;
  wire f_arrdiv16_fs92_and1;
  wire f_arrdiv16_fs92_or0;
  wire f_arrdiv16_fs93_xor0;
  wire f_arrdiv16_fs93_not0;
  wire f_arrdiv16_fs93_and0;
  wire f_arrdiv16_fs93_xor1;
  wire f_arrdiv16_fs93_not1;
  wire f_arrdiv16_fs93_and1;
  wire f_arrdiv16_fs93_or0;
  wire f_arrdiv16_fs94_xor0;
  wire f_arrdiv16_fs94_not0;
  wire f_arrdiv16_fs94_and0;
  wire f_arrdiv16_fs94_xor1;
  wire f_arrdiv16_fs94_not1;
  wire f_arrdiv16_fs94_and1;
  wire f_arrdiv16_fs94_or0;
  wire f_arrdiv16_fs95_xor0;
  wire f_arrdiv16_fs95_not0;
  wire f_arrdiv16_fs95_and0;
  wire f_arrdiv16_fs95_xor1;
  wire f_arrdiv16_fs95_not1;
  wire f_arrdiv16_fs95_and1;
  wire f_arrdiv16_fs95_or0;
  wire f_arrdiv16_mux2to175_and0;
  wire f_arrdiv16_mux2to175_not0;
  wire f_arrdiv16_mux2to175_and1;
  wire f_arrdiv16_mux2to175_xor0;
  wire f_arrdiv16_mux2to176_and0;
  wire f_arrdiv16_mux2to176_not0;
  wire f_arrdiv16_mux2to176_and1;
  wire f_arrdiv16_mux2to176_xor0;
  wire f_arrdiv16_mux2to177_and0;
  wire f_arrdiv16_mux2to177_not0;
  wire f_arrdiv16_mux2to177_and1;
  wire f_arrdiv16_mux2to177_xor0;
  wire f_arrdiv16_mux2to178_and0;
  wire f_arrdiv16_mux2to178_not0;
  wire f_arrdiv16_mux2to178_and1;
  wire f_arrdiv16_mux2to178_xor0;
  wire f_arrdiv16_mux2to179_and0;
  wire f_arrdiv16_mux2to179_not0;
  wire f_arrdiv16_mux2to179_and1;
  wire f_arrdiv16_mux2to179_xor0;
  wire f_arrdiv16_mux2to180_and0;
  wire f_arrdiv16_mux2to180_not0;
  wire f_arrdiv16_mux2to180_and1;
  wire f_arrdiv16_mux2to180_xor0;
  wire f_arrdiv16_mux2to181_and0;
  wire f_arrdiv16_mux2to181_not0;
  wire f_arrdiv16_mux2to181_and1;
  wire f_arrdiv16_mux2to181_xor0;
  wire f_arrdiv16_mux2to182_and0;
  wire f_arrdiv16_mux2to182_not0;
  wire f_arrdiv16_mux2to182_and1;
  wire f_arrdiv16_mux2to182_xor0;
  wire f_arrdiv16_mux2to183_and0;
  wire f_arrdiv16_mux2to183_not0;
  wire f_arrdiv16_mux2to183_and1;
  wire f_arrdiv16_mux2to183_xor0;
  wire f_arrdiv16_mux2to184_and0;
  wire f_arrdiv16_mux2to184_not0;
  wire f_arrdiv16_mux2to184_and1;
  wire f_arrdiv16_mux2to184_xor0;
  wire f_arrdiv16_mux2to185_and0;
  wire f_arrdiv16_mux2to185_not0;
  wire f_arrdiv16_mux2to185_and1;
  wire f_arrdiv16_mux2to185_xor0;
  wire f_arrdiv16_mux2to186_and0;
  wire f_arrdiv16_mux2to186_not0;
  wire f_arrdiv16_mux2to186_and1;
  wire f_arrdiv16_mux2to186_xor0;
  wire f_arrdiv16_mux2to187_and0;
  wire f_arrdiv16_mux2to187_not0;
  wire f_arrdiv16_mux2to187_and1;
  wire f_arrdiv16_mux2to187_xor0;
  wire f_arrdiv16_mux2to188_and0;
  wire f_arrdiv16_mux2to188_not0;
  wire f_arrdiv16_mux2to188_and1;
  wire f_arrdiv16_mux2to188_xor0;
  wire f_arrdiv16_mux2to189_and0;
  wire f_arrdiv16_mux2to189_not0;
  wire f_arrdiv16_mux2to189_and1;
  wire f_arrdiv16_mux2to189_xor0;
  wire f_arrdiv16_not5;
  wire f_arrdiv16_fs96_xor0;
  wire f_arrdiv16_fs96_not0;
  wire f_arrdiv16_fs96_and0;
  wire f_arrdiv16_fs96_not1;
  wire f_arrdiv16_fs97_xor0;
  wire f_arrdiv16_fs97_not0;
  wire f_arrdiv16_fs97_and0;
  wire f_arrdiv16_fs97_xor1;
  wire f_arrdiv16_fs97_not1;
  wire f_arrdiv16_fs97_and1;
  wire f_arrdiv16_fs97_or0;
  wire f_arrdiv16_fs98_xor0;
  wire f_arrdiv16_fs98_not0;
  wire f_arrdiv16_fs98_and0;
  wire f_arrdiv16_fs98_xor1;
  wire f_arrdiv16_fs98_not1;
  wire f_arrdiv16_fs98_and1;
  wire f_arrdiv16_fs98_or0;
  wire f_arrdiv16_fs99_xor0;
  wire f_arrdiv16_fs99_not0;
  wire f_arrdiv16_fs99_and0;
  wire f_arrdiv16_fs99_xor1;
  wire f_arrdiv16_fs99_not1;
  wire f_arrdiv16_fs99_and1;
  wire f_arrdiv16_fs99_or0;
  wire f_arrdiv16_fs100_xor0;
  wire f_arrdiv16_fs100_not0;
  wire f_arrdiv16_fs100_and0;
  wire f_arrdiv16_fs100_xor1;
  wire f_arrdiv16_fs100_not1;
  wire f_arrdiv16_fs100_and1;
  wire f_arrdiv16_fs100_or0;
  wire f_arrdiv16_fs101_xor0;
  wire f_arrdiv16_fs101_not0;
  wire f_arrdiv16_fs101_and0;
  wire f_arrdiv16_fs101_xor1;
  wire f_arrdiv16_fs101_not1;
  wire f_arrdiv16_fs101_and1;
  wire f_arrdiv16_fs101_or0;
  wire f_arrdiv16_fs102_xor0;
  wire f_arrdiv16_fs102_not0;
  wire f_arrdiv16_fs102_and0;
  wire f_arrdiv16_fs102_xor1;
  wire f_arrdiv16_fs102_not1;
  wire f_arrdiv16_fs102_and1;
  wire f_arrdiv16_fs102_or0;
  wire f_arrdiv16_fs103_xor0;
  wire f_arrdiv16_fs103_not0;
  wire f_arrdiv16_fs103_and0;
  wire f_arrdiv16_fs103_xor1;
  wire f_arrdiv16_fs103_not1;
  wire f_arrdiv16_fs103_and1;
  wire f_arrdiv16_fs103_or0;
  wire f_arrdiv16_fs104_xor0;
  wire f_arrdiv16_fs104_not0;
  wire f_arrdiv16_fs104_and0;
  wire f_arrdiv16_fs104_xor1;
  wire f_arrdiv16_fs104_not1;
  wire f_arrdiv16_fs104_and1;
  wire f_arrdiv16_fs104_or0;
  wire f_arrdiv16_fs105_xor0;
  wire f_arrdiv16_fs105_not0;
  wire f_arrdiv16_fs105_and0;
  wire f_arrdiv16_fs105_xor1;
  wire f_arrdiv16_fs105_not1;
  wire f_arrdiv16_fs105_and1;
  wire f_arrdiv16_fs105_or0;
  wire f_arrdiv16_fs106_xor0;
  wire f_arrdiv16_fs106_not0;
  wire f_arrdiv16_fs106_and0;
  wire f_arrdiv16_fs106_xor1;
  wire f_arrdiv16_fs106_not1;
  wire f_arrdiv16_fs106_and1;
  wire f_arrdiv16_fs106_or0;
  wire f_arrdiv16_fs107_xor0;
  wire f_arrdiv16_fs107_not0;
  wire f_arrdiv16_fs107_and0;
  wire f_arrdiv16_fs107_xor1;
  wire f_arrdiv16_fs107_not1;
  wire f_arrdiv16_fs107_and1;
  wire f_arrdiv16_fs107_or0;
  wire f_arrdiv16_fs108_xor0;
  wire f_arrdiv16_fs108_not0;
  wire f_arrdiv16_fs108_and0;
  wire f_arrdiv16_fs108_xor1;
  wire f_arrdiv16_fs108_not1;
  wire f_arrdiv16_fs108_and1;
  wire f_arrdiv16_fs108_or0;
  wire f_arrdiv16_fs109_xor0;
  wire f_arrdiv16_fs109_not0;
  wire f_arrdiv16_fs109_and0;
  wire f_arrdiv16_fs109_xor1;
  wire f_arrdiv16_fs109_not1;
  wire f_arrdiv16_fs109_and1;
  wire f_arrdiv16_fs109_or0;
  wire f_arrdiv16_fs110_xor0;
  wire f_arrdiv16_fs110_not0;
  wire f_arrdiv16_fs110_and0;
  wire f_arrdiv16_fs110_xor1;
  wire f_arrdiv16_fs110_not1;
  wire f_arrdiv16_fs110_and1;
  wire f_arrdiv16_fs110_or0;
  wire f_arrdiv16_fs111_xor0;
  wire f_arrdiv16_fs111_not0;
  wire f_arrdiv16_fs111_and0;
  wire f_arrdiv16_fs111_xor1;
  wire f_arrdiv16_fs111_not1;
  wire f_arrdiv16_fs111_and1;
  wire f_arrdiv16_fs111_or0;
  wire f_arrdiv16_mux2to190_and0;
  wire f_arrdiv16_mux2to190_not0;
  wire f_arrdiv16_mux2to190_and1;
  wire f_arrdiv16_mux2to190_xor0;
  wire f_arrdiv16_mux2to191_and0;
  wire f_arrdiv16_mux2to191_not0;
  wire f_arrdiv16_mux2to191_and1;
  wire f_arrdiv16_mux2to191_xor0;
  wire f_arrdiv16_mux2to192_and0;
  wire f_arrdiv16_mux2to192_not0;
  wire f_arrdiv16_mux2to192_and1;
  wire f_arrdiv16_mux2to192_xor0;
  wire f_arrdiv16_mux2to193_and0;
  wire f_arrdiv16_mux2to193_not0;
  wire f_arrdiv16_mux2to193_and1;
  wire f_arrdiv16_mux2to193_xor0;
  wire f_arrdiv16_mux2to194_and0;
  wire f_arrdiv16_mux2to194_not0;
  wire f_arrdiv16_mux2to194_and1;
  wire f_arrdiv16_mux2to194_xor0;
  wire f_arrdiv16_mux2to195_and0;
  wire f_arrdiv16_mux2to195_not0;
  wire f_arrdiv16_mux2to195_and1;
  wire f_arrdiv16_mux2to195_xor0;
  wire f_arrdiv16_mux2to196_and0;
  wire f_arrdiv16_mux2to196_not0;
  wire f_arrdiv16_mux2to196_and1;
  wire f_arrdiv16_mux2to196_xor0;
  wire f_arrdiv16_mux2to197_and0;
  wire f_arrdiv16_mux2to197_not0;
  wire f_arrdiv16_mux2to197_and1;
  wire f_arrdiv16_mux2to197_xor0;
  wire f_arrdiv16_mux2to198_and0;
  wire f_arrdiv16_mux2to198_not0;
  wire f_arrdiv16_mux2to198_and1;
  wire f_arrdiv16_mux2to198_xor0;
  wire f_arrdiv16_mux2to199_and0;
  wire f_arrdiv16_mux2to199_not0;
  wire f_arrdiv16_mux2to199_and1;
  wire f_arrdiv16_mux2to199_xor0;
  wire f_arrdiv16_mux2to1100_and0;
  wire f_arrdiv16_mux2to1100_not0;
  wire f_arrdiv16_mux2to1100_and1;
  wire f_arrdiv16_mux2to1100_xor0;
  wire f_arrdiv16_mux2to1101_and0;
  wire f_arrdiv16_mux2to1101_not0;
  wire f_arrdiv16_mux2to1101_and1;
  wire f_arrdiv16_mux2to1101_xor0;
  wire f_arrdiv16_mux2to1102_and0;
  wire f_arrdiv16_mux2to1102_not0;
  wire f_arrdiv16_mux2to1102_and1;
  wire f_arrdiv16_mux2to1102_xor0;
  wire f_arrdiv16_mux2to1103_and0;
  wire f_arrdiv16_mux2to1103_not0;
  wire f_arrdiv16_mux2to1103_and1;
  wire f_arrdiv16_mux2to1103_xor0;
  wire f_arrdiv16_mux2to1104_and0;
  wire f_arrdiv16_mux2to1104_not0;
  wire f_arrdiv16_mux2to1104_and1;
  wire f_arrdiv16_mux2to1104_xor0;
  wire f_arrdiv16_not6;
  wire f_arrdiv16_fs112_xor0;
  wire f_arrdiv16_fs112_not0;
  wire f_arrdiv16_fs112_and0;
  wire f_arrdiv16_fs112_not1;
  wire f_arrdiv16_fs113_xor0;
  wire f_arrdiv16_fs113_not0;
  wire f_arrdiv16_fs113_and0;
  wire f_arrdiv16_fs113_xor1;
  wire f_arrdiv16_fs113_not1;
  wire f_arrdiv16_fs113_and1;
  wire f_arrdiv16_fs113_or0;
  wire f_arrdiv16_fs114_xor0;
  wire f_arrdiv16_fs114_not0;
  wire f_arrdiv16_fs114_and0;
  wire f_arrdiv16_fs114_xor1;
  wire f_arrdiv16_fs114_not1;
  wire f_arrdiv16_fs114_and1;
  wire f_arrdiv16_fs114_or0;
  wire f_arrdiv16_fs115_xor0;
  wire f_arrdiv16_fs115_not0;
  wire f_arrdiv16_fs115_and0;
  wire f_arrdiv16_fs115_xor1;
  wire f_arrdiv16_fs115_not1;
  wire f_arrdiv16_fs115_and1;
  wire f_arrdiv16_fs115_or0;
  wire f_arrdiv16_fs116_xor0;
  wire f_arrdiv16_fs116_not0;
  wire f_arrdiv16_fs116_and0;
  wire f_arrdiv16_fs116_xor1;
  wire f_arrdiv16_fs116_not1;
  wire f_arrdiv16_fs116_and1;
  wire f_arrdiv16_fs116_or0;
  wire f_arrdiv16_fs117_xor0;
  wire f_arrdiv16_fs117_not0;
  wire f_arrdiv16_fs117_and0;
  wire f_arrdiv16_fs117_xor1;
  wire f_arrdiv16_fs117_not1;
  wire f_arrdiv16_fs117_and1;
  wire f_arrdiv16_fs117_or0;
  wire f_arrdiv16_fs118_xor0;
  wire f_arrdiv16_fs118_not0;
  wire f_arrdiv16_fs118_and0;
  wire f_arrdiv16_fs118_xor1;
  wire f_arrdiv16_fs118_not1;
  wire f_arrdiv16_fs118_and1;
  wire f_arrdiv16_fs118_or0;
  wire f_arrdiv16_fs119_xor0;
  wire f_arrdiv16_fs119_not0;
  wire f_arrdiv16_fs119_and0;
  wire f_arrdiv16_fs119_xor1;
  wire f_arrdiv16_fs119_not1;
  wire f_arrdiv16_fs119_and1;
  wire f_arrdiv16_fs119_or0;
  wire f_arrdiv16_fs120_xor0;
  wire f_arrdiv16_fs120_not0;
  wire f_arrdiv16_fs120_and0;
  wire f_arrdiv16_fs120_xor1;
  wire f_arrdiv16_fs120_not1;
  wire f_arrdiv16_fs120_and1;
  wire f_arrdiv16_fs120_or0;
  wire f_arrdiv16_fs121_xor0;
  wire f_arrdiv16_fs121_not0;
  wire f_arrdiv16_fs121_and0;
  wire f_arrdiv16_fs121_xor1;
  wire f_arrdiv16_fs121_not1;
  wire f_arrdiv16_fs121_and1;
  wire f_arrdiv16_fs121_or0;
  wire f_arrdiv16_fs122_xor0;
  wire f_arrdiv16_fs122_not0;
  wire f_arrdiv16_fs122_and0;
  wire f_arrdiv16_fs122_xor1;
  wire f_arrdiv16_fs122_not1;
  wire f_arrdiv16_fs122_and1;
  wire f_arrdiv16_fs122_or0;
  wire f_arrdiv16_fs123_xor0;
  wire f_arrdiv16_fs123_not0;
  wire f_arrdiv16_fs123_and0;
  wire f_arrdiv16_fs123_xor1;
  wire f_arrdiv16_fs123_not1;
  wire f_arrdiv16_fs123_and1;
  wire f_arrdiv16_fs123_or0;
  wire f_arrdiv16_fs124_xor0;
  wire f_arrdiv16_fs124_not0;
  wire f_arrdiv16_fs124_and0;
  wire f_arrdiv16_fs124_xor1;
  wire f_arrdiv16_fs124_not1;
  wire f_arrdiv16_fs124_and1;
  wire f_arrdiv16_fs124_or0;
  wire f_arrdiv16_fs125_xor0;
  wire f_arrdiv16_fs125_not0;
  wire f_arrdiv16_fs125_and0;
  wire f_arrdiv16_fs125_xor1;
  wire f_arrdiv16_fs125_not1;
  wire f_arrdiv16_fs125_and1;
  wire f_arrdiv16_fs125_or0;
  wire f_arrdiv16_fs126_xor0;
  wire f_arrdiv16_fs126_not0;
  wire f_arrdiv16_fs126_and0;
  wire f_arrdiv16_fs126_xor1;
  wire f_arrdiv16_fs126_not1;
  wire f_arrdiv16_fs126_and1;
  wire f_arrdiv16_fs126_or0;
  wire f_arrdiv16_fs127_xor0;
  wire f_arrdiv16_fs127_not0;
  wire f_arrdiv16_fs127_and0;
  wire f_arrdiv16_fs127_xor1;
  wire f_arrdiv16_fs127_not1;
  wire f_arrdiv16_fs127_and1;
  wire f_arrdiv16_fs127_or0;
  wire f_arrdiv16_mux2to1105_and0;
  wire f_arrdiv16_mux2to1105_not0;
  wire f_arrdiv16_mux2to1105_and1;
  wire f_arrdiv16_mux2to1105_xor0;
  wire f_arrdiv16_mux2to1106_and0;
  wire f_arrdiv16_mux2to1106_not0;
  wire f_arrdiv16_mux2to1106_and1;
  wire f_arrdiv16_mux2to1106_xor0;
  wire f_arrdiv16_mux2to1107_and0;
  wire f_arrdiv16_mux2to1107_not0;
  wire f_arrdiv16_mux2to1107_and1;
  wire f_arrdiv16_mux2to1107_xor0;
  wire f_arrdiv16_mux2to1108_and0;
  wire f_arrdiv16_mux2to1108_not0;
  wire f_arrdiv16_mux2to1108_and1;
  wire f_arrdiv16_mux2to1108_xor0;
  wire f_arrdiv16_mux2to1109_and0;
  wire f_arrdiv16_mux2to1109_not0;
  wire f_arrdiv16_mux2to1109_and1;
  wire f_arrdiv16_mux2to1109_xor0;
  wire f_arrdiv16_mux2to1110_and0;
  wire f_arrdiv16_mux2to1110_not0;
  wire f_arrdiv16_mux2to1110_and1;
  wire f_arrdiv16_mux2to1110_xor0;
  wire f_arrdiv16_mux2to1111_and0;
  wire f_arrdiv16_mux2to1111_not0;
  wire f_arrdiv16_mux2to1111_and1;
  wire f_arrdiv16_mux2to1111_xor0;
  wire f_arrdiv16_mux2to1112_and0;
  wire f_arrdiv16_mux2to1112_not0;
  wire f_arrdiv16_mux2to1112_and1;
  wire f_arrdiv16_mux2to1112_xor0;
  wire f_arrdiv16_mux2to1113_and0;
  wire f_arrdiv16_mux2to1113_not0;
  wire f_arrdiv16_mux2to1113_and1;
  wire f_arrdiv16_mux2to1113_xor0;
  wire f_arrdiv16_mux2to1114_and0;
  wire f_arrdiv16_mux2to1114_not0;
  wire f_arrdiv16_mux2to1114_and1;
  wire f_arrdiv16_mux2to1114_xor0;
  wire f_arrdiv16_mux2to1115_and0;
  wire f_arrdiv16_mux2to1115_not0;
  wire f_arrdiv16_mux2to1115_and1;
  wire f_arrdiv16_mux2to1115_xor0;
  wire f_arrdiv16_mux2to1116_and0;
  wire f_arrdiv16_mux2to1116_not0;
  wire f_arrdiv16_mux2to1116_and1;
  wire f_arrdiv16_mux2to1116_xor0;
  wire f_arrdiv16_mux2to1117_and0;
  wire f_arrdiv16_mux2to1117_not0;
  wire f_arrdiv16_mux2to1117_and1;
  wire f_arrdiv16_mux2to1117_xor0;
  wire f_arrdiv16_mux2to1118_and0;
  wire f_arrdiv16_mux2to1118_not0;
  wire f_arrdiv16_mux2to1118_and1;
  wire f_arrdiv16_mux2to1118_xor0;
  wire f_arrdiv16_mux2to1119_and0;
  wire f_arrdiv16_mux2to1119_not0;
  wire f_arrdiv16_mux2to1119_and1;
  wire f_arrdiv16_mux2to1119_xor0;
  wire f_arrdiv16_not7;
  wire f_arrdiv16_fs128_xor0;
  wire f_arrdiv16_fs128_not0;
  wire f_arrdiv16_fs128_and0;
  wire f_arrdiv16_fs128_not1;
  wire f_arrdiv16_fs129_xor0;
  wire f_arrdiv16_fs129_not0;
  wire f_arrdiv16_fs129_and0;
  wire f_arrdiv16_fs129_xor1;
  wire f_arrdiv16_fs129_not1;
  wire f_arrdiv16_fs129_and1;
  wire f_arrdiv16_fs129_or0;
  wire f_arrdiv16_fs130_xor0;
  wire f_arrdiv16_fs130_not0;
  wire f_arrdiv16_fs130_and0;
  wire f_arrdiv16_fs130_xor1;
  wire f_arrdiv16_fs130_not1;
  wire f_arrdiv16_fs130_and1;
  wire f_arrdiv16_fs130_or0;
  wire f_arrdiv16_fs131_xor0;
  wire f_arrdiv16_fs131_not0;
  wire f_arrdiv16_fs131_and0;
  wire f_arrdiv16_fs131_xor1;
  wire f_arrdiv16_fs131_not1;
  wire f_arrdiv16_fs131_and1;
  wire f_arrdiv16_fs131_or0;
  wire f_arrdiv16_fs132_xor0;
  wire f_arrdiv16_fs132_not0;
  wire f_arrdiv16_fs132_and0;
  wire f_arrdiv16_fs132_xor1;
  wire f_arrdiv16_fs132_not1;
  wire f_arrdiv16_fs132_and1;
  wire f_arrdiv16_fs132_or0;
  wire f_arrdiv16_fs133_xor0;
  wire f_arrdiv16_fs133_not0;
  wire f_arrdiv16_fs133_and0;
  wire f_arrdiv16_fs133_xor1;
  wire f_arrdiv16_fs133_not1;
  wire f_arrdiv16_fs133_and1;
  wire f_arrdiv16_fs133_or0;
  wire f_arrdiv16_fs134_xor0;
  wire f_arrdiv16_fs134_not0;
  wire f_arrdiv16_fs134_and0;
  wire f_arrdiv16_fs134_xor1;
  wire f_arrdiv16_fs134_not1;
  wire f_arrdiv16_fs134_and1;
  wire f_arrdiv16_fs134_or0;
  wire f_arrdiv16_fs135_xor0;
  wire f_arrdiv16_fs135_not0;
  wire f_arrdiv16_fs135_and0;
  wire f_arrdiv16_fs135_xor1;
  wire f_arrdiv16_fs135_not1;
  wire f_arrdiv16_fs135_and1;
  wire f_arrdiv16_fs135_or0;
  wire f_arrdiv16_fs136_xor0;
  wire f_arrdiv16_fs136_not0;
  wire f_arrdiv16_fs136_and0;
  wire f_arrdiv16_fs136_xor1;
  wire f_arrdiv16_fs136_not1;
  wire f_arrdiv16_fs136_and1;
  wire f_arrdiv16_fs136_or0;
  wire f_arrdiv16_fs137_xor0;
  wire f_arrdiv16_fs137_not0;
  wire f_arrdiv16_fs137_and0;
  wire f_arrdiv16_fs137_xor1;
  wire f_arrdiv16_fs137_not1;
  wire f_arrdiv16_fs137_and1;
  wire f_arrdiv16_fs137_or0;
  wire f_arrdiv16_fs138_xor0;
  wire f_arrdiv16_fs138_not0;
  wire f_arrdiv16_fs138_and0;
  wire f_arrdiv16_fs138_xor1;
  wire f_arrdiv16_fs138_not1;
  wire f_arrdiv16_fs138_and1;
  wire f_arrdiv16_fs138_or0;
  wire f_arrdiv16_fs139_xor0;
  wire f_arrdiv16_fs139_not0;
  wire f_arrdiv16_fs139_and0;
  wire f_arrdiv16_fs139_xor1;
  wire f_arrdiv16_fs139_not1;
  wire f_arrdiv16_fs139_and1;
  wire f_arrdiv16_fs139_or0;
  wire f_arrdiv16_fs140_xor0;
  wire f_arrdiv16_fs140_not0;
  wire f_arrdiv16_fs140_and0;
  wire f_arrdiv16_fs140_xor1;
  wire f_arrdiv16_fs140_not1;
  wire f_arrdiv16_fs140_and1;
  wire f_arrdiv16_fs140_or0;
  wire f_arrdiv16_fs141_xor0;
  wire f_arrdiv16_fs141_not0;
  wire f_arrdiv16_fs141_and0;
  wire f_arrdiv16_fs141_xor1;
  wire f_arrdiv16_fs141_not1;
  wire f_arrdiv16_fs141_and1;
  wire f_arrdiv16_fs141_or0;
  wire f_arrdiv16_fs142_xor0;
  wire f_arrdiv16_fs142_not0;
  wire f_arrdiv16_fs142_and0;
  wire f_arrdiv16_fs142_xor1;
  wire f_arrdiv16_fs142_not1;
  wire f_arrdiv16_fs142_and1;
  wire f_arrdiv16_fs142_or0;
  wire f_arrdiv16_fs143_xor0;
  wire f_arrdiv16_fs143_not0;
  wire f_arrdiv16_fs143_and0;
  wire f_arrdiv16_fs143_xor1;
  wire f_arrdiv16_fs143_not1;
  wire f_arrdiv16_fs143_and1;
  wire f_arrdiv16_fs143_or0;
  wire f_arrdiv16_mux2to1120_and0;
  wire f_arrdiv16_mux2to1120_not0;
  wire f_arrdiv16_mux2to1120_and1;
  wire f_arrdiv16_mux2to1120_xor0;
  wire f_arrdiv16_mux2to1121_and0;
  wire f_arrdiv16_mux2to1121_not0;
  wire f_arrdiv16_mux2to1121_and1;
  wire f_arrdiv16_mux2to1121_xor0;
  wire f_arrdiv16_mux2to1122_and0;
  wire f_arrdiv16_mux2to1122_not0;
  wire f_arrdiv16_mux2to1122_and1;
  wire f_arrdiv16_mux2to1122_xor0;
  wire f_arrdiv16_mux2to1123_and0;
  wire f_arrdiv16_mux2to1123_not0;
  wire f_arrdiv16_mux2to1123_and1;
  wire f_arrdiv16_mux2to1123_xor0;
  wire f_arrdiv16_mux2to1124_and0;
  wire f_arrdiv16_mux2to1124_not0;
  wire f_arrdiv16_mux2to1124_and1;
  wire f_arrdiv16_mux2to1124_xor0;
  wire f_arrdiv16_mux2to1125_and0;
  wire f_arrdiv16_mux2to1125_not0;
  wire f_arrdiv16_mux2to1125_and1;
  wire f_arrdiv16_mux2to1125_xor0;
  wire f_arrdiv16_mux2to1126_and0;
  wire f_arrdiv16_mux2to1126_not0;
  wire f_arrdiv16_mux2to1126_and1;
  wire f_arrdiv16_mux2to1126_xor0;
  wire f_arrdiv16_mux2to1127_and0;
  wire f_arrdiv16_mux2to1127_not0;
  wire f_arrdiv16_mux2to1127_and1;
  wire f_arrdiv16_mux2to1127_xor0;
  wire f_arrdiv16_mux2to1128_and0;
  wire f_arrdiv16_mux2to1128_not0;
  wire f_arrdiv16_mux2to1128_and1;
  wire f_arrdiv16_mux2to1128_xor0;
  wire f_arrdiv16_mux2to1129_and0;
  wire f_arrdiv16_mux2to1129_not0;
  wire f_arrdiv16_mux2to1129_and1;
  wire f_arrdiv16_mux2to1129_xor0;
  wire f_arrdiv16_mux2to1130_and0;
  wire f_arrdiv16_mux2to1130_not0;
  wire f_arrdiv16_mux2to1130_and1;
  wire f_arrdiv16_mux2to1130_xor0;
  wire f_arrdiv16_mux2to1131_and0;
  wire f_arrdiv16_mux2to1131_not0;
  wire f_arrdiv16_mux2to1131_and1;
  wire f_arrdiv16_mux2to1131_xor0;
  wire f_arrdiv16_mux2to1132_and0;
  wire f_arrdiv16_mux2to1132_not0;
  wire f_arrdiv16_mux2to1132_and1;
  wire f_arrdiv16_mux2to1132_xor0;
  wire f_arrdiv16_mux2to1133_and0;
  wire f_arrdiv16_mux2to1133_not0;
  wire f_arrdiv16_mux2to1133_and1;
  wire f_arrdiv16_mux2to1133_xor0;
  wire f_arrdiv16_mux2to1134_and0;
  wire f_arrdiv16_mux2to1134_not0;
  wire f_arrdiv16_mux2to1134_and1;
  wire f_arrdiv16_mux2to1134_xor0;
  wire f_arrdiv16_not8;
  wire f_arrdiv16_fs144_xor0;
  wire f_arrdiv16_fs144_not0;
  wire f_arrdiv16_fs144_and0;
  wire f_arrdiv16_fs144_not1;
  wire f_arrdiv16_fs145_xor0;
  wire f_arrdiv16_fs145_not0;
  wire f_arrdiv16_fs145_and0;
  wire f_arrdiv16_fs145_xor1;
  wire f_arrdiv16_fs145_not1;
  wire f_arrdiv16_fs145_and1;
  wire f_arrdiv16_fs145_or0;
  wire f_arrdiv16_fs146_xor0;
  wire f_arrdiv16_fs146_not0;
  wire f_arrdiv16_fs146_and0;
  wire f_arrdiv16_fs146_xor1;
  wire f_arrdiv16_fs146_not1;
  wire f_arrdiv16_fs146_and1;
  wire f_arrdiv16_fs146_or0;
  wire f_arrdiv16_fs147_xor0;
  wire f_arrdiv16_fs147_not0;
  wire f_arrdiv16_fs147_and0;
  wire f_arrdiv16_fs147_xor1;
  wire f_arrdiv16_fs147_not1;
  wire f_arrdiv16_fs147_and1;
  wire f_arrdiv16_fs147_or0;
  wire f_arrdiv16_fs148_xor0;
  wire f_arrdiv16_fs148_not0;
  wire f_arrdiv16_fs148_and0;
  wire f_arrdiv16_fs148_xor1;
  wire f_arrdiv16_fs148_not1;
  wire f_arrdiv16_fs148_and1;
  wire f_arrdiv16_fs148_or0;
  wire f_arrdiv16_fs149_xor0;
  wire f_arrdiv16_fs149_not0;
  wire f_arrdiv16_fs149_and0;
  wire f_arrdiv16_fs149_xor1;
  wire f_arrdiv16_fs149_not1;
  wire f_arrdiv16_fs149_and1;
  wire f_arrdiv16_fs149_or0;
  wire f_arrdiv16_fs150_xor0;
  wire f_arrdiv16_fs150_not0;
  wire f_arrdiv16_fs150_and0;
  wire f_arrdiv16_fs150_xor1;
  wire f_arrdiv16_fs150_not1;
  wire f_arrdiv16_fs150_and1;
  wire f_arrdiv16_fs150_or0;
  wire f_arrdiv16_fs151_xor0;
  wire f_arrdiv16_fs151_not0;
  wire f_arrdiv16_fs151_and0;
  wire f_arrdiv16_fs151_xor1;
  wire f_arrdiv16_fs151_not1;
  wire f_arrdiv16_fs151_and1;
  wire f_arrdiv16_fs151_or0;
  wire f_arrdiv16_fs152_xor0;
  wire f_arrdiv16_fs152_not0;
  wire f_arrdiv16_fs152_and0;
  wire f_arrdiv16_fs152_xor1;
  wire f_arrdiv16_fs152_not1;
  wire f_arrdiv16_fs152_and1;
  wire f_arrdiv16_fs152_or0;
  wire f_arrdiv16_fs153_xor0;
  wire f_arrdiv16_fs153_not0;
  wire f_arrdiv16_fs153_and0;
  wire f_arrdiv16_fs153_xor1;
  wire f_arrdiv16_fs153_not1;
  wire f_arrdiv16_fs153_and1;
  wire f_arrdiv16_fs153_or0;
  wire f_arrdiv16_fs154_xor0;
  wire f_arrdiv16_fs154_not0;
  wire f_arrdiv16_fs154_and0;
  wire f_arrdiv16_fs154_xor1;
  wire f_arrdiv16_fs154_not1;
  wire f_arrdiv16_fs154_and1;
  wire f_arrdiv16_fs154_or0;
  wire f_arrdiv16_fs155_xor0;
  wire f_arrdiv16_fs155_not0;
  wire f_arrdiv16_fs155_and0;
  wire f_arrdiv16_fs155_xor1;
  wire f_arrdiv16_fs155_not1;
  wire f_arrdiv16_fs155_and1;
  wire f_arrdiv16_fs155_or0;
  wire f_arrdiv16_fs156_xor0;
  wire f_arrdiv16_fs156_not0;
  wire f_arrdiv16_fs156_and0;
  wire f_arrdiv16_fs156_xor1;
  wire f_arrdiv16_fs156_not1;
  wire f_arrdiv16_fs156_and1;
  wire f_arrdiv16_fs156_or0;
  wire f_arrdiv16_fs157_xor0;
  wire f_arrdiv16_fs157_not0;
  wire f_arrdiv16_fs157_and0;
  wire f_arrdiv16_fs157_xor1;
  wire f_arrdiv16_fs157_not1;
  wire f_arrdiv16_fs157_and1;
  wire f_arrdiv16_fs157_or0;
  wire f_arrdiv16_fs158_xor0;
  wire f_arrdiv16_fs158_not0;
  wire f_arrdiv16_fs158_and0;
  wire f_arrdiv16_fs158_xor1;
  wire f_arrdiv16_fs158_not1;
  wire f_arrdiv16_fs158_and1;
  wire f_arrdiv16_fs158_or0;
  wire f_arrdiv16_fs159_xor0;
  wire f_arrdiv16_fs159_not0;
  wire f_arrdiv16_fs159_and0;
  wire f_arrdiv16_fs159_xor1;
  wire f_arrdiv16_fs159_not1;
  wire f_arrdiv16_fs159_and1;
  wire f_arrdiv16_fs159_or0;
  wire f_arrdiv16_mux2to1135_and0;
  wire f_arrdiv16_mux2to1135_not0;
  wire f_arrdiv16_mux2to1135_and1;
  wire f_arrdiv16_mux2to1135_xor0;
  wire f_arrdiv16_mux2to1136_and0;
  wire f_arrdiv16_mux2to1136_not0;
  wire f_arrdiv16_mux2to1136_and1;
  wire f_arrdiv16_mux2to1136_xor0;
  wire f_arrdiv16_mux2to1137_and0;
  wire f_arrdiv16_mux2to1137_not0;
  wire f_arrdiv16_mux2to1137_and1;
  wire f_arrdiv16_mux2to1137_xor0;
  wire f_arrdiv16_mux2to1138_and0;
  wire f_arrdiv16_mux2to1138_not0;
  wire f_arrdiv16_mux2to1138_and1;
  wire f_arrdiv16_mux2to1138_xor0;
  wire f_arrdiv16_mux2to1139_and0;
  wire f_arrdiv16_mux2to1139_not0;
  wire f_arrdiv16_mux2to1139_and1;
  wire f_arrdiv16_mux2to1139_xor0;
  wire f_arrdiv16_mux2to1140_and0;
  wire f_arrdiv16_mux2to1140_not0;
  wire f_arrdiv16_mux2to1140_and1;
  wire f_arrdiv16_mux2to1140_xor0;
  wire f_arrdiv16_mux2to1141_and0;
  wire f_arrdiv16_mux2to1141_not0;
  wire f_arrdiv16_mux2to1141_and1;
  wire f_arrdiv16_mux2to1141_xor0;
  wire f_arrdiv16_mux2to1142_and0;
  wire f_arrdiv16_mux2to1142_not0;
  wire f_arrdiv16_mux2to1142_and1;
  wire f_arrdiv16_mux2to1142_xor0;
  wire f_arrdiv16_mux2to1143_and0;
  wire f_arrdiv16_mux2to1143_not0;
  wire f_arrdiv16_mux2to1143_and1;
  wire f_arrdiv16_mux2to1143_xor0;
  wire f_arrdiv16_mux2to1144_and0;
  wire f_arrdiv16_mux2to1144_not0;
  wire f_arrdiv16_mux2to1144_and1;
  wire f_arrdiv16_mux2to1144_xor0;
  wire f_arrdiv16_mux2to1145_and0;
  wire f_arrdiv16_mux2to1145_not0;
  wire f_arrdiv16_mux2to1145_and1;
  wire f_arrdiv16_mux2to1145_xor0;
  wire f_arrdiv16_mux2to1146_and0;
  wire f_arrdiv16_mux2to1146_not0;
  wire f_arrdiv16_mux2to1146_and1;
  wire f_arrdiv16_mux2to1146_xor0;
  wire f_arrdiv16_mux2to1147_and0;
  wire f_arrdiv16_mux2to1147_not0;
  wire f_arrdiv16_mux2to1147_and1;
  wire f_arrdiv16_mux2to1147_xor0;
  wire f_arrdiv16_mux2to1148_and0;
  wire f_arrdiv16_mux2to1148_not0;
  wire f_arrdiv16_mux2to1148_and1;
  wire f_arrdiv16_mux2to1148_xor0;
  wire f_arrdiv16_mux2to1149_and0;
  wire f_arrdiv16_mux2to1149_not0;
  wire f_arrdiv16_mux2to1149_and1;
  wire f_arrdiv16_mux2to1149_xor0;
  wire f_arrdiv16_not9;
  wire f_arrdiv16_fs160_xor0;
  wire f_arrdiv16_fs160_not0;
  wire f_arrdiv16_fs160_and0;
  wire f_arrdiv16_fs160_not1;
  wire f_arrdiv16_fs161_xor0;
  wire f_arrdiv16_fs161_not0;
  wire f_arrdiv16_fs161_and0;
  wire f_arrdiv16_fs161_xor1;
  wire f_arrdiv16_fs161_not1;
  wire f_arrdiv16_fs161_and1;
  wire f_arrdiv16_fs161_or0;
  wire f_arrdiv16_fs162_xor0;
  wire f_arrdiv16_fs162_not0;
  wire f_arrdiv16_fs162_and0;
  wire f_arrdiv16_fs162_xor1;
  wire f_arrdiv16_fs162_not1;
  wire f_arrdiv16_fs162_and1;
  wire f_arrdiv16_fs162_or0;
  wire f_arrdiv16_fs163_xor0;
  wire f_arrdiv16_fs163_not0;
  wire f_arrdiv16_fs163_and0;
  wire f_arrdiv16_fs163_xor1;
  wire f_arrdiv16_fs163_not1;
  wire f_arrdiv16_fs163_and1;
  wire f_arrdiv16_fs163_or0;
  wire f_arrdiv16_fs164_xor0;
  wire f_arrdiv16_fs164_not0;
  wire f_arrdiv16_fs164_and0;
  wire f_arrdiv16_fs164_xor1;
  wire f_arrdiv16_fs164_not1;
  wire f_arrdiv16_fs164_and1;
  wire f_arrdiv16_fs164_or0;
  wire f_arrdiv16_fs165_xor0;
  wire f_arrdiv16_fs165_not0;
  wire f_arrdiv16_fs165_and0;
  wire f_arrdiv16_fs165_xor1;
  wire f_arrdiv16_fs165_not1;
  wire f_arrdiv16_fs165_and1;
  wire f_arrdiv16_fs165_or0;
  wire f_arrdiv16_fs166_xor0;
  wire f_arrdiv16_fs166_not0;
  wire f_arrdiv16_fs166_and0;
  wire f_arrdiv16_fs166_xor1;
  wire f_arrdiv16_fs166_not1;
  wire f_arrdiv16_fs166_and1;
  wire f_arrdiv16_fs166_or0;
  wire f_arrdiv16_fs167_xor0;
  wire f_arrdiv16_fs167_not0;
  wire f_arrdiv16_fs167_and0;
  wire f_arrdiv16_fs167_xor1;
  wire f_arrdiv16_fs167_not1;
  wire f_arrdiv16_fs167_and1;
  wire f_arrdiv16_fs167_or0;
  wire f_arrdiv16_fs168_xor0;
  wire f_arrdiv16_fs168_not0;
  wire f_arrdiv16_fs168_and0;
  wire f_arrdiv16_fs168_xor1;
  wire f_arrdiv16_fs168_not1;
  wire f_arrdiv16_fs168_and1;
  wire f_arrdiv16_fs168_or0;
  wire f_arrdiv16_fs169_xor0;
  wire f_arrdiv16_fs169_not0;
  wire f_arrdiv16_fs169_and0;
  wire f_arrdiv16_fs169_xor1;
  wire f_arrdiv16_fs169_not1;
  wire f_arrdiv16_fs169_and1;
  wire f_arrdiv16_fs169_or0;
  wire f_arrdiv16_fs170_xor0;
  wire f_arrdiv16_fs170_not0;
  wire f_arrdiv16_fs170_and0;
  wire f_arrdiv16_fs170_xor1;
  wire f_arrdiv16_fs170_not1;
  wire f_arrdiv16_fs170_and1;
  wire f_arrdiv16_fs170_or0;
  wire f_arrdiv16_fs171_xor0;
  wire f_arrdiv16_fs171_not0;
  wire f_arrdiv16_fs171_and0;
  wire f_arrdiv16_fs171_xor1;
  wire f_arrdiv16_fs171_not1;
  wire f_arrdiv16_fs171_and1;
  wire f_arrdiv16_fs171_or0;
  wire f_arrdiv16_fs172_xor0;
  wire f_arrdiv16_fs172_not0;
  wire f_arrdiv16_fs172_and0;
  wire f_arrdiv16_fs172_xor1;
  wire f_arrdiv16_fs172_not1;
  wire f_arrdiv16_fs172_and1;
  wire f_arrdiv16_fs172_or0;
  wire f_arrdiv16_fs173_xor0;
  wire f_arrdiv16_fs173_not0;
  wire f_arrdiv16_fs173_and0;
  wire f_arrdiv16_fs173_xor1;
  wire f_arrdiv16_fs173_not1;
  wire f_arrdiv16_fs173_and1;
  wire f_arrdiv16_fs173_or0;
  wire f_arrdiv16_fs174_xor0;
  wire f_arrdiv16_fs174_not0;
  wire f_arrdiv16_fs174_and0;
  wire f_arrdiv16_fs174_xor1;
  wire f_arrdiv16_fs174_not1;
  wire f_arrdiv16_fs174_and1;
  wire f_arrdiv16_fs174_or0;
  wire f_arrdiv16_fs175_xor0;
  wire f_arrdiv16_fs175_not0;
  wire f_arrdiv16_fs175_and0;
  wire f_arrdiv16_fs175_xor1;
  wire f_arrdiv16_fs175_not1;
  wire f_arrdiv16_fs175_and1;
  wire f_arrdiv16_fs175_or0;
  wire f_arrdiv16_mux2to1150_and0;
  wire f_arrdiv16_mux2to1150_not0;
  wire f_arrdiv16_mux2to1150_and1;
  wire f_arrdiv16_mux2to1150_xor0;
  wire f_arrdiv16_mux2to1151_and0;
  wire f_arrdiv16_mux2to1151_not0;
  wire f_arrdiv16_mux2to1151_and1;
  wire f_arrdiv16_mux2to1151_xor0;
  wire f_arrdiv16_mux2to1152_and0;
  wire f_arrdiv16_mux2to1152_not0;
  wire f_arrdiv16_mux2to1152_and1;
  wire f_arrdiv16_mux2to1152_xor0;
  wire f_arrdiv16_mux2to1153_and0;
  wire f_arrdiv16_mux2to1153_not0;
  wire f_arrdiv16_mux2to1153_and1;
  wire f_arrdiv16_mux2to1153_xor0;
  wire f_arrdiv16_mux2to1154_and0;
  wire f_arrdiv16_mux2to1154_not0;
  wire f_arrdiv16_mux2to1154_and1;
  wire f_arrdiv16_mux2to1154_xor0;
  wire f_arrdiv16_mux2to1155_and0;
  wire f_arrdiv16_mux2to1155_not0;
  wire f_arrdiv16_mux2to1155_and1;
  wire f_arrdiv16_mux2to1155_xor0;
  wire f_arrdiv16_mux2to1156_and0;
  wire f_arrdiv16_mux2to1156_not0;
  wire f_arrdiv16_mux2to1156_and1;
  wire f_arrdiv16_mux2to1156_xor0;
  wire f_arrdiv16_mux2to1157_and0;
  wire f_arrdiv16_mux2to1157_not0;
  wire f_arrdiv16_mux2to1157_and1;
  wire f_arrdiv16_mux2to1157_xor0;
  wire f_arrdiv16_mux2to1158_and0;
  wire f_arrdiv16_mux2to1158_not0;
  wire f_arrdiv16_mux2to1158_and1;
  wire f_arrdiv16_mux2to1158_xor0;
  wire f_arrdiv16_mux2to1159_and0;
  wire f_arrdiv16_mux2to1159_not0;
  wire f_arrdiv16_mux2to1159_and1;
  wire f_arrdiv16_mux2to1159_xor0;
  wire f_arrdiv16_mux2to1160_and0;
  wire f_arrdiv16_mux2to1160_not0;
  wire f_arrdiv16_mux2to1160_and1;
  wire f_arrdiv16_mux2to1160_xor0;
  wire f_arrdiv16_mux2to1161_and0;
  wire f_arrdiv16_mux2to1161_not0;
  wire f_arrdiv16_mux2to1161_and1;
  wire f_arrdiv16_mux2to1161_xor0;
  wire f_arrdiv16_mux2to1162_and0;
  wire f_arrdiv16_mux2to1162_not0;
  wire f_arrdiv16_mux2to1162_and1;
  wire f_arrdiv16_mux2to1162_xor0;
  wire f_arrdiv16_mux2to1163_and0;
  wire f_arrdiv16_mux2to1163_not0;
  wire f_arrdiv16_mux2to1163_and1;
  wire f_arrdiv16_mux2to1163_xor0;
  wire f_arrdiv16_mux2to1164_and0;
  wire f_arrdiv16_mux2to1164_not0;
  wire f_arrdiv16_mux2to1164_and1;
  wire f_arrdiv16_mux2to1164_xor0;
  wire f_arrdiv16_not10;
  wire f_arrdiv16_fs176_xor0;
  wire f_arrdiv16_fs176_not0;
  wire f_arrdiv16_fs176_and0;
  wire f_arrdiv16_fs176_not1;
  wire f_arrdiv16_fs177_xor0;
  wire f_arrdiv16_fs177_not0;
  wire f_arrdiv16_fs177_and0;
  wire f_arrdiv16_fs177_xor1;
  wire f_arrdiv16_fs177_not1;
  wire f_arrdiv16_fs177_and1;
  wire f_arrdiv16_fs177_or0;
  wire f_arrdiv16_fs178_xor0;
  wire f_arrdiv16_fs178_not0;
  wire f_arrdiv16_fs178_and0;
  wire f_arrdiv16_fs178_xor1;
  wire f_arrdiv16_fs178_not1;
  wire f_arrdiv16_fs178_and1;
  wire f_arrdiv16_fs178_or0;
  wire f_arrdiv16_fs179_xor0;
  wire f_arrdiv16_fs179_not0;
  wire f_arrdiv16_fs179_and0;
  wire f_arrdiv16_fs179_xor1;
  wire f_arrdiv16_fs179_not1;
  wire f_arrdiv16_fs179_and1;
  wire f_arrdiv16_fs179_or0;
  wire f_arrdiv16_fs180_xor0;
  wire f_arrdiv16_fs180_not0;
  wire f_arrdiv16_fs180_and0;
  wire f_arrdiv16_fs180_xor1;
  wire f_arrdiv16_fs180_not1;
  wire f_arrdiv16_fs180_and1;
  wire f_arrdiv16_fs180_or0;
  wire f_arrdiv16_fs181_xor0;
  wire f_arrdiv16_fs181_not0;
  wire f_arrdiv16_fs181_and0;
  wire f_arrdiv16_fs181_xor1;
  wire f_arrdiv16_fs181_not1;
  wire f_arrdiv16_fs181_and1;
  wire f_arrdiv16_fs181_or0;
  wire f_arrdiv16_fs182_xor0;
  wire f_arrdiv16_fs182_not0;
  wire f_arrdiv16_fs182_and0;
  wire f_arrdiv16_fs182_xor1;
  wire f_arrdiv16_fs182_not1;
  wire f_arrdiv16_fs182_and1;
  wire f_arrdiv16_fs182_or0;
  wire f_arrdiv16_fs183_xor0;
  wire f_arrdiv16_fs183_not0;
  wire f_arrdiv16_fs183_and0;
  wire f_arrdiv16_fs183_xor1;
  wire f_arrdiv16_fs183_not1;
  wire f_arrdiv16_fs183_and1;
  wire f_arrdiv16_fs183_or0;
  wire f_arrdiv16_fs184_xor0;
  wire f_arrdiv16_fs184_not0;
  wire f_arrdiv16_fs184_and0;
  wire f_arrdiv16_fs184_xor1;
  wire f_arrdiv16_fs184_not1;
  wire f_arrdiv16_fs184_and1;
  wire f_arrdiv16_fs184_or0;
  wire f_arrdiv16_fs185_xor0;
  wire f_arrdiv16_fs185_not0;
  wire f_arrdiv16_fs185_and0;
  wire f_arrdiv16_fs185_xor1;
  wire f_arrdiv16_fs185_not1;
  wire f_arrdiv16_fs185_and1;
  wire f_arrdiv16_fs185_or0;
  wire f_arrdiv16_fs186_xor0;
  wire f_arrdiv16_fs186_not0;
  wire f_arrdiv16_fs186_and0;
  wire f_arrdiv16_fs186_xor1;
  wire f_arrdiv16_fs186_not1;
  wire f_arrdiv16_fs186_and1;
  wire f_arrdiv16_fs186_or0;
  wire f_arrdiv16_fs187_xor0;
  wire f_arrdiv16_fs187_not0;
  wire f_arrdiv16_fs187_and0;
  wire f_arrdiv16_fs187_xor1;
  wire f_arrdiv16_fs187_not1;
  wire f_arrdiv16_fs187_and1;
  wire f_arrdiv16_fs187_or0;
  wire f_arrdiv16_fs188_xor0;
  wire f_arrdiv16_fs188_not0;
  wire f_arrdiv16_fs188_and0;
  wire f_arrdiv16_fs188_xor1;
  wire f_arrdiv16_fs188_not1;
  wire f_arrdiv16_fs188_and1;
  wire f_arrdiv16_fs188_or0;
  wire f_arrdiv16_fs189_xor0;
  wire f_arrdiv16_fs189_not0;
  wire f_arrdiv16_fs189_and0;
  wire f_arrdiv16_fs189_xor1;
  wire f_arrdiv16_fs189_not1;
  wire f_arrdiv16_fs189_and1;
  wire f_arrdiv16_fs189_or0;
  wire f_arrdiv16_fs190_xor0;
  wire f_arrdiv16_fs190_not0;
  wire f_arrdiv16_fs190_and0;
  wire f_arrdiv16_fs190_xor1;
  wire f_arrdiv16_fs190_not1;
  wire f_arrdiv16_fs190_and1;
  wire f_arrdiv16_fs190_or0;
  wire f_arrdiv16_fs191_xor0;
  wire f_arrdiv16_fs191_not0;
  wire f_arrdiv16_fs191_and0;
  wire f_arrdiv16_fs191_xor1;
  wire f_arrdiv16_fs191_not1;
  wire f_arrdiv16_fs191_and1;
  wire f_arrdiv16_fs191_or0;
  wire f_arrdiv16_mux2to1165_and0;
  wire f_arrdiv16_mux2to1165_not0;
  wire f_arrdiv16_mux2to1165_and1;
  wire f_arrdiv16_mux2to1165_xor0;
  wire f_arrdiv16_mux2to1166_and0;
  wire f_arrdiv16_mux2to1166_not0;
  wire f_arrdiv16_mux2to1166_and1;
  wire f_arrdiv16_mux2to1166_xor0;
  wire f_arrdiv16_mux2to1167_and0;
  wire f_arrdiv16_mux2to1167_not0;
  wire f_arrdiv16_mux2to1167_and1;
  wire f_arrdiv16_mux2to1167_xor0;
  wire f_arrdiv16_mux2to1168_and0;
  wire f_arrdiv16_mux2to1168_not0;
  wire f_arrdiv16_mux2to1168_and1;
  wire f_arrdiv16_mux2to1168_xor0;
  wire f_arrdiv16_mux2to1169_and0;
  wire f_arrdiv16_mux2to1169_not0;
  wire f_arrdiv16_mux2to1169_and1;
  wire f_arrdiv16_mux2to1169_xor0;
  wire f_arrdiv16_mux2to1170_and0;
  wire f_arrdiv16_mux2to1170_not0;
  wire f_arrdiv16_mux2to1170_and1;
  wire f_arrdiv16_mux2to1170_xor0;
  wire f_arrdiv16_mux2to1171_and0;
  wire f_arrdiv16_mux2to1171_not0;
  wire f_arrdiv16_mux2to1171_and1;
  wire f_arrdiv16_mux2to1171_xor0;
  wire f_arrdiv16_mux2to1172_and0;
  wire f_arrdiv16_mux2to1172_not0;
  wire f_arrdiv16_mux2to1172_and1;
  wire f_arrdiv16_mux2to1172_xor0;
  wire f_arrdiv16_mux2to1173_and0;
  wire f_arrdiv16_mux2to1173_not0;
  wire f_arrdiv16_mux2to1173_and1;
  wire f_arrdiv16_mux2to1173_xor0;
  wire f_arrdiv16_mux2to1174_and0;
  wire f_arrdiv16_mux2to1174_not0;
  wire f_arrdiv16_mux2to1174_and1;
  wire f_arrdiv16_mux2to1174_xor0;
  wire f_arrdiv16_mux2to1175_and0;
  wire f_arrdiv16_mux2to1175_not0;
  wire f_arrdiv16_mux2to1175_and1;
  wire f_arrdiv16_mux2to1175_xor0;
  wire f_arrdiv16_mux2to1176_and0;
  wire f_arrdiv16_mux2to1176_not0;
  wire f_arrdiv16_mux2to1176_and1;
  wire f_arrdiv16_mux2to1176_xor0;
  wire f_arrdiv16_mux2to1177_and0;
  wire f_arrdiv16_mux2to1177_not0;
  wire f_arrdiv16_mux2to1177_and1;
  wire f_arrdiv16_mux2to1177_xor0;
  wire f_arrdiv16_mux2to1178_and0;
  wire f_arrdiv16_mux2to1178_not0;
  wire f_arrdiv16_mux2to1178_and1;
  wire f_arrdiv16_mux2to1178_xor0;
  wire f_arrdiv16_mux2to1179_and0;
  wire f_arrdiv16_mux2to1179_not0;
  wire f_arrdiv16_mux2to1179_and1;
  wire f_arrdiv16_mux2to1179_xor0;
  wire f_arrdiv16_not11;
  wire f_arrdiv16_fs192_xor0;
  wire f_arrdiv16_fs192_not0;
  wire f_arrdiv16_fs192_and0;
  wire f_arrdiv16_fs192_not1;
  wire f_arrdiv16_fs193_xor0;
  wire f_arrdiv16_fs193_not0;
  wire f_arrdiv16_fs193_and0;
  wire f_arrdiv16_fs193_xor1;
  wire f_arrdiv16_fs193_not1;
  wire f_arrdiv16_fs193_and1;
  wire f_arrdiv16_fs193_or0;
  wire f_arrdiv16_fs194_xor0;
  wire f_arrdiv16_fs194_not0;
  wire f_arrdiv16_fs194_and0;
  wire f_arrdiv16_fs194_xor1;
  wire f_arrdiv16_fs194_not1;
  wire f_arrdiv16_fs194_and1;
  wire f_arrdiv16_fs194_or0;
  wire f_arrdiv16_fs195_xor0;
  wire f_arrdiv16_fs195_not0;
  wire f_arrdiv16_fs195_and0;
  wire f_arrdiv16_fs195_xor1;
  wire f_arrdiv16_fs195_not1;
  wire f_arrdiv16_fs195_and1;
  wire f_arrdiv16_fs195_or0;
  wire f_arrdiv16_fs196_xor0;
  wire f_arrdiv16_fs196_not0;
  wire f_arrdiv16_fs196_and0;
  wire f_arrdiv16_fs196_xor1;
  wire f_arrdiv16_fs196_not1;
  wire f_arrdiv16_fs196_and1;
  wire f_arrdiv16_fs196_or0;
  wire f_arrdiv16_fs197_xor0;
  wire f_arrdiv16_fs197_not0;
  wire f_arrdiv16_fs197_and0;
  wire f_arrdiv16_fs197_xor1;
  wire f_arrdiv16_fs197_not1;
  wire f_arrdiv16_fs197_and1;
  wire f_arrdiv16_fs197_or0;
  wire f_arrdiv16_fs198_xor0;
  wire f_arrdiv16_fs198_not0;
  wire f_arrdiv16_fs198_and0;
  wire f_arrdiv16_fs198_xor1;
  wire f_arrdiv16_fs198_not1;
  wire f_arrdiv16_fs198_and1;
  wire f_arrdiv16_fs198_or0;
  wire f_arrdiv16_fs199_xor0;
  wire f_arrdiv16_fs199_not0;
  wire f_arrdiv16_fs199_and0;
  wire f_arrdiv16_fs199_xor1;
  wire f_arrdiv16_fs199_not1;
  wire f_arrdiv16_fs199_and1;
  wire f_arrdiv16_fs199_or0;
  wire f_arrdiv16_fs200_xor0;
  wire f_arrdiv16_fs200_not0;
  wire f_arrdiv16_fs200_and0;
  wire f_arrdiv16_fs200_xor1;
  wire f_arrdiv16_fs200_not1;
  wire f_arrdiv16_fs200_and1;
  wire f_arrdiv16_fs200_or0;
  wire f_arrdiv16_fs201_xor0;
  wire f_arrdiv16_fs201_not0;
  wire f_arrdiv16_fs201_and0;
  wire f_arrdiv16_fs201_xor1;
  wire f_arrdiv16_fs201_not1;
  wire f_arrdiv16_fs201_and1;
  wire f_arrdiv16_fs201_or0;
  wire f_arrdiv16_fs202_xor0;
  wire f_arrdiv16_fs202_not0;
  wire f_arrdiv16_fs202_and0;
  wire f_arrdiv16_fs202_xor1;
  wire f_arrdiv16_fs202_not1;
  wire f_arrdiv16_fs202_and1;
  wire f_arrdiv16_fs202_or0;
  wire f_arrdiv16_fs203_xor0;
  wire f_arrdiv16_fs203_not0;
  wire f_arrdiv16_fs203_and0;
  wire f_arrdiv16_fs203_xor1;
  wire f_arrdiv16_fs203_not1;
  wire f_arrdiv16_fs203_and1;
  wire f_arrdiv16_fs203_or0;
  wire f_arrdiv16_fs204_xor0;
  wire f_arrdiv16_fs204_not0;
  wire f_arrdiv16_fs204_and0;
  wire f_arrdiv16_fs204_xor1;
  wire f_arrdiv16_fs204_not1;
  wire f_arrdiv16_fs204_and1;
  wire f_arrdiv16_fs204_or0;
  wire f_arrdiv16_fs205_xor0;
  wire f_arrdiv16_fs205_not0;
  wire f_arrdiv16_fs205_and0;
  wire f_arrdiv16_fs205_xor1;
  wire f_arrdiv16_fs205_not1;
  wire f_arrdiv16_fs205_and1;
  wire f_arrdiv16_fs205_or0;
  wire f_arrdiv16_fs206_xor0;
  wire f_arrdiv16_fs206_not0;
  wire f_arrdiv16_fs206_and0;
  wire f_arrdiv16_fs206_xor1;
  wire f_arrdiv16_fs206_not1;
  wire f_arrdiv16_fs206_and1;
  wire f_arrdiv16_fs206_or0;
  wire f_arrdiv16_fs207_xor0;
  wire f_arrdiv16_fs207_not0;
  wire f_arrdiv16_fs207_and0;
  wire f_arrdiv16_fs207_xor1;
  wire f_arrdiv16_fs207_not1;
  wire f_arrdiv16_fs207_and1;
  wire f_arrdiv16_fs207_or0;
  wire f_arrdiv16_mux2to1180_and0;
  wire f_arrdiv16_mux2to1180_not0;
  wire f_arrdiv16_mux2to1180_and1;
  wire f_arrdiv16_mux2to1180_xor0;
  wire f_arrdiv16_mux2to1181_and0;
  wire f_arrdiv16_mux2to1181_not0;
  wire f_arrdiv16_mux2to1181_and1;
  wire f_arrdiv16_mux2to1181_xor0;
  wire f_arrdiv16_mux2to1182_and0;
  wire f_arrdiv16_mux2to1182_not0;
  wire f_arrdiv16_mux2to1182_and1;
  wire f_arrdiv16_mux2to1182_xor0;
  wire f_arrdiv16_mux2to1183_and0;
  wire f_arrdiv16_mux2to1183_not0;
  wire f_arrdiv16_mux2to1183_and1;
  wire f_arrdiv16_mux2to1183_xor0;
  wire f_arrdiv16_mux2to1184_and0;
  wire f_arrdiv16_mux2to1184_not0;
  wire f_arrdiv16_mux2to1184_and1;
  wire f_arrdiv16_mux2to1184_xor0;
  wire f_arrdiv16_mux2to1185_and0;
  wire f_arrdiv16_mux2to1185_not0;
  wire f_arrdiv16_mux2to1185_and1;
  wire f_arrdiv16_mux2to1185_xor0;
  wire f_arrdiv16_mux2to1186_and0;
  wire f_arrdiv16_mux2to1186_not0;
  wire f_arrdiv16_mux2to1186_and1;
  wire f_arrdiv16_mux2to1186_xor0;
  wire f_arrdiv16_mux2to1187_and0;
  wire f_arrdiv16_mux2to1187_not0;
  wire f_arrdiv16_mux2to1187_and1;
  wire f_arrdiv16_mux2to1187_xor0;
  wire f_arrdiv16_mux2to1188_and0;
  wire f_arrdiv16_mux2to1188_not0;
  wire f_arrdiv16_mux2to1188_and1;
  wire f_arrdiv16_mux2to1188_xor0;
  wire f_arrdiv16_mux2to1189_and0;
  wire f_arrdiv16_mux2to1189_not0;
  wire f_arrdiv16_mux2to1189_and1;
  wire f_arrdiv16_mux2to1189_xor0;
  wire f_arrdiv16_mux2to1190_and0;
  wire f_arrdiv16_mux2to1190_not0;
  wire f_arrdiv16_mux2to1190_and1;
  wire f_arrdiv16_mux2to1190_xor0;
  wire f_arrdiv16_mux2to1191_and0;
  wire f_arrdiv16_mux2to1191_not0;
  wire f_arrdiv16_mux2to1191_and1;
  wire f_arrdiv16_mux2to1191_xor0;
  wire f_arrdiv16_mux2to1192_and0;
  wire f_arrdiv16_mux2to1192_not0;
  wire f_arrdiv16_mux2to1192_and1;
  wire f_arrdiv16_mux2to1192_xor0;
  wire f_arrdiv16_mux2to1193_and0;
  wire f_arrdiv16_mux2to1193_not0;
  wire f_arrdiv16_mux2to1193_and1;
  wire f_arrdiv16_mux2to1193_xor0;
  wire f_arrdiv16_mux2to1194_and0;
  wire f_arrdiv16_mux2to1194_not0;
  wire f_arrdiv16_mux2to1194_and1;
  wire f_arrdiv16_mux2to1194_xor0;
  wire f_arrdiv16_not12;
  wire f_arrdiv16_fs208_xor0;
  wire f_arrdiv16_fs208_not0;
  wire f_arrdiv16_fs208_and0;
  wire f_arrdiv16_fs208_not1;
  wire f_arrdiv16_fs209_xor0;
  wire f_arrdiv16_fs209_not0;
  wire f_arrdiv16_fs209_and0;
  wire f_arrdiv16_fs209_xor1;
  wire f_arrdiv16_fs209_not1;
  wire f_arrdiv16_fs209_and1;
  wire f_arrdiv16_fs209_or0;
  wire f_arrdiv16_fs210_xor0;
  wire f_arrdiv16_fs210_not0;
  wire f_arrdiv16_fs210_and0;
  wire f_arrdiv16_fs210_xor1;
  wire f_arrdiv16_fs210_not1;
  wire f_arrdiv16_fs210_and1;
  wire f_arrdiv16_fs210_or0;
  wire f_arrdiv16_fs211_xor0;
  wire f_arrdiv16_fs211_not0;
  wire f_arrdiv16_fs211_and0;
  wire f_arrdiv16_fs211_xor1;
  wire f_arrdiv16_fs211_not1;
  wire f_arrdiv16_fs211_and1;
  wire f_arrdiv16_fs211_or0;
  wire f_arrdiv16_fs212_xor0;
  wire f_arrdiv16_fs212_not0;
  wire f_arrdiv16_fs212_and0;
  wire f_arrdiv16_fs212_xor1;
  wire f_arrdiv16_fs212_not1;
  wire f_arrdiv16_fs212_and1;
  wire f_arrdiv16_fs212_or0;
  wire f_arrdiv16_fs213_xor0;
  wire f_arrdiv16_fs213_not0;
  wire f_arrdiv16_fs213_and0;
  wire f_arrdiv16_fs213_xor1;
  wire f_arrdiv16_fs213_not1;
  wire f_arrdiv16_fs213_and1;
  wire f_arrdiv16_fs213_or0;
  wire f_arrdiv16_fs214_xor0;
  wire f_arrdiv16_fs214_not0;
  wire f_arrdiv16_fs214_and0;
  wire f_arrdiv16_fs214_xor1;
  wire f_arrdiv16_fs214_not1;
  wire f_arrdiv16_fs214_and1;
  wire f_arrdiv16_fs214_or0;
  wire f_arrdiv16_fs215_xor0;
  wire f_arrdiv16_fs215_not0;
  wire f_arrdiv16_fs215_and0;
  wire f_arrdiv16_fs215_xor1;
  wire f_arrdiv16_fs215_not1;
  wire f_arrdiv16_fs215_and1;
  wire f_arrdiv16_fs215_or0;
  wire f_arrdiv16_fs216_xor0;
  wire f_arrdiv16_fs216_not0;
  wire f_arrdiv16_fs216_and0;
  wire f_arrdiv16_fs216_xor1;
  wire f_arrdiv16_fs216_not1;
  wire f_arrdiv16_fs216_and1;
  wire f_arrdiv16_fs216_or0;
  wire f_arrdiv16_fs217_xor0;
  wire f_arrdiv16_fs217_not0;
  wire f_arrdiv16_fs217_and0;
  wire f_arrdiv16_fs217_xor1;
  wire f_arrdiv16_fs217_not1;
  wire f_arrdiv16_fs217_and1;
  wire f_arrdiv16_fs217_or0;
  wire f_arrdiv16_fs218_xor0;
  wire f_arrdiv16_fs218_not0;
  wire f_arrdiv16_fs218_and0;
  wire f_arrdiv16_fs218_xor1;
  wire f_arrdiv16_fs218_not1;
  wire f_arrdiv16_fs218_and1;
  wire f_arrdiv16_fs218_or0;
  wire f_arrdiv16_fs219_xor0;
  wire f_arrdiv16_fs219_not0;
  wire f_arrdiv16_fs219_and0;
  wire f_arrdiv16_fs219_xor1;
  wire f_arrdiv16_fs219_not1;
  wire f_arrdiv16_fs219_and1;
  wire f_arrdiv16_fs219_or0;
  wire f_arrdiv16_fs220_xor0;
  wire f_arrdiv16_fs220_not0;
  wire f_arrdiv16_fs220_and0;
  wire f_arrdiv16_fs220_xor1;
  wire f_arrdiv16_fs220_not1;
  wire f_arrdiv16_fs220_and1;
  wire f_arrdiv16_fs220_or0;
  wire f_arrdiv16_fs221_xor0;
  wire f_arrdiv16_fs221_not0;
  wire f_arrdiv16_fs221_and0;
  wire f_arrdiv16_fs221_xor1;
  wire f_arrdiv16_fs221_not1;
  wire f_arrdiv16_fs221_and1;
  wire f_arrdiv16_fs221_or0;
  wire f_arrdiv16_fs222_xor0;
  wire f_arrdiv16_fs222_not0;
  wire f_arrdiv16_fs222_and0;
  wire f_arrdiv16_fs222_xor1;
  wire f_arrdiv16_fs222_not1;
  wire f_arrdiv16_fs222_and1;
  wire f_arrdiv16_fs222_or0;
  wire f_arrdiv16_fs223_xor0;
  wire f_arrdiv16_fs223_not0;
  wire f_arrdiv16_fs223_and0;
  wire f_arrdiv16_fs223_xor1;
  wire f_arrdiv16_fs223_not1;
  wire f_arrdiv16_fs223_and1;
  wire f_arrdiv16_fs223_or0;
  wire f_arrdiv16_mux2to1195_and0;
  wire f_arrdiv16_mux2to1195_not0;
  wire f_arrdiv16_mux2to1195_and1;
  wire f_arrdiv16_mux2to1195_xor0;
  wire f_arrdiv16_mux2to1196_and0;
  wire f_arrdiv16_mux2to1196_not0;
  wire f_arrdiv16_mux2to1196_and1;
  wire f_arrdiv16_mux2to1196_xor0;
  wire f_arrdiv16_mux2to1197_and0;
  wire f_arrdiv16_mux2to1197_not0;
  wire f_arrdiv16_mux2to1197_and1;
  wire f_arrdiv16_mux2to1197_xor0;
  wire f_arrdiv16_mux2to1198_and0;
  wire f_arrdiv16_mux2to1198_not0;
  wire f_arrdiv16_mux2to1198_and1;
  wire f_arrdiv16_mux2to1198_xor0;
  wire f_arrdiv16_mux2to1199_and0;
  wire f_arrdiv16_mux2to1199_not0;
  wire f_arrdiv16_mux2to1199_and1;
  wire f_arrdiv16_mux2to1199_xor0;
  wire f_arrdiv16_mux2to1200_and0;
  wire f_arrdiv16_mux2to1200_not0;
  wire f_arrdiv16_mux2to1200_and1;
  wire f_arrdiv16_mux2to1200_xor0;
  wire f_arrdiv16_mux2to1201_and0;
  wire f_arrdiv16_mux2to1201_not0;
  wire f_arrdiv16_mux2to1201_and1;
  wire f_arrdiv16_mux2to1201_xor0;
  wire f_arrdiv16_mux2to1202_and0;
  wire f_arrdiv16_mux2to1202_not0;
  wire f_arrdiv16_mux2to1202_and1;
  wire f_arrdiv16_mux2to1202_xor0;
  wire f_arrdiv16_mux2to1203_and0;
  wire f_arrdiv16_mux2to1203_not0;
  wire f_arrdiv16_mux2to1203_and1;
  wire f_arrdiv16_mux2to1203_xor0;
  wire f_arrdiv16_mux2to1204_and0;
  wire f_arrdiv16_mux2to1204_not0;
  wire f_arrdiv16_mux2to1204_and1;
  wire f_arrdiv16_mux2to1204_xor0;
  wire f_arrdiv16_mux2to1205_and0;
  wire f_arrdiv16_mux2to1205_not0;
  wire f_arrdiv16_mux2to1205_and1;
  wire f_arrdiv16_mux2to1205_xor0;
  wire f_arrdiv16_mux2to1206_and0;
  wire f_arrdiv16_mux2to1206_not0;
  wire f_arrdiv16_mux2to1206_and1;
  wire f_arrdiv16_mux2to1206_xor0;
  wire f_arrdiv16_mux2to1207_and0;
  wire f_arrdiv16_mux2to1207_not0;
  wire f_arrdiv16_mux2to1207_and1;
  wire f_arrdiv16_mux2to1207_xor0;
  wire f_arrdiv16_mux2to1208_and0;
  wire f_arrdiv16_mux2to1208_not0;
  wire f_arrdiv16_mux2to1208_and1;
  wire f_arrdiv16_mux2to1208_xor0;
  wire f_arrdiv16_mux2to1209_and0;
  wire f_arrdiv16_mux2to1209_not0;
  wire f_arrdiv16_mux2to1209_and1;
  wire f_arrdiv16_mux2to1209_xor0;
  wire f_arrdiv16_not13;
  wire f_arrdiv16_fs224_xor0;
  wire f_arrdiv16_fs224_not0;
  wire f_arrdiv16_fs224_and0;
  wire f_arrdiv16_fs224_not1;
  wire f_arrdiv16_fs225_xor0;
  wire f_arrdiv16_fs225_not0;
  wire f_arrdiv16_fs225_and0;
  wire f_arrdiv16_fs225_xor1;
  wire f_arrdiv16_fs225_not1;
  wire f_arrdiv16_fs225_and1;
  wire f_arrdiv16_fs225_or0;
  wire f_arrdiv16_fs226_xor0;
  wire f_arrdiv16_fs226_not0;
  wire f_arrdiv16_fs226_and0;
  wire f_arrdiv16_fs226_xor1;
  wire f_arrdiv16_fs226_not1;
  wire f_arrdiv16_fs226_and1;
  wire f_arrdiv16_fs226_or0;
  wire f_arrdiv16_fs227_xor0;
  wire f_arrdiv16_fs227_not0;
  wire f_arrdiv16_fs227_and0;
  wire f_arrdiv16_fs227_xor1;
  wire f_arrdiv16_fs227_not1;
  wire f_arrdiv16_fs227_and1;
  wire f_arrdiv16_fs227_or0;
  wire f_arrdiv16_fs228_xor0;
  wire f_arrdiv16_fs228_not0;
  wire f_arrdiv16_fs228_and0;
  wire f_arrdiv16_fs228_xor1;
  wire f_arrdiv16_fs228_not1;
  wire f_arrdiv16_fs228_and1;
  wire f_arrdiv16_fs228_or0;
  wire f_arrdiv16_fs229_xor0;
  wire f_arrdiv16_fs229_not0;
  wire f_arrdiv16_fs229_and0;
  wire f_arrdiv16_fs229_xor1;
  wire f_arrdiv16_fs229_not1;
  wire f_arrdiv16_fs229_and1;
  wire f_arrdiv16_fs229_or0;
  wire f_arrdiv16_fs230_xor0;
  wire f_arrdiv16_fs230_not0;
  wire f_arrdiv16_fs230_and0;
  wire f_arrdiv16_fs230_xor1;
  wire f_arrdiv16_fs230_not1;
  wire f_arrdiv16_fs230_and1;
  wire f_arrdiv16_fs230_or0;
  wire f_arrdiv16_fs231_xor0;
  wire f_arrdiv16_fs231_not0;
  wire f_arrdiv16_fs231_and0;
  wire f_arrdiv16_fs231_xor1;
  wire f_arrdiv16_fs231_not1;
  wire f_arrdiv16_fs231_and1;
  wire f_arrdiv16_fs231_or0;
  wire f_arrdiv16_fs232_xor0;
  wire f_arrdiv16_fs232_not0;
  wire f_arrdiv16_fs232_and0;
  wire f_arrdiv16_fs232_xor1;
  wire f_arrdiv16_fs232_not1;
  wire f_arrdiv16_fs232_and1;
  wire f_arrdiv16_fs232_or0;
  wire f_arrdiv16_fs233_xor0;
  wire f_arrdiv16_fs233_not0;
  wire f_arrdiv16_fs233_and0;
  wire f_arrdiv16_fs233_xor1;
  wire f_arrdiv16_fs233_not1;
  wire f_arrdiv16_fs233_and1;
  wire f_arrdiv16_fs233_or0;
  wire f_arrdiv16_fs234_xor0;
  wire f_arrdiv16_fs234_not0;
  wire f_arrdiv16_fs234_and0;
  wire f_arrdiv16_fs234_xor1;
  wire f_arrdiv16_fs234_not1;
  wire f_arrdiv16_fs234_and1;
  wire f_arrdiv16_fs234_or0;
  wire f_arrdiv16_fs235_xor0;
  wire f_arrdiv16_fs235_not0;
  wire f_arrdiv16_fs235_and0;
  wire f_arrdiv16_fs235_xor1;
  wire f_arrdiv16_fs235_not1;
  wire f_arrdiv16_fs235_and1;
  wire f_arrdiv16_fs235_or0;
  wire f_arrdiv16_fs236_xor0;
  wire f_arrdiv16_fs236_not0;
  wire f_arrdiv16_fs236_and0;
  wire f_arrdiv16_fs236_xor1;
  wire f_arrdiv16_fs236_not1;
  wire f_arrdiv16_fs236_and1;
  wire f_arrdiv16_fs236_or0;
  wire f_arrdiv16_fs237_xor0;
  wire f_arrdiv16_fs237_not0;
  wire f_arrdiv16_fs237_and0;
  wire f_arrdiv16_fs237_xor1;
  wire f_arrdiv16_fs237_not1;
  wire f_arrdiv16_fs237_and1;
  wire f_arrdiv16_fs237_or0;
  wire f_arrdiv16_fs238_xor0;
  wire f_arrdiv16_fs238_not0;
  wire f_arrdiv16_fs238_and0;
  wire f_arrdiv16_fs238_xor1;
  wire f_arrdiv16_fs238_not1;
  wire f_arrdiv16_fs238_and1;
  wire f_arrdiv16_fs238_or0;
  wire f_arrdiv16_fs239_xor0;
  wire f_arrdiv16_fs239_not0;
  wire f_arrdiv16_fs239_and0;
  wire f_arrdiv16_fs239_xor1;
  wire f_arrdiv16_fs239_not1;
  wire f_arrdiv16_fs239_and1;
  wire f_arrdiv16_fs239_or0;
  wire f_arrdiv16_mux2to1210_and0;
  wire f_arrdiv16_mux2to1210_not0;
  wire f_arrdiv16_mux2to1210_and1;
  wire f_arrdiv16_mux2to1210_xor0;
  wire f_arrdiv16_mux2to1211_and0;
  wire f_arrdiv16_mux2to1211_not0;
  wire f_arrdiv16_mux2to1211_and1;
  wire f_arrdiv16_mux2to1211_xor0;
  wire f_arrdiv16_mux2to1212_and0;
  wire f_arrdiv16_mux2to1212_not0;
  wire f_arrdiv16_mux2to1212_and1;
  wire f_arrdiv16_mux2to1212_xor0;
  wire f_arrdiv16_mux2to1213_and0;
  wire f_arrdiv16_mux2to1213_not0;
  wire f_arrdiv16_mux2to1213_and1;
  wire f_arrdiv16_mux2to1213_xor0;
  wire f_arrdiv16_mux2to1214_and0;
  wire f_arrdiv16_mux2to1214_not0;
  wire f_arrdiv16_mux2to1214_and1;
  wire f_arrdiv16_mux2to1214_xor0;
  wire f_arrdiv16_mux2to1215_and0;
  wire f_arrdiv16_mux2to1215_not0;
  wire f_arrdiv16_mux2to1215_and1;
  wire f_arrdiv16_mux2to1215_xor0;
  wire f_arrdiv16_mux2to1216_and0;
  wire f_arrdiv16_mux2to1216_not0;
  wire f_arrdiv16_mux2to1216_and1;
  wire f_arrdiv16_mux2to1216_xor0;
  wire f_arrdiv16_mux2to1217_and0;
  wire f_arrdiv16_mux2to1217_not0;
  wire f_arrdiv16_mux2to1217_and1;
  wire f_arrdiv16_mux2to1217_xor0;
  wire f_arrdiv16_mux2to1218_and0;
  wire f_arrdiv16_mux2to1218_not0;
  wire f_arrdiv16_mux2to1218_and1;
  wire f_arrdiv16_mux2to1218_xor0;
  wire f_arrdiv16_mux2to1219_and0;
  wire f_arrdiv16_mux2to1219_not0;
  wire f_arrdiv16_mux2to1219_and1;
  wire f_arrdiv16_mux2to1219_xor0;
  wire f_arrdiv16_mux2to1220_and0;
  wire f_arrdiv16_mux2to1220_not0;
  wire f_arrdiv16_mux2to1220_and1;
  wire f_arrdiv16_mux2to1220_xor0;
  wire f_arrdiv16_mux2to1221_and0;
  wire f_arrdiv16_mux2to1221_not0;
  wire f_arrdiv16_mux2to1221_and1;
  wire f_arrdiv16_mux2to1221_xor0;
  wire f_arrdiv16_mux2to1222_and0;
  wire f_arrdiv16_mux2to1222_not0;
  wire f_arrdiv16_mux2to1222_and1;
  wire f_arrdiv16_mux2to1222_xor0;
  wire f_arrdiv16_mux2to1223_and0;
  wire f_arrdiv16_mux2to1223_not0;
  wire f_arrdiv16_mux2to1223_and1;
  wire f_arrdiv16_mux2to1223_xor0;
  wire f_arrdiv16_mux2to1224_and0;
  wire f_arrdiv16_mux2to1224_not0;
  wire f_arrdiv16_mux2to1224_and1;
  wire f_arrdiv16_mux2to1224_xor0;
  wire f_arrdiv16_not14;
  wire f_arrdiv16_fs240_xor0;
  wire f_arrdiv16_fs240_not0;
  wire f_arrdiv16_fs240_and0;
  wire f_arrdiv16_fs240_not1;
  wire f_arrdiv16_fs241_xor0;
  wire f_arrdiv16_fs241_not0;
  wire f_arrdiv16_fs241_and0;
  wire f_arrdiv16_fs241_xor1;
  wire f_arrdiv16_fs241_not1;
  wire f_arrdiv16_fs241_and1;
  wire f_arrdiv16_fs241_or0;
  wire f_arrdiv16_fs242_xor0;
  wire f_arrdiv16_fs242_not0;
  wire f_arrdiv16_fs242_and0;
  wire f_arrdiv16_fs242_xor1;
  wire f_arrdiv16_fs242_not1;
  wire f_arrdiv16_fs242_and1;
  wire f_arrdiv16_fs242_or0;
  wire f_arrdiv16_fs243_xor0;
  wire f_arrdiv16_fs243_not0;
  wire f_arrdiv16_fs243_and0;
  wire f_arrdiv16_fs243_xor1;
  wire f_arrdiv16_fs243_not1;
  wire f_arrdiv16_fs243_and1;
  wire f_arrdiv16_fs243_or0;
  wire f_arrdiv16_fs244_xor0;
  wire f_arrdiv16_fs244_not0;
  wire f_arrdiv16_fs244_and0;
  wire f_arrdiv16_fs244_xor1;
  wire f_arrdiv16_fs244_not1;
  wire f_arrdiv16_fs244_and1;
  wire f_arrdiv16_fs244_or0;
  wire f_arrdiv16_fs245_xor0;
  wire f_arrdiv16_fs245_not0;
  wire f_arrdiv16_fs245_and0;
  wire f_arrdiv16_fs245_xor1;
  wire f_arrdiv16_fs245_not1;
  wire f_arrdiv16_fs245_and1;
  wire f_arrdiv16_fs245_or0;
  wire f_arrdiv16_fs246_xor0;
  wire f_arrdiv16_fs246_not0;
  wire f_arrdiv16_fs246_and0;
  wire f_arrdiv16_fs246_xor1;
  wire f_arrdiv16_fs246_not1;
  wire f_arrdiv16_fs246_and1;
  wire f_arrdiv16_fs246_or0;
  wire f_arrdiv16_fs247_xor0;
  wire f_arrdiv16_fs247_not0;
  wire f_arrdiv16_fs247_and0;
  wire f_arrdiv16_fs247_xor1;
  wire f_arrdiv16_fs247_not1;
  wire f_arrdiv16_fs247_and1;
  wire f_arrdiv16_fs247_or0;
  wire f_arrdiv16_fs248_xor0;
  wire f_arrdiv16_fs248_not0;
  wire f_arrdiv16_fs248_and0;
  wire f_arrdiv16_fs248_xor1;
  wire f_arrdiv16_fs248_not1;
  wire f_arrdiv16_fs248_and1;
  wire f_arrdiv16_fs248_or0;
  wire f_arrdiv16_fs249_xor0;
  wire f_arrdiv16_fs249_not0;
  wire f_arrdiv16_fs249_and0;
  wire f_arrdiv16_fs249_xor1;
  wire f_arrdiv16_fs249_not1;
  wire f_arrdiv16_fs249_and1;
  wire f_arrdiv16_fs249_or0;
  wire f_arrdiv16_fs250_xor0;
  wire f_arrdiv16_fs250_not0;
  wire f_arrdiv16_fs250_and0;
  wire f_arrdiv16_fs250_xor1;
  wire f_arrdiv16_fs250_not1;
  wire f_arrdiv16_fs250_and1;
  wire f_arrdiv16_fs250_or0;
  wire f_arrdiv16_fs251_xor0;
  wire f_arrdiv16_fs251_not0;
  wire f_arrdiv16_fs251_and0;
  wire f_arrdiv16_fs251_xor1;
  wire f_arrdiv16_fs251_not1;
  wire f_arrdiv16_fs251_and1;
  wire f_arrdiv16_fs251_or0;
  wire f_arrdiv16_fs252_xor0;
  wire f_arrdiv16_fs252_not0;
  wire f_arrdiv16_fs252_and0;
  wire f_arrdiv16_fs252_xor1;
  wire f_arrdiv16_fs252_not1;
  wire f_arrdiv16_fs252_and1;
  wire f_arrdiv16_fs252_or0;
  wire f_arrdiv16_fs253_xor0;
  wire f_arrdiv16_fs253_not0;
  wire f_arrdiv16_fs253_and0;
  wire f_arrdiv16_fs253_xor1;
  wire f_arrdiv16_fs253_not1;
  wire f_arrdiv16_fs253_and1;
  wire f_arrdiv16_fs253_or0;
  wire f_arrdiv16_fs254_xor0;
  wire f_arrdiv16_fs254_not0;
  wire f_arrdiv16_fs254_and0;
  wire f_arrdiv16_fs254_xor1;
  wire f_arrdiv16_fs254_not1;
  wire f_arrdiv16_fs254_and1;
  wire f_arrdiv16_fs254_or0;
  wire f_arrdiv16_fs255_xor0;
  wire f_arrdiv16_fs255_not0;
  wire f_arrdiv16_fs255_and0;
  wire f_arrdiv16_fs255_xor1;
  wire f_arrdiv16_fs255_not1;
  wire f_arrdiv16_fs255_and1;
  wire f_arrdiv16_fs255_or0;
  wire f_arrdiv16_not15;

  assign f_arrdiv16_fs0_xor0 = a[15] ^ b[0];
  assign f_arrdiv16_fs0_not0 = ~a[15];
  assign f_arrdiv16_fs0_and0 = f_arrdiv16_fs0_not0 & b[0];
  assign f_arrdiv16_fs0_not1 = ~f_arrdiv16_fs0_xor0;
  assign f_arrdiv16_fs1_xor1 = f_arrdiv16_fs0_and0 ^ b[1];
  assign f_arrdiv16_fs1_not1 = ~b[1];
  assign f_arrdiv16_fs1_and1 = f_arrdiv16_fs1_not1 & f_arrdiv16_fs0_and0;
  assign f_arrdiv16_fs1_or0 = f_arrdiv16_fs1_and1 | b[1];
  assign f_arrdiv16_fs2_xor1 = f_arrdiv16_fs1_or0 ^ b[2];
  assign f_arrdiv16_fs2_not1 = ~b[2];
  assign f_arrdiv16_fs2_and1 = f_arrdiv16_fs2_not1 & f_arrdiv16_fs1_or0;
  assign f_arrdiv16_fs2_or0 = f_arrdiv16_fs2_and1 | b[2];
  assign f_arrdiv16_fs3_xor1 = f_arrdiv16_fs2_or0 ^ b[3];
  assign f_arrdiv16_fs3_not1 = ~b[3];
  assign f_arrdiv16_fs3_and1 = f_arrdiv16_fs3_not1 & f_arrdiv16_fs2_or0;
  assign f_arrdiv16_fs3_or0 = f_arrdiv16_fs3_and1 | b[3];
  assign f_arrdiv16_fs4_xor1 = f_arrdiv16_fs3_or0 ^ b[4];
  assign f_arrdiv16_fs4_not1 = ~b[4];
  assign f_arrdiv16_fs4_and1 = f_arrdiv16_fs4_not1 & f_arrdiv16_fs3_or0;
  assign f_arrdiv16_fs4_or0 = f_arrdiv16_fs4_and1 | b[4];
  assign f_arrdiv16_fs5_xor1 = f_arrdiv16_fs4_or0 ^ b[5];
  assign f_arrdiv16_fs5_not1 = ~b[5];
  assign f_arrdiv16_fs5_and1 = f_arrdiv16_fs5_not1 & f_arrdiv16_fs4_or0;
  assign f_arrdiv16_fs5_or0 = f_arrdiv16_fs5_and1 | b[5];
  assign f_arrdiv16_fs6_xor1 = f_arrdiv16_fs5_or0 ^ b[6];
  assign f_arrdiv16_fs6_not1 = ~b[6];
  assign f_arrdiv16_fs6_and1 = f_arrdiv16_fs6_not1 & f_arrdiv16_fs5_or0;
  assign f_arrdiv16_fs6_or0 = f_arrdiv16_fs6_and1 | b[6];
  assign f_arrdiv16_fs7_xor1 = f_arrdiv16_fs6_or0 ^ b[7];
  assign f_arrdiv16_fs7_not1 = ~b[7];
  assign f_arrdiv16_fs7_and1 = f_arrdiv16_fs7_not1 & f_arrdiv16_fs6_or0;
  assign f_arrdiv16_fs7_or0 = f_arrdiv16_fs7_and1 | b[7];
  assign f_arrdiv16_fs8_xor1 = f_arrdiv16_fs7_or0 ^ b[8];
  assign f_arrdiv16_fs8_not1 = ~b[8];
  assign f_arrdiv16_fs8_and1 = f_arrdiv16_fs8_not1 & f_arrdiv16_fs7_or0;
  assign f_arrdiv16_fs8_or0 = f_arrdiv16_fs8_and1 | b[8];
  assign f_arrdiv16_fs9_xor1 = f_arrdiv16_fs8_or0 ^ b[9];
  assign f_arrdiv16_fs9_not1 = ~b[9];
  assign f_arrdiv16_fs9_and1 = f_arrdiv16_fs9_not1 & f_arrdiv16_fs8_or0;
  assign f_arrdiv16_fs9_or0 = f_arrdiv16_fs9_and1 | b[9];
  assign f_arrdiv16_fs10_xor1 = f_arrdiv16_fs9_or0 ^ b[10];
  assign f_arrdiv16_fs10_not1 = ~b[10];
  assign f_arrdiv16_fs10_and1 = f_arrdiv16_fs10_not1 & f_arrdiv16_fs9_or0;
  assign f_arrdiv16_fs10_or0 = f_arrdiv16_fs10_and1 | b[10];
  assign f_arrdiv16_fs11_xor1 = f_arrdiv16_fs10_or0 ^ b[11];
  assign f_arrdiv16_fs11_not1 = ~b[11];
  assign f_arrdiv16_fs11_and1 = f_arrdiv16_fs11_not1 & f_arrdiv16_fs10_or0;
  assign f_arrdiv16_fs11_or0 = f_arrdiv16_fs11_and1 | b[11];
  assign f_arrdiv16_fs12_xor1 = f_arrdiv16_fs11_or0 ^ b[12];
  assign f_arrdiv16_fs12_not1 = ~b[12];
  assign f_arrdiv16_fs12_and1 = f_arrdiv16_fs12_not1 & f_arrdiv16_fs11_or0;
  assign f_arrdiv16_fs12_or0 = f_arrdiv16_fs12_and1 | b[12];
  assign f_arrdiv16_fs13_xor1 = f_arrdiv16_fs12_or0 ^ b[13];
  assign f_arrdiv16_fs13_not1 = ~b[13];
  assign f_arrdiv16_fs13_and1 = f_arrdiv16_fs13_not1 & f_arrdiv16_fs12_or0;
  assign f_arrdiv16_fs13_or0 = f_arrdiv16_fs13_and1 | b[13];
  assign f_arrdiv16_fs14_xor1 = f_arrdiv16_fs13_or0 ^ b[14];
  assign f_arrdiv16_fs14_not1 = ~b[14];
  assign f_arrdiv16_fs14_and1 = f_arrdiv16_fs14_not1 & f_arrdiv16_fs13_or0;
  assign f_arrdiv16_fs14_or0 = f_arrdiv16_fs14_and1 | b[14];
  assign f_arrdiv16_fs15_xor1 = f_arrdiv16_fs14_or0 ^ b[15];
  assign f_arrdiv16_fs15_not1 = ~b[15];
  assign f_arrdiv16_fs15_and1 = f_arrdiv16_fs15_not1 & f_arrdiv16_fs14_or0;
  assign f_arrdiv16_fs15_or0 = f_arrdiv16_fs15_and1 | b[15];
  assign f_arrdiv16_mux2to10_and0 = a[15] & f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to10_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to10_and1 = f_arrdiv16_fs0_xor0 & f_arrdiv16_mux2to10_not0;
  assign f_arrdiv16_mux2to10_xor0 = f_arrdiv16_mux2to10_and0 ^ f_arrdiv16_mux2to10_and1;
  assign f_arrdiv16_mux2to11_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to11_and1 = f_arrdiv16_fs1_xor1 & f_arrdiv16_mux2to11_not0;
  assign f_arrdiv16_mux2to12_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to12_and1 = f_arrdiv16_fs2_xor1 & f_arrdiv16_mux2to12_not0;
  assign f_arrdiv16_mux2to13_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to13_and1 = f_arrdiv16_fs3_xor1 & f_arrdiv16_mux2to13_not0;
  assign f_arrdiv16_mux2to14_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to14_and1 = f_arrdiv16_fs4_xor1 & f_arrdiv16_mux2to14_not0;
  assign f_arrdiv16_mux2to15_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to15_and1 = f_arrdiv16_fs5_xor1 & f_arrdiv16_mux2to15_not0;
  assign f_arrdiv16_mux2to16_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to16_and1 = f_arrdiv16_fs6_xor1 & f_arrdiv16_mux2to16_not0;
  assign f_arrdiv16_mux2to17_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to17_and1 = f_arrdiv16_fs7_xor1 & f_arrdiv16_mux2to17_not0;
  assign f_arrdiv16_mux2to18_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to18_and1 = f_arrdiv16_fs8_xor1 & f_arrdiv16_mux2to18_not0;
  assign f_arrdiv16_mux2to19_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to19_and1 = f_arrdiv16_fs9_xor1 & f_arrdiv16_mux2to19_not0;
  assign f_arrdiv16_mux2to110_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to110_and1 = f_arrdiv16_fs10_xor1 & f_arrdiv16_mux2to110_not0;
  assign f_arrdiv16_mux2to111_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to111_and1 = f_arrdiv16_fs11_xor1 & f_arrdiv16_mux2to111_not0;
  assign f_arrdiv16_mux2to112_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to112_and1 = f_arrdiv16_fs12_xor1 & f_arrdiv16_mux2to112_not0;
  assign f_arrdiv16_mux2to113_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to113_and1 = f_arrdiv16_fs13_xor1 & f_arrdiv16_mux2to113_not0;
  assign f_arrdiv16_mux2to114_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_mux2to114_and1 = f_arrdiv16_fs14_xor1 & f_arrdiv16_mux2to114_not0;
  assign f_arrdiv16_not0 = ~f_arrdiv16_fs15_or0;
  assign f_arrdiv16_fs16_xor0 = a[14] ^ b[0];
  assign f_arrdiv16_fs16_not0 = ~a[14];
  assign f_arrdiv16_fs16_and0 = f_arrdiv16_fs16_not0 & b[0];
  assign f_arrdiv16_fs16_not1 = ~f_arrdiv16_fs16_xor0;
  assign f_arrdiv16_fs17_xor0 = f_arrdiv16_mux2to10_xor0 ^ b[1];
  assign f_arrdiv16_fs17_not0 = ~f_arrdiv16_mux2to10_xor0;
  assign f_arrdiv16_fs17_and0 = f_arrdiv16_fs17_not0 & b[1];
  assign f_arrdiv16_fs17_xor1 = f_arrdiv16_fs16_and0 ^ f_arrdiv16_fs17_xor0;
  assign f_arrdiv16_fs17_not1 = ~f_arrdiv16_fs17_xor0;
  assign f_arrdiv16_fs17_and1 = f_arrdiv16_fs17_not1 & f_arrdiv16_fs16_and0;
  assign f_arrdiv16_fs17_or0 = f_arrdiv16_fs17_and1 | f_arrdiv16_fs17_and0;
  assign f_arrdiv16_fs18_xor0 = f_arrdiv16_mux2to11_and1 ^ b[2];
  assign f_arrdiv16_fs18_not0 = ~f_arrdiv16_mux2to11_and1;
  assign f_arrdiv16_fs18_and0 = f_arrdiv16_fs18_not0 & b[2];
  assign f_arrdiv16_fs18_xor1 = f_arrdiv16_fs17_or0 ^ f_arrdiv16_fs18_xor0;
  assign f_arrdiv16_fs18_not1 = ~f_arrdiv16_fs18_xor0;
  assign f_arrdiv16_fs18_and1 = f_arrdiv16_fs18_not1 & f_arrdiv16_fs17_or0;
  assign f_arrdiv16_fs18_or0 = f_arrdiv16_fs18_and1 | f_arrdiv16_fs18_and0;
  assign f_arrdiv16_fs19_xor0 = f_arrdiv16_mux2to12_and1 ^ b[3];
  assign f_arrdiv16_fs19_not0 = ~f_arrdiv16_mux2to12_and1;
  assign f_arrdiv16_fs19_and0 = f_arrdiv16_fs19_not0 & b[3];
  assign f_arrdiv16_fs19_xor1 = f_arrdiv16_fs18_or0 ^ f_arrdiv16_fs19_xor0;
  assign f_arrdiv16_fs19_not1 = ~f_arrdiv16_fs19_xor0;
  assign f_arrdiv16_fs19_and1 = f_arrdiv16_fs19_not1 & f_arrdiv16_fs18_or0;
  assign f_arrdiv16_fs19_or0 = f_arrdiv16_fs19_and1 | f_arrdiv16_fs19_and0;
  assign f_arrdiv16_fs20_xor0 = f_arrdiv16_mux2to13_and1 ^ b[4];
  assign f_arrdiv16_fs20_not0 = ~f_arrdiv16_mux2to13_and1;
  assign f_arrdiv16_fs20_and0 = f_arrdiv16_fs20_not0 & b[4];
  assign f_arrdiv16_fs20_xor1 = f_arrdiv16_fs19_or0 ^ f_arrdiv16_fs20_xor0;
  assign f_arrdiv16_fs20_not1 = ~f_arrdiv16_fs20_xor0;
  assign f_arrdiv16_fs20_and1 = f_arrdiv16_fs20_not1 & f_arrdiv16_fs19_or0;
  assign f_arrdiv16_fs20_or0 = f_arrdiv16_fs20_and1 | f_arrdiv16_fs20_and0;
  assign f_arrdiv16_fs21_xor0 = f_arrdiv16_mux2to14_and1 ^ b[5];
  assign f_arrdiv16_fs21_not0 = ~f_arrdiv16_mux2to14_and1;
  assign f_arrdiv16_fs21_and0 = f_arrdiv16_fs21_not0 & b[5];
  assign f_arrdiv16_fs21_xor1 = f_arrdiv16_fs20_or0 ^ f_arrdiv16_fs21_xor0;
  assign f_arrdiv16_fs21_not1 = ~f_arrdiv16_fs21_xor0;
  assign f_arrdiv16_fs21_and1 = f_arrdiv16_fs21_not1 & f_arrdiv16_fs20_or0;
  assign f_arrdiv16_fs21_or0 = f_arrdiv16_fs21_and1 | f_arrdiv16_fs21_and0;
  assign f_arrdiv16_fs22_xor0 = f_arrdiv16_mux2to15_and1 ^ b[6];
  assign f_arrdiv16_fs22_not0 = ~f_arrdiv16_mux2to15_and1;
  assign f_arrdiv16_fs22_and0 = f_arrdiv16_fs22_not0 & b[6];
  assign f_arrdiv16_fs22_xor1 = f_arrdiv16_fs21_or0 ^ f_arrdiv16_fs22_xor0;
  assign f_arrdiv16_fs22_not1 = ~f_arrdiv16_fs22_xor0;
  assign f_arrdiv16_fs22_and1 = f_arrdiv16_fs22_not1 & f_arrdiv16_fs21_or0;
  assign f_arrdiv16_fs22_or0 = f_arrdiv16_fs22_and1 | f_arrdiv16_fs22_and0;
  assign f_arrdiv16_fs23_xor0 = f_arrdiv16_mux2to16_and1 ^ b[7];
  assign f_arrdiv16_fs23_not0 = ~f_arrdiv16_mux2to16_and1;
  assign f_arrdiv16_fs23_and0 = f_arrdiv16_fs23_not0 & b[7];
  assign f_arrdiv16_fs23_xor1 = f_arrdiv16_fs22_or0 ^ f_arrdiv16_fs23_xor0;
  assign f_arrdiv16_fs23_not1 = ~f_arrdiv16_fs23_xor0;
  assign f_arrdiv16_fs23_and1 = f_arrdiv16_fs23_not1 & f_arrdiv16_fs22_or0;
  assign f_arrdiv16_fs23_or0 = f_arrdiv16_fs23_and1 | f_arrdiv16_fs23_and0;
  assign f_arrdiv16_fs24_xor0 = f_arrdiv16_mux2to17_and1 ^ b[8];
  assign f_arrdiv16_fs24_not0 = ~f_arrdiv16_mux2to17_and1;
  assign f_arrdiv16_fs24_and0 = f_arrdiv16_fs24_not0 & b[8];
  assign f_arrdiv16_fs24_xor1 = f_arrdiv16_fs23_or0 ^ f_arrdiv16_fs24_xor0;
  assign f_arrdiv16_fs24_not1 = ~f_arrdiv16_fs24_xor0;
  assign f_arrdiv16_fs24_and1 = f_arrdiv16_fs24_not1 & f_arrdiv16_fs23_or0;
  assign f_arrdiv16_fs24_or0 = f_arrdiv16_fs24_and1 | f_arrdiv16_fs24_and0;
  assign f_arrdiv16_fs25_xor0 = f_arrdiv16_mux2to18_and1 ^ b[9];
  assign f_arrdiv16_fs25_not0 = ~f_arrdiv16_mux2to18_and1;
  assign f_arrdiv16_fs25_and0 = f_arrdiv16_fs25_not0 & b[9];
  assign f_arrdiv16_fs25_xor1 = f_arrdiv16_fs24_or0 ^ f_arrdiv16_fs25_xor0;
  assign f_arrdiv16_fs25_not1 = ~f_arrdiv16_fs25_xor0;
  assign f_arrdiv16_fs25_and1 = f_arrdiv16_fs25_not1 & f_arrdiv16_fs24_or0;
  assign f_arrdiv16_fs25_or0 = f_arrdiv16_fs25_and1 | f_arrdiv16_fs25_and0;
  assign f_arrdiv16_fs26_xor0 = f_arrdiv16_mux2to19_and1 ^ b[10];
  assign f_arrdiv16_fs26_not0 = ~f_arrdiv16_mux2to19_and1;
  assign f_arrdiv16_fs26_and0 = f_arrdiv16_fs26_not0 & b[10];
  assign f_arrdiv16_fs26_xor1 = f_arrdiv16_fs25_or0 ^ f_arrdiv16_fs26_xor0;
  assign f_arrdiv16_fs26_not1 = ~f_arrdiv16_fs26_xor0;
  assign f_arrdiv16_fs26_and1 = f_arrdiv16_fs26_not1 & f_arrdiv16_fs25_or0;
  assign f_arrdiv16_fs26_or0 = f_arrdiv16_fs26_and1 | f_arrdiv16_fs26_and0;
  assign f_arrdiv16_fs27_xor0 = f_arrdiv16_mux2to110_and1 ^ b[11];
  assign f_arrdiv16_fs27_not0 = ~f_arrdiv16_mux2to110_and1;
  assign f_arrdiv16_fs27_and0 = f_arrdiv16_fs27_not0 & b[11];
  assign f_arrdiv16_fs27_xor1 = f_arrdiv16_fs26_or0 ^ f_arrdiv16_fs27_xor0;
  assign f_arrdiv16_fs27_not1 = ~f_arrdiv16_fs27_xor0;
  assign f_arrdiv16_fs27_and1 = f_arrdiv16_fs27_not1 & f_arrdiv16_fs26_or0;
  assign f_arrdiv16_fs27_or0 = f_arrdiv16_fs27_and1 | f_arrdiv16_fs27_and0;
  assign f_arrdiv16_fs28_xor0 = f_arrdiv16_mux2to111_and1 ^ b[12];
  assign f_arrdiv16_fs28_not0 = ~f_arrdiv16_mux2to111_and1;
  assign f_arrdiv16_fs28_and0 = f_arrdiv16_fs28_not0 & b[12];
  assign f_arrdiv16_fs28_xor1 = f_arrdiv16_fs27_or0 ^ f_arrdiv16_fs28_xor0;
  assign f_arrdiv16_fs28_not1 = ~f_arrdiv16_fs28_xor0;
  assign f_arrdiv16_fs28_and1 = f_arrdiv16_fs28_not1 & f_arrdiv16_fs27_or0;
  assign f_arrdiv16_fs28_or0 = f_arrdiv16_fs28_and1 | f_arrdiv16_fs28_and0;
  assign f_arrdiv16_fs29_xor0 = f_arrdiv16_mux2to112_and1 ^ b[13];
  assign f_arrdiv16_fs29_not0 = ~f_arrdiv16_mux2to112_and1;
  assign f_arrdiv16_fs29_and0 = f_arrdiv16_fs29_not0 & b[13];
  assign f_arrdiv16_fs29_xor1 = f_arrdiv16_fs28_or0 ^ f_arrdiv16_fs29_xor0;
  assign f_arrdiv16_fs29_not1 = ~f_arrdiv16_fs29_xor0;
  assign f_arrdiv16_fs29_and1 = f_arrdiv16_fs29_not1 & f_arrdiv16_fs28_or0;
  assign f_arrdiv16_fs29_or0 = f_arrdiv16_fs29_and1 | f_arrdiv16_fs29_and0;
  assign f_arrdiv16_fs30_xor0 = f_arrdiv16_mux2to113_and1 ^ b[14];
  assign f_arrdiv16_fs30_not0 = ~f_arrdiv16_mux2to113_and1;
  assign f_arrdiv16_fs30_and0 = f_arrdiv16_fs30_not0 & b[14];
  assign f_arrdiv16_fs30_xor1 = f_arrdiv16_fs29_or0 ^ f_arrdiv16_fs30_xor0;
  assign f_arrdiv16_fs30_not1 = ~f_arrdiv16_fs30_xor0;
  assign f_arrdiv16_fs30_and1 = f_arrdiv16_fs30_not1 & f_arrdiv16_fs29_or0;
  assign f_arrdiv16_fs30_or0 = f_arrdiv16_fs30_and1 | f_arrdiv16_fs30_and0;
  assign f_arrdiv16_fs31_xor0 = f_arrdiv16_mux2to114_and1 ^ b[15];
  assign f_arrdiv16_fs31_not0 = ~f_arrdiv16_mux2to114_and1;
  assign f_arrdiv16_fs31_and0 = f_arrdiv16_fs31_not0 & b[15];
  assign f_arrdiv16_fs31_xor1 = f_arrdiv16_fs30_or0 ^ f_arrdiv16_fs31_xor0;
  assign f_arrdiv16_fs31_not1 = ~f_arrdiv16_fs31_xor0;
  assign f_arrdiv16_fs31_and1 = f_arrdiv16_fs31_not1 & f_arrdiv16_fs30_or0;
  assign f_arrdiv16_fs31_or0 = f_arrdiv16_fs31_and1 | f_arrdiv16_fs31_and0;
  assign f_arrdiv16_mux2to115_and0 = a[14] & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to115_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to115_and1 = f_arrdiv16_fs16_xor0 & f_arrdiv16_mux2to115_not0;
  assign f_arrdiv16_mux2to115_xor0 = f_arrdiv16_mux2to115_and0 ^ f_arrdiv16_mux2to115_and1;
  assign f_arrdiv16_mux2to116_and0 = f_arrdiv16_mux2to10_xor0 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to116_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to116_and1 = f_arrdiv16_fs17_xor1 & f_arrdiv16_mux2to116_not0;
  assign f_arrdiv16_mux2to116_xor0 = f_arrdiv16_mux2to116_and0 ^ f_arrdiv16_mux2to116_and1;
  assign f_arrdiv16_mux2to117_and0 = f_arrdiv16_mux2to11_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to117_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to117_and1 = f_arrdiv16_fs18_xor1 & f_arrdiv16_mux2to117_not0;
  assign f_arrdiv16_mux2to117_xor0 = f_arrdiv16_mux2to117_and0 ^ f_arrdiv16_mux2to117_and1;
  assign f_arrdiv16_mux2to118_and0 = f_arrdiv16_mux2to12_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to118_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to118_and1 = f_arrdiv16_fs19_xor1 & f_arrdiv16_mux2to118_not0;
  assign f_arrdiv16_mux2to118_xor0 = f_arrdiv16_mux2to118_and0 ^ f_arrdiv16_mux2to118_and1;
  assign f_arrdiv16_mux2to119_and0 = f_arrdiv16_mux2to13_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to119_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to119_and1 = f_arrdiv16_fs20_xor1 & f_arrdiv16_mux2to119_not0;
  assign f_arrdiv16_mux2to119_xor0 = f_arrdiv16_mux2to119_and0 ^ f_arrdiv16_mux2to119_and1;
  assign f_arrdiv16_mux2to120_and0 = f_arrdiv16_mux2to14_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to120_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to120_and1 = f_arrdiv16_fs21_xor1 & f_arrdiv16_mux2to120_not0;
  assign f_arrdiv16_mux2to120_xor0 = f_arrdiv16_mux2to120_and0 ^ f_arrdiv16_mux2to120_and1;
  assign f_arrdiv16_mux2to121_and0 = f_arrdiv16_mux2to15_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to121_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to121_and1 = f_arrdiv16_fs22_xor1 & f_arrdiv16_mux2to121_not0;
  assign f_arrdiv16_mux2to121_xor0 = f_arrdiv16_mux2to121_and0 ^ f_arrdiv16_mux2to121_and1;
  assign f_arrdiv16_mux2to122_and0 = f_arrdiv16_mux2to16_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to122_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to122_and1 = f_arrdiv16_fs23_xor1 & f_arrdiv16_mux2to122_not0;
  assign f_arrdiv16_mux2to122_xor0 = f_arrdiv16_mux2to122_and0 ^ f_arrdiv16_mux2to122_and1;
  assign f_arrdiv16_mux2to123_and0 = f_arrdiv16_mux2to17_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to123_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to123_and1 = f_arrdiv16_fs24_xor1 & f_arrdiv16_mux2to123_not0;
  assign f_arrdiv16_mux2to123_xor0 = f_arrdiv16_mux2to123_and0 ^ f_arrdiv16_mux2to123_and1;
  assign f_arrdiv16_mux2to124_and0 = f_arrdiv16_mux2to18_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to124_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to124_and1 = f_arrdiv16_fs25_xor1 & f_arrdiv16_mux2to124_not0;
  assign f_arrdiv16_mux2to124_xor0 = f_arrdiv16_mux2to124_and0 ^ f_arrdiv16_mux2to124_and1;
  assign f_arrdiv16_mux2to125_and0 = f_arrdiv16_mux2to19_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to125_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to125_and1 = f_arrdiv16_fs26_xor1 & f_arrdiv16_mux2to125_not0;
  assign f_arrdiv16_mux2to125_xor0 = f_arrdiv16_mux2to125_and0 ^ f_arrdiv16_mux2to125_and1;
  assign f_arrdiv16_mux2to126_and0 = f_arrdiv16_mux2to110_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to126_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to126_and1 = f_arrdiv16_fs27_xor1 & f_arrdiv16_mux2to126_not0;
  assign f_arrdiv16_mux2to126_xor0 = f_arrdiv16_mux2to126_and0 ^ f_arrdiv16_mux2to126_and1;
  assign f_arrdiv16_mux2to127_and0 = f_arrdiv16_mux2to111_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to127_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to127_and1 = f_arrdiv16_fs28_xor1 & f_arrdiv16_mux2to127_not0;
  assign f_arrdiv16_mux2to127_xor0 = f_arrdiv16_mux2to127_and0 ^ f_arrdiv16_mux2to127_and1;
  assign f_arrdiv16_mux2to128_and0 = f_arrdiv16_mux2to112_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to128_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to128_and1 = f_arrdiv16_fs29_xor1 & f_arrdiv16_mux2to128_not0;
  assign f_arrdiv16_mux2to128_xor0 = f_arrdiv16_mux2to128_and0 ^ f_arrdiv16_mux2to128_and1;
  assign f_arrdiv16_mux2to129_and0 = f_arrdiv16_mux2to113_and1 & f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to129_not0 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_mux2to129_and1 = f_arrdiv16_fs30_xor1 & f_arrdiv16_mux2to129_not0;
  assign f_arrdiv16_mux2to129_xor0 = f_arrdiv16_mux2to129_and0 ^ f_arrdiv16_mux2to129_and1;
  assign f_arrdiv16_not1 = ~f_arrdiv16_fs31_or0;
  assign f_arrdiv16_fs32_xor0 = a[13] ^ b[0];
  assign f_arrdiv16_fs32_not0 = ~a[13];
  assign f_arrdiv16_fs32_and0 = f_arrdiv16_fs32_not0 & b[0];
  assign f_arrdiv16_fs32_not1 = ~f_arrdiv16_fs32_xor0;
  assign f_arrdiv16_fs33_xor0 = f_arrdiv16_mux2to115_xor0 ^ b[1];
  assign f_arrdiv16_fs33_not0 = ~f_arrdiv16_mux2to115_xor0;
  assign f_arrdiv16_fs33_and0 = f_arrdiv16_fs33_not0 & b[1];
  assign f_arrdiv16_fs33_xor1 = f_arrdiv16_fs32_and0 ^ f_arrdiv16_fs33_xor0;
  assign f_arrdiv16_fs33_not1 = ~f_arrdiv16_fs33_xor0;
  assign f_arrdiv16_fs33_and1 = f_arrdiv16_fs33_not1 & f_arrdiv16_fs32_and0;
  assign f_arrdiv16_fs33_or0 = f_arrdiv16_fs33_and1 | f_arrdiv16_fs33_and0;
  assign f_arrdiv16_fs34_xor0 = f_arrdiv16_mux2to116_xor0 ^ b[2];
  assign f_arrdiv16_fs34_not0 = ~f_arrdiv16_mux2to116_xor0;
  assign f_arrdiv16_fs34_and0 = f_arrdiv16_fs34_not0 & b[2];
  assign f_arrdiv16_fs34_xor1 = f_arrdiv16_fs33_or0 ^ f_arrdiv16_fs34_xor0;
  assign f_arrdiv16_fs34_not1 = ~f_arrdiv16_fs34_xor0;
  assign f_arrdiv16_fs34_and1 = f_arrdiv16_fs34_not1 & f_arrdiv16_fs33_or0;
  assign f_arrdiv16_fs34_or0 = f_arrdiv16_fs34_and1 | f_arrdiv16_fs34_and0;
  assign f_arrdiv16_fs35_xor0 = f_arrdiv16_mux2to117_xor0 ^ b[3];
  assign f_arrdiv16_fs35_not0 = ~f_arrdiv16_mux2to117_xor0;
  assign f_arrdiv16_fs35_and0 = f_arrdiv16_fs35_not0 & b[3];
  assign f_arrdiv16_fs35_xor1 = f_arrdiv16_fs34_or0 ^ f_arrdiv16_fs35_xor0;
  assign f_arrdiv16_fs35_not1 = ~f_arrdiv16_fs35_xor0;
  assign f_arrdiv16_fs35_and1 = f_arrdiv16_fs35_not1 & f_arrdiv16_fs34_or0;
  assign f_arrdiv16_fs35_or0 = f_arrdiv16_fs35_and1 | f_arrdiv16_fs35_and0;
  assign f_arrdiv16_fs36_xor0 = f_arrdiv16_mux2to118_xor0 ^ b[4];
  assign f_arrdiv16_fs36_not0 = ~f_arrdiv16_mux2to118_xor0;
  assign f_arrdiv16_fs36_and0 = f_arrdiv16_fs36_not0 & b[4];
  assign f_arrdiv16_fs36_xor1 = f_arrdiv16_fs35_or0 ^ f_arrdiv16_fs36_xor0;
  assign f_arrdiv16_fs36_not1 = ~f_arrdiv16_fs36_xor0;
  assign f_arrdiv16_fs36_and1 = f_arrdiv16_fs36_not1 & f_arrdiv16_fs35_or0;
  assign f_arrdiv16_fs36_or0 = f_arrdiv16_fs36_and1 | f_arrdiv16_fs36_and0;
  assign f_arrdiv16_fs37_xor0 = f_arrdiv16_mux2to119_xor0 ^ b[5];
  assign f_arrdiv16_fs37_not0 = ~f_arrdiv16_mux2to119_xor0;
  assign f_arrdiv16_fs37_and0 = f_arrdiv16_fs37_not0 & b[5];
  assign f_arrdiv16_fs37_xor1 = f_arrdiv16_fs36_or0 ^ f_arrdiv16_fs37_xor0;
  assign f_arrdiv16_fs37_not1 = ~f_arrdiv16_fs37_xor0;
  assign f_arrdiv16_fs37_and1 = f_arrdiv16_fs37_not1 & f_arrdiv16_fs36_or0;
  assign f_arrdiv16_fs37_or0 = f_arrdiv16_fs37_and1 | f_arrdiv16_fs37_and0;
  assign f_arrdiv16_fs38_xor0 = f_arrdiv16_mux2to120_xor0 ^ b[6];
  assign f_arrdiv16_fs38_not0 = ~f_arrdiv16_mux2to120_xor0;
  assign f_arrdiv16_fs38_and0 = f_arrdiv16_fs38_not0 & b[6];
  assign f_arrdiv16_fs38_xor1 = f_arrdiv16_fs37_or0 ^ f_arrdiv16_fs38_xor0;
  assign f_arrdiv16_fs38_not1 = ~f_arrdiv16_fs38_xor0;
  assign f_arrdiv16_fs38_and1 = f_arrdiv16_fs38_not1 & f_arrdiv16_fs37_or0;
  assign f_arrdiv16_fs38_or0 = f_arrdiv16_fs38_and1 | f_arrdiv16_fs38_and0;
  assign f_arrdiv16_fs39_xor0 = f_arrdiv16_mux2to121_xor0 ^ b[7];
  assign f_arrdiv16_fs39_not0 = ~f_arrdiv16_mux2to121_xor0;
  assign f_arrdiv16_fs39_and0 = f_arrdiv16_fs39_not0 & b[7];
  assign f_arrdiv16_fs39_xor1 = f_arrdiv16_fs38_or0 ^ f_arrdiv16_fs39_xor0;
  assign f_arrdiv16_fs39_not1 = ~f_arrdiv16_fs39_xor0;
  assign f_arrdiv16_fs39_and1 = f_arrdiv16_fs39_not1 & f_arrdiv16_fs38_or0;
  assign f_arrdiv16_fs39_or0 = f_arrdiv16_fs39_and1 | f_arrdiv16_fs39_and0;
  assign f_arrdiv16_fs40_xor0 = f_arrdiv16_mux2to122_xor0 ^ b[8];
  assign f_arrdiv16_fs40_not0 = ~f_arrdiv16_mux2to122_xor0;
  assign f_arrdiv16_fs40_and0 = f_arrdiv16_fs40_not0 & b[8];
  assign f_arrdiv16_fs40_xor1 = f_arrdiv16_fs39_or0 ^ f_arrdiv16_fs40_xor0;
  assign f_arrdiv16_fs40_not1 = ~f_arrdiv16_fs40_xor0;
  assign f_arrdiv16_fs40_and1 = f_arrdiv16_fs40_not1 & f_arrdiv16_fs39_or0;
  assign f_arrdiv16_fs40_or0 = f_arrdiv16_fs40_and1 | f_arrdiv16_fs40_and0;
  assign f_arrdiv16_fs41_xor0 = f_arrdiv16_mux2to123_xor0 ^ b[9];
  assign f_arrdiv16_fs41_not0 = ~f_arrdiv16_mux2to123_xor0;
  assign f_arrdiv16_fs41_and0 = f_arrdiv16_fs41_not0 & b[9];
  assign f_arrdiv16_fs41_xor1 = f_arrdiv16_fs40_or0 ^ f_arrdiv16_fs41_xor0;
  assign f_arrdiv16_fs41_not1 = ~f_arrdiv16_fs41_xor0;
  assign f_arrdiv16_fs41_and1 = f_arrdiv16_fs41_not1 & f_arrdiv16_fs40_or0;
  assign f_arrdiv16_fs41_or0 = f_arrdiv16_fs41_and1 | f_arrdiv16_fs41_and0;
  assign f_arrdiv16_fs42_xor0 = f_arrdiv16_mux2to124_xor0 ^ b[10];
  assign f_arrdiv16_fs42_not0 = ~f_arrdiv16_mux2to124_xor0;
  assign f_arrdiv16_fs42_and0 = f_arrdiv16_fs42_not0 & b[10];
  assign f_arrdiv16_fs42_xor1 = f_arrdiv16_fs41_or0 ^ f_arrdiv16_fs42_xor0;
  assign f_arrdiv16_fs42_not1 = ~f_arrdiv16_fs42_xor0;
  assign f_arrdiv16_fs42_and1 = f_arrdiv16_fs42_not1 & f_arrdiv16_fs41_or0;
  assign f_arrdiv16_fs42_or0 = f_arrdiv16_fs42_and1 | f_arrdiv16_fs42_and0;
  assign f_arrdiv16_fs43_xor0 = f_arrdiv16_mux2to125_xor0 ^ b[11];
  assign f_arrdiv16_fs43_not0 = ~f_arrdiv16_mux2to125_xor0;
  assign f_arrdiv16_fs43_and0 = f_arrdiv16_fs43_not0 & b[11];
  assign f_arrdiv16_fs43_xor1 = f_arrdiv16_fs42_or0 ^ f_arrdiv16_fs43_xor0;
  assign f_arrdiv16_fs43_not1 = ~f_arrdiv16_fs43_xor0;
  assign f_arrdiv16_fs43_and1 = f_arrdiv16_fs43_not1 & f_arrdiv16_fs42_or0;
  assign f_arrdiv16_fs43_or0 = f_arrdiv16_fs43_and1 | f_arrdiv16_fs43_and0;
  assign f_arrdiv16_fs44_xor0 = f_arrdiv16_mux2to126_xor0 ^ b[12];
  assign f_arrdiv16_fs44_not0 = ~f_arrdiv16_mux2to126_xor0;
  assign f_arrdiv16_fs44_and0 = f_arrdiv16_fs44_not0 & b[12];
  assign f_arrdiv16_fs44_xor1 = f_arrdiv16_fs43_or0 ^ f_arrdiv16_fs44_xor0;
  assign f_arrdiv16_fs44_not1 = ~f_arrdiv16_fs44_xor0;
  assign f_arrdiv16_fs44_and1 = f_arrdiv16_fs44_not1 & f_arrdiv16_fs43_or0;
  assign f_arrdiv16_fs44_or0 = f_arrdiv16_fs44_and1 | f_arrdiv16_fs44_and0;
  assign f_arrdiv16_fs45_xor0 = f_arrdiv16_mux2to127_xor0 ^ b[13];
  assign f_arrdiv16_fs45_not0 = ~f_arrdiv16_mux2to127_xor0;
  assign f_arrdiv16_fs45_and0 = f_arrdiv16_fs45_not0 & b[13];
  assign f_arrdiv16_fs45_xor1 = f_arrdiv16_fs44_or0 ^ f_arrdiv16_fs45_xor0;
  assign f_arrdiv16_fs45_not1 = ~f_arrdiv16_fs45_xor0;
  assign f_arrdiv16_fs45_and1 = f_arrdiv16_fs45_not1 & f_arrdiv16_fs44_or0;
  assign f_arrdiv16_fs45_or0 = f_arrdiv16_fs45_and1 | f_arrdiv16_fs45_and0;
  assign f_arrdiv16_fs46_xor0 = f_arrdiv16_mux2to128_xor0 ^ b[14];
  assign f_arrdiv16_fs46_not0 = ~f_arrdiv16_mux2to128_xor0;
  assign f_arrdiv16_fs46_and0 = f_arrdiv16_fs46_not0 & b[14];
  assign f_arrdiv16_fs46_xor1 = f_arrdiv16_fs45_or0 ^ f_arrdiv16_fs46_xor0;
  assign f_arrdiv16_fs46_not1 = ~f_arrdiv16_fs46_xor0;
  assign f_arrdiv16_fs46_and1 = f_arrdiv16_fs46_not1 & f_arrdiv16_fs45_or0;
  assign f_arrdiv16_fs46_or0 = f_arrdiv16_fs46_and1 | f_arrdiv16_fs46_and0;
  assign f_arrdiv16_fs47_xor0 = f_arrdiv16_mux2to129_xor0 ^ b[15];
  assign f_arrdiv16_fs47_not0 = ~f_arrdiv16_mux2to129_xor0;
  assign f_arrdiv16_fs47_and0 = f_arrdiv16_fs47_not0 & b[15];
  assign f_arrdiv16_fs47_xor1 = f_arrdiv16_fs46_or0 ^ f_arrdiv16_fs47_xor0;
  assign f_arrdiv16_fs47_not1 = ~f_arrdiv16_fs47_xor0;
  assign f_arrdiv16_fs47_and1 = f_arrdiv16_fs47_not1 & f_arrdiv16_fs46_or0;
  assign f_arrdiv16_fs47_or0 = f_arrdiv16_fs47_and1 | f_arrdiv16_fs47_and0;
  assign f_arrdiv16_mux2to130_and0 = a[13] & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to130_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to130_and1 = f_arrdiv16_fs32_xor0 & f_arrdiv16_mux2to130_not0;
  assign f_arrdiv16_mux2to130_xor0 = f_arrdiv16_mux2to130_and0 ^ f_arrdiv16_mux2to130_and1;
  assign f_arrdiv16_mux2to131_and0 = f_arrdiv16_mux2to115_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to131_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to131_and1 = f_arrdiv16_fs33_xor1 & f_arrdiv16_mux2to131_not0;
  assign f_arrdiv16_mux2to131_xor0 = f_arrdiv16_mux2to131_and0 ^ f_arrdiv16_mux2to131_and1;
  assign f_arrdiv16_mux2to132_and0 = f_arrdiv16_mux2to116_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to132_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to132_and1 = f_arrdiv16_fs34_xor1 & f_arrdiv16_mux2to132_not0;
  assign f_arrdiv16_mux2to132_xor0 = f_arrdiv16_mux2to132_and0 ^ f_arrdiv16_mux2to132_and1;
  assign f_arrdiv16_mux2to133_and0 = f_arrdiv16_mux2to117_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to133_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to133_and1 = f_arrdiv16_fs35_xor1 & f_arrdiv16_mux2to133_not0;
  assign f_arrdiv16_mux2to133_xor0 = f_arrdiv16_mux2to133_and0 ^ f_arrdiv16_mux2to133_and1;
  assign f_arrdiv16_mux2to134_and0 = f_arrdiv16_mux2to118_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to134_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to134_and1 = f_arrdiv16_fs36_xor1 & f_arrdiv16_mux2to134_not0;
  assign f_arrdiv16_mux2to134_xor0 = f_arrdiv16_mux2to134_and0 ^ f_arrdiv16_mux2to134_and1;
  assign f_arrdiv16_mux2to135_and0 = f_arrdiv16_mux2to119_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to135_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to135_and1 = f_arrdiv16_fs37_xor1 & f_arrdiv16_mux2to135_not0;
  assign f_arrdiv16_mux2to135_xor0 = f_arrdiv16_mux2to135_and0 ^ f_arrdiv16_mux2to135_and1;
  assign f_arrdiv16_mux2to136_and0 = f_arrdiv16_mux2to120_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to136_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to136_and1 = f_arrdiv16_fs38_xor1 & f_arrdiv16_mux2to136_not0;
  assign f_arrdiv16_mux2to136_xor0 = f_arrdiv16_mux2to136_and0 ^ f_arrdiv16_mux2to136_and1;
  assign f_arrdiv16_mux2to137_and0 = f_arrdiv16_mux2to121_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to137_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to137_and1 = f_arrdiv16_fs39_xor1 & f_arrdiv16_mux2to137_not0;
  assign f_arrdiv16_mux2to137_xor0 = f_arrdiv16_mux2to137_and0 ^ f_arrdiv16_mux2to137_and1;
  assign f_arrdiv16_mux2to138_and0 = f_arrdiv16_mux2to122_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to138_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to138_and1 = f_arrdiv16_fs40_xor1 & f_arrdiv16_mux2to138_not0;
  assign f_arrdiv16_mux2to138_xor0 = f_arrdiv16_mux2to138_and0 ^ f_arrdiv16_mux2to138_and1;
  assign f_arrdiv16_mux2to139_and0 = f_arrdiv16_mux2to123_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to139_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to139_and1 = f_arrdiv16_fs41_xor1 & f_arrdiv16_mux2to139_not0;
  assign f_arrdiv16_mux2to139_xor0 = f_arrdiv16_mux2to139_and0 ^ f_arrdiv16_mux2to139_and1;
  assign f_arrdiv16_mux2to140_and0 = f_arrdiv16_mux2to124_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to140_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to140_and1 = f_arrdiv16_fs42_xor1 & f_arrdiv16_mux2to140_not0;
  assign f_arrdiv16_mux2to140_xor0 = f_arrdiv16_mux2to140_and0 ^ f_arrdiv16_mux2to140_and1;
  assign f_arrdiv16_mux2to141_and0 = f_arrdiv16_mux2to125_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to141_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to141_and1 = f_arrdiv16_fs43_xor1 & f_arrdiv16_mux2to141_not0;
  assign f_arrdiv16_mux2to141_xor0 = f_arrdiv16_mux2to141_and0 ^ f_arrdiv16_mux2to141_and1;
  assign f_arrdiv16_mux2to142_and0 = f_arrdiv16_mux2to126_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to142_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to142_and1 = f_arrdiv16_fs44_xor1 & f_arrdiv16_mux2to142_not0;
  assign f_arrdiv16_mux2to142_xor0 = f_arrdiv16_mux2to142_and0 ^ f_arrdiv16_mux2to142_and1;
  assign f_arrdiv16_mux2to143_and0 = f_arrdiv16_mux2to127_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to143_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to143_and1 = f_arrdiv16_fs45_xor1 & f_arrdiv16_mux2to143_not0;
  assign f_arrdiv16_mux2to143_xor0 = f_arrdiv16_mux2to143_and0 ^ f_arrdiv16_mux2to143_and1;
  assign f_arrdiv16_mux2to144_and0 = f_arrdiv16_mux2to128_xor0 & f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to144_not0 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_mux2to144_and1 = f_arrdiv16_fs46_xor1 & f_arrdiv16_mux2to144_not0;
  assign f_arrdiv16_mux2to144_xor0 = f_arrdiv16_mux2to144_and0 ^ f_arrdiv16_mux2to144_and1;
  assign f_arrdiv16_not2 = ~f_arrdiv16_fs47_or0;
  assign f_arrdiv16_fs48_xor0 = a[12] ^ b[0];
  assign f_arrdiv16_fs48_not0 = ~a[12];
  assign f_arrdiv16_fs48_and0 = f_arrdiv16_fs48_not0 & b[0];
  assign f_arrdiv16_fs48_not1 = ~f_arrdiv16_fs48_xor0;
  assign f_arrdiv16_fs49_xor0 = f_arrdiv16_mux2to130_xor0 ^ b[1];
  assign f_arrdiv16_fs49_not0 = ~f_arrdiv16_mux2to130_xor0;
  assign f_arrdiv16_fs49_and0 = f_arrdiv16_fs49_not0 & b[1];
  assign f_arrdiv16_fs49_xor1 = f_arrdiv16_fs48_and0 ^ f_arrdiv16_fs49_xor0;
  assign f_arrdiv16_fs49_not1 = ~f_arrdiv16_fs49_xor0;
  assign f_arrdiv16_fs49_and1 = f_arrdiv16_fs49_not1 & f_arrdiv16_fs48_and0;
  assign f_arrdiv16_fs49_or0 = f_arrdiv16_fs49_and1 | f_arrdiv16_fs49_and0;
  assign f_arrdiv16_fs50_xor0 = f_arrdiv16_mux2to131_xor0 ^ b[2];
  assign f_arrdiv16_fs50_not0 = ~f_arrdiv16_mux2to131_xor0;
  assign f_arrdiv16_fs50_and0 = f_arrdiv16_fs50_not0 & b[2];
  assign f_arrdiv16_fs50_xor1 = f_arrdiv16_fs49_or0 ^ f_arrdiv16_fs50_xor0;
  assign f_arrdiv16_fs50_not1 = ~f_arrdiv16_fs50_xor0;
  assign f_arrdiv16_fs50_and1 = f_arrdiv16_fs50_not1 & f_arrdiv16_fs49_or0;
  assign f_arrdiv16_fs50_or0 = f_arrdiv16_fs50_and1 | f_arrdiv16_fs50_and0;
  assign f_arrdiv16_fs51_xor0 = f_arrdiv16_mux2to132_xor0 ^ b[3];
  assign f_arrdiv16_fs51_not0 = ~f_arrdiv16_mux2to132_xor0;
  assign f_arrdiv16_fs51_and0 = f_arrdiv16_fs51_not0 & b[3];
  assign f_arrdiv16_fs51_xor1 = f_arrdiv16_fs50_or0 ^ f_arrdiv16_fs51_xor0;
  assign f_arrdiv16_fs51_not1 = ~f_arrdiv16_fs51_xor0;
  assign f_arrdiv16_fs51_and1 = f_arrdiv16_fs51_not1 & f_arrdiv16_fs50_or0;
  assign f_arrdiv16_fs51_or0 = f_arrdiv16_fs51_and1 | f_arrdiv16_fs51_and0;
  assign f_arrdiv16_fs52_xor0 = f_arrdiv16_mux2to133_xor0 ^ b[4];
  assign f_arrdiv16_fs52_not0 = ~f_arrdiv16_mux2to133_xor0;
  assign f_arrdiv16_fs52_and0 = f_arrdiv16_fs52_not0 & b[4];
  assign f_arrdiv16_fs52_xor1 = f_arrdiv16_fs51_or0 ^ f_arrdiv16_fs52_xor0;
  assign f_arrdiv16_fs52_not1 = ~f_arrdiv16_fs52_xor0;
  assign f_arrdiv16_fs52_and1 = f_arrdiv16_fs52_not1 & f_arrdiv16_fs51_or0;
  assign f_arrdiv16_fs52_or0 = f_arrdiv16_fs52_and1 | f_arrdiv16_fs52_and0;
  assign f_arrdiv16_fs53_xor0 = f_arrdiv16_mux2to134_xor0 ^ b[5];
  assign f_arrdiv16_fs53_not0 = ~f_arrdiv16_mux2to134_xor0;
  assign f_arrdiv16_fs53_and0 = f_arrdiv16_fs53_not0 & b[5];
  assign f_arrdiv16_fs53_xor1 = f_arrdiv16_fs52_or0 ^ f_arrdiv16_fs53_xor0;
  assign f_arrdiv16_fs53_not1 = ~f_arrdiv16_fs53_xor0;
  assign f_arrdiv16_fs53_and1 = f_arrdiv16_fs53_not1 & f_arrdiv16_fs52_or0;
  assign f_arrdiv16_fs53_or0 = f_arrdiv16_fs53_and1 | f_arrdiv16_fs53_and0;
  assign f_arrdiv16_fs54_xor0 = f_arrdiv16_mux2to135_xor0 ^ b[6];
  assign f_arrdiv16_fs54_not0 = ~f_arrdiv16_mux2to135_xor0;
  assign f_arrdiv16_fs54_and0 = f_arrdiv16_fs54_not0 & b[6];
  assign f_arrdiv16_fs54_xor1 = f_arrdiv16_fs53_or0 ^ f_arrdiv16_fs54_xor0;
  assign f_arrdiv16_fs54_not1 = ~f_arrdiv16_fs54_xor0;
  assign f_arrdiv16_fs54_and1 = f_arrdiv16_fs54_not1 & f_arrdiv16_fs53_or0;
  assign f_arrdiv16_fs54_or0 = f_arrdiv16_fs54_and1 | f_arrdiv16_fs54_and0;
  assign f_arrdiv16_fs55_xor0 = f_arrdiv16_mux2to136_xor0 ^ b[7];
  assign f_arrdiv16_fs55_not0 = ~f_arrdiv16_mux2to136_xor0;
  assign f_arrdiv16_fs55_and0 = f_arrdiv16_fs55_not0 & b[7];
  assign f_arrdiv16_fs55_xor1 = f_arrdiv16_fs54_or0 ^ f_arrdiv16_fs55_xor0;
  assign f_arrdiv16_fs55_not1 = ~f_arrdiv16_fs55_xor0;
  assign f_arrdiv16_fs55_and1 = f_arrdiv16_fs55_not1 & f_arrdiv16_fs54_or0;
  assign f_arrdiv16_fs55_or0 = f_arrdiv16_fs55_and1 | f_arrdiv16_fs55_and0;
  assign f_arrdiv16_fs56_xor0 = f_arrdiv16_mux2to137_xor0 ^ b[8];
  assign f_arrdiv16_fs56_not0 = ~f_arrdiv16_mux2to137_xor0;
  assign f_arrdiv16_fs56_and0 = f_arrdiv16_fs56_not0 & b[8];
  assign f_arrdiv16_fs56_xor1 = f_arrdiv16_fs55_or0 ^ f_arrdiv16_fs56_xor0;
  assign f_arrdiv16_fs56_not1 = ~f_arrdiv16_fs56_xor0;
  assign f_arrdiv16_fs56_and1 = f_arrdiv16_fs56_not1 & f_arrdiv16_fs55_or0;
  assign f_arrdiv16_fs56_or0 = f_arrdiv16_fs56_and1 | f_arrdiv16_fs56_and0;
  assign f_arrdiv16_fs57_xor0 = f_arrdiv16_mux2to138_xor0 ^ b[9];
  assign f_arrdiv16_fs57_not0 = ~f_arrdiv16_mux2to138_xor0;
  assign f_arrdiv16_fs57_and0 = f_arrdiv16_fs57_not0 & b[9];
  assign f_arrdiv16_fs57_xor1 = f_arrdiv16_fs56_or0 ^ f_arrdiv16_fs57_xor0;
  assign f_arrdiv16_fs57_not1 = ~f_arrdiv16_fs57_xor0;
  assign f_arrdiv16_fs57_and1 = f_arrdiv16_fs57_not1 & f_arrdiv16_fs56_or0;
  assign f_arrdiv16_fs57_or0 = f_arrdiv16_fs57_and1 | f_arrdiv16_fs57_and0;
  assign f_arrdiv16_fs58_xor0 = f_arrdiv16_mux2to139_xor0 ^ b[10];
  assign f_arrdiv16_fs58_not0 = ~f_arrdiv16_mux2to139_xor0;
  assign f_arrdiv16_fs58_and0 = f_arrdiv16_fs58_not0 & b[10];
  assign f_arrdiv16_fs58_xor1 = f_arrdiv16_fs57_or0 ^ f_arrdiv16_fs58_xor0;
  assign f_arrdiv16_fs58_not1 = ~f_arrdiv16_fs58_xor0;
  assign f_arrdiv16_fs58_and1 = f_arrdiv16_fs58_not1 & f_arrdiv16_fs57_or0;
  assign f_arrdiv16_fs58_or0 = f_arrdiv16_fs58_and1 | f_arrdiv16_fs58_and0;
  assign f_arrdiv16_fs59_xor0 = f_arrdiv16_mux2to140_xor0 ^ b[11];
  assign f_arrdiv16_fs59_not0 = ~f_arrdiv16_mux2to140_xor0;
  assign f_arrdiv16_fs59_and0 = f_arrdiv16_fs59_not0 & b[11];
  assign f_arrdiv16_fs59_xor1 = f_arrdiv16_fs58_or0 ^ f_arrdiv16_fs59_xor0;
  assign f_arrdiv16_fs59_not1 = ~f_arrdiv16_fs59_xor0;
  assign f_arrdiv16_fs59_and1 = f_arrdiv16_fs59_not1 & f_arrdiv16_fs58_or0;
  assign f_arrdiv16_fs59_or0 = f_arrdiv16_fs59_and1 | f_arrdiv16_fs59_and0;
  assign f_arrdiv16_fs60_xor0 = f_arrdiv16_mux2to141_xor0 ^ b[12];
  assign f_arrdiv16_fs60_not0 = ~f_arrdiv16_mux2to141_xor0;
  assign f_arrdiv16_fs60_and0 = f_arrdiv16_fs60_not0 & b[12];
  assign f_arrdiv16_fs60_xor1 = f_arrdiv16_fs59_or0 ^ f_arrdiv16_fs60_xor0;
  assign f_arrdiv16_fs60_not1 = ~f_arrdiv16_fs60_xor0;
  assign f_arrdiv16_fs60_and1 = f_arrdiv16_fs60_not1 & f_arrdiv16_fs59_or0;
  assign f_arrdiv16_fs60_or0 = f_arrdiv16_fs60_and1 | f_arrdiv16_fs60_and0;
  assign f_arrdiv16_fs61_xor0 = f_arrdiv16_mux2to142_xor0 ^ b[13];
  assign f_arrdiv16_fs61_not0 = ~f_arrdiv16_mux2to142_xor0;
  assign f_arrdiv16_fs61_and0 = f_arrdiv16_fs61_not0 & b[13];
  assign f_arrdiv16_fs61_xor1 = f_arrdiv16_fs60_or0 ^ f_arrdiv16_fs61_xor0;
  assign f_arrdiv16_fs61_not1 = ~f_arrdiv16_fs61_xor0;
  assign f_arrdiv16_fs61_and1 = f_arrdiv16_fs61_not1 & f_arrdiv16_fs60_or0;
  assign f_arrdiv16_fs61_or0 = f_arrdiv16_fs61_and1 | f_arrdiv16_fs61_and0;
  assign f_arrdiv16_fs62_xor0 = f_arrdiv16_mux2to143_xor0 ^ b[14];
  assign f_arrdiv16_fs62_not0 = ~f_arrdiv16_mux2to143_xor0;
  assign f_arrdiv16_fs62_and0 = f_arrdiv16_fs62_not0 & b[14];
  assign f_arrdiv16_fs62_xor1 = f_arrdiv16_fs61_or0 ^ f_arrdiv16_fs62_xor0;
  assign f_arrdiv16_fs62_not1 = ~f_arrdiv16_fs62_xor0;
  assign f_arrdiv16_fs62_and1 = f_arrdiv16_fs62_not1 & f_arrdiv16_fs61_or0;
  assign f_arrdiv16_fs62_or0 = f_arrdiv16_fs62_and1 | f_arrdiv16_fs62_and0;
  assign f_arrdiv16_fs63_xor0 = f_arrdiv16_mux2to144_xor0 ^ b[15];
  assign f_arrdiv16_fs63_not0 = ~f_arrdiv16_mux2to144_xor0;
  assign f_arrdiv16_fs63_and0 = f_arrdiv16_fs63_not0 & b[15];
  assign f_arrdiv16_fs63_xor1 = f_arrdiv16_fs62_or0 ^ f_arrdiv16_fs63_xor0;
  assign f_arrdiv16_fs63_not1 = ~f_arrdiv16_fs63_xor0;
  assign f_arrdiv16_fs63_and1 = f_arrdiv16_fs63_not1 & f_arrdiv16_fs62_or0;
  assign f_arrdiv16_fs63_or0 = f_arrdiv16_fs63_and1 | f_arrdiv16_fs63_and0;
  assign f_arrdiv16_mux2to145_and0 = a[12] & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to145_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to145_and1 = f_arrdiv16_fs48_xor0 & f_arrdiv16_mux2to145_not0;
  assign f_arrdiv16_mux2to145_xor0 = f_arrdiv16_mux2to145_and0 ^ f_arrdiv16_mux2to145_and1;
  assign f_arrdiv16_mux2to146_and0 = f_arrdiv16_mux2to130_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to146_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to146_and1 = f_arrdiv16_fs49_xor1 & f_arrdiv16_mux2to146_not0;
  assign f_arrdiv16_mux2to146_xor0 = f_arrdiv16_mux2to146_and0 ^ f_arrdiv16_mux2to146_and1;
  assign f_arrdiv16_mux2to147_and0 = f_arrdiv16_mux2to131_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to147_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to147_and1 = f_arrdiv16_fs50_xor1 & f_arrdiv16_mux2to147_not0;
  assign f_arrdiv16_mux2to147_xor0 = f_arrdiv16_mux2to147_and0 ^ f_arrdiv16_mux2to147_and1;
  assign f_arrdiv16_mux2to148_and0 = f_arrdiv16_mux2to132_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to148_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to148_and1 = f_arrdiv16_fs51_xor1 & f_arrdiv16_mux2to148_not0;
  assign f_arrdiv16_mux2to148_xor0 = f_arrdiv16_mux2to148_and0 ^ f_arrdiv16_mux2to148_and1;
  assign f_arrdiv16_mux2to149_and0 = f_arrdiv16_mux2to133_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to149_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to149_and1 = f_arrdiv16_fs52_xor1 & f_arrdiv16_mux2to149_not0;
  assign f_arrdiv16_mux2to149_xor0 = f_arrdiv16_mux2to149_and0 ^ f_arrdiv16_mux2to149_and1;
  assign f_arrdiv16_mux2to150_and0 = f_arrdiv16_mux2to134_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to150_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to150_and1 = f_arrdiv16_fs53_xor1 & f_arrdiv16_mux2to150_not0;
  assign f_arrdiv16_mux2to150_xor0 = f_arrdiv16_mux2to150_and0 ^ f_arrdiv16_mux2to150_and1;
  assign f_arrdiv16_mux2to151_and0 = f_arrdiv16_mux2to135_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to151_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to151_and1 = f_arrdiv16_fs54_xor1 & f_arrdiv16_mux2to151_not0;
  assign f_arrdiv16_mux2to151_xor0 = f_arrdiv16_mux2to151_and0 ^ f_arrdiv16_mux2to151_and1;
  assign f_arrdiv16_mux2to152_and0 = f_arrdiv16_mux2to136_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to152_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to152_and1 = f_arrdiv16_fs55_xor1 & f_arrdiv16_mux2to152_not0;
  assign f_arrdiv16_mux2to152_xor0 = f_arrdiv16_mux2to152_and0 ^ f_arrdiv16_mux2to152_and1;
  assign f_arrdiv16_mux2to153_and0 = f_arrdiv16_mux2to137_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to153_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to153_and1 = f_arrdiv16_fs56_xor1 & f_arrdiv16_mux2to153_not0;
  assign f_arrdiv16_mux2to153_xor0 = f_arrdiv16_mux2to153_and0 ^ f_arrdiv16_mux2to153_and1;
  assign f_arrdiv16_mux2to154_and0 = f_arrdiv16_mux2to138_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to154_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to154_and1 = f_arrdiv16_fs57_xor1 & f_arrdiv16_mux2to154_not0;
  assign f_arrdiv16_mux2to154_xor0 = f_arrdiv16_mux2to154_and0 ^ f_arrdiv16_mux2to154_and1;
  assign f_arrdiv16_mux2to155_and0 = f_arrdiv16_mux2to139_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to155_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to155_and1 = f_arrdiv16_fs58_xor1 & f_arrdiv16_mux2to155_not0;
  assign f_arrdiv16_mux2to155_xor0 = f_arrdiv16_mux2to155_and0 ^ f_arrdiv16_mux2to155_and1;
  assign f_arrdiv16_mux2to156_and0 = f_arrdiv16_mux2to140_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to156_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to156_and1 = f_arrdiv16_fs59_xor1 & f_arrdiv16_mux2to156_not0;
  assign f_arrdiv16_mux2to156_xor0 = f_arrdiv16_mux2to156_and0 ^ f_arrdiv16_mux2to156_and1;
  assign f_arrdiv16_mux2to157_and0 = f_arrdiv16_mux2to141_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to157_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to157_and1 = f_arrdiv16_fs60_xor1 & f_arrdiv16_mux2to157_not0;
  assign f_arrdiv16_mux2to157_xor0 = f_arrdiv16_mux2to157_and0 ^ f_arrdiv16_mux2to157_and1;
  assign f_arrdiv16_mux2to158_and0 = f_arrdiv16_mux2to142_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to158_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to158_and1 = f_arrdiv16_fs61_xor1 & f_arrdiv16_mux2to158_not0;
  assign f_arrdiv16_mux2to158_xor0 = f_arrdiv16_mux2to158_and0 ^ f_arrdiv16_mux2to158_and1;
  assign f_arrdiv16_mux2to159_and0 = f_arrdiv16_mux2to143_xor0 & f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to159_not0 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_mux2to159_and1 = f_arrdiv16_fs62_xor1 & f_arrdiv16_mux2to159_not0;
  assign f_arrdiv16_mux2to159_xor0 = f_arrdiv16_mux2to159_and0 ^ f_arrdiv16_mux2to159_and1;
  assign f_arrdiv16_not3 = ~f_arrdiv16_fs63_or0;
  assign f_arrdiv16_fs64_xor0 = a[11] ^ b[0];
  assign f_arrdiv16_fs64_not0 = ~a[11];
  assign f_arrdiv16_fs64_and0 = f_arrdiv16_fs64_not0 & b[0];
  assign f_arrdiv16_fs64_not1 = ~f_arrdiv16_fs64_xor0;
  assign f_arrdiv16_fs65_xor0 = f_arrdiv16_mux2to145_xor0 ^ b[1];
  assign f_arrdiv16_fs65_not0 = ~f_arrdiv16_mux2to145_xor0;
  assign f_arrdiv16_fs65_and0 = f_arrdiv16_fs65_not0 & b[1];
  assign f_arrdiv16_fs65_xor1 = f_arrdiv16_fs64_and0 ^ f_arrdiv16_fs65_xor0;
  assign f_arrdiv16_fs65_not1 = ~f_arrdiv16_fs65_xor0;
  assign f_arrdiv16_fs65_and1 = f_arrdiv16_fs65_not1 & f_arrdiv16_fs64_and0;
  assign f_arrdiv16_fs65_or0 = f_arrdiv16_fs65_and1 | f_arrdiv16_fs65_and0;
  assign f_arrdiv16_fs66_xor0 = f_arrdiv16_mux2to146_xor0 ^ b[2];
  assign f_arrdiv16_fs66_not0 = ~f_arrdiv16_mux2to146_xor0;
  assign f_arrdiv16_fs66_and0 = f_arrdiv16_fs66_not0 & b[2];
  assign f_arrdiv16_fs66_xor1 = f_arrdiv16_fs65_or0 ^ f_arrdiv16_fs66_xor0;
  assign f_arrdiv16_fs66_not1 = ~f_arrdiv16_fs66_xor0;
  assign f_arrdiv16_fs66_and1 = f_arrdiv16_fs66_not1 & f_arrdiv16_fs65_or0;
  assign f_arrdiv16_fs66_or0 = f_arrdiv16_fs66_and1 | f_arrdiv16_fs66_and0;
  assign f_arrdiv16_fs67_xor0 = f_arrdiv16_mux2to147_xor0 ^ b[3];
  assign f_arrdiv16_fs67_not0 = ~f_arrdiv16_mux2to147_xor0;
  assign f_arrdiv16_fs67_and0 = f_arrdiv16_fs67_not0 & b[3];
  assign f_arrdiv16_fs67_xor1 = f_arrdiv16_fs66_or0 ^ f_arrdiv16_fs67_xor0;
  assign f_arrdiv16_fs67_not1 = ~f_arrdiv16_fs67_xor0;
  assign f_arrdiv16_fs67_and1 = f_arrdiv16_fs67_not1 & f_arrdiv16_fs66_or0;
  assign f_arrdiv16_fs67_or0 = f_arrdiv16_fs67_and1 | f_arrdiv16_fs67_and0;
  assign f_arrdiv16_fs68_xor0 = f_arrdiv16_mux2to148_xor0 ^ b[4];
  assign f_arrdiv16_fs68_not0 = ~f_arrdiv16_mux2to148_xor0;
  assign f_arrdiv16_fs68_and0 = f_arrdiv16_fs68_not0 & b[4];
  assign f_arrdiv16_fs68_xor1 = f_arrdiv16_fs67_or0 ^ f_arrdiv16_fs68_xor0;
  assign f_arrdiv16_fs68_not1 = ~f_arrdiv16_fs68_xor0;
  assign f_arrdiv16_fs68_and1 = f_arrdiv16_fs68_not1 & f_arrdiv16_fs67_or0;
  assign f_arrdiv16_fs68_or0 = f_arrdiv16_fs68_and1 | f_arrdiv16_fs68_and0;
  assign f_arrdiv16_fs69_xor0 = f_arrdiv16_mux2to149_xor0 ^ b[5];
  assign f_arrdiv16_fs69_not0 = ~f_arrdiv16_mux2to149_xor0;
  assign f_arrdiv16_fs69_and0 = f_arrdiv16_fs69_not0 & b[5];
  assign f_arrdiv16_fs69_xor1 = f_arrdiv16_fs68_or0 ^ f_arrdiv16_fs69_xor0;
  assign f_arrdiv16_fs69_not1 = ~f_arrdiv16_fs69_xor0;
  assign f_arrdiv16_fs69_and1 = f_arrdiv16_fs69_not1 & f_arrdiv16_fs68_or0;
  assign f_arrdiv16_fs69_or0 = f_arrdiv16_fs69_and1 | f_arrdiv16_fs69_and0;
  assign f_arrdiv16_fs70_xor0 = f_arrdiv16_mux2to150_xor0 ^ b[6];
  assign f_arrdiv16_fs70_not0 = ~f_arrdiv16_mux2to150_xor0;
  assign f_arrdiv16_fs70_and0 = f_arrdiv16_fs70_not0 & b[6];
  assign f_arrdiv16_fs70_xor1 = f_arrdiv16_fs69_or0 ^ f_arrdiv16_fs70_xor0;
  assign f_arrdiv16_fs70_not1 = ~f_arrdiv16_fs70_xor0;
  assign f_arrdiv16_fs70_and1 = f_arrdiv16_fs70_not1 & f_arrdiv16_fs69_or0;
  assign f_arrdiv16_fs70_or0 = f_arrdiv16_fs70_and1 | f_arrdiv16_fs70_and0;
  assign f_arrdiv16_fs71_xor0 = f_arrdiv16_mux2to151_xor0 ^ b[7];
  assign f_arrdiv16_fs71_not0 = ~f_arrdiv16_mux2to151_xor0;
  assign f_arrdiv16_fs71_and0 = f_arrdiv16_fs71_not0 & b[7];
  assign f_arrdiv16_fs71_xor1 = f_arrdiv16_fs70_or0 ^ f_arrdiv16_fs71_xor0;
  assign f_arrdiv16_fs71_not1 = ~f_arrdiv16_fs71_xor0;
  assign f_arrdiv16_fs71_and1 = f_arrdiv16_fs71_not1 & f_arrdiv16_fs70_or0;
  assign f_arrdiv16_fs71_or0 = f_arrdiv16_fs71_and1 | f_arrdiv16_fs71_and0;
  assign f_arrdiv16_fs72_xor0 = f_arrdiv16_mux2to152_xor0 ^ b[8];
  assign f_arrdiv16_fs72_not0 = ~f_arrdiv16_mux2to152_xor0;
  assign f_arrdiv16_fs72_and0 = f_arrdiv16_fs72_not0 & b[8];
  assign f_arrdiv16_fs72_xor1 = f_arrdiv16_fs71_or0 ^ f_arrdiv16_fs72_xor0;
  assign f_arrdiv16_fs72_not1 = ~f_arrdiv16_fs72_xor0;
  assign f_arrdiv16_fs72_and1 = f_arrdiv16_fs72_not1 & f_arrdiv16_fs71_or0;
  assign f_arrdiv16_fs72_or0 = f_arrdiv16_fs72_and1 | f_arrdiv16_fs72_and0;
  assign f_arrdiv16_fs73_xor0 = f_arrdiv16_mux2to153_xor0 ^ b[9];
  assign f_arrdiv16_fs73_not0 = ~f_arrdiv16_mux2to153_xor0;
  assign f_arrdiv16_fs73_and0 = f_arrdiv16_fs73_not0 & b[9];
  assign f_arrdiv16_fs73_xor1 = f_arrdiv16_fs72_or0 ^ f_arrdiv16_fs73_xor0;
  assign f_arrdiv16_fs73_not1 = ~f_arrdiv16_fs73_xor0;
  assign f_arrdiv16_fs73_and1 = f_arrdiv16_fs73_not1 & f_arrdiv16_fs72_or0;
  assign f_arrdiv16_fs73_or0 = f_arrdiv16_fs73_and1 | f_arrdiv16_fs73_and0;
  assign f_arrdiv16_fs74_xor0 = f_arrdiv16_mux2to154_xor0 ^ b[10];
  assign f_arrdiv16_fs74_not0 = ~f_arrdiv16_mux2to154_xor0;
  assign f_arrdiv16_fs74_and0 = f_arrdiv16_fs74_not0 & b[10];
  assign f_arrdiv16_fs74_xor1 = f_arrdiv16_fs73_or0 ^ f_arrdiv16_fs74_xor0;
  assign f_arrdiv16_fs74_not1 = ~f_arrdiv16_fs74_xor0;
  assign f_arrdiv16_fs74_and1 = f_arrdiv16_fs74_not1 & f_arrdiv16_fs73_or0;
  assign f_arrdiv16_fs74_or0 = f_arrdiv16_fs74_and1 | f_arrdiv16_fs74_and0;
  assign f_arrdiv16_fs75_xor0 = f_arrdiv16_mux2to155_xor0 ^ b[11];
  assign f_arrdiv16_fs75_not0 = ~f_arrdiv16_mux2to155_xor0;
  assign f_arrdiv16_fs75_and0 = f_arrdiv16_fs75_not0 & b[11];
  assign f_arrdiv16_fs75_xor1 = f_arrdiv16_fs74_or0 ^ f_arrdiv16_fs75_xor0;
  assign f_arrdiv16_fs75_not1 = ~f_arrdiv16_fs75_xor0;
  assign f_arrdiv16_fs75_and1 = f_arrdiv16_fs75_not1 & f_arrdiv16_fs74_or0;
  assign f_arrdiv16_fs75_or0 = f_arrdiv16_fs75_and1 | f_arrdiv16_fs75_and0;
  assign f_arrdiv16_fs76_xor0 = f_arrdiv16_mux2to156_xor0 ^ b[12];
  assign f_arrdiv16_fs76_not0 = ~f_arrdiv16_mux2to156_xor0;
  assign f_arrdiv16_fs76_and0 = f_arrdiv16_fs76_not0 & b[12];
  assign f_arrdiv16_fs76_xor1 = f_arrdiv16_fs75_or0 ^ f_arrdiv16_fs76_xor0;
  assign f_arrdiv16_fs76_not1 = ~f_arrdiv16_fs76_xor0;
  assign f_arrdiv16_fs76_and1 = f_arrdiv16_fs76_not1 & f_arrdiv16_fs75_or0;
  assign f_arrdiv16_fs76_or0 = f_arrdiv16_fs76_and1 | f_arrdiv16_fs76_and0;
  assign f_arrdiv16_fs77_xor0 = f_arrdiv16_mux2to157_xor0 ^ b[13];
  assign f_arrdiv16_fs77_not0 = ~f_arrdiv16_mux2to157_xor0;
  assign f_arrdiv16_fs77_and0 = f_arrdiv16_fs77_not0 & b[13];
  assign f_arrdiv16_fs77_xor1 = f_arrdiv16_fs76_or0 ^ f_arrdiv16_fs77_xor0;
  assign f_arrdiv16_fs77_not1 = ~f_arrdiv16_fs77_xor0;
  assign f_arrdiv16_fs77_and1 = f_arrdiv16_fs77_not1 & f_arrdiv16_fs76_or0;
  assign f_arrdiv16_fs77_or0 = f_arrdiv16_fs77_and1 | f_arrdiv16_fs77_and0;
  assign f_arrdiv16_fs78_xor0 = f_arrdiv16_mux2to158_xor0 ^ b[14];
  assign f_arrdiv16_fs78_not0 = ~f_arrdiv16_mux2to158_xor0;
  assign f_arrdiv16_fs78_and0 = f_arrdiv16_fs78_not0 & b[14];
  assign f_arrdiv16_fs78_xor1 = f_arrdiv16_fs77_or0 ^ f_arrdiv16_fs78_xor0;
  assign f_arrdiv16_fs78_not1 = ~f_arrdiv16_fs78_xor0;
  assign f_arrdiv16_fs78_and1 = f_arrdiv16_fs78_not1 & f_arrdiv16_fs77_or0;
  assign f_arrdiv16_fs78_or0 = f_arrdiv16_fs78_and1 | f_arrdiv16_fs78_and0;
  assign f_arrdiv16_fs79_xor0 = f_arrdiv16_mux2to159_xor0 ^ b[15];
  assign f_arrdiv16_fs79_not0 = ~f_arrdiv16_mux2to159_xor0;
  assign f_arrdiv16_fs79_and0 = f_arrdiv16_fs79_not0 & b[15];
  assign f_arrdiv16_fs79_xor1 = f_arrdiv16_fs78_or0 ^ f_arrdiv16_fs79_xor0;
  assign f_arrdiv16_fs79_not1 = ~f_arrdiv16_fs79_xor0;
  assign f_arrdiv16_fs79_and1 = f_arrdiv16_fs79_not1 & f_arrdiv16_fs78_or0;
  assign f_arrdiv16_fs79_or0 = f_arrdiv16_fs79_and1 | f_arrdiv16_fs79_and0;
  assign f_arrdiv16_mux2to160_and0 = a[11] & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to160_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to160_and1 = f_arrdiv16_fs64_xor0 & f_arrdiv16_mux2to160_not0;
  assign f_arrdiv16_mux2to160_xor0 = f_arrdiv16_mux2to160_and0 ^ f_arrdiv16_mux2to160_and1;
  assign f_arrdiv16_mux2to161_and0 = f_arrdiv16_mux2to145_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to161_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to161_and1 = f_arrdiv16_fs65_xor1 & f_arrdiv16_mux2to161_not0;
  assign f_arrdiv16_mux2to161_xor0 = f_arrdiv16_mux2to161_and0 ^ f_arrdiv16_mux2to161_and1;
  assign f_arrdiv16_mux2to162_and0 = f_arrdiv16_mux2to146_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to162_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to162_and1 = f_arrdiv16_fs66_xor1 & f_arrdiv16_mux2to162_not0;
  assign f_arrdiv16_mux2to162_xor0 = f_arrdiv16_mux2to162_and0 ^ f_arrdiv16_mux2to162_and1;
  assign f_arrdiv16_mux2to163_and0 = f_arrdiv16_mux2to147_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to163_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to163_and1 = f_arrdiv16_fs67_xor1 & f_arrdiv16_mux2to163_not0;
  assign f_arrdiv16_mux2to163_xor0 = f_arrdiv16_mux2to163_and0 ^ f_arrdiv16_mux2to163_and1;
  assign f_arrdiv16_mux2to164_and0 = f_arrdiv16_mux2to148_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to164_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to164_and1 = f_arrdiv16_fs68_xor1 & f_arrdiv16_mux2to164_not0;
  assign f_arrdiv16_mux2to164_xor0 = f_arrdiv16_mux2to164_and0 ^ f_arrdiv16_mux2to164_and1;
  assign f_arrdiv16_mux2to165_and0 = f_arrdiv16_mux2to149_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to165_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to165_and1 = f_arrdiv16_fs69_xor1 & f_arrdiv16_mux2to165_not0;
  assign f_arrdiv16_mux2to165_xor0 = f_arrdiv16_mux2to165_and0 ^ f_arrdiv16_mux2to165_and1;
  assign f_arrdiv16_mux2to166_and0 = f_arrdiv16_mux2to150_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to166_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to166_and1 = f_arrdiv16_fs70_xor1 & f_arrdiv16_mux2to166_not0;
  assign f_arrdiv16_mux2to166_xor0 = f_arrdiv16_mux2to166_and0 ^ f_arrdiv16_mux2to166_and1;
  assign f_arrdiv16_mux2to167_and0 = f_arrdiv16_mux2to151_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to167_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to167_and1 = f_arrdiv16_fs71_xor1 & f_arrdiv16_mux2to167_not0;
  assign f_arrdiv16_mux2to167_xor0 = f_arrdiv16_mux2to167_and0 ^ f_arrdiv16_mux2to167_and1;
  assign f_arrdiv16_mux2to168_and0 = f_arrdiv16_mux2to152_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to168_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to168_and1 = f_arrdiv16_fs72_xor1 & f_arrdiv16_mux2to168_not0;
  assign f_arrdiv16_mux2to168_xor0 = f_arrdiv16_mux2to168_and0 ^ f_arrdiv16_mux2to168_and1;
  assign f_arrdiv16_mux2to169_and0 = f_arrdiv16_mux2to153_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to169_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to169_and1 = f_arrdiv16_fs73_xor1 & f_arrdiv16_mux2to169_not0;
  assign f_arrdiv16_mux2to169_xor0 = f_arrdiv16_mux2to169_and0 ^ f_arrdiv16_mux2to169_and1;
  assign f_arrdiv16_mux2to170_and0 = f_arrdiv16_mux2to154_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to170_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to170_and1 = f_arrdiv16_fs74_xor1 & f_arrdiv16_mux2to170_not0;
  assign f_arrdiv16_mux2to170_xor0 = f_arrdiv16_mux2to170_and0 ^ f_arrdiv16_mux2to170_and1;
  assign f_arrdiv16_mux2to171_and0 = f_arrdiv16_mux2to155_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to171_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to171_and1 = f_arrdiv16_fs75_xor1 & f_arrdiv16_mux2to171_not0;
  assign f_arrdiv16_mux2to171_xor0 = f_arrdiv16_mux2to171_and0 ^ f_arrdiv16_mux2to171_and1;
  assign f_arrdiv16_mux2to172_and0 = f_arrdiv16_mux2to156_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to172_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to172_and1 = f_arrdiv16_fs76_xor1 & f_arrdiv16_mux2to172_not0;
  assign f_arrdiv16_mux2to172_xor0 = f_arrdiv16_mux2to172_and0 ^ f_arrdiv16_mux2to172_and1;
  assign f_arrdiv16_mux2to173_and0 = f_arrdiv16_mux2to157_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to173_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to173_and1 = f_arrdiv16_fs77_xor1 & f_arrdiv16_mux2to173_not0;
  assign f_arrdiv16_mux2to173_xor0 = f_arrdiv16_mux2to173_and0 ^ f_arrdiv16_mux2to173_and1;
  assign f_arrdiv16_mux2to174_and0 = f_arrdiv16_mux2to158_xor0 & f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to174_not0 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_mux2to174_and1 = f_arrdiv16_fs78_xor1 & f_arrdiv16_mux2to174_not0;
  assign f_arrdiv16_mux2to174_xor0 = f_arrdiv16_mux2to174_and0 ^ f_arrdiv16_mux2to174_and1;
  assign f_arrdiv16_not4 = ~f_arrdiv16_fs79_or0;
  assign f_arrdiv16_fs80_xor0 = a[10] ^ b[0];
  assign f_arrdiv16_fs80_not0 = ~a[10];
  assign f_arrdiv16_fs80_and0 = f_arrdiv16_fs80_not0 & b[0];
  assign f_arrdiv16_fs80_not1 = ~f_arrdiv16_fs80_xor0;
  assign f_arrdiv16_fs81_xor0 = f_arrdiv16_mux2to160_xor0 ^ b[1];
  assign f_arrdiv16_fs81_not0 = ~f_arrdiv16_mux2to160_xor0;
  assign f_arrdiv16_fs81_and0 = f_arrdiv16_fs81_not0 & b[1];
  assign f_arrdiv16_fs81_xor1 = f_arrdiv16_fs80_and0 ^ f_arrdiv16_fs81_xor0;
  assign f_arrdiv16_fs81_not1 = ~f_arrdiv16_fs81_xor0;
  assign f_arrdiv16_fs81_and1 = f_arrdiv16_fs81_not1 & f_arrdiv16_fs80_and0;
  assign f_arrdiv16_fs81_or0 = f_arrdiv16_fs81_and1 | f_arrdiv16_fs81_and0;
  assign f_arrdiv16_fs82_xor0 = f_arrdiv16_mux2to161_xor0 ^ b[2];
  assign f_arrdiv16_fs82_not0 = ~f_arrdiv16_mux2to161_xor0;
  assign f_arrdiv16_fs82_and0 = f_arrdiv16_fs82_not0 & b[2];
  assign f_arrdiv16_fs82_xor1 = f_arrdiv16_fs81_or0 ^ f_arrdiv16_fs82_xor0;
  assign f_arrdiv16_fs82_not1 = ~f_arrdiv16_fs82_xor0;
  assign f_arrdiv16_fs82_and1 = f_arrdiv16_fs82_not1 & f_arrdiv16_fs81_or0;
  assign f_arrdiv16_fs82_or0 = f_arrdiv16_fs82_and1 | f_arrdiv16_fs82_and0;
  assign f_arrdiv16_fs83_xor0 = f_arrdiv16_mux2to162_xor0 ^ b[3];
  assign f_arrdiv16_fs83_not0 = ~f_arrdiv16_mux2to162_xor0;
  assign f_arrdiv16_fs83_and0 = f_arrdiv16_fs83_not0 & b[3];
  assign f_arrdiv16_fs83_xor1 = f_arrdiv16_fs82_or0 ^ f_arrdiv16_fs83_xor0;
  assign f_arrdiv16_fs83_not1 = ~f_arrdiv16_fs83_xor0;
  assign f_arrdiv16_fs83_and1 = f_arrdiv16_fs83_not1 & f_arrdiv16_fs82_or0;
  assign f_arrdiv16_fs83_or0 = f_arrdiv16_fs83_and1 | f_arrdiv16_fs83_and0;
  assign f_arrdiv16_fs84_xor0 = f_arrdiv16_mux2to163_xor0 ^ b[4];
  assign f_arrdiv16_fs84_not0 = ~f_arrdiv16_mux2to163_xor0;
  assign f_arrdiv16_fs84_and0 = f_arrdiv16_fs84_not0 & b[4];
  assign f_arrdiv16_fs84_xor1 = f_arrdiv16_fs83_or0 ^ f_arrdiv16_fs84_xor0;
  assign f_arrdiv16_fs84_not1 = ~f_arrdiv16_fs84_xor0;
  assign f_arrdiv16_fs84_and1 = f_arrdiv16_fs84_not1 & f_arrdiv16_fs83_or0;
  assign f_arrdiv16_fs84_or0 = f_arrdiv16_fs84_and1 | f_arrdiv16_fs84_and0;
  assign f_arrdiv16_fs85_xor0 = f_arrdiv16_mux2to164_xor0 ^ b[5];
  assign f_arrdiv16_fs85_not0 = ~f_arrdiv16_mux2to164_xor0;
  assign f_arrdiv16_fs85_and0 = f_arrdiv16_fs85_not0 & b[5];
  assign f_arrdiv16_fs85_xor1 = f_arrdiv16_fs84_or0 ^ f_arrdiv16_fs85_xor0;
  assign f_arrdiv16_fs85_not1 = ~f_arrdiv16_fs85_xor0;
  assign f_arrdiv16_fs85_and1 = f_arrdiv16_fs85_not1 & f_arrdiv16_fs84_or0;
  assign f_arrdiv16_fs85_or0 = f_arrdiv16_fs85_and1 | f_arrdiv16_fs85_and0;
  assign f_arrdiv16_fs86_xor0 = f_arrdiv16_mux2to165_xor0 ^ b[6];
  assign f_arrdiv16_fs86_not0 = ~f_arrdiv16_mux2to165_xor0;
  assign f_arrdiv16_fs86_and0 = f_arrdiv16_fs86_not0 & b[6];
  assign f_arrdiv16_fs86_xor1 = f_arrdiv16_fs85_or0 ^ f_arrdiv16_fs86_xor0;
  assign f_arrdiv16_fs86_not1 = ~f_arrdiv16_fs86_xor0;
  assign f_arrdiv16_fs86_and1 = f_arrdiv16_fs86_not1 & f_arrdiv16_fs85_or0;
  assign f_arrdiv16_fs86_or0 = f_arrdiv16_fs86_and1 | f_arrdiv16_fs86_and0;
  assign f_arrdiv16_fs87_xor0 = f_arrdiv16_mux2to166_xor0 ^ b[7];
  assign f_arrdiv16_fs87_not0 = ~f_arrdiv16_mux2to166_xor0;
  assign f_arrdiv16_fs87_and0 = f_arrdiv16_fs87_not0 & b[7];
  assign f_arrdiv16_fs87_xor1 = f_arrdiv16_fs86_or0 ^ f_arrdiv16_fs87_xor0;
  assign f_arrdiv16_fs87_not1 = ~f_arrdiv16_fs87_xor0;
  assign f_arrdiv16_fs87_and1 = f_arrdiv16_fs87_not1 & f_arrdiv16_fs86_or0;
  assign f_arrdiv16_fs87_or0 = f_arrdiv16_fs87_and1 | f_arrdiv16_fs87_and0;
  assign f_arrdiv16_fs88_xor0 = f_arrdiv16_mux2to167_xor0 ^ b[8];
  assign f_arrdiv16_fs88_not0 = ~f_arrdiv16_mux2to167_xor0;
  assign f_arrdiv16_fs88_and0 = f_arrdiv16_fs88_not0 & b[8];
  assign f_arrdiv16_fs88_xor1 = f_arrdiv16_fs87_or0 ^ f_arrdiv16_fs88_xor0;
  assign f_arrdiv16_fs88_not1 = ~f_arrdiv16_fs88_xor0;
  assign f_arrdiv16_fs88_and1 = f_arrdiv16_fs88_not1 & f_arrdiv16_fs87_or0;
  assign f_arrdiv16_fs88_or0 = f_arrdiv16_fs88_and1 | f_arrdiv16_fs88_and0;
  assign f_arrdiv16_fs89_xor0 = f_arrdiv16_mux2to168_xor0 ^ b[9];
  assign f_arrdiv16_fs89_not0 = ~f_arrdiv16_mux2to168_xor0;
  assign f_arrdiv16_fs89_and0 = f_arrdiv16_fs89_not0 & b[9];
  assign f_arrdiv16_fs89_xor1 = f_arrdiv16_fs88_or0 ^ f_arrdiv16_fs89_xor0;
  assign f_arrdiv16_fs89_not1 = ~f_arrdiv16_fs89_xor0;
  assign f_arrdiv16_fs89_and1 = f_arrdiv16_fs89_not1 & f_arrdiv16_fs88_or0;
  assign f_arrdiv16_fs89_or0 = f_arrdiv16_fs89_and1 | f_arrdiv16_fs89_and0;
  assign f_arrdiv16_fs90_xor0 = f_arrdiv16_mux2to169_xor0 ^ b[10];
  assign f_arrdiv16_fs90_not0 = ~f_arrdiv16_mux2to169_xor0;
  assign f_arrdiv16_fs90_and0 = f_arrdiv16_fs90_not0 & b[10];
  assign f_arrdiv16_fs90_xor1 = f_arrdiv16_fs89_or0 ^ f_arrdiv16_fs90_xor0;
  assign f_arrdiv16_fs90_not1 = ~f_arrdiv16_fs90_xor0;
  assign f_arrdiv16_fs90_and1 = f_arrdiv16_fs90_not1 & f_arrdiv16_fs89_or0;
  assign f_arrdiv16_fs90_or0 = f_arrdiv16_fs90_and1 | f_arrdiv16_fs90_and0;
  assign f_arrdiv16_fs91_xor0 = f_arrdiv16_mux2to170_xor0 ^ b[11];
  assign f_arrdiv16_fs91_not0 = ~f_arrdiv16_mux2to170_xor0;
  assign f_arrdiv16_fs91_and0 = f_arrdiv16_fs91_not0 & b[11];
  assign f_arrdiv16_fs91_xor1 = f_arrdiv16_fs90_or0 ^ f_arrdiv16_fs91_xor0;
  assign f_arrdiv16_fs91_not1 = ~f_arrdiv16_fs91_xor0;
  assign f_arrdiv16_fs91_and1 = f_arrdiv16_fs91_not1 & f_arrdiv16_fs90_or0;
  assign f_arrdiv16_fs91_or0 = f_arrdiv16_fs91_and1 | f_arrdiv16_fs91_and0;
  assign f_arrdiv16_fs92_xor0 = f_arrdiv16_mux2to171_xor0 ^ b[12];
  assign f_arrdiv16_fs92_not0 = ~f_arrdiv16_mux2to171_xor0;
  assign f_arrdiv16_fs92_and0 = f_arrdiv16_fs92_not0 & b[12];
  assign f_arrdiv16_fs92_xor1 = f_arrdiv16_fs91_or0 ^ f_arrdiv16_fs92_xor0;
  assign f_arrdiv16_fs92_not1 = ~f_arrdiv16_fs92_xor0;
  assign f_arrdiv16_fs92_and1 = f_arrdiv16_fs92_not1 & f_arrdiv16_fs91_or0;
  assign f_arrdiv16_fs92_or0 = f_arrdiv16_fs92_and1 | f_arrdiv16_fs92_and0;
  assign f_arrdiv16_fs93_xor0 = f_arrdiv16_mux2to172_xor0 ^ b[13];
  assign f_arrdiv16_fs93_not0 = ~f_arrdiv16_mux2to172_xor0;
  assign f_arrdiv16_fs93_and0 = f_arrdiv16_fs93_not0 & b[13];
  assign f_arrdiv16_fs93_xor1 = f_arrdiv16_fs92_or0 ^ f_arrdiv16_fs93_xor0;
  assign f_arrdiv16_fs93_not1 = ~f_arrdiv16_fs93_xor0;
  assign f_arrdiv16_fs93_and1 = f_arrdiv16_fs93_not1 & f_arrdiv16_fs92_or0;
  assign f_arrdiv16_fs93_or0 = f_arrdiv16_fs93_and1 | f_arrdiv16_fs93_and0;
  assign f_arrdiv16_fs94_xor0 = f_arrdiv16_mux2to173_xor0 ^ b[14];
  assign f_arrdiv16_fs94_not0 = ~f_arrdiv16_mux2to173_xor0;
  assign f_arrdiv16_fs94_and0 = f_arrdiv16_fs94_not0 & b[14];
  assign f_arrdiv16_fs94_xor1 = f_arrdiv16_fs93_or0 ^ f_arrdiv16_fs94_xor0;
  assign f_arrdiv16_fs94_not1 = ~f_arrdiv16_fs94_xor0;
  assign f_arrdiv16_fs94_and1 = f_arrdiv16_fs94_not1 & f_arrdiv16_fs93_or0;
  assign f_arrdiv16_fs94_or0 = f_arrdiv16_fs94_and1 | f_arrdiv16_fs94_and0;
  assign f_arrdiv16_fs95_xor0 = f_arrdiv16_mux2to174_xor0 ^ b[15];
  assign f_arrdiv16_fs95_not0 = ~f_arrdiv16_mux2to174_xor0;
  assign f_arrdiv16_fs95_and0 = f_arrdiv16_fs95_not0 & b[15];
  assign f_arrdiv16_fs95_xor1 = f_arrdiv16_fs94_or0 ^ f_arrdiv16_fs95_xor0;
  assign f_arrdiv16_fs95_not1 = ~f_arrdiv16_fs95_xor0;
  assign f_arrdiv16_fs95_and1 = f_arrdiv16_fs95_not1 & f_arrdiv16_fs94_or0;
  assign f_arrdiv16_fs95_or0 = f_arrdiv16_fs95_and1 | f_arrdiv16_fs95_and0;
  assign f_arrdiv16_mux2to175_and0 = a[10] & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to175_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to175_and1 = f_arrdiv16_fs80_xor0 & f_arrdiv16_mux2to175_not0;
  assign f_arrdiv16_mux2to175_xor0 = f_arrdiv16_mux2to175_and0 ^ f_arrdiv16_mux2to175_and1;
  assign f_arrdiv16_mux2to176_and0 = f_arrdiv16_mux2to160_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to176_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to176_and1 = f_arrdiv16_fs81_xor1 & f_arrdiv16_mux2to176_not0;
  assign f_arrdiv16_mux2to176_xor0 = f_arrdiv16_mux2to176_and0 ^ f_arrdiv16_mux2to176_and1;
  assign f_arrdiv16_mux2to177_and0 = f_arrdiv16_mux2to161_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to177_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to177_and1 = f_arrdiv16_fs82_xor1 & f_arrdiv16_mux2to177_not0;
  assign f_arrdiv16_mux2to177_xor0 = f_arrdiv16_mux2to177_and0 ^ f_arrdiv16_mux2to177_and1;
  assign f_arrdiv16_mux2to178_and0 = f_arrdiv16_mux2to162_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to178_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to178_and1 = f_arrdiv16_fs83_xor1 & f_arrdiv16_mux2to178_not0;
  assign f_arrdiv16_mux2to178_xor0 = f_arrdiv16_mux2to178_and0 ^ f_arrdiv16_mux2to178_and1;
  assign f_arrdiv16_mux2to179_and0 = f_arrdiv16_mux2to163_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to179_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to179_and1 = f_arrdiv16_fs84_xor1 & f_arrdiv16_mux2to179_not0;
  assign f_arrdiv16_mux2to179_xor0 = f_arrdiv16_mux2to179_and0 ^ f_arrdiv16_mux2to179_and1;
  assign f_arrdiv16_mux2to180_and0 = f_arrdiv16_mux2to164_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to180_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to180_and1 = f_arrdiv16_fs85_xor1 & f_arrdiv16_mux2to180_not0;
  assign f_arrdiv16_mux2to180_xor0 = f_arrdiv16_mux2to180_and0 ^ f_arrdiv16_mux2to180_and1;
  assign f_arrdiv16_mux2to181_and0 = f_arrdiv16_mux2to165_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to181_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to181_and1 = f_arrdiv16_fs86_xor1 & f_arrdiv16_mux2to181_not0;
  assign f_arrdiv16_mux2to181_xor0 = f_arrdiv16_mux2to181_and0 ^ f_arrdiv16_mux2to181_and1;
  assign f_arrdiv16_mux2to182_and0 = f_arrdiv16_mux2to166_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to182_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to182_and1 = f_arrdiv16_fs87_xor1 & f_arrdiv16_mux2to182_not0;
  assign f_arrdiv16_mux2to182_xor0 = f_arrdiv16_mux2to182_and0 ^ f_arrdiv16_mux2to182_and1;
  assign f_arrdiv16_mux2to183_and0 = f_arrdiv16_mux2to167_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to183_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to183_and1 = f_arrdiv16_fs88_xor1 & f_arrdiv16_mux2to183_not0;
  assign f_arrdiv16_mux2to183_xor0 = f_arrdiv16_mux2to183_and0 ^ f_arrdiv16_mux2to183_and1;
  assign f_arrdiv16_mux2to184_and0 = f_arrdiv16_mux2to168_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to184_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to184_and1 = f_arrdiv16_fs89_xor1 & f_arrdiv16_mux2to184_not0;
  assign f_arrdiv16_mux2to184_xor0 = f_arrdiv16_mux2to184_and0 ^ f_arrdiv16_mux2to184_and1;
  assign f_arrdiv16_mux2to185_and0 = f_arrdiv16_mux2to169_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to185_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to185_and1 = f_arrdiv16_fs90_xor1 & f_arrdiv16_mux2to185_not0;
  assign f_arrdiv16_mux2to185_xor0 = f_arrdiv16_mux2to185_and0 ^ f_arrdiv16_mux2to185_and1;
  assign f_arrdiv16_mux2to186_and0 = f_arrdiv16_mux2to170_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to186_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to186_and1 = f_arrdiv16_fs91_xor1 & f_arrdiv16_mux2to186_not0;
  assign f_arrdiv16_mux2to186_xor0 = f_arrdiv16_mux2to186_and0 ^ f_arrdiv16_mux2to186_and1;
  assign f_arrdiv16_mux2to187_and0 = f_arrdiv16_mux2to171_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to187_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to187_and1 = f_arrdiv16_fs92_xor1 & f_arrdiv16_mux2to187_not0;
  assign f_arrdiv16_mux2to187_xor0 = f_arrdiv16_mux2to187_and0 ^ f_arrdiv16_mux2to187_and1;
  assign f_arrdiv16_mux2to188_and0 = f_arrdiv16_mux2to172_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to188_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to188_and1 = f_arrdiv16_fs93_xor1 & f_arrdiv16_mux2to188_not0;
  assign f_arrdiv16_mux2to188_xor0 = f_arrdiv16_mux2to188_and0 ^ f_arrdiv16_mux2to188_and1;
  assign f_arrdiv16_mux2to189_and0 = f_arrdiv16_mux2to173_xor0 & f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to189_not0 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_mux2to189_and1 = f_arrdiv16_fs94_xor1 & f_arrdiv16_mux2to189_not0;
  assign f_arrdiv16_mux2to189_xor0 = f_arrdiv16_mux2to189_and0 ^ f_arrdiv16_mux2to189_and1;
  assign f_arrdiv16_not5 = ~f_arrdiv16_fs95_or0;
  assign f_arrdiv16_fs96_xor0 = a[9] ^ b[0];
  assign f_arrdiv16_fs96_not0 = ~a[9];
  assign f_arrdiv16_fs96_and0 = f_arrdiv16_fs96_not0 & b[0];
  assign f_arrdiv16_fs96_not1 = ~f_arrdiv16_fs96_xor0;
  assign f_arrdiv16_fs97_xor0 = f_arrdiv16_mux2to175_xor0 ^ b[1];
  assign f_arrdiv16_fs97_not0 = ~f_arrdiv16_mux2to175_xor0;
  assign f_arrdiv16_fs97_and0 = f_arrdiv16_fs97_not0 & b[1];
  assign f_arrdiv16_fs97_xor1 = f_arrdiv16_fs96_and0 ^ f_arrdiv16_fs97_xor0;
  assign f_arrdiv16_fs97_not1 = ~f_arrdiv16_fs97_xor0;
  assign f_arrdiv16_fs97_and1 = f_arrdiv16_fs97_not1 & f_arrdiv16_fs96_and0;
  assign f_arrdiv16_fs97_or0 = f_arrdiv16_fs97_and1 | f_arrdiv16_fs97_and0;
  assign f_arrdiv16_fs98_xor0 = f_arrdiv16_mux2to176_xor0 ^ b[2];
  assign f_arrdiv16_fs98_not0 = ~f_arrdiv16_mux2to176_xor0;
  assign f_arrdiv16_fs98_and0 = f_arrdiv16_fs98_not0 & b[2];
  assign f_arrdiv16_fs98_xor1 = f_arrdiv16_fs97_or0 ^ f_arrdiv16_fs98_xor0;
  assign f_arrdiv16_fs98_not1 = ~f_arrdiv16_fs98_xor0;
  assign f_arrdiv16_fs98_and1 = f_arrdiv16_fs98_not1 & f_arrdiv16_fs97_or0;
  assign f_arrdiv16_fs98_or0 = f_arrdiv16_fs98_and1 | f_arrdiv16_fs98_and0;
  assign f_arrdiv16_fs99_xor0 = f_arrdiv16_mux2to177_xor0 ^ b[3];
  assign f_arrdiv16_fs99_not0 = ~f_arrdiv16_mux2to177_xor0;
  assign f_arrdiv16_fs99_and0 = f_arrdiv16_fs99_not0 & b[3];
  assign f_arrdiv16_fs99_xor1 = f_arrdiv16_fs98_or0 ^ f_arrdiv16_fs99_xor0;
  assign f_arrdiv16_fs99_not1 = ~f_arrdiv16_fs99_xor0;
  assign f_arrdiv16_fs99_and1 = f_arrdiv16_fs99_not1 & f_arrdiv16_fs98_or0;
  assign f_arrdiv16_fs99_or0 = f_arrdiv16_fs99_and1 | f_arrdiv16_fs99_and0;
  assign f_arrdiv16_fs100_xor0 = f_arrdiv16_mux2to178_xor0 ^ b[4];
  assign f_arrdiv16_fs100_not0 = ~f_arrdiv16_mux2to178_xor0;
  assign f_arrdiv16_fs100_and0 = f_arrdiv16_fs100_not0 & b[4];
  assign f_arrdiv16_fs100_xor1 = f_arrdiv16_fs99_or0 ^ f_arrdiv16_fs100_xor0;
  assign f_arrdiv16_fs100_not1 = ~f_arrdiv16_fs100_xor0;
  assign f_arrdiv16_fs100_and1 = f_arrdiv16_fs100_not1 & f_arrdiv16_fs99_or0;
  assign f_arrdiv16_fs100_or0 = f_arrdiv16_fs100_and1 | f_arrdiv16_fs100_and0;
  assign f_arrdiv16_fs101_xor0 = f_arrdiv16_mux2to179_xor0 ^ b[5];
  assign f_arrdiv16_fs101_not0 = ~f_arrdiv16_mux2to179_xor0;
  assign f_arrdiv16_fs101_and0 = f_arrdiv16_fs101_not0 & b[5];
  assign f_arrdiv16_fs101_xor1 = f_arrdiv16_fs100_or0 ^ f_arrdiv16_fs101_xor0;
  assign f_arrdiv16_fs101_not1 = ~f_arrdiv16_fs101_xor0;
  assign f_arrdiv16_fs101_and1 = f_arrdiv16_fs101_not1 & f_arrdiv16_fs100_or0;
  assign f_arrdiv16_fs101_or0 = f_arrdiv16_fs101_and1 | f_arrdiv16_fs101_and0;
  assign f_arrdiv16_fs102_xor0 = f_arrdiv16_mux2to180_xor0 ^ b[6];
  assign f_arrdiv16_fs102_not0 = ~f_arrdiv16_mux2to180_xor0;
  assign f_arrdiv16_fs102_and0 = f_arrdiv16_fs102_not0 & b[6];
  assign f_arrdiv16_fs102_xor1 = f_arrdiv16_fs101_or0 ^ f_arrdiv16_fs102_xor0;
  assign f_arrdiv16_fs102_not1 = ~f_arrdiv16_fs102_xor0;
  assign f_arrdiv16_fs102_and1 = f_arrdiv16_fs102_not1 & f_arrdiv16_fs101_or0;
  assign f_arrdiv16_fs102_or0 = f_arrdiv16_fs102_and1 | f_arrdiv16_fs102_and0;
  assign f_arrdiv16_fs103_xor0 = f_arrdiv16_mux2to181_xor0 ^ b[7];
  assign f_arrdiv16_fs103_not0 = ~f_arrdiv16_mux2to181_xor0;
  assign f_arrdiv16_fs103_and0 = f_arrdiv16_fs103_not0 & b[7];
  assign f_arrdiv16_fs103_xor1 = f_arrdiv16_fs102_or0 ^ f_arrdiv16_fs103_xor0;
  assign f_arrdiv16_fs103_not1 = ~f_arrdiv16_fs103_xor0;
  assign f_arrdiv16_fs103_and1 = f_arrdiv16_fs103_not1 & f_arrdiv16_fs102_or0;
  assign f_arrdiv16_fs103_or0 = f_arrdiv16_fs103_and1 | f_arrdiv16_fs103_and0;
  assign f_arrdiv16_fs104_xor0 = f_arrdiv16_mux2to182_xor0 ^ b[8];
  assign f_arrdiv16_fs104_not0 = ~f_arrdiv16_mux2to182_xor0;
  assign f_arrdiv16_fs104_and0 = f_arrdiv16_fs104_not0 & b[8];
  assign f_arrdiv16_fs104_xor1 = f_arrdiv16_fs103_or0 ^ f_arrdiv16_fs104_xor0;
  assign f_arrdiv16_fs104_not1 = ~f_arrdiv16_fs104_xor0;
  assign f_arrdiv16_fs104_and1 = f_arrdiv16_fs104_not1 & f_arrdiv16_fs103_or0;
  assign f_arrdiv16_fs104_or0 = f_arrdiv16_fs104_and1 | f_arrdiv16_fs104_and0;
  assign f_arrdiv16_fs105_xor0 = f_arrdiv16_mux2to183_xor0 ^ b[9];
  assign f_arrdiv16_fs105_not0 = ~f_arrdiv16_mux2to183_xor0;
  assign f_arrdiv16_fs105_and0 = f_arrdiv16_fs105_not0 & b[9];
  assign f_arrdiv16_fs105_xor1 = f_arrdiv16_fs104_or0 ^ f_arrdiv16_fs105_xor0;
  assign f_arrdiv16_fs105_not1 = ~f_arrdiv16_fs105_xor0;
  assign f_arrdiv16_fs105_and1 = f_arrdiv16_fs105_not1 & f_arrdiv16_fs104_or0;
  assign f_arrdiv16_fs105_or0 = f_arrdiv16_fs105_and1 | f_arrdiv16_fs105_and0;
  assign f_arrdiv16_fs106_xor0 = f_arrdiv16_mux2to184_xor0 ^ b[10];
  assign f_arrdiv16_fs106_not0 = ~f_arrdiv16_mux2to184_xor0;
  assign f_arrdiv16_fs106_and0 = f_arrdiv16_fs106_not0 & b[10];
  assign f_arrdiv16_fs106_xor1 = f_arrdiv16_fs105_or0 ^ f_arrdiv16_fs106_xor0;
  assign f_arrdiv16_fs106_not1 = ~f_arrdiv16_fs106_xor0;
  assign f_arrdiv16_fs106_and1 = f_arrdiv16_fs106_not1 & f_arrdiv16_fs105_or0;
  assign f_arrdiv16_fs106_or0 = f_arrdiv16_fs106_and1 | f_arrdiv16_fs106_and0;
  assign f_arrdiv16_fs107_xor0 = f_arrdiv16_mux2to185_xor0 ^ b[11];
  assign f_arrdiv16_fs107_not0 = ~f_arrdiv16_mux2to185_xor0;
  assign f_arrdiv16_fs107_and0 = f_arrdiv16_fs107_not0 & b[11];
  assign f_arrdiv16_fs107_xor1 = f_arrdiv16_fs106_or0 ^ f_arrdiv16_fs107_xor0;
  assign f_arrdiv16_fs107_not1 = ~f_arrdiv16_fs107_xor0;
  assign f_arrdiv16_fs107_and1 = f_arrdiv16_fs107_not1 & f_arrdiv16_fs106_or0;
  assign f_arrdiv16_fs107_or0 = f_arrdiv16_fs107_and1 | f_arrdiv16_fs107_and0;
  assign f_arrdiv16_fs108_xor0 = f_arrdiv16_mux2to186_xor0 ^ b[12];
  assign f_arrdiv16_fs108_not0 = ~f_arrdiv16_mux2to186_xor0;
  assign f_arrdiv16_fs108_and0 = f_arrdiv16_fs108_not0 & b[12];
  assign f_arrdiv16_fs108_xor1 = f_arrdiv16_fs107_or0 ^ f_arrdiv16_fs108_xor0;
  assign f_arrdiv16_fs108_not1 = ~f_arrdiv16_fs108_xor0;
  assign f_arrdiv16_fs108_and1 = f_arrdiv16_fs108_not1 & f_arrdiv16_fs107_or0;
  assign f_arrdiv16_fs108_or0 = f_arrdiv16_fs108_and1 | f_arrdiv16_fs108_and0;
  assign f_arrdiv16_fs109_xor0 = f_arrdiv16_mux2to187_xor0 ^ b[13];
  assign f_arrdiv16_fs109_not0 = ~f_arrdiv16_mux2to187_xor0;
  assign f_arrdiv16_fs109_and0 = f_arrdiv16_fs109_not0 & b[13];
  assign f_arrdiv16_fs109_xor1 = f_arrdiv16_fs108_or0 ^ f_arrdiv16_fs109_xor0;
  assign f_arrdiv16_fs109_not1 = ~f_arrdiv16_fs109_xor0;
  assign f_arrdiv16_fs109_and1 = f_arrdiv16_fs109_not1 & f_arrdiv16_fs108_or0;
  assign f_arrdiv16_fs109_or0 = f_arrdiv16_fs109_and1 | f_arrdiv16_fs109_and0;
  assign f_arrdiv16_fs110_xor0 = f_arrdiv16_mux2to188_xor0 ^ b[14];
  assign f_arrdiv16_fs110_not0 = ~f_arrdiv16_mux2to188_xor0;
  assign f_arrdiv16_fs110_and0 = f_arrdiv16_fs110_not0 & b[14];
  assign f_arrdiv16_fs110_xor1 = f_arrdiv16_fs109_or0 ^ f_arrdiv16_fs110_xor0;
  assign f_arrdiv16_fs110_not1 = ~f_arrdiv16_fs110_xor0;
  assign f_arrdiv16_fs110_and1 = f_arrdiv16_fs110_not1 & f_arrdiv16_fs109_or0;
  assign f_arrdiv16_fs110_or0 = f_arrdiv16_fs110_and1 | f_arrdiv16_fs110_and0;
  assign f_arrdiv16_fs111_xor0 = f_arrdiv16_mux2to189_xor0 ^ b[15];
  assign f_arrdiv16_fs111_not0 = ~f_arrdiv16_mux2to189_xor0;
  assign f_arrdiv16_fs111_and0 = f_arrdiv16_fs111_not0 & b[15];
  assign f_arrdiv16_fs111_xor1 = f_arrdiv16_fs110_or0 ^ f_arrdiv16_fs111_xor0;
  assign f_arrdiv16_fs111_not1 = ~f_arrdiv16_fs111_xor0;
  assign f_arrdiv16_fs111_and1 = f_arrdiv16_fs111_not1 & f_arrdiv16_fs110_or0;
  assign f_arrdiv16_fs111_or0 = f_arrdiv16_fs111_and1 | f_arrdiv16_fs111_and0;
  assign f_arrdiv16_mux2to190_and0 = a[9] & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to190_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to190_and1 = f_arrdiv16_fs96_xor0 & f_arrdiv16_mux2to190_not0;
  assign f_arrdiv16_mux2to190_xor0 = f_arrdiv16_mux2to190_and0 ^ f_arrdiv16_mux2to190_and1;
  assign f_arrdiv16_mux2to191_and0 = f_arrdiv16_mux2to175_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to191_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to191_and1 = f_arrdiv16_fs97_xor1 & f_arrdiv16_mux2to191_not0;
  assign f_arrdiv16_mux2to191_xor0 = f_arrdiv16_mux2to191_and0 ^ f_arrdiv16_mux2to191_and1;
  assign f_arrdiv16_mux2to192_and0 = f_arrdiv16_mux2to176_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to192_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to192_and1 = f_arrdiv16_fs98_xor1 & f_arrdiv16_mux2to192_not0;
  assign f_arrdiv16_mux2to192_xor0 = f_arrdiv16_mux2to192_and0 ^ f_arrdiv16_mux2to192_and1;
  assign f_arrdiv16_mux2to193_and0 = f_arrdiv16_mux2to177_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to193_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to193_and1 = f_arrdiv16_fs99_xor1 & f_arrdiv16_mux2to193_not0;
  assign f_arrdiv16_mux2to193_xor0 = f_arrdiv16_mux2to193_and0 ^ f_arrdiv16_mux2to193_and1;
  assign f_arrdiv16_mux2to194_and0 = f_arrdiv16_mux2to178_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to194_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to194_and1 = f_arrdiv16_fs100_xor1 & f_arrdiv16_mux2to194_not0;
  assign f_arrdiv16_mux2to194_xor0 = f_arrdiv16_mux2to194_and0 ^ f_arrdiv16_mux2to194_and1;
  assign f_arrdiv16_mux2to195_and0 = f_arrdiv16_mux2to179_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to195_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to195_and1 = f_arrdiv16_fs101_xor1 & f_arrdiv16_mux2to195_not0;
  assign f_arrdiv16_mux2to195_xor0 = f_arrdiv16_mux2to195_and0 ^ f_arrdiv16_mux2to195_and1;
  assign f_arrdiv16_mux2to196_and0 = f_arrdiv16_mux2to180_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to196_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to196_and1 = f_arrdiv16_fs102_xor1 & f_arrdiv16_mux2to196_not0;
  assign f_arrdiv16_mux2to196_xor0 = f_arrdiv16_mux2to196_and0 ^ f_arrdiv16_mux2to196_and1;
  assign f_arrdiv16_mux2to197_and0 = f_arrdiv16_mux2to181_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to197_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to197_and1 = f_arrdiv16_fs103_xor1 & f_arrdiv16_mux2to197_not0;
  assign f_arrdiv16_mux2to197_xor0 = f_arrdiv16_mux2to197_and0 ^ f_arrdiv16_mux2to197_and1;
  assign f_arrdiv16_mux2to198_and0 = f_arrdiv16_mux2to182_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to198_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to198_and1 = f_arrdiv16_fs104_xor1 & f_arrdiv16_mux2to198_not0;
  assign f_arrdiv16_mux2to198_xor0 = f_arrdiv16_mux2to198_and0 ^ f_arrdiv16_mux2to198_and1;
  assign f_arrdiv16_mux2to199_and0 = f_arrdiv16_mux2to183_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to199_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to199_and1 = f_arrdiv16_fs105_xor1 & f_arrdiv16_mux2to199_not0;
  assign f_arrdiv16_mux2to199_xor0 = f_arrdiv16_mux2to199_and0 ^ f_arrdiv16_mux2to199_and1;
  assign f_arrdiv16_mux2to1100_and0 = f_arrdiv16_mux2to184_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1100_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1100_and1 = f_arrdiv16_fs106_xor1 & f_arrdiv16_mux2to1100_not0;
  assign f_arrdiv16_mux2to1100_xor0 = f_arrdiv16_mux2to1100_and0 ^ f_arrdiv16_mux2to1100_and1;
  assign f_arrdiv16_mux2to1101_and0 = f_arrdiv16_mux2to185_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1101_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1101_and1 = f_arrdiv16_fs107_xor1 & f_arrdiv16_mux2to1101_not0;
  assign f_arrdiv16_mux2to1101_xor0 = f_arrdiv16_mux2to1101_and0 ^ f_arrdiv16_mux2to1101_and1;
  assign f_arrdiv16_mux2to1102_and0 = f_arrdiv16_mux2to186_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1102_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1102_and1 = f_arrdiv16_fs108_xor1 & f_arrdiv16_mux2to1102_not0;
  assign f_arrdiv16_mux2to1102_xor0 = f_arrdiv16_mux2to1102_and0 ^ f_arrdiv16_mux2to1102_and1;
  assign f_arrdiv16_mux2to1103_and0 = f_arrdiv16_mux2to187_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1103_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1103_and1 = f_arrdiv16_fs109_xor1 & f_arrdiv16_mux2to1103_not0;
  assign f_arrdiv16_mux2to1103_xor0 = f_arrdiv16_mux2to1103_and0 ^ f_arrdiv16_mux2to1103_and1;
  assign f_arrdiv16_mux2to1104_and0 = f_arrdiv16_mux2to188_xor0 & f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1104_not0 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_mux2to1104_and1 = f_arrdiv16_fs110_xor1 & f_arrdiv16_mux2to1104_not0;
  assign f_arrdiv16_mux2to1104_xor0 = f_arrdiv16_mux2to1104_and0 ^ f_arrdiv16_mux2to1104_and1;
  assign f_arrdiv16_not6 = ~f_arrdiv16_fs111_or0;
  assign f_arrdiv16_fs112_xor0 = a[8] ^ b[0];
  assign f_arrdiv16_fs112_not0 = ~a[8];
  assign f_arrdiv16_fs112_and0 = f_arrdiv16_fs112_not0 & b[0];
  assign f_arrdiv16_fs112_not1 = ~f_arrdiv16_fs112_xor0;
  assign f_arrdiv16_fs113_xor0 = f_arrdiv16_mux2to190_xor0 ^ b[1];
  assign f_arrdiv16_fs113_not0 = ~f_arrdiv16_mux2to190_xor0;
  assign f_arrdiv16_fs113_and0 = f_arrdiv16_fs113_not0 & b[1];
  assign f_arrdiv16_fs113_xor1 = f_arrdiv16_fs112_and0 ^ f_arrdiv16_fs113_xor0;
  assign f_arrdiv16_fs113_not1 = ~f_arrdiv16_fs113_xor0;
  assign f_arrdiv16_fs113_and1 = f_arrdiv16_fs113_not1 & f_arrdiv16_fs112_and0;
  assign f_arrdiv16_fs113_or0 = f_arrdiv16_fs113_and1 | f_arrdiv16_fs113_and0;
  assign f_arrdiv16_fs114_xor0 = f_arrdiv16_mux2to191_xor0 ^ b[2];
  assign f_arrdiv16_fs114_not0 = ~f_arrdiv16_mux2to191_xor0;
  assign f_arrdiv16_fs114_and0 = f_arrdiv16_fs114_not0 & b[2];
  assign f_arrdiv16_fs114_xor1 = f_arrdiv16_fs113_or0 ^ f_arrdiv16_fs114_xor0;
  assign f_arrdiv16_fs114_not1 = ~f_arrdiv16_fs114_xor0;
  assign f_arrdiv16_fs114_and1 = f_arrdiv16_fs114_not1 & f_arrdiv16_fs113_or0;
  assign f_arrdiv16_fs114_or0 = f_arrdiv16_fs114_and1 | f_arrdiv16_fs114_and0;
  assign f_arrdiv16_fs115_xor0 = f_arrdiv16_mux2to192_xor0 ^ b[3];
  assign f_arrdiv16_fs115_not0 = ~f_arrdiv16_mux2to192_xor0;
  assign f_arrdiv16_fs115_and0 = f_arrdiv16_fs115_not0 & b[3];
  assign f_arrdiv16_fs115_xor1 = f_arrdiv16_fs114_or0 ^ f_arrdiv16_fs115_xor0;
  assign f_arrdiv16_fs115_not1 = ~f_arrdiv16_fs115_xor0;
  assign f_arrdiv16_fs115_and1 = f_arrdiv16_fs115_not1 & f_arrdiv16_fs114_or0;
  assign f_arrdiv16_fs115_or0 = f_arrdiv16_fs115_and1 | f_arrdiv16_fs115_and0;
  assign f_arrdiv16_fs116_xor0 = f_arrdiv16_mux2to193_xor0 ^ b[4];
  assign f_arrdiv16_fs116_not0 = ~f_arrdiv16_mux2to193_xor0;
  assign f_arrdiv16_fs116_and0 = f_arrdiv16_fs116_not0 & b[4];
  assign f_arrdiv16_fs116_xor1 = f_arrdiv16_fs115_or0 ^ f_arrdiv16_fs116_xor0;
  assign f_arrdiv16_fs116_not1 = ~f_arrdiv16_fs116_xor0;
  assign f_arrdiv16_fs116_and1 = f_arrdiv16_fs116_not1 & f_arrdiv16_fs115_or0;
  assign f_arrdiv16_fs116_or0 = f_arrdiv16_fs116_and1 | f_arrdiv16_fs116_and0;
  assign f_arrdiv16_fs117_xor0 = f_arrdiv16_mux2to194_xor0 ^ b[5];
  assign f_arrdiv16_fs117_not0 = ~f_arrdiv16_mux2to194_xor0;
  assign f_arrdiv16_fs117_and0 = f_arrdiv16_fs117_not0 & b[5];
  assign f_arrdiv16_fs117_xor1 = f_arrdiv16_fs116_or0 ^ f_arrdiv16_fs117_xor0;
  assign f_arrdiv16_fs117_not1 = ~f_arrdiv16_fs117_xor0;
  assign f_arrdiv16_fs117_and1 = f_arrdiv16_fs117_not1 & f_arrdiv16_fs116_or0;
  assign f_arrdiv16_fs117_or0 = f_arrdiv16_fs117_and1 | f_arrdiv16_fs117_and0;
  assign f_arrdiv16_fs118_xor0 = f_arrdiv16_mux2to195_xor0 ^ b[6];
  assign f_arrdiv16_fs118_not0 = ~f_arrdiv16_mux2to195_xor0;
  assign f_arrdiv16_fs118_and0 = f_arrdiv16_fs118_not0 & b[6];
  assign f_arrdiv16_fs118_xor1 = f_arrdiv16_fs117_or0 ^ f_arrdiv16_fs118_xor0;
  assign f_arrdiv16_fs118_not1 = ~f_arrdiv16_fs118_xor0;
  assign f_arrdiv16_fs118_and1 = f_arrdiv16_fs118_not1 & f_arrdiv16_fs117_or0;
  assign f_arrdiv16_fs118_or0 = f_arrdiv16_fs118_and1 | f_arrdiv16_fs118_and0;
  assign f_arrdiv16_fs119_xor0 = f_arrdiv16_mux2to196_xor0 ^ b[7];
  assign f_arrdiv16_fs119_not0 = ~f_arrdiv16_mux2to196_xor0;
  assign f_arrdiv16_fs119_and0 = f_arrdiv16_fs119_not0 & b[7];
  assign f_arrdiv16_fs119_xor1 = f_arrdiv16_fs118_or0 ^ f_arrdiv16_fs119_xor0;
  assign f_arrdiv16_fs119_not1 = ~f_arrdiv16_fs119_xor0;
  assign f_arrdiv16_fs119_and1 = f_arrdiv16_fs119_not1 & f_arrdiv16_fs118_or0;
  assign f_arrdiv16_fs119_or0 = f_arrdiv16_fs119_and1 | f_arrdiv16_fs119_and0;
  assign f_arrdiv16_fs120_xor0 = f_arrdiv16_mux2to197_xor0 ^ b[8];
  assign f_arrdiv16_fs120_not0 = ~f_arrdiv16_mux2to197_xor0;
  assign f_arrdiv16_fs120_and0 = f_arrdiv16_fs120_not0 & b[8];
  assign f_arrdiv16_fs120_xor1 = f_arrdiv16_fs119_or0 ^ f_arrdiv16_fs120_xor0;
  assign f_arrdiv16_fs120_not1 = ~f_arrdiv16_fs120_xor0;
  assign f_arrdiv16_fs120_and1 = f_arrdiv16_fs120_not1 & f_arrdiv16_fs119_or0;
  assign f_arrdiv16_fs120_or0 = f_arrdiv16_fs120_and1 | f_arrdiv16_fs120_and0;
  assign f_arrdiv16_fs121_xor0 = f_arrdiv16_mux2to198_xor0 ^ b[9];
  assign f_arrdiv16_fs121_not0 = ~f_arrdiv16_mux2to198_xor0;
  assign f_arrdiv16_fs121_and0 = f_arrdiv16_fs121_not0 & b[9];
  assign f_arrdiv16_fs121_xor1 = f_arrdiv16_fs120_or0 ^ f_arrdiv16_fs121_xor0;
  assign f_arrdiv16_fs121_not1 = ~f_arrdiv16_fs121_xor0;
  assign f_arrdiv16_fs121_and1 = f_arrdiv16_fs121_not1 & f_arrdiv16_fs120_or0;
  assign f_arrdiv16_fs121_or0 = f_arrdiv16_fs121_and1 | f_arrdiv16_fs121_and0;
  assign f_arrdiv16_fs122_xor0 = f_arrdiv16_mux2to199_xor0 ^ b[10];
  assign f_arrdiv16_fs122_not0 = ~f_arrdiv16_mux2to199_xor0;
  assign f_arrdiv16_fs122_and0 = f_arrdiv16_fs122_not0 & b[10];
  assign f_arrdiv16_fs122_xor1 = f_arrdiv16_fs121_or0 ^ f_arrdiv16_fs122_xor0;
  assign f_arrdiv16_fs122_not1 = ~f_arrdiv16_fs122_xor0;
  assign f_arrdiv16_fs122_and1 = f_arrdiv16_fs122_not1 & f_arrdiv16_fs121_or0;
  assign f_arrdiv16_fs122_or0 = f_arrdiv16_fs122_and1 | f_arrdiv16_fs122_and0;
  assign f_arrdiv16_fs123_xor0 = f_arrdiv16_mux2to1100_xor0 ^ b[11];
  assign f_arrdiv16_fs123_not0 = ~f_arrdiv16_mux2to1100_xor0;
  assign f_arrdiv16_fs123_and0 = f_arrdiv16_fs123_not0 & b[11];
  assign f_arrdiv16_fs123_xor1 = f_arrdiv16_fs122_or0 ^ f_arrdiv16_fs123_xor0;
  assign f_arrdiv16_fs123_not1 = ~f_arrdiv16_fs123_xor0;
  assign f_arrdiv16_fs123_and1 = f_arrdiv16_fs123_not1 & f_arrdiv16_fs122_or0;
  assign f_arrdiv16_fs123_or0 = f_arrdiv16_fs123_and1 | f_arrdiv16_fs123_and0;
  assign f_arrdiv16_fs124_xor0 = f_arrdiv16_mux2to1101_xor0 ^ b[12];
  assign f_arrdiv16_fs124_not0 = ~f_arrdiv16_mux2to1101_xor0;
  assign f_arrdiv16_fs124_and0 = f_arrdiv16_fs124_not0 & b[12];
  assign f_arrdiv16_fs124_xor1 = f_arrdiv16_fs123_or0 ^ f_arrdiv16_fs124_xor0;
  assign f_arrdiv16_fs124_not1 = ~f_arrdiv16_fs124_xor0;
  assign f_arrdiv16_fs124_and1 = f_arrdiv16_fs124_not1 & f_arrdiv16_fs123_or0;
  assign f_arrdiv16_fs124_or0 = f_arrdiv16_fs124_and1 | f_arrdiv16_fs124_and0;
  assign f_arrdiv16_fs125_xor0 = f_arrdiv16_mux2to1102_xor0 ^ b[13];
  assign f_arrdiv16_fs125_not0 = ~f_arrdiv16_mux2to1102_xor0;
  assign f_arrdiv16_fs125_and0 = f_arrdiv16_fs125_not0 & b[13];
  assign f_arrdiv16_fs125_xor1 = f_arrdiv16_fs124_or0 ^ f_arrdiv16_fs125_xor0;
  assign f_arrdiv16_fs125_not1 = ~f_arrdiv16_fs125_xor0;
  assign f_arrdiv16_fs125_and1 = f_arrdiv16_fs125_not1 & f_arrdiv16_fs124_or0;
  assign f_arrdiv16_fs125_or0 = f_arrdiv16_fs125_and1 | f_arrdiv16_fs125_and0;
  assign f_arrdiv16_fs126_xor0 = f_arrdiv16_mux2to1103_xor0 ^ b[14];
  assign f_arrdiv16_fs126_not0 = ~f_arrdiv16_mux2to1103_xor0;
  assign f_arrdiv16_fs126_and0 = f_arrdiv16_fs126_not0 & b[14];
  assign f_arrdiv16_fs126_xor1 = f_arrdiv16_fs125_or0 ^ f_arrdiv16_fs126_xor0;
  assign f_arrdiv16_fs126_not1 = ~f_arrdiv16_fs126_xor0;
  assign f_arrdiv16_fs126_and1 = f_arrdiv16_fs126_not1 & f_arrdiv16_fs125_or0;
  assign f_arrdiv16_fs126_or0 = f_arrdiv16_fs126_and1 | f_arrdiv16_fs126_and0;
  assign f_arrdiv16_fs127_xor0 = f_arrdiv16_mux2to1104_xor0 ^ b[15];
  assign f_arrdiv16_fs127_not0 = ~f_arrdiv16_mux2to1104_xor0;
  assign f_arrdiv16_fs127_and0 = f_arrdiv16_fs127_not0 & b[15];
  assign f_arrdiv16_fs127_xor1 = f_arrdiv16_fs126_or0 ^ f_arrdiv16_fs127_xor0;
  assign f_arrdiv16_fs127_not1 = ~f_arrdiv16_fs127_xor0;
  assign f_arrdiv16_fs127_and1 = f_arrdiv16_fs127_not1 & f_arrdiv16_fs126_or0;
  assign f_arrdiv16_fs127_or0 = f_arrdiv16_fs127_and1 | f_arrdiv16_fs127_and0;
  assign f_arrdiv16_mux2to1105_and0 = a[8] & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1105_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1105_and1 = f_arrdiv16_fs112_xor0 & f_arrdiv16_mux2to1105_not0;
  assign f_arrdiv16_mux2to1105_xor0 = f_arrdiv16_mux2to1105_and0 ^ f_arrdiv16_mux2to1105_and1;
  assign f_arrdiv16_mux2to1106_and0 = f_arrdiv16_mux2to190_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1106_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1106_and1 = f_arrdiv16_fs113_xor1 & f_arrdiv16_mux2to1106_not0;
  assign f_arrdiv16_mux2to1106_xor0 = f_arrdiv16_mux2to1106_and0 ^ f_arrdiv16_mux2to1106_and1;
  assign f_arrdiv16_mux2to1107_and0 = f_arrdiv16_mux2to191_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1107_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1107_and1 = f_arrdiv16_fs114_xor1 & f_arrdiv16_mux2to1107_not0;
  assign f_arrdiv16_mux2to1107_xor0 = f_arrdiv16_mux2to1107_and0 ^ f_arrdiv16_mux2to1107_and1;
  assign f_arrdiv16_mux2to1108_and0 = f_arrdiv16_mux2to192_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1108_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1108_and1 = f_arrdiv16_fs115_xor1 & f_arrdiv16_mux2to1108_not0;
  assign f_arrdiv16_mux2to1108_xor0 = f_arrdiv16_mux2to1108_and0 ^ f_arrdiv16_mux2to1108_and1;
  assign f_arrdiv16_mux2to1109_and0 = f_arrdiv16_mux2to193_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1109_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1109_and1 = f_arrdiv16_fs116_xor1 & f_arrdiv16_mux2to1109_not0;
  assign f_arrdiv16_mux2to1109_xor0 = f_arrdiv16_mux2to1109_and0 ^ f_arrdiv16_mux2to1109_and1;
  assign f_arrdiv16_mux2to1110_and0 = f_arrdiv16_mux2to194_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1110_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1110_and1 = f_arrdiv16_fs117_xor1 & f_arrdiv16_mux2to1110_not0;
  assign f_arrdiv16_mux2to1110_xor0 = f_arrdiv16_mux2to1110_and0 ^ f_arrdiv16_mux2to1110_and1;
  assign f_arrdiv16_mux2to1111_and0 = f_arrdiv16_mux2to195_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1111_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1111_and1 = f_arrdiv16_fs118_xor1 & f_arrdiv16_mux2to1111_not0;
  assign f_arrdiv16_mux2to1111_xor0 = f_arrdiv16_mux2to1111_and0 ^ f_arrdiv16_mux2to1111_and1;
  assign f_arrdiv16_mux2to1112_and0 = f_arrdiv16_mux2to196_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1112_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1112_and1 = f_arrdiv16_fs119_xor1 & f_arrdiv16_mux2to1112_not0;
  assign f_arrdiv16_mux2to1112_xor0 = f_arrdiv16_mux2to1112_and0 ^ f_arrdiv16_mux2to1112_and1;
  assign f_arrdiv16_mux2to1113_and0 = f_arrdiv16_mux2to197_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1113_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1113_and1 = f_arrdiv16_fs120_xor1 & f_arrdiv16_mux2to1113_not0;
  assign f_arrdiv16_mux2to1113_xor0 = f_arrdiv16_mux2to1113_and0 ^ f_arrdiv16_mux2to1113_and1;
  assign f_arrdiv16_mux2to1114_and0 = f_arrdiv16_mux2to198_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1114_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1114_and1 = f_arrdiv16_fs121_xor1 & f_arrdiv16_mux2to1114_not0;
  assign f_arrdiv16_mux2to1114_xor0 = f_arrdiv16_mux2to1114_and0 ^ f_arrdiv16_mux2to1114_and1;
  assign f_arrdiv16_mux2to1115_and0 = f_arrdiv16_mux2to199_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1115_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1115_and1 = f_arrdiv16_fs122_xor1 & f_arrdiv16_mux2to1115_not0;
  assign f_arrdiv16_mux2to1115_xor0 = f_arrdiv16_mux2to1115_and0 ^ f_arrdiv16_mux2to1115_and1;
  assign f_arrdiv16_mux2to1116_and0 = f_arrdiv16_mux2to1100_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1116_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1116_and1 = f_arrdiv16_fs123_xor1 & f_arrdiv16_mux2to1116_not0;
  assign f_arrdiv16_mux2to1116_xor0 = f_arrdiv16_mux2to1116_and0 ^ f_arrdiv16_mux2to1116_and1;
  assign f_arrdiv16_mux2to1117_and0 = f_arrdiv16_mux2to1101_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1117_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1117_and1 = f_arrdiv16_fs124_xor1 & f_arrdiv16_mux2to1117_not0;
  assign f_arrdiv16_mux2to1117_xor0 = f_arrdiv16_mux2to1117_and0 ^ f_arrdiv16_mux2to1117_and1;
  assign f_arrdiv16_mux2to1118_and0 = f_arrdiv16_mux2to1102_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1118_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1118_and1 = f_arrdiv16_fs125_xor1 & f_arrdiv16_mux2to1118_not0;
  assign f_arrdiv16_mux2to1118_xor0 = f_arrdiv16_mux2to1118_and0 ^ f_arrdiv16_mux2to1118_and1;
  assign f_arrdiv16_mux2to1119_and0 = f_arrdiv16_mux2to1103_xor0 & f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1119_not0 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_mux2to1119_and1 = f_arrdiv16_fs126_xor1 & f_arrdiv16_mux2to1119_not0;
  assign f_arrdiv16_mux2to1119_xor0 = f_arrdiv16_mux2to1119_and0 ^ f_arrdiv16_mux2to1119_and1;
  assign f_arrdiv16_not7 = ~f_arrdiv16_fs127_or0;
  assign f_arrdiv16_fs128_xor0 = a[7] ^ b[0];
  assign f_arrdiv16_fs128_not0 = ~a[7];
  assign f_arrdiv16_fs128_and0 = f_arrdiv16_fs128_not0 & b[0];
  assign f_arrdiv16_fs128_not1 = ~f_arrdiv16_fs128_xor0;
  assign f_arrdiv16_fs129_xor0 = f_arrdiv16_mux2to1105_xor0 ^ b[1];
  assign f_arrdiv16_fs129_not0 = ~f_arrdiv16_mux2to1105_xor0;
  assign f_arrdiv16_fs129_and0 = f_arrdiv16_fs129_not0 & b[1];
  assign f_arrdiv16_fs129_xor1 = f_arrdiv16_fs128_and0 ^ f_arrdiv16_fs129_xor0;
  assign f_arrdiv16_fs129_not1 = ~f_arrdiv16_fs129_xor0;
  assign f_arrdiv16_fs129_and1 = f_arrdiv16_fs129_not1 & f_arrdiv16_fs128_and0;
  assign f_arrdiv16_fs129_or0 = f_arrdiv16_fs129_and1 | f_arrdiv16_fs129_and0;
  assign f_arrdiv16_fs130_xor0 = f_arrdiv16_mux2to1106_xor0 ^ b[2];
  assign f_arrdiv16_fs130_not0 = ~f_arrdiv16_mux2to1106_xor0;
  assign f_arrdiv16_fs130_and0 = f_arrdiv16_fs130_not0 & b[2];
  assign f_arrdiv16_fs130_xor1 = f_arrdiv16_fs129_or0 ^ f_arrdiv16_fs130_xor0;
  assign f_arrdiv16_fs130_not1 = ~f_arrdiv16_fs130_xor0;
  assign f_arrdiv16_fs130_and1 = f_arrdiv16_fs130_not1 & f_arrdiv16_fs129_or0;
  assign f_arrdiv16_fs130_or0 = f_arrdiv16_fs130_and1 | f_arrdiv16_fs130_and0;
  assign f_arrdiv16_fs131_xor0 = f_arrdiv16_mux2to1107_xor0 ^ b[3];
  assign f_arrdiv16_fs131_not0 = ~f_arrdiv16_mux2to1107_xor0;
  assign f_arrdiv16_fs131_and0 = f_arrdiv16_fs131_not0 & b[3];
  assign f_arrdiv16_fs131_xor1 = f_arrdiv16_fs130_or0 ^ f_arrdiv16_fs131_xor0;
  assign f_arrdiv16_fs131_not1 = ~f_arrdiv16_fs131_xor0;
  assign f_arrdiv16_fs131_and1 = f_arrdiv16_fs131_not1 & f_arrdiv16_fs130_or0;
  assign f_arrdiv16_fs131_or0 = f_arrdiv16_fs131_and1 | f_arrdiv16_fs131_and0;
  assign f_arrdiv16_fs132_xor0 = f_arrdiv16_mux2to1108_xor0 ^ b[4];
  assign f_arrdiv16_fs132_not0 = ~f_arrdiv16_mux2to1108_xor0;
  assign f_arrdiv16_fs132_and0 = f_arrdiv16_fs132_not0 & b[4];
  assign f_arrdiv16_fs132_xor1 = f_arrdiv16_fs131_or0 ^ f_arrdiv16_fs132_xor0;
  assign f_arrdiv16_fs132_not1 = ~f_arrdiv16_fs132_xor0;
  assign f_arrdiv16_fs132_and1 = f_arrdiv16_fs132_not1 & f_arrdiv16_fs131_or0;
  assign f_arrdiv16_fs132_or0 = f_arrdiv16_fs132_and1 | f_arrdiv16_fs132_and0;
  assign f_arrdiv16_fs133_xor0 = f_arrdiv16_mux2to1109_xor0 ^ b[5];
  assign f_arrdiv16_fs133_not0 = ~f_arrdiv16_mux2to1109_xor0;
  assign f_arrdiv16_fs133_and0 = f_arrdiv16_fs133_not0 & b[5];
  assign f_arrdiv16_fs133_xor1 = f_arrdiv16_fs132_or0 ^ f_arrdiv16_fs133_xor0;
  assign f_arrdiv16_fs133_not1 = ~f_arrdiv16_fs133_xor0;
  assign f_arrdiv16_fs133_and1 = f_arrdiv16_fs133_not1 & f_arrdiv16_fs132_or0;
  assign f_arrdiv16_fs133_or0 = f_arrdiv16_fs133_and1 | f_arrdiv16_fs133_and0;
  assign f_arrdiv16_fs134_xor0 = f_arrdiv16_mux2to1110_xor0 ^ b[6];
  assign f_arrdiv16_fs134_not0 = ~f_arrdiv16_mux2to1110_xor0;
  assign f_arrdiv16_fs134_and0 = f_arrdiv16_fs134_not0 & b[6];
  assign f_arrdiv16_fs134_xor1 = f_arrdiv16_fs133_or0 ^ f_arrdiv16_fs134_xor0;
  assign f_arrdiv16_fs134_not1 = ~f_arrdiv16_fs134_xor0;
  assign f_arrdiv16_fs134_and1 = f_arrdiv16_fs134_not1 & f_arrdiv16_fs133_or0;
  assign f_arrdiv16_fs134_or0 = f_arrdiv16_fs134_and1 | f_arrdiv16_fs134_and0;
  assign f_arrdiv16_fs135_xor0 = f_arrdiv16_mux2to1111_xor0 ^ b[7];
  assign f_arrdiv16_fs135_not0 = ~f_arrdiv16_mux2to1111_xor0;
  assign f_arrdiv16_fs135_and0 = f_arrdiv16_fs135_not0 & b[7];
  assign f_arrdiv16_fs135_xor1 = f_arrdiv16_fs134_or0 ^ f_arrdiv16_fs135_xor0;
  assign f_arrdiv16_fs135_not1 = ~f_arrdiv16_fs135_xor0;
  assign f_arrdiv16_fs135_and1 = f_arrdiv16_fs135_not1 & f_arrdiv16_fs134_or0;
  assign f_arrdiv16_fs135_or0 = f_arrdiv16_fs135_and1 | f_arrdiv16_fs135_and0;
  assign f_arrdiv16_fs136_xor0 = f_arrdiv16_mux2to1112_xor0 ^ b[8];
  assign f_arrdiv16_fs136_not0 = ~f_arrdiv16_mux2to1112_xor0;
  assign f_arrdiv16_fs136_and0 = f_arrdiv16_fs136_not0 & b[8];
  assign f_arrdiv16_fs136_xor1 = f_arrdiv16_fs135_or0 ^ f_arrdiv16_fs136_xor0;
  assign f_arrdiv16_fs136_not1 = ~f_arrdiv16_fs136_xor0;
  assign f_arrdiv16_fs136_and1 = f_arrdiv16_fs136_not1 & f_arrdiv16_fs135_or0;
  assign f_arrdiv16_fs136_or0 = f_arrdiv16_fs136_and1 | f_arrdiv16_fs136_and0;
  assign f_arrdiv16_fs137_xor0 = f_arrdiv16_mux2to1113_xor0 ^ b[9];
  assign f_arrdiv16_fs137_not0 = ~f_arrdiv16_mux2to1113_xor0;
  assign f_arrdiv16_fs137_and0 = f_arrdiv16_fs137_not0 & b[9];
  assign f_arrdiv16_fs137_xor1 = f_arrdiv16_fs136_or0 ^ f_arrdiv16_fs137_xor0;
  assign f_arrdiv16_fs137_not1 = ~f_arrdiv16_fs137_xor0;
  assign f_arrdiv16_fs137_and1 = f_arrdiv16_fs137_not1 & f_arrdiv16_fs136_or0;
  assign f_arrdiv16_fs137_or0 = f_arrdiv16_fs137_and1 | f_arrdiv16_fs137_and0;
  assign f_arrdiv16_fs138_xor0 = f_arrdiv16_mux2to1114_xor0 ^ b[10];
  assign f_arrdiv16_fs138_not0 = ~f_arrdiv16_mux2to1114_xor0;
  assign f_arrdiv16_fs138_and0 = f_arrdiv16_fs138_not0 & b[10];
  assign f_arrdiv16_fs138_xor1 = f_arrdiv16_fs137_or0 ^ f_arrdiv16_fs138_xor0;
  assign f_arrdiv16_fs138_not1 = ~f_arrdiv16_fs138_xor0;
  assign f_arrdiv16_fs138_and1 = f_arrdiv16_fs138_not1 & f_arrdiv16_fs137_or0;
  assign f_arrdiv16_fs138_or0 = f_arrdiv16_fs138_and1 | f_arrdiv16_fs138_and0;
  assign f_arrdiv16_fs139_xor0 = f_arrdiv16_mux2to1115_xor0 ^ b[11];
  assign f_arrdiv16_fs139_not0 = ~f_arrdiv16_mux2to1115_xor0;
  assign f_arrdiv16_fs139_and0 = f_arrdiv16_fs139_not0 & b[11];
  assign f_arrdiv16_fs139_xor1 = f_arrdiv16_fs138_or0 ^ f_arrdiv16_fs139_xor0;
  assign f_arrdiv16_fs139_not1 = ~f_arrdiv16_fs139_xor0;
  assign f_arrdiv16_fs139_and1 = f_arrdiv16_fs139_not1 & f_arrdiv16_fs138_or0;
  assign f_arrdiv16_fs139_or0 = f_arrdiv16_fs139_and1 | f_arrdiv16_fs139_and0;
  assign f_arrdiv16_fs140_xor0 = f_arrdiv16_mux2to1116_xor0 ^ b[12];
  assign f_arrdiv16_fs140_not0 = ~f_arrdiv16_mux2to1116_xor0;
  assign f_arrdiv16_fs140_and0 = f_arrdiv16_fs140_not0 & b[12];
  assign f_arrdiv16_fs140_xor1 = f_arrdiv16_fs139_or0 ^ f_arrdiv16_fs140_xor0;
  assign f_arrdiv16_fs140_not1 = ~f_arrdiv16_fs140_xor0;
  assign f_arrdiv16_fs140_and1 = f_arrdiv16_fs140_not1 & f_arrdiv16_fs139_or0;
  assign f_arrdiv16_fs140_or0 = f_arrdiv16_fs140_and1 | f_arrdiv16_fs140_and0;
  assign f_arrdiv16_fs141_xor0 = f_arrdiv16_mux2to1117_xor0 ^ b[13];
  assign f_arrdiv16_fs141_not0 = ~f_arrdiv16_mux2to1117_xor0;
  assign f_arrdiv16_fs141_and0 = f_arrdiv16_fs141_not0 & b[13];
  assign f_arrdiv16_fs141_xor1 = f_arrdiv16_fs140_or0 ^ f_arrdiv16_fs141_xor0;
  assign f_arrdiv16_fs141_not1 = ~f_arrdiv16_fs141_xor0;
  assign f_arrdiv16_fs141_and1 = f_arrdiv16_fs141_not1 & f_arrdiv16_fs140_or0;
  assign f_arrdiv16_fs141_or0 = f_arrdiv16_fs141_and1 | f_arrdiv16_fs141_and0;
  assign f_arrdiv16_fs142_xor0 = f_arrdiv16_mux2to1118_xor0 ^ b[14];
  assign f_arrdiv16_fs142_not0 = ~f_arrdiv16_mux2to1118_xor0;
  assign f_arrdiv16_fs142_and0 = f_arrdiv16_fs142_not0 & b[14];
  assign f_arrdiv16_fs142_xor1 = f_arrdiv16_fs141_or0 ^ f_arrdiv16_fs142_xor0;
  assign f_arrdiv16_fs142_not1 = ~f_arrdiv16_fs142_xor0;
  assign f_arrdiv16_fs142_and1 = f_arrdiv16_fs142_not1 & f_arrdiv16_fs141_or0;
  assign f_arrdiv16_fs142_or0 = f_arrdiv16_fs142_and1 | f_arrdiv16_fs142_and0;
  assign f_arrdiv16_fs143_xor0 = f_arrdiv16_mux2to1119_xor0 ^ b[15];
  assign f_arrdiv16_fs143_not0 = ~f_arrdiv16_mux2to1119_xor0;
  assign f_arrdiv16_fs143_and0 = f_arrdiv16_fs143_not0 & b[15];
  assign f_arrdiv16_fs143_xor1 = f_arrdiv16_fs142_or0 ^ f_arrdiv16_fs143_xor0;
  assign f_arrdiv16_fs143_not1 = ~f_arrdiv16_fs143_xor0;
  assign f_arrdiv16_fs143_and1 = f_arrdiv16_fs143_not1 & f_arrdiv16_fs142_or0;
  assign f_arrdiv16_fs143_or0 = f_arrdiv16_fs143_and1 | f_arrdiv16_fs143_and0;
  assign f_arrdiv16_mux2to1120_and0 = a[7] & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1120_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1120_and1 = f_arrdiv16_fs128_xor0 & f_arrdiv16_mux2to1120_not0;
  assign f_arrdiv16_mux2to1120_xor0 = f_arrdiv16_mux2to1120_and0 ^ f_arrdiv16_mux2to1120_and1;
  assign f_arrdiv16_mux2to1121_and0 = f_arrdiv16_mux2to1105_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1121_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1121_and1 = f_arrdiv16_fs129_xor1 & f_arrdiv16_mux2to1121_not0;
  assign f_arrdiv16_mux2to1121_xor0 = f_arrdiv16_mux2to1121_and0 ^ f_arrdiv16_mux2to1121_and1;
  assign f_arrdiv16_mux2to1122_and0 = f_arrdiv16_mux2to1106_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1122_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1122_and1 = f_arrdiv16_fs130_xor1 & f_arrdiv16_mux2to1122_not0;
  assign f_arrdiv16_mux2to1122_xor0 = f_arrdiv16_mux2to1122_and0 ^ f_arrdiv16_mux2to1122_and1;
  assign f_arrdiv16_mux2to1123_and0 = f_arrdiv16_mux2to1107_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1123_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1123_and1 = f_arrdiv16_fs131_xor1 & f_arrdiv16_mux2to1123_not0;
  assign f_arrdiv16_mux2to1123_xor0 = f_arrdiv16_mux2to1123_and0 ^ f_arrdiv16_mux2to1123_and1;
  assign f_arrdiv16_mux2to1124_and0 = f_arrdiv16_mux2to1108_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1124_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1124_and1 = f_arrdiv16_fs132_xor1 & f_arrdiv16_mux2to1124_not0;
  assign f_arrdiv16_mux2to1124_xor0 = f_arrdiv16_mux2to1124_and0 ^ f_arrdiv16_mux2to1124_and1;
  assign f_arrdiv16_mux2to1125_and0 = f_arrdiv16_mux2to1109_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1125_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1125_and1 = f_arrdiv16_fs133_xor1 & f_arrdiv16_mux2to1125_not0;
  assign f_arrdiv16_mux2to1125_xor0 = f_arrdiv16_mux2to1125_and0 ^ f_arrdiv16_mux2to1125_and1;
  assign f_arrdiv16_mux2to1126_and0 = f_arrdiv16_mux2to1110_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1126_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1126_and1 = f_arrdiv16_fs134_xor1 & f_arrdiv16_mux2to1126_not0;
  assign f_arrdiv16_mux2to1126_xor0 = f_arrdiv16_mux2to1126_and0 ^ f_arrdiv16_mux2to1126_and1;
  assign f_arrdiv16_mux2to1127_and0 = f_arrdiv16_mux2to1111_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1127_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1127_and1 = f_arrdiv16_fs135_xor1 & f_arrdiv16_mux2to1127_not0;
  assign f_arrdiv16_mux2to1127_xor0 = f_arrdiv16_mux2to1127_and0 ^ f_arrdiv16_mux2to1127_and1;
  assign f_arrdiv16_mux2to1128_and0 = f_arrdiv16_mux2to1112_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1128_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1128_and1 = f_arrdiv16_fs136_xor1 & f_arrdiv16_mux2to1128_not0;
  assign f_arrdiv16_mux2to1128_xor0 = f_arrdiv16_mux2to1128_and0 ^ f_arrdiv16_mux2to1128_and1;
  assign f_arrdiv16_mux2to1129_and0 = f_arrdiv16_mux2to1113_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1129_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1129_and1 = f_arrdiv16_fs137_xor1 & f_arrdiv16_mux2to1129_not0;
  assign f_arrdiv16_mux2to1129_xor0 = f_arrdiv16_mux2to1129_and0 ^ f_arrdiv16_mux2to1129_and1;
  assign f_arrdiv16_mux2to1130_and0 = f_arrdiv16_mux2to1114_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1130_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1130_and1 = f_arrdiv16_fs138_xor1 & f_arrdiv16_mux2to1130_not0;
  assign f_arrdiv16_mux2to1130_xor0 = f_arrdiv16_mux2to1130_and0 ^ f_arrdiv16_mux2to1130_and1;
  assign f_arrdiv16_mux2to1131_and0 = f_arrdiv16_mux2to1115_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1131_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1131_and1 = f_arrdiv16_fs139_xor1 & f_arrdiv16_mux2to1131_not0;
  assign f_arrdiv16_mux2to1131_xor0 = f_arrdiv16_mux2to1131_and0 ^ f_arrdiv16_mux2to1131_and1;
  assign f_arrdiv16_mux2to1132_and0 = f_arrdiv16_mux2to1116_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1132_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1132_and1 = f_arrdiv16_fs140_xor1 & f_arrdiv16_mux2to1132_not0;
  assign f_arrdiv16_mux2to1132_xor0 = f_arrdiv16_mux2to1132_and0 ^ f_arrdiv16_mux2to1132_and1;
  assign f_arrdiv16_mux2to1133_and0 = f_arrdiv16_mux2to1117_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1133_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1133_and1 = f_arrdiv16_fs141_xor1 & f_arrdiv16_mux2to1133_not0;
  assign f_arrdiv16_mux2to1133_xor0 = f_arrdiv16_mux2to1133_and0 ^ f_arrdiv16_mux2to1133_and1;
  assign f_arrdiv16_mux2to1134_and0 = f_arrdiv16_mux2to1118_xor0 & f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1134_not0 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_mux2to1134_and1 = f_arrdiv16_fs142_xor1 & f_arrdiv16_mux2to1134_not0;
  assign f_arrdiv16_mux2to1134_xor0 = f_arrdiv16_mux2to1134_and0 ^ f_arrdiv16_mux2to1134_and1;
  assign f_arrdiv16_not8 = ~f_arrdiv16_fs143_or0;
  assign f_arrdiv16_fs144_xor0 = a[6] ^ b[0];
  assign f_arrdiv16_fs144_not0 = ~a[6];
  assign f_arrdiv16_fs144_and0 = f_arrdiv16_fs144_not0 & b[0];
  assign f_arrdiv16_fs144_not1 = ~f_arrdiv16_fs144_xor0;
  assign f_arrdiv16_fs145_xor0 = f_arrdiv16_mux2to1120_xor0 ^ b[1];
  assign f_arrdiv16_fs145_not0 = ~f_arrdiv16_mux2to1120_xor0;
  assign f_arrdiv16_fs145_and0 = f_arrdiv16_fs145_not0 & b[1];
  assign f_arrdiv16_fs145_xor1 = f_arrdiv16_fs144_and0 ^ f_arrdiv16_fs145_xor0;
  assign f_arrdiv16_fs145_not1 = ~f_arrdiv16_fs145_xor0;
  assign f_arrdiv16_fs145_and1 = f_arrdiv16_fs145_not1 & f_arrdiv16_fs144_and0;
  assign f_arrdiv16_fs145_or0 = f_arrdiv16_fs145_and1 | f_arrdiv16_fs145_and0;
  assign f_arrdiv16_fs146_xor0 = f_arrdiv16_mux2to1121_xor0 ^ b[2];
  assign f_arrdiv16_fs146_not0 = ~f_arrdiv16_mux2to1121_xor0;
  assign f_arrdiv16_fs146_and0 = f_arrdiv16_fs146_not0 & b[2];
  assign f_arrdiv16_fs146_xor1 = f_arrdiv16_fs145_or0 ^ f_arrdiv16_fs146_xor0;
  assign f_arrdiv16_fs146_not1 = ~f_arrdiv16_fs146_xor0;
  assign f_arrdiv16_fs146_and1 = f_arrdiv16_fs146_not1 & f_arrdiv16_fs145_or0;
  assign f_arrdiv16_fs146_or0 = f_arrdiv16_fs146_and1 | f_arrdiv16_fs146_and0;
  assign f_arrdiv16_fs147_xor0 = f_arrdiv16_mux2to1122_xor0 ^ b[3];
  assign f_arrdiv16_fs147_not0 = ~f_arrdiv16_mux2to1122_xor0;
  assign f_arrdiv16_fs147_and0 = f_arrdiv16_fs147_not0 & b[3];
  assign f_arrdiv16_fs147_xor1 = f_arrdiv16_fs146_or0 ^ f_arrdiv16_fs147_xor0;
  assign f_arrdiv16_fs147_not1 = ~f_arrdiv16_fs147_xor0;
  assign f_arrdiv16_fs147_and1 = f_arrdiv16_fs147_not1 & f_arrdiv16_fs146_or0;
  assign f_arrdiv16_fs147_or0 = f_arrdiv16_fs147_and1 | f_arrdiv16_fs147_and0;
  assign f_arrdiv16_fs148_xor0 = f_arrdiv16_mux2to1123_xor0 ^ b[4];
  assign f_arrdiv16_fs148_not0 = ~f_arrdiv16_mux2to1123_xor0;
  assign f_arrdiv16_fs148_and0 = f_arrdiv16_fs148_not0 & b[4];
  assign f_arrdiv16_fs148_xor1 = f_arrdiv16_fs147_or0 ^ f_arrdiv16_fs148_xor0;
  assign f_arrdiv16_fs148_not1 = ~f_arrdiv16_fs148_xor0;
  assign f_arrdiv16_fs148_and1 = f_arrdiv16_fs148_not1 & f_arrdiv16_fs147_or0;
  assign f_arrdiv16_fs148_or0 = f_arrdiv16_fs148_and1 | f_arrdiv16_fs148_and0;
  assign f_arrdiv16_fs149_xor0 = f_arrdiv16_mux2to1124_xor0 ^ b[5];
  assign f_arrdiv16_fs149_not0 = ~f_arrdiv16_mux2to1124_xor0;
  assign f_arrdiv16_fs149_and0 = f_arrdiv16_fs149_not0 & b[5];
  assign f_arrdiv16_fs149_xor1 = f_arrdiv16_fs148_or0 ^ f_arrdiv16_fs149_xor0;
  assign f_arrdiv16_fs149_not1 = ~f_arrdiv16_fs149_xor0;
  assign f_arrdiv16_fs149_and1 = f_arrdiv16_fs149_not1 & f_arrdiv16_fs148_or0;
  assign f_arrdiv16_fs149_or0 = f_arrdiv16_fs149_and1 | f_arrdiv16_fs149_and0;
  assign f_arrdiv16_fs150_xor0 = f_arrdiv16_mux2to1125_xor0 ^ b[6];
  assign f_arrdiv16_fs150_not0 = ~f_arrdiv16_mux2to1125_xor0;
  assign f_arrdiv16_fs150_and0 = f_arrdiv16_fs150_not0 & b[6];
  assign f_arrdiv16_fs150_xor1 = f_arrdiv16_fs149_or0 ^ f_arrdiv16_fs150_xor0;
  assign f_arrdiv16_fs150_not1 = ~f_arrdiv16_fs150_xor0;
  assign f_arrdiv16_fs150_and1 = f_arrdiv16_fs150_not1 & f_arrdiv16_fs149_or0;
  assign f_arrdiv16_fs150_or0 = f_arrdiv16_fs150_and1 | f_arrdiv16_fs150_and0;
  assign f_arrdiv16_fs151_xor0 = f_arrdiv16_mux2to1126_xor0 ^ b[7];
  assign f_arrdiv16_fs151_not0 = ~f_arrdiv16_mux2to1126_xor0;
  assign f_arrdiv16_fs151_and0 = f_arrdiv16_fs151_not0 & b[7];
  assign f_arrdiv16_fs151_xor1 = f_arrdiv16_fs150_or0 ^ f_arrdiv16_fs151_xor0;
  assign f_arrdiv16_fs151_not1 = ~f_arrdiv16_fs151_xor0;
  assign f_arrdiv16_fs151_and1 = f_arrdiv16_fs151_not1 & f_arrdiv16_fs150_or0;
  assign f_arrdiv16_fs151_or0 = f_arrdiv16_fs151_and1 | f_arrdiv16_fs151_and0;
  assign f_arrdiv16_fs152_xor0 = f_arrdiv16_mux2to1127_xor0 ^ b[8];
  assign f_arrdiv16_fs152_not0 = ~f_arrdiv16_mux2to1127_xor0;
  assign f_arrdiv16_fs152_and0 = f_arrdiv16_fs152_not0 & b[8];
  assign f_arrdiv16_fs152_xor1 = f_arrdiv16_fs151_or0 ^ f_arrdiv16_fs152_xor0;
  assign f_arrdiv16_fs152_not1 = ~f_arrdiv16_fs152_xor0;
  assign f_arrdiv16_fs152_and1 = f_arrdiv16_fs152_not1 & f_arrdiv16_fs151_or0;
  assign f_arrdiv16_fs152_or0 = f_arrdiv16_fs152_and1 | f_arrdiv16_fs152_and0;
  assign f_arrdiv16_fs153_xor0 = f_arrdiv16_mux2to1128_xor0 ^ b[9];
  assign f_arrdiv16_fs153_not0 = ~f_arrdiv16_mux2to1128_xor0;
  assign f_arrdiv16_fs153_and0 = f_arrdiv16_fs153_not0 & b[9];
  assign f_arrdiv16_fs153_xor1 = f_arrdiv16_fs152_or0 ^ f_arrdiv16_fs153_xor0;
  assign f_arrdiv16_fs153_not1 = ~f_arrdiv16_fs153_xor0;
  assign f_arrdiv16_fs153_and1 = f_arrdiv16_fs153_not1 & f_arrdiv16_fs152_or0;
  assign f_arrdiv16_fs153_or0 = f_arrdiv16_fs153_and1 | f_arrdiv16_fs153_and0;
  assign f_arrdiv16_fs154_xor0 = f_arrdiv16_mux2to1129_xor0 ^ b[10];
  assign f_arrdiv16_fs154_not0 = ~f_arrdiv16_mux2to1129_xor0;
  assign f_arrdiv16_fs154_and0 = f_arrdiv16_fs154_not0 & b[10];
  assign f_arrdiv16_fs154_xor1 = f_arrdiv16_fs153_or0 ^ f_arrdiv16_fs154_xor0;
  assign f_arrdiv16_fs154_not1 = ~f_arrdiv16_fs154_xor0;
  assign f_arrdiv16_fs154_and1 = f_arrdiv16_fs154_not1 & f_arrdiv16_fs153_or0;
  assign f_arrdiv16_fs154_or0 = f_arrdiv16_fs154_and1 | f_arrdiv16_fs154_and0;
  assign f_arrdiv16_fs155_xor0 = f_arrdiv16_mux2to1130_xor0 ^ b[11];
  assign f_arrdiv16_fs155_not0 = ~f_arrdiv16_mux2to1130_xor0;
  assign f_arrdiv16_fs155_and0 = f_arrdiv16_fs155_not0 & b[11];
  assign f_arrdiv16_fs155_xor1 = f_arrdiv16_fs154_or0 ^ f_arrdiv16_fs155_xor0;
  assign f_arrdiv16_fs155_not1 = ~f_arrdiv16_fs155_xor0;
  assign f_arrdiv16_fs155_and1 = f_arrdiv16_fs155_not1 & f_arrdiv16_fs154_or0;
  assign f_arrdiv16_fs155_or0 = f_arrdiv16_fs155_and1 | f_arrdiv16_fs155_and0;
  assign f_arrdiv16_fs156_xor0 = f_arrdiv16_mux2to1131_xor0 ^ b[12];
  assign f_arrdiv16_fs156_not0 = ~f_arrdiv16_mux2to1131_xor0;
  assign f_arrdiv16_fs156_and0 = f_arrdiv16_fs156_not0 & b[12];
  assign f_arrdiv16_fs156_xor1 = f_arrdiv16_fs155_or0 ^ f_arrdiv16_fs156_xor0;
  assign f_arrdiv16_fs156_not1 = ~f_arrdiv16_fs156_xor0;
  assign f_arrdiv16_fs156_and1 = f_arrdiv16_fs156_not1 & f_arrdiv16_fs155_or0;
  assign f_arrdiv16_fs156_or0 = f_arrdiv16_fs156_and1 | f_arrdiv16_fs156_and0;
  assign f_arrdiv16_fs157_xor0 = f_arrdiv16_mux2to1132_xor0 ^ b[13];
  assign f_arrdiv16_fs157_not0 = ~f_arrdiv16_mux2to1132_xor0;
  assign f_arrdiv16_fs157_and0 = f_arrdiv16_fs157_not0 & b[13];
  assign f_arrdiv16_fs157_xor1 = f_arrdiv16_fs156_or0 ^ f_arrdiv16_fs157_xor0;
  assign f_arrdiv16_fs157_not1 = ~f_arrdiv16_fs157_xor0;
  assign f_arrdiv16_fs157_and1 = f_arrdiv16_fs157_not1 & f_arrdiv16_fs156_or0;
  assign f_arrdiv16_fs157_or0 = f_arrdiv16_fs157_and1 | f_arrdiv16_fs157_and0;
  assign f_arrdiv16_fs158_xor0 = f_arrdiv16_mux2to1133_xor0 ^ b[14];
  assign f_arrdiv16_fs158_not0 = ~f_arrdiv16_mux2to1133_xor0;
  assign f_arrdiv16_fs158_and0 = f_arrdiv16_fs158_not0 & b[14];
  assign f_arrdiv16_fs158_xor1 = f_arrdiv16_fs157_or0 ^ f_arrdiv16_fs158_xor0;
  assign f_arrdiv16_fs158_not1 = ~f_arrdiv16_fs158_xor0;
  assign f_arrdiv16_fs158_and1 = f_arrdiv16_fs158_not1 & f_arrdiv16_fs157_or0;
  assign f_arrdiv16_fs158_or0 = f_arrdiv16_fs158_and1 | f_arrdiv16_fs158_and0;
  assign f_arrdiv16_fs159_xor0 = f_arrdiv16_mux2to1134_xor0 ^ b[15];
  assign f_arrdiv16_fs159_not0 = ~f_arrdiv16_mux2to1134_xor0;
  assign f_arrdiv16_fs159_and0 = f_arrdiv16_fs159_not0 & b[15];
  assign f_arrdiv16_fs159_xor1 = f_arrdiv16_fs158_or0 ^ f_arrdiv16_fs159_xor0;
  assign f_arrdiv16_fs159_not1 = ~f_arrdiv16_fs159_xor0;
  assign f_arrdiv16_fs159_and1 = f_arrdiv16_fs159_not1 & f_arrdiv16_fs158_or0;
  assign f_arrdiv16_fs159_or0 = f_arrdiv16_fs159_and1 | f_arrdiv16_fs159_and0;
  assign f_arrdiv16_mux2to1135_and0 = a[6] & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1135_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1135_and1 = f_arrdiv16_fs144_xor0 & f_arrdiv16_mux2to1135_not0;
  assign f_arrdiv16_mux2to1135_xor0 = f_arrdiv16_mux2to1135_and0 ^ f_arrdiv16_mux2to1135_and1;
  assign f_arrdiv16_mux2to1136_and0 = f_arrdiv16_mux2to1120_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1136_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1136_and1 = f_arrdiv16_fs145_xor1 & f_arrdiv16_mux2to1136_not0;
  assign f_arrdiv16_mux2to1136_xor0 = f_arrdiv16_mux2to1136_and0 ^ f_arrdiv16_mux2to1136_and1;
  assign f_arrdiv16_mux2to1137_and0 = f_arrdiv16_mux2to1121_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1137_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1137_and1 = f_arrdiv16_fs146_xor1 & f_arrdiv16_mux2to1137_not0;
  assign f_arrdiv16_mux2to1137_xor0 = f_arrdiv16_mux2to1137_and0 ^ f_arrdiv16_mux2to1137_and1;
  assign f_arrdiv16_mux2to1138_and0 = f_arrdiv16_mux2to1122_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1138_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1138_and1 = f_arrdiv16_fs147_xor1 & f_arrdiv16_mux2to1138_not0;
  assign f_arrdiv16_mux2to1138_xor0 = f_arrdiv16_mux2to1138_and0 ^ f_arrdiv16_mux2to1138_and1;
  assign f_arrdiv16_mux2to1139_and0 = f_arrdiv16_mux2to1123_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1139_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1139_and1 = f_arrdiv16_fs148_xor1 & f_arrdiv16_mux2to1139_not0;
  assign f_arrdiv16_mux2to1139_xor0 = f_arrdiv16_mux2to1139_and0 ^ f_arrdiv16_mux2to1139_and1;
  assign f_arrdiv16_mux2to1140_and0 = f_arrdiv16_mux2to1124_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1140_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1140_and1 = f_arrdiv16_fs149_xor1 & f_arrdiv16_mux2to1140_not0;
  assign f_arrdiv16_mux2to1140_xor0 = f_arrdiv16_mux2to1140_and0 ^ f_arrdiv16_mux2to1140_and1;
  assign f_arrdiv16_mux2to1141_and0 = f_arrdiv16_mux2to1125_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1141_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1141_and1 = f_arrdiv16_fs150_xor1 & f_arrdiv16_mux2to1141_not0;
  assign f_arrdiv16_mux2to1141_xor0 = f_arrdiv16_mux2to1141_and0 ^ f_arrdiv16_mux2to1141_and1;
  assign f_arrdiv16_mux2to1142_and0 = f_arrdiv16_mux2to1126_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1142_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1142_and1 = f_arrdiv16_fs151_xor1 & f_arrdiv16_mux2to1142_not0;
  assign f_arrdiv16_mux2to1142_xor0 = f_arrdiv16_mux2to1142_and0 ^ f_arrdiv16_mux2to1142_and1;
  assign f_arrdiv16_mux2to1143_and0 = f_arrdiv16_mux2to1127_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1143_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1143_and1 = f_arrdiv16_fs152_xor1 & f_arrdiv16_mux2to1143_not0;
  assign f_arrdiv16_mux2to1143_xor0 = f_arrdiv16_mux2to1143_and0 ^ f_arrdiv16_mux2to1143_and1;
  assign f_arrdiv16_mux2to1144_and0 = f_arrdiv16_mux2to1128_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1144_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1144_and1 = f_arrdiv16_fs153_xor1 & f_arrdiv16_mux2to1144_not0;
  assign f_arrdiv16_mux2to1144_xor0 = f_arrdiv16_mux2to1144_and0 ^ f_arrdiv16_mux2to1144_and1;
  assign f_arrdiv16_mux2to1145_and0 = f_arrdiv16_mux2to1129_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1145_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1145_and1 = f_arrdiv16_fs154_xor1 & f_arrdiv16_mux2to1145_not0;
  assign f_arrdiv16_mux2to1145_xor0 = f_arrdiv16_mux2to1145_and0 ^ f_arrdiv16_mux2to1145_and1;
  assign f_arrdiv16_mux2to1146_and0 = f_arrdiv16_mux2to1130_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1146_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1146_and1 = f_arrdiv16_fs155_xor1 & f_arrdiv16_mux2to1146_not0;
  assign f_arrdiv16_mux2to1146_xor0 = f_arrdiv16_mux2to1146_and0 ^ f_arrdiv16_mux2to1146_and1;
  assign f_arrdiv16_mux2to1147_and0 = f_arrdiv16_mux2to1131_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1147_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1147_and1 = f_arrdiv16_fs156_xor1 & f_arrdiv16_mux2to1147_not0;
  assign f_arrdiv16_mux2to1147_xor0 = f_arrdiv16_mux2to1147_and0 ^ f_arrdiv16_mux2to1147_and1;
  assign f_arrdiv16_mux2to1148_and0 = f_arrdiv16_mux2to1132_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1148_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1148_and1 = f_arrdiv16_fs157_xor1 & f_arrdiv16_mux2to1148_not0;
  assign f_arrdiv16_mux2to1148_xor0 = f_arrdiv16_mux2to1148_and0 ^ f_arrdiv16_mux2to1148_and1;
  assign f_arrdiv16_mux2to1149_and0 = f_arrdiv16_mux2to1133_xor0 & f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1149_not0 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_mux2to1149_and1 = f_arrdiv16_fs158_xor1 & f_arrdiv16_mux2to1149_not0;
  assign f_arrdiv16_mux2to1149_xor0 = f_arrdiv16_mux2to1149_and0 ^ f_arrdiv16_mux2to1149_and1;
  assign f_arrdiv16_not9 = ~f_arrdiv16_fs159_or0;
  assign f_arrdiv16_fs160_xor0 = a[5] ^ b[0];
  assign f_arrdiv16_fs160_not0 = ~a[5];
  assign f_arrdiv16_fs160_and0 = f_arrdiv16_fs160_not0 & b[0];
  assign f_arrdiv16_fs160_not1 = ~f_arrdiv16_fs160_xor0;
  assign f_arrdiv16_fs161_xor0 = f_arrdiv16_mux2to1135_xor0 ^ b[1];
  assign f_arrdiv16_fs161_not0 = ~f_arrdiv16_mux2to1135_xor0;
  assign f_arrdiv16_fs161_and0 = f_arrdiv16_fs161_not0 & b[1];
  assign f_arrdiv16_fs161_xor1 = f_arrdiv16_fs160_and0 ^ f_arrdiv16_fs161_xor0;
  assign f_arrdiv16_fs161_not1 = ~f_arrdiv16_fs161_xor0;
  assign f_arrdiv16_fs161_and1 = f_arrdiv16_fs161_not1 & f_arrdiv16_fs160_and0;
  assign f_arrdiv16_fs161_or0 = f_arrdiv16_fs161_and1 | f_arrdiv16_fs161_and0;
  assign f_arrdiv16_fs162_xor0 = f_arrdiv16_mux2to1136_xor0 ^ b[2];
  assign f_arrdiv16_fs162_not0 = ~f_arrdiv16_mux2to1136_xor0;
  assign f_arrdiv16_fs162_and0 = f_arrdiv16_fs162_not0 & b[2];
  assign f_arrdiv16_fs162_xor1 = f_arrdiv16_fs161_or0 ^ f_arrdiv16_fs162_xor0;
  assign f_arrdiv16_fs162_not1 = ~f_arrdiv16_fs162_xor0;
  assign f_arrdiv16_fs162_and1 = f_arrdiv16_fs162_not1 & f_arrdiv16_fs161_or0;
  assign f_arrdiv16_fs162_or0 = f_arrdiv16_fs162_and1 | f_arrdiv16_fs162_and0;
  assign f_arrdiv16_fs163_xor0 = f_arrdiv16_mux2to1137_xor0 ^ b[3];
  assign f_arrdiv16_fs163_not0 = ~f_arrdiv16_mux2to1137_xor0;
  assign f_arrdiv16_fs163_and0 = f_arrdiv16_fs163_not0 & b[3];
  assign f_arrdiv16_fs163_xor1 = f_arrdiv16_fs162_or0 ^ f_arrdiv16_fs163_xor0;
  assign f_arrdiv16_fs163_not1 = ~f_arrdiv16_fs163_xor0;
  assign f_arrdiv16_fs163_and1 = f_arrdiv16_fs163_not1 & f_arrdiv16_fs162_or0;
  assign f_arrdiv16_fs163_or0 = f_arrdiv16_fs163_and1 | f_arrdiv16_fs163_and0;
  assign f_arrdiv16_fs164_xor0 = f_arrdiv16_mux2to1138_xor0 ^ b[4];
  assign f_arrdiv16_fs164_not0 = ~f_arrdiv16_mux2to1138_xor0;
  assign f_arrdiv16_fs164_and0 = f_arrdiv16_fs164_not0 & b[4];
  assign f_arrdiv16_fs164_xor1 = f_arrdiv16_fs163_or0 ^ f_arrdiv16_fs164_xor0;
  assign f_arrdiv16_fs164_not1 = ~f_arrdiv16_fs164_xor0;
  assign f_arrdiv16_fs164_and1 = f_arrdiv16_fs164_not1 & f_arrdiv16_fs163_or0;
  assign f_arrdiv16_fs164_or0 = f_arrdiv16_fs164_and1 | f_arrdiv16_fs164_and0;
  assign f_arrdiv16_fs165_xor0 = f_arrdiv16_mux2to1139_xor0 ^ b[5];
  assign f_arrdiv16_fs165_not0 = ~f_arrdiv16_mux2to1139_xor0;
  assign f_arrdiv16_fs165_and0 = f_arrdiv16_fs165_not0 & b[5];
  assign f_arrdiv16_fs165_xor1 = f_arrdiv16_fs164_or0 ^ f_arrdiv16_fs165_xor0;
  assign f_arrdiv16_fs165_not1 = ~f_arrdiv16_fs165_xor0;
  assign f_arrdiv16_fs165_and1 = f_arrdiv16_fs165_not1 & f_arrdiv16_fs164_or0;
  assign f_arrdiv16_fs165_or0 = f_arrdiv16_fs165_and1 | f_arrdiv16_fs165_and0;
  assign f_arrdiv16_fs166_xor0 = f_arrdiv16_mux2to1140_xor0 ^ b[6];
  assign f_arrdiv16_fs166_not0 = ~f_arrdiv16_mux2to1140_xor0;
  assign f_arrdiv16_fs166_and0 = f_arrdiv16_fs166_not0 & b[6];
  assign f_arrdiv16_fs166_xor1 = f_arrdiv16_fs165_or0 ^ f_arrdiv16_fs166_xor0;
  assign f_arrdiv16_fs166_not1 = ~f_arrdiv16_fs166_xor0;
  assign f_arrdiv16_fs166_and1 = f_arrdiv16_fs166_not1 & f_arrdiv16_fs165_or0;
  assign f_arrdiv16_fs166_or0 = f_arrdiv16_fs166_and1 | f_arrdiv16_fs166_and0;
  assign f_arrdiv16_fs167_xor0 = f_arrdiv16_mux2to1141_xor0 ^ b[7];
  assign f_arrdiv16_fs167_not0 = ~f_arrdiv16_mux2to1141_xor0;
  assign f_arrdiv16_fs167_and0 = f_arrdiv16_fs167_not0 & b[7];
  assign f_arrdiv16_fs167_xor1 = f_arrdiv16_fs166_or0 ^ f_arrdiv16_fs167_xor0;
  assign f_arrdiv16_fs167_not1 = ~f_arrdiv16_fs167_xor0;
  assign f_arrdiv16_fs167_and1 = f_arrdiv16_fs167_not1 & f_arrdiv16_fs166_or0;
  assign f_arrdiv16_fs167_or0 = f_arrdiv16_fs167_and1 | f_arrdiv16_fs167_and0;
  assign f_arrdiv16_fs168_xor0 = f_arrdiv16_mux2to1142_xor0 ^ b[8];
  assign f_arrdiv16_fs168_not0 = ~f_arrdiv16_mux2to1142_xor0;
  assign f_arrdiv16_fs168_and0 = f_arrdiv16_fs168_not0 & b[8];
  assign f_arrdiv16_fs168_xor1 = f_arrdiv16_fs167_or0 ^ f_arrdiv16_fs168_xor0;
  assign f_arrdiv16_fs168_not1 = ~f_arrdiv16_fs168_xor0;
  assign f_arrdiv16_fs168_and1 = f_arrdiv16_fs168_not1 & f_arrdiv16_fs167_or0;
  assign f_arrdiv16_fs168_or0 = f_arrdiv16_fs168_and1 | f_arrdiv16_fs168_and0;
  assign f_arrdiv16_fs169_xor0 = f_arrdiv16_mux2to1143_xor0 ^ b[9];
  assign f_arrdiv16_fs169_not0 = ~f_arrdiv16_mux2to1143_xor0;
  assign f_arrdiv16_fs169_and0 = f_arrdiv16_fs169_not0 & b[9];
  assign f_arrdiv16_fs169_xor1 = f_arrdiv16_fs168_or0 ^ f_arrdiv16_fs169_xor0;
  assign f_arrdiv16_fs169_not1 = ~f_arrdiv16_fs169_xor0;
  assign f_arrdiv16_fs169_and1 = f_arrdiv16_fs169_not1 & f_arrdiv16_fs168_or0;
  assign f_arrdiv16_fs169_or0 = f_arrdiv16_fs169_and1 | f_arrdiv16_fs169_and0;
  assign f_arrdiv16_fs170_xor0 = f_arrdiv16_mux2to1144_xor0 ^ b[10];
  assign f_arrdiv16_fs170_not0 = ~f_arrdiv16_mux2to1144_xor0;
  assign f_arrdiv16_fs170_and0 = f_arrdiv16_fs170_not0 & b[10];
  assign f_arrdiv16_fs170_xor1 = f_arrdiv16_fs169_or0 ^ f_arrdiv16_fs170_xor0;
  assign f_arrdiv16_fs170_not1 = ~f_arrdiv16_fs170_xor0;
  assign f_arrdiv16_fs170_and1 = f_arrdiv16_fs170_not1 & f_arrdiv16_fs169_or0;
  assign f_arrdiv16_fs170_or0 = f_arrdiv16_fs170_and1 | f_arrdiv16_fs170_and0;
  assign f_arrdiv16_fs171_xor0 = f_arrdiv16_mux2to1145_xor0 ^ b[11];
  assign f_arrdiv16_fs171_not0 = ~f_arrdiv16_mux2to1145_xor0;
  assign f_arrdiv16_fs171_and0 = f_arrdiv16_fs171_not0 & b[11];
  assign f_arrdiv16_fs171_xor1 = f_arrdiv16_fs170_or0 ^ f_arrdiv16_fs171_xor0;
  assign f_arrdiv16_fs171_not1 = ~f_arrdiv16_fs171_xor0;
  assign f_arrdiv16_fs171_and1 = f_arrdiv16_fs171_not1 & f_arrdiv16_fs170_or0;
  assign f_arrdiv16_fs171_or0 = f_arrdiv16_fs171_and1 | f_arrdiv16_fs171_and0;
  assign f_arrdiv16_fs172_xor0 = f_arrdiv16_mux2to1146_xor0 ^ b[12];
  assign f_arrdiv16_fs172_not0 = ~f_arrdiv16_mux2to1146_xor0;
  assign f_arrdiv16_fs172_and0 = f_arrdiv16_fs172_not0 & b[12];
  assign f_arrdiv16_fs172_xor1 = f_arrdiv16_fs171_or0 ^ f_arrdiv16_fs172_xor0;
  assign f_arrdiv16_fs172_not1 = ~f_arrdiv16_fs172_xor0;
  assign f_arrdiv16_fs172_and1 = f_arrdiv16_fs172_not1 & f_arrdiv16_fs171_or0;
  assign f_arrdiv16_fs172_or0 = f_arrdiv16_fs172_and1 | f_arrdiv16_fs172_and0;
  assign f_arrdiv16_fs173_xor0 = f_arrdiv16_mux2to1147_xor0 ^ b[13];
  assign f_arrdiv16_fs173_not0 = ~f_arrdiv16_mux2to1147_xor0;
  assign f_arrdiv16_fs173_and0 = f_arrdiv16_fs173_not0 & b[13];
  assign f_arrdiv16_fs173_xor1 = f_arrdiv16_fs172_or0 ^ f_arrdiv16_fs173_xor0;
  assign f_arrdiv16_fs173_not1 = ~f_arrdiv16_fs173_xor0;
  assign f_arrdiv16_fs173_and1 = f_arrdiv16_fs173_not1 & f_arrdiv16_fs172_or0;
  assign f_arrdiv16_fs173_or0 = f_arrdiv16_fs173_and1 | f_arrdiv16_fs173_and0;
  assign f_arrdiv16_fs174_xor0 = f_arrdiv16_mux2to1148_xor0 ^ b[14];
  assign f_arrdiv16_fs174_not0 = ~f_arrdiv16_mux2to1148_xor0;
  assign f_arrdiv16_fs174_and0 = f_arrdiv16_fs174_not0 & b[14];
  assign f_arrdiv16_fs174_xor1 = f_arrdiv16_fs173_or0 ^ f_arrdiv16_fs174_xor0;
  assign f_arrdiv16_fs174_not1 = ~f_arrdiv16_fs174_xor0;
  assign f_arrdiv16_fs174_and1 = f_arrdiv16_fs174_not1 & f_arrdiv16_fs173_or0;
  assign f_arrdiv16_fs174_or0 = f_arrdiv16_fs174_and1 | f_arrdiv16_fs174_and0;
  assign f_arrdiv16_fs175_xor0 = f_arrdiv16_mux2to1149_xor0 ^ b[15];
  assign f_arrdiv16_fs175_not0 = ~f_arrdiv16_mux2to1149_xor0;
  assign f_arrdiv16_fs175_and0 = f_arrdiv16_fs175_not0 & b[15];
  assign f_arrdiv16_fs175_xor1 = f_arrdiv16_fs174_or0 ^ f_arrdiv16_fs175_xor0;
  assign f_arrdiv16_fs175_not1 = ~f_arrdiv16_fs175_xor0;
  assign f_arrdiv16_fs175_and1 = f_arrdiv16_fs175_not1 & f_arrdiv16_fs174_or0;
  assign f_arrdiv16_fs175_or0 = f_arrdiv16_fs175_and1 | f_arrdiv16_fs175_and0;
  assign f_arrdiv16_mux2to1150_and0 = a[5] & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1150_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1150_and1 = f_arrdiv16_fs160_xor0 & f_arrdiv16_mux2to1150_not0;
  assign f_arrdiv16_mux2to1150_xor0 = f_arrdiv16_mux2to1150_and0 ^ f_arrdiv16_mux2to1150_and1;
  assign f_arrdiv16_mux2to1151_and0 = f_arrdiv16_mux2to1135_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1151_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1151_and1 = f_arrdiv16_fs161_xor1 & f_arrdiv16_mux2to1151_not0;
  assign f_arrdiv16_mux2to1151_xor0 = f_arrdiv16_mux2to1151_and0 ^ f_arrdiv16_mux2to1151_and1;
  assign f_arrdiv16_mux2to1152_and0 = f_arrdiv16_mux2to1136_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1152_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1152_and1 = f_arrdiv16_fs162_xor1 & f_arrdiv16_mux2to1152_not0;
  assign f_arrdiv16_mux2to1152_xor0 = f_arrdiv16_mux2to1152_and0 ^ f_arrdiv16_mux2to1152_and1;
  assign f_arrdiv16_mux2to1153_and0 = f_arrdiv16_mux2to1137_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1153_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1153_and1 = f_arrdiv16_fs163_xor1 & f_arrdiv16_mux2to1153_not0;
  assign f_arrdiv16_mux2to1153_xor0 = f_arrdiv16_mux2to1153_and0 ^ f_arrdiv16_mux2to1153_and1;
  assign f_arrdiv16_mux2to1154_and0 = f_arrdiv16_mux2to1138_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1154_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1154_and1 = f_arrdiv16_fs164_xor1 & f_arrdiv16_mux2to1154_not0;
  assign f_arrdiv16_mux2to1154_xor0 = f_arrdiv16_mux2to1154_and0 ^ f_arrdiv16_mux2to1154_and1;
  assign f_arrdiv16_mux2to1155_and0 = f_arrdiv16_mux2to1139_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1155_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1155_and1 = f_arrdiv16_fs165_xor1 & f_arrdiv16_mux2to1155_not0;
  assign f_arrdiv16_mux2to1155_xor0 = f_arrdiv16_mux2to1155_and0 ^ f_arrdiv16_mux2to1155_and1;
  assign f_arrdiv16_mux2to1156_and0 = f_arrdiv16_mux2to1140_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1156_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1156_and1 = f_arrdiv16_fs166_xor1 & f_arrdiv16_mux2to1156_not0;
  assign f_arrdiv16_mux2to1156_xor0 = f_arrdiv16_mux2to1156_and0 ^ f_arrdiv16_mux2to1156_and1;
  assign f_arrdiv16_mux2to1157_and0 = f_arrdiv16_mux2to1141_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1157_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1157_and1 = f_arrdiv16_fs167_xor1 & f_arrdiv16_mux2to1157_not0;
  assign f_arrdiv16_mux2to1157_xor0 = f_arrdiv16_mux2to1157_and0 ^ f_arrdiv16_mux2to1157_and1;
  assign f_arrdiv16_mux2to1158_and0 = f_arrdiv16_mux2to1142_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1158_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1158_and1 = f_arrdiv16_fs168_xor1 & f_arrdiv16_mux2to1158_not0;
  assign f_arrdiv16_mux2to1158_xor0 = f_arrdiv16_mux2to1158_and0 ^ f_arrdiv16_mux2to1158_and1;
  assign f_arrdiv16_mux2to1159_and0 = f_arrdiv16_mux2to1143_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1159_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1159_and1 = f_arrdiv16_fs169_xor1 & f_arrdiv16_mux2to1159_not0;
  assign f_arrdiv16_mux2to1159_xor0 = f_arrdiv16_mux2to1159_and0 ^ f_arrdiv16_mux2to1159_and1;
  assign f_arrdiv16_mux2to1160_and0 = f_arrdiv16_mux2to1144_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1160_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1160_and1 = f_arrdiv16_fs170_xor1 & f_arrdiv16_mux2to1160_not0;
  assign f_arrdiv16_mux2to1160_xor0 = f_arrdiv16_mux2to1160_and0 ^ f_arrdiv16_mux2to1160_and1;
  assign f_arrdiv16_mux2to1161_and0 = f_arrdiv16_mux2to1145_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1161_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1161_and1 = f_arrdiv16_fs171_xor1 & f_arrdiv16_mux2to1161_not0;
  assign f_arrdiv16_mux2to1161_xor0 = f_arrdiv16_mux2to1161_and0 ^ f_arrdiv16_mux2to1161_and1;
  assign f_arrdiv16_mux2to1162_and0 = f_arrdiv16_mux2to1146_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1162_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1162_and1 = f_arrdiv16_fs172_xor1 & f_arrdiv16_mux2to1162_not0;
  assign f_arrdiv16_mux2to1162_xor0 = f_arrdiv16_mux2to1162_and0 ^ f_arrdiv16_mux2to1162_and1;
  assign f_arrdiv16_mux2to1163_and0 = f_arrdiv16_mux2to1147_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1163_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1163_and1 = f_arrdiv16_fs173_xor1 & f_arrdiv16_mux2to1163_not0;
  assign f_arrdiv16_mux2to1163_xor0 = f_arrdiv16_mux2to1163_and0 ^ f_arrdiv16_mux2to1163_and1;
  assign f_arrdiv16_mux2to1164_and0 = f_arrdiv16_mux2to1148_xor0 & f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1164_not0 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_mux2to1164_and1 = f_arrdiv16_fs174_xor1 & f_arrdiv16_mux2to1164_not0;
  assign f_arrdiv16_mux2to1164_xor0 = f_arrdiv16_mux2to1164_and0 ^ f_arrdiv16_mux2to1164_and1;
  assign f_arrdiv16_not10 = ~f_arrdiv16_fs175_or0;
  assign f_arrdiv16_fs176_xor0 = a[4] ^ b[0];
  assign f_arrdiv16_fs176_not0 = ~a[4];
  assign f_arrdiv16_fs176_and0 = f_arrdiv16_fs176_not0 & b[0];
  assign f_arrdiv16_fs176_not1 = ~f_arrdiv16_fs176_xor0;
  assign f_arrdiv16_fs177_xor0 = f_arrdiv16_mux2to1150_xor0 ^ b[1];
  assign f_arrdiv16_fs177_not0 = ~f_arrdiv16_mux2to1150_xor0;
  assign f_arrdiv16_fs177_and0 = f_arrdiv16_fs177_not0 & b[1];
  assign f_arrdiv16_fs177_xor1 = f_arrdiv16_fs176_and0 ^ f_arrdiv16_fs177_xor0;
  assign f_arrdiv16_fs177_not1 = ~f_arrdiv16_fs177_xor0;
  assign f_arrdiv16_fs177_and1 = f_arrdiv16_fs177_not1 & f_arrdiv16_fs176_and0;
  assign f_arrdiv16_fs177_or0 = f_arrdiv16_fs177_and1 | f_arrdiv16_fs177_and0;
  assign f_arrdiv16_fs178_xor0 = f_arrdiv16_mux2to1151_xor0 ^ b[2];
  assign f_arrdiv16_fs178_not0 = ~f_arrdiv16_mux2to1151_xor0;
  assign f_arrdiv16_fs178_and0 = f_arrdiv16_fs178_not0 & b[2];
  assign f_arrdiv16_fs178_xor1 = f_arrdiv16_fs177_or0 ^ f_arrdiv16_fs178_xor0;
  assign f_arrdiv16_fs178_not1 = ~f_arrdiv16_fs178_xor0;
  assign f_arrdiv16_fs178_and1 = f_arrdiv16_fs178_not1 & f_arrdiv16_fs177_or0;
  assign f_arrdiv16_fs178_or0 = f_arrdiv16_fs178_and1 | f_arrdiv16_fs178_and0;
  assign f_arrdiv16_fs179_xor0 = f_arrdiv16_mux2to1152_xor0 ^ b[3];
  assign f_arrdiv16_fs179_not0 = ~f_arrdiv16_mux2to1152_xor0;
  assign f_arrdiv16_fs179_and0 = f_arrdiv16_fs179_not0 & b[3];
  assign f_arrdiv16_fs179_xor1 = f_arrdiv16_fs178_or0 ^ f_arrdiv16_fs179_xor0;
  assign f_arrdiv16_fs179_not1 = ~f_arrdiv16_fs179_xor0;
  assign f_arrdiv16_fs179_and1 = f_arrdiv16_fs179_not1 & f_arrdiv16_fs178_or0;
  assign f_arrdiv16_fs179_or0 = f_arrdiv16_fs179_and1 | f_arrdiv16_fs179_and0;
  assign f_arrdiv16_fs180_xor0 = f_arrdiv16_mux2to1153_xor0 ^ b[4];
  assign f_arrdiv16_fs180_not0 = ~f_arrdiv16_mux2to1153_xor0;
  assign f_arrdiv16_fs180_and0 = f_arrdiv16_fs180_not0 & b[4];
  assign f_arrdiv16_fs180_xor1 = f_arrdiv16_fs179_or0 ^ f_arrdiv16_fs180_xor0;
  assign f_arrdiv16_fs180_not1 = ~f_arrdiv16_fs180_xor0;
  assign f_arrdiv16_fs180_and1 = f_arrdiv16_fs180_not1 & f_arrdiv16_fs179_or0;
  assign f_arrdiv16_fs180_or0 = f_arrdiv16_fs180_and1 | f_arrdiv16_fs180_and0;
  assign f_arrdiv16_fs181_xor0 = f_arrdiv16_mux2to1154_xor0 ^ b[5];
  assign f_arrdiv16_fs181_not0 = ~f_arrdiv16_mux2to1154_xor0;
  assign f_arrdiv16_fs181_and0 = f_arrdiv16_fs181_not0 & b[5];
  assign f_arrdiv16_fs181_xor1 = f_arrdiv16_fs180_or0 ^ f_arrdiv16_fs181_xor0;
  assign f_arrdiv16_fs181_not1 = ~f_arrdiv16_fs181_xor0;
  assign f_arrdiv16_fs181_and1 = f_arrdiv16_fs181_not1 & f_arrdiv16_fs180_or0;
  assign f_arrdiv16_fs181_or0 = f_arrdiv16_fs181_and1 | f_arrdiv16_fs181_and0;
  assign f_arrdiv16_fs182_xor0 = f_arrdiv16_mux2to1155_xor0 ^ b[6];
  assign f_arrdiv16_fs182_not0 = ~f_arrdiv16_mux2to1155_xor0;
  assign f_arrdiv16_fs182_and0 = f_arrdiv16_fs182_not0 & b[6];
  assign f_arrdiv16_fs182_xor1 = f_arrdiv16_fs181_or0 ^ f_arrdiv16_fs182_xor0;
  assign f_arrdiv16_fs182_not1 = ~f_arrdiv16_fs182_xor0;
  assign f_arrdiv16_fs182_and1 = f_arrdiv16_fs182_not1 & f_arrdiv16_fs181_or0;
  assign f_arrdiv16_fs182_or0 = f_arrdiv16_fs182_and1 | f_arrdiv16_fs182_and0;
  assign f_arrdiv16_fs183_xor0 = f_arrdiv16_mux2to1156_xor0 ^ b[7];
  assign f_arrdiv16_fs183_not0 = ~f_arrdiv16_mux2to1156_xor0;
  assign f_arrdiv16_fs183_and0 = f_arrdiv16_fs183_not0 & b[7];
  assign f_arrdiv16_fs183_xor1 = f_arrdiv16_fs182_or0 ^ f_arrdiv16_fs183_xor0;
  assign f_arrdiv16_fs183_not1 = ~f_arrdiv16_fs183_xor0;
  assign f_arrdiv16_fs183_and1 = f_arrdiv16_fs183_not1 & f_arrdiv16_fs182_or0;
  assign f_arrdiv16_fs183_or0 = f_arrdiv16_fs183_and1 | f_arrdiv16_fs183_and0;
  assign f_arrdiv16_fs184_xor0 = f_arrdiv16_mux2to1157_xor0 ^ b[8];
  assign f_arrdiv16_fs184_not0 = ~f_arrdiv16_mux2to1157_xor0;
  assign f_arrdiv16_fs184_and0 = f_arrdiv16_fs184_not0 & b[8];
  assign f_arrdiv16_fs184_xor1 = f_arrdiv16_fs183_or0 ^ f_arrdiv16_fs184_xor0;
  assign f_arrdiv16_fs184_not1 = ~f_arrdiv16_fs184_xor0;
  assign f_arrdiv16_fs184_and1 = f_arrdiv16_fs184_not1 & f_arrdiv16_fs183_or0;
  assign f_arrdiv16_fs184_or0 = f_arrdiv16_fs184_and1 | f_arrdiv16_fs184_and0;
  assign f_arrdiv16_fs185_xor0 = f_arrdiv16_mux2to1158_xor0 ^ b[9];
  assign f_arrdiv16_fs185_not0 = ~f_arrdiv16_mux2to1158_xor0;
  assign f_arrdiv16_fs185_and0 = f_arrdiv16_fs185_not0 & b[9];
  assign f_arrdiv16_fs185_xor1 = f_arrdiv16_fs184_or0 ^ f_arrdiv16_fs185_xor0;
  assign f_arrdiv16_fs185_not1 = ~f_arrdiv16_fs185_xor0;
  assign f_arrdiv16_fs185_and1 = f_arrdiv16_fs185_not1 & f_arrdiv16_fs184_or0;
  assign f_arrdiv16_fs185_or0 = f_arrdiv16_fs185_and1 | f_arrdiv16_fs185_and0;
  assign f_arrdiv16_fs186_xor0 = f_arrdiv16_mux2to1159_xor0 ^ b[10];
  assign f_arrdiv16_fs186_not0 = ~f_arrdiv16_mux2to1159_xor0;
  assign f_arrdiv16_fs186_and0 = f_arrdiv16_fs186_not0 & b[10];
  assign f_arrdiv16_fs186_xor1 = f_arrdiv16_fs185_or0 ^ f_arrdiv16_fs186_xor0;
  assign f_arrdiv16_fs186_not1 = ~f_arrdiv16_fs186_xor0;
  assign f_arrdiv16_fs186_and1 = f_arrdiv16_fs186_not1 & f_arrdiv16_fs185_or0;
  assign f_arrdiv16_fs186_or0 = f_arrdiv16_fs186_and1 | f_arrdiv16_fs186_and0;
  assign f_arrdiv16_fs187_xor0 = f_arrdiv16_mux2to1160_xor0 ^ b[11];
  assign f_arrdiv16_fs187_not0 = ~f_arrdiv16_mux2to1160_xor0;
  assign f_arrdiv16_fs187_and0 = f_arrdiv16_fs187_not0 & b[11];
  assign f_arrdiv16_fs187_xor1 = f_arrdiv16_fs186_or0 ^ f_arrdiv16_fs187_xor0;
  assign f_arrdiv16_fs187_not1 = ~f_arrdiv16_fs187_xor0;
  assign f_arrdiv16_fs187_and1 = f_arrdiv16_fs187_not1 & f_arrdiv16_fs186_or0;
  assign f_arrdiv16_fs187_or0 = f_arrdiv16_fs187_and1 | f_arrdiv16_fs187_and0;
  assign f_arrdiv16_fs188_xor0 = f_arrdiv16_mux2to1161_xor0 ^ b[12];
  assign f_arrdiv16_fs188_not0 = ~f_arrdiv16_mux2to1161_xor0;
  assign f_arrdiv16_fs188_and0 = f_arrdiv16_fs188_not0 & b[12];
  assign f_arrdiv16_fs188_xor1 = f_arrdiv16_fs187_or0 ^ f_arrdiv16_fs188_xor0;
  assign f_arrdiv16_fs188_not1 = ~f_arrdiv16_fs188_xor0;
  assign f_arrdiv16_fs188_and1 = f_arrdiv16_fs188_not1 & f_arrdiv16_fs187_or0;
  assign f_arrdiv16_fs188_or0 = f_arrdiv16_fs188_and1 | f_arrdiv16_fs188_and0;
  assign f_arrdiv16_fs189_xor0 = f_arrdiv16_mux2to1162_xor0 ^ b[13];
  assign f_arrdiv16_fs189_not0 = ~f_arrdiv16_mux2to1162_xor0;
  assign f_arrdiv16_fs189_and0 = f_arrdiv16_fs189_not0 & b[13];
  assign f_arrdiv16_fs189_xor1 = f_arrdiv16_fs188_or0 ^ f_arrdiv16_fs189_xor0;
  assign f_arrdiv16_fs189_not1 = ~f_arrdiv16_fs189_xor0;
  assign f_arrdiv16_fs189_and1 = f_arrdiv16_fs189_not1 & f_arrdiv16_fs188_or0;
  assign f_arrdiv16_fs189_or0 = f_arrdiv16_fs189_and1 | f_arrdiv16_fs189_and0;
  assign f_arrdiv16_fs190_xor0 = f_arrdiv16_mux2to1163_xor0 ^ b[14];
  assign f_arrdiv16_fs190_not0 = ~f_arrdiv16_mux2to1163_xor0;
  assign f_arrdiv16_fs190_and0 = f_arrdiv16_fs190_not0 & b[14];
  assign f_arrdiv16_fs190_xor1 = f_arrdiv16_fs189_or0 ^ f_arrdiv16_fs190_xor0;
  assign f_arrdiv16_fs190_not1 = ~f_arrdiv16_fs190_xor0;
  assign f_arrdiv16_fs190_and1 = f_arrdiv16_fs190_not1 & f_arrdiv16_fs189_or0;
  assign f_arrdiv16_fs190_or0 = f_arrdiv16_fs190_and1 | f_arrdiv16_fs190_and0;
  assign f_arrdiv16_fs191_xor0 = f_arrdiv16_mux2to1164_xor0 ^ b[15];
  assign f_arrdiv16_fs191_not0 = ~f_arrdiv16_mux2to1164_xor0;
  assign f_arrdiv16_fs191_and0 = f_arrdiv16_fs191_not0 & b[15];
  assign f_arrdiv16_fs191_xor1 = f_arrdiv16_fs190_or0 ^ f_arrdiv16_fs191_xor0;
  assign f_arrdiv16_fs191_not1 = ~f_arrdiv16_fs191_xor0;
  assign f_arrdiv16_fs191_and1 = f_arrdiv16_fs191_not1 & f_arrdiv16_fs190_or0;
  assign f_arrdiv16_fs191_or0 = f_arrdiv16_fs191_and1 | f_arrdiv16_fs191_and0;
  assign f_arrdiv16_mux2to1165_and0 = a[4] & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1165_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1165_and1 = f_arrdiv16_fs176_xor0 & f_arrdiv16_mux2to1165_not0;
  assign f_arrdiv16_mux2to1165_xor0 = f_arrdiv16_mux2to1165_and0 ^ f_arrdiv16_mux2to1165_and1;
  assign f_arrdiv16_mux2to1166_and0 = f_arrdiv16_mux2to1150_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1166_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1166_and1 = f_arrdiv16_fs177_xor1 & f_arrdiv16_mux2to1166_not0;
  assign f_arrdiv16_mux2to1166_xor0 = f_arrdiv16_mux2to1166_and0 ^ f_arrdiv16_mux2to1166_and1;
  assign f_arrdiv16_mux2to1167_and0 = f_arrdiv16_mux2to1151_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1167_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1167_and1 = f_arrdiv16_fs178_xor1 & f_arrdiv16_mux2to1167_not0;
  assign f_arrdiv16_mux2to1167_xor0 = f_arrdiv16_mux2to1167_and0 ^ f_arrdiv16_mux2to1167_and1;
  assign f_arrdiv16_mux2to1168_and0 = f_arrdiv16_mux2to1152_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1168_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1168_and1 = f_arrdiv16_fs179_xor1 & f_arrdiv16_mux2to1168_not0;
  assign f_arrdiv16_mux2to1168_xor0 = f_arrdiv16_mux2to1168_and0 ^ f_arrdiv16_mux2to1168_and1;
  assign f_arrdiv16_mux2to1169_and0 = f_arrdiv16_mux2to1153_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1169_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1169_and1 = f_arrdiv16_fs180_xor1 & f_arrdiv16_mux2to1169_not0;
  assign f_arrdiv16_mux2to1169_xor0 = f_arrdiv16_mux2to1169_and0 ^ f_arrdiv16_mux2to1169_and1;
  assign f_arrdiv16_mux2to1170_and0 = f_arrdiv16_mux2to1154_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1170_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1170_and1 = f_arrdiv16_fs181_xor1 & f_arrdiv16_mux2to1170_not0;
  assign f_arrdiv16_mux2to1170_xor0 = f_arrdiv16_mux2to1170_and0 ^ f_arrdiv16_mux2to1170_and1;
  assign f_arrdiv16_mux2to1171_and0 = f_arrdiv16_mux2to1155_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1171_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1171_and1 = f_arrdiv16_fs182_xor1 & f_arrdiv16_mux2to1171_not0;
  assign f_arrdiv16_mux2to1171_xor0 = f_arrdiv16_mux2to1171_and0 ^ f_arrdiv16_mux2to1171_and1;
  assign f_arrdiv16_mux2to1172_and0 = f_arrdiv16_mux2to1156_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1172_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1172_and1 = f_arrdiv16_fs183_xor1 & f_arrdiv16_mux2to1172_not0;
  assign f_arrdiv16_mux2to1172_xor0 = f_arrdiv16_mux2to1172_and0 ^ f_arrdiv16_mux2to1172_and1;
  assign f_arrdiv16_mux2to1173_and0 = f_arrdiv16_mux2to1157_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1173_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1173_and1 = f_arrdiv16_fs184_xor1 & f_arrdiv16_mux2to1173_not0;
  assign f_arrdiv16_mux2to1173_xor0 = f_arrdiv16_mux2to1173_and0 ^ f_arrdiv16_mux2to1173_and1;
  assign f_arrdiv16_mux2to1174_and0 = f_arrdiv16_mux2to1158_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1174_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1174_and1 = f_arrdiv16_fs185_xor1 & f_arrdiv16_mux2to1174_not0;
  assign f_arrdiv16_mux2to1174_xor0 = f_arrdiv16_mux2to1174_and0 ^ f_arrdiv16_mux2to1174_and1;
  assign f_arrdiv16_mux2to1175_and0 = f_arrdiv16_mux2to1159_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1175_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1175_and1 = f_arrdiv16_fs186_xor1 & f_arrdiv16_mux2to1175_not0;
  assign f_arrdiv16_mux2to1175_xor0 = f_arrdiv16_mux2to1175_and0 ^ f_arrdiv16_mux2to1175_and1;
  assign f_arrdiv16_mux2to1176_and0 = f_arrdiv16_mux2to1160_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1176_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1176_and1 = f_arrdiv16_fs187_xor1 & f_arrdiv16_mux2to1176_not0;
  assign f_arrdiv16_mux2to1176_xor0 = f_arrdiv16_mux2to1176_and0 ^ f_arrdiv16_mux2to1176_and1;
  assign f_arrdiv16_mux2to1177_and0 = f_arrdiv16_mux2to1161_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1177_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1177_and1 = f_arrdiv16_fs188_xor1 & f_arrdiv16_mux2to1177_not0;
  assign f_arrdiv16_mux2to1177_xor0 = f_arrdiv16_mux2to1177_and0 ^ f_arrdiv16_mux2to1177_and1;
  assign f_arrdiv16_mux2to1178_and0 = f_arrdiv16_mux2to1162_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1178_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1178_and1 = f_arrdiv16_fs189_xor1 & f_arrdiv16_mux2to1178_not0;
  assign f_arrdiv16_mux2to1178_xor0 = f_arrdiv16_mux2to1178_and0 ^ f_arrdiv16_mux2to1178_and1;
  assign f_arrdiv16_mux2to1179_and0 = f_arrdiv16_mux2to1163_xor0 & f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1179_not0 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_mux2to1179_and1 = f_arrdiv16_fs190_xor1 & f_arrdiv16_mux2to1179_not0;
  assign f_arrdiv16_mux2to1179_xor0 = f_arrdiv16_mux2to1179_and0 ^ f_arrdiv16_mux2to1179_and1;
  assign f_arrdiv16_not11 = ~f_arrdiv16_fs191_or0;
  assign f_arrdiv16_fs192_xor0 = a[3] ^ b[0];
  assign f_arrdiv16_fs192_not0 = ~a[3];
  assign f_arrdiv16_fs192_and0 = f_arrdiv16_fs192_not0 & b[0];
  assign f_arrdiv16_fs192_not1 = ~f_arrdiv16_fs192_xor0;
  assign f_arrdiv16_fs193_xor0 = f_arrdiv16_mux2to1165_xor0 ^ b[1];
  assign f_arrdiv16_fs193_not0 = ~f_arrdiv16_mux2to1165_xor0;
  assign f_arrdiv16_fs193_and0 = f_arrdiv16_fs193_not0 & b[1];
  assign f_arrdiv16_fs193_xor1 = f_arrdiv16_fs192_and0 ^ f_arrdiv16_fs193_xor0;
  assign f_arrdiv16_fs193_not1 = ~f_arrdiv16_fs193_xor0;
  assign f_arrdiv16_fs193_and1 = f_arrdiv16_fs193_not1 & f_arrdiv16_fs192_and0;
  assign f_arrdiv16_fs193_or0 = f_arrdiv16_fs193_and1 | f_arrdiv16_fs193_and0;
  assign f_arrdiv16_fs194_xor0 = f_arrdiv16_mux2to1166_xor0 ^ b[2];
  assign f_arrdiv16_fs194_not0 = ~f_arrdiv16_mux2to1166_xor0;
  assign f_arrdiv16_fs194_and0 = f_arrdiv16_fs194_not0 & b[2];
  assign f_arrdiv16_fs194_xor1 = f_arrdiv16_fs193_or0 ^ f_arrdiv16_fs194_xor0;
  assign f_arrdiv16_fs194_not1 = ~f_arrdiv16_fs194_xor0;
  assign f_arrdiv16_fs194_and1 = f_arrdiv16_fs194_not1 & f_arrdiv16_fs193_or0;
  assign f_arrdiv16_fs194_or0 = f_arrdiv16_fs194_and1 | f_arrdiv16_fs194_and0;
  assign f_arrdiv16_fs195_xor0 = f_arrdiv16_mux2to1167_xor0 ^ b[3];
  assign f_arrdiv16_fs195_not0 = ~f_arrdiv16_mux2to1167_xor0;
  assign f_arrdiv16_fs195_and0 = f_arrdiv16_fs195_not0 & b[3];
  assign f_arrdiv16_fs195_xor1 = f_arrdiv16_fs194_or0 ^ f_arrdiv16_fs195_xor0;
  assign f_arrdiv16_fs195_not1 = ~f_arrdiv16_fs195_xor0;
  assign f_arrdiv16_fs195_and1 = f_arrdiv16_fs195_not1 & f_arrdiv16_fs194_or0;
  assign f_arrdiv16_fs195_or0 = f_arrdiv16_fs195_and1 | f_arrdiv16_fs195_and0;
  assign f_arrdiv16_fs196_xor0 = f_arrdiv16_mux2to1168_xor0 ^ b[4];
  assign f_arrdiv16_fs196_not0 = ~f_arrdiv16_mux2to1168_xor0;
  assign f_arrdiv16_fs196_and0 = f_arrdiv16_fs196_not0 & b[4];
  assign f_arrdiv16_fs196_xor1 = f_arrdiv16_fs195_or0 ^ f_arrdiv16_fs196_xor0;
  assign f_arrdiv16_fs196_not1 = ~f_arrdiv16_fs196_xor0;
  assign f_arrdiv16_fs196_and1 = f_arrdiv16_fs196_not1 & f_arrdiv16_fs195_or0;
  assign f_arrdiv16_fs196_or0 = f_arrdiv16_fs196_and1 | f_arrdiv16_fs196_and0;
  assign f_arrdiv16_fs197_xor0 = f_arrdiv16_mux2to1169_xor0 ^ b[5];
  assign f_arrdiv16_fs197_not0 = ~f_arrdiv16_mux2to1169_xor0;
  assign f_arrdiv16_fs197_and0 = f_arrdiv16_fs197_not0 & b[5];
  assign f_arrdiv16_fs197_xor1 = f_arrdiv16_fs196_or0 ^ f_arrdiv16_fs197_xor0;
  assign f_arrdiv16_fs197_not1 = ~f_arrdiv16_fs197_xor0;
  assign f_arrdiv16_fs197_and1 = f_arrdiv16_fs197_not1 & f_arrdiv16_fs196_or0;
  assign f_arrdiv16_fs197_or0 = f_arrdiv16_fs197_and1 | f_arrdiv16_fs197_and0;
  assign f_arrdiv16_fs198_xor0 = f_arrdiv16_mux2to1170_xor0 ^ b[6];
  assign f_arrdiv16_fs198_not0 = ~f_arrdiv16_mux2to1170_xor0;
  assign f_arrdiv16_fs198_and0 = f_arrdiv16_fs198_not0 & b[6];
  assign f_arrdiv16_fs198_xor1 = f_arrdiv16_fs197_or0 ^ f_arrdiv16_fs198_xor0;
  assign f_arrdiv16_fs198_not1 = ~f_arrdiv16_fs198_xor0;
  assign f_arrdiv16_fs198_and1 = f_arrdiv16_fs198_not1 & f_arrdiv16_fs197_or0;
  assign f_arrdiv16_fs198_or0 = f_arrdiv16_fs198_and1 | f_arrdiv16_fs198_and0;
  assign f_arrdiv16_fs199_xor0 = f_arrdiv16_mux2to1171_xor0 ^ b[7];
  assign f_arrdiv16_fs199_not0 = ~f_arrdiv16_mux2to1171_xor0;
  assign f_arrdiv16_fs199_and0 = f_arrdiv16_fs199_not0 & b[7];
  assign f_arrdiv16_fs199_xor1 = f_arrdiv16_fs198_or0 ^ f_arrdiv16_fs199_xor0;
  assign f_arrdiv16_fs199_not1 = ~f_arrdiv16_fs199_xor0;
  assign f_arrdiv16_fs199_and1 = f_arrdiv16_fs199_not1 & f_arrdiv16_fs198_or0;
  assign f_arrdiv16_fs199_or0 = f_arrdiv16_fs199_and1 | f_arrdiv16_fs199_and0;
  assign f_arrdiv16_fs200_xor0 = f_arrdiv16_mux2to1172_xor0 ^ b[8];
  assign f_arrdiv16_fs200_not0 = ~f_arrdiv16_mux2to1172_xor0;
  assign f_arrdiv16_fs200_and0 = f_arrdiv16_fs200_not0 & b[8];
  assign f_arrdiv16_fs200_xor1 = f_arrdiv16_fs199_or0 ^ f_arrdiv16_fs200_xor0;
  assign f_arrdiv16_fs200_not1 = ~f_arrdiv16_fs200_xor0;
  assign f_arrdiv16_fs200_and1 = f_arrdiv16_fs200_not1 & f_arrdiv16_fs199_or0;
  assign f_arrdiv16_fs200_or0 = f_arrdiv16_fs200_and1 | f_arrdiv16_fs200_and0;
  assign f_arrdiv16_fs201_xor0 = f_arrdiv16_mux2to1173_xor0 ^ b[9];
  assign f_arrdiv16_fs201_not0 = ~f_arrdiv16_mux2to1173_xor0;
  assign f_arrdiv16_fs201_and0 = f_arrdiv16_fs201_not0 & b[9];
  assign f_arrdiv16_fs201_xor1 = f_arrdiv16_fs200_or0 ^ f_arrdiv16_fs201_xor0;
  assign f_arrdiv16_fs201_not1 = ~f_arrdiv16_fs201_xor0;
  assign f_arrdiv16_fs201_and1 = f_arrdiv16_fs201_not1 & f_arrdiv16_fs200_or0;
  assign f_arrdiv16_fs201_or0 = f_arrdiv16_fs201_and1 | f_arrdiv16_fs201_and0;
  assign f_arrdiv16_fs202_xor0 = f_arrdiv16_mux2to1174_xor0 ^ b[10];
  assign f_arrdiv16_fs202_not0 = ~f_arrdiv16_mux2to1174_xor0;
  assign f_arrdiv16_fs202_and0 = f_arrdiv16_fs202_not0 & b[10];
  assign f_arrdiv16_fs202_xor1 = f_arrdiv16_fs201_or0 ^ f_arrdiv16_fs202_xor0;
  assign f_arrdiv16_fs202_not1 = ~f_arrdiv16_fs202_xor0;
  assign f_arrdiv16_fs202_and1 = f_arrdiv16_fs202_not1 & f_arrdiv16_fs201_or0;
  assign f_arrdiv16_fs202_or0 = f_arrdiv16_fs202_and1 | f_arrdiv16_fs202_and0;
  assign f_arrdiv16_fs203_xor0 = f_arrdiv16_mux2to1175_xor0 ^ b[11];
  assign f_arrdiv16_fs203_not0 = ~f_arrdiv16_mux2to1175_xor0;
  assign f_arrdiv16_fs203_and0 = f_arrdiv16_fs203_not0 & b[11];
  assign f_arrdiv16_fs203_xor1 = f_arrdiv16_fs202_or0 ^ f_arrdiv16_fs203_xor0;
  assign f_arrdiv16_fs203_not1 = ~f_arrdiv16_fs203_xor0;
  assign f_arrdiv16_fs203_and1 = f_arrdiv16_fs203_not1 & f_arrdiv16_fs202_or0;
  assign f_arrdiv16_fs203_or0 = f_arrdiv16_fs203_and1 | f_arrdiv16_fs203_and0;
  assign f_arrdiv16_fs204_xor0 = f_arrdiv16_mux2to1176_xor0 ^ b[12];
  assign f_arrdiv16_fs204_not0 = ~f_arrdiv16_mux2to1176_xor0;
  assign f_arrdiv16_fs204_and0 = f_arrdiv16_fs204_not0 & b[12];
  assign f_arrdiv16_fs204_xor1 = f_arrdiv16_fs203_or0 ^ f_arrdiv16_fs204_xor0;
  assign f_arrdiv16_fs204_not1 = ~f_arrdiv16_fs204_xor0;
  assign f_arrdiv16_fs204_and1 = f_arrdiv16_fs204_not1 & f_arrdiv16_fs203_or0;
  assign f_arrdiv16_fs204_or0 = f_arrdiv16_fs204_and1 | f_arrdiv16_fs204_and0;
  assign f_arrdiv16_fs205_xor0 = f_arrdiv16_mux2to1177_xor0 ^ b[13];
  assign f_arrdiv16_fs205_not0 = ~f_arrdiv16_mux2to1177_xor0;
  assign f_arrdiv16_fs205_and0 = f_arrdiv16_fs205_not0 & b[13];
  assign f_arrdiv16_fs205_xor1 = f_arrdiv16_fs204_or0 ^ f_arrdiv16_fs205_xor0;
  assign f_arrdiv16_fs205_not1 = ~f_arrdiv16_fs205_xor0;
  assign f_arrdiv16_fs205_and1 = f_arrdiv16_fs205_not1 & f_arrdiv16_fs204_or0;
  assign f_arrdiv16_fs205_or0 = f_arrdiv16_fs205_and1 | f_arrdiv16_fs205_and0;
  assign f_arrdiv16_fs206_xor0 = f_arrdiv16_mux2to1178_xor0 ^ b[14];
  assign f_arrdiv16_fs206_not0 = ~f_arrdiv16_mux2to1178_xor0;
  assign f_arrdiv16_fs206_and0 = f_arrdiv16_fs206_not0 & b[14];
  assign f_arrdiv16_fs206_xor1 = f_arrdiv16_fs205_or0 ^ f_arrdiv16_fs206_xor0;
  assign f_arrdiv16_fs206_not1 = ~f_arrdiv16_fs206_xor0;
  assign f_arrdiv16_fs206_and1 = f_arrdiv16_fs206_not1 & f_arrdiv16_fs205_or0;
  assign f_arrdiv16_fs206_or0 = f_arrdiv16_fs206_and1 | f_arrdiv16_fs206_and0;
  assign f_arrdiv16_fs207_xor0 = f_arrdiv16_mux2to1179_xor0 ^ b[15];
  assign f_arrdiv16_fs207_not0 = ~f_arrdiv16_mux2to1179_xor0;
  assign f_arrdiv16_fs207_and0 = f_arrdiv16_fs207_not0 & b[15];
  assign f_arrdiv16_fs207_xor1 = f_arrdiv16_fs206_or0 ^ f_arrdiv16_fs207_xor0;
  assign f_arrdiv16_fs207_not1 = ~f_arrdiv16_fs207_xor0;
  assign f_arrdiv16_fs207_and1 = f_arrdiv16_fs207_not1 & f_arrdiv16_fs206_or0;
  assign f_arrdiv16_fs207_or0 = f_arrdiv16_fs207_and1 | f_arrdiv16_fs207_and0;
  assign f_arrdiv16_mux2to1180_and0 = a[3] & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1180_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1180_and1 = f_arrdiv16_fs192_xor0 & f_arrdiv16_mux2to1180_not0;
  assign f_arrdiv16_mux2to1180_xor0 = f_arrdiv16_mux2to1180_and0 ^ f_arrdiv16_mux2to1180_and1;
  assign f_arrdiv16_mux2to1181_and0 = f_arrdiv16_mux2to1165_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1181_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1181_and1 = f_arrdiv16_fs193_xor1 & f_arrdiv16_mux2to1181_not0;
  assign f_arrdiv16_mux2to1181_xor0 = f_arrdiv16_mux2to1181_and0 ^ f_arrdiv16_mux2to1181_and1;
  assign f_arrdiv16_mux2to1182_and0 = f_arrdiv16_mux2to1166_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1182_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1182_and1 = f_arrdiv16_fs194_xor1 & f_arrdiv16_mux2to1182_not0;
  assign f_arrdiv16_mux2to1182_xor0 = f_arrdiv16_mux2to1182_and0 ^ f_arrdiv16_mux2to1182_and1;
  assign f_arrdiv16_mux2to1183_and0 = f_arrdiv16_mux2to1167_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1183_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1183_and1 = f_arrdiv16_fs195_xor1 & f_arrdiv16_mux2to1183_not0;
  assign f_arrdiv16_mux2to1183_xor0 = f_arrdiv16_mux2to1183_and0 ^ f_arrdiv16_mux2to1183_and1;
  assign f_arrdiv16_mux2to1184_and0 = f_arrdiv16_mux2to1168_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1184_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1184_and1 = f_arrdiv16_fs196_xor1 & f_arrdiv16_mux2to1184_not0;
  assign f_arrdiv16_mux2to1184_xor0 = f_arrdiv16_mux2to1184_and0 ^ f_arrdiv16_mux2to1184_and1;
  assign f_arrdiv16_mux2to1185_and0 = f_arrdiv16_mux2to1169_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1185_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1185_and1 = f_arrdiv16_fs197_xor1 & f_arrdiv16_mux2to1185_not0;
  assign f_arrdiv16_mux2to1185_xor0 = f_arrdiv16_mux2to1185_and0 ^ f_arrdiv16_mux2to1185_and1;
  assign f_arrdiv16_mux2to1186_and0 = f_arrdiv16_mux2to1170_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1186_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1186_and1 = f_arrdiv16_fs198_xor1 & f_arrdiv16_mux2to1186_not0;
  assign f_arrdiv16_mux2to1186_xor0 = f_arrdiv16_mux2to1186_and0 ^ f_arrdiv16_mux2to1186_and1;
  assign f_arrdiv16_mux2to1187_and0 = f_arrdiv16_mux2to1171_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1187_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1187_and1 = f_arrdiv16_fs199_xor1 & f_arrdiv16_mux2to1187_not0;
  assign f_arrdiv16_mux2to1187_xor0 = f_arrdiv16_mux2to1187_and0 ^ f_arrdiv16_mux2to1187_and1;
  assign f_arrdiv16_mux2to1188_and0 = f_arrdiv16_mux2to1172_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1188_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1188_and1 = f_arrdiv16_fs200_xor1 & f_arrdiv16_mux2to1188_not0;
  assign f_arrdiv16_mux2to1188_xor0 = f_arrdiv16_mux2to1188_and0 ^ f_arrdiv16_mux2to1188_and1;
  assign f_arrdiv16_mux2to1189_and0 = f_arrdiv16_mux2to1173_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1189_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1189_and1 = f_arrdiv16_fs201_xor1 & f_arrdiv16_mux2to1189_not0;
  assign f_arrdiv16_mux2to1189_xor0 = f_arrdiv16_mux2to1189_and0 ^ f_arrdiv16_mux2to1189_and1;
  assign f_arrdiv16_mux2to1190_and0 = f_arrdiv16_mux2to1174_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1190_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1190_and1 = f_arrdiv16_fs202_xor1 & f_arrdiv16_mux2to1190_not0;
  assign f_arrdiv16_mux2to1190_xor0 = f_arrdiv16_mux2to1190_and0 ^ f_arrdiv16_mux2to1190_and1;
  assign f_arrdiv16_mux2to1191_and0 = f_arrdiv16_mux2to1175_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1191_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1191_and1 = f_arrdiv16_fs203_xor1 & f_arrdiv16_mux2to1191_not0;
  assign f_arrdiv16_mux2to1191_xor0 = f_arrdiv16_mux2to1191_and0 ^ f_arrdiv16_mux2to1191_and1;
  assign f_arrdiv16_mux2to1192_and0 = f_arrdiv16_mux2to1176_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1192_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1192_and1 = f_arrdiv16_fs204_xor1 & f_arrdiv16_mux2to1192_not0;
  assign f_arrdiv16_mux2to1192_xor0 = f_arrdiv16_mux2to1192_and0 ^ f_arrdiv16_mux2to1192_and1;
  assign f_arrdiv16_mux2to1193_and0 = f_arrdiv16_mux2to1177_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1193_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1193_and1 = f_arrdiv16_fs205_xor1 & f_arrdiv16_mux2to1193_not0;
  assign f_arrdiv16_mux2to1193_xor0 = f_arrdiv16_mux2to1193_and0 ^ f_arrdiv16_mux2to1193_and1;
  assign f_arrdiv16_mux2to1194_and0 = f_arrdiv16_mux2to1178_xor0 & f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1194_not0 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_mux2to1194_and1 = f_arrdiv16_fs206_xor1 & f_arrdiv16_mux2to1194_not0;
  assign f_arrdiv16_mux2to1194_xor0 = f_arrdiv16_mux2to1194_and0 ^ f_arrdiv16_mux2to1194_and1;
  assign f_arrdiv16_not12 = ~f_arrdiv16_fs207_or0;
  assign f_arrdiv16_fs208_xor0 = a[2] ^ b[0];
  assign f_arrdiv16_fs208_not0 = ~a[2];
  assign f_arrdiv16_fs208_and0 = f_arrdiv16_fs208_not0 & b[0];
  assign f_arrdiv16_fs208_not1 = ~f_arrdiv16_fs208_xor0;
  assign f_arrdiv16_fs209_xor0 = f_arrdiv16_mux2to1180_xor0 ^ b[1];
  assign f_arrdiv16_fs209_not0 = ~f_arrdiv16_mux2to1180_xor0;
  assign f_arrdiv16_fs209_and0 = f_arrdiv16_fs209_not0 & b[1];
  assign f_arrdiv16_fs209_xor1 = f_arrdiv16_fs208_and0 ^ f_arrdiv16_fs209_xor0;
  assign f_arrdiv16_fs209_not1 = ~f_arrdiv16_fs209_xor0;
  assign f_arrdiv16_fs209_and1 = f_arrdiv16_fs209_not1 & f_arrdiv16_fs208_and0;
  assign f_arrdiv16_fs209_or0 = f_arrdiv16_fs209_and1 | f_arrdiv16_fs209_and0;
  assign f_arrdiv16_fs210_xor0 = f_arrdiv16_mux2to1181_xor0 ^ b[2];
  assign f_arrdiv16_fs210_not0 = ~f_arrdiv16_mux2to1181_xor0;
  assign f_arrdiv16_fs210_and0 = f_arrdiv16_fs210_not0 & b[2];
  assign f_arrdiv16_fs210_xor1 = f_arrdiv16_fs209_or0 ^ f_arrdiv16_fs210_xor0;
  assign f_arrdiv16_fs210_not1 = ~f_arrdiv16_fs210_xor0;
  assign f_arrdiv16_fs210_and1 = f_arrdiv16_fs210_not1 & f_arrdiv16_fs209_or0;
  assign f_arrdiv16_fs210_or0 = f_arrdiv16_fs210_and1 | f_arrdiv16_fs210_and0;
  assign f_arrdiv16_fs211_xor0 = f_arrdiv16_mux2to1182_xor0 ^ b[3];
  assign f_arrdiv16_fs211_not0 = ~f_arrdiv16_mux2to1182_xor0;
  assign f_arrdiv16_fs211_and0 = f_arrdiv16_fs211_not0 & b[3];
  assign f_arrdiv16_fs211_xor1 = f_arrdiv16_fs210_or0 ^ f_arrdiv16_fs211_xor0;
  assign f_arrdiv16_fs211_not1 = ~f_arrdiv16_fs211_xor0;
  assign f_arrdiv16_fs211_and1 = f_arrdiv16_fs211_not1 & f_arrdiv16_fs210_or0;
  assign f_arrdiv16_fs211_or0 = f_arrdiv16_fs211_and1 | f_arrdiv16_fs211_and0;
  assign f_arrdiv16_fs212_xor0 = f_arrdiv16_mux2to1183_xor0 ^ b[4];
  assign f_arrdiv16_fs212_not0 = ~f_arrdiv16_mux2to1183_xor0;
  assign f_arrdiv16_fs212_and0 = f_arrdiv16_fs212_not0 & b[4];
  assign f_arrdiv16_fs212_xor1 = f_arrdiv16_fs211_or0 ^ f_arrdiv16_fs212_xor0;
  assign f_arrdiv16_fs212_not1 = ~f_arrdiv16_fs212_xor0;
  assign f_arrdiv16_fs212_and1 = f_arrdiv16_fs212_not1 & f_arrdiv16_fs211_or0;
  assign f_arrdiv16_fs212_or0 = f_arrdiv16_fs212_and1 | f_arrdiv16_fs212_and0;
  assign f_arrdiv16_fs213_xor0 = f_arrdiv16_mux2to1184_xor0 ^ b[5];
  assign f_arrdiv16_fs213_not0 = ~f_arrdiv16_mux2to1184_xor0;
  assign f_arrdiv16_fs213_and0 = f_arrdiv16_fs213_not0 & b[5];
  assign f_arrdiv16_fs213_xor1 = f_arrdiv16_fs212_or0 ^ f_arrdiv16_fs213_xor0;
  assign f_arrdiv16_fs213_not1 = ~f_arrdiv16_fs213_xor0;
  assign f_arrdiv16_fs213_and1 = f_arrdiv16_fs213_not1 & f_arrdiv16_fs212_or0;
  assign f_arrdiv16_fs213_or0 = f_arrdiv16_fs213_and1 | f_arrdiv16_fs213_and0;
  assign f_arrdiv16_fs214_xor0 = f_arrdiv16_mux2to1185_xor0 ^ b[6];
  assign f_arrdiv16_fs214_not0 = ~f_arrdiv16_mux2to1185_xor0;
  assign f_arrdiv16_fs214_and0 = f_arrdiv16_fs214_not0 & b[6];
  assign f_arrdiv16_fs214_xor1 = f_arrdiv16_fs213_or0 ^ f_arrdiv16_fs214_xor0;
  assign f_arrdiv16_fs214_not1 = ~f_arrdiv16_fs214_xor0;
  assign f_arrdiv16_fs214_and1 = f_arrdiv16_fs214_not1 & f_arrdiv16_fs213_or0;
  assign f_arrdiv16_fs214_or0 = f_arrdiv16_fs214_and1 | f_arrdiv16_fs214_and0;
  assign f_arrdiv16_fs215_xor0 = f_arrdiv16_mux2to1186_xor0 ^ b[7];
  assign f_arrdiv16_fs215_not0 = ~f_arrdiv16_mux2to1186_xor0;
  assign f_arrdiv16_fs215_and0 = f_arrdiv16_fs215_not0 & b[7];
  assign f_arrdiv16_fs215_xor1 = f_arrdiv16_fs214_or0 ^ f_arrdiv16_fs215_xor0;
  assign f_arrdiv16_fs215_not1 = ~f_arrdiv16_fs215_xor0;
  assign f_arrdiv16_fs215_and1 = f_arrdiv16_fs215_not1 & f_arrdiv16_fs214_or0;
  assign f_arrdiv16_fs215_or0 = f_arrdiv16_fs215_and1 | f_arrdiv16_fs215_and0;
  assign f_arrdiv16_fs216_xor0 = f_arrdiv16_mux2to1187_xor0 ^ b[8];
  assign f_arrdiv16_fs216_not0 = ~f_arrdiv16_mux2to1187_xor0;
  assign f_arrdiv16_fs216_and0 = f_arrdiv16_fs216_not0 & b[8];
  assign f_arrdiv16_fs216_xor1 = f_arrdiv16_fs215_or0 ^ f_arrdiv16_fs216_xor0;
  assign f_arrdiv16_fs216_not1 = ~f_arrdiv16_fs216_xor0;
  assign f_arrdiv16_fs216_and1 = f_arrdiv16_fs216_not1 & f_arrdiv16_fs215_or0;
  assign f_arrdiv16_fs216_or0 = f_arrdiv16_fs216_and1 | f_arrdiv16_fs216_and0;
  assign f_arrdiv16_fs217_xor0 = f_arrdiv16_mux2to1188_xor0 ^ b[9];
  assign f_arrdiv16_fs217_not0 = ~f_arrdiv16_mux2to1188_xor0;
  assign f_arrdiv16_fs217_and0 = f_arrdiv16_fs217_not0 & b[9];
  assign f_arrdiv16_fs217_xor1 = f_arrdiv16_fs216_or0 ^ f_arrdiv16_fs217_xor0;
  assign f_arrdiv16_fs217_not1 = ~f_arrdiv16_fs217_xor0;
  assign f_arrdiv16_fs217_and1 = f_arrdiv16_fs217_not1 & f_arrdiv16_fs216_or0;
  assign f_arrdiv16_fs217_or0 = f_arrdiv16_fs217_and1 | f_arrdiv16_fs217_and0;
  assign f_arrdiv16_fs218_xor0 = f_arrdiv16_mux2to1189_xor0 ^ b[10];
  assign f_arrdiv16_fs218_not0 = ~f_arrdiv16_mux2to1189_xor0;
  assign f_arrdiv16_fs218_and0 = f_arrdiv16_fs218_not0 & b[10];
  assign f_arrdiv16_fs218_xor1 = f_arrdiv16_fs217_or0 ^ f_arrdiv16_fs218_xor0;
  assign f_arrdiv16_fs218_not1 = ~f_arrdiv16_fs218_xor0;
  assign f_arrdiv16_fs218_and1 = f_arrdiv16_fs218_not1 & f_arrdiv16_fs217_or0;
  assign f_arrdiv16_fs218_or0 = f_arrdiv16_fs218_and1 | f_arrdiv16_fs218_and0;
  assign f_arrdiv16_fs219_xor0 = f_arrdiv16_mux2to1190_xor0 ^ b[11];
  assign f_arrdiv16_fs219_not0 = ~f_arrdiv16_mux2to1190_xor0;
  assign f_arrdiv16_fs219_and0 = f_arrdiv16_fs219_not0 & b[11];
  assign f_arrdiv16_fs219_xor1 = f_arrdiv16_fs218_or0 ^ f_arrdiv16_fs219_xor0;
  assign f_arrdiv16_fs219_not1 = ~f_arrdiv16_fs219_xor0;
  assign f_arrdiv16_fs219_and1 = f_arrdiv16_fs219_not1 & f_arrdiv16_fs218_or0;
  assign f_arrdiv16_fs219_or0 = f_arrdiv16_fs219_and1 | f_arrdiv16_fs219_and0;
  assign f_arrdiv16_fs220_xor0 = f_arrdiv16_mux2to1191_xor0 ^ b[12];
  assign f_arrdiv16_fs220_not0 = ~f_arrdiv16_mux2to1191_xor0;
  assign f_arrdiv16_fs220_and0 = f_arrdiv16_fs220_not0 & b[12];
  assign f_arrdiv16_fs220_xor1 = f_arrdiv16_fs219_or0 ^ f_arrdiv16_fs220_xor0;
  assign f_arrdiv16_fs220_not1 = ~f_arrdiv16_fs220_xor0;
  assign f_arrdiv16_fs220_and1 = f_arrdiv16_fs220_not1 & f_arrdiv16_fs219_or0;
  assign f_arrdiv16_fs220_or0 = f_arrdiv16_fs220_and1 | f_arrdiv16_fs220_and0;
  assign f_arrdiv16_fs221_xor0 = f_arrdiv16_mux2to1192_xor0 ^ b[13];
  assign f_arrdiv16_fs221_not0 = ~f_arrdiv16_mux2to1192_xor0;
  assign f_arrdiv16_fs221_and0 = f_arrdiv16_fs221_not0 & b[13];
  assign f_arrdiv16_fs221_xor1 = f_arrdiv16_fs220_or0 ^ f_arrdiv16_fs221_xor0;
  assign f_arrdiv16_fs221_not1 = ~f_arrdiv16_fs221_xor0;
  assign f_arrdiv16_fs221_and1 = f_arrdiv16_fs221_not1 & f_arrdiv16_fs220_or0;
  assign f_arrdiv16_fs221_or0 = f_arrdiv16_fs221_and1 | f_arrdiv16_fs221_and0;
  assign f_arrdiv16_fs222_xor0 = f_arrdiv16_mux2to1193_xor0 ^ b[14];
  assign f_arrdiv16_fs222_not0 = ~f_arrdiv16_mux2to1193_xor0;
  assign f_arrdiv16_fs222_and0 = f_arrdiv16_fs222_not0 & b[14];
  assign f_arrdiv16_fs222_xor1 = f_arrdiv16_fs221_or0 ^ f_arrdiv16_fs222_xor0;
  assign f_arrdiv16_fs222_not1 = ~f_arrdiv16_fs222_xor0;
  assign f_arrdiv16_fs222_and1 = f_arrdiv16_fs222_not1 & f_arrdiv16_fs221_or0;
  assign f_arrdiv16_fs222_or0 = f_arrdiv16_fs222_and1 | f_arrdiv16_fs222_and0;
  assign f_arrdiv16_fs223_xor0 = f_arrdiv16_mux2to1194_xor0 ^ b[15];
  assign f_arrdiv16_fs223_not0 = ~f_arrdiv16_mux2to1194_xor0;
  assign f_arrdiv16_fs223_and0 = f_arrdiv16_fs223_not0 & b[15];
  assign f_arrdiv16_fs223_xor1 = f_arrdiv16_fs222_or0 ^ f_arrdiv16_fs223_xor0;
  assign f_arrdiv16_fs223_not1 = ~f_arrdiv16_fs223_xor0;
  assign f_arrdiv16_fs223_and1 = f_arrdiv16_fs223_not1 & f_arrdiv16_fs222_or0;
  assign f_arrdiv16_fs223_or0 = f_arrdiv16_fs223_and1 | f_arrdiv16_fs223_and0;
  assign f_arrdiv16_mux2to1195_and0 = a[2] & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1195_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1195_and1 = f_arrdiv16_fs208_xor0 & f_arrdiv16_mux2to1195_not0;
  assign f_arrdiv16_mux2to1195_xor0 = f_arrdiv16_mux2to1195_and0 ^ f_arrdiv16_mux2to1195_and1;
  assign f_arrdiv16_mux2to1196_and0 = f_arrdiv16_mux2to1180_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1196_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1196_and1 = f_arrdiv16_fs209_xor1 & f_arrdiv16_mux2to1196_not0;
  assign f_arrdiv16_mux2to1196_xor0 = f_arrdiv16_mux2to1196_and0 ^ f_arrdiv16_mux2to1196_and1;
  assign f_arrdiv16_mux2to1197_and0 = f_arrdiv16_mux2to1181_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1197_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1197_and1 = f_arrdiv16_fs210_xor1 & f_arrdiv16_mux2to1197_not0;
  assign f_arrdiv16_mux2to1197_xor0 = f_arrdiv16_mux2to1197_and0 ^ f_arrdiv16_mux2to1197_and1;
  assign f_arrdiv16_mux2to1198_and0 = f_arrdiv16_mux2to1182_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1198_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1198_and1 = f_arrdiv16_fs211_xor1 & f_arrdiv16_mux2to1198_not0;
  assign f_arrdiv16_mux2to1198_xor0 = f_arrdiv16_mux2to1198_and0 ^ f_arrdiv16_mux2to1198_and1;
  assign f_arrdiv16_mux2to1199_and0 = f_arrdiv16_mux2to1183_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1199_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1199_and1 = f_arrdiv16_fs212_xor1 & f_arrdiv16_mux2to1199_not0;
  assign f_arrdiv16_mux2to1199_xor0 = f_arrdiv16_mux2to1199_and0 ^ f_arrdiv16_mux2to1199_and1;
  assign f_arrdiv16_mux2to1200_and0 = f_arrdiv16_mux2to1184_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1200_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1200_and1 = f_arrdiv16_fs213_xor1 & f_arrdiv16_mux2to1200_not0;
  assign f_arrdiv16_mux2to1200_xor0 = f_arrdiv16_mux2to1200_and0 ^ f_arrdiv16_mux2to1200_and1;
  assign f_arrdiv16_mux2to1201_and0 = f_arrdiv16_mux2to1185_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1201_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1201_and1 = f_arrdiv16_fs214_xor1 & f_arrdiv16_mux2to1201_not0;
  assign f_arrdiv16_mux2to1201_xor0 = f_arrdiv16_mux2to1201_and0 ^ f_arrdiv16_mux2to1201_and1;
  assign f_arrdiv16_mux2to1202_and0 = f_arrdiv16_mux2to1186_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1202_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1202_and1 = f_arrdiv16_fs215_xor1 & f_arrdiv16_mux2to1202_not0;
  assign f_arrdiv16_mux2to1202_xor0 = f_arrdiv16_mux2to1202_and0 ^ f_arrdiv16_mux2to1202_and1;
  assign f_arrdiv16_mux2to1203_and0 = f_arrdiv16_mux2to1187_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1203_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1203_and1 = f_arrdiv16_fs216_xor1 & f_arrdiv16_mux2to1203_not0;
  assign f_arrdiv16_mux2to1203_xor0 = f_arrdiv16_mux2to1203_and0 ^ f_arrdiv16_mux2to1203_and1;
  assign f_arrdiv16_mux2to1204_and0 = f_arrdiv16_mux2to1188_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1204_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1204_and1 = f_arrdiv16_fs217_xor1 & f_arrdiv16_mux2to1204_not0;
  assign f_arrdiv16_mux2to1204_xor0 = f_arrdiv16_mux2to1204_and0 ^ f_arrdiv16_mux2to1204_and1;
  assign f_arrdiv16_mux2to1205_and0 = f_arrdiv16_mux2to1189_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1205_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1205_and1 = f_arrdiv16_fs218_xor1 & f_arrdiv16_mux2to1205_not0;
  assign f_arrdiv16_mux2to1205_xor0 = f_arrdiv16_mux2to1205_and0 ^ f_arrdiv16_mux2to1205_and1;
  assign f_arrdiv16_mux2to1206_and0 = f_arrdiv16_mux2to1190_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1206_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1206_and1 = f_arrdiv16_fs219_xor1 & f_arrdiv16_mux2to1206_not0;
  assign f_arrdiv16_mux2to1206_xor0 = f_arrdiv16_mux2to1206_and0 ^ f_arrdiv16_mux2to1206_and1;
  assign f_arrdiv16_mux2to1207_and0 = f_arrdiv16_mux2to1191_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1207_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1207_and1 = f_arrdiv16_fs220_xor1 & f_arrdiv16_mux2to1207_not0;
  assign f_arrdiv16_mux2to1207_xor0 = f_arrdiv16_mux2to1207_and0 ^ f_arrdiv16_mux2to1207_and1;
  assign f_arrdiv16_mux2to1208_and0 = f_arrdiv16_mux2to1192_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1208_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1208_and1 = f_arrdiv16_fs221_xor1 & f_arrdiv16_mux2to1208_not0;
  assign f_arrdiv16_mux2to1208_xor0 = f_arrdiv16_mux2to1208_and0 ^ f_arrdiv16_mux2to1208_and1;
  assign f_arrdiv16_mux2to1209_and0 = f_arrdiv16_mux2to1193_xor0 & f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1209_not0 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_mux2to1209_and1 = f_arrdiv16_fs222_xor1 & f_arrdiv16_mux2to1209_not0;
  assign f_arrdiv16_mux2to1209_xor0 = f_arrdiv16_mux2to1209_and0 ^ f_arrdiv16_mux2to1209_and1;
  assign f_arrdiv16_not13 = ~f_arrdiv16_fs223_or0;
  assign f_arrdiv16_fs224_xor0 = a[1] ^ b[0];
  assign f_arrdiv16_fs224_not0 = ~a[1];
  assign f_arrdiv16_fs224_and0 = f_arrdiv16_fs224_not0 & b[0];
  assign f_arrdiv16_fs224_not1 = ~f_arrdiv16_fs224_xor0;
  assign f_arrdiv16_fs225_xor0 = f_arrdiv16_mux2to1195_xor0 ^ b[1];
  assign f_arrdiv16_fs225_not0 = ~f_arrdiv16_mux2to1195_xor0;
  assign f_arrdiv16_fs225_and0 = f_arrdiv16_fs225_not0 & b[1];
  assign f_arrdiv16_fs225_xor1 = f_arrdiv16_fs224_and0 ^ f_arrdiv16_fs225_xor0;
  assign f_arrdiv16_fs225_not1 = ~f_arrdiv16_fs225_xor0;
  assign f_arrdiv16_fs225_and1 = f_arrdiv16_fs225_not1 & f_arrdiv16_fs224_and0;
  assign f_arrdiv16_fs225_or0 = f_arrdiv16_fs225_and1 | f_arrdiv16_fs225_and0;
  assign f_arrdiv16_fs226_xor0 = f_arrdiv16_mux2to1196_xor0 ^ b[2];
  assign f_arrdiv16_fs226_not0 = ~f_arrdiv16_mux2to1196_xor0;
  assign f_arrdiv16_fs226_and0 = f_arrdiv16_fs226_not0 & b[2];
  assign f_arrdiv16_fs226_xor1 = f_arrdiv16_fs225_or0 ^ f_arrdiv16_fs226_xor0;
  assign f_arrdiv16_fs226_not1 = ~f_arrdiv16_fs226_xor0;
  assign f_arrdiv16_fs226_and1 = f_arrdiv16_fs226_not1 & f_arrdiv16_fs225_or0;
  assign f_arrdiv16_fs226_or0 = f_arrdiv16_fs226_and1 | f_arrdiv16_fs226_and0;
  assign f_arrdiv16_fs227_xor0 = f_arrdiv16_mux2to1197_xor0 ^ b[3];
  assign f_arrdiv16_fs227_not0 = ~f_arrdiv16_mux2to1197_xor0;
  assign f_arrdiv16_fs227_and0 = f_arrdiv16_fs227_not0 & b[3];
  assign f_arrdiv16_fs227_xor1 = f_arrdiv16_fs226_or0 ^ f_arrdiv16_fs227_xor0;
  assign f_arrdiv16_fs227_not1 = ~f_arrdiv16_fs227_xor0;
  assign f_arrdiv16_fs227_and1 = f_arrdiv16_fs227_not1 & f_arrdiv16_fs226_or0;
  assign f_arrdiv16_fs227_or0 = f_arrdiv16_fs227_and1 | f_arrdiv16_fs227_and0;
  assign f_arrdiv16_fs228_xor0 = f_arrdiv16_mux2to1198_xor0 ^ b[4];
  assign f_arrdiv16_fs228_not0 = ~f_arrdiv16_mux2to1198_xor0;
  assign f_arrdiv16_fs228_and0 = f_arrdiv16_fs228_not0 & b[4];
  assign f_arrdiv16_fs228_xor1 = f_arrdiv16_fs227_or0 ^ f_arrdiv16_fs228_xor0;
  assign f_arrdiv16_fs228_not1 = ~f_arrdiv16_fs228_xor0;
  assign f_arrdiv16_fs228_and1 = f_arrdiv16_fs228_not1 & f_arrdiv16_fs227_or0;
  assign f_arrdiv16_fs228_or0 = f_arrdiv16_fs228_and1 | f_arrdiv16_fs228_and0;
  assign f_arrdiv16_fs229_xor0 = f_arrdiv16_mux2to1199_xor0 ^ b[5];
  assign f_arrdiv16_fs229_not0 = ~f_arrdiv16_mux2to1199_xor0;
  assign f_arrdiv16_fs229_and0 = f_arrdiv16_fs229_not0 & b[5];
  assign f_arrdiv16_fs229_xor1 = f_arrdiv16_fs228_or0 ^ f_arrdiv16_fs229_xor0;
  assign f_arrdiv16_fs229_not1 = ~f_arrdiv16_fs229_xor0;
  assign f_arrdiv16_fs229_and1 = f_arrdiv16_fs229_not1 & f_arrdiv16_fs228_or0;
  assign f_arrdiv16_fs229_or0 = f_arrdiv16_fs229_and1 | f_arrdiv16_fs229_and0;
  assign f_arrdiv16_fs230_xor0 = f_arrdiv16_mux2to1200_xor0 ^ b[6];
  assign f_arrdiv16_fs230_not0 = ~f_arrdiv16_mux2to1200_xor0;
  assign f_arrdiv16_fs230_and0 = f_arrdiv16_fs230_not0 & b[6];
  assign f_arrdiv16_fs230_xor1 = f_arrdiv16_fs229_or0 ^ f_arrdiv16_fs230_xor0;
  assign f_arrdiv16_fs230_not1 = ~f_arrdiv16_fs230_xor0;
  assign f_arrdiv16_fs230_and1 = f_arrdiv16_fs230_not1 & f_arrdiv16_fs229_or0;
  assign f_arrdiv16_fs230_or0 = f_arrdiv16_fs230_and1 | f_arrdiv16_fs230_and0;
  assign f_arrdiv16_fs231_xor0 = f_arrdiv16_mux2to1201_xor0 ^ b[7];
  assign f_arrdiv16_fs231_not0 = ~f_arrdiv16_mux2to1201_xor0;
  assign f_arrdiv16_fs231_and0 = f_arrdiv16_fs231_not0 & b[7];
  assign f_arrdiv16_fs231_xor1 = f_arrdiv16_fs230_or0 ^ f_arrdiv16_fs231_xor0;
  assign f_arrdiv16_fs231_not1 = ~f_arrdiv16_fs231_xor0;
  assign f_arrdiv16_fs231_and1 = f_arrdiv16_fs231_not1 & f_arrdiv16_fs230_or0;
  assign f_arrdiv16_fs231_or0 = f_arrdiv16_fs231_and1 | f_arrdiv16_fs231_and0;
  assign f_arrdiv16_fs232_xor0 = f_arrdiv16_mux2to1202_xor0 ^ b[8];
  assign f_arrdiv16_fs232_not0 = ~f_arrdiv16_mux2to1202_xor0;
  assign f_arrdiv16_fs232_and0 = f_arrdiv16_fs232_not0 & b[8];
  assign f_arrdiv16_fs232_xor1 = f_arrdiv16_fs231_or0 ^ f_arrdiv16_fs232_xor0;
  assign f_arrdiv16_fs232_not1 = ~f_arrdiv16_fs232_xor0;
  assign f_arrdiv16_fs232_and1 = f_arrdiv16_fs232_not1 & f_arrdiv16_fs231_or0;
  assign f_arrdiv16_fs232_or0 = f_arrdiv16_fs232_and1 | f_arrdiv16_fs232_and0;
  assign f_arrdiv16_fs233_xor0 = f_arrdiv16_mux2to1203_xor0 ^ b[9];
  assign f_arrdiv16_fs233_not0 = ~f_arrdiv16_mux2to1203_xor0;
  assign f_arrdiv16_fs233_and0 = f_arrdiv16_fs233_not0 & b[9];
  assign f_arrdiv16_fs233_xor1 = f_arrdiv16_fs232_or0 ^ f_arrdiv16_fs233_xor0;
  assign f_arrdiv16_fs233_not1 = ~f_arrdiv16_fs233_xor0;
  assign f_arrdiv16_fs233_and1 = f_arrdiv16_fs233_not1 & f_arrdiv16_fs232_or0;
  assign f_arrdiv16_fs233_or0 = f_arrdiv16_fs233_and1 | f_arrdiv16_fs233_and0;
  assign f_arrdiv16_fs234_xor0 = f_arrdiv16_mux2to1204_xor0 ^ b[10];
  assign f_arrdiv16_fs234_not0 = ~f_arrdiv16_mux2to1204_xor0;
  assign f_arrdiv16_fs234_and0 = f_arrdiv16_fs234_not0 & b[10];
  assign f_arrdiv16_fs234_xor1 = f_arrdiv16_fs233_or0 ^ f_arrdiv16_fs234_xor0;
  assign f_arrdiv16_fs234_not1 = ~f_arrdiv16_fs234_xor0;
  assign f_arrdiv16_fs234_and1 = f_arrdiv16_fs234_not1 & f_arrdiv16_fs233_or0;
  assign f_arrdiv16_fs234_or0 = f_arrdiv16_fs234_and1 | f_arrdiv16_fs234_and0;
  assign f_arrdiv16_fs235_xor0 = f_arrdiv16_mux2to1205_xor0 ^ b[11];
  assign f_arrdiv16_fs235_not0 = ~f_arrdiv16_mux2to1205_xor0;
  assign f_arrdiv16_fs235_and0 = f_arrdiv16_fs235_not0 & b[11];
  assign f_arrdiv16_fs235_xor1 = f_arrdiv16_fs234_or0 ^ f_arrdiv16_fs235_xor0;
  assign f_arrdiv16_fs235_not1 = ~f_arrdiv16_fs235_xor0;
  assign f_arrdiv16_fs235_and1 = f_arrdiv16_fs235_not1 & f_arrdiv16_fs234_or0;
  assign f_arrdiv16_fs235_or0 = f_arrdiv16_fs235_and1 | f_arrdiv16_fs235_and0;
  assign f_arrdiv16_fs236_xor0 = f_arrdiv16_mux2to1206_xor0 ^ b[12];
  assign f_arrdiv16_fs236_not0 = ~f_arrdiv16_mux2to1206_xor0;
  assign f_arrdiv16_fs236_and0 = f_arrdiv16_fs236_not0 & b[12];
  assign f_arrdiv16_fs236_xor1 = f_arrdiv16_fs235_or0 ^ f_arrdiv16_fs236_xor0;
  assign f_arrdiv16_fs236_not1 = ~f_arrdiv16_fs236_xor0;
  assign f_arrdiv16_fs236_and1 = f_arrdiv16_fs236_not1 & f_arrdiv16_fs235_or0;
  assign f_arrdiv16_fs236_or0 = f_arrdiv16_fs236_and1 | f_arrdiv16_fs236_and0;
  assign f_arrdiv16_fs237_xor0 = f_arrdiv16_mux2to1207_xor0 ^ b[13];
  assign f_arrdiv16_fs237_not0 = ~f_arrdiv16_mux2to1207_xor0;
  assign f_arrdiv16_fs237_and0 = f_arrdiv16_fs237_not0 & b[13];
  assign f_arrdiv16_fs237_xor1 = f_arrdiv16_fs236_or0 ^ f_arrdiv16_fs237_xor0;
  assign f_arrdiv16_fs237_not1 = ~f_arrdiv16_fs237_xor0;
  assign f_arrdiv16_fs237_and1 = f_arrdiv16_fs237_not1 & f_arrdiv16_fs236_or0;
  assign f_arrdiv16_fs237_or0 = f_arrdiv16_fs237_and1 | f_arrdiv16_fs237_and0;
  assign f_arrdiv16_fs238_xor0 = f_arrdiv16_mux2to1208_xor0 ^ b[14];
  assign f_arrdiv16_fs238_not0 = ~f_arrdiv16_mux2to1208_xor0;
  assign f_arrdiv16_fs238_and0 = f_arrdiv16_fs238_not0 & b[14];
  assign f_arrdiv16_fs238_xor1 = f_arrdiv16_fs237_or0 ^ f_arrdiv16_fs238_xor0;
  assign f_arrdiv16_fs238_not1 = ~f_arrdiv16_fs238_xor0;
  assign f_arrdiv16_fs238_and1 = f_arrdiv16_fs238_not1 & f_arrdiv16_fs237_or0;
  assign f_arrdiv16_fs238_or0 = f_arrdiv16_fs238_and1 | f_arrdiv16_fs238_and0;
  assign f_arrdiv16_fs239_xor0 = f_arrdiv16_mux2to1209_xor0 ^ b[15];
  assign f_arrdiv16_fs239_not0 = ~f_arrdiv16_mux2to1209_xor0;
  assign f_arrdiv16_fs239_and0 = f_arrdiv16_fs239_not0 & b[15];
  assign f_arrdiv16_fs239_xor1 = f_arrdiv16_fs238_or0 ^ f_arrdiv16_fs239_xor0;
  assign f_arrdiv16_fs239_not1 = ~f_arrdiv16_fs239_xor0;
  assign f_arrdiv16_fs239_and1 = f_arrdiv16_fs239_not1 & f_arrdiv16_fs238_or0;
  assign f_arrdiv16_fs239_or0 = f_arrdiv16_fs239_and1 | f_arrdiv16_fs239_and0;
  assign f_arrdiv16_mux2to1210_and0 = a[1] & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1210_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1210_and1 = f_arrdiv16_fs224_xor0 & f_arrdiv16_mux2to1210_not0;
  assign f_arrdiv16_mux2to1210_xor0 = f_arrdiv16_mux2to1210_and0 ^ f_arrdiv16_mux2to1210_and1;
  assign f_arrdiv16_mux2to1211_and0 = f_arrdiv16_mux2to1195_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1211_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1211_and1 = f_arrdiv16_fs225_xor1 & f_arrdiv16_mux2to1211_not0;
  assign f_arrdiv16_mux2to1211_xor0 = f_arrdiv16_mux2to1211_and0 ^ f_arrdiv16_mux2to1211_and1;
  assign f_arrdiv16_mux2to1212_and0 = f_arrdiv16_mux2to1196_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1212_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1212_and1 = f_arrdiv16_fs226_xor1 & f_arrdiv16_mux2to1212_not0;
  assign f_arrdiv16_mux2to1212_xor0 = f_arrdiv16_mux2to1212_and0 ^ f_arrdiv16_mux2to1212_and1;
  assign f_arrdiv16_mux2to1213_and0 = f_arrdiv16_mux2to1197_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1213_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1213_and1 = f_arrdiv16_fs227_xor1 & f_arrdiv16_mux2to1213_not0;
  assign f_arrdiv16_mux2to1213_xor0 = f_arrdiv16_mux2to1213_and0 ^ f_arrdiv16_mux2to1213_and1;
  assign f_arrdiv16_mux2to1214_and0 = f_arrdiv16_mux2to1198_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1214_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1214_and1 = f_arrdiv16_fs228_xor1 & f_arrdiv16_mux2to1214_not0;
  assign f_arrdiv16_mux2to1214_xor0 = f_arrdiv16_mux2to1214_and0 ^ f_arrdiv16_mux2to1214_and1;
  assign f_arrdiv16_mux2to1215_and0 = f_arrdiv16_mux2to1199_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1215_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1215_and1 = f_arrdiv16_fs229_xor1 & f_arrdiv16_mux2to1215_not0;
  assign f_arrdiv16_mux2to1215_xor0 = f_arrdiv16_mux2to1215_and0 ^ f_arrdiv16_mux2to1215_and1;
  assign f_arrdiv16_mux2to1216_and0 = f_arrdiv16_mux2to1200_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1216_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1216_and1 = f_arrdiv16_fs230_xor1 & f_arrdiv16_mux2to1216_not0;
  assign f_arrdiv16_mux2to1216_xor0 = f_arrdiv16_mux2to1216_and0 ^ f_arrdiv16_mux2to1216_and1;
  assign f_arrdiv16_mux2to1217_and0 = f_arrdiv16_mux2to1201_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1217_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1217_and1 = f_arrdiv16_fs231_xor1 & f_arrdiv16_mux2to1217_not0;
  assign f_arrdiv16_mux2to1217_xor0 = f_arrdiv16_mux2to1217_and0 ^ f_arrdiv16_mux2to1217_and1;
  assign f_arrdiv16_mux2to1218_and0 = f_arrdiv16_mux2to1202_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1218_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1218_and1 = f_arrdiv16_fs232_xor1 & f_arrdiv16_mux2to1218_not0;
  assign f_arrdiv16_mux2to1218_xor0 = f_arrdiv16_mux2to1218_and0 ^ f_arrdiv16_mux2to1218_and1;
  assign f_arrdiv16_mux2to1219_and0 = f_arrdiv16_mux2to1203_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1219_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1219_and1 = f_arrdiv16_fs233_xor1 & f_arrdiv16_mux2to1219_not0;
  assign f_arrdiv16_mux2to1219_xor0 = f_arrdiv16_mux2to1219_and0 ^ f_arrdiv16_mux2to1219_and1;
  assign f_arrdiv16_mux2to1220_and0 = f_arrdiv16_mux2to1204_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1220_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1220_and1 = f_arrdiv16_fs234_xor1 & f_arrdiv16_mux2to1220_not0;
  assign f_arrdiv16_mux2to1220_xor0 = f_arrdiv16_mux2to1220_and0 ^ f_arrdiv16_mux2to1220_and1;
  assign f_arrdiv16_mux2to1221_and0 = f_arrdiv16_mux2to1205_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1221_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1221_and1 = f_arrdiv16_fs235_xor1 & f_arrdiv16_mux2to1221_not0;
  assign f_arrdiv16_mux2to1221_xor0 = f_arrdiv16_mux2to1221_and0 ^ f_arrdiv16_mux2to1221_and1;
  assign f_arrdiv16_mux2to1222_and0 = f_arrdiv16_mux2to1206_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1222_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1222_and1 = f_arrdiv16_fs236_xor1 & f_arrdiv16_mux2to1222_not0;
  assign f_arrdiv16_mux2to1222_xor0 = f_arrdiv16_mux2to1222_and0 ^ f_arrdiv16_mux2to1222_and1;
  assign f_arrdiv16_mux2to1223_and0 = f_arrdiv16_mux2to1207_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1223_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1223_and1 = f_arrdiv16_fs237_xor1 & f_arrdiv16_mux2to1223_not0;
  assign f_arrdiv16_mux2to1223_xor0 = f_arrdiv16_mux2to1223_and0 ^ f_arrdiv16_mux2to1223_and1;
  assign f_arrdiv16_mux2to1224_and0 = f_arrdiv16_mux2to1208_xor0 & f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1224_not0 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_mux2to1224_and1 = f_arrdiv16_fs238_xor1 & f_arrdiv16_mux2to1224_not0;
  assign f_arrdiv16_mux2to1224_xor0 = f_arrdiv16_mux2to1224_and0 ^ f_arrdiv16_mux2to1224_and1;
  assign f_arrdiv16_not14 = ~f_arrdiv16_fs239_or0;
  assign f_arrdiv16_fs240_xor0 = a[0] ^ b[0];
  assign f_arrdiv16_fs240_not0 = ~a[0];
  assign f_arrdiv16_fs240_and0 = f_arrdiv16_fs240_not0 & b[0];
  assign f_arrdiv16_fs240_not1 = ~f_arrdiv16_fs240_xor0;
  assign f_arrdiv16_fs241_xor0 = f_arrdiv16_mux2to1210_xor0 ^ b[1];
  assign f_arrdiv16_fs241_not0 = ~f_arrdiv16_mux2to1210_xor0;
  assign f_arrdiv16_fs241_and0 = f_arrdiv16_fs241_not0 & b[1];
  assign f_arrdiv16_fs241_xor1 = f_arrdiv16_fs240_and0 ^ f_arrdiv16_fs241_xor0;
  assign f_arrdiv16_fs241_not1 = ~f_arrdiv16_fs241_xor0;
  assign f_arrdiv16_fs241_and1 = f_arrdiv16_fs241_not1 & f_arrdiv16_fs240_and0;
  assign f_arrdiv16_fs241_or0 = f_arrdiv16_fs241_and1 | f_arrdiv16_fs241_and0;
  assign f_arrdiv16_fs242_xor0 = f_arrdiv16_mux2to1211_xor0 ^ b[2];
  assign f_arrdiv16_fs242_not0 = ~f_arrdiv16_mux2to1211_xor0;
  assign f_arrdiv16_fs242_and0 = f_arrdiv16_fs242_not0 & b[2];
  assign f_arrdiv16_fs242_xor1 = f_arrdiv16_fs241_or0 ^ f_arrdiv16_fs242_xor0;
  assign f_arrdiv16_fs242_not1 = ~f_arrdiv16_fs242_xor0;
  assign f_arrdiv16_fs242_and1 = f_arrdiv16_fs242_not1 & f_arrdiv16_fs241_or0;
  assign f_arrdiv16_fs242_or0 = f_arrdiv16_fs242_and1 | f_arrdiv16_fs242_and0;
  assign f_arrdiv16_fs243_xor0 = f_arrdiv16_mux2to1212_xor0 ^ b[3];
  assign f_arrdiv16_fs243_not0 = ~f_arrdiv16_mux2to1212_xor0;
  assign f_arrdiv16_fs243_and0 = f_arrdiv16_fs243_not0 & b[3];
  assign f_arrdiv16_fs243_xor1 = f_arrdiv16_fs242_or0 ^ f_arrdiv16_fs243_xor0;
  assign f_arrdiv16_fs243_not1 = ~f_arrdiv16_fs243_xor0;
  assign f_arrdiv16_fs243_and1 = f_arrdiv16_fs243_not1 & f_arrdiv16_fs242_or0;
  assign f_arrdiv16_fs243_or0 = f_arrdiv16_fs243_and1 | f_arrdiv16_fs243_and0;
  assign f_arrdiv16_fs244_xor0 = f_arrdiv16_mux2to1213_xor0 ^ b[4];
  assign f_arrdiv16_fs244_not0 = ~f_arrdiv16_mux2to1213_xor0;
  assign f_arrdiv16_fs244_and0 = f_arrdiv16_fs244_not0 & b[4];
  assign f_arrdiv16_fs244_xor1 = f_arrdiv16_fs243_or0 ^ f_arrdiv16_fs244_xor0;
  assign f_arrdiv16_fs244_not1 = ~f_arrdiv16_fs244_xor0;
  assign f_arrdiv16_fs244_and1 = f_arrdiv16_fs244_not1 & f_arrdiv16_fs243_or0;
  assign f_arrdiv16_fs244_or0 = f_arrdiv16_fs244_and1 | f_arrdiv16_fs244_and0;
  assign f_arrdiv16_fs245_xor0 = f_arrdiv16_mux2to1214_xor0 ^ b[5];
  assign f_arrdiv16_fs245_not0 = ~f_arrdiv16_mux2to1214_xor0;
  assign f_arrdiv16_fs245_and0 = f_arrdiv16_fs245_not0 & b[5];
  assign f_arrdiv16_fs245_xor1 = f_arrdiv16_fs244_or0 ^ f_arrdiv16_fs245_xor0;
  assign f_arrdiv16_fs245_not1 = ~f_arrdiv16_fs245_xor0;
  assign f_arrdiv16_fs245_and1 = f_arrdiv16_fs245_not1 & f_arrdiv16_fs244_or0;
  assign f_arrdiv16_fs245_or0 = f_arrdiv16_fs245_and1 | f_arrdiv16_fs245_and0;
  assign f_arrdiv16_fs246_xor0 = f_arrdiv16_mux2to1215_xor0 ^ b[6];
  assign f_arrdiv16_fs246_not0 = ~f_arrdiv16_mux2to1215_xor0;
  assign f_arrdiv16_fs246_and0 = f_arrdiv16_fs246_not0 & b[6];
  assign f_arrdiv16_fs246_xor1 = f_arrdiv16_fs245_or0 ^ f_arrdiv16_fs246_xor0;
  assign f_arrdiv16_fs246_not1 = ~f_arrdiv16_fs246_xor0;
  assign f_arrdiv16_fs246_and1 = f_arrdiv16_fs246_not1 & f_arrdiv16_fs245_or0;
  assign f_arrdiv16_fs246_or0 = f_arrdiv16_fs246_and1 | f_arrdiv16_fs246_and0;
  assign f_arrdiv16_fs247_xor0 = f_arrdiv16_mux2to1216_xor0 ^ b[7];
  assign f_arrdiv16_fs247_not0 = ~f_arrdiv16_mux2to1216_xor0;
  assign f_arrdiv16_fs247_and0 = f_arrdiv16_fs247_not0 & b[7];
  assign f_arrdiv16_fs247_xor1 = f_arrdiv16_fs246_or0 ^ f_arrdiv16_fs247_xor0;
  assign f_arrdiv16_fs247_not1 = ~f_arrdiv16_fs247_xor0;
  assign f_arrdiv16_fs247_and1 = f_arrdiv16_fs247_not1 & f_arrdiv16_fs246_or0;
  assign f_arrdiv16_fs247_or0 = f_arrdiv16_fs247_and1 | f_arrdiv16_fs247_and0;
  assign f_arrdiv16_fs248_xor0 = f_arrdiv16_mux2to1217_xor0 ^ b[8];
  assign f_arrdiv16_fs248_not0 = ~f_arrdiv16_mux2to1217_xor0;
  assign f_arrdiv16_fs248_and0 = f_arrdiv16_fs248_not0 & b[8];
  assign f_arrdiv16_fs248_xor1 = f_arrdiv16_fs247_or0 ^ f_arrdiv16_fs248_xor0;
  assign f_arrdiv16_fs248_not1 = ~f_arrdiv16_fs248_xor0;
  assign f_arrdiv16_fs248_and1 = f_arrdiv16_fs248_not1 & f_arrdiv16_fs247_or0;
  assign f_arrdiv16_fs248_or0 = f_arrdiv16_fs248_and1 | f_arrdiv16_fs248_and0;
  assign f_arrdiv16_fs249_xor0 = f_arrdiv16_mux2to1218_xor0 ^ b[9];
  assign f_arrdiv16_fs249_not0 = ~f_arrdiv16_mux2to1218_xor0;
  assign f_arrdiv16_fs249_and0 = f_arrdiv16_fs249_not0 & b[9];
  assign f_arrdiv16_fs249_xor1 = f_arrdiv16_fs248_or0 ^ f_arrdiv16_fs249_xor0;
  assign f_arrdiv16_fs249_not1 = ~f_arrdiv16_fs249_xor0;
  assign f_arrdiv16_fs249_and1 = f_arrdiv16_fs249_not1 & f_arrdiv16_fs248_or0;
  assign f_arrdiv16_fs249_or0 = f_arrdiv16_fs249_and1 | f_arrdiv16_fs249_and0;
  assign f_arrdiv16_fs250_xor0 = f_arrdiv16_mux2to1219_xor0 ^ b[10];
  assign f_arrdiv16_fs250_not0 = ~f_arrdiv16_mux2to1219_xor0;
  assign f_arrdiv16_fs250_and0 = f_arrdiv16_fs250_not0 & b[10];
  assign f_arrdiv16_fs250_xor1 = f_arrdiv16_fs249_or0 ^ f_arrdiv16_fs250_xor0;
  assign f_arrdiv16_fs250_not1 = ~f_arrdiv16_fs250_xor0;
  assign f_arrdiv16_fs250_and1 = f_arrdiv16_fs250_not1 & f_arrdiv16_fs249_or0;
  assign f_arrdiv16_fs250_or0 = f_arrdiv16_fs250_and1 | f_arrdiv16_fs250_and0;
  assign f_arrdiv16_fs251_xor0 = f_arrdiv16_mux2to1220_xor0 ^ b[11];
  assign f_arrdiv16_fs251_not0 = ~f_arrdiv16_mux2to1220_xor0;
  assign f_arrdiv16_fs251_and0 = f_arrdiv16_fs251_not0 & b[11];
  assign f_arrdiv16_fs251_xor1 = f_arrdiv16_fs250_or0 ^ f_arrdiv16_fs251_xor0;
  assign f_arrdiv16_fs251_not1 = ~f_arrdiv16_fs251_xor0;
  assign f_arrdiv16_fs251_and1 = f_arrdiv16_fs251_not1 & f_arrdiv16_fs250_or0;
  assign f_arrdiv16_fs251_or0 = f_arrdiv16_fs251_and1 | f_arrdiv16_fs251_and0;
  assign f_arrdiv16_fs252_xor0 = f_arrdiv16_mux2to1221_xor0 ^ b[12];
  assign f_arrdiv16_fs252_not0 = ~f_arrdiv16_mux2to1221_xor0;
  assign f_arrdiv16_fs252_and0 = f_arrdiv16_fs252_not0 & b[12];
  assign f_arrdiv16_fs252_xor1 = f_arrdiv16_fs251_or0 ^ f_arrdiv16_fs252_xor0;
  assign f_arrdiv16_fs252_not1 = ~f_arrdiv16_fs252_xor0;
  assign f_arrdiv16_fs252_and1 = f_arrdiv16_fs252_not1 & f_arrdiv16_fs251_or0;
  assign f_arrdiv16_fs252_or0 = f_arrdiv16_fs252_and1 | f_arrdiv16_fs252_and0;
  assign f_arrdiv16_fs253_xor0 = f_arrdiv16_mux2to1222_xor0 ^ b[13];
  assign f_arrdiv16_fs253_not0 = ~f_arrdiv16_mux2to1222_xor0;
  assign f_arrdiv16_fs253_and0 = f_arrdiv16_fs253_not0 & b[13];
  assign f_arrdiv16_fs253_xor1 = f_arrdiv16_fs252_or0 ^ f_arrdiv16_fs253_xor0;
  assign f_arrdiv16_fs253_not1 = ~f_arrdiv16_fs253_xor0;
  assign f_arrdiv16_fs253_and1 = f_arrdiv16_fs253_not1 & f_arrdiv16_fs252_or0;
  assign f_arrdiv16_fs253_or0 = f_arrdiv16_fs253_and1 | f_arrdiv16_fs253_and0;
  assign f_arrdiv16_fs254_xor0 = f_arrdiv16_mux2to1223_xor0 ^ b[14];
  assign f_arrdiv16_fs254_not0 = ~f_arrdiv16_mux2to1223_xor0;
  assign f_arrdiv16_fs254_and0 = f_arrdiv16_fs254_not0 & b[14];
  assign f_arrdiv16_fs254_xor1 = f_arrdiv16_fs253_or0 ^ f_arrdiv16_fs254_xor0;
  assign f_arrdiv16_fs254_not1 = ~f_arrdiv16_fs254_xor0;
  assign f_arrdiv16_fs254_and1 = f_arrdiv16_fs254_not1 & f_arrdiv16_fs253_or0;
  assign f_arrdiv16_fs254_or0 = f_arrdiv16_fs254_and1 | f_arrdiv16_fs254_and0;
  assign f_arrdiv16_fs255_xor0 = f_arrdiv16_mux2to1224_xor0 ^ b[15];
  assign f_arrdiv16_fs255_not0 = ~f_arrdiv16_mux2to1224_xor0;
  assign f_arrdiv16_fs255_and0 = f_arrdiv16_fs255_not0 & b[15];
  assign f_arrdiv16_fs255_xor1 = f_arrdiv16_fs254_or0 ^ f_arrdiv16_fs255_xor0;
  assign f_arrdiv16_fs255_not1 = ~f_arrdiv16_fs255_xor0;
  assign f_arrdiv16_fs255_and1 = f_arrdiv16_fs255_not1 & f_arrdiv16_fs254_or0;
  assign f_arrdiv16_fs255_or0 = f_arrdiv16_fs255_and1 | f_arrdiv16_fs255_and0;
  assign f_arrdiv16_not15 = ~f_arrdiv16_fs255_or0;

  assign f_arrdiv16_out[0] = f_arrdiv16_not15;
  assign f_arrdiv16_out[1] = f_arrdiv16_not14;
  assign f_arrdiv16_out[2] = f_arrdiv16_not13;
  assign f_arrdiv16_out[3] = f_arrdiv16_not12;
  assign f_arrdiv16_out[4] = f_arrdiv16_not11;
  assign f_arrdiv16_out[5] = f_arrdiv16_not10;
  assign f_arrdiv16_out[6] = f_arrdiv16_not9;
  assign f_arrdiv16_out[7] = f_arrdiv16_not8;
  assign f_arrdiv16_out[8] = f_arrdiv16_not7;
  assign f_arrdiv16_out[9] = f_arrdiv16_not6;
  assign f_arrdiv16_out[10] = f_arrdiv16_not5;
  assign f_arrdiv16_out[11] = f_arrdiv16_not4;
  assign f_arrdiv16_out[12] = f_arrdiv16_not3;
  assign f_arrdiv16_out[13] = f_arrdiv16_not2;
  assign f_arrdiv16_out[14] = f_arrdiv16_not1;
  assign f_arrdiv16_out[15] = f_arrdiv16_not0;
endmodule