module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module u_cska62(input [61:0] a, input [61:0] b, output [62:0] u_cska62_out);
  wire [0:0] u_cska62_xor0;
  wire [0:0] u_cska62_ha0_xor0;
  wire [0:0] u_cska62_ha0_and0;
  wire [0:0] u_cska62_xor1;
  wire [0:0] u_cska62_fa0_xor1;
  wire [0:0] u_cska62_fa0_or0;
  wire [0:0] u_cska62_xor2;
  wire [0:0] u_cska62_fa1_xor1;
  wire [0:0] u_cska62_fa1_or0;
  wire [0:0] u_cska62_xor3;
  wire [0:0] u_cska62_fa2_xor1;
  wire [0:0] u_cska62_fa2_or0;
  wire [0:0] u_cska62_and_propagate00;
  wire [0:0] u_cska62_and_propagate01;
  wire [0:0] u_cska62_and_propagate02;
  wire [0:0] u_cska62_mux2to10_and1;
  wire [0:0] u_cska62_xor4;
  wire [0:0] u_cska62_fa3_xor1;
  wire [0:0] u_cska62_fa3_or0;
  wire [0:0] u_cska62_xor5;
  wire [0:0] u_cska62_fa4_xor1;
  wire [0:0] u_cska62_fa4_or0;
  wire [0:0] u_cska62_xor6;
  wire [0:0] u_cska62_fa5_xor1;
  wire [0:0] u_cska62_fa5_or0;
  wire [0:0] u_cska62_xor7;
  wire [0:0] u_cska62_fa6_xor1;
  wire [0:0] u_cska62_fa6_or0;
  wire [0:0] u_cska62_and_propagate13;
  wire [0:0] u_cska62_and_propagate14;
  wire [0:0] u_cska62_and_propagate15;
  wire [0:0] u_cska62_mux2to11_xor0;
  wire [0:0] u_cska62_xor8;
  wire [0:0] u_cska62_fa7_xor1;
  wire [0:0] u_cska62_fa7_or0;
  wire [0:0] u_cska62_xor9;
  wire [0:0] u_cska62_fa8_xor1;
  wire [0:0] u_cska62_fa8_or0;
  wire [0:0] u_cska62_xor10;
  wire [0:0] u_cska62_fa9_xor1;
  wire [0:0] u_cska62_fa9_or0;
  wire [0:0] u_cska62_xor11;
  wire [0:0] u_cska62_fa10_xor1;
  wire [0:0] u_cska62_fa10_or0;
  wire [0:0] u_cska62_and_propagate26;
  wire [0:0] u_cska62_and_propagate27;
  wire [0:0] u_cska62_and_propagate28;
  wire [0:0] u_cska62_mux2to12_xor0;
  wire [0:0] u_cska62_xor12;
  wire [0:0] u_cska62_fa11_xor1;
  wire [0:0] u_cska62_fa11_or0;
  wire [0:0] u_cska62_xor13;
  wire [0:0] u_cska62_fa12_xor1;
  wire [0:0] u_cska62_fa12_or0;
  wire [0:0] u_cska62_xor14;
  wire [0:0] u_cska62_fa13_xor1;
  wire [0:0] u_cska62_fa13_or0;
  wire [0:0] u_cska62_xor15;
  wire [0:0] u_cska62_fa14_xor1;
  wire [0:0] u_cska62_fa14_or0;
  wire [0:0] u_cska62_and_propagate39;
  wire [0:0] u_cska62_and_propagate310;
  wire [0:0] u_cska62_and_propagate311;
  wire [0:0] u_cska62_mux2to13_xor0;
  wire [0:0] u_cska62_xor16;
  wire [0:0] u_cska62_fa15_xor1;
  wire [0:0] u_cska62_fa15_or0;
  wire [0:0] u_cska62_xor17;
  wire [0:0] u_cska62_fa16_xor1;
  wire [0:0] u_cska62_fa16_or0;
  wire [0:0] u_cska62_xor18;
  wire [0:0] u_cska62_fa17_xor1;
  wire [0:0] u_cska62_fa17_or0;
  wire [0:0] u_cska62_xor19;
  wire [0:0] u_cska62_fa18_xor1;
  wire [0:0] u_cska62_fa18_or0;
  wire [0:0] u_cska62_and_propagate412;
  wire [0:0] u_cska62_and_propagate413;
  wire [0:0] u_cska62_and_propagate414;
  wire [0:0] u_cska62_mux2to14_xor0;
  wire [0:0] u_cska62_xor20;
  wire [0:0] u_cska62_fa19_xor1;
  wire [0:0] u_cska62_fa19_or0;
  wire [0:0] u_cska62_xor21;
  wire [0:0] u_cska62_fa20_xor1;
  wire [0:0] u_cska62_fa20_or0;
  wire [0:0] u_cska62_xor22;
  wire [0:0] u_cska62_fa21_xor1;
  wire [0:0] u_cska62_fa21_or0;
  wire [0:0] u_cska62_xor23;
  wire [0:0] u_cska62_fa22_xor1;
  wire [0:0] u_cska62_fa22_or0;
  wire [0:0] u_cska62_and_propagate515;
  wire [0:0] u_cska62_and_propagate516;
  wire [0:0] u_cska62_and_propagate517;
  wire [0:0] u_cska62_mux2to15_xor0;
  wire [0:0] u_cska62_xor24;
  wire [0:0] u_cska62_fa23_xor1;
  wire [0:0] u_cska62_fa23_or0;
  wire [0:0] u_cska62_xor25;
  wire [0:0] u_cska62_fa24_xor1;
  wire [0:0] u_cska62_fa24_or0;
  wire [0:0] u_cska62_xor26;
  wire [0:0] u_cska62_fa25_xor1;
  wire [0:0] u_cska62_fa25_or0;
  wire [0:0] u_cska62_xor27;
  wire [0:0] u_cska62_fa26_xor1;
  wire [0:0] u_cska62_fa26_or0;
  wire [0:0] u_cska62_and_propagate618;
  wire [0:0] u_cska62_and_propagate619;
  wire [0:0] u_cska62_and_propagate620;
  wire [0:0] u_cska62_mux2to16_xor0;
  wire [0:0] u_cska62_xor28;
  wire [0:0] u_cska62_fa27_xor1;
  wire [0:0] u_cska62_fa27_or0;
  wire [0:0] u_cska62_xor29;
  wire [0:0] u_cska62_fa28_xor1;
  wire [0:0] u_cska62_fa28_or0;
  wire [0:0] u_cska62_xor30;
  wire [0:0] u_cska62_fa29_xor1;
  wire [0:0] u_cska62_fa29_or0;
  wire [0:0] u_cska62_xor31;
  wire [0:0] u_cska62_fa30_xor1;
  wire [0:0] u_cska62_fa30_or0;
  wire [0:0] u_cska62_and_propagate721;
  wire [0:0] u_cska62_and_propagate722;
  wire [0:0] u_cska62_and_propagate723;
  wire [0:0] u_cska62_mux2to17_xor0;
  wire [0:0] u_cska62_xor32;
  wire [0:0] u_cska62_fa31_xor1;
  wire [0:0] u_cska62_fa31_or0;
  wire [0:0] u_cska62_xor33;
  wire [0:0] u_cska62_fa32_xor1;
  wire [0:0] u_cska62_fa32_or0;
  wire [0:0] u_cska62_xor34;
  wire [0:0] u_cska62_fa33_xor1;
  wire [0:0] u_cska62_fa33_or0;
  wire [0:0] u_cska62_xor35;
  wire [0:0] u_cska62_fa34_xor1;
  wire [0:0] u_cska62_fa34_or0;
  wire [0:0] u_cska62_and_propagate824;
  wire [0:0] u_cska62_and_propagate825;
  wire [0:0] u_cska62_and_propagate826;
  wire [0:0] u_cska62_mux2to18_xor0;
  wire [0:0] u_cska62_xor36;
  wire [0:0] u_cska62_fa35_xor1;
  wire [0:0] u_cska62_fa35_or0;
  wire [0:0] u_cska62_xor37;
  wire [0:0] u_cska62_fa36_xor1;
  wire [0:0] u_cska62_fa36_or0;
  wire [0:0] u_cska62_xor38;
  wire [0:0] u_cska62_fa37_xor1;
  wire [0:0] u_cska62_fa37_or0;
  wire [0:0] u_cska62_xor39;
  wire [0:0] u_cska62_fa38_xor1;
  wire [0:0] u_cska62_fa38_or0;
  wire [0:0] u_cska62_and_propagate927;
  wire [0:0] u_cska62_and_propagate928;
  wire [0:0] u_cska62_and_propagate929;
  wire [0:0] u_cska62_mux2to19_xor0;
  wire [0:0] u_cska62_xor40;
  wire [0:0] u_cska62_fa39_xor1;
  wire [0:0] u_cska62_fa39_or0;
  wire [0:0] u_cska62_xor41;
  wire [0:0] u_cska62_fa40_xor1;
  wire [0:0] u_cska62_fa40_or0;
  wire [0:0] u_cska62_xor42;
  wire [0:0] u_cska62_fa41_xor1;
  wire [0:0] u_cska62_fa41_or0;
  wire [0:0] u_cska62_xor43;
  wire [0:0] u_cska62_fa42_xor1;
  wire [0:0] u_cska62_fa42_or0;
  wire [0:0] u_cska62_and_propagate1030;
  wire [0:0] u_cska62_and_propagate1031;
  wire [0:0] u_cska62_and_propagate1032;
  wire [0:0] u_cska62_mux2to110_xor0;
  wire [0:0] u_cska62_xor44;
  wire [0:0] u_cska62_fa43_xor1;
  wire [0:0] u_cska62_fa43_or0;
  wire [0:0] u_cska62_xor45;
  wire [0:0] u_cska62_fa44_xor1;
  wire [0:0] u_cska62_fa44_or0;
  wire [0:0] u_cska62_xor46;
  wire [0:0] u_cska62_fa45_xor1;
  wire [0:0] u_cska62_fa45_or0;
  wire [0:0] u_cska62_xor47;
  wire [0:0] u_cska62_fa46_xor1;
  wire [0:0] u_cska62_fa46_or0;
  wire [0:0] u_cska62_and_propagate1133;
  wire [0:0] u_cska62_and_propagate1134;
  wire [0:0] u_cska62_and_propagate1135;
  wire [0:0] u_cska62_mux2to111_xor0;
  wire [0:0] u_cska62_xor48;
  wire [0:0] u_cska62_fa47_xor1;
  wire [0:0] u_cska62_fa47_or0;
  wire [0:0] u_cska62_xor49;
  wire [0:0] u_cska62_fa48_xor1;
  wire [0:0] u_cska62_fa48_or0;
  wire [0:0] u_cska62_xor50;
  wire [0:0] u_cska62_fa49_xor1;
  wire [0:0] u_cska62_fa49_or0;
  wire [0:0] u_cska62_xor51;
  wire [0:0] u_cska62_fa50_xor1;
  wire [0:0] u_cska62_fa50_or0;
  wire [0:0] u_cska62_and_propagate1236;
  wire [0:0] u_cska62_and_propagate1237;
  wire [0:0] u_cska62_and_propagate1238;
  wire [0:0] u_cska62_mux2to112_xor0;
  wire [0:0] u_cska62_xor52;
  wire [0:0] u_cska62_fa51_xor1;
  wire [0:0] u_cska62_fa51_or0;
  wire [0:0] u_cska62_xor53;
  wire [0:0] u_cska62_fa52_xor1;
  wire [0:0] u_cska62_fa52_or0;
  wire [0:0] u_cska62_xor54;
  wire [0:0] u_cska62_fa53_xor1;
  wire [0:0] u_cska62_fa53_or0;
  wire [0:0] u_cska62_xor55;
  wire [0:0] u_cska62_fa54_xor1;
  wire [0:0] u_cska62_fa54_or0;
  wire [0:0] u_cska62_and_propagate1339;
  wire [0:0] u_cska62_and_propagate1340;
  wire [0:0] u_cska62_and_propagate1341;
  wire [0:0] u_cska62_mux2to113_xor0;
  wire [0:0] u_cska62_xor56;
  wire [0:0] u_cska62_fa55_xor1;
  wire [0:0] u_cska62_fa55_or0;
  wire [0:0] u_cska62_xor57;
  wire [0:0] u_cska62_fa56_xor1;
  wire [0:0] u_cska62_fa56_or0;
  wire [0:0] u_cska62_xor58;
  wire [0:0] u_cska62_fa57_xor1;
  wire [0:0] u_cska62_fa57_or0;
  wire [0:0] u_cska62_xor59;
  wire [0:0] u_cska62_fa58_xor1;
  wire [0:0] u_cska62_fa58_or0;
  wire [0:0] u_cska62_and_propagate1442;
  wire [0:0] u_cska62_and_propagate1443;
  wire [0:0] u_cska62_and_propagate1444;
  wire [0:0] u_cska62_mux2to114_xor0;
  wire [0:0] u_cska62_xor60;
  wire [0:0] u_cska62_fa59_xor1;
  wire [0:0] u_cska62_fa59_or0;
  wire [0:0] u_cska62_xor61;
  wire [0:0] u_cska62_fa60_xor1;
  wire [0:0] u_cska62_fa60_or0;
  wire [0:0] u_cska62_and_propagate1545;
  wire [0:0] u_cska62_mux2to115_xor0;

  xor_gate xor_gate_u_cska62_xor0(.a(a[0]), .b(b[0]), .out(u_cska62_xor0));
  ha ha_u_cska62_ha0_out(.a(a[0]), .b(b[0]), .ha_xor0(u_cska62_ha0_xor0), .ha_and0(u_cska62_ha0_and0));
  xor_gate xor_gate_u_cska62_xor1(.a(a[1]), .b(b[1]), .out(u_cska62_xor1));
  fa fa_u_cska62_fa0_out(.a(a[1]), .b(b[1]), .cin(u_cska62_ha0_and0[0]), .fa_xor1(u_cska62_fa0_xor1), .fa_or0(u_cska62_fa0_or0));
  xor_gate xor_gate_u_cska62_xor2(.a(a[2]), .b(b[2]), .out(u_cska62_xor2));
  fa fa_u_cska62_fa1_out(.a(a[2]), .b(b[2]), .cin(u_cska62_fa0_or0[0]), .fa_xor1(u_cska62_fa1_xor1), .fa_or0(u_cska62_fa1_or0));
  xor_gate xor_gate_u_cska62_xor3(.a(a[3]), .b(b[3]), .out(u_cska62_xor3));
  fa fa_u_cska62_fa2_out(.a(a[3]), .b(b[3]), .cin(u_cska62_fa1_or0[0]), .fa_xor1(u_cska62_fa2_xor1), .fa_or0(u_cska62_fa2_or0));
  and_gate and_gate_u_cska62_and_propagate00(.a(u_cska62_xor0[0]), .b(u_cska62_xor2[0]), .out(u_cska62_and_propagate00));
  and_gate and_gate_u_cska62_and_propagate01(.a(u_cska62_xor1[0]), .b(u_cska62_xor3[0]), .out(u_cska62_and_propagate01));
  and_gate and_gate_u_cska62_and_propagate02(.a(u_cska62_and_propagate00[0]), .b(u_cska62_and_propagate01[0]), .out(u_cska62_and_propagate02));
  mux2to1 mux2to1_u_cska62_mux2to10_out(.d0(u_cska62_fa2_or0[0]), .d1(1'b0), .sel(u_cska62_and_propagate02[0]), .mux2to1_xor0(u_cska62_mux2to10_and1));
  xor_gate xor_gate_u_cska62_xor4(.a(a[4]), .b(b[4]), .out(u_cska62_xor4));
  fa fa_u_cska62_fa3_out(.a(a[4]), .b(b[4]), .cin(u_cska62_mux2to10_and1[0]), .fa_xor1(u_cska62_fa3_xor1), .fa_or0(u_cska62_fa3_or0));
  xor_gate xor_gate_u_cska62_xor5(.a(a[5]), .b(b[5]), .out(u_cska62_xor5));
  fa fa_u_cska62_fa4_out(.a(a[5]), .b(b[5]), .cin(u_cska62_fa3_or0[0]), .fa_xor1(u_cska62_fa4_xor1), .fa_or0(u_cska62_fa4_or0));
  xor_gate xor_gate_u_cska62_xor6(.a(a[6]), .b(b[6]), .out(u_cska62_xor6));
  fa fa_u_cska62_fa5_out(.a(a[6]), .b(b[6]), .cin(u_cska62_fa4_or0[0]), .fa_xor1(u_cska62_fa5_xor1), .fa_or0(u_cska62_fa5_or0));
  xor_gate xor_gate_u_cska62_xor7(.a(a[7]), .b(b[7]), .out(u_cska62_xor7));
  fa fa_u_cska62_fa6_out(.a(a[7]), .b(b[7]), .cin(u_cska62_fa5_or0[0]), .fa_xor1(u_cska62_fa6_xor1), .fa_or0(u_cska62_fa6_or0));
  and_gate and_gate_u_cska62_and_propagate13(.a(u_cska62_xor4[0]), .b(u_cska62_xor6[0]), .out(u_cska62_and_propagate13));
  and_gate and_gate_u_cska62_and_propagate14(.a(u_cska62_xor5[0]), .b(u_cska62_xor7[0]), .out(u_cska62_and_propagate14));
  and_gate and_gate_u_cska62_and_propagate15(.a(u_cska62_and_propagate13[0]), .b(u_cska62_and_propagate14[0]), .out(u_cska62_and_propagate15));
  mux2to1 mux2to1_u_cska62_mux2to11_out(.d0(u_cska62_fa6_or0[0]), .d1(u_cska62_mux2to10_and1[0]), .sel(u_cska62_and_propagate15[0]), .mux2to1_xor0(u_cska62_mux2to11_xor0));
  xor_gate xor_gate_u_cska62_xor8(.a(a[8]), .b(b[8]), .out(u_cska62_xor8));
  fa fa_u_cska62_fa7_out(.a(a[8]), .b(b[8]), .cin(u_cska62_mux2to11_xor0[0]), .fa_xor1(u_cska62_fa7_xor1), .fa_or0(u_cska62_fa7_or0));
  xor_gate xor_gate_u_cska62_xor9(.a(a[9]), .b(b[9]), .out(u_cska62_xor9));
  fa fa_u_cska62_fa8_out(.a(a[9]), .b(b[9]), .cin(u_cska62_fa7_or0[0]), .fa_xor1(u_cska62_fa8_xor1), .fa_or0(u_cska62_fa8_or0));
  xor_gate xor_gate_u_cska62_xor10(.a(a[10]), .b(b[10]), .out(u_cska62_xor10));
  fa fa_u_cska62_fa9_out(.a(a[10]), .b(b[10]), .cin(u_cska62_fa8_or0[0]), .fa_xor1(u_cska62_fa9_xor1), .fa_or0(u_cska62_fa9_or0));
  xor_gate xor_gate_u_cska62_xor11(.a(a[11]), .b(b[11]), .out(u_cska62_xor11));
  fa fa_u_cska62_fa10_out(.a(a[11]), .b(b[11]), .cin(u_cska62_fa9_or0[0]), .fa_xor1(u_cska62_fa10_xor1), .fa_or0(u_cska62_fa10_or0));
  and_gate and_gate_u_cska62_and_propagate26(.a(u_cska62_xor8[0]), .b(u_cska62_xor10[0]), .out(u_cska62_and_propagate26));
  and_gate and_gate_u_cska62_and_propagate27(.a(u_cska62_xor9[0]), .b(u_cska62_xor11[0]), .out(u_cska62_and_propagate27));
  and_gate and_gate_u_cska62_and_propagate28(.a(u_cska62_and_propagate26[0]), .b(u_cska62_and_propagate27[0]), .out(u_cska62_and_propagate28));
  mux2to1 mux2to1_u_cska62_mux2to12_out(.d0(u_cska62_fa10_or0[0]), .d1(u_cska62_mux2to11_xor0[0]), .sel(u_cska62_and_propagate28[0]), .mux2to1_xor0(u_cska62_mux2to12_xor0));
  xor_gate xor_gate_u_cska62_xor12(.a(a[12]), .b(b[12]), .out(u_cska62_xor12));
  fa fa_u_cska62_fa11_out(.a(a[12]), .b(b[12]), .cin(u_cska62_mux2to12_xor0[0]), .fa_xor1(u_cska62_fa11_xor1), .fa_or0(u_cska62_fa11_or0));
  xor_gate xor_gate_u_cska62_xor13(.a(a[13]), .b(b[13]), .out(u_cska62_xor13));
  fa fa_u_cska62_fa12_out(.a(a[13]), .b(b[13]), .cin(u_cska62_fa11_or0[0]), .fa_xor1(u_cska62_fa12_xor1), .fa_or0(u_cska62_fa12_or0));
  xor_gate xor_gate_u_cska62_xor14(.a(a[14]), .b(b[14]), .out(u_cska62_xor14));
  fa fa_u_cska62_fa13_out(.a(a[14]), .b(b[14]), .cin(u_cska62_fa12_or0[0]), .fa_xor1(u_cska62_fa13_xor1), .fa_or0(u_cska62_fa13_or0));
  xor_gate xor_gate_u_cska62_xor15(.a(a[15]), .b(b[15]), .out(u_cska62_xor15));
  fa fa_u_cska62_fa14_out(.a(a[15]), .b(b[15]), .cin(u_cska62_fa13_or0[0]), .fa_xor1(u_cska62_fa14_xor1), .fa_or0(u_cska62_fa14_or0));
  and_gate and_gate_u_cska62_and_propagate39(.a(u_cska62_xor12[0]), .b(u_cska62_xor14[0]), .out(u_cska62_and_propagate39));
  and_gate and_gate_u_cska62_and_propagate310(.a(u_cska62_xor13[0]), .b(u_cska62_xor15[0]), .out(u_cska62_and_propagate310));
  and_gate and_gate_u_cska62_and_propagate311(.a(u_cska62_and_propagate39[0]), .b(u_cska62_and_propagate310[0]), .out(u_cska62_and_propagate311));
  mux2to1 mux2to1_u_cska62_mux2to13_out(.d0(u_cska62_fa14_or0[0]), .d1(u_cska62_mux2to12_xor0[0]), .sel(u_cska62_and_propagate311[0]), .mux2to1_xor0(u_cska62_mux2to13_xor0));
  xor_gate xor_gate_u_cska62_xor16(.a(a[16]), .b(b[16]), .out(u_cska62_xor16));
  fa fa_u_cska62_fa15_out(.a(a[16]), .b(b[16]), .cin(u_cska62_mux2to13_xor0[0]), .fa_xor1(u_cska62_fa15_xor1), .fa_or0(u_cska62_fa15_or0));
  xor_gate xor_gate_u_cska62_xor17(.a(a[17]), .b(b[17]), .out(u_cska62_xor17));
  fa fa_u_cska62_fa16_out(.a(a[17]), .b(b[17]), .cin(u_cska62_fa15_or0[0]), .fa_xor1(u_cska62_fa16_xor1), .fa_or0(u_cska62_fa16_or0));
  xor_gate xor_gate_u_cska62_xor18(.a(a[18]), .b(b[18]), .out(u_cska62_xor18));
  fa fa_u_cska62_fa17_out(.a(a[18]), .b(b[18]), .cin(u_cska62_fa16_or0[0]), .fa_xor1(u_cska62_fa17_xor1), .fa_or0(u_cska62_fa17_or0));
  xor_gate xor_gate_u_cska62_xor19(.a(a[19]), .b(b[19]), .out(u_cska62_xor19));
  fa fa_u_cska62_fa18_out(.a(a[19]), .b(b[19]), .cin(u_cska62_fa17_or0[0]), .fa_xor1(u_cska62_fa18_xor1), .fa_or0(u_cska62_fa18_or0));
  and_gate and_gate_u_cska62_and_propagate412(.a(u_cska62_xor16[0]), .b(u_cska62_xor18[0]), .out(u_cska62_and_propagate412));
  and_gate and_gate_u_cska62_and_propagate413(.a(u_cska62_xor17[0]), .b(u_cska62_xor19[0]), .out(u_cska62_and_propagate413));
  and_gate and_gate_u_cska62_and_propagate414(.a(u_cska62_and_propagate412[0]), .b(u_cska62_and_propagate413[0]), .out(u_cska62_and_propagate414));
  mux2to1 mux2to1_u_cska62_mux2to14_out(.d0(u_cska62_fa18_or0[0]), .d1(u_cska62_mux2to13_xor0[0]), .sel(u_cska62_and_propagate414[0]), .mux2to1_xor0(u_cska62_mux2to14_xor0));
  xor_gate xor_gate_u_cska62_xor20(.a(a[20]), .b(b[20]), .out(u_cska62_xor20));
  fa fa_u_cska62_fa19_out(.a(a[20]), .b(b[20]), .cin(u_cska62_mux2to14_xor0[0]), .fa_xor1(u_cska62_fa19_xor1), .fa_or0(u_cska62_fa19_or0));
  xor_gate xor_gate_u_cska62_xor21(.a(a[21]), .b(b[21]), .out(u_cska62_xor21));
  fa fa_u_cska62_fa20_out(.a(a[21]), .b(b[21]), .cin(u_cska62_fa19_or0[0]), .fa_xor1(u_cska62_fa20_xor1), .fa_or0(u_cska62_fa20_or0));
  xor_gate xor_gate_u_cska62_xor22(.a(a[22]), .b(b[22]), .out(u_cska62_xor22));
  fa fa_u_cska62_fa21_out(.a(a[22]), .b(b[22]), .cin(u_cska62_fa20_or0[0]), .fa_xor1(u_cska62_fa21_xor1), .fa_or0(u_cska62_fa21_or0));
  xor_gate xor_gate_u_cska62_xor23(.a(a[23]), .b(b[23]), .out(u_cska62_xor23));
  fa fa_u_cska62_fa22_out(.a(a[23]), .b(b[23]), .cin(u_cska62_fa21_or0[0]), .fa_xor1(u_cska62_fa22_xor1), .fa_or0(u_cska62_fa22_or0));
  and_gate and_gate_u_cska62_and_propagate515(.a(u_cska62_xor20[0]), .b(u_cska62_xor22[0]), .out(u_cska62_and_propagate515));
  and_gate and_gate_u_cska62_and_propagate516(.a(u_cska62_xor21[0]), .b(u_cska62_xor23[0]), .out(u_cska62_and_propagate516));
  and_gate and_gate_u_cska62_and_propagate517(.a(u_cska62_and_propagate515[0]), .b(u_cska62_and_propagate516[0]), .out(u_cska62_and_propagate517));
  mux2to1 mux2to1_u_cska62_mux2to15_out(.d0(u_cska62_fa22_or0[0]), .d1(u_cska62_mux2to14_xor0[0]), .sel(u_cska62_and_propagate517[0]), .mux2to1_xor0(u_cska62_mux2to15_xor0));
  xor_gate xor_gate_u_cska62_xor24(.a(a[24]), .b(b[24]), .out(u_cska62_xor24));
  fa fa_u_cska62_fa23_out(.a(a[24]), .b(b[24]), .cin(u_cska62_mux2to15_xor0[0]), .fa_xor1(u_cska62_fa23_xor1), .fa_or0(u_cska62_fa23_or0));
  xor_gate xor_gate_u_cska62_xor25(.a(a[25]), .b(b[25]), .out(u_cska62_xor25));
  fa fa_u_cska62_fa24_out(.a(a[25]), .b(b[25]), .cin(u_cska62_fa23_or0[0]), .fa_xor1(u_cska62_fa24_xor1), .fa_or0(u_cska62_fa24_or0));
  xor_gate xor_gate_u_cska62_xor26(.a(a[26]), .b(b[26]), .out(u_cska62_xor26));
  fa fa_u_cska62_fa25_out(.a(a[26]), .b(b[26]), .cin(u_cska62_fa24_or0[0]), .fa_xor1(u_cska62_fa25_xor1), .fa_or0(u_cska62_fa25_or0));
  xor_gate xor_gate_u_cska62_xor27(.a(a[27]), .b(b[27]), .out(u_cska62_xor27));
  fa fa_u_cska62_fa26_out(.a(a[27]), .b(b[27]), .cin(u_cska62_fa25_or0[0]), .fa_xor1(u_cska62_fa26_xor1), .fa_or0(u_cska62_fa26_or0));
  and_gate and_gate_u_cska62_and_propagate618(.a(u_cska62_xor24[0]), .b(u_cska62_xor26[0]), .out(u_cska62_and_propagate618));
  and_gate and_gate_u_cska62_and_propagate619(.a(u_cska62_xor25[0]), .b(u_cska62_xor27[0]), .out(u_cska62_and_propagate619));
  and_gate and_gate_u_cska62_and_propagate620(.a(u_cska62_and_propagate618[0]), .b(u_cska62_and_propagate619[0]), .out(u_cska62_and_propagate620));
  mux2to1 mux2to1_u_cska62_mux2to16_out(.d0(u_cska62_fa26_or0[0]), .d1(u_cska62_mux2to15_xor0[0]), .sel(u_cska62_and_propagate620[0]), .mux2to1_xor0(u_cska62_mux2to16_xor0));
  xor_gate xor_gate_u_cska62_xor28(.a(a[28]), .b(b[28]), .out(u_cska62_xor28));
  fa fa_u_cska62_fa27_out(.a(a[28]), .b(b[28]), .cin(u_cska62_mux2to16_xor0[0]), .fa_xor1(u_cska62_fa27_xor1), .fa_or0(u_cska62_fa27_or0));
  xor_gate xor_gate_u_cska62_xor29(.a(a[29]), .b(b[29]), .out(u_cska62_xor29));
  fa fa_u_cska62_fa28_out(.a(a[29]), .b(b[29]), .cin(u_cska62_fa27_or0[0]), .fa_xor1(u_cska62_fa28_xor1), .fa_or0(u_cska62_fa28_or0));
  xor_gate xor_gate_u_cska62_xor30(.a(a[30]), .b(b[30]), .out(u_cska62_xor30));
  fa fa_u_cska62_fa29_out(.a(a[30]), .b(b[30]), .cin(u_cska62_fa28_or0[0]), .fa_xor1(u_cska62_fa29_xor1), .fa_or0(u_cska62_fa29_or0));
  xor_gate xor_gate_u_cska62_xor31(.a(a[31]), .b(b[31]), .out(u_cska62_xor31));
  fa fa_u_cska62_fa30_out(.a(a[31]), .b(b[31]), .cin(u_cska62_fa29_or0[0]), .fa_xor1(u_cska62_fa30_xor1), .fa_or0(u_cska62_fa30_or0));
  and_gate and_gate_u_cska62_and_propagate721(.a(u_cska62_xor28[0]), .b(u_cska62_xor30[0]), .out(u_cska62_and_propagate721));
  and_gate and_gate_u_cska62_and_propagate722(.a(u_cska62_xor29[0]), .b(u_cska62_xor31[0]), .out(u_cska62_and_propagate722));
  and_gate and_gate_u_cska62_and_propagate723(.a(u_cska62_and_propagate721[0]), .b(u_cska62_and_propagate722[0]), .out(u_cska62_and_propagate723));
  mux2to1 mux2to1_u_cska62_mux2to17_out(.d0(u_cska62_fa30_or0[0]), .d1(u_cska62_mux2to16_xor0[0]), .sel(u_cska62_and_propagate723[0]), .mux2to1_xor0(u_cska62_mux2to17_xor0));
  xor_gate xor_gate_u_cska62_xor32(.a(a[32]), .b(b[32]), .out(u_cska62_xor32));
  fa fa_u_cska62_fa31_out(.a(a[32]), .b(b[32]), .cin(u_cska62_mux2to17_xor0[0]), .fa_xor1(u_cska62_fa31_xor1), .fa_or0(u_cska62_fa31_or0));
  xor_gate xor_gate_u_cska62_xor33(.a(a[33]), .b(b[33]), .out(u_cska62_xor33));
  fa fa_u_cska62_fa32_out(.a(a[33]), .b(b[33]), .cin(u_cska62_fa31_or0[0]), .fa_xor1(u_cska62_fa32_xor1), .fa_or0(u_cska62_fa32_or0));
  xor_gate xor_gate_u_cska62_xor34(.a(a[34]), .b(b[34]), .out(u_cska62_xor34));
  fa fa_u_cska62_fa33_out(.a(a[34]), .b(b[34]), .cin(u_cska62_fa32_or0[0]), .fa_xor1(u_cska62_fa33_xor1), .fa_or0(u_cska62_fa33_or0));
  xor_gate xor_gate_u_cska62_xor35(.a(a[35]), .b(b[35]), .out(u_cska62_xor35));
  fa fa_u_cska62_fa34_out(.a(a[35]), .b(b[35]), .cin(u_cska62_fa33_or0[0]), .fa_xor1(u_cska62_fa34_xor1), .fa_or0(u_cska62_fa34_or0));
  and_gate and_gate_u_cska62_and_propagate824(.a(u_cska62_xor32[0]), .b(u_cska62_xor34[0]), .out(u_cska62_and_propagate824));
  and_gate and_gate_u_cska62_and_propagate825(.a(u_cska62_xor33[0]), .b(u_cska62_xor35[0]), .out(u_cska62_and_propagate825));
  and_gate and_gate_u_cska62_and_propagate826(.a(u_cska62_and_propagate824[0]), .b(u_cska62_and_propagate825[0]), .out(u_cska62_and_propagate826));
  mux2to1 mux2to1_u_cska62_mux2to18_out(.d0(u_cska62_fa34_or0[0]), .d1(u_cska62_mux2to17_xor0[0]), .sel(u_cska62_and_propagate826[0]), .mux2to1_xor0(u_cska62_mux2to18_xor0));
  xor_gate xor_gate_u_cska62_xor36(.a(a[36]), .b(b[36]), .out(u_cska62_xor36));
  fa fa_u_cska62_fa35_out(.a(a[36]), .b(b[36]), .cin(u_cska62_mux2to18_xor0[0]), .fa_xor1(u_cska62_fa35_xor1), .fa_or0(u_cska62_fa35_or0));
  xor_gate xor_gate_u_cska62_xor37(.a(a[37]), .b(b[37]), .out(u_cska62_xor37));
  fa fa_u_cska62_fa36_out(.a(a[37]), .b(b[37]), .cin(u_cska62_fa35_or0[0]), .fa_xor1(u_cska62_fa36_xor1), .fa_or0(u_cska62_fa36_or0));
  xor_gate xor_gate_u_cska62_xor38(.a(a[38]), .b(b[38]), .out(u_cska62_xor38));
  fa fa_u_cska62_fa37_out(.a(a[38]), .b(b[38]), .cin(u_cska62_fa36_or0[0]), .fa_xor1(u_cska62_fa37_xor1), .fa_or0(u_cska62_fa37_or0));
  xor_gate xor_gate_u_cska62_xor39(.a(a[39]), .b(b[39]), .out(u_cska62_xor39));
  fa fa_u_cska62_fa38_out(.a(a[39]), .b(b[39]), .cin(u_cska62_fa37_or0[0]), .fa_xor1(u_cska62_fa38_xor1), .fa_or0(u_cska62_fa38_or0));
  and_gate and_gate_u_cska62_and_propagate927(.a(u_cska62_xor36[0]), .b(u_cska62_xor38[0]), .out(u_cska62_and_propagate927));
  and_gate and_gate_u_cska62_and_propagate928(.a(u_cska62_xor37[0]), .b(u_cska62_xor39[0]), .out(u_cska62_and_propagate928));
  and_gate and_gate_u_cska62_and_propagate929(.a(u_cska62_and_propagate927[0]), .b(u_cska62_and_propagate928[0]), .out(u_cska62_and_propagate929));
  mux2to1 mux2to1_u_cska62_mux2to19_out(.d0(u_cska62_fa38_or0[0]), .d1(u_cska62_mux2to18_xor0[0]), .sel(u_cska62_and_propagate929[0]), .mux2to1_xor0(u_cska62_mux2to19_xor0));
  xor_gate xor_gate_u_cska62_xor40(.a(a[40]), .b(b[40]), .out(u_cska62_xor40));
  fa fa_u_cska62_fa39_out(.a(a[40]), .b(b[40]), .cin(u_cska62_mux2to19_xor0[0]), .fa_xor1(u_cska62_fa39_xor1), .fa_or0(u_cska62_fa39_or0));
  xor_gate xor_gate_u_cska62_xor41(.a(a[41]), .b(b[41]), .out(u_cska62_xor41));
  fa fa_u_cska62_fa40_out(.a(a[41]), .b(b[41]), .cin(u_cska62_fa39_or0[0]), .fa_xor1(u_cska62_fa40_xor1), .fa_or0(u_cska62_fa40_or0));
  xor_gate xor_gate_u_cska62_xor42(.a(a[42]), .b(b[42]), .out(u_cska62_xor42));
  fa fa_u_cska62_fa41_out(.a(a[42]), .b(b[42]), .cin(u_cska62_fa40_or0[0]), .fa_xor1(u_cska62_fa41_xor1), .fa_or0(u_cska62_fa41_or0));
  xor_gate xor_gate_u_cska62_xor43(.a(a[43]), .b(b[43]), .out(u_cska62_xor43));
  fa fa_u_cska62_fa42_out(.a(a[43]), .b(b[43]), .cin(u_cska62_fa41_or0[0]), .fa_xor1(u_cska62_fa42_xor1), .fa_or0(u_cska62_fa42_or0));
  and_gate and_gate_u_cska62_and_propagate1030(.a(u_cska62_xor40[0]), .b(u_cska62_xor42[0]), .out(u_cska62_and_propagate1030));
  and_gate and_gate_u_cska62_and_propagate1031(.a(u_cska62_xor41[0]), .b(u_cska62_xor43[0]), .out(u_cska62_and_propagate1031));
  and_gate and_gate_u_cska62_and_propagate1032(.a(u_cska62_and_propagate1030[0]), .b(u_cska62_and_propagate1031[0]), .out(u_cska62_and_propagate1032));
  mux2to1 mux2to1_u_cska62_mux2to110_out(.d0(u_cska62_fa42_or0[0]), .d1(u_cska62_mux2to19_xor0[0]), .sel(u_cska62_and_propagate1032[0]), .mux2to1_xor0(u_cska62_mux2to110_xor0));
  xor_gate xor_gate_u_cska62_xor44(.a(a[44]), .b(b[44]), .out(u_cska62_xor44));
  fa fa_u_cska62_fa43_out(.a(a[44]), .b(b[44]), .cin(u_cska62_mux2to110_xor0[0]), .fa_xor1(u_cska62_fa43_xor1), .fa_or0(u_cska62_fa43_or0));
  xor_gate xor_gate_u_cska62_xor45(.a(a[45]), .b(b[45]), .out(u_cska62_xor45));
  fa fa_u_cska62_fa44_out(.a(a[45]), .b(b[45]), .cin(u_cska62_fa43_or0[0]), .fa_xor1(u_cska62_fa44_xor1), .fa_or0(u_cska62_fa44_or0));
  xor_gate xor_gate_u_cska62_xor46(.a(a[46]), .b(b[46]), .out(u_cska62_xor46));
  fa fa_u_cska62_fa45_out(.a(a[46]), .b(b[46]), .cin(u_cska62_fa44_or0[0]), .fa_xor1(u_cska62_fa45_xor1), .fa_or0(u_cska62_fa45_or0));
  xor_gate xor_gate_u_cska62_xor47(.a(a[47]), .b(b[47]), .out(u_cska62_xor47));
  fa fa_u_cska62_fa46_out(.a(a[47]), .b(b[47]), .cin(u_cska62_fa45_or0[0]), .fa_xor1(u_cska62_fa46_xor1), .fa_or0(u_cska62_fa46_or0));
  and_gate and_gate_u_cska62_and_propagate1133(.a(u_cska62_xor44[0]), .b(u_cska62_xor46[0]), .out(u_cska62_and_propagate1133));
  and_gate and_gate_u_cska62_and_propagate1134(.a(u_cska62_xor45[0]), .b(u_cska62_xor47[0]), .out(u_cska62_and_propagate1134));
  and_gate and_gate_u_cska62_and_propagate1135(.a(u_cska62_and_propagate1133[0]), .b(u_cska62_and_propagate1134[0]), .out(u_cska62_and_propagate1135));
  mux2to1 mux2to1_u_cska62_mux2to111_out(.d0(u_cska62_fa46_or0[0]), .d1(u_cska62_mux2to110_xor0[0]), .sel(u_cska62_and_propagate1135[0]), .mux2to1_xor0(u_cska62_mux2to111_xor0));
  xor_gate xor_gate_u_cska62_xor48(.a(a[48]), .b(b[48]), .out(u_cska62_xor48));
  fa fa_u_cska62_fa47_out(.a(a[48]), .b(b[48]), .cin(u_cska62_mux2to111_xor0[0]), .fa_xor1(u_cska62_fa47_xor1), .fa_or0(u_cska62_fa47_or0));
  xor_gate xor_gate_u_cska62_xor49(.a(a[49]), .b(b[49]), .out(u_cska62_xor49));
  fa fa_u_cska62_fa48_out(.a(a[49]), .b(b[49]), .cin(u_cska62_fa47_or0[0]), .fa_xor1(u_cska62_fa48_xor1), .fa_or0(u_cska62_fa48_or0));
  xor_gate xor_gate_u_cska62_xor50(.a(a[50]), .b(b[50]), .out(u_cska62_xor50));
  fa fa_u_cska62_fa49_out(.a(a[50]), .b(b[50]), .cin(u_cska62_fa48_or0[0]), .fa_xor1(u_cska62_fa49_xor1), .fa_or0(u_cska62_fa49_or0));
  xor_gate xor_gate_u_cska62_xor51(.a(a[51]), .b(b[51]), .out(u_cska62_xor51));
  fa fa_u_cska62_fa50_out(.a(a[51]), .b(b[51]), .cin(u_cska62_fa49_or0[0]), .fa_xor1(u_cska62_fa50_xor1), .fa_or0(u_cska62_fa50_or0));
  and_gate and_gate_u_cska62_and_propagate1236(.a(u_cska62_xor48[0]), .b(u_cska62_xor50[0]), .out(u_cska62_and_propagate1236));
  and_gate and_gate_u_cska62_and_propagate1237(.a(u_cska62_xor49[0]), .b(u_cska62_xor51[0]), .out(u_cska62_and_propagate1237));
  and_gate and_gate_u_cska62_and_propagate1238(.a(u_cska62_and_propagate1236[0]), .b(u_cska62_and_propagate1237[0]), .out(u_cska62_and_propagate1238));
  mux2to1 mux2to1_u_cska62_mux2to112_out(.d0(u_cska62_fa50_or0[0]), .d1(u_cska62_mux2to111_xor0[0]), .sel(u_cska62_and_propagate1238[0]), .mux2to1_xor0(u_cska62_mux2to112_xor0));
  xor_gate xor_gate_u_cska62_xor52(.a(a[52]), .b(b[52]), .out(u_cska62_xor52));
  fa fa_u_cska62_fa51_out(.a(a[52]), .b(b[52]), .cin(u_cska62_mux2to112_xor0[0]), .fa_xor1(u_cska62_fa51_xor1), .fa_or0(u_cska62_fa51_or0));
  xor_gate xor_gate_u_cska62_xor53(.a(a[53]), .b(b[53]), .out(u_cska62_xor53));
  fa fa_u_cska62_fa52_out(.a(a[53]), .b(b[53]), .cin(u_cska62_fa51_or0[0]), .fa_xor1(u_cska62_fa52_xor1), .fa_or0(u_cska62_fa52_or0));
  xor_gate xor_gate_u_cska62_xor54(.a(a[54]), .b(b[54]), .out(u_cska62_xor54));
  fa fa_u_cska62_fa53_out(.a(a[54]), .b(b[54]), .cin(u_cska62_fa52_or0[0]), .fa_xor1(u_cska62_fa53_xor1), .fa_or0(u_cska62_fa53_or0));
  xor_gate xor_gate_u_cska62_xor55(.a(a[55]), .b(b[55]), .out(u_cska62_xor55));
  fa fa_u_cska62_fa54_out(.a(a[55]), .b(b[55]), .cin(u_cska62_fa53_or0[0]), .fa_xor1(u_cska62_fa54_xor1), .fa_or0(u_cska62_fa54_or0));
  and_gate and_gate_u_cska62_and_propagate1339(.a(u_cska62_xor52[0]), .b(u_cska62_xor54[0]), .out(u_cska62_and_propagate1339));
  and_gate and_gate_u_cska62_and_propagate1340(.a(u_cska62_xor53[0]), .b(u_cska62_xor55[0]), .out(u_cska62_and_propagate1340));
  and_gate and_gate_u_cska62_and_propagate1341(.a(u_cska62_and_propagate1339[0]), .b(u_cska62_and_propagate1340[0]), .out(u_cska62_and_propagate1341));
  mux2to1 mux2to1_u_cska62_mux2to113_out(.d0(u_cska62_fa54_or0[0]), .d1(u_cska62_mux2to112_xor0[0]), .sel(u_cska62_and_propagate1341[0]), .mux2to1_xor0(u_cska62_mux2to113_xor0));
  xor_gate xor_gate_u_cska62_xor56(.a(a[56]), .b(b[56]), .out(u_cska62_xor56));
  fa fa_u_cska62_fa55_out(.a(a[56]), .b(b[56]), .cin(u_cska62_mux2to113_xor0[0]), .fa_xor1(u_cska62_fa55_xor1), .fa_or0(u_cska62_fa55_or0));
  xor_gate xor_gate_u_cska62_xor57(.a(a[57]), .b(b[57]), .out(u_cska62_xor57));
  fa fa_u_cska62_fa56_out(.a(a[57]), .b(b[57]), .cin(u_cska62_fa55_or0[0]), .fa_xor1(u_cska62_fa56_xor1), .fa_or0(u_cska62_fa56_or0));
  xor_gate xor_gate_u_cska62_xor58(.a(a[58]), .b(b[58]), .out(u_cska62_xor58));
  fa fa_u_cska62_fa57_out(.a(a[58]), .b(b[58]), .cin(u_cska62_fa56_or0[0]), .fa_xor1(u_cska62_fa57_xor1), .fa_or0(u_cska62_fa57_or0));
  xor_gate xor_gate_u_cska62_xor59(.a(a[59]), .b(b[59]), .out(u_cska62_xor59));
  fa fa_u_cska62_fa58_out(.a(a[59]), .b(b[59]), .cin(u_cska62_fa57_or0[0]), .fa_xor1(u_cska62_fa58_xor1), .fa_or0(u_cska62_fa58_or0));
  and_gate and_gate_u_cska62_and_propagate1442(.a(u_cska62_xor56[0]), .b(u_cska62_xor58[0]), .out(u_cska62_and_propagate1442));
  and_gate and_gate_u_cska62_and_propagate1443(.a(u_cska62_xor57[0]), .b(u_cska62_xor59[0]), .out(u_cska62_and_propagate1443));
  and_gate and_gate_u_cska62_and_propagate1444(.a(u_cska62_and_propagate1442[0]), .b(u_cska62_and_propagate1443[0]), .out(u_cska62_and_propagate1444));
  mux2to1 mux2to1_u_cska62_mux2to114_out(.d0(u_cska62_fa58_or0[0]), .d1(u_cska62_mux2to113_xor0[0]), .sel(u_cska62_and_propagate1444[0]), .mux2to1_xor0(u_cska62_mux2to114_xor0));
  xor_gate xor_gate_u_cska62_xor60(.a(a[60]), .b(b[60]), .out(u_cska62_xor60));
  fa fa_u_cska62_fa59_out(.a(a[60]), .b(b[60]), .cin(u_cska62_mux2to114_xor0[0]), .fa_xor1(u_cska62_fa59_xor1), .fa_or0(u_cska62_fa59_or0));
  xor_gate xor_gate_u_cska62_xor61(.a(a[61]), .b(b[61]), .out(u_cska62_xor61));
  fa fa_u_cska62_fa60_out(.a(a[61]), .b(b[61]), .cin(u_cska62_fa59_or0[0]), .fa_xor1(u_cska62_fa60_xor1), .fa_or0(u_cska62_fa60_or0));
  and_gate and_gate_u_cska62_and_propagate1545(.a(u_cska62_xor60[0]), .b(u_cska62_xor61[0]), .out(u_cska62_and_propagate1545));
  mux2to1 mux2to1_u_cska62_mux2to115_out(.d0(u_cska62_fa60_or0[0]), .d1(u_cska62_mux2to114_xor0[0]), .sel(u_cska62_and_propagate1545[0]), .mux2to1_xor0(u_cska62_mux2to115_xor0));

  assign u_cska62_out[0] = u_cska62_ha0_xor0[0];
  assign u_cska62_out[1] = u_cska62_fa0_xor1[0];
  assign u_cska62_out[2] = u_cska62_fa1_xor1[0];
  assign u_cska62_out[3] = u_cska62_fa2_xor1[0];
  assign u_cska62_out[4] = u_cska62_fa3_xor1[0];
  assign u_cska62_out[5] = u_cska62_fa4_xor1[0];
  assign u_cska62_out[6] = u_cska62_fa5_xor1[0];
  assign u_cska62_out[7] = u_cska62_fa6_xor1[0];
  assign u_cska62_out[8] = u_cska62_fa7_xor1[0];
  assign u_cska62_out[9] = u_cska62_fa8_xor1[0];
  assign u_cska62_out[10] = u_cska62_fa9_xor1[0];
  assign u_cska62_out[11] = u_cska62_fa10_xor1[0];
  assign u_cska62_out[12] = u_cska62_fa11_xor1[0];
  assign u_cska62_out[13] = u_cska62_fa12_xor1[0];
  assign u_cska62_out[14] = u_cska62_fa13_xor1[0];
  assign u_cska62_out[15] = u_cska62_fa14_xor1[0];
  assign u_cska62_out[16] = u_cska62_fa15_xor1[0];
  assign u_cska62_out[17] = u_cska62_fa16_xor1[0];
  assign u_cska62_out[18] = u_cska62_fa17_xor1[0];
  assign u_cska62_out[19] = u_cska62_fa18_xor1[0];
  assign u_cska62_out[20] = u_cska62_fa19_xor1[0];
  assign u_cska62_out[21] = u_cska62_fa20_xor1[0];
  assign u_cska62_out[22] = u_cska62_fa21_xor1[0];
  assign u_cska62_out[23] = u_cska62_fa22_xor1[0];
  assign u_cska62_out[24] = u_cska62_fa23_xor1[0];
  assign u_cska62_out[25] = u_cska62_fa24_xor1[0];
  assign u_cska62_out[26] = u_cska62_fa25_xor1[0];
  assign u_cska62_out[27] = u_cska62_fa26_xor1[0];
  assign u_cska62_out[28] = u_cska62_fa27_xor1[0];
  assign u_cska62_out[29] = u_cska62_fa28_xor1[0];
  assign u_cska62_out[30] = u_cska62_fa29_xor1[0];
  assign u_cska62_out[31] = u_cska62_fa30_xor1[0];
  assign u_cska62_out[32] = u_cska62_fa31_xor1[0];
  assign u_cska62_out[33] = u_cska62_fa32_xor1[0];
  assign u_cska62_out[34] = u_cska62_fa33_xor1[0];
  assign u_cska62_out[35] = u_cska62_fa34_xor1[0];
  assign u_cska62_out[36] = u_cska62_fa35_xor1[0];
  assign u_cska62_out[37] = u_cska62_fa36_xor1[0];
  assign u_cska62_out[38] = u_cska62_fa37_xor1[0];
  assign u_cska62_out[39] = u_cska62_fa38_xor1[0];
  assign u_cska62_out[40] = u_cska62_fa39_xor1[0];
  assign u_cska62_out[41] = u_cska62_fa40_xor1[0];
  assign u_cska62_out[42] = u_cska62_fa41_xor1[0];
  assign u_cska62_out[43] = u_cska62_fa42_xor1[0];
  assign u_cska62_out[44] = u_cska62_fa43_xor1[0];
  assign u_cska62_out[45] = u_cska62_fa44_xor1[0];
  assign u_cska62_out[46] = u_cska62_fa45_xor1[0];
  assign u_cska62_out[47] = u_cska62_fa46_xor1[0];
  assign u_cska62_out[48] = u_cska62_fa47_xor1[0];
  assign u_cska62_out[49] = u_cska62_fa48_xor1[0];
  assign u_cska62_out[50] = u_cska62_fa49_xor1[0];
  assign u_cska62_out[51] = u_cska62_fa50_xor1[0];
  assign u_cska62_out[52] = u_cska62_fa51_xor1[0];
  assign u_cska62_out[53] = u_cska62_fa52_xor1[0];
  assign u_cska62_out[54] = u_cska62_fa53_xor1[0];
  assign u_cska62_out[55] = u_cska62_fa54_xor1[0];
  assign u_cska62_out[56] = u_cska62_fa55_xor1[0];
  assign u_cska62_out[57] = u_cska62_fa56_xor1[0];
  assign u_cska62_out[58] = u_cska62_fa57_xor1[0];
  assign u_cska62_out[59] = u_cska62_fa58_xor1[0];
  assign u_cska62_out[60] = u_cska62_fa59_xor1[0];
  assign u_cska62_out[61] = u_cska62_fa60_xor1[0];
  assign u_cska62_out[62] = u_cska62_mux2to115_xor0[0];
endmodule

module s_wallace_cska32(input [31:0] a, input [31:0] b, output [63:0] s_wallace_cska32_out);
  wire [0:0] s_wallace_cska32_and_2_0;
  wire [0:0] s_wallace_cska32_and_1_1;
  wire [0:0] s_wallace_cska32_ha0_xor0;
  wire [0:0] s_wallace_cska32_ha0_and0;
  wire [0:0] s_wallace_cska32_and_3_0;
  wire [0:0] s_wallace_cska32_and_2_1;
  wire [0:0] s_wallace_cska32_fa0_xor1;
  wire [0:0] s_wallace_cska32_fa0_or0;
  wire [0:0] s_wallace_cska32_and_4_0;
  wire [0:0] s_wallace_cska32_and_3_1;
  wire [0:0] s_wallace_cska32_fa1_xor1;
  wire [0:0] s_wallace_cska32_fa1_or0;
  wire [0:0] s_wallace_cska32_and_5_0;
  wire [0:0] s_wallace_cska32_and_4_1;
  wire [0:0] s_wallace_cska32_fa2_xor1;
  wire [0:0] s_wallace_cska32_fa2_or0;
  wire [0:0] s_wallace_cska32_and_6_0;
  wire [0:0] s_wallace_cska32_and_5_1;
  wire [0:0] s_wallace_cska32_fa3_xor1;
  wire [0:0] s_wallace_cska32_fa3_or0;
  wire [0:0] s_wallace_cska32_and_7_0;
  wire [0:0] s_wallace_cska32_and_6_1;
  wire [0:0] s_wallace_cska32_fa4_xor1;
  wire [0:0] s_wallace_cska32_fa4_or0;
  wire [0:0] s_wallace_cska32_and_8_0;
  wire [0:0] s_wallace_cska32_and_7_1;
  wire [0:0] s_wallace_cska32_fa5_xor1;
  wire [0:0] s_wallace_cska32_fa5_or0;
  wire [0:0] s_wallace_cska32_and_9_0;
  wire [0:0] s_wallace_cska32_and_8_1;
  wire [0:0] s_wallace_cska32_fa6_xor1;
  wire [0:0] s_wallace_cska32_fa6_or0;
  wire [0:0] s_wallace_cska32_and_10_0;
  wire [0:0] s_wallace_cska32_and_9_1;
  wire [0:0] s_wallace_cska32_fa7_xor1;
  wire [0:0] s_wallace_cska32_fa7_or0;
  wire [0:0] s_wallace_cska32_and_11_0;
  wire [0:0] s_wallace_cska32_and_10_1;
  wire [0:0] s_wallace_cska32_fa8_xor1;
  wire [0:0] s_wallace_cska32_fa8_or0;
  wire [0:0] s_wallace_cska32_and_12_0;
  wire [0:0] s_wallace_cska32_and_11_1;
  wire [0:0] s_wallace_cska32_fa9_xor1;
  wire [0:0] s_wallace_cska32_fa9_or0;
  wire [0:0] s_wallace_cska32_and_13_0;
  wire [0:0] s_wallace_cska32_and_12_1;
  wire [0:0] s_wallace_cska32_fa10_xor1;
  wire [0:0] s_wallace_cska32_fa10_or0;
  wire [0:0] s_wallace_cska32_and_14_0;
  wire [0:0] s_wallace_cska32_and_13_1;
  wire [0:0] s_wallace_cska32_fa11_xor1;
  wire [0:0] s_wallace_cska32_fa11_or0;
  wire [0:0] s_wallace_cska32_and_15_0;
  wire [0:0] s_wallace_cska32_and_14_1;
  wire [0:0] s_wallace_cska32_fa12_xor1;
  wire [0:0] s_wallace_cska32_fa12_or0;
  wire [0:0] s_wallace_cska32_and_16_0;
  wire [0:0] s_wallace_cska32_and_15_1;
  wire [0:0] s_wallace_cska32_fa13_xor1;
  wire [0:0] s_wallace_cska32_fa13_or0;
  wire [0:0] s_wallace_cska32_and_17_0;
  wire [0:0] s_wallace_cska32_and_16_1;
  wire [0:0] s_wallace_cska32_fa14_xor1;
  wire [0:0] s_wallace_cska32_fa14_or0;
  wire [0:0] s_wallace_cska32_and_18_0;
  wire [0:0] s_wallace_cska32_and_17_1;
  wire [0:0] s_wallace_cska32_fa15_xor1;
  wire [0:0] s_wallace_cska32_fa15_or0;
  wire [0:0] s_wallace_cska32_and_19_0;
  wire [0:0] s_wallace_cska32_and_18_1;
  wire [0:0] s_wallace_cska32_fa16_xor1;
  wire [0:0] s_wallace_cska32_fa16_or0;
  wire [0:0] s_wallace_cska32_and_20_0;
  wire [0:0] s_wallace_cska32_and_19_1;
  wire [0:0] s_wallace_cska32_fa17_xor1;
  wire [0:0] s_wallace_cska32_fa17_or0;
  wire [0:0] s_wallace_cska32_and_21_0;
  wire [0:0] s_wallace_cska32_and_20_1;
  wire [0:0] s_wallace_cska32_fa18_xor1;
  wire [0:0] s_wallace_cska32_fa18_or0;
  wire [0:0] s_wallace_cska32_and_22_0;
  wire [0:0] s_wallace_cska32_and_21_1;
  wire [0:0] s_wallace_cska32_fa19_xor1;
  wire [0:0] s_wallace_cska32_fa19_or0;
  wire [0:0] s_wallace_cska32_and_23_0;
  wire [0:0] s_wallace_cska32_and_22_1;
  wire [0:0] s_wallace_cska32_fa20_xor1;
  wire [0:0] s_wallace_cska32_fa20_or0;
  wire [0:0] s_wallace_cska32_and_24_0;
  wire [0:0] s_wallace_cska32_and_23_1;
  wire [0:0] s_wallace_cska32_fa21_xor1;
  wire [0:0] s_wallace_cska32_fa21_or0;
  wire [0:0] s_wallace_cska32_and_25_0;
  wire [0:0] s_wallace_cska32_and_24_1;
  wire [0:0] s_wallace_cska32_fa22_xor1;
  wire [0:0] s_wallace_cska32_fa22_or0;
  wire [0:0] s_wallace_cska32_and_26_0;
  wire [0:0] s_wallace_cska32_and_25_1;
  wire [0:0] s_wallace_cska32_fa23_xor1;
  wire [0:0] s_wallace_cska32_fa23_or0;
  wire [0:0] s_wallace_cska32_and_27_0;
  wire [0:0] s_wallace_cska32_and_26_1;
  wire [0:0] s_wallace_cska32_fa24_xor1;
  wire [0:0] s_wallace_cska32_fa24_or0;
  wire [0:0] s_wallace_cska32_and_28_0;
  wire [0:0] s_wallace_cska32_and_27_1;
  wire [0:0] s_wallace_cska32_fa25_xor1;
  wire [0:0] s_wallace_cska32_fa25_or0;
  wire [0:0] s_wallace_cska32_and_29_0;
  wire [0:0] s_wallace_cska32_and_28_1;
  wire [0:0] s_wallace_cska32_fa26_xor1;
  wire [0:0] s_wallace_cska32_fa26_or0;
  wire [0:0] s_wallace_cska32_and_30_0;
  wire [0:0] s_wallace_cska32_and_29_1;
  wire [0:0] s_wallace_cska32_fa27_xor1;
  wire [0:0] s_wallace_cska32_fa27_or0;
  wire [0:0] s_wallace_cska32_nand_31_0;
  wire [0:0] s_wallace_cska32_and_30_1;
  wire [0:0] s_wallace_cska32_fa28_xor1;
  wire [0:0] s_wallace_cska32_fa28_or0;
  wire [0:0] s_wallace_cska32_nand_31_1;
  wire [0:0] s_wallace_cska32_fa29_xor1;
  wire [0:0] s_wallace_cska32_fa29_or0;
  wire [0:0] s_wallace_cska32_nand_31_2;
  wire [0:0] s_wallace_cska32_and_30_3;
  wire [0:0] s_wallace_cska32_fa30_xor1;
  wire [0:0] s_wallace_cska32_fa30_or0;
  wire [0:0] s_wallace_cska32_nand_31_3;
  wire [0:0] s_wallace_cska32_and_30_4;
  wire [0:0] s_wallace_cska32_fa31_xor1;
  wire [0:0] s_wallace_cska32_fa31_or0;
  wire [0:0] s_wallace_cska32_nand_31_4;
  wire [0:0] s_wallace_cska32_and_30_5;
  wire [0:0] s_wallace_cska32_fa32_xor1;
  wire [0:0] s_wallace_cska32_fa32_or0;
  wire [0:0] s_wallace_cska32_nand_31_5;
  wire [0:0] s_wallace_cska32_and_30_6;
  wire [0:0] s_wallace_cska32_fa33_xor1;
  wire [0:0] s_wallace_cska32_fa33_or0;
  wire [0:0] s_wallace_cska32_nand_31_6;
  wire [0:0] s_wallace_cska32_and_30_7;
  wire [0:0] s_wallace_cska32_fa34_xor1;
  wire [0:0] s_wallace_cska32_fa34_or0;
  wire [0:0] s_wallace_cska32_nand_31_7;
  wire [0:0] s_wallace_cska32_and_30_8;
  wire [0:0] s_wallace_cska32_fa35_xor1;
  wire [0:0] s_wallace_cska32_fa35_or0;
  wire [0:0] s_wallace_cska32_nand_31_8;
  wire [0:0] s_wallace_cska32_and_30_9;
  wire [0:0] s_wallace_cska32_fa36_xor1;
  wire [0:0] s_wallace_cska32_fa36_or0;
  wire [0:0] s_wallace_cska32_nand_31_9;
  wire [0:0] s_wallace_cska32_and_30_10;
  wire [0:0] s_wallace_cska32_fa37_xor1;
  wire [0:0] s_wallace_cska32_fa37_or0;
  wire [0:0] s_wallace_cska32_nand_31_10;
  wire [0:0] s_wallace_cska32_and_30_11;
  wire [0:0] s_wallace_cska32_fa38_xor1;
  wire [0:0] s_wallace_cska32_fa38_or0;
  wire [0:0] s_wallace_cska32_nand_31_11;
  wire [0:0] s_wallace_cska32_and_30_12;
  wire [0:0] s_wallace_cska32_fa39_xor1;
  wire [0:0] s_wallace_cska32_fa39_or0;
  wire [0:0] s_wallace_cska32_nand_31_12;
  wire [0:0] s_wallace_cska32_and_30_13;
  wire [0:0] s_wallace_cska32_fa40_xor1;
  wire [0:0] s_wallace_cska32_fa40_or0;
  wire [0:0] s_wallace_cska32_nand_31_13;
  wire [0:0] s_wallace_cska32_and_30_14;
  wire [0:0] s_wallace_cska32_fa41_xor1;
  wire [0:0] s_wallace_cska32_fa41_or0;
  wire [0:0] s_wallace_cska32_nand_31_14;
  wire [0:0] s_wallace_cska32_and_30_15;
  wire [0:0] s_wallace_cska32_fa42_xor1;
  wire [0:0] s_wallace_cska32_fa42_or0;
  wire [0:0] s_wallace_cska32_nand_31_15;
  wire [0:0] s_wallace_cska32_and_30_16;
  wire [0:0] s_wallace_cska32_fa43_xor1;
  wire [0:0] s_wallace_cska32_fa43_or0;
  wire [0:0] s_wallace_cska32_nand_31_16;
  wire [0:0] s_wallace_cska32_and_30_17;
  wire [0:0] s_wallace_cska32_fa44_xor1;
  wire [0:0] s_wallace_cska32_fa44_or0;
  wire [0:0] s_wallace_cska32_nand_31_17;
  wire [0:0] s_wallace_cska32_and_30_18;
  wire [0:0] s_wallace_cska32_fa45_xor1;
  wire [0:0] s_wallace_cska32_fa45_or0;
  wire [0:0] s_wallace_cska32_nand_31_18;
  wire [0:0] s_wallace_cska32_and_30_19;
  wire [0:0] s_wallace_cska32_fa46_xor1;
  wire [0:0] s_wallace_cska32_fa46_or0;
  wire [0:0] s_wallace_cska32_nand_31_19;
  wire [0:0] s_wallace_cska32_and_30_20;
  wire [0:0] s_wallace_cska32_fa47_xor1;
  wire [0:0] s_wallace_cska32_fa47_or0;
  wire [0:0] s_wallace_cska32_nand_31_20;
  wire [0:0] s_wallace_cska32_and_30_21;
  wire [0:0] s_wallace_cska32_fa48_xor1;
  wire [0:0] s_wallace_cska32_fa48_or0;
  wire [0:0] s_wallace_cska32_nand_31_21;
  wire [0:0] s_wallace_cska32_and_30_22;
  wire [0:0] s_wallace_cska32_fa49_xor1;
  wire [0:0] s_wallace_cska32_fa49_or0;
  wire [0:0] s_wallace_cska32_nand_31_22;
  wire [0:0] s_wallace_cska32_and_30_23;
  wire [0:0] s_wallace_cska32_fa50_xor1;
  wire [0:0] s_wallace_cska32_fa50_or0;
  wire [0:0] s_wallace_cska32_nand_31_23;
  wire [0:0] s_wallace_cska32_and_30_24;
  wire [0:0] s_wallace_cska32_fa51_xor1;
  wire [0:0] s_wallace_cska32_fa51_or0;
  wire [0:0] s_wallace_cska32_nand_31_24;
  wire [0:0] s_wallace_cska32_and_30_25;
  wire [0:0] s_wallace_cska32_fa52_xor1;
  wire [0:0] s_wallace_cska32_fa52_or0;
  wire [0:0] s_wallace_cska32_nand_31_25;
  wire [0:0] s_wallace_cska32_and_30_26;
  wire [0:0] s_wallace_cska32_fa53_xor1;
  wire [0:0] s_wallace_cska32_fa53_or0;
  wire [0:0] s_wallace_cska32_nand_31_26;
  wire [0:0] s_wallace_cska32_and_30_27;
  wire [0:0] s_wallace_cska32_fa54_xor1;
  wire [0:0] s_wallace_cska32_fa54_or0;
  wire [0:0] s_wallace_cska32_nand_31_27;
  wire [0:0] s_wallace_cska32_and_30_28;
  wire [0:0] s_wallace_cska32_fa55_xor1;
  wire [0:0] s_wallace_cska32_fa55_or0;
  wire [0:0] s_wallace_cska32_nand_31_28;
  wire [0:0] s_wallace_cska32_and_30_29;
  wire [0:0] s_wallace_cska32_fa56_xor1;
  wire [0:0] s_wallace_cska32_fa56_or0;
  wire [0:0] s_wallace_cska32_nand_31_29;
  wire [0:0] s_wallace_cska32_and_30_30;
  wire [0:0] s_wallace_cska32_fa57_xor1;
  wire [0:0] s_wallace_cska32_fa57_or0;
  wire [0:0] s_wallace_cska32_and_1_2;
  wire [0:0] s_wallace_cska32_and_0_3;
  wire [0:0] s_wallace_cska32_ha1_xor0;
  wire [0:0] s_wallace_cska32_ha1_and0;
  wire [0:0] s_wallace_cska32_and_2_2;
  wire [0:0] s_wallace_cska32_and_1_3;
  wire [0:0] s_wallace_cska32_fa58_xor1;
  wire [0:0] s_wallace_cska32_fa58_or0;
  wire [0:0] s_wallace_cska32_and_3_2;
  wire [0:0] s_wallace_cska32_and_2_3;
  wire [0:0] s_wallace_cska32_fa59_xor1;
  wire [0:0] s_wallace_cska32_fa59_or0;
  wire [0:0] s_wallace_cska32_and_4_2;
  wire [0:0] s_wallace_cska32_and_3_3;
  wire [0:0] s_wallace_cska32_fa60_xor1;
  wire [0:0] s_wallace_cska32_fa60_or0;
  wire [0:0] s_wallace_cska32_and_5_2;
  wire [0:0] s_wallace_cska32_and_4_3;
  wire [0:0] s_wallace_cska32_fa61_xor1;
  wire [0:0] s_wallace_cska32_fa61_or0;
  wire [0:0] s_wallace_cska32_and_6_2;
  wire [0:0] s_wallace_cska32_and_5_3;
  wire [0:0] s_wallace_cska32_fa62_xor1;
  wire [0:0] s_wallace_cska32_fa62_or0;
  wire [0:0] s_wallace_cska32_and_7_2;
  wire [0:0] s_wallace_cska32_and_6_3;
  wire [0:0] s_wallace_cska32_fa63_xor1;
  wire [0:0] s_wallace_cska32_fa63_or0;
  wire [0:0] s_wallace_cska32_and_8_2;
  wire [0:0] s_wallace_cska32_and_7_3;
  wire [0:0] s_wallace_cska32_fa64_xor1;
  wire [0:0] s_wallace_cska32_fa64_or0;
  wire [0:0] s_wallace_cska32_and_9_2;
  wire [0:0] s_wallace_cska32_and_8_3;
  wire [0:0] s_wallace_cska32_fa65_xor1;
  wire [0:0] s_wallace_cska32_fa65_or0;
  wire [0:0] s_wallace_cska32_and_10_2;
  wire [0:0] s_wallace_cska32_and_9_3;
  wire [0:0] s_wallace_cska32_fa66_xor1;
  wire [0:0] s_wallace_cska32_fa66_or0;
  wire [0:0] s_wallace_cska32_and_11_2;
  wire [0:0] s_wallace_cska32_and_10_3;
  wire [0:0] s_wallace_cska32_fa67_xor1;
  wire [0:0] s_wallace_cska32_fa67_or0;
  wire [0:0] s_wallace_cska32_and_12_2;
  wire [0:0] s_wallace_cska32_and_11_3;
  wire [0:0] s_wallace_cska32_fa68_xor1;
  wire [0:0] s_wallace_cska32_fa68_or0;
  wire [0:0] s_wallace_cska32_and_13_2;
  wire [0:0] s_wallace_cska32_and_12_3;
  wire [0:0] s_wallace_cska32_fa69_xor1;
  wire [0:0] s_wallace_cska32_fa69_or0;
  wire [0:0] s_wallace_cska32_and_14_2;
  wire [0:0] s_wallace_cska32_and_13_3;
  wire [0:0] s_wallace_cska32_fa70_xor1;
  wire [0:0] s_wallace_cska32_fa70_or0;
  wire [0:0] s_wallace_cska32_and_15_2;
  wire [0:0] s_wallace_cska32_and_14_3;
  wire [0:0] s_wallace_cska32_fa71_xor1;
  wire [0:0] s_wallace_cska32_fa71_or0;
  wire [0:0] s_wallace_cska32_and_16_2;
  wire [0:0] s_wallace_cska32_and_15_3;
  wire [0:0] s_wallace_cska32_fa72_xor1;
  wire [0:0] s_wallace_cska32_fa72_or0;
  wire [0:0] s_wallace_cska32_and_17_2;
  wire [0:0] s_wallace_cska32_and_16_3;
  wire [0:0] s_wallace_cska32_fa73_xor1;
  wire [0:0] s_wallace_cska32_fa73_or0;
  wire [0:0] s_wallace_cska32_and_18_2;
  wire [0:0] s_wallace_cska32_and_17_3;
  wire [0:0] s_wallace_cska32_fa74_xor1;
  wire [0:0] s_wallace_cska32_fa74_or0;
  wire [0:0] s_wallace_cska32_and_19_2;
  wire [0:0] s_wallace_cska32_and_18_3;
  wire [0:0] s_wallace_cska32_fa75_xor1;
  wire [0:0] s_wallace_cska32_fa75_or0;
  wire [0:0] s_wallace_cska32_and_20_2;
  wire [0:0] s_wallace_cska32_and_19_3;
  wire [0:0] s_wallace_cska32_fa76_xor1;
  wire [0:0] s_wallace_cska32_fa76_or0;
  wire [0:0] s_wallace_cska32_and_21_2;
  wire [0:0] s_wallace_cska32_and_20_3;
  wire [0:0] s_wallace_cska32_fa77_xor1;
  wire [0:0] s_wallace_cska32_fa77_or0;
  wire [0:0] s_wallace_cska32_and_22_2;
  wire [0:0] s_wallace_cska32_and_21_3;
  wire [0:0] s_wallace_cska32_fa78_xor1;
  wire [0:0] s_wallace_cska32_fa78_or0;
  wire [0:0] s_wallace_cska32_and_23_2;
  wire [0:0] s_wallace_cska32_and_22_3;
  wire [0:0] s_wallace_cska32_fa79_xor1;
  wire [0:0] s_wallace_cska32_fa79_or0;
  wire [0:0] s_wallace_cska32_and_24_2;
  wire [0:0] s_wallace_cska32_and_23_3;
  wire [0:0] s_wallace_cska32_fa80_xor1;
  wire [0:0] s_wallace_cska32_fa80_or0;
  wire [0:0] s_wallace_cska32_and_25_2;
  wire [0:0] s_wallace_cska32_and_24_3;
  wire [0:0] s_wallace_cska32_fa81_xor1;
  wire [0:0] s_wallace_cska32_fa81_or0;
  wire [0:0] s_wallace_cska32_and_26_2;
  wire [0:0] s_wallace_cska32_and_25_3;
  wire [0:0] s_wallace_cska32_fa82_xor1;
  wire [0:0] s_wallace_cska32_fa82_or0;
  wire [0:0] s_wallace_cska32_and_27_2;
  wire [0:0] s_wallace_cska32_and_26_3;
  wire [0:0] s_wallace_cska32_fa83_xor1;
  wire [0:0] s_wallace_cska32_fa83_or0;
  wire [0:0] s_wallace_cska32_and_28_2;
  wire [0:0] s_wallace_cska32_and_27_3;
  wire [0:0] s_wallace_cska32_fa84_xor1;
  wire [0:0] s_wallace_cska32_fa84_or0;
  wire [0:0] s_wallace_cska32_and_29_2;
  wire [0:0] s_wallace_cska32_and_28_3;
  wire [0:0] s_wallace_cska32_fa85_xor1;
  wire [0:0] s_wallace_cska32_fa85_or0;
  wire [0:0] s_wallace_cska32_and_30_2;
  wire [0:0] s_wallace_cska32_and_29_3;
  wire [0:0] s_wallace_cska32_fa86_xor1;
  wire [0:0] s_wallace_cska32_fa86_or0;
  wire [0:0] s_wallace_cska32_and_29_4;
  wire [0:0] s_wallace_cska32_and_28_5;
  wire [0:0] s_wallace_cska32_fa87_xor1;
  wire [0:0] s_wallace_cska32_fa87_or0;
  wire [0:0] s_wallace_cska32_and_29_5;
  wire [0:0] s_wallace_cska32_and_28_6;
  wire [0:0] s_wallace_cska32_fa88_xor1;
  wire [0:0] s_wallace_cska32_fa88_or0;
  wire [0:0] s_wallace_cska32_and_29_6;
  wire [0:0] s_wallace_cska32_and_28_7;
  wire [0:0] s_wallace_cska32_fa89_xor1;
  wire [0:0] s_wallace_cska32_fa89_or0;
  wire [0:0] s_wallace_cska32_and_29_7;
  wire [0:0] s_wallace_cska32_and_28_8;
  wire [0:0] s_wallace_cska32_fa90_xor1;
  wire [0:0] s_wallace_cska32_fa90_or0;
  wire [0:0] s_wallace_cska32_and_29_8;
  wire [0:0] s_wallace_cska32_and_28_9;
  wire [0:0] s_wallace_cska32_fa91_xor1;
  wire [0:0] s_wallace_cska32_fa91_or0;
  wire [0:0] s_wallace_cska32_and_29_9;
  wire [0:0] s_wallace_cska32_and_28_10;
  wire [0:0] s_wallace_cska32_fa92_xor1;
  wire [0:0] s_wallace_cska32_fa92_or0;
  wire [0:0] s_wallace_cska32_and_29_10;
  wire [0:0] s_wallace_cska32_and_28_11;
  wire [0:0] s_wallace_cska32_fa93_xor1;
  wire [0:0] s_wallace_cska32_fa93_or0;
  wire [0:0] s_wallace_cska32_and_29_11;
  wire [0:0] s_wallace_cska32_and_28_12;
  wire [0:0] s_wallace_cska32_fa94_xor1;
  wire [0:0] s_wallace_cska32_fa94_or0;
  wire [0:0] s_wallace_cska32_and_29_12;
  wire [0:0] s_wallace_cska32_and_28_13;
  wire [0:0] s_wallace_cska32_fa95_xor1;
  wire [0:0] s_wallace_cska32_fa95_or0;
  wire [0:0] s_wallace_cska32_and_29_13;
  wire [0:0] s_wallace_cska32_and_28_14;
  wire [0:0] s_wallace_cska32_fa96_xor1;
  wire [0:0] s_wallace_cska32_fa96_or0;
  wire [0:0] s_wallace_cska32_and_29_14;
  wire [0:0] s_wallace_cska32_and_28_15;
  wire [0:0] s_wallace_cska32_fa97_xor1;
  wire [0:0] s_wallace_cska32_fa97_or0;
  wire [0:0] s_wallace_cska32_and_29_15;
  wire [0:0] s_wallace_cska32_and_28_16;
  wire [0:0] s_wallace_cska32_fa98_xor1;
  wire [0:0] s_wallace_cska32_fa98_or0;
  wire [0:0] s_wallace_cska32_and_29_16;
  wire [0:0] s_wallace_cska32_and_28_17;
  wire [0:0] s_wallace_cska32_fa99_xor1;
  wire [0:0] s_wallace_cska32_fa99_or0;
  wire [0:0] s_wallace_cska32_and_29_17;
  wire [0:0] s_wallace_cska32_and_28_18;
  wire [0:0] s_wallace_cska32_fa100_xor1;
  wire [0:0] s_wallace_cska32_fa100_or0;
  wire [0:0] s_wallace_cska32_and_29_18;
  wire [0:0] s_wallace_cska32_and_28_19;
  wire [0:0] s_wallace_cska32_fa101_xor1;
  wire [0:0] s_wallace_cska32_fa101_or0;
  wire [0:0] s_wallace_cska32_and_29_19;
  wire [0:0] s_wallace_cska32_and_28_20;
  wire [0:0] s_wallace_cska32_fa102_xor1;
  wire [0:0] s_wallace_cska32_fa102_or0;
  wire [0:0] s_wallace_cska32_and_29_20;
  wire [0:0] s_wallace_cska32_and_28_21;
  wire [0:0] s_wallace_cska32_fa103_xor1;
  wire [0:0] s_wallace_cska32_fa103_or0;
  wire [0:0] s_wallace_cska32_and_29_21;
  wire [0:0] s_wallace_cska32_and_28_22;
  wire [0:0] s_wallace_cska32_fa104_xor1;
  wire [0:0] s_wallace_cska32_fa104_or0;
  wire [0:0] s_wallace_cska32_and_29_22;
  wire [0:0] s_wallace_cska32_and_28_23;
  wire [0:0] s_wallace_cska32_fa105_xor1;
  wire [0:0] s_wallace_cska32_fa105_or0;
  wire [0:0] s_wallace_cska32_and_29_23;
  wire [0:0] s_wallace_cska32_and_28_24;
  wire [0:0] s_wallace_cska32_fa106_xor1;
  wire [0:0] s_wallace_cska32_fa106_or0;
  wire [0:0] s_wallace_cska32_and_29_24;
  wire [0:0] s_wallace_cska32_and_28_25;
  wire [0:0] s_wallace_cska32_fa107_xor1;
  wire [0:0] s_wallace_cska32_fa107_or0;
  wire [0:0] s_wallace_cska32_and_29_25;
  wire [0:0] s_wallace_cska32_and_28_26;
  wire [0:0] s_wallace_cska32_fa108_xor1;
  wire [0:0] s_wallace_cska32_fa108_or0;
  wire [0:0] s_wallace_cska32_and_29_26;
  wire [0:0] s_wallace_cska32_and_28_27;
  wire [0:0] s_wallace_cska32_fa109_xor1;
  wire [0:0] s_wallace_cska32_fa109_or0;
  wire [0:0] s_wallace_cska32_and_29_27;
  wire [0:0] s_wallace_cska32_and_28_28;
  wire [0:0] s_wallace_cska32_fa110_xor1;
  wire [0:0] s_wallace_cska32_fa110_or0;
  wire [0:0] s_wallace_cska32_and_29_28;
  wire [0:0] s_wallace_cska32_and_28_29;
  wire [0:0] s_wallace_cska32_fa111_xor1;
  wire [0:0] s_wallace_cska32_fa111_or0;
  wire [0:0] s_wallace_cska32_and_29_29;
  wire [0:0] s_wallace_cska32_and_28_30;
  wire [0:0] s_wallace_cska32_fa112_xor1;
  wire [0:0] s_wallace_cska32_fa112_or0;
  wire [0:0] s_wallace_cska32_and_29_30;
  wire [0:0] s_wallace_cska32_nand_28_31;
  wire [0:0] s_wallace_cska32_fa113_xor1;
  wire [0:0] s_wallace_cska32_fa113_or0;
  wire [0:0] s_wallace_cska32_and_0_4;
  wire [0:0] s_wallace_cska32_ha2_xor0;
  wire [0:0] s_wallace_cska32_ha2_and0;
  wire [0:0] s_wallace_cska32_and_1_4;
  wire [0:0] s_wallace_cska32_and_0_5;
  wire [0:0] s_wallace_cska32_fa114_xor1;
  wire [0:0] s_wallace_cska32_fa114_or0;
  wire [0:0] s_wallace_cska32_and_2_4;
  wire [0:0] s_wallace_cska32_and_1_5;
  wire [0:0] s_wallace_cska32_fa115_xor1;
  wire [0:0] s_wallace_cska32_fa115_or0;
  wire [0:0] s_wallace_cska32_and_3_4;
  wire [0:0] s_wallace_cska32_and_2_5;
  wire [0:0] s_wallace_cska32_fa116_xor1;
  wire [0:0] s_wallace_cska32_fa116_or0;
  wire [0:0] s_wallace_cska32_and_4_4;
  wire [0:0] s_wallace_cska32_and_3_5;
  wire [0:0] s_wallace_cska32_fa117_xor1;
  wire [0:0] s_wallace_cska32_fa117_or0;
  wire [0:0] s_wallace_cska32_and_5_4;
  wire [0:0] s_wallace_cska32_and_4_5;
  wire [0:0] s_wallace_cska32_fa118_xor1;
  wire [0:0] s_wallace_cska32_fa118_or0;
  wire [0:0] s_wallace_cska32_and_6_4;
  wire [0:0] s_wallace_cska32_and_5_5;
  wire [0:0] s_wallace_cska32_fa119_xor1;
  wire [0:0] s_wallace_cska32_fa119_or0;
  wire [0:0] s_wallace_cska32_and_7_4;
  wire [0:0] s_wallace_cska32_and_6_5;
  wire [0:0] s_wallace_cska32_fa120_xor1;
  wire [0:0] s_wallace_cska32_fa120_or0;
  wire [0:0] s_wallace_cska32_and_8_4;
  wire [0:0] s_wallace_cska32_and_7_5;
  wire [0:0] s_wallace_cska32_fa121_xor1;
  wire [0:0] s_wallace_cska32_fa121_or0;
  wire [0:0] s_wallace_cska32_and_9_4;
  wire [0:0] s_wallace_cska32_and_8_5;
  wire [0:0] s_wallace_cska32_fa122_xor1;
  wire [0:0] s_wallace_cska32_fa122_or0;
  wire [0:0] s_wallace_cska32_and_10_4;
  wire [0:0] s_wallace_cska32_and_9_5;
  wire [0:0] s_wallace_cska32_fa123_xor1;
  wire [0:0] s_wallace_cska32_fa123_or0;
  wire [0:0] s_wallace_cska32_and_11_4;
  wire [0:0] s_wallace_cska32_and_10_5;
  wire [0:0] s_wallace_cska32_fa124_xor1;
  wire [0:0] s_wallace_cska32_fa124_or0;
  wire [0:0] s_wallace_cska32_and_12_4;
  wire [0:0] s_wallace_cska32_and_11_5;
  wire [0:0] s_wallace_cska32_fa125_xor1;
  wire [0:0] s_wallace_cska32_fa125_or0;
  wire [0:0] s_wallace_cska32_and_13_4;
  wire [0:0] s_wallace_cska32_and_12_5;
  wire [0:0] s_wallace_cska32_fa126_xor1;
  wire [0:0] s_wallace_cska32_fa126_or0;
  wire [0:0] s_wallace_cska32_and_14_4;
  wire [0:0] s_wallace_cska32_and_13_5;
  wire [0:0] s_wallace_cska32_fa127_xor1;
  wire [0:0] s_wallace_cska32_fa127_or0;
  wire [0:0] s_wallace_cska32_and_15_4;
  wire [0:0] s_wallace_cska32_and_14_5;
  wire [0:0] s_wallace_cska32_fa128_xor1;
  wire [0:0] s_wallace_cska32_fa128_or0;
  wire [0:0] s_wallace_cska32_and_16_4;
  wire [0:0] s_wallace_cska32_and_15_5;
  wire [0:0] s_wallace_cska32_fa129_xor1;
  wire [0:0] s_wallace_cska32_fa129_or0;
  wire [0:0] s_wallace_cska32_and_17_4;
  wire [0:0] s_wallace_cska32_and_16_5;
  wire [0:0] s_wallace_cska32_fa130_xor1;
  wire [0:0] s_wallace_cska32_fa130_or0;
  wire [0:0] s_wallace_cska32_and_18_4;
  wire [0:0] s_wallace_cska32_and_17_5;
  wire [0:0] s_wallace_cska32_fa131_xor1;
  wire [0:0] s_wallace_cska32_fa131_or0;
  wire [0:0] s_wallace_cska32_and_19_4;
  wire [0:0] s_wallace_cska32_and_18_5;
  wire [0:0] s_wallace_cska32_fa132_xor1;
  wire [0:0] s_wallace_cska32_fa132_or0;
  wire [0:0] s_wallace_cska32_and_20_4;
  wire [0:0] s_wallace_cska32_and_19_5;
  wire [0:0] s_wallace_cska32_fa133_xor1;
  wire [0:0] s_wallace_cska32_fa133_or0;
  wire [0:0] s_wallace_cska32_and_21_4;
  wire [0:0] s_wallace_cska32_and_20_5;
  wire [0:0] s_wallace_cska32_fa134_xor1;
  wire [0:0] s_wallace_cska32_fa134_or0;
  wire [0:0] s_wallace_cska32_and_22_4;
  wire [0:0] s_wallace_cska32_and_21_5;
  wire [0:0] s_wallace_cska32_fa135_xor1;
  wire [0:0] s_wallace_cska32_fa135_or0;
  wire [0:0] s_wallace_cska32_and_23_4;
  wire [0:0] s_wallace_cska32_and_22_5;
  wire [0:0] s_wallace_cska32_fa136_xor1;
  wire [0:0] s_wallace_cska32_fa136_or0;
  wire [0:0] s_wallace_cska32_and_24_4;
  wire [0:0] s_wallace_cska32_and_23_5;
  wire [0:0] s_wallace_cska32_fa137_xor1;
  wire [0:0] s_wallace_cska32_fa137_or0;
  wire [0:0] s_wallace_cska32_and_25_4;
  wire [0:0] s_wallace_cska32_and_24_5;
  wire [0:0] s_wallace_cska32_fa138_xor1;
  wire [0:0] s_wallace_cska32_fa138_or0;
  wire [0:0] s_wallace_cska32_and_26_4;
  wire [0:0] s_wallace_cska32_and_25_5;
  wire [0:0] s_wallace_cska32_fa139_xor1;
  wire [0:0] s_wallace_cska32_fa139_or0;
  wire [0:0] s_wallace_cska32_and_27_4;
  wire [0:0] s_wallace_cska32_and_26_5;
  wire [0:0] s_wallace_cska32_fa140_xor1;
  wire [0:0] s_wallace_cska32_fa140_or0;
  wire [0:0] s_wallace_cska32_and_28_4;
  wire [0:0] s_wallace_cska32_and_27_5;
  wire [0:0] s_wallace_cska32_fa141_xor1;
  wire [0:0] s_wallace_cska32_fa141_or0;
  wire [0:0] s_wallace_cska32_and_27_6;
  wire [0:0] s_wallace_cska32_and_26_7;
  wire [0:0] s_wallace_cska32_fa142_xor1;
  wire [0:0] s_wallace_cska32_fa142_or0;
  wire [0:0] s_wallace_cska32_and_27_7;
  wire [0:0] s_wallace_cska32_and_26_8;
  wire [0:0] s_wallace_cska32_fa143_xor1;
  wire [0:0] s_wallace_cska32_fa143_or0;
  wire [0:0] s_wallace_cska32_and_27_8;
  wire [0:0] s_wallace_cska32_and_26_9;
  wire [0:0] s_wallace_cska32_fa144_xor1;
  wire [0:0] s_wallace_cska32_fa144_or0;
  wire [0:0] s_wallace_cska32_and_27_9;
  wire [0:0] s_wallace_cska32_and_26_10;
  wire [0:0] s_wallace_cska32_fa145_xor1;
  wire [0:0] s_wallace_cska32_fa145_or0;
  wire [0:0] s_wallace_cska32_and_27_10;
  wire [0:0] s_wallace_cska32_and_26_11;
  wire [0:0] s_wallace_cska32_fa146_xor1;
  wire [0:0] s_wallace_cska32_fa146_or0;
  wire [0:0] s_wallace_cska32_and_27_11;
  wire [0:0] s_wallace_cska32_and_26_12;
  wire [0:0] s_wallace_cska32_fa147_xor1;
  wire [0:0] s_wallace_cska32_fa147_or0;
  wire [0:0] s_wallace_cska32_and_27_12;
  wire [0:0] s_wallace_cska32_and_26_13;
  wire [0:0] s_wallace_cska32_fa148_xor1;
  wire [0:0] s_wallace_cska32_fa148_or0;
  wire [0:0] s_wallace_cska32_and_27_13;
  wire [0:0] s_wallace_cska32_and_26_14;
  wire [0:0] s_wallace_cska32_fa149_xor1;
  wire [0:0] s_wallace_cska32_fa149_or0;
  wire [0:0] s_wallace_cska32_and_27_14;
  wire [0:0] s_wallace_cska32_and_26_15;
  wire [0:0] s_wallace_cska32_fa150_xor1;
  wire [0:0] s_wallace_cska32_fa150_or0;
  wire [0:0] s_wallace_cska32_and_27_15;
  wire [0:0] s_wallace_cska32_and_26_16;
  wire [0:0] s_wallace_cska32_fa151_xor1;
  wire [0:0] s_wallace_cska32_fa151_or0;
  wire [0:0] s_wallace_cska32_and_27_16;
  wire [0:0] s_wallace_cska32_and_26_17;
  wire [0:0] s_wallace_cska32_fa152_xor1;
  wire [0:0] s_wallace_cska32_fa152_or0;
  wire [0:0] s_wallace_cska32_and_27_17;
  wire [0:0] s_wallace_cska32_and_26_18;
  wire [0:0] s_wallace_cska32_fa153_xor1;
  wire [0:0] s_wallace_cska32_fa153_or0;
  wire [0:0] s_wallace_cska32_and_27_18;
  wire [0:0] s_wallace_cska32_and_26_19;
  wire [0:0] s_wallace_cska32_fa154_xor1;
  wire [0:0] s_wallace_cska32_fa154_or0;
  wire [0:0] s_wallace_cska32_and_27_19;
  wire [0:0] s_wallace_cska32_and_26_20;
  wire [0:0] s_wallace_cska32_fa155_xor1;
  wire [0:0] s_wallace_cska32_fa155_or0;
  wire [0:0] s_wallace_cska32_and_27_20;
  wire [0:0] s_wallace_cska32_and_26_21;
  wire [0:0] s_wallace_cska32_fa156_xor1;
  wire [0:0] s_wallace_cska32_fa156_or0;
  wire [0:0] s_wallace_cska32_and_27_21;
  wire [0:0] s_wallace_cska32_and_26_22;
  wire [0:0] s_wallace_cska32_fa157_xor1;
  wire [0:0] s_wallace_cska32_fa157_or0;
  wire [0:0] s_wallace_cska32_and_27_22;
  wire [0:0] s_wallace_cska32_and_26_23;
  wire [0:0] s_wallace_cska32_fa158_xor1;
  wire [0:0] s_wallace_cska32_fa158_or0;
  wire [0:0] s_wallace_cska32_and_27_23;
  wire [0:0] s_wallace_cska32_and_26_24;
  wire [0:0] s_wallace_cska32_fa159_xor1;
  wire [0:0] s_wallace_cska32_fa159_or0;
  wire [0:0] s_wallace_cska32_and_27_24;
  wire [0:0] s_wallace_cska32_and_26_25;
  wire [0:0] s_wallace_cska32_fa160_xor1;
  wire [0:0] s_wallace_cska32_fa160_or0;
  wire [0:0] s_wallace_cska32_and_27_25;
  wire [0:0] s_wallace_cska32_and_26_26;
  wire [0:0] s_wallace_cska32_fa161_xor1;
  wire [0:0] s_wallace_cska32_fa161_or0;
  wire [0:0] s_wallace_cska32_and_27_26;
  wire [0:0] s_wallace_cska32_and_26_27;
  wire [0:0] s_wallace_cska32_fa162_xor1;
  wire [0:0] s_wallace_cska32_fa162_or0;
  wire [0:0] s_wallace_cska32_and_27_27;
  wire [0:0] s_wallace_cska32_and_26_28;
  wire [0:0] s_wallace_cska32_fa163_xor1;
  wire [0:0] s_wallace_cska32_fa163_or0;
  wire [0:0] s_wallace_cska32_and_27_28;
  wire [0:0] s_wallace_cska32_and_26_29;
  wire [0:0] s_wallace_cska32_fa164_xor1;
  wire [0:0] s_wallace_cska32_fa164_or0;
  wire [0:0] s_wallace_cska32_and_27_29;
  wire [0:0] s_wallace_cska32_and_26_30;
  wire [0:0] s_wallace_cska32_fa165_xor1;
  wire [0:0] s_wallace_cska32_fa165_or0;
  wire [0:0] s_wallace_cska32_and_27_30;
  wire [0:0] s_wallace_cska32_nand_26_31;
  wire [0:0] s_wallace_cska32_fa166_xor1;
  wire [0:0] s_wallace_cska32_fa166_or0;
  wire [0:0] s_wallace_cska32_nand_27_31;
  wire [0:0] s_wallace_cska32_fa167_xor1;
  wire [0:0] s_wallace_cska32_fa167_or0;
  wire [0:0] s_wallace_cska32_ha3_xor0;
  wire [0:0] s_wallace_cska32_ha3_and0;
  wire [0:0] s_wallace_cska32_and_0_6;
  wire [0:0] s_wallace_cska32_fa168_xor1;
  wire [0:0] s_wallace_cska32_fa168_or0;
  wire [0:0] s_wallace_cska32_and_1_6;
  wire [0:0] s_wallace_cska32_and_0_7;
  wire [0:0] s_wallace_cska32_fa169_xor1;
  wire [0:0] s_wallace_cska32_fa169_or0;
  wire [0:0] s_wallace_cska32_and_2_6;
  wire [0:0] s_wallace_cska32_and_1_7;
  wire [0:0] s_wallace_cska32_fa170_xor1;
  wire [0:0] s_wallace_cska32_fa170_or0;
  wire [0:0] s_wallace_cska32_and_3_6;
  wire [0:0] s_wallace_cska32_and_2_7;
  wire [0:0] s_wallace_cska32_fa171_xor1;
  wire [0:0] s_wallace_cska32_fa171_or0;
  wire [0:0] s_wallace_cska32_and_4_6;
  wire [0:0] s_wallace_cska32_and_3_7;
  wire [0:0] s_wallace_cska32_fa172_xor1;
  wire [0:0] s_wallace_cska32_fa172_or0;
  wire [0:0] s_wallace_cska32_and_5_6;
  wire [0:0] s_wallace_cska32_and_4_7;
  wire [0:0] s_wallace_cska32_fa173_xor1;
  wire [0:0] s_wallace_cska32_fa173_or0;
  wire [0:0] s_wallace_cska32_and_6_6;
  wire [0:0] s_wallace_cska32_and_5_7;
  wire [0:0] s_wallace_cska32_fa174_xor1;
  wire [0:0] s_wallace_cska32_fa174_or0;
  wire [0:0] s_wallace_cska32_and_7_6;
  wire [0:0] s_wallace_cska32_and_6_7;
  wire [0:0] s_wallace_cska32_fa175_xor1;
  wire [0:0] s_wallace_cska32_fa175_or0;
  wire [0:0] s_wallace_cska32_and_8_6;
  wire [0:0] s_wallace_cska32_and_7_7;
  wire [0:0] s_wallace_cska32_fa176_xor1;
  wire [0:0] s_wallace_cska32_fa176_or0;
  wire [0:0] s_wallace_cska32_and_9_6;
  wire [0:0] s_wallace_cska32_and_8_7;
  wire [0:0] s_wallace_cska32_fa177_xor1;
  wire [0:0] s_wallace_cska32_fa177_or0;
  wire [0:0] s_wallace_cska32_and_10_6;
  wire [0:0] s_wallace_cska32_and_9_7;
  wire [0:0] s_wallace_cska32_fa178_xor1;
  wire [0:0] s_wallace_cska32_fa178_or0;
  wire [0:0] s_wallace_cska32_and_11_6;
  wire [0:0] s_wallace_cska32_and_10_7;
  wire [0:0] s_wallace_cska32_fa179_xor1;
  wire [0:0] s_wallace_cska32_fa179_or0;
  wire [0:0] s_wallace_cska32_and_12_6;
  wire [0:0] s_wallace_cska32_and_11_7;
  wire [0:0] s_wallace_cska32_fa180_xor1;
  wire [0:0] s_wallace_cska32_fa180_or0;
  wire [0:0] s_wallace_cska32_and_13_6;
  wire [0:0] s_wallace_cska32_and_12_7;
  wire [0:0] s_wallace_cska32_fa181_xor1;
  wire [0:0] s_wallace_cska32_fa181_or0;
  wire [0:0] s_wallace_cska32_and_14_6;
  wire [0:0] s_wallace_cska32_and_13_7;
  wire [0:0] s_wallace_cska32_fa182_xor1;
  wire [0:0] s_wallace_cska32_fa182_or0;
  wire [0:0] s_wallace_cska32_and_15_6;
  wire [0:0] s_wallace_cska32_and_14_7;
  wire [0:0] s_wallace_cska32_fa183_xor1;
  wire [0:0] s_wallace_cska32_fa183_or0;
  wire [0:0] s_wallace_cska32_and_16_6;
  wire [0:0] s_wallace_cska32_and_15_7;
  wire [0:0] s_wallace_cska32_fa184_xor1;
  wire [0:0] s_wallace_cska32_fa184_or0;
  wire [0:0] s_wallace_cska32_and_17_6;
  wire [0:0] s_wallace_cska32_and_16_7;
  wire [0:0] s_wallace_cska32_fa185_xor1;
  wire [0:0] s_wallace_cska32_fa185_or0;
  wire [0:0] s_wallace_cska32_and_18_6;
  wire [0:0] s_wallace_cska32_and_17_7;
  wire [0:0] s_wallace_cska32_fa186_xor1;
  wire [0:0] s_wallace_cska32_fa186_or0;
  wire [0:0] s_wallace_cska32_and_19_6;
  wire [0:0] s_wallace_cska32_and_18_7;
  wire [0:0] s_wallace_cska32_fa187_xor1;
  wire [0:0] s_wallace_cska32_fa187_or0;
  wire [0:0] s_wallace_cska32_and_20_6;
  wire [0:0] s_wallace_cska32_and_19_7;
  wire [0:0] s_wallace_cska32_fa188_xor1;
  wire [0:0] s_wallace_cska32_fa188_or0;
  wire [0:0] s_wallace_cska32_and_21_6;
  wire [0:0] s_wallace_cska32_and_20_7;
  wire [0:0] s_wallace_cska32_fa189_xor1;
  wire [0:0] s_wallace_cska32_fa189_or0;
  wire [0:0] s_wallace_cska32_and_22_6;
  wire [0:0] s_wallace_cska32_and_21_7;
  wire [0:0] s_wallace_cska32_fa190_xor1;
  wire [0:0] s_wallace_cska32_fa190_or0;
  wire [0:0] s_wallace_cska32_and_23_6;
  wire [0:0] s_wallace_cska32_and_22_7;
  wire [0:0] s_wallace_cska32_fa191_xor1;
  wire [0:0] s_wallace_cska32_fa191_or0;
  wire [0:0] s_wallace_cska32_and_24_6;
  wire [0:0] s_wallace_cska32_and_23_7;
  wire [0:0] s_wallace_cska32_fa192_xor1;
  wire [0:0] s_wallace_cska32_fa192_or0;
  wire [0:0] s_wallace_cska32_and_25_6;
  wire [0:0] s_wallace_cska32_and_24_7;
  wire [0:0] s_wallace_cska32_fa193_xor1;
  wire [0:0] s_wallace_cska32_fa193_or0;
  wire [0:0] s_wallace_cska32_and_26_6;
  wire [0:0] s_wallace_cska32_and_25_7;
  wire [0:0] s_wallace_cska32_fa194_xor1;
  wire [0:0] s_wallace_cska32_fa194_or0;
  wire [0:0] s_wallace_cska32_and_25_8;
  wire [0:0] s_wallace_cska32_and_24_9;
  wire [0:0] s_wallace_cska32_fa195_xor1;
  wire [0:0] s_wallace_cska32_fa195_or0;
  wire [0:0] s_wallace_cska32_and_25_9;
  wire [0:0] s_wallace_cska32_and_24_10;
  wire [0:0] s_wallace_cska32_fa196_xor1;
  wire [0:0] s_wallace_cska32_fa196_or0;
  wire [0:0] s_wallace_cska32_and_25_10;
  wire [0:0] s_wallace_cska32_and_24_11;
  wire [0:0] s_wallace_cska32_fa197_xor1;
  wire [0:0] s_wallace_cska32_fa197_or0;
  wire [0:0] s_wallace_cska32_and_25_11;
  wire [0:0] s_wallace_cska32_and_24_12;
  wire [0:0] s_wallace_cska32_fa198_xor1;
  wire [0:0] s_wallace_cska32_fa198_or0;
  wire [0:0] s_wallace_cska32_and_25_12;
  wire [0:0] s_wallace_cska32_and_24_13;
  wire [0:0] s_wallace_cska32_fa199_xor1;
  wire [0:0] s_wallace_cska32_fa199_or0;
  wire [0:0] s_wallace_cska32_and_25_13;
  wire [0:0] s_wallace_cska32_and_24_14;
  wire [0:0] s_wallace_cska32_fa200_xor1;
  wire [0:0] s_wallace_cska32_fa200_or0;
  wire [0:0] s_wallace_cska32_and_25_14;
  wire [0:0] s_wallace_cska32_and_24_15;
  wire [0:0] s_wallace_cska32_fa201_xor1;
  wire [0:0] s_wallace_cska32_fa201_or0;
  wire [0:0] s_wallace_cska32_and_25_15;
  wire [0:0] s_wallace_cska32_and_24_16;
  wire [0:0] s_wallace_cska32_fa202_xor1;
  wire [0:0] s_wallace_cska32_fa202_or0;
  wire [0:0] s_wallace_cska32_and_25_16;
  wire [0:0] s_wallace_cska32_and_24_17;
  wire [0:0] s_wallace_cska32_fa203_xor1;
  wire [0:0] s_wallace_cska32_fa203_or0;
  wire [0:0] s_wallace_cska32_and_25_17;
  wire [0:0] s_wallace_cska32_and_24_18;
  wire [0:0] s_wallace_cska32_fa204_xor1;
  wire [0:0] s_wallace_cska32_fa204_or0;
  wire [0:0] s_wallace_cska32_and_25_18;
  wire [0:0] s_wallace_cska32_and_24_19;
  wire [0:0] s_wallace_cska32_fa205_xor1;
  wire [0:0] s_wallace_cska32_fa205_or0;
  wire [0:0] s_wallace_cska32_and_25_19;
  wire [0:0] s_wallace_cska32_and_24_20;
  wire [0:0] s_wallace_cska32_fa206_xor1;
  wire [0:0] s_wallace_cska32_fa206_or0;
  wire [0:0] s_wallace_cska32_and_25_20;
  wire [0:0] s_wallace_cska32_and_24_21;
  wire [0:0] s_wallace_cska32_fa207_xor1;
  wire [0:0] s_wallace_cska32_fa207_or0;
  wire [0:0] s_wallace_cska32_and_25_21;
  wire [0:0] s_wallace_cska32_and_24_22;
  wire [0:0] s_wallace_cska32_fa208_xor1;
  wire [0:0] s_wallace_cska32_fa208_or0;
  wire [0:0] s_wallace_cska32_and_25_22;
  wire [0:0] s_wallace_cska32_and_24_23;
  wire [0:0] s_wallace_cska32_fa209_xor1;
  wire [0:0] s_wallace_cska32_fa209_or0;
  wire [0:0] s_wallace_cska32_and_25_23;
  wire [0:0] s_wallace_cska32_and_24_24;
  wire [0:0] s_wallace_cska32_fa210_xor1;
  wire [0:0] s_wallace_cska32_fa210_or0;
  wire [0:0] s_wallace_cska32_and_25_24;
  wire [0:0] s_wallace_cska32_and_24_25;
  wire [0:0] s_wallace_cska32_fa211_xor1;
  wire [0:0] s_wallace_cska32_fa211_or0;
  wire [0:0] s_wallace_cska32_and_25_25;
  wire [0:0] s_wallace_cska32_and_24_26;
  wire [0:0] s_wallace_cska32_fa212_xor1;
  wire [0:0] s_wallace_cska32_fa212_or0;
  wire [0:0] s_wallace_cska32_and_25_26;
  wire [0:0] s_wallace_cska32_and_24_27;
  wire [0:0] s_wallace_cska32_fa213_xor1;
  wire [0:0] s_wallace_cska32_fa213_or0;
  wire [0:0] s_wallace_cska32_and_25_27;
  wire [0:0] s_wallace_cska32_and_24_28;
  wire [0:0] s_wallace_cska32_fa214_xor1;
  wire [0:0] s_wallace_cska32_fa214_or0;
  wire [0:0] s_wallace_cska32_and_25_28;
  wire [0:0] s_wallace_cska32_and_24_29;
  wire [0:0] s_wallace_cska32_fa215_xor1;
  wire [0:0] s_wallace_cska32_fa215_or0;
  wire [0:0] s_wallace_cska32_and_25_29;
  wire [0:0] s_wallace_cska32_and_24_30;
  wire [0:0] s_wallace_cska32_fa216_xor1;
  wire [0:0] s_wallace_cska32_fa216_or0;
  wire [0:0] s_wallace_cska32_and_25_30;
  wire [0:0] s_wallace_cska32_nand_24_31;
  wire [0:0] s_wallace_cska32_fa217_xor1;
  wire [0:0] s_wallace_cska32_fa217_or0;
  wire [0:0] s_wallace_cska32_nand_25_31;
  wire [0:0] s_wallace_cska32_fa218_xor1;
  wire [0:0] s_wallace_cska32_fa218_or0;
  wire [0:0] s_wallace_cska32_fa219_xor1;
  wire [0:0] s_wallace_cska32_fa219_or0;
  wire [0:0] s_wallace_cska32_ha4_xor0;
  wire [0:0] s_wallace_cska32_ha4_and0;
  wire [0:0] s_wallace_cska32_fa220_xor1;
  wire [0:0] s_wallace_cska32_fa220_or0;
  wire [0:0] s_wallace_cska32_and_0_8;
  wire [0:0] s_wallace_cska32_fa221_xor1;
  wire [0:0] s_wallace_cska32_fa221_or0;
  wire [0:0] s_wallace_cska32_and_1_8;
  wire [0:0] s_wallace_cska32_and_0_9;
  wire [0:0] s_wallace_cska32_fa222_xor1;
  wire [0:0] s_wallace_cska32_fa222_or0;
  wire [0:0] s_wallace_cska32_and_2_8;
  wire [0:0] s_wallace_cska32_and_1_9;
  wire [0:0] s_wallace_cska32_fa223_xor1;
  wire [0:0] s_wallace_cska32_fa223_or0;
  wire [0:0] s_wallace_cska32_and_3_8;
  wire [0:0] s_wallace_cska32_and_2_9;
  wire [0:0] s_wallace_cska32_fa224_xor1;
  wire [0:0] s_wallace_cska32_fa224_or0;
  wire [0:0] s_wallace_cska32_and_4_8;
  wire [0:0] s_wallace_cska32_and_3_9;
  wire [0:0] s_wallace_cska32_fa225_xor1;
  wire [0:0] s_wallace_cska32_fa225_or0;
  wire [0:0] s_wallace_cska32_and_5_8;
  wire [0:0] s_wallace_cska32_and_4_9;
  wire [0:0] s_wallace_cska32_fa226_xor1;
  wire [0:0] s_wallace_cska32_fa226_or0;
  wire [0:0] s_wallace_cska32_and_6_8;
  wire [0:0] s_wallace_cska32_and_5_9;
  wire [0:0] s_wallace_cska32_fa227_xor1;
  wire [0:0] s_wallace_cska32_fa227_or0;
  wire [0:0] s_wallace_cska32_and_7_8;
  wire [0:0] s_wallace_cska32_and_6_9;
  wire [0:0] s_wallace_cska32_fa228_xor1;
  wire [0:0] s_wallace_cska32_fa228_or0;
  wire [0:0] s_wallace_cska32_and_8_8;
  wire [0:0] s_wallace_cska32_and_7_9;
  wire [0:0] s_wallace_cska32_fa229_xor1;
  wire [0:0] s_wallace_cska32_fa229_or0;
  wire [0:0] s_wallace_cska32_and_9_8;
  wire [0:0] s_wallace_cska32_and_8_9;
  wire [0:0] s_wallace_cska32_fa230_xor1;
  wire [0:0] s_wallace_cska32_fa230_or0;
  wire [0:0] s_wallace_cska32_and_10_8;
  wire [0:0] s_wallace_cska32_and_9_9;
  wire [0:0] s_wallace_cska32_fa231_xor1;
  wire [0:0] s_wallace_cska32_fa231_or0;
  wire [0:0] s_wallace_cska32_and_11_8;
  wire [0:0] s_wallace_cska32_and_10_9;
  wire [0:0] s_wallace_cska32_fa232_xor1;
  wire [0:0] s_wallace_cska32_fa232_or0;
  wire [0:0] s_wallace_cska32_and_12_8;
  wire [0:0] s_wallace_cska32_and_11_9;
  wire [0:0] s_wallace_cska32_fa233_xor1;
  wire [0:0] s_wallace_cska32_fa233_or0;
  wire [0:0] s_wallace_cska32_and_13_8;
  wire [0:0] s_wallace_cska32_and_12_9;
  wire [0:0] s_wallace_cska32_fa234_xor1;
  wire [0:0] s_wallace_cska32_fa234_or0;
  wire [0:0] s_wallace_cska32_and_14_8;
  wire [0:0] s_wallace_cska32_and_13_9;
  wire [0:0] s_wallace_cska32_fa235_xor1;
  wire [0:0] s_wallace_cska32_fa235_or0;
  wire [0:0] s_wallace_cska32_and_15_8;
  wire [0:0] s_wallace_cska32_and_14_9;
  wire [0:0] s_wallace_cska32_fa236_xor1;
  wire [0:0] s_wallace_cska32_fa236_or0;
  wire [0:0] s_wallace_cska32_and_16_8;
  wire [0:0] s_wallace_cska32_and_15_9;
  wire [0:0] s_wallace_cska32_fa237_xor1;
  wire [0:0] s_wallace_cska32_fa237_or0;
  wire [0:0] s_wallace_cska32_and_17_8;
  wire [0:0] s_wallace_cska32_and_16_9;
  wire [0:0] s_wallace_cska32_fa238_xor1;
  wire [0:0] s_wallace_cska32_fa238_or0;
  wire [0:0] s_wallace_cska32_and_18_8;
  wire [0:0] s_wallace_cska32_and_17_9;
  wire [0:0] s_wallace_cska32_fa239_xor1;
  wire [0:0] s_wallace_cska32_fa239_or0;
  wire [0:0] s_wallace_cska32_and_19_8;
  wire [0:0] s_wallace_cska32_and_18_9;
  wire [0:0] s_wallace_cska32_fa240_xor1;
  wire [0:0] s_wallace_cska32_fa240_or0;
  wire [0:0] s_wallace_cska32_and_20_8;
  wire [0:0] s_wallace_cska32_and_19_9;
  wire [0:0] s_wallace_cska32_fa241_xor1;
  wire [0:0] s_wallace_cska32_fa241_or0;
  wire [0:0] s_wallace_cska32_and_21_8;
  wire [0:0] s_wallace_cska32_and_20_9;
  wire [0:0] s_wallace_cska32_fa242_xor1;
  wire [0:0] s_wallace_cska32_fa242_or0;
  wire [0:0] s_wallace_cska32_and_22_8;
  wire [0:0] s_wallace_cska32_and_21_9;
  wire [0:0] s_wallace_cska32_fa243_xor1;
  wire [0:0] s_wallace_cska32_fa243_or0;
  wire [0:0] s_wallace_cska32_and_23_8;
  wire [0:0] s_wallace_cska32_and_22_9;
  wire [0:0] s_wallace_cska32_fa244_xor1;
  wire [0:0] s_wallace_cska32_fa244_or0;
  wire [0:0] s_wallace_cska32_and_24_8;
  wire [0:0] s_wallace_cska32_and_23_9;
  wire [0:0] s_wallace_cska32_fa245_xor1;
  wire [0:0] s_wallace_cska32_fa245_or0;
  wire [0:0] s_wallace_cska32_and_23_10;
  wire [0:0] s_wallace_cska32_and_22_11;
  wire [0:0] s_wallace_cska32_fa246_xor1;
  wire [0:0] s_wallace_cska32_fa246_or0;
  wire [0:0] s_wallace_cska32_and_23_11;
  wire [0:0] s_wallace_cska32_and_22_12;
  wire [0:0] s_wallace_cska32_fa247_xor1;
  wire [0:0] s_wallace_cska32_fa247_or0;
  wire [0:0] s_wallace_cska32_and_23_12;
  wire [0:0] s_wallace_cska32_and_22_13;
  wire [0:0] s_wallace_cska32_fa248_xor1;
  wire [0:0] s_wallace_cska32_fa248_or0;
  wire [0:0] s_wallace_cska32_and_23_13;
  wire [0:0] s_wallace_cska32_and_22_14;
  wire [0:0] s_wallace_cska32_fa249_xor1;
  wire [0:0] s_wallace_cska32_fa249_or0;
  wire [0:0] s_wallace_cska32_and_23_14;
  wire [0:0] s_wallace_cska32_and_22_15;
  wire [0:0] s_wallace_cska32_fa250_xor1;
  wire [0:0] s_wallace_cska32_fa250_or0;
  wire [0:0] s_wallace_cska32_and_23_15;
  wire [0:0] s_wallace_cska32_and_22_16;
  wire [0:0] s_wallace_cska32_fa251_xor1;
  wire [0:0] s_wallace_cska32_fa251_or0;
  wire [0:0] s_wallace_cska32_and_23_16;
  wire [0:0] s_wallace_cska32_and_22_17;
  wire [0:0] s_wallace_cska32_fa252_xor1;
  wire [0:0] s_wallace_cska32_fa252_or0;
  wire [0:0] s_wallace_cska32_and_23_17;
  wire [0:0] s_wallace_cska32_and_22_18;
  wire [0:0] s_wallace_cska32_fa253_xor1;
  wire [0:0] s_wallace_cska32_fa253_or0;
  wire [0:0] s_wallace_cska32_and_23_18;
  wire [0:0] s_wallace_cska32_and_22_19;
  wire [0:0] s_wallace_cska32_fa254_xor1;
  wire [0:0] s_wallace_cska32_fa254_or0;
  wire [0:0] s_wallace_cska32_and_23_19;
  wire [0:0] s_wallace_cska32_and_22_20;
  wire [0:0] s_wallace_cska32_fa255_xor1;
  wire [0:0] s_wallace_cska32_fa255_or0;
  wire [0:0] s_wallace_cska32_and_23_20;
  wire [0:0] s_wallace_cska32_and_22_21;
  wire [0:0] s_wallace_cska32_fa256_xor1;
  wire [0:0] s_wallace_cska32_fa256_or0;
  wire [0:0] s_wallace_cska32_and_23_21;
  wire [0:0] s_wallace_cska32_and_22_22;
  wire [0:0] s_wallace_cska32_fa257_xor1;
  wire [0:0] s_wallace_cska32_fa257_or0;
  wire [0:0] s_wallace_cska32_and_23_22;
  wire [0:0] s_wallace_cska32_and_22_23;
  wire [0:0] s_wallace_cska32_fa258_xor1;
  wire [0:0] s_wallace_cska32_fa258_or0;
  wire [0:0] s_wallace_cska32_and_23_23;
  wire [0:0] s_wallace_cska32_and_22_24;
  wire [0:0] s_wallace_cska32_fa259_xor1;
  wire [0:0] s_wallace_cska32_fa259_or0;
  wire [0:0] s_wallace_cska32_and_23_24;
  wire [0:0] s_wallace_cska32_and_22_25;
  wire [0:0] s_wallace_cska32_fa260_xor1;
  wire [0:0] s_wallace_cska32_fa260_or0;
  wire [0:0] s_wallace_cska32_and_23_25;
  wire [0:0] s_wallace_cska32_and_22_26;
  wire [0:0] s_wallace_cska32_fa261_xor1;
  wire [0:0] s_wallace_cska32_fa261_or0;
  wire [0:0] s_wallace_cska32_and_23_26;
  wire [0:0] s_wallace_cska32_and_22_27;
  wire [0:0] s_wallace_cska32_fa262_xor1;
  wire [0:0] s_wallace_cska32_fa262_or0;
  wire [0:0] s_wallace_cska32_and_23_27;
  wire [0:0] s_wallace_cska32_and_22_28;
  wire [0:0] s_wallace_cska32_fa263_xor1;
  wire [0:0] s_wallace_cska32_fa263_or0;
  wire [0:0] s_wallace_cska32_and_23_28;
  wire [0:0] s_wallace_cska32_and_22_29;
  wire [0:0] s_wallace_cska32_fa264_xor1;
  wire [0:0] s_wallace_cska32_fa264_or0;
  wire [0:0] s_wallace_cska32_and_23_29;
  wire [0:0] s_wallace_cska32_and_22_30;
  wire [0:0] s_wallace_cska32_fa265_xor1;
  wire [0:0] s_wallace_cska32_fa265_or0;
  wire [0:0] s_wallace_cska32_and_23_30;
  wire [0:0] s_wallace_cska32_nand_22_31;
  wire [0:0] s_wallace_cska32_fa266_xor1;
  wire [0:0] s_wallace_cska32_fa266_or0;
  wire [0:0] s_wallace_cska32_nand_23_31;
  wire [0:0] s_wallace_cska32_fa267_xor1;
  wire [0:0] s_wallace_cska32_fa267_or0;
  wire [0:0] s_wallace_cska32_fa268_xor1;
  wire [0:0] s_wallace_cska32_fa268_or0;
  wire [0:0] s_wallace_cska32_fa269_xor1;
  wire [0:0] s_wallace_cska32_fa269_or0;
  wire [0:0] s_wallace_cska32_ha5_xor0;
  wire [0:0] s_wallace_cska32_ha5_and0;
  wire [0:0] s_wallace_cska32_fa270_xor1;
  wire [0:0] s_wallace_cska32_fa270_or0;
  wire [0:0] s_wallace_cska32_fa271_xor1;
  wire [0:0] s_wallace_cska32_fa271_or0;
  wire [0:0] s_wallace_cska32_and_0_10;
  wire [0:0] s_wallace_cska32_fa272_xor1;
  wire [0:0] s_wallace_cska32_fa272_or0;
  wire [0:0] s_wallace_cska32_and_1_10;
  wire [0:0] s_wallace_cska32_and_0_11;
  wire [0:0] s_wallace_cska32_fa273_xor1;
  wire [0:0] s_wallace_cska32_fa273_or0;
  wire [0:0] s_wallace_cska32_and_2_10;
  wire [0:0] s_wallace_cska32_and_1_11;
  wire [0:0] s_wallace_cska32_fa274_xor1;
  wire [0:0] s_wallace_cska32_fa274_or0;
  wire [0:0] s_wallace_cska32_and_3_10;
  wire [0:0] s_wallace_cska32_and_2_11;
  wire [0:0] s_wallace_cska32_fa275_xor1;
  wire [0:0] s_wallace_cska32_fa275_or0;
  wire [0:0] s_wallace_cska32_and_4_10;
  wire [0:0] s_wallace_cska32_and_3_11;
  wire [0:0] s_wallace_cska32_fa276_xor1;
  wire [0:0] s_wallace_cska32_fa276_or0;
  wire [0:0] s_wallace_cska32_and_5_10;
  wire [0:0] s_wallace_cska32_and_4_11;
  wire [0:0] s_wallace_cska32_fa277_xor1;
  wire [0:0] s_wallace_cska32_fa277_or0;
  wire [0:0] s_wallace_cska32_and_6_10;
  wire [0:0] s_wallace_cska32_and_5_11;
  wire [0:0] s_wallace_cska32_fa278_xor1;
  wire [0:0] s_wallace_cska32_fa278_or0;
  wire [0:0] s_wallace_cska32_and_7_10;
  wire [0:0] s_wallace_cska32_and_6_11;
  wire [0:0] s_wallace_cska32_fa279_xor1;
  wire [0:0] s_wallace_cska32_fa279_or0;
  wire [0:0] s_wallace_cska32_and_8_10;
  wire [0:0] s_wallace_cska32_and_7_11;
  wire [0:0] s_wallace_cska32_fa280_xor1;
  wire [0:0] s_wallace_cska32_fa280_or0;
  wire [0:0] s_wallace_cska32_and_9_10;
  wire [0:0] s_wallace_cska32_and_8_11;
  wire [0:0] s_wallace_cska32_fa281_xor1;
  wire [0:0] s_wallace_cska32_fa281_or0;
  wire [0:0] s_wallace_cska32_and_10_10;
  wire [0:0] s_wallace_cska32_and_9_11;
  wire [0:0] s_wallace_cska32_fa282_xor1;
  wire [0:0] s_wallace_cska32_fa282_or0;
  wire [0:0] s_wallace_cska32_and_11_10;
  wire [0:0] s_wallace_cska32_and_10_11;
  wire [0:0] s_wallace_cska32_fa283_xor1;
  wire [0:0] s_wallace_cska32_fa283_or0;
  wire [0:0] s_wallace_cska32_and_12_10;
  wire [0:0] s_wallace_cska32_and_11_11;
  wire [0:0] s_wallace_cska32_fa284_xor1;
  wire [0:0] s_wallace_cska32_fa284_or0;
  wire [0:0] s_wallace_cska32_and_13_10;
  wire [0:0] s_wallace_cska32_and_12_11;
  wire [0:0] s_wallace_cska32_fa285_xor1;
  wire [0:0] s_wallace_cska32_fa285_or0;
  wire [0:0] s_wallace_cska32_and_14_10;
  wire [0:0] s_wallace_cska32_and_13_11;
  wire [0:0] s_wallace_cska32_fa286_xor1;
  wire [0:0] s_wallace_cska32_fa286_or0;
  wire [0:0] s_wallace_cska32_and_15_10;
  wire [0:0] s_wallace_cska32_and_14_11;
  wire [0:0] s_wallace_cska32_fa287_xor1;
  wire [0:0] s_wallace_cska32_fa287_or0;
  wire [0:0] s_wallace_cska32_and_16_10;
  wire [0:0] s_wallace_cska32_and_15_11;
  wire [0:0] s_wallace_cska32_fa288_xor1;
  wire [0:0] s_wallace_cska32_fa288_or0;
  wire [0:0] s_wallace_cska32_and_17_10;
  wire [0:0] s_wallace_cska32_and_16_11;
  wire [0:0] s_wallace_cska32_fa289_xor1;
  wire [0:0] s_wallace_cska32_fa289_or0;
  wire [0:0] s_wallace_cska32_and_18_10;
  wire [0:0] s_wallace_cska32_and_17_11;
  wire [0:0] s_wallace_cska32_fa290_xor1;
  wire [0:0] s_wallace_cska32_fa290_or0;
  wire [0:0] s_wallace_cska32_and_19_10;
  wire [0:0] s_wallace_cska32_and_18_11;
  wire [0:0] s_wallace_cska32_fa291_xor1;
  wire [0:0] s_wallace_cska32_fa291_or0;
  wire [0:0] s_wallace_cska32_and_20_10;
  wire [0:0] s_wallace_cska32_and_19_11;
  wire [0:0] s_wallace_cska32_fa292_xor1;
  wire [0:0] s_wallace_cska32_fa292_or0;
  wire [0:0] s_wallace_cska32_and_21_10;
  wire [0:0] s_wallace_cska32_and_20_11;
  wire [0:0] s_wallace_cska32_fa293_xor1;
  wire [0:0] s_wallace_cska32_fa293_or0;
  wire [0:0] s_wallace_cska32_and_22_10;
  wire [0:0] s_wallace_cska32_and_21_11;
  wire [0:0] s_wallace_cska32_fa294_xor1;
  wire [0:0] s_wallace_cska32_fa294_or0;
  wire [0:0] s_wallace_cska32_and_21_12;
  wire [0:0] s_wallace_cska32_and_20_13;
  wire [0:0] s_wallace_cska32_fa295_xor1;
  wire [0:0] s_wallace_cska32_fa295_or0;
  wire [0:0] s_wallace_cska32_and_21_13;
  wire [0:0] s_wallace_cska32_and_20_14;
  wire [0:0] s_wallace_cska32_fa296_xor1;
  wire [0:0] s_wallace_cska32_fa296_or0;
  wire [0:0] s_wallace_cska32_and_21_14;
  wire [0:0] s_wallace_cska32_and_20_15;
  wire [0:0] s_wallace_cska32_fa297_xor1;
  wire [0:0] s_wallace_cska32_fa297_or0;
  wire [0:0] s_wallace_cska32_and_21_15;
  wire [0:0] s_wallace_cska32_and_20_16;
  wire [0:0] s_wallace_cska32_fa298_xor1;
  wire [0:0] s_wallace_cska32_fa298_or0;
  wire [0:0] s_wallace_cska32_and_21_16;
  wire [0:0] s_wallace_cska32_and_20_17;
  wire [0:0] s_wallace_cska32_fa299_xor1;
  wire [0:0] s_wallace_cska32_fa299_or0;
  wire [0:0] s_wallace_cska32_and_21_17;
  wire [0:0] s_wallace_cska32_and_20_18;
  wire [0:0] s_wallace_cska32_fa300_xor1;
  wire [0:0] s_wallace_cska32_fa300_or0;
  wire [0:0] s_wallace_cska32_and_21_18;
  wire [0:0] s_wallace_cska32_and_20_19;
  wire [0:0] s_wallace_cska32_fa301_xor1;
  wire [0:0] s_wallace_cska32_fa301_or0;
  wire [0:0] s_wallace_cska32_and_21_19;
  wire [0:0] s_wallace_cska32_and_20_20;
  wire [0:0] s_wallace_cska32_fa302_xor1;
  wire [0:0] s_wallace_cska32_fa302_or0;
  wire [0:0] s_wallace_cska32_and_21_20;
  wire [0:0] s_wallace_cska32_and_20_21;
  wire [0:0] s_wallace_cska32_fa303_xor1;
  wire [0:0] s_wallace_cska32_fa303_or0;
  wire [0:0] s_wallace_cska32_and_21_21;
  wire [0:0] s_wallace_cska32_and_20_22;
  wire [0:0] s_wallace_cska32_fa304_xor1;
  wire [0:0] s_wallace_cska32_fa304_or0;
  wire [0:0] s_wallace_cska32_and_21_22;
  wire [0:0] s_wallace_cska32_and_20_23;
  wire [0:0] s_wallace_cska32_fa305_xor1;
  wire [0:0] s_wallace_cska32_fa305_or0;
  wire [0:0] s_wallace_cska32_and_21_23;
  wire [0:0] s_wallace_cska32_and_20_24;
  wire [0:0] s_wallace_cska32_fa306_xor1;
  wire [0:0] s_wallace_cska32_fa306_or0;
  wire [0:0] s_wallace_cska32_and_21_24;
  wire [0:0] s_wallace_cska32_and_20_25;
  wire [0:0] s_wallace_cska32_fa307_xor1;
  wire [0:0] s_wallace_cska32_fa307_or0;
  wire [0:0] s_wallace_cska32_and_21_25;
  wire [0:0] s_wallace_cska32_and_20_26;
  wire [0:0] s_wallace_cska32_fa308_xor1;
  wire [0:0] s_wallace_cska32_fa308_or0;
  wire [0:0] s_wallace_cska32_and_21_26;
  wire [0:0] s_wallace_cska32_and_20_27;
  wire [0:0] s_wallace_cska32_fa309_xor1;
  wire [0:0] s_wallace_cska32_fa309_or0;
  wire [0:0] s_wallace_cska32_and_21_27;
  wire [0:0] s_wallace_cska32_and_20_28;
  wire [0:0] s_wallace_cska32_fa310_xor1;
  wire [0:0] s_wallace_cska32_fa310_or0;
  wire [0:0] s_wallace_cska32_and_21_28;
  wire [0:0] s_wallace_cska32_and_20_29;
  wire [0:0] s_wallace_cska32_fa311_xor1;
  wire [0:0] s_wallace_cska32_fa311_or0;
  wire [0:0] s_wallace_cska32_and_21_29;
  wire [0:0] s_wallace_cska32_and_20_30;
  wire [0:0] s_wallace_cska32_fa312_xor1;
  wire [0:0] s_wallace_cska32_fa312_or0;
  wire [0:0] s_wallace_cska32_and_21_30;
  wire [0:0] s_wallace_cska32_nand_20_31;
  wire [0:0] s_wallace_cska32_fa313_xor1;
  wire [0:0] s_wallace_cska32_fa313_or0;
  wire [0:0] s_wallace_cska32_nand_21_31;
  wire [0:0] s_wallace_cska32_fa314_xor1;
  wire [0:0] s_wallace_cska32_fa314_or0;
  wire [0:0] s_wallace_cska32_fa315_xor1;
  wire [0:0] s_wallace_cska32_fa315_or0;
  wire [0:0] s_wallace_cska32_fa316_xor1;
  wire [0:0] s_wallace_cska32_fa316_or0;
  wire [0:0] s_wallace_cska32_fa317_xor1;
  wire [0:0] s_wallace_cska32_fa317_or0;
  wire [0:0] s_wallace_cska32_ha6_xor0;
  wire [0:0] s_wallace_cska32_ha6_and0;
  wire [0:0] s_wallace_cska32_fa318_xor1;
  wire [0:0] s_wallace_cska32_fa318_or0;
  wire [0:0] s_wallace_cska32_fa319_xor1;
  wire [0:0] s_wallace_cska32_fa319_or0;
  wire [0:0] s_wallace_cska32_fa320_xor1;
  wire [0:0] s_wallace_cska32_fa320_or0;
  wire [0:0] s_wallace_cska32_and_0_12;
  wire [0:0] s_wallace_cska32_fa321_xor1;
  wire [0:0] s_wallace_cska32_fa321_or0;
  wire [0:0] s_wallace_cska32_and_1_12;
  wire [0:0] s_wallace_cska32_and_0_13;
  wire [0:0] s_wallace_cska32_fa322_xor1;
  wire [0:0] s_wallace_cska32_fa322_or0;
  wire [0:0] s_wallace_cska32_and_2_12;
  wire [0:0] s_wallace_cska32_and_1_13;
  wire [0:0] s_wallace_cska32_fa323_xor1;
  wire [0:0] s_wallace_cska32_fa323_or0;
  wire [0:0] s_wallace_cska32_and_3_12;
  wire [0:0] s_wallace_cska32_and_2_13;
  wire [0:0] s_wallace_cska32_fa324_xor1;
  wire [0:0] s_wallace_cska32_fa324_or0;
  wire [0:0] s_wallace_cska32_and_4_12;
  wire [0:0] s_wallace_cska32_and_3_13;
  wire [0:0] s_wallace_cska32_fa325_xor1;
  wire [0:0] s_wallace_cska32_fa325_or0;
  wire [0:0] s_wallace_cska32_and_5_12;
  wire [0:0] s_wallace_cska32_and_4_13;
  wire [0:0] s_wallace_cska32_fa326_xor1;
  wire [0:0] s_wallace_cska32_fa326_or0;
  wire [0:0] s_wallace_cska32_and_6_12;
  wire [0:0] s_wallace_cska32_and_5_13;
  wire [0:0] s_wallace_cska32_fa327_xor1;
  wire [0:0] s_wallace_cska32_fa327_or0;
  wire [0:0] s_wallace_cska32_and_7_12;
  wire [0:0] s_wallace_cska32_and_6_13;
  wire [0:0] s_wallace_cska32_fa328_xor1;
  wire [0:0] s_wallace_cska32_fa328_or0;
  wire [0:0] s_wallace_cska32_and_8_12;
  wire [0:0] s_wallace_cska32_and_7_13;
  wire [0:0] s_wallace_cska32_fa329_xor1;
  wire [0:0] s_wallace_cska32_fa329_or0;
  wire [0:0] s_wallace_cska32_and_9_12;
  wire [0:0] s_wallace_cska32_and_8_13;
  wire [0:0] s_wallace_cska32_fa330_xor1;
  wire [0:0] s_wallace_cska32_fa330_or0;
  wire [0:0] s_wallace_cska32_and_10_12;
  wire [0:0] s_wallace_cska32_and_9_13;
  wire [0:0] s_wallace_cska32_fa331_xor1;
  wire [0:0] s_wallace_cska32_fa331_or0;
  wire [0:0] s_wallace_cska32_and_11_12;
  wire [0:0] s_wallace_cska32_and_10_13;
  wire [0:0] s_wallace_cska32_fa332_xor1;
  wire [0:0] s_wallace_cska32_fa332_or0;
  wire [0:0] s_wallace_cska32_and_12_12;
  wire [0:0] s_wallace_cska32_and_11_13;
  wire [0:0] s_wallace_cska32_fa333_xor1;
  wire [0:0] s_wallace_cska32_fa333_or0;
  wire [0:0] s_wallace_cska32_and_13_12;
  wire [0:0] s_wallace_cska32_and_12_13;
  wire [0:0] s_wallace_cska32_fa334_xor1;
  wire [0:0] s_wallace_cska32_fa334_or0;
  wire [0:0] s_wallace_cska32_and_14_12;
  wire [0:0] s_wallace_cska32_and_13_13;
  wire [0:0] s_wallace_cska32_fa335_xor1;
  wire [0:0] s_wallace_cska32_fa335_or0;
  wire [0:0] s_wallace_cska32_and_15_12;
  wire [0:0] s_wallace_cska32_and_14_13;
  wire [0:0] s_wallace_cska32_fa336_xor1;
  wire [0:0] s_wallace_cska32_fa336_or0;
  wire [0:0] s_wallace_cska32_and_16_12;
  wire [0:0] s_wallace_cska32_and_15_13;
  wire [0:0] s_wallace_cska32_fa337_xor1;
  wire [0:0] s_wallace_cska32_fa337_or0;
  wire [0:0] s_wallace_cska32_and_17_12;
  wire [0:0] s_wallace_cska32_and_16_13;
  wire [0:0] s_wallace_cska32_fa338_xor1;
  wire [0:0] s_wallace_cska32_fa338_or0;
  wire [0:0] s_wallace_cska32_and_18_12;
  wire [0:0] s_wallace_cska32_and_17_13;
  wire [0:0] s_wallace_cska32_fa339_xor1;
  wire [0:0] s_wallace_cska32_fa339_or0;
  wire [0:0] s_wallace_cska32_and_19_12;
  wire [0:0] s_wallace_cska32_and_18_13;
  wire [0:0] s_wallace_cska32_fa340_xor1;
  wire [0:0] s_wallace_cska32_fa340_or0;
  wire [0:0] s_wallace_cska32_and_20_12;
  wire [0:0] s_wallace_cska32_and_19_13;
  wire [0:0] s_wallace_cska32_fa341_xor1;
  wire [0:0] s_wallace_cska32_fa341_or0;
  wire [0:0] s_wallace_cska32_and_19_14;
  wire [0:0] s_wallace_cska32_and_18_15;
  wire [0:0] s_wallace_cska32_fa342_xor1;
  wire [0:0] s_wallace_cska32_fa342_or0;
  wire [0:0] s_wallace_cska32_and_19_15;
  wire [0:0] s_wallace_cska32_and_18_16;
  wire [0:0] s_wallace_cska32_fa343_xor1;
  wire [0:0] s_wallace_cska32_fa343_or0;
  wire [0:0] s_wallace_cska32_and_19_16;
  wire [0:0] s_wallace_cska32_and_18_17;
  wire [0:0] s_wallace_cska32_fa344_xor1;
  wire [0:0] s_wallace_cska32_fa344_or0;
  wire [0:0] s_wallace_cska32_and_19_17;
  wire [0:0] s_wallace_cska32_and_18_18;
  wire [0:0] s_wallace_cska32_fa345_xor1;
  wire [0:0] s_wallace_cska32_fa345_or0;
  wire [0:0] s_wallace_cska32_and_19_18;
  wire [0:0] s_wallace_cska32_and_18_19;
  wire [0:0] s_wallace_cska32_fa346_xor1;
  wire [0:0] s_wallace_cska32_fa346_or0;
  wire [0:0] s_wallace_cska32_and_19_19;
  wire [0:0] s_wallace_cska32_and_18_20;
  wire [0:0] s_wallace_cska32_fa347_xor1;
  wire [0:0] s_wallace_cska32_fa347_or0;
  wire [0:0] s_wallace_cska32_and_19_20;
  wire [0:0] s_wallace_cska32_and_18_21;
  wire [0:0] s_wallace_cska32_fa348_xor1;
  wire [0:0] s_wallace_cska32_fa348_or0;
  wire [0:0] s_wallace_cska32_and_19_21;
  wire [0:0] s_wallace_cska32_and_18_22;
  wire [0:0] s_wallace_cska32_fa349_xor1;
  wire [0:0] s_wallace_cska32_fa349_or0;
  wire [0:0] s_wallace_cska32_and_19_22;
  wire [0:0] s_wallace_cska32_and_18_23;
  wire [0:0] s_wallace_cska32_fa350_xor1;
  wire [0:0] s_wallace_cska32_fa350_or0;
  wire [0:0] s_wallace_cska32_and_19_23;
  wire [0:0] s_wallace_cska32_and_18_24;
  wire [0:0] s_wallace_cska32_fa351_xor1;
  wire [0:0] s_wallace_cska32_fa351_or0;
  wire [0:0] s_wallace_cska32_and_19_24;
  wire [0:0] s_wallace_cska32_and_18_25;
  wire [0:0] s_wallace_cska32_fa352_xor1;
  wire [0:0] s_wallace_cska32_fa352_or0;
  wire [0:0] s_wallace_cska32_and_19_25;
  wire [0:0] s_wallace_cska32_and_18_26;
  wire [0:0] s_wallace_cska32_fa353_xor1;
  wire [0:0] s_wallace_cska32_fa353_or0;
  wire [0:0] s_wallace_cska32_and_19_26;
  wire [0:0] s_wallace_cska32_and_18_27;
  wire [0:0] s_wallace_cska32_fa354_xor1;
  wire [0:0] s_wallace_cska32_fa354_or0;
  wire [0:0] s_wallace_cska32_and_19_27;
  wire [0:0] s_wallace_cska32_and_18_28;
  wire [0:0] s_wallace_cska32_fa355_xor1;
  wire [0:0] s_wallace_cska32_fa355_or0;
  wire [0:0] s_wallace_cska32_and_19_28;
  wire [0:0] s_wallace_cska32_and_18_29;
  wire [0:0] s_wallace_cska32_fa356_xor1;
  wire [0:0] s_wallace_cska32_fa356_or0;
  wire [0:0] s_wallace_cska32_and_19_29;
  wire [0:0] s_wallace_cska32_and_18_30;
  wire [0:0] s_wallace_cska32_fa357_xor1;
  wire [0:0] s_wallace_cska32_fa357_or0;
  wire [0:0] s_wallace_cska32_and_19_30;
  wire [0:0] s_wallace_cska32_nand_18_31;
  wire [0:0] s_wallace_cska32_fa358_xor1;
  wire [0:0] s_wallace_cska32_fa358_or0;
  wire [0:0] s_wallace_cska32_nand_19_31;
  wire [0:0] s_wallace_cska32_fa359_xor1;
  wire [0:0] s_wallace_cska32_fa359_or0;
  wire [0:0] s_wallace_cska32_fa360_xor1;
  wire [0:0] s_wallace_cska32_fa360_or0;
  wire [0:0] s_wallace_cska32_fa361_xor1;
  wire [0:0] s_wallace_cska32_fa361_or0;
  wire [0:0] s_wallace_cska32_fa362_xor1;
  wire [0:0] s_wallace_cska32_fa362_or0;
  wire [0:0] s_wallace_cska32_fa363_xor1;
  wire [0:0] s_wallace_cska32_fa363_or0;
  wire [0:0] s_wallace_cska32_ha7_xor0;
  wire [0:0] s_wallace_cska32_ha7_and0;
  wire [0:0] s_wallace_cska32_fa364_xor1;
  wire [0:0] s_wallace_cska32_fa364_or0;
  wire [0:0] s_wallace_cska32_fa365_xor1;
  wire [0:0] s_wallace_cska32_fa365_or0;
  wire [0:0] s_wallace_cska32_fa366_xor1;
  wire [0:0] s_wallace_cska32_fa366_or0;
  wire [0:0] s_wallace_cska32_fa367_xor1;
  wire [0:0] s_wallace_cska32_fa367_or0;
  wire [0:0] s_wallace_cska32_and_0_14;
  wire [0:0] s_wallace_cska32_fa368_xor1;
  wire [0:0] s_wallace_cska32_fa368_or0;
  wire [0:0] s_wallace_cska32_and_1_14;
  wire [0:0] s_wallace_cska32_and_0_15;
  wire [0:0] s_wallace_cska32_fa369_xor1;
  wire [0:0] s_wallace_cska32_fa369_or0;
  wire [0:0] s_wallace_cska32_and_2_14;
  wire [0:0] s_wallace_cska32_and_1_15;
  wire [0:0] s_wallace_cska32_fa370_xor1;
  wire [0:0] s_wallace_cska32_fa370_or0;
  wire [0:0] s_wallace_cska32_and_3_14;
  wire [0:0] s_wallace_cska32_and_2_15;
  wire [0:0] s_wallace_cska32_fa371_xor1;
  wire [0:0] s_wallace_cska32_fa371_or0;
  wire [0:0] s_wallace_cska32_and_4_14;
  wire [0:0] s_wallace_cska32_and_3_15;
  wire [0:0] s_wallace_cska32_fa372_xor1;
  wire [0:0] s_wallace_cska32_fa372_or0;
  wire [0:0] s_wallace_cska32_and_5_14;
  wire [0:0] s_wallace_cska32_and_4_15;
  wire [0:0] s_wallace_cska32_fa373_xor1;
  wire [0:0] s_wallace_cska32_fa373_or0;
  wire [0:0] s_wallace_cska32_and_6_14;
  wire [0:0] s_wallace_cska32_and_5_15;
  wire [0:0] s_wallace_cska32_fa374_xor1;
  wire [0:0] s_wallace_cska32_fa374_or0;
  wire [0:0] s_wallace_cska32_and_7_14;
  wire [0:0] s_wallace_cska32_and_6_15;
  wire [0:0] s_wallace_cska32_fa375_xor1;
  wire [0:0] s_wallace_cska32_fa375_or0;
  wire [0:0] s_wallace_cska32_and_8_14;
  wire [0:0] s_wallace_cska32_and_7_15;
  wire [0:0] s_wallace_cska32_fa376_xor1;
  wire [0:0] s_wallace_cska32_fa376_or0;
  wire [0:0] s_wallace_cska32_and_9_14;
  wire [0:0] s_wallace_cska32_and_8_15;
  wire [0:0] s_wallace_cska32_fa377_xor1;
  wire [0:0] s_wallace_cska32_fa377_or0;
  wire [0:0] s_wallace_cska32_and_10_14;
  wire [0:0] s_wallace_cska32_and_9_15;
  wire [0:0] s_wallace_cska32_fa378_xor1;
  wire [0:0] s_wallace_cska32_fa378_or0;
  wire [0:0] s_wallace_cska32_and_11_14;
  wire [0:0] s_wallace_cska32_and_10_15;
  wire [0:0] s_wallace_cska32_fa379_xor1;
  wire [0:0] s_wallace_cska32_fa379_or0;
  wire [0:0] s_wallace_cska32_and_12_14;
  wire [0:0] s_wallace_cska32_and_11_15;
  wire [0:0] s_wallace_cska32_fa380_xor1;
  wire [0:0] s_wallace_cska32_fa380_or0;
  wire [0:0] s_wallace_cska32_and_13_14;
  wire [0:0] s_wallace_cska32_and_12_15;
  wire [0:0] s_wallace_cska32_fa381_xor1;
  wire [0:0] s_wallace_cska32_fa381_or0;
  wire [0:0] s_wallace_cska32_and_14_14;
  wire [0:0] s_wallace_cska32_and_13_15;
  wire [0:0] s_wallace_cska32_fa382_xor1;
  wire [0:0] s_wallace_cska32_fa382_or0;
  wire [0:0] s_wallace_cska32_and_15_14;
  wire [0:0] s_wallace_cska32_and_14_15;
  wire [0:0] s_wallace_cska32_fa383_xor1;
  wire [0:0] s_wallace_cska32_fa383_or0;
  wire [0:0] s_wallace_cska32_and_16_14;
  wire [0:0] s_wallace_cska32_and_15_15;
  wire [0:0] s_wallace_cska32_fa384_xor1;
  wire [0:0] s_wallace_cska32_fa384_or0;
  wire [0:0] s_wallace_cska32_and_17_14;
  wire [0:0] s_wallace_cska32_and_16_15;
  wire [0:0] s_wallace_cska32_fa385_xor1;
  wire [0:0] s_wallace_cska32_fa385_or0;
  wire [0:0] s_wallace_cska32_and_18_14;
  wire [0:0] s_wallace_cska32_and_17_15;
  wire [0:0] s_wallace_cska32_fa386_xor1;
  wire [0:0] s_wallace_cska32_fa386_or0;
  wire [0:0] s_wallace_cska32_and_17_16;
  wire [0:0] s_wallace_cska32_and_16_17;
  wire [0:0] s_wallace_cska32_fa387_xor1;
  wire [0:0] s_wallace_cska32_fa387_or0;
  wire [0:0] s_wallace_cska32_and_17_17;
  wire [0:0] s_wallace_cska32_and_16_18;
  wire [0:0] s_wallace_cska32_fa388_xor1;
  wire [0:0] s_wallace_cska32_fa388_or0;
  wire [0:0] s_wallace_cska32_and_17_18;
  wire [0:0] s_wallace_cska32_and_16_19;
  wire [0:0] s_wallace_cska32_fa389_xor1;
  wire [0:0] s_wallace_cska32_fa389_or0;
  wire [0:0] s_wallace_cska32_and_17_19;
  wire [0:0] s_wallace_cska32_and_16_20;
  wire [0:0] s_wallace_cska32_fa390_xor1;
  wire [0:0] s_wallace_cska32_fa390_or0;
  wire [0:0] s_wallace_cska32_and_17_20;
  wire [0:0] s_wallace_cska32_and_16_21;
  wire [0:0] s_wallace_cska32_fa391_xor1;
  wire [0:0] s_wallace_cska32_fa391_or0;
  wire [0:0] s_wallace_cska32_and_17_21;
  wire [0:0] s_wallace_cska32_and_16_22;
  wire [0:0] s_wallace_cska32_fa392_xor1;
  wire [0:0] s_wallace_cska32_fa392_or0;
  wire [0:0] s_wallace_cska32_and_17_22;
  wire [0:0] s_wallace_cska32_and_16_23;
  wire [0:0] s_wallace_cska32_fa393_xor1;
  wire [0:0] s_wallace_cska32_fa393_or0;
  wire [0:0] s_wallace_cska32_and_17_23;
  wire [0:0] s_wallace_cska32_and_16_24;
  wire [0:0] s_wallace_cska32_fa394_xor1;
  wire [0:0] s_wallace_cska32_fa394_or0;
  wire [0:0] s_wallace_cska32_and_17_24;
  wire [0:0] s_wallace_cska32_and_16_25;
  wire [0:0] s_wallace_cska32_fa395_xor1;
  wire [0:0] s_wallace_cska32_fa395_or0;
  wire [0:0] s_wallace_cska32_and_17_25;
  wire [0:0] s_wallace_cska32_and_16_26;
  wire [0:0] s_wallace_cska32_fa396_xor1;
  wire [0:0] s_wallace_cska32_fa396_or0;
  wire [0:0] s_wallace_cska32_and_17_26;
  wire [0:0] s_wallace_cska32_and_16_27;
  wire [0:0] s_wallace_cska32_fa397_xor1;
  wire [0:0] s_wallace_cska32_fa397_or0;
  wire [0:0] s_wallace_cska32_and_17_27;
  wire [0:0] s_wallace_cska32_and_16_28;
  wire [0:0] s_wallace_cska32_fa398_xor1;
  wire [0:0] s_wallace_cska32_fa398_or0;
  wire [0:0] s_wallace_cska32_and_17_28;
  wire [0:0] s_wallace_cska32_and_16_29;
  wire [0:0] s_wallace_cska32_fa399_xor1;
  wire [0:0] s_wallace_cska32_fa399_or0;
  wire [0:0] s_wallace_cska32_and_17_29;
  wire [0:0] s_wallace_cska32_and_16_30;
  wire [0:0] s_wallace_cska32_fa400_xor1;
  wire [0:0] s_wallace_cska32_fa400_or0;
  wire [0:0] s_wallace_cska32_and_17_30;
  wire [0:0] s_wallace_cska32_nand_16_31;
  wire [0:0] s_wallace_cska32_fa401_xor1;
  wire [0:0] s_wallace_cska32_fa401_or0;
  wire [0:0] s_wallace_cska32_nand_17_31;
  wire [0:0] s_wallace_cska32_fa402_xor1;
  wire [0:0] s_wallace_cska32_fa402_or0;
  wire [0:0] s_wallace_cska32_fa403_xor1;
  wire [0:0] s_wallace_cska32_fa403_or0;
  wire [0:0] s_wallace_cska32_fa404_xor1;
  wire [0:0] s_wallace_cska32_fa404_or0;
  wire [0:0] s_wallace_cska32_fa405_xor1;
  wire [0:0] s_wallace_cska32_fa405_or0;
  wire [0:0] s_wallace_cska32_fa406_xor1;
  wire [0:0] s_wallace_cska32_fa406_or0;
  wire [0:0] s_wallace_cska32_fa407_xor1;
  wire [0:0] s_wallace_cska32_fa407_or0;
  wire [0:0] s_wallace_cska32_ha8_xor0;
  wire [0:0] s_wallace_cska32_ha8_and0;
  wire [0:0] s_wallace_cska32_fa408_xor1;
  wire [0:0] s_wallace_cska32_fa408_or0;
  wire [0:0] s_wallace_cska32_fa409_xor1;
  wire [0:0] s_wallace_cska32_fa409_or0;
  wire [0:0] s_wallace_cska32_fa410_xor1;
  wire [0:0] s_wallace_cska32_fa410_or0;
  wire [0:0] s_wallace_cska32_fa411_xor1;
  wire [0:0] s_wallace_cska32_fa411_or0;
  wire [0:0] s_wallace_cska32_fa412_xor1;
  wire [0:0] s_wallace_cska32_fa412_or0;
  wire [0:0] s_wallace_cska32_and_0_16;
  wire [0:0] s_wallace_cska32_fa413_xor1;
  wire [0:0] s_wallace_cska32_fa413_or0;
  wire [0:0] s_wallace_cska32_and_1_16;
  wire [0:0] s_wallace_cska32_and_0_17;
  wire [0:0] s_wallace_cska32_fa414_xor1;
  wire [0:0] s_wallace_cska32_fa414_or0;
  wire [0:0] s_wallace_cska32_and_2_16;
  wire [0:0] s_wallace_cska32_and_1_17;
  wire [0:0] s_wallace_cska32_fa415_xor1;
  wire [0:0] s_wallace_cska32_fa415_or0;
  wire [0:0] s_wallace_cska32_and_3_16;
  wire [0:0] s_wallace_cska32_and_2_17;
  wire [0:0] s_wallace_cska32_fa416_xor1;
  wire [0:0] s_wallace_cska32_fa416_or0;
  wire [0:0] s_wallace_cska32_and_4_16;
  wire [0:0] s_wallace_cska32_and_3_17;
  wire [0:0] s_wallace_cska32_fa417_xor1;
  wire [0:0] s_wallace_cska32_fa417_or0;
  wire [0:0] s_wallace_cska32_and_5_16;
  wire [0:0] s_wallace_cska32_and_4_17;
  wire [0:0] s_wallace_cska32_fa418_xor1;
  wire [0:0] s_wallace_cska32_fa418_or0;
  wire [0:0] s_wallace_cska32_and_6_16;
  wire [0:0] s_wallace_cska32_and_5_17;
  wire [0:0] s_wallace_cska32_fa419_xor1;
  wire [0:0] s_wallace_cska32_fa419_or0;
  wire [0:0] s_wallace_cska32_and_7_16;
  wire [0:0] s_wallace_cska32_and_6_17;
  wire [0:0] s_wallace_cska32_fa420_xor1;
  wire [0:0] s_wallace_cska32_fa420_or0;
  wire [0:0] s_wallace_cska32_and_8_16;
  wire [0:0] s_wallace_cska32_and_7_17;
  wire [0:0] s_wallace_cska32_fa421_xor1;
  wire [0:0] s_wallace_cska32_fa421_or0;
  wire [0:0] s_wallace_cska32_and_9_16;
  wire [0:0] s_wallace_cska32_and_8_17;
  wire [0:0] s_wallace_cska32_fa422_xor1;
  wire [0:0] s_wallace_cska32_fa422_or0;
  wire [0:0] s_wallace_cska32_and_10_16;
  wire [0:0] s_wallace_cska32_and_9_17;
  wire [0:0] s_wallace_cska32_fa423_xor1;
  wire [0:0] s_wallace_cska32_fa423_or0;
  wire [0:0] s_wallace_cska32_and_11_16;
  wire [0:0] s_wallace_cska32_and_10_17;
  wire [0:0] s_wallace_cska32_fa424_xor1;
  wire [0:0] s_wallace_cska32_fa424_or0;
  wire [0:0] s_wallace_cska32_and_12_16;
  wire [0:0] s_wallace_cska32_and_11_17;
  wire [0:0] s_wallace_cska32_fa425_xor1;
  wire [0:0] s_wallace_cska32_fa425_or0;
  wire [0:0] s_wallace_cska32_and_13_16;
  wire [0:0] s_wallace_cska32_and_12_17;
  wire [0:0] s_wallace_cska32_fa426_xor1;
  wire [0:0] s_wallace_cska32_fa426_or0;
  wire [0:0] s_wallace_cska32_and_14_16;
  wire [0:0] s_wallace_cska32_and_13_17;
  wire [0:0] s_wallace_cska32_fa427_xor1;
  wire [0:0] s_wallace_cska32_fa427_or0;
  wire [0:0] s_wallace_cska32_and_15_16;
  wire [0:0] s_wallace_cska32_and_14_17;
  wire [0:0] s_wallace_cska32_fa428_xor1;
  wire [0:0] s_wallace_cska32_fa428_or0;
  wire [0:0] s_wallace_cska32_and_16_16;
  wire [0:0] s_wallace_cska32_and_15_17;
  wire [0:0] s_wallace_cska32_fa429_xor1;
  wire [0:0] s_wallace_cska32_fa429_or0;
  wire [0:0] s_wallace_cska32_and_15_18;
  wire [0:0] s_wallace_cska32_and_14_19;
  wire [0:0] s_wallace_cska32_fa430_xor1;
  wire [0:0] s_wallace_cska32_fa430_or0;
  wire [0:0] s_wallace_cska32_and_15_19;
  wire [0:0] s_wallace_cska32_and_14_20;
  wire [0:0] s_wallace_cska32_fa431_xor1;
  wire [0:0] s_wallace_cska32_fa431_or0;
  wire [0:0] s_wallace_cska32_and_15_20;
  wire [0:0] s_wallace_cska32_and_14_21;
  wire [0:0] s_wallace_cska32_fa432_xor1;
  wire [0:0] s_wallace_cska32_fa432_or0;
  wire [0:0] s_wallace_cska32_and_15_21;
  wire [0:0] s_wallace_cska32_and_14_22;
  wire [0:0] s_wallace_cska32_fa433_xor1;
  wire [0:0] s_wallace_cska32_fa433_or0;
  wire [0:0] s_wallace_cska32_and_15_22;
  wire [0:0] s_wallace_cska32_and_14_23;
  wire [0:0] s_wallace_cska32_fa434_xor1;
  wire [0:0] s_wallace_cska32_fa434_or0;
  wire [0:0] s_wallace_cska32_and_15_23;
  wire [0:0] s_wallace_cska32_and_14_24;
  wire [0:0] s_wallace_cska32_fa435_xor1;
  wire [0:0] s_wallace_cska32_fa435_or0;
  wire [0:0] s_wallace_cska32_and_15_24;
  wire [0:0] s_wallace_cska32_and_14_25;
  wire [0:0] s_wallace_cska32_fa436_xor1;
  wire [0:0] s_wallace_cska32_fa436_or0;
  wire [0:0] s_wallace_cska32_and_15_25;
  wire [0:0] s_wallace_cska32_and_14_26;
  wire [0:0] s_wallace_cska32_fa437_xor1;
  wire [0:0] s_wallace_cska32_fa437_or0;
  wire [0:0] s_wallace_cska32_and_15_26;
  wire [0:0] s_wallace_cska32_and_14_27;
  wire [0:0] s_wallace_cska32_fa438_xor1;
  wire [0:0] s_wallace_cska32_fa438_or0;
  wire [0:0] s_wallace_cska32_and_15_27;
  wire [0:0] s_wallace_cska32_and_14_28;
  wire [0:0] s_wallace_cska32_fa439_xor1;
  wire [0:0] s_wallace_cska32_fa439_or0;
  wire [0:0] s_wallace_cska32_and_15_28;
  wire [0:0] s_wallace_cska32_and_14_29;
  wire [0:0] s_wallace_cska32_fa440_xor1;
  wire [0:0] s_wallace_cska32_fa440_or0;
  wire [0:0] s_wallace_cska32_and_15_29;
  wire [0:0] s_wallace_cska32_and_14_30;
  wire [0:0] s_wallace_cska32_fa441_xor1;
  wire [0:0] s_wallace_cska32_fa441_or0;
  wire [0:0] s_wallace_cska32_and_15_30;
  wire [0:0] s_wallace_cska32_nand_14_31;
  wire [0:0] s_wallace_cska32_fa442_xor1;
  wire [0:0] s_wallace_cska32_fa442_or0;
  wire [0:0] s_wallace_cska32_nand_15_31;
  wire [0:0] s_wallace_cska32_fa443_xor1;
  wire [0:0] s_wallace_cska32_fa443_or0;
  wire [0:0] s_wallace_cska32_fa444_xor1;
  wire [0:0] s_wallace_cska32_fa444_or0;
  wire [0:0] s_wallace_cska32_fa445_xor1;
  wire [0:0] s_wallace_cska32_fa445_or0;
  wire [0:0] s_wallace_cska32_fa446_xor1;
  wire [0:0] s_wallace_cska32_fa446_or0;
  wire [0:0] s_wallace_cska32_fa447_xor1;
  wire [0:0] s_wallace_cska32_fa447_or0;
  wire [0:0] s_wallace_cska32_fa448_xor1;
  wire [0:0] s_wallace_cska32_fa448_or0;
  wire [0:0] s_wallace_cska32_fa449_xor1;
  wire [0:0] s_wallace_cska32_fa449_or0;
  wire [0:0] s_wallace_cska32_ha9_xor0;
  wire [0:0] s_wallace_cska32_ha9_and0;
  wire [0:0] s_wallace_cska32_fa450_xor1;
  wire [0:0] s_wallace_cska32_fa450_or0;
  wire [0:0] s_wallace_cska32_fa451_xor1;
  wire [0:0] s_wallace_cska32_fa451_or0;
  wire [0:0] s_wallace_cska32_fa452_xor1;
  wire [0:0] s_wallace_cska32_fa452_or0;
  wire [0:0] s_wallace_cska32_fa453_xor1;
  wire [0:0] s_wallace_cska32_fa453_or0;
  wire [0:0] s_wallace_cska32_fa454_xor1;
  wire [0:0] s_wallace_cska32_fa454_or0;
  wire [0:0] s_wallace_cska32_fa455_xor1;
  wire [0:0] s_wallace_cska32_fa455_or0;
  wire [0:0] s_wallace_cska32_and_0_18;
  wire [0:0] s_wallace_cska32_fa456_xor1;
  wire [0:0] s_wallace_cska32_fa456_or0;
  wire [0:0] s_wallace_cska32_and_1_18;
  wire [0:0] s_wallace_cska32_and_0_19;
  wire [0:0] s_wallace_cska32_fa457_xor1;
  wire [0:0] s_wallace_cska32_fa457_or0;
  wire [0:0] s_wallace_cska32_and_2_18;
  wire [0:0] s_wallace_cska32_and_1_19;
  wire [0:0] s_wallace_cska32_fa458_xor1;
  wire [0:0] s_wallace_cska32_fa458_or0;
  wire [0:0] s_wallace_cska32_and_3_18;
  wire [0:0] s_wallace_cska32_and_2_19;
  wire [0:0] s_wallace_cska32_fa459_xor1;
  wire [0:0] s_wallace_cska32_fa459_or0;
  wire [0:0] s_wallace_cska32_and_4_18;
  wire [0:0] s_wallace_cska32_and_3_19;
  wire [0:0] s_wallace_cska32_fa460_xor1;
  wire [0:0] s_wallace_cska32_fa460_or0;
  wire [0:0] s_wallace_cska32_and_5_18;
  wire [0:0] s_wallace_cska32_and_4_19;
  wire [0:0] s_wallace_cska32_fa461_xor1;
  wire [0:0] s_wallace_cska32_fa461_or0;
  wire [0:0] s_wallace_cska32_and_6_18;
  wire [0:0] s_wallace_cska32_and_5_19;
  wire [0:0] s_wallace_cska32_fa462_xor1;
  wire [0:0] s_wallace_cska32_fa462_or0;
  wire [0:0] s_wallace_cska32_and_7_18;
  wire [0:0] s_wallace_cska32_and_6_19;
  wire [0:0] s_wallace_cska32_fa463_xor1;
  wire [0:0] s_wallace_cska32_fa463_or0;
  wire [0:0] s_wallace_cska32_and_8_18;
  wire [0:0] s_wallace_cska32_and_7_19;
  wire [0:0] s_wallace_cska32_fa464_xor1;
  wire [0:0] s_wallace_cska32_fa464_or0;
  wire [0:0] s_wallace_cska32_and_9_18;
  wire [0:0] s_wallace_cska32_and_8_19;
  wire [0:0] s_wallace_cska32_fa465_xor1;
  wire [0:0] s_wallace_cska32_fa465_or0;
  wire [0:0] s_wallace_cska32_and_10_18;
  wire [0:0] s_wallace_cska32_and_9_19;
  wire [0:0] s_wallace_cska32_fa466_xor1;
  wire [0:0] s_wallace_cska32_fa466_or0;
  wire [0:0] s_wallace_cska32_and_11_18;
  wire [0:0] s_wallace_cska32_and_10_19;
  wire [0:0] s_wallace_cska32_fa467_xor1;
  wire [0:0] s_wallace_cska32_fa467_or0;
  wire [0:0] s_wallace_cska32_and_12_18;
  wire [0:0] s_wallace_cska32_and_11_19;
  wire [0:0] s_wallace_cska32_fa468_xor1;
  wire [0:0] s_wallace_cska32_fa468_or0;
  wire [0:0] s_wallace_cska32_and_13_18;
  wire [0:0] s_wallace_cska32_and_12_19;
  wire [0:0] s_wallace_cska32_fa469_xor1;
  wire [0:0] s_wallace_cska32_fa469_or0;
  wire [0:0] s_wallace_cska32_and_14_18;
  wire [0:0] s_wallace_cska32_and_13_19;
  wire [0:0] s_wallace_cska32_fa470_xor1;
  wire [0:0] s_wallace_cska32_fa470_or0;
  wire [0:0] s_wallace_cska32_and_13_20;
  wire [0:0] s_wallace_cska32_and_12_21;
  wire [0:0] s_wallace_cska32_fa471_xor1;
  wire [0:0] s_wallace_cska32_fa471_or0;
  wire [0:0] s_wallace_cska32_and_13_21;
  wire [0:0] s_wallace_cska32_and_12_22;
  wire [0:0] s_wallace_cska32_fa472_xor1;
  wire [0:0] s_wallace_cska32_fa472_or0;
  wire [0:0] s_wallace_cska32_and_13_22;
  wire [0:0] s_wallace_cska32_and_12_23;
  wire [0:0] s_wallace_cska32_fa473_xor1;
  wire [0:0] s_wallace_cska32_fa473_or0;
  wire [0:0] s_wallace_cska32_and_13_23;
  wire [0:0] s_wallace_cska32_and_12_24;
  wire [0:0] s_wallace_cska32_fa474_xor1;
  wire [0:0] s_wallace_cska32_fa474_or0;
  wire [0:0] s_wallace_cska32_and_13_24;
  wire [0:0] s_wallace_cska32_and_12_25;
  wire [0:0] s_wallace_cska32_fa475_xor1;
  wire [0:0] s_wallace_cska32_fa475_or0;
  wire [0:0] s_wallace_cska32_and_13_25;
  wire [0:0] s_wallace_cska32_and_12_26;
  wire [0:0] s_wallace_cska32_fa476_xor1;
  wire [0:0] s_wallace_cska32_fa476_or0;
  wire [0:0] s_wallace_cska32_and_13_26;
  wire [0:0] s_wallace_cska32_and_12_27;
  wire [0:0] s_wallace_cska32_fa477_xor1;
  wire [0:0] s_wallace_cska32_fa477_or0;
  wire [0:0] s_wallace_cska32_and_13_27;
  wire [0:0] s_wallace_cska32_and_12_28;
  wire [0:0] s_wallace_cska32_fa478_xor1;
  wire [0:0] s_wallace_cska32_fa478_or0;
  wire [0:0] s_wallace_cska32_and_13_28;
  wire [0:0] s_wallace_cska32_and_12_29;
  wire [0:0] s_wallace_cska32_fa479_xor1;
  wire [0:0] s_wallace_cska32_fa479_or0;
  wire [0:0] s_wallace_cska32_and_13_29;
  wire [0:0] s_wallace_cska32_and_12_30;
  wire [0:0] s_wallace_cska32_fa480_xor1;
  wire [0:0] s_wallace_cska32_fa480_or0;
  wire [0:0] s_wallace_cska32_and_13_30;
  wire [0:0] s_wallace_cska32_nand_12_31;
  wire [0:0] s_wallace_cska32_fa481_xor1;
  wire [0:0] s_wallace_cska32_fa481_or0;
  wire [0:0] s_wallace_cska32_nand_13_31;
  wire [0:0] s_wallace_cska32_fa482_xor1;
  wire [0:0] s_wallace_cska32_fa482_or0;
  wire [0:0] s_wallace_cska32_fa483_xor1;
  wire [0:0] s_wallace_cska32_fa483_or0;
  wire [0:0] s_wallace_cska32_fa484_xor1;
  wire [0:0] s_wallace_cska32_fa484_or0;
  wire [0:0] s_wallace_cska32_fa485_xor1;
  wire [0:0] s_wallace_cska32_fa485_or0;
  wire [0:0] s_wallace_cska32_fa486_xor1;
  wire [0:0] s_wallace_cska32_fa486_or0;
  wire [0:0] s_wallace_cska32_fa487_xor1;
  wire [0:0] s_wallace_cska32_fa487_or0;
  wire [0:0] s_wallace_cska32_fa488_xor1;
  wire [0:0] s_wallace_cska32_fa488_or0;
  wire [0:0] s_wallace_cska32_fa489_xor1;
  wire [0:0] s_wallace_cska32_fa489_or0;
  wire [0:0] s_wallace_cska32_ha10_xor0;
  wire [0:0] s_wallace_cska32_ha10_and0;
  wire [0:0] s_wallace_cska32_fa490_xor1;
  wire [0:0] s_wallace_cska32_fa490_or0;
  wire [0:0] s_wallace_cska32_fa491_xor1;
  wire [0:0] s_wallace_cska32_fa491_or0;
  wire [0:0] s_wallace_cska32_fa492_xor1;
  wire [0:0] s_wallace_cska32_fa492_or0;
  wire [0:0] s_wallace_cska32_fa493_xor1;
  wire [0:0] s_wallace_cska32_fa493_or0;
  wire [0:0] s_wallace_cska32_fa494_xor1;
  wire [0:0] s_wallace_cska32_fa494_or0;
  wire [0:0] s_wallace_cska32_fa495_xor1;
  wire [0:0] s_wallace_cska32_fa495_or0;
  wire [0:0] s_wallace_cska32_fa496_xor1;
  wire [0:0] s_wallace_cska32_fa496_or0;
  wire [0:0] s_wallace_cska32_and_0_20;
  wire [0:0] s_wallace_cska32_fa497_xor1;
  wire [0:0] s_wallace_cska32_fa497_or0;
  wire [0:0] s_wallace_cska32_and_1_20;
  wire [0:0] s_wallace_cska32_and_0_21;
  wire [0:0] s_wallace_cska32_fa498_xor1;
  wire [0:0] s_wallace_cska32_fa498_or0;
  wire [0:0] s_wallace_cska32_and_2_20;
  wire [0:0] s_wallace_cska32_and_1_21;
  wire [0:0] s_wallace_cska32_fa499_xor1;
  wire [0:0] s_wallace_cska32_fa499_or0;
  wire [0:0] s_wallace_cska32_and_3_20;
  wire [0:0] s_wallace_cska32_and_2_21;
  wire [0:0] s_wallace_cska32_fa500_xor1;
  wire [0:0] s_wallace_cska32_fa500_or0;
  wire [0:0] s_wallace_cska32_and_4_20;
  wire [0:0] s_wallace_cska32_and_3_21;
  wire [0:0] s_wallace_cska32_fa501_xor1;
  wire [0:0] s_wallace_cska32_fa501_or0;
  wire [0:0] s_wallace_cska32_and_5_20;
  wire [0:0] s_wallace_cska32_and_4_21;
  wire [0:0] s_wallace_cska32_fa502_xor1;
  wire [0:0] s_wallace_cska32_fa502_or0;
  wire [0:0] s_wallace_cska32_and_6_20;
  wire [0:0] s_wallace_cska32_and_5_21;
  wire [0:0] s_wallace_cska32_fa503_xor1;
  wire [0:0] s_wallace_cska32_fa503_or0;
  wire [0:0] s_wallace_cska32_and_7_20;
  wire [0:0] s_wallace_cska32_and_6_21;
  wire [0:0] s_wallace_cska32_fa504_xor1;
  wire [0:0] s_wallace_cska32_fa504_or0;
  wire [0:0] s_wallace_cska32_and_8_20;
  wire [0:0] s_wallace_cska32_and_7_21;
  wire [0:0] s_wallace_cska32_fa505_xor1;
  wire [0:0] s_wallace_cska32_fa505_or0;
  wire [0:0] s_wallace_cska32_and_9_20;
  wire [0:0] s_wallace_cska32_and_8_21;
  wire [0:0] s_wallace_cska32_fa506_xor1;
  wire [0:0] s_wallace_cska32_fa506_or0;
  wire [0:0] s_wallace_cska32_and_10_20;
  wire [0:0] s_wallace_cska32_and_9_21;
  wire [0:0] s_wallace_cska32_fa507_xor1;
  wire [0:0] s_wallace_cska32_fa507_or0;
  wire [0:0] s_wallace_cska32_and_11_20;
  wire [0:0] s_wallace_cska32_and_10_21;
  wire [0:0] s_wallace_cska32_fa508_xor1;
  wire [0:0] s_wallace_cska32_fa508_or0;
  wire [0:0] s_wallace_cska32_and_12_20;
  wire [0:0] s_wallace_cska32_and_11_21;
  wire [0:0] s_wallace_cska32_fa509_xor1;
  wire [0:0] s_wallace_cska32_fa509_or0;
  wire [0:0] s_wallace_cska32_and_11_22;
  wire [0:0] s_wallace_cska32_and_10_23;
  wire [0:0] s_wallace_cska32_fa510_xor1;
  wire [0:0] s_wallace_cska32_fa510_or0;
  wire [0:0] s_wallace_cska32_and_11_23;
  wire [0:0] s_wallace_cska32_and_10_24;
  wire [0:0] s_wallace_cska32_fa511_xor1;
  wire [0:0] s_wallace_cska32_fa511_or0;
  wire [0:0] s_wallace_cska32_and_11_24;
  wire [0:0] s_wallace_cska32_and_10_25;
  wire [0:0] s_wallace_cska32_fa512_xor1;
  wire [0:0] s_wallace_cska32_fa512_or0;
  wire [0:0] s_wallace_cska32_and_11_25;
  wire [0:0] s_wallace_cska32_and_10_26;
  wire [0:0] s_wallace_cska32_fa513_xor1;
  wire [0:0] s_wallace_cska32_fa513_or0;
  wire [0:0] s_wallace_cska32_and_11_26;
  wire [0:0] s_wallace_cska32_and_10_27;
  wire [0:0] s_wallace_cska32_fa514_xor1;
  wire [0:0] s_wallace_cska32_fa514_or0;
  wire [0:0] s_wallace_cska32_and_11_27;
  wire [0:0] s_wallace_cska32_and_10_28;
  wire [0:0] s_wallace_cska32_fa515_xor1;
  wire [0:0] s_wallace_cska32_fa515_or0;
  wire [0:0] s_wallace_cska32_and_11_28;
  wire [0:0] s_wallace_cska32_and_10_29;
  wire [0:0] s_wallace_cska32_fa516_xor1;
  wire [0:0] s_wallace_cska32_fa516_or0;
  wire [0:0] s_wallace_cska32_and_11_29;
  wire [0:0] s_wallace_cska32_and_10_30;
  wire [0:0] s_wallace_cska32_fa517_xor1;
  wire [0:0] s_wallace_cska32_fa517_or0;
  wire [0:0] s_wallace_cska32_and_11_30;
  wire [0:0] s_wallace_cska32_nand_10_31;
  wire [0:0] s_wallace_cska32_fa518_xor1;
  wire [0:0] s_wallace_cska32_fa518_or0;
  wire [0:0] s_wallace_cska32_nand_11_31;
  wire [0:0] s_wallace_cska32_fa519_xor1;
  wire [0:0] s_wallace_cska32_fa519_or0;
  wire [0:0] s_wallace_cska32_fa520_xor1;
  wire [0:0] s_wallace_cska32_fa520_or0;
  wire [0:0] s_wallace_cska32_fa521_xor1;
  wire [0:0] s_wallace_cska32_fa521_or0;
  wire [0:0] s_wallace_cska32_fa522_xor1;
  wire [0:0] s_wallace_cska32_fa522_or0;
  wire [0:0] s_wallace_cska32_fa523_xor1;
  wire [0:0] s_wallace_cska32_fa523_or0;
  wire [0:0] s_wallace_cska32_fa524_xor1;
  wire [0:0] s_wallace_cska32_fa524_or0;
  wire [0:0] s_wallace_cska32_fa525_xor1;
  wire [0:0] s_wallace_cska32_fa525_or0;
  wire [0:0] s_wallace_cska32_fa526_xor1;
  wire [0:0] s_wallace_cska32_fa526_or0;
  wire [0:0] s_wallace_cska32_fa527_xor1;
  wire [0:0] s_wallace_cska32_fa527_or0;
  wire [0:0] s_wallace_cska32_ha11_xor0;
  wire [0:0] s_wallace_cska32_ha11_and0;
  wire [0:0] s_wallace_cska32_fa528_xor1;
  wire [0:0] s_wallace_cska32_fa528_or0;
  wire [0:0] s_wallace_cska32_fa529_xor1;
  wire [0:0] s_wallace_cska32_fa529_or0;
  wire [0:0] s_wallace_cska32_fa530_xor1;
  wire [0:0] s_wallace_cska32_fa530_or0;
  wire [0:0] s_wallace_cska32_fa531_xor1;
  wire [0:0] s_wallace_cska32_fa531_or0;
  wire [0:0] s_wallace_cska32_fa532_xor1;
  wire [0:0] s_wallace_cska32_fa532_or0;
  wire [0:0] s_wallace_cska32_fa533_xor1;
  wire [0:0] s_wallace_cska32_fa533_or0;
  wire [0:0] s_wallace_cska32_fa534_xor1;
  wire [0:0] s_wallace_cska32_fa534_or0;
  wire [0:0] s_wallace_cska32_fa535_xor1;
  wire [0:0] s_wallace_cska32_fa535_or0;
  wire [0:0] s_wallace_cska32_and_0_22;
  wire [0:0] s_wallace_cska32_fa536_xor1;
  wire [0:0] s_wallace_cska32_fa536_or0;
  wire [0:0] s_wallace_cska32_and_1_22;
  wire [0:0] s_wallace_cska32_and_0_23;
  wire [0:0] s_wallace_cska32_fa537_xor1;
  wire [0:0] s_wallace_cska32_fa537_or0;
  wire [0:0] s_wallace_cska32_and_2_22;
  wire [0:0] s_wallace_cska32_and_1_23;
  wire [0:0] s_wallace_cska32_fa538_xor1;
  wire [0:0] s_wallace_cska32_fa538_or0;
  wire [0:0] s_wallace_cska32_and_3_22;
  wire [0:0] s_wallace_cska32_and_2_23;
  wire [0:0] s_wallace_cska32_fa539_xor1;
  wire [0:0] s_wallace_cska32_fa539_or0;
  wire [0:0] s_wallace_cska32_and_4_22;
  wire [0:0] s_wallace_cska32_and_3_23;
  wire [0:0] s_wallace_cska32_fa540_xor1;
  wire [0:0] s_wallace_cska32_fa540_or0;
  wire [0:0] s_wallace_cska32_and_5_22;
  wire [0:0] s_wallace_cska32_and_4_23;
  wire [0:0] s_wallace_cska32_fa541_xor1;
  wire [0:0] s_wallace_cska32_fa541_or0;
  wire [0:0] s_wallace_cska32_and_6_22;
  wire [0:0] s_wallace_cska32_and_5_23;
  wire [0:0] s_wallace_cska32_fa542_xor1;
  wire [0:0] s_wallace_cska32_fa542_or0;
  wire [0:0] s_wallace_cska32_and_7_22;
  wire [0:0] s_wallace_cska32_and_6_23;
  wire [0:0] s_wallace_cska32_fa543_xor1;
  wire [0:0] s_wallace_cska32_fa543_or0;
  wire [0:0] s_wallace_cska32_and_8_22;
  wire [0:0] s_wallace_cska32_and_7_23;
  wire [0:0] s_wallace_cska32_fa544_xor1;
  wire [0:0] s_wallace_cska32_fa544_or0;
  wire [0:0] s_wallace_cska32_and_9_22;
  wire [0:0] s_wallace_cska32_and_8_23;
  wire [0:0] s_wallace_cska32_fa545_xor1;
  wire [0:0] s_wallace_cska32_fa545_or0;
  wire [0:0] s_wallace_cska32_and_10_22;
  wire [0:0] s_wallace_cska32_and_9_23;
  wire [0:0] s_wallace_cska32_fa546_xor1;
  wire [0:0] s_wallace_cska32_fa546_or0;
  wire [0:0] s_wallace_cska32_and_9_24;
  wire [0:0] s_wallace_cska32_and_8_25;
  wire [0:0] s_wallace_cska32_fa547_xor1;
  wire [0:0] s_wallace_cska32_fa547_or0;
  wire [0:0] s_wallace_cska32_and_9_25;
  wire [0:0] s_wallace_cska32_and_8_26;
  wire [0:0] s_wallace_cska32_fa548_xor1;
  wire [0:0] s_wallace_cska32_fa548_or0;
  wire [0:0] s_wallace_cska32_and_9_26;
  wire [0:0] s_wallace_cska32_and_8_27;
  wire [0:0] s_wallace_cska32_fa549_xor1;
  wire [0:0] s_wallace_cska32_fa549_or0;
  wire [0:0] s_wallace_cska32_and_9_27;
  wire [0:0] s_wallace_cska32_and_8_28;
  wire [0:0] s_wallace_cska32_fa550_xor1;
  wire [0:0] s_wallace_cska32_fa550_or0;
  wire [0:0] s_wallace_cska32_and_9_28;
  wire [0:0] s_wallace_cska32_and_8_29;
  wire [0:0] s_wallace_cska32_fa551_xor1;
  wire [0:0] s_wallace_cska32_fa551_or0;
  wire [0:0] s_wallace_cska32_and_9_29;
  wire [0:0] s_wallace_cska32_and_8_30;
  wire [0:0] s_wallace_cska32_fa552_xor1;
  wire [0:0] s_wallace_cska32_fa552_or0;
  wire [0:0] s_wallace_cska32_and_9_30;
  wire [0:0] s_wallace_cska32_nand_8_31;
  wire [0:0] s_wallace_cska32_fa553_xor1;
  wire [0:0] s_wallace_cska32_fa553_or0;
  wire [0:0] s_wallace_cska32_nand_9_31;
  wire [0:0] s_wallace_cska32_fa554_xor1;
  wire [0:0] s_wallace_cska32_fa554_or0;
  wire [0:0] s_wallace_cska32_fa555_xor1;
  wire [0:0] s_wallace_cska32_fa555_or0;
  wire [0:0] s_wallace_cska32_fa556_xor1;
  wire [0:0] s_wallace_cska32_fa556_or0;
  wire [0:0] s_wallace_cska32_fa557_xor1;
  wire [0:0] s_wallace_cska32_fa557_or0;
  wire [0:0] s_wallace_cska32_fa558_xor1;
  wire [0:0] s_wallace_cska32_fa558_or0;
  wire [0:0] s_wallace_cska32_fa559_xor1;
  wire [0:0] s_wallace_cska32_fa559_or0;
  wire [0:0] s_wallace_cska32_fa560_xor1;
  wire [0:0] s_wallace_cska32_fa560_or0;
  wire [0:0] s_wallace_cska32_fa561_xor1;
  wire [0:0] s_wallace_cska32_fa561_or0;
  wire [0:0] s_wallace_cska32_fa562_xor1;
  wire [0:0] s_wallace_cska32_fa562_or0;
  wire [0:0] s_wallace_cska32_fa563_xor1;
  wire [0:0] s_wallace_cska32_fa563_or0;
  wire [0:0] s_wallace_cska32_ha12_xor0;
  wire [0:0] s_wallace_cska32_ha12_and0;
  wire [0:0] s_wallace_cska32_fa564_xor1;
  wire [0:0] s_wallace_cska32_fa564_or0;
  wire [0:0] s_wallace_cska32_fa565_xor1;
  wire [0:0] s_wallace_cska32_fa565_or0;
  wire [0:0] s_wallace_cska32_fa566_xor1;
  wire [0:0] s_wallace_cska32_fa566_or0;
  wire [0:0] s_wallace_cska32_fa567_xor1;
  wire [0:0] s_wallace_cska32_fa567_or0;
  wire [0:0] s_wallace_cska32_fa568_xor1;
  wire [0:0] s_wallace_cska32_fa568_or0;
  wire [0:0] s_wallace_cska32_fa569_xor1;
  wire [0:0] s_wallace_cska32_fa569_or0;
  wire [0:0] s_wallace_cska32_fa570_xor1;
  wire [0:0] s_wallace_cska32_fa570_or0;
  wire [0:0] s_wallace_cska32_fa571_xor1;
  wire [0:0] s_wallace_cska32_fa571_or0;
  wire [0:0] s_wallace_cska32_fa572_xor1;
  wire [0:0] s_wallace_cska32_fa572_or0;
  wire [0:0] s_wallace_cska32_and_0_24;
  wire [0:0] s_wallace_cska32_fa573_xor1;
  wire [0:0] s_wallace_cska32_fa573_or0;
  wire [0:0] s_wallace_cska32_and_1_24;
  wire [0:0] s_wallace_cska32_and_0_25;
  wire [0:0] s_wallace_cska32_fa574_xor1;
  wire [0:0] s_wallace_cska32_fa574_or0;
  wire [0:0] s_wallace_cska32_and_2_24;
  wire [0:0] s_wallace_cska32_and_1_25;
  wire [0:0] s_wallace_cska32_fa575_xor1;
  wire [0:0] s_wallace_cska32_fa575_or0;
  wire [0:0] s_wallace_cska32_and_3_24;
  wire [0:0] s_wallace_cska32_and_2_25;
  wire [0:0] s_wallace_cska32_fa576_xor1;
  wire [0:0] s_wallace_cska32_fa576_or0;
  wire [0:0] s_wallace_cska32_and_4_24;
  wire [0:0] s_wallace_cska32_and_3_25;
  wire [0:0] s_wallace_cska32_fa577_xor1;
  wire [0:0] s_wallace_cska32_fa577_or0;
  wire [0:0] s_wallace_cska32_and_5_24;
  wire [0:0] s_wallace_cska32_and_4_25;
  wire [0:0] s_wallace_cska32_fa578_xor1;
  wire [0:0] s_wallace_cska32_fa578_or0;
  wire [0:0] s_wallace_cska32_and_6_24;
  wire [0:0] s_wallace_cska32_and_5_25;
  wire [0:0] s_wallace_cska32_fa579_xor1;
  wire [0:0] s_wallace_cska32_fa579_or0;
  wire [0:0] s_wallace_cska32_and_7_24;
  wire [0:0] s_wallace_cska32_and_6_25;
  wire [0:0] s_wallace_cska32_fa580_xor1;
  wire [0:0] s_wallace_cska32_fa580_or0;
  wire [0:0] s_wallace_cska32_and_8_24;
  wire [0:0] s_wallace_cska32_and_7_25;
  wire [0:0] s_wallace_cska32_fa581_xor1;
  wire [0:0] s_wallace_cska32_fa581_or0;
  wire [0:0] s_wallace_cska32_and_7_26;
  wire [0:0] s_wallace_cska32_and_6_27;
  wire [0:0] s_wallace_cska32_fa582_xor1;
  wire [0:0] s_wallace_cska32_fa582_or0;
  wire [0:0] s_wallace_cska32_and_7_27;
  wire [0:0] s_wallace_cska32_and_6_28;
  wire [0:0] s_wallace_cska32_fa583_xor1;
  wire [0:0] s_wallace_cska32_fa583_or0;
  wire [0:0] s_wallace_cska32_and_7_28;
  wire [0:0] s_wallace_cska32_and_6_29;
  wire [0:0] s_wallace_cska32_fa584_xor1;
  wire [0:0] s_wallace_cska32_fa584_or0;
  wire [0:0] s_wallace_cska32_and_7_29;
  wire [0:0] s_wallace_cska32_and_6_30;
  wire [0:0] s_wallace_cska32_fa585_xor1;
  wire [0:0] s_wallace_cska32_fa585_or0;
  wire [0:0] s_wallace_cska32_and_7_30;
  wire [0:0] s_wallace_cska32_nand_6_31;
  wire [0:0] s_wallace_cska32_fa586_xor1;
  wire [0:0] s_wallace_cska32_fa586_or0;
  wire [0:0] s_wallace_cska32_nand_7_31;
  wire [0:0] s_wallace_cska32_fa587_xor1;
  wire [0:0] s_wallace_cska32_fa587_or0;
  wire [0:0] s_wallace_cska32_fa588_xor1;
  wire [0:0] s_wallace_cska32_fa588_or0;
  wire [0:0] s_wallace_cska32_fa589_xor1;
  wire [0:0] s_wallace_cska32_fa589_or0;
  wire [0:0] s_wallace_cska32_fa590_xor1;
  wire [0:0] s_wallace_cska32_fa590_or0;
  wire [0:0] s_wallace_cska32_fa591_xor1;
  wire [0:0] s_wallace_cska32_fa591_or0;
  wire [0:0] s_wallace_cska32_fa592_xor1;
  wire [0:0] s_wallace_cska32_fa592_or0;
  wire [0:0] s_wallace_cska32_fa593_xor1;
  wire [0:0] s_wallace_cska32_fa593_or0;
  wire [0:0] s_wallace_cska32_fa594_xor1;
  wire [0:0] s_wallace_cska32_fa594_or0;
  wire [0:0] s_wallace_cska32_fa595_xor1;
  wire [0:0] s_wallace_cska32_fa595_or0;
  wire [0:0] s_wallace_cska32_fa596_xor1;
  wire [0:0] s_wallace_cska32_fa596_or0;
  wire [0:0] s_wallace_cska32_fa597_xor1;
  wire [0:0] s_wallace_cska32_fa597_or0;
  wire [0:0] s_wallace_cska32_ha13_xor0;
  wire [0:0] s_wallace_cska32_ha13_and0;
  wire [0:0] s_wallace_cska32_fa598_xor1;
  wire [0:0] s_wallace_cska32_fa598_or0;
  wire [0:0] s_wallace_cska32_fa599_xor1;
  wire [0:0] s_wallace_cska32_fa599_or0;
  wire [0:0] s_wallace_cska32_fa600_xor1;
  wire [0:0] s_wallace_cska32_fa600_or0;
  wire [0:0] s_wallace_cska32_fa601_xor1;
  wire [0:0] s_wallace_cska32_fa601_or0;
  wire [0:0] s_wallace_cska32_fa602_xor1;
  wire [0:0] s_wallace_cska32_fa602_or0;
  wire [0:0] s_wallace_cska32_fa603_xor1;
  wire [0:0] s_wallace_cska32_fa603_or0;
  wire [0:0] s_wallace_cska32_fa604_xor1;
  wire [0:0] s_wallace_cska32_fa604_or0;
  wire [0:0] s_wallace_cska32_fa605_xor1;
  wire [0:0] s_wallace_cska32_fa605_or0;
  wire [0:0] s_wallace_cska32_fa606_xor1;
  wire [0:0] s_wallace_cska32_fa606_or0;
  wire [0:0] s_wallace_cska32_fa607_xor1;
  wire [0:0] s_wallace_cska32_fa607_or0;
  wire [0:0] s_wallace_cska32_and_0_26;
  wire [0:0] s_wallace_cska32_fa608_xor1;
  wire [0:0] s_wallace_cska32_fa608_or0;
  wire [0:0] s_wallace_cska32_and_1_26;
  wire [0:0] s_wallace_cska32_and_0_27;
  wire [0:0] s_wallace_cska32_fa609_xor1;
  wire [0:0] s_wallace_cska32_fa609_or0;
  wire [0:0] s_wallace_cska32_and_2_26;
  wire [0:0] s_wallace_cska32_and_1_27;
  wire [0:0] s_wallace_cska32_fa610_xor1;
  wire [0:0] s_wallace_cska32_fa610_or0;
  wire [0:0] s_wallace_cska32_and_3_26;
  wire [0:0] s_wallace_cska32_and_2_27;
  wire [0:0] s_wallace_cska32_fa611_xor1;
  wire [0:0] s_wallace_cska32_fa611_or0;
  wire [0:0] s_wallace_cska32_and_4_26;
  wire [0:0] s_wallace_cska32_and_3_27;
  wire [0:0] s_wallace_cska32_fa612_xor1;
  wire [0:0] s_wallace_cska32_fa612_or0;
  wire [0:0] s_wallace_cska32_and_5_26;
  wire [0:0] s_wallace_cska32_and_4_27;
  wire [0:0] s_wallace_cska32_fa613_xor1;
  wire [0:0] s_wallace_cska32_fa613_or0;
  wire [0:0] s_wallace_cska32_and_6_26;
  wire [0:0] s_wallace_cska32_and_5_27;
  wire [0:0] s_wallace_cska32_fa614_xor1;
  wire [0:0] s_wallace_cska32_fa614_or0;
  wire [0:0] s_wallace_cska32_and_5_28;
  wire [0:0] s_wallace_cska32_and_4_29;
  wire [0:0] s_wallace_cska32_fa615_xor1;
  wire [0:0] s_wallace_cska32_fa615_or0;
  wire [0:0] s_wallace_cska32_and_5_29;
  wire [0:0] s_wallace_cska32_and_4_30;
  wire [0:0] s_wallace_cska32_fa616_xor1;
  wire [0:0] s_wallace_cska32_fa616_or0;
  wire [0:0] s_wallace_cska32_and_5_30;
  wire [0:0] s_wallace_cska32_nand_4_31;
  wire [0:0] s_wallace_cska32_fa617_xor1;
  wire [0:0] s_wallace_cska32_fa617_or0;
  wire [0:0] s_wallace_cska32_nand_5_31;
  wire [0:0] s_wallace_cska32_fa618_xor1;
  wire [0:0] s_wallace_cska32_fa618_or0;
  wire [0:0] s_wallace_cska32_fa619_xor1;
  wire [0:0] s_wallace_cska32_fa619_or0;
  wire [0:0] s_wallace_cska32_fa620_xor1;
  wire [0:0] s_wallace_cska32_fa620_or0;
  wire [0:0] s_wallace_cska32_fa621_xor1;
  wire [0:0] s_wallace_cska32_fa621_or0;
  wire [0:0] s_wallace_cska32_fa622_xor1;
  wire [0:0] s_wallace_cska32_fa622_or0;
  wire [0:0] s_wallace_cska32_fa623_xor1;
  wire [0:0] s_wallace_cska32_fa623_or0;
  wire [0:0] s_wallace_cska32_fa624_xor1;
  wire [0:0] s_wallace_cska32_fa624_or0;
  wire [0:0] s_wallace_cska32_fa625_xor1;
  wire [0:0] s_wallace_cska32_fa625_or0;
  wire [0:0] s_wallace_cska32_fa626_xor1;
  wire [0:0] s_wallace_cska32_fa626_or0;
  wire [0:0] s_wallace_cska32_fa627_xor1;
  wire [0:0] s_wallace_cska32_fa627_or0;
  wire [0:0] s_wallace_cska32_fa628_xor1;
  wire [0:0] s_wallace_cska32_fa628_or0;
  wire [0:0] s_wallace_cska32_fa629_xor1;
  wire [0:0] s_wallace_cska32_fa629_or0;
  wire [0:0] s_wallace_cska32_ha14_xor0;
  wire [0:0] s_wallace_cska32_ha14_and0;
  wire [0:0] s_wallace_cska32_fa630_xor1;
  wire [0:0] s_wallace_cska32_fa630_or0;
  wire [0:0] s_wallace_cska32_fa631_xor1;
  wire [0:0] s_wallace_cska32_fa631_or0;
  wire [0:0] s_wallace_cska32_fa632_xor1;
  wire [0:0] s_wallace_cska32_fa632_or0;
  wire [0:0] s_wallace_cska32_fa633_xor1;
  wire [0:0] s_wallace_cska32_fa633_or0;
  wire [0:0] s_wallace_cska32_fa634_xor1;
  wire [0:0] s_wallace_cska32_fa634_or0;
  wire [0:0] s_wallace_cska32_fa635_xor1;
  wire [0:0] s_wallace_cska32_fa635_or0;
  wire [0:0] s_wallace_cska32_fa636_xor1;
  wire [0:0] s_wallace_cska32_fa636_or0;
  wire [0:0] s_wallace_cska32_fa637_xor1;
  wire [0:0] s_wallace_cska32_fa637_or0;
  wire [0:0] s_wallace_cska32_fa638_xor1;
  wire [0:0] s_wallace_cska32_fa638_or0;
  wire [0:0] s_wallace_cska32_fa639_xor1;
  wire [0:0] s_wallace_cska32_fa639_or0;
  wire [0:0] s_wallace_cska32_fa640_xor1;
  wire [0:0] s_wallace_cska32_fa640_or0;
  wire [0:0] s_wallace_cska32_and_0_28;
  wire [0:0] s_wallace_cska32_fa641_xor1;
  wire [0:0] s_wallace_cska32_fa641_or0;
  wire [0:0] s_wallace_cska32_and_1_28;
  wire [0:0] s_wallace_cska32_and_0_29;
  wire [0:0] s_wallace_cska32_fa642_xor1;
  wire [0:0] s_wallace_cska32_fa642_or0;
  wire [0:0] s_wallace_cska32_and_2_28;
  wire [0:0] s_wallace_cska32_and_1_29;
  wire [0:0] s_wallace_cska32_fa643_xor1;
  wire [0:0] s_wallace_cska32_fa643_or0;
  wire [0:0] s_wallace_cska32_and_3_28;
  wire [0:0] s_wallace_cska32_and_2_29;
  wire [0:0] s_wallace_cska32_fa644_xor1;
  wire [0:0] s_wallace_cska32_fa644_or0;
  wire [0:0] s_wallace_cska32_and_4_28;
  wire [0:0] s_wallace_cska32_and_3_29;
  wire [0:0] s_wallace_cska32_fa645_xor1;
  wire [0:0] s_wallace_cska32_fa645_or0;
  wire [0:0] s_wallace_cska32_and_3_30;
  wire [0:0] s_wallace_cska32_nand_2_31;
  wire [0:0] s_wallace_cska32_fa646_xor1;
  wire [0:0] s_wallace_cska32_fa646_or0;
  wire [0:0] s_wallace_cska32_nand_3_31;
  wire [0:0] s_wallace_cska32_fa647_xor1;
  wire [0:0] s_wallace_cska32_fa647_or0;
  wire [0:0] s_wallace_cska32_fa648_xor1;
  wire [0:0] s_wallace_cska32_fa648_or0;
  wire [0:0] s_wallace_cska32_fa649_xor1;
  wire [0:0] s_wallace_cska32_fa649_or0;
  wire [0:0] s_wallace_cska32_fa650_xor1;
  wire [0:0] s_wallace_cska32_fa650_or0;
  wire [0:0] s_wallace_cska32_fa651_xor1;
  wire [0:0] s_wallace_cska32_fa651_or0;
  wire [0:0] s_wallace_cska32_fa652_xor1;
  wire [0:0] s_wallace_cska32_fa652_or0;
  wire [0:0] s_wallace_cska32_fa653_xor1;
  wire [0:0] s_wallace_cska32_fa653_or0;
  wire [0:0] s_wallace_cska32_fa654_xor1;
  wire [0:0] s_wallace_cska32_fa654_or0;
  wire [0:0] s_wallace_cska32_fa655_xor1;
  wire [0:0] s_wallace_cska32_fa655_or0;
  wire [0:0] s_wallace_cska32_fa656_xor1;
  wire [0:0] s_wallace_cska32_fa656_or0;
  wire [0:0] s_wallace_cska32_fa657_xor1;
  wire [0:0] s_wallace_cska32_fa657_or0;
  wire [0:0] s_wallace_cska32_fa658_xor1;
  wire [0:0] s_wallace_cska32_fa658_or0;
  wire [0:0] s_wallace_cska32_fa659_xor1;
  wire [0:0] s_wallace_cska32_fa659_or0;
  wire [0:0] s_wallace_cska32_ha15_xor0;
  wire [0:0] s_wallace_cska32_ha15_and0;
  wire [0:0] s_wallace_cska32_fa660_xor1;
  wire [0:0] s_wallace_cska32_fa660_or0;
  wire [0:0] s_wallace_cska32_fa661_xor1;
  wire [0:0] s_wallace_cska32_fa661_or0;
  wire [0:0] s_wallace_cska32_fa662_xor1;
  wire [0:0] s_wallace_cska32_fa662_or0;
  wire [0:0] s_wallace_cska32_fa663_xor1;
  wire [0:0] s_wallace_cska32_fa663_or0;
  wire [0:0] s_wallace_cska32_fa664_xor1;
  wire [0:0] s_wallace_cska32_fa664_or0;
  wire [0:0] s_wallace_cska32_fa665_xor1;
  wire [0:0] s_wallace_cska32_fa665_or0;
  wire [0:0] s_wallace_cska32_fa666_xor1;
  wire [0:0] s_wallace_cska32_fa666_or0;
  wire [0:0] s_wallace_cska32_fa667_xor1;
  wire [0:0] s_wallace_cska32_fa667_or0;
  wire [0:0] s_wallace_cska32_fa668_xor1;
  wire [0:0] s_wallace_cska32_fa668_or0;
  wire [0:0] s_wallace_cska32_fa669_xor1;
  wire [0:0] s_wallace_cska32_fa669_or0;
  wire [0:0] s_wallace_cska32_fa670_xor1;
  wire [0:0] s_wallace_cska32_fa670_or0;
  wire [0:0] s_wallace_cska32_fa671_xor1;
  wire [0:0] s_wallace_cska32_fa671_or0;
  wire [0:0] s_wallace_cska32_and_0_30;
  wire [0:0] s_wallace_cska32_fa672_xor1;
  wire [0:0] s_wallace_cska32_fa672_or0;
  wire [0:0] s_wallace_cska32_and_1_30;
  wire [0:0] s_wallace_cska32_nand_0_31;
  wire [0:0] s_wallace_cska32_fa673_xor1;
  wire [0:0] s_wallace_cska32_fa673_or0;
  wire [0:0] s_wallace_cska32_and_2_30;
  wire [0:0] s_wallace_cska32_nand_1_31;
  wire [0:0] s_wallace_cska32_fa674_xor1;
  wire [0:0] s_wallace_cska32_fa674_or0;
  wire [0:0] s_wallace_cska32_fa675_xor1;
  wire [0:0] s_wallace_cska32_fa675_or0;
  wire [0:0] s_wallace_cska32_fa676_xor1;
  wire [0:0] s_wallace_cska32_fa676_or0;
  wire [0:0] s_wallace_cska32_fa677_xor1;
  wire [0:0] s_wallace_cska32_fa677_or0;
  wire [0:0] s_wallace_cska32_fa678_xor1;
  wire [0:0] s_wallace_cska32_fa678_or0;
  wire [0:0] s_wallace_cska32_fa679_xor1;
  wire [0:0] s_wallace_cska32_fa679_or0;
  wire [0:0] s_wallace_cska32_fa680_xor1;
  wire [0:0] s_wallace_cska32_fa680_or0;
  wire [0:0] s_wallace_cska32_fa681_xor1;
  wire [0:0] s_wallace_cska32_fa681_or0;
  wire [0:0] s_wallace_cska32_fa682_xor1;
  wire [0:0] s_wallace_cska32_fa682_or0;
  wire [0:0] s_wallace_cska32_fa683_xor1;
  wire [0:0] s_wallace_cska32_fa683_or0;
  wire [0:0] s_wallace_cska32_fa684_xor1;
  wire [0:0] s_wallace_cska32_fa684_or0;
  wire [0:0] s_wallace_cska32_fa685_xor1;
  wire [0:0] s_wallace_cska32_fa685_or0;
  wire [0:0] s_wallace_cska32_fa686_xor1;
  wire [0:0] s_wallace_cska32_fa686_or0;
  wire [0:0] s_wallace_cska32_fa687_xor1;
  wire [0:0] s_wallace_cska32_fa687_or0;
  wire [0:0] s_wallace_cska32_ha16_xor0;
  wire [0:0] s_wallace_cska32_ha16_and0;
  wire [0:0] s_wallace_cska32_fa688_xor1;
  wire [0:0] s_wallace_cska32_fa688_or0;
  wire [0:0] s_wallace_cska32_fa689_xor1;
  wire [0:0] s_wallace_cska32_fa689_or0;
  wire [0:0] s_wallace_cska32_fa690_xor1;
  wire [0:0] s_wallace_cska32_fa690_or0;
  wire [0:0] s_wallace_cska32_fa691_xor1;
  wire [0:0] s_wallace_cska32_fa691_or0;
  wire [0:0] s_wallace_cska32_fa692_xor1;
  wire [0:0] s_wallace_cska32_fa692_or0;
  wire [0:0] s_wallace_cska32_fa693_xor1;
  wire [0:0] s_wallace_cska32_fa693_or0;
  wire [0:0] s_wallace_cska32_fa694_xor1;
  wire [0:0] s_wallace_cska32_fa694_or0;
  wire [0:0] s_wallace_cska32_fa695_xor1;
  wire [0:0] s_wallace_cska32_fa695_or0;
  wire [0:0] s_wallace_cska32_fa696_xor1;
  wire [0:0] s_wallace_cska32_fa696_or0;
  wire [0:0] s_wallace_cska32_fa697_xor1;
  wire [0:0] s_wallace_cska32_fa697_or0;
  wire [0:0] s_wallace_cska32_fa698_xor1;
  wire [0:0] s_wallace_cska32_fa698_or0;
  wire [0:0] s_wallace_cska32_fa699_xor1;
  wire [0:0] s_wallace_cska32_fa699_or0;
  wire [0:0] s_wallace_cska32_fa700_xor1;
  wire [0:0] s_wallace_cska32_fa700_or0;
  wire [0:0] s_wallace_cska32_fa701_xor1;
  wire [0:0] s_wallace_cska32_fa701_or0;
  wire [0:0] s_wallace_cska32_fa702_xor1;
  wire [0:0] s_wallace_cska32_fa702_or0;
  wire [0:0] s_wallace_cska32_fa703_xor1;
  wire [0:0] s_wallace_cska32_fa703_or0;
  wire [0:0] s_wallace_cska32_fa704_xor1;
  wire [0:0] s_wallace_cska32_fa704_or0;
  wire [0:0] s_wallace_cska32_fa705_xor1;
  wire [0:0] s_wallace_cska32_fa705_or0;
  wire [0:0] s_wallace_cska32_fa706_xor1;
  wire [0:0] s_wallace_cska32_fa706_or0;
  wire [0:0] s_wallace_cska32_fa707_xor1;
  wire [0:0] s_wallace_cska32_fa707_or0;
  wire [0:0] s_wallace_cska32_fa708_xor1;
  wire [0:0] s_wallace_cska32_fa708_or0;
  wire [0:0] s_wallace_cska32_fa709_xor1;
  wire [0:0] s_wallace_cska32_fa709_or0;
  wire [0:0] s_wallace_cska32_fa710_xor1;
  wire [0:0] s_wallace_cska32_fa710_or0;
  wire [0:0] s_wallace_cska32_fa711_xor1;
  wire [0:0] s_wallace_cska32_fa711_or0;
  wire [0:0] s_wallace_cska32_fa712_xor1;
  wire [0:0] s_wallace_cska32_fa712_or0;
  wire [0:0] s_wallace_cska32_fa713_xor1;
  wire [0:0] s_wallace_cska32_fa713_or0;
  wire [0:0] s_wallace_cska32_ha17_xor0;
  wire [0:0] s_wallace_cska32_ha17_and0;
  wire [0:0] s_wallace_cska32_fa714_xor1;
  wire [0:0] s_wallace_cska32_fa714_or0;
  wire [0:0] s_wallace_cska32_fa715_xor1;
  wire [0:0] s_wallace_cska32_fa715_or0;
  wire [0:0] s_wallace_cska32_fa716_xor1;
  wire [0:0] s_wallace_cska32_fa716_or0;
  wire [0:0] s_wallace_cska32_fa717_xor1;
  wire [0:0] s_wallace_cska32_fa717_or0;
  wire [0:0] s_wallace_cska32_fa718_xor1;
  wire [0:0] s_wallace_cska32_fa718_or0;
  wire [0:0] s_wallace_cska32_fa719_xor1;
  wire [0:0] s_wallace_cska32_fa719_or0;
  wire [0:0] s_wallace_cska32_fa720_xor1;
  wire [0:0] s_wallace_cska32_fa720_or0;
  wire [0:0] s_wallace_cska32_fa721_xor1;
  wire [0:0] s_wallace_cska32_fa721_or0;
  wire [0:0] s_wallace_cska32_fa722_xor1;
  wire [0:0] s_wallace_cska32_fa722_or0;
  wire [0:0] s_wallace_cska32_fa723_xor1;
  wire [0:0] s_wallace_cska32_fa723_or0;
  wire [0:0] s_wallace_cska32_fa724_xor1;
  wire [0:0] s_wallace_cska32_fa724_or0;
  wire [0:0] s_wallace_cska32_fa725_xor1;
  wire [0:0] s_wallace_cska32_fa725_or0;
  wire [0:0] s_wallace_cska32_fa726_xor1;
  wire [0:0] s_wallace_cska32_fa726_or0;
  wire [0:0] s_wallace_cska32_fa727_xor1;
  wire [0:0] s_wallace_cska32_fa727_or0;
  wire [0:0] s_wallace_cska32_fa728_xor1;
  wire [0:0] s_wallace_cska32_fa728_or0;
  wire [0:0] s_wallace_cska32_fa729_xor1;
  wire [0:0] s_wallace_cska32_fa729_or0;
  wire [0:0] s_wallace_cska32_fa730_xor1;
  wire [0:0] s_wallace_cska32_fa730_or0;
  wire [0:0] s_wallace_cska32_fa731_xor1;
  wire [0:0] s_wallace_cska32_fa731_or0;
  wire [0:0] s_wallace_cska32_fa732_xor1;
  wire [0:0] s_wallace_cska32_fa732_or0;
  wire [0:0] s_wallace_cska32_fa733_xor1;
  wire [0:0] s_wallace_cska32_fa733_or0;
  wire [0:0] s_wallace_cska32_fa734_xor1;
  wire [0:0] s_wallace_cska32_fa734_or0;
  wire [0:0] s_wallace_cska32_fa735_xor1;
  wire [0:0] s_wallace_cska32_fa735_or0;
  wire [0:0] s_wallace_cska32_fa736_xor1;
  wire [0:0] s_wallace_cska32_fa736_or0;
  wire [0:0] s_wallace_cska32_fa737_xor1;
  wire [0:0] s_wallace_cska32_fa737_or0;
  wire [0:0] s_wallace_cska32_ha18_xor0;
  wire [0:0] s_wallace_cska32_ha18_and0;
  wire [0:0] s_wallace_cska32_fa738_xor1;
  wire [0:0] s_wallace_cska32_fa738_or0;
  wire [0:0] s_wallace_cska32_fa739_xor1;
  wire [0:0] s_wallace_cska32_fa739_or0;
  wire [0:0] s_wallace_cska32_fa740_xor1;
  wire [0:0] s_wallace_cska32_fa740_or0;
  wire [0:0] s_wallace_cska32_fa741_xor1;
  wire [0:0] s_wallace_cska32_fa741_or0;
  wire [0:0] s_wallace_cska32_fa742_xor1;
  wire [0:0] s_wallace_cska32_fa742_or0;
  wire [0:0] s_wallace_cska32_fa743_xor1;
  wire [0:0] s_wallace_cska32_fa743_or0;
  wire [0:0] s_wallace_cska32_fa744_xor1;
  wire [0:0] s_wallace_cska32_fa744_or0;
  wire [0:0] s_wallace_cska32_fa745_xor1;
  wire [0:0] s_wallace_cska32_fa745_or0;
  wire [0:0] s_wallace_cska32_fa746_xor1;
  wire [0:0] s_wallace_cska32_fa746_or0;
  wire [0:0] s_wallace_cska32_fa747_xor1;
  wire [0:0] s_wallace_cska32_fa747_or0;
  wire [0:0] s_wallace_cska32_fa748_xor1;
  wire [0:0] s_wallace_cska32_fa748_or0;
  wire [0:0] s_wallace_cska32_fa749_xor1;
  wire [0:0] s_wallace_cska32_fa749_or0;
  wire [0:0] s_wallace_cska32_fa750_xor1;
  wire [0:0] s_wallace_cska32_fa750_or0;
  wire [0:0] s_wallace_cska32_fa751_xor1;
  wire [0:0] s_wallace_cska32_fa751_or0;
  wire [0:0] s_wallace_cska32_fa752_xor1;
  wire [0:0] s_wallace_cska32_fa752_or0;
  wire [0:0] s_wallace_cska32_fa753_xor1;
  wire [0:0] s_wallace_cska32_fa753_or0;
  wire [0:0] s_wallace_cska32_fa754_xor1;
  wire [0:0] s_wallace_cska32_fa754_or0;
  wire [0:0] s_wallace_cska32_fa755_xor1;
  wire [0:0] s_wallace_cska32_fa755_or0;
  wire [0:0] s_wallace_cska32_fa756_xor1;
  wire [0:0] s_wallace_cska32_fa756_or0;
  wire [0:0] s_wallace_cska32_fa757_xor1;
  wire [0:0] s_wallace_cska32_fa757_or0;
  wire [0:0] s_wallace_cska32_fa758_xor1;
  wire [0:0] s_wallace_cska32_fa758_or0;
  wire [0:0] s_wallace_cska32_fa759_xor1;
  wire [0:0] s_wallace_cska32_fa759_or0;
  wire [0:0] s_wallace_cska32_ha19_xor0;
  wire [0:0] s_wallace_cska32_ha19_and0;
  wire [0:0] s_wallace_cska32_fa760_xor1;
  wire [0:0] s_wallace_cska32_fa760_or0;
  wire [0:0] s_wallace_cska32_fa761_xor1;
  wire [0:0] s_wallace_cska32_fa761_or0;
  wire [0:0] s_wallace_cska32_fa762_xor1;
  wire [0:0] s_wallace_cska32_fa762_or0;
  wire [0:0] s_wallace_cska32_fa763_xor1;
  wire [0:0] s_wallace_cska32_fa763_or0;
  wire [0:0] s_wallace_cska32_fa764_xor1;
  wire [0:0] s_wallace_cska32_fa764_or0;
  wire [0:0] s_wallace_cska32_fa765_xor1;
  wire [0:0] s_wallace_cska32_fa765_or0;
  wire [0:0] s_wallace_cska32_fa766_xor1;
  wire [0:0] s_wallace_cska32_fa766_or0;
  wire [0:0] s_wallace_cska32_fa767_xor1;
  wire [0:0] s_wallace_cska32_fa767_or0;
  wire [0:0] s_wallace_cska32_fa768_xor1;
  wire [0:0] s_wallace_cska32_fa768_or0;
  wire [0:0] s_wallace_cska32_fa769_xor1;
  wire [0:0] s_wallace_cska32_fa769_or0;
  wire [0:0] s_wallace_cska32_fa770_xor1;
  wire [0:0] s_wallace_cska32_fa770_or0;
  wire [0:0] s_wallace_cska32_fa771_xor1;
  wire [0:0] s_wallace_cska32_fa771_or0;
  wire [0:0] s_wallace_cska32_fa772_xor1;
  wire [0:0] s_wallace_cska32_fa772_or0;
  wire [0:0] s_wallace_cska32_fa773_xor1;
  wire [0:0] s_wallace_cska32_fa773_or0;
  wire [0:0] s_wallace_cska32_fa774_xor1;
  wire [0:0] s_wallace_cska32_fa774_or0;
  wire [0:0] s_wallace_cska32_fa775_xor1;
  wire [0:0] s_wallace_cska32_fa775_or0;
  wire [0:0] s_wallace_cska32_fa776_xor1;
  wire [0:0] s_wallace_cska32_fa776_or0;
  wire [0:0] s_wallace_cska32_fa777_xor1;
  wire [0:0] s_wallace_cska32_fa777_or0;
  wire [0:0] s_wallace_cska32_fa778_xor1;
  wire [0:0] s_wallace_cska32_fa778_or0;
  wire [0:0] s_wallace_cska32_fa779_xor1;
  wire [0:0] s_wallace_cska32_fa779_or0;
  wire [0:0] s_wallace_cska32_ha20_xor0;
  wire [0:0] s_wallace_cska32_ha20_and0;
  wire [0:0] s_wallace_cska32_fa780_xor1;
  wire [0:0] s_wallace_cska32_fa780_or0;
  wire [0:0] s_wallace_cska32_fa781_xor1;
  wire [0:0] s_wallace_cska32_fa781_or0;
  wire [0:0] s_wallace_cska32_fa782_xor1;
  wire [0:0] s_wallace_cska32_fa782_or0;
  wire [0:0] s_wallace_cska32_fa783_xor1;
  wire [0:0] s_wallace_cska32_fa783_or0;
  wire [0:0] s_wallace_cska32_fa784_xor1;
  wire [0:0] s_wallace_cska32_fa784_or0;
  wire [0:0] s_wallace_cska32_fa785_xor1;
  wire [0:0] s_wallace_cska32_fa785_or0;
  wire [0:0] s_wallace_cska32_fa786_xor1;
  wire [0:0] s_wallace_cska32_fa786_or0;
  wire [0:0] s_wallace_cska32_fa787_xor1;
  wire [0:0] s_wallace_cska32_fa787_or0;
  wire [0:0] s_wallace_cska32_fa788_xor1;
  wire [0:0] s_wallace_cska32_fa788_or0;
  wire [0:0] s_wallace_cska32_fa789_xor1;
  wire [0:0] s_wallace_cska32_fa789_or0;
  wire [0:0] s_wallace_cska32_fa790_xor1;
  wire [0:0] s_wallace_cska32_fa790_or0;
  wire [0:0] s_wallace_cska32_fa791_xor1;
  wire [0:0] s_wallace_cska32_fa791_or0;
  wire [0:0] s_wallace_cska32_fa792_xor1;
  wire [0:0] s_wallace_cska32_fa792_or0;
  wire [0:0] s_wallace_cska32_fa793_xor1;
  wire [0:0] s_wallace_cska32_fa793_or0;
  wire [0:0] s_wallace_cska32_fa794_xor1;
  wire [0:0] s_wallace_cska32_fa794_or0;
  wire [0:0] s_wallace_cska32_fa795_xor1;
  wire [0:0] s_wallace_cska32_fa795_or0;
  wire [0:0] s_wallace_cska32_fa796_xor1;
  wire [0:0] s_wallace_cska32_fa796_or0;
  wire [0:0] s_wallace_cska32_fa797_xor1;
  wire [0:0] s_wallace_cska32_fa797_or0;
  wire [0:0] s_wallace_cska32_ha21_xor0;
  wire [0:0] s_wallace_cska32_ha21_and0;
  wire [0:0] s_wallace_cska32_fa798_xor1;
  wire [0:0] s_wallace_cska32_fa798_or0;
  wire [0:0] s_wallace_cska32_fa799_xor1;
  wire [0:0] s_wallace_cska32_fa799_or0;
  wire [0:0] s_wallace_cska32_fa800_xor1;
  wire [0:0] s_wallace_cska32_fa800_or0;
  wire [0:0] s_wallace_cska32_fa801_xor1;
  wire [0:0] s_wallace_cska32_fa801_or0;
  wire [0:0] s_wallace_cska32_fa802_xor1;
  wire [0:0] s_wallace_cska32_fa802_or0;
  wire [0:0] s_wallace_cska32_fa803_xor1;
  wire [0:0] s_wallace_cska32_fa803_or0;
  wire [0:0] s_wallace_cska32_fa804_xor1;
  wire [0:0] s_wallace_cska32_fa804_or0;
  wire [0:0] s_wallace_cska32_fa805_xor1;
  wire [0:0] s_wallace_cska32_fa805_or0;
  wire [0:0] s_wallace_cska32_fa806_xor1;
  wire [0:0] s_wallace_cska32_fa806_or0;
  wire [0:0] s_wallace_cska32_fa807_xor1;
  wire [0:0] s_wallace_cska32_fa807_or0;
  wire [0:0] s_wallace_cska32_fa808_xor1;
  wire [0:0] s_wallace_cska32_fa808_or0;
  wire [0:0] s_wallace_cska32_fa809_xor1;
  wire [0:0] s_wallace_cska32_fa809_or0;
  wire [0:0] s_wallace_cska32_fa810_xor1;
  wire [0:0] s_wallace_cska32_fa810_or0;
  wire [0:0] s_wallace_cska32_fa811_xor1;
  wire [0:0] s_wallace_cska32_fa811_or0;
  wire [0:0] s_wallace_cska32_fa812_xor1;
  wire [0:0] s_wallace_cska32_fa812_or0;
  wire [0:0] s_wallace_cska32_fa813_xor1;
  wire [0:0] s_wallace_cska32_fa813_or0;
  wire [0:0] s_wallace_cska32_ha22_xor0;
  wire [0:0] s_wallace_cska32_ha22_and0;
  wire [0:0] s_wallace_cska32_fa814_xor1;
  wire [0:0] s_wallace_cska32_fa814_or0;
  wire [0:0] s_wallace_cska32_fa815_xor1;
  wire [0:0] s_wallace_cska32_fa815_or0;
  wire [0:0] s_wallace_cska32_fa816_xor1;
  wire [0:0] s_wallace_cska32_fa816_or0;
  wire [0:0] s_wallace_cska32_fa817_xor1;
  wire [0:0] s_wallace_cska32_fa817_or0;
  wire [0:0] s_wallace_cska32_fa818_xor1;
  wire [0:0] s_wallace_cska32_fa818_or0;
  wire [0:0] s_wallace_cska32_fa819_xor1;
  wire [0:0] s_wallace_cska32_fa819_or0;
  wire [0:0] s_wallace_cska32_fa820_xor1;
  wire [0:0] s_wallace_cska32_fa820_or0;
  wire [0:0] s_wallace_cska32_fa821_xor1;
  wire [0:0] s_wallace_cska32_fa821_or0;
  wire [0:0] s_wallace_cska32_fa822_xor1;
  wire [0:0] s_wallace_cska32_fa822_or0;
  wire [0:0] s_wallace_cska32_fa823_xor1;
  wire [0:0] s_wallace_cska32_fa823_or0;
  wire [0:0] s_wallace_cska32_fa824_xor1;
  wire [0:0] s_wallace_cska32_fa824_or0;
  wire [0:0] s_wallace_cska32_fa825_xor1;
  wire [0:0] s_wallace_cska32_fa825_or0;
  wire [0:0] s_wallace_cska32_fa826_xor1;
  wire [0:0] s_wallace_cska32_fa826_or0;
  wire [0:0] s_wallace_cska32_fa827_xor1;
  wire [0:0] s_wallace_cska32_fa827_or0;
  wire [0:0] s_wallace_cska32_ha23_xor0;
  wire [0:0] s_wallace_cska32_ha23_and0;
  wire [0:0] s_wallace_cska32_fa828_xor1;
  wire [0:0] s_wallace_cska32_fa828_or0;
  wire [0:0] s_wallace_cska32_fa829_xor1;
  wire [0:0] s_wallace_cska32_fa829_or0;
  wire [0:0] s_wallace_cska32_fa830_xor1;
  wire [0:0] s_wallace_cska32_fa830_or0;
  wire [0:0] s_wallace_cska32_fa831_xor1;
  wire [0:0] s_wallace_cska32_fa831_or0;
  wire [0:0] s_wallace_cska32_fa832_xor1;
  wire [0:0] s_wallace_cska32_fa832_or0;
  wire [0:0] s_wallace_cska32_fa833_xor1;
  wire [0:0] s_wallace_cska32_fa833_or0;
  wire [0:0] s_wallace_cska32_fa834_xor1;
  wire [0:0] s_wallace_cska32_fa834_or0;
  wire [0:0] s_wallace_cska32_fa835_xor1;
  wire [0:0] s_wallace_cska32_fa835_or0;
  wire [0:0] s_wallace_cska32_fa836_xor1;
  wire [0:0] s_wallace_cska32_fa836_or0;
  wire [0:0] s_wallace_cska32_fa837_xor1;
  wire [0:0] s_wallace_cska32_fa837_or0;
  wire [0:0] s_wallace_cska32_fa838_xor1;
  wire [0:0] s_wallace_cska32_fa838_or0;
  wire [0:0] s_wallace_cska32_fa839_xor1;
  wire [0:0] s_wallace_cska32_fa839_or0;
  wire [0:0] s_wallace_cska32_ha24_xor0;
  wire [0:0] s_wallace_cska32_ha24_and0;
  wire [0:0] s_wallace_cska32_fa840_xor1;
  wire [0:0] s_wallace_cska32_fa840_or0;
  wire [0:0] s_wallace_cska32_fa841_xor1;
  wire [0:0] s_wallace_cska32_fa841_or0;
  wire [0:0] s_wallace_cska32_fa842_xor1;
  wire [0:0] s_wallace_cska32_fa842_or0;
  wire [0:0] s_wallace_cska32_fa843_xor1;
  wire [0:0] s_wallace_cska32_fa843_or0;
  wire [0:0] s_wallace_cska32_fa844_xor1;
  wire [0:0] s_wallace_cska32_fa844_or0;
  wire [0:0] s_wallace_cska32_fa845_xor1;
  wire [0:0] s_wallace_cska32_fa845_or0;
  wire [0:0] s_wallace_cska32_fa846_xor1;
  wire [0:0] s_wallace_cska32_fa846_or0;
  wire [0:0] s_wallace_cska32_fa847_xor1;
  wire [0:0] s_wallace_cska32_fa847_or0;
  wire [0:0] s_wallace_cska32_fa848_xor1;
  wire [0:0] s_wallace_cska32_fa848_or0;
  wire [0:0] s_wallace_cska32_fa849_xor1;
  wire [0:0] s_wallace_cska32_fa849_or0;
  wire [0:0] s_wallace_cska32_ha25_xor0;
  wire [0:0] s_wallace_cska32_ha25_and0;
  wire [0:0] s_wallace_cska32_fa850_xor1;
  wire [0:0] s_wallace_cska32_fa850_or0;
  wire [0:0] s_wallace_cska32_fa851_xor1;
  wire [0:0] s_wallace_cska32_fa851_or0;
  wire [0:0] s_wallace_cska32_fa852_xor1;
  wire [0:0] s_wallace_cska32_fa852_or0;
  wire [0:0] s_wallace_cska32_fa853_xor1;
  wire [0:0] s_wallace_cska32_fa853_or0;
  wire [0:0] s_wallace_cska32_fa854_xor1;
  wire [0:0] s_wallace_cska32_fa854_or0;
  wire [0:0] s_wallace_cska32_fa855_xor1;
  wire [0:0] s_wallace_cska32_fa855_or0;
  wire [0:0] s_wallace_cska32_fa856_xor1;
  wire [0:0] s_wallace_cska32_fa856_or0;
  wire [0:0] s_wallace_cska32_fa857_xor1;
  wire [0:0] s_wallace_cska32_fa857_or0;
  wire [0:0] s_wallace_cska32_ha26_xor0;
  wire [0:0] s_wallace_cska32_ha26_and0;
  wire [0:0] s_wallace_cska32_fa858_xor1;
  wire [0:0] s_wallace_cska32_fa858_or0;
  wire [0:0] s_wallace_cska32_fa859_xor1;
  wire [0:0] s_wallace_cska32_fa859_or0;
  wire [0:0] s_wallace_cska32_fa860_xor1;
  wire [0:0] s_wallace_cska32_fa860_or0;
  wire [0:0] s_wallace_cska32_fa861_xor1;
  wire [0:0] s_wallace_cska32_fa861_or0;
  wire [0:0] s_wallace_cska32_fa862_xor1;
  wire [0:0] s_wallace_cska32_fa862_or0;
  wire [0:0] s_wallace_cska32_fa863_xor1;
  wire [0:0] s_wallace_cska32_fa863_or0;
  wire [0:0] s_wallace_cska32_ha27_xor0;
  wire [0:0] s_wallace_cska32_ha27_and0;
  wire [0:0] s_wallace_cska32_fa864_xor1;
  wire [0:0] s_wallace_cska32_fa864_or0;
  wire [0:0] s_wallace_cska32_fa865_xor1;
  wire [0:0] s_wallace_cska32_fa865_or0;
  wire [0:0] s_wallace_cska32_fa866_xor1;
  wire [0:0] s_wallace_cska32_fa866_or0;
  wire [0:0] s_wallace_cska32_fa867_xor1;
  wire [0:0] s_wallace_cska32_fa867_or0;
  wire [0:0] s_wallace_cska32_ha28_xor0;
  wire [0:0] s_wallace_cska32_ha28_and0;
  wire [0:0] s_wallace_cska32_fa868_xor1;
  wire [0:0] s_wallace_cska32_fa868_or0;
  wire [0:0] s_wallace_cska32_fa869_xor1;
  wire [0:0] s_wallace_cska32_fa869_or0;
  wire [0:0] s_wallace_cska32_ha29_xor0;
  wire [0:0] s_wallace_cska32_ha29_and0;
  wire [0:0] s_wallace_cska32_fa870_xor1;
  wire [0:0] s_wallace_cska32_fa870_or0;
  wire [0:0] s_wallace_cska32_fa871_xor1;
  wire [0:0] s_wallace_cska32_fa871_or0;
  wire [0:0] s_wallace_cska32_fa872_xor1;
  wire [0:0] s_wallace_cska32_fa872_or0;
  wire [0:0] s_wallace_cska32_fa873_xor1;
  wire [0:0] s_wallace_cska32_fa873_or0;
  wire [0:0] s_wallace_cska32_fa874_xor1;
  wire [0:0] s_wallace_cska32_fa874_or0;
  wire [0:0] s_wallace_cska32_fa875_xor1;
  wire [0:0] s_wallace_cska32_fa875_or0;
  wire [0:0] s_wallace_cska32_fa876_xor1;
  wire [0:0] s_wallace_cska32_fa876_or0;
  wire [0:0] s_wallace_cska32_fa877_xor1;
  wire [0:0] s_wallace_cska32_fa877_or0;
  wire [0:0] s_wallace_cska32_fa878_xor1;
  wire [0:0] s_wallace_cska32_fa878_or0;
  wire [0:0] s_wallace_cska32_fa879_xor1;
  wire [0:0] s_wallace_cska32_fa879_or0;
  wire [0:0] s_wallace_cska32_fa880_xor1;
  wire [0:0] s_wallace_cska32_fa880_or0;
  wire [0:0] s_wallace_cska32_fa881_xor1;
  wire [0:0] s_wallace_cska32_fa881_or0;
  wire [0:0] s_wallace_cska32_fa882_xor1;
  wire [0:0] s_wallace_cska32_fa882_or0;
  wire [0:0] s_wallace_cska32_fa883_xor1;
  wire [0:0] s_wallace_cska32_fa883_or0;
  wire [0:0] s_wallace_cska32_fa884_xor1;
  wire [0:0] s_wallace_cska32_fa884_or0;
  wire [0:0] s_wallace_cska32_fa885_xor1;
  wire [0:0] s_wallace_cska32_fa885_or0;
  wire [0:0] s_wallace_cska32_fa886_xor1;
  wire [0:0] s_wallace_cska32_fa886_or0;
  wire [0:0] s_wallace_cska32_fa887_xor1;
  wire [0:0] s_wallace_cska32_fa887_or0;
  wire [0:0] s_wallace_cska32_fa888_xor1;
  wire [0:0] s_wallace_cska32_fa888_or0;
  wire [0:0] s_wallace_cska32_fa889_xor1;
  wire [0:0] s_wallace_cska32_fa889_or0;
  wire [0:0] s_wallace_cska32_fa890_xor1;
  wire [0:0] s_wallace_cska32_fa890_or0;
  wire [0:0] s_wallace_cska32_fa891_xor1;
  wire [0:0] s_wallace_cska32_fa891_or0;
  wire [0:0] s_wallace_cska32_fa892_xor1;
  wire [0:0] s_wallace_cska32_fa892_or0;
  wire [0:0] s_wallace_cska32_fa893_xor1;
  wire [0:0] s_wallace_cska32_fa893_or0;
  wire [0:0] s_wallace_cska32_fa894_xor1;
  wire [0:0] s_wallace_cska32_fa894_or0;
  wire [0:0] s_wallace_cska32_fa895_xor1;
  wire [0:0] s_wallace_cska32_fa895_or0;
  wire [0:0] s_wallace_cska32_fa896_xor1;
  wire [0:0] s_wallace_cska32_fa896_or0;
  wire [0:0] s_wallace_cska32_fa897_xor1;
  wire [0:0] s_wallace_cska32_fa897_or0;
  wire [0:0] s_wallace_cska32_nand_29_31;
  wire [0:0] s_wallace_cska32_fa898_xor1;
  wire [0:0] s_wallace_cska32_fa898_or0;
  wire [0:0] s_wallace_cska32_nand_31_30;
  wire [0:0] s_wallace_cska32_fa899_xor1;
  wire [0:0] s_wallace_cska32_fa899_or0;
  wire [0:0] s_wallace_cska32_and_0_0;
  wire [0:0] s_wallace_cska32_and_1_0;
  wire [0:0] s_wallace_cska32_and_0_2;
  wire [0:0] s_wallace_cska32_nand_30_31;
  wire [0:0] s_wallace_cska32_and_0_1;
  wire [0:0] s_wallace_cska32_and_31_31;
  wire [61:0] s_wallace_cska32_u_cska62_a;
  wire [61:0] s_wallace_cska32_u_cska62_b;
  wire [62:0] s_wallace_cska32_u_cska62_out;
  wire [0:0] s_wallace_cska32_xor0;

  and_gate and_gate_s_wallace_cska32_and_2_0(.a(a[2]), .b(b[0]), .out(s_wallace_cska32_and_2_0));
  and_gate and_gate_s_wallace_cska32_and_1_1(.a(a[1]), .b(b[1]), .out(s_wallace_cska32_and_1_1));
  ha ha_s_wallace_cska32_ha0_out(.a(s_wallace_cska32_and_2_0[0]), .b(s_wallace_cska32_and_1_1[0]), .ha_xor0(s_wallace_cska32_ha0_xor0), .ha_and0(s_wallace_cska32_ha0_and0));
  and_gate and_gate_s_wallace_cska32_and_3_0(.a(a[3]), .b(b[0]), .out(s_wallace_cska32_and_3_0));
  and_gate and_gate_s_wallace_cska32_and_2_1(.a(a[2]), .b(b[1]), .out(s_wallace_cska32_and_2_1));
  fa fa_s_wallace_cska32_fa0_out(.a(s_wallace_cska32_ha0_and0[0]), .b(s_wallace_cska32_and_3_0[0]), .cin(s_wallace_cska32_and_2_1[0]), .fa_xor1(s_wallace_cska32_fa0_xor1), .fa_or0(s_wallace_cska32_fa0_or0));
  and_gate and_gate_s_wallace_cska32_and_4_0(.a(a[4]), .b(b[0]), .out(s_wallace_cska32_and_4_0));
  and_gate and_gate_s_wallace_cska32_and_3_1(.a(a[3]), .b(b[1]), .out(s_wallace_cska32_and_3_1));
  fa fa_s_wallace_cska32_fa1_out(.a(s_wallace_cska32_fa0_or0[0]), .b(s_wallace_cska32_and_4_0[0]), .cin(s_wallace_cska32_and_3_1[0]), .fa_xor1(s_wallace_cska32_fa1_xor1), .fa_or0(s_wallace_cska32_fa1_or0));
  and_gate and_gate_s_wallace_cska32_and_5_0(.a(a[5]), .b(b[0]), .out(s_wallace_cska32_and_5_0));
  and_gate and_gate_s_wallace_cska32_and_4_1(.a(a[4]), .b(b[1]), .out(s_wallace_cska32_and_4_1));
  fa fa_s_wallace_cska32_fa2_out(.a(s_wallace_cska32_fa1_or0[0]), .b(s_wallace_cska32_and_5_0[0]), .cin(s_wallace_cska32_and_4_1[0]), .fa_xor1(s_wallace_cska32_fa2_xor1), .fa_or0(s_wallace_cska32_fa2_or0));
  and_gate and_gate_s_wallace_cska32_and_6_0(.a(a[6]), .b(b[0]), .out(s_wallace_cska32_and_6_0));
  and_gate and_gate_s_wallace_cska32_and_5_1(.a(a[5]), .b(b[1]), .out(s_wallace_cska32_and_5_1));
  fa fa_s_wallace_cska32_fa3_out(.a(s_wallace_cska32_fa2_or0[0]), .b(s_wallace_cska32_and_6_0[0]), .cin(s_wallace_cska32_and_5_1[0]), .fa_xor1(s_wallace_cska32_fa3_xor1), .fa_or0(s_wallace_cska32_fa3_or0));
  and_gate and_gate_s_wallace_cska32_and_7_0(.a(a[7]), .b(b[0]), .out(s_wallace_cska32_and_7_0));
  and_gate and_gate_s_wallace_cska32_and_6_1(.a(a[6]), .b(b[1]), .out(s_wallace_cska32_and_6_1));
  fa fa_s_wallace_cska32_fa4_out(.a(s_wallace_cska32_fa3_or0[0]), .b(s_wallace_cska32_and_7_0[0]), .cin(s_wallace_cska32_and_6_1[0]), .fa_xor1(s_wallace_cska32_fa4_xor1), .fa_or0(s_wallace_cska32_fa4_or0));
  and_gate and_gate_s_wallace_cska32_and_8_0(.a(a[8]), .b(b[0]), .out(s_wallace_cska32_and_8_0));
  and_gate and_gate_s_wallace_cska32_and_7_1(.a(a[7]), .b(b[1]), .out(s_wallace_cska32_and_7_1));
  fa fa_s_wallace_cska32_fa5_out(.a(s_wallace_cska32_fa4_or0[0]), .b(s_wallace_cska32_and_8_0[0]), .cin(s_wallace_cska32_and_7_1[0]), .fa_xor1(s_wallace_cska32_fa5_xor1), .fa_or0(s_wallace_cska32_fa5_or0));
  and_gate and_gate_s_wallace_cska32_and_9_0(.a(a[9]), .b(b[0]), .out(s_wallace_cska32_and_9_0));
  and_gate and_gate_s_wallace_cska32_and_8_1(.a(a[8]), .b(b[1]), .out(s_wallace_cska32_and_8_1));
  fa fa_s_wallace_cska32_fa6_out(.a(s_wallace_cska32_fa5_or0[0]), .b(s_wallace_cska32_and_9_0[0]), .cin(s_wallace_cska32_and_8_1[0]), .fa_xor1(s_wallace_cska32_fa6_xor1), .fa_or0(s_wallace_cska32_fa6_or0));
  and_gate and_gate_s_wallace_cska32_and_10_0(.a(a[10]), .b(b[0]), .out(s_wallace_cska32_and_10_0));
  and_gate and_gate_s_wallace_cska32_and_9_1(.a(a[9]), .b(b[1]), .out(s_wallace_cska32_and_9_1));
  fa fa_s_wallace_cska32_fa7_out(.a(s_wallace_cska32_fa6_or0[0]), .b(s_wallace_cska32_and_10_0[0]), .cin(s_wallace_cska32_and_9_1[0]), .fa_xor1(s_wallace_cska32_fa7_xor1), .fa_or0(s_wallace_cska32_fa7_or0));
  and_gate and_gate_s_wallace_cska32_and_11_0(.a(a[11]), .b(b[0]), .out(s_wallace_cska32_and_11_0));
  and_gate and_gate_s_wallace_cska32_and_10_1(.a(a[10]), .b(b[1]), .out(s_wallace_cska32_and_10_1));
  fa fa_s_wallace_cska32_fa8_out(.a(s_wallace_cska32_fa7_or0[0]), .b(s_wallace_cska32_and_11_0[0]), .cin(s_wallace_cska32_and_10_1[0]), .fa_xor1(s_wallace_cska32_fa8_xor1), .fa_or0(s_wallace_cska32_fa8_or0));
  and_gate and_gate_s_wallace_cska32_and_12_0(.a(a[12]), .b(b[0]), .out(s_wallace_cska32_and_12_0));
  and_gate and_gate_s_wallace_cska32_and_11_1(.a(a[11]), .b(b[1]), .out(s_wallace_cska32_and_11_1));
  fa fa_s_wallace_cska32_fa9_out(.a(s_wallace_cska32_fa8_or0[0]), .b(s_wallace_cska32_and_12_0[0]), .cin(s_wallace_cska32_and_11_1[0]), .fa_xor1(s_wallace_cska32_fa9_xor1), .fa_or0(s_wallace_cska32_fa9_or0));
  and_gate and_gate_s_wallace_cska32_and_13_0(.a(a[13]), .b(b[0]), .out(s_wallace_cska32_and_13_0));
  and_gate and_gate_s_wallace_cska32_and_12_1(.a(a[12]), .b(b[1]), .out(s_wallace_cska32_and_12_1));
  fa fa_s_wallace_cska32_fa10_out(.a(s_wallace_cska32_fa9_or0[0]), .b(s_wallace_cska32_and_13_0[0]), .cin(s_wallace_cska32_and_12_1[0]), .fa_xor1(s_wallace_cska32_fa10_xor1), .fa_or0(s_wallace_cska32_fa10_or0));
  and_gate and_gate_s_wallace_cska32_and_14_0(.a(a[14]), .b(b[0]), .out(s_wallace_cska32_and_14_0));
  and_gate and_gate_s_wallace_cska32_and_13_1(.a(a[13]), .b(b[1]), .out(s_wallace_cska32_and_13_1));
  fa fa_s_wallace_cska32_fa11_out(.a(s_wallace_cska32_fa10_or0[0]), .b(s_wallace_cska32_and_14_0[0]), .cin(s_wallace_cska32_and_13_1[0]), .fa_xor1(s_wallace_cska32_fa11_xor1), .fa_or0(s_wallace_cska32_fa11_or0));
  and_gate and_gate_s_wallace_cska32_and_15_0(.a(a[15]), .b(b[0]), .out(s_wallace_cska32_and_15_0));
  and_gate and_gate_s_wallace_cska32_and_14_1(.a(a[14]), .b(b[1]), .out(s_wallace_cska32_and_14_1));
  fa fa_s_wallace_cska32_fa12_out(.a(s_wallace_cska32_fa11_or0[0]), .b(s_wallace_cska32_and_15_0[0]), .cin(s_wallace_cska32_and_14_1[0]), .fa_xor1(s_wallace_cska32_fa12_xor1), .fa_or0(s_wallace_cska32_fa12_or0));
  and_gate and_gate_s_wallace_cska32_and_16_0(.a(a[16]), .b(b[0]), .out(s_wallace_cska32_and_16_0));
  and_gate and_gate_s_wallace_cska32_and_15_1(.a(a[15]), .b(b[1]), .out(s_wallace_cska32_and_15_1));
  fa fa_s_wallace_cska32_fa13_out(.a(s_wallace_cska32_fa12_or0[0]), .b(s_wallace_cska32_and_16_0[0]), .cin(s_wallace_cska32_and_15_1[0]), .fa_xor1(s_wallace_cska32_fa13_xor1), .fa_or0(s_wallace_cska32_fa13_or0));
  and_gate and_gate_s_wallace_cska32_and_17_0(.a(a[17]), .b(b[0]), .out(s_wallace_cska32_and_17_0));
  and_gate and_gate_s_wallace_cska32_and_16_1(.a(a[16]), .b(b[1]), .out(s_wallace_cska32_and_16_1));
  fa fa_s_wallace_cska32_fa14_out(.a(s_wallace_cska32_fa13_or0[0]), .b(s_wallace_cska32_and_17_0[0]), .cin(s_wallace_cska32_and_16_1[0]), .fa_xor1(s_wallace_cska32_fa14_xor1), .fa_or0(s_wallace_cska32_fa14_or0));
  and_gate and_gate_s_wallace_cska32_and_18_0(.a(a[18]), .b(b[0]), .out(s_wallace_cska32_and_18_0));
  and_gate and_gate_s_wallace_cska32_and_17_1(.a(a[17]), .b(b[1]), .out(s_wallace_cska32_and_17_1));
  fa fa_s_wallace_cska32_fa15_out(.a(s_wallace_cska32_fa14_or0[0]), .b(s_wallace_cska32_and_18_0[0]), .cin(s_wallace_cska32_and_17_1[0]), .fa_xor1(s_wallace_cska32_fa15_xor1), .fa_or0(s_wallace_cska32_fa15_or0));
  and_gate and_gate_s_wallace_cska32_and_19_0(.a(a[19]), .b(b[0]), .out(s_wallace_cska32_and_19_0));
  and_gate and_gate_s_wallace_cska32_and_18_1(.a(a[18]), .b(b[1]), .out(s_wallace_cska32_and_18_1));
  fa fa_s_wallace_cska32_fa16_out(.a(s_wallace_cska32_fa15_or0[0]), .b(s_wallace_cska32_and_19_0[0]), .cin(s_wallace_cska32_and_18_1[0]), .fa_xor1(s_wallace_cska32_fa16_xor1), .fa_or0(s_wallace_cska32_fa16_or0));
  and_gate and_gate_s_wallace_cska32_and_20_0(.a(a[20]), .b(b[0]), .out(s_wallace_cska32_and_20_0));
  and_gate and_gate_s_wallace_cska32_and_19_1(.a(a[19]), .b(b[1]), .out(s_wallace_cska32_and_19_1));
  fa fa_s_wallace_cska32_fa17_out(.a(s_wallace_cska32_fa16_or0[0]), .b(s_wallace_cska32_and_20_0[0]), .cin(s_wallace_cska32_and_19_1[0]), .fa_xor1(s_wallace_cska32_fa17_xor1), .fa_or0(s_wallace_cska32_fa17_or0));
  and_gate and_gate_s_wallace_cska32_and_21_0(.a(a[21]), .b(b[0]), .out(s_wallace_cska32_and_21_0));
  and_gate and_gate_s_wallace_cska32_and_20_1(.a(a[20]), .b(b[1]), .out(s_wallace_cska32_and_20_1));
  fa fa_s_wallace_cska32_fa18_out(.a(s_wallace_cska32_fa17_or0[0]), .b(s_wallace_cska32_and_21_0[0]), .cin(s_wallace_cska32_and_20_1[0]), .fa_xor1(s_wallace_cska32_fa18_xor1), .fa_or0(s_wallace_cska32_fa18_or0));
  and_gate and_gate_s_wallace_cska32_and_22_0(.a(a[22]), .b(b[0]), .out(s_wallace_cska32_and_22_0));
  and_gate and_gate_s_wallace_cska32_and_21_1(.a(a[21]), .b(b[1]), .out(s_wallace_cska32_and_21_1));
  fa fa_s_wallace_cska32_fa19_out(.a(s_wallace_cska32_fa18_or0[0]), .b(s_wallace_cska32_and_22_0[0]), .cin(s_wallace_cska32_and_21_1[0]), .fa_xor1(s_wallace_cska32_fa19_xor1), .fa_or0(s_wallace_cska32_fa19_or0));
  and_gate and_gate_s_wallace_cska32_and_23_0(.a(a[23]), .b(b[0]), .out(s_wallace_cska32_and_23_0));
  and_gate and_gate_s_wallace_cska32_and_22_1(.a(a[22]), .b(b[1]), .out(s_wallace_cska32_and_22_1));
  fa fa_s_wallace_cska32_fa20_out(.a(s_wallace_cska32_fa19_or0[0]), .b(s_wallace_cska32_and_23_0[0]), .cin(s_wallace_cska32_and_22_1[0]), .fa_xor1(s_wallace_cska32_fa20_xor1), .fa_or0(s_wallace_cska32_fa20_or0));
  and_gate and_gate_s_wallace_cska32_and_24_0(.a(a[24]), .b(b[0]), .out(s_wallace_cska32_and_24_0));
  and_gate and_gate_s_wallace_cska32_and_23_1(.a(a[23]), .b(b[1]), .out(s_wallace_cska32_and_23_1));
  fa fa_s_wallace_cska32_fa21_out(.a(s_wallace_cska32_fa20_or0[0]), .b(s_wallace_cska32_and_24_0[0]), .cin(s_wallace_cska32_and_23_1[0]), .fa_xor1(s_wallace_cska32_fa21_xor1), .fa_or0(s_wallace_cska32_fa21_or0));
  and_gate and_gate_s_wallace_cska32_and_25_0(.a(a[25]), .b(b[0]), .out(s_wallace_cska32_and_25_0));
  and_gate and_gate_s_wallace_cska32_and_24_1(.a(a[24]), .b(b[1]), .out(s_wallace_cska32_and_24_1));
  fa fa_s_wallace_cska32_fa22_out(.a(s_wallace_cska32_fa21_or0[0]), .b(s_wallace_cska32_and_25_0[0]), .cin(s_wallace_cska32_and_24_1[0]), .fa_xor1(s_wallace_cska32_fa22_xor1), .fa_or0(s_wallace_cska32_fa22_or0));
  and_gate and_gate_s_wallace_cska32_and_26_0(.a(a[26]), .b(b[0]), .out(s_wallace_cska32_and_26_0));
  and_gate and_gate_s_wallace_cska32_and_25_1(.a(a[25]), .b(b[1]), .out(s_wallace_cska32_and_25_1));
  fa fa_s_wallace_cska32_fa23_out(.a(s_wallace_cska32_fa22_or0[0]), .b(s_wallace_cska32_and_26_0[0]), .cin(s_wallace_cska32_and_25_1[0]), .fa_xor1(s_wallace_cska32_fa23_xor1), .fa_or0(s_wallace_cska32_fa23_or0));
  and_gate and_gate_s_wallace_cska32_and_27_0(.a(a[27]), .b(b[0]), .out(s_wallace_cska32_and_27_0));
  and_gate and_gate_s_wallace_cska32_and_26_1(.a(a[26]), .b(b[1]), .out(s_wallace_cska32_and_26_1));
  fa fa_s_wallace_cska32_fa24_out(.a(s_wallace_cska32_fa23_or0[0]), .b(s_wallace_cska32_and_27_0[0]), .cin(s_wallace_cska32_and_26_1[0]), .fa_xor1(s_wallace_cska32_fa24_xor1), .fa_or0(s_wallace_cska32_fa24_or0));
  and_gate and_gate_s_wallace_cska32_and_28_0(.a(a[28]), .b(b[0]), .out(s_wallace_cska32_and_28_0));
  and_gate and_gate_s_wallace_cska32_and_27_1(.a(a[27]), .b(b[1]), .out(s_wallace_cska32_and_27_1));
  fa fa_s_wallace_cska32_fa25_out(.a(s_wallace_cska32_fa24_or0[0]), .b(s_wallace_cska32_and_28_0[0]), .cin(s_wallace_cska32_and_27_1[0]), .fa_xor1(s_wallace_cska32_fa25_xor1), .fa_or0(s_wallace_cska32_fa25_or0));
  and_gate and_gate_s_wallace_cska32_and_29_0(.a(a[29]), .b(b[0]), .out(s_wallace_cska32_and_29_0));
  and_gate and_gate_s_wallace_cska32_and_28_1(.a(a[28]), .b(b[1]), .out(s_wallace_cska32_and_28_1));
  fa fa_s_wallace_cska32_fa26_out(.a(s_wallace_cska32_fa25_or0[0]), .b(s_wallace_cska32_and_29_0[0]), .cin(s_wallace_cska32_and_28_1[0]), .fa_xor1(s_wallace_cska32_fa26_xor1), .fa_or0(s_wallace_cska32_fa26_or0));
  and_gate and_gate_s_wallace_cska32_and_30_0(.a(a[30]), .b(b[0]), .out(s_wallace_cska32_and_30_0));
  and_gate and_gate_s_wallace_cska32_and_29_1(.a(a[29]), .b(b[1]), .out(s_wallace_cska32_and_29_1));
  fa fa_s_wallace_cska32_fa27_out(.a(s_wallace_cska32_fa26_or0[0]), .b(s_wallace_cska32_and_30_0[0]), .cin(s_wallace_cska32_and_29_1[0]), .fa_xor1(s_wallace_cska32_fa27_xor1), .fa_or0(s_wallace_cska32_fa27_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_0(.a(a[31]), .b(b[0]), .out(s_wallace_cska32_nand_31_0));
  and_gate and_gate_s_wallace_cska32_and_30_1(.a(a[30]), .b(b[1]), .out(s_wallace_cska32_and_30_1));
  fa fa_s_wallace_cska32_fa28_out(.a(s_wallace_cska32_fa27_or0[0]), .b(s_wallace_cska32_nand_31_0[0]), .cin(s_wallace_cska32_and_30_1[0]), .fa_xor1(s_wallace_cska32_fa28_xor1), .fa_or0(s_wallace_cska32_fa28_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_1(.a(a[31]), .b(b[1]), .out(s_wallace_cska32_nand_31_1));
  fa fa_s_wallace_cska32_fa29_out(.a(s_wallace_cska32_fa28_or0[0]), .b(1'b1), .cin(s_wallace_cska32_nand_31_1[0]), .fa_xor1(s_wallace_cska32_fa29_xor1), .fa_or0(s_wallace_cska32_fa29_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_2(.a(a[31]), .b(b[2]), .out(s_wallace_cska32_nand_31_2));
  and_gate and_gate_s_wallace_cska32_and_30_3(.a(a[30]), .b(b[3]), .out(s_wallace_cska32_and_30_3));
  fa fa_s_wallace_cska32_fa30_out(.a(s_wallace_cska32_fa29_or0[0]), .b(s_wallace_cska32_nand_31_2[0]), .cin(s_wallace_cska32_and_30_3[0]), .fa_xor1(s_wallace_cska32_fa30_xor1), .fa_or0(s_wallace_cska32_fa30_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_3(.a(a[31]), .b(b[3]), .out(s_wallace_cska32_nand_31_3));
  and_gate and_gate_s_wallace_cska32_and_30_4(.a(a[30]), .b(b[4]), .out(s_wallace_cska32_and_30_4));
  fa fa_s_wallace_cska32_fa31_out(.a(s_wallace_cska32_fa30_or0[0]), .b(s_wallace_cska32_nand_31_3[0]), .cin(s_wallace_cska32_and_30_4[0]), .fa_xor1(s_wallace_cska32_fa31_xor1), .fa_or0(s_wallace_cska32_fa31_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_4(.a(a[31]), .b(b[4]), .out(s_wallace_cska32_nand_31_4));
  and_gate and_gate_s_wallace_cska32_and_30_5(.a(a[30]), .b(b[5]), .out(s_wallace_cska32_and_30_5));
  fa fa_s_wallace_cska32_fa32_out(.a(s_wallace_cska32_fa31_or0[0]), .b(s_wallace_cska32_nand_31_4[0]), .cin(s_wallace_cska32_and_30_5[0]), .fa_xor1(s_wallace_cska32_fa32_xor1), .fa_or0(s_wallace_cska32_fa32_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_5(.a(a[31]), .b(b[5]), .out(s_wallace_cska32_nand_31_5));
  and_gate and_gate_s_wallace_cska32_and_30_6(.a(a[30]), .b(b[6]), .out(s_wallace_cska32_and_30_6));
  fa fa_s_wallace_cska32_fa33_out(.a(s_wallace_cska32_fa32_or0[0]), .b(s_wallace_cska32_nand_31_5[0]), .cin(s_wallace_cska32_and_30_6[0]), .fa_xor1(s_wallace_cska32_fa33_xor1), .fa_or0(s_wallace_cska32_fa33_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_6(.a(a[31]), .b(b[6]), .out(s_wallace_cska32_nand_31_6));
  and_gate and_gate_s_wallace_cska32_and_30_7(.a(a[30]), .b(b[7]), .out(s_wallace_cska32_and_30_7));
  fa fa_s_wallace_cska32_fa34_out(.a(s_wallace_cska32_fa33_or0[0]), .b(s_wallace_cska32_nand_31_6[0]), .cin(s_wallace_cska32_and_30_7[0]), .fa_xor1(s_wallace_cska32_fa34_xor1), .fa_or0(s_wallace_cska32_fa34_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_7(.a(a[31]), .b(b[7]), .out(s_wallace_cska32_nand_31_7));
  and_gate and_gate_s_wallace_cska32_and_30_8(.a(a[30]), .b(b[8]), .out(s_wallace_cska32_and_30_8));
  fa fa_s_wallace_cska32_fa35_out(.a(s_wallace_cska32_fa34_or0[0]), .b(s_wallace_cska32_nand_31_7[0]), .cin(s_wallace_cska32_and_30_8[0]), .fa_xor1(s_wallace_cska32_fa35_xor1), .fa_or0(s_wallace_cska32_fa35_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_8(.a(a[31]), .b(b[8]), .out(s_wallace_cska32_nand_31_8));
  and_gate and_gate_s_wallace_cska32_and_30_9(.a(a[30]), .b(b[9]), .out(s_wallace_cska32_and_30_9));
  fa fa_s_wallace_cska32_fa36_out(.a(s_wallace_cska32_fa35_or0[0]), .b(s_wallace_cska32_nand_31_8[0]), .cin(s_wallace_cska32_and_30_9[0]), .fa_xor1(s_wallace_cska32_fa36_xor1), .fa_or0(s_wallace_cska32_fa36_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_9(.a(a[31]), .b(b[9]), .out(s_wallace_cska32_nand_31_9));
  and_gate and_gate_s_wallace_cska32_and_30_10(.a(a[30]), .b(b[10]), .out(s_wallace_cska32_and_30_10));
  fa fa_s_wallace_cska32_fa37_out(.a(s_wallace_cska32_fa36_or0[0]), .b(s_wallace_cska32_nand_31_9[0]), .cin(s_wallace_cska32_and_30_10[0]), .fa_xor1(s_wallace_cska32_fa37_xor1), .fa_or0(s_wallace_cska32_fa37_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_10(.a(a[31]), .b(b[10]), .out(s_wallace_cska32_nand_31_10));
  and_gate and_gate_s_wallace_cska32_and_30_11(.a(a[30]), .b(b[11]), .out(s_wallace_cska32_and_30_11));
  fa fa_s_wallace_cska32_fa38_out(.a(s_wallace_cska32_fa37_or0[0]), .b(s_wallace_cska32_nand_31_10[0]), .cin(s_wallace_cska32_and_30_11[0]), .fa_xor1(s_wallace_cska32_fa38_xor1), .fa_or0(s_wallace_cska32_fa38_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_11(.a(a[31]), .b(b[11]), .out(s_wallace_cska32_nand_31_11));
  and_gate and_gate_s_wallace_cska32_and_30_12(.a(a[30]), .b(b[12]), .out(s_wallace_cska32_and_30_12));
  fa fa_s_wallace_cska32_fa39_out(.a(s_wallace_cska32_fa38_or0[0]), .b(s_wallace_cska32_nand_31_11[0]), .cin(s_wallace_cska32_and_30_12[0]), .fa_xor1(s_wallace_cska32_fa39_xor1), .fa_or0(s_wallace_cska32_fa39_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_12(.a(a[31]), .b(b[12]), .out(s_wallace_cska32_nand_31_12));
  and_gate and_gate_s_wallace_cska32_and_30_13(.a(a[30]), .b(b[13]), .out(s_wallace_cska32_and_30_13));
  fa fa_s_wallace_cska32_fa40_out(.a(s_wallace_cska32_fa39_or0[0]), .b(s_wallace_cska32_nand_31_12[0]), .cin(s_wallace_cska32_and_30_13[0]), .fa_xor1(s_wallace_cska32_fa40_xor1), .fa_or0(s_wallace_cska32_fa40_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_13(.a(a[31]), .b(b[13]), .out(s_wallace_cska32_nand_31_13));
  and_gate and_gate_s_wallace_cska32_and_30_14(.a(a[30]), .b(b[14]), .out(s_wallace_cska32_and_30_14));
  fa fa_s_wallace_cska32_fa41_out(.a(s_wallace_cska32_fa40_or0[0]), .b(s_wallace_cska32_nand_31_13[0]), .cin(s_wallace_cska32_and_30_14[0]), .fa_xor1(s_wallace_cska32_fa41_xor1), .fa_or0(s_wallace_cska32_fa41_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_14(.a(a[31]), .b(b[14]), .out(s_wallace_cska32_nand_31_14));
  and_gate and_gate_s_wallace_cska32_and_30_15(.a(a[30]), .b(b[15]), .out(s_wallace_cska32_and_30_15));
  fa fa_s_wallace_cska32_fa42_out(.a(s_wallace_cska32_fa41_or0[0]), .b(s_wallace_cska32_nand_31_14[0]), .cin(s_wallace_cska32_and_30_15[0]), .fa_xor1(s_wallace_cska32_fa42_xor1), .fa_or0(s_wallace_cska32_fa42_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_15(.a(a[31]), .b(b[15]), .out(s_wallace_cska32_nand_31_15));
  and_gate and_gate_s_wallace_cska32_and_30_16(.a(a[30]), .b(b[16]), .out(s_wallace_cska32_and_30_16));
  fa fa_s_wallace_cska32_fa43_out(.a(s_wallace_cska32_fa42_or0[0]), .b(s_wallace_cska32_nand_31_15[0]), .cin(s_wallace_cska32_and_30_16[0]), .fa_xor1(s_wallace_cska32_fa43_xor1), .fa_or0(s_wallace_cska32_fa43_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_16(.a(a[31]), .b(b[16]), .out(s_wallace_cska32_nand_31_16));
  and_gate and_gate_s_wallace_cska32_and_30_17(.a(a[30]), .b(b[17]), .out(s_wallace_cska32_and_30_17));
  fa fa_s_wallace_cska32_fa44_out(.a(s_wallace_cska32_fa43_or0[0]), .b(s_wallace_cska32_nand_31_16[0]), .cin(s_wallace_cska32_and_30_17[0]), .fa_xor1(s_wallace_cska32_fa44_xor1), .fa_or0(s_wallace_cska32_fa44_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_17(.a(a[31]), .b(b[17]), .out(s_wallace_cska32_nand_31_17));
  and_gate and_gate_s_wallace_cska32_and_30_18(.a(a[30]), .b(b[18]), .out(s_wallace_cska32_and_30_18));
  fa fa_s_wallace_cska32_fa45_out(.a(s_wallace_cska32_fa44_or0[0]), .b(s_wallace_cska32_nand_31_17[0]), .cin(s_wallace_cska32_and_30_18[0]), .fa_xor1(s_wallace_cska32_fa45_xor1), .fa_or0(s_wallace_cska32_fa45_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_18(.a(a[31]), .b(b[18]), .out(s_wallace_cska32_nand_31_18));
  and_gate and_gate_s_wallace_cska32_and_30_19(.a(a[30]), .b(b[19]), .out(s_wallace_cska32_and_30_19));
  fa fa_s_wallace_cska32_fa46_out(.a(s_wallace_cska32_fa45_or0[0]), .b(s_wallace_cska32_nand_31_18[0]), .cin(s_wallace_cska32_and_30_19[0]), .fa_xor1(s_wallace_cska32_fa46_xor1), .fa_or0(s_wallace_cska32_fa46_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_19(.a(a[31]), .b(b[19]), .out(s_wallace_cska32_nand_31_19));
  and_gate and_gate_s_wallace_cska32_and_30_20(.a(a[30]), .b(b[20]), .out(s_wallace_cska32_and_30_20));
  fa fa_s_wallace_cska32_fa47_out(.a(s_wallace_cska32_fa46_or0[0]), .b(s_wallace_cska32_nand_31_19[0]), .cin(s_wallace_cska32_and_30_20[0]), .fa_xor1(s_wallace_cska32_fa47_xor1), .fa_or0(s_wallace_cska32_fa47_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_20(.a(a[31]), .b(b[20]), .out(s_wallace_cska32_nand_31_20));
  and_gate and_gate_s_wallace_cska32_and_30_21(.a(a[30]), .b(b[21]), .out(s_wallace_cska32_and_30_21));
  fa fa_s_wallace_cska32_fa48_out(.a(s_wallace_cska32_fa47_or0[0]), .b(s_wallace_cska32_nand_31_20[0]), .cin(s_wallace_cska32_and_30_21[0]), .fa_xor1(s_wallace_cska32_fa48_xor1), .fa_or0(s_wallace_cska32_fa48_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_21(.a(a[31]), .b(b[21]), .out(s_wallace_cska32_nand_31_21));
  and_gate and_gate_s_wallace_cska32_and_30_22(.a(a[30]), .b(b[22]), .out(s_wallace_cska32_and_30_22));
  fa fa_s_wallace_cska32_fa49_out(.a(s_wallace_cska32_fa48_or0[0]), .b(s_wallace_cska32_nand_31_21[0]), .cin(s_wallace_cska32_and_30_22[0]), .fa_xor1(s_wallace_cska32_fa49_xor1), .fa_or0(s_wallace_cska32_fa49_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_22(.a(a[31]), .b(b[22]), .out(s_wallace_cska32_nand_31_22));
  and_gate and_gate_s_wallace_cska32_and_30_23(.a(a[30]), .b(b[23]), .out(s_wallace_cska32_and_30_23));
  fa fa_s_wallace_cska32_fa50_out(.a(s_wallace_cska32_fa49_or0[0]), .b(s_wallace_cska32_nand_31_22[0]), .cin(s_wallace_cska32_and_30_23[0]), .fa_xor1(s_wallace_cska32_fa50_xor1), .fa_or0(s_wallace_cska32_fa50_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_23(.a(a[31]), .b(b[23]), .out(s_wallace_cska32_nand_31_23));
  and_gate and_gate_s_wallace_cska32_and_30_24(.a(a[30]), .b(b[24]), .out(s_wallace_cska32_and_30_24));
  fa fa_s_wallace_cska32_fa51_out(.a(s_wallace_cska32_fa50_or0[0]), .b(s_wallace_cska32_nand_31_23[0]), .cin(s_wallace_cska32_and_30_24[0]), .fa_xor1(s_wallace_cska32_fa51_xor1), .fa_or0(s_wallace_cska32_fa51_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_24(.a(a[31]), .b(b[24]), .out(s_wallace_cska32_nand_31_24));
  and_gate and_gate_s_wallace_cska32_and_30_25(.a(a[30]), .b(b[25]), .out(s_wallace_cska32_and_30_25));
  fa fa_s_wallace_cska32_fa52_out(.a(s_wallace_cska32_fa51_or0[0]), .b(s_wallace_cska32_nand_31_24[0]), .cin(s_wallace_cska32_and_30_25[0]), .fa_xor1(s_wallace_cska32_fa52_xor1), .fa_or0(s_wallace_cska32_fa52_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_25(.a(a[31]), .b(b[25]), .out(s_wallace_cska32_nand_31_25));
  and_gate and_gate_s_wallace_cska32_and_30_26(.a(a[30]), .b(b[26]), .out(s_wallace_cska32_and_30_26));
  fa fa_s_wallace_cska32_fa53_out(.a(s_wallace_cska32_fa52_or0[0]), .b(s_wallace_cska32_nand_31_25[0]), .cin(s_wallace_cska32_and_30_26[0]), .fa_xor1(s_wallace_cska32_fa53_xor1), .fa_or0(s_wallace_cska32_fa53_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_26(.a(a[31]), .b(b[26]), .out(s_wallace_cska32_nand_31_26));
  and_gate and_gate_s_wallace_cska32_and_30_27(.a(a[30]), .b(b[27]), .out(s_wallace_cska32_and_30_27));
  fa fa_s_wallace_cska32_fa54_out(.a(s_wallace_cska32_fa53_or0[0]), .b(s_wallace_cska32_nand_31_26[0]), .cin(s_wallace_cska32_and_30_27[0]), .fa_xor1(s_wallace_cska32_fa54_xor1), .fa_or0(s_wallace_cska32_fa54_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_27(.a(a[31]), .b(b[27]), .out(s_wallace_cska32_nand_31_27));
  and_gate and_gate_s_wallace_cska32_and_30_28(.a(a[30]), .b(b[28]), .out(s_wallace_cska32_and_30_28));
  fa fa_s_wallace_cska32_fa55_out(.a(s_wallace_cska32_fa54_or0[0]), .b(s_wallace_cska32_nand_31_27[0]), .cin(s_wallace_cska32_and_30_28[0]), .fa_xor1(s_wallace_cska32_fa55_xor1), .fa_or0(s_wallace_cska32_fa55_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_28(.a(a[31]), .b(b[28]), .out(s_wallace_cska32_nand_31_28));
  and_gate and_gate_s_wallace_cska32_and_30_29(.a(a[30]), .b(b[29]), .out(s_wallace_cska32_and_30_29));
  fa fa_s_wallace_cska32_fa56_out(.a(s_wallace_cska32_fa55_or0[0]), .b(s_wallace_cska32_nand_31_28[0]), .cin(s_wallace_cska32_and_30_29[0]), .fa_xor1(s_wallace_cska32_fa56_xor1), .fa_or0(s_wallace_cska32_fa56_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_29(.a(a[31]), .b(b[29]), .out(s_wallace_cska32_nand_31_29));
  and_gate and_gate_s_wallace_cska32_and_30_30(.a(a[30]), .b(b[30]), .out(s_wallace_cska32_and_30_30));
  fa fa_s_wallace_cska32_fa57_out(.a(s_wallace_cska32_fa56_or0[0]), .b(s_wallace_cska32_nand_31_29[0]), .cin(s_wallace_cska32_and_30_30[0]), .fa_xor1(s_wallace_cska32_fa57_xor1), .fa_or0(s_wallace_cska32_fa57_or0));
  and_gate and_gate_s_wallace_cska32_and_1_2(.a(a[1]), .b(b[2]), .out(s_wallace_cska32_and_1_2));
  and_gate and_gate_s_wallace_cska32_and_0_3(.a(a[0]), .b(b[3]), .out(s_wallace_cska32_and_0_3));
  ha ha_s_wallace_cska32_ha1_out(.a(s_wallace_cska32_and_1_2[0]), .b(s_wallace_cska32_and_0_3[0]), .ha_xor0(s_wallace_cska32_ha1_xor0), .ha_and0(s_wallace_cska32_ha1_and0));
  and_gate and_gate_s_wallace_cska32_and_2_2(.a(a[2]), .b(b[2]), .out(s_wallace_cska32_and_2_2));
  and_gate and_gate_s_wallace_cska32_and_1_3(.a(a[1]), .b(b[3]), .out(s_wallace_cska32_and_1_3));
  fa fa_s_wallace_cska32_fa58_out(.a(s_wallace_cska32_ha1_and0[0]), .b(s_wallace_cska32_and_2_2[0]), .cin(s_wallace_cska32_and_1_3[0]), .fa_xor1(s_wallace_cska32_fa58_xor1), .fa_or0(s_wallace_cska32_fa58_or0));
  and_gate and_gate_s_wallace_cska32_and_3_2(.a(a[3]), .b(b[2]), .out(s_wallace_cska32_and_3_2));
  and_gate and_gate_s_wallace_cska32_and_2_3(.a(a[2]), .b(b[3]), .out(s_wallace_cska32_and_2_3));
  fa fa_s_wallace_cska32_fa59_out(.a(s_wallace_cska32_fa58_or0[0]), .b(s_wallace_cska32_and_3_2[0]), .cin(s_wallace_cska32_and_2_3[0]), .fa_xor1(s_wallace_cska32_fa59_xor1), .fa_or0(s_wallace_cska32_fa59_or0));
  and_gate and_gate_s_wallace_cska32_and_4_2(.a(a[4]), .b(b[2]), .out(s_wallace_cska32_and_4_2));
  and_gate and_gate_s_wallace_cska32_and_3_3(.a(a[3]), .b(b[3]), .out(s_wallace_cska32_and_3_3));
  fa fa_s_wallace_cska32_fa60_out(.a(s_wallace_cska32_fa59_or0[0]), .b(s_wallace_cska32_and_4_2[0]), .cin(s_wallace_cska32_and_3_3[0]), .fa_xor1(s_wallace_cska32_fa60_xor1), .fa_or0(s_wallace_cska32_fa60_or0));
  and_gate and_gate_s_wallace_cska32_and_5_2(.a(a[5]), .b(b[2]), .out(s_wallace_cska32_and_5_2));
  and_gate and_gate_s_wallace_cska32_and_4_3(.a(a[4]), .b(b[3]), .out(s_wallace_cska32_and_4_3));
  fa fa_s_wallace_cska32_fa61_out(.a(s_wallace_cska32_fa60_or0[0]), .b(s_wallace_cska32_and_5_2[0]), .cin(s_wallace_cska32_and_4_3[0]), .fa_xor1(s_wallace_cska32_fa61_xor1), .fa_or0(s_wallace_cska32_fa61_or0));
  and_gate and_gate_s_wallace_cska32_and_6_2(.a(a[6]), .b(b[2]), .out(s_wallace_cska32_and_6_2));
  and_gate and_gate_s_wallace_cska32_and_5_3(.a(a[5]), .b(b[3]), .out(s_wallace_cska32_and_5_3));
  fa fa_s_wallace_cska32_fa62_out(.a(s_wallace_cska32_fa61_or0[0]), .b(s_wallace_cska32_and_6_2[0]), .cin(s_wallace_cska32_and_5_3[0]), .fa_xor1(s_wallace_cska32_fa62_xor1), .fa_or0(s_wallace_cska32_fa62_or0));
  and_gate and_gate_s_wallace_cska32_and_7_2(.a(a[7]), .b(b[2]), .out(s_wallace_cska32_and_7_2));
  and_gate and_gate_s_wallace_cska32_and_6_3(.a(a[6]), .b(b[3]), .out(s_wallace_cska32_and_6_3));
  fa fa_s_wallace_cska32_fa63_out(.a(s_wallace_cska32_fa62_or0[0]), .b(s_wallace_cska32_and_7_2[0]), .cin(s_wallace_cska32_and_6_3[0]), .fa_xor1(s_wallace_cska32_fa63_xor1), .fa_or0(s_wallace_cska32_fa63_or0));
  and_gate and_gate_s_wallace_cska32_and_8_2(.a(a[8]), .b(b[2]), .out(s_wallace_cska32_and_8_2));
  and_gate and_gate_s_wallace_cska32_and_7_3(.a(a[7]), .b(b[3]), .out(s_wallace_cska32_and_7_3));
  fa fa_s_wallace_cska32_fa64_out(.a(s_wallace_cska32_fa63_or0[0]), .b(s_wallace_cska32_and_8_2[0]), .cin(s_wallace_cska32_and_7_3[0]), .fa_xor1(s_wallace_cska32_fa64_xor1), .fa_or0(s_wallace_cska32_fa64_or0));
  and_gate and_gate_s_wallace_cska32_and_9_2(.a(a[9]), .b(b[2]), .out(s_wallace_cska32_and_9_2));
  and_gate and_gate_s_wallace_cska32_and_8_3(.a(a[8]), .b(b[3]), .out(s_wallace_cska32_and_8_3));
  fa fa_s_wallace_cska32_fa65_out(.a(s_wallace_cska32_fa64_or0[0]), .b(s_wallace_cska32_and_9_2[0]), .cin(s_wallace_cska32_and_8_3[0]), .fa_xor1(s_wallace_cska32_fa65_xor1), .fa_or0(s_wallace_cska32_fa65_or0));
  and_gate and_gate_s_wallace_cska32_and_10_2(.a(a[10]), .b(b[2]), .out(s_wallace_cska32_and_10_2));
  and_gate and_gate_s_wallace_cska32_and_9_3(.a(a[9]), .b(b[3]), .out(s_wallace_cska32_and_9_3));
  fa fa_s_wallace_cska32_fa66_out(.a(s_wallace_cska32_fa65_or0[0]), .b(s_wallace_cska32_and_10_2[0]), .cin(s_wallace_cska32_and_9_3[0]), .fa_xor1(s_wallace_cska32_fa66_xor1), .fa_or0(s_wallace_cska32_fa66_or0));
  and_gate and_gate_s_wallace_cska32_and_11_2(.a(a[11]), .b(b[2]), .out(s_wallace_cska32_and_11_2));
  and_gate and_gate_s_wallace_cska32_and_10_3(.a(a[10]), .b(b[3]), .out(s_wallace_cska32_and_10_3));
  fa fa_s_wallace_cska32_fa67_out(.a(s_wallace_cska32_fa66_or0[0]), .b(s_wallace_cska32_and_11_2[0]), .cin(s_wallace_cska32_and_10_3[0]), .fa_xor1(s_wallace_cska32_fa67_xor1), .fa_or0(s_wallace_cska32_fa67_or0));
  and_gate and_gate_s_wallace_cska32_and_12_2(.a(a[12]), .b(b[2]), .out(s_wallace_cska32_and_12_2));
  and_gate and_gate_s_wallace_cska32_and_11_3(.a(a[11]), .b(b[3]), .out(s_wallace_cska32_and_11_3));
  fa fa_s_wallace_cska32_fa68_out(.a(s_wallace_cska32_fa67_or0[0]), .b(s_wallace_cska32_and_12_2[0]), .cin(s_wallace_cska32_and_11_3[0]), .fa_xor1(s_wallace_cska32_fa68_xor1), .fa_or0(s_wallace_cska32_fa68_or0));
  and_gate and_gate_s_wallace_cska32_and_13_2(.a(a[13]), .b(b[2]), .out(s_wallace_cska32_and_13_2));
  and_gate and_gate_s_wallace_cska32_and_12_3(.a(a[12]), .b(b[3]), .out(s_wallace_cska32_and_12_3));
  fa fa_s_wallace_cska32_fa69_out(.a(s_wallace_cska32_fa68_or0[0]), .b(s_wallace_cska32_and_13_2[0]), .cin(s_wallace_cska32_and_12_3[0]), .fa_xor1(s_wallace_cska32_fa69_xor1), .fa_or0(s_wallace_cska32_fa69_or0));
  and_gate and_gate_s_wallace_cska32_and_14_2(.a(a[14]), .b(b[2]), .out(s_wallace_cska32_and_14_2));
  and_gate and_gate_s_wallace_cska32_and_13_3(.a(a[13]), .b(b[3]), .out(s_wallace_cska32_and_13_3));
  fa fa_s_wallace_cska32_fa70_out(.a(s_wallace_cska32_fa69_or0[0]), .b(s_wallace_cska32_and_14_2[0]), .cin(s_wallace_cska32_and_13_3[0]), .fa_xor1(s_wallace_cska32_fa70_xor1), .fa_or0(s_wallace_cska32_fa70_or0));
  and_gate and_gate_s_wallace_cska32_and_15_2(.a(a[15]), .b(b[2]), .out(s_wallace_cska32_and_15_2));
  and_gate and_gate_s_wallace_cska32_and_14_3(.a(a[14]), .b(b[3]), .out(s_wallace_cska32_and_14_3));
  fa fa_s_wallace_cska32_fa71_out(.a(s_wallace_cska32_fa70_or0[0]), .b(s_wallace_cska32_and_15_2[0]), .cin(s_wallace_cska32_and_14_3[0]), .fa_xor1(s_wallace_cska32_fa71_xor1), .fa_or0(s_wallace_cska32_fa71_or0));
  and_gate and_gate_s_wallace_cska32_and_16_2(.a(a[16]), .b(b[2]), .out(s_wallace_cska32_and_16_2));
  and_gate and_gate_s_wallace_cska32_and_15_3(.a(a[15]), .b(b[3]), .out(s_wallace_cska32_and_15_3));
  fa fa_s_wallace_cska32_fa72_out(.a(s_wallace_cska32_fa71_or0[0]), .b(s_wallace_cska32_and_16_2[0]), .cin(s_wallace_cska32_and_15_3[0]), .fa_xor1(s_wallace_cska32_fa72_xor1), .fa_or0(s_wallace_cska32_fa72_or0));
  and_gate and_gate_s_wallace_cska32_and_17_2(.a(a[17]), .b(b[2]), .out(s_wallace_cska32_and_17_2));
  and_gate and_gate_s_wallace_cska32_and_16_3(.a(a[16]), .b(b[3]), .out(s_wallace_cska32_and_16_3));
  fa fa_s_wallace_cska32_fa73_out(.a(s_wallace_cska32_fa72_or0[0]), .b(s_wallace_cska32_and_17_2[0]), .cin(s_wallace_cska32_and_16_3[0]), .fa_xor1(s_wallace_cska32_fa73_xor1), .fa_or0(s_wallace_cska32_fa73_or0));
  and_gate and_gate_s_wallace_cska32_and_18_2(.a(a[18]), .b(b[2]), .out(s_wallace_cska32_and_18_2));
  and_gate and_gate_s_wallace_cska32_and_17_3(.a(a[17]), .b(b[3]), .out(s_wallace_cska32_and_17_3));
  fa fa_s_wallace_cska32_fa74_out(.a(s_wallace_cska32_fa73_or0[0]), .b(s_wallace_cska32_and_18_2[0]), .cin(s_wallace_cska32_and_17_3[0]), .fa_xor1(s_wallace_cska32_fa74_xor1), .fa_or0(s_wallace_cska32_fa74_or0));
  and_gate and_gate_s_wallace_cska32_and_19_2(.a(a[19]), .b(b[2]), .out(s_wallace_cska32_and_19_2));
  and_gate and_gate_s_wallace_cska32_and_18_3(.a(a[18]), .b(b[3]), .out(s_wallace_cska32_and_18_3));
  fa fa_s_wallace_cska32_fa75_out(.a(s_wallace_cska32_fa74_or0[0]), .b(s_wallace_cska32_and_19_2[0]), .cin(s_wallace_cska32_and_18_3[0]), .fa_xor1(s_wallace_cska32_fa75_xor1), .fa_or0(s_wallace_cska32_fa75_or0));
  and_gate and_gate_s_wallace_cska32_and_20_2(.a(a[20]), .b(b[2]), .out(s_wallace_cska32_and_20_2));
  and_gate and_gate_s_wallace_cska32_and_19_3(.a(a[19]), .b(b[3]), .out(s_wallace_cska32_and_19_3));
  fa fa_s_wallace_cska32_fa76_out(.a(s_wallace_cska32_fa75_or0[0]), .b(s_wallace_cska32_and_20_2[0]), .cin(s_wallace_cska32_and_19_3[0]), .fa_xor1(s_wallace_cska32_fa76_xor1), .fa_or0(s_wallace_cska32_fa76_or0));
  and_gate and_gate_s_wallace_cska32_and_21_2(.a(a[21]), .b(b[2]), .out(s_wallace_cska32_and_21_2));
  and_gate and_gate_s_wallace_cska32_and_20_3(.a(a[20]), .b(b[3]), .out(s_wallace_cska32_and_20_3));
  fa fa_s_wallace_cska32_fa77_out(.a(s_wallace_cska32_fa76_or0[0]), .b(s_wallace_cska32_and_21_2[0]), .cin(s_wallace_cska32_and_20_3[0]), .fa_xor1(s_wallace_cska32_fa77_xor1), .fa_or0(s_wallace_cska32_fa77_or0));
  and_gate and_gate_s_wallace_cska32_and_22_2(.a(a[22]), .b(b[2]), .out(s_wallace_cska32_and_22_2));
  and_gate and_gate_s_wallace_cska32_and_21_3(.a(a[21]), .b(b[3]), .out(s_wallace_cska32_and_21_3));
  fa fa_s_wallace_cska32_fa78_out(.a(s_wallace_cska32_fa77_or0[0]), .b(s_wallace_cska32_and_22_2[0]), .cin(s_wallace_cska32_and_21_3[0]), .fa_xor1(s_wallace_cska32_fa78_xor1), .fa_or0(s_wallace_cska32_fa78_or0));
  and_gate and_gate_s_wallace_cska32_and_23_2(.a(a[23]), .b(b[2]), .out(s_wallace_cska32_and_23_2));
  and_gate and_gate_s_wallace_cska32_and_22_3(.a(a[22]), .b(b[3]), .out(s_wallace_cska32_and_22_3));
  fa fa_s_wallace_cska32_fa79_out(.a(s_wallace_cska32_fa78_or0[0]), .b(s_wallace_cska32_and_23_2[0]), .cin(s_wallace_cska32_and_22_3[0]), .fa_xor1(s_wallace_cska32_fa79_xor1), .fa_or0(s_wallace_cska32_fa79_or0));
  and_gate and_gate_s_wallace_cska32_and_24_2(.a(a[24]), .b(b[2]), .out(s_wallace_cska32_and_24_2));
  and_gate and_gate_s_wallace_cska32_and_23_3(.a(a[23]), .b(b[3]), .out(s_wallace_cska32_and_23_3));
  fa fa_s_wallace_cska32_fa80_out(.a(s_wallace_cska32_fa79_or0[0]), .b(s_wallace_cska32_and_24_2[0]), .cin(s_wallace_cska32_and_23_3[0]), .fa_xor1(s_wallace_cska32_fa80_xor1), .fa_or0(s_wallace_cska32_fa80_or0));
  and_gate and_gate_s_wallace_cska32_and_25_2(.a(a[25]), .b(b[2]), .out(s_wallace_cska32_and_25_2));
  and_gate and_gate_s_wallace_cska32_and_24_3(.a(a[24]), .b(b[3]), .out(s_wallace_cska32_and_24_3));
  fa fa_s_wallace_cska32_fa81_out(.a(s_wallace_cska32_fa80_or0[0]), .b(s_wallace_cska32_and_25_2[0]), .cin(s_wallace_cska32_and_24_3[0]), .fa_xor1(s_wallace_cska32_fa81_xor1), .fa_or0(s_wallace_cska32_fa81_or0));
  and_gate and_gate_s_wallace_cska32_and_26_2(.a(a[26]), .b(b[2]), .out(s_wallace_cska32_and_26_2));
  and_gate and_gate_s_wallace_cska32_and_25_3(.a(a[25]), .b(b[3]), .out(s_wallace_cska32_and_25_3));
  fa fa_s_wallace_cska32_fa82_out(.a(s_wallace_cska32_fa81_or0[0]), .b(s_wallace_cska32_and_26_2[0]), .cin(s_wallace_cska32_and_25_3[0]), .fa_xor1(s_wallace_cska32_fa82_xor1), .fa_or0(s_wallace_cska32_fa82_or0));
  and_gate and_gate_s_wallace_cska32_and_27_2(.a(a[27]), .b(b[2]), .out(s_wallace_cska32_and_27_2));
  and_gate and_gate_s_wallace_cska32_and_26_3(.a(a[26]), .b(b[3]), .out(s_wallace_cska32_and_26_3));
  fa fa_s_wallace_cska32_fa83_out(.a(s_wallace_cska32_fa82_or0[0]), .b(s_wallace_cska32_and_27_2[0]), .cin(s_wallace_cska32_and_26_3[0]), .fa_xor1(s_wallace_cska32_fa83_xor1), .fa_or0(s_wallace_cska32_fa83_or0));
  and_gate and_gate_s_wallace_cska32_and_28_2(.a(a[28]), .b(b[2]), .out(s_wallace_cska32_and_28_2));
  and_gate and_gate_s_wallace_cska32_and_27_3(.a(a[27]), .b(b[3]), .out(s_wallace_cska32_and_27_3));
  fa fa_s_wallace_cska32_fa84_out(.a(s_wallace_cska32_fa83_or0[0]), .b(s_wallace_cska32_and_28_2[0]), .cin(s_wallace_cska32_and_27_3[0]), .fa_xor1(s_wallace_cska32_fa84_xor1), .fa_or0(s_wallace_cska32_fa84_or0));
  and_gate and_gate_s_wallace_cska32_and_29_2(.a(a[29]), .b(b[2]), .out(s_wallace_cska32_and_29_2));
  and_gate and_gate_s_wallace_cska32_and_28_3(.a(a[28]), .b(b[3]), .out(s_wallace_cska32_and_28_3));
  fa fa_s_wallace_cska32_fa85_out(.a(s_wallace_cska32_fa84_or0[0]), .b(s_wallace_cska32_and_29_2[0]), .cin(s_wallace_cska32_and_28_3[0]), .fa_xor1(s_wallace_cska32_fa85_xor1), .fa_or0(s_wallace_cska32_fa85_or0));
  and_gate and_gate_s_wallace_cska32_and_30_2(.a(a[30]), .b(b[2]), .out(s_wallace_cska32_and_30_2));
  and_gate and_gate_s_wallace_cska32_and_29_3(.a(a[29]), .b(b[3]), .out(s_wallace_cska32_and_29_3));
  fa fa_s_wallace_cska32_fa86_out(.a(s_wallace_cska32_fa85_or0[0]), .b(s_wallace_cska32_and_30_2[0]), .cin(s_wallace_cska32_and_29_3[0]), .fa_xor1(s_wallace_cska32_fa86_xor1), .fa_or0(s_wallace_cska32_fa86_or0));
  and_gate and_gate_s_wallace_cska32_and_29_4(.a(a[29]), .b(b[4]), .out(s_wallace_cska32_and_29_4));
  and_gate and_gate_s_wallace_cska32_and_28_5(.a(a[28]), .b(b[5]), .out(s_wallace_cska32_and_28_5));
  fa fa_s_wallace_cska32_fa87_out(.a(s_wallace_cska32_fa86_or0[0]), .b(s_wallace_cska32_and_29_4[0]), .cin(s_wallace_cska32_and_28_5[0]), .fa_xor1(s_wallace_cska32_fa87_xor1), .fa_or0(s_wallace_cska32_fa87_or0));
  and_gate and_gate_s_wallace_cska32_and_29_5(.a(a[29]), .b(b[5]), .out(s_wallace_cska32_and_29_5));
  and_gate and_gate_s_wallace_cska32_and_28_6(.a(a[28]), .b(b[6]), .out(s_wallace_cska32_and_28_6));
  fa fa_s_wallace_cska32_fa88_out(.a(s_wallace_cska32_fa87_or0[0]), .b(s_wallace_cska32_and_29_5[0]), .cin(s_wallace_cska32_and_28_6[0]), .fa_xor1(s_wallace_cska32_fa88_xor1), .fa_or0(s_wallace_cska32_fa88_or0));
  and_gate and_gate_s_wallace_cska32_and_29_6(.a(a[29]), .b(b[6]), .out(s_wallace_cska32_and_29_6));
  and_gate and_gate_s_wallace_cska32_and_28_7(.a(a[28]), .b(b[7]), .out(s_wallace_cska32_and_28_7));
  fa fa_s_wallace_cska32_fa89_out(.a(s_wallace_cska32_fa88_or0[0]), .b(s_wallace_cska32_and_29_6[0]), .cin(s_wallace_cska32_and_28_7[0]), .fa_xor1(s_wallace_cska32_fa89_xor1), .fa_or0(s_wallace_cska32_fa89_or0));
  and_gate and_gate_s_wallace_cska32_and_29_7(.a(a[29]), .b(b[7]), .out(s_wallace_cska32_and_29_7));
  and_gate and_gate_s_wallace_cska32_and_28_8(.a(a[28]), .b(b[8]), .out(s_wallace_cska32_and_28_8));
  fa fa_s_wallace_cska32_fa90_out(.a(s_wallace_cska32_fa89_or0[0]), .b(s_wallace_cska32_and_29_7[0]), .cin(s_wallace_cska32_and_28_8[0]), .fa_xor1(s_wallace_cska32_fa90_xor1), .fa_or0(s_wallace_cska32_fa90_or0));
  and_gate and_gate_s_wallace_cska32_and_29_8(.a(a[29]), .b(b[8]), .out(s_wallace_cska32_and_29_8));
  and_gate and_gate_s_wallace_cska32_and_28_9(.a(a[28]), .b(b[9]), .out(s_wallace_cska32_and_28_9));
  fa fa_s_wallace_cska32_fa91_out(.a(s_wallace_cska32_fa90_or0[0]), .b(s_wallace_cska32_and_29_8[0]), .cin(s_wallace_cska32_and_28_9[0]), .fa_xor1(s_wallace_cska32_fa91_xor1), .fa_or0(s_wallace_cska32_fa91_or0));
  and_gate and_gate_s_wallace_cska32_and_29_9(.a(a[29]), .b(b[9]), .out(s_wallace_cska32_and_29_9));
  and_gate and_gate_s_wallace_cska32_and_28_10(.a(a[28]), .b(b[10]), .out(s_wallace_cska32_and_28_10));
  fa fa_s_wallace_cska32_fa92_out(.a(s_wallace_cska32_fa91_or0[0]), .b(s_wallace_cska32_and_29_9[0]), .cin(s_wallace_cska32_and_28_10[0]), .fa_xor1(s_wallace_cska32_fa92_xor1), .fa_or0(s_wallace_cska32_fa92_or0));
  and_gate and_gate_s_wallace_cska32_and_29_10(.a(a[29]), .b(b[10]), .out(s_wallace_cska32_and_29_10));
  and_gate and_gate_s_wallace_cska32_and_28_11(.a(a[28]), .b(b[11]), .out(s_wallace_cska32_and_28_11));
  fa fa_s_wallace_cska32_fa93_out(.a(s_wallace_cska32_fa92_or0[0]), .b(s_wallace_cska32_and_29_10[0]), .cin(s_wallace_cska32_and_28_11[0]), .fa_xor1(s_wallace_cska32_fa93_xor1), .fa_or0(s_wallace_cska32_fa93_or0));
  and_gate and_gate_s_wallace_cska32_and_29_11(.a(a[29]), .b(b[11]), .out(s_wallace_cska32_and_29_11));
  and_gate and_gate_s_wallace_cska32_and_28_12(.a(a[28]), .b(b[12]), .out(s_wallace_cska32_and_28_12));
  fa fa_s_wallace_cska32_fa94_out(.a(s_wallace_cska32_fa93_or0[0]), .b(s_wallace_cska32_and_29_11[0]), .cin(s_wallace_cska32_and_28_12[0]), .fa_xor1(s_wallace_cska32_fa94_xor1), .fa_or0(s_wallace_cska32_fa94_or0));
  and_gate and_gate_s_wallace_cska32_and_29_12(.a(a[29]), .b(b[12]), .out(s_wallace_cska32_and_29_12));
  and_gate and_gate_s_wallace_cska32_and_28_13(.a(a[28]), .b(b[13]), .out(s_wallace_cska32_and_28_13));
  fa fa_s_wallace_cska32_fa95_out(.a(s_wallace_cska32_fa94_or0[0]), .b(s_wallace_cska32_and_29_12[0]), .cin(s_wallace_cska32_and_28_13[0]), .fa_xor1(s_wallace_cska32_fa95_xor1), .fa_or0(s_wallace_cska32_fa95_or0));
  and_gate and_gate_s_wallace_cska32_and_29_13(.a(a[29]), .b(b[13]), .out(s_wallace_cska32_and_29_13));
  and_gate and_gate_s_wallace_cska32_and_28_14(.a(a[28]), .b(b[14]), .out(s_wallace_cska32_and_28_14));
  fa fa_s_wallace_cska32_fa96_out(.a(s_wallace_cska32_fa95_or0[0]), .b(s_wallace_cska32_and_29_13[0]), .cin(s_wallace_cska32_and_28_14[0]), .fa_xor1(s_wallace_cska32_fa96_xor1), .fa_or0(s_wallace_cska32_fa96_or0));
  and_gate and_gate_s_wallace_cska32_and_29_14(.a(a[29]), .b(b[14]), .out(s_wallace_cska32_and_29_14));
  and_gate and_gate_s_wallace_cska32_and_28_15(.a(a[28]), .b(b[15]), .out(s_wallace_cska32_and_28_15));
  fa fa_s_wallace_cska32_fa97_out(.a(s_wallace_cska32_fa96_or0[0]), .b(s_wallace_cska32_and_29_14[0]), .cin(s_wallace_cska32_and_28_15[0]), .fa_xor1(s_wallace_cska32_fa97_xor1), .fa_or0(s_wallace_cska32_fa97_or0));
  and_gate and_gate_s_wallace_cska32_and_29_15(.a(a[29]), .b(b[15]), .out(s_wallace_cska32_and_29_15));
  and_gate and_gate_s_wallace_cska32_and_28_16(.a(a[28]), .b(b[16]), .out(s_wallace_cska32_and_28_16));
  fa fa_s_wallace_cska32_fa98_out(.a(s_wallace_cska32_fa97_or0[0]), .b(s_wallace_cska32_and_29_15[0]), .cin(s_wallace_cska32_and_28_16[0]), .fa_xor1(s_wallace_cska32_fa98_xor1), .fa_or0(s_wallace_cska32_fa98_or0));
  and_gate and_gate_s_wallace_cska32_and_29_16(.a(a[29]), .b(b[16]), .out(s_wallace_cska32_and_29_16));
  and_gate and_gate_s_wallace_cska32_and_28_17(.a(a[28]), .b(b[17]), .out(s_wallace_cska32_and_28_17));
  fa fa_s_wallace_cska32_fa99_out(.a(s_wallace_cska32_fa98_or0[0]), .b(s_wallace_cska32_and_29_16[0]), .cin(s_wallace_cska32_and_28_17[0]), .fa_xor1(s_wallace_cska32_fa99_xor1), .fa_or0(s_wallace_cska32_fa99_or0));
  and_gate and_gate_s_wallace_cska32_and_29_17(.a(a[29]), .b(b[17]), .out(s_wallace_cska32_and_29_17));
  and_gate and_gate_s_wallace_cska32_and_28_18(.a(a[28]), .b(b[18]), .out(s_wallace_cska32_and_28_18));
  fa fa_s_wallace_cska32_fa100_out(.a(s_wallace_cska32_fa99_or0[0]), .b(s_wallace_cska32_and_29_17[0]), .cin(s_wallace_cska32_and_28_18[0]), .fa_xor1(s_wallace_cska32_fa100_xor1), .fa_or0(s_wallace_cska32_fa100_or0));
  and_gate and_gate_s_wallace_cska32_and_29_18(.a(a[29]), .b(b[18]), .out(s_wallace_cska32_and_29_18));
  and_gate and_gate_s_wallace_cska32_and_28_19(.a(a[28]), .b(b[19]), .out(s_wallace_cska32_and_28_19));
  fa fa_s_wallace_cska32_fa101_out(.a(s_wallace_cska32_fa100_or0[0]), .b(s_wallace_cska32_and_29_18[0]), .cin(s_wallace_cska32_and_28_19[0]), .fa_xor1(s_wallace_cska32_fa101_xor1), .fa_or0(s_wallace_cska32_fa101_or0));
  and_gate and_gate_s_wallace_cska32_and_29_19(.a(a[29]), .b(b[19]), .out(s_wallace_cska32_and_29_19));
  and_gate and_gate_s_wallace_cska32_and_28_20(.a(a[28]), .b(b[20]), .out(s_wallace_cska32_and_28_20));
  fa fa_s_wallace_cska32_fa102_out(.a(s_wallace_cska32_fa101_or0[0]), .b(s_wallace_cska32_and_29_19[0]), .cin(s_wallace_cska32_and_28_20[0]), .fa_xor1(s_wallace_cska32_fa102_xor1), .fa_or0(s_wallace_cska32_fa102_or0));
  and_gate and_gate_s_wallace_cska32_and_29_20(.a(a[29]), .b(b[20]), .out(s_wallace_cska32_and_29_20));
  and_gate and_gate_s_wallace_cska32_and_28_21(.a(a[28]), .b(b[21]), .out(s_wallace_cska32_and_28_21));
  fa fa_s_wallace_cska32_fa103_out(.a(s_wallace_cska32_fa102_or0[0]), .b(s_wallace_cska32_and_29_20[0]), .cin(s_wallace_cska32_and_28_21[0]), .fa_xor1(s_wallace_cska32_fa103_xor1), .fa_or0(s_wallace_cska32_fa103_or0));
  and_gate and_gate_s_wallace_cska32_and_29_21(.a(a[29]), .b(b[21]), .out(s_wallace_cska32_and_29_21));
  and_gate and_gate_s_wallace_cska32_and_28_22(.a(a[28]), .b(b[22]), .out(s_wallace_cska32_and_28_22));
  fa fa_s_wallace_cska32_fa104_out(.a(s_wallace_cska32_fa103_or0[0]), .b(s_wallace_cska32_and_29_21[0]), .cin(s_wallace_cska32_and_28_22[0]), .fa_xor1(s_wallace_cska32_fa104_xor1), .fa_or0(s_wallace_cska32_fa104_or0));
  and_gate and_gate_s_wallace_cska32_and_29_22(.a(a[29]), .b(b[22]), .out(s_wallace_cska32_and_29_22));
  and_gate and_gate_s_wallace_cska32_and_28_23(.a(a[28]), .b(b[23]), .out(s_wallace_cska32_and_28_23));
  fa fa_s_wallace_cska32_fa105_out(.a(s_wallace_cska32_fa104_or0[0]), .b(s_wallace_cska32_and_29_22[0]), .cin(s_wallace_cska32_and_28_23[0]), .fa_xor1(s_wallace_cska32_fa105_xor1), .fa_or0(s_wallace_cska32_fa105_or0));
  and_gate and_gate_s_wallace_cska32_and_29_23(.a(a[29]), .b(b[23]), .out(s_wallace_cska32_and_29_23));
  and_gate and_gate_s_wallace_cska32_and_28_24(.a(a[28]), .b(b[24]), .out(s_wallace_cska32_and_28_24));
  fa fa_s_wallace_cska32_fa106_out(.a(s_wallace_cska32_fa105_or0[0]), .b(s_wallace_cska32_and_29_23[0]), .cin(s_wallace_cska32_and_28_24[0]), .fa_xor1(s_wallace_cska32_fa106_xor1), .fa_or0(s_wallace_cska32_fa106_or0));
  and_gate and_gate_s_wallace_cska32_and_29_24(.a(a[29]), .b(b[24]), .out(s_wallace_cska32_and_29_24));
  and_gate and_gate_s_wallace_cska32_and_28_25(.a(a[28]), .b(b[25]), .out(s_wallace_cska32_and_28_25));
  fa fa_s_wallace_cska32_fa107_out(.a(s_wallace_cska32_fa106_or0[0]), .b(s_wallace_cska32_and_29_24[0]), .cin(s_wallace_cska32_and_28_25[0]), .fa_xor1(s_wallace_cska32_fa107_xor1), .fa_or0(s_wallace_cska32_fa107_or0));
  and_gate and_gate_s_wallace_cska32_and_29_25(.a(a[29]), .b(b[25]), .out(s_wallace_cska32_and_29_25));
  and_gate and_gate_s_wallace_cska32_and_28_26(.a(a[28]), .b(b[26]), .out(s_wallace_cska32_and_28_26));
  fa fa_s_wallace_cska32_fa108_out(.a(s_wallace_cska32_fa107_or0[0]), .b(s_wallace_cska32_and_29_25[0]), .cin(s_wallace_cska32_and_28_26[0]), .fa_xor1(s_wallace_cska32_fa108_xor1), .fa_or0(s_wallace_cska32_fa108_or0));
  and_gate and_gate_s_wallace_cska32_and_29_26(.a(a[29]), .b(b[26]), .out(s_wallace_cska32_and_29_26));
  and_gate and_gate_s_wallace_cska32_and_28_27(.a(a[28]), .b(b[27]), .out(s_wallace_cska32_and_28_27));
  fa fa_s_wallace_cska32_fa109_out(.a(s_wallace_cska32_fa108_or0[0]), .b(s_wallace_cska32_and_29_26[0]), .cin(s_wallace_cska32_and_28_27[0]), .fa_xor1(s_wallace_cska32_fa109_xor1), .fa_or0(s_wallace_cska32_fa109_or0));
  and_gate and_gate_s_wallace_cska32_and_29_27(.a(a[29]), .b(b[27]), .out(s_wallace_cska32_and_29_27));
  and_gate and_gate_s_wallace_cska32_and_28_28(.a(a[28]), .b(b[28]), .out(s_wallace_cska32_and_28_28));
  fa fa_s_wallace_cska32_fa110_out(.a(s_wallace_cska32_fa109_or0[0]), .b(s_wallace_cska32_and_29_27[0]), .cin(s_wallace_cska32_and_28_28[0]), .fa_xor1(s_wallace_cska32_fa110_xor1), .fa_or0(s_wallace_cska32_fa110_or0));
  and_gate and_gate_s_wallace_cska32_and_29_28(.a(a[29]), .b(b[28]), .out(s_wallace_cska32_and_29_28));
  and_gate and_gate_s_wallace_cska32_and_28_29(.a(a[28]), .b(b[29]), .out(s_wallace_cska32_and_28_29));
  fa fa_s_wallace_cska32_fa111_out(.a(s_wallace_cska32_fa110_or0[0]), .b(s_wallace_cska32_and_29_28[0]), .cin(s_wallace_cska32_and_28_29[0]), .fa_xor1(s_wallace_cska32_fa111_xor1), .fa_or0(s_wallace_cska32_fa111_or0));
  and_gate and_gate_s_wallace_cska32_and_29_29(.a(a[29]), .b(b[29]), .out(s_wallace_cska32_and_29_29));
  and_gate and_gate_s_wallace_cska32_and_28_30(.a(a[28]), .b(b[30]), .out(s_wallace_cska32_and_28_30));
  fa fa_s_wallace_cska32_fa112_out(.a(s_wallace_cska32_fa111_or0[0]), .b(s_wallace_cska32_and_29_29[0]), .cin(s_wallace_cska32_and_28_30[0]), .fa_xor1(s_wallace_cska32_fa112_xor1), .fa_or0(s_wallace_cska32_fa112_or0));
  and_gate and_gate_s_wallace_cska32_and_29_30(.a(a[29]), .b(b[30]), .out(s_wallace_cska32_and_29_30));
  nand_gate nand_gate_s_wallace_cska32_nand_28_31(.a(a[28]), .b(b[31]), .out(s_wallace_cska32_nand_28_31));
  fa fa_s_wallace_cska32_fa113_out(.a(s_wallace_cska32_fa112_or0[0]), .b(s_wallace_cska32_and_29_30[0]), .cin(s_wallace_cska32_nand_28_31[0]), .fa_xor1(s_wallace_cska32_fa113_xor1), .fa_or0(s_wallace_cska32_fa113_or0));
  and_gate and_gate_s_wallace_cska32_and_0_4(.a(a[0]), .b(b[4]), .out(s_wallace_cska32_and_0_4));
  ha ha_s_wallace_cska32_ha2_out(.a(s_wallace_cska32_and_0_4[0]), .b(s_wallace_cska32_fa1_xor1[0]), .ha_xor0(s_wallace_cska32_ha2_xor0), .ha_and0(s_wallace_cska32_ha2_and0));
  and_gate and_gate_s_wallace_cska32_and_1_4(.a(a[1]), .b(b[4]), .out(s_wallace_cska32_and_1_4));
  and_gate and_gate_s_wallace_cska32_and_0_5(.a(a[0]), .b(b[5]), .out(s_wallace_cska32_and_0_5));
  fa fa_s_wallace_cska32_fa114_out(.a(s_wallace_cska32_ha2_and0[0]), .b(s_wallace_cska32_and_1_4[0]), .cin(s_wallace_cska32_and_0_5[0]), .fa_xor1(s_wallace_cska32_fa114_xor1), .fa_or0(s_wallace_cska32_fa114_or0));
  and_gate and_gate_s_wallace_cska32_and_2_4(.a(a[2]), .b(b[4]), .out(s_wallace_cska32_and_2_4));
  and_gate and_gate_s_wallace_cska32_and_1_5(.a(a[1]), .b(b[5]), .out(s_wallace_cska32_and_1_5));
  fa fa_s_wallace_cska32_fa115_out(.a(s_wallace_cska32_fa114_or0[0]), .b(s_wallace_cska32_and_2_4[0]), .cin(s_wallace_cska32_and_1_5[0]), .fa_xor1(s_wallace_cska32_fa115_xor1), .fa_or0(s_wallace_cska32_fa115_or0));
  and_gate and_gate_s_wallace_cska32_and_3_4(.a(a[3]), .b(b[4]), .out(s_wallace_cska32_and_3_4));
  and_gate and_gate_s_wallace_cska32_and_2_5(.a(a[2]), .b(b[5]), .out(s_wallace_cska32_and_2_5));
  fa fa_s_wallace_cska32_fa116_out(.a(s_wallace_cska32_fa115_or0[0]), .b(s_wallace_cska32_and_3_4[0]), .cin(s_wallace_cska32_and_2_5[0]), .fa_xor1(s_wallace_cska32_fa116_xor1), .fa_or0(s_wallace_cska32_fa116_or0));
  and_gate and_gate_s_wallace_cska32_and_4_4(.a(a[4]), .b(b[4]), .out(s_wallace_cska32_and_4_4));
  and_gate and_gate_s_wallace_cska32_and_3_5(.a(a[3]), .b(b[5]), .out(s_wallace_cska32_and_3_5));
  fa fa_s_wallace_cska32_fa117_out(.a(s_wallace_cska32_fa116_or0[0]), .b(s_wallace_cska32_and_4_4[0]), .cin(s_wallace_cska32_and_3_5[0]), .fa_xor1(s_wallace_cska32_fa117_xor1), .fa_or0(s_wallace_cska32_fa117_or0));
  and_gate and_gate_s_wallace_cska32_and_5_4(.a(a[5]), .b(b[4]), .out(s_wallace_cska32_and_5_4));
  and_gate and_gate_s_wallace_cska32_and_4_5(.a(a[4]), .b(b[5]), .out(s_wallace_cska32_and_4_5));
  fa fa_s_wallace_cska32_fa118_out(.a(s_wallace_cska32_fa117_or0[0]), .b(s_wallace_cska32_and_5_4[0]), .cin(s_wallace_cska32_and_4_5[0]), .fa_xor1(s_wallace_cska32_fa118_xor1), .fa_or0(s_wallace_cska32_fa118_or0));
  and_gate and_gate_s_wallace_cska32_and_6_4(.a(a[6]), .b(b[4]), .out(s_wallace_cska32_and_6_4));
  and_gate and_gate_s_wallace_cska32_and_5_5(.a(a[5]), .b(b[5]), .out(s_wallace_cska32_and_5_5));
  fa fa_s_wallace_cska32_fa119_out(.a(s_wallace_cska32_fa118_or0[0]), .b(s_wallace_cska32_and_6_4[0]), .cin(s_wallace_cska32_and_5_5[0]), .fa_xor1(s_wallace_cska32_fa119_xor1), .fa_or0(s_wallace_cska32_fa119_or0));
  and_gate and_gate_s_wallace_cska32_and_7_4(.a(a[7]), .b(b[4]), .out(s_wallace_cska32_and_7_4));
  and_gate and_gate_s_wallace_cska32_and_6_5(.a(a[6]), .b(b[5]), .out(s_wallace_cska32_and_6_5));
  fa fa_s_wallace_cska32_fa120_out(.a(s_wallace_cska32_fa119_or0[0]), .b(s_wallace_cska32_and_7_4[0]), .cin(s_wallace_cska32_and_6_5[0]), .fa_xor1(s_wallace_cska32_fa120_xor1), .fa_or0(s_wallace_cska32_fa120_or0));
  and_gate and_gate_s_wallace_cska32_and_8_4(.a(a[8]), .b(b[4]), .out(s_wallace_cska32_and_8_4));
  and_gate and_gate_s_wallace_cska32_and_7_5(.a(a[7]), .b(b[5]), .out(s_wallace_cska32_and_7_5));
  fa fa_s_wallace_cska32_fa121_out(.a(s_wallace_cska32_fa120_or0[0]), .b(s_wallace_cska32_and_8_4[0]), .cin(s_wallace_cska32_and_7_5[0]), .fa_xor1(s_wallace_cska32_fa121_xor1), .fa_or0(s_wallace_cska32_fa121_or0));
  and_gate and_gate_s_wallace_cska32_and_9_4(.a(a[9]), .b(b[4]), .out(s_wallace_cska32_and_9_4));
  and_gate and_gate_s_wallace_cska32_and_8_5(.a(a[8]), .b(b[5]), .out(s_wallace_cska32_and_8_5));
  fa fa_s_wallace_cska32_fa122_out(.a(s_wallace_cska32_fa121_or0[0]), .b(s_wallace_cska32_and_9_4[0]), .cin(s_wallace_cska32_and_8_5[0]), .fa_xor1(s_wallace_cska32_fa122_xor1), .fa_or0(s_wallace_cska32_fa122_or0));
  and_gate and_gate_s_wallace_cska32_and_10_4(.a(a[10]), .b(b[4]), .out(s_wallace_cska32_and_10_4));
  and_gate and_gate_s_wallace_cska32_and_9_5(.a(a[9]), .b(b[5]), .out(s_wallace_cska32_and_9_5));
  fa fa_s_wallace_cska32_fa123_out(.a(s_wallace_cska32_fa122_or0[0]), .b(s_wallace_cska32_and_10_4[0]), .cin(s_wallace_cska32_and_9_5[0]), .fa_xor1(s_wallace_cska32_fa123_xor1), .fa_or0(s_wallace_cska32_fa123_or0));
  and_gate and_gate_s_wallace_cska32_and_11_4(.a(a[11]), .b(b[4]), .out(s_wallace_cska32_and_11_4));
  and_gate and_gate_s_wallace_cska32_and_10_5(.a(a[10]), .b(b[5]), .out(s_wallace_cska32_and_10_5));
  fa fa_s_wallace_cska32_fa124_out(.a(s_wallace_cska32_fa123_or0[0]), .b(s_wallace_cska32_and_11_4[0]), .cin(s_wallace_cska32_and_10_5[0]), .fa_xor1(s_wallace_cska32_fa124_xor1), .fa_or0(s_wallace_cska32_fa124_or0));
  and_gate and_gate_s_wallace_cska32_and_12_4(.a(a[12]), .b(b[4]), .out(s_wallace_cska32_and_12_4));
  and_gate and_gate_s_wallace_cska32_and_11_5(.a(a[11]), .b(b[5]), .out(s_wallace_cska32_and_11_5));
  fa fa_s_wallace_cska32_fa125_out(.a(s_wallace_cska32_fa124_or0[0]), .b(s_wallace_cska32_and_12_4[0]), .cin(s_wallace_cska32_and_11_5[0]), .fa_xor1(s_wallace_cska32_fa125_xor1), .fa_or0(s_wallace_cska32_fa125_or0));
  and_gate and_gate_s_wallace_cska32_and_13_4(.a(a[13]), .b(b[4]), .out(s_wallace_cska32_and_13_4));
  and_gate and_gate_s_wallace_cska32_and_12_5(.a(a[12]), .b(b[5]), .out(s_wallace_cska32_and_12_5));
  fa fa_s_wallace_cska32_fa126_out(.a(s_wallace_cska32_fa125_or0[0]), .b(s_wallace_cska32_and_13_4[0]), .cin(s_wallace_cska32_and_12_5[0]), .fa_xor1(s_wallace_cska32_fa126_xor1), .fa_or0(s_wallace_cska32_fa126_or0));
  and_gate and_gate_s_wallace_cska32_and_14_4(.a(a[14]), .b(b[4]), .out(s_wallace_cska32_and_14_4));
  and_gate and_gate_s_wallace_cska32_and_13_5(.a(a[13]), .b(b[5]), .out(s_wallace_cska32_and_13_5));
  fa fa_s_wallace_cska32_fa127_out(.a(s_wallace_cska32_fa126_or0[0]), .b(s_wallace_cska32_and_14_4[0]), .cin(s_wallace_cska32_and_13_5[0]), .fa_xor1(s_wallace_cska32_fa127_xor1), .fa_or0(s_wallace_cska32_fa127_or0));
  and_gate and_gate_s_wallace_cska32_and_15_4(.a(a[15]), .b(b[4]), .out(s_wallace_cska32_and_15_4));
  and_gate and_gate_s_wallace_cska32_and_14_5(.a(a[14]), .b(b[5]), .out(s_wallace_cska32_and_14_5));
  fa fa_s_wallace_cska32_fa128_out(.a(s_wallace_cska32_fa127_or0[0]), .b(s_wallace_cska32_and_15_4[0]), .cin(s_wallace_cska32_and_14_5[0]), .fa_xor1(s_wallace_cska32_fa128_xor1), .fa_or0(s_wallace_cska32_fa128_or0));
  and_gate and_gate_s_wallace_cska32_and_16_4(.a(a[16]), .b(b[4]), .out(s_wallace_cska32_and_16_4));
  and_gate and_gate_s_wallace_cska32_and_15_5(.a(a[15]), .b(b[5]), .out(s_wallace_cska32_and_15_5));
  fa fa_s_wallace_cska32_fa129_out(.a(s_wallace_cska32_fa128_or0[0]), .b(s_wallace_cska32_and_16_4[0]), .cin(s_wallace_cska32_and_15_5[0]), .fa_xor1(s_wallace_cska32_fa129_xor1), .fa_or0(s_wallace_cska32_fa129_or0));
  and_gate and_gate_s_wallace_cska32_and_17_4(.a(a[17]), .b(b[4]), .out(s_wallace_cska32_and_17_4));
  and_gate and_gate_s_wallace_cska32_and_16_5(.a(a[16]), .b(b[5]), .out(s_wallace_cska32_and_16_5));
  fa fa_s_wallace_cska32_fa130_out(.a(s_wallace_cska32_fa129_or0[0]), .b(s_wallace_cska32_and_17_4[0]), .cin(s_wallace_cska32_and_16_5[0]), .fa_xor1(s_wallace_cska32_fa130_xor1), .fa_or0(s_wallace_cska32_fa130_or0));
  and_gate and_gate_s_wallace_cska32_and_18_4(.a(a[18]), .b(b[4]), .out(s_wallace_cska32_and_18_4));
  and_gate and_gate_s_wallace_cska32_and_17_5(.a(a[17]), .b(b[5]), .out(s_wallace_cska32_and_17_5));
  fa fa_s_wallace_cska32_fa131_out(.a(s_wallace_cska32_fa130_or0[0]), .b(s_wallace_cska32_and_18_4[0]), .cin(s_wallace_cska32_and_17_5[0]), .fa_xor1(s_wallace_cska32_fa131_xor1), .fa_or0(s_wallace_cska32_fa131_or0));
  and_gate and_gate_s_wallace_cska32_and_19_4(.a(a[19]), .b(b[4]), .out(s_wallace_cska32_and_19_4));
  and_gate and_gate_s_wallace_cska32_and_18_5(.a(a[18]), .b(b[5]), .out(s_wallace_cska32_and_18_5));
  fa fa_s_wallace_cska32_fa132_out(.a(s_wallace_cska32_fa131_or0[0]), .b(s_wallace_cska32_and_19_4[0]), .cin(s_wallace_cska32_and_18_5[0]), .fa_xor1(s_wallace_cska32_fa132_xor1), .fa_or0(s_wallace_cska32_fa132_or0));
  and_gate and_gate_s_wallace_cska32_and_20_4(.a(a[20]), .b(b[4]), .out(s_wallace_cska32_and_20_4));
  and_gate and_gate_s_wallace_cska32_and_19_5(.a(a[19]), .b(b[5]), .out(s_wallace_cska32_and_19_5));
  fa fa_s_wallace_cska32_fa133_out(.a(s_wallace_cska32_fa132_or0[0]), .b(s_wallace_cska32_and_20_4[0]), .cin(s_wallace_cska32_and_19_5[0]), .fa_xor1(s_wallace_cska32_fa133_xor1), .fa_or0(s_wallace_cska32_fa133_or0));
  and_gate and_gate_s_wallace_cska32_and_21_4(.a(a[21]), .b(b[4]), .out(s_wallace_cska32_and_21_4));
  and_gate and_gate_s_wallace_cska32_and_20_5(.a(a[20]), .b(b[5]), .out(s_wallace_cska32_and_20_5));
  fa fa_s_wallace_cska32_fa134_out(.a(s_wallace_cska32_fa133_or0[0]), .b(s_wallace_cska32_and_21_4[0]), .cin(s_wallace_cska32_and_20_5[0]), .fa_xor1(s_wallace_cska32_fa134_xor1), .fa_or0(s_wallace_cska32_fa134_or0));
  and_gate and_gate_s_wallace_cska32_and_22_4(.a(a[22]), .b(b[4]), .out(s_wallace_cska32_and_22_4));
  and_gate and_gate_s_wallace_cska32_and_21_5(.a(a[21]), .b(b[5]), .out(s_wallace_cska32_and_21_5));
  fa fa_s_wallace_cska32_fa135_out(.a(s_wallace_cska32_fa134_or0[0]), .b(s_wallace_cska32_and_22_4[0]), .cin(s_wallace_cska32_and_21_5[0]), .fa_xor1(s_wallace_cska32_fa135_xor1), .fa_or0(s_wallace_cska32_fa135_or0));
  and_gate and_gate_s_wallace_cska32_and_23_4(.a(a[23]), .b(b[4]), .out(s_wallace_cska32_and_23_4));
  and_gate and_gate_s_wallace_cska32_and_22_5(.a(a[22]), .b(b[5]), .out(s_wallace_cska32_and_22_5));
  fa fa_s_wallace_cska32_fa136_out(.a(s_wallace_cska32_fa135_or0[0]), .b(s_wallace_cska32_and_23_4[0]), .cin(s_wallace_cska32_and_22_5[0]), .fa_xor1(s_wallace_cska32_fa136_xor1), .fa_or0(s_wallace_cska32_fa136_or0));
  and_gate and_gate_s_wallace_cska32_and_24_4(.a(a[24]), .b(b[4]), .out(s_wallace_cska32_and_24_4));
  and_gate and_gate_s_wallace_cska32_and_23_5(.a(a[23]), .b(b[5]), .out(s_wallace_cska32_and_23_5));
  fa fa_s_wallace_cska32_fa137_out(.a(s_wallace_cska32_fa136_or0[0]), .b(s_wallace_cska32_and_24_4[0]), .cin(s_wallace_cska32_and_23_5[0]), .fa_xor1(s_wallace_cska32_fa137_xor1), .fa_or0(s_wallace_cska32_fa137_or0));
  and_gate and_gate_s_wallace_cska32_and_25_4(.a(a[25]), .b(b[4]), .out(s_wallace_cska32_and_25_4));
  and_gate and_gate_s_wallace_cska32_and_24_5(.a(a[24]), .b(b[5]), .out(s_wallace_cska32_and_24_5));
  fa fa_s_wallace_cska32_fa138_out(.a(s_wallace_cska32_fa137_or0[0]), .b(s_wallace_cska32_and_25_4[0]), .cin(s_wallace_cska32_and_24_5[0]), .fa_xor1(s_wallace_cska32_fa138_xor1), .fa_or0(s_wallace_cska32_fa138_or0));
  and_gate and_gate_s_wallace_cska32_and_26_4(.a(a[26]), .b(b[4]), .out(s_wallace_cska32_and_26_4));
  and_gate and_gate_s_wallace_cska32_and_25_5(.a(a[25]), .b(b[5]), .out(s_wallace_cska32_and_25_5));
  fa fa_s_wallace_cska32_fa139_out(.a(s_wallace_cska32_fa138_or0[0]), .b(s_wallace_cska32_and_26_4[0]), .cin(s_wallace_cska32_and_25_5[0]), .fa_xor1(s_wallace_cska32_fa139_xor1), .fa_or0(s_wallace_cska32_fa139_or0));
  and_gate and_gate_s_wallace_cska32_and_27_4(.a(a[27]), .b(b[4]), .out(s_wallace_cska32_and_27_4));
  and_gate and_gate_s_wallace_cska32_and_26_5(.a(a[26]), .b(b[5]), .out(s_wallace_cska32_and_26_5));
  fa fa_s_wallace_cska32_fa140_out(.a(s_wallace_cska32_fa139_or0[0]), .b(s_wallace_cska32_and_27_4[0]), .cin(s_wallace_cska32_and_26_5[0]), .fa_xor1(s_wallace_cska32_fa140_xor1), .fa_or0(s_wallace_cska32_fa140_or0));
  and_gate and_gate_s_wallace_cska32_and_28_4(.a(a[28]), .b(b[4]), .out(s_wallace_cska32_and_28_4));
  and_gate and_gate_s_wallace_cska32_and_27_5(.a(a[27]), .b(b[5]), .out(s_wallace_cska32_and_27_5));
  fa fa_s_wallace_cska32_fa141_out(.a(s_wallace_cska32_fa140_or0[0]), .b(s_wallace_cska32_and_28_4[0]), .cin(s_wallace_cska32_and_27_5[0]), .fa_xor1(s_wallace_cska32_fa141_xor1), .fa_or0(s_wallace_cska32_fa141_or0));
  and_gate and_gate_s_wallace_cska32_and_27_6(.a(a[27]), .b(b[6]), .out(s_wallace_cska32_and_27_6));
  and_gate and_gate_s_wallace_cska32_and_26_7(.a(a[26]), .b(b[7]), .out(s_wallace_cska32_and_26_7));
  fa fa_s_wallace_cska32_fa142_out(.a(s_wallace_cska32_fa141_or0[0]), .b(s_wallace_cska32_and_27_6[0]), .cin(s_wallace_cska32_and_26_7[0]), .fa_xor1(s_wallace_cska32_fa142_xor1), .fa_or0(s_wallace_cska32_fa142_or0));
  and_gate and_gate_s_wallace_cska32_and_27_7(.a(a[27]), .b(b[7]), .out(s_wallace_cska32_and_27_7));
  and_gate and_gate_s_wallace_cska32_and_26_8(.a(a[26]), .b(b[8]), .out(s_wallace_cska32_and_26_8));
  fa fa_s_wallace_cska32_fa143_out(.a(s_wallace_cska32_fa142_or0[0]), .b(s_wallace_cska32_and_27_7[0]), .cin(s_wallace_cska32_and_26_8[0]), .fa_xor1(s_wallace_cska32_fa143_xor1), .fa_or0(s_wallace_cska32_fa143_or0));
  and_gate and_gate_s_wallace_cska32_and_27_8(.a(a[27]), .b(b[8]), .out(s_wallace_cska32_and_27_8));
  and_gate and_gate_s_wallace_cska32_and_26_9(.a(a[26]), .b(b[9]), .out(s_wallace_cska32_and_26_9));
  fa fa_s_wallace_cska32_fa144_out(.a(s_wallace_cska32_fa143_or0[0]), .b(s_wallace_cska32_and_27_8[0]), .cin(s_wallace_cska32_and_26_9[0]), .fa_xor1(s_wallace_cska32_fa144_xor1), .fa_or0(s_wallace_cska32_fa144_or0));
  and_gate and_gate_s_wallace_cska32_and_27_9(.a(a[27]), .b(b[9]), .out(s_wallace_cska32_and_27_9));
  and_gate and_gate_s_wallace_cska32_and_26_10(.a(a[26]), .b(b[10]), .out(s_wallace_cska32_and_26_10));
  fa fa_s_wallace_cska32_fa145_out(.a(s_wallace_cska32_fa144_or0[0]), .b(s_wallace_cska32_and_27_9[0]), .cin(s_wallace_cska32_and_26_10[0]), .fa_xor1(s_wallace_cska32_fa145_xor1), .fa_or0(s_wallace_cska32_fa145_or0));
  and_gate and_gate_s_wallace_cska32_and_27_10(.a(a[27]), .b(b[10]), .out(s_wallace_cska32_and_27_10));
  and_gate and_gate_s_wallace_cska32_and_26_11(.a(a[26]), .b(b[11]), .out(s_wallace_cska32_and_26_11));
  fa fa_s_wallace_cska32_fa146_out(.a(s_wallace_cska32_fa145_or0[0]), .b(s_wallace_cska32_and_27_10[0]), .cin(s_wallace_cska32_and_26_11[0]), .fa_xor1(s_wallace_cska32_fa146_xor1), .fa_or0(s_wallace_cska32_fa146_or0));
  and_gate and_gate_s_wallace_cska32_and_27_11(.a(a[27]), .b(b[11]), .out(s_wallace_cska32_and_27_11));
  and_gate and_gate_s_wallace_cska32_and_26_12(.a(a[26]), .b(b[12]), .out(s_wallace_cska32_and_26_12));
  fa fa_s_wallace_cska32_fa147_out(.a(s_wallace_cska32_fa146_or0[0]), .b(s_wallace_cska32_and_27_11[0]), .cin(s_wallace_cska32_and_26_12[0]), .fa_xor1(s_wallace_cska32_fa147_xor1), .fa_or0(s_wallace_cska32_fa147_or0));
  and_gate and_gate_s_wallace_cska32_and_27_12(.a(a[27]), .b(b[12]), .out(s_wallace_cska32_and_27_12));
  and_gate and_gate_s_wallace_cska32_and_26_13(.a(a[26]), .b(b[13]), .out(s_wallace_cska32_and_26_13));
  fa fa_s_wallace_cska32_fa148_out(.a(s_wallace_cska32_fa147_or0[0]), .b(s_wallace_cska32_and_27_12[0]), .cin(s_wallace_cska32_and_26_13[0]), .fa_xor1(s_wallace_cska32_fa148_xor1), .fa_or0(s_wallace_cska32_fa148_or0));
  and_gate and_gate_s_wallace_cska32_and_27_13(.a(a[27]), .b(b[13]), .out(s_wallace_cska32_and_27_13));
  and_gate and_gate_s_wallace_cska32_and_26_14(.a(a[26]), .b(b[14]), .out(s_wallace_cska32_and_26_14));
  fa fa_s_wallace_cska32_fa149_out(.a(s_wallace_cska32_fa148_or0[0]), .b(s_wallace_cska32_and_27_13[0]), .cin(s_wallace_cska32_and_26_14[0]), .fa_xor1(s_wallace_cska32_fa149_xor1), .fa_or0(s_wallace_cska32_fa149_or0));
  and_gate and_gate_s_wallace_cska32_and_27_14(.a(a[27]), .b(b[14]), .out(s_wallace_cska32_and_27_14));
  and_gate and_gate_s_wallace_cska32_and_26_15(.a(a[26]), .b(b[15]), .out(s_wallace_cska32_and_26_15));
  fa fa_s_wallace_cska32_fa150_out(.a(s_wallace_cska32_fa149_or0[0]), .b(s_wallace_cska32_and_27_14[0]), .cin(s_wallace_cska32_and_26_15[0]), .fa_xor1(s_wallace_cska32_fa150_xor1), .fa_or0(s_wallace_cska32_fa150_or0));
  and_gate and_gate_s_wallace_cska32_and_27_15(.a(a[27]), .b(b[15]), .out(s_wallace_cska32_and_27_15));
  and_gate and_gate_s_wallace_cska32_and_26_16(.a(a[26]), .b(b[16]), .out(s_wallace_cska32_and_26_16));
  fa fa_s_wallace_cska32_fa151_out(.a(s_wallace_cska32_fa150_or0[0]), .b(s_wallace_cska32_and_27_15[0]), .cin(s_wallace_cska32_and_26_16[0]), .fa_xor1(s_wallace_cska32_fa151_xor1), .fa_or0(s_wallace_cska32_fa151_or0));
  and_gate and_gate_s_wallace_cska32_and_27_16(.a(a[27]), .b(b[16]), .out(s_wallace_cska32_and_27_16));
  and_gate and_gate_s_wallace_cska32_and_26_17(.a(a[26]), .b(b[17]), .out(s_wallace_cska32_and_26_17));
  fa fa_s_wallace_cska32_fa152_out(.a(s_wallace_cska32_fa151_or0[0]), .b(s_wallace_cska32_and_27_16[0]), .cin(s_wallace_cska32_and_26_17[0]), .fa_xor1(s_wallace_cska32_fa152_xor1), .fa_or0(s_wallace_cska32_fa152_or0));
  and_gate and_gate_s_wallace_cska32_and_27_17(.a(a[27]), .b(b[17]), .out(s_wallace_cska32_and_27_17));
  and_gate and_gate_s_wallace_cska32_and_26_18(.a(a[26]), .b(b[18]), .out(s_wallace_cska32_and_26_18));
  fa fa_s_wallace_cska32_fa153_out(.a(s_wallace_cska32_fa152_or0[0]), .b(s_wallace_cska32_and_27_17[0]), .cin(s_wallace_cska32_and_26_18[0]), .fa_xor1(s_wallace_cska32_fa153_xor1), .fa_or0(s_wallace_cska32_fa153_or0));
  and_gate and_gate_s_wallace_cska32_and_27_18(.a(a[27]), .b(b[18]), .out(s_wallace_cska32_and_27_18));
  and_gate and_gate_s_wallace_cska32_and_26_19(.a(a[26]), .b(b[19]), .out(s_wallace_cska32_and_26_19));
  fa fa_s_wallace_cska32_fa154_out(.a(s_wallace_cska32_fa153_or0[0]), .b(s_wallace_cska32_and_27_18[0]), .cin(s_wallace_cska32_and_26_19[0]), .fa_xor1(s_wallace_cska32_fa154_xor1), .fa_or0(s_wallace_cska32_fa154_or0));
  and_gate and_gate_s_wallace_cska32_and_27_19(.a(a[27]), .b(b[19]), .out(s_wallace_cska32_and_27_19));
  and_gate and_gate_s_wallace_cska32_and_26_20(.a(a[26]), .b(b[20]), .out(s_wallace_cska32_and_26_20));
  fa fa_s_wallace_cska32_fa155_out(.a(s_wallace_cska32_fa154_or0[0]), .b(s_wallace_cska32_and_27_19[0]), .cin(s_wallace_cska32_and_26_20[0]), .fa_xor1(s_wallace_cska32_fa155_xor1), .fa_or0(s_wallace_cska32_fa155_or0));
  and_gate and_gate_s_wallace_cska32_and_27_20(.a(a[27]), .b(b[20]), .out(s_wallace_cska32_and_27_20));
  and_gate and_gate_s_wallace_cska32_and_26_21(.a(a[26]), .b(b[21]), .out(s_wallace_cska32_and_26_21));
  fa fa_s_wallace_cska32_fa156_out(.a(s_wallace_cska32_fa155_or0[0]), .b(s_wallace_cska32_and_27_20[0]), .cin(s_wallace_cska32_and_26_21[0]), .fa_xor1(s_wallace_cska32_fa156_xor1), .fa_or0(s_wallace_cska32_fa156_or0));
  and_gate and_gate_s_wallace_cska32_and_27_21(.a(a[27]), .b(b[21]), .out(s_wallace_cska32_and_27_21));
  and_gate and_gate_s_wallace_cska32_and_26_22(.a(a[26]), .b(b[22]), .out(s_wallace_cska32_and_26_22));
  fa fa_s_wallace_cska32_fa157_out(.a(s_wallace_cska32_fa156_or0[0]), .b(s_wallace_cska32_and_27_21[0]), .cin(s_wallace_cska32_and_26_22[0]), .fa_xor1(s_wallace_cska32_fa157_xor1), .fa_or0(s_wallace_cska32_fa157_or0));
  and_gate and_gate_s_wallace_cska32_and_27_22(.a(a[27]), .b(b[22]), .out(s_wallace_cska32_and_27_22));
  and_gate and_gate_s_wallace_cska32_and_26_23(.a(a[26]), .b(b[23]), .out(s_wallace_cska32_and_26_23));
  fa fa_s_wallace_cska32_fa158_out(.a(s_wallace_cska32_fa157_or0[0]), .b(s_wallace_cska32_and_27_22[0]), .cin(s_wallace_cska32_and_26_23[0]), .fa_xor1(s_wallace_cska32_fa158_xor1), .fa_or0(s_wallace_cska32_fa158_or0));
  and_gate and_gate_s_wallace_cska32_and_27_23(.a(a[27]), .b(b[23]), .out(s_wallace_cska32_and_27_23));
  and_gate and_gate_s_wallace_cska32_and_26_24(.a(a[26]), .b(b[24]), .out(s_wallace_cska32_and_26_24));
  fa fa_s_wallace_cska32_fa159_out(.a(s_wallace_cska32_fa158_or0[0]), .b(s_wallace_cska32_and_27_23[0]), .cin(s_wallace_cska32_and_26_24[0]), .fa_xor1(s_wallace_cska32_fa159_xor1), .fa_or0(s_wallace_cska32_fa159_or0));
  and_gate and_gate_s_wallace_cska32_and_27_24(.a(a[27]), .b(b[24]), .out(s_wallace_cska32_and_27_24));
  and_gate and_gate_s_wallace_cska32_and_26_25(.a(a[26]), .b(b[25]), .out(s_wallace_cska32_and_26_25));
  fa fa_s_wallace_cska32_fa160_out(.a(s_wallace_cska32_fa159_or0[0]), .b(s_wallace_cska32_and_27_24[0]), .cin(s_wallace_cska32_and_26_25[0]), .fa_xor1(s_wallace_cska32_fa160_xor1), .fa_or0(s_wallace_cska32_fa160_or0));
  and_gate and_gate_s_wallace_cska32_and_27_25(.a(a[27]), .b(b[25]), .out(s_wallace_cska32_and_27_25));
  and_gate and_gate_s_wallace_cska32_and_26_26(.a(a[26]), .b(b[26]), .out(s_wallace_cska32_and_26_26));
  fa fa_s_wallace_cska32_fa161_out(.a(s_wallace_cska32_fa160_or0[0]), .b(s_wallace_cska32_and_27_25[0]), .cin(s_wallace_cska32_and_26_26[0]), .fa_xor1(s_wallace_cska32_fa161_xor1), .fa_or0(s_wallace_cska32_fa161_or0));
  and_gate and_gate_s_wallace_cska32_and_27_26(.a(a[27]), .b(b[26]), .out(s_wallace_cska32_and_27_26));
  and_gate and_gate_s_wallace_cska32_and_26_27(.a(a[26]), .b(b[27]), .out(s_wallace_cska32_and_26_27));
  fa fa_s_wallace_cska32_fa162_out(.a(s_wallace_cska32_fa161_or0[0]), .b(s_wallace_cska32_and_27_26[0]), .cin(s_wallace_cska32_and_26_27[0]), .fa_xor1(s_wallace_cska32_fa162_xor1), .fa_or0(s_wallace_cska32_fa162_or0));
  and_gate and_gate_s_wallace_cska32_and_27_27(.a(a[27]), .b(b[27]), .out(s_wallace_cska32_and_27_27));
  and_gate and_gate_s_wallace_cska32_and_26_28(.a(a[26]), .b(b[28]), .out(s_wallace_cska32_and_26_28));
  fa fa_s_wallace_cska32_fa163_out(.a(s_wallace_cska32_fa162_or0[0]), .b(s_wallace_cska32_and_27_27[0]), .cin(s_wallace_cska32_and_26_28[0]), .fa_xor1(s_wallace_cska32_fa163_xor1), .fa_or0(s_wallace_cska32_fa163_or0));
  and_gate and_gate_s_wallace_cska32_and_27_28(.a(a[27]), .b(b[28]), .out(s_wallace_cska32_and_27_28));
  and_gate and_gate_s_wallace_cska32_and_26_29(.a(a[26]), .b(b[29]), .out(s_wallace_cska32_and_26_29));
  fa fa_s_wallace_cska32_fa164_out(.a(s_wallace_cska32_fa163_or0[0]), .b(s_wallace_cska32_and_27_28[0]), .cin(s_wallace_cska32_and_26_29[0]), .fa_xor1(s_wallace_cska32_fa164_xor1), .fa_or0(s_wallace_cska32_fa164_or0));
  and_gate and_gate_s_wallace_cska32_and_27_29(.a(a[27]), .b(b[29]), .out(s_wallace_cska32_and_27_29));
  and_gate and_gate_s_wallace_cska32_and_26_30(.a(a[26]), .b(b[30]), .out(s_wallace_cska32_and_26_30));
  fa fa_s_wallace_cska32_fa165_out(.a(s_wallace_cska32_fa164_or0[0]), .b(s_wallace_cska32_and_27_29[0]), .cin(s_wallace_cska32_and_26_30[0]), .fa_xor1(s_wallace_cska32_fa165_xor1), .fa_or0(s_wallace_cska32_fa165_or0));
  and_gate and_gate_s_wallace_cska32_and_27_30(.a(a[27]), .b(b[30]), .out(s_wallace_cska32_and_27_30));
  nand_gate nand_gate_s_wallace_cska32_nand_26_31(.a(a[26]), .b(b[31]), .out(s_wallace_cska32_nand_26_31));
  fa fa_s_wallace_cska32_fa166_out(.a(s_wallace_cska32_fa165_or0[0]), .b(s_wallace_cska32_and_27_30[0]), .cin(s_wallace_cska32_nand_26_31[0]), .fa_xor1(s_wallace_cska32_fa166_xor1), .fa_or0(s_wallace_cska32_fa166_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_27_31(.a(a[27]), .b(b[31]), .out(s_wallace_cska32_nand_27_31));
  fa fa_s_wallace_cska32_fa167_out(.a(s_wallace_cska32_fa166_or0[0]), .b(s_wallace_cska32_nand_27_31[0]), .cin(s_wallace_cska32_fa55_xor1[0]), .fa_xor1(s_wallace_cska32_fa167_xor1), .fa_or0(s_wallace_cska32_fa167_or0));
  ha ha_s_wallace_cska32_ha3_out(.a(s_wallace_cska32_fa2_xor1[0]), .b(s_wallace_cska32_fa59_xor1[0]), .ha_xor0(s_wallace_cska32_ha3_xor0), .ha_and0(s_wallace_cska32_ha3_and0));
  and_gate and_gate_s_wallace_cska32_and_0_6(.a(a[0]), .b(b[6]), .out(s_wallace_cska32_and_0_6));
  fa fa_s_wallace_cska32_fa168_out(.a(s_wallace_cska32_ha3_and0[0]), .b(s_wallace_cska32_and_0_6[0]), .cin(s_wallace_cska32_fa3_xor1[0]), .fa_xor1(s_wallace_cska32_fa168_xor1), .fa_or0(s_wallace_cska32_fa168_or0));
  and_gate and_gate_s_wallace_cska32_and_1_6(.a(a[1]), .b(b[6]), .out(s_wallace_cska32_and_1_6));
  and_gate and_gate_s_wallace_cska32_and_0_7(.a(a[0]), .b(b[7]), .out(s_wallace_cska32_and_0_7));
  fa fa_s_wallace_cska32_fa169_out(.a(s_wallace_cska32_fa168_or0[0]), .b(s_wallace_cska32_and_1_6[0]), .cin(s_wallace_cska32_and_0_7[0]), .fa_xor1(s_wallace_cska32_fa169_xor1), .fa_or0(s_wallace_cska32_fa169_or0));
  and_gate and_gate_s_wallace_cska32_and_2_6(.a(a[2]), .b(b[6]), .out(s_wallace_cska32_and_2_6));
  and_gate and_gate_s_wallace_cska32_and_1_7(.a(a[1]), .b(b[7]), .out(s_wallace_cska32_and_1_7));
  fa fa_s_wallace_cska32_fa170_out(.a(s_wallace_cska32_fa169_or0[0]), .b(s_wallace_cska32_and_2_6[0]), .cin(s_wallace_cska32_and_1_7[0]), .fa_xor1(s_wallace_cska32_fa170_xor1), .fa_or0(s_wallace_cska32_fa170_or0));
  and_gate and_gate_s_wallace_cska32_and_3_6(.a(a[3]), .b(b[6]), .out(s_wallace_cska32_and_3_6));
  and_gate and_gate_s_wallace_cska32_and_2_7(.a(a[2]), .b(b[7]), .out(s_wallace_cska32_and_2_7));
  fa fa_s_wallace_cska32_fa171_out(.a(s_wallace_cska32_fa170_or0[0]), .b(s_wallace_cska32_and_3_6[0]), .cin(s_wallace_cska32_and_2_7[0]), .fa_xor1(s_wallace_cska32_fa171_xor1), .fa_or0(s_wallace_cska32_fa171_or0));
  and_gate and_gate_s_wallace_cska32_and_4_6(.a(a[4]), .b(b[6]), .out(s_wallace_cska32_and_4_6));
  and_gate and_gate_s_wallace_cska32_and_3_7(.a(a[3]), .b(b[7]), .out(s_wallace_cska32_and_3_7));
  fa fa_s_wallace_cska32_fa172_out(.a(s_wallace_cska32_fa171_or0[0]), .b(s_wallace_cska32_and_4_6[0]), .cin(s_wallace_cska32_and_3_7[0]), .fa_xor1(s_wallace_cska32_fa172_xor1), .fa_or0(s_wallace_cska32_fa172_or0));
  and_gate and_gate_s_wallace_cska32_and_5_6(.a(a[5]), .b(b[6]), .out(s_wallace_cska32_and_5_6));
  and_gate and_gate_s_wallace_cska32_and_4_7(.a(a[4]), .b(b[7]), .out(s_wallace_cska32_and_4_7));
  fa fa_s_wallace_cska32_fa173_out(.a(s_wallace_cska32_fa172_or0[0]), .b(s_wallace_cska32_and_5_6[0]), .cin(s_wallace_cska32_and_4_7[0]), .fa_xor1(s_wallace_cska32_fa173_xor1), .fa_or0(s_wallace_cska32_fa173_or0));
  and_gate and_gate_s_wallace_cska32_and_6_6(.a(a[6]), .b(b[6]), .out(s_wallace_cska32_and_6_6));
  and_gate and_gate_s_wallace_cska32_and_5_7(.a(a[5]), .b(b[7]), .out(s_wallace_cska32_and_5_7));
  fa fa_s_wallace_cska32_fa174_out(.a(s_wallace_cska32_fa173_or0[0]), .b(s_wallace_cska32_and_6_6[0]), .cin(s_wallace_cska32_and_5_7[0]), .fa_xor1(s_wallace_cska32_fa174_xor1), .fa_or0(s_wallace_cska32_fa174_or0));
  and_gate and_gate_s_wallace_cska32_and_7_6(.a(a[7]), .b(b[6]), .out(s_wallace_cska32_and_7_6));
  and_gate and_gate_s_wallace_cska32_and_6_7(.a(a[6]), .b(b[7]), .out(s_wallace_cska32_and_6_7));
  fa fa_s_wallace_cska32_fa175_out(.a(s_wallace_cska32_fa174_or0[0]), .b(s_wallace_cska32_and_7_6[0]), .cin(s_wallace_cska32_and_6_7[0]), .fa_xor1(s_wallace_cska32_fa175_xor1), .fa_or0(s_wallace_cska32_fa175_or0));
  and_gate and_gate_s_wallace_cska32_and_8_6(.a(a[8]), .b(b[6]), .out(s_wallace_cska32_and_8_6));
  and_gate and_gate_s_wallace_cska32_and_7_7(.a(a[7]), .b(b[7]), .out(s_wallace_cska32_and_7_7));
  fa fa_s_wallace_cska32_fa176_out(.a(s_wallace_cska32_fa175_or0[0]), .b(s_wallace_cska32_and_8_6[0]), .cin(s_wallace_cska32_and_7_7[0]), .fa_xor1(s_wallace_cska32_fa176_xor1), .fa_or0(s_wallace_cska32_fa176_or0));
  and_gate and_gate_s_wallace_cska32_and_9_6(.a(a[9]), .b(b[6]), .out(s_wallace_cska32_and_9_6));
  and_gate and_gate_s_wallace_cska32_and_8_7(.a(a[8]), .b(b[7]), .out(s_wallace_cska32_and_8_7));
  fa fa_s_wallace_cska32_fa177_out(.a(s_wallace_cska32_fa176_or0[0]), .b(s_wallace_cska32_and_9_6[0]), .cin(s_wallace_cska32_and_8_7[0]), .fa_xor1(s_wallace_cska32_fa177_xor1), .fa_or0(s_wallace_cska32_fa177_or0));
  and_gate and_gate_s_wallace_cska32_and_10_6(.a(a[10]), .b(b[6]), .out(s_wallace_cska32_and_10_6));
  and_gate and_gate_s_wallace_cska32_and_9_7(.a(a[9]), .b(b[7]), .out(s_wallace_cska32_and_9_7));
  fa fa_s_wallace_cska32_fa178_out(.a(s_wallace_cska32_fa177_or0[0]), .b(s_wallace_cska32_and_10_6[0]), .cin(s_wallace_cska32_and_9_7[0]), .fa_xor1(s_wallace_cska32_fa178_xor1), .fa_or0(s_wallace_cska32_fa178_or0));
  and_gate and_gate_s_wallace_cska32_and_11_6(.a(a[11]), .b(b[6]), .out(s_wallace_cska32_and_11_6));
  and_gate and_gate_s_wallace_cska32_and_10_7(.a(a[10]), .b(b[7]), .out(s_wallace_cska32_and_10_7));
  fa fa_s_wallace_cska32_fa179_out(.a(s_wallace_cska32_fa178_or0[0]), .b(s_wallace_cska32_and_11_6[0]), .cin(s_wallace_cska32_and_10_7[0]), .fa_xor1(s_wallace_cska32_fa179_xor1), .fa_or0(s_wallace_cska32_fa179_or0));
  and_gate and_gate_s_wallace_cska32_and_12_6(.a(a[12]), .b(b[6]), .out(s_wallace_cska32_and_12_6));
  and_gate and_gate_s_wallace_cska32_and_11_7(.a(a[11]), .b(b[7]), .out(s_wallace_cska32_and_11_7));
  fa fa_s_wallace_cska32_fa180_out(.a(s_wallace_cska32_fa179_or0[0]), .b(s_wallace_cska32_and_12_6[0]), .cin(s_wallace_cska32_and_11_7[0]), .fa_xor1(s_wallace_cska32_fa180_xor1), .fa_or0(s_wallace_cska32_fa180_or0));
  and_gate and_gate_s_wallace_cska32_and_13_6(.a(a[13]), .b(b[6]), .out(s_wallace_cska32_and_13_6));
  and_gate and_gate_s_wallace_cska32_and_12_7(.a(a[12]), .b(b[7]), .out(s_wallace_cska32_and_12_7));
  fa fa_s_wallace_cska32_fa181_out(.a(s_wallace_cska32_fa180_or0[0]), .b(s_wallace_cska32_and_13_6[0]), .cin(s_wallace_cska32_and_12_7[0]), .fa_xor1(s_wallace_cska32_fa181_xor1), .fa_or0(s_wallace_cska32_fa181_or0));
  and_gate and_gate_s_wallace_cska32_and_14_6(.a(a[14]), .b(b[6]), .out(s_wallace_cska32_and_14_6));
  and_gate and_gate_s_wallace_cska32_and_13_7(.a(a[13]), .b(b[7]), .out(s_wallace_cska32_and_13_7));
  fa fa_s_wallace_cska32_fa182_out(.a(s_wallace_cska32_fa181_or0[0]), .b(s_wallace_cska32_and_14_6[0]), .cin(s_wallace_cska32_and_13_7[0]), .fa_xor1(s_wallace_cska32_fa182_xor1), .fa_or0(s_wallace_cska32_fa182_or0));
  and_gate and_gate_s_wallace_cska32_and_15_6(.a(a[15]), .b(b[6]), .out(s_wallace_cska32_and_15_6));
  and_gate and_gate_s_wallace_cska32_and_14_7(.a(a[14]), .b(b[7]), .out(s_wallace_cska32_and_14_7));
  fa fa_s_wallace_cska32_fa183_out(.a(s_wallace_cska32_fa182_or0[0]), .b(s_wallace_cska32_and_15_6[0]), .cin(s_wallace_cska32_and_14_7[0]), .fa_xor1(s_wallace_cska32_fa183_xor1), .fa_or0(s_wallace_cska32_fa183_or0));
  and_gate and_gate_s_wallace_cska32_and_16_6(.a(a[16]), .b(b[6]), .out(s_wallace_cska32_and_16_6));
  and_gate and_gate_s_wallace_cska32_and_15_7(.a(a[15]), .b(b[7]), .out(s_wallace_cska32_and_15_7));
  fa fa_s_wallace_cska32_fa184_out(.a(s_wallace_cska32_fa183_or0[0]), .b(s_wallace_cska32_and_16_6[0]), .cin(s_wallace_cska32_and_15_7[0]), .fa_xor1(s_wallace_cska32_fa184_xor1), .fa_or0(s_wallace_cska32_fa184_or0));
  and_gate and_gate_s_wallace_cska32_and_17_6(.a(a[17]), .b(b[6]), .out(s_wallace_cska32_and_17_6));
  and_gate and_gate_s_wallace_cska32_and_16_7(.a(a[16]), .b(b[7]), .out(s_wallace_cska32_and_16_7));
  fa fa_s_wallace_cska32_fa185_out(.a(s_wallace_cska32_fa184_or0[0]), .b(s_wallace_cska32_and_17_6[0]), .cin(s_wallace_cska32_and_16_7[0]), .fa_xor1(s_wallace_cska32_fa185_xor1), .fa_or0(s_wallace_cska32_fa185_or0));
  and_gate and_gate_s_wallace_cska32_and_18_6(.a(a[18]), .b(b[6]), .out(s_wallace_cska32_and_18_6));
  and_gate and_gate_s_wallace_cska32_and_17_7(.a(a[17]), .b(b[7]), .out(s_wallace_cska32_and_17_7));
  fa fa_s_wallace_cska32_fa186_out(.a(s_wallace_cska32_fa185_or0[0]), .b(s_wallace_cska32_and_18_6[0]), .cin(s_wallace_cska32_and_17_7[0]), .fa_xor1(s_wallace_cska32_fa186_xor1), .fa_or0(s_wallace_cska32_fa186_or0));
  and_gate and_gate_s_wallace_cska32_and_19_6(.a(a[19]), .b(b[6]), .out(s_wallace_cska32_and_19_6));
  and_gate and_gate_s_wallace_cska32_and_18_7(.a(a[18]), .b(b[7]), .out(s_wallace_cska32_and_18_7));
  fa fa_s_wallace_cska32_fa187_out(.a(s_wallace_cska32_fa186_or0[0]), .b(s_wallace_cska32_and_19_6[0]), .cin(s_wallace_cska32_and_18_7[0]), .fa_xor1(s_wallace_cska32_fa187_xor1), .fa_or0(s_wallace_cska32_fa187_or0));
  and_gate and_gate_s_wallace_cska32_and_20_6(.a(a[20]), .b(b[6]), .out(s_wallace_cska32_and_20_6));
  and_gate and_gate_s_wallace_cska32_and_19_7(.a(a[19]), .b(b[7]), .out(s_wallace_cska32_and_19_7));
  fa fa_s_wallace_cska32_fa188_out(.a(s_wallace_cska32_fa187_or0[0]), .b(s_wallace_cska32_and_20_6[0]), .cin(s_wallace_cska32_and_19_7[0]), .fa_xor1(s_wallace_cska32_fa188_xor1), .fa_or0(s_wallace_cska32_fa188_or0));
  and_gate and_gate_s_wallace_cska32_and_21_6(.a(a[21]), .b(b[6]), .out(s_wallace_cska32_and_21_6));
  and_gate and_gate_s_wallace_cska32_and_20_7(.a(a[20]), .b(b[7]), .out(s_wallace_cska32_and_20_7));
  fa fa_s_wallace_cska32_fa189_out(.a(s_wallace_cska32_fa188_or0[0]), .b(s_wallace_cska32_and_21_6[0]), .cin(s_wallace_cska32_and_20_7[0]), .fa_xor1(s_wallace_cska32_fa189_xor1), .fa_or0(s_wallace_cska32_fa189_or0));
  and_gate and_gate_s_wallace_cska32_and_22_6(.a(a[22]), .b(b[6]), .out(s_wallace_cska32_and_22_6));
  and_gate and_gate_s_wallace_cska32_and_21_7(.a(a[21]), .b(b[7]), .out(s_wallace_cska32_and_21_7));
  fa fa_s_wallace_cska32_fa190_out(.a(s_wallace_cska32_fa189_or0[0]), .b(s_wallace_cska32_and_22_6[0]), .cin(s_wallace_cska32_and_21_7[0]), .fa_xor1(s_wallace_cska32_fa190_xor1), .fa_or0(s_wallace_cska32_fa190_or0));
  and_gate and_gate_s_wallace_cska32_and_23_6(.a(a[23]), .b(b[6]), .out(s_wallace_cska32_and_23_6));
  and_gate and_gate_s_wallace_cska32_and_22_7(.a(a[22]), .b(b[7]), .out(s_wallace_cska32_and_22_7));
  fa fa_s_wallace_cska32_fa191_out(.a(s_wallace_cska32_fa190_or0[0]), .b(s_wallace_cska32_and_23_6[0]), .cin(s_wallace_cska32_and_22_7[0]), .fa_xor1(s_wallace_cska32_fa191_xor1), .fa_or0(s_wallace_cska32_fa191_or0));
  and_gate and_gate_s_wallace_cska32_and_24_6(.a(a[24]), .b(b[6]), .out(s_wallace_cska32_and_24_6));
  and_gate and_gate_s_wallace_cska32_and_23_7(.a(a[23]), .b(b[7]), .out(s_wallace_cska32_and_23_7));
  fa fa_s_wallace_cska32_fa192_out(.a(s_wallace_cska32_fa191_or0[0]), .b(s_wallace_cska32_and_24_6[0]), .cin(s_wallace_cska32_and_23_7[0]), .fa_xor1(s_wallace_cska32_fa192_xor1), .fa_or0(s_wallace_cska32_fa192_or0));
  and_gate and_gate_s_wallace_cska32_and_25_6(.a(a[25]), .b(b[6]), .out(s_wallace_cska32_and_25_6));
  and_gate and_gate_s_wallace_cska32_and_24_7(.a(a[24]), .b(b[7]), .out(s_wallace_cska32_and_24_7));
  fa fa_s_wallace_cska32_fa193_out(.a(s_wallace_cska32_fa192_or0[0]), .b(s_wallace_cska32_and_25_6[0]), .cin(s_wallace_cska32_and_24_7[0]), .fa_xor1(s_wallace_cska32_fa193_xor1), .fa_or0(s_wallace_cska32_fa193_or0));
  and_gate and_gate_s_wallace_cska32_and_26_6(.a(a[26]), .b(b[6]), .out(s_wallace_cska32_and_26_6));
  and_gate and_gate_s_wallace_cska32_and_25_7(.a(a[25]), .b(b[7]), .out(s_wallace_cska32_and_25_7));
  fa fa_s_wallace_cska32_fa194_out(.a(s_wallace_cska32_fa193_or0[0]), .b(s_wallace_cska32_and_26_6[0]), .cin(s_wallace_cska32_and_25_7[0]), .fa_xor1(s_wallace_cska32_fa194_xor1), .fa_or0(s_wallace_cska32_fa194_or0));
  and_gate and_gate_s_wallace_cska32_and_25_8(.a(a[25]), .b(b[8]), .out(s_wallace_cska32_and_25_8));
  and_gate and_gate_s_wallace_cska32_and_24_9(.a(a[24]), .b(b[9]), .out(s_wallace_cska32_and_24_9));
  fa fa_s_wallace_cska32_fa195_out(.a(s_wallace_cska32_fa194_or0[0]), .b(s_wallace_cska32_and_25_8[0]), .cin(s_wallace_cska32_and_24_9[0]), .fa_xor1(s_wallace_cska32_fa195_xor1), .fa_or0(s_wallace_cska32_fa195_or0));
  and_gate and_gate_s_wallace_cska32_and_25_9(.a(a[25]), .b(b[9]), .out(s_wallace_cska32_and_25_9));
  and_gate and_gate_s_wallace_cska32_and_24_10(.a(a[24]), .b(b[10]), .out(s_wallace_cska32_and_24_10));
  fa fa_s_wallace_cska32_fa196_out(.a(s_wallace_cska32_fa195_or0[0]), .b(s_wallace_cska32_and_25_9[0]), .cin(s_wallace_cska32_and_24_10[0]), .fa_xor1(s_wallace_cska32_fa196_xor1), .fa_or0(s_wallace_cska32_fa196_or0));
  and_gate and_gate_s_wallace_cska32_and_25_10(.a(a[25]), .b(b[10]), .out(s_wallace_cska32_and_25_10));
  and_gate and_gate_s_wallace_cska32_and_24_11(.a(a[24]), .b(b[11]), .out(s_wallace_cska32_and_24_11));
  fa fa_s_wallace_cska32_fa197_out(.a(s_wallace_cska32_fa196_or0[0]), .b(s_wallace_cska32_and_25_10[0]), .cin(s_wallace_cska32_and_24_11[0]), .fa_xor1(s_wallace_cska32_fa197_xor1), .fa_or0(s_wallace_cska32_fa197_or0));
  and_gate and_gate_s_wallace_cska32_and_25_11(.a(a[25]), .b(b[11]), .out(s_wallace_cska32_and_25_11));
  and_gate and_gate_s_wallace_cska32_and_24_12(.a(a[24]), .b(b[12]), .out(s_wallace_cska32_and_24_12));
  fa fa_s_wallace_cska32_fa198_out(.a(s_wallace_cska32_fa197_or0[0]), .b(s_wallace_cska32_and_25_11[0]), .cin(s_wallace_cska32_and_24_12[0]), .fa_xor1(s_wallace_cska32_fa198_xor1), .fa_or0(s_wallace_cska32_fa198_or0));
  and_gate and_gate_s_wallace_cska32_and_25_12(.a(a[25]), .b(b[12]), .out(s_wallace_cska32_and_25_12));
  and_gate and_gate_s_wallace_cska32_and_24_13(.a(a[24]), .b(b[13]), .out(s_wallace_cska32_and_24_13));
  fa fa_s_wallace_cska32_fa199_out(.a(s_wallace_cska32_fa198_or0[0]), .b(s_wallace_cska32_and_25_12[0]), .cin(s_wallace_cska32_and_24_13[0]), .fa_xor1(s_wallace_cska32_fa199_xor1), .fa_or0(s_wallace_cska32_fa199_or0));
  and_gate and_gate_s_wallace_cska32_and_25_13(.a(a[25]), .b(b[13]), .out(s_wallace_cska32_and_25_13));
  and_gate and_gate_s_wallace_cska32_and_24_14(.a(a[24]), .b(b[14]), .out(s_wallace_cska32_and_24_14));
  fa fa_s_wallace_cska32_fa200_out(.a(s_wallace_cska32_fa199_or0[0]), .b(s_wallace_cska32_and_25_13[0]), .cin(s_wallace_cska32_and_24_14[0]), .fa_xor1(s_wallace_cska32_fa200_xor1), .fa_or0(s_wallace_cska32_fa200_or0));
  and_gate and_gate_s_wallace_cska32_and_25_14(.a(a[25]), .b(b[14]), .out(s_wallace_cska32_and_25_14));
  and_gate and_gate_s_wallace_cska32_and_24_15(.a(a[24]), .b(b[15]), .out(s_wallace_cska32_and_24_15));
  fa fa_s_wallace_cska32_fa201_out(.a(s_wallace_cska32_fa200_or0[0]), .b(s_wallace_cska32_and_25_14[0]), .cin(s_wallace_cska32_and_24_15[0]), .fa_xor1(s_wallace_cska32_fa201_xor1), .fa_or0(s_wallace_cska32_fa201_or0));
  and_gate and_gate_s_wallace_cska32_and_25_15(.a(a[25]), .b(b[15]), .out(s_wallace_cska32_and_25_15));
  and_gate and_gate_s_wallace_cska32_and_24_16(.a(a[24]), .b(b[16]), .out(s_wallace_cska32_and_24_16));
  fa fa_s_wallace_cska32_fa202_out(.a(s_wallace_cska32_fa201_or0[0]), .b(s_wallace_cska32_and_25_15[0]), .cin(s_wallace_cska32_and_24_16[0]), .fa_xor1(s_wallace_cska32_fa202_xor1), .fa_or0(s_wallace_cska32_fa202_or0));
  and_gate and_gate_s_wallace_cska32_and_25_16(.a(a[25]), .b(b[16]), .out(s_wallace_cska32_and_25_16));
  and_gate and_gate_s_wallace_cska32_and_24_17(.a(a[24]), .b(b[17]), .out(s_wallace_cska32_and_24_17));
  fa fa_s_wallace_cska32_fa203_out(.a(s_wallace_cska32_fa202_or0[0]), .b(s_wallace_cska32_and_25_16[0]), .cin(s_wallace_cska32_and_24_17[0]), .fa_xor1(s_wallace_cska32_fa203_xor1), .fa_or0(s_wallace_cska32_fa203_or0));
  and_gate and_gate_s_wallace_cska32_and_25_17(.a(a[25]), .b(b[17]), .out(s_wallace_cska32_and_25_17));
  and_gate and_gate_s_wallace_cska32_and_24_18(.a(a[24]), .b(b[18]), .out(s_wallace_cska32_and_24_18));
  fa fa_s_wallace_cska32_fa204_out(.a(s_wallace_cska32_fa203_or0[0]), .b(s_wallace_cska32_and_25_17[0]), .cin(s_wallace_cska32_and_24_18[0]), .fa_xor1(s_wallace_cska32_fa204_xor1), .fa_or0(s_wallace_cska32_fa204_or0));
  and_gate and_gate_s_wallace_cska32_and_25_18(.a(a[25]), .b(b[18]), .out(s_wallace_cska32_and_25_18));
  and_gate and_gate_s_wallace_cska32_and_24_19(.a(a[24]), .b(b[19]), .out(s_wallace_cska32_and_24_19));
  fa fa_s_wallace_cska32_fa205_out(.a(s_wallace_cska32_fa204_or0[0]), .b(s_wallace_cska32_and_25_18[0]), .cin(s_wallace_cska32_and_24_19[0]), .fa_xor1(s_wallace_cska32_fa205_xor1), .fa_or0(s_wallace_cska32_fa205_or0));
  and_gate and_gate_s_wallace_cska32_and_25_19(.a(a[25]), .b(b[19]), .out(s_wallace_cska32_and_25_19));
  and_gate and_gate_s_wallace_cska32_and_24_20(.a(a[24]), .b(b[20]), .out(s_wallace_cska32_and_24_20));
  fa fa_s_wallace_cska32_fa206_out(.a(s_wallace_cska32_fa205_or0[0]), .b(s_wallace_cska32_and_25_19[0]), .cin(s_wallace_cska32_and_24_20[0]), .fa_xor1(s_wallace_cska32_fa206_xor1), .fa_or0(s_wallace_cska32_fa206_or0));
  and_gate and_gate_s_wallace_cska32_and_25_20(.a(a[25]), .b(b[20]), .out(s_wallace_cska32_and_25_20));
  and_gate and_gate_s_wallace_cska32_and_24_21(.a(a[24]), .b(b[21]), .out(s_wallace_cska32_and_24_21));
  fa fa_s_wallace_cska32_fa207_out(.a(s_wallace_cska32_fa206_or0[0]), .b(s_wallace_cska32_and_25_20[0]), .cin(s_wallace_cska32_and_24_21[0]), .fa_xor1(s_wallace_cska32_fa207_xor1), .fa_or0(s_wallace_cska32_fa207_or0));
  and_gate and_gate_s_wallace_cska32_and_25_21(.a(a[25]), .b(b[21]), .out(s_wallace_cska32_and_25_21));
  and_gate and_gate_s_wallace_cska32_and_24_22(.a(a[24]), .b(b[22]), .out(s_wallace_cska32_and_24_22));
  fa fa_s_wallace_cska32_fa208_out(.a(s_wallace_cska32_fa207_or0[0]), .b(s_wallace_cska32_and_25_21[0]), .cin(s_wallace_cska32_and_24_22[0]), .fa_xor1(s_wallace_cska32_fa208_xor1), .fa_or0(s_wallace_cska32_fa208_or0));
  and_gate and_gate_s_wallace_cska32_and_25_22(.a(a[25]), .b(b[22]), .out(s_wallace_cska32_and_25_22));
  and_gate and_gate_s_wallace_cska32_and_24_23(.a(a[24]), .b(b[23]), .out(s_wallace_cska32_and_24_23));
  fa fa_s_wallace_cska32_fa209_out(.a(s_wallace_cska32_fa208_or0[0]), .b(s_wallace_cska32_and_25_22[0]), .cin(s_wallace_cska32_and_24_23[0]), .fa_xor1(s_wallace_cska32_fa209_xor1), .fa_or0(s_wallace_cska32_fa209_or0));
  and_gate and_gate_s_wallace_cska32_and_25_23(.a(a[25]), .b(b[23]), .out(s_wallace_cska32_and_25_23));
  and_gate and_gate_s_wallace_cska32_and_24_24(.a(a[24]), .b(b[24]), .out(s_wallace_cska32_and_24_24));
  fa fa_s_wallace_cska32_fa210_out(.a(s_wallace_cska32_fa209_or0[0]), .b(s_wallace_cska32_and_25_23[0]), .cin(s_wallace_cska32_and_24_24[0]), .fa_xor1(s_wallace_cska32_fa210_xor1), .fa_or0(s_wallace_cska32_fa210_or0));
  and_gate and_gate_s_wallace_cska32_and_25_24(.a(a[25]), .b(b[24]), .out(s_wallace_cska32_and_25_24));
  and_gate and_gate_s_wallace_cska32_and_24_25(.a(a[24]), .b(b[25]), .out(s_wallace_cska32_and_24_25));
  fa fa_s_wallace_cska32_fa211_out(.a(s_wallace_cska32_fa210_or0[0]), .b(s_wallace_cska32_and_25_24[0]), .cin(s_wallace_cska32_and_24_25[0]), .fa_xor1(s_wallace_cska32_fa211_xor1), .fa_or0(s_wallace_cska32_fa211_or0));
  and_gate and_gate_s_wallace_cska32_and_25_25(.a(a[25]), .b(b[25]), .out(s_wallace_cska32_and_25_25));
  and_gate and_gate_s_wallace_cska32_and_24_26(.a(a[24]), .b(b[26]), .out(s_wallace_cska32_and_24_26));
  fa fa_s_wallace_cska32_fa212_out(.a(s_wallace_cska32_fa211_or0[0]), .b(s_wallace_cska32_and_25_25[0]), .cin(s_wallace_cska32_and_24_26[0]), .fa_xor1(s_wallace_cska32_fa212_xor1), .fa_or0(s_wallace_cska32_fa212_or0));
  and_gate and_gate_s_wallace_cska32_and_25_26(.a(a[25]), .b(b[26]), .out(s_wallace_cska32_and_25_26));
  and_gate and_gate_s_wallace_cska32_and_24_27(.a(a[24]), .b(b[27]), .out(s_wallace_cska32_and_24_27));
  fa fa_s_wallace_cska32_fa213_out(.a(s_wallace_cska32_fa212_or0[0]), .b(s_wallace_cska32_and_25_26[0]), .cin(s_wallace_cska32_and_24_27[0]), .fa_xor1(s_wallace_cska32_fa213_xor1), .fa_or0(s_wallace_cska32_fa213_or0));
  and_gate and_gate_s_wallace_cska32_and_25_27(.a(a[25]), .b(b[27]), .out(s_wallace_cska32_and_25_27));
  and_gate and_gate_s_wallace_cska32_and_24_28(.a(a[24]), .b(b[28]), .out(s_wallace_cska32_and_24_28));
  fa fa_s_wallace_cska32_fa214_out(.a(s_wallace_cska32_fa213_or0[0]), .b(s_wallace_cska32_and_25_27[0]), .cin(s_wallace_cska32_and_24_28[0]), .fa_xor1(s_wallace_cska32_fa214_xor1), .fa_or0(s_wallace_cska32_fa214_or0));
  and_gate and_gate_s_wallace_cska32_and_25_28(.a(a[25]), .b(b[28]), .out(s_wallace_cska32_and_25_28));
  and_gate and_gate_s_wallace_cska32_and_24_29(.a(a[24]), .b(b[29]), .out(s_wallace_cska32_and_24_29));
  fa fa_s_wallace_cska32_fa215_out(.a(s_wallace_cska32_fa214_or0[0]), .b(s_wallace_cska32_and_25_28[0]), .cin(s_wallace_cska32_and_24_29[0]), .fa_xor1(s_wallace_cska32_fa215_xor1), .fa_or0(s_wallace_cska32_fa215_or0));
  and_gate and_gate_s_wallace_cska32_and_25_29(.a(a[25]), .b(b[29]), .out(s_wallace_cska32_and_25_29));
  and_gate and_gate_s_wallace_cska32_and_24_30(.a(a[24]), .b(b[30]), .out(s_wallace_cska32_and_24_30));
  fa fa_s_wallace_cska32_fa216_out(.a(s_wallace_cska32_fa215_or0[0]), .b(s_wallace_cska32_and_25_29[0]), .cin(s_wallace_cska32_and_24_30[0]), .fa_xor1(s_wallace_cska32_fa216_xor1), .fa_or0(s_wallace_cska32_fa216_or0));
  and_gate and_gate_s_wallace_cska32_and_25_30(.a(a[25]), .b(b[30]), .out(s_wallace_cska32_and_25_30));
  nand_gate nand_gate_s_wallace_cska32_nand_24_31(.a(a[24]), .b(b[31]), .out(s_wallace_cska32_nand_24_31));
  fa fa_s_wallace_cska32_fa217_out(.a(s_wallace_cska32_fa216_or0[0]), .b(s_wallace_cska32_and_25_30[0]), .cin(s_wallace_cska32_nand_24_31[0]), .fa_xor1(s_wallace_cska32_fa217_xor1), .fa_or0(s_wallace_cska32_fa217_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_25_31(.a(a[25]), .b(b[31]), .out(s_wallace_cska32_nand_25_31));
  fa fa_s_wallace_cska32_fa218_out(.a(s_wallace_cska32_fa217_or0[0]), .b(s_wallace_cska32_nand_25_31[0]), .cin(s_wallace_cska32_fa53_xor1[0]), .fa_xor1(s_wallace_cska32_fa218_xor1), .fa_or0(s_wallace_cska32_fa218_or0));
  fa fa_s_wallace_cska32_fa219_out(.a(s_wallace_cska32_fa218_or0[0]), .b(s_wallace_cska32_fa54_xor1[0]), .cin(s_wallace_cska32_fa111_xor1[0]), .fa_xor1(s_wallace_cska32_fa219_xor1), .fa_or0(s_wallace_cska32_fa219_or0));
  ha ha_s_wallace_cska32_ha4_out(.a(s_wallace_cska32_fa60_xor1[0]), .b(s_wallace_cska32_fa115_xor1[0]), .ha_xor0(s_wallace_cska32_ha4_xor0), .ha_and0(s_wallace_cska32_ha4_and0));
  fa fa_s_wallace_cska32_fa220_out(.a(s_wallace_cska32_ha4_and0[0]), .b(s_wallace_cska32_fa4_xor1[0]), .cin(s_wallace_cska32_fa61_xor1[0]), .fa_xor1(s_wallace_cska32_fa220_xor1), .fa_or0(s_wallace_cska32_fa220_or0));
  and_gate and_gate_s_wallace_cska32_and_0_8(.a(a[0]), .b(b[8]), .out(s_wallace_cska32_and_0_8));
  fa fa_s_wallace_cska32_fa221_out(.a(s_wallace_cska32_fa220_or0[0]), .b(s_wallace_cska32_and_0_8[0]), .cin(s_wallace_cska32_fa5_xor1[0]), .fa_xor1(s_wallace_cska32_fa221_xor1), .fa_or0(s_wallace_cska32_fa221_or0));
  and_gate and_gate_s_wallace_cska32_and_1_8(.a(a[1]), .b(b[8]), .out(s_wallace_cska32_and_1_8));
  and_gate and_gate_s_wallace_cska32_and_0_9(.a(a[0]), .b(b[9]), .out(s_wallace_cska32_and_0_9));
  fa fa_s_wallace_cska32_fa222_out(.a(s_wallace_cska32_fa221_or0[0]), .b(s_wallace_cska32_and_1_8[0]), .cin(s_wallace_cska32_and_0_9[0]), .fa_xor1(s_wallace_cska32_fa222_xor1), .fa_or0(s_wallace_cska32_fa222_or0));
  and_gate and_gate_s_wallace_cska32_and_2_8(.a(a[2]), .b(b[8]), .out(s_wallace_cska32_and_2_8));
  and_gate and_gate_s_wallace_cska32_and_1_9(.a(a[1]), .b(b[9]), .out(s_wallace_cska32_and_1_9));
  fa fa_s_wallace_cska32_fa223_out(.a(s_wallace_cska32_fa222_or0[0]), .b(s_wallace_cska32_and_2_8[0]), .cin(s_wallace_cska32_and_1_9[0]), .fa_xor1(s_wallace_cska32_fa223_xor1), .fa_or0(s_wallace_cska32_fa223_or0));
  and_gate and_gate_s_wallace_cska32_and_3_8(.a(a[3]), .b(b[8]), .out(s_wallace_cska32_and_3_8));
  and_gate and_gate_s_wallace_cska32_and_2_9(.a(a[2]), .b(b[9]), .out(s_wallace_cska32_and_2_9));
  fa fa_s_wallace_cska32_fa224_out(.a(s_wallace_cska32_fa223_or0[0]), .b(s_wallace_cska32_and_3_8[0]), .cin(s_wallace_cska32_and_2_9[0]), .fa_xor1(s_wallace_cska32_fa224_xor1), .fa_or0(s_wallace_cska32_fa224_or0));
  and_gate and_gate_s_wallace_cska32_and_4_8(.a(a[4]), .b(b[8]), .out(s_wallace_cska32_and_4_8));
  and_gate and_gate_s_wallace_cska32_and_3_9(.a(a[3]), .b(b[9]), .out(s_wallace_cska32_and_3_9));
  fa fa_s_wallace_cska32_fa225_out(.a(s_wallace_cska32_fa224_or0[0]), .b(s_wallace_cska32_and_4_8[0]), .cin(s_wallace_cska32_and_3_9[0]), .fa_xor1(s_wallace_cska32_fa225_xor1), .fa_or0(s_wallace_cska32_fa225_or0));
  and_gate and_gate_s_wallace_cska32_and_5_8(.a(a[5]), .b(b[8]), .out(s_wallace_cska32_and_5_8));
  and_gate and_gate_s_wallace_cska32_and_4_9(.a(a[4]), .b(b[9]), .out(s_wallace_cska32_and_4_9));
  fa fa_s_wallace_cska32_fa226_out(.a(s_wallace_cska32_fa225_or0[0]), .b(s_wallace_cska32_and_5_8[0]), .cin(s_wallace_cska32_and_4_9[0]), .fa_xor1(s_wallace_cska32_fa226_xor1), .fa_or0(s_wallace_cska32_fa226_or0));
  and_gate and_gate_s_wallace_cska32_and_6_8(.a(a[6]), .b(b[8]), .out(s_wallace_cska32_and_6_8));
  and_gate and_gate_s_wallace_cska32_and_5_9(.a(a[5]), .b(b[9]), .out(s_wallace_cska32_and_5_9));
  fa fa_s_wallace_cska32_fa227_out(.a(s_wallace_cska32_fa226_or0[0]), .b(s_wallace_cska32_and_6_8[0]), .cin(s_wallace_cska32_and_5_9[0]), .fa_xor1(s_wallace_cska32_fa227_xor1), .fa_or0(s_wallace_cska32_fa227_or0));
  and_gate and_gate_s_wallace_cska32_and_7_8(.a(a[7]), .b(b[8]), .out(s_wallace_cska32_and_7_8));
  and_gate and_gate_s_wallace_cska32_and_6_9(.a(a[6]), .b(b[9]), .out(s_wallace_cska32_and_6_9));
  fa fa_s_wallace_cska32_fa228_out(.a(s_wallace_cska32_fa227_or0[0]), .b(s_wallace_cska32_and_7_8[0]), .cin(s_wallace_cska32_and_6_9[0]), .fa_xor1(s_wallace_cska32_fa228_xor1), .fa_or0(s_wallace_cska32_fa228_or0));
  and_gate and_gate_s_wallace_cska32_and_8_8(.a(a[8]), .b(b[8]), .out(s_wallace_cska32_and_8_8));
  and_gate and_gate_s_wallace_cska32_and_7_9(.a(a[7]), .b(b[9]), .out(s_wallace_cska32_and_7_9));
  fa fa_s_wallace_cska32_fa229_out(.a(s_wallace_cska32_fa228_or0[0]), .b(s_wallace_cska32_and_8_8[0]), .cin(s_wallace_cska32_and_7_9[0]), .fa_xor1(s_wallace_cska32_fa229_xor1), .fa_or0(s_wallace_cska32_fa229_or0));
  and_gate and_gate_s_wallace_cska32_and_9_8(.a(a[9]), .b(b[8]), .out(s_wallace_cska32_and_9_8));
  and_gate and_gate_s_wallace_cska32_and_8_9(.a(a[8]), .b(b[9]), .out(s_wallace_cska32_and_8_9));
  fa fa_s_wallace_cska32_fa230_out(.a(s_wallace_cska32_fa229_or0[0]), .b(s_wallace_cska32_and_9_8[0]), .cin(s_wallace_cska32_and_8_9[0]), .fa_xor1(s_wallace_cska32_fa230_xor1), .fa_or0(s_wallace_cska32_fa230_or0));
  and_gate and_gate_s_wallace_cska32_and_10_8(.a(a[10]), .b(b[8]), .out(s_wallace_cska32_and_10_8));
  and_gate and_gate_s_wallace_cska32_and_9_9(.a(a[9]), .b(b[9]), .out(s_wallace_cska32_and_9_9));
  fa fa_s_wallace_cska32_fa231_out(.a(s_wallace_cska32_fa230_or0[0]), .b(s_wallace_cska32_and_10_8[0]), .cin(s_wallace_cska32_and_9_9[0]), .fa_xor1(s_wallace_cska32_fa231_xor1), .fa_or0(s_wallace_cska32_fa231_or0));
  and_gate and_gate_s_wallace_cska32_and_11_8(.a(a[11]), .b(b[8]), .out(s_wallace_cska32_and_11_8));
  and_gate and_gate_s_wallace_cska32_and_10_9(.a(a[10]), .b(b[9]), .out(s_wallace_cska32_and_10_9));
  fa fa_s_wallace_cska32_fa232_out(.a(s_wallace_cska32_fa231_or0[0]), .b(s_wallace_cska32_and_11_8[0]), .cin(s_wallace_cska32_and_10_9[0]), .fa_xor1(s_wallace_cska32_fa232_xor1), .fa_or0(s_wallace_cska32_fa232_or0));
  and_gate and_gate_s_wallace_cska32_and_12_8(.a(a[12]), .b(b[8]), .out(s_wallace_cska32_and_12_8));
  and_gate and_gate_s_wallace_cska32_and_11_9(.a(a[11]), .b(b[9]), .out(s_wallace_cska32_and_11_9));
  fa fa_s_wallace_cska32_fa233_out(.a(s_wallace_cska32_fa232_or0[0]), .b(s_wallace_cska32_and_12_8[0]), .cin(s_wallace_cska32_and_11_9[0]), .fa_xor1(s_wallace_cska32_fa233_xor1), .fa_or0(s_wallace_cska32_fa233_or0));
  and_gate and_gate_s_wallace_cska32_and_13_8(.a(a[13]), .b(b[8]), .out(s_wallace_cska32_and_13_8));
  and_gate and_gate_s_wallace_cska32_and_12_9(.a(a[12]), .b(b[9]), .out(s_wallace_cska32_and_12_9));
  fa fa_s_wallace_cska32_fa234_out(.a(s_wallace_cska32_fa233_or0[0]), .b(s_wallace_cska32_and_13_8[0]), .cin(s_wallace_cska32_and_12_9[0]), .fa_xor1(s_wallace_cska32_fa234_xor1), .fa_or0(s_wallace_cska32_fa234_or0));
  and_gate and_gate_s_wallace_cska32_and_14_8(.a(a[14]), .b(b[8]), .out(s_wallace_cska32_and_14_8));
  and_gate and_gate_s_wallace_cska32_and_13_9(.a(a[13]), .b(b[9]), .out(s_wallace_cska32_and_13_9));
  fa fa_s_wallace_cska32_fa235_out(.a(s_wallace_cska32_fa234_or0[0]), .b(s_wallace_cska32_and_14_8[0]), .cin(s_wallace_cska32_and_13_9[0]), .fa_xor1(s_wallace_cska32_fa235_xor1), .fa_or0(s_wallace_cska32_fa235_or0));
  and_gate and_gate_s_wallace_cska32_and_15_8(.a(a[15]), .b(b[8]), .out(s_wallace_cska32_and_15_8));
  and_gate and_gate_s_wallace_cska32_and_14_9(.a(a[14]), .b(b[9]), .out(s_wallace_cska32_and_14_9));
  fa fa_s_wallace_cska32_fa236_out(.a(s_wallace_cska32_fa235_or0[0]), .b(s_wallace_cska32_and_15_8[0]), .cin(s_wallace_cska32_and_14_9[0]), .fa_xor1(s_wallace_cska32_fa236_xor1), .fa_or0(s_wallace_cska32_fa236_or0));
  and_gate and_gate_s_wallace_cska32_and_16_8(.a(a[16]), .b(b[8]), .out(s_wallace_cska32_and_16_8));
  and_gate and_gate_s_wallace_cska32_and_15_9(.a(a[15]), .b(b[9]), .out(s_wallace_cska32_and_15_9));
  fa fa_s_wallace_cska32_fa237_out(.a(s_wallace_cska32_fa236_or0[0]), .b(s_wallace_cska32_and_16_8[0]), .cin(s_wallace_cska32_and_15_9[0]), .fa_xor1(s_wallace_cska32_fa237_xor1), .fa_or0(s_wallace_cska32_fa237_or0));
  and_gate and_gate_s_wallace_cska32_and_17_8(.a(a[17]), .b(b[8]), .out(s_wallace_cska32_and_17_8));
  and_gate and_gate_s_wallace_cska32_and_16_9(.a(a[16]), .b(b[9]), .out(s_wallace_cska32_and_16_9));
  fa fa_s_wallace_cska32_fa238_out(.a(s_wallace_cska32_fa237_or0[0]), .b(s_wallace_cska32_and_17_8[0]), .cin(s_wallace_cska32_and_16_9[0]), .fa_xor1(s_wallace_cska32_fa238_xor1), .fa_or0(s_wallace_cska32_fa238_or0));
  and_gate and_gate_s_wallace_cska32_and_18_8(.a(a[18]), .b(b[8]), .out(s_wallace_cska32_and_18_8));
  and_gate and_gate_s_wallace_cska32_and_17_9(.a(a[17]), .b(b[9]), .out(s_wallace_cska32_and_17_9));
  fa fa_s_wallace_cska32_fa239_out(.a(s_wallace_cska32_fa238_or0[0]), .b(s_wallace_cska32_and_18_8[0]), .cin(s_wallace_cska32_and_17_9[0]), .fa_xor1(s_wallace_cska32_fa239_xor1), .fa_or0(s_wallace_cska32_fa239_or0));
  and_gate and_gate_s_wallace_cska32_and_19_8(.a(a[19]), .b(b[8]), .out(s_wallace_cska32_and_19_8));
  and_gate and_gate_s_wallace_cska32_and_18_9(.a(a[18]), .b(b[9]), .out(s_wallace_cska32_and_18_9));
  fa fa_s_wallace_cska32_fa240_out(.a(s_wallace_cska32_fa239_or0[0]), .b(s_wallace_cska32_and_19_8[0]), .cin(s_wallace_cska32_and_18_9[0]), .fa_xor1(s_wallace_cska32_fa240_xor1), .fa_or0(s_wallace_cska32_fa240_or0));
  and_gate and_gate_s_wallace_cska32_and_20_8(.a(a[20]), .b(b[8]), .out(s_wallace_cska32_and_20_8));
  and_gate and_gate_s_wallace_cska32_and_19_9(.a(a[19]), .b(b[9]), .out(s_wallace_cska32_and_19_9));
  fa fa_s_wallace_cska32_fa241_out(.a(s_wallace_cska32_fa240_or0[0]), .b(s_wallace_cska32_and_20_8[0]), .cin(s_wallace_cska32_and_19_9[0]), .fa_xor1(s_wallace_cska32_fa241_xor1), .fa_or0(s_wallace_cska32_fa241_or0));
  and_gate and_gate_s_wallace_cska32_and_21_8(.a(a[21]), .b(b[8]), .out(s_wallace_cska32_and_21_8));
  and_gate and_gate_s_wallace_cska32_and_20_9(.a(a[20]), .b(b[9]), .out(s_wallace_cska32_and_20_9));
  fa fa_s_wallace_cska32_fa242_out(.a(s_wallace_cska32_fa241_or0[0]), .b(s_wallace_cska32_and_21_8[0]), .cin(s_wallace_cska32_and_20_9[0]), .fa_xor1(s_wallace_cska32_fa242_xor1), .fa_or0(s_wallace_cska32_fa242_or0));
  and_gate and_gate_s_wallace_cska32_and_22_8(.a(a[22]), .b(b[8]), .out(s_wallace_cska32_and_22_8));
  and_gate and_gate_s_wallace_cska32_and_21_9(.a(a[21]), .b(b[9]), .out(s_wallace_cska32_and_21_9));
  fa fa_s_wallace_cska32_fa243_out(.a(s_wallace_cska32_fa242_or0[0]), .b(s_wallace_cska32_and_22_8[0]), .cin(s_wallace_cska32_and_21_9[0]), .fa_xor1(s_wallace_cska32_fa243_xor1), .fa_or0(s_wallace_cska32_fa243_or0));
  and_gate and_gate_s_wallace_cska32_and_23_8(.a(a[23]), .b(b[8]), .out(s_wallace_cska32_and_23_8));
  and_gate and_gate_s_wallace_cska32_and_22_9(.a(a[22]), .b(b[9]), .out(s_wallace_cska32_and_22_9));
  fa fa_s_wallace_cska32_fa244_out(.a(s_wallace_cska32_fa243_or0[0]), .b(s_wallace_cska32_and_23_8[0]), .cin(s_wallace_cska32_and_22_9[0]), .fa_xor1(s_wallace_cska32_fa244_xor1), .fa_or0(s_wallace_cska32_fa244_or0));
  and_gate and_gate_s_wallace_cska32_and_24_8(.a(a[24]), .b(b[8]), .out(s_wallace_cska32_and_24_8));
  and_gate and_gate_s_wallace_cska32_and_23_9(.a(a[23]), .b(b[9]), .out(s_wallace_cska32_and_23_9));
  fa fa_s_wallace_cska32_fa245_out(.a(s_wallace_cska32_fa244_or0[0]), .b(s_wallace_cska32_and_24_8[0]), .cin(s_wallace_cska32_and_23_9[0]), .fa_xor1(s_wallace_cska32_fa245_xor1), .fa_or0(s_wallace_cska32_fa245_or0));
  and_gate and_gate_s_wallace_cska32_and_23_10(.a(a[23]), .b(b[10]), .out(s_wallace_cska32_and_23_10));
  and_gate and_gate_s_wallace_cska32_and_22_11(.a(a[22]), .b(b[11]), .out(s_wallace_cska32_and_22_11));
  fa fa_s_wallace_cska32_fa246_out(.a(s_wallace_cska32_fa245_or0[0]), .b(s_wallace_cska32_and_23_10[0]), .cin(s_wallace_cska32_and_22_11[0]), .fa_xor1(s_wallace_cska32_fa246_xor1), .fa_or0(s_wallace_cska32_fa246_or0));
  and_gate and_gate_s_wallace_cska32_and_23_11(.a(a[23]), .b(b[11]), .out(s_wallace_cska32_and_23_11));
  and_gate and_gate_s_wallace_cska32_and_22_12(.a(a[22]), .b(b[12]), .out(s_wallace_cska32_and_22_12));
  fa fa_s_wallace_cska32_fa247_out(.a(s_wallace_cska32_fa246_or0[0]), .b(s_wallace_cska32_and_23_11[0]), .cin(s_wallace_cska32_and_22_12[0]), .fa_xor1(s_wallace_cska32_fa247_xor1), .fa_or0(s_wallace_cska32_fa247_or0));
  and_gate and_gate_s_wallace_cska32_and_23_12(.a(a[23]), .b(b[12]), .out(s_wallace_cska32_and_23_12));
  and_gate and_gate_s_wallace_cska32_and_22_13(.a(a[22]), .b(b[13]), .out(s_wallace_cska32_and_22_13));
  fa fa_s_wallace_cska32_fa248_out(.a(s_wallace_cska32_fa247_or0[0]), .b(s_wallace_cska32_and_23_12[0]), .cin(s_wallace_cska32_and_22_13[0]), .fa_xor1(s_wallace_cska32_fa248_xor1), .fa_or0(s_wallace_cska32_fa248_or0));
  and_gate and_gate_s_wallace_cska32_and_23_13(.a(a[23]), .b(b[13]), .out(s_wallace_cska32_and_23_13));
  and_gate and_gate_s_wallace_cska32_and_22_14(.a(a[22]), .b(b[14]), .out(s_wallace_cska32_and_22_14));
  fa fa_s_wallace_cska32_fa249_out(.a(s_wallace_cska32_fa248_or0[0]), .b(s_wallace_cska32_and_23_13[0]), .cin(s_wallace_cska32_and_22_14[0]), .fa_xor1(s_wallace_cska32_fa249_xor1), .fa_or0(s_wallace_cska32_fa249_or0));
  and_gate and_gate_s_wallace_cska32_and_23_14(.a(a[23]), .b(b[14]), .out(s_wallace_cska32_and_23_14));
  and_gate and_gate_s_wallace_cska32_and_22_15(.a(a[22]), .b(b[15]), .out(s_wallace_cska32_and_22_15));
  fa fa_s_wallace_cska32_fa250_out(.a(s_wallace_cska32_fa249_or0[0]), .b(s_wallace_cska32_and_23_14[0]), .cin(s_wallace_cska32_and_22_15[0]), .fa_xor1(s_wallace_cska32_fa250_xor1), .fa_or0(s_wallace_cska32_fa250_or0));
  and_gate and_gate_s_wallace_cska32_and_23_15(.a(a[23]), .b(b[15]), .out(s_wallace_cska32_and_23_15));
  and_gate and_gate_s_wallace_cska32_and_22_16(.a(a[22]), .b(b[16]), .out(s_wallace_cska32_and_22_16));
  fa fa_s_wallace_cska32_fa251_out(.a(s_wallace_cska32_fa250_or0[0]), .b(s_wallace_cska32_and_23_15[0]), .cin(s_wallace_cska32_and_22_16[0]), .fa_xor1(s_wallace_cska32_fa251_xor1), .fa_or0(s_wallace_cska32_fa251_or0));
  and_gate and_gate_s_wallace_cska32_and_23_16(.a(a[23]), .b(b[16]), .out(s_wallace_cska32_and_23_16));
  and_gate and_gate_s_wallace_cska32_and_22_17(.a(a[22]), .b(b[17]), .out(s_wallace_cska32_and_22_17));
  fa fa_s_wallace_cska32_fa252_out(.a(s_wallace_cska32_fa251_or0[0]), .b(s_wallace_cska32_and_23_16[0]), .cin(s_wallace_cska32_and_22_17[0]), .fa_xor1(s_wallace_cska32_fa252_xor1), .fa_or0(s_wallace_cska32_fa252_or0));
  and_gate and_gate_s_wallace_cska32_and_23_17(.a(a[23]), .b(b[17]), .out(s_wallace_cska32_and_23_17));
  and_gate and_gate_s_wallace_cska32_and_22_18(.a(a[22]), .b(b[18]), .out(s_wallace_cska32_and_22_18));
  fa fa_s_wallace_cska32_fa253_out(.a(s_wallace_cska32_fa252_or0[0]), .b(s_wallace_cska32_and_23_17[0]), .cin(s_wallace_cska32_and_22_18[0]), .fa_xor1(s_wallace_cska32_fa253_xor1), .fa_or0(s_wallace_cska32_fa253_or0));
  and_gate and_gate_s_wallace_cska32_and_23_18(.a(a[23]), .b(b[18]), .out(s_wallace_cska32_and_23_18));
  and_gate and_gate_s_wallace_cska32_and_22_19(.a(a[22]), .b(b[19]), .out(s_wallace_cska32_and_22_19));
  fa fa_s_wallace_cska32_fa254_out(.a(s_wallace_cska32_fa253_or0[0]), .b(s_wallace_cska32_and_23_18[0]), .cin(s_wallace_cska32_and_22_19[0]), .fa_xor1(s_wallace_cska32_fa254_xor1), .fa_or0(s_wallace_cska32_fa254_or0));
  and_gate and_gate_s_wallace_cska32_and_23_19(.a(a[23]), .b(b[19]), .out(s_wallace_cska32_and_23_19));
  and_gate and_gate_s_wallace_cska32_and_22_20(.a(a[22]), .b(b[20]), .out(s_wallace_cska32_and_22_20));
  fa fa_s_wallace_cska32_fa255_out(.a(s_wallace_cska32_fa254_or0[0]), .b(s_wallace_cska32_and_23_19[0]), .cin(s_wallace_cska32_and_22_20[0]), .fa_xor1(s_wallace_cska32_fa255_xor1), .fa_or0(s_wallace_cska32_fa255_or0));
  and_gate and_gate_s_wallace_cska32_and_23_20(.a(a[23]), .b(b[20]), .out(s_wallace_cska32_and_23_20));
  and_gate and_gate_s_wallace_cska32_and_22_21(.a(a[22]), .b(b[21]), .out(s_wallace_cska32_and_22_21));
  fa fa_s_wallace_cska32_fa256_out(.a(s_wallace_cska32_fa255_or0[0]), .b(s_wallace_cska32_and_23_20[0]), .cin(s_wallace_cska32_and_22_21[0]), .fa_xor1(s_wallace_cska32_fa256_xor1), .fa_or0(s_wallace_cska32_fa256_or0));
  and_gate and_gate_s_wallace_cska32_and_23_21(.a(a[23]), .b(b[21]), .out(s_wallace_cska32_and_23_21));
  and_gate and_gate_s_wallace_cska32_and_22_22(.a(a[22]), .b(b[22]), .out(s_wallace_cska32_and_22_22));
  fa fa_s_wallace_cska32_fa257_out(.a(s_wallace_cska32_fa256_or0[0]), .b(s_wallace_cska32_and_23_21[0]), .cin(s_wallace_cska32_and_22_22[0]), .fa_xor1(s_wallace_cska32_fa257_xor1), .fa_or0(s_wallace_cska32_fa257_or0));
  and_gate and_gate_s_wallace_cska32_and_23_22(.a(a[23]), .b(b[22]), .out(s_wallace_cska32_and_23_22));
  and_gate and_gate_s_wallace_cska32_and_22_23(.a(a[22]), .b(b[23]), .out(s_wallace_cska32_and_22_23));
  fa fa_s_wallace_cska32_fa258_out(.a(s_wallace_cska32_fa257_or0[0]), .b(s_wallace_cska32_and_23_22[0]), .cin(s_wallace_cska32_and_22_23[0]), .fa_xor1(s_wallace_cska32_fa258_xor1), .fa_or0(s_wallace_cska32_fa258_or0));
  and_gate and_gate_s_wallace_cska32_and_23_23(.a(a[23]), .b(b[23]), .out(s_wallace_cska32_and_23_23));
  and_gate and_gate_s_wallace_cska32_and_22_24(.a(a[22]), .b(b[24]), .out(s_wallace_cska32_and_22_24));
  fa fa_s_wallace_cska32_fa259_out(.a(s_wallace_cska32_fa258_or0[0]), .b(s_wallace_cska32_and_23_23[0]), .cin(s_wallace_cska32_and_22_24[0]), .fa_xor1(s_wallace_cska32_fa259_xor1), .fa_or0(s_wallace_cska32_fa259_or0));
  and_gate and_gate_s_wallace_cska32_and_23_24(.a(a[23]), .b(b[24]), .out(s_wallace_cska32_and_23_24));
  and_gate and_gate_s_wallace_cska32_and_22_25(.a(a[22]), .b(b[25]), .out(s_wallace_cska32_and_22_25));
  fa fa_s_wallace_cska32_fa260_out(.a(s_wallace_cska32_fa259_or0[0]), .b(s_wallace_cska32_and_23_24[0]), .cin(s_wallace_cska32_and_22_25[0]), .fa_xor1(s_wallace_cska32_fa260_xor1), .fa_or0(s_wallace_cska32_fa260_or0));
  and_gate and_gate_s_wallace_cska32_and_23_25(.a(a[23]), .b(b[25]), .out(s_wallace_cska32_and_23_25));
  and_gate and_gate_s_wallace_cska32_and_22_26(.a(a[22]), .b(b[26]), .out(s_wallace_cska32_and_22_26));
  fa fa_s_wallace_cska32_fa261_out(.a(s_wallace_cska32_fa260_or0[0]), .b(s_wallace_cska32_and_23_25[0]), .cin(s_wallace_cska32_and_22_26[0]), .fa_xor1(s_wallace_cska32_fa261_xor1), .fa_or0(s_wallace_cska32_fa261_or0));
  and_gate and_gate_s_wallace_cska32_and_23_26(.a(a[23]), .b(b[26]), .out(s_wallace_cska32_and_23_26));
  and_gate and_gate_s_wallace_cska32_and_22_27(.a(a[22]), .b(b[27]), .out(s_wallace_cska32_and_22_27));
  fa fa_s_wallace_cska32_fa262_out(.a(s_wallace_cska32_fa261_or0[0]), .b(s_wallace_cska32_and_23_26[0]), .cin(s_wallace_cska32_and_22_27[0]), .fa_xor1(s_wallace_cska32_fa262_xor1), .fa_or0(s_wallace_cska32_fa262_or0));
  and_gate and_gate_s_wallace_cska32_and_23_27(.a(a[23]), .b(b[27]), .out(s_wallace_cska32_and_23_27));
  and_gate and_gate_s_wallace_cska32_and_22_28(.a(a[22]), .b(b[28]), .out(s_wallace_cska32_and_22_28));
  fa fa_s_wallace_cska32_fa263_out(.a(s_wallace_cska32_fa262_or0[0]), .b(s_wallace_cska32_and_23_27[0]), .cin(s_wallace_cska32_and_22_28[0]), .fa_xor1(s_wallace_cska32_fa263_xor1), .fa_or0(s_wallace_cska32_fa263_or0));
  and_gate and_gate_s_wallace_cska32_and_23_28(.a(a[23]), .b(b[28]), .out(s_wallace_cska32_and_23_28));
  and_gate and_gate_s_wallace_cska32_and_22_29(.a(a[22]), .b(b[29]), .out(s_wallace_cska32_and_22_29));
  fa fa_s_wallace_cska32_fa264_out(.a(s_wallace_cska32_fa263_or0[0]), .b(s_wallace_cska32_and_23_28[0]), .cin(s_wallace_cska32_and_22_29[0]), .fa_xor1(s_wallace_cska32_fa264_xor1), .fa_or0(s_wallace_cska32_fa264_or0));
  and_gate and_gate_s_wallace_cska32_and_23_29(.a(a[23]), .b(b[29]), .out(s_wallace_cska32_and_23_29));
  and_gate and_gate_s_wallace_cska32_and_22_30(.a(a[22]), .b(b[30]), .out(s_wallace_cska32_and_22_30));
  fa fa_s_wallace_cska32_fa265_out(.a(s_wallace_cska32_fa264_or0[0]), .b(s_wallace_cska32_and_23_29[0]), .cin(s_wallace_cska32_and_22_30[0]), .fa_xor1(s_wallace_cska32_fa265_xor1), .fa_or0(s_wallace_cska32_fa265_or0));
  and_gate and_gate_s_wallace_cska32_and_23_30(.a(a[23]), .b(b[30]), .out(s_wallace_cska32_and_23_30));
  nand_gate nand_gate_s_wallace_cska32_nand_22_31(.a(a[22]), .b(b[31]), .out(s_wallace_cska32_nand_22_31));
  fa fa_s_wallace_cska32_fa266_out(.a(s_wallace_cska32_fa265_or0[0]), .b(s_wallace_cska32_and_23_30[0]), .cin(s_wallace_cska32_nand_22_31[0]), .fa_xor1(s_wallace_cska32_fa266_xor1), .fa_or0(s_wallace_cska32_fa266_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_23_31(.a(a[23]), .b(b[31]), .out(s_wallace_cska32_nand_23_31));
  fa fa_s_wallace_cska32_fa267_out(.a(s_wallace_cska32_fa266_or0[0]), .b(s_wallace_cska32_nand_23_31[0]), .cin(s_wallace_cska32_fa51_xor1[0]), .fa_xor1(s_wallace_cska32_fa267_xor1), .fa_or0(s_wallace_cska32_fa267_or0));
  fa fa_s_wallace_cska32_fa268_out(.a(s_wallace_cska32_fa267_or0[0]), .b(s_wallace_cska32_fa52_xor1[0]), .cin(s_wallace_cska32_fa109_xor1[0]), .fa_xor1(s_wallace_cska32_fa268_xor1), .fa_or0(s_wallace_cska32_fa268_or0));
  fa fa_s_wallace_cska32_fa269_out(.a(s_wallace_cska32_fa268_or0[0]), .b(s_wallace_cska32_fa110_xor1[0]), .cin(s_wallace_cska32_fa165_xor1[0]), .fa_xor1(s_wallace_cska32_fa269_xor1), .fa_or0(s_wallace_cska32_fa269_or0));
  ha ha_s_wallace_cska32_ha5_out(.a(s_wallace_cska32_fa116_xor1[0]), .b(s_wallace_cska32_fa169_xor1[0]), .ha_xor0(s_wallace_cska32_ha5_xor0), .ha_and0(s_wallace_cska32_ha5_and0));
  fa fa_s_wallace_cska32_fa270_out(.a(s_wallace_cska32_ha5_and0[0]), .b(s_wallace_cska32_fa62_xor1[0]), .cin(s_wallace_cska32_fa117_xor1[0]), .fa_xor1(s_wallace_cska32_fa270_xor1), .fa_or0(s_wallace_cska32_fa270_or0));
  fa fa_s_wallace_cska32_fa271_out(.a(s_wallace_cska32_fa270_or0[0]), .b(s_wallace_cska32_fa6_xor1[0]), .cin(s_wallace_cska32_fa63_xor1[0]), .fa_xor1(s_wallace_cska32_fa271_xor1), .fa_or0(s_wallace_cska32_fa271_or0));
  and_gate and_gate_s_wallace_cska32_and_0_10(.a(a[0]), .b(b[10]), .out(s_wallace_cska32_and_0_10));
  fa fa_s_wallace_cska32_fa272_out(.a(s_wallace_cska32_fa271_or0[0]), .b(s_wallace_cska32_and_0_10[0]), .cin(s_wallace_cska32_fa7_xor1[0]), .fa_xor1(s_wallace_cska32_fa272_xor1), .fa_or0(s_wallace_cska32_fa272_or0));
  and_gate and_gate_s_wallace_cska32_and_1_10(.a(a[1]), .b(b[10]), .out(s_wallace_cska32_and_1_10));
  and_gate and_gate_s_wallace_cska32_and_0_11(.a(a[0]), .b(b[11]), .out(s_wallace_cska32_and_0_11));
  fa fa_s_wallace_cska32_fa273_out(.a(s_wallace_cska32_fa272_or0[0]), .b(s_wallace_cska32_and_1_10[0]), .cin(s_wallace_cska32_and_0_11[0]), .fa_xor1(s_wallace_cska32_fa273_xor1), .fa_or0(s_wallace_cska32_fa273_or0));
  and_gate and_gate_s_wallace_cska32_and_2_10(.a(a[2]), .b(b[10]), .out(s_wallace_cska32_and_2_10));
  and_gate and_gate_s_wallace_cska32_and_1_11(.a(a[1]), .b(b[11]), .out(s_wallace_cska32_and_1_11));
  fa fa_s_wallace_cska32_fa274_out(.a(s_wallace_cska32_fa273_or0[0]), .b(s_wallace_cska32_and_2_10[0]), .cin(s_wallace_cska32_and_1_11[0]), .fa_xor1(s_wallace_cska32_fa274_xor1), .fa_or0(s_wallace_cska32_fa274_or0));
  and_gate and_gate_s_wallace_cska32_and_3_10(.a(a[3]), .b(b[10]), .out(s_wallace_cska32_and_3_10));
  and_gate and_gate_s_wallace_cska32_and_2_11(.a(a[2]), .b(b[11]), .out(s_wallace_cska32_and_2_11));
  fa fa_s_wallace_cska32_fa275_out(.a(s_wallace_cska32_fa274_or0[0]), .b(s_wallace_cska32_and_3_10[0]), .cin(s_wallace_cska32_and_2_11[0]), .fa_xor1(s_wallace_cska32_fa275_xor1), .fa_or0(s_wallace_cska32_fa275_or0));
  and_gate and_gate_s_wallace_cska32_and_4_10(.a(a[4]), .b(b[10]), .out(s_wallace_cska32_and_4_10));
  and_gate and_gate_s_wallace_cska32_and_3_11(.a(a[3]), .b(b[11]), .out(s_wallace_cska32_and_3_11));
  fa fa_s_wallace_cska32_fa276_out(.a(s_wallace_cska32_fa275_or0[0]), .b(s_wallace_cska32_and_4_10[0]), .cin(s_wallace_cska32_and_3_11[0]), .fa_xor1(s_wallace_cska32_fa276_xor1), .fa_or0(s_wallace_cska32_fa276_or0));
  and_gate and_gate_s_wallace_cska32_and_5_10(.a(a[5]), .b(b[10]), .out(s_wallace_cska32_and_5_10));
  and_gate and_gate_s_wallace_cska32_and_4_11(.a(a[4]), .b(b[11]), .out(s_wallace_cska32_and_4_11));
  fa fa_s_wallace_cska32_fa277_out(.a(s_wallace_cska32_fa276_or0[0]), .b(s_wallace_cska32_and_5_10[0]), .cin(s_wallace_cska32_and_4_11[0]), .fa_xor1(s_wallace_cska32_fa277_xor1), .fa_or0(s_wallace_cska32_fa277_or0));
  and_gate and_gate_s_wallace_cska32_and_6_10(.a(a[6]), .b(b[10]), .out(s_wallace_cska32_and_6_10));
  and_gate and_gate_s_wallace_cska32_and_5_11(.a(a[5]), .b(b[11]), .out(s_wallace_cska32_and_5_11));
  fa fa_s_wallace_cska32_fa278_out(.a(s_wallace_cska32_fa277_or0[0]), .b(s_wallace_cska32_and_6_10[0]), .cin(s_wallace_cska32_and_5_11[0]), .fa_xor1(s_wallace_cska32_fa278_xor1), .fa_or0(s_wallace_cska32_fa278_or0));
  and_gate and_gate_s_wallace_cska32_and_7_10(.a(a[7]), .b(b[10]), .out(s_wallace_cska32_and_7_10));
  and_gate and_gate_s_wallace_cska32_and_6_11(.a(a[6]), .b(b[11]), .out(s_wallace_cska32_and_6_11));
  fa fa_s_wallace_cska32_fa279_out(.a(s_wallace_cska32_fa278_or0[0]), .b(s_wallace_cska32_and_7_10[0]), .cin(s_wallace_cska32_and_6_11[0]), .fa_xor1(s_wallace_cska32_fa279_xor1), .fa_or0(s_wallace_cska32_fa279_or0));
  and_gate and_gate_s_wallace_cska32_and_8_10(.a(a[8]), .b(b[10]), .out(s_wallace_cska32_and_8_10));
  and_gate and_gate_s_wallace_cska32_and_7_11(.a(a[7]), .b(b[11]), .out(s_wallace_cska32_and_7_11));
  fa fa_s_wallace_cska32_fa280_out(.a(s_wallace_cska32_fa279_or0[0]), .b(s_wallace_cska32_and_8_10[0]), .cin(s_wallace_cska32_and_7_11[0]), .fa_xor1(s_wallace_cska32_fa280_xor1), .fa_or0(s_wallace_cska32_fa280_or0));
  and_gate and_gate_s_wallace_cska32_and_9_10(.a(a[9]), .b(b[10]), .out(s_wallace_cska32_and_9_10));
  and_gate and_gate_s_wallace_cska32_and_8_11(.a(a[8]), .b(b[11]), .out(s_wallace_cska32_and_8_11));
  fa fa_s_wallace_cska32_fa281_out(.a(s_wallace_cska32_fa280_or0[0]), .b(s_wallace_cska32_and_9_10[0]), .cin(s_wallace_cska32_and_8_11[0]), .fa_xor1(s_wallace_cska32_fa281_xor1), .fa_or0(s_wallace_cska32_fa281_or0));
  and_gate and_gate_s_wallace_cska32_and_10_10(.a(a[10]), .b(b[10]), .out(s_wallace_cska32_and_10_10));
  and_gate and_gate_s_wallace_cska32_and_9_11(.a(a[9]), .b(b[11]), .out(s_wallace_cska32_and_9_11));
  fa fa_s_wallace_cska32_fa282_out(.a(s_wallace_cska32_fa281_or0[0]), .b(s_wallace_cska32_and_10_10[0]), .cin(s_wallace_cska32_and_9_11[0]), .fa_xor1(s_wallace_cska32_fa282_xor1), .fa_or0(s_wallace_cska32_fa282_or0));
  and_gate and_gate_s_wallace_cska32_and_11_10(.a(a[11]), .b(b[10]), .out(s_wallace_cska32_and_11_10));
  and_gate and_gate_s_wallace_cska32_and_10_11(.a(a[10]), .b(b[11]), .out(s_wallace_cska32_and_10_11));
  fa fa_s_wallace_cska32_fa283_out(.a(s_wallace_cska32_fa282_or0[0]), .b(s_wallace_cska32_and_11_10[0]), .cin(s_wallace_cska32_and_10_11[0]), .fa_xor1(s_wallace_cska32_fa283_xor1), .fa_or0(s_wallace_cska32_fa283_or0));
  and_gate and_gate_s_wallace_cska32_and_12_10(.a(a[12]), .b(b[10]), .out(s_wallace_cska32_and_12_10));
  and_gate and_gate_s_wallace_cska32_and_11_11(.a(a[11]), .b(b[11]), .out(s_wallace_cska32_and_11_11));
  fa fa_s_wallace_cska32_fa284_out(.a(s_wallace_cska32_fa283_or0[0]), .b(s_wallace_cska32_and_12_10[0]), .cin(s_wallace_cska32_and_11_11[0]), .fa_xor1(s_wallace_cska32_fa284_xor1), .fa_or0(s_wallace_cska32_fa284_or0));
  and_gate and_gate_s_wallace_cska32_and_13_10(.a(a[13]), .b(b[10]), .out(s_wallace_cska32_and_13_10));
  and_gate and_gate_s_wallace_cska32_and_12_11(.a(a[12]), .b(b[11]), .out(s_wallace_cska32_and_12_11));
  fa fa_s_wallace_cska32_fa285_out(.a(s_wallace_cska32_fa284_or0[0]), .b(s_wallace_cska32_and_13_10[0]), .cin(s_wallace_cska32_and_12_11[0]), .fa_xor1(s_wallace_cska32_fa285_xor1), .fa_or0(s_wallace_cska32_fa285_or0));
  and_gate and_gate_s_wallace_cska32_and_14_10(.a(a[14]), .b(b[10]), .out(s_wallace_cska32_and_14_10));
  and_gate and_gate_s_wallace_cska32_and_13_11(.a(a[13]), .b(b[11]), .out(s_wallace_cska32_and_13_11));
  fa fa_s_wallace_cska32_fa286_out(.a(s_wallace_cska32_fa285_or0[0]), .b(s_wallace_cska32_and_14_10[0]), .cin(s_wallace_cska32_and_13_11[0]), .fa_xor1(s_wallace_cska32_fa286_xor1), .fa_or0(s_wallace_cska32_fa286_or0));
  and_gate and_gate_s_wallace_cska32_and_15_10(.a(a[15]), .b(b[10]), .out(s_wallace_cska32_and_15_10));
  and_gate and_gate_s_wallace_cska32_and_14_11(.a(a[14]), .b(b[11]), .out(s_wallace_cska32_and_14_11));
  fa fa_s_wallace_cska32_fa287_out(.a(s_wallace_cska32_fa286_or0[0]), .b(s_wallace_cska32_and_15_10[0]), .cin(s_wallace_cska32_and_14_11[0]), .fa_xor1(s_wallace_cska32_fa287_xor1), .fa_or0(s_wallace_cska32_fa287_or0));
  and_gate and_gate_s_wallace_cska32_and_16_10(.a(a[16]), .b(b[10]), .out(s_wallace_cska32_and_16_10));
  and_gate and_gate_s_wallace_cska32_and_15_11(.a(a[15]), .b(b[11]), .out(s_wallace_cska32_and_15_11));
  fa fa_s_wallace_cska32_fa288_out(.a(s_wallace_cska32_fa287_or0[0]), .b(s_wallace_cska32_and_16_10[0]), .cin(s_wallace_cska32_and_15_11[0]), .fa_xor1(s_wallace_cska32_fa288_xor1), .fa_or0(s_wallace_cska32_fa288_or0));
  and_gate and_gate_s_wallace_cska32_and_17_10(.a(a[17]), .b(b[10]), .out(s_wallace_cska32_and_17_10));
  and_gate and_gate_s_wallace_cska32_and_16_11(.a(a[16]), .b(b[11]), .out(s_wallace_cska32_and_16_11));
  fa fa_s_wallace_cska32_fa289_out(.a(s_wallace_cska32_fa288_or0[0]), .b(s_wallace_cska32_and_17_10[0]), .cin(s_wallace_cska32_and_16_11[0]), .fa_xor1(s_wallace_cska32_fa289_xor1), .fa_or0(s_wallace_cska32_fa289_or0));
  and_gate and_gate_s_wallace_cska32_and_18_10(.a(a[18]), .b(b[10]), .out(s_wallace_cska32_and_18_10));
  and_gate and_gate_s_wallace_cska32_and_17_11(.a(a[17]), .b(b[11]), .out(s_wallace_cska32_and_17_11));
  fa fa_s_wallace_cska32_fa290_out(.a(s_wallace_cska32_fa289_or0[0]), .b(s_wallace_cska32_and_18_10[0]), .cin(s_wallace_cska32_and_17_11[0]), .fa_xor1(s_wallace_cska32_fa290_xor1), .fa_or0(s_wallace_cska32_fa290_or0));
  and_gate and_gate_s_wallace_cska32_and_19_10(.a(a[19]), .b(b[10]), .out(s_wallace_cska32_and_19_10));
  and_gate and_gate_s_wallace_cska32_and_18_11(.a(a[18]), .b(b[11]), .out(s_wallace_cska32_and_18_11));
  fa fa_s_wallace_cska32_fa291_out(.a(s_wallace_cska32_fa290_or0[0]), .b(s_wallace_cska32_and_19_10[0]), .cin(s_wallace_cska32_and_18_11[0]), .fa_xor1(s_wallace_cska32_fa291_xor1), .fa_or0(s_wallace_cska32_fa291_or0));
  and_gate and_gate_s_wallace_cska32_and_20_10(.a(a[20]), .b(b[10]), .out(s_wallace_cska32_and_20_10));
  and_gate and_gate_s_wallace_cska32_and_19_11(.a(a[19]), .b(b[11]), .out(s_wallace_cska32_and_19_11));
  fa fa_s_wallace_cska32_fa292_out(.a(s_wallace_cska32_fa291_or0[0]), .b(s_wallace_cska32_and_20_10[0]), .cin(s_wallace_cska32_and_19_11[0]), .fa_xor1(s_wallace_cska32_fa292_xor1), .fa_or0(s_wallace_cska32_fa292_or0));
  and_gate and_gate_s_wallace_cska32_and_21_10(.a(a[21]), .b(b[10]), .out(s_wallace_cska32_and_21_10));
  and_gate and_gate_s_wallace_cska32_and_20_11(.a(a[20]), .b(b[11]), .out(s_wallace_cska32_and_20_11));
  fa fa_s_wallace_cska32_fa293_out(.a(s_wallace_cska32_fa292_or0[0]), .b(s_wallace_cska32_and_21_10[0]), .cin(s_wallace_cska32_and_20_11[0]), .fa_xor1(s_wallace_cska32_fa293_xor1), .fa_or0(s_wallace_cska32_fa293_or0));
  and_gate and_gate_s_wallace_cska32_and_22_10(.a(a[22]), .b(b[10]), .out(s_wallace_cska32_and_22_10));
  and_gate and_gate_s_wallace_cska32_and_21_11(.a(a[21]), .b(b[11]), .out(s_wallace_cska32_and_21_11));
  fa fa_s_wallace_cska32_fa294_out(.a(s_wallace_cska32_fa293_or0[0]), .b(s_wallace_cska32_and_22_10[0]), .cin(s_wallace_cska32_and_21_11[0]), .fa_xor1(s_wallace_cska32_fa294_xor1), .fa_or0(s_wallace_cska32_fa294_or0));
  and_gate and_gate_s_wallace_cska32_and_21_12(.a(a[21]), .b(b[12]), .out(s_wallace_cska32_and_21_12));
  and_gate and_gate_s_wallace_cska32_and_20_13(.a(a[20]), .b(b[13]), .out(s_wallace_cska32_and_20_13));
  fa fa_s_wallace_cska32_fa295_out(.a(s_wallace_cska32_fa294_or0[0]), .b(s_wallace_cska32_and_21_12[0]), .cin(s_wallace_cska32_and_20_13[0]), .fa_xor1(s_wallace_cska32_fa295_xor1), .fa_or0(s_wallace_cska32_fa295_or0));
  and_gate and_gate_s_wallace_cska32_and_21_13(.a(a[21]), .b(b[13]), .out(s_wallace_cska32_and_21_13));
  and_gate and_gate_s_wallace_cska32_and_20_14(.a(a[20]), .b(b[14]), .out(s_wallace_cska32_and_20_14));
  fa fa_s_wallace_cska32_fa296_out(.a(s_wallace_cska32_fa295_or0[0]), .b(s_wallace_cska32_and_21_13[0]), .cin(s_wallace_cska32_and_20_14[0]), .fa_xor1(s_wallace_cska32_fa296_xor1), .fa_or0(s_wallace_cska32_fa296_or0));
  and_gate and_gate_s_wallace_cska32_and_21_14(.a(a[21]), .b(b[14]), .out(s_wallace_cska32_and_21_14));
  and_gate and_gate_s_wallace_cska32_and_20_15(.a(a[20]), .b(b[15]), .out(s_wallace_cska32_and_20_15));
  fa fa_s_wallace_cska32_fa297_out(.a(s_wallace_cska32_fa296_or0[0]), .b(s_wallace_cska32_and_21_14[0]), .cin(s_wallace_cska32_and_20_15[0]), .fa_xor1(s_wallace_cska32_fa297_xor1), .fa_or0(s_wallace_cska32_fa297_or0));
  and_gate and_gate_s_wallace_cska32_and_21_15(.a(a[21]), .b(b[15]), .out(s_wallace_cska32_and_21_15));
  and_gate and_gate_s_wallace_cska32_and_20_16(.a(a[20]), .b(b[16]), .out(s_wallace_cska32_and_20_16));
  fa fa_s_wallace_cska32_fa298_out(.a(s_wallace_cska32_fa297_or0[0]), .b(s_wallace_cska32_and_21_15[0]), .cin(s_wallace_cska32_and_20_16[0]), .fa_xor1(s_wallace_cska32_fa298_xor1), .fa_or0(s_wallace_cska32_fa298_or0));
  and_gate and_gate_s_wallace_cska32_and_21_16(.a(a[21]), .b(b[16]), .out(s_wallace_cska32_and_21_16));
  and_gate and_gate_s_wallace_cska32_and_20_17(.a(a[20]), .b(b[17]), .out(s_wallace_cska32_and_20_17));
  fa fa_s_wallace_cska32_fa299_out(.a(s_wallace_cska32_fa298_or0[0]), .b(s_wallace_cska32_and_21_16[0]), .cin(s_wallace_cska32_and_20_17[0]), .fa_xor1(s_wallace_cska32_fa299_xor1), .fa_or0(s_wallace_cska32_fa299_or0));
  and_gate and_gate_s_wallace_cska32_and_21_17(.a(a[21]), .b(b[17]), .out(s_wallace_cska32_and_21_17));
  and_gate and_gate_s_wallace_cska32_and_20_18(.a(a[20]), .b(b[18]), .out(s_wallace_cska32_and_20_18));
  fa fa_s_wallace_cska32_fa300_out(.a(s_wallace_cska32_fa299_or0[0]), .b(s_wallace_cska32_and_21_17[0]), .cin(s_wallace_cska32_and_20_18[0]), .fa_xor1(s_wallace_cska32_fa300_xor1), .fa_or0(s_wallace_cska32_fa300_or0));
  and_gate and_gate_s_wallace_cska32_and_21_18(.a(a[21]), .b(b[18]), .out(s_wallace_cska32_and_21_18));
  and_gate and_gate_s_wallace_cska32_and_20_19(.a(a[20]), .b(b[19]), .out(s_wallace_cska32_and_20_19));
  fa fa_s_wallace_cska32_fa301_out(.a(s_wallace_cska32_fa300_or0[0]), .b(s_wallace_cska32_and_21_18[0]), .cin(s_wallace_cska32_and_20_19[0]), .fa_xor1(s_wallace_cska32_fa301_xor1), .fa_or0(s_wallace_cska32_fa301_or0));
  and_gate and_gate_s_wallace_cska32_and_21_19(.a(a[21]), .b(b[19]), .out(s_wallace_cska32_and_21_19));
  and_gate and_gate_s_wallace_cska32_and_20_20(.a(a[20]), .b(b[20]), .out(s_wallace_cska32_and_20_20));
  fa fa_s_wallace_cska32_fa302_out(.a(s_wallace_cska32_fa301_or0[0]), .b(s_wallace_cska32_and_21_19[0]), .cin(s_wallace_cska32_and_20_20[0]), .fa_xor1(s_wallace_cska32_fa302_xor1), .fa_or0(s_wallace_cska32_fa302_or0));
  and_gate and_gate_s_wallace_cska32_and_21_20(.a(a[21]), .b(b[20]), .out(s_wallace_cska32_and_21_20));
  and_gate and_gate_s_wallace_cska32_and_20_21(.a(a[20]), .b(b[21]), .out(s_wallace_cska32_and_20_21));
  fa fa_s_wallace_cska32_fa303_out(.a(s_wallace_cska32_fa302_or0[0]), .b(s_wallace_cska32_and_21_20[0]), .cin(s_wallace_cska32_and_20_21[0]), .fa_xor1(s_wallace_cska32_fa303_xor1), .fa_or0(s_wallace_cska32_fa303_or0));
  and_gate and_gate_s_wallace_cska32_and_21_21(.a(a[21]), .b(b[21]), .out(s_wallace_cska32_and_21_21));
  and_gate and_gate_s_wallace_cska32_and_20_22(.a(a[20]), .b(b[22]), .out(s_wallace_cska32_and_20_22));
  fa fa_s_wallace_cska32_fa304_out(.a(s_wallace_cska32_fa303_or0[0]), .b(s_wallace_cska32_and_21_21[0]), .cin(s_wallace_cska32_and_20_22[0]), .fa_xor1(s_wallace_cska32_fa304_xor1), .fa_or0(s_wallace_cska32_fa304_or0));
  and_gate and_gate_s_wallace_cska32_and_21_22(.a(a[21]), .b(b[22]), .out(s_wallace_cska32_and_21_22));
  and_gate and_gate_s_wallace_cska32_and_20_23(.a(a[20]), .b(b[23]), .out(s_wallace_cska32_and_20_23));
  fa fa_s_wallace_cska32_fa305_out(.a(s_wallace_cska32_fa304_or0[0]), .b(s_wallace_cska32_and_21_22[0]), .cin(s_wallace_cska32_and_20_23[0]), .fa_xor1(s_wallace_cska32_fa305_xor1), .fa_or0(s_wallace_cska32_fa305_or0));
  and_gate and_gate_s_wallace_cska32_and_21_23(.a(a[21]), .b(b[23]), .out(s_wallace_cska32_and_21_23));
  and_gate and_gate_s_wallace_cska32_and_20_24(.a(a[20]), .b(b[24]), .out(s_wallace_cska32_and_20_24));
  fa fa_s_wallace_cska32_fa306_out(.a(s_wallace_cska32_fa305_or0[0]), .b(s_wallace_cska32_and_21_23[0]), .cin(s_wallace_cska32_and_20_24[0]), .fa_xor1(s_wallace_cska32_fa306_xor1), .fa_or0(s_wallace_cska32_fa306_or0));
  and_gate and_gate_s_wallace_cska32_and_21_24(.a(a[21]), .b(b[24]), .out(s_wallace_cska32_and_21_24));
  and_gate and_gate_s_wallace_cska32_and_20_25(.a(a[20]), .b(b[25]), .out(s_wallace_cska32_and_20_25));
  fa fa_s_wallace_cska32_fa307_out(.a(s_wallace_cska32_fa306_or0[0]), .b(s_wallace_cska32_and_21_24[0]), .cin(s_wallace_cska32_and_20_25[0]), .fa_xor1(s_wallace_cska32_fa307_xor1), .fa_or0(s_wallace_cska32_fa307_or0));
  and_gate and_gate_s_wallace_cska32_and_21_25(.a(a[21]), .b(b[25]), .out(s_wallace_cska32_and_21_25));
  and_gate and_gate_s_wallace_cska32_and_20_26(.a(a[20]), .b(b[26]), .out(s_wallace_cska32_and_20_26));
  fa fa_s_wallace_cska32_fa308_out(.a(s_wallace_cska32_fa307_or0[0]), .b(s_wallace_cska32_and_21_25[0]), .cin(s_wallace_cska32_and_20_26[0]), .fa_xor1(s_wallace_cska32_fa308_xor1), .fa_or0(s_wallace_cska32_fa308_or0));
  and_gate and_gate_s_wallace_cska32_and_21_26(.a(a[21]), .b(b[26]), .out(s_wallace_cska32_and_21_26));
  and_gate and_gate_s_wallace_cska32_and_20_27(.a(a[20]), .b(b[27]), .out(s_wallace_cska32_and_20_27));
  fa fa_s_wallace_cska32_fa309_out(.a(s_wallace_cska32_fa308_or0[0]), .b(s_wallace_cska32_and_21_26[0]), .cin(s_wallace_cska32_and_20_27[0]), .fa_xor1(s_wallace_cska32_fa309_xor1), .fa_or0(s_wallace_cska32_fa309_or0));
  and_gate and_gate_s_wallace_cska32_and_21_27(.a(a[21]), .b(b[27]), .out(s_wallace_cska32_and_21_27));
  and_gate and_gate_s_wallace_cska32_and_20_28(.a(a[20]), .b(b[28]), .out(s_wallace_cska32_and_20_28));
  fa fa_s_wallace_cska32_fa310_out(.a(s_wallace_cska32_fa309_or0[0]), .b(s_wallace_cska32_and_21_27[0]), .cin(s_wallace_cska32_and_20_28[0]), .fa_xor1(s_wallace_cska32_fa310_xor1), .fa_or0(s_wallace_cska32_fa310_or0));
  and_gate and_gate_s_wallace_cska32_and_21_28(.a(a[21]), .b(b[28]), .out(s_wallace_cska32_and_21_28));
  and_gate and_gate_s_wallace_cska32_and_20_29(.a(a[20]), .b(b[29]), .out(s_wallace_cska32_and_20_29));
  fa fa_s_wallace_cska32_fa311_out(.a(s_wallace_cska32_fa310_or0[0]), .b(s_wallace_cska32_and_21_28[0]), .cin(s_wallace_cska32_and_20_29[0]), .fa_xor1(s_wallace_cska32_fa311_xor1), .fa_or0(s_wallace_cska32_fa311_or0));
  and_gate and_gate_s_wallace_cska32_and_21_29(.a(a[21]), .b(b[29]), .out(s_wallace_cska32_and_21_29));
  and_gate and_gate_s_wallace_cska32_and_20_30(.a(a[20]), .b(b[30]), .out(s_wallace_cska32_and_20_30));
  fa fa_s_wallace_cska32_fa312_out(.a(s_wallace_cska32_fa311_or0[0]), .b(s_wallace_cska32_and_21_29[0]), .cin(s_wallace_cska32_and_20_30[0]), .fa_xor1(s_wallace_cska32_fa312_xor1), .fa_or0(s_wallace_cska32_fa312_or0));
  and_gate and_gate_s_wallace_cska32_and_21_30(.a(a[21]), .b(b[30]), .out(s_wallace_cska32_and_21_30));
  nand_gate nand_gate_s_wallace_cska32_nand_20_31(.a(a[20]), .b(b[31]), .out(s_wallace_cska32_nand_20_31));
  fa fa_s_wallace_cska32_fa313_out(.a(s_wallace_cska32_fa312_or0[0]), .b(s_wallace_cska32_and_21_30[0]), .cin(s_wallace_cska32_nand_20_31[0]), .fa_xor1(s_wallace_cska32_fa313_xor1), .fa_or0(s_wallace_cska32_fa313_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_21_31(.a(a[21]), .b(b[31]), .out(s_wallace_cska32_nand_21_31));
  fa fa_s_wallace_cska32_fa314_out(.a(s_wallace_cska32_fa313_or0[0]), .b(s_wallace_cska32_nand_21_31[0]), .cin(s_wallace_cska32_fa49_xor1[0]), .fa_xor1(s_wallace_cska32_fa314_xor1), .fa_or0(s_wallace_cska32_fa314_or0));
  fa fa_s_wallace_cska32_fa315_out(.a(s_wallace_cska32_fa314_or0[0]), .b(s_wallace_cska32_fa50_xor1[0]), .cin(s_wallace_cska32_fa107_xor1[0]), .fa_xor1(s_wallace_cska32_fa315_xor1), .fa_or0(s_wallace_cska32_fa315_or0));
  fa fa_s_wallace_cska32_fa316_out(.a(s_wallace_cska32_fa315_or0[0]), .b(s_wallace_cska32_fa108_xor1[0]), .cin(s_wallace_cska32_fa163_xor1[0]), .fa_xor1(s_wallace_cska32_fa316_xor1), .fa_or0(s_wallace_cska32_fa316_or0));
  fa fa_s_wallace_cska32_fa317_out(.a(s_wallace_cska32_fa316_or0[0]), .b(s_wallace_cska32_fa164_xor1[0]), .cin(s_wallace_cska32_fa217_xor1[0]), .fa_xor1(s_wallace_cska32_fa317_xor1), .fa_or0(s_wallace_cska32_fa317_or0));
  ha ha_s_wallace_cska32_ha6_out(.a(s_wallace_cska32_fa170_xor1[0]), .b(s_wallace_cska32_fa221_xor1[0]), .ha_xor0(s_wallace_cska32_ha6_xor0), .ha_and0(s_wallace_cska32_ha6_and0));
  fa fa_s_wallace_cska32_fa318_out(.a(s_wallace_cska32_ha6_and0[0]), .b(s_wallace_cska32_fa118_xor1[0]), .cin(s_wallace_cska32_fa171_xor1[0]), .fa_xor1(s_wallace_cska32_fa318_xor1), .fa_or0(s_wallace_cska32_fa318_or0));
  fa fa_s_wallace_cska32_fa319_out(.a(s_wallace_cska32_fa318_or0[0]), .b(s_wallace_cska32_fa64_xor1[0]), .cin(s_wallace_cska32_fa119_xor1[0]), .fa_xor1(s_wallace_cska32_fa319_xor1), .fa_or0(s_wallace_cska32_fa319_or0));
  fa fa_s_wallace_cska32_fa320_out(.a(s_wallace_cska32_fa319_or0[0]), .b(s_wallace_cska32_fa8_xor1[0]), .cin(s_wallace_cska32_fa65_xor1[0]), .fa_xor1(s_wallace_cska32_fa320_xor1), .fa_or0(s_wallace_cska32_fa320_or0));
  and_gate and_gate_s_wallace_cska32_and_0_12(.a(a[0]), .b(b[12]), .out(s_wallace_cska32_and_0_12));
  fa fa_s_wallace_cska32_fa321_out(.a(s_wallace_cska32_fa320_or0[0]), .b(s_wallace_cska32_and_0_12[0]), .cin(s_wallace_cska32_fa9_xor1[0]), .fa_xor1(s_wallace_cska32_fa321_xor1), .fa_or0(s_wallace_cska32_fa321_or0));
  and_gate and_gate_s_wallace_cska32_and_1_12(.a(a[1]), .b(b[12]), .out(s_wallace_cska32_and_1_12));
  and_gate and_gate_s_wallace_cska32_and_0_13(.a(a[0]), .b(b[13]), .out(s_wallace_cska32_and_0_13));
  fa fa_s_wallace_cska32_fa322_out(.a(s_wallace_cska32_fa321_or0[0]), .b(s_wallace_cska32_and_1_12[0]), .cin(s_wallace_cska32_and_0_13[0]), .fa_xor1(s_wallace_cska32_fa322_xor1), .fa_or0(s_wallace_cska32_fa322_or0));
  and_gate and_gate_s_wallace_cska32_and_2_12(.a(a[2]), .b(b[12]), .out(s_wallace_cska32_and_2_12));
  and_gate and_gate_s_wallace_cska32_and_1_13(.a(a[1]), .b(b[13]), .out(s_wallace_cska32_and_1_13));
  fa fa_s_wallace_cska32_fa323_out(.a(s_wallace_cska32_fa322_or0[0]), .b(s_wallace_cska32_and_2_12[0]), .cin(s_wallace_cska32_and_1_13[0]), .fa_xor1(s_wallace_cska32_fa323_xor1), .fa_or0(s_wallace_cska32_fa323_or0));
  and_gate and_gate_s_wallace_cska32_and_3_12(.a(a[3]), .b(b[12]), .out(s_wallace_cska32_and_3_12));
  and_gate and_gate_s_wallace_cska32_and_2_13(.a(a[2]), .b(b[13]), .out(s_wallace_cska32_and_2_13));
  fa fa_s_wallace_cska32_fa324_out(.a(s_wallace_cska32_fa323_or0[0]), .b(s_wallace_cska32_and_3_12[0]), .cin(s_wallace_cska32_and_2_13[0]), .fa_xor1(s_wallace_cska32_fa324_xor1), .fa_or0(s_wallace_cska32_fa324_or0));
  and_gate and_gate_s_wallace_cska32_and_4_12(.a(a[4]), .b(b[12]), .out(s_wallace_cska32_and_4_12));
  and_gate and_gate_s_wallace_cska32_and_3_13(.a(a[3]), .b(b[13]), .out(s_wallace_cska32_and_3_13));
  fa fa_s_wallace_cska32_fa325_out(.a(s_wallace_cska32_fa324_or0[0]), .b(s_wallace_cska32_and_4_12[0]), .cin(s_wallace_cska32_and_3_13[0]), .fa_xor1(s_wallace_cska32_fa325_xor1), .fa_or0(s_wallace_cska32_fa325_or0));
  and_gate and_gate_s_wallace_cska32_and_5_12(.a(a[5]), .b(b[12]), .out(s_wallace_cska32_and_5_12));
  and_gate and_gate_s_wallace_cska32_and_4_13(.a(a[4]), .b(b[13]), .out(s_wallace_cska32_and_4_13));
  fa fa_s_wallace_cska32_fa326_out(.a(s_wallace_cska32_fa325_or0[0]), .b(s_wallace_cska32_and_5_12[0]), .cin(s_wallace_cska32_and_4_13[0]), .fa_xor1(s_wallace_cska32_fa326_xor1), .fa_or0(s_wallace_cska32_fa326_or0));
  and_gate and_gate_s_wallace_cska32_and_6_12(.a(a[6]), .b(b[12]), .out(s_wallace_cska32_and_6_12));
  and_gate and_gate_s_wallace_cska32_and_5_13(.a(a[5]), .b(b[13]), .out(s_wallace_cska32_and_5_13));
  fa fa_s_wallace_cska32_fa327_out(.a(s_wallace_cska32_fa326_or0[0]), .b(s_wallace_cska32_and_6_12[0]), .cin(s_wallace_cska32_and_5_13[0]), .fa_xor1(s_wallace_cska32_fa327_xor1), .fa_or0(s_wallace_cska32_fa327_or0));
  and_gate and_gate_s_wallace_cska32_and_7_12(.a(a[7]), .b(b[12]), .out(s_wallace_cska32_and_7_12));
  and_gate and_gate_s_wallace_cska32_and_6_13(.a(a[6]), .b(b[13]), .out(s_wallace_cska32_and_6_13));
  fa fa_s_wallace_cska32_fa328_out(.a(s_wallace_cska32_fa327_or0[0]), .b(s_wallace_cska32_and_7_12[0]), .cin(s_wallace_cska32_and_6_13[0]), .fa_xor1(s_wallace_cska32_fa328_xor1), .fa_or0(s_wallace_cska32_fa328_or0));
  and_gate and_gate_s_wallace_cska32_and_8_12(.a(a[8]), .b(b[12]), .out(s_wallace_cska32_and_8_12));
  and_gate and_gate_s_wallace_cska32_and_7_13(.a(a[7]), .b(b[13]), .out(s_wallace_cska32_and_7_13));
  fa fa_s_wallace_cska32_fa329_out(.a(s_wallace_cska32_fa328_or0[0]), .b(s_wallace_cska32_and_8_12[0]), .cin(s_wallace_cska32_and_7_13[0]), .fa_xor1(s_wallace_cska32_fa329_xor1), .fa_or0(s_wallace_cska32_fa329_or0));
  and_gate and_gate_s_wallace_cska32_and_9_12(.a(a[9]), .b(b[12]), .out(s_wallace_cska32_and_9_12));
  and_gate and_gate_s_wallace_cska32_and_8_13(.a(a[8]), .b(b[13]), .out(s_wallace_cska32_and_8_13));
  fa fa_s_wallace_cska32_fa330_out(.a(s_wallace_cska32_fa329_or0[0]), .b(s_wallace_cska32_and_9_12[0]), .cin(s_wallace_cska32_and_8_13[0]), .fa_xor1(s_wallace_cska32_fa330_xor1), .fa_or0(s_wallace_cska32_fa330_or0));
  and_gate and_gate_s_wallace_cska32_and_10_12(.a(a[10]), .b(b[12]), .out(s_wallace_cska32_and_10_12));
  and_gate and_gate_s_wallace_cska32_and_9_13(.a(a[9]), .b(b[13]), .out(s_wallace_cska32_and_9_13));
  fa fa_s_wallace_cska32_fa331_out(.a(s_wallace_cska32_fa330_or0[0]), .b(s_wallace_cska32_and_10_12[0]), .cin(s_wallace_cska32_and_9_13[0]), .fa_xor1(s_wallace_cska32_fa331_xor1), .fa_or0(s_wallace_cska32_fa331_or0));
  and_gate and_gate_s_wallace_cska32_and_11_12(.a(a[11]), .b(b[12]), .out(s_wallace_cska32_and_11_12));
  and_gate and_gate_s_wallace_cska32_and_10_13(.a(a[10]), .b(b[13]), .out(s_wallace_cska32_and_10_13));
  fa fa_s_wallace_cska32_fa332_out(.a(s_wallace_cska32_fa331_or0[0]), .b(s_wallace_cska32_and_11_12[0]), .cin(s_wallace_cska32_and_10_13[0]), .fa_xor1(s_wallace_cska32_fa332_xor1), .fa_or0(s_wallace_cska32_fa332_or0));
  and_gate and_gate_s_wallace_cska32_and_12_12(.a(a[12]), .b(b[12]), .out(s_wallace_cska32_and_12_12));
  and_gate and_gate_s_wallace_cska32_and_11_13(.a(a[11]), .b(b[13]), .out(s_wallace_cska32_and_11_13));
  fa fa_s_wallace_cska32_fa333_out(.a(s_wallace_cska32_fa332_or0[0]), .b(s_wallace_cska32_and_12_12[0]), .cin(s_wallace_cska32_and_11_13[0]), .fa_xor1(s_wallace_cska32_fa333_xor1), .fa_or0(s_wallace_cska32_fa333_or0));
  and_gate and_gate_s_wallace_cska32_and_13_12(.a(a[13]), .b(b[12]), .out(s_wallace_cska32_and_13_12));
  and_gate and_gate_s_wallace_cska32_and_12_13(.a(a[12]), .b(b[13]), .out(s_wallace_cska32_and_12_13));
  fa fa_s_wallace_cska32_fa334_out(.a(s_wallace_cska32_fa333_or0[0]), .b(s_wallace_cska32_and_13_12[0]), .cin(s_wallace_cska32_and_12_13[0]), .fa_xor1(s_wallace_cska32_fa334_xor1), .fa_or0(s_wallace_cska32_fa334_or0));
  and_gate and_gate_s_wallace_cska32_and_14_12(.a(a[14]), .b(b[12]), .out(s_wallace_cska32_and_14_12));
  and_gate and_gate_s_wallace_cska32_and_13_13(.a(a[13]), .b(b[13]), .out(s_wallace_cska32_and_13_13));
  fa fa_s_wallace_cska32_fa335_out(.a(s_wallace_cska32_fa334_or0[0]), .b(s_wallace_cska32_and_14_12[0]), .cin(s_wallace_cska32_and_13_13[0]), .fa_xor1(s_wallace_cska32_fa335_xor1), .fa_or0(s_wallace_cska32_fa335_or0));
  and_gate and_gate_s_wallace_cska32_and_15_12(.a(a[15]), .b(b[12]), .out(s_wallace_cska32_and_15_12));
  and_gate and_gate_s_wallace_cska32_and_14_13(.a(a[14]), .b(b[13]), .out(s_wallace_cska32_and_14_13));
  fa fa_s_wallace_cska32_fa336_out(.a(s_wallace_cska32_fa335_or0[0]), .b(s_wallace_cska32_and_15_12[0]), .cin(s_wallace_cska32_and_14_13[0]), .fa_xor1(s_wallace_cska32_fa336_xor1), .fa_or0(s_wallace_cska32_fa336_or0));
  and_gate and_gate_s_wallace_cska32_and_16_12(.a(a[16]), .b(b[12]), .out(s_wallace_cska32_and_16_12));
  and_gate and_gate_s_wallace_cska32_and_15_13(.a(a[15]), .b(b[13]), .out(s_wallace_cska32_and_15_13));
  fa fa_s_wallace_cska32_fa337_out(.a(s_wallace_cska32_fa336_or0[0]), .b(s_wallace_cska32_and_16_12[0]), .cin(s_wallace_cska32_and_15_13[0]), .fa_xor1(s_wallace_cska32_fa337_xor1), .fa_or0(s_wallace_cska32_fa337_or0));
  and_gate and_gate_s_wallace_cska32_and_17_12(.a(a[17]), .b(b[12]), .out(s_wallace_cska32_and_17_12));
  and_gate and_gate_s_wallace_cska32_and_16_13(.a(a[16]), .b(b[13]), .out(s_wallace_cska32_and_16_13));
  fa fa_s_wallace_cska32_fa338_out(.a(s_wallace_cska32_fa337_or0[0]), .b(s_wallace_cska32_and_17_12[0]), .cin(s_wallace_cska32_and_16_13[0]), .fa_xor1(s_wallace_cska32_fa338_xor1), .fa_or0(s_wallace_cska32_fa338_or0));
  and_gate and_gate_s_wallace_cska32_and_18_12(.a(a[18]), .b(b[12]), .out(s_wallace_cska32_and_18_12));
  and_gate and_gate_s_wallace_cska32_and_17_13(.a(a[17]), .b(b[13]), .out(s_wallace_cska32_and_17_13));
  fa fa_s_wallace_cska32_fa339_out(.a(s_wallace_cska32_fa338_or0[0]), .b(s_wallace_cska32_and_18_12[0]), .cin(s_wallace_cska32_and_17_13[0]), .fa_xor1(s_wallace_cska32_fa339_xor1), .fa_or0(s_wallace_cska32_fa339_or0));
  and_gate and_gate_s_wallace_cska32_and_19_12(.a(a[19]), .b(b[12]), .out(s_wallace_cska32_and_19_12));
  and_gate and_gate_s_wallace_cska32_and_18_13(.a(a[18]), .b(b[13]), .out(s_wallace_cska32_and_18_13));
  fa fa_s_wallace_cska32_fa340_out(.a(s_wallace_cska32_fa339_or0[0]), .b(s_wallace_cska32_and_19_12[0]), .cin(s_wallace_cska32_and_18_13[0]), .fa_xor1(s_wallace_cska32_fa340_xor1), .fa_or0(s_wallace_cska32_fa340_or0));
  and_gate and_gate_s_wallace_cska32_and_20_12(.a(a[20]), .b(b[12]), .out(s_wallace_cska32_and_20_12));
  and_gate and_gate_s_wallace_cska32_and_19_13(.a(a[19]), .b(b[13]), .out(s_wallace_cska32_and_19_13));
  fa fa_s_wallace_cska32_fa341_out(.a(s_wallace_cska32_fa340_or0[0]), .b(s_wallace_cska32_and_20_12[0]), .cin(s_wallace_cska32_and_19_13[0]), .fa_xor1(s_wallace_cska32_fa341_xor1), .fa_or0(s_wallace_cska32_fa341_or0));
  and_gate and_gate_s_wallace_cska32_and_19_14(.a(a[19]), .b(b[14]), .out(s_wallace_cska32_and_19_14));
  and_gate and_gate_s_wallace_cska32_and_18_15(.a(a[18]), .b(b[15]), .out(s_wallace_cska32_and_18_15));
  fa fa_s_wallace_cska32_fa342_out(.a(s_wallace_cska32_fa341_or0[0]), .b(s_wallace_cska32_and_19_14[0]), .cin(s_wallace_cska32_and_18_15[0]), .fa_xor1(s_wallace_cska32_fa342_xor1), .fa_or0(s_wallace_cska32_fa342_or0));
  and_gate and_gate_s_wallace_cska32_and_19_15(.a(a[19]), .b(b[15]), .out(s_wallace_cska32_and_19_15));
  and_gate and_gate_s_wallace_cska32_and_18_16(.a(a[18]), .b(b[16]), .out(s_wallace_cska32_and_18_16));
  fa fa_s_wallace_cska32_fa343_out(.a(s_wallace_cska32_fa342_or0[0]), .b(s_wallace_cska32_and_19_15[0]), .cin(s_wallace_cska32_and_18_16[0]), .fa_xor1(s_wallace_cska32_fa343_xor1), .fa_or0(s_wallace_cska32_fa343_or0));
  and_gate and_gate_s_wallace_cska32_and_19_16(.a(a[19]), .b(b[16]), .out(s_wallace_cska32_and_19_16));
  and_gate and_gate_s_wallace_cska32_and_18_17(.a(a[18]), .b(b[17]), .out(s_wallace_cska32_and_18_17));
  fa fa_s_wallace_cska32_fa344_out(.a(s_wallace_cska32_fa343_or0[0]), .b(s_wallace_cska32_and_19_16[0]), .cin(s_wallace_cska32_and_18_17[0]), .fa_xor1(s_wallace_cska32_fa344_xor1), .fa_or0(s_wallace_cska32_fa344_or0));
  and_gate and_gate_s_wallace_cska32_and_19_17(.a(a[19]), .b(b[17]), .out(s_wallace_cska32_and_19_17));
  and_gate and_gate_s_wallace_cska32_and_18_18(.a(a[18]), .b(b[18]), .out(s_wallace_cska32_and_18_18));
  fa fa_s_wallace_cska32_fa345_out(.a(s_wallace_cska32_fa344_or0[0]), .b(s_wallace_cska32_and_19_17[0]), .cin(s_wallace_cska32_and_18_18[0]), .fa_xor1(s_wallace_cska32_fa345_xor1), .fa_or0(s_wallace_cska32_fa345_or0));
  and_gate and_gate_s_wallace_cska32_and_19_18(.a(a[19]), .b(b[18]), .out(s_wallace_cska32_and_19_18));
  and_gate and_gate_s_wallace_cska32_and_18_19(.a(a[18]), .b(b[19]), .out(s_wallace_cska32_and_18_19));
  fa fa_s_wallace_cska32_fa346_out(.a(s_wallace_cska32_fa345_or0[0]), .b(s_wallace_cska32_and_19_18[0]), .cin(s_wallace_cska32_and_18_19[0]), .fa_xor1(s_wallace_cska32_fa346_xor1), .fa_or0(s_wallace_cska32_fa346_or0));
  and_gate and_gate_s_wallace_cska32_and_19_19(.a(a[19]), .b(b[19]), .out(s_wallace_cska32_and_19_19));
  and_gate and_gate_s_wallace_cska32_and_18_20(.a(a[18]), .b(b[20]), .out(s_wallace_cska32_and_18_20));
  fa fa_s_wallace_cska32_fa347_out(.a(s_wallace_cska32_fa346_or0[0]), .b(s_wallace_cska32_and_19_19[0]), .cin(s_wallace_cska32_and_18_20[0]), .fa_xor1(s_wallace_cska32_fa347_xor1), .fa_or0(s_wallace_cska32_fa347_or0));
  and_gate and_gate_s_wallace_cska32_and_19_20(.a(a[19]), .b(b[20]), .out(s_wallace_cska32_and_19_20));
  and_gate and_gate_s_wallace_cska32_and_18_21(.a(a[18]), .b(b[21]), .out(s_wallace_cska32_and_18_21));
  fa fa_s_wallace_cska32_fa348_out(.a(s_wallace_cska32_fa347_or0[0]), .b(s_wallace_cska32_and_19_20[0]), .cin(s_wallace_cska32_and_18_21[0]), .fa_xor1(s_wallace_cska32_fa348_xor1), .fa_or0(s_wallace_cska32_fa348_or0));
  and_gate and_gate_s_wallace_cska32_and_19_21(.a(a[19]), .b(b[21]), .out(s_wallace_cska32_and_19_21));
  and_gate and_gate_s_wallace_cska32_and_18_22(.a(a[18]), .b(b[22]), .out(s_wallace_cska32_and_18_22));
  fa fa_s_wallace_cska32_fa349_out(.a(s_wallace_cska32_fa348_or0[0]), .b(s_wallace_cska32_and_19_21[0]), .cin(s_wallace_cska32_and_18_22[0]), .fa_xor1(s_wallace_cska32_fa349_xor1), .fa_or0(s_wallace_cska32_fa349_or0));
  and_gate and_gate_s_wallace_cska32_and_19_22(.a(a[19]), .b(b[22]), .out(s_wallace_cska32_and_19_22));
  and_gate and_gate_s_wallace_cska32_and_18_23(.a(a[18]), .b(b[23]), .out(s_wallace_cska32_and_18_23));
  fa fa_s_wallace_cska32_fa350_out(.a(s_wallace_cska32_fa349_or0[0]), .b(s_wallace_cska32_and_19_22[0]), .cin(s_wallace_cska32_and_18_23[0]), .fa_xor1(s_wallace_cska32_fa350_xor1), .fa_or0(s_wallace_cska32_fa350_or0));
  and_gate and_gate_s_wallace_cska32_and_19_23(.a(a[19]), .b(b[23]), .out(s_wallace_cska32_and_19_23));
  and_gate and_gate_s_wallace_cska32_and_18_24(.a(a[18]), .b(b[24]), .out(s_wallace_cska32_and_18_24));
  fa fa_s_wallace_cska32_fa351_out(.a(s_wallace_cska32_fa350_or0[0]), .b(s_wallace_cska32_and_19_23[0]), .cin(s_wallace_cska32_and_18_24[0]), .fa_xor1(s_wallace_cska32_fa351_xor1), .fa_or0(s_wallace_cska32_fa351_or0));
  and_gate and_gate_s_wallace_cska32_and_19_24(.a(a[19]), .b(b[24]), .out(s_wallace_cska32_and_19_24));
  and_gate and_gate_s_wallace_cska32_and_18_25(.a(a[18]), .b(b[25]), .out(s_wallace_cska32_and_18_25));
  fa fa_s_wallace_cska32_fa352_out(.a(s_wallace_cska32_fa351_or0[0]), .b(s_wallace_cska32_and_19_24[0]), .cin(s_wallace_cska32_and_18_25[0]), .fa_xor1(s_wallace_cska32_fa352_xor1), .fa_or0(s_wallace_cska32_fa352_or0));
  and_gate and_gate_s_wallace_cska32_and_19_25(.a(a[19]), .b(b[25]), .out(s_wallace_cska32_and_19_25));
  and_gate and_gate_s_wallace_cska32_and_18_26(.a(a[18]), .b(b[26]), .out(s_wallace_cska32_and_18_26));
  fa fa_s_wallace_cska32_fa353_out(.a(s_wallace_cska32_fa352_or0[0]), .b(s_wallace_cska32_and_19_25[0]), .cin(s_wallace_cska32_and_18_26[0]), .fa_xor1(s_wallace_cska32_fa353_xor1), .fa_or0(s_wallace_cska32_fa353_or0));
  and_gate and_gate_s_wallace_cska32_and_19_26(.a(a[19]), .b(b[26]), .out(s_wallace_cska32_and_19_26));
  and_gate and_gate_s_wallace_cska32_and_18_27(.a(a[18]), .b(b[27]), .out(s_wallace_cska32_and_18_27));
  fa fa_s_wallace_cska32_fa354_out(.a(s_wallace_cska32_fa353_or0[0]), .b(s_wallace_cska32_and_19_26[0]), .cin(s_wallace_cska32_and_18_27[0]), .fa_xor1(s_wallace_cska32_fa354_xor1), .fa_or0(s_wallace_cska32_fa354_or0));
  and_gate and_gate_s_wallace_cska32_and_19_27(.a(a[19]), .b(b[27]), .out(s_wallace_cska32_and_19_27));
  and_gate and_gate_s_wallace_cska32_and_18_28(.a(a[18]), .b(b[28]), .out(s_wallace_cska32_and_18_28));
  fa fa_s_wallace_cska32_fa355_out(.a(s_wallace_cska32_fa354_or0[0]), .b(s_wallace_cska32_and_19_27[0]), .cin(s_wallace_cska32_and_18_28[0]), .fa_xor1(s_wallace_cska32_fa355_xor1), .fa_or0(s_wallace_cska32_fa355_or0));
  and_gate and_gate_s_wallace_cska32_and_19_28(.a(a[19]), .b(b[28]), .out(s_wallace_cska32_and_19_28));
  and_gate and_gate_s_wallace_cska32_and_18_29(.a(a[18]), .b(b[29]), .out(s_wallace_cska32_and_18_29));
  fa fa_s_wallace_cska32_fa356_out(.a(s_wallace_cska32_fa355_or0[0]), .b(s_wallace_cska32_and_19_28[0]), .cin(s_wallace_cska32_and_18_29[0]), .fa_xor1(s_wallace_cska32_fa356_xor1), .fa_or0(s_wallace_cska32_fa356_or0));
  and_gate and_gate_s_wallace_cska32_and_19_29(.a(a[19]), .b(b[29]), .out(s_wallace_cska32_and_19_29));
  and_gate and_gate_s_wallace_cska32_and_18_30(.a(a[18]), .b(b[30]), .out(s_wallace_cska32_and_18_30));
  fa fa_s_wallace_cska32_fa357_out(.a(s_wallace_cska32_fa356_or0[0]), .b(s_wallace_cska32_and_19_29[0]), .cin(s_wallace_cska32_and_18_30[0]), .fa_xor1(s_wallace_cska32_fa357_xor1), .fa_or0(s_wallace_cska32_fa357_or0));
  and_gate and_gate_s_wallace_cska32_and_19_30(.a(a[19]), .b(b[30]), .out(s_wallace_cska32_and_19_30));
  nand_gate nand_gate_s_wallace_cska32_nand_18_31(.a(a[18]), .b(b[31]), .out(s_wallace_cska32_nand_18_31));
  fa fa_s_wallace_cska32_fa358_out(.a(s_wallace_cska32_fa357_or0[0]), .b(s_wallace_cska32_and_19_30[0]), .cin(s_wallace_cska32_nand_18_31[0]), .fa_xor1(s_wallace_cska32_fa358_xor1), .fa_or0(s_wallace_cska32_fa358_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_19_31(.a(a[19]), .b(b[31]), .out(s_wallace_cska32_nand_19_31));
  fa fa_s_wallace_cska32_fa359_out(.a(s_wallace_cska32_fa358_or0[0]), .b(s_wallace_cska32_nand_19_31[0]), .cin(s_wallace_cska32_fa47_xor1[0]), .fa_xor1(s_wallace_cska32_fa359_xor1), .fa_or0(s_wallace_cska32_fa359_or0));
  fa fa_s_wallace_cska32_fa360_out(.a(s_wallace_cska32_fa359_or0[0]), .b(s_wallace_cska32_fa48_xor1[0]), .cin(s_wallace_cska32_fa105_xor1[0]), .fa_xor1(s_wallace_cska32_fa360_xor1), .fa_or0(s_wallace_cska32_fa360_or0));
  fa fa_s_wallace_cska32_fa361_out(.a(s_wallace_cska32_fa360_or0[0]), .b(s_wallace_cska32_fa106_xor1[0]), .cin(s_wallace_cska32_fa161_xor1[0]), .fa_xor1(s_wallace_cska32_fa361_xor1), .fa_or0(s_wallace_cska32_fa361_or0));
  fa fa_s_wallace_cska32_fa362_out(.a(s_wallace_cska32_fa361_or0[0]), .b(s_wallace_cska32_fa162_xor1[0]), .cin(s_wallace_cska32_fa215_xor1[0]), .fa_xor1(s_wallace_cska32_fa362_xor1), .fa_or0(s_wallace_cska32_fa362_or0));
  fa fa_s_wallace_cska32_fa363_out(.a(s_wallace_cska32_fa362_or0[0]), .b(s_wallace_cska32_fa216_xor1[0]), .cin(s_wallace_cska32_fa267_xor1[0]), .fa_xor1(s_wallace_cska32_fa363_xor1), .fa_or0(s_wallace_cska32_fa363_or0));
  ha ha_s_wallace_cska32_ha7_out(.a(s_wallace_cska32_fa222_xor1[0]), .b(s_wallace_cska32_fa271_xor1[0]), .ha_xor0(s_wallace_cska32_ha7_xor0), .ha_and0(s_wallace_cska32_ha7_and0));
  fa fa_s_wallace_cska32_fa364_out(.a(s_wallace_cska32_ha7_and0[0]), .b(s_wallace_cska32_fa172_xor1[0]), .cin(s_wallace_cska32_fa223_xor1[0]), .fa_xor1(s_wallace_cska32_fa364_xor1), .fa_or0(s_wallace_cska32_fa364_or0));
  fa fa_s_wallace_cska32_fa365_out(.a(s_wallace_cska32_fa364_or0[0]), .b(s_wallace_cska32_fa120_xor1[0]), .cin(s_wallace_cska32_fa173_xor1[0]), .fa_xor1(s_wallace_cska32_fa365_xor1), .fa_or0(s_wallace_cska32_fa365_or0));
  fa fa_s_wallace_cska32_fa366_out(.a(s_wallace_cska32_fa365_or0[0]), .b(s_wallace_cska32_fa66_xor1[0]), .cin(s_wallace_cska32_fa121_xor1[0]), .fa_xor1(s_wallace_cska32_fa366_xor1), .fa_or0(s_wallace_cska32_fa366_or0));
  fa fa_s_wallace_cska32_fa367_out(.a(s_wallace_cska32_fa366_or0[0]), .b(s_wallace_cska32_fa10_xor1[0]), .cin(s_wallace_cska32_fa67_xor1[0]), .fa_xor1(s_wallace_cska32_fa367_xor1), .fa_or0(s_wallace_cska32_fa367_or0));
  and_gate and_gate_s_wallace_cska32_and_0_14(.a(a[0]), .b(b[14]), .out(s_wallace_cska32_and_0_14));
  fa fa_s_wallace_cska32_fa368_out(.a(s_wallace_cska32_fa367_or0[0]), .b(s_wallace_cska32_and_0_14[0]), .cin(s_wallace_cska32_fa11_xor1[0]), .fa_xor1(s_wallace_cska32_fa368_xor1), .fa_or0(s_wallace_cska32_fa368_or0));
  and_gate and_gate_s_wallace_cska32_and_1_14(.a(a[1]), .b(b[14]), .out(s_wallace_cska32_and_1_14));
  and_gate and_gate_s_wallace_cska32_and_0_15(.a(a[0]), .b(b[15]), .out(s_wallace_cska32_and_0_15));
  fa fa_s_wallace_cska32_fa369_out(.a(s_wallace_cska32_fa368_or0[0]), .b(s_wallace_cska32_and_1_14[0]), .cin(s_wallace_cska32_and_0_15[0]), .fa_xor1(s_wallace_cska32_fa369_xor1), .fa_or0(s_wallace_cska32_fa369_or0));
  and_gate and_gate_s_wallace_cska32_and_2_14(.a(a[2]), .b(b[14]), .out(s_wallace_cska32_and_2_14));
  and_gate and_gate_s_wallace_cska32_and_1_15(.a(a[1]), .b(b[15]), .out(s_wallace_cska32_and_1_15));
  fa fa_s_wallace_cska32_fa370_out(.a(s_wallace_cska32_fa369_or0[0]), .b(s_wallace_cska32_and_2_14[0]), .cin(s_wallace_cska32_and_1_15[0]), .fa_xor1(s_wallace_cska32_fa370_xor1), .fa_or0(s_wallace_cska32_fa370_or0));
  and_gate and_gate_s_wallace_cska32_and_3_14(.a(a[3]), .b(b[14]), .out(s_wallace_cska32_and_3_14));
  and_gate and_gate_s_wallace_cska32_and_2_15(.a(a[2]), .b(b[15]), .out(s_wallace_cska32_and_2_15));
  fa fa_s_wallace_cska32_fa371_out(.a(s_wallace_cska32_fa370_or0[0]), .b(s_wallace_cska32_and_3_14[0]), .cin(s_wallace_cska32_and_2_15[0]), .fa_xor1(s_wallace_cska32_fa371_xor1), .fa_or0(s_wallace_cska32_fa371_or0));
  and_gate and_gate_s_wallace_cska32_and_4_14(.a(a[4]), .b(b[14]), .out(s_wallace_cska32_and_4_14));
  and_gate and_gate_s_wallace_cska32_and_3_15(.a(a[3]), .b(b[15]), .out(s_wallace_cska32_and_3_15));
  fa fa_s_wallace_cska32_fa372_out(.a(s_wallace_cska32_fa371_or0[0]), .b(s_wallace_cska32_and_4_14[0]), .cin(s_wallace_cska32_and_3_15[0]), .fa_xor1(s_wallace_cska32_fa372_xor1), .fa_or0(s_wallace_cska32_fa372_or0));
  and_gate and_gate_s_wallace_cska32_and_5_14(.a(a[5]), .b(b[14]), .out(s_wallace_cska32_and_5_14));
  and_gate and_gate_s_wallace_cska32_and_4_15(.a(a[4]), .b(b[15]), .out(s_wallace_cska32_and_4_15));
  fa fa_s_wallace_cska32_fa373_out(.a(s_wallace_cska32_fa372_or0[0]), .b(s_wallace_cska32_and_5_14[0]), .cin(s_wallace_cska32_and_4_15[0]), .fa_xor1(s_wallace_cska32_fa373_xor1), .fa_or0(s_wallace_cska32_fa373_or0));
  and_gate and_gate_s_wallace_cska32_and_6_14(.a(a[6]), .b(b[14]), .out(s_wallace_cska32_and_6_14));
  and_gate and_gate_s_wallace_cska32_and_5_15(.a(a[5]), .b(b[15]), .out(s_wallace_cska32_and_5_15));
  fa fa_s_wallace_cska32_fa374_out(.a(s_wallace_cska32_fa373_or0[0]), .b(s_wallace_cska32_and_6_14[0]), .cin(s_wallace_cska32_and_5_15[0]), .fa_xor1(s_wallace_cska32_fa374_xor1), .fa_or0(s_wallace_cska32_fa374_or0));
  and_gate and_gate_s_wallace_cska32_and_7_14(.a(a[7]), .b(b[14]), .out(s_wallace_cska32_and_7_14));
  and_gate and_gate_s_wallace_cska32_and_6_15(.a(a[6]), .b(b[15]), .out(s_wallace_cska32_and_6_15));
  fa fa_s_wallace_cska32_fa375_out(.a(s_wallace_cska32_fa374_or0[0]), .b(s_wallace_cska32_and_7_14[0]), .cin(s_wallace_cska32_and_6_15[0]), .fa_xor1(s_wallace_cska32_fa375_xor1), .fa_or0(s_wallace_cska32_fa375_or0));
  and_gate and_gate_s_wallace_cska32_and_8_14(.a(a[8]), .b(b[14]), .out(s_wallace_cska32_and_8_14));
  and_gate and_gate_s_wallace_cska32_and_7_15(.a(a[7]), .b(b[15]), .out(s_wallace_cska32_and_7_15));
  fa fa_s_wallace_cska32_fa376_out(.a(s_wallace_cska32_fa375_or0[0]), .b(s_wallace_cska32_and_8_14[0]), .cin(s_wallace_cska32_and_7_15[0]), .fa_xor1(s_wallace_cska32_fa376_xor1), .fa_or0(s_wallace_cska32_fa376_or0));
  and_gate and_gate_s_wallace_cska32_and_9_14(.a(a[9]), .b(b[14]), .out(s_wallace_cska32_and_9_14));
  and_gate and_gate_s_wallace_cska32_and_8_15(.a(a[8]), .b(b[15]), .out(s_wallace_cska32_and_8_15));
  fa fa_s_wallace_cska32_fa377_out(.a(s_wallace_cska32_fa376_or0[0]), .b(s_wallace_cska32_and_9_14[0]), .cin(s_wallace_cska32_and_8_15[0]), .fa_xor1(s_wallace_cska32_fa377_xor1), .fa_or0(s_wallace_cska32_fa377_or0));
  and_gate and_gate_s_wallace_cska32_and_10_14(.a(a[10]), .b(b[14]), .out(s_wallace_cska32_and_10_14));
  and_gate and_gate_s_wallace_cska32_and_9_15(.a(a[9]), .b(b[15]), .out(s_wallace_cska32_and_9_15));
  fa fa_s_wallace_cska32_fa378_out(.a(s_wallace_cska32_fa377_or0[0]), .b(s_wallace_cska32_and_10_14[0]), .cin(s_wallace_cska32_and_9_15[0]), .fa_xor1(s_wallace_cska32_fa378_xor1), .fa_or0(s_wallace_cska32_fa378_or0));
  and_gate and_gate_s_wallace_cska32_and_11_14(.a(a[11]), .b(b[14]), .out(s_wallace_cska32_and_11_14));
  and_gate and_gate_s_wallace_cska32_and_10_15(.a(a[10]), .b(b[15]), .out(s_wallace_cska32_and_10_15));
  fa fa_s_wallace_cska32_fa379_out(.a(s_wallace_cska32_fa378_or0[0]), .b(s_wallace_cska32_and_11_14[0]), .cin(s_wallace_cska32_and_10_15[0]), .fa_xor1(s_wallace_cska32_fa379_xor1), .fa_or0(s_wallace_cska32_fa379_or0));
  and_gate and_gate_s_wallace_cska32_and_12_14(.a(a[12]), .b(b[14]), .out(s_wallace_cska32_and_12_14));
  and_gate and_gate_s_wallace_cska32_and_11_15(.a(a[11]), .b(b[15]), .out(s_wallace_cska32_and_11_15));
  fa fa_s_wallace_cska32_fa380_out(.a(s_wallace_cska32_fa379_or0[0]), .b(s_wallace_cska32_and_12_14[0]), .cin(s_wallace_cska32_and_11_15[0]), .fa_xor1(s_wallace_cska32_fa380_xor1), .fa_or0(s_wallace_cska32_fa380_or0));
  and_gate and_gate_s_wallace_cska32_and_13_14(.a(a[13]), .b(b[14]), .out(s_wallace_cska32_and_13_14));
  and_gate and_gate_s_wallace_cska32_and_12_15(.a(a[12]), .b(b[15]), .out(s_wallace_cska32_and_12_15));
  fa fa_s_wallace_cska32_fa381_out(.a(s_wallace_cska32_fa380_or0[0]), .b(s_wallace_cska32_and_13_14[0]), .cin(s_wallace_cska32_and_12_15[0]), .fa_xor1(s_wallace_cska32_fa381_xor1), .fa_or0(s_wallace_cska32_fa381_or0));
  and_gate and_gate_s_wallace_cska32_and_14_14(.a(a[14]), .b(b[14]), .out(s_wallace_cska32_and_14_14));
  and_gate and_gate_s_wallace_cska32_and_13_15(.a(a[13]), .b(b[15]), .out(s_wallace_cska32_and_13_15));
  fa fa_s_wallace_cska32_fa382_out(.a(s_wallace_cska32_fa381_or0[0]), .b(s_wallace_cska32_and_14_14[0]), .cin(s_wallace_cska32_and_13_15[0]), .fa_xor1(s_wallace_cska32_fa382_xor1), .fa_or0(s_wallace_cska32_fa382_or0));
  and_gate and_gate_s_wallace_cska32_and_15_14(.a(a[15]), .b(b[14]), .out(s_wallace_cska32_and_15_14));
  and_gate and_gate_s_wallace_cska32_and_14_15(.a(a[14]), .b(b[15]), .out(s_wallace_cska32_and_14_15));
  fa fa_s_wallace_cska32_fa383_out(.a(s_wallace_cska32_fa382_or0[0]), .b(s_wallace_cska32_and_15_14[0]), .cin(s_wallace_cska32_and_14_15[0]), .fa_xor1(s_wallace_cska32_fa383_xor1), .fa_or0(s_wallace_cska32_fa383_or0));
  and_gate and_gate_s_wallace_cska32_and_16_14(.a(a[16]), .b(b[14]), .out(s_wallace_cska32_and_16_14));
  and_gate and_gate_s_wallace_cska32_and_15_15(.a(a[15]), .b(b[15]), .out(s_wallace_cska32_and_15_15));
  fa fa_s_wallace_cska32_fa384_out(.a(s_wallace_cska32_fa383_or0[0]), .b(s_wallace_cska32_and_16_14[0]), .cin(s_wallace_cska32_and_15_15[0]), .fa_xor1(s_wallace_cska32_fa384_xor1), .fa_or0(s_wallace_cska32_fa384_or0));
  and_gate and_gate_s_wallace_cska32_and_17_14(.a(a[17]), .b(b[14]), .out(s_wallace_cska32_and_17_14));
  and_gate and_gate_s_wallace_cska32_and_16_15(.a(a[16]), .b(b[15]), .out(s_wallace_cska32_and_16_15));
  fa fa_s_wallace_cska32_fa385_out(.a(s_wallace_cska32_fa384_or0[0]), .b(s_wallace_cska32_and_17_14[0]), .cin(s_wallace_cska32_and_16_15[0]), .fa_xor1(s_wallace_cska32_fa385_xor1), .fa_or0(s_wallace_cska32_fa385_or0));
  and_gate and_gate_s_wallace_cska32_and_18_14(.a(a[18]), .b(b[14]), .out(s_wallace_cska32_and_18_14));
  and_gate and_gate_s_wallace_cska32_and_17_15(.a(a[17]), .b(b[15]), .out(s_wallace_cska32_and_17_15));
  fa fa_s_wallace_cska32_fa386_out(.a(s_wallace_cska32_fa385_or0[0]), .b(s_wallace_cska32_and_18_14[0]), .cin(s_wallace_cska32_and_17_15[0]), .fa_xor1(s_wallace_cska32_fa386_xor1), .fa_or0(s_wallace_cska32_fa386_or0));
  and_gate and_gate_s_wallace_cska32_and_17_16(.a(a[17]), .b(b[16]), .out(s_wallace_cska32_and_17_16));
  and_gate and_gate_s_wallace_cska32_and_16_17(.a(a[16]), .b(b[17]), .out(s_wallace_cska32_and_16_17));
  fa fa_s_wallace_cska32_fa387_out(.a(s_wallace_cska32_fa386_or0[0]), .b(s_wallace_cska32_and_17_16[0]), .cin(s_wallace_cska32_and_16_17[0]), .fa_xor1(s_wallace_cska32_fa387_xor1), .fa_or0(s_wallace_cska32_fa387_or0));
  and_gate and_gate_s_wallace_cska32_and_17_17(.a(a[17]), .b(b[17]), .out(s_wallace_cska32_and_17_17));
  and_gate and_gate_s_wallace_cska32_and_16_18(.a(a[16]), .b(b[18]), .out(s_wallace_cska32_and_16_18));
  fa fa_s_wallace_cska32_fa388_out(.a(s_wallace_cska32_fa387_or0[0]), .b(s_wallace_cska32_and_17_17[0]), .cin(s_wallace_cska32_and_16_18[0]), .fa_xor1(s_wallace_cska32_fa388_xor1), .fa_or0(s_wallace_cska32_fa388_or0));
  and_gate and_gate_s_wallace_cska32_and_17_18(.a(a[17]), .b(b[18]), .out(s_wallace_cska32_and_17_18));
  and_gate and_gate_s_wallace_cska32_and_16_19(.a(a[16]), .b(b[19]), .out(s_wallace_cska32_and_16_19));
  fa fa_s_wallace_cska32_fa389_out(.a(s_wallace_cska32_fa388_or0[0]), .b(s_wallace_cska32_and_17_18[0]), .cin(s_wallace_cska32_and_16_19[0]), .fa_xor1(s_wallace_cska32_fa389_xor1), .fa_or0(s_wallace_cska32_fa389_or0));
  and_gate and_gate_s_wallace_cska32_and_17_19(.a(a[17]), .b(b[19]), .out(s_wallace_cska32_and_17_19));
  and_gate and_gate_s_wallace_cska32_and_16_20(.a(a[16]), .b(b[20]), .out(s_wallace_cska32_and_16_20));
  fa fa_s_wallace_cska32_fa390_out(.a(s_wallace_cska32_fa389_or0[0]), .b(s_wallace_cska32_and_17_19[0]), .cin(s_wallace_cska32_and_16_20[0]), .fa_xor1(s_wallace_cska32_fa390_xor1), .fa_or0(s_wallace_cska32_fa390_or0));
  and_gate and_gate_s_wallace_cska32_and_17_20(.a(a[17]), .b(b[20]), .out(s_wallace_cska32_and_17_20));
  and_gate and_gate_s_wallace_cska32_and_16_21(.a(a[16]), .b(b[21]), .out(s_wallace_cska32_and_16_21));
  fa fa_s_wallace_cska32_fa391_out(.a(s_wallace_cska32_fa390_or0[0]), .b(s_wallace_cska32_and_17_20[0]), .cin(s_wallace_cska32_and_16_21[0]), .fa_xor1(s_wallace_cska32_fa391_xor1), .fa_or0(s_wallace_cska32_fa391_or0));
  and_gate and_gate_s_wallace_cska32_and_17_21(.a(a[17]), .b(b[21]), .out(s_wallace_cska32_and_17_21));
  and_gate and_gate_s_wallace_cska32_and_16_22(.a(a[16]), .b(b[22]), .out(s_wallace_cska32_and_16_22));
  fa fa_s_wallace_cska32_fa392_out(.a(s_wallace_cska32_fa391_or0[0]), .b(s_wallace_cska32_and_17_21[0]), .cin(s_wallace_cska32_and_16_22[0]), .fa_xor1(s_wallace_cska32_fa392_xor1), .fa_or0(s_wallace_cska32_fa392_or0));
  and_gate and_gate_s_wallace_cska32_and_17_22(.a(a[17]), .b(b[22]), .out(s_wallace_cska32_and_17_22));
  and_gate and_gate_s_wallace_cska32_and_16_23(.a(a[16]), .b(b[23]), .out(s_wallace_cska32_and_16_23));
  fa fa_s_wallace_cska32_fa393_out(.a(s_wallace_cska32_fa392_or0[0]), .b(s_wallace_cska32_and_17_22[0]), .cin(s_wallace_cska32_and_16_23[0]), .fa_xor1(s_wallace_cska32_fa393_xor1), .fa_or0(s_wallace_cska32_fa393_or0));
  and_gate and_gate_s_wallace_cska32_and_17_23(.a(a[17]), .b(b[23]), .out(s_wallace_cska32_and_17_23));
  and_gate and_gate_s_wallace_cska32_and_16_24(.a(a[16]), .b(b[24]), .out(s_wallace_cska32_and_16_24));
  fa fa_s_wallace_cska32_fa394_out(.a(s_wallace_cska32_fa393_or0[0]), .b(s_wallace_cska32_and_17_23[0]), .cin(s_wallace_cska32_and_16_24[0]), .fa_xor1(s_wallace_cska32_fa394_xor1), .fa_or0(s_wallace_cska32_fa394_or0));
  and_gate and_gate_s_wallace_cska32_and_17_24(.a(a[17]), .b(b[24]), .out(s_wallace_cska32_and_17_24));
  and_gate and_gate_s_wallace_cska32_and_16_25(.a(a[16]), .b(b[25]), .out(s_wallace_cska32_and_16_25));
  fa fa_s_wallace_cska32_fa395_out(.a(s_wallace_cska32_fa394_or0[0]), .b(s_wallace_cska32_and_17_24[0]), .cin(s_wallace_cska32_and_16_25[0]), .fa_xor1(s_wallace_cska32_fa395_xor1), .fa_or0(s_wallace_cska32_fa395_or0));
  and_gate and_gate_s_wallace_cska32_and_17_25(.a(a[17]), .b(b[25]), .out(s_wallace_cska32_and_17_25));
  and_gate and_gate_s_wallace_cska32_and_16_26(.a(a[16]), .b(b[26]), .out(s_wallace_cska32_and_16_26));
  fa fa_s_wallace_cska32_fa396_out(.a(s_wallace_cska32_fa395_or0[0]), .b(s_wallace_cska32_and_17_25[0]), .cin(s_wallace_cska32_and_16_26[0]), .fa_xor1(s_wallace_cska32_fa396_xor1), .fa_or0(s_wallace_cska32_fa396_or0));
  and_gate and_gate_s_wallace_cska32_and_17_26(.a(a[17]), .b(b[26]), .out(s_wallace_cska32_and_17_26));
  and_gate and_gate_s_wallace_cska32_and_16_27(.a(a[16]), .b(b[27]), .out(s_wallace_cska32_and_16_27));
  fa fa_s_wallace_cska32_fa397_out(.a(s_wallace_cska32_fa396_or0[0]), .b(s_wallace_cska32_and_17_26[0]), .cin(s_wallace_cska32_and_16_27[0]), .fa_xor1(s_wallace_cska32_fa397_xor1), .fa_or0(s_wallace_cska32_fa397_or0));
  and_gate and_gate_s_wallace_cska32_and_17_27(.a(a[17]), .b(b[27]), .out(s_wallace_cska32_and_17_27));
  and_gate and_gate_s_wallace_cska32_and_16_28(.a(a[16]), .b(b[28]), .out(s_wallace_cska32_and_16_28));
  fa fa_s_wallace_cska32_fa398_out(.a(s_wallace_cska32_fa397_or0[0]), .b(s_wallace_cska32_and_17_27[0]), .cin(s_wallace_cska32_and_16_28[0]), .fa_xor1(s_wallace_cska32_fa398_xor1), .fa_or0(s_wallace_cska32_fa398_or0));
  and_gate and_gate_s_wallace_cska32_and_17_28(.a(a[17]), .b(b[28]), .out(s_wallace_cska32_and_17_28));
  and_gate and_gate_s_wallace_cska32_and_16_29(.a(a[16]), .b(b[29]), .out(s_wallace_cska32_and_16_29));
  fa fa_s_wallace_cska32_fa399_out(.a(s_wallace_cska32_fa398_or0[0]), .b(s_wallace_cska32_and_17_28[0]), .cin(s_wallace_cska32_and_16_29[0]), .fa_xor1(s_wallace_cska32_fa399_xor1), .fa_or0(s_wallace_cska32_fa399_or0));
  and_gate and_gate_s_wallace_cska32_and_17_29(.a(a[17]), .b(b[29]), .out(s_wallace_cska32_and_17_29));
  and_gate and_gate_s_wallace_cska32_and_16_30(.a(a[16]), .b(b[30]), .out(s_wallace_cska32_and_16_30));
  fa fa_s_wallace_cska32_fa400_out(.a(s_wallace_cska32_fa399_or0[0]), .b(s_wallace_cska32_and_17_29[0]), .cin(s_wallace_cska32_and_16_30[0]), .fa_xor1(s_wallace_cska32_fa400_xor1), .fa_or0(s_wallace_cska32_fa400_or0));
  and_gate and_gate_s_wallace_cska32_and_17_30(.a(a[17]), .b(b[30]), .out(s_wallace_cska32_and_17_30));
  nand_gate nand_gate_s_wallace_cska32_nand_16_31(.a(a[16]), .b(b[31]), .out(s_wallace_cska32_nand_16_31));
  fa fa_s_wallace_cska32_fa401_out(.a(s_wallace_cska32_fa400_or0[0]), .b(s_wallace_cska32_and_17_30[0]), .cin(s_wallace_cska32_nand_16_31[0]), .fa_xor1(s_wallace_cska32_fa401_xor1), .fa_or0(s_wallace_cska32_fa401_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_17_31(.a(a[17]), .b(b[31]), .out(s_wallace_cska32_nand_17_31));
  fa fa_s_wallace_cska32_fa402_out(.a(s_wallace_cska32_fa401_or0[0]), .b(s_wallace_cska32_nand_17_31[0]), .cin(s_wallace_cska32_fa45_xor1[0]), .fa_xor1(s_wallace_cska32_fa402_xor1), .fa_or0(s_wallace_cska32_fa402_or0));
  fa fa_s_wallace_cska32_fa403_out(.a(s_wallace_cska32_fa402_or0[0]), .b(s_wallace_cska32_fa46_xor1[0]), .cin(s_wallace_cska32_fa103_xor1[0]), .fa_xor1(s_wallace_cska32_fa403_xor1), .fa_or0(s_wallace_cska32_fa403_or0));
  fa fa_s_wallace_cska32_fa404_out(.a(s_wallace_cska32_fa403_or0[0]), .b(s_wallace_cska32_fa104_xor1[0]), .cin(s_wallace_cska32_fa159_xor1[0]), .fa_xor1(s_wallace_cska32_fa404_xor1), .fa_or0(s_wallace_cska32_fa404_or0));
  fa fa_s_wallace_cska32_fa405_out(.a(s_wallace_cska32_fa404_or0[0]), .b(s_wallace_cska32_fa160_xor1[0]), .cin(s_wallace_cska32_fa213_xor1[0]), .fa_xor1(s_wallace_cska32_fa405_xor1), .fa_or0(s_wallace_cska32_fa405_or0));
  fa fa_s_wallace_cska32_fa406_out(.a(s_wallace_cska32_fa405_or0[0]), .b(s_wallace_cska32_fa214_xor1[0]), .cin(s_wallace_cska32_fa265_xor1[0]), .fa_xor1(s_wallace_cska32_fa406_xor1), .fa_or0(s_wallace_cska32_fa406_or0));
  fa fa_s_wallace_cska32_fa407_out(.a(s_wallace_cska32_fa406_or0[0]), .b(s_wallace_cska32_fa266_xor1[0]), .cin(s_wallace_cska32_fa315_xor1[0]), .fa_xor1(s_wallace_cska32_fa407_xor1), .fa_or0(s_wallace_cska32_fa407_or0));
  ha ha_s_wallace_cska32_ha8_out(.a(s_wallace_cska32_fa272_xor1[0]), .b(s_wallace_cska32_fa319_xor1[0]), .ha_xor0(s_wallace_cska32_ha8_xor0), .ha_and0(s_wallace_cska32_ha8_and0));
  fa fa_s_wallace_cska32_fa408_out(.a(s_wallace_cska32_ha8_and0[0]), .b(s_wallace_cska32_fa224_xor1[0]), .cin(s_wallace_cska32_fa273_xor1[0]), .fa_xor1(s_wallace_cska32_fa408_xor1), .fa_or0(s_wallace_cska32_fa408_or0));
  fa fa_s_wallace_cska32_fa409_out(.a(s_wallace_cska32_fa408_or0[0]), .b(s_wallace_cska32_fa174_xor1[0]), .cin(s_wallace_cska32_fa225_xor1[0]), .fa_xor1(s_wallace_cska32_fa409_xor1), .fa_or0(s_wallace_cska32_fa409_or0));
  fa fa_s_wallace_cska32_fa410_out(.a(s_wallace_cska32_fa409_or0[0]), .b(s_wallace_cska32_fa122_xor1[0]), .cin(s_wallace_cska32_fa175_xor1[0]), .fa_xor1(s_wallace_cska32_fa410_xor1), .fa_or0(s_wallace_cska32_fa410_or0));
  fa fa_s_wallace_cska32_fa411_out(.a(s_wallace_cska32_fa410_or0[0]), .b(s_wallace_cska32_fa68_xor1[0]), .cin(s_wallace_cska32_fa123_xor1[0]), .fa_xor1(s_wallace_cska32_fa411_xor1), .fa_or0(s_wallace_cska32_fa411_or0));
  fa fa_s_wallace_cska32_fa412_out(.a(s_wallace_cska32_fa411_or0[0]), .b(s_wallace_cska32_fa12_xor1[0]), .cin(s_wallace_cska32_fa69_xor1[0]), .fa_xor1(s_wallace_cska32_fa412_xor1), .fa_or0(s_wallace_cska32_fa412_or0));
  and_gate and_gate_s_wallace_cska32_and_0_16(.a(a[0]), .b(b[16]), .out(s_wallace_cska32_and_0_16));
  fa fa_s_wallace_cska32_fa413_out(.a(s_wallace_cska32_fa412_or0[0]), .b(s_wallace_cska32_and_0_16[0]), .cin(s_wallace_cska32_fa13_xor1[0]), .fa_xor1(s_wallace_cska32_fa413_xor1), .fa_or0(s_wallace_cska32_fa413_or0));
  and_gate and_gate_s_wallace_cska32_and_1_16(.a(a[1]), .b(b[16]), .out(s_wallace_cska32_and_1_16));
  and_gate and_gate_s_wallace_cska32_and_0_17(.a(a[0]), .b(b[17]), .out(s_wallace_cska32_and_0_17));
  fa fa_s_wallace_cska32_fa414_out(.a(s_wallace_cska32_fa413_or0[0]), .b(s_wallace_cska32_and_1_16[0]), .cin(s_wallace_cska32_and_0_17[0]), .fa_xor1(s_wallace_cska32_fa414_xor1), .fa_or0(s_wallace_cska32_fa414_or0));
  and_gate and_gate_s_wallace_cska32_and_2_16(.a(a[2]), .b(b[16]), .out(s_wallace_cska32_and_2_16));
  and_gate and_gate_s_wallace_cska32_and_1_17(.a(a[1]), .b(b[17]), .out(s_wallace_cska32_and_1_17));
  fa fa_s_wallace_cska32_fa415_out(.a(s_wallace_cska32_fa414_or0[0]), .b(s_wallace_cska32_and_2_16[0]), .cin(s_wallace_cska32_and_1_17[0]), .fa_xor1(s_wallace_cska32_fa415_xor1), .fa_or0(s_wallace_cska32_fa415_or0));
  and_gate and_gate_s_wallace_cska32_and_3_16(.a(a[3]), .b(b[16]), .out(s_wallace_cska32_and_3_16));
  and_gate and_gate_s_wallace_cska32_and_2_17(.a(a[2]), .b(b[17]), .out(s_wallace_cska32_and_2_17));
  fa fa_s_wallace_cska32_fa416_out(.a(s_wallace_cska32_fa415_or0[0]), .b(s_wallace_cska32_and_3_16[0]), .cin(s_wallace_cska32_and_2_17[0]), .fa_xor1(s_wallace_cska32_fa416_xor1), .fa_or0(s_wallace_cska32_fa416_or0));
  and_gate and_gate_s_wallace_cska32_and_4_16(.a(a[4]), .b(b[16]), .out(s_wallace_cska32_and_4_16));
  and_gate and_gate_s_wallace_cska32_and_3_17(.a(a[3]), .b(b[17]), .out(s_wallace_cska32_and_3_17));
  fa fa_s_wallace_cska32_fa417_out(.a(s_wallace_cska32_fa416_or0[0]), .b(s_wallace_cska32_and_4_16[0]), .cin(s_wallace_cska32_and_3_17[0]), .fa_xor1(s_wallace_cska32_fa417_xor1), .fa_or0(s_wallace_cska32_fa417_or0));
  and_gate and_gate_s_wallace_cska32_and_5_16(.a(a[5]), .b(b[16]), .out(s_wallace_cska32_and_5_16));
  and_gate and_gate_s_wallace_cska32_and_4_17(.a(a[4]), .b(b[17]), .out(s_wallace_cska32_and_4_17));
  fa fa_s_wallace_cska32_fa418_out(.a(s_wallace_cska32_fa417_or0[0]), .b(s_wallace_cska32_and_5_16[0]), .cin(s_wallace_cska32_and_4_17[0]), .fa_xor1(s_wallace_cska32_fa418_xor1), .fa_or0(s_wallace_cska32_fa418_or0));
  and_gate and_gate_s_wallace_cska32_and_6_16(.a(a[6]), .b(b[16]), .out(s_wallace_cska32_and_6_16));
  and_gate and_gate_s_wallace_cska32_and_5_17(.a(a[5]), .b(b[17]), .out(s_wallace_cska32_and_5_17));
  fa fa_s_wallace_cska32_fa419_out(.a(s_wallace_cska32_fa418_or0[0]), .b(s_wallace_cska32_and_6_16[0]), .cin(s_wallace_cska32_and_5_17[0]), .fa_xor1(s_wallace_cska32_fa419_xor1), .fa_or0(s_wallace_cska32_fa419_or0));
  and_gate and_gate_s_wallace_cska32_and_7_16(.a(a[7]), .b(b[16]), .out(s_wallace_cska32_and_7_16));
  and_gate and_gate_s_wallace_cska32_and_6_17(.a(a[6]), .b(b[17]), .out(s_wallace_cska32_and_6_17));
  fa fa_s_wallace_cska32_fa420_out(.a(s_wallace_cska32_fa419_or0[0]), .b(s_wallace_cska32_and_7_16[0]), .cin(s_wallace_cska32_and_6_17[0]), .fa_xor1(s_wallace_cska32_fa420_xor1), .fa_or0(s_wallace_cska32_fa420_or0));
  and_gate and_gate_s_wallace_cska32_and_8_16(.a(a[8]), .b(b[16]), .out(s_wallace_cska32_and_8_16));
  and_gate and_gate_s_wallace_cska32_and_7_17(.a(a[7]), .b(b[17]), .out(s_wallace_cska32_and_7_17));
  fa fa_s_wallace_cska32_fa421_out(.a(s_wallace_cska32_fa420_or0[0]), .b(s_wallace_cska32_and_8_16[0]), .cin(s_wallace_cska32_and_7_17[0]), .fa_xor1(s_wallace_cska32_fa421_xor1), .fa_or0(s_wallace_cska32_fa421_or0));
  and_gate and_gate_s_wallace_cska32_and_9_16(.a(a[9]), .b(b[16]), .out(s_wallace_cska32_and_9_16));
  and_gate and_gate_s_wallace_cska32_and_8_17(.a(a[8]), .b(b[17]), .out(s_wallace_cska32_and_8_17));
  fa fa_s_wallace_cska32_fa422_out(.a(s_wallace_cska32_fa421_or0[0]), .b(s_wallace_cska32_and_9_16[0]), .cin(s_wallace_cska32_and_8_17[0]), .fa_xor1(s_wallace_cska32_fa422_xor1), .fa_or0(s_wallace_cska32_fa422_or0));
  and_gate and_gate_s_wallace_cska32_and_10_16(.a(a[10]), .b(b[16]), .out(s_wallace_cska32_and_10_16));
  and_gate and_gate_s_wallace_cska32_and_9_17(.a(a[9]), .b(b[17]), .out(s_wallace_cska32_and_9_17));
  fa fa_s_wallace_cska32_fa423_out(.a(s_wallace_cska32_fa422_or0[0]), .b(s_wallace_cska32_and_10_16[0]), .cin(s_wallace_cska32_and_9_17[0]), .fa_xor1(s_wallace_cska32_fa423_xor1), .fa_or0(s_wallace_cska32_fa423_or0));
  and_gate and_gate_s_wallace_cska32_and_11_16(.a(a[11]), .b(b[16]), .out(s_wallace_cska32_and_11_16));
  and_gate and_gate_s_wallace_cska32_and_10_17(.a(a[10]), .b(b[17]), .out(s_wallace_cska32_and_10_17));
  fa fa_s_wallace_cska32_fa424_out(.a(s_wallace_cska32_fa423_or0[0]), .b(s_wallace_cska32_and_11_16[0]), .cin(s_wallace_cska32_and_10_17[0]), .fa_xor1(s_wallace_cska32_fa424_xor1), .fa_or0(s_wallace_cska32_fa424_or0));
  and_gate and_gate_s_wallace_cska32_and_12_16(.a(a[12]), .b(b[16]), .out(s_wallace_cska32_and_12_16));
  and_gate and_gate_s_wallace_cska32_and_11_17(.a(a[11]), .b(b[17]), .out(s_wallace_cska32_and_11_17));
  fa fa_s_wallace_cska32_fa425_out(.a(s_wallace_cska32_fa424_or0[0]), .b(s_wallace_cska32_and_12_16[0]), .cin(s_wallace_cska32_and_11_17[0]), .fa_xor1(s_wallace_cska32_fa425_xor1), .fa_or0(s_wallace_cska32_fa425_or0));
  and_gate and_gate_s_wallace_cska32_and_13_16(.a(a[13]), .b(b[16]), .out(s_wallace_cska32_and_13_16));
  and_gate and_gate_s_wallace_cska32_and_12_17(.a(a[12]), .b(b[17]), .out(s_wallace_cska32_and_12_17));
  fa fa_s_wallace_cska32_fa426_out(.a(s_wallace_cska32_fa425_or0[0]), .b(s_wallace_cska32_and_13_16[0]), .cin(s_wallace_cska32_and_12_17[0]), .fa_xor1(s_wallace_cska32_fa426_xor1), .fa_or0(s_wallace_cska32_fa426_or0));
  and_gate and_gate_s_wallace_cska32_and_14_16(.a(a[14]), .b(b[16]), .out(s_wallace_cska32_and_14_16));
  and_gate and_gate_s_wallace_cska32_and_13_17(.a(a[13]), .b(b[17]), .out(s_wallace_cska32_and_13_17));
  fa fa_s_wallace_cska32_fa427_out(.a(s_wallace_cska32_fa426_or0[0]), .b(s_wallace_cska32_and_14_16[0]), .cin(s_wallace_cska32_and_13_17[0]), .fa_xor1(s_wallace_cska32_fa427_xor1), .fa_or0(s_wallace_cska32_fa427_or0));
  and_gate and_gate_s_wallace_cska32_and_15_16(.a(a[15]), .b(b[16]), .out(s_wallace_cska32_and_15_16));
  and_gate and_gate_s_wallace_cska32_and_14_17(.a(a[14]), .b(b[17]), .out(s_wallace_cska32_and_14_17));
  fa fa_s_wallace_cska32_fa428_out(.a(s_wallace_cska32_fa427_or0[0]), .b(s_wallace_cska32_and_15_16[0]), .cin(s_wallace_cska32_and_14_17[0]), .fa_xor1(s_wallace_cska32_fa428_xor1), .fa_or0(s_wallace_cska32_fa428_or0));
  and_gate and_gate_s_wallace_cska32_and_16_16(.a(a[16]), .b(b[16]), .out(s_wallace_cska32_and_16_16));
  and_gate and_gate_s_wallace_cska32_and_15_17(.a(a[15]), .b(b[17]), .out(s_wallace_cska32_and_15_17));
  fa fa_s_wallace_cska32_fa429_out(.a(s_wallace_cska32_fa428_or0[0]), .b(s_wallace_cska32_and_16_16[0]), .cin(s_wallace_cska32_and_15_17[0]), .fa_xor1(s_wallace_cska32_fa429_xor1), .fa_or0(s_wallace_cska32_fa429_or0));
  and_gate and_gate_s_wallace_cska32_and_15_18(.a(a[15]), .b(b[18]), .out(s_wallace_cska32_and_15_18));
  and_gate and_gate_s_wallace_cska32_and_14_19(.a(a[14]), .b(b[19]), .out(s_wallace_cska32_and_14_19));
  fa fa_s_wallace_cska32_fa430_out(.a(s_wallace_cska32_fa429_or0[0]), .b(s_wallace_cska32_and_15_18[0]), .cin(s_wallace_cska32_and_14_19[0]), .fa_xor1(s_wallace_cska32_fa430_xor1), .fa_or0(s_wallace_cska32_fa430_or0));
  and_gate and_gate_s_wallace_cska32_and_15_19(.a(a[15]), .b(b[19]), .out(s_wallace_cska32_and_15_19));
  and_gate and_gate_s_wallace_cska32_and_14_20(.a(a[14]), .b(b[20]), .out(s_wallace_cska32_and_14_20));
  fa fa_s_wallace_cska32_fa431_out(.a(s_wallace_cska32_fa430_or0[0]), .b(s_wallace_cska32_and_15_19[0]), .cin(s_wallace_cska32_and_14_20[0]), .fa_xor1(s_wallace_cska32_fa431_xor1), .fa_or0(s_wallace_cska32_fa431_or0));
  and_gate and_gate_s_wallace_cska32_and_15_20(.a(a[15]), .b(b[20]), .out(s_wallace_cska32_and_15_20));
  and_gate and_gate_s_wallace_cska32_and_14_21(.a(a[14]), .b(b[21]), .out(s_wallace_cska32_and_14_21));
  fa fa_s_wallace_cska32_fa432_out(.a(s_wallace_cska32_fa431_or0[0]), .b(s_wallace_cska32_and_15_20[0]), .cin(s_wallace_cska32_and_14_21[0]), .fa_xor1(s_wallace_cska32_fa432_xor1), .fa_or0(s_wallace_cska32_fa432_or0));
  and_gate and_gate_s_wallace_cska32_and_15_21(.a(a[15]), .b(b[21]), .out(s_wallace_cska32_and_15_21));
  and_gate and_gate_s_wallace_cska32_and_14_22(.a(a[14]), .b(b[22]), .out(s_wallace_cska32_and_14_22));
  fa fa_s_wallace_cska32_fa433_out(.a(s_wallace_cska32_fa432_or0[0]), .b(s_wallace_cska32_and_15_21[0]), .cin(s_wallace_cska32_and_14_22[0]), .fa_xor1(s_wallace_cska32_fa433_xor1), .fa_or0(s_wallace_cska32_fa433_or0));
  and_gate and_gate_s_wallace_cska32_and_15_22(.a(a[15]), .b(b[22]), .out(s_wallace_cska32_and_15_22));
  and_gate and_gate_s_wallace_cska32_and_14_23(.a(a[14]), .b(b[23]), .out(s_wallace_cska32_and_14_23));
  fa fa_s_wallace_cska32_fa434_out(.a(s_wallace_cska32_fa433_or0[0]), .b(s_wallace_cska32_and_15_22[0]), .cin(s_wallace_cska32_and_14_23[0]), .fa_xor1(s_wallace_cska32_fa434_xor1), .fa_or0(s_wallace_cska32_fa434_or0));
  and_gate and_gate_s_wallace_cska32_and_15_23(.a(a[15]), .b(b[23]), .out(s_wallace_cska32_and_15_23));
  and_gate and_gate_s_wallace_cska32_and_14_24(.a(a[14]), .b(b[24]), .out(s_wallace_cska32_and_14_24));
  fa fa_s_wallace_cska32_fa435_out(.a(s_wallace_cska32_fa434_or0[0]), .b(s_wallace_cska32_and_15_23[0]), .cin(s_wallace_cska32_and_14_24[0]), .fa_xor1(s_wallace_cska32_fa435_xor1), .fa_or0(s_wallace_cska32_fa435_or0));
  and_gate and_gate_s_wallace_cska32_and_15_24(.a(a[15]), .b(b[24]), .out(s_wallace_cska32_and_15_24));
  and_gate and_gate_s_wallace_cska32_and_14_25(.a(a[14]), .b(b[25]), .out(s_wallace_cska32_and_14_25));
  fa fa_s_wallace_cska32_fa436_out(.a(s_wallace_cska32_fa435_or0[0]), .b(s_wallace_cska32_and_15_24[0]), .cin(s_wallace_cska32_and_14_25[0]), .fa_xor1(s_wallace_cska32_fa436_xor1), .fa_or0(s_wallace_cska32_fa436_or0));
  and_gate and_gate_s_wallace_cska32_and_15_25(.a(a[15]), .b(b[25]), .out(s_wallace_cska32_and_15_25));
  and_gate and_gate_s_wallace_cska32_and_14_26(.a(a[14]), .b(b[26]), .out(s_wallace_cska32_and_14_26));
  fa fa_s_wallace_cska32_fa437_out(.a(s_wallace_cska32_fa436_or0[0]), .b(s_wallace_cska32_and_15_25[0]), .cin(s_wallace_cska32_and_14_26[0]), .fa_xor1(s_wallace_cska32_fa437_xor1), .fa_or0(s_wallace_cska32_fa437_or0));
  and_gate and_gate_s_wallace_cska32_and_15_26(.a(a[15]), .b(b[26]), .out(s_wallace_cska32_and_15_26));
  and_gate and_gate_s_wallace_cska32_and_14_27(.a(a[14]), .b(b[27]), .out(s_wallace_cska32_and_14_27));
  fa fa_s_wallace_cska32_fa438_out(.a(s_wallace_cska32_fa437_or0[0]), .b(s_wallace_cska32_and_15_26[0]), .cin(s_wallace_cska32_and_14_27[0]), .fa_xor1(s_wallace_cska32_fa438_xor1), .fa_or0(s_wallace_cska32_fa438_or0));
  and_gate and_gate_s_wallace_cska32_and_15_27(.a(a[15]), .b(b[27]), .out(s_wallace_cska32_and_15_27));
  and_gate and_gate_s_wallace_cska32_and_14_28(.a(a[14]), .b(b[28]), .out(s_wallace_cska32_and_14_28));
  fa fa_s_wallace_cska32_fa439_out(.a(s_wallace_cska32_fa438_or0[0]), .b(s_wallace_cska32_and_15_27[0]), .cin(s_wallace_cska32_and_14_28[0]), .fa_xor1(s_wallace_cska32_fa439_xor1), .fa_or0(s_wallace_cska32_fa439_or0));
  and_gate and_gate_s_wallace_cska32_and_15_28(.a(a[15]), .b(b[28]), .out(s_wallace_cska32_and_15_28));
  and_gate and_gate_s_wallace_cska32_and_14_29(.a(a[14]), .b(b[29]), .out(s_wallace_cska32_and_14_29));
  fa fa_s_wallace_cska32_fa440_out(.a(s_wallace_cska32_fa439_or0[0]), .b(s_wallace_cska32_and_15_28[0]), .cin(s_wallace_cska32_and_14_29[0]), .fa_xor1(s_wallace_cska32_fa440_xor1), .fa_or0(s_wallace_cska32_fa440_or0));
  and_gate and_gate_s_wallace_cska32_and_15_29(.a(a[15]), .b(b[29]), .out(s_wallace_cska32_and_15_29));
  and_gate and_gate_s_wallace_cska32_and_14_30(.a(a[14]), .b(b[30]), .out(s_wallace_cska32_and_14_30));
  fa fa_s_wallace_cska32_fa441_out(.a(s_wallace_cska32_fa440_or0[0]), .b(s_wallace_cska32_and_15_29[0]), .cin(s_wallace_cska32_and_14_30[0]), .fa_xor1(s_wallace_cska32_fa441_xor1), .fa_or0(s_wallace_cska32_fa441_or0));
  and_gate and_gate_s_wallace_cska32_and_15_30(.a(a[15]), .b(b[30]), .out(s_wallace_cska32_and_15_30));
  nand_gate nand_gate_s_wallace_cska32_nand_14_31(.a(a[14]), .b(b[31]), .out(s_wallace_cska32_nand_14_31));
  fa fa_s_wallace_cska32_fa442_out(.a(s_wallace_cska32_fa441_or0[0]), .b(s_wallace_cska32_and_15_30[0]), .cin(s_wallace_cska32_nand_14_31[0]), .fa_xor1(s_wallace_cska32_fa442_xor1), .fa_or0(s_wallace_cska32_fa442_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_15_31(.a(a[15]), .b(b[31]), .out(s_wallace_cska32_nand_15_31));
  fa fa_s_wallace_cska32_fa443_out(.a(s_wallace_cska32_fa442_or0[0]), .b(s_wallace_cska32_nand_15_31[0]), .cin(s_wallace_cska32_fa43_xor1[0]), .fa_xor1(s_wallace_cska32_fa443_xor1), .fa_or0(s_wallace_cska32_fa443_or0));
  fa fa_s_wallace_cska32_fa444_out(.a(s_wallace_cska32_fa443_or0[0]), .b(s_wallace_cska32_fa44_xor1[0]), .cin(s_wallace_cska32_fa101_xor1[0]), .fa_xor1(s_wallace_cska32_fa444_xor1), .fa_or0(s_wallace_cska32_fa444_or0));
  fa fa_s_wallace_cska32_fa445_out(.a(s_wallace_cska32_fa444_or0[0]), .b(s_wallace_cska32_fa102_xor1[0]), .cin(s_wallace_cska32_fa157_xor1[0]), .fa_xor1(s_wallace_cska32_fa445_xor1), .fa_or0(s_wallace_cska32_fa445_or0));
  fa fa_s_wallace_cska32_fa446_out(.a(s_wallace_cska32_fa445_or0[0]), .b(s_wallace_cska32_fa158_xor1[0]), .cin(s_wallace_cska32_fa211_xor1[0]), .fa_xor1(s_wallace_cska32_fa446_xor1), .fa_or0(s_wallace_cska32_fa446_or0));
  fa fa_s_wallace_cska32_fa447_out(.a(s_wallace_cska32_fa446_or0[0]), .b(s_wallace_cska32_fa212_xor1[0]), .cin(s_wallace_cska32_fa263_xor1[0]), .fa_xor1(s_wallace_cska32_fa447_xor1), .fa_or0(s_wallace_cska32_fa447_or0));
  fa fa_s_wallace_cska32_fa448_out(.a(s_wallace_cska32_fa447_or0[0]), .b(s_wallace_cska32_fa264_xor1[0]), .cin(s_wallace_cska32_fa313_xor1[0]), .fa_xor1(s_wallace_cska32_fa448_xor1), .fa_or0(s_wallace_cska32_fa448_or0));
  fa fa_s_wallace_cska32_fa449_out(.a(s_wallace_cska32_fa448_or0[0]), .b(s_wallace_cska32_fa314_xor1[0]), .cin(s_wallace_cska32_fa361_xor1[0]), .fa_xor1(s_wallace_cska32_fa449_xor1), .fa_or0(s_wallace_cska32_fa449_or0));
  ha ha_s_wallace_cska32_ha9_out(.a(s_wallace_cska32_fa320_xor1[0]), .b(s_wallace_cska32_fa365_xor1[0]), .ha_xor0(s_wallace_cska32_ha9_xor0), .ha_and0(s_wallace_cska32_ha9_and0));
  fa fa_s_wallace_cska32_fa450_out(.a(s_wallace_cska32_ha9_and0[0]), .b(s_wallace_cska32_fa274_xor1[0]), .cin(s_wallace_cska32_fa321_xor1[0]), .fa_xor1(s_wallace_cska32_fa450_xor1), .fa_or0(s_wallace_cska32_fa450_or0));
  fa fa_s_wallace_cska32_fa451_out(.a(s_wallace_cska32_fa450_or0[0]), .b(s_wallace_cska32_fa226_xor1[0]), .cin(s_wallace_cska32_fa275_xor1[0]), .fa_xor1(s_wallace_cska32_fa451_xor1), .fa_or0(s_wallace_cska32_fa451_or0));
  fa fa_s_wallace_cska32_fa452_out(.a(s_wallace_cska32_fa451_or0[0]), .b(s_wallace_cska32_fa176_xor1[0]), .cin(s_wallace_cska32_fa227_xor1[0]), .fa_xor1(s_wallace_cska32_fa452_xor1), .fa_or0(s_wallace_cska32_fa452_or0));
  fa fa_s_wallace_cska32_fa453_out(.a(s_wallace_cska32_fa452_or0[0]), .b(s_wallace_cska32_fa124_xor1[0]), .cin(s_wallace_cska32_fa177_xor1[0]), .fa_xor1(s_wallace_cska32_fa453_xor1), .fa_or0(s_wallace_cska32_fa453_or0));
  fa fa_s_wallace_cska32_fa454_out(.a(s_wallace_cska32_fa453_or0[0]), .b(s_wallace_cska32_fa70_xor1[0]), .cin(s_wallace_cska32_fa125_xor1[0]), .fa_xor1(s_wallace_cska32_fa454_xor1), .fa_or0(s_wallace_cska32_fa454_or0));
  fa fa_s_wallace_cska32_fa455_out(.a(s_wallace_cska32_fa454_or0[0]), .b(s_wallace_cska32_fa14_xor1[0]), .cin(s_wallace_cska32_fa71_xor1[0]), .fa_xor1(s_wallace_cska32_fa455_xor1), .fa_or0(s_wallace_cska32_fa455_or0));
  and_gate and_gate_s_wallace_cska32_and_0_18(.a(a[0]), .b(b[18]), .out(s_wallace_cska32_and_0_18));
  fa fa_s_wallace_cska32_fa456_out(.a(s_wallace_cska32_fa455_or0[0]), .b(s_wallace_cska32_and_0_18[0]), .cin(s_wallace_cska32_fa15_xor1[0]), .fa_xor1(s_wallace_cska32_fa456_xor1), .fa_or0(s_wallace_cska32_fa456_or0));
  and_gate and_gate_s_wallace_cska32_and_1_18(.a(a[1]), .b(b[18]), .out(s_wallace_cska32_and_1_18));
  and_gate and_gate_s_wallace_cska32_and_0_19(.a(a[0]), .b(b[19]), .out(s_wallace_cska32_and_0_19));
  fa fa_s_wallace_cska32_fa457_out(.a(s_wallace_cska32_fa456_or0[0]), .b(s_wallace_cska32_and_1_18[0]), .cin(s_wallace_cska32_and_0_19[0]), .fa_xor1(s_wallace_cska32_fa457_xor1), .fa_or0(s_wallace_cska32_fa457_or0));
  and_gate and_gate_s_wallace_cska32_and_2_18(.a(a[2]), .b(b[18]), .out(s_wallace_cska32_and_2_18));
  and_gate and_gate_s_wallace_cska32_and_1_19(.a(a[1]), .b(b[19]), .out(s_wallace_cska32_and_1_19));
  fa fa_s_wallace_cska32_fa458_out(.a(s_wallace_cska32_fa457_or0[0]), .b(s_wallace_cska32_and_2_18[0]), .cin(s_wallace_cska32_and_1_19[0]), .fa_xor1(s_wallace_cska32_fa458_xor1), .fa_or0(s_wallace_cska32_fa458_or0));
  and_gate and_gate_s_wallace_cska32_and_3_18(.a(a[3]), .b(b[18]), .out(s_wallace_cska32_and_3_18));
  and_gate and_gate_s_wallace_cska32_and_2_19(.a(a[2]), .b(b[19]), .out(s_wallace_cska32_and_2_19));
  fa fa_s_wallace_cska32_fa459_out(.a(s_wallace_cska32_fa458_or0[0]), .b(s_wallace_cska32_and_3_18[0]), .cin(s_wallace_cska32_and_2_19[0]), .fa_xor1(s_wallace_cska32_fa459_xor1), .fa_or0(s_wallace_cska32_fa459_or0));
  and_gate and_gate_s_wallace_cska32_and_4_18(.a(a[4]), .b(b[18]), .out(s_wallace_cska32_and_4_18));
  and_gate and_gate_s_wallace_cska32_and_3_19(.a(a[3]), .b(b[19]), .out(s_wallace_cska32_and_3_19));
  fa fa_s_wallace_cska32_fa460_out(.a(s_wallace_cska32_fa459_or0[0]), .b(s_wallace_cska32_and_4_18[0]), .cin(s_wallace_cska32_and_3_19[0]), .fa_xor1(s_wallace_cska32_fa460_xor1), .fa_or0(s_wallace_cska32_fa460_or0));
  and_gate and_gate_s_wallace_cska32_and_5_18(.a(a[5]), .b(b[18]), .out(s_wallace_cska32_and_5_18));
  and_gate and_gate_s_wallace_cska32_and_4_19(.a(a[4]), .b(b[19]), .out(s_wallace_cska32_and_4_19));
  fa fa_s_wallace_cska32_fa461_out(.a(s_wallace_cska32_fa460_or0[0]), .b(s_wallace_cska32_and_5_18[0]), .cin(s_wallace_cska32_and_4_19[0]), .fa_xor1(s_wallace_cska32_fa461_xor1), .fa_or0(s_wallace_cska32_fa461_or0));
  and_gate and_gate_s_wallace_cska32_and_6_18(.a(a[6]), .b(b[18]), .out(s_wallace_cska32_and_6_18));
  and_gate and_gate_s_wallace_cska32_and_5_19(.a(a[5]), .b(b[19]), .out(s_wallace_cska32_and_5_19));
  fa fa_s_wallace_cska32_fa462_out(.a(s_wallace_cska32_fa461_or0[0]), .b(s_wallace_cska32_and_6_18[0]), .cin(s_wallace_cska32_and_5_19[0]), .fa_xor1(s_wallace_cska32_fa462_xor1), .fa_or0(s_wallace_cska32_fa462_or0));
  and_gate and_gate_s_wallace_cska32_and_7_18(.a(a[7]), .b(b[18]), .out(s_wallace_cska32_and_7_18));
  and_gate and_gate_s_wallace_cska32_and_6_19(.a(a[6]), .b(b[19]), .out(s_wallace_cska32_and_6_19));
  fa fa_s_wallace_cska32_fa463_out(.a(s_wallace_cska32_fa462_or0[0]), .b(s_wallace_cska32_and_7_18[0]), .cin(s_wallace_cska32_and_6_19[0]), .fa_xor1(s_wallace_cska32_fa463_xor1), .fa_or0(s_wallace_cska32_fa463_or0));
  and_gate and_gate_s_wallace_cska32_and_8_18(.a(a[8]), .b(b[18]), .out(s_wallace_cska32_and_8_18));
  and_gate and_gate_s_wallace_cska32_and_7_19(.a(a[7]), .b(b[19]), .out(s_wallace_cska32_and_7_19));
  fa fa_s_wallace_cska32_fa464_out(.a(s_wallace_cska32_fa463_or0[0]), .b(s_wallace_cska32_and_8_18[0]), .cin(s_wallace_cska32_and_7_19[0]), .fa_xor1(s_wallace_cska32_fa464_xor1), .fa_or0(s_wallace_cska32_fa464_or0));
  and_gate and_gate_s_wallace_cska32_and_9_18(.a(a[9]), .b(b[18]), .out(s_wallace_cska32_and_9_18));
  and_gate and_gate_s_wallace_cska32_and_8_19(.a(a[8]), .b(b[19]), .out(s_wallace_cska32_and_8_19));
  fa fa_s_wallace_cska32_fa465_out(.a(s_wallace_cska32_fa464_or0[0]), .b(s_wallace_cska32_and_9_18[0]), .cin(s_wallace_cska32_and_8_19[0]), .fa_xor1(s_wallace_cska32_fa465_xor1), .fa_or0(s_wallace_cska32_fa465_or0));
  and_gate and_gate_s_wallace_cska32_and_10_18(.a(a[10]), .b(b[18]), .out(s_wallace_cska32_and_10_18));
  and_gate and_gate_s_wallace_cska32_and_9_19(.a(a[9]), .b(b[19]), .out(s_wallace_cska32_and_9_19));
  fa fa_s_wallace_cska32_fa466_out(.a(s_wallace_cska32_fa465_or0[0]), .b(s_wallace_cska32_and_10_18[0]), .cin(s_wallace_cska32_and_9_19[0]), .fa_xor1(s_wallace_cska32_fa466_xor1), .fa_or0(s_wallace_cska32_fa466_or0));
  and_gate and_gate_s_wallace_cska32_and_11_18(.a(a[11]), .b(b[18]), .out(s_wallace_cska32_and_11_18));
  and_gate and_gate_s_wallace_cska32_and_10_19(.a(a[10]), .b(b[19]), .out(s_wallace_cska32_and_10_19));
  fa fa_s_wallace_cska32_fa467_out(.a(s_wallace_cska32_fa466_or0[0]), .b(s_wallace_cska32_and_11_18[0]), .cin(s_wallace_cska32_and_10_19[0]), .fa_xor1(s_wallace_cska32_fa467_xor1), .fa_or0(s_wallace_cska32_fa467_or0));
  and_gate and_gate_s_wallace_cska32_and_12_18(.a(a[12]), .b(b[18]), .out(s_wallace_cska32_and_12_18));
  and_gate and_gate_s_wallace_cska32_and_11_19(.a(a[11]), .b(b[19]), .out(s_wallace_cska32_and_11_19));
  fa fa_s_wallace_cska32_fa468_out(.a(s_wallace_cska32_fa467_or0[0]), .b(s_wallace_cska32_and_12_18[0]), .cin(s_wallace_cska32_and_11_19[0]), .fa_xor1(s_wallace_cska32_fa468_xor1), .fa_or0(s_wallace_cska32_fa468_or0));
  and_gate and_gate_s_wallace_cska32_and_13_18(.a(a[13]), .b(b[18]), .out(s_wallace_cska32_and_13_18));
  and_gate and_gate_s_wallace_cska32_and_12_19(.a(a[12]), .b(b[19]), .out(s_wallace_cska32_and_12_19));
  fa fa_s_wallace_cska32_fa469_out(.a(s_wallace_cska32_fa468_or0[0]), .b(s_wallace_cska32_and_13_18[0]), .cin(s_wallace_cska32_and_12_19[0]), .fa_xor1(s_wallace_cska32_fa469_xor1), .fa_or0(s_wallace_cska32_fa469_or0));
  and_gate and_gate_s_wallace_cska32_and_14_18(.a(a[14]), .b(b[18]), .out(s_wallace_cska32_and_14_18));
  and_gate and_gate_s_wallace_cska32_and_13_19(.a(a[13]), .b(b[19]), .out(s_wallace_cska32_and_13_19));
  fa fa_s_wallace_cska32_fa470_out(.a(s_wallace_cska32_fa469_or0[0]), .b(s_wallace_cska32_and_14_18[0]), .cin(s_wallace_cska32_and_13_19[0]), .fa_xor1(s_wallace_cska32_fa470_xor1), .fa_or0(s_wallace_cska32_fa470_or0));
  and_gate and_gate_s_wallace_cska32_and_13_20(.a(a[13]), .b(b[20]), .out(s_wallace_cska32_and_13_20));
  and_gate and_gate_s_wallace_cska32_and_12_21(.a(a[12]), .b(b[21]), .out(s_wallace_cska32_and_12_21));
  fa fa_s_wallace_cska32_fa471_out(.a(s_wallace_cska32_fa470_or0[0]), .b(s_wallace_cska32_and_13_20[0]), .cin(s_wallace_cska32_and_12_21[0]), .fa_xor1(s_wallace_cska32_fa471_xor1), .fa_or0(s_wallace_cska32_fa471_or0));
  and_gate and_gate_s_wallace_cska32_and_13_21(.a(a[13]), .b(b[21]), .out(s_wallace_cska32_and_13_21));
  and_gate and_gate_s_wallace_cska32_and_12_22(.a(a[12]), .b(b[22]), .out(s_wallace_cska32_and_12_22));
  fa fa_s_wallace_cska32_fa472_out(.a(s_wallace_cska32_fa471_or0[0]), .b(s_wallace_cska32_and_13_21[0]), .cin(s_wallace_cska32_and_12_22[0]), .fa_xor1(s_wallace_cska32_fa472_xor1), .fa_or0(s_wallace_cska32_fa472_or0));
  and_gate and_gate_s_wallace_cska32_and_13_22(.a(a[13]), .b(b[22]), .out(s_wallace_cska32_and_13_22));
  and_gate and_gate_s_wallace_cska32_and_12_23(.a(a[12]), .b(b[23]), .out(s_wallace_cska32_and_12_23));
  fa fa_s_wallace_cska32_fa473_out(.a(s_wallace_cska32_fa472_or0[0]), .b(s_wallace_cska32_and_13_22[0]), .cin(s_wallace_cska32_and_12_23[0]), .fa_xor1(s_wallace_cska32_fa473_xor1), .fa_or0(s_wallace_cska32_fa473_or0));
  and_gate and_gate_s_wallace_cska32_and_13_23(.a(a[13]), .b(b[23]), .out(s_wallace_cska32_and_13_23));
  and_gate and_gate_s_wallace_cska32_and_12_24(.a(a[12]), .b(b[24]), .out(s_wallace_cska32_and_12_24));
  fa fa_s_wallace_cska32_fa474_out(.a(s_wallace_cska32_fa473_or0[0]), .b(s_wallace_cska32_and_13_23[0]), .cin(s_wallace_cska32_and_12_24[0]), .fa_xor1(s_wallace_cska32_fa474_xor1), .fa_or0(s_wallace_cska32_fa474_or0));
  and_gate and_gate_s_wallace_cska32_and_13_24(.a(a[13]), .b(b[24]), .out(s_wallace_cska32_and_13_24));
  and_gate and_gate_s_wallace_cska32_and_12_25(.a(a[12]), .b(b[25]), .out(s_wallace_cska32_and_12_25));
  fa fa_s_wallace_cska32_fa475_out(.a(s_wallace_cska32_fa474_or0[0]), .b(s_wallace_cska32_and_13_24[0]), .cin(s_wallace_cska32_and_12_25[0]), .fa_xor1(s_wallace_cska32_fa475_xor1), .fa_or0(s_wallace_cska32_fa475_or0));
  and_gate and_gate_s_wallace_cska32_and_13_25(.a(a[13]), .b(b[25]), .out(s_wallace_cska32_and_13_25));
  and_gate and_gate_s_wallace_cska32_and_12_26(.a(a[12]), .b(b[26]), .out(s_wallace_cska32_and_12_26));
  fa fa_s_wallace_cska32_fa476_out(.a(s_wallace_cska32_fa475_or0[0]), .b(s_wallace_cska32_and_13_25[0]), .cin(s_wallace_cska32_and_12_26[0]), .fa_xor1(s_wallace_cska32_fa476_xor1), .fa_or0(s_wallace_cska32_fa476_or0));
  and_gate and_gate_s_wallace_cska32_and_13_26(.a(a[13]), .b(b[26]), .out(s_wallace_cska32_and_13_26));
  and_gate and_gate_s_wallace_cska32_and_12_27(.a(a[12]), .b(b[27]), .out(s_wallace_cska32_and_12_27));
  fa fa_s_wallace_cska32_fa477_out(.a(s_wallace_cska32_fa476_or0[0]), .b(s_wallace_cska32_and_13_26[0]), .cin(s_wallace_cska32_and_12_27[0]), .fa_xor1(s_wallace_cska32_fa477_xor1), .fa_or0(s_wallace_cska32_fa477_or0));
  and_gate and_gate_s_wallace_cska32_and_13_27(.a(a[13]), .b(b[27]), .out(s_wallace_cska32_and_13_27));
  and_gate and_gate_s_wallace_cska32_and_12_28(.a(a[12]), .b(b[28]), .out(s_wallace_cska32_and_12_28));
  fa fa_s_wallace_cska32_fa478_out(.a(s_wallace_cska32_fa477_or0[0]), .b(s_wallace_cska32_and_13_27[0]), .cin(s_wallace_cska32_and_12_28[0]), .fa_xor1(s_wallace_cska32_fa478_xor1), .fa_or0(s_wallace_cska32_fa478_or0));
  and_gate and_gate_s_wallace_cska32_and_13_28(.a(a[13]), .b(b[28]), .out(s_wallace_cska32_and_13_28));
  and_gate and_gate_s_wallace_cska32_and_12_29(.a(a[12]), .b(b[29]), .out(s_wallace_cska32_and_12_29));
  fa fa_s_wallace_cska32_fa479_out(.a(s_wallace_cska32_fa478_or0[0]), .b(s_wallace_cska32_and_13_28[0]), .cin(s_wallace_cska32_and_12_29[0]), .fa_xor1(s_wallace_cska32_fa479_xor1), .fa_or0(s_wallace_cska32_fa479_or0));
  and_gate and_gate_s_wallace_cska32_and_13_29(.a(a[13]), .b(b[29]), .out(s_wallace_cska32_and_13_29));
  and_gate and_gate_s_wallace_cska32_and_12_30(.a(a[12]), .b(b[30]), .out(s_wallace_cska32_and_12_30));
  fa fa_s_wallace_cska32_fa480_out(.a(s_wallace_cska32_fa479_or0[0]), .b(s_wallace_cska32_and_13_29[0]), .cin(s_wallace_cska32_and_12_30[0]), .fa_xor1(s_wallace_cska32_fa480_xor1), .fa_or0(s_wallace_cska32_fa480_or0));
  and_gate and_gate_s_wallace_cska32_and_13_30(.a(a[13]), .b(b[30]), .out(s_wallace_cska32_and_13_30));
  nand_gate nand_gate_s_wallace_cska32_nand_12_31(.a(a[12]), .b(b[31]), .out(s_wallace_cska32_nand_12_31));
  fa fa_s_wallace_cska32_fa481_out(.a(s_wallace_cska32_fa480_or0[0]), .b(s_wallace_cska32_and_13_30[0]), .cin(s_wallace_cska32_nand_12_31[0]), .fa_xor1(s_wallace_cska32_fa481_xor1), .fa_or0(s_wallace_cska32_fa481_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_13_31(.a(a[13]), .b(b[31]), .out(s_wallace_cska32_nand_13_31));
  fa fa_s_wallace_cska32_fa482_out(.a(s_wallace_cska32_fa481_or0[0]), .b(s_wallace_cska32_nand_13_31[0]), .cin(s_wallace_cska32_fa41_xor1[0]), .fa_xor1(s_wallace_cska32_fa482_xor1), .fa_or0(s_wallace_cska32_fa482_or0));
  fa fa_s_wallace_cska32_fa483_out(.a(s_wallace_cska32_fa482_or0[0]), .b(s_wallace_cska32_fa42_xor1[0]), .cin(s_wallace_cska32_fa99_xor1[0]), .fa_xor1(s_wallace_cska32_fa483_xor1), .fa_or0(s_wallace_cska32_fa483_or0));
  fa fa_s_wallace_cska32_fa484_out(.a(s_wallace_cska32_fa483_or0[0]), .b(s_wallace_cska32_fa100_xor1[0]), .cin(s_wallace_cska32_fa155_xor1[0]), .fa_xor1(s_wallace_cska32_fa484_xor1), .fa_or0(s_wallace_cska32_fa484_or0));
  fa fa_s_wallace_cska32_fa485_out(.a(s_wallace_cska32_fa484_or0[0]), .b(s_wallace_cska32_fa156_xor1[0]), .cin(s_wallace_cska32_fa209_xor1[0]), .fa_xor1(s_wallace_cska32_fa485_xor1), .fa_or0(s_wallace_cska32_fa485_or0));
  fa fa_s_wallace_cska32_fa486_out(.a(s_wallace_cska32_fa485_or0[0]), .b(s_wallace_cska32_fa210_xor1[0]), .cin(s_wallace_cska32_fa261_xor1[0]), .fa_xor1(s_wallace_cska32_fa486_xor1), .fa_or0(s_wallace_cska32_fa486_or0));
  fa fa_s_wallace_cska32_fa487_out(.a(s_wallace_cska32_fa486_or0[0]), .b(s_wallace_cska32_fa262_xor1[0]), .cin(s_wallace_cska32_fa311_xor1[0]), .fa_xor1(s_wallace_cska32_fa487_xor1), .fa_or0(s_wallace_cska32_fa487_or0));
  fa fa_s_wallace_cska32_fa488_out(.a(s_wallace_cska32_fa487_or0[0]), .b(s_wallace_cska32_fa312_xor1[0]), .cin(s_wallace_cska32_fa359_xor1[0]), .fa_xor1(s_wallace_cska32_fa488_xor1), .fa_or0(s_wallace_cska32_fa488_or0));
  fa fa_s_wallace_cska32_fa489_out(.a(s_wallace_cska32_fa488_or0[0]), .b(s_wallace_cska32_fa360_xor1[0]), .cin(s_wallace_cska32_fa405_xor1[0]), .fa_xor1(s_wallace_cska32_fa489_xor1), .fa_or0(s_wallace_cska32_fa489_or0));
  ha ha_s_wallace_cska32_ha10_out(.a(s_wallace_cska32_fa366_xor1[0]), .b(s_wallace_cska32_fa409_xor1[0]), .ha_xor0(s_wallace_cska32_ha10_xor0), .ha_and0(s_wallace_cska32_ha10_and0));
  fa fa_s_wallace_cska32_fa490_out(.a(s_wallace_cska32_ha10_and0[0]), .b(s_wallace_cska32_fa322_xor1[0]), .cin(s_wallace_cska32_fa367_xor1[0]), .fa_xor1(s_wallace_cska32_fa490_xor1), .fa_or0(s_wallace_cska32_fa490_or0));
  fa fa_s_wallace_cska32_fa491_out(.a(s_wallace_cska32_fa490_or0[0]), .b(s_wallace_cska32_fa276_xor1[0]), .cin(s_wallace_cska32_fa323_xor1[0]), .fa_xor1(s_wallace_cska32_fa491_xor1), .fa_or0(s_wallace_cska32_fa491_or0));
  fa fa_s_wallace_cska32_fa492_out(.a(s_wallace_cska32_fa491_or0[0]), .b(s_wallace_cska32_fa228_xor1[0]), .cin(s_wallace_cska32_fa277_xor1[0]), .fa_xor1(s_wallace_cska32_fa492_xor1), .fa_or0(s_wallace_cska32_fa492_or0));
  fa fa_s_wallace_cska32_fa493_out(.a(s_wallace_cska32_fa492_or0[0]), .b(s_wallace_cska32_fa178_xor1[0]), .cin(s_wallace_cska32_fa229_xor1[0]), .fa_xor1(s_wallace_cska32_fa493_xor1), .fa_or0(s_wallace_cska32_fa493_or0));
  fa fa_s_wallace_cska32_fa494_out(.a(s_wallace_cska32_fa493_or0[0]), .b(s_wallace_cska32_fa126_xor1[0]), .cin(s_wallace_cska32_fa179_xor1[0]), .fa_xor1(s_wallace_cska32_fa494_xor1), .fa_or0(s_wallace_cska32_fa494_or0));
  fa fa_s_wallace_cska32_fa495_out(.a(s_wallace_cska32_fa494_or0[0]), .b(s_wallace_cska32_fa72_xor1[0]), .cin(s_wallace_cska32_fa127_xor1[0]), .fa_xor1(s_wallace_cska32_fa495_xor1), .fa_or0(s_wallace_cska32_fa495_or0));
  fa fa_s_wallace_cska32_fa496_out(.a(s_wallace_cska32_fa495_or0[0]), .b(s_wallace_cska32_fa16_xor1[0]), .cin(s_wallace_cska32_fa73_xor1[0]), .fa_xor1(s_wallace_cska32_fa496_xor1), .fa_or0(s_wallace_cska32_fa496_or0));
  and_gate and_gate_s_wallace_cska32_and_0_20(.a(a[0]), .b(b[20]), .out(s_wallace_cska32_and_0_20));
  fa fa_s_wallace_cska32_fa497_out(.a(s_wallace_cska32_fa496_or0[0]), .b(s_wallace_cska32_and_0_20[0]), .cin(s_wallace_cska32_fa17_xor1[0]), .fa_xor1(s_wallace_cska32_fa497_xor1), .fa_or0(s_wallace_cska32_fa497_or0));
  and_gate and_gate_s_wallace_cska32_and_1_20(.a(a[1]), .b(b[20]), .out(s_wallace_cska32_and_1_20));
  and_gate and_gate_s_wallace_cska32_and_0_21(.a(a[0]), .b(b[21]), .out(s_wallace_cska32_and_0_21));
  fa fa_s_wallace_cska32_fa498_out(.a(s_wallace_cska32_fa497_or0[0]), .b(s_wallace_cska32_and_1_20[0]), .cin(s_wallace_cska32_and_0_21[0]), .fa_xor1(s_wallace_cska32_fa498_xor1), .fa_or0(s_wallace_cska32_fa498_or0));
  and_gate and_gate_s_wallace_cska32_and_2_20(.a(a[2]), .b(b[20]), .out(s_wallace_cska32_and_2_20));
  and_gate and_gate_s_wallace_cska32_and_1_21(.a(a[1]), .b(b[21]), .out(s_wallace_cska32_and_1_21));
  fa fa_s_wallace_cska32_fa499_out(.a(s_wallace_cska32_fa498_or0[0]), .b(s_wallace_cska32_and_2_20[0]), .cin(s_wallace_cska32_and_1_21[0]), .fa_xor1(s_wallace_cska32_fa499_xor1), .fa_or0(s_wallace_cska32_fa499_or0));
  and_gate and_gate_s_wallace_cska32_and_3_20(.a(a[3]), .b(b[20]), .out(s_wallace_cska32_and_3_20));
  and_gate and_gate_s_wallace_cska32_and_2_21(.a(a[2]), .b(b[21]), .out(s_wallace_cska32_and_2_21));
  fa fa_s_wallace_cska32_fa500_out(.a(s_wallace_cska32_fa499_or0[0]), .b(s_wallace_cska32_and_3_20[0]), .cin(s_wallace_cska32_and_2_21[0]), .fa_xor1(s_wallace_cska32_fa500_xor1), .fa_or0(s_wallace_cska32_fa500_or0));
  and_gate and_gate_s_wallace_cska32_and_4_20(.a(a[4]), .b(b[20]), .out(s_wallace_cska32_and_4_20));
  and_gate and_gate_s_wallace_cska32_and_3_21(.a(a[3]), .b(b[21]), .out(s_wallace_cska32_and_3_21));
  fa fa_s_wallace_cska32_fa501_out(.a(s_wallace_cska32_fa500_or0[0]), .b(s_wallace_cska32_and_4_20[0]), .cin(s_wallace_cska32_and_3_21[0]), .fa_xor1(s_wallace_cska32_fa501_xor1), .fa_or0(s_wallace_cska32_fa501_or0));
  and_gate and_gate_s_wallace_cska32_and_5_20(.a(a[5]), .b(b[20]), .out(s_wallace_cska32_and_5_20));
  and_gate and_gate_s_wallace_cska32_and_4_21(.a(a[4]), .b(b[21]), .out(s_wallace_cska32_and_4_21));
  fa fa_s_wallace_cska32_fa502_out(.a(s_wallace_cska32_fa501_or0[0]), .b(s_wallace_cska32_and_5_20[0]), .cin(s_wallace_cska32_and_4_21[0]), .fa_xor1(s_wallace_cska32_fa502_xor1), .fa_or0(s_wallace_cska32_fa502_or0));
  and_gate and_gate_s_wallace_cska32_and_6_20(.a(a[6]), .b(b[20]), .out(s_wallace_cska32_and_6_20));
  and_gate and_gate_s_wallace_cska32_and_5_21(.a(a[5]), .b(b[21]), .out(s_wallace_cska32_and_5_21));
  fa fa_s_wallace_cska32_fa503_out(.a(s_wallace_cska32_fa502_or0[0]), .b(s_wallace_cska32_and_6_20[0]), .cin(s_wallace_cska32_and_5_21[0]), .fa_xor1(s_wallace_cska32_fa503_xor1), .fa_or0(s_wallace_cska32_fa503_or0));
  and_gate and_gate_s_wallace_cska32_and_7_20(.a(a[7]), .b(b[20]), .out(s_wallace_cska32_and_7_20));
  and_gate and_gate_s_wallace_cska32_and_6_21(.a(a[6]), .b(b[21]), .out(s_wallace_cska32_and_6_21));
  fa fa_s_wallace_cska32_fa504_out(.a(s_wallace_cska32_fa503_or0[0]), .b(s_wallace_cska32_and_7_20[0]), .cin(s_wallace_cska32_and_6_21[0]), .fa_xor1(s_wallace_cska32_fa504_xor1), .fa_or0(s_wallace_cska32_fa504_or0));
  and_gate and_gate_s_wallace_cska32_and_8_20(.a(a[8]), .b(b[20]), .out(s_wallace_cska32_and_8_20));
  and_gate and_gate_s_wallace_cska32_and_7_21(.a(a[7]), .b(b[21]), .out(s_wallace_cska32_and_7_21));
  fa fa_s_wallace_cska32_fa505_out(.a(s_wallace_cska32_fa504_or0[0]), .b(s_wallace_cska32_and_8_20[0]), .cin(s_wallace_cska32_and_7_21[0]), .fa_xor1(s_wallace_cska32_fa505_xor1), .fa_or0(s_wallace_cska32_fa505_or0));
  and_gate and_gate_s_wallace_cska32_and_9_20(.a(a[9]), .b(b[20]), .out(s_wallace_cska32_and_9_20));
  and_gate and_gate_s_wallace_cska32_and_8_21(.a(a[8]), .b(b[21]), .out(s_wallace_cska32_and_8_21));
  fa fa_s_wallace_cska32_fa506_out(.a(s_wallace_cska32_fa505_or0[0]), .b(s_wallace_cska32_and_9_20[0]), .cin(s_wallace_cska32_and_8_21[0]), .fa_xor1(s_wallace_cska32_fa506_xor1), .fa_or0(s_wallace_cska32_fa506_or0));
  and_gate and_gate_s_wallace_cska32_and_10_20(.a(a[10]), .b(b[20]), .out(s_wallace_cska32_and_10_20));
  and_gate and_gate_s_wallace_cska32_and_9_21(.a(a[9]), .b(b[21]), .out(s_wallace_cska32_and_9_21));
  fa fa_s_wallace_cska32_fa507_out(.a(s_wallace_cska32_fa506_or0[0]), .b(s_wallace_cska32_and_10_20[0]), .cin(s_wallace_cska32_and_9_21[0]), .fa_xor1(s_wallace_cska32_fa507_xor1), .fa_or0(s_wallace_cska32_fa507_or0));
  and_gate and_gate_s_wallace_cska32_and_11_20(.a(a[11]), .b(b[20]), .out(s_wallace_cska32_and_11_20));
  and_gate and_gate_s_wallace_cska32_and_10_21(.a(a[10]), .b(b[21]), .out(s_wallace_cska32_and_10_21));
  fa fa_s_wallace_cska32_fa508_out(.a(s_wallace_cska32_fa507_or0[0]), .b(s_wallace_cska32_and_11_20[0]), .cin(s_wallace_cska32_and_10_21[0]), .fa_xor1(s_wallace_cska32_fa508_xor1), .fa_or0(s_wallace_cska32_fa508_or0));
  and_gate and_gate_s_wallace_cska32_and_12_20(.a(a[12]), .b(b[20]), .out(s_wallace_cska32_and_12_20));
  and_gate and_gate_s_wallace_cska32_and_11_21(.a(a[11]), .b(b[21]), .out(s_wallace_cska32_and_11_21));
  fa fa_s_wallace_cska32_fa509_out(.a(s_wallace_cska32_fa508_or0[0]), .b(s_wallace_cska32_and_12_20[0]), .cin(s_wallace_cska32_and_11_21[0]), .fa_xor1(s_wallace_cska32_fa509_xor1), .fa_or0(s_wallace_cska32_fa509_or0));
  and_gate and_gate_s_wallace_cska32_and_11_22(.a(a[11]), .b(b[22]), .out(s_wallace_cska32_and_11_22));
  and_gate and_gate_s_wallace_cska32_and_10_23(.a(a[10]), .b(b[23]), .out(s_wallace_cska32_and_10_23));
  fa fa_s_wallace_cska32_fa510_out(.a(s_wallace_cska32_fa509_or0[0]), .b(s_wallace_cska32_and_11_22[0]), .cin(s_wallace_cska32_and_10_23[0]), .fa_xor1(s_wallace_cska32_fa510_xor1), .fa_or0(s_wallace_cska32_fa510_or0));
  and_gate and_gate_s_wallace_cska32_and_11_23(.a(a[11]), .b(b[23]), .out(s_wallace_cska32_and_11_23));
  and_gate and_gate_s_wallace_cska32_and_10_24(.a(a[10]), .b(b[24]), .out(s_wallace_cska32_and_10_24));
  fa fa_s_wallace_cska32_fa511_out(.a(s_wallace_cska32_fa510_or0[0]), .b(s_wallace_cska32_and_11_23[0]), .cin(s_wallace_cska32_and_10_24[0]), .fa_xor1(s_wallace_cska32_fa511_xor1), .fa_or0(s_wallace_cska32_fa511_or0));
  and_gate and_gate_s_wallace_cska32_and_11_24(.a(a[11]), .b(b[24]), .out(s_wallace_cska32_and_11_24));
  and_gate and_gate_s_wallace_cska32_and_10_25(.a(a[10]), .b(b[25]), .out(s_wallace_cska32_and_10_25));
  fa fa_s_wallace_cska32_fa512_out(.a(s_wallace_cska32_fa511_or0[0]), .b(s_wallace_cska32_and_11_24[0]), .cin(s_wallace_cska32_and_10_25[0]), .fa_xor1(s_wallace_cska32_fa512_xor1), .fa_or0(s_wallace_cska32_fa512_or0));
  and_gate and_gate_s_wallace_cska32_and_11_25(.a(a[11]), .b(b[25]), .out(s_wallace_cska32_and_11_25));
  and_gate and_gate_s_wallace_cska32_and_10_26(.a(a[10]), .b(b[26]), .out(s_wallace_cska32_and_10_26));
  fa fa_s_wallace_cska32_fa513_out(.a(s_wallace_cska32_fa512_or0[0]), .b(s_wallace_cska32_and_11_25[0]), .cin(s_wallace_cska32_and_10_26[0]), .fa_xor1(s_wallace_cska32_fa513_xor1), .fa_or0(s_wallace_cska32_fa513_or0));
  and_gate and_gate_s_wallace_cska32_and_11_26(.a(a[11]), .b(b[26]), .out(s_wallace_cska32_and_11_26));
  and_gate and_gate_s_wallace_cska32_and_10_27(.a(a[10]), .b(b[27]), .out(s_wallace_cska32_and_10_27));
  fa fa_s_wallace_cska32_fa514_out(.a(s_wallace_cska32_fa513_or0[0]), .b(s_wallace_cska32_and_11_26[0]), .cin(s_wallace_cska32_and_10_27[0]), .fa_xor1(s_wallace_cska32_fa514_xor1), .fa_or0(s_wallace_cska32_fa514_or0));
  and_gate and_gate_s_wallace_cska32_and_11_27(.a(a[11]), .b(b[27]), .out(s_wallace_cska32_and_11_27));
  and_gate and_gate_s_wallace_cska32_and_10_28(.a(a[10]), .b(b[28]), .out(s_wallace_cska32_and_10_28));
  fa fa_s_wallace_cska32_fa515_out(.a(s_wallace_cska32_fa514_or0[0]), .b(s_wallace_cska32_and_11_27[0]), .cin(s_wallace_cska32_and_10_28[0]), .fa_xor1(s_wallace_cska32_fa515_xor1), .fa_or0(s_wallace_cska32_fa515_or0));
  and_gate and_gate_s_wallace_cska32_and_11_28(.a(a[11]), .b(b[28]), .out(s_wallace_cska32_and_11_28));
  and_gate and_gate_s_wallace_cska32_and_10_29(.a(a[10]), .b(b[29]), .out(s_wallace_cska32_and_10_29));
  fa fa_s_wallace_cska32_fa516_out(.a(s_wallace_cska32_fa515_or0[0]), .b(s_wallace_cska32_and_11_28[0]), .cin(s_wallace_cska32_and_10_29[0]), .fa_xor1(s_wallace_cska32_fa516_xor1), .fa_or0(s_wallace_cska32_fa516_or0));
  and_gate and_gate_s_wallace_cska32_and_11_29(.a(a[11]), .b(b[29]), .out(s_wallace_cska32_and_11_29));
  and_gate and_gate_s_wallace_cska32_and_10_30(.a(a[10]), .b(b[30]), .out(s_wallace_cska32_and_10_30));
  fa fa_s_wallace_cska32_fa517_out(.a(s_wallace_cska32_fa516_or0[0]), .b(s_wallace_cska32_and_11_29[0]), .cin(s_wallace_cska32_and_10_30[0]), .fa_xor1(s_wallace_cska32_fa517_xor1), .fa_or0(s_wallace_cska32_fa517_or0));
  and_gate and_gate_s_wallace_cska32_and_11_30(.a(a[11]), .b(b[30]), .out(s_wallace_cska32_and_11_30));
  nand_gate nand_gate_s_wallace_cska32_nand_10_31(.a(a[10]), .b(b[31]), .out(s_wallace_cska32_nand_10_31));
  fa fa_s_wallace_cska32_fa518_out(.a(s_wallace_cska32_fa517_or0[0]), .b(s_wallace_cska32_and_11_30[0]), .cin(s_wallace_cska32_nand_10_31[0]), .fa_xor1(s_wallace_cska32_fa518_xor1), .fa_or0(s_wallace_cska32_fa518_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_11_31(.a(a[11]), .b(b[31]), .out(s_wallace_cska32_nand_11_31));
  fa fa_s_wallace_cska32_fa519_out(.a(s_wallace_cska32_fa518_or0[0]), .b(s_wallace_cska32_nand_11_31[0]), .cin(s_wallace_cska32_fa39_xor1[0]), .fa_xor1(s_wallace_cska32_fa519_xor1), .fa_or0(s_wallace_cska32_fa519_or0));
  fa fa_s_wallace_cska32_fa520_out(.a(s_wallace_cska32_fa519_or0[0]), .b(s_wallace_cska32_fa40_xor1[0]), .cin(s_wallace_cska32_fa97_xor1[0]), .fa_xor1(s_wallace_cska32_fa520_xor1), .fa_or0(s_wallace_cska32_fa520_or0));
  fa fa_s_wallace_cska32_fa521_out(.a(s_wallace_cska32_fa520_or0[0]), .b(s_wallace_cska32_fa98_xor1[0]), .cin(s_wallace_cska32_fa153_xor1[0]), .fa_xor1(s_wallace_cska32_fa521_xor1), .fa_or0(s_wallace_cska32_fa521_or0));
  fa fa_s_wallace_cska32_fa522_out(.a(s_wallace_cska32_fa521_or0[0]), .b(s_wallace_cska32_fa154_xor1[0]), .cin(s_wallace_cska32_fa207_xor1[0]), .fa_xor1(s_wallace_cska32_fa522_xor1), .fa_or0(s_wallace_cska32_fa522_or0));
  fa fa_s_wallace_cska32_fa523_out(.a(s_wallace_cska32_fa522_or0[0]), .b(s_wallace_cska32_fa208_xor1[0]), .cin(s_wallace_cska32_fa259_xor1[0]), .fa_xor1(s_wallace_cska32_fa523_xor1), .fa_or0(s_wallace_cska32_fa523_or0));
  fa fa_s_wallace_cska32_fa524_out(.a(s_wallace_cska32_fa523_or0[0]), .b(s_wallace_cska32_fa260_xor1[0]), .cin(s_wallace_cska32_fa309_xor1[0]), .fa_xor1(s_wallace_cska32_fa524_xor1), .fa_or0(s_wallace_cska32_fa524_or0));
  fa fa_s_wallace_cska32_fa525_out(.a(s_wallace_cska32_fa524_or0[0]), .b(s_wallace_cska32_fa310_xor1[0]), .cin(s_wallace_cska32_fa357_xor1[0]), .fa_xor1(s_wallace_cska32_fa525_xor1), .fa_or0(s_wallace_cska32_fa525_or0));
  fa fa_s_wallace_cska32_fa526_out(.a(s_wallace_cska32_fa525_or0[0]), .b(s_wallace_cska32_fa358_xor1[0]), .cin(s_wallace_cska32_fa403_xor1[0]), .fa_xor1(s_wallace_cska32_fa526_xor1), .fa_or0(s_wallace_cska32_fa526_or0));
  fa fa_s_wallace_cska32_fa527_out(.a(s_wallace_cska32_fa526_or0[0]), .b(s_wallace_cska32_fa404_xor1[0]), .cin(s_wallace_cska32_fa447_xor1[0]), .fa_xor1(s_wallace_cska32_fa527_xor1), .fa_or0(s_wallace_cska32_fa527_or0));
  ha ha_s_wallace_cska32_ha11_out(.a(s_wallace_cska32_fa410_xor1[0]), .b(s_wallace_cska32_fa451_xor1[0]), .ha_xor0(s_wallace_cska32_ha11_xor0), .ha_and0(s_wallace_cska32_ha11_and0));
  fa fa_s_wallace_cska32_fa528_out(.a(s_wallace_cska32_ha11_and0[0]), .b(s_wallace_cska32_fa368_xor1[0]), .cin(s_wallace_cska32_fa411_xor1[0]), .fa_xor1(s_wallace_cska32_fa528_xor1), .fa_or0(s_wallace_cska32_fa528_or0));
  fa fa_s_wallace_cska32_fa529_out(.a(s_wallace_cska32_fa528_or0[0]), .b(s_wallace_cska32_fa324_xor1[0]), .cin(s_wallace_cska32_fa369_xor1[0]), .fa_xor1(s_wallace_cska32_fa529_xor1), .fa_or0(s_wallace_cska32_fa529_or0));
  fa fa_s_wallace_cska32_fa530_out(.a(s_wallace_cska32_fa529_or0[0]), .b(s_wallace_cska32_fa278_xor1[0]), .cin(s_wallace_cska32_fa325_xor1[0]), .fa_xor1(s_wallace_cska32_fa530_xor1), .fa_or0(s_wallace_cska32_fa530_or0));
  fa fa_s_wallace_cska32_fa531_out(.a(s_wallace_cska32_fa530_or0[0]), .b(s_wallace_cska32_fa230_xor1[0]), .cin(s_wallace_cska32_fa279_xor1[0]), .fa_xor1(s_wallace_cska32_fa531_xor1), .fa_or0(s_wallace_cska32_fa531_or0));
  fa fa_s_wallace_cska32_fa532_out(.a(s_wallace_cska32_fa531_or0[0]), .b(s_wallace_cska32_fa180_xor1[0]), .cin(s_wallace_cska32_fa231_xor1[0]), .fa_xor1(s_wallace_cska32_fa532_xor1), .fa_or0(s_wallace_cska32_fa532_or0));
  fa fa_s_wallace_cska32_fa533_out(.a(s_wallace_cska32_fa532_or0[0]), .b(s_wallace_cska32_fa128_xor1[0]), .cin(s_wallace_cska32_fa181_xor1[0]), .fa_xor1(s_wallace_cska32_fa533_xor1), .fa_or0(s_wallace_cska32_fa533_or0));
  fa fa_s_wallace_cska32_fa534_out(.a(s_wallace_cska32_fa533_or0[0]), .b(s_wallace_cska32_fa74_xor1[0]), .cin(s_wallace_cska32_fa129_xor1[0]), .fa_xor1(s_wallace_cska32_fa534_xor1), .fa_or0(s_wallace_cska32_fa534_or0));
  fa fa_s_wallace_cska32_fa535_out(.a(s_wallace_cska32_fa534_or0[0]), .b(s_wallace_cska32_fa18_xor1[0]), .cin(s_wallace_cska32_fa75_xor1[0]), .fa_xor1(s_wallace_cska32_fa535_xor1), .fa_or0(s_wallace_cska32_fa535_or0));
  and_gate and_gate_s_wallace_cska32_and_0_22(.a(a[0]), .b(b[22]), .out(s_wallace_cska32_and_0_22));
  fa fa_s_wallace_cska32_fa536_out(.a(s_wallace_cska32_fa535_or0[0]), .b(s_wallace_cska32_and_0_22[0]), .cin(s_wallace_cska32_fa19_xor1[0]), .fa_xor1(s_wallace_cska32_fa536_xor1), .fa_or0(s_wallace_cska32_fa536_or0));
  and_gate and_gate_s_wallace_cska32_and_1_22(.a(a[1]), .b(b[22]), .out(s_wallace_cska32_and_1_22));
  and_gate and_gate_s_wallace_cska32_and_0_23(.a(a[0]), .b(b[23]), .out(s_wallace_cska32_and_0_23));
  fa fa_s_wallace_cska32_fa537_out(.a(s_wallace_cska32_fa536_or0[0]), .b(s_wallace_cska32_and_1_22[0]), .cin(s_wallace_cska32_and_0_23[0]), .fa_xor1(s_wallace_cska32_fa537_xor1), .fa_or0(s_wallace_cska32_fa537_or0));
  and_gate and_gate_s_wallace_cska32_and_2_22(.a(a[2]), .b(b[22]), .out(s_wallace_cska32_and_2_22));
  and_gate and_gate_s_wallace_cska32_and_1_23(.a(a[1]), .b(b[23]), .out(s_wallace_cska32_and_1_23));
  fa fa_s_wallace_cska32_fa538_out(.a(s_wallace_cska32_fa537_or0[0]), .b(s_wallace_cska32_and_2_22[0]), .cin(s_wallace_cska32_and_1_23[0]), .fa_xor1(s_wallace_cska32_fa538_xor1), .fa_or0(s_wallace_cska32_fa538_or0));
  and_gate and_gate_s_wallace_cska32_and_3_22(.a(a[3]), .b(b[22]), .out(s_wallace_cska32_and_3_22));
  and_gate and_gate_s_wallace_cska32_and_2_23(.a(a[2]), .b(b[23]), .out(s_wallace_cska32_and_2_23));
  fa fa_s_wallace_cska32_fa539_out(.a(s_wallace_cska32_fa538_or0[0]), .b(s_wallace_cska32_and_3_22[0]), .cin(s_wallace_cska32_and_2_23[0]), .fa_xor1(s_wallace_cska32_fa539_xor1), .fa_or0(s_wallace_cska32_fa539_or0));
  and_gate and_gate_s_wallace_cska32_and_4_22(.a(a[4]), .b(b[22]), .out(s_wallace_cska32_and_4_22));
  and_gate and_gate_s_wallace_cska32_and_3_23(.a(a[3]), .b(b[23]), .out(s_wallace_cska32_and_3_23));
  fa fa_s_wallace_cska32_fa540_out(.a(s_wallace_cska32_fa539_or0[0]), .b(s_wallace_cska32_and_4_22[0]), .cin(s_wallace_cska32_and_3_23[0]), .fa_xor1(s_wallace_cska32_fa540_xor1), .fa_or0(s_wallace_cska32_fa540_or0));
  and_gate and_gate_s_wallace_cska32_and_5_22(.a(a[5]), .b(b[22]), .out(s_wallace_cska32_and_5_22));
  and_gate and_gate_s_wallace_cska32_and_4_23(.a(a[4]), .b(b[23]), .out(s_wallace_cska32_and_4_23));
  fa fa_s_wallace_cska32_fa541_out(.a(s_wallace_cska32_fa540_or0[0]), .b(s_wallace_cska32_and_5_22[0]), .cin(s_wallace_cska32_and_4_23[0]), .fa_xor1(s_wallace_cska32_fa541_xor1), .fa_or0(s_wallace_cska32_fa541_or0));
  and_gate and_gate_s_wallace_cska32_and_6_22(.a(a[6]), .b(b[22]), .out(s_wallace_cska32_and_6_22));
  and_gate and_gate_s_wallace_cska32_and_5_23(.a(a[5]), .b(b[23]), .out(s_wallace_cska32_and_5_23));
  fa fa_s_wallace_cska32_fa542_out(.a(s_wallace_cska32_fa541_or0[0]), .b(s_wallace_cska32_and_6_22[0]), .cin(s_wallace_cska32_and_5_23[0]), .fa_xor1(s_wallace_cska32_fa542_xor1), .fa_or0(s_wallace_cska32_fa542_or0));
  and_gate and_gate_s_wallace_cska32_and_7_22(.a(a[7]), .b(b[22]), .out(s_wallace_cska32_and_7_22));
  and_gate and_gate_s_wallace_cska32_and_6_23(.a(a[6]), .b(b[23]), .out(s_wallace_cska32_and_6_23));
  fa fa_s_wallace_cska32_fa543_out(.a(s_wallace_cska32_fa542_or0[0]), .b(s_wallace_cska32_and_7_22[0]), .cin(s_wallace_cska32_and_6_23[0]), .fa_xor1(s_wallace_cska32_fa543_xor1), .fa_or0(s_wallace_cska32_fa543_or0));
  and_gate and_gate_s_wallace_cska32_and_8_22(.a(a[8]), .b(b[22]), .out(s_wallace_cska32_and_8_22));
  and_gate and_gate_s_wallace_cska32_and_7_23(.a(a[7]), .b(b[23]), .out(s_wallace_cska32_and_7_23));
  fa fa_s_wallace_cska32_fa544_out(.a(s_wallace_cska32_fa543_or0[0]), .b(s_wallace_cska32_and_8_22[0]), .cin(s_wallace_cska32_and_7_23[0]), .fa_xor1(s_wallace_cska32_fa544_xor1), .fa_or0(s_wallace_cska32_fa544_or0));
  and_gate and_gate_s_wallace_cska32_and_9_22(.a(a[9]), .b(b[22]), .out(s_wallace_cska32_and_9_22));
  and_gate and_gate_s_wallace_cska32_and_8_23(.a(a[8]), .b(b[23]), .out(s_wallace_cska32_and_8_23));
  fa fa_s_wallace_cska32_fa545_out(.a(s_wallace_cska32_fa544_or0[0]), .b(s_wallace_cska32_and_9_22[0]), .cin(s_wallace_cska32_and_8_23[0]), .fa_xor1(s_wallace_cska32_fa545_xor1), .fa_or0(s_wallace_cska32_fa545_or0));
  and_gate and_gate_s_wallace_cska32_and_10_22(.a(a[10]), .b(b[22]), .out(s_wallace_cska32_and_10_22));
  and_gate and_gate_s_wallace_cska32_and_9_23(.a(a[9]), .b(b[23]), .out(s_wallace_cska32_and_9_23));
  fa fa_s_wallace_cska32_fa546_out(.a(s_wallace_cska32_fa545_or0[0]), .b(s_wallace_cska32_and_10_22[0]), .cin(s_wallace_cska32_and_9_23[0]), .fa_xor1(s_wallace_cska32_fa546_xor1), .fa_or0(s_wallace_cska32_fa546_or0));
  and_gate and_gate_s_wallace_cska32_and_9_24(.a(a[9]), .b(b[24]), .out(s_wallace_cska32_and_9_24));
  and_gate and_gate_s_wallace_cska32_and_8_25(.a(a[8]), .b(b[25]), .out(s_wallace_cska32_and_8_25));
  fa fa_s_wallace_cska32_fa547_out(.a(s_wallace_cska32_fa546_or0[0]), .b(s_wallace_cska32_and_9_24[0]), .cin(s_wallace_cska32_and_8_25[0]), .fa_xor1(s_wallace_cska32_fa547_xor1), .fa_or0(s_wallace_cska32_fa547_or0));
  and_gate and_gate_s_wallace_cska32_and_9_25(.a(a[9]), .b(b[25]), .out(s_wallace_cska32_and_9_25));
  and_gate and_gate_s_wallace_cska32_and_8_26(.a(a[8]), .b(b[26]), .out(s_wallace_cska32_and_8_26));
  fa fa_s_wallace_cska32_fa548_out(.a(s_wallace_cska32_fa547_or0[0]), .b(s_wallace_cska32_and_9_25[0]), .cin(s_wallace_cska32_and_8_26[0]), .fa_xor1(s_wallace_cska32_fa548_xor1), .fa_or0(s_wallace_cska32_fa548_or0));
  and_gate and_gate_s_wallace_cska32_and_9_26(.a(a[9]), .b(b[26]), .out(s_wallace_cska32_and_9_26));
  and_gate and_gate_s_wallace_cska32_and_8_27(.a(a[8]), .b(b[27]), .out(s_wallace_cska32_and_8_27));
  fa fa_s_wallace_cska32_fa549_out(.a(s_wallace_cska32_fa548_or0[0]), .b(s_wallace_cska32_and_9_26[0]), .cin(s_wallace_cska32_and_8_27[0]), .fa_xor1(s_wallace_cska32_fa549_xor1), .fa_or0(s_wallace_cska32_fa549_or0));
  and_gate and_gate_s_wallace_cska32_and_9_27(.a(a[9]), .b(b[27]), .out(s_wallace_cska32_and_9_27));
  and_gate and_gate_s_wallace_cska32_and_8_28(.a(a[8]), .b(b[28]), .out(s_wallace_cska32_and_8_28));
  fa fa_s_wallace_cska32_fa550_out(.a(s_wallace_cska32_fa549_or0[0]), .b(s_wallace_cska32_and_9_27[0]), .cin(s_wallace_cska32_and_8_28[0]), .fa_xor1(s_wallace_cska32_fa550_xor1), .fa_or0(s_wallace_cska32_fa550_or0));
  and_gate and_gate_s_wallace_cska32_and_9_28(.a(a[9]), .b(b[28]), .out(s_wallace_cska32_and_9_28));
  and_gate and_gate_s_wallace_cska32_and_8_29(.a(a[8]), .b(b[29]), .out(s_wallace_cska32_and_8_29));
  fa fa_s_wallace_cska32_fa551_out(.a(s_wallace_cska32_fa550_or0[0]), .b(s_wallace_cska32_and_9_28[0]), .cin(s_wallace_cska32_and_8_29[0]), .fa_xor1(s_wallace_cska32_fa551_xor1), .fa_or0(s_wallace_cska32_fa551_or0));
  and_gate and_gate_s_wallace_cska32_and_9_29(.a(a[9]), .b(b[29]), .out(s_wallace_cska32_and_9_29));
  and_gate and_gate_s_wallace_cska32_and_8_30(.a(a[8]), .b(b[30]), .out(s_wallace_cska32_and_8_30));
  fa fa_s_wallace_cska32_fa552_out(.a(s_wallace_cska32_fa551_or0[0]), .b(s_wallace_cska32_and_9_29[0]), .cin(s_wallace_cska32_and_8_30[0]), .fa_xor1(s_wallace_cska32_fa552_xor1), .fa_or0(s_wallace_cska32_fa552_or0));
  and_gate and_gate_s_wallace_cska32_and_9_30(.a(a[9]), .b(b[30]), .out(s_wallace_cska32_and_9_30));
  nand_gate nand_gate_s_wallace_cska32_nand_8_31(.a(a[8]), .b(b[31]), .out(s_wallace_cska32_nand_8_31));
  fa fa_s_wallace_cska32_fa553_out(.a(s_wallace_cska32_fa552_or0[0]), .b(s_wallace_cska32_and_9_30[0]), .cin(s_wallace_cska32_nand_8_31[0]), .fa_xor1(s_wallace_cska32_fa553_xor1), .fa_or0(s_wallace_cska32_fa553_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_9_31(.a(a[9]), .b(b[31]), .out(s_wallace_cska32_nand_9_31));
  fa fa_s_wallace_cska32_fa554_out(.a(s_wallace_cska32_fa553_or0[0]), .b(s_wallace_cska32_nand_9_31[0]), .cin(s_wallace_cska32_fa37_xor1[0]), .fa_xor1(s_wallace_cska32_fa554_xor1), .fa_or0(s_wallace_cska32_fa554_or0));
  fa fa_s_wallace_cska32_fa555_out(.a(s_wallace_cska32_fa554_or0[0]), .b(s_wallace_cska32_fa38_xor1[0]), .cin(s_wallace_cska32_fa95_xor1[0]), .fa_xor1(s_wallace_cska32_fa555_xor1), .fa_or0(s_wallace_cska32_fa555_or0));
  fa fa_s_wallace_cska32_fa556_out(.a(s_wallace_cska32_fa555_or0[0]), .b(s_wallace_cska32_fa96_xor1[0]), .cin(s_wallace_cska32_fa151_xor1[0]), .fa_xor1(s_wallace_cska32_fa556_xor1), .fa_or0(s_wallace_cska32_fa556_or0));
  fa fa_s_wallace_cska32_fa557_out(.a(s_wallace_cska32_fa556_or0[0]), .b(s_wallace_cska32_fa152_xor1[0]), .cin(s_wallace_cska32_fa205_xor1[0]), .fa_xor1(s_wallace_cska32_fa557_xor1), .fa_or0(s_wallace_cska32_fa557_or0));
  fa fa_s_wallace_cska32_fa558_out(.a(s_wallace_cska32_fa557_or0[0]), .b(s_wallace_cska32_fa206_xor1[0]), .cin(s_wallace_cska32_fa257_xor1[0]), .fa_xor1(s_wallace_cska32_fa558_xor1), .fa_or0(s_wallace_cska32_fa558_or0));
  fa fa_s_wallace_cska32_fa559_out(.a(s_wallace_cska32_fa558_or0[0]), .b(s_wallace_cska32_fa258_xor1[0]), .cin(s_wallace_cska32_fa307_xor1[0]), .fa_xor1(s_wallace_cska32_fa559_xor1), .fa_or0(s_wallace_cska32_fa559_or0));
  fa fa_s_wallace_cska32_fa560_out(.a(s_wallace_cska32_fa559_or0[0]), .b(s_wallace_cska32_fa308_xor1[0]), .cin(s_wallace_cska32_fa355_xor1[0]), .fa_xor1(s_wallace_cska32_fa560_xor1), .fa_or0(s_wallace_cska32_fa560_or0));
  fa fa_s_wallace_cska32_fa561_out(.a(s_wallace_cska32_fa560_or0[0]), .b(s_wallace_cska32_fa356_xor1[0]), .cin(s_wallace_cska32_fa401_xor1[0]), .fa_xor1(s_wallace_cska32_fa561_xor1), .fa_or0(s_wallace_cska32_fa561_or0));
  fa fa_s_wallace_cska32_fa562_out(.a(s_wallace_cska32_fa561_or0[0]), .b(s_wallace_cska32_fa402_xor1[0]), .cin(s_wallace_cska32_fa445_xor1[0]), .fa_xor1(s_wallace_cska32_fa562_xor1), .fa_or0(s_wallace_cska32_fa562_or0));
  fa fa_s_wallace_cska32_fa563_out(.a(s_wallace_cska32_fa562_or0[0]), .b(s_wallace_cska32_fa446_xor1[0]), .cin(s_wallace_cska32_fa487_xor1[0]), .fa_xor1(s_wallace_cska32_fa563_xor1), .fa_or0(s_wallace_cska32_fa563_or0));
  ha ha_s_wallace_cska32_ha12_out(.a(s_wallace_cska32_fa452_xor1[0]), .b(s_wallace_cska32_fa491_xor1[0]), .ha_xor0(s_wallace_cska32_ha12_xor0), .ha_and0(s_wallace_cska32_ha12_and0));
  fa fa_s_wallace_cska32_fa564_out(.a(s_wallace_cska32_ha12_and0[0]), .b(s_wallace_cska32_fa412_xor1[0]), .cin(s_wallace_cska32_fa453_xor1[0]), .fa_xor1(s_wallace_cska32_fa564_xor1), .fa_or0(s_wallace_cska32_fa564_or0));
  fa fa_s_wallace_cska32_fa565_out(.a(s_wallace_cska32_fa564_or0[0]), .b(s_wallace_cska32_fa370_xor1[0]), .cin(s_wallace_cska32_fa413_xor1[0]), .fa_xor1(s_wallace_cska32_fa565_xor1), .fa_or0(s_wallace_cska32_fa565_or0));
  fa fa_s_wallace_cska32_fa566_out(.a(s_wallace_cska32_fa565_or0[0]), .b(s_wallace_cska32_fa326_xor1[0]), .cin(s_wallace_cska32_fa371_xor1[0]), .fa_xor1(s_wallace_cska32_fa566_xor1), .fa_or0(s_wallace_cska32_fa566_or0));
  fa fa_s_wallace_cska32_fa567_out(.a(s_wallace_cska32_fa566_or0[0]), .b(s_wallace_cska32_fa280_xor1[0]), .cin(s_wallace_cska32_fa327_xor1[0]), .fa_xor1(s_wallace_cska32_fa567_xor1), .fa_or0(s_wallace_cska32_fa567_or0));
  fa fa_s_wallace_cska32_fa568_out(.a(s_wallace_cska32_fa567_or0[0]), .b(s_wallace_cska32_fa232_xor1[0]), .cin(s_wallace_cska32_fa281_xor1[0]), .fa_xor1(s_wallace_cska32_fa568_xor1), .fa_or0(s_wallace_cska32_fa568_or0));
  fa fa_s_wallace_cska32_fa569_out(.a(s_wallace_cska32_fa568_or0[0]), .b(s_wallace_cska32_fa182_xor1[0]), .cin(s_wallace_cska32_fa233_xor1[0]), .fa_xor1(s_wallace_cska32_fa569_xor1), .fa_or0(s_wallace_cska32_fa569_or0));
  fa fa_s_wallace_cska32_fa570_out(.a(s_wallace_cska32_fa569_or0[0]), .b(s_wallace_cska32_fa130_xor1[0]), .cin(s_wallace_cska32_fa183_xor1[0]), .fa_xor1(s_wallace_cska32_fa570_xor1), .fa_or0(s_wallace_cska32_fa570_or0));
  fa fa_s_wallace_cska32_fa571_out(.a(s_wallace_cska32_fa570_or0[0]), .b(s_wallace_cska32_fa76_xor1[0]), .cin(s_wallace_cska32_fa131_xor1[0]), .fa_xor1(s_wallace_cska32_fa571_xor1), .fa_or0(s_wallace_cska32_fa571_or0));
  fa fa_s_wallace_cska32_fa572_out(.a(s_wallace_cska32_fa571_or0[0]), .b(s_wallace_cska32_fa20_xor1[0]), .cin(s_wallace_cska32_fa77_xor1[0]), .fa_xor1(s_wallace_cska32_fa572_xor1), .fa_or0(s_wallace_cska32_fa572_or0));
  and_gate and_gate_s_wallace_cska32_and_0_24(.a(a[0]), .b(b[24]), .out(s_wallace_cska32_and_0_24));
  fa fa_s_wallace_cska32_fa573_out(.a(s_wallace_cska32_fa572_or0[0]), .b(s_wallace_cska32_and_0_24[0]), .cin(s_wallace_cska32_fa21_xor1[0]), .fa_xor1(s_wallace_cska32_fa573_xor1), .fa_or0(s_wallace_cska32_fa573_or0));
  and_gate and_gate_s_wallace_cska32_and_1_24(.a(a[1]), .b(b[24]), .out(s_wallace_cska32_and_1_24));
  and_gate and_gate_s_wallace_cska32_and_0_25(.a(a[0]), .b(b[25]), .out(s_wallace_cska32_and_0_25));
  fa fa_s_wallace_cska32_fa574_out(.a(s_wallace_cska32_fa573_or0[0]), .b(s_wallace_cska32_and_1_24[0]), .cin(s_wallace_cska32_and_0_25[0]), .fa_xor1(s_wallace_cska32_fa574_xor1), .fa_or0(s_wallace_cska32_fa574_or0));
  and_gate and_gate_s_wallace_cska32_and_2_24(.a(a[2]), .b(b[24]), .out(s_wallace_cska32_and_2_24));
  and_gate and_gate_s_wallace_cska32_and_1_25(.a(a[1]), .b(b[25]), .out(s_wallace_cska32_and_1_25));
  fa fa_s_wallace_cska32_fa575_out(.a(s_wallace_cska32_fa574_or0[0]), .b(s_wallace_cska32_and_2_24[0]), .cin(s_wallace_cska32_and_1_25[0]), .fa_xor1(s_wallace_cska32_fa575_xor1), .fa_or0(s_wallace_cska32_fa575_or0));
  and_gate and_gate_s_wallace_cska32_and_3_24(.a(a[3]), .b(b[24]), .out(s_wallace_cska32_and_3_24));
  and_gate and_gate_s_wallace_cska32_and_2_25(.a(a[2]), .b(b[25]), .out(s_wallace_cska32_and_2_25));
  fa fa_s_wallace_cska32_fa576_out(.a(s_wallace_cska32_fa575_or0[0]), .b(s_wallace_cska32_and_3_24[0]), .cin(s_wallace_cska32_and_2_25[0]), .fa_xor1(s_wallace_cska32_fa576_xor1), .fa_or0(s_wallace_cska32_fa576_or0));
  and_gate and_gate_s_wallace_cska32_and_4_24(.a(a[4]), .b(b[24]), .out(s_wallace_cska32_and_4_24));
  and_gate and_gate_s_wallace_cska32_and_3_25(.a(a[3]), .b(b[25]), .out(s_wallace_cska32_and_3_25));
  fa fa_s_wallace_cska32_fa577_out(.a(s_wallace_cska32_fa576_or0[0]), .b(s_wallace_cska32_and_4_24[0]), .cin(s_wallace_cska32_and_3_25[0]), .fa_xor1(s_wallace_cska32_fa577_xor1), .fa_or0(s_wallace_cska32_fa577_or0));
  and_gate and_gate_s_wallace_cska32_and_5_24(.a(a[5]), .b(b[24]), .out(s_wallace_cska32_and_5_24));
  and_gate and_gate_s_wallace_cska32_and_4_25(.a(a[4]), .b(b[25]), .out(s_wallace_cska32_and_4_25));
  fa fa_s_wallace_cska32_fa578_out(.a(s_wallace_cska32_fa577_or0[0]), .b(s_wallace_cska32_and_5_24[0]), .cin(s_wallace_cska32_and_4_25[0]), .fa_xor1(s_wallace_cska32_fa578_xor1), .fa_or0(s_wallace_cska32_fa578_or0));
  and_gate and_gate_s_wallace_cska32_and_6_24(.a(a[6]), .b(b[24]), .out(s_wallace_cska32_and_6_24));
  and_gate and_gate_s_wallace_cska32_and_5_25(.a(a[5]), .b(b[25]), .out(s_wallace_cska32_and_5_25));
  fa fa_s_wallace_cska32_fa579_out(.a(s_wallace_cska32_fa578_or0[0]), .b(s_wallace_cska32_and_6_24[0]), .cin(s_wallace_cska32_and_5_25[0]), .fa_xor1(s_wallace_cska32_fa579_xor1), .fa_or0(s_wallace_cska32_fa579_or0));
  and_gate and_gate_s_wallace_cska32_and_7_24(.a(a[7]), .b(b[24]), .out(s_wallace_cska32_and_7_24));
  and_gate and_gate_s_wallace_cska32_and_6_25(.a(a[6]), .b(b[25]), .out(s_wallace_cska32_and_6_25));
  fa fa_s_wallace_cska32_fa580_out(.a(s_wallace_cska32_fa579_or0[0]), .b(s_wallace_cska32_and_7_24[0]), .cin(s_wallace_cska32_and_6_25[0]), .fa_xor1(s_wallace_cska32_fa580_xor1), .fa_or0(s_wallace_cska32_fa580_or0));
  and_gate and_gate_s_wallace_cska32_and_8_24(.a(a[8]), .b(b[24]), .out(s_wallace_cska32_and_8_24));
  and_gate and_gate_s_wallace_cska32_and_7_25(.a(a[7]), .b(b[25]), .out(s_wallace_cska32_and_7_25));
  fa fa_s_wallace_cska32_fa581_out(.a(s_wallace_cska32_fa580_or0[0]), .b(s_wallace_cska32_and_8_24[0]), .cin(s_wallace_cska32_and_7_25[0]), .fa_xor1(s_wallace_cska32_fa581_xor1), .fa_or0(s_wallace_cska32_fa581_or0));
  and_gate and_gate_s_wallace_cska32_and_7_26(.a(a[7]), .b(b[26]), .out(s_wallace_cska32_and_7_26));
  and_gate and_gate_s_wallace_cska32_and_6_27(.a(a[6]), .b(b[27]), .out(s_wallace_cska32_and_6_27));
  fa fa_s_wallace_cska32_fa582_out(.a(s_wallace_cska32_fa581_or0[0]), .b(s_wallace_cska32_and_7_26[0]), .cin(s_wallace_cska32_and_6_27[0]), .fa_xor1(s_wallace_cska32_fa582_xor1), .fa_or0(s_wallace_cska32_fa582_or0));
  and_gate and_gate_s_wallace_cska32_and_7_27(.a(a[7]), .b(b[27]), .out(s_wallace_cska32_and_7_27));
  and_gate and_gate_s_wallace_cska32_and_6_28(.a(a[6]), .b(b[28]), .out(s_wallace_cska32_and_6_28));
  fa fa_s_wallace_cska32_fa583_out(.a(s_wallace_cska32_fa582_or0[0]), .b(s_wallace_cska32_and_7_27[0]), .cin(s_wallace_cska32_and_6_28[0]), .fa_xor1(s_wallace_cska32_fa583_xor1), .fa_or0(s_wallace_cska32_fa583_or0));
  and_gate and_gate_s_wallace_cska32_and_7_28(.a(a[7]), .b(b[28]), .out(s_wallace_cska32_and_7_28));
  and_gate and_gate_s_wallace_cska32_and_6_29(.a(a[6]), .b(b[29]), .out(s_wallace_cska32_and_6_29));
  fa fa_s_wallace_cska32_fa584_out(.a(s_wallace_cska32_fa583_or0[0]), .b(s_wallace_cska32_and_7_28[0]), .cin(s_wallace_cska32_and_6_29[0]), .fa_xor1(s_wallace_cska32_fa584_xor1), .fa_or0(s_wallace_cska32_fa584_or0));
  and_gate and_gate_s_wallace_cska32_and_7_29(.a(a[7]), .b(b[29]), .out(s_wallace_cska32_and_7_29));
  and_gate and_gate_s_wallace_cska32_and_6_30(.a(a[6]), .b(b[30]), .out(s_wallace_cska32_and_6_30));
  fa fa_s_wallace_cska32_fa585_out(.a(s_wallace_cska32_fa584_or0[0]), .b(s_wallace_cska32_and_7_29[0]), .cin(s_wallace_cska32_and_6_30[0]), .fa_xor1(s_wallace_cska32_fa585_xor1), .fa_or0(s_wallace_cska32_fa585_or0));
  and_gate and_gate_s_wallace_cska32_and_7_30(.a(a[7]), .b(b[30]), .out(s_wallace_cska32_and_7_30));
  nand_gate nand_gate_s_wallace_cska32_nand_6_31(.a(a[6]), .b(b[31]), .out(s_wallace_cska32_nand_6_31));
  fa fa_s_wallace_cska32_fa586_out(.a(s_wallace_cska32_fa585_or0[0]), .b(s_wallace_cska32_and_7_30[0]), .cin(s_wallace_cska32_nand_6_31[0]), .fa_xor1(s_wallace_cska32_fa586_xor1), .fa_or0(s_wallace_cska32_fa586_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_7_31(.a(a[7]), .b(b[31]), .out(s_wallace_cska32_nand_7_31));
  fa fa_s_wallace_cska32_fa587_out(.a(s_wallace_cska32_fa586_or0[0]), .b(s_wallace_cska32_nand_7_31[0]), .cin(s_wallace_cska32_fa35_xor1[0]), .fa_xor1(s_wallace_cska32_fa587_xor1), .fa_or0(s_wallace_cska32_fa587_or0));
  fa fa_s_wallace_cska32_fa588_out(.a(s_wallace_cska32_fa587_or0[0]), .b(s_wallace_cska32_fa36_xor1[0]), .cin(s_wallace_cska32_fa93_xor1[0]), .fa_xor1(s_wallace_cska32_fa588_xor1), .fa_or0(s_wallace_cska32_fa588_or0));
  fa fa_s_wallace_cska32_fa589_out(.a(s_wallace_cska32_fa588_or0[0]), .b(s_wallace_cska32_fa94_xor1[0]), .cin(s_wallace_cska32_fa149_xor1[0]), .fa_xor1(s_wallace_cska32_fa589_xor1), .fa_or0(s_wallace_cska32_fa589_or0));
  fa fa_s_wallace_cska32_fa590_out(.a(s_wallace_cska32_fa589_or0[0]), .b(s_wallace_cska32_fa150_xor1[0]), .cin(s_wallace_cska32_fa203_xor1[0]), .fa_xor1(s_wallace_cska32_fa590_xor1), .fa_or0(s_wallace_cska32_fa590_or0));
  fa fa_s_wallace_cska32_fa591_out(.a(s_wallace_cska32_fa590_or0[0]), .b(s_wallace_cska32_fa204_xor1[0]), .cin(s_wallace_cska32_fa255_xor1[0]), .fa_xor1(s_wallace_cska32_fa591_xor1), .fa_or0(s_wallace_cska32_fa591_or0));
  fa fa_s_wallace_cska32_fa592_out(.a(s_wallace_cska32_fa591_or0[0]), .b(s_wallace_cska32_fa256_xor1[0]), .cin(s_wallace_cska32_fa305_xor1[0]), .fa_xor1(s_wallace_cska32_fa592_xor1), .fa_or0(s_wallace_cska32_fa592_or0));
  fa fa_s_wallace_cska32_fa593_out(.a(s_wallace_cska32_fa592_or0[0]), .b(s_wallace_cska32_fa306_xor1[0]), .cin(s_wallace_cska32_fa353_xor1[0]), .fa_xor1(s_wallace_cska32_fa593_xor1), .fa_or0(s_wallace_cska32_fa593_or0));
  fa fa_s_wallace_cska32_fa594_out(.a(s_wallace_cska32_fa593_or0[0]), .b(s_wallace_cska32_fa354_xor1[0]), .cin(s_wallace_cska32_fa399_xor1[0]), .fa_xor1(s_wallace_cska32_fa594_xor1), .fa_or0(s_wallace_cska32_fa594_or0));
  fa fa_s_wallace_cska32_fa595_out(.a(s_wallace_cska32_fa594_or0[0]), .b(s_wallace_cska32_fa400_xor1[0]), .cin(s_wallace_cska32_fa443_xor1[0]), .fa_xor1(s_wallace_cska32_fa595_xor1), .fa_or0(s_wallace_cska32_fa595_or0));
  fa fa_s_wallace_cska32_fa596_out(.a(s_wallace_cska32_fa595_or0[0]), .b(s_wallace_cska32_fa444_xor1[0]), .cin(s_wallace_cska32_fa485_xor1[0]), .fa_xor1(s_wallace_cska32_fa596_xor1), .fa_or0(s_wallace_cska32_fa596_or0));
  fa fa_s_wallace_cska32_fa597_out(.a(s_wallace_cska32_fa596_or0[0]), .b(s_wallace_cska32_fa486_xor1[0]), .cin(s_wallace_cska32_fa525_xor1[0]), .fa_xor1(s_wallace_cska32_fa597_xor1), .fa_or0(s_wallace_cska32_fa597_or0));
  ha ha_s_wallace_cska32_ha13_out(.a(s_wallace_cska32_fa492_xor1[0]), .b(s_wallace_cska32_fa529_xor1[0]), .ha_xor0(s_wallace_cska32_ha13_xor0), .ha_and0(s_wallace_cska32_ha13_and0));
  fa fa_s_wallace_cska32_fa598_out(.a(s_wallace_cska32_ha13_and0[0]), .b(s_wallace_cska32_fa454_xor1[0]), .cin(s_wallace_cska32_fa493_xor1[0]), .fa_xor1(s_wallace_cska32_fa598_xor1), .fa_or0(s_wallace_cska32_fa598_or0));
  fa fa_s_wallace_cska32_fa599_out(.a(s_wallace_cska32_fa598_or0[0]), .b(s_wallace_cska32_fa414_xor1[0]), .cin(s_wallace_cska32_fa455_xor1[0]), .fa_xor1(s_wallace_cska32_fa599_xor1), .fa_or0(s_wallace_cska32_fa599_or0));
  fa fa_s_wallace_cska32_fa600_out(.a(s_wallace_cska32_fa599_or0[0]), .b(s_wallace_cska32_fa372_xor1[0]), .cin(s_wallace_cska32_fa415_xor1[0]), .fa_xor1(s_wallace_cska32_fa600_xor1), .fa_or0(s_wallace_cska32_fa600_or0));
  fa fa_s_wallace_cska32_fa601_out(.a(s_wallace_cska32_fa600_or0[0]), .b(s_wallace_cska32_fa328_xor1[0]), .cin(s_wallace_cska32_fa373_xor1[0]), .fa_xor1(s_wallace_cska32_fa601_xor1), .fa_or0(s_wallace_cska32_fa601_or0));
  fa fa_s_wallace_cska32_fa602_out(.a(s_wallace_cska32_fa601_or0[0]), .b(s_wallace_cska32_fa282_xor1[0]), .cin(s_wallace_cska32_fa329_xor1[0]), .fa_xor1(s_wallace_cska32_fa602_xor1), .fa_or0(s_wallace_cska32_fa602_or0));
  fa fa_s_wallace_cska32_fa603_out(.a(s_wallace_cska32_fa602_or0[0]), .b(s_wallace_cska32_fa234_xor1[0]), .cin(s_wallace_cska32_fa283_xor1[0]), .fa_xor1(s_wallace_cska32_fa603_xor1), .fa_or0(s_wallace_cska32_fa603_or0));
  fa fa_s_wallace_cska32_fa604_out(.a(s_wallace_cska32_fa603_or0[0]), .b(s_wallace_cska32_fa184_xor1[0]), .cin(s_wallace_cska32_fa235_xor1[0]), .fa_xor1(s_wallace_cska32_fa604_xor1), .fa_or0(s_wallace_cska32_fa604_or0));
  fa fa_s_wallace_cska32_fa605_out(.a(s_wallace_cska32_fa604_or0[0]), .b(s_wallace_cska32_fa132_xor1[0]), .cin(s_wallace_cska32_fa185_xor1[0]), .fa_xor1(s_wallace_cska32_fa605_xor1), .fa_or0(s_wallace_cska32_fa605_or0));
  fa fa_s_wallace_cska32_fa606_out(.a(s_wallace_cska32_fa605_or0[0]), .b(s_wallace_cska32_fa78_xor1[0]), .cin(s_wallace_cska32_fa133_xor1[0]), .fa_xor1(s_wallace_cska32_fa606_xor1), .fa_or0(s_wallace_cska32_fa606_or0));
  fa fa_s_wallace_cska32_fa607_out(.a(s_wallace_cska32_fa606_or0[0]), .b(s_wallace_cska32_fa22_xor1[0]), .cin(s_wallace_cska32_fa79_xor1[0]), .fa_xor1(s_wallace_cska32_fa607_xor1), .fa_or0(s_wallace_cska32_fa607_or0));
  and_gate and_gate_s_wallace_cska32_and_0_26(.a(a[0]), .b(b[26]), .out(s_wallace_cska32_and_0_26));
  fa fa_s_wallace_cska32_fa608_out(.a(s_wallace_cska32_fa607_or0[0]), .b(s_wallace_cska32_and_0_26[0]), .cin(s_wallace_cska32_fa23_xor1[0]), .fa_xor1(s_wallace_cska32_fa608_xor1), .fa_or0(s_wallace_cska32_fa608_or0));
  and_gate and_gate_s_wallace_cska32_and_1_26(.a(a[1]), .b(b[26]), .out(s_wallace_cska32_and_1_26));
  and_gate and_gate_s_wallace_cska32_and_0_27(.a(a[0]), .b(b[27]), .out(s_wallace_cska32_and_0_27));
  fa fa_s_wallace_cska32_fa609_out(.a(s_wallace_cska32_fa608_or0[0]), .b(s_wallace_cska32_and_1_26[0]), .cin(s_wallace_cska32_and_0_27[0]), .fa_xor1(s_wallace_cska32_fa609_xor1), .fa_or0(s_wallace_cska32_fa609_or0));
  and_gate and_gate_s_wallace_cska32_and_2_26(.a(a[2]), .b(b[26]), .out(s_wallace_cska32_and_2_26));
  and_gate and_gate_s_wallace_cska32_and_1_27(.a(a[1]), .b(b[27]), .out(s_wallace_cska32_and_1_27));
  fa fa_s_wallace_cska32_fa610_out(.a(s_wallace_cska32_fa609_or0[0]), .b(s_wallace_cska32_and_2_26[0]), .cin(s_wallace_cska32_and_1_27[0]), .fa_xor1(s_wallace_cska32_fa610_xor1), .fa_or0(s_wallace_cska32_fa610_or0));
  and_gate and_gate_s_wallace_cska32_and_3_26(.a(a[3]), .b(b[26]), .out(s_wallace_cska32_and_3_26));
  and_gate and_gate_s_wallace_cska32_and_2_27(.a(a[2]), .b(b[27]), .out(s_wallace_cska32_and_2_27));
  fa fa_s_wallace_cska32_fa611_out(.a(s_wallace_cska32_fa610_or0[0]), .b(s_wallace_cska32_and_3_26[0]), .cin(s_wallace_cska32_and_2_27[0]), .fa_xor1(s_wallace_cska32_fa611_xor1), .fa_or0(s_wallace_cska32_fa611_or0));
  and_gate and_gate_s_wallace_cska32_and_4_26(.a(a[4]), .b(b[26]), .out(s_wallace_cska32_and_4_26));
  and_gate and_gate_s_wallace_cska32_and_3_27(.a(a[3]), .b(b[27]), .out(s_wallace_cska32_and_3_27));
  fa fa_s_wallace_cska32_fa612_out(.a(s_wallace_cska32_fa611_or0[0]), .b(s_wallace_cska32_and_4_26[0]), .cin(s_wallace_cska32_and_3_27[0]), .fa_xor1(s_wallace_cska32_fa612_xor1), .fa_or0(s_wallace_cska32_fa612_or0));
  and_gate and_gate_s_wallace_cska32_and_5_26(.a(a[5]), .b(b[26]), .out(s_wallace_cska32_and_5_26));
  and_gate and_gate_s_wallace_cska32_and_4_27(.a(a[4]), .b(b[27]), .out(s_wallace_cska32_and_4_27));
  fa fa_s_wallace_cska32_fa613_out(.a(s_wallace_cska32_fa612_or0[0]), .b(s_wallace_cska32_and_5_26[0]), .cin(s_wallace_cska32_and_4_27[0]), .fa_xor1(s_wallace_cska32_fa613_xor1), .fa_or0(s_wallace_cska32_fa613_or0));
  and_gate and_gate_s_wallace_cska32_and_6_26(.a(a[6]), .b(b[26]), .out(s_wallace_cska32_and_6_26));
  and_gate and_gate_s_wallace_cska32_and_5_27(.a(a[5]), .b(b[27]), .out(s_wallace_cska32_and_5_27));
  fa fa_s_wallace_cska32_fa614_out(.a(s_wallace_cska32_fa613_or0[0]), .b(s_wallace_cska32_and_6_26[0]), .cin(s_wallace_cska32_and_5_27[0]), .fa_xor1(s_wallace_cska32_fa614_xor1), .fa_or0(s_wallace_cska32_fa614_or0));
  and_gate and_gate_s_wallace_cska32_and_5_28(.a(a[5]), .b(b[28]), .out(s_wallace_cska32_and_5_28));
  and_gate and_gate_s_wallace_cska32_and_4_29(.a(a[4]), .b(b[29]), .out(s_wallace_cska32_and_4_29));
  fa fa_s_wallace_cska32_fa615_out(.a(s_wallace_cska32_fa614_or0[0]), .b(s_wallace_cska32_and_5_28[0]), .cin(s_wallace_cska32_and_4_29[0]), .fa_xor1(s_wallace_cska32_fa615_xor1), .fa_or0(s_wallace_cska32_fa615_or0));
  and_gate and_gate_s_wallace_cska32_and_5_29(.a(a[5]), .b(b[29]), .out(s_wallace_cska32_and_5_29));
  and_gate and_gate_s_wallace_cska32_and_4_30(.a(a[4]), .b(b[30]), .out(s_wallace_cska32_and_4_30));
  fa fa_s_wallace_cska32_fa616_out(.a(s_wallace_cska32_fa615_or0[0]), .b(s_wallace_cska32_and_5_29[0]), .cin(s_wallace_cska32_and_4_30[0]), .fa_xor1(s_wallace_cska32_fa616_xor1), .fa_or0(s_wallace_cska32_fa616_or0));
  and_gate and_gate_s_wallace_cska32_and_5_30(.a(a[5]), .b(b[30]), .out(s_wallace_cska32_and_5_30));
  nand_gate nand_gate_s_wallace_cska32_nand_4_31(.a(a[4]), .b(b[31]), .out(s_wallace_cska32_nand_4_31));
  fa fa_s_wallace_cska32_fa617_out(.a(s_wallace_cska32_fa616_or0[0]), .b(s_wallace_cska32_and_5_30[0]), .cin(s_wallace_cska32_nand_4_31[0]), .fa_xor1(s_wallace_cska32_fa617_xor1), .fa_or0(s_wallace_cska32_fa617_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_5_31(.a(a[5]), .b(b[31]), .out(s_wallace_cska32_nand_5_31));
  fa fa_s_wallace_cska32_fa618_out(.a(s_wallace_cska32_fa617_or0[0]), .b(s_wallace_cska32_nand_5_31[0]), .cin(s_wallace_cska32_fa33_xor1[0]), .fa_xor1(s_wallace_cska32_fa618_xor1), .fa_or0(s_wallace_cska32_fa618_or0));
  fa fa_s_wallace_cska32_fa619_out(.a(s_wallace_cska32_fa618_or0[0]), .b(s_wallace_cska32_fa34_xor1[0]), .cin(s_wallace_cska32_fa91_xor1[0]), .fa_xor1(s_wallace_cska32_fa619_xor1), .fa_or0(s_wallace_cska32_fa619_or0));
  fa fa_s_wallace_cska32_fa620_out(.a(s_wallace_cska32_fa619_or0[0]), .b(s_wallace_cska32_fa92_xor1[0]), .cin(s_wallace_cska32_fa147_xor1[0]), .fa_xor1(s_wallace_cska32_fa620_xor1), .fa_or0(s_wallace_cska32_fa620_or0));
  fa fa_s_wallace_cska32_fa621_out(.a(s_wallace_cska32_fa620_or0[0]), .b(s_wallace_cska32_fa148_xor1[0]), .cin(s_wallace_cska32_fa201_xor1[0]), .fa_xor1(s_wallace_cska32_fa621_xor1), .fa_or0(s_wallace_cska32_fa621_or0));
  fa fa_s_wallace_cska32_fa622_out(.a(s_wallace_cska32_fa621_or0[0]), .b(s_wallace_cska32_fa202_xor1[0]), .cin(s_wallace_cska32_fa253_xor1[0]), .fa_xor1(s_wallace_cska32_fa622_xor1), .fa_or0(s_wallace_cska32_fa622_or0));
  fa fa_s_wallace_cska32_fa623_out(.a(s_wallace_cska32_fa622_or0[0]), .b(s_wallace_cska32_fa254_xor1[0]), .cin(s_wallace_cska32_fa303_xor1[0]), .fa_xor1(s_wallace_cska32_fa623_xor1), .fa_or0(s_wallace_cska32_fa623_or0));
  fa fa_s_wallace_cska32_fa624_out(.a(s_wallace_cska32_fa623_or0[0]), .b(s_wallace_cska32_fa304_xor1[0]), .cin(s_wallace_cska32_fa351_xor1[0]), .fa_xor1(s_wallace_cska32_fa624_xor1), .fa_or0(s_wallace_cska32_fa624_or0));
  fa fa_s_wallace_cska32_fa625_out(.a(s_wallace_cska32_fa624_or0[0]), .b(s_wallace_cska32_fa352_xor1[0]), .cin(s_wallace_cska32_fa397_xor1[0]), .fa_xor1(s_wallace_cska32_fa625_xor1), .fa_or0(s_wallace_cska32_fa625_or0));
  fa fa_s_wallace_cska32_fa626_out(.a(s_wallace_cska32_fa625_or0[0]), .b(s_wallace_cska32_fa398_xor1[0]), .cin(s_wallace_cska32_fa441_xor1[0]), .fa_xor1(s_wallace_cska32_fa626_xor1), .fa_or0(s_wallace_cska32_fa626_or0));
  fa fa_s_wallace_cska32_fa627_out(.a(s_wallace_cska32_fa626_or0[0]), .b(s_wallace_cska32_fa442_xor1[0]), .cin(s_wallace_cska32_fa483_xor1[0]), .fa_xor1(s_wallace_cska32_fa627_xor1), .fa_or0(s_wallace_cska32_fa627_or0));
  fa fa_s_wallace_cska32_fa628_out(.a(s_wallace_cska32_fa627_or0[0]), .b(s_wallace_cska32_fa484_xor1[0]), .cin(s_wallace_cska32_fa523_xor1[0]), .fa_xor1(s_wallace_cska32_fa628_xor1), .fa_or0(s_wallace_cska32_fa628_or0));
  fa fa_s_wallace_cska32_fa629_out(.a(s_wallace_cska32_fa628_or0[0]), .b(s_wallace_cska32_fa524_xor1[0]), .cin(s_wallace_cska32_fa561_xor1[0]), .fa_xor1(s_wallace_cska32_fa629_xor1), .fa_or0(s_wallace_cska32_fa629_or0));
  ha ha_s_wallace_cska32_ha14_out(.a(s_wallace_cska32_fa530_xor1[0]), .b(s_wallace_cska32_fa565_xor1[0]), .ha_xor0(s_wallace_cska32_ha14_xor0), .ha_and0(s_wallace_cska32_ha14_and0));
  fa fa_s_wallace_cska32_fa630_out(.a(s_wallace_cska32_ha14_and0[0]), .b(s_wallace_cska32_fa494_xor1[0]), .cin(s_wallace_cska32_fa531_xor1[0]), .fa_xor1(s_wallace_cska32_fa630_xor1), .fa_or0(s_wallace_cska32_fa630_or0));
  fa fa_s_wallace_cska32_fa631_out(.a(s_wallace_cska32_fa630_or0[0]), .b(s_wallace_cska32_fa456_xor1[0]), .cin(s_wallace_cska32_fa495_xor1[0]), .fa_xor1(s_wallace_cska32_fa631_xor1), .fa_or0(s_wallace_cska32_fa631_or0));
  fa fa_s_wallace_cska32_fa632_out(.a(s_wallace_cska32_fa631_or0[0]), .b(s_wallace_cska32_fa416_xor1[0]), .cin(s_wallace_cska32_fa457_xor1[0]), .fa_xor1(s_wallace_cska32_fa632_xor1), .fa_or0(s_wallace_cska32_fa632_or0));
  fa fa_s_wallace_cska32_fa633_out(.a(s_wallace_cska32_fa632_or0[0]), .b(s_wallace_cska32_fa374_xor1[0]), .cin(s_wallace_cska32_fa417_xor1[0]), .fa_xor1(s_wallace_cska32_fa633_xor1), .fa_or0(s_wallace_cska32_fa633_or0));
  fa fa_s_wallace_cska32_fa634_out(.a(s_wallace_cska32_fa633_or0[0]), .b(s_wallace_cska32_fa330_xor1[0]), .cin(s_wallace_cska32_fa375_xor1[0]), .fa_xor1(s_wallace_cska32_fa634_xor1), .fa_or0(s_wallace_cska32_fa634_or0));
  fa fa_s_wallace_cska32_fa635_out(.a(s_wallace_cska32_fa634_or0[0]), .b(s_wallace_cska32_fa284_xor1[0]), .cin(s_wallace_cska32_fa331_xor1[0]), .fa_xor1(s_wallace_cska32_fa635_xor1), .fa_or0(s_wallace_cska32_fa635_or0));
  fa fa_s_wallace_cska32_fa636_out(.a(s_wallace_cska32_fa635_or0[0]), .b(s_wallace_cska32_fa236_xor1[0]), .cin(s_wallace_cska32_fa285_xor1[0]), .fa_xor1(s_wallace_cska32_fa636_xor1), .fa_or0(s_wallace_cska32_fa636_or0));
  fa fa_s_wallace_cska32_fa637_out(.a(s_wallace_cska32_fa636_or0[0]), .b(s_wallace_cska32_fa186_xor1[0]), .cin(s_wallace_cska32_fa237_xor1[0]), .fa_xor1(s_wallace_cska32_fa637_xor1), .fa_or0(s_wallace_cska32_fa637_or0));
  fa fa_s_wallace_cska32_fa638_out(.a(s_wallace_cska32_fa637_or0[0]), .b(s_wallace_cska32_fa134_xor1[0]), .cin(s_wallace_cska32_fa187_xor1[0]), .fa_xor1(s_wallace_cska32_fa638_xor1), .fa_or0(s_wallace_cska32_fa638_or0));
  fa fa_s_wallace_cska32_fa639_out(.a(s_wallace_cska32_fa638_or0[0]), .b(s_wallace_cska32_fa80_xor1[0]), .cin(s_wallace_cska32_fa135_xor1[0]), .fa_xor1(s_wallace_cska32_fa639_xor1), .fa_or0(s_wallace_cska32_fa639_or0));
  fa fa_s_wallace_cska32_fa640_out(.a(s_wallace_cska32_fa639_or0[0]), .b(s_wallace_cska32_fa24_xor1[0]), .cin(s_wallace_cska32_fa81_xor1[0]), .fa_xor1(s_wallace_cska32_fa640_xor1), .fa_or0(s_wallace_cska32_fa640_or0));
  and_gate and_gate_s_wallace_cska32_and_0_28(.a(a[0]), .b(b[28]), .out(s_wallace_cska32_and_0_28));
  fa fa_s_wallace_cska32_fa641_out(.a(s_wallace_cska32_fa640_or0[0]), .b(s_wallace_cska32_and_0_28[0]), .cin(s_wallace_cska32_fa25_xor1[0]), .fa_xor1(s_wallace_cska32_fa641_xor1), .fa_or0(s_wallace_cska32_fa641_or0));
  and_gate and_gate_s_wallace_cska32_and_1_28(.a(a[1]), .b(b[28]), .out(s_wallace_cska32_and_1_28));
  and_gate and_gate_s_wallace_cska32_and_0_29(.a(a[0]), .b(b[29]), .out(s_wallace_cska32_and_0_29));
  fa fa_s_wallace_cska32_fa642_out(.a(s_wallace_cska32_fa641_or0[0]), .b(s_wallace_cska32_and_1_28[0]), .cin(s_wallace_cska32_and_0_29[0]), .fa_xor1(s_wallace_cska32_fa642_xor1), .fa_or0(s_wallace_cska32_fa642_or0));
  and_gate and_gate_s_wallace_cska32_and_2_28(.a(a[2]), .b(b[28]), .out(s_wallace_cska32_and_2_28));
  and_gate and_gate_s_wallace_cska32_and_1_29(.a(a[1]), .b(b[29]), .out(s_wallace_cska32_and_1_29));
  fa fa_s_wallace_cska32_fa643_out(.a(s_wallace_cska32_fa642_or0[0]), .b(s_wallace_cska32_and_2_28[0]), .cin(s_wallace_cska32_and_1_29[0]), .fa_xor1(s_wallace_cska32_fa643_xor1), .fa_or0(s_wallace_cska32_fa643_or0));
  and_gate and_gate_s_wallace_cska32_and_3_28(.a(a[3]), .b(b[28]), .out(s_wallace_cska32_and_3_28));
  and_gate and_gate_s_wallace_cska32_and_2_29(.a(a[2]), .b(b[29]), .out(s_wallace_cska32_and_2_29));
  fa fa_s_wallace_cska32_fa644_out(.a(s_wallace_cska32_fa643_or0[0]), .b(s_wallace_cska32_and_3_28[0]), .cin(s_wallace_cska32_and_2_29[0]), .fa_xor1(s_wallace_cska32_fa644_xor1), .fa_or0(s_wallace_cska32_fa644_or0));
  and_gate and_gate_s_wallace_cska32_and_4_28(.a(a[4]), .b(b[28]), .out(s_wallace_cska32_and_4_28));
  and_gate and_gate_s_wallace_cska32_and_3_29(.a(a[3]), .b(b[29]), .out(s_wallace_cska32_and_3_29));
  fa fa_s_wallace_cska32_fa645_out(.a(s_wallace_cska32_fa644_or0[0]), .b(s_wallace_cska32_and_4_28[0]), .cin(s_wallace_cska32_and_3_29[0]), .fa_xor1(s_wallace_cska32_fa645_xor1), .fa_or0(s_wallace_cska32_fa645_or0));
  and_gate and_gate_s_wallace_cska32_and_3_30(.a(a[3]), .b(b[30]), .out(s_wallace_cska32_and_3_30));
  nand_gate nand_gate_s_wallace_cska32_nand_2_31(.a(a[2]), .b(b[31]), .out(s_wallace_cska32_nand_2_31));
  fa fa_s_wallace_cska32_fa646_out(.a(s_wallace_cska32_fa645_or0[0]), .b(s_wallace_cska32_and_3_30[0]), .cin(s_wallace_cska32_nand_2_31[0]), .fa_xor1(s_wallace_cska32_fa646_xor1), .fa_or0(s_wallace_cska32_fa646_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_3_31(.a(a[3]), .b(b[31]), .out(s_wallace_cska32_nand_3_31));
  fa fa_s_wallace_cska32_fa647_out(.a(s_wallace_cska32_fa646_or0[0]), .b(s_wallace_cska32_nand_3_31[0]), .cin(s_wallace_cska32_fa31_xor1[0]), .fa_xor1(s_wallace_cska32_fa647_xor1), .fa_or0(s_wallace_cska32_fa647_or0));
  fa fa_s_wallace_cska32_fa648_out(.a(s_wallace_cska32_fa647_or0[0]), .b(s_wallace_cska32_fa32_xor1[0]), .cin(s_wallace_cska32_fa89_xor1[0]), .fa_xor1(s_wallace_cska32_fa648_xor1), .fa_or0(s_wallace_cska32_fa648_or0));
  fa fa_s_wallace_cska32_fa649_out(.a(s_wallace_cska32_fa648_or0[0]), .b(s_wallace_cska32_fa90_xor1[0]), .cin(s_wallace_cska32_fa145_xor1[0]), .fa_xor1(s_wallace_cska32_fa649_xor1), .fa_or0(s_wallace_cska32_fa649_or0));
  fa fa_s_wallace_cska32_fa650_out(.a(s_wallace_cska32_fa649_or0[0]), .b(s_wallace_cska32_fa146_xor1[0]), .cin(s_wallace_cska32_fa199_xor1[0]), .fa_xor1(s_wallace_cska32_fa650_xor1), .fa_or0(s_wallace_cska32_fa650_or0));
  fa fa_s_wallace_cska32_fa651_out(.a(s_wallace_cska32_fa650_or0[0]), .b(s_wallace_cska32_fa200_xor1[0]), .cin(s_wallace_cska32_fa251_xor1[0]), .fa_xor1(s_wallace_cska32_fa651_xor1), .fa_or0(s_wallace_cska32_fa651_or0));
  fa fa_s_wallace_cska32_fa652_out(.a(s_wallace_cska32_fa651_or0[0]), .b(s_wallace_cska32_fa252_xor1[0]), .cin(s_wallace_cska32_fa301_xor1[0]), .fa_xor1(s_wallace_cska32_fa652_xor1), .fa_or0(s_wallace_cska32_fa652_or0));
  fa fa_s_wallace_cska32_fa653_out(.a(s_wallace_cska32_fa652_or0[0]), .b(s_wallace_cska32_fa302_xor1[0]), .cin(s_wallace_cska32_fa349_xor1[0]), .fa_xor1(s_wallace_cska32_fa653_xor1), .fa_or0(s_wallace_cska32_fa653_or0));
  fa fa_s_wallace_cska32_fa654_out(.a(s_wallace_cska32_fa653_or0[0]), .b(s_wallace_cska32_fa350_xor1[0]), .cin(s_wallace_cska32_fa395_xor1[0]), .fa_xor1(s_wallace_cska32_fa654_xor1), .fa_or0(s_wallace_cska32_fa654_or0));
  fa fa_s_wallace_cska32_fa655_out(.a(s_wallace_cska32_fa654_or0[0]), .b(s_wallace_cska32_fa396_xor1[0]), .cin(s_wallace_cska32_fa439_xor1[0]), .fa_xor1(s_wallace_cska32_fa655_xor1), .fa_or0(s_wallace_cska32_fa655_or0));
  fa fa_s_wallace_cska32_fa656_out(.a(s_wallace_cska32_fa655_or0[0]), .b(s_wallace_cska32_fa440_xor1[0]), .cin(s_wallace_cska32_fa481_xor1[0]), .fa_xor1(s_wallace_cska32_fa656_xor1), .fa_or0(s_wallace_cska32_fa656_or0));
  fa fa_s_wallace_cska32_fa657_out(.a(s_wallace_cska32_fa656_or0[0]), .b(s_wallace_cska32_fa482_xor1[0]), .cin(s_wallace_cska32_fa521_xor1[0]), .fa_xor1(s_wallace_cska32_fa657_xor1), .fa_or0(s_wallace_cska32_fa657_or0));
  fa fa_s_wallace_cska32_fa658_out(.a(s_wallace_cska32_fa657_or0[0]), .b(s_wallace_cska32_fa522_xor1[0]), .cin(s_wallace_cska32_fa559_xor1[0]), .fa_xor1(s_wallace_cska32_fa658_xor1), .fa_or0(s_wallace_cska32_fa658_or0));
  fa fa_s_wallace_cska32_fa659_out(.a(s_wallace_cska32_fa658_or0[0]), .b(s_wallace_cska32_fa560_xor1[0]), .cin(s_wallace_cska32_fa595_xor1[0]), .fa_xor1(s_wallace_cska32_fa659_xor1), .fa_or0(s_wallace_cska32_fa659_or0));
  ha ha_s_wallace_cska32_ha15_out(.a(s_wallace_cska32_fa566_xor1[0]), .b(s_wallace_cska32_fa599_xor1[0]), .ha_xor0(s_wallace_cska32_ha15_xor0), .ha_and0(s_wallace_cska32_ha15_and0));
  fa fa_s_wallace_cska32_fa660_out(.a(s_wallace_cska32_ha15_and0[0]), .b(s_wallace_cska32_fa532_xor1[0]), .cin(s_wallace_cska32_fa567_xor1[0]), .fa_xor1(s_wallace_cska32_fa660_xor1), .fa_or0(s_wallace_cska32_fa660_or0));
  fa fa_s_wallace_cska32_fa661_out(.a(s_wallace_cska32_fa660_or0[0]), .b(s_wallace_cska32_fa496_xor1[0]), .cin(s_wallace_cska32_fa533_xor1[0]), .fa_xor1(s_wallace_cska32_fa661_xor1), .fa_or0(s_wallace_cska32_fa661_or0));
  fa fa_s_wallace_cska32_fa662_out(.a(s_wallace_cska32_fa661_or0[0]), .b(s_wallace_cska32_fa458_xor1[0]), .cin(s_wallace_cska32_fa497_xor1[0]), .fa_xor1(s_wallace_cska32_fa662_xor1), .fa_or0(s_wallace_cska32_fa662_or0));
  fa fa_s_wallace_cska32_fa663_out(.a(s_wallace_cska32_fa662_or0[0]), .b(s_wallace_cska32_fa418_xor1[0]), .cin(s_wallace_cska32_fa459_xor1[0]), .fa_xor1(s_wallace_cska32_fa663_xor1), .fa_or0(s_wallace_cska32_fa663_or0));
  fa fa_s_wallace_cska32_fa664_out(.a(s_wallace_cska32_fa663_or0[0]), .b(s_wallace_cska32_fa376_xor1[0]), .cin(s_wallace_cska32_fa419_xor1[0]), .fa_xor1(s_wallace_cska32_fa664_xor1), .fa_or0(s_wallace_cska32_fa664_or0));
  fa fa_s_wallace_cska32_fa665_out(.a(s_wallace_cska32_fa664_or0[0]), .b(s_wallace_cska32_fa332_xor1[0]), .cin(s_wallace_cska32_fa377_xor1[0]), .fa_xor1(s_wallace_cska32_fa665_xor1), .fa_or0(s_wallace_cska32_fa665_or0));
  fa fa_s_wallace_cska32_fa666_out(.a(s_wallace_cska32_fa665_or0[0]), .b(s_wallace_cska32_fa286_xor1[0]), .cin(s_wallace_cska32_fa333_xor1[0]), .fa_xor1(s_wallace_cska32_fa666_xor1), .fa_or0(s_wallace_cska32_fa666_or0));
  fa fa_s_wallace_cska32_fa667_out(.a(s_wallace_cska32_fa666_or0[0]), .b(s_wallace_cska32_fa238_xor1[0]), .cin(s_wallace_cska32_fa287_xor1[0]), .fa_xor1(s_wallace_cska32_fa667_xor1), .fa_or0(s_wallace_cska32_fa667_or0));
  fa fa_s_wallace_cska32_fa668_out(.a(s_wallace_cska32_fa667_or0[0]), .b(s_wallace_cska32_fa188_xor1[0]), .cin(s_wallace_cska32_fa239_xor1[0]), .fa_xor1(s_wallace_cska32_fa668_xor1), .fa_or0(s_wallace_cska32_fa668_or0));
  fa fa_s_wallace_cska32_fa669_out(.a(s_wallace_cska32_fa668_or0[0]), .b(s_wallace_cska32_fa136_xor1[0]), .cin(s_wallace_cska32_fa189_xor1[0]), .fa_xor1(s_wallace_cska32_fa669_xor1), .fa_or0(s_wallace_cska32_fa669_or0));
  fa fa_s_wallace_cska32_fa670_out(.a(s_wallace_cska32_fa669_or0[0]), .b(s_wallace_cska32_fa82_xor1[0]), .cin(s_wallace_cska32_fa137_xor1[0]), .fa_xor1(s_wallace_cska32_fa670_xor1), .fa_or0(s_wallace_cska32_fa670_or0));
  fa fa_s_wallace_cska32_fa671_out(.a(s_wallace_cska32_fa670_or0[0]), .b(s_wallace_cska32_fa26_xor1[0]), .cin(s_wallace_cska32_fa83_xor1[0]), .fa_xor1(s_wallace_cska32_fa671_xor1), .fa_or0(s_wallace_cska32_fa671_or0));
  and_gate and_gate_s_wallace_cska32_and_0_30(.a(a[0]), .b(b[30]), .out(s_wallace_cska32_and_0_30));
  fa fa_s_wallace_cska32_fa672_out(.a(s_wallace_cska32_fa671_or0[0]), .b(s_wallace_cska32_and_0_30[0]), .cin(s_wallace_cska32_fa27_xor1[0]), .fa_xor1(s_wallace_cska32_fa672_xor1), .fa_or0(s_wallace_cska32_fa672_or0));
  and_gate and_gate_s_wallace_cska32_and_1_30(.a(a[1]), .b(b[30]), .out(s_wallace_cska32_and_1_30));
  nand_gate nand_gate_s_wallace_cska32_nand_0_31(.a(a[0]), .b(b[31]), .out(s_wallace_cska32_nand_0_31));
  fa fa_s_wallace_cska32_fa673_out(.a(s_wallace_cska32_fa672_or0[0]), .b(s_wallace_cska32_and_1_30[0]), .cin(s_wallace_cska32_nand_0_31[0]), .fa_xor1(s_wallace_cska32_fa673_xor1), .fa_or0(s_wallace_cska32_fa673_or0));
  and_gate and_gate_s_wallace_cska32_and_2_30(.a(a[2]), .b(b[30]), .out(s_wallace_cska32_and_2_30));
  nand_gate nand_gate_s_wallace_cska32_nand_1_31(.a(a[1]), .b(b[31]), .out(s_wallace_cska32_nand_1_31));
  fa fa_s_wallace_cska32_fa674_out(.a(s_wallace_cska32_fa673_or0[0]), .b(s_wallace_cska32_and_2_30[0]), .cin(s_wallace_cska32_nand_1_31[0]), .fa_xor1(s_wallace_cska32_fa674_xor1), .fa_or0(s_wallace_cska32_fa674_or0));
  fa fa_s_wallace_cska32_fa675_out(.a(s_wallace_cska32_fa674_or0[0]), .b(s_wallace_cska32_fa30_xor1[0]), .cin(s_wallace_cska32_fa87_xor1[0]), .fa_xor1(s_wallace_cska32_fa675_xor1), .fa_or0(s_wallace_cska32_fa675_or0));
  fa fa_s_wallace_cska32_fa676_out(.a(s_wallace_cska32_fa675_or0[0]), .b(s_wallace_cska32_fa88_xor1[0]), .cin(s_wallace_cska32_fa143_xor1[0]), .fa_xor1(s_wallace_cska32_fa676_xor1), .fa_or0(s_wallace_cska32_fa676_or0));
  fa fa_s_wallace_cska32_fa677_out(.a(s_wallace_cska32_fa676_or0[0]), .b(s_wallace_cska32_fa144_xor1[0]), .cin(s_wallace_cska32_fa197_xor1[0]), .fa_xor1(s_wallace_cska32_fa677_xor1), .fa_or0(s_wallace_cska32_fa677_or0));
  fa fa_s_wallace_cska32_fa678_out(.a(s_wallace_cska32_fa677_or0[0]), .b(s_wallace_cska32_fa198_xor1[0]), .cin(s_wallace_cska32_fa249_xor1[0]), .fa_xor1(s_wallace_cska32_fa678_xor1), .fa_or0(s_wallace_cska32_fa678_or0));
  fa fa_s_wallace_cska32_fa679_out(.a(s_wallace_cska32_fa678_or0[0]), .b(s_wallace_cska32_fa250_xor1[0]), .cin(s_wallace_cska32_fa299_xor1[0]), .fa_xor1(s_wallace_cska32_fa679_xor1), .fa_or0(s_wallace_cska32_fa679_or0));
  fa fa_s_wallace_cska32_fa680_out(.a(s_wallace_cska32_fa679_or0[0]), .b(s_wallace_cska32_fa300_xor1[0]), .cin(s_wallace_cska32_fa347_xor1[0]), .fa_xor1(s_wallace_cska32_fa680_xor1), .fa_or0(s_wallace_cska32_fa680_or0));
  fa fa_s_wallace_cska32_fa681_out(.a(s_wallace_cska32_fa680_or0[0]), .b(s_wallace_cska32_fa348_xor1[0]), .cin(s_wallace_cska32_fa393_xor1[0]), .fa_xor1(s_wallace_cska32_fa681_xor1), .fa_or0(s_wallace_cska32_fa681_or0));
  fa fa_s_wallace_cska32_fa682_out(.a(s_wallace_cska32_fa681_or0[0]), .b(s_wallace_cska32_fa394_xor1[0]), .cin(s_wallace_cska32_fa437_xor1[0]), .fa_xor1(s_wallace_cska32_fa682_xor1), .fa_or0(s_wallace_cska32_fa682_or0));
  fa fa_s_wallace_cska32_fa683_out(.a(s_wallace_cska32_fa682_or0[0]), .b(s_wallace_cska32_fa438_xor1[0]), .cin(s_wallace_cska32_fa479_xor1[0]), .fa_xor1(s_wallace_cska32_fa683_xor1), .fa_or0(s_wallace_cska32_fa683_or0));
  fa fa_s_wallace_cska32_fa684_out(.a(s_wallace_cska32_fa683_or0[0]), .b(s_wallace_cska32_fa480_xor1[0]), .cin(s_wallace_cska32_fa519_xor1[0]), .fa_xor1(s_wallace_cska32_fa684_xor1), .fa_or0(s_wallace_cska32_fa684_or0));
  fa fa_s_wallace_cska32_fa685_out(.a(s_wallace_cska32_fa684_or0[0]), .b(s_wallace_cska32_fa520_xor1[0]), .cin(s_wallace_cska32_fa557_xor1[0]), .fa_xor1(s_wallace_cska32_fa685_xor1), .fa_or0(s_wallace_cska32_fa685_or0));
  fa fa_s_wallace_cska32_fa686_out(.a(s_wallace_cska32_fa685_or0[0]), .b(s_wallace_cska32_fa558_xor1[0]), .cin(s_wallace_cska32_fa593_xor1[0]), .fa_xor1(s_wallace_cska32_fa686_xor1), .fa_or0(s_wallace_cska32_fa686_or0));
  fa fa_s_wallace_cska32_fa687_out(.a(s_wallace_cska32_fa686_or0[0]), .b(s_wallace_cska32_fa594_xor1[0]), .cin(s_wallace_cska32_fa627_xor1[0]), .fa_xor1(s_wallace_cska32_fa687_xor1), .fa_or0(s_wallace_cska32_fa687_or0));
  ha ha_s_wallace_cska32_ha16_out(.a(s_wallace_cska32_fa600_xor1[0]), .b(s_wallace_cska32_fa631_xor1[0]), .ha_xor0(s_wallace_cska32_ha16_xor0), .ha_and0(s_wallace_cska32_ha16_and0));
  fa fa_s_wallace_cska32_fa688_out(.a(s_wallace_cska32_ha16_and0[0]), .b(s_wallace_cska32_fa568_xor1[0]), .cin(s_wallace_cska32_fa601_xor1[0]), .fa_xor1(s_wallace_cska32_fa688_xor1), .fa_or0(s_wallace_cska32_fa688_or0));
  fa fa_s_wallace_cska32_fa689_out(.a(s_wallace_cska32_fa688_or0[0]), .b(s_wallace_cska32_fa534_xor1[0]), .cin(s_wallace_cska32_fa569_xor1[0]), .fa_xor1(s_wallace_cska32_fa689_xor1), .fa_or0(s_wallace_cska32_fa689_or0));
  fa fa_s_wallace_cska32_fa690_out(.a(s_wallace_cska32_fa689_or0[0]), .b(s_wallace_cska32_fa498_xor1[0]), .cin(s_wallace_cska32_fa535_xor1[0]), .fa_xor1(s_wallace_cska32_fa690_xor1), .fa_or0(s_wallace_cska32_fa690_or0));
  fa fa_s_wallace_cska32_fa691_out(.a(s_wallace_cska32_fa690_or0[0]), .b(s_wallace_cska32_fa460_xor1[0]), .cin(s_wallace_cska32_fa499_xor1[0]), .fa_xor1(s_wallace_cska32_fa691_xor1), .fa_or0(s_wallace_cska32_fa691_or0));
  fa fa_s_wallace_cska32_fa692_out(.a(s_wallace_cska32_fa691_or0[0]), .b(s_wallace_cska32_fa420_xor1[0]), .cin(s_wallace_cska32_fa461_xor1[0]), .fa_xor1(s_wallace_cska32_fa692_xor1), .fa_or0(s_wallace_cska32_fa692_or0));
  fa fa_s_wallace_cska32_fa693_out(.a(s_wallace_cska32_fa692_or0[0]), .b(s_wallace_cska32_fa378_xor1[0]), .cin(s_wallace_cska32_fa421_xor1[0]), .fa_xor1(s_wallace_cska32_fa693_xor1), .fa_or0(s_wallace_cska32_fa693_or0));
  fa fa_s_wallace_cska32_fa694_out(.a(s_wallace_cska32_fa693_or0[0]), .b(s_wallace_cska32_fa334_xor1[0]), .cin(s_wallace_cska32_fa379_xor1[0]), .fa_xor1(s_wallace_cska32_fa694_xor1), .fa_or0(s_wallace_cska32_fa694_or0));
  fa fa_s_wallace_cska32_fa695_out(.a(s_wallace_cska32_fa694_or0[0]), .b(s_wallace_cska32_fa288_xor1[0]), .cin(s_wallace_cska32_fa335_xor1[0]), .fa_xor1(s_wallace_cska32_fa695_xor1), .fa_or0(s_wallace_cska32_fa695_or0));
  fa fa_s_wallace_cska32_fa696_out(.a(s_wallace_cska32_fa695_or0[0]), .b(s_wallace_cska32_fa240_xor1[0]), .cin(s_wallace_cska32_fa289_xor1[0]), .fa_xor1(s_wallace_cska32_fa696_xor1), .fa_or0(s_wallace_cska32_fa696_or0));
  fa fa_s_wallace_cska32_fa697_out(.a(s_wallace_cska32_fa696_or0[0]), .b(s_wallace_cska32_fa190_xor1[0]), .cin(s_wallace_cska32_fa241_xor1[0]), .fa_xor1(s_wallace_cska32_fa697_xor1), .fa_or0(s_wallace_cska32_fa697_or0));
  fa fa_s_wallace_cska32_fa698_out(.a(s_wallace_cska32_fa697_or0[0]), .b(s_wallace_cska32_fa138_xor1[0]), .cin(s_wallace_cska32_fa191_xor1[0]), .fa_xor1(s_wallace_cska32_fa698_xor1), .fa_or0(s_wallace_cska32_fa698_or0));
  fa fa_s_wallace_cska32_fa699_out(.a(s_wallace_cska32_fa698_or0[0]), .b(s_wallace_cska32_fa84_xor1[0]), .cin(s_wallace_cska32_fa139_xor1[0]), .fa_xor1(s_wallace_cska32_fa699_xor1), .fa_or0(s_wallace_cska32_fa699_or0));
  fa fa_s_wallace_cska32_fa700_out(.a(s_wallace_cska32_fa699_or0[0]), .b(s_wallace_cska32_fa28_xor1[0]), .cin(s_wallace_cska32_fa85_xor1[0]), .fa_xor1(s_wallace_cska32_fa700_xor1), .fa_or0(s_wallace_cska32_fa700_or0));
  fa fa_s_wallace_cska32_fa701_out(.a(s_wallace_cska32_fa700_or0[0]), .b(s_wallace_cska32_fa29_xor1[0]), .cin(s_wallace_cska32_fa86_xor1[0]), .fa_xor1(s_wallace_cska32_fa701_xor1), .fa_or0(s_wallace_cska32_fa701_or0));
  fa fa_s_wallace_cska32_fa702_out(.a(s_wallace_cska32_fa701_or0[0]), .b(s_wallace_cska32_fa142_xor1[0]), .cin(s_wallace_cska32_fa195_xor1[0]), .fa_xor1(s_wallace_cska32_fa702_xor1), .fa_or0(s_wallace_cska32_fa702_or0));
  fa fa_s_wallace_cska32_fa703_out(.a(s_wallace_cska32_fa702_or0[0]), .b(s_wallace_cska32_fa196_xor1[0]), .cin(s_wallace_cska32_fa247_xor1[0]), .fa_xor1(s_wallace_cska32_fa703_xor1), .fa_or0(s_wallace_cska32_fa703_or0));
  fa fa_s_wallace_cska32_fa704_out(.a(s_wallace_cska32_fa703_or0[0]), .b(s_wallace_cska32_fa248_xor1[0]), .cin(s_wallace_cska32_fa297_xor1[0]), .fa_xor1(s_wallace_cska32_fa704_xor1), .fa_or0(s_wallace_cska32_fa704_or0));
  fa fa_s_wallace_cska32_fa705_out(.a(s_wallace_cska32_fa704_or0[0]), .b(s_wallace_cska32_fa298_xor1[0]), .cin(s_wallace_cska32_fa345_xor1[0]), .fa_xor1(s_wallace_cska32_fa705_xor1), .fa_or0(s_wallace_cska32_fa705_or0));
  fa fa_s_wallace_cska32_fa706_out(.a(s_wallace_cska32_fa705_or0[0]), .b(s_wallace_cska32_fa346_xor1[0]), .cin(s_wallace_cska32_fa391_xor1[0]), .fa_xor1(s_wallace_cska32_fa706_xor1), .fa_or0(s_wallace_cska32_fa706_or0));
  fa fa_s_wallace_cska32_fa707_out(.a(s_wallace_cska32_fa706_or0[0]), .b(s_wallace_cska32_fa392_xor1[0]), .cin(s_wallace_cska32_fa435_xor1[0]), .fa_xor1(s_wallace_cska32_fa707_xor1), .fa_or0(s_wallace_cska32_fa707_or0));
  fa fa_s_wallace_cska32_fa708_out(.a(s_wallace_cska32_fa707_or0[0]), .b(s_wallace_cska32_fa436_xor1[0]), .cin(s_wallace_cska32_fa477_xor1[0]), .fa_xor1(s_wallace_cska32_fa708_xor1), .fa_or0(s_wallace_cska32_fa708_or0));
  fa fa_s_wallace_cska32_fa709_out(.a(s_wallace_cska32_fa708_or0[0]), .b(s_wallace_cska32_fa478_xor1[0]), .cin(s_wallace_cska32_fa517_xor1[0]), .fa_xor1(s_wallace_cska32_fa709_xor1), .fa_or0(s_wallace_cska32_fa709_or0));
  fa fa_s_wallace_cska32_fa710_out(.a(s_wallace_cska32_fa709_or0[0]), .b(s_wallace_cska32_fa518_xor1[0]), .cin(s_wallace_cska32_fa555_xor1[0]), .fa_xor1(s_wallace_cska32_fa710_xor1), .fa_or0(s_wallace_cska32_fa710_or0));
  fa fa_s_wallace_cska32_fa711_out(.a(s_wallace_cska32_fa710_or0[0]), .b(s_wallace_cska32_fa556_xor1[0]), .cin(s_wallace_cska32_fa591_xor1[0]), .fa_xor1(s_wallace_cska32_fa711_xor1), .fa_or0(s_wallace_cska32_fa711_or0));
  fa fa_s_wallace_cska32_fa712_out(.a(s_wallace_cska32_fa711_or0[0]), .b(s_wallace_cska32_fa592_xor1[0]), .cin(s_wallace_cska32_fa625_xor1[0]), .fa_xor1(s_wallace_cska32_fa712_xor1), .fa_or0(s_wallace_cska32_fa712_or0));
  fa fa_s_wallace_cska32_fa713_out(.a(s_wallace_cska32_fa712_or0[0]), .b(s_wallace_cska32_fa626_xor1[0]), .cin(s_wallace_cska32_fa657_xor1[0]), .fa_xor1(s_wallace_cska32_fa713_xor1), .fa_or0(s_wallace_cska32_fa713_or0));
  ha ha_s_wallace_cska32_ha17_out(.a(s_wallace_cska32_fa632_xor1[0]), .b(s_wallace_cska32_fa661_xor1[0]), .ha_xor0(s_wallace_cska32_ha17_xor0), .ha_and0(s_wallace_cska32_ha17_and0));
  fa fa_s_wallace_cska32_fa714_out(.a(s_wallace_cska32_ha17_and0[0]), .b(s_wallace_cska32_fa602_xor1[0]), .cin(s_wallace_cska32_fa633_xor1[0]), .fa_xor1(s_wallace_cska32_fa714_xor1), .fa_or0(s_wallace_cska32_fa714_or0));
  fa fa_s_wallace_cska32_fa715_out(.a(s_wallace_cska32_fa714_or0[0]), .b(s_wallace_cska32_fa570_xor1[0]), .cin(s_wallace_cska32_fa603_xor1[0]), .fa_xor1(s_wallace_cska32_fa715_xor1), .fa_or0(s_wallace_cska32_fa715_or0));
  fa fa_s_wallace_cska32_fa716_out(.a(s_wallace_cska32_fa715_or0[0]), .b(s_wallace_cska32_fa536_xor1[0]), .cin(s_wallace_cska32_fa571_xor1[0]), .fa_xor1(s_wallace_cska32_fa716_xor1), .fa_or0(s_wallace_cska32_fa716_or0));
  fa fa_s_wallace_cska32_fa717_out(.a(s_wallace_cska32_fa716_or0[0]), .b(s_wallace_cska32_fa500_xor1[0]), .cin(s_wallace_cska32_fa537_xor1[0]), .fa_xor1(s_wallace_cska32_fa717_xor1), .fa_or0(s_wallace_cska32_fa717_or0));
  fa fa_s_wallace_cska32_fa718_out(.a(s_wallace_cska32_fa717_or0[0]), .b(s_wallace_cska32_fa462_xor1[0]), .cin(s_wallace_cska32_fa501_xor1[0]), .fa_xor1(s_wallace_cska32_fa718_xor1), .fa_or0(s_wallace_cska32_fa718_or0));
  fa fa_s_wallace_cska32_fa719_out(.a(s_wallace_cska32_fa718_or0[0]), .b(s_wallace_cska32_fa422_xor1[0]), .cin(s_wallace_cska32_fa463_xor1[0]), .fa_xor1(s_wallace_cska32_fa719_xor1), .fa_or0(s_wallace_cska32_fa719_or0));
  fa fa_s_wallace_cska32_fa720_out(.a(s_wallace_cska32_fa719_or0[0]), .b(s_wallace_cska32_fa380_xor1[0]), .cin(s_wallace_cska32_fa423_xor1[0]), .fa_xor1(s_wallace_cska32_fa720_xor1), .fa_or0(s_wallace_cska32_fa720_or0));
  fa fa_s_wallace_cska32_fa721_out(.a(s_wallace_cska32_fa720_or0[0]), .b(s_wallace_cska32_fa336_xor1[0]), .cin(s_wallace_cska32_fa381_xor1[0]), .fa_xor1(s_wallace_cska32_fa721_xor1), .fa_or0(s_wallace_cska32_fa721_or0));
  fa fa_s_wallace_cska32_fa722_out(.a(s_wallace_cska32_fa721_or0[0]), .b(s_wallace_cska32_fa290_xor1[0]), .cin(s_wallace_cska32_fa337_xor1[0]), .fa_xor1(s_wallace_cska32_fa722_xor1), .fa_or0(s_wallace_cska32_fa722_or0));
  fa fa_s_wallace_cska32_fa723_out(.a(s_wallace_cska32_fa722_or0[0]), .b(s_wallace_cska32_fa242_xor1[0]), .cin(s_wallace_cska32_fa291_xor1[0]), .fa_xor1(s_wallace_cska32_fa723_xor1), .fa_or0(s_wallace_cska32_fa723_or0));
  fa fa_s_wallace_cska32_fa724_out(.a(s_wallace_cska32_fa723_or0[0]), .b(s_wallace_cska32_fa192_xor1[0]), .cin(s_wallace_cska32_fa243_xor1[0]), .fa_xor1(s_wallace_cska32_fa724_xor1), .fa_or0(s_wallace_cska32_fa724_or0));
  fa fa_s_wallace_cska32_fa725_out(.a(s_wallace_cska32_fa724_or0[0]), .b(s_wallace_cska32_fa140_xor1[0]), .cin(s_wallace_cska32_fa193_xor1[0]), .fa_xor1(s_wallace_cska32_fa725_xor1), .fa_or0(s_wallace_cska32_fa725_or0));
  fa fa_s_wallace_cska32_fa726_out(.a(s_wallace_cska32_fa725_or0[0]), .b(s_wallace_cska32_fa141_xor1[0]), .cin(s_wallace_cska32_fa194_xor1[0]), .fa_xor1(s_wallace_cska32_fa726_xor1), .fa_or0(s_wallace_cska32_fa726_or0));
  fa fa_s_wallace_cska32_fa727_out(.a(s_wallace_cska32_fa726_or0[0]), .b(s_wallace_cska32_fa246_xor1[0]), .cin(s_wallace_cska32_fa295_xor1[0]), .fa_xor1(s_wallace_cska32_fa727_xor1), .fa_or0(s_wallace_cska32_fa727_or0));
  fa fa_s_wallace_cska32_fa728_out(.a(s_wallace_cska32_fa727_or0[0]), .b(s_wallace_cska32_fa296_xor1[0]), .cin(s_wallace_cska32_fa343_xor1[0]), .fa_xor1(s_wallace_cska32_fa728_xor1), .fa_or0(s_wallace_cska32_fa728_or0));
  fa fa_s_wallace_cska32_fa729_out(.a(s_wallace_cska32_fa728_or0[0]), .b(s_wallace_cska32_fa344_xor1[0]), .cin(s_wallace_cska32_fa389_xor1[0]), .fa_xor1(s_wallace_cska32_fa729_xor1), .fa_or0(s_wallace_cska32_fa729_or0));
  fa fa_s_wallace_cska32_fa730_out(.a(s_wallace_cska32_fa729_or0[0]), .b(s_wallace_cska32_fa390_xor1[0]), .cin(s_wallace_cska32_fa433_xor1[0]), .fa_xor1(s_wallace_cska32_fa730_xor1), .fa_or0(s_wallace_cska32_fa730_or0));
  fa fa_s_wallace_cska32_fa731_out(.a(s_wallace_cska32_fa730_or0[0]), .b(s_wallace_cska32_fa434_xor1[0]), .cin(s_wallace_cska32_fa475_xor1[0]), .fa_xor1(s_wallace_cska32_fa731_xor1), .fa_or0(s_wallace_cska32_fa731_or0));
  fa fa_s_wallace_cska32_fa732_out(.a(s_wallace_cska32_fa731_or0[0]), .b(s_wallace_cska32_fa476_xor1[0]), .cin(s_wallace_cska32_fa515_xor1[0]), .fa_xor1(s_wallace_cska32_fa732_xor1), .fa_or0(s_wallace_cska32_fa732_or0));
  fa fa_s_wallace_cska32_fa733_out(.a(s_wallace_cska32_fa732_or0[0]), .b(s_wallace_cska32_fa516_xor1[0]), .cin(s_wallace_cska32_fa553_xor1[0]), .fa_xor1(s_wallace_cska32_fa733_xor1), .fa_or0(s_wallace_cska32_fa733_or0));
  fa fa_s_wallace_cska32_fa734_out(.a(s_wallace_cska32_fa733_or0[0]), .b(s_wallace_cska32_fa554_xor1[0]), .cin(s_wallace_cska32_fa589_xor1[0]), .fa_xor1(s_wallace_cska32_fa734_xor1), .fa_or0(s_wallace_cska32_fa734_or0));
  fa fa_s_wallace_cska32_fa735_out(.a(s_wallace_cska32_fa734_or0[0]), .b(s_wallace_cska32_fa590_xor1[0]), .cin(s_wallace_cska32_fa623_xor1[0]), .fa_xor1(s_wallace_cska32_fa735_xor1), .fa_or0(s_wallace_cska32_fa735_or0));
  fa fa_s_wallace_cska32_fa736_out(.a(s_wallace_cska32_fa735_or0[0]), .b(s_wallace_cska32_fa624_xor1[0]), .cin(s_wallace_cska32_fa655_xor1[0]), .fa_xor1(s_wallace_cska32_fa736_xor1), .fa_or0(s_wallace_cska32_fa736_or0));
  fa fa_s_wallace_cska32_fa737_out(.a(s_wallace_cska32_fa736_or0[0]), .b(s_wallace_cska32_fa656_xor1[0]), .cin(s_wallace_cska32_fa685_xor1[0]), .fa_xor1(s_wallace_cska32_fa737_xor1), .fa_or0(s_wallace_cska32_fa737_or0));
  ha ha_s_wallace_cska32_ha18_out(.a(s_wallace_cska32_fa662_xor1[0]), .b(s_wallace_cska32_fa689_xor1[0]), .ha_xor0(s_wallace_cska32_ha18_xor0), .ha_and0(s_wallace_cska32_ha18_and0));
  fa fa_s_wallace_cska32_fa738_out(.a(s_wallace_cska32_ha18_and0[0]), .b(s_wallace_cska32_fa634_xor1[0]), .cin(s_wallace_cska32_fa663_xor1[0]), .fa_xor1(s_wallace_cska32_fa738_xor1), .fa_or0(s_wallace_cska32_fa738_or0));
  fa fa_s_wallace_cska32_fa739_out(.a(s_wallace_cska32_fa738_or0[0]), .b(s_wallace_cska32_fa604_xor1[0]), .cin(s_wallace_cska32_fa635_xor1[0]), .fa_xor1(s_wallace_cska32_fa739_xor1), .fa_or0(s_wallace_cska32_fa739_or0));
  fa fa_s_wallace_cska32_fa740_out(.a(s_wallace_cska32_fa739_or0[0]), .b(s_wallace_cska32_fa572_xor1[0]), .cin(s_wallace_cska32_fa605_xor1[0]), .fa_xor1(s_wallace_cska32_fa740_xor1), .fa_or0(s_wallace_cska32_fa740_or0));
  fa fa_s_wallace_cska32_fa741_out(.a(s_wallace_cska32_fa740_or0[0]), .b(s_wallace_cska32_fa538_xor1[0]), .cin(s_wallace_cska32_fa573_xor1[0]), .fa_xor1(s_wallace_cska32_fa741_xor1), .fa_or0(s_wallace_cska32_fa741_or0));
  fa fa_s_wallace_cska32_fa742_out(.a(s_wallace_cska32_fa741_or0[0]), .b(s_wallace_cska32_fa502_xor1[0]), .cin(s_wallace_cska32_fa539_xor1[0]), .fa_xor1(s_wallace_cska32_fa742_xor1), .fa_or0(s_wallace_cska32_fa742_or0));
  fa fa_s_wallace_cska32_fa743_out(.a(s_wallace_cska32_fa742_or0[0]), .b(s_wallace_cska32_fa464_xor1[0]), .cin(s_wallace_cska32_fa503_xor1[0]), .fa_xor1(s_wallace_cska32_fa743_xor1), .fa_or0(s_wallace_cska32_fa743_or0));
  fa fa_s_wallace_cska32_fa744_out(.a(s_wallace_cska32_fa743_or0[0]), .b(s_wallace_cska32_fa424_xor1[0]), .cin(s_wallace_cska32_fa465_xor1[0]), .fa_xor1(s_wallace_cska32_fa744_xor1), .fa_or0(s_wallace_cska32_fa744_or0));
  fa fa_s_wallace_cska32_fa745_out(.a(s_wallace_cska32_fa744_or0[0]), .b(s_wallace_cska32_fa382_xor1[0]), .cin(s_wallace_cska32_fa425_xor1[0]), .fa_xor1(s_wallace_cska32_fa745_xor1), .fa_or0(s_wallace_cska32_fa745_or0));
  fa fa_s_wallace_cska32_fa746_out(.a(s_wallace_cska32_fa745_or0[0]), .b(s_wallace_cska32_fa338_xor1[0]), .cin(s_wallace_cska32_fa383_xor1[0]), .fa_xor1(s_wallace_cska32_fa746_xor1), .fa_or0(s_wallace_cska32_fa746_or0));
  fa fa_s_wallace_cska32_fa747_out(.a(s_wallace_cska32_fa746_or0[0]), .b(s_wallace_cska32_fa292_xor1[0]), .cin(s_wallace_cska32_fa339_xor1[0]), .fa_xor1(s_wallace_cska32_fa747_xor1), .fa_or0(s_wallace_cska32_fa747_or0));
  fa fa_s_wallace_cska32_fa748_out(.a(s_wallace_cska32_fa747_or0[0]), .b(s_wallace_cska32_fa244_xor1[0]), .cin(s_wallace_cska32_fa293_xor1[0]), .fa_xor1(s_wallace_cska32_fa748_xor1), .fa_or0(s_wallace_cska32_fa748_or0));
  fa fa_s_wallace_cska32_fa749_out(.a(s_wallace_cska32_fa748_or0[0]), .b(s_wallace_cska32_fa245_xor1[0]), .cin(s_wallace_cska32_fa294_xor1[0]), .fa_xor1(s_wallace_cska32_fa749_xor1), .fa_or0(s_wallace_cska32_fa749_or0));
  fa fa_s_wallace_cska32_fa750_out(.a(s_wallace_cska32_fa749_or0[0]), .b(s_wallace_cska32_fa342_xor1[0]), .cin(s_wallace_cska32_fa387_xor1[0]), .fa_xor1(s_wallace_cska32_fa750_xor1), .fa_or0(s_wallace_cska32_fa750_or0));
  fa fa_s_wallace_cska32_fa751_out(.a(s_wallace_cska32_fa750_or0[0]), .b(s_wallace_cska32_fa388_xor1[0]), .cin(s_wallace_cska32_fa431_xor1[0]), .fa_xor1(s_wallace_cska32_fa751_xor1), .fa_or0(s_wallace_cska32_fa751_or0));
  fa fa_s_wallace_cska32_fa752_out(.a(s_wallace_cska32_fa751_or0[0]), .b(s_wallace_cska32_fa432_xor1[0]), .cin(s_wallace_cska32_fa473_xor1[0]), .fa_xor1(s_wallace_cska32_fa752_xor1), .fa_or0(s_wallace_cska32_fa752_or0));
  fa fa_s_wallace_cska32_fa753_out(.a(s_wallace_cska32_fa752_or0[0]), .b(s_wallace_cska32_fa474_xor1[0]), .cin(s_wallace_cska32_fa513_xor1[0]), .fa_xor1(s_wallace_cska32_fa753_xor1), .fa_or0(s_wallace_cska32_fa753_or0));
  fa fa_s_wallace_cska32_fa754_out(.a(s_wallace_cska32_fa753_or0[0]), .b(s_wallace_cska32_fa514_xor1[0]), .cin(s_wallace_cska32_fa551_xor1[0]), .fa_xor1(s_wallace_cska32_fa754_xor1), .fa_or0(s_wallace_cska32_fa754_or0));
  fa fa_s_wallace_cska32_fa755_out(.a(s_wallace_cska32_fa754_or0[0]), .b(s_wallace_cska32_fa552_xor1[0]), .cin(s_wallace_cska32_fa587_xor1[0]), .fa_xor1(s_wallace_cska32_fa755_xor1), .fa_or0(s_wallace_cska32_fa755_or0));
  fa fa_s_wallace_cska32_fa756_out(.a(s_wallace_cska32_fa755_or0[0]), .b(s_wallace_cska32_fa588_xor1[0]), .cin(s_wallace_cska32_fa621_xor1[0]), .fa_xor1(s_wallace_cska32_fa756_xor1), .fa_or0(s_wallace_cska32_fa756_or0));
  fa fa_s_wallace_cska32_fa757_out(.a(s_wallace_cska32_fa756_or0[0]), .b(s_wallace_cska32_fa622_xor1[0]), .cin(s_wallace_cska32_fa653_xor1[0]), .fa_xor1(s_wallace_cska32_fa757_xor1), .fa_or0(s_wallace_cska32_fa757_or0));
  fa fa_s_wallace_cska32_fa758_out(.a(s_wallace_cska32_fa757_or0[0]), .b(s_wallace_cska32_fa654_xor1[0]), .cin(s_wallace_cska32_fa683_xor1[0]), .fa_xor1(s_wallace_cska32_fa758_xor1), .fa_or0(s_wallace_cska32_fa758_or0));
  fa fa_s_wallace_cska32_fa759_out(.a(s_wallace_cska32_fa758_or0[0]), .b(s_wallace_cska32_fa684_xor1[0]), .cin(s_wallace_cska32_fa711_xor1[0]), .fa_xor1(s_wallace_cska32_fa759_xor1), .fa_or0(s_wallace_cska32_fa759_or0));
  ha ha_s_wallace_cska32_ha19_out(.a(s_wallace_cska32_fa690_xor1[0]), .b(s_wallace_cska32_fa715_xor1[0]), .ha_xor0(s_wallace_cska32_ha19_xor0), .ha_and0(s_wallace_cska32_ha19_and0));
  fa fa_s_wallace_cska32_fa760_out(.a(s_wallace_cska32_ha19_and0[0]), .b(s_wallace_cska32_fa664_xor1[0]), .cin(s_wallace_cska32_fa691_xor1[0]), .fa_xor1(s_wallace_cska32_fa760_xor1), .fa_or0(s_wallace_cska32_fa760_or0));
  fa fa_s_wallace_cska32_fa761_out(.a(s_wallace_cska32_fa760_or0[0]), .b(s_wallace_cska32_fa636_xor1[0]), .cin(s_wallace_cska32_fa665_xor1[0]), .fa_xor1(s_wallace_cska32_fa761_xor1), .fa_or0(s_wallace_cska32_fa761_or0));
  fa fa_s_wallace_cska32_fa762_out(.a(s_wallace_cska32_fa761_or0[0]), .b(s_wallace_cska32_fa606_xor1[0]), .cin(s_wallace_cska32_fa637_xor1[0]), .fa_xor1(s_wallace_cska32_fa762_xor1), .fa_or0(s_wallace_cska32_fa762_or0));
  fa fa_s_wallace_cska32_fa763_out(.a(s_wallace_cska32_fa762_or0[0]), .b(s_wallace_cska32_fa574_xor1[0]), .cin(s_wallace_cska32_fa607_xor1[0]), .fa_xor1(s_wallace_cska32_fa763_xor1), .fa_or0(s_wallace_cska32_fa763_or0));
  fa fa_s_wallace_cska32_fa764_out(.a(s_wallace_cska32_fa763_or0[0]), .b(s_wallace_cska32_fa540_xor1[0]), .cin(s_wallace_cska32_fa575_xor1[0]), .fa_xor1(s_wallace_cska32_fa764_xor1), .fa_or0(s_wallace_cska32_fa764_or0));
  fa fa_s_wallace_cska32_fa765_out(.a(s_wallace_cska32_fa764_or0[0]), .b(s_wallace_cska32_fa504_xor1[0]), .cin(s_wallace_cska32_fa541_xor1[0]), .fa_xor1(s_wallace_cska32_fa765_xor1), .fa_or0(s_wallace_cska32_fa765_or0));
  fa fa_s_wallace_cska32_fa766_out(.a(s_wallace_cska32_fa765_or0[0]), .b(s_wallace_cska32_fa466_xor1[0]), .cin(s_wallace_cska32_fa505_xor1[0]), .fa_xor1(s_wallace_cska32_fa766_xor1), .fa_or0(s_wallace_cska32_fa766_or0));
  fa fa_s_wallace_cska32_fa767_out(.a(s_wallace_cska32_fa766_or0[0]), .b(s_wallace_cska32_fa426_xor1[0]), .cin(s_wallace_cska32_fa467_xor1[0]), .fa_xor1(s_wallace_cska32_fa767_xor1), .fa_or0(s_wallace_cska32_fa767_or0));
  fa fa_s_wallace_cska32_fa768_out(.a(s_wallace_cska32_fa767_or0[0]), .b(s_wallace_cska32_fa384_xor1[0]), .cin(s_wallace_cska32_fa427_xor1[0]), .fa_xor1(s_wallace_cska32_fa768_xor1), .fa_or0(s_wallace_cska32_fa768_or0));
  fa fa_s_wallace_cska32_fa769_out(.a(s_wallace_cska32_fa768_or0[0]), .b(s_wallace_cska32_fa340_xor1[0]), .cin(s_wallace_cska32_fa385_xor1[0]), .fa_xor1(s_wallace_cska32_fa769_xor1), .fa_or0(s_wallace_cska32_fa769_or0));
  fa fa_s_wallace_cska32_fa770_out(.a(s_wallace_cska32_fa769_or0[0]), .b(s_wallace_cska32_fa341_xor1[0]), .cin(s_wallace_cska32_fa386_xor1[0]), .fa_xor1(s_wallace_cska32_fa770_xor1), .fa_or0(s_wallace_cska32_fa770_or0));
  fa fa_s_wallace_cska32_fa771_out(.a(s_wallace_cska32_fa770_or0[0]), .b(s_wallace_cska32_fa430_xor1[0]), .cin(s_wallace_cska32_fa471_xor1[0]), .fa_xor1(s_wallace_cska32_fa771_xor1), .fa_or0(s_wallace_cska32_fa771_or0));
  fa fa_s_wallace_cska32_fa772_out(.a(s_wallace_cska32_fa771_or0[0]), .b(s_wallace_cska32_fa472_xor1[0]), .cin(s_wallace_cska32_fa511_xor1[0]), .fa_xor1(s_wallace_cska32_fa772_xor1), .fa_or0(s_wallace_cska32_fa772_or0));
  fa fa_s_wallace_cska32_fa773_out(.a(s_wallace_cska32_fa772_or0[0]), .b(s_wallace_cska32_fa512_xor1[0]), .cin(s_wallace_cska32_fa549_xor1[0]), .fa_xor1(s_wallace_cska32_fa773_xor1), .fa_or0(s_wallace_cska32_fa773_or0));
  fa fa_s_wallace_cska32_fa774_out(.a(s_wallace_cska32_fa773_or0[0]), .b(s_wallace_cska32_fa550_xor1[0]), .cin(s_wallace_cska32_fa585_xor1[0]), .fa_xor1(s_wallace_cska32_fa774_xor1), .fa_or0(s_wallace_cska32_fa774_or0));
  fa fa_s_wallace_cska32_fa775_out(.a(s_wallace_cska32_fa774_or0[0]), .b(s_wallace_cska32_fa586_xor1[0]), .cin(s_wallace_cska32_fa619_xor1[0]), .fa_xor1(s_wallace_cska32_fa775_xor1), .fa_or0(s_wallace_cska32_fa775_or0));
  fa fa_s_wallace_cska32_fa776_out(.a(s_wallace_cska32_fa775_or0[0]), .b(s_wallace_cska32_fa620_xor1[0]), .cin(s_wallace_cska32_fa651_xor1[0]), .fa_xor1(s_wallace_cska32_fa776_xor1), .fa_or0(s_wallace_cska32_fa776_or0));
  fa fa_s_wallace_cska32_fa777_out(.a(s_wallace_cska32_fa776_or0[0]), .b(s_wallace_cska32_fa652_xor1[0]), .cin(s_wallace_cska32_fa681_xor1[0]), .fa_xor1(s_wallace_cska32_fa777_xor1), .fa_or0(s_wallace_cska32_fa777_or0));
  fa fa_s_wallace_cska32_fa778_out(.a(s_wallace_cska32_fa777_or0[0]), .b(s_wallace_cska32_fa682_xor1[0]), .cin(s_wallace_cska32_fa709_xor1[0]), .fa_xor1(s_wallace_cska32_fa778_xor1), .fa_or0(s_wallace_cska32_fa778_or0));
  fa fa_s_wallace_cska32_fa779_out(.a(s_wallace_cska32_fa778_or0[0]), .b(s_wallace_cska32_fa710_xor1[0]), .cin(s_wallace_cska32_fa735_xor1[0]), .fa_xor1(s_wallace_cska32_fa779_xor1), .fa_or0(s_wallace_cska32_fa779_or0));
  ha ha_s_wallace_cska32_ha20_out(.a(s_wallace_cska32_fa716_xor1[0]), .b(s_wallace_cska32_fa739_xor1[0]), .ha_xor0(s_wallace_cska32_ha20_xor0), .ha_and0(s_wallace_cska32_ha20_and0));
  fa fa_s_wallace_cska32_fa780_out(.a(s_wallace_cska32_ha20_and0[0]), .b(s_wallace_cska32_fa692_xor1[0]), .cin(s_wallace_cska32_fa717_xor1[0]), .fa_xor1(s_wallace_cska32_fa780_xor1), .fa_or0(s_wallace_cska32_fa780_or0));
  fa fa_s_wallace_cska32_fa781_out(.a(s_wallace_cska32_fa780_or0[0]), .b(s_wallace_cska32_fa666_xor1[0]), .cin(s_wallace_cska32_fa693_xor1[0]), .fa_xor1(s_wallace_cska32_fa781_xor1), .fa_or0(s_wallace_cska32_fa781_or0));
  fa fa_s_wallace_cska32_fa782_out(.a(s_wallace_cska32_fa781_or0[0]), .b(s_wallace_cska32_fa638_xor1[0]), .cin(s_wallace_cska32_fa667_xor1[0]), .fa_xor1(s_wallace_cska32_fa782_xor1), .fa_or0(s_wallace_cska32_fa782_or0));
  fa fa_s_wallace_cska32_fa783_out(.a(s_wallace_cska32_fa782_or0[0]), .b(s_wallace_cska32_fa608_xor1[0]), .cin(s_wallace_cska32_fa639_xor1[0]), .fa_xor1(s_wallace_cska32_fa783_xor1), .fa_or0(s_wallace_cska32_fa783_or0));
  fa fa_s_wallace_cska32_fa784_out(.a(s_wallace_cska32_fa783_or0[0]), .b(s_wallace_cska32_fa576_xor1[0]), .cin(s_wallace_cska32_fa609_xor1[0]), .fa_xor1(s_wallace_cska32_fa784_xor1), .fa_or0(s_wallace_cska32_fa784_or0));
  fa fa_s_wallace_cska32_fa785_out(.a(s_wallace_cska32_fa784_or0[0]), .b(s_wallace_cska32_fa542_xor1[0]), .cin(s_wallace_cska32_fa577_xor1[0]), .fa_xor1(s_wallace_cska32_fa785_xor1), .fa_or0(s_wallace_cska32_fa785_or0));
  fa fa_s_wallace_cska32_fa786_out(.a(s_wallace_cska32_fa785_or0[0]), .b(s_wallace_cska32_fa506_xor1[0]), .cin(s_wallace_cska32_fa543_xor1[0]), .fa_xor1(s_wallace_cska32_fa786_xor1), .fa_or0(s_wallace_cska32_fa786_or0));
  fa fa_s_wallace_cska32_fa787_out(.a(s_wallace_cska32_fa786_or0[0]), .b(s_wallace_cska32_fa468_xor1[0]), .cin(s_wallace_cska32_fa507_xor1[0]), .fa_xor1(s_wallace_cska32_fa787_xor1), .fa_or0(s_wallace_cska32_fa787_or0));
  fa fa_s_wallace_cska32_fa788_out(.a(s_wallace_cska32_fa787_or0[0]), .b(s_wallace_cska32_fa428_xor1[0]), .cin(s_wallace_cska32_fa469_xor1[0]), .fa_xor1(s_wallace_cska32_fa788_xor1), .fa_or0(s_wallace_cska32_fa788_or0));
  fa fa_s_wallace_cska32_fa789_out(.a(s_wallace_cska32_fa788_or0[0]), .b(s_wallace_cska32_fa429_xor1[0]), .cin(s_wallace_cska32_fa470_xor1[0]), .fa_xor1(s_wallace_cska32_fa789_xor1), .fa_or0(s_wallace_cska32_fa789_or0));
  fa fa_s_wallace_cska32_fa790_out(.a(s_wallace_cska32_fa789_or0[0]), .b(s_wallace_cska32_fa510_xor1[0]), .cin(s_wallace_cska32_fa547_xor1[0]), .fa_xor1(s_wallace_cska32_fa790_xor1), .fa_or0(s_wallace_cska32_fa790_or0));
  fa fa_s_wallace_cska32_fa791_out(.a(s_wallace_cska32_fa790_or0[0]), .b(s_wallace_cska32_fa548_xor1[0]), .cin(s_wallace_cska32_fa583_xor1[0]), .fa_xor1(s_wallace_cska32_fa791_xor1), .fa_or0(s_wallace_cska32_fa791_or0));
  fa fa_s_wallace_cska32_fa792_out(.a(s_wallace_cska32_fa791_or0[0]), .b(s_wallace_cska32_fa584_xor1[0]), .cin(s_wallace_cska32_fa617_xor1[0]), .fa_xor1(s_wallace_cska32_fa792_xor1), .fa_or0(s_wallace_cska32_fa792_or0));
  fa fa_s_wallace_cska32_fa793_out(.a(s_wallace_cska32_fa792_or0[0]), .b(s_wallace_cska32_fa618_xor1[0]), .cin(s_wallace_cska32_fa649_xor1[0]), .fa_xor1(s_wallace_cska32_fa793_xor1), .fa_or0(s_wallace_cska32_fa793_or0));
  fa fa_s_wallace_cska32_fa794_out(.a(s_wallace_cska32_fa793_or0[0]), .b(s_wallace_cska32_fa650_xor1[0]), .cin(s_wallace_cska32_fa679_xor1[0]), .fa_xor1(s_wallace_cska32_fa794_xor1), .fa_or0(s_wallace_cska32_fa794_or0));
  fa fa_s_wallace_cska32_fa795_out(.a(s_wallace_cska32_fa794_or0[0]), .b(s_wallace_cska32_fa680_xor1[0]), .cin(s_wallace_cska32_fa707_xor1[0]), .fa_xor1(s_wallace_cska32_fa795_xor1), .fa_or0(s_wallace_cska32_fa795_or0));
  fa fa_s_wallace_cska32_fa796_out(.a(s_wallace_cska32_fa795_or0[0]), .b(s_wallace_cska32_fa708_xor1[0]), .cin(s_wallace_cska32_fa733_xor1[0]), .fa_xor1(s_wallace_cska32_fa796_xor1), .fa_or0(s_wallace_cska32_fa796_or0));
  fa fa_s_wallace_cska32_fa797_out(.a(s_wallace_cska32_fa796_or0[0]), .b(s_wallace_cska32_fa734_xor1[0]), .cin(s_wallace_cska32_fa757_xor1[0]), .fa_xor1(s_wallace_cska32_fa797_xor1), .fa_or0(s_wallace_cska32_fa797_or0));
  ha ha_s_wallace_cska32_ha21_out(.a(s_wallace_cska32_fa740_xor1[0]), .b(s_wallace_cska32_fa761_xor1[0]), .ha_xor0(s_wallace_cska32_ha21_xor0), .ha_and0(s_wallace_cska32_ha21_and0));
  fa fa_s_wallace_cska32_fa798_out(.a(s_wallace_cska32_ha21_and0[0]), .b(s_wallace_cska32_fa718_xor1[0]), .cin(s_wallace_cska32_fa741_xor1[0]), .fa_xor1(s_wallace_cska32_fa798_xor1), .fa_or0(s_wallace_cska32_fa798_or0));
  fa fa_s_wallace_cska32_fa799_out(.a(s_wallace_cska32_fa798_or0[0]), .b(s_wallace_cska32_fa694_xor1[0]), .cin(s_wallace_cska32_fa719_xor1[0]), .fa_xor1(s_wallace_cska32_fa799_xor1), .fa_or0(s_wallace_cska32_fa799_or0));
  fa fa_s_wallace_cska32_fa800_out(.a(s_wallace_cska32_fa799_or0[0]), .b(s_wallace_cska32_fa668_xor1[0]), .cin(s_wallace_cska32_fa695_xor1[0]), .fa_xor1(s_wallace_cska32_fa800_xor1), .fa_or0(s_wallace_cska32_fa800_or0));
  fa fa_s_wallace_cska32_fa801_out(.a(s_wallace_cska32_fa800_or0[0]), .b(s_wallace_cska32_fa640_xor1[0]), .cin(s_wallace_cska32_fa669_xor1[0]), .fa_xor1(s_wallace_cska32_fa801_xor1), .fa_or0(s_wallace_cska32_fa801_or0));
  fa fa_s_wallace_cska32_fa802_out(.a(s_wallace_cska32_fa801_or0[0]), .b(s_wallace_cska32_fa610_xor1[0]), .cin(s_wallace_cska32_fa641_xor1[0]), .fa_xor1(s_wallace_cska32_fa802_xor1), .fa_or0(s_wallace_cska32_fa802_or0));
  fa fa_s_wallace_cska32_fa803_out(.a(s_wallace_cska32_fa802_or0[0]), .b(s_wallace_cska32_fa578_xor1[0]), .cin(s_wallace_cska32_fa611_xor1[0]), .fa_xor1(s_wallace_cska32_fa803_xor1), .fa_or0(s_wallace_cska32_fa803_or0));
  fa fa_s_wallace_cska32_fa804_out(.a(s_wallace_cska32_fa803_or0[0]), .b(s_wallace_cska32_fa544_xor1[0]), .cin(s_wallace_cska32_fa579_xor1[0]), .fa_xor1(s_wallace_cska32_fa804_xor1), .fa_or0(s_wallace_cska32_fa804_or0));
  fa fa_s_wallace_cska32_fa805_out(.a(s_wallace_cska32_fa804_or0[0]), .b(s_wallace_cska32_fa508_xor1[0]), .cin(s_wallace_cska32_fa545_xor1[0]), .fa_xor1(s_wallace_cska32_fa805_xor1), .fa_or0(s_wallace_cska32_fa805_or0));
  fa fa_s_wallace_cska32_fa806_out(.a(s_wallace_cska32_fa805_or0[0]), .b(s_wallace_cska32_fa509_xor1[0]), .cin(s_wallace_cska32_fa546_xor1[0]), .fa_xor1(s_wallace_cska32_fa806_xor1), .fa_or0(s_wallace_cska32_fa806_or0));
  fa fa_s_wallace_cska32_fa807_out(.a(s_wallace_cska32_fa806_or0[0]), .b(s_wallace_cska32_fa582_xor1[0]), .cin(s_wallace_cska32_fa615_xor1[0]), .fa_xor1(s_wallace_cska32_fa807_xor1), .fa_or0(s_wallace_cska32_fa807_or0));
  fa fa_s_wallace_cska32_fa808_out(.a(s_wallace_cska32_fa807_or0[0]), .b(s_wallace_cska32_fa616_xor1[0]), .cin(s_wallace_cska32_fa647_xor1[0]), .fa_xor1(s_wallace_cska32_fa808_xor1), .fa_or0(s_wallace_cska32_fa808_or0));
  fa fa_s_wallace_cska32_fa809_out(.a(s_wallace_cska32_fa808_or0[0]), .b(s_wallace_cska32_fa648_xor1[0]), .cin(s_wallace_cska32_fa677_xor1[0]), .fa_xor1(s_wallace_cska32_fa809_xor1), .fa_or0(s_wallace_cska32_fa809_or0));
  fa fa_s_wallace_cska32_fa810_out(.a(s_wallace_cska32_fa809_or0[0]), .b(s_wallace_cska32_fa678_xor1[0]), .cin(s_wallace_cska32_fa705_xor1[0]), .fa_xor1(s_wallace_cska32_fa810_xor1), .fa_or0(s_wallace_cska32_fa810_or0));
  fa fa_s_wallace_cska32_fa811_out(.a(s_wallace_cska32_fa810_or0[0]), .b(s_wallace_cska32_fa706_xor1[0]), .cin(s_wallace_cska32_fa731_xor1[0]), .fa_xor1(s_wallace_cska32_fa811_xor1), .fa_or0(s_wallace_cska32_fa811_or0));
  fa fa_s_wallace_cska32_fa812_out(.a(s_wallace_cska32_fa811_or0[0]), .b(s_wallace_cska32_fa732_xor1[0]), .cin(s_wallace_cska32_fa755_xor1[0]), .fa_xor1(s_wallace_cska32_fa812_xor1), .fa_or0(s_wallace_cska32_fa812_or0));
  fa fa_s_wallace_cska32_fa813_out(.a(s_wallace_cska32_fa812_or0[0]), .b(s_wallace_cska32_fa756_xor1[0]), .cin(s_wallace_cska32_fa777_xor1[0]), .fa_xor1(s_wallace_cska32_fa813_xor1), .fa_or0(s_wallace_cska32_fa813_or0));
  ha ha_s_wallace_cska32_ha22_out(.a(s_wallace_cska32_fa762_xor1[0]), .b(s_wallace_cska32_fa781_xor1[0]), .ha_xor0(s_wallace_cska32_ha22_xor0), .ha_and0(s_wallace_cska32_ha22_and0));
  fa fa_s_wallace_cska32_fa814_out(.a(s_wallace_cska32_ha22_and0[0]), .b(s_wallace_cska32_fa742_xor1[0]), .cin(s_wallace_cska32_fa763_xor1[0]), .fa_xor1(s_wallace_cska32_fa814_xor1), .fa_or0(s_wallace_cska32_fa814_or0));
  fa fa_s_wallace_cska32_fa815_out(.a(s_wallace_cska32_fa814_or0[0]), .b(s_wallace_cska32_fa720_xor1[0]), .cin(s_wallace_cska32_fa743_xor1[0]), .fa_xor1(s_wallace_cska32_fa815_xor1), .fa_or0(s_wallace_cska32_fa815_or0));
  fa fa_s_wallace_cska32_fa816_out(.a(s_wallace_cska32_fa815_or0[0]), .b(s_wallace_cska32_fa696_xor1[0]), .cin(s_wallace_cska32_fa721_xor1[0]), .fa_xor1(s_wallace_cska32_fa816_xor1), .fa_or0(s_wallace_cska32_fa816_or0));
  fa fa_s_wallace_cska32_fa817_out(.a(s_wallace_cska32_fa816_or0[0]), .b(s_wallace_cska32_fa670_xor1[0]), .cin(s_wallace_cska32_fa697_xor1[0]), .fa_xor1(s_wallace_cska32_fa817_xor1), .fa_or0(s_wallace_cska32_fa817_or0));
  fa fa_s_wallace_cska32_fa818_out(.a(s_wallace_cska32_fa817_or0[0]), .b(s_wallace_cska32_fa642_xor1[0]), .cin(s_wallace_cska32_fa671_xor1[0]), .fa_xor1(s_wallace_cska32_fa818_xor1), .fa_or0(s_wallace_cska32_fa818_or0));
  fa fa_s_wallace_cska32_fa819_out(.a(s_wallace_cska32_fa818_or0[0]), .b(s_wallace_cska32_fa612_xor1[0]), .cin(s_wallace_cska32_fa643_xor1[0]), .fa_xor1(s_wallace_cska32_fa819_xor1), .fa_or0(s_wallace_cska32_fa819_or0));
  fa fa_s_wallace_cska32_fa820_out(.a(s_wallace_cska32_fa819_or0[0]), .b(s_wallace_cska32_fa580_xor1[0]), .cin(s_wallace_cska32_fa613_xor1[0]), .fa_xor1(s_wallace_cska32_fa820_xor1), .fa_or0(s_wallace_cska32_fa820_or0));
  fa fa_s_wallace_cska32_fa821_out(.a(s_wallace_cska32_fa820_or0[0]), .b(s_wallace_cska32_fa581_xor1[0]), .cin(s_wallace_cska32_fa614_xor1[0]), .fa_xor1(s_wallace_cska32_fa821_xor1), .fa_or0(s_wallace_cska32_fa821_or0));
  fa fa_s_wallace_cska32_fa822_out(.a(s_wallace_cska32_fa821_or0[0]), .b(s_wallace_cska32_fa646_xor1[0]), .cin(s_wallace_cska32_fa675_xor1[0]), .fa_xor1(s_wallace_cska32_fa822_xor1), .fa_or0(s_wallace_cska32_fa822_or0));
  fa fa_s_wallace_cska32_fa823_out(.a(s_wallace_cska32_fa822_or0[0]), .b(s_wallace_cska32_fa676_xor1[0]), .cin(s_wallace_cska32_fa703_xor1[0]), .fa_xor1(s_wallace_cska32_fa823_xor1), .fa_or0(s_wallace_cska32_fa823_or0));
  fa fa_s_wallace_cska32_fa824_out(.a(s_wallace_cska32_fa823_or0[0]), .b(s_wallace_cska32_fa704_xor1[0]), .cin(s_wallace_cska32_fa729_xor1[0]), .fa_xor1(s_wallace_cska32_fa824_xor1), .fa_or0(s_wallace_cska32_fa824_or0));
  fa fa_s_wallace_cska32_fa825_out(.a(s_wallace_cska32_fa824_or0[0]), .b(s_wallace_cska32_fa730_xor1[0]), .cin(s_wallace_cska32_fa753_xor1[0]), .fa_xor1(s_wallace_cska32_fa825_xor1), .fa_or0(s_wallace_cska32_fa825_or0));
  fa fa_s_wallace_cska32_fa826_out(.a(s_wallace_cska32_fa825_or0[0]), .b(s_wallace_cska32_fa754_xor1[0]), .cin(s_wallace_cska32_fa775_xor1[0]), .fa_xor1(s_wallace_cska32_fa826_xor1), .fa_or0(s_wallace_cska32_fa826_or0));
  fa fa_s_wallace_cska32_fa827_out(.a(s_wallace_cska32_fa826_or0[0]), .b(s_wallace_cska32_fa776_xor1[0]), .cin(s_wallace_cska32_fa795_xor1[0]), .fa_xor1(s_wallace_cska32_fa827_xor1), .fa_or0(s_wallace_cska32_fa827_or0));
  ha ha_s_wallace_cska32_ha23_out(.a(s_wallace_cska32_fa782_xor1[0]), .b(s_wallace_cska32_fa799_xor1[0]), .ha_xor0(s_wallace_cska32_ha23_xor0), .ha_and0(s_wallace_cska32_ha23_and0));
  fa fa_s_wallace_cska32_fa828_out(.a(s_wallace_cska32_ha23_and0[0]), .b(s_wallace_cska32_fa764_xor1[0]), .cin(s_wallace_cska32_fa783_xor1[0]), .fa_xor1(s_wallace_cska32_fa828_xor1), .fa_or0(s_wallace_cska32_fa828_or0));
  fa fa_s_wallace_cska32_fa829_out(.a(s_wallace_cska32_fa828_or0[0]), .b(s_wallace_cska32_fa744_xor1[0]), .cin(s_wallace_cska32_fa765_xor1[0]), .fa_xor1(s_wallace_cska32_fa829_xor1), .fa_or0(s_wallace_cska32_fa829_or0));
  fa fa_s_wallace_cska32_fa830_out(.a(s_wallace_cska32_fa829_or0[0]), .b(s_wallace_cska32_fa722_xor1[0]), .cin(s_wallace_cska32_fa745_xor1[0]), .fa_xor1(s_wallace_cska32_fa830_xor1), .fa_or0(s_wallace_cska32_fa830_or0));
  fa fa_s_wallace_cska32_fa831_out(.a(s_wallace_cska32_fa830_or0[0]), .b(s_wallace_cska32_fa698_xor1[0]), .cin(s_wallace_cska32_fa723_xor1[0]), .fa_xor1(s_wallace_cska32_fa831_xor1), .fa_or0(s_wallace_cska32_fa831_or0));
  fa fa_s_wallace_cska32_fa832_out(.a(s_wallace_cska32_fa831_or0[0]), .b(s_wallace_cska32_fa672_xor1[0]), .cin(s_wallace_cska32_fa699_xor1[0]), .fa_xor1(s_wallace_cska32_fa832_xor1), .fa_or0(s_wallace_cska32_fa832_or0));
  fa fa_s_wallace_cska32_fa833_out(.a(s_wallace_cska32_fa832_or0[0]), .b(s_wallace_cska32_fa644_xor1[0]), .cin(s_wallace_cska32_fa673_xor1[0]), .fa_xor1(s_wallace_cska32_fa833_xor1), .fa_or0(s_wallace_cska32_fa833_or0));
  fa fa_s_wallace_cska32_fa834_out(.a(s_wallace_cska32_fa833_or0[0]), .b(s_wallace_cska32_fa645_xor1[0]), .cin(s_wallace_cska32_fa674_xor1[0]), .fa_xor1(s_wallace_cska32_fa834_xor1), .fa_or0(s_wallace_cska32_fa834_or0));
  fa fa_s_wallace_cska32_fa835_out(.a(s_wallace_cska32_fa834_or0[0]), .b(s_wallace_cska32_fa702_xor1[0]), .cin(s_wallace_cska32_fa727_xor1[0]), .fa_xor1(s_wallace_cska32_fa835_xor1), .fa_or0(s_wallace_cska32_fa835_or0));
  fa fa_s_wallace_cska32_fa836_out(.a(s_wallace_cska32_fa835_or0[0]), .b(s_wallace_cska32_fa728_xor1[0]), .cin(s_wallace_cska32_fa751_xor1[0]), .fa_xor1(s_wallace_cska32_fa836_xor1), .fa_or0(s_wallace_cska32_fa836_or0));
  fa fa_s_wallace_cska32_fa837_out(.a(s_wallace_cska32_fa836_or0[0]), .b(s_wallace_cska32_fa752_xor1[0]), .cin(s_wallace_cska32_fa773_xor1[0]), .fa_xor1(s_wallace_cska32_fa837_xor1), .fa_or0(s_wallace_cska32_fa837_or0));
  fa fa_s_wallace_cska32_fa838_out(.a(s_wallace_cska32_fa837_or0[0]), .b(s_wallace_cska32_fa774_xor1[0]), .cin(s_wallace_cska32_fa793_xor1[0]), .fa_xor1(s_wallace_cska32_fa838_xor1), .fa_or0(s_wallace_cska32_fa838_or0));
  fa fa_s_wallace_cska32_fa839_out(.a(s_wallace_cska32_fa838_or0[0]), .b(s_wallace_cska32_fa794_xor1[0]), .cin(s_wallace_cska32_fa811_xor1[0]), .fa_xor1(s_wallace_cska32_fa839_xor1), .fa_or0(s_wallace_cska32_fa839_or0));
  ha ha_s_wallace_cska32_ha24_out(.a(s_wallace_cska32_fa800_xor1[0]), .b(s_wallace_cska32_fa815_xor1[0]), .ha_xor0(s_wallace_cska32_ha24_xor0), .ha_and0(s_wallace_cska32_ha24_and0));
  fa fa_s_wallace_cska32_fa840_out(.a(s_wallace_cska32_ha24_and0[0]), .b(s_wallace_cska32_fa784_xor1[0]), .cin(s_wallace_cska32_fa801_xor1[0]), .fa_xor1(s_wallace_cska32_fa840_xor1), .fa_or0(s_wallace_cska32_fa840_or0));
  fa fa_s_wallace_cska32_fa841_out(.a(s_wallace_cska32_fa840_or0[0]), .b(s_wallace_cska32_fa766_xor1[0]), .cin(s_wallace_cska32_fa785_xor1[0]), .fa_xor1(s_wallace_cska32_fa841_xor1), .fa_or0(s_wallace_cska32_fa841_or0));
  fa fa_s_wallace_cska32_fa842_out(.a(s_wallace_cska32_fa841_or0[0]), .b(s_wallace_cska32_fa746_xor1[0]), .cin(s_wallace_cska32_fa767_xor1[0]), .fa_xor1(s_wallace_cska32_fa842_xor1), .fa_or0(s_wallace_cska32_fa842_or0));
  fa fa_s_wallace_cska32_fa843_out(.a(s_wallace_cska32_fa842_or0[0]), .b(s_wallace_cska32_fa724_xor1[0]), .cin(s_wallace_cska32_fa747_xor1[0]), .fa_xor1(s_wallace_cska32_fa843_xor1), .fa_or0(s_wallace_cska32_fa843_or0));
  fa fa_s_wallace_cska32_fa844_out(.a(s_wallace_cska32_fa843_or0[0]), .b(s_wallace_cska32_fa700_xor1[0]), .cin(s_wallace_cska32_fa725_xor1[0]), .fa_xor1(s_wallace_cska32_fa844_xor1), .fa_or0(s_wallace_cska32_fa844_or0));
  fa fa_s_wallace_cska32_fa845_out(.a(s_wallace_cska32_fa844_or0[0]), .b(s_wallace_cska32_fa701_xor1[0]), .cin(s_wallace_cska32_fa726_xor1[0]), .fa_xor1(s_wallace_cska32_fa845_xor1), .fa_or0(s_wallace_cska32_fa845_or0));
  fa fa_s_wallace_cska32_fa846_out(.a(s_wallace_cska32_fa845_or0[0]), .b(s_wallace_cska32_fa750_xor1[0]), .cin(s_wallace_cska32_fa771_xor1[0]), .fa_xor1(s_wallace_cska32_fa846_xor1), .fa_or0(s_wallace_cska32_fa846_or0));
  fa fa_s_wallace_cska32_fa847_out(.a(s_wallace_cska32_fa846_or0[0]), .b(s_wallace_cska32_fa772_xor1[0]), .cin(s_wallace_cska32_fa791_xor1[0]), .fa_xor1(s_wallace_cska32_fa847_xor1), .fa_or0(s_wallace_cska32_fa847_or0));
  fa fa_s_wallace_cska32_fa848_out(.a(s_wallace_cska32_fa847_or0[0]), .b(s_wallace_cska32_fa792_xor1[0]), .cin(s_wallace_cska32_fa809_xor1[0]), .fa_xor1(s_wallace_cska32_fa848_xor1), .fa_or0(s_wallace_cska32_fa848_or0));
  fa fa_s_wallace_cska32_fa849_out(.a(s_wallace_cska32_fa848_or0[0]), .b(s_wallace_cska32_fa810_xor1[0]), .cin(s_wallace_cska32_fa825_xor1[0]), .fa_xor1(s_wallace_cska32_fa849_xor1), .fa_or0(s_wallace_cska32_fa849_or0));
  ha ha_s_wallace_cska32_ha25_out(.a(s_wallace_cska32_fa816_xor1[0]), .b(s_wallace_cska32_fa829_xor1[0]), .ha_xor0(s_wallace_cska32_ha25_xor0), .ha_and0(s_wallace_cska32_ha25_and0));
  fa fa_s_wallace_cska32_fa850_out(.a(s_wallace_cska32_ha25_and0[0]), .b(s_wallace_cska32_fa802_xor1[0]), .cin(s_wallace_cska32_fa817_xor1[0]), .fa_xor1(s_wallace_cska32_fa850_xor1), .fa_or0(s_wallace_cska32_fa850_or0));
  fa fa_s_wallace_cska32_fa851_out(.a(s_wallace_cska32_fa850_or0[0]), .b(s_wallace_cska32_fa786_xor1[0]), .cin(s_wallace_cska32_fa803_xor1[0]), .fa_xor1(s_wallace_cska32_fa851_xor1), .fa_or0(s_wallace_cska32_fa851_or0));
  fa fa_s_wallace_cska32_fa852_out(.a(s_wallace_cska32_fa851_or0[0]), .b(s_wallace_cska32_fa768_xor1[0]), .cin(s_wallace_cska32_fa787_xor1[0]), .fa_xor1(s_wallace_cska32_fa852_xor1), .fa_or0(s_wallace_cska32_fa852_or0));
  fa fa_s_wallace_cska32_fa853_out(.a(s_wallace_cska32_fa852_or0[0]), .b(s_wallace_cska32_fa748_xor1[0]), .cin(s_wallace_cska32_fa769_xor1[0]), .fa_xor1(s_wallace_cska32_fa853_xor1), .fa_or0(s_wallace_cska32_fa853_or0));
  fa fa_s_wallace_cska32_fa854_out(.a(s_wallace_cska32_fa853_or0[0]), .b(s_wallace_cska32_fa749_xor1[0]), .cin(s_wallace_cska32_fa770_xor1[0]), .fa_xor1(s_wallace_cska32_fa854_xor1), .fa_or0(s_wallace_cska32_fa854_or0));
  fa fa_s_wallace_cska32_fa855_out(.a(s_wallace_cska32_fa854_or0[0]), .b(s_wallace_cska32_fa790_xor1[0]), .cin(s_wallace_cska32_fa807_xor1[0]), .fa_xor1(s_wallace_cska32_fa855_xor1), .fa_or0(s_wallace_cska32_fa855_or0));
  fa fa_s_wallace_cska32_fa856_out(.a(s_wallace_cska32_fa855_or0[0]), .b(s_wallace_cska32_fa808_xor1[0]), .cin(s_wallace_cska32_fa823_xor1[0]), .fa_xor1(s_wallace_cska32_fa856_xor1), .fa_or0(s_wallace_cska32_fa856_or0));
  fa fa_s_wallace_cska32_fa857_out(.a(s_wallace_cska32_fa856_or0[0]), .b(s_wallace_cska32_fa824_xor1[0]), .cin(s_wallace_cska32_fa837_xor1[0]), .fa_xor1(s_wallace_cska32_fa857_xor1), .fa_or0(s_wallace_cska32_fa857_or0));
  ha ha_s_wallace_cska32_ha26_out(.a(s_wallace_cska32_fa830_xor1[0]), .b(s_wallace_cska32_fa841_xor1[0]), .ha_xor0(s_wallace_cska32_ha26_xor0), .ha_and0(s_wallace_cska32_ha26_and0));
  fa fa_s_wallace_cska32_fa858_out(.a(s_wallace_cska32_ha26_and0[0]), .b(s_wallace_cska32_fa818_xor1[0]), .cin(s_wallace_cska32_fa831_xor1[0]), .fa_xor1(s_wallace_cska32_fa858_xor1), .fa_or0(s_wallace_cska32_fa858_or0));
  fa fa_s_wallace_cska32_fa859_out(.a(s_wallace_cska32_fa858_or0[0]), .b(s_wallace_cska32_fa804_xor1[0]), .cin(s_wallace_cska32_fa819_xor1[0]), .fa_xor1(s_wallace_cska32_fa859_xor1), .fa_or0(s_wallace_cska32_fa859_or0));
  fa fa_s_wallace_cska32_fa860_out(.a(s_wallace_cska32_fa859_or0[0]), .b(s_wallace_cska32_fa788_xor1[0]), .cin(s_wallace_cska32_fa805_xor1[0]), .fa_xor1(s_wallace_cska32_fa860_xor1), .fa_or0(s_wallace_cska32_fa860_or0));
  fa fa_s_wallace_cska32_fa861_out(.a(s_wallace_cska32_fa860_or0[0]), .b(s_wallace_cska32_fa789_xor1[0]), .cin(s_wallace_cska32_fa806_xor1[0]), .fa_xor1(s_wallace_cska32_fa861_xor1), .fa_or0(s_wallace_cska32_fa861_or0));
  fa fa_s_wallace_cska32_fa862_out(.a(s_wallace_cska32_fa861_or0[0]), .b(s_wallace_cska32_fa822_xor1[0]), .cin(s_wallace_cska32_fa835_xor1[0]), .fa_xor1(s_wallace_cska32_fa862_xor1), .fa_or0(s_wallace_cska32_fa862_or0));
  fa fa_s_wallace_cska32_fa863_out(.a(s_wallace_cska32_fa862_or0[0]), .b(s_wallace_cska32_fa836_xor1[0]), .cin(s_wallace_cska32_fa847_xor1[0]), .fa_xor1(s_wallace_cska32_fa863_xor1), .fa_or0(s_wallace_cska32_fa863_or0));
  ha ha_s_wallace_cska32_ha27_out(.a(s_wallace_cska32_fa842_xor1[0]), .b(s_wallace_cska32_fa851_xor1[0]), .ha_xor0(s_wallace_cska32_ha27_xor0), .ha_and0(s_wallace_cska32_ha27_and0));
  fa fa_s_wallace_cska32_fa864_out(.a(s_wallace_cska32_ha27_and0[0]), .b(s_wallace_cska32_fa832_xor1[0]), .cin(s_wallace_cska32_fa843_xor1[0]), .fa_xor1(s_wallace_cska32_fa864_xor1), .fa_or0(s_wallace_cska32_fa864_or0));
  fa fa_s_wallace_cska32_fa865_out(.a(s_wallace_cska32_fa864_or0[0]), .b(s_wallace_cska32_fa820_xor1[0]), .cin(s_wallace_cska32_fa833_xor1[0]), .fa_xor1(s_wallace_cska32_fa865_xor1), .fa_or0(s_wallace_cska32_fa865_or0));
  fa fa_s_wallace_cska32_fa866_out(.a(s_wallace_cska32_fa865_or0[0]), .b(s_wallace_cska32_fa821_xor1[0]), .cin(s_wallace_cska32_fa834_xor1[0]), .fa_xor1(s_wallace_cska32_fa866_xor1), .fa_or0(s_wallace_cska32_fa866_or0));
  fa fa_s_wallace_cska32_fa867_out(.a(s_wallace_cska32_fa866_or0[0]), .b(s_wallace_cska32_fa846_xor1[0]), .cin(s_wallace_cska32_fa855_xor1[0]), .fa_xor1(s_wallace_cska32_fa867_xor1), .fa_or0(s_wallace_cska32_fa867_or0));
  ha ha_s_wallace_cska32_ha28_out(.a(s_wallace_cska32_fa852_xor1[0]), .b(s_wallace_cska32_fa859_xor1[0]), .ha_xor0(s_wallace_cska32_ha28_xor0), .ha_and0(s_wallace_cska32_ha28_and0));
  fa fa_s_wallace_cska32_fa868_out(.a(s_wallace_cska32_ha28_and0[0]), .b(s_wallace_cska32_fa844_xor1[0]), .cin(s_wallace_cska32_fa853_xor1[0]), .fa_xor1(s_wallace_cska32_fa868_xor1), .fa_or0(s_wallace_cska32_fa868_or0));
  fa fa_s_wallace_cska32_fa869_out(.a(s_wallace_cska32_fa868_or0[0]), .b(s_wallace_cska32_fa845_xor1[0]), .cin(s_wallace_cska32_fa854_xor1[0]), .fa_xor1(s_wallace_cska32_fa869_xor1), .fa_or0(s_wallace_cska32_fa869_or0));
  ha ha_s_wallace_cska32_ha29_out(.a(s_wallace_cska32_fa860_xor1[0]), .b(s_wallace_cska32_fa865_xor1[0]), .ha_xor0(s_wallace_cska32_ha29_xor0), .ha_and0(s_wallace_cska32_ha29_and0));
  fa fa_s_wallace_cska32_fa870_out(.a(s_wallace_cska32_ha29_and0[0]), .b(s_wallace_cska32_fa861_xor1[0]), .cin(s_wallace_cska32_fa866_xor1[0]), .fa_xor1(s_wallace_cska32_fa870_xor1), .fa_or0(s_wallace_cska32_fa870_or0));
  fa fa_s_wallace_cska32_fa871_out(.a(s_wallace_cska32_fa870_or0[0]), .b(s_wallace_cska32_fa869_or0[0]), .cin(s_wallace_cska32_fa862_xor1[0]), .fa_xor1(s_wallace_cska32_fa871_xor1), .fa_or0(s_wallace_cska32_fa871_or0));
  fa fa_s_wallace_cska32_fa872_out(.a(s_wallace_cska32_fa871_or0[0]), .b(s_wallace_cska32_fa867_or0[0]), .cin(s_wallace_cska32_fa856_xor1[0]), .fa_xor1(s_wallace_cska32_fa872_xor1), .fa_or0(s_wallace_cska32_fa872_or0));
  fa fa_s_wallace_cska32_fa873_out(.a(s_wallace_cska32_fa872_or0[0]), .b(s_wallace_cska32_fa863_or0[0]), .cin(s_wallace_cska32_fa848_xor1[0]), .fa_xor1(s_wallace_cska32_fa873_xor1), .fa_or0(s_wallace_cska32_fa873_or0));
  fa fa_s_wallace_cska32_fa874_out(.a(s_wallace_cska32_fa873_or0[0]), .b(s_wallace_cska32_fa857_or0[0]), .cin(s_wallace_cska32_fa838_xor1[0]), .fa_xor1(s_wallace_cska32_fa874_xor1), .fa_or0(s_wallace_cska32_fa874_or0));
  fa fa_s_wallace_cska32_fa875_out(.a(s_wallace_cska32_fa874_or0[0]), .b(s_wallace_cska32_fa849_or0[0]), .cin(s_wallace_cska32_fa826_xor1[0]), .fa_xor1(s_wallace_cska32_fa875_xor1), .fa_or0(s_wallace_cska32_fa875_or0));
  fa fa_s_wallace_cska32_fa876_out(.a(s_wallace_cska32_fa875_or0[0]), .b(s_wallace_cska32_fa839_or0[0]), .cin(s_wallace_cska32_fa812_xor1[0]), .fa_xor1(s_wallace_cska32_fa876_xor1), .fa_or0(s_wallace_cska32_fa876_or0));
  fa fa_s_wallace_cska32_fa877_out(.a(s_wallace_cska32_fa876_or0[0]), .b(s_wallace_cska32_fa827_or0[0]), .cin(s_wallace_cska32_fa796_xor1[0]), .fa_xor1(s_wallace_cska32_fa877_xor1), .fa_or0(s_wallace_cska32_fa877_or0));
  fa fa_s_wallace_cska32_fa878_out(.a(s_wallace_cska32_fa877_or0[0]), .b(s_wallace_cska32_fa813_or0[0]), .cin(s_wallace_cska32_fa778_xor1[0]), .fa_xor1(s_wallace_cska32_fa878_xor1), .fa_or0(s_wallace_cska32_fa878_or0));
  fa fa_s_wallace_cska32_fa879_out(.a(s_wallace_cska32_fa878_or0[0]), .b(s_wallace_cska32_fa797_or0[0]), .cin(s_wallace_cska32_fa758_xor1[0]), .fa_xor1(s_wallace_cska32_fa879_xor1), .fa_or0(s_wallace_cska32_fa879_or0));
  fa fa_s_wallace_cska32_fa880_out(.a(s_wallace_cska32_fa879_or0[0]), .b(s_wallace_cska32_fa779_or0[0]), .cin(s_wallace_cska32_fa736_xor1[0]), .fa_xor1(s_wallace_cska32_fa880_xor1), .fa_or0(s_wallace_cska32_fa880_or0));
  fa fa_s_wallace_cska32_fa881_out(.a(s_wallace_cska32_fa880_or0[0]), .b(s_wallace_cska32_fa759_or0[0]), .cin(s_wallace_cska32_fa712_xor1[0]), .fa_xor1(s_wallace_cska32_fa881_xor1), .fa_or0(s_wallace_cska32_fa881_or0));
  fa fa_s_wallace_cska32_fa882_out(.a(s_wallace_cska32_fa881_or0[0]), .b(s_wallace_cska32_fa737_or0[0]), .cin(s_wallace_cska32_fa686_xor1[0]), .fa_xor1(s_wallace_cska32_fa882_xor1), .fa_or0(s_wallace_cska32_fa882_or0));
  fa fa_s_wallace_cska32_fa883_out(.a(s_wallace_cska32_fa882_or0[0]), .b(s_wallace_cska32_fa713_or0[0]), .cin(s_wallace_cska32_fa658_xor1[0]), .fa_xor1(s_wallace_cska32_fa883_xor1), .fa_or0(s_wallace_cska32_fa883_or0));
  fa fa_s_wallace_cska32_fa884_out(.a(s_wallace_cska32_fa883_or0[0]), .b(s_wallace_cska32_fa687_or0[0]), .cin(s_wallace_cska32_fa628_xor1[0]), .fa_xor1(s_wallace_cska32_fa884_xor1), .fa_or0(s_wallace_cska32_fa884_or0));
  fa fa_s_wallace_cska32_fa885_out(.a(s_wallace_cska32_fa884_or0[0]), .b(s_wallace_cska32_fa659_or0[0]), .cin(s_wallace_cska32_fa596_xor1[0]), .fa_xor1(s_wallace_cska32_fa885_xor1), .fa_or0(s_wallace_cska32_fa885_or0));
  fa fa_s_wallace_cska32_fa886_out(.a(s_wallace_cska32_fa885_or0[0]), .b(s_wallace_cska32_fa629_or0[0]), .cin(s_wallace_cska32_fa562_xor1[0]), .fa_xor1(s_wallace_cska32_fa886_xor1), .fa_or0(s_wallace_cska32_fa886_or0));
  fa fa_s_wallace_cska32_fa887_out(.a(s_wallace_cska32_fa886_or0[0]), .b(s_wallace_cska32_fa597_or0[0]), .cin(s_wallace_cska32_fa526_xor1[0]), .fa_xor1(s_wallace_cska32_fa887_xor1), .fa_or0(s_wallace_cska32_fa887_or0));
  fa fa_s_wallace_cska32_fa888_out(.a(s_wallace_cska32_fa887_or0[0]), .b(s_wallace_cska32_fa563_or0[0]), .cin(s_wallace_cska32_fa488_xor1[0]), .fa_xor1(s_wallace_cska32_fa888_xor1), .fa_or0(s_wallace_cska32_fa888_or0));
  fa fa_s_wallace_cska32_fa889_out(.a(s_wallace_cska32_fa888_or0[0]), .b(s_wallace_cska32_fa527_or0[0]), .cin(s_wallace_cska32_fa448_xor1[0]), .fa_xor1(s_wallace_cska32_fa889_xor1), .fa_or0(s_wallace_cska32_fa889_or0));
  fa fa_s_wallace_cska32_fa890_out(.a(s_wallace_cska32_fa889_or0[0]), .b(s_wallace_cska32_fa489_or0[0]), .cin(s_wallace_cska32_fa406_xor1[0]), .fa_xor1(s_wallace_cska32_fa890_xor1), .fa_or0(s_wallace_cska32_fa890_or0));
  fa fa_s_wallace_cska32_fa891_out(.a(s_wallace_cska32_fa890_or0[0]), .b(s_wallace_cska32_fa449_or0[0]), .cin(s_wallace_cska32_fa362_xor1[0]), .fa_xor1(s_wallace_cska32_fa891_xor1), .fa_or0(s_wallace_cska32_fa891_or0));
  fa fa_s_wallace_cska32_fa892_out(.a(s_wallace_cska32_fa891_or0[0]), .b(s_wallace_cska32_fa407_or0[0]), .cin(s_wallace_cska32_fa316_xor1[0]), .fa_xor1(s_wallace_cska32_fa892_xor1), .fa_or0(s_wallace_cska32_fa892_or0));
  fa fa_s_wallace_cska32_fa893_out(.a(s_wallace_cska32_fa892_or0[0]), .b(s_wallace_cska32_fa363_or0[0]), .cin(s_wallace_cska32_fa268_xor1[0]), .fa_xor1(s_wallace_cska32_fa893_xor1), .fa_or0(s_wallace_cska32_fa893_or0));
  fa fa_s_wallace_cska32_fa894_out(.a(s_wallace_cska32_fa893_or0[0]), .b(s_wallace_cska32_fa317_or0[0]), .cin(s_wallace_cska32_fa218_xor1[0]), .fa_xor1(s_wallace_cska32_fa894_xor1), .fa_or0(s_wallace_cska32_fa894_or0));
  fa fa_s_wallace_cska32_fa895_out(.a(s_wallace_cska32_fa894_or0[0]), .b(s_wallace_cska32_fa269_or0[0]), .cin(s_wallace_cska32_fa166_xor1[0]), .fa_xor1(s_wallace_cska32_fa895_xor1), .fa_or0(s_wallace_cska32_fa895_or0));
  fa fa_s_wallace_cska32_fa896_out(.a(s_wallace_cska32_fa895_or0[0]), .b(s_wallace_cska32_fa219_or0[0]), .cin(s_wallace_cska32_fa112_xor1[0]), .fa_xor1(s_wallace_cska32_fa896_xor1), .fa_or0(s_wallace_cska32_fa896_or0));
  fa fa_s_wallace_cska32_fa897_out(.a(s_wallace_cska32_fa896_or0[0]), .b(s_wallace_cska32_fa167_or0[0]), .cin(s_wallace_cska32_fa56_xor1[0]), .fa_xor1(s_wallace_cska32_fa897_xor1), .fa_or0(s_wallace_cska32_fa897_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_29_31(.a(a[29]), .b(b[31]), .out(s_wallace_cska32_nand_29_31));
  fa fa_s_wallace_cska32_fa898_out(.a(s_wallace_cska32_fa897_or0[0]), .b(s_wallace_cska32_fa113_or0[0]), .cin(s_wallace_cska32_nand_29_31[0]), .fa_xor1(s_wallace_cska32_fa898_xor1), .fa_or0(s_wallace_cska32_fa898_or0));
  nand_gate nand_gate_s_wallace_cska32_nand_31_30(.a(a[31]), .b(b[30]), .out(s_wallace_cska32_nand_31_30));
  fa fa_s_wallace_cska32_fa899_out(.a(s_wallace_cska32_fa898_or0[0]), .b(s_wallace_cska32_fa57_or0[0]), .cin(s_wallace_cska32_nand_31_30[0]), .fa_xor1(s_wallace_cska32_fa899_xor1), .fa_or0(s_wallace_cska32_fa899_or0));
  and_gate and_gate_s_wallace_cska32_and_0_0(.a(a[0]), .b(b[0]), .out(s_wallace_cska32_and_0_0));
  and_gate and_gate_s_wallace_cska32_and_1_0(.a(a[1]), .b(b[0]), .out(s_wallace_cska32_and_1_0));
  and_gate and_gate_s_wallace_cska32_and_0_2(.a(a[0]), .b(b[2]), .out(s_wallace_cska32_and_0_2));
  nand_gate nand_gate_s_wallace_cska32_nand_30_31(.a(a[30]), .b(b[31]), .out(s_wallace_cska32_nand_30_31));
  and_gate and_gate_s_wallace_cska32_and_0_1(.a(a[0]), .b(b[1]), .out(s_wallace_cska32_and_0_1));
  and_gate and_gate_s_wallace_cska32_and_31_31(.a(a[31]), .b(b[31]), .out(s_wallace_cska32_and_31_31));
  assign s_wallace_cska32_u_cska62_a[0] = s_wallace_cska32_and_1_0[0];
  assign s_wallace_cska32_u_cska62_a[1] = s_wallace_cska32_and_0_2[0];
  assign s_wallace_cska32_u_cska62_a[2] = s_wallace_cska32_fa0_xor1[0];
  assign s_wallace_cska32_u_cska62_a[3] = s_wallace_cska32_fa58_xor1[0];
  assign s_wallace_cska32_u_cska62_a[4] = s_wallace_cska32_fa114_xor1[0];
  assign s_wallace_cska32_u_cska62_a[5] = s_wallace_cska32_fa168_xor1[0];
  assign s_wallace_cska32_u_cska62_a[6] = s_wallace_cska32_fa220_xor1[0];
  assign s_wallace_cska32_u_cska62_a[7] = s_wallace_cska32_fa270_xor1[0];
  assign s_wallace_cska32_u_cska62_a[8] = s_wallace_cska32_fa318_xor1[0];
  assign s_wallace_cska32_u_cska62_a[9] = s_wallace_cska32_fa364_xor1[0];
  assign s_wallace_cska32_u_cska62_a[10] = s_wallace_cska32_fa408_xor1[0];
  assign s_wallace_cska32_u_cska62_a[11] = s_wallace_cska32_fa450_xor1[0];
  assign s_wallace_cska32_u_cska62_a[12] = s_wallace_cska32_fa490_xor1[0];
  assign s_wallace_cska32_u_cska62_a[13] = s_wallace_cska32_fa528_xor1[0];
  assign s_wallace_cska32_u_cska62_a[14] = s_wallace_cska32_fa564_xor1[0];
  assign s_wallace_cska32_u_cska62_a[15] = s_wallace_cska32_fa598_xor1[0];
  assign s_wallace_cska32_u_cska62_a[16] = s_wallace_cska32_fa630_xor1[0];
  assign s_wallace_cska32_u_cska62_a[17] = s_wallace_cska32_fa660_xor1[0];
  assign s_wallace_cska32_u_cska62_a[18] = s_wallace_cska32_fa688_xor1[0];
  assign s_wallace_cska32_u_cska62_a[19] = s_wallace_cska32_fa714_xor1[0];
  assign s_wallace_cska32_u_cska62_a[20] = s_wallace_cska32_fa738_xor1[0];
  assign s_wallace_cska32_u_cska62_a[21] = s_wallace_cska32_fa760_xor1[0];
  assign s_wallace_cska32_u_cska62_a[22] = s_wallace_cska32_fa780_xor1[0];
  assign s_wallace_cska32_u_cska62_a[23] = s_wallace_cska32_fa798_xor1[0];
  assign s_wallace_cska32_u_cska62_a[24] = s_wallace_cska32_fa814_xor1[0];
  assign s_wallace_cska32_u_cska62_a[25] = s_wallace_cska32_fa828_xor1[0];
  assign s_wallace_cska32_u_cska62_a[26] = s_wallace_cska32_fa840_xor1[0];
  assign s_wallace_cska32_u_cska62_a[27] = s_wallace_cska32_fa850_xor1[0];
  assign s_wallace_cska32_u_cska62_a[28] = s_wallace_cska32_fa858_xor1[0];
  assign s_wallace_cska32_u_cska62_a[29] = s_wallace_cska32_fa864_xor1[0];
  assign s_wallace_cska32_u_cska62_a[30] = s_wallace_cska32_fa868_xor1[0];
  assign s_wallace_cska32_u_cska62_a[31] = s_wallace_cska32_fa869_xor1[0];
  assign s_wallace_cska32_u_cska62_a[32] = s_wallace_cska32_fa867_xor1[0];
  assign s_wallace_cska32_u_cska62_a[33] = s_wallace_cska32_fa863_xor1[0];
  assign s_wallace_cska32_u_cska62_a[34] = s_wallace_cska32_fa857_xor1[0];
  assign s_wallace_cska32_u_cska62_a[35] = s_wallace_cska32_fa849_xor1[0];
  assign s_wallace_cska32_u_cska62_a[36] = s_wallace_cska32_fa839_xor1[0];
  assign s_wallace_cska32_u_cska62_a[37] = s_wallace_cska32_fa827_xor1[0];
  assign s_wallace_cska32_u_cska62_a[38] = s_wallace_cska32_fa813_xor1[0];
  assign s_wallace_cska32_u_cska62_a[39] = s_wallace_cska32_fa797_xor1[0];
  assign s_wallace_cska32_u_cska62_a[40] = s_wallace_cska32_fa779_xor1[0];
  assign s_wallace_cska32_u_cska62_a[41] = s_wallace_cska32_fa759_xor1[0];
  assign s_wallace_cska32_u_cska62_a[42] = s_wallace_cska32_fa737_xor1[0];
  assign s_wallace_cska32_u_cska62_a[43] = s_wallace_cska32_fa713_xor1[0];
  assign s_wallace_cska32_u_cska62_a[44] = s_wallace_cska32_fa687_xor1[0];
  assign s_wallace_cska32_u_cska62_a[45] = s_wallace_cska32_fa659_xor1[0];
  assign s_wallace_cska32_u_cska62_a[46] = s_wallace_cska32_fa629_xor1[0];
  assign s_wallace_cska32_u_cska62_a[47] = s_wallace_cska32_fa597_xor1[0];
  assign s_wallace_cska32_u_cska62_a[48] = s_wallace_cska32_fa563_xor1[0];
  assign s_wallace_cska32_u_cska62_a[49] = s_wallace_cska32_fa527_xor1[0];
  assign s_wallace_cska32_u_cska62_a[50] = s_wallace_cska32_fa489_xor1[0];
  assign s_wallace_cska32_u_cska62_a[51] = s_wallace_cska32_fa449_xor1[0];
  assign s_wallace_cska32_u_cska62_a[52] = s_wallace_cska32_fa407_xor1[0];
  assign s_wallace_cska32_u_cska62_a[53] = s_wallace_cska32_fa363_xor1[0];
  assign s_wallace_cska32_u_cska62_a[54] = s_wallace_cska32_fa317_xor1[0];
  assign s_wallace_cska32_u_cska62_a[55] = s_wallace_cska32_fa269_xor1[0];
  assign s_wallace_cska32_u_cska62_a[56] = s_wallace_cska32_fa219_xor1[0];
  assign s_wallace_cska32_u_cska62_a[57] = s_wallace_cska32_fa167_xor1[0];
  assign s_wallace_cska32_u_cska62_a[58] = s_wallace_cska32_fa113_xor1[0];
  assign s_wallace_cska32_u_cska62_a[59] = s_wallace_cska32_fa57_xor1[0];
  assign s_wallace_cska32_u_cska62_a[60] = s_wallace_cska32_nand_30_31[0];
  assign s_wallace_cska32_u_cska62_a[61] = s_wallace_cska32_fa899_or0[0];
  assign s_wallace_cska32_u_cska62_b[0] = s_wallace_cska32_and_0_1[0];
  assign s_wallace_cska32_u_cska62_b[1] = s_wallace_cska32_ha0_xor0[0];
  assign s_wallace_cska32_u_cska62_b[2] = s_wallace_cska32_ha1_xor0[0];
  assign s_wallace_cska32_u_cska62_b[3] = s_wallace_cska32_ha2_xor0[0];
  assign s_wallace_cska32_u_cska62_b[4] = s_wallace_cska32_ha3_xor0[0];
  assign s_wallace_cska32_u_cska62_b[5] = s_wallace_cska32_ha4_xor0[0];
  assign s_wallace_cska32_u_cska62_b[6] = s_wallace_cska32_ha5_xor0[0];
  assign s_wallace_cska32_u_cska62_b[7] = s_wallace_cska32_ha6_xor0[0];
  assign s_wallace_cska32_u_cska62_b[8] = s_wallace_cska32_ha7_xor0[0];
  assign s_wallace_cska32_u_cska62_b[9] = s_wallace_cska32_ha8_xor0[0];
  assign s_wallace_cska32_u_cska62_b[10] = s_wallace_cska32_ha9_xor0[0];
  assign s_wallace_cska32_u_cska62_b[11] = s_wallace_cska32_ha10_xor0[0];
  assign s_wallace_cska32_u_cska62_b[12] = s_wallace_cska32_ha11_xor0[0];
  assign s_wallace_cska32_u_cska62_b[13] = s_wallace_cska32_ha12_xor0[0];
  assign s_wallace_cska32_u_cska62_b[14] = s_wallace_cska32_ha13_xor0[0];
  assign s_wallace_cska32_u_cska62_b[15] = s_wallace_cska32_ha14_xor0[0];
  assign s_wallace_cska32_u_cska62_b[16] = s_wallace_cska32_ha15_xor0[0];
  assign s_wallace_cska32_u_cska62_b[17] = s_wallace_cska32_ha16_xor0[0];
  assign s_wallace_cska32_u_cska62_b[18] = s_wallace_cska32_ha17_xor0[0];
  assign s_wallace_cska32_u_cska62_b[19] = s_wallace_cska32_ha18_xor0[0];
  assign s_wallace_cska32_u_cska62_b[20] = s_wallace_cska32_ha19_xor0[0];
  assign s_wallace_cska32_u_cska62_b[21] = s_wallace_cska32_ha20_xor0[0];
  assign s_wallace_cska32_u_cska62_b[22] = s_wallace_cska32_ha21_xor0[0];
  assign s_wallace_cska32_u_cska62_b[23] = s_wallace_cska32_ha22_xor0[0];
  assign s_wallace_cska32_u_cska62_b[24] = s_wallace_cska32_ha23_xor0[0];
  assign s_wallace_cska32_u_cska62_b[25] = s_wallace_cska32_ha24_xor0[0];
  assign s_wallace_cska32_u_cska62_b[26] = s_wallace_cska32_ha25_xor0[0];
  assign s_wallace_cska32_u_cska62_b[27] = s_wallace_cska32_ha26_xor0[0];
  assign s_wallace_cska32_u_cska62_b[28] = s_wallace_cska32_ha27_xor0[0];
  assign s_wallace_cska32_u_cska62_b[29] = s_wallace_cska32_ha28_xor0[0];
  assign s_wallace_cska32_u_cska62_b[30] = s_wallace_cska32_ha29_xor0[0];
  assign s_wallace_cska32_u_cska62_b[31] = s_wallace_cska32_fa870_xor1[0];
  assign s_wallace_cska32_u_cska62_b[32] = s_wallace_cska32_fa871_xor1[0];
  assign s_wallace_cska32_u_cska62_b[33] = s_wallace_cska32_fa872_xor1[0];
  assign s_wallace_cska32_u_cska62_b[34] = s_wallace_cska32_fa873_xor1[0];
  assign s_wallace_cska32_u_cska62_b[35] = s_wallace_cska32_fa874_xor1[0];
  assign s_wallace_cska32_u_cska62_b[36] = s_wallace_cska32_fa875_xor1[0];
  assign s_wallace_cska32_u_cska62_b[37] = s_wallace_cska32_fa876_xor1[0];
  assign s_wallace_cska32_u_cska62_b[38] = s_wallace_cska32_fa877_xor1[0];
  assign s_wallace_cska32_u_cska62_b[39] = s_wallace_cska32_fa878_xor1[0];
  assign s_wallace_cska32_u_cska62_b[40] = s_wallace_cska32_fa879_xor1[0];
  assign s_wallace_cska32_u_cska62_b[41] = s_wallace_cska32_fa880_xor1[0];
  assign s_wallace_cska32_u_cska62_b[42] = s_wallace_cska32_fa881_xor1[0];
  assign s_wallace_cska32_u_cska62_b[43] = s_wallace_cska32_fa882_xor1[0];
  assign s_wallace_cska32_u_cska62_b[44] = s_wallace_cska32_fa883_xor1[0];
  assign s_wallace_cska32_u_cska62_b[45] = s_wallace_cska32_fa884_xor1[0];
  assign s_wallace_cska32_u_cska62_b[46] = s_wallace_cska32_fa885_xor1[0];
  assign s_wallace_cska32_u_cska62_b[47] = s_wallace_cska32_fa886_xor1[0];
  assign s_wallace_cska32_u_cska62_b[48] = s_wallace_cska32_fa887_xor1[0];
  assign s_wallace_cska32_u_cska62_b[49] = s_wallace_cska32_fa888_xor1[0];
  assign s_wallace_cska32_u_cska62_b[50] = s_wallace_cska32_fa889_xor1[0];
  assign s_wallace_cska32_u_cska62_b[51] = s_wallace_cska32_fa890_xor1[0];
  assign s_wallace_cska32_u_cska62_b[52] = s_wallace_cska32_fa891_xor1[0];
  assign s_wallace_cska32_u_cska62_b[53] = s_wallace_cska32_fa892_xor1[0];
  assign s_wallace_cska32_u_cska62_b[54] = s_wallace_cska32_fa893_xor1[0];
  assign s_wallace_cska32_u_cska62_b[55] = s_wallace_cska32_fa894_xor1[0];
  assign s_wallace_cska32_u_cska62_b[56] = s_wallace_cska32_fa895_xor1[0];
  assign s_wallace_cska32_u_cska62_b[57] = s_wallace_cska32_fa896_xor1[0];
  assign s_wallace_cska32_u_cska62_b[58] = s_wallace_cska32_fa897_xor1[0];
  assign s_wallace_cska32_u_cska62_b[59] = s_wallace_cska32_fa898_xor1[0];
  assign s_wallace_cska32_u_cska62_b[60] = s_wallace_cska32_fa899_xor1[0];
  assign s_wallace_cska32_u_cska62_b[61] = s_wallace_cska32_and_31_31[0];
  u_cska62 u_cska62_s_wallace_cska32_u_cska62_out(.a(s_wallace_cska32_u_cska62_a), .b(s_wallace_cska32_u_cska62_b), .u_cska62_out(s_wallace_cska32_u_cska62_out));
  not_gate not_gate_s_wallace_cska32_xor0(.a(s_wallace_cska32_u_cska62_out[62]), .out(s_wallace_cska32_xor0));

  assign s_wallace_cska32_out[0] = s_wallace_cska32_and_0_0[0];
  assign s_wallace_cska32_out[1] = s_wallace_cska32_u_cska62_out[0];
  assign s_wallace_cska32_out[2] = s_wallace_cska32_u_cska62_out[1];
  assign s_wallace_cska32_out[3] = s_wallace_cska32_u_cska62_out[2];
  assign s_wallace_cska32_out[4] = s_wallace_cska32_u_cska62_out[3];
  assign s_wallace_cska32_out[5] = s_wallace_cska32_u_cska62_out[4];
  assign s_wallace_cska32_out[6] = s_wallace_cska32_u_cska62_out[5];
  assign s_wallace_cska32_out[7] = s_wallace_cska32_u_cska62_out[6];
  assign s_wallace_cska32_out[8] = s_wallace_cska32_u_cska62_out[7];
  assign s_wallace_cska32_out[9] = s_wallace_cska32_u_cska62_out[8];
  assign s_wallace_cska32_out[10] = s_wallace_cska32_u_cska62_out[9];
  assign s_wallace_cska32_out[11] = s_wallace_cska32_u_cska62_out[10];
  assign s_wallace_cska32_out[12] = s_wallace_cska32_u_cska62_out[11];
  assign s_wallace_cska32_out[13] = s_wallace_cska32_u_cska62_out[12];
  assign s_wallace_cska32_out[14] = s_wallace_cska32_u_cska62_out[13];
  assign s_wallace_cska32_out[15] = s_wallace_cska32_u_cska62_out[14];
  assign s_wallace_cska32_out[16] = s_wallace_cska32_u_cska62_out[15];
  assign s_wallace_cska32_out[17] = s_wallace_cska32_u_cska62_out[16];
  assign s_wallace_cska32_out[18] = s_wallace_cska32_u_cska62_out[17];
  assign s_wallace_cska32_out[19] = s_wallace_cska32_u_cska62_out[18];
  assign s_wallace_cska32_out[20] = s_wallace_cska32_u_cska62_out[19];
  assign s_wallace_cska32_out[21] = s_wallace_cska32_u_cska62_out[20];
  assign s_wallace_cska32_out[22] = s_wallace_cska32_u_cska62_out[21];
  assign s_wallace_cska32_out[23] = s_wallace_cska32_u_cska62_out[22];
  assign s_wallace_cska32_out[24] = s_wallace_cska32_u_cska62_out[23];
  assign s_wallace_cska32_out[25] = s_wallace_cska32_u_cska62_out[24];
  assign s_wallace_cska32_out[26] = s_wallace_cska32_u_cska62_out[25];
  assign s_wallace_cska32_out[27] = s_wallace_cska32_u_cska62_out[26];
  assign s_wallace_cska32_out[28] = s_wallace_cska32_u_cska62_out[27];
  assign s_wallace_cska32_out[29] = s_wallace_cska32_u_cska62_out[28];
  assign s_wallace_cska32_out[30] = s_wallace_cska32_u_cska62_out[29];
  assign s_wallace_cska32_out[31] = s_wallace_cska32_u_cska62_out[30];
  assign s_wallace_cska32_out[32] = s_wallace_cska32_u_cska62_out[31];
  assign s_wallace_cska32_out[33] = s_wallace_cska32_u_cska62_out[32];
  assign s_wallace_cska32_out[34] = s_wallace_cska32_u_cska62_out[33];
  assign s_wallace_cska32_out[35] = s_wallace_cska32_u_cska62_out[34];
  assign s_wallace_cska32_out[36] = s_wallace_cska32_u_cska62_out[35];
  assign s_wallace_cska32_out[37] = s_wallace_cska32_u_cska62_out[36];
  assign s_wallace_cska32_out[38] = s_wallace_cska32_u_cska62_out[37];
  assign s_wallace_cska32_out[39] = s_wallace_cska32_u_cska62_out[38];
  assign s_wallace_cska32_out[40] = s_wallace_cska32_u_cska62_out[39];
  assign s_wallace_cska32_out[41] = s_wallace_cska32_u_cska62_out[40];
  assign s_wallace_cska32_out[42] = s_wallace_cska32_u_cska62_out[41];
  assign s_wallace_cska32_out[43] = s_wallace_cska32_u_cska62_out[42];
  assign s_wallace_cska32_out[44] = s_wallace_cska32_u_cska62_out[43];
  assign s_wallace_cska32_out[45] = s_wallace_cska32_u_cska62_out[44];
  assign s_wallace_cska32_out[46] = s_wallace_cska32_u_cska62_out[45];
  assign s_wallace_cska32_out[47] = s_wallace_cska32_u_cska62_out[46];
  assign s_wallace_cska32_out[48] = s_wallace_cska32_u_cska62_out[47];
  assign s_wallace_cska32_out[49] = s_wallace_cska32_u_cska62_out[48];
  assign s_wallace_cska32_out[50] = s_wallace_cska32_u_cska62_out[49];
  assign s_wallace_cska32_out[51] = s_wallace_cska32_u_cska62_out[50];
  assign s_wallace_cska32_out[52] = s_wallace_cska32_u_cska62_out[51];
  assign s_wallace_cska32_out[53] = s_wallace_cska32_u_cska62_out[52];
  assign s_wallace_cska32_out[54] = s_wallace_cska32_u_cska62_out[53];
  assign s_wallace_cska32_out[55] = s_wallace_cska32_u_cska62_out[54];
  assign s_wallace_cska32_out[56] = s_wallace_cska32_u_cska62_out[55];
  assign s_wallace_cska32_out[57] = s_wallace_cska32_u_cska62_out[56];
  assign s_wallace_cska32_out[58] = s_wallace_cska32_u_cska62_out[57];
  assign s_wallace_cska32_out[59] = s_wallace_cska32_u_cska62_out[58];
  assign s_wallace_cska32_out[60] = s_wallace_cska32_u_cska62_out[59];
  assign s_wallace_cska32_out[61] = s_wallace_cska32_u_cska62_out[60];
  assign s_wallace_cska32_out[62] = s_wallace_cska32_u_cska62_out[61];
  assign s_wallace_cska32_out[63] = s_wallace_cska32_xor0[0];
endmodule