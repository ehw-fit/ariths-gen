module f_u_arr_mul3(input [2:0] a, input [2:0] b, output [5:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire b_0;
  wire b_1;
  wire b_2;
  wire f_u_arr_mul3_and_0_0_a_0;
  wire f_u_arr_mul3_and_0_0_b_0;
  wire f_u_arr_mul3_and_0_0_y0;
  wire f_u_arr_mul3_and_1_0_a_1;
  wire f_u_arr_mul3_and_1_0_b_0;
  wire f_u_arr_mul3_and_1_0_y0;
  wire f_u_arr_mul3_and_2_0_a_2;
  wire f_u_arr_mul3_and_2_0_b_0;
  wire f_u_arr_mul3_and_2_0_y0;
  wire f_u_arr_mul3_and_0_1_a_0;
  wire f_u_arr_mul3_and_0_1_b_1;
  wire f_u_arr_mul3_and_0_1_y0;
  wire f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_0_1_y0;
  wire f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_1_0_y0;
  wire f_u_arr_mul3_ha_0_1_y0;
  wire f_u_arr_mul3_ha_0_1_y1;
  wire f_u_arr_mul3_and_1_1_a_1;
  wire f_u_arr_mul3_and_1_1_b_1;
  wire f_u_arr_mul3_and_1_1_y0;
  wire f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_1_1_y0;
  wire f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_2_0_y0;
  wire f_u_arr_mul3_fa_1_1_y0;
  wire f_u_arr_mul3_fa_1_1_y1;
  wire f_u_arr_mul3_fa_1_1_f_u_arr_mul3_ha_0_1_y1;
  wire f_u_arr_mul3_fa_1_1_y2;
  wire f_u_arr_mul3_fa_1_1_y3;
  wire f_u_arr_mul3_fa_1_1_y4;
  wire f_u_arr_mul3_and_2_1_a_2;
  wire f_u_arr_mul3_and_2_1_b_1;
  wire f_u_arr_mul3_and_2_1_y0;
  wire f_u_arr_mul3_ha_2_1_f_u_arr_mul3_and_2_1_y0;
  wire f_u_arr_mul3_ha_2_1_f_u_arr_mul3_fa_1_1_y4;
  wire f_u_arr_mul3_ha_2_1_y0;
  wire f_u_arr_mul3_ha_2_1_y1;
  wire f_u_arr_mul3_and_0_2_a_0;
  wire f_u_arr_mul3_and_0_2_b_2;
  wire f_u_arr_mul3_and_0_2_y0;
  wire f_u_arr_mul3_ha_0_2_f_u_arr_mul3_and_0_2_y0;
  wire f_u_arr_mul3_ha_0_2_f_u_arr_mul3_fa_1_1_y2;
  wire f_u_arr_mul3_ha_0_2_y0;
  wire f_u_arr_mul3_ha_0_2_y1;
  wire f_u_arr_mul3_and_1_2_a_1;
  wire f_u_arr_mul3_and_1_2_b_2;
  wire f_u_arr_mul3_and_1_2_y0;
  wire f_u_arr_mul3_fa_1_2_f_u_arr_mul3_and_1_2_y0;
  wire f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_2_1_y0;
  wire f_u_arr_mul3_fa_1_2_y0;
  wire f_u_arr_mul3_fa_1_2_y1;
  wire f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_0_2_y1;
  wire f_u_arr_mul3_fa_1_2_y2;
  wire f_u_arr_mul3_fa_1_2_y3;
  wire f_u_arr_mul3_fa_1_2_y4;
  wire f_u_arr_mul3_and_2_2_a_2;
  wire f_u_arr_mul3_and_2_2_b_2;
  wire f_u_arr_mul3_and_2_2_y0;
  wire f_u_arr_mul3_fa_2_2_f_u_arr_mul3_and_2_2_y0;
  wire f_u_arr_mul3_fa_2_2_f_u_arr_mul3_ha_2_1_y1;
  wire f_u_arr_mul3_fa_2_2_y0;
  wire f_u_arr_mul3_fa_2_2_y1;
  wire f_u_arr_mul3_fa_2_2_f_u_arr_mul3_fa_1_2_y4;
  wire f_u_arr_mul3_fa_2_2_y2;
  wire f_u_arr_mul3_fa_2_2_y3;
  wire f_u_arr_mul3_fa_2_2_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign f_u_arr_mul3_and_0_0_a_0 = a_0;
  assign f_u_arr_mul3_and_0_0_b_0 = b_0;
  assign f_u_arr_mul3_and_0_0_y0 = f_u_arr_mul3_and_0_0_a_0 & f_u_arr_mul3_and_0_0_b_0;
  assign f_u_arr_mul3_and_1_0_a_1 = a_1;
  assign f_u_arr_mul3_and_1_0_b_0 = b_0;
  assign f_u_arr_mul3_and_1_0_y0 = f_u_arr_mul3_and_1_0_a_1 & f_u_arr_mul3_and_1_0_b_0;
  assign f_u_arr_mul3_and_2_0_a_2 = a_2;
  assign f_u_arr_mul3_and_2_0_b_0 = b_0;
  assign f_u_arr_mul3_and_2_0_y0 = f_u_arr_mul3_and_2_0_a_2 & f_u_arr_mul3_and_2_0_b_0;
  assign f_u_arr_mul3_and_0_1_a_0 = a_0;
  assign f_u_arr_mul3_and_0_1_b_1 = b_1;
  assign f_u_arr_mul3_and_0_1_y0 = f_u_arr_mul3_and_0_1_a_0 & f_u_arr_mul3_and_0_1_b_1;
  assign f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_0_1_y0 = f_u_arr_mul3_and_0_1_y0;
  assign f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_1_0_y0 = f_u_arr_mul3_and_1_0_y0;
  assign f_u_arr_mul3_ha_0_1_y0 = f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_0_1_y0 ^ f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_1_0_y0;
  assign f_u_arr_mul3_ha_0_1_y1 = f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_0_1_y0 & f_u_arr_mul3_ha_0_1_f_u_arr_mul3_and_1_0_y0;
  assign f_u_arr_mul3_and_1_1_a_1 = a_1;
  assign f_u_arr_mul3_and_1_1_b_1 = b_1;
  assign f_u_arr_mul3_and_1_1_y0 = f_u_arr_mul3_and_1_1_a_1 & f_u_arr_mul3_and_1_1_b_1;
  assign f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_1_1_y0 = f_u_arr_mul3_and_1_1_y0;
  assign f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_2_0_y0 = f_u_arr_mul3_and_2_0_y0;
  assign f_u_arr_mul3_fa_1_1_f_u_arr_mul3_ha_0_1_y1 = f_u_arr_mul3_ha_0_1_y1;
  assign f_u_arr_mul3_fa_1_1_y0 = f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_1_1_y0 ^ f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_2_0_y0;
  assign f_u_arr_mul3_fa_1_1_y1 = f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_1_1_y0 & f_u_arr_mul3_fa_1_1_f_u_arr_mul3_and_2_0_y0;
  assign f_u_arr_mul3_fa_1_1_y2 = f_u_arr_mul3_fa_1_1_y0 ^ f_u_arr_mul3_fa_1_1_f_u_arr_mul3_ha_0_1_y1;
  assign f_u_arr_mul3_fa_1_1_y3 = f_u_arr_mul3_fa_1_1_y0 & f_u_arr_mul3_fa_1_1_f_u_arr_mul3_ha_0_1_y1;
  assign f_u_arr_mul3_fa_1_1_y4 = f_u_arr_mul3_fa_1_1_y1 | f_u_arr_mul3_fa_1_1_y3;
  assign f_u_arr_mul3_and_2_1_a_2 = a_2;
  assign f_u_arr_mul3_and_2_1_b_1 = b_1;
  assign f_u_arr_mul3_and_2_1_y0 = f_u_arr_mul3_and_2_1_a_2 & f_u_arr_mul3_and_2_1_b_1;
  assign f_u_arr_mul3_ha_2_1_f_u_arr_mul3_and_2_1_y0 = f_u_arr_mul3_and_2_1_y0;
  assign f_u_arr_mul3_ha_2_1_f_u_arr_mul3_fa_1_1_y4 = f_u_arr_mul3_fa_1_1_y4;
  assign f_u_arr_mul3_ha_2_1_y0 = f_u_arr_mul3_ha_2_1_f_u_arr_mul3_and_2_1_y0 ^ f_u_arr_mul3_ha_2_1_f_u_arr_mul3_fa_1_1_y4;
  assign f_u_arr_mul3_ha_2_1_y1 = f_u_arr_mul3_ha_2_1_f_u_arr_mul3_and_2_1_y0 & f_u_arr_mul3_ha_2_1_f_u_arr_mul3_fa_1_1_y4;
  assign f_u_arr_mul3_and_0_2_a_0 = a_0;
  assign f_u_arr_mul3_and_0_2_b_2 = b_2;
  assign f_u_arr_mul3_and_0_2_y0 = f_u_arr_mul3_and_0_2_a_0 & f_u_arr_mul3_and_0_2_b_2;
  assign f_u_arr_mul3_ha_0_2_f_u_arr_mul3_and_0_2_y0 = f_u_arr_mul3_and_0_2_y0;
  assign f_u_arr_mul3_ha_0_2_f_u_arr_mul3_fa_1_1_y2 = f_u_arr_mul3_fa_1_1_y2;
  assign f_u_arr_mul3_ha_0_2_y0 = f_u_arr_mul3_ha_0_2_f_u_arr_mul3_and_0_2_y0 ^ f_u_arr_mul3_ha_0_2_f_u_arr_mul3_fa_1_1_y2;
  assign f_u_arr_mul3_ha_0_2_y1 = f_u_arr_mul3_ha_0_2_f_u_arr_mul3_and_0_2_y0 & f_u_arr_mul3_ha_0_2_f_u_arr_mul3_fa_1_1_y2;
  assign f_u_arr_mul3_and_1_2_a_1 = a_1;
  assign f_u_arr_mul3_and_1_2_b_2 = b_2;
  assign f_u_arr_mul3_and_1_2_y0 = f_u_arr_mul3_and_1_2_a_1 & f_u_arr_mul3_and_1_2_b_2;
  assign f_u_arr_mul3_fa_1_2_f_u_arr_mul3_and_1_2_y0 = f_u_arr_mul3_and_1_2_y0;
  assign f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_2_1_y0 = f_u_arr_mul3_ha_2_1_y0;
  assign f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_0_2_y1 = f_u_arr_mul3_ha_0_2_y1;
  assign f_u_arr_mul3_fa_1_2_y0 = f_u_arr_mul3_fa_1_2_f_u_arr_mul3_and_1_2_y0 ^ f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_2_1_y0;
  assign f_u_arr_mul3_fa_1_2_y1 = f_u_arr_mul3_fa_1_2_f_u_arr_mul3_and_1_2_y0 & f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_2_1_y0;
  assign f_u_arr_mul3_fa_1_2_y2 = f_u_arr_mul3_fa_1_2_y0 ^ f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_0_2_y1;
  assign f_u_arr_mul3_fa_1_2_y3 = f_u_arr_mul3_fa_1_2_y0 & f_u_arr_mul3_fa_1_2_f_u_arr_mul3_ha_0_2_y1;
  assign f_u_arr_mul3_fa_1_2_y4 = f_u_arr_mul3_fa_1_2_y1 | f_u_arr_mul3_fa_1_2_y3;
  assign f_u_arr_mul3_and_2_2_a_2 = a_2;
  assign f_u_arr_mul3_and_2_2_b_2 = b_2;
  assign f_u_arr_mul3_and_2_2_y0 = f_u_arr_mul3_and_2_2_a_2 & f_u_arr_mul3_and_2_2_b_2;
  assign f_u_arr_mul3_fa_2_2_f_u_arr_mul3_and_2_2_y0 = f_u_arr_mul3_and_2_2_y0;
  assign f_u_arr_mul3_fa_2_2_f_u_arr_mul3_ha_2_1_y1 = f_u_arr_mul3_ha_2_1_y1;
  assign f_u_arr_mul3_fa_2_2_f_u_arr_mul3_fa_1_2_y4 = f_u_arr_mul3_fa_1_2_y4;
  assign f_u_arr_mul3_fa_2_2_y0 = f_u_arr_mul3_fa_2_2_f_u_arr_mul3_and_2_2_y0 ^ f_u_arr_mul3_fa_2_2_f_u_arr_mul3_ha_2_1_y1;
  assign f_u_arr_mul3_fa_2_2_y1 = f_u_arr_mul3_fa_2_2_f_u_arr_mul3_and_2_2_y0 & f_u_arr_mul3_fa_2_2_f_u_arr_mul3_ha_2_1_y1;
  assign f_u_arr_mul3_fa_2_2_y2 = f_u_arr_mul3_fa_2_2_y0 ^ f_u_arr_mul3_fa_2_2_f_u_arr_mul3_fa_1_2_y4;
  assign f_u_arr_mul3_fa_2_2_y3 = f_u_arr_mul3_fa_2_2_y0 & f_u_arr_mul3_fa_2_2_f_u_arr_mul3_fa_1_2_y4;
  assign f_u_arr_mul3_fa_2_2_y4 = f_u_arr_mul3_fa_2_2_y1 | f_u_arr_mul3_fa_2_2_y3;

  assign out[0] = f_u_arr_mul3_and_0_0_y0;
  assign out[1] = f_u_arr_mul3_ha_0_1_y0;
  assign out[2] = f_u_arr_mul3_ha_0_2_y0;
  assign out[3] = f_u_arr_mul3_fa_1_2_y2;
  assign out[4] = f_u_arr_mul3_fa_2_2_y2;
  assign out[5] = f_u_arr_mul3_fa_2_2_y4;
endmodule