module s_cla8(input [7:0] a, input [7:0] b, output [8:0] s_cla8_out);
  wire s_cla8_pg_logic0_or0;
  wire s_cla8_pg_logic0_and0;
  wire s_cla8_pg_logic0_xor0;
  wire s_cla8_pg_logic1_or0;
  wire s_cla8_pg_logic1_and0;
  wire s_cla8_pg_logic1_xor0;
  wire s_cla8_xor1;
  wire s_cla8_and0;
  wire s_cla8_or0;
  wire s_cla8_pg_logic2_or0;
  wire s_cla8_pg_logic2_and0;
  wire s_cla8_pg_logic2_xor0;
  wire s_cla8_xor2;
  wire s_cla8_and1;
  wire s_cla8_and2;
  wire s_cla8_and3;
  wire s_cla8_and4;
  wire s_cla8_or1;
  wire s_cla8_or2;
  wire s_cla8_pg_logic3_or0;
  wire s_cla8_pg_logic3_and0;
  wire s_cla8_pg_logic3_xor0;
  wire s_cla8_xor3;
  wire s_cla8_and5;
  wire s_cla8_and6;
  wire s_cla8_and7;
  wire s_cla8_and8;
  wire s_cla8_and9;
  wire s_cla8_and10;
  wire s_cla8_and11;
  wire s_cla8_or3;
  wire s_cla8_or4;
  wire s_cla8_or5;
  wire s_cla8_pg_logic4_or0;
  wire s_cla8_pg_logic4_and0;
  wire s_cla8_pg_logic4_xor0;
  wire s_cla8_xor4;
  wire s_cla8_and12;
  wire s_cla8_or6;
  wire s_cla8_pg_logic5_or0;
  wire s_cla8_pg_logic5_and0;
  wire s_cla8_pg_logic5_xor0;
  wire s_cla8_xor5;
  wire s_cla8_and13;
  wire s_cla8_and14;
  wire s_cla8_and15;
  wire s_cla8_or7;
  wire s_cla8_or8;
  wire s_cla8_pg_logic6_or0;
  wire s_cla8_pg_logic6_and0;
  wire s_cla8_pg_logic6_xor0;
  wire s_cla8_xor6;
  wire s_cla8_and16;
  wire s_cla8_and17;
  wire s_cla8_and18;
  wire s_cla8_and19;
  wire s_cla8_and20;
  wire s_cla8_and21;
  wire s_cla8_or9;
  wire s_cla8_or10;
  wire s_cla8_or11;
  wire s_cla8_pg_logic7_or0;
  wire s_cla8_pg_logic7_and0;
  wire s_cla8_pg_logic7_xor0;
  wire s_cla8_xor7;
  wire s_cla8_and22;
  wire s_cla8_and23;
  wire s_cla8_and24;
  wire s_cla8_and25;
  wire s_cla8_and26;
  wire s_cla8_and27;
  wire s_cla8_and28;
  wire s_cla8_and29;
  wire s_cla8_and30;
  wire s_cla8_and31;
  wire s_cla8_or12;
  wire s_cla8_or13;
  wire s_cla8_or14;
  wire s_cla8_or15;
  wire s_cla8_xor8;
  wire s_cla8_xor9;

  assign s_cla8_pg_logic0_or0 = a[0] | b[0];
  assign s_cla8_pg_logic0_and0 = a[0] & b[0];
  assign s_cla8_pg_logic0_xor0 = a[0] ^ b[0];
  assign s_cla8_pg_logic1_or0 = a[1] | b[1];
  assign s_cla8_pg_logic1_and0 = a[1] & b[1];
  assign s_cla8_pg_logic1_xor0 = a[1] ^ b[1];
  assign s_cla8_xor1 = s_cla8_pg_logic1_xor0 ^ s_cla8_pg_logic0_and0;
  assign s_cla8_and0 = s_cla8_pg_logic0_and0 & s_cla8_pg_logic1_or0;
  assign s_cla8_or0 = s_cla8_pg_logic1_and0 | s_cla8_and0;
  assign s_cla8_pg_logic2_or0 = a[2] | b[2];
  assign s_cla8_pg_logic2_and0 = a[2] & b[2];
  assign s_cla8_pg_logic2_xor0 = a[2] ^ b[2];
  assign s_cla8_xor2 = s_cla8_pg_logic2_xor0 ^ s_cla8_or0;
  assign s_cla8_and1 = s_cla8_pg_logic2_or0 & s_cla8_pg_logic0_or0;
  assign s_cla8_and2 = s_cla8_pg_logic0_and0 & s_cla8_pg_logic2_or0;
  assign s_cla8_and3 = s_cla8_and2 & s_cla8_pg_logic1_or0;
  assign s_cla8_and4 = s_cla8_pg_logic1_and0 & s_cla8_pg_logic2_or0;
  assign s_cla8_or1 = s_cla8_and3 | s_cla8_and4;
  assign s_cla8_or2 = s_cla8_pg_logic2_and0 | s_cla8_or1;
  assign s_cla8_pg_logic3_or0 = a[3] | b[3];
  assign s_cla8_pg_logic3_and0 = a[3] & b[3];
  assign s_cla8_pg_logic3_xor0 = a[3] ^ b[3];
  assign s_cla8_xor3 = s_cla8_pg_logic3_xor0 ^ s_cla8_or2;
  assign s_cla8_and5 = s_cla8_pg_logic3_or0 & s_cla8_pg_logic1_or0;
  assign s_cla8_and6 = s_cla8_pg_logic0_and0 & s_cla8_pg_logic2_or0;
  assign s_cla8_and7 = s_cla8_pg_logic3_or0 & s_cla8_pg_logic1_or0;
  assign s_cla8_and8 = s_cla8_and6 & s_cla8_and7;
  assign s_cla8_and9 = s_cla8_pg_logic1_and0 & s_cla8_pg_logic3_or0;
  assign s_cla8_and10 = s_cla8_and9 & s_cla8_pg_logic2_or0;
  assign s_cla8_and11 = s_cla8_pg_logic2_and0 & s_cla8_pg_logic3_or0;
  assign s_cla8_or3 = s_cla8_and8 | s_cla8_and11;
  assign s_cla8_or4 = s_cla8_and10 | s_cla8_or3;
  assign s_cla8_or5 = s_cla8_pg_logic3_and0 | s_cla8_or4;
  assign s_cla8_pg_logic4_or0 = a[4] | b[4];
  assign s_cla8_pg_logic4_and0 = a[4] & b[4];
  assign s_cla8_pg_logic4_xor0 = a[4] ^ b[4];
  assign s_cla8_xor4 = s_cla8_pg_logic4_xor0 ^ s_cla8_or5;
  assign s_cla8_and12 = s_cla8_or5 & s_cla8_pg_logic4_or0;
  assign s_cla8_or6 = s_cla8_pg_logic4_and0 | s_cla8_and12;
  assign s_cla8_pg_logic5_or0 = a[5] | b[5];
  assign s_cla8_pg_logic5_and0 = a[5] & b[5];
  assign s_cla8_pg_logic5_xor0 = a[5] ^ b[5];
  assign s_cla8_xor5 = s_cla8_pg_logic5_xor0 ^ s_cla8_or6;
  assign s_cla8_and13 = s_cla8_or5 & s_cla8_pg_logic5_or0;
  assign s_cla8_and14 = s_cla8_and13 & s_cla8_pg_logic4_or0;
  assign s_cla8_and15 = s_cla8_pg_logic4_and0 & s_cla8_pg_logic5_or0;
  assign s_cla8_or7 = s_cla8_and14 | s_cla8_and15;
  assign s_cla8_or8 = s_cla8_pg_logic5_and0 | s_cla8_or7;
  assign s_cla8_pg_logic6_or0 = a[6] | b[6];
  assign s_cla8_pg_logic6_and0 = a[6] & b[6];
  assign s_cla8_pg_logic6_xor0 = a[6] ^ b[6];
  assign s_cla8_xor6 = s_cla8_pg_logic6_xor0 ^ s_cla8_or8;
  assign s_cla8_and16 = s_cla8_or5 & s_cla8_pg_logic5_or0;
  assign s_cla8_and17 = s_cla8_pg_logic6_or0 & s_cla8_pg_logic4_or0;
  assign s_cla8_and18 = s_cla8_and16 & s_cla8_and17;
  assign s_cla8_and19 = s_cla8_pg_logic4_and0 & s_cla8_pg_logic6_or0;
  assign s_cla8_and20 = s_cla8_and19 & s_cla8_pg_logic5_or0;
  assign s_cla8_and21 = s_cla8_pg_logic5_and0 & s_cla8_pg_logic6_or0;
  assign s_cla8_or9 = s_cla8_and18 | s_cla8_and20;
  assign s_cla8_or10 = s_cla8_or9 | s_cla8_and21;
  assign s_cla8_or11 = s_cla8_pg_logic6_and0 | s_cla8_or10;
  assign s_cla8_pg_logic7_or0 = a[7] | b[7];
  assign s_cla8_pg_logic7_and0 = a[7] & b[7];
  assign s_cla8_pg_logic7_xor0 = a[7] ^ b[7];
  assign s_cla8_xor7 = s_cla8_pg_logic7_xor0 ^ s_cla8_or11;
  assign s_cla8_and22 = s_cla8_or5 & s_cla8_pg_logic6_or0;
  assign s_cla8_and23 = s_cla8_pg_logic7_or0 & s_cla8_pg_logic5_or0;
  assign s_cla8_and24 = s_cla8_and22 & s_cla8_and23;
  assign s_cla8_and25 = s_cla8_and24 & s_cla8_pg_logic4_or0;
  assign s_cla8_and26 = s_cla8_pg_logic4_and0 & s_cla8_pg_logic6_or0;
  assign s_cla8_and27 = s_cla8_pg_logic7_or0 & s_cla8_pg_logic5_or0;
  assign s_cla8_and28 = s_cla8_and26 & s_cla8_and27;
  assign s_cla8_and29 = s_cla8_pg_logic5_and0 & s_cla8_pg_logic7_or0;
  assign s_cla8_and30 = s_cla8_and29 & s_cla8_pg_logic6_or0;
  assign s_cla8_and31 = s_cla8_pg_logic6_and0 & s_cla8_pg_logic7_or0;
  assign s_cla8_or12 = s_cla8_and25 | s_cla8_and30;
  assign s_cla8_or13 = s_cla8_and28 | s_cla8_and31;
  assign s_cla8_or14 = s_cla8_or12 | s_cla8_or13;
  assign s_cla8_or15 = s_cla8_pg_logic7_and0 | s_cla8_or14;
  assign s_cla8_xor8 = a[7] ^ b[7];
  assign s_cla8_xor9 = s_cla8_xor8 ^ s_cla8_or15;

  assign s_cla8_out[0] = s_cla8_pg_logic0_xor0;
  assign s_cla8_out[1] = s_cla8_xor1;
  assign s_cla8_out[2] = s_cla8_xor2;
  assign s_cla8_out[3] = s_cla8_xor3;
  assign s_cla8_out[4] = s_cla8_xor4;
  assign s_cla8_out[5] = s_cla8_xor5;
  assign s_cla8_out[6] = s_cla8_xor6;
  assign s_cla8_out[7] = s_cla8_xor7;
  assign s_cla8_out[8] = s_cla8_xor9;
endmodule