module _and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule