module and_gate(input a, input b, output and_gate);
  assign and_gate = a & b;
endmodule