module f_arrdiv8(input [7:0] a, input [7:0] b, output [7:0] f_arrdiv8_out);
  wire f_arrdiv8_fs0_xor0;
  wire f_arrdiv8_fs0_not0;
  wire f_arrdiv8_fs0_and0;
  wire f_arrdiv8_fs0_not1;
  wire f_arrdiv8_fs1_xor1;
  wire f_arrdiv8_fs1_not1;
  wire f_arrdiv8_fs1_and1;
  wire f_arrdiv8_fs1_or0;
  wire f_arrdiv8_fs2_xor1;
  wire f_arrdiv8_fs2_not1;
  wire f_arrdiv8_fs2_and1;
  wire f_arrdiv8_fs2_or0;
  wire f_arrdiv8_fs3_xor1;
  wire f_arrdiv8_fs3_not1;
  wire f_arrdiv8_fs3_and1;
  wire f_arrdiv8_fs3_or0;
  wire f_arrdiv8_fs4_xor1;
  wire f_arrdiv8_fs4_not1;
  wire f_arrdiv8_fs4_and1;
  wire f_arrdiv8_fs4_or0;
  wire f_arrdiv8_fs5_xor1;
  wire f_arrdiv8_fs5_not1;
  wire f_arrdiv8_fs5_and1;
  wire f_arrdiv8_fs5_or0;
  wire f_arrdiv8_fs6_xor1;
  wire f_arrdiv8_fs6_not1;
  wire f_arrdiv8_fs6_and1;
  wire f_arrdiv8_fs6_or0;
  wire f_arrdiv8_fs7_xor1;
  wire f_arrdiv8_fs7_not1;
  wire f_arrdiv8_fs7_and1;
  wire f_arrdiv8_fs7_or0;
  wire f_arrdiv8_mux2to10_and0;
  wire f_arrdiv8_mux2to10_not0;
  wire f_arrdiv8_mux2to10_and1;
  wire f_arrdiv8_mux2to10_xor0;
  wire f_arrdiv8_mux2to11_not0;
  wire f_arrdiv8_mux2to11_and1;
  wire f_arrdiv8_mux2to12_not0;
  wire f_arrdiv8_mux2to12_and1;
  wire f_arrdiv8_mux2to13_not0;
  wire f_arrdiv8_mux2to13_and1;
  wire f_arrdiv8_mux2to14_not0;
  wire f_arrdiv8_mux2to14_and1;
  wire f_arrdiv8_mux2to15_not0;
  wire f_arrdiv8_mux2to15_and1;
  wire f_arrdiv8_mux2to16_not0;
  wire f_arrdiv8_mux2to16_and1;
  wire f_arrdiv8_not0;
  wire f_arrdiv8_fs8_xor0;
  wire f_arrdiv8_fs8_not0;
  wire f_arrdiv8_fs8_and0;
  wire f_arrdiv8_fs8_not1;
  wire f_arrdiv8_fs9_xor0;
  wire f_arrdiv8_fs9_not0;
  wire f_arrdiv8_fs9_and0;
  wire f_arrdiv8_fs9_xor1;
  wire f_arrdiv8_fs9_not1;
  wire f_arrdiv8_fs9_and1;
  wire f_arrdiv8_fs9_or0;
  wire f_arrdiv8_fs10_xor0;
  wire f_arrdiv8_fs10_not0;
  wire f_arrdiv8_fs10_and0;
  wire f_arrdiv8_fs10_xor1;
  wire f_arrdiv8_fs10_not1;
  wire f_arrdiv8_fs10_and1;
  wire f_arrdiv8_fs10_or0;
  wire f_arrdiv8_fs11_xor0;
  wire f_arrdiv8_fs11_not0;
  wire f_arrdiv8_fs11_and0;
  wire f_arrdiv8_fs11_xor1;
  wire f_arrdiv8_fs11_not1;
  wire f_arrdiv8_fs11_and1;
  wire f_arrdiv8_fs11_or0;
  wire f_arrdiv8_fs12_xor0;
  wire f_arrdiv8_fs12_not0;
  wire f_arrdiv8_fs12_and0;
  wire f_arrdiv8_fs12_xor1;
  wire f_arrdiv8_fs12_not1;
  wire f_arrdiv8_fs12_and1;
  wire f_arrdiv8_fs12_or0;
  wire f_arrdiv8_fs13_xor0;
  wire f_arrdiv8_fs13_not0;
  wire f_arrdiv8_fs13_and0;
  wire f_arrdiv8_fs13_xor1;
  wire f_arrdiv8_fs13_not1;
  wire f_arrdiv8_fs13_and1;
  wire f_arrdiv8_fs13_or0;
  wire f_arrdiv8_fs14_xor0;
  wire f_arrdiv8_fs14_not0;
  wire f_arrdiv8_fs14_and0;
  wire f_arrdiv8_fs14_xor1;
  wire f_arrdiv8_fs14_not1;
  wire f_arrdiv8_fs14_and1;
  wire f_arrdiv8_fs14_or0;
  wire f_arrdiv8_fs15_xor0;
  wire f_arrdiv8_fs15_not0;
  wire f_arrdiv8_fs15_and0;
  wire f_arrdiv8_fs15_xor1;
  wire f_arrdiv8_fs15_not1;
  wire f_arrdiv8_fs15_and1;
  wire f_arrdiv8_fs15_or0;
  wire f_arrdiv8_mux2to17_and0;
  wire f_arrdiv8_mux2to17_not0;
  wire f_arrdiv8_mux2to17_and1;
  wire f_arrdiv8_mux2to17_xor0;
  wire f_arrdiv8_mux2to18_and0;
  wire f_arrdiv8_mux2to18_not0;
  wire f_arrdiv8_mux2to18_and1;
  wire f_arrdiv8_mux2to18_xor0;
  wire f_arrdiv8_mux2to19_and0;
  wire f_arrdiv8_mux2to19_not0;
  wire f_arrdiv8_mux2to19_and1;
  wire f_arrdiv8_mux2to19_xor0;
  wire f_arrdiv8_mux2to110_and0;
  wire f_arrdiv8_mux2to110_not0;
  wire f_arrdiv8_mux2to110_and1;
  wire f_arrdiv8_mux2to110_xor0;
  wire f_arrdiv8_mux2to111_and0;
  wire f_arrdiv8_mux2to111_not0;
  wire f_arrdiv8_mux2to111_and1;
  wire f_arrdiv8_mux2to111_xor0;
  wire f_arrdiv8_mux2to112_and0;
  wire f_arrdiv8_mux2to112_not0;
  wire f_arrdiv8_mux2to112_and1;
  wire f_arrdiv8_mux2to112_xor0;
  wire f_arrdiv8_mux2to113_and0;
  wire f_arrdiv8_mux2to113_not0;
  wire f_arrdiv8_mux2to113_and1;
  wire f_arrdiv8_mux2to113_xor0;
  wire f_arrdiv8_not1;
  wire f_arrdiv8_fs16_xor0;
  wire f_arrdiv8_fs16_not0;
  wire f_arrdiv8_fs16_and0;
  wire f_arrdiv8_fs16_not1;
  wire f_arrdiv8_fs17_xor0;
  wire f_arrdiv8_fs17_not0;
  wire f_arrdiv8_fs17_and0;
  wire f_arrdiv8_fs17_xor1;
  wire f_arrdiv8_fs17_not1;
  wire f_arrdiv8_fs17_and1;
  wire f_arrdiv8_fs17_or0;
  wire f_arrdiv8_fs18_xor0;
  wire f_arrdiv8_fs18_not0;
  wire f_arrdiv8_fs18_and0;
  wire f_arrdiv8_fs18_xor1;
  wire f_arrdiv8_fs18_not1;
  wire f_arrdiv8_fs18_and1;
  wire f_arrdiv8_fs18_or0;
  wire f_arrdiv8_fs19_xor0;
  wire f_arrdiv8_fs19_not0;
  wire f_arrdiv8_fs19_and0;
  wire f_arrdiv8_fs19_xor1;
  wire f_arrdiv8_fs19_not1;
  wire f_arrdiv8_fs19_and1;
  wire f_arrdiv8_fs19_or0;
  wire f_arrdiv8_fs20_xor0;
  wire f_arrdiv8_fs20_not0;
  wire f_arrdiv8_fs20_and0;
  wire f_arrdiv8_fs20_xor1;
  wire f_arrdiv8_fs20_not1;
  wire f_arrdiv8_fs20_and1;
  wire f_arrdiv8_fs20_or0;
  wire f_arrdiv8_fs21_xor0;
  wire f_arrdiv8_fs21_not0;
  wire f_arrdiv8_fs21_and0;
  wire f_arrdiv8_fs21_xor1;
  wire f_arrdiv8_fs21_not1;
  wire f_arrdiv8_fs21_and1;
  wire f_arrdiv8_fs21_or0;
  wire f_arrdiv8_fs22_xor0;
  wire f_arrdiv8_fs22_not0;
  wire f_arrdiv8_fs22_and0;
  wire f_arrdiv8_fs22_xor1;
  wire f_arrdiv8_fs22_not1;
  wire f_arrdiv8_fs22_and1;
  wire f_arrdiv8_fs22_or0;
  wire f_arrdiv8_fs23_xor0;
  wire f_arrdiv8_fs23_not0;
  wire f_arrdiv8_fs23_and0;
  wire f_arrdiv8_fs23_xor1;
  wire f_arrdiv8_fs23_not1;
  wire f_arrdiv8_fs23_and1;
  wire f_arrdiv8_fs23_or0;
  wire f_arrdiv8_mux2to114_and0;
  wire f_arrdiv8_mux2to114_not0;
  wire f_arrdiv8_mux2to114_and1;
  wire f_arrdiv8_mux2to114_xor0;
  wire f_arrdiv8_mux2to115_and0;
  wire f_arrdiv8_mux2to115_not0;
  wire f_arrdiv8_mux2to115_and1;
  wire f_arrdiv8_mux2to115_xor0;
  wire f_arrdiv8_mux2to116_and0;
  wire f_arrdiv8_mux2to116_not0;
  wire f_arrdiv8_mux2to116_and1;
  wire f_arrdiv8_mux2to116_xor0;
  wire f_arrdiv8_mux2to117_and0;
  wire f_arrdiv8_mux2to117_not0;
  wire f_arrdiv8_mux2to117_and1;
  wire f_arrdiv8_mux2to117_xor0;
  wire f_arrdiv8_mux2to118_and0;
  wire f_arrdiv8_mux2to118_not0;
  wire f_arrdiv8_mux2to118_and1;
  wire f_arrdiv8_mux2to118_xor0;
  wire f_arrdiv8_mux2to119_and0;
  wire f_arrdiv8_mux2to119_not0;
  wire f_arrdiv8_mux2to119_and1;
  wire f_arrdiv8_mux2to119_xor0;
  wire f_arrdiv8_mux2to120_and0;
  wire f_arrdiv8_mux2to120_not0;
  wire f_arrdiv8_mux2to120_and1;
  wire f_arrdiv8_mux2to120_xor0;
  wire f_arrdiv8_not2;
  wire f_arrdiv8_fs24_xor0;
  wire f_arrdiv8_fs24_not0;
  wire f_arrdiv8_fs24_and0;
  wire f_arrdiv8_fs24_not1;
  wire f_arrdiv8_fs25_xor0;
  wire f_arrdiv8_fs25_not0;
  wire f_arrdiv8_fs25_and0;
  wire f_arrdiv8_fs25_xor1;
  wire f_arrdiv8_fs25_not1;
  wire f_arrdiv8_fs25_and1;
  wire f_arrdiv8_fs25_or0;
  wire f_arrdiv8_fs26_xor0;
  wire f_arrdiv8_fs26_not0;
  wire f_arrdiv8_fs26_and0;
  wire f_arrdiv8_fs26_xor1;
  wire f_arrdiv8_fs26_not1;
  wire f_arrdiv8_fs26_and1;
  wire f_arrdiv8_fs26_or0;
  wire f_arrdiv8_fs27_xor0;
  wire f_arrdiv8_fs27_not0;
  wire f_arrdiv8_fs27_and0;
  wire f_arrdiv8_fs27_xor1;
  wire f_arrdiv8_fs27_not1;
  wire f_arrdiv8_fs27_and1;
  wire f_arrdiv8_fs27_or0;
  wire f_arrdiv8_fs28_xor0;
  wire f_arrdiv8_fs28_not0;
  wire f_arrdiv8_fs28_and0;
  wire f_arrdiv8_fs28_xor1;
  wire f_arrdiv8_fs28_not1;
  wire f_arrdiv8_fs28_and1;
  wire f_arrdiv8_fs28_or0;
  wire f_arrdiv8_fs29_xor0;
  wire f_arrdiv8_fs29_not0;
  wire f_arrdiv8_fs29_and0;
  wire f_arrdiv8_fs29_xor1;
  wire f_arrdiv8_fs29_not1;
  wire f_arrdiv8_fs29_and1;
  wire f_arrdiv8_fs29_or0;
  wire f_arrdiv8_fs30_xor0;
  wire f_arrdiv8_fs30_not0;
  wire f_arrdiv8_fs30_and0;
  wire f_arrdiv8_fs30_xor1;
  wire f_arrdiv8_fs30_not1;
  wire f_arrdiv8_fs30_and1;
  wire f_arrdiv8_fs30_or0;
  wire f_arrdiv8_fs31_xor0;
  wire f_arrdiv8_fs31_not0;
  wire f_arrdiv8_fs31_and0;
  wire f_arrdiv8_fs31_xor1;
  wire f_arrdiv8_fs31_not1;
  wire f_arrdiv8_fs31_and1;
  wire f_arrdiv8_fs31_or0;
  wire f_arrdiv8_mux2to121_and0;
  wire f_arrdiv8_mux2to121_not0;
  wire f_arrdiv8_mux2to121_and1;
  wire f_arrdiv8_mux2to121_xor0;
  wire f_arrdiv8_mux2to122_and0;
  wire f_arrdiv8_mux2to122_not0;
  wire f_arrdiv8_mux2to122_and1;
  wire f_arrdiv8_mux2to122_xor0;
  wire f_arrdiv8_mux2to123_and0;
  wire f_arrdiv8_mux2to123_not0;
  wire f_arrdiv8_mux2to123_and1;
  wire f_arrdiv8_mux2to123_xor0;
  wire f_arrdiv8_mux2to124_and0;
  wire f_arrdiv8_mux2to124_not0;
  wire f_arrdiv8_mux2to124_and1;
  wire f_arrdiv8_mux2to124_xor0;
  wire f_arrdiv8_mux2to125_and0;
  wire f_arrdiv8_mux2to125_not0;
  wire f_arrdiv8_mux2to125_and1;
  wire f_arrdiv8_mux2to125_xor0;
  wire f_arrdiv8_mux2to126_and0;
  wire f_arrdiv8_mux2to126_not0;
  wire f_arrdiv8_mux2to126_and1;
  wire f_arrdiv8_mux2to126_xor0;
  wire f_arrdiv8_mux2to127_and0;
  wire f_arrdiv8_mux2to127_not0;
  wire f_arrdiv8_mux2to127_and1;
  wire f_arrdiv8_mux2to127_xor0;
  wire f_arrdiv8_not3;
  wire f_arrdiv8_fs32_xor0;
  wire f_arrdiv8_fs32_not0;
  wire f_arrdiv8_fs32_and0;
  wire f_arrdiv8_fs32_not1;
  wire f_arrdiv8_fs33_xor0;
  wire f_arrdiv8_fs33_not0;
  wire f_arrdiv8_fs33_and0;
  wire f_arrdiv8_fs33_xor1;
  wire f_arrdiv8_fs33_not1;
  wire f_arrdiv8_fs33_and1;
  wire f_arrdiv8_fs33_or0;
  wire f_arrdiv8_fs34_xor0;
  wire f_arrdiv8_fs34_not0;
  wire f_arrdiv8_fs34_and0;
  wire f_arrdiv8_fs34_xor1;
  wire f_arrdiv8_fs34_not1;
  wire f_arrdiv8_fs34_and1;
  wire f_arrdiv8_fs34_or0;
  wire f_arrdiv8_fs35_xor0;
  wire f_arrdiv8_fs35_not0;
  wire f_arrdiv8_fs35_and0;
  wire f_arrdiv8_fs35_xor1;
  wire f_arrdiv8_fs35_not1;
  wire f_arrdiv8_fs35_and1;
  wire f_arrdiv8_fs35_or0;
  wire f_arrdiv8_fs36_xor0;
  wire f_arrdiv8_fs36_not0;
  wire f_arrdiv8_fs36_and0;
  wire f_arrdiv8_fs36_xor1;
  wire f_arrdiv8_fs36_not1;
  wire f_arrdiv8_fs36_and1;
  wire f_arrdiv8_fs36_or0;
  wire f_arrdiv8_fs37_xor0;
  wire f_arrdiv8_fs37_not0;
  wire f_arrdiv8_fs37_and0;
  wire f_arrdiv8_fs37_xor1;
  wire f_arrdiv8_fs37_not1;
  wire f_arrdiv8_fs37_and1;
  wire f_arrdiv8_fs37_or0;
  wire f_arrdiv8_fs38_xor0;
  wire f_arrdiv8_fs38_not0;
  wire f_arrdiv8_fs38_and0;
  wire f_arrdiv8_fs38_xor1;
  wire f_arrdiv8_fs38_not1;
  wire f_arrdiv8_fs38_and1;
  wire f_arrdiv8_fs38_or0;
  wire f_arrdiv8_fs39_xor0;
  wire f_arrdiv8_fs39_not0;
  wire f_arrdiv8_fs39_and0;
  wire f_arrdiv8_fs39_xor1;
  wire f_arrdiv8_fs39_not1;
  wire f_arrdiv8_fs39_and1;
  wire f_arrdiv8_fs39_or0;
  wire f_arrdiv8_mux2to128_and0;
  wire f_arrdiv8_mux2to128_not0;
  wire f_arrdiv8_mux2to128_and1;
  wire f_arrdiv8_mux2to128_xor0;
  wire f_arrdiv8_mux2to129_and0;
  wire f_arrdiv8_mux2to129_not0;
  wire f_arrdiv8_mux2to129_and1;
  wire f_arrdiv8_mux2to129_xor0;
  wire f_arrdiv8_mux2to130_and0;
  wire f_arrdiv8_mux2to130_not0;
  wire f_arrdiv8_mux2to130_and1;
  wire f_arrdiv8_mux2to130_xor0;
  wire f_arrdiv8_mux2to131_and0;
  wire f_arrdiv8_mux2to131_not0;
  wire f_arrdiv8_mux2to131_and1;
  wire f_arrdiv8_mux2to131_xor0;
  wire f_arrdiv8_mux2to132_and0;
  wire f_arrdiv8_mux2to132_not0;
  wire f_arrdiv8_mux2to132_and1;
  wire f_arrdiv8_mux2to132_xor0;
  wire f_arrdiv8_mux2to133_and0;
  wire f_arrdiv8_mux2to133_not0;
  wire f_arrdiv8_mux2to133_and1;
  wire f_arrdiv8_mux2to133_xor0;
  wire f_arrdiv8_mux2to134_and0;
  wire f_arrdiv8_mux2to134_not0;
  wire f_arrdiv8_mux2to134_and1;
  wire f_arrdiv8_mux2to134_xor0;
  wire f_arrdiv8_not4;
  wire f_arrdiv8_fs40_xor0;
  wire f_arrdiv8_fs40_not0;
  wire f_arrdiv8_fs40_and0;
  wire f_arrdiv8_fs40_not1;
  wire f_arrdiv8_fs41_xor0;
  wire f_arrdiv8_fs41_not0;
  wire f_arrdiv8_fs41_and0;
  wire f_arrdiv8_fs41_xor1;
  wire f_arrdiv8_fs41_not1;
  wire f_arrdiv8_fs41_and1;
  wire f_arrdiv8_fs41_or0;
  wire f_arrdiv8_fs42_xor0;
  wire f_arrdiv8_fs42_not0;
  wire f_arrdiv8_fs42_and0;
  wire f_arrdiv8_fs42_xor1;
  wire f_arrdiv8_fs42_not1;
  wire f_arrdiv8_fs42_and1;
  wire f_arrdiv8_fs42_or0;
  wire f_arrdiv8_fs43_xor0;
  wire f_arrdiv8_fs43_not0;
  wire f_arrdiv8_fs43_and0;
  wire f_arrdiv8_fs43_xor1;
  wire f_arrdiv8_fs43_not1;
  wire f_arrdiv8_fs43_and1;
  wire f_arrdiv8_fs43_or0;
  wire f_arrdiv8_fs44_xor0;
  wire f_arrdiv8_fs44_not0;
  wire f_arrdiv8_fs44_and0;
  wire f_arrdiv8_fs44_xor1;
  wire f_arrdiv8_fs44_not1;
  wire f_arrdiv8_fs44_and1;
  wire f_arrdiv8_fs44_or0;
  wire f_arrdiv8_fs45_xor0;
  wire f_arrdiv8_fs45_not0;
  wire f_arrdiv8_fs45_and0;
  wire f_arrdiv8_fs45_xor1;
  wire f_arrdiv8_fs45_not1;
  wire f_arrdiv8_fs45_and1;
  wire f_arrdiv8_fs45_or0;
  wire f_arrdiv8_fs46_xor0;
  wire f_arrdiv8_fs46_not0;
  wire f_arrdiv8_fs46_and0;
  wire f_arrdiv8_fs46_xor1;
  wire f_arrdiv8_fs46_not1;
  wire f_arrdiv8_fs46_and1;
  wire f_arrdiv8_fs46_or0;
  wire f_arrdiv8_fs47_xor0;
  wire f_arrdiv8_fs47_not0;
  wire f_arrdiv8_fs47_and0;
  wire f_arrdiv8_fs47_xor1;
  wire f_arrdiv8_fs47_not1;
  wire f_arrdiv8_fs47_and1;
  wire f_arrdiv8_fs47_or0;
  wire f_arrdiv8_mux2to135_and0;
  wire f_arrdiv8_mux2to135_not0;
  wire f_arrdiv8_mux2to135_and1;
  wire f_arrdiv8_mux2to135_xor0;
  wire f_arrdiv8_mux2to136_and0;
  wire f_arrdiv8_mux2to136_not0;
  wire f_arrdiv8_mux2to136_and1;
  wire f_arrdiv8_mux2to136_xor0;
  wire f_arrdiv8_mux2to137_and0;
  wire f_arrdiv8_mux2to137_not0;
  wire f_arrdiv8_mux2to137_and1;
  wire f_arrdiv8_mux2to137_xor0;
  wire f_arrdiv8_mux2to138_and0;
  wire f_arrdiv8_mux2to138_not0;
  wire f_arrdiv8_mux2to138_and1;
  wire f_arrdiv8_mux2to138_xor0;
  wire f_arrdiv8_mux2to139_and0;
  wire f_arrdiv8_mux2to139_not0;
  wire f_arrdiv8_mux2to139_and1;
  wire f_arrdiv8_mux2to139_xor0;
  wire f_arrdiv8_mux2to140_and0;
  wire f_arrdiv8_mux2to140_not0;
  wire f_arrdiv8_mux2to140_and1;
  wire f_arrdiv8_mux2to140_xor0;
  wire f_arrdiv8_mux2to141_and0;
  wire f_arrdiv8_mux2to141_not0;
  wire f_arrdiv8_mux2to141_and1;
  wire f_arrdiv8_mux2to141_xor0;
  wire f_arrdiv8_not5;
  wire f_arrdiv8_fs48_xor0;
  wire f_arrdiv8_fs48_not0;
  wire f_arrdiv8_fs48_and0;
  wire f_arrdiv8_fs48_not1;
  wire f_arrdiv8_fs49_xor0;
  wire f_arrdiv8_fs49_not0;
  wire f_arrdiv8_fs49_and0;
  wire f_arrdiv8_fs49_xor1;
  wire f_arrdiv8_fs49_not1;
  wire f_arrdiv8_fs49_and1;
  wire f_arrdiv8_fs49_or0;
  wire f_arrdiv8_fs50_xor0;
  wire f_arrdiv8_fs50_not0;
  wire f_arrdiv8_fs50_and0;
  wire f_arrdiv8_fs50_xor1;
  wire f_arrdiv8_fs50_not1;
  wire f_arrdiv8_fs50_and1;
  wire f_arrdiv8_fs50_or0;
  wire f_arrdiv8_fs51_xor0;
  wire f_arrdiv8_fs51_not0;
  wire f_arrdiv8_fs51_and0;
  wire f_arrdiv8_fs51_xor1;
  wire f_arrdiv8_fs51_not1;
  wire f_arrdiv8_fs51_and1;
  wire f_arrdiv8_fs51_or0;
  wire f_arrdiv8_fs52_xor0;
  wire f_arrdiv8_fs52_not0;
  wire f_arrdiv8_fs52_and0;
  wire f_arrdiv8_fs52_xor1;
  wire f_arrdiv8_fs52_not1;
  wire f_arrdiv8_fs52_and1;
  wire f_arrdiv8_fs52_or0;
  wire f_arrdiv8_fs53_xor0;
  wire f_arrdiv8_fs53_not0;
  wire f_arrdiv8_fs53_and0;
  wire f_arrdiv8_fs53_xor1;
  wire f_arrdiv8_fs53_not1;
  wire f_arrdiv8_fs53_and1;
  wire f_arrdiv8_fs53_or0;
  wire f_arrdiv8_fs54_xor0;
  wire f_arrdiv8_fs54_not0;
  wire f_arrdiv8_fs54_and0;
  wire f_arrdiv8_fs54_xor1;
  wire f_arrdiv8_fs54_not1;
  wire f_arrdiv8_fs54_and1;
  wire f_arrdiv8_fs54_or0;
  wire f_arrdiv8_fs55_xor0;
  wire f_arrdiv8_fs55_not0;
  wire f_arrdiv8_fs55_and0;
  wire f_arrdiv8_fs55_xor1;
  wire f_arrdiv8_fs55_not1;
  wire f_arrdiv8_fs55_and1;
  wire f_arrdiv8_fs55_or0;
  wire f_arrdiv8_mux2to142_and0;
  wire f_arrdiv8_mux2to142_not0;
  wire f_arrdiv8_mux2to142_and1;
  wire f_arrdiv8_mux2to142_xor0;
  wire f_arrdiv8_mux2to143_and0;
  wire f_arrdiv8_mux2to143_not0;
  wire f_arrdiv8_mux2to143_and1;
  wire f_arrdiv8_mux2to143_xor0;
  wire f_arrdiv8_mux2to144_and0;
  wire f_arrdiv8_mux2to144_not0;
  wire f_arrdiv8_mux2to144_and1;
  wire f_arrdiv8_mux2to144_xor0;
  wire f_arrdiv8_mux2to145_and0;
  wire f_arrdiv8_mux2to145_not0;
  wire f_arrdiv8_mux2to145_and1;
  wire f_arrdiv8_mux2to145_xor0;
  wire f_arrdiv8_mux2to146_and0;
  wire f_arrdiv8_mux2to146_not0;
  wire f_arrdiv8_mux2to146_and1;
  wire f_arrdiv8_mux2to146_xor0;
  wire f_arrdiv8_mux2to147_and0;
  wire f_arrdiv8_mux2to147_not0;
  wire f_arrdiv8_mux2to147_and1;
  wire f_arrdiv8_mux2to147_xor0;
  wire f_arrdiv8_mux2to148_and0;
  wire f_arrdiv8_mux2to148_not0;
  wire f_arrdiv8_mux2to148_and1;
  wire f_arrdiv8_mux2to148_xor0;
  wire f_arrdiv8_not6;
  wire f_arrdiv8_fs56_xor0;
  wire f_arrdiv8_fs56_not0;
  wire f_arrdiv8_fs56_and0;
  wire f_arrdiv8_fs56_not1;
  wire f_arrdiv8_fs57_xor0;
  wire f_arrdiv8_fs57_not0;
  wire f_arrdiv8_fs57_and0;
  wire f_arrdiv8_fs57_xor1;
  wire f_arrdiv8_fs57_not1;
  wire f_arrdiv8_fs57_and1;
  wire f_arrdiv8_fs57_or0;
  wire f_arrdiv8_fs58_xor0;
  wire f_arrdiv8_fs58_not0;
  wire f_arrdiv8_fs58_and0;
  wire f_arrdiv8_fs58_xor1;
  wire f_arrdiv8_fs58_not1;
  wire f_arrdiv8_fs58_and1;
  wire f_arrdiv8_fs58_or0;
  wire f_arrdiv8_fs59_xor0;
  wire f_arrdiv8_fs59_not0;
  wire f_arrdiv8_fs59_and0;
  wire f_arrdiv8_fs59_xor1;
  wire f_arrdiv8_fs59_not1;
  wire f_arrdiv8_fs59_and1;
  wire f_arrdiv8_fs59_or0;
  wire f_arrdiv8_fs60_xor0;
  wire f_arrdiv8_fs60_not0;
  wire f_arrdiv8_fs60_and0;
  wire f_arrdiv8_fs60_xor1;
  wire f_arrdiv8_fs60_not1;
  wire f_arrdiv8_fs60_and1;
  wire f_arrdiv8_fs60_or0;
  wire f_arrdiv8_fs61_xor0;
  wire f_arrdiv8_fs61_not0;
  wire f_arrdiv8_fs61_and0;
  wire f_arrdiv8_fs61_xor1;
  wire f_arrdiv8_fs61_not1;
  wire f_arrdiv8_fs61_and1;
  wire f_arrdiv8_fs61_or0;
  wire f_arrdiv8_fs62_xor0;
  wire f_arrdiv8_fs62_not0;
  wire f_arrdiv8_fs62_and0;
  wire f_arrdiv8_fs62_xor1;
  wire f_arrdiv8_fs62_not1;
  wire f_arrdiv8_fs62_and1;
  wire f_arrdiv8_fs62_or0;
  wire f_arrdiv8_fs63_xor0;
  wire f_arrdiv8_fs63_not0;
  wire f_arrdiv8_fs63_and0;
  wire f_arrdiv8_fs63_xor1;
  wire f_arrdiv8_fs63_not1;
  wire f_arrdiv8_fs63_and1;
  wire f_arrdiv8_fs63_or0;
  wire f_arrdiv8_not7;

  assign f_arrdiv8_fs0_xor0 = a[7] ^ b[0];
  assign f_arrdiv8_fs0_not0 = ~a[7];
  assign f_arrdiv8_fs0_and0 = f_arrdiv8_fs0_not0 & b[0];
  assign f_arrdiv8_fs0_not1 = ~f_arrdiv8_fs0_xor0;
  assign f_arrdiv8_fs1_xor1 = f_arrdiv8_fs0_and0 ^ b[1];
  assign f_arrdiv8_fs1_not1 = ~b[1];
  assign f_arrdiv8_fs1_and1 = f_arrdiv8_fs1_not1 & f_arrdiv8_fs0_and0;
  assign f_arrdiv8_fs1_or0 = f_arrdiv8_fs1_and1 | b[1];
  assign f_arrdiv8_fs2_xor1 = f_arrdiv8_fs1_or0 ^ b[2];
  assign f_arrdiv8_fs2_not1 = ~b[2];
  assign f_arrdiv8_fs2_and1 = f_arrdiv8_fs2_not1 & f_arrdiv8_fs1_or0;
  assign f_arrdiv8_fs2_or0 = f_arrdiv8_fs2_and1 | b[2];
  assign f_arrdiv8_fs3_xor1 = f_arrdiv8_fs2_or0 ^ b[3];
  assign f_arrdiv8_fs3_not1 = ~b[3];
  assign f_arrdiv8_fs3_and1 = f_arrdiv8_fs3_not1 & f_arrdiv8_fs2_or0;
  assign f_arrdiv8_fs3_or0 = f_arrdiv8_fs3_and1 | b[3];
  assign f_arrdiv8_fs4_xor1 = f_arrdiv8_fs3_or0 ^ b[4];
  assign f_arrdiv8_fs4_not1 = ~b[4];
  assign f_arrdiv8_fs4_and1 = f_arrdiv8_fs4_not1 & f_arrdiv8_fs3_or0;
  assign f_arrdiv8_fs4_or0 = f_arrdiv8_fs4_and1 | b[4];
  assign f_arrdiv8_fs5_xor1 = f_arrdiv8_fs4_or0 ^ b[5];
  assign f_arrdiv8_fs5_not1 = ~b[5];
  assign f_arrdiv8_fs5_and1 = f_arrdiv8_fs5_not1 & f_arrdiv8_fs4_or0;
  assign f_arrdiv8_fs5_or0 = f_arrdiv8_fs5_and1 | b[5];
  assign f_arrdiv8_fs6_xor1 = f_arrdiv8_fs5_or0 ^ b[6];
  assign f_arrdiv8_fs6_not1 = ~b[6];
  assign f_arrdiv8_fs6_and1 = f_arrdiv8_fs6_not1 & f_arrdiv8_fs5_or0;
  assign f_arrdiv8_fs6_or0 = f_arrdiv8_fs6_and1 | b[6];
  assign f_arrdiv8_fs7_xor1 = f_arrdiv8_fs6_or0 ^ b[7];
  assign f_arrdiv8_fs7_not1 = ~b[7];
  assign f_arrdiv8_fs7_and1 = f_arrdiv8_fs7_not1 & f_arrdiv8_fs6_or0;
  assign f_arrdiv8_fs7_or0 = f_arrdiv8_fs7_and1 | b[7];
  assign f_arrdiv8_mux2to10_and0 = a[7] & f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to10_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to10_and1 = f_arrdiv8_fs0_xor0 & f_arrdiv8_mux2to10_not0;
  assign f_arrdiv8_mux2to10_xor0 = f_arrdiv8_mux2to10_and0 ^ f_arrdiv8_mux2to10_and1;
  assign f_arrdiv8_mux2to11_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to11_and1 = f_arrdiv8_fs1_xor1 & f_arrdiv8_mux2to11_not0;
  assign f_arrdiv8_mux2to12_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to12_and1 = f_arrdiv8_fs2_xor1 & f_arrdiv8_mux2to12_not0;
  assign f_arrdiv8_mux2to13_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to13_and1 = f_arrdiv8_fs3_xor1 & f_arrdiv8_mux2to13_not0;
  assign f_arrdiv8_mux2to14_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to14_and1 = f_arrdiv8_fs4_xor1 & f_arrdiv8_mux2to14_not0;
  assign f_arrdiv8_mux2to15_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to15_and1 = f_arrdiv8_fs5_xor1 & f_arrdiv8_mux2to15_not0;
  assign f_arrdiv8_mux2to16_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_mux2to16_and1 = f_arrdiv8_fs6_xor1 & f_arrdiv8_mux2to16_not0;
  assign f_arrdiv8_not0 = ~f_arrdiv8_fs7_or0;
  assign f_arrdiv8_fs8_xor0 = a[6] ^ b[0];
  assign f_arrdiv8_fs8_not0 = ~a[6];
  assign f_arrdiv8_fs8_and0 = f_arrdiv8_fs8_not0 & b[0];
  assign f_arrdiv8_fs8_not1 = ~f_arrdiv8_fs8_xor0;
  assign f_arrdiv8_fs9_xor0 = f_arrdiv8_mux2to10_xor0 ^ b[1];
  assign f_arrdiv8_fs9_not0 = ~f_arrdiv8_mux2to10_xor0;
  assign f_arrdiv8_fs9_and0 = f_arrdiv8_fs9_not0 & b[1];
  assign f_arrdiv8_fs9_xor1 = f_arrdiv8_fs8_and0 ^ f_arrdiv8_fs9_xor0;
  assign f_arrdiv8_fs9_not1 = ~f_arrdiv8_fs9_xor0;
  assign f_arrdiv8_fs9_and1 = f_arrdiv8_fs9_not1 & f_arrdiv8_fs8_and0;
  assign f_arrdiv8_fs9_or0 = f_arrdiv8_fs9_and1 | f_arrdiv8_fs9_and0;
  assign f_arrdiv8_fs10_xor0 = f_arrdiv8_mux2to11_and1 ^ b[2];
  assign f_arrdiv8_fs10_not0 = ~f_arrdiv8_mux2to11_and1;
  assign f_arrdiv8_fs10_and0 = f_arrdiv8_fs10_not0 & b[2];
  assign f_arrdiv8_fs10_xor1 = f_arrdiv8_fs9_or0 ^ f_arrdiv8_fs10_xor0;
  assign f_arrdiv8_fs10_not1 = ~f_arrdiv8_fs10_xor0;
  assign f_arrdiv8_fs10_and1 = f_arrdiv8_fs10_not1 & f_arrdiv8_fs9_or0;
  assign f_arrdiv8_fs10_or0 = f_arrdiv8_fs10_and1 | f_arrdiv8_fs10_and0;
  assign f_arrdiv8_fs11_xor0 = f_arrdiv8_mux2to12_and1 ^ b[3];
  assign f_arrdiv8_fs11_not0 = ~f_arrdiv8_mux2to12_and1;
  assign f_arrdiv8_fs11_and0 = f_arrdiv8_fs11_not0 & b[3];
  assign f_arrdiv8_fs11_xor1 = f_arrdiv8_fs10_or0 ^ f_arrdiv8_fs11_xor0;
  assign f_arrdiv8_fs11_not1 = ~f_arrdiv8_fs11_xor0;
  assign f_arrdiv8_fs11_and1 = f_arrdiv8_fs11_not1 & f_arrdiv8_fs10_or0;
  assign f_arrdiv8_fs11_or0 = f_arrdiv8_fs11_and1 | f_arrdiv8_fs11_and0;
  assign f_arrdiv8_fs12_xor0 = f_arrdiv8_mux2to13_and1 ^ b[4];
  assign f_arrdiv8_fs12_not0 = ~f_arrdiv8_mux2to13_and1;
  assign f_arrdiv8_fs12_and0 = f_arrdiv8_fs12_not0 & b[4];
  assign f_arrdiv8_fs12_xor1 = f_arrdiv8_fs11_or0 ^ f_arrdiv8_fs12_xor0;
  assign f_arrdiv8_fs12_not1 = ~f_arrdiv8_fs12_xor0;
  assign f_arrdiv8_fs12_and1 = f_arrdiv8_fs12_not1 & f_arrdiv8_fs11_or0;
  assign f_arrdiv8_fs12_or0 = f_arrdiv8_fs12_and1 | f_arrdiv8_fs12_and0;
  assign f_arrdiv8_fs13_xor0 = f_arrdiv8_mux2to14_and1 ^ b[5];
  assign f_arrdiv8_fs13_not0 = ~f_arrdiv8_mux2to14_and1;
  assign f_arrdiv8_fs13_and0 = f_arrdiv8_fs13_not0 & b[5];
  assign f_arrdiv8_fs13_xor1 = f_arrdiv8_fs12_or0 ^ f_arrdiv8_fs13_xor0;
  assign f_arrdiv8_fs13_not1 = ~f_arrdiv8_fs13_xor0;
  assign f_arrdiv8_fs13_and1 = f_arrdiv8_fs13_not1 & f_arrdiv8_fs12_or0;
  assign f_arrdiv8_fs13_or0 = f_arrdiv8_fs13_and1 | f_arrdiv8_fs13_and0;
  assign f_arrdiv8_fs14_xor0 = f_arrdiv8_mux2to15_and1 ^ b[6];
  assign f_arrdiv8_fs14_not0 = ~f_arrdiv8_mux2to15_and1;
  assign f_arrdiv8_fs14_and0 = f_arrdiv8_fs14_not0 & b[6];
  assign f_arrdiv8_fs14_xor1 = f_arrdiv8_fs13_or0 ^ f_arrdiv8_fs14_xor0;
  assign f_arrdiv8_fs14_not1 = ~f_arrdiv8_fs14_xor0;
  assign f_arrdiv8_fs14_and1 = f_arrdiv8_fs14_not1 & f_arrdiv8_fs13_or0;
  assign f_arrdiv8_fs14_or0 = f_arrdiv8_fs14_and1 | f_arrdiv8_fs14_and0;
  assign f_arrdiv8_fs15_xor0 = f_arrdiv8_mux2to16_and1 ^ b[7];
  assign f_arrdiv8_fs15_not0 = ~f_arrdiv8_mux2to16_and1;
  assign f_arrdiv8_fs15_and0 = f_arrdiv8_fs15_not0 & b[7];
  assign f_arrdiv8_fs15_xor1 = f_arrdiv8_fs14_or0 ^ f_arrdiv8_fs15_xor0;
  assign f_arrdiv8_fs15_not1 = ~f_arrdiv8_fs15_xor0;
  assign f_arrdiv8_fs15_and1 = f_arrdiv8_fs15_not1 & f_arrdiv8_fs14_or0;
  assign f_arrdiv8_fs15_or0 = f_arrdiv8_fs15_and1 | f_arrdiv8_fs15_and0;
  assign f_arrdiv8_mux2to17_and0 = a[6] & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to17_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to17_and1 = f_arrdiv8_fs8_xor0 & f_arrdiv8_mux2to17_not0;
  assign f_arrdiv8_mux2to17_xor0 = f_arrdiv8_mux2to17_and0 ^ f_arrdiv8_mux2to17_and1;
  assign f_arrdiv8_mux2to18_and0 = f_arrdiv8_mux2to10_xor0 & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to18_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to18_and1 = f_arrdiv8_fs9_xor1 & f_arrdiv8_mux2to18_not0;
  assign f_arrdiv8_mux2to18_xor0 = f_arrdiv8_mux2to18_and0 ^ f_arrdiv8_mux2to18_and1;
  assign f_arrdiv8_mux2to19_and0 = f_arrdiv8_mux2to11_and1 & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to19_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to19_and1 = f_arrdiv8_fs10_xor1 & f_arrdiv8_mux2to19_not0;
  assign f_arrdiv8_mux2to19_xor0 = f_arrdiv8_mux2to19_and0 ^ f_arrdiv8_mux2to19_and1;
  assign f_arrdiv8_mux2to110_and0 = f_arrdiv8_mux2to12_and1 & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to110_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to110_and1 = f_arrdiv8_fs11_xor1 & f_arrdiv8_mux2to110_not0;
  assign f_arrdiv8_mux2to110_xor0 = f_arrdiv8_mux2to110_and0 ^ f_arrdiv8_mux2to110_and1;
  assign f_arrdiv8_mux2to111_and0 = f_arrdiv8_mux2to13_and1 & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to111_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to111_and1 = f_arrdiv8_fs12_xor1 & f_arrdiv8_mux2to111_not0;
  assign f_arrdiv8_mux2to111_xor0 = f_arrdiv8_mux2to111_and0 ^ f_arrdiv8_mux2to111_and1;
  assign f_arrdiv8_mux2to112_and0 = f_arrdiv8_mux2to14_and1 & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to112_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to112_and1 = f_arrdiv8_fs13_xor1 & f_arrdiv8_mux2to112_not0;
  assign f_arrdiv8_mux2to112_xor0 = f_arrdiv8_mux2to112_and0 ^ f_arrdiv8_mux2to112_and1;
  assign f_arrdiv8_mux2to113_and0 = f_arrdiv8_mux2to15_and1 & f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to113_not0 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_mux2to113_and1 = f_arrdiv8_fs14_xor1 & f_arrdiv8_mux2to113_not0;
  assign f_arrdiv8_mux2to113_xor0 = f_arrdiv8_mux2to113_and0 ^ f_arrdiv8_mux2to113_and1;
  assign f_arrdiv8_not1 = ~f_arrdiv8_fs15_or0;
  assign f_arrdiv8_fs16_xor0 = a[5] ^ b[0];
  assign f_arrdiv8_fs16_not0 = ~a[5];
  assign f_arrdiv8_fs16_and0 = f_arrdiv8_fs16_not0 & b[0];
  assign f_arrdiv8_fs16_not1 = ~f_arrdiv8_fs16_xor0;
  assign f_arrdiv8_fs17_xor0 = f_arrdiv8_mux2to17_xor0 ^ b[1];
  assign f_arrdiv8_fs17_not0 = ~f_arrdiv8_mux2to17_xor0;
  assign f_arrdiv8_fs17_and0 = f_arrdiv8_fs17_not0 & b[1];
  assign f_arrdiv8_fs17_xor1 = f_arrdiv8_fs16_and0 ^ f_arrdiv8_fs17_xor0;
  assign f_arrdiv8_fs17_not1 = ~f_arrdiv8_fs17_xor0;
  assign f_arrdiv8_fs17_and1 = f_arrdiv8_fs17_not1 & f_arrdiv8_fs16_and0;
  assign f_arrdiv8_fs17_or0 = f_arrdiv8_fs17_and1 | f_arrdiv8_fs17_and0;
  assign f_arrdiv8_fs18_xor0 = f_arrdiv8_mux2to18_xor0 ^ b[2];
  assign f_arrdiv8_fs18_not0 = ~f_arrdiv8_mux2to18_xor0;
  assign f_arrdiv8_fs18_and0 = f_arrdiv8_fs18_not0 & b[2];
  assign f_arrdiv8_fs18_xor1 = f_arrdiv8_fs17_or0 ^ f_arrdiv8_fs18_xor0;
  assign f_arrdiv8_fs18_not1 = ~f_arrdiv8_fs18_xor0;
  assign f_arrdiv8_fs18_and1 = f_arrdiv8_fs18_not1 & f_arrdiv8_fs17_or0;
  assign f_arrdiv8_fs18_or0 = f_arrdiv8_fs18_and1 | f_arrdiv8_fs18_and0;
  assign f_arrdiv8_fs19_xor0 = f_arrdiv8_mux2to19_xor0 ^ b[3];
  assign f_arrdiv8_fs19_not0 = ~f_arrdiv8_mux2to19_xor0;
  assign f_arrdiv8_fs19_and0 = f_arrdiv8_fs19_not0 & b[3];
  assign f_arrdiv8_fs19_xor1 = f_arrdiv8_fs18_or0 ^ f_arrdiv8_fs19_xor0;
  assign f_arrdiv8_fs19_not1 = ~f_arrdiv8_fs19_xor0;
  assign f_arrdiv8_fs19_and1 = f_arrdiv8_fs19_not1 & f_arrdiv8_fs18_or0;
  assign f_arrdiv8_fs19_or0 = f_arrdiv8_fs19_and1 | f_arrdiv8_fs19_and0;
  assign f_arrdiv8_fs20_xor0 = f_arrdiv8_mux2to110_xor0 ^ b[4];
  assign f_arrdiv8_fs20_not0 = ~f_arrdiv8_mux2to110_xor0;
  assign f_arrdiv8_fs20_and0 = f_arrdiv8_fs20_not0 & b[4];
  assign f_arrdiv8_fs20_xor1 = f_arrdiv8_fs19_or0 ^ f_arrdiv8_fs20_xor0;
  assign f_arrdiv8_fs20_not1 = ~f_arrdiv8_fs20_xor0;
  assign f_arrdiv8_fs20_and1 = f_arrdiv8_fs20_not1 & f_arrdiv8_fs19_or0;
  assign f_arrdiv8_fs20_or0 = f_arrdiv8_fs20_and1 | f_arrdiv8_fs20_and0;
  assign f_arrdiv8_fs21_xor0 = f_arrdiv8_mux2to111_xor0 ^ b[5];
  assign f_arrdiv8_fs21_not0 = ~f_arrdiv8_mux2to111_xor0;
  assign f_arrdiv8_fs21_and0 = f_arrdiv8_fs21_not0 & b[5];
  assign f_arrdiv8_fs21_xor1 = f_arrdiv8_fs20_or0 ^ f_arrdiv8_fs21_xor0;
  assign f_arrdiv8_fs21_not1 = ~f_arrdiv8_fs21_xor0;
  assign f_arrdiv8_fs21_and1 = f_arrdiv8_fs21_not1 & f_arrdiv8_fs20_or0;
  assign f_arrdiv8_fs21_or0 = f_arrdiv8_fs21_and1 | f_arrdiv8_fs21_and0;
  assign f_arrdiv8_fs22_xor0 = f_arrdiv8_mux2to112_xor0 ^ b[6];
  assign f_arrdiv8_fs22_not0 = ~f_arrdiv8_mux2to112_xor0;
  assign f_arrdiv8_fs22_and0 = f_arrdiv8_fs22_not0 & b[6];
  assign f_arrdiv8_fs22_xor1 = f_arrdiv8_fs21_or0 ^ f_arrdiv8_fs22_xor0;
  assign f_arrdiv8_fs22_not1 = ~f_arrdiv8_fs22_xor0;
  assign f_arrdiv8_fs22_and1 = f_arrdiv8_fs22_not1 & f_arrdiv8_fs21_or0;
  assign f_arrdiv8_fs22_or0 = f_arrdiv8_fs22_and1 | f_arrdiv8_fs22_and0;
  assign f_arrdiv8_fs23_xor0 = f_arrdiv8_mux2to113_xor0 ^ b[7];
  assign f_arrdiv8_fs23_not0 = ~f_arrdiv8_mux2to113_xor0;
  assign f_arrdiv8_fs23_and0 = f_arrdiv8_fs23_not0 & b[7];
  assign f_arrdiv8_fs23_xor1 = f_arrdiv8_fs22_or0 ^ f_arrdiv8_fs23_xor0;
  assign f_arrdiv8_fs23_not1 = ~f_arrdiv8_fs23_xor0;
  assign f_arrdiv8_fs23_and1 = f_arrdiv8_fs23_not1 & f_arrdiv8_fs22_or0;
  assign f_arrdiv8_fs23_or0 = f_arrdiv8_fs23_and1 | f_arrdiv8_fs23_and0;
  assign f_arrdiv8_mux2to114_and0 = a[5] & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to114_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to114_and1 = f_arrdiv8_fs16_xor0 & f_arrdiv8_mux2to114_not0;
  assign f_arrdiv8_mux2to114_xor0 = f_arrdiv8_mux2to114_and0 ^ f_arrdiv8_mux2to114_and1;
  assign f_arrdiv8_mux2to115_and0 = f_arrdiv8_mux2to17_xor0 & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to115_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to115_and1 = f_arrdiv8_fs17_xor1 & f_arrdiv8_mux2to115_not0;
  assign f_arrdiv8_mux2to115_xor0 = f_arrdiv8_mux2to115_and0 ^ f_arrdiv8_mux2to115_and1;
  assign f_arrdiv8_mux2to116_and0 = f_arrdiv8_mux2to18_xor0 & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to116_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to116_and1 = f_arrdiv8_fs18_xor1 & f_arrdiv8_mux2to116_not0;
  assign f_arrdiv8_mux2to116_xor0 = f_arrdiv8_mux2to116_and0 ^ f_arrdiv8_mux2to116_and1;
  assign f_arrdiv8_mux2to117_and0 = f_arrdiv8_mux2to19_xor0 & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to117_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to117_and1 = f_arrdiv8_fs19_xor1 & f_arrdiv8_mux2to117_not0;
  assign f_arrdiv8_mux2to117_xor0 = f_arrdiv8_mux2to117_and0 ^ f_arrdiv8_mux2to117_and1;
  assign f_arrdiv8_mux2to118_and0 = f_arrdiv8_mux2to110_xor0 & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to118_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to118_and1 = f_arrdiv8_fs20_xor1 & f_arrdiv8_mux2to118_not0;
  assign f_arrdiv8_mux2to118_xor0 = f_arrdiv8_mux2to118_and0 ^ f_arrdiv8_mux2to118_and1;
  assign f_arrdiv8_mux2to119_and0 = f_arrdiv8_mux2to111_xor0 & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to119_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to119_and1 = f_arrdiv8_fs21_xor1 & f_arrdiv8_mux2to119_not0;
  assign f_arrdiv8_mux2to119_xor0 = f_arrdiv8_mux2to119_and0 ^ f_arrdiv8_mux2to119_and1;
  assign f_arrdiv8_mux2to120_and0 = f_arrdiv8_mux2to112_xor0 & f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to120_not0 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_mux2to120_and1 = f_arrdiv8_fs22_xor1 & f_arrdiv8_mux2to120_not0;
  assign f_arrdiv8_mux2to120_xor0 = f_arrdiv8_mux2to120_and0 ^ f_arrdiv8_mux2to120_and1;
  assign f_arrdiv8_not2 = ~f_arrdiv8_fs23_or0;
  assign f_arrdiv8_fs24_xor0 = a[4] ^ b[0];
  assign f_arrdiv8_fs24_not0 = ~a[4];
  assign f_arrdiv8_fs24_and0 = f_arrdiv8_fs24_not0 & b[0];
  assign f_arrdiv8_fs24_not1 = ~f_arrdiv8_fs24_xor0;
  assign f_arrdiv8_fs25_xor0 = f_arrdiv8_mux2to114_xor0 ^ b[1];
  assign f_arrdiv8_fs25_not0 = ~f_arrdiv8_mux2to114_xor0;
  assign f_arrdiv8_fs25_and0 = f_arrdiv8_fs25_not0 & b[1];
  assign f_arrdiv8_fs25_xor1 = f_arrdiv8_fs24_and0 ^ f_arrdiv8_fs25_xor0;
  assign f_arrdiv8_fs25_not1 = ~f_arrdiv8_fs25_xor0;
  assign f_arrdiv8_fs25_and1 = f_arrdiv8_fs25_not1 & f_arrdiv8_fs24_and0;
  assign f_arrdiv8_fs25_or0 = f_arrdiv8_fs25_and1 | f_arrdiv8_fs25_and0;
  assign f_arrdiv8_fs26_xor0 = f_arrdiv8_mux2to115_xor0 ^ b[2];
  assign f_arrdiv8_fs26_not0 = ~f_arrdiv8_mux2to115_xor0;
  assign f_arrdiv8_fs26_and0 = f_arrdiv8_fs26_not0 & b[2];
  assign f_arrdiv8_fs26_xor1 = f_arrdiv8_fs25_or0 ^ f_arrdiv8_fs26_xor0;
  assign f_arrdiv8_fs26_not1 = ~f_arrdiv8_fs26_xor0;
  assign f_arrdiv8_fs26_and1 = f_arrdiv8_fs26_not1 & f_arrdiv8_fs25_or0;
  assign f_arrdiv8_fs26_or0 = f_arrdiv8_fs26_and1 | f_arrdiv8_fs26_and0;
  assign f_arrdiv8_fs27_xor0 = f_arrdiv8_mux2to116_xor0 ^ b[3];
  assign f_arrdiv8_fs27_not0 = ~f_arrdiv8_mux2to116_xor0;
  assign f_arrdiv8_fs27_and0 = f_arrdiv8_fs27_not0 & b[3];
  assign f_arrdiv8_fs27_xor1 = f_arrdiv8_fs26_or0 ^ f_arrdiv8_fs27_xor0;
  assign f_arrdiv8_fs27_not1 = ~f_arrdiv8_fs27_xor0;
  assign f_arrdiv8_fs27_and1 = f_arrdiv8_fs27_not1 & f_arrdiv8_fs26_or0;
  assign f_arrdiv8_fs27_or0 = f_arrdiv8_fs27_and1 | f_arrdiv8_fs27_and0;
  assign f_arrdiv8_fs28_xor0 = f_arrdiv8_mux2to117_xor0 ^ b[4];
  assign f_arrdiv8_fs28_not0 = ~f_arrdiv8_mux2to117_xor0;
  assign f_arrdiv8_fs28_and0 = f_arrdiv8_fs28_not0 & b[4];
  assign f_arrdiv8_fs28_xor1 = f_arrdiv8_fs27_or0 ^ f_arrdiv8_fs28_xor0;
  assign f_arrdiv8_fs28_not1 = ~f_arrdiv8_fs28_xor0;
  assign f_arrdiv8_fs28_and1 = f_arrdiv8_fs28_not1 & f_arrdiv8_fs27_or0;
  assign f_arrdiv8_fs28_or0 = f_arrdiv8_fs28_and1 | f_arrdiv8_fs28_and0;
  assign f_arrdiv8_fs29_xor0 = f_arrdiv8_mux2to118_xor0 ^ b[5];
  assign f_arrdiv8_fs29_not0 = ~f_arrdiv8_mux2to118_xor0;
  assign f_arrdiv8_fs29_and0 = f_arrdiv8_fs29_not0 & b[5];
  assign f_arrdiv8_fs29_xor1 = f_arrdiv8_fs28_or0 ^ f_arrdiv8_fs29_xor0;
  assign f_arrdiv8_fs29_not1 = ~f_arrdiv8_fs29_xor0;
  assign f_arrdiv8_fs29_and1 = f_arrdiv8_fs29_not1 & f_arrdiv8_fs28_or0;
  assign f_arrdiv8_fs29_or0 = f_arrdiv8_fs29_and1 | f_arrdiv8_fs29_and0;
  assign f_arrdiv8_fs30_xor0 = f_arrdiv8_mux2to119_xor0 ^ b[6];
  assign f_arrdiv8_fs30_not0 = ~f_arrdiv8_mux2to119_xor0;
  assign f_arrdiv8_fs30_and0 = f_arrdiv8_fs30_not0 & b[6];
  assign f_arrdiv8_fs30_xor1 = f_arrdiv8_fs29_or0 ^ f_arrdiv8_fs30_xor0;
  assign f_arrdiv8_fs30_not1 = ~f_arrdiv8_fs30_xor0;
  assign f_arrdiv8_fs30_and1 = f_arrdiv8_fs30_not1 & f_arrdiv8_fs29_or0;
  assign f_arrdiv8_fs30_or0 = f_arrdiv8_fs30_and1 | f_arrdiv8_fs30_and0;
  assign f_arrdiv8_fs31_xor0 = f_arrdiv8_mux2to120_xor0 ^ b[7];
  assign f_arrdiv8_fs31_not0 = ~f_arrdiv8_mux2to120_xor0;
  assign f_arrdiv8_fs31_and0 = f_arrdiv8_fs31_not0 & b[7];
  assign f_arrdiv8_fs31_xor1 = f_arrdiv8_fs30_or0 ^ f_arrdiv8_fs31_xor0;
  assign f_arrdiv8_fs31_not1 = ~f_arrdiv8_fs31_xor0;
  assign f_arrdiv8_fs31_and1 = f_arrdiv8_fs31_not1 & f_arrdiv8_fs30_or0;
  assign f_arrdiv8_fs31_or0 = f_arrdiv8_fs31_and1 | f_arrdiv8_fs31_and0;
  assign f_arrdiv8_mux2to121_and0 = a[4] & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to121_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to121_and1 = f_arrdiv8_fs24_xor0 & f_arrdiv8_mux2to121_not0;
  assign f_arrdiv8_mux2to121_xor0 = f_arrdiv8_mux2to121_and0 ^ f_arrdiv8_mux2to121_and1;
  assign f_arrdiv8_mux2to122_and0 = f_arrdiv8_mux2to114_xor0 & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to122_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to122_and1 = f_arrdiv8_fs25_xor1 & f_arrdiv8_mux2to122_not0;
  assign f_arrdiv8_mux2to122_xor0 = f_arrdiv8_mux2to122_and0 ^ f_arrdiv8_mux2to122_and1;
  assign f_arrdiv8_mux2to123_and0 = f_arrdiv8_mux2to115_xor0 & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to123_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to123_and1 = f_arrdiv8_fs26_xor1 & f_arrdiv8_mux2to123_not0;
  assign f_arrdiv8_mux2to123_xor0 = f_arrdiv8_mux2to123_and0 ^ f_arrdiv8_mux2to123_and1;
  assign f_arrdiv8_mux2to124_and0 = f_arrdiv8_mux2to116_xor0 & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to124_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to124_and1 = f_arrdiv8_fs27_xor1 & f_arrdiv8_mux2to124_not0;
  assign f_arrdiv8_mux2to124_xor0 = f_arrdiv8_mux2to124_and0 ^ f_arrdiv8_mux2to124_and1;
  assign f_arrdiv8_mux2to125_and0 = f_arrdiv8_mux2to117_xor0 & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to125_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to125_and1 = f_arrdiv8_fs28_xor1 & f_arrdiv8_mux2to125_not0;
  assign f_arrdiv8_mux2to125_xor0 = f_arrdiv8_mux2to125_and0 ^ f_arrdiv8_mux2to125_and1;
  assign f_arrdiv8_mux2to126_and0 = f_arrdiv8_mux2to118_xor0 & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to126_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to126_and1 = f_arrdiv8_fs29_xor1 & f_arrdiv8_mux2to126_not0;
  assign f_arrdiv8_mux2to126_xor0 = f_arrdiv8_mux2to126_and0 ^ f_arrdiv8_mux2to126_and1;
  assign f_arrdiv8_mux2to127_and0 = f_arrdiv8_mux2to119_xor0 & f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to127_not0 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_mux2to127_and1 = f_arrdiv8_fs30_xor1 & f_arrdiv8_mux2to127_not0;
  assign f_arrdiv8_mux2to127_xor0 = f_arrdiv8_mux2to127_and0 ^ f_arrdiv8_mux2to127_and1;
  assign f_arrdiv8_not3 = ~f_arrdiv8_fs31_or0;
  assign f_arrdiv8_fs32_xor0 = a[3] ^ b[0];
  assign f_arrdiv8_fs32_not0 = ~a[3];
  assign f_arrdiv8_fs32_and0 = f_arrdiv8_fs32_not0 & b[0];
  assign f_arrdiv8_fs32_not1 = ~f_arrdiv8_fs32_xor0;
  assign f_arrdiv8_fs33_xor0 = f_arrdiv8_mux2to121_xor0 ^ b[1];
  assign f_arrdiv8_fs33_not0 = ~f_arrdiv8_mux2to121_xor0;
  assign f_arrdiv8_fs33_and0 = f_arrdiv8_fs33_not0 & b[1];
  assign f_arrdiv8_fs33_xor1 = f_arrdiv8_fs32_and0 ^ f_arrdiv8_fs33_xor0;
  assign f_arrdiv8_fs33_not1 = ~f_arrdiv8_fs33_xor0;
  assign f_arrdiv8_fs33_and1 = f_arrdiv8_fs33_not1 & f_arrdiv8_fs32_and0;
  assign f_arrdiv8_fs33_or0 = f_arrdiv8_fs33_and1 | f_arrdiv8_fs33_and0;
  assign f_arrdiv8_fs34_xor0 = f_arrdiv8_mux2to122_xor0 ^ b[2];
  assign f_arrdiv8_fs34_not0 = ~f_arrdiv8_mux2to122_xor0;
  assign f_arrdiv8_fs34_and0 = f_arrdiv8_fs34_not0 & b[2];
  assign f_arrdiv8_fs34_xor1 = f_arrdiv8_fs33_or0 ^ f_arrdiv8_fs34_xor0;
  assign f_arrdiv8_fs34_not1 = ~f_arrdiv8_fs34_xor0;
  assign f_arrdiv8_fs34_and1 = f_arrdiv8_fs34_not1 & f_arrdiv8_fs33_or0;
  assign f_arrdiv8_fs34_or0 = f_arrdiv8_fs34_and1 | f_arrdiv8_fs34_and0;
  assign f_arrdiv8_fs35_xor0 = f_arrdiv8_mux2to123_xor0 ^ b[3];
  assign f_arrdiv8_fs35_not0 = ~f_arrdiv8_mux2to123_xor0;
  assign f_arrdiv8_fs35_and0 = f_arrdiv8_fs35_not0 & b[3];
  assign f_arrdiv8_fs35_xor1 = f_arrdiv8_fs34_or0 ^ f_arrdiv8_fs35_xor0;
  assign f_arrdiv8_fs35_not1 = ~f_arrdiv8_fs35_xor0;
  assign f_arrdiv8_fs35_and1 = f_arrdiv8_fs35_not1 & f_arrdiv8_fs34_or0;
  assign f_arrdiv8_fs35_or0 = f_arrdiv8_fs35_and1 | f_arrdiv8_fs35_and0;
  assign f_arrdiv8_fs36_xor0 = f_arrdiv8_mux2to124_xor0 ^ b[4];
  assign f_arrdiv8_fs36_not0 = ~f_arrdiv8_mux2to124_xor0;
  assign f_arrdiv8_fs36_and0 = f_arrdiv8_fs36_not0 & b[4];
  assign f_arrdiv8_fs36_xor1 = f_arrdiv8_fs35_or0 ^ f_arrdiv8_fs36_xor0;
  assign f_arrdiv8_fs36_not1 = ~f_arrdiv8_fs36_xor0;
  assign f_arrdiv8_fs36_and1 = f_arrdiv8_fs36_not1 & f_arrdiv8_fs35_or0;
  assign f_arrdiv8_fs36_or0 = f_arrdiv8_fs36_and1 | f_arrdiv8_fs36_and0;
  assign f_arrdiv8_fs37_xor0 = f_arrdiv8_mux2to125_xor0 ^ b[5];
  assign f_arrdiv8_fs37_not0 = ~f_arrdiv8_mux2to125_xor0;
  assign f_arrdiv8_fs37_and0 = f_arrdiv8_fs37_not0 & b[5];
  assign f_arrdiv8_fs37_xor1 = f_arrdiv8_fs36_or0 ^ f_arrdiv8_fs37_xor0;
  assign f_arrdiv8_fs37_not1 = ~f_arrdiv8_fs37_xor0;
  assign f_arrdiv8_fs37_and1 = f_arrdiv8_fs37_not1 & f_arrdiv8_fs36_or0;
  assign f_arrdiv8_fs37_or0 = f_arrdiv8_fs37_and1 | f_arrdiv8_fs37_and0;
  assign f_arrdiv8_fs38_xor0 = f_arrdiv8_mux2to126_xor0 ^ b[6];
  assign f_arrdiv8_fs38_not0 = ~f_arrdiv8_mux2to126_xor0;
  assign f_arrdiv8_fs38_and0 = f_arrdiv8_fs38_not0 & b[6];
  assign f_arrdiv8_fs38_xor1 = f_arrdiv8_fs37_or0 ^ f_arrdiv8_fs38_xor0;
  assign f_arrdiv8_fs38_not1 = ~f_arrdiv8_fs38_xor0;
  assign f_arrdiv8_fs38_and1 = f_arrdiv8_fs38_not1 & f_arrdiv8_fs37_or0;
  assign f_arrdiv8_fs38_or0 = f_arrdiv8_fs38_and1 | f_arrdiv8_fs38_and0;
  assign f_arrdiv8_fs39_xor0 = f_arrdiv8_mux2to127_xor0 ^ b[7];
  assign f_arrdiv8_fs39_not0 = ~f_arrdiv8_mux2to127_xor0;
  assign f_arrdiv8_fs39_and0 = f_arrdiv8_fs39_not0 & b[7];
  assign f_arrdiv8_fs39_xor1 = f_arrdiv8_fs38_or0 ^ f_arrdiv8_fs39_xor0;
  assign f_arrdiv8_fs39_not1 = ~f_arrdiv8_fs39_xor0;
  assign f_arrdiv8_fs39_and1 = f_arrdiv8_fs39_not1 & f_arrdiv8_fs38_or0;
  assign f_arrdiv8_fs39_or0 = f_arrdiv8_fs39_and1 | f_arrdiv8_fs39_and0;
  assign f_arrdiv8_mux2to128_and0 = a[3] & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to128_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to128_and1 = f_arrdiv8_fs32_xor0 & f_arrdiv8_mux2to128_not0;
  assign f_arrdiv8_mux2to128_xor0 = f_arrdiv8_mux2to128_and0 ^ f_arrdiv8_mux2to128_and1;
  assign f_arrdiv8_mux2to129_and0 = f_arrdiv8_mux2to121_xor0 & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to129_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to129_and1 = f_arrdiv8_fs33_xor1 & f_arrdiv8_mux2to129_not0;
  assign f_arrdiv8_mux2to129_xor0 = f_arrdiv8_mux2to129_and0 ^ f_arrdiv8_mux2to129_and1;
  assign f_arrdiv8_mux2to130_and0 = f_arrdiv8_mux2to122_xor0 & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to130_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to130_and1 = f_arrdiv8_fs34_xor1 & f_arrdiv8_mux2to130_not0;
  assign f_arrdiv8_mux2to130_xor0 = f_arrdiv8_mux2to130_and0 ^ f_arrdiv8_mux2to130_and1;
  assign f_arrdiv8_mux2to131_and0 = f_arrdiv8_mux2to123_xor0 & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to131_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to131_and1 = f_arrdiv8_fs35_xor1 & f_arrdiv8_mux2to131_not0;
  assign f_arrdiv8_mux2to131_xor0 = f_arrdiv8_mux2to131_and0 ^ f_arrdiv8_mux2to131_and1;
  assign f_arrdiv8_mux2to132_and0 = f_arrdiv8_mux2to124_xor0 & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to132_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to132_and1 = f_arrdiv8_fs36_xor1 & f_arrdiv8_mux2to132_not0;
  assign f_arrdiv8_mux2to132_xor0 = f_arrdiv8_mux2to132_and0 ^ f_arrdiv8_mux2to132_and1;
  assign f_arrdiv8_mux2to133_and0 = f_arrdiv8_mux2to125_xor0 & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to133_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to133_and1 = f_arrdiv8_fs37_xor1 & f_arrdiv8_mux2to133_not0;
  assign f_arrdiv8_mux2to133_xor0 = f_arrdiv8_mux2to133_and0 ^ f_arrdiv8_mux2to133_and1;
  assign f_arrdiv8_mux2to134_and0 = f_arrdiv8_mux2to126_xor0 & f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to134_not0 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_mux2to134_and1 = f_arrdiv8_fs38_xor1 & f_arrdiv8_mux2to134_not0;
  assign f_arrdiv8_mux2to134_xor0 = f_arrdiv8_mux2to134_and0 ^ f_arrdiv8_mux2to134_and1;
  assign f_arrdiv8_not4 = ~f_arrdiv8_fs39_or0;
  assign f_arrdiv8_fs40_xor0 = a[2] ^ b[0];
  assign f_arrdiv8_fs40_not0 = ~a[2];
  assign f_arrdiv8_fs40_and0 = f_arrdiv8_fs40_not0 & b[0];
  assign f_arrdiv8_fs40_not1 = ~f_arrdiv8_fs40_xor0;
  assign f_arrdiv8_fs41_xor0 = f_arrdiv8_mux2to128_xor0 ^ b[1];
  assign f_arrdiv8_fs41_not0 = ~f_arrdiv8_mux2to128_xor0;
  assign f_arrdiv8_fs41_and0 = f_arrdiv8_fs41_not0 & b[1];
  assign f_arrdiv8_fs41_xor1 = f_arrdiv8_fs40_and0 ^ f_arrdiv8_fs41_xor0;
  assign f_arrdiv8_fs41_not1 = ~f_arrdiv8_fs41_xor0;
  assign f_arrdiv8_fs41_and1 = f_arrdiv8_fs41_not1 & f_arrdiv8_fs40_and0;
  assign f_arrdiv8_fs41_or0 = f_arrdiv8_fs41_and1 | f_arrdiv8_fs41_and0;
  assign f_arrdiv8_fs42_xor0 = f_arrdiv8_mux2to129_xor0 ^ b[2];
  assign f_arrdiv8_fs42_not0 = ~f_arrdiv8_mux2to129_xor0;
  assign f_arrdiv8_fs42_and0 = f_arrdiv8_fs42_not0 & b[2];
  assign f_arrdiv8_fs42_xor1 = f_arrdiv8_fs41_or0 ^ f_arrdiv8_fs42_xor0;
  assign f_arrdiv8_fs42_not1 = ~f_arrdiv8_fs42_xor0;
  assign f_arrdiv8_fs42_and1 = f_arrdiv8_fs42_not1 & f_arrdiv8_fs41_or0;
  assign f_arrdiv8_fs42_or0 = f_arrdiv8_fs42_and1 | f_arrdiv8_fs42_and0;
  assign f_arrdiv8_fs43_xor0 = f_arrdiv8_mux2to130_xor0 ^ b[3];
  assign f_arrdiv8_fs43_not0 = ~f_arrdiv8_mux2to130_xor0;
  assign f_arrdiv8_fs43_and0 = f_arrdiv8_fs43_not0 & b[3];
  assign f_arrdiv8_fs43_xor1 = f_arrdiv8_fs42_or0 ^ f_arrdiv8_fs43_xor0;
  assign f_arrdiv8_fs43_not1 = ~f_arrdiv8_fs43_xor0;
  assign f_arrdiv8_fs43_and1 = f_arrdiv8_fs43_not1 & f_arrdiv8_fs42_or0;
  assign f_arrdiv8_fs43_or0 = f_arrdiv8_fs43_and1 | f_arrdiv8_fs43_and0;
  assign f_arrdiv8_fs44_xor0 = f_arrdiv8_mux2to131_xor0 ^ b[4];
  assign f_arrdiv8_fs44_not0 = ~f_arrdiv8_mux2to131_xor0;
  assign f_arrdiv8_fs44_and0 = f_arrdiv8_fs44_not0 & b[4];
  assign f_arrdiv8_fs44_xor1 = f_arrdiv8_fs43_or0 ^ f_arrdiv8_fs44_xor0;
  assign f_arrdiv8_fs44_not1 = ~f_arrdiv8_fs44_xor0;
  assign f_arrdiv8_fs44_and1 = f_arrdiv8_fs44_not1 & f_arrdiv8_fs43_or0;
  assign f_arrdiv8_fs44_or0 = f_arrdiv8_fs44_and1 | f_arrdiv8_fs44_and0;
  assign f_arrdiv8_fs45_xor0 = f_arrdiv8_mux2to132_xor0 ^ b[5];
  assign f_arrdiv8_fs45_not0 = ~f_arrdiv8_mux2to132_xor0;
  assign f_arrdiv8_fs45_and0 = f_arrdiv8_fs45_not0 & b[5];
  assign f_arrdiv8_fs45_xor1 = f_arrdiv8_fs44_or0 ^ f_arrdiv8_fs45_xor0;
  assign f_arrdiv8_fs45_not1 = ~f_arrdiv8_fs45_xor0;
  assign f_arrdiv8_fs45_and1 = f_arrdiv8_fs45_not1 & f_arrdiv8_fs44_or0;
  assign f_arrdiv8_fs45_or0 = f_arrdiv8_fs45_and1 | f_arrdiv8_fs45_and0;
  assign f_arrdiv8_fs46_xor0 = f_arrdiv8_mux2to133_xor0 ^ b[6];
  assign f_arrdiv8_fs46_not0 = ~f_arrdiv8_mux2to133_xor0;
  assign f_arrdiv8_fs46_and0 = f_arrdiv8_fs46_not0 & b[6];
  assign f_arrdiv8_fs46_xor1 = f_arrdiv8_fs45_or0 ^ f_arrdiv8_fs46_xor0;
  assign f_arrdiv8_fs46_not1 = ~f_arrdiv8_fs46_xor0;
  assign f_arrdiv8_fs46_and1 = f_arrdiv8_fs46_not1 & f_arrdiv8_fs45_or0;
  assign f_arrdiv8_fs46_or0 = f_arrdiv8_fs46_and1 | f_arrdiv8_fs46_and0;
  assign f_arrdiv8_fs47_xor0 = f_arrdiv8_mux2to134_xor0 ^ b[7];
  assign f_arrdiv8_fs47_not0 = ~f_arrdiv8_mux2to134_xor0;
  assign f_arrdiv8_fs47_and0 = f_arrdiv8_fs47_not0 & b[7];
  assign f_arrdiv8_fs47_xor1 = f_arrdiv8_fs46_or0 ^ f_arrdiv8_fs47_xor0;
  assign f_arrdiv8_fs47_not1 = ~f_arrdiv8_fs47_xor0;
  assign f_arrdiv8_fs47_and1 = f_arrdiv8_fs47_not1 & f_arrdiv8_fs46_or0;
  assign f_arrdiv8_fs47_or0 = f_arrdiv8_fs47_and1 | f_arrdiv8_fs47_and0;
  assign f_arrdiv8_mux2to135_and0 = a[2] & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to135_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to135_and1 = f_arrdiv8_fs40_xor0 & f_arrdiv8_mux2to135_not0;
  assign f_arrdiv8_mux2to135_xor0 = f_arrdiv8_mux2to135_and0 ^ f_arrdiv8_mux2to135_and1;
  assign f_arrdiv8_mux2to136_and0 = f_arrdiv8_mux2to128_xor0 & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to136_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to136_and1 = f_arrdiv8_fs41_xor1 & f_arrdiv8_mux2to136_not0;
  assign f_arrdiv8_mux2to136_xor0 = f_arrdiv8_mux2to136_and0 ^ f_arrdiv8_mux2to136_and1;
  assign f_arrdiv8_mux2to137_and0 = f_arrdiv8_mux2to129_xor0 & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to137_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to137_and1 = f_arrdiv8_fs42_xor1 & f_arrdiv8_mux2to137_not0;
  assign f_arrdiv8_mux2to137_xor0 = f_arrdiv8_mux2to137_and0 ^ f_arrdiv8_mux2to137_and1;
  assign f_arrdiv8_mux2to138_and0 = f_arrdiv8_mux2to130_xor0 & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to138_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to138_and1 = f_arrdiv8_fs43_xor1 & f_arrdiv8_mux2to138_not0;
  assign f_arrdiv8_mux2to138_xor0 = f_arrdiv8_mux2to138_and0 ^ f_arrdiv8_mux2to138_and1;
  assign f_arrdiv8_mux2to139_and0 = f_arrdiv8_mux2to131_xor0 & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to139_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to139_and1 = f_arrdiv8_fs44_xor1 & f_arrdiv8_mux2to139_not0;
  assign f_arrdiv8_mux2to139_xor0 = f_arrdiv8_mux2to139_and0 ^ f_arrdiv8_mux2to139_and1;
  assign f_arrdiv8_mux2to140_and0 = f_arrdiv8_mux2to132_xor0 & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to140_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to140_and1 = f_arrdiv8_fs45_xor1 & f_arrdiv8_mux2to140_not0;
  assign f_arrdiv8_mux2to140_xor0 = f_arrdiv8_mux2to140_and0 ^ f_arrdiv8_mux2to140_and1;
  assign f_arrdiv8_mux2to141_and0 = f_arrdiv8_mux2to133_xor0 & f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to141_not0 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_mux2to141_and1 = f_arrdiv8_fs46_xor1 & f_arrdiv8_mux2to141_not0;
  assign f_arrdiv8_mux2to141_xor0 = f_arrdiv8_mux2to141_and0 ^ f_arrdiv8_mux2to141_and1;
  assign f_arrdiv8_not5 = ~f_arrdiv8_fs47_or0;
  assign f_arrdiv8_fs48_xor0 = a[1] ^ b[0];
  assign f_arrdiv8_fs48_not0 = ~a[1];
  assign f_arrdiv8_fs48_and0 = f_arrdiv8_fs48_not0 & b[0];
  assign f_arrdiv8_fs48_not1 = ~f_arrdiv8_fs48_xor0;
  assign f_arrdiv8_fs49_xor0 = f_arrdiv8_mux2to135_xor0 ^ b[1];
  assign f_arrdiv8_fs49_not0 = ~f_arrdiv8_mux2to135_xor0;
  assign f_arrdiv8_fs49_and0 = f_arrdiv8_fs49_not0 & b[1];
  assign f_arrdiv8_fs49_xor1 = f_arrdiv8_fs48_and0 ^ f_arrdiv8_fs49_xor0;
  assign f_arrdiv8_fs49_not1 = ~f_arrdiv8_fs49_xor0;
  assign f_arrdiv8_fs49_and1 = f_arrdiv8_fs49_not1 & f_arrdiv8_fs48_and0;
  assign f_arrdiv8_fs49_or0 = f_arrdiv8_fs49_and1 | f_arrdiv8_fs49_and0;
  assign f_arrdiv8_fs50_xor0 = f_arrdiv8_mux2to136_xor0 ^ b[2];
  assign f_arrdiv8_fs50_not0 = ~f_arrdiv8_mux2to136_xor0;
  assign f_arrdiv8_fs50_and0 = f_arrdiv8_fs50_not0 & b[2];
  assign f_arrdiv8_fs50_xor1 = f_arrdiv8_fs49_or0 ^ f_arrdiv8_fs50_xor0;
  assign f_arrdiv8_fs50_not1 = ~f_arrdiv8_fs50_xor0;
  assign f_arrdiv8_fs50_and1 = f_arrdiv8_fs50_not1 & f_arrdiv8_fs49_or0;
  assign f_arrdiv8_fs50_or0 = f_arrdiv8_fs50_and1 | f_arrdiv8_fs50_and0;
  assign f_arrdiv8_fs51_xor0 = f_arrdiv8_mux2to137_xor0 ^ b[3];
  assign f_arrdiv8_fs51_not0 = ~f_arrdiv8_mux2to137_xor0;
  assign f_arrdiv8_fs51_and0 = f_arrdiv8_fs51_not0 & b[3];
  assign f_arrdiv8_fs51_xor1 = f_arrdiv8_fs50_or0 ^ f_arrdiv8_fs51_xor0;
  assign f_arrdiv8_fs51_not1 = ~f_arrdiv8_fs51_xor0;
  assign f_arrdiv8_fs51_and1 = f_arrdiv8_fs51_not1 & f_arrdiv8_fs50_or0;
  assign f_arrdiv8_fs51_or0 = f_arrdiv8_fs51_and1 | f_arrdiv8_fs51_and0;
  assign f_arrdiv8_fs52_xor0 = f_arrdiv8_mux2to138_xor0 ^ b[4];
  assign f_arrdiv8_fs52_not0 = ~f_arrdiv8_mux2to138_xor0;
  assign f_arrdiv8_fs52_and0 = f_arrdiv8_fs52_not0 & b[4];
  assign f_arrdiv8_fs52_xor1 = f_arrdiv8_fs51_or0 ^ f_arrdiv8_fs52_xor0;
  assign f_arrdiv8_fs52_not1 = ~f_arrdiv8_fs52_xor0;
  assign f_arrdiv8_fs52_and1 = f_arrdiv8_fs52_not1 & f_arrdiv8_fs51_or0;
  assign f_arrdiv8_fs52_or0 = f_arrdiv8_fs52_and1 | f_arrdiv8_fs52_and0;
  assign f_arrdiv8_fs53_xor0 = f_arrdiv8_mux2to139_xor0 ^ b[5];
  assign f_arrdiv8_fs53_not0 = ~f_arrdiv8_mux2to139_xor0;
  assign f_arrdiv8_fs53_and0 = f_arrdiv8_fs53_not0 & b[5];
  assign f_arrdiv8_fs53_xor1 = f_arrdiv8_fs52_or0 ^ f_arrdiv8_fs53_xor0;
  assign f_arrdiv8_fs53_not1 = ~f_arrdiv8_fs53_xor0;
  assign f_arrdiv8_fs53_and1 = f_arrdiv8_fs53_not1 & f_arrdiv8_fs52_or0;
  assign f_arrdiv8_fs53_or0 = f_arrdiv8_fs53_and1 | f_arrdiv8_fs53_and0;
  assign f_arrdiv8_fs54_xor0 = f_arrdiv8_mux2to140_xor0 ^ b[6];
  assign f_arrdiv8_fs54_not0 = ~f_arrdiv8_mux2to140_xor0;
  assign f_arrdiv8_fs54_and0 = f_arrdiv8_fs54_not0 & b[6];
  assign f_arrdiv8_fs54_xor1 = f_arrdiv8_fs53_or0 ^ f_arrdiv8_fs54_xor0;
  assign f_arrdiv8_fs54_not1 = ~f_arrdiv8_fs54_xor0;
  assign f_arrdiv8_fs54_and1 = f_arrdiv8_fs54_not1 & f_arrdiv8_fs53_or0;
  assign f_arrdiv8_fs54_or0 = f_arrdiv8_fs54_and1 | f_arrdiv8_fs54_and0;
  assign f_arrdiv8_fs55_xor0 = f_arrdiv8_mux2to141_xor0 ^ b[7];
  assign f_arrdiv8_fs55_not0 = ~f_arrdiv8_mux2to141_xor0;
  assign f_arrdiv8_fs55_and0 = f_arrdiv8_fs55_not0 & b[7];
  assign f_arrdiv8_fs55_xor1 = f_arrdiv8_fs54_or0 ^ f_arrdiv8_fs55_xor0;
  assign f_arrdiv8_fs55_not1 = ~f_arrdiv8_fs55_xor0;
  assign f_arrdiv8_fs55_and1 = f_arrdiv8_fs55_not1 & f_arrdiv8_fs54_or0;
  assign f_arrdiv8_fs55_or0 = f_arrdiv8_fs55_and1 | f_arrdiv8_fs55_and0;
  assign f_arrdiv8_mux2to142_and0 = a[1] & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to142_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to142_and1 = f_arrdiv8_fs48_xor0 & f_arrdiv8_mux2to142_not0;
  assign f_arrdiv8_mux2to142_xor0 = f_arrdiv8_mux2to142_and0 ^ f_arrdiv8_mux2to142_and1;
  assign f_arrdiv8_mux2to143_and0 = f_arrdiv8_mux2to135_xor0 & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to143_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to143_and1 = f_arrdiv8_fs49_xor1 & f_arrdiv8_mux2to143_not0;
  assign f_arrdiv8_mux2to143_xor0 = f_arrdiv8_mux2to143_and0 ^ f_arrdiv8_mux2to143_and1;
  assign f_arrdiv8_mux2to144_and0 = f_arrdiv8_mux2to136_xor0 & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to144_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to144_and1 = f_arrdiv8_fs50_xor1 & f_arrdiv8_mux2to144_not0;
  assign f_arrdiv8_mux2to144_xor0 = f_arrdiv8_mux2to144_and0 ^ f_arrdiv8_mux2to144_and1;
  assign f_arrdiv8_mux2to145_and0 = f_arrdiv8_mux2to137_xor0 & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to145_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to145_and1 = f_arrdiv8_fs51_xor1 & f_arrdiv8_mux2to145_not0;
  assign f_arrdiv8_mux2to145_xor0 = f_arrdiv8_mux2to145_and0 ^ f_arrdiv8_mux2to145_and1;
  assign f_arrdiv8_mux2to146_and0 = f_arrdiv8_mux2to138_xor0 & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to146_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to146_and1 = f_arrdiv8_fs52_xor1 & f_arrdiv8_mux2to146_not0;
  assign f_arrdiv8_mux2to146_xor0 = f_arrdiv8_mux2to146_and0 ^ f_arrdiv8_mux2to146_and1;
  assign f_arrdiv8_mux2to147_and0 = f_arrdiv8_mux2to139_xor0 & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to147_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to147_and1 = f_arrdiv8_fs53_xor1 & f_arrdiv8_mux2to147_not0;
  assign f_arrdiv8_mux2to147_xor0 = f_arrdiv8_mux2to147_and0 ^ f_arrdiv8_mux2to147_and1;
  assign f_arrdiv8_mux2to148_and0 = f_arrdiv8_mux2to140_xor0 & f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to148_not0 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_mux2to148_and1 = f_arrdiv8_fs54_xor1 & f_arrdiv8_mux2to148_not0;
  assign f_arrdiv8_mux2to148_xor0 = f_arrdiv8_mux2to148_and0 ^ f_arrdiv8_mux2to148_and1;
  assign f_arrdiv8_not6 = ~f_arrdiv8_fs55_or0;
  assign f_arrdiv8_fs56_xor0 = a[0] ^ b[0];
  assign f_arrdiv8_fs56_not0 = ~a[0];
  assign f_arrdiv8_fs56_and0 = f_arrdiv8_fs56_not0 & b[0];
  assign f_arrdiv8_fs56_not1 = ~f_arrdiv8_fs56_xor0;
  assign f_arrdiv8_fs57_xor0 = f_arrdiv8_mux2to142_xor0 ^ b[1];
  assign f_arrdiv8_fs57_not0 = ~f_arrdiv8_mux2to142_xor0;
  assign f_arrdiv8_fs57_and0 = f_arrdiv8_fs57_not0 & b[1];
  assign f_arrdiv8_fs57_xor1 = f_arrdiv8_fs56_and0 ^ f_arrdiv8_fs57_xor0;
  assign f_arrdiv8_fs57_not1 = ~f_arrdiv8_fs57_xor0;
  assign f_arrdiv8_fs57_and1 = f_arrdiv8_fs57_not1 & f_arrdiv8_fs56_and0;
  assign f_arrdiv8_fs57_or0 = f_arrdiv8_fs57_and1 | f_arrdiv8_fs57_and0;
  assign f_arrdiv8_fs58_xor0 = f_arrdiv8_mux2to143_xor0 ^ b[2];
  assign f_arrdiv8_fs58_not0 = ~f_arrdiv8_mux2to143_xor0;
  assign f_arrdiv8_fs58_and0 = f_arrdiv8_fs58_not0 & b[2];
  assign f_arrdiv8_fs58_xor1 = f_arrdiv8_fs57_or0 ^ f_arrdiv8_fs58_xor0;
  assign f_arrdiv8_fs58_not1 = ~f_arrdiv8_fs58_xor0;
  assign f_arrdiv8_fs58_and1 = f_arrdiv8_fs58_not1 & f_arrdiv8_fs57_or0;
  assign f_arrdiv8_fs58_or0 = f_arrdiv8_fs58_and1 | f_arrdiv8_fs58_and0;
  assign f_arrdiv8_fs59_xor0 = f_arrdiv8_mux2to144_xor0 ^ b[3];
  assign f_arrdiv8_fs59_not0 = ~f_arrdiv8_mux2to144_xor0;
  assign f_arrdiv8_fs59_and0 = f_arrdiv8_fs59_not0 & b[3];
  assign f_arrdiv8_fs59_xor1 = f_arrdiv8_fs58_or0 ^ f_arrdiv8_fs59_xor0;
  assign f_arrdiv8_fs59_not1 = ~f_arrdiv8_fs59_xor0;
  assign f_arrdiv8_fs59_and1 = f_arrdiv8_fs59_not1 & f_arrdiv8_fs58_or0;
  assign f_arrdiv8_fs59_or0 = f_arrdiv8_fs59_and1 | f_arrdiv8_fs59_and0;
  assign f_arrdiv8_fs60_xor0 = f_arrdiv8_mux2to145_xor0 ^ b[4];
  assign f_arrdiv8_fs60_not0 = ~f_arrdiv8_mux2to145_xor0;
  assign f_arrdiv8_fs60_and0 = f_arrdiv8_fs60_not0 & b[4];
  assign f_arrdiv8_fs60_xor1 = f_arrdiv8_fs59_or0 ^ f_arrdiv8_fs60_xor0;
  assign f_arrdiv8_fs60_not1 = ~f_arrdiv8_fs60_xor0;
  assign f_arrdiv8_fs60_and1 = f_arrdiv8_fs60_not1 & f_arrdiv8_fs59_or0;
  assign f_arrdiv8_fs60_or0 = f_arrdiv8_fs60_and1 | f_arrdiv8_fs60_and0;
  assign f_arrdiv8_fs61_xor0 = f_arrdiv8_mux2to146_xor0 ^ b[5];
  assign f_arrdiv8_fs61_not0 = ~f_arrdiv8_mux2to146_xor0;
  assign f_arrdiv8_fs61_and0 = f_arrdiv8_fs61_not0 & b[5];
  assign f_arrdiv8_fs61_xor1 = f_arrdiv8_fs60_or0 ^ f_arrdiv8_fs61_xor0;
  assign f_arrdiv8_fs61_not1 = ~f_arrdiv8_fs61_xor0;
  assign f_arrdiv8_fs61_and1 = f_arrdiv8_fs61_not1 & f_arrdiv8_fs60_or0;
  assign f_arrdiv8_fs61_or0 = f_arrdiv8_fs61_and1 | f_arrdiv8_fs61_and0;
  assign f_arrdiv8_fs62_xor0 = f_arrdiv8_mux2to147_xor0 ^ b[6];
  assign f_arrdiv8_fs62_not0 = ~f_arrdiv8_mux2to147_xor0;
  assign f_arrdiv8_fs62_and0 = f_arrdiv8_fs62_not0 & b[6];
  assign f_arrdiv8_fs62_xor1 = f_arrdiv8_fs61_or0 ^ f_arrdiv8_fs62_xor0;
  assign f_arrdiv8_fs62_not1 = ~f_arrdiv8_fs62_xor0;
  assign f_arrdiv8_fs62_and1 = f_arrdiv8_fs62_not1 & f_arrdiv8_fs61_or0;
  assign f_arrdiv8_fs62_or0 = f_arrdiv8_fs62_and1 | f_arrdiv8_fs62_and0;
  assign f_arrdiv8_fs63_xor0 = f_arrdiv8_mux2to148_xor0 ^ b[7];
  assign f_arrdiv8_fs63_not0 = ~f_arrdiv8_mux2to148_xor0;
  assign f_arrdiv8_fs63_and0 = f_arrdiv8_fs63_not0 & b[7];
  assign f_arrdiv8_fs63_xor1 = f_arrdiv8_fs62_or0 ^ f_arrdiv8_fs63_xor0;
  assign f_arrdiv8_fs63_not1 = ~f_arrdiv8_fs63_xor0;
  assign f_arrdiv8_fs63_and1 = f_arrdiv8_fs63_not1 & f_arrdiv8_fs62_or0;
  assign f_arrdiv8_fs63_or0 = f_arrdiv8_fs63_and1 | f_arrdiv8_fs63_and0;
  assign f_arrdiv8_not7 = ~f_arrdiv8_fs63_or0;

  assign f_arrdiv8_out[0] = f_arrdiv8_not7;
  assign f_arrdiv8_out[1] = f_arrdiv8_not6;
  assign f_arrdiv8_out[2] = f_arrdiv8_not5;
  assign f_arrdiv8_out[3] = f_arrdiv8_not4;
  assign f_arrdiv8_out[4] = f_arrdiv8_not3;
  assign f_arrdiv8_out[5] = f_arrdiv8_not2;
  assign f_arrdiv8_out[6] = f_arrdiv8_not1;
  assign f_arrdiv8_out[7] = f_arrdiv8_not0;
endmodule