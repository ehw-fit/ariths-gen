module f_u_pg_rca4(input [3:0] a, input [3:0] b, output [4:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire constant_wire_value_0_a_0;
  wire constant_wire_value_0_b_0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_u_pg_rca4_fa0_a_0;
  wire f_u_pg_rca4_fa0_b_0;
  wire f_u_pg_rca4_fa0_y0;
  wire f_u_pg_rca4_fa0_y1;
  wire f_u_pg_rca4_fa0_constant_wire_0;
  wire f_u_pg_rca4_fa0_y2;
  wire f_u_pg_rca4_and0_constant_wire_0;
  wire f_u_pg_rca4_and0_f_u_pg_rca4_fa0_y0;
  wire f_u_pg_rca4_and0_y0;
  wire f_u_pg_rca4_or0_f_u_pg_rca4_and0_y0;
  wire f_u_pg_rca4_or0_f_u_pg_rca4_fa0_y1;
  wire f_u_pg_rca4_or0_y0;
  wire f_u_pg_rca4_fa1_a_1;
  wire f_u_pg_rca4_fa1_b_1;
  wire f_u_pg_rca4_fa1_y0;
  wire f_u_pg_rca4_fa1_y1;
  wire f_u_pg_rca4_fa1_f_u_pg_rca4_or0_y0;
  wire f_u_pg_rca4_fa1_y2;
  wire f_u_pg_rca4_and1_f_u_pg_rca4_or0_y0;
  wire f_u_pg_rca4_and1_f_u_pg_rca4_fa1_y0;
  wire f_u_pg_rca4_and1_y0;
  wire f_u_pg_rca4_or1_f_u_pg_rca4_and1_y0;
  wire f_u_pg_rca4_or1_f_u_pg_rca4_fa1_y1;
  wire f_u_pg_rca4_or1_y0;
  wire f_u_pg_rca4_fa2_a_2;
  wire f_u_pg_rca4_fa2_b_2;
  wire f_u_pg_rca4_fa2_y0;
  wire f_u_pg_rca4_fa2_y1;
  wire f_u_pg_rca4_fa2_f_u_pg_rca4_or1_y0;
  wire f_u_pg_rca4_fa2_y2;
  wire f_u_pg_rca4_and2_f_u_pg_rca4_or1_y0;
  wire f_u_pg_rca4_and2_f_u_pg_rca4_fa2_y0;
  wire f_u_pg_rca4_and2_y0;
  wire f_u_pg_rca4_or2_f_u_pg_rca4_and2_y0;
  wire f_u_pg_rca4_or2_f_u_pg_rca4_fa2_y1;
  wire f_u_pg_rca4_or2_y0;
  wire f_u_pg_rca4_fa3_a_3;
  wire f_u_pg_rca4_fa3_b_3;
  wire f_u_pg_rca4_fa3_y0;
  wire f_u_pg_rca4_fa3_y1;
  wire f_u_pg_rca4_fa3_f_u_pg_rca4_or2_y0;
  wire f_u_pg_rca4_fa3_y2;
  wire f_u_pg_rca4_and3_f_u_pg_rca4_or2_y0;
  wire f_u_pg_rca4_and3_f_u_pg_rca4_fa3_y0;
  wire f_u_pg_rca4_and3_y0;
  wire f_u_pg_rca4_or3_f_u_pg_rca4_and3_y0;
  wire f_u_pg_rca4_or3_f_u_pg_rca4_fa3_y1;
  wire f_u_pg_rca4_or3_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign constant_wire_value_0_a_0 = a_0;
  assign constant_wire_value_0_b_0 = b_0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_u_pg_rca4_fa0_a_0 = a_0;
  assign f_u_pg_rca4_fa0_b_0 = b_0;
  assign f_u_pg_rca4_fa0_constant_wire_0 = constant_wire_0;
  assign f_u_pg_rca4_fa0_y0 = f_u_pg_rca4_fa0_a_0 ^ f_u_pg_rca4_fa0_b_0;
  assign f_u_pg_rca4_fa0_y1 = f_u_pg_rca4_fa0_a_0 & f_u_pg_rca4_fa0_b_0;
  assign f_u_pg_rca4_fa0_y2 = f_u_pg_rca4_fa0_y0 ^ f_u_pg_rca4_fa0_constant_wire_0;
  assign f_u_pg_rca4_and0_constant_wire_0 = constant_wire_0;
  assign f_u_pg_rca4_and0_f_u_pg_rca4_fa0_y0 = f_u_pg_rca4_fa0_y0;
  assign f_u_pg_rca4_and0_y0 = f_u_pg_rca4_and0_constant_wire_0 & f_u_pg_rca4_and0_f_u_pg_rca4_fa0_y0;
  assign f_u_pg_rca4_or0_f_u_pg_rca4_and0_y0 = f_u_pg_rca4_and0_y0;
  assign f_u_pg_rca4_or0_f_u_pg_rca4_fa0_y1 = f_u_pg_rca4_fa0_y1;
  assign f_u_pg_rca4_or0_y0 = f_u_pg_rca4_or0_f_u_pg_rca4_and0_y0 | f_u_pg_rca4_or0_f_u_pg_rca4_fa0_y1;
  assign f_u_pg_rca4_fa1_a_1 = a_1;
  assign f_u_pg_rca4_fa1_b_1 = b_1;
  assign f_u_pg_rca4_fa1_f_u_pg_rca4_or0_y0 = f_u_pg_rca4_or0_y0;
  assign f_u_pg_rca4_fa1_y0 = f_u_pg_rca4_fa1_a_1 ^ f_u_pg_rca4_fa1_b_1;
  assign f_u_pg_rca4_fa1_y1 = f_u_pg_rca4_fa1_a_1 & f_u_pg_rca4_fa1_b_1;
  assign f_u_pg_rca4_fa1_y2 = f_u_pg_rca4_fa1_y0 ^ f_u_pg_rca4_fa1_f_u_pg_rca4_or0_y0;
  assign f_u_pg_rca4_and1_f_u_pg_rca4_or0_y0 = f_u_pg_rca4_or0_y0;
  assign f_u_pg_rca4_and1_f_u_pg_rca4_fa1_y0 = f_u_pg_rca4_fa1_y0;
  assign f_u_pg_rca4_and1_y0 = f_u_pg_rca4_and1_f_u_pg_rca4_or0_y0 & f_u_pg_rca4_and1_f_u_pg_rca4_fa1_y0;
  assign f_u_pg_rca4_or1_f_u_pg_rca4_and1_y0 = f_u_pg_rca4_and1_y0;
  assign f_u_pg_rca4_or1_f_u_pg_rca4_fa1_y1 = f_u_pg_rca4_fa1_y1;
  assign f_u_pg_rca4_or1_y0 = f_u_pg_rca4_or1_f_u_pg_rca4_and1_y0 | f_u_pg_rca4_or1_f_u_pg_rca4_fa1_y1;
  assign f_u_pg_rca4_fa2_a_2 = a_2;
  assign f_u_pg_rca4_fa2_b_2 = b_2;
  assign f_u_pg_rca4_fa2_f_u_pg_rca4_or1_y0 = f_u_pg_rca4_or1_y0;
  assign f_u_pg_rca4_fa2_y0 = f_u_pg_rca4_fa2_a_2 ^ f_u_pg_rca4_fa2_b_2;
  assign f_u_pg_rca4_fa2_y1 = f_u_pg_rca4_fa2_a_2 & f_u_pg_rca4_fa2_b_2;
  assign f_u_pg_rca4_fa2_y2 = f_u_pg_rca4_fa2_y0 ^ f_u_pg_rca4_fa2_f_u_pg_rca4_or1_y0;
  assign f_u_pg_rca4_and2_f_u_pg_rca4_or1_y0 = f_u_pg_rca4_or1_y0;
  assign f_u_pg_rca4_and2_f_u_pg_rca4_fa2_y0 = f_u_pg_rca4_fa2_y0;
  assign f_u_pg_rca4_and2_y0 = f_u_pg_rca4_and2_f_u_pg_rca4_or1_y0 & f_u_pg_rca4_and2_f_u_pg_rca4_fa2_y0;
  assign f_u_pg_rca4_or2_f_u_pg_rca4_and2_y0 = f_u_pg_rca4_and2_y0;
  assign f_u_pg_rca4_or2_f_u_pg_rca4_fa2_y1 = f_u_pg_rca4_fa2_y1;
  assign f_u_pg_rca4_or2_y0 = f_u_pg_rca4_or2_f_u_pg_rca4_and2_y0 | f_u_pg_rca4_or2_f_u_pg_rca4_fa2_y1;
  assign f_u_pg_rca4_fa3_a_3 = a_3;
  assign f_u_pg_rca4_fa3_b_3 = b_3;
  assign f_u_pg_rca4_fa3_f_u_pg_rca4_or2_y0 = f_u_pg_rca4_or2_y0;
  assign f_u_pg_rca4_fa3_y0 = f_u_pg_rca4_fa3_a_3 ^ f_u_pg_rca4_fa3_b_3;
  assign f_u_pg_rca4_fa3_y1 = f_u_pg_rca4_fa3_a_3 & f_u_pg_rca4_fa3_b_3;
  assign f_u_pg_rca4_fa3_y2 = f_u_pg_rca4_fa3_y0 ^ f_u_pg_rca4_fa3_f_u_pg_rca4_or2_y0;
  assign f_u_pg_rca4_and3_f_u_pg_rca4_or2_y0 = f_u_pg_rca4_or2_y0;
  assign f_u_pg_rca4_and3_f_u_pg_rca4_fa3_y0 = f_u_pg_rca4_fa3_y0;
  assign f_u_pg_rca4_and3_y0 = f_u_pg_rca4_and3_f_u_pg_rca4_or2_y0 & f_u_pg_rca4_and3_f_u_pg_rca4_fa3_y0;
  assign f_u_pg_rca4_or3_f_u_pg_rca4_and3_y0 = f_u_pg_rca4_and3_y0;
  assign f_u_pg_rca4_or3_f_u_pg_rca4_fa3_y1 = f_u_pg_rca4_fa3_y1;
  assign f_u_pg_rca4_or3_y0 = f_u_pg_rca4_or3_f_u_pg_rca4_and3_y0 | f_u_pg_rca4_or3_f_u_pg_rca4_fa3_y1;

  assign out[0] = f_u_pg_rca4_fa0_y2;
  assign out[1] = f_u_pg_rca4_fa1_y2;
  assign out[2] = f_u_pg_rca4_fa2_y2;
  assign out[3] = f_u_pg_rca4_fa3_y2;
  assign out[4] = f_u_pg_rca4_or3_y0;
endmodule