module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fs(input [0:0] a, input [0:0] b, input [0:0] bin, output [0:0] fs_xor1, output [0:0] fs_or0);
  wire [0:0] fs_xor0;
  wire [0:0] fs_not0;
  wire [0:0] fs_and0;
  wire [0:0] fs_not1;
  wire [0:0] fs_and1;
  xor_gate xor_gate_fs_xor0(.a(a[0]), .b(b[0]), .out(fs_xor0));
  not_gate not_gate_fs_not0(.a(a[0]), .out(fs_not0));
  and_gate and_gate_fs_and0(.a(fs_not0[0]), .b(b[0]), .out(fs_and0));
  xor_gate xor_gate_fs_xor1(.a(bin[0]), .b(fs_xor0[0]), .out(fs_xor1));
  not_gate not_gate_fs_not1(.a(fs_xor0[0]), .out(fs_not1));
  and_gate and_gate_fs_and1(.a(fs_not1[0]), .b(bin[0]), .out(fs_and1));
  or_gate or_gate_fs_or0(.a(fs_and1[0]), .b(fs_and0[0]), .out(fs_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module arrdiv12(input [11:0] a, input [11:0] b, output [11:0] arrdiv12_out);
  wire [0:0] arrdiv12_fs0_xor0;
  wire [0:0] arrdiv12_fs0_and0;
  wire [0:0] arrdiv12_fs1_xor1;
  wire [0:0] arrdiv12_fs1_or0;
  wire [0:0] arrdiv12_fs2_xor1;
  wire [0:0] arrdiv12_fs2_or0;
  wire [0:0] arrdiv12_fs3_xor1;
  wire [0:0] arrdiv12_fs3_or0;
  wire [0:0] arrdiv12_fs4_xor1;
  wire [0:0] arrdiv12_fs4_or0;
  wire [0:0] arrdiv12_fs5_xor1;
  wire [0:0] arrdiv12_fs5_or0;
  wire [0:0] arrdiv12_fs6_xor1;
  wire [0:0] arrdiv12_fs6_or0;
  wire [0:0] arrdiv12_fs7_xor1;
  wire [0:0] arrdiv12_fs7_or0;
  wire [0:0] arrdiv12_fs8_xor1;
  wire [0:0] arrdiv12_fs8_or0;
  wire [0:0] arrdiv12_fs9_xor1;
  wire [0:0] arrdiv12_fs9_or0;
  wire [0:0] arrdiv12_fs10_xor1;
  wire [0:0] arrdiv12_fs10_or0;
  wire [0:0] arrdiv12_fs11_xor1;
  wire [0:0] arrdiv12_fs11_or0;
  wire [0:0] arrdiv12_mux2to10_xor0;
  wire [0:0] arrdiv12_mux2to11_and1;
  wire [0:0] arrdiv12_mux2to12_and1;
  wire [0:0] arrdiv12_mux2to13_and1;
  wire [0:0] arrdiv12_mux2to14_and1;
  wire [0:0] arrdiv12_mux2to15_and1;
  wire [0:0] arrdiv12_mux2to16_and1;
  wire [0:0] arrdiv12_mux2to17_and1;
  wire [0:0] arrdiv12_mux2to18_and1;
  wire [0:0] arrdiv12_mux2to19_and1;
  wire [0:0] arrdiv12_mux2to110_and1;
  wire [0:0] arrdiv12_not0;
  wire [0:0] arrdiv12_fs12_xor0;
  wire [0:0] arrdiv12_fs12_and0;
  wire [0:0] arrdiv12_fs13_xor1;
  wire [0:0] arrdiv12_fs13_or0;
  wire [0:0] arrdiv12_fs14_xor1;
  wire [0:0] arrdiv12_fs14_or0;
  wire [0:0] arrdiv12_fs15_xor1;
  wire [0:0] arrdiv12_fs15_or0;
  wire [0:0] arrdiv12_fs16_xor1;
  wire [0:0] arrdiv12_fs16_or0;
  wire [0:0] arrdiv12_fs17_xor1;
  wire [0:0] arrdiv12_fs17_or0;
  wire [0:0] arrdiv12_fs18_xor1;
  wire [0:0] arrdiv12_fs18_or0;
  wire [0:0] arrdiv12_fs19_xor1;
  wire [0:0] arrdiv12_fs19_or0;
  wire [0:0] arrdiv12_fs20_xor1;
  wire [0:0] arrdiv12_fs20_or0;
  wire [0:0] arrdiv12_fs21_xor1;
  wire [0:0] arrdiv12_fs21_or0;
  wire [0:0] arrdiv12_fs22_xor1;
  wire [0:0] arrdiv12_fs22_or0;
  wire [0:0] arrdiv12_fs23_xor1;
  wire [0:0] arrdiv12_fs23_or0;
  wire [0:0] arrdiv12_mux2to111_xor0;
  wire [0:0] arrdiv12_mux2to112_xor0;
  wire [0:0] arrdiv12_mux2to113_xor0;
  wire [0:0] arrdiv12_mux2to114_xor0;
  wire [0:0] arrdiv12_mux2to115_xor0;
  wire [0:0] arrdiv12_mux2to116_xor0;
  wire [0:0] arrdiv12_mux2to117_xor0;
  wire [0:0] arrdiv12_mux2to118_xor0;
  wire [0:0] arrdiv12_mux2to119_xor0;
  wire [0:0] arrdiv12_mux2to120_xor0;
  wire [0:0] arrdiv12_mux2to121_xor0;
  wire [0:0] arrdiv12_not1;
  wire [0:0] arrdiv12_fs24_xor0;
  wire [0:0] arrdiv12_fs24_and0;
  wire [0:0] arrdiv12_fs25_xor1;
  wire [0:0] arrdiv12_fs25_or0;
  wire [0:0] arrdiv12_fs26_xor1;
  wire [0:0] arrdiv12_fs26_or0;
  wire [0:0] arrdiv12_fs27_xor1;
  wire [0:0] arrdiv12_fs27_or0;
  wire [0:0] arrdiv12_fs28_xor1;
  wire [0:0] arrdiv12_fs28_or0;
  wire [0:0] arrdiv12_fs29_xor1;
  wire [0:0] arrdiv12_fs29_or0;
  wire [0:0] arrdiv12_fs30_xor1;
  wire [0:0] arrdiv12_fs30_or0;
  wire [0:0] arrdiv12_fs31_xor1;
  wire [0:0] arrdiv12_fs31_or0;
  wire [0:0] arrdiv12_fs32_xor1;
  wire [0:0] arrdiv12_fs32_or0;
  wire [0:0] arrdiv12_fs33_xor1;
  wire [0:0] arrdiv12_fs33_or0;
  wire [0:0] arrdiv12_fs34_xor1;
  wire [0:0] arrdiv12_fs34_or0;
  wire [0:0] arrdiv12_fs35_xor1;
  wire [0:0] arrdiv12_fs35_or0;
  wire [0:0] arrdiv12_mux2to122_xor0;
  wire [0:0] arrdiv12_mux2to123_xor0;
  wire [0:0] arrdiv12_mux2to124_xor0;
  wire [0:0] arrdiv12_mux2to125_xor0;
  wire [0:0] arrdiv12_mux2to126_xor0;
  wire [0:0] arrdiv12_mux2to127_xor0;
  wire [0:0] arrdiv12_mux2to128_xor0;
  wire [0:0] arrdiv12_mux2to129_xor0;
  wire [0:0] arrdiv12_mux2to130_xor0;
  wire [0:0] arrdiv12_mux2to131_xor0;
  wire [0:0] arrdiv12_mux2to132_xor0;
  wire [0:0] arrdiv12_not2;
  wire [0:0] arrdiv12_fs36_xor0;
  wire [0:0] arrdiv12_fs36_and0;
  wire [0:0] arrdiv12_fs37_xor1;
  wire [0:0] arrdiv12_fs37_or0;
  wire [0:0] arrdiv12_fs38_xor1;
  wire [0:0] arrdiv12_fs38_or0;
  wire [0:0] arrdiv12_fs39_xor1;
  wire [0:0] arrdiv12_fs39_or0;
  wire [0:0] arrdiv12_fs40_xor1;
  wire [0:0] arrdiv12_fs40_or0;
  wire [0:0] arrdiv12_fs41_xor1;
  wire [0:0] arrdiv12_fs41_or0;
  wire [0:0] arrdiv12_fs42_xor1;
  wire [0:0] arrdiv12_fs42_or0;
  wire [0:0] arrdiv12_fs43_xor1;
  wire [0:0] arrdiv12_fs43_or0;
  wire [0:0] arrdiv12_fs44_xor1;
  wire [0:0] arrdiv12_fs44_or0;
  wire [0:0] arrdiv12_fs45_xor1;
  wire [0:0] arrdiv12_fs45_or0;
  wire [0:0] arrdiv12_fs46_xor1;
  wire [0:0] arrdiv12_fs46_or0;
  wire [0:0] arrdiv12_fs47_xor1;
  wire [0:0] arrdiv12_fs47_or0;
  wire [0:0] arrdiv12_mux2to133_xor0;
  wire [0:0] arrdiv12_mux2to134_xor0;
  wire [0:0] arrdiv12_mux2to135_xor0;
  wire [0:0] arrdiv12_mux2to136_xor0;
  wire [0:0] arrdiv12_mux2to137_xor0;
  wire [0:0] arrdiv12_mux2to138_xor0;
  wire [0:0] arrdiv12_mux2to139_xor0;
  wire [0:0] arrdiv12_mux2to140_xor0;
  wire [0:0] arrdiv12_mux2to141_xor0;
  wire [0:0] arrdiv12_mux2to142_xor0;
  wire [0:0] arrdiv12_mux2to143_xor0;
  wire [0:0] arrdiv12_not3;
  wire [0:0] arrdiv12_fs48_xor0;
  wire [0:0] arrdiv12_fs48_and0;
  wire [0:0] arrdiv12_fs49_xor1;
  wire [0:0] arrdiv12_fs49_or0;
  wire [0:0] arrdiv12_fs50_xor1;
  wire [0:0] arrdiv12_fs50_or0;
  wire [0:0] arrdiv12_fs51_xor1;
  wire [0:0] arrdiv12_fs51_or0;
  wire [0:0] arrdiv12_fs52_xor1;
  wire [0:0] arrdiv12_fs52_or0;
  wire [0:0] arrdiv12_fs53_xor1;
  wire [0:0] arrdiv12_fs53_or0;
  wire [0:0] arrdiv12_fs54_xor1;
  wire [0:0] arrdiv12_fs54_or0;
  wire [0:0] arrdiv12_fs55_xor1;
  wire [0:0] arrdiv12_fs55_or0;
  wire [0:0] arrdiv12_fs56_xor1;
  wire [0:0] arrdiv12_fs56_or0;
  wire [0:0] arrdiv12_fs57_xor1;
  wire [0:0] arrdiv12_fs57_or0;
  wire [0:0] arrdiv12_fs58_xor1;
  wire [0:0] arrdiv12_fs58_or0;
  wire [0:0] arrdiv12_fs59_xor1;
  wire [0:0] arrdiv12_fs59_or0;
  wire [0:0] arrdiv12_mux2to144_xor0;
  wire [0:0] arrdiv12_mux2to145_xor0;
  wire [0:0] arrdiv12_mux2to146_xor0;
  wire [0:0] arrdiv12_mux2to147_xor0;
  wire [0:0] arrdiv12_mux2to148_xor0;
  wire [0:0] arrdiv12_mux2to149_xor0;
  wire [0:0] arrdiv12_mux2to150_xor0;
  wire [0:0] arrdiv12_mux2to151_xor0;
  wire [0:0] arrdiv12_mux2to152_xor0;
  wire [0:0] arrdiv12_mux2to153_xor0;
  wire [0:0] arrdiv12_mux2to154_xor0;
  wire [0:0] arrdiv12_not4;
  wire [0:0] arrdiv12_fs60_xor0;
  wire [0:0] arrdiv12_fs60_and0;
  wire [0:0] arrdiv12_fs61_xor1;
  wire [0:0] arrdiv12_fs61_or0;
  wire [0:0] arrdiv12_fs62_xor1;
  wire [0:0] arrdiv12_fs62_or0;
  wire [0:0] arrdiv12_fs63_xor1;
  wire [0:0] arrdiv12_fs63_or0;
  wire [0:0] arrdiv12_fs64_xor1;
  wire [0:0] arrdiv12_fs64_or0;
  wire [0:0] arrdiv12_fs65_xor1;
  wire [0:0] arrdiv12_fs65_or0;
  wire [0:0] arrdiv12_fs66_xor1;
  wire [0:0] arrdiv12_fs66_or0;
  wire [0:0] arrdiv12_fs67_xor1;
  wire [0:0] arrdiv12_fs67_or0;
  wire [0:0] arrdiv12_fs68_xor1;
  wire [0:0] arrdiv12_fs68_or0;
  wire [0:0] arrdiv12_fs69_xor1;
  wire [0:0] arrdiv12_fs69_or0;
  wire [0:0] arrdiv12_fs70_xor1;
  wire [0:0] arrdiv12_fs70_or0;
  wire [0:0] arrdiv12_fs71_xor1;
  wire [0:0] arrdiv12_fs71_or0;
  wire [0:0] arrdiv12_mux2to155_xor0;
  wire [0:0] arrdiv12_mux2to156_xor0;
  wire [0:0] arrdiv12_mux2to157_xor0;
  wire [0:0] arrdiv12_mux2to158_xor0;
  wire [0:0] arrdiv12_mux2to159_xor0;
  wire [0:0] arrdiv12_mux2to160_xor0;
  wire [0:0] arrdiv12_mux2to161_xor0;
  wire [0:0] arrdiv12_mux2to162_xor0;
  wire [0:0] arrdiv12_mux2to163_xor0;
  wire [0:0] arrdiv12_mux2to164_xor0;
  wire [0:0] arrdiv12_mux2to165_xor0;
  wire [0:0] arrdiv12_not5;
  wire [0:0] arrdiv12_fs72_xor0;
  wire [0:0] arrdiv12_fs72_and0;
  wire [0:0] arrdiv12_fs73_xor1;
  wire [0:0] arrdiv12_fs73_or0;
  wire [0:0] arrdiv12_fs74_xor1;
  wire [0:0] arrdiv12_fs74_or0;
  wire [0:0] arrdiv12_fs75_xor1;
  wire [0:0] arrdiv12_fs75_or0;
  wire [0:0] arrdiv12_fs76_xor1;
  wire [0:0] arrdiv12_fs76_or0;
  wire [0:0] arrdiv12_fs77_xor1;
  wire [0:0] arrdiv12_fs77_or0;
  wire [0:0] arrdiv12_fs78_xor1;
  wire [0:0] arrdiv12_fs78_or0;
  wire [0:0] arrdiv12_fs79_xor1;
  wire [0:0] arrdiv12_fs79_or0;
  wire [0:0] arrdiv12_fs80_xor1;
  wire [0:0] arrdiv12_fs80_or0;
  wire [0:0] arrdiv12_fs81_xor1;
  wire [0:0] arrdiv12_fs81_or0;
  wire [0:0] arrdiv12_fs82_xor1;
  wire [0:0] arrdiv12_fs82_or0;
  wire [0:0] arrdiv12_fs83_xor1;
  wire [0:0] arrdiv12_fs83_or0;
  wire [0:0] arrdiv12_mux2to166_xor0;
  wire [0:0] arrdiv12_mux2to167_xor0;
  wire [0:0] arrdiv12_mux2to168_xor0;
  wire [0:0] arrdiv12_mux2to169_xor0;
  wire [0:0] arrdiv12_mux2to170_xor0;
  wire [0:0] arrdiv12_mux2to171_xor0;
  wire [0:0] arrdiv12_mux2to172_xor0;
  wire [0:0] arrdiv12_mux2to173_xor0;
  wire [0:0] arrdiv12_mux2to174_xor0;
  wire [0:0] arrdiv12_mux2to175_xor0;
  wire [0:0] arrdiv12_mux2to176_xor0;
  wire [0:0] arrdiv12_not6;
  wire [0:0] arrdiv12_fs84_xor0;
  wire [0:0] arrdiv12_fs84_and0;
  wire [0:0] arrdiv12_fs85_xor1;
  wire [0:0] arrdiv12_fs85_or0;
  wire [0:0] arrdiv12_fs86_xor1;
  wire [0:0] arrdiv12_fs86_or0;
  wire [0:0] arrdiv12_fs87_xor1;
  wire [0:0] arrdiv12_fs87_or0;
  wire [0:0] arrdiv12_fs88_xor1;
  wire [0:0] arrdiv12_fs88_or0;
  wire [0:0] arrdiv12_fs89_xor1;
  wire [0:0] arrdiv12_fs89_or0;
  wire [0:0] arrdiv12_fs90_xor1;
  wire [0:0] arrdiv12_fs90_or0;
  wire [0:0] arrdiv12_fs91_xor1;
  wire [0:0] arrdiv12_fs91_or0;
  wire [0:0] arrdiv12_fs92_xor1;
  wire [0:0] arrdiv12_fs92_or0;
  wire [0:0] arrdiv12_fs93_xor1;
  wire [0:0] arrdiv12_fs93_or0;
  wire [0:0] arrdiv12_fs94_xor1;
  wire [0:0] arrdiv12_fs94_or0;
  wire [0:0] arrdiv12_fs95_xor1;
  wire [0:0] arrdiv12_fs95_or0;
  wire [0:0] arrdiv12_mux2to177_xor0;
  wire [0:0] arrdiv12_mux2to178_xor0;
  wire [0:0] arrdiv12_mux2to179_xor0;
  wire [0:0] arrdiv12_mux2to180_xor0;
  wire [0:0] arrdiv12_mux2to181_xor0;
  wire [0:0] arrdiv12_mux2to182_xor0;
  wire [0:0] arrdiv12_mux2to183_xor0;
  wire [0:0] arrdiv12_mux2to184_xor0;
  wire [0:0] arrdiv12_mux2to185_xor0;
  wire [0:0] arrdiv12_mux2to186_xor0;
  wire [0:0] arrdiv12_mux2to187_xor0;
  wire [0:0] arrdiv12_not7;
  wire [0:0] arrdiv12_fs96_xor0;
  wire [0:0] arrdiv12_fs96_and0;
  wire [0:0] arrdiv12_fs97_xor1;
  wire [0:0] arrdiv12_fs97_or0;
  wire [0:0] arrdiv12_fs98_xor1;
  wire [0:0] arrdiv12_fs98_or0;
  wire [0:0] arrdiv12_fs99_xor1;
  wire [0:0] arrdiv12_fs99_or0;
  wire [0:0] arrdiv12_fs100_xor1;
  wire [0:0] arrdiv12_fs100_or0;
  wire [0:0] arrdiv12_fs101_xor1;
  wire [0:0] arrdiv12_fs101_or0;
  wire [0:0] arrdiv12_fs102_xor1;
  wire [0:0] arrdiv12_fs102_or0;
  wire [0:0] arrdiv12_fs103_xor1;
  wire [0:0] arrdiv12_fs103_or0;
  wire [0:0] arrdiv12_fs104_xor1;
  wire [0:0] arrdiv12_fs104_or0;
  wire [0:0] arrdiv12_fs105_xor1;
  wire [0:0] arrdiv12_fs105_or0;
  wire [0:0] arrdiv12_fs106_xor1;
  wire [0:0] arrdiv12_fs106_or0;
  wire [0:0] arrdiv12_fs107_xor1;
  wire [0:0] arrdiv12_fs107_or0;
  wire [0:0] arrdiv12_mux2to188_xor0;
  wire [0:0] arrdiv12_mux2to189_xor0;
  wire [0:0] arrdiv12_mux2to190_xor0;
  wire [0:0] arrdiv12_mux2to191_xor0;
  wire [0:0] arrdiv12_mux2to192_xor0;
  wire [0:0] arrdiv12_mux2to193_xor0;
  wire [0:0] arrdiv12_mux2to194_xor0;
  wire [0:0] arrdiv12_mux2to195_xor0;
  wire [0:0] arrdiv12_mux2to196_xor0;
  wire [0:0] arrdiv12_mux2to197_xor0;
  wire [0:0] arrdiv12_mux2to198_xor0;
  wire [0:0] arrdiv12_not8;
  wire [0:0] arrdiv12_fs108_xor0;
  wire [0:0] arrdiv12_fs108_and0;
  wire [0:0] arrdiv12_fs109_xor1;
  wire [0:0] arrdiv12_fs109_or0;
  wire [0:0] arrdiv12_fs110_xor1;
  wire [0:0] arrdiv12_fs110_or0;
  wire [0:0] arrdiv12_fs111_xor1;
  wire [0:0] arrdiv12_fs111_or0;
  wire [0:0] arrdiv12_fs112_xor1;
  wire [0:0] arrdiv12_fs112_or0;
  wire [0:0] arrdiv12_fs113_xor1;
  wire [0:0] arrdiv12_fs113_or0;
  wire [0:0] arrdiv12_fs114_xor1;
  wire [0:0] arrdiv12_fs114_or0;
  wire [0:0] arrdiv12_fs115_xor1;
  wire [0:0] arrdiv12_fs115_or0;
  wire [0:0] arrdiv12_fs116_xor1;
  wire [0:0] arrdiv12_fs116_or0;
  wire [0:0] arrdiv12_fs117_xor1;
  wire [0:0] arrdiv12_fs117_or0;
  wire [0:0] arrdiv12_fs118_xor1;
  wire [0:0] arrdiv12_fs118_or0;
  wire [0:0] arrdiv12_fs119_xor1;
  wire [0:0] arrdiv12_fs119_or0;
  wire [0:0] arrdiv12_mux2to199_xor0;
  wire [0:0] arrdiv12_mux2to1100_xor0;
  wire [0:0] arrdiv12_mux2to1101_xor0;
  wire [0:0] arrdiv12_mux2to1102_xor0;
  wire [0:0] arrdiv12_mux2to1103_xor0;
  wire [0:0] arrdiv12_mux2to1104_xor0;
  wire [0:0] arrdiv12_mux2to1105_xor0;
  wire [0:0] arrdiv12_mux2to1106_xor0;
  wire [0:0] arrdiv12_mux2to1107_xor0;
  wire [0:0] arrdiv12_mux2to1108_xor0;
  wire [0:0] arrdiv12_mux2to1109_xor0;
  wire [0:0] arrdiv12_not9;
  wire [0:0] arrdiv12_fs120_xor0;
  wire [0:0] arrdiv12_fs120_and0;
  wire [0:0] arrdiv12_fs121_xor1;
  wire [0:0] arrdiv12_fs121_or0;
  wire [0:0] arrdiv12_fs122_xor1;
  wire [0:0] arrdiv12_fs122_or0;
  wire [0:0] arrdiv12_fs123_xor1;
  wire [0:0] arrdiv12_fs123_or0;
  wire [0:0] arrdiv12_fs124_xor1;
  wire [0:0] arrdiv12_fs124_or0;
  wire [0:0] arrdiv12_fs125_xor1;
  wire [0:0] arrdiv12_fs125_or0;
  wire [0:0] arrdiv12_fs126_xor1;
  wire [0:0] arrdiv12_fs126_or0;
  wire [0:0] arrdiv12_fs127_xor1;
  wire [0:0] arrdiv12_fs127_or0;
  wire [0:0] arrdiv12_fs128_xor1;
  wire [0:0] arrdiv12_fs128_or0;
  wire [0:0] arrdiv12_fs129_xor1;
  wire [0:0] arrdiv12_fs129_or0;
  wire [0:0] arrdiv12_fs130_xor1;
  wire [0:0] arrdiv12_fs130_or0;
  wire [0:0] arrdiv12_fs131_xor1;
  wire [0:0] arrdiv12_fs131_or0;
  wire [0:0] arrdiv12_mux2to1110_xor0;
  wire [0:0] arrdiv12_mux2to1111_xor0;
  wire [0:0] arrdiv12_mux2to1112_xor0;
  wire [0:0] arrdiv12_mux2to1113_xor0;
  wire [0:0] arrdiv12_mux2to1114_xor0;
  wire [0:0] arrdiv12_mux2to1115_xor0;
  wire [0:0] arrdiv12_mux2to1116_xor0;
  wire [0:0] arrdiv12_mux2to1117_xor0;
  wire [0:0] arrdiv12_mux2to1118_xor0;
  wire [0:0] arrdiv12_mux2to1119_xor0;
  wire [0:0] arrdiv12_mux2to1120_xor0;
  wire [0:0] arrdiv12_not10;
  wire [0:0] arrdiv12_fs132_xor0;
  wire [0:0] arrdiv12_fs132_and0;
  wire [0:0] arrdiv12_fs133_xor1;
  wire [0:0] arrdiv12_fs133_or0;
  wire [0:0] arrdiv12_fs134_xor1;
  wire [0:0] arrdiv12_fs134_or0;
  wire [0:0] arrdiv12_fs135_xor1;
  wire [0:0] arrdiv12_fs135_or0;
  wire [0:0] arrdiv12_fs136_xor1;
  wire [0:0] arrdiv12_fs136_or0;
  wire [0:0] arrdiv12_fs137_xor1;
  wire [0:0] arrdiv12_fs137_or0;
  wire [0:0] arrdiv12_fs138_xor1;
  wire [0:0] arrdiv12_fs138_or0;
  wire [0:0] arrdiv12_fs139_xor1;
  wire [0:0] arrdiv12_fs139_or0;
  wire [0:0] arrdiv12_fs140_xor1;
  wire [0:0] arrdiv12_fs140_or0;
  wire [0:0] arrdiv12_fs141_xor1;
  wire [0:0] arrdiv12_fs141_or0;
  wire [0:0] arrdiv12_fs142_xor1;
  wire [0:0] arrdiv12_fs142_or0;
  wire [0:0] arrdiv12_fs143_xor1;
  wire [0:0] arrdiv12_fs143_or0;
  wire [0:0] arrdiv12_not11;

  fs fs_arrdiv12_fs0_out(.a(a[11]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs0_xor0), .fs_or0(arrdiv12_fs0_and0));
  fs fs_arrdiv12_fs1_out(.a(1'b0), .b(b[1]), .bin(arrdiv12_fs0_and0[0]), .fs_xor1(arrdiv12_fs1_xor1), .fs_or0(arrdiv12_fs1_or0));
  fs fs_arrdiv12_fs2_out(.a(1'b0), .b(b[2]), .bin(arrdiv12_fs1_or0[0]), .fs_xor1(arrdiv12_fs2_xor1), .fs_or0(arrdiv12_fs2_or0));
  fs fs_arrdiv12_fs3_out(.a(1'b0), .b(b[3]), .bin(arrdiv12_fs2_or0[0]), .fs_xor1(arrdiv12_fs3_xor1), .fs_or0(arrdiv12_fs3_or0));
  fs fs_arrdiv12_fs4_out(.a(1'b0), .b(b[4]), .bin(arrdiv12_fs3_or0[0]), .fs_xor1(arrdiv12_fs4_xor1), .fs_or0(arrdiv12_fs4_or0));
  fs fs_arrdiv12_fs5_out(.a(1'b0), .b(b[5]), .bin(arrdiv12_fs4_or0[0]), .fs_xor1(arrdiv12_fs5_xor1), .fs_or0(arrdiv12_fs5_or0));
  fs fs_arrdiv12_fs6_out(.a(1'b0), .b(b[6]), .bin(arrdiv12_fs5_or0[0]), .fs_xor1(arrdiv12_fs6_xor1), .fs_or0(arrdiv12_fs6_or0));
  fs fs_arrdiv12_fs7_out(.a(1'b0), .b(b[7]), .bin(arrdiv12_fs6_or0[0]), .fs_xor1(arrdiv12_fs7_xor1), .fs_or0(arrdiv12_fs7_or0));
  fs fs_arrdiv12_fs8_out(.a(1'b0), .b(b[8]), .bin(arrdiv12_fs7_or0[0]), .fs_xor1(arrdiv12_fs8_xor1), .fs_or0(arrdiv12_fs8_or0));
  fs fs_arrdiv12_fs9_out(.a(1'b0), .b(b[9]), .bin(arrdiv12_fs8_or0[0]), .fs_xor1(arrdiv12_fs9_xor1), .fs_or0(arrdiv12_fs9_or0));
  fs fs_arrdiv12_fs10_out(.a(1'b0), .b(b[10]), .bin(arrdiv12_fs9_or0[0]), .fs_xor1(arrdiv12_fs10_xor1), .fs_or0(arrdiv12_fs10_or0));
  fs fs_arrdiv12_fs11_out(.a(1'b0), .b(b[11]), .bin(arrdiv12_fs10_or0[0]), .fs_xor1(arrdiv12_fs11_xor1), .fs_or0(arrdiv12_fs11_or0));
  mux2to1 mux2to1_arrdiv12_mux2to10_out(.d0(arrdiv12_fs0_xor0[0]), .d1(a[11]), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to10_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to11_out(.d0(arrdiv12_fs1_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to11_and1));
  mux2to1 mux2to1_arrdiv12_mux2to12_out(.d0(arrdiv12_fs2_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to12_and1));
  mux2to1 mux2to1_arrdiv12_mux2to13_out(.d0(arrdiv12_fs3_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to13_and1));
  mux2to1 mux2to1_arrdiv12_mux2to14_out(.d0(arrdiv12_fs4_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to14_and1));
  mux2to1 mux2to1_arrdiv12_mux2to15_out(.d0(arrdiv12_fs5_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to15_and1));
  mux2to1 mux2to1_arrdiv12_mux2to16_out(.d0(arrdiv12_fs6_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to16_and1));
  mux2to1 mux2to1_arrdiv12_mux2to17_out(.d0(arrdiv12_fs7_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to17_and1));
  mux2to1 mux2to1_arrdiv12_mux2to18_out(.d0(arrdiv12_fs8_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to18_and1));
  mux2to1 mux2to1_arrdiv12_mux2to19_out(.d0(arrdiv12_fs9_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to19_and1));
  mux2to1 mux2to1_arrdiv12_mux2to110_out(.d0(arrdiv12_fs10_xor1[0]), .d1(1'b0), .sel(arrdiv12_fs11_or0[0]), .mux2to1_xor0(arrdiv12_mux2to110_and1));
  not_gate not_gate_arrdiv12_not0(.a(arrdiv12_fs11_or0[0]), .out(arrdiv12_not0));
  fs fs_arrdiv12_fs12_out(.a(a[10]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs12_xor0), .fs_or0(arrdiv12_fs12_and0));
  fs fs_arrdiv12_fs13_out(.a(arrdiv12_mux2to10_xor0[0]), .b(b[1]), .bin(arrdiv12_fs12_and0[0]), .fs_xor1(arrdiv12_fs13_xor1), .fs_or0(arrdiv12_fs13_or0));
  fs fs_arrdiv12_fs14_out(.a(arrdiv12_mux2to11_and1[0]), .b(b[2]), .bin(arrdiv12_fs13_or0[0]), .fs_xor1(arrdiv12_fs14_xor1), .fs_or0(arrdiv12_fs14_or0));
  fs fs_arrdiv12_fs15_out(.a(arrdiv12_mux2to12_and1[0]), .b(b[3]), .bin(arrdiv12_fs14_or0[0]), .fs_xor1(arrdiv12_fs15_xor1), .fs_or0(arrdiv12_fs15_or0));
  fs fs_arrdiv12_fs16_out(.a(arrdiv12_mux2to13_and1[0]), .b(b[4]), .bin(arrdiv12_fs15_or0[0]), .fs_xor1(arrdiv12_fs16_xor1), .fs_or0(arrdiv12_fs16_or0));
  fs fs_arrdiv12_fs17_out(.a(arrdiv12_mux2to14_and1[0]), .b(b[5]), .bin(arrdiv12_fs16_or0[0]), .fs_xor1(arrdiv12_fs17_xor1), .fs_or0(arrdiv12_fs17_or0));
  fs fs_arrdiv12_fs18_out(.a(arrdiv12_mux2to15_and1[0]), .b(b[6]), .bin(arrdiv12_fs17_or0[0]), .fs_xor1(arrdiv12_fs18_xor1), .fs_or0(arrdiv12_fs18_or0));
  fs fs_arrdiv12_fs19_out(.a(arrdiv12_mux2to16_and1[0]), .b(b[7]), .bin(arrdiv12_fs18_or0[0]), .fs_xor1(arrdiv12_fs19_xor1), .fs_or0(arrdiv12_fs19_or0));
  fs fs_arrdiv12_fs20_out(.a(arrdiv12_mux2to17_and1[0]), .b(b[8]), .bin(arrdiv12_fs19_or0[0]), .fs_xor1(arrdiv12_fs20_xor1), .fs_or0(arrdiv12_fs20_or0));
  fs fs_arrdiv12_fs21_out(.a(arrdiv12_mux2to18_and1[0]), .b(b[9]), .bin(arrdiv12_fs20_or0[0]), .fs_xor1(arrdiv12_fs21_xor1), .fs_or0(arrdiv12_fs21_or0));
  fs fs_arrdiv12_fs22_out(.a(arrdiv12_mux2to19_and1[0]), .b(b[10]), .bin(arrdiv12_fs21_or0[0]), .fs_xor1(arrdiv12_fs22_xor1), .fs_or0(arrdiv12_fs22_or0));
  fs fs_arrdiv12_fs23_out(.a(arrdiv12_mux2to110_and1[0]), .b(b[11]), .bin(arrdiv12_fs22_or0[0]), .fs_xor1(arrdiv12_fs23_xor1), .fs_or0(arrdiv12_fs23_or0));
  mux2to1 mux2to1_arrdiv12_mux2to111_out(.d0(arrdiv12_fs12_xor0[0]), .d1(a[10]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to111_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to112_out(.d0(arrdiv12_fs13_xor1[0]), .d1(arrdiv12_mux2to10_xor0[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to112_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to113_out(.d0(arrdiv12_fs14_xor1[0]), .d1(arrdiv12_mux2to11_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to113_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to114_out(.d0(arrdiv12_fs15_xor1[0]), .d1(arrdiv12_mux2to12_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to114_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to115_out(.d0(arrdiv12_fs16_xor1[0]), .d1(arrdiv12_mux2to13_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to115_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to116_out(.d0(arrdiv12_fs17_xor1[0]), .d1(arrdiv12_mux2to14_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to116_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to117_out(.d0(arrdiv12_fs18_xor1[0]), .d1(arrdiv12_mux2to15_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to117_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to118_out(.d0(arrdiv12_fs19_xor1[0]), .d1(arrdiv12_mux2to16_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to118_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to119_out(.d0(arrdiv12_fs20_xor1[0]), .d1(arrdiv12_mux2to17_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to119_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to120_out(.d0(arrdiv12_fs21_xor1[0]), .d1(arrdiv12_mux2to18_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to120_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to121_out(.d0(arrdiv12_fs22_xor1[0]), .d1(arrdiv12_mux2to19_and1[0]), .sel(arrdiv12_fs23_or0[0]), .mux2to1_xor0(arrdiv12_mux2to121_xor0));
  not_gate not_gate_arrdiv12_not1(.a(arrdiv12_fs23_or0[0]), .out(arrdiv12_not1));
  fs fs_arrdiv12_fs24_out(.a(a[9]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs24_xor0), .fs_or0(arrdiv12_fs24_and0));
  fs fs_arrdiv12_fs25_out(.a(arrdiv12_mux2to111_xor0[0]), .b(b[1]), .bin(arrdiv12_fs24_and0[0]), .fs_xor1(arrdiv12_fs25_xor1), .fs_or0(arrdiv12_fs25_or0));
  fs fs_arrdiv12_fs26_out(.a(arrdiv12_mux2to112_xor0[0]), .b(b[2]), .bin(arrdiv12_fs25_or0[0]), .fs_xor1(arrdiv12_fs26_xor1), .fs_or0(arrdiv12_fs26_or0));
  fs fs_arrdiv12_fs27_out(.a(arrdiv12_mux2to113_xor0[0]), .b(b[3]), .bin(arrdiv12_fs26_or0[0]), .fs_xor1(arrdiv12_fs27_xor1), .fs_or0(arrdiv12_fs27_or0));
  fs fs_arrdiv12_fs28_out(.a(arrdiv12_mux2to114_xor0[0]), .b(b[4]), .bin(arrdiv12_fs27_or0[0]), .fs_xor1(arrdiv12_fs28_xor1), .fs_or0(arrdiv12_fs28_or0));
  fs fs_arrdiv12_fs29_out(.a(arrdiv12_mux2to115_xor0[0]), .b(b[5]), .bin(arrdiv12_fs28_or0[0]), .fs_xor1(arrdiv12_fs29_xor1), .fs_or0(arrdiv12_fs29_or0));
  fs fs_arrdiv12_fs30_out(.a(arrdiv12_mux2to116_xor0[0]), .b(b[6]), .bin(arrdiv12_fs29_or0[0]), .fs_xor1(arrdiv12_fs30_xor1), .fs_or0(arrdiv12_fs30_or0));
  fs fs_arrdiv12_fs31_out(.a(arrdiv12_mux2to117_xor0[0]), .b(b[7]), .bin(arrdiv12_fs30_or0[0]), .fs_xor1(arrdiv12_fs31_xor1), .fs_or0(arrdiv12_fs31_or0));
  fs fs_arrdiv12_fs32_out(.a(arrdiv12_mux2to118_xor0[0]), .b(b[8]), .bin(arrdiv12_fs31_or0[0]), .fs_xor1(arrdiv12_fs32_xor1), .fs_or0(arrdiv12_fs32_or0));
  fs fs_arrdiv12_fs33_out(.a(arrdiv12_mux2to119_xor0[0]), .b(b[9]), .bin(arrdiv12_fs32_or0[0]), .fs_xor1(arrdiv12_fs33_xor1), .fs_or0(arrdiv12_fs33_or0));
  fs fs_arrdiv12_fs34_out(.a(arrdiv12_mux2to120_xor0[0]), .b(b[10]), .bin(arrdiv12_fs33_or0[0]), .fs_xor1(arrdiv12_fs34_xor1), .fs_or0(arrdiv12_fs34_or0));
  fs fs_arrdiv12_fs35_out(.a(arrdiv12_mux2to121_xor0[0]), .b(b[11]), .bin(arrdiv12_fs34_or0[0]), .fs_xor1(arrdiv12_fs35_xor1), .fs_or0(arrdiv12_fs35_or0));
  mux2to1 mux2to1_arrdiv12_mux2to122_out(.d0(arrdiv12_fs24_xor0[0]), .d1(a[9]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to122_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to123_out(.d0(arrdiv12_fs25_xor1[0]), .d1(arrdiv12_mux2to111_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to123_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to124_out(.d0(arrdiv12_fs26_xor1[0]), .d1(arrdiv12_mux2to112_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to124_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to125_out(.d0(arrdiv12_fs27_xor1[0]), .d1(arrdiv12_mux2to113_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to125_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to126_out(.d0(arrdiv12_fs28_xor1[0]), .d1(arrdiv12_mux2to114_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to126_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to127_out(.d0(arrdiv12_fs29_xor1[0]), .d1(arrdiv12_mux2to115_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to127_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to128_out(.d0(arrdiv12_fs30_xor1[0]), .d1(arrdiv12_mux2to116_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to128_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to129_out(.d0(arrdiv12_fs31_xor1[0]), .d1(arrdiv12_mux2to117_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to129_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to130_out(.d0(arrdiv12_fs32_xor1[0]), .d1(arrdiv12_mux2to118_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to130_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to131_out(.d0(arrdiv12_fs33_xor1[0]), .d1(arrdiv12_mux2to119_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to131_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to132_out(.d0(arrdiv12_fs34_xor1[0]), .d1(arrdiv12_mux2to120_xor0[0]), .sel(arrdiv12_fs35_or0[0]), .mux2to1_xor0(arrdiv12_mux2to132_xor0));
  not_gate not_gate_arrdiv12_not2(.a(arrdiv12_fs35_or0[0]), .out(arrdiv12_not2));
  fs fs_arrdiv12_fs36_out(.a(a[8]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs36_xor0), .fs_or0(arrdiv12_fs36_and0));
  fs fs_arrdiv12_fs37_out(.a(arrdiv12_mux2to122_xor0[0]), .b(b[1]), .bin(arrdiv12_fs36_and0[0]), .fs_xor1(arrdiv12_fs37_xor1), .fs_or0(arrdiv12_fs37_or0));
  fs fs_arrdiv12_fs38_out(.a(arrdiv12_mux2to123_xor0[0]), .b(b[2]), .bin(arrdiv12_fs37_or0[0]), .fs_xor1(arrdiv12_fs38_xor1), .fs_or0(arrdiv12_fs38_or0));
  fs fs_arrdiv12_fs39_out(.a(arrdiv12_mux2to124_xor0[0]), .b(b[3]), .bin(arrdiv12_fs38_or0[0]), .fs_xor1(arrdiv12_fs39_xor1), .fs_or0(arrdiv12_fs39_or0));
  fs fs_arrdiv12_fs40_out(.a(arrdiv12_mux2to125_xor0[0]), .b(b[4]), .bin(arrdiv12_fs39_or0[0]), .fs_xor1(arrdiv12_fs40_xor1), .fs_or0(arrdiv12_fs40_or0));
  fs fs_arrdiv12_fs41_out(.a(arrdiv12_mux2to126_xor0[0]), .b(b[5]), .bin(arrdiv12_fs40_or0[0]), .fs_xor1(arrdiv12_fs41_xor1), .fs_or0(arrdiv12_fs41_or0));
  fs fs_arrdiv12_fs42_out(.a(arrdiv12_mux2to127_xor0[0]), .b(b[6]), .bin(arrdiv12_fs41_or0[0]), .fs_xor1(arrdiv12_fs42_xor1), .fs_or0(arrdiv12_fs42_or0));
  fs fs_arrdiv12_fs43_out(.a(arrdiv12_mux2to128_xor0[0]), .b(b[7]), .bin(arrdiv12_fs42_or0[0]), .fs_xor1(arrdiv12_fs43_xor1), .fs_or0(arrdiv12_fs43_or0));
  fs fs_arrdiv12_fs44_out(.a(arrdiv12_mux2to129_xor0[0]), .b(b[8]), .bin(arrdiv12_fs43_or0[0]), .fs_xor1(arrdiv12_fs44_xor1), .fs_or0(arrdiv12_fs44_or0));
  fs fs_arrdiv12_fs45_out(.a(arrdiv12_mux2to130_xor0[0]), .b(b[9]), .bin(arrdiv12_fs44_or0[0]), .fs_xor1(arrdiv12_fs45_xor1), .fs_or0(arrdiv12_fs45_or0));
  fs fs_arrdiv12_fs46_out(.a(arrdiv12_mux2to131_xor0[0]), .b(b[10]), .bin(arrdiv12_fs45_or0[0]), .fs_xor1(arrdiv12_fs46_xor1), .fs_or0(arrdiv12_fs46_or0));
  fs fs_arrdiv12_fs47_out(.a(arrdiv12_mux2to132_xor0[0]), .b(b[11]), .bin(arrdiv12_fs46_or0[0]), .fs_xor1(arrdiv12_fs47_xor1), .fs_or0(arrdiv12_fs47_or0));
  mux2to1 mux2to1_arrdiv12_mux2to133_out(.d0(arrdiv12_fs36_xor0[0]), .d1(a[8]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to133_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to134_out(.d0(arrdiv12_fs37_xor1[0]), .d1(arrdiv12_mux2to122_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to134_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to135_out(.d0(arrdiv12_fs38_xor1[0]), .d1(arrdiv12_mux2to123_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to135_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to136_out(.d0(arrdiv12_fs39_xor1[0]), .d1(arrdiv12_mux2to124_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to136_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to137_out(.d0(arrdiv12_fs40_xor1[0]), .d1(arrdiv12_mux2to125_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to137_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to138_out(.d0(arrdiv12_fs41_xor1[0]), .d1(arrdiv12_mux2to126_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to138_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to139_out(.d0(arrdiv12_fs42_xor1[0]), .d1(arrdiv12_mux2to127_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to139_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to140_out(.d0(arrdiv12_fs43_xor1[0]), .d1(arrdiv12_mux2to128_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to140_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to141_out(.d0(arrdiv12_fs44_xor1[0]), .d1(arrdiv12_mux2to129_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to141_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to142_out(.d0(arrdiv12_fs45_xor1[0]), .d1(arrdiv12_mux2to130_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to142_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to143_out(.d0(arrdiv12_fs46_xor1[0]), .d1(arrdiv12_mux2to131_xor0[0]), .sel(arrdiv12_fs47_or0[0]), .mux2to1_xor0(arrdiv12_mux2to143_xor0));
  not_gate not_gate_arrdiv12_not3(.a(arrdiv12_fs47_or0[0]), .out(arrdiv12_not3));
  fs fs_arrdiv12_fs48_out(.a(a[7]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs48_xor0), .fs_or0(arrdiv12_fs48_and0));
  fs fs_arrdiv12_fs49_out(.a(arrdiv12_mux2to133_xor0[0]), .b(b[1]), .bin(arrdiv12_fs48_and0[0]), .fs_xor1(arrdiv12_fs49_xor1), .fs_or0(arrdiv12_fs49_or0));
  fs fs_arrdiv12_fs50_out(.a(arrdiv12_mux2to134_xor0[0]), .b(b[2]), .bin(arrdiv12_fs49_or0[0]), .fs_xor1(arrdiv12_fs50_xor1), .fs_or0(arrdiv12_fs50_or0));
  fs fs_arrdiv12_fs51_out(.a(arrdiv12_mux2to135_xor0[0]), .b(b[3]), .bin(arrdiv12_fs50_or0[0]), .fs_xor1(arrdiv12_fs51_xor1), .fs_or0(arrdiv12_fs51_or0));
  fs fs_arrdiv12_fs52_out(.a(arrdiv12_mux2to136_xor0[0]), .b(b[4]), .bin(arrdiv12_fs51_or0[0]), .fs_xor1(arrdiv12_fs52_xor1), .fs_or0(arrdiv12_fs52_or0));
  fs fs_arrdiv12_fs53_out(.a(arrdiv12_mux2to137_xor0[0]), .b(b[5]), .bin(arrdiv12_fs52_or0[0]), .fs_xor1(arrdiv12_fs53_xor1), .fs_or0(arrdiv12_fs53_or0));
  fs fs_arrdiv12_fs54_out(.a(arrdiv12_mux2to138_xor0[0]), .b(b[6]), .bin(arrdiv12_fs53_or0[0]), .fs_xor1(arrdiv12_fs54_xor1), .fs_or0(arrdiv12_fs54_or0));
  fs fs_arrdiv12_fs55_out(.a(arrdiv12_mux2to139_xor0[0]), .b(b[7]), .bin(arrdiv12_fs54_or0[0]), .fs_xor1(arrdiv12_fs55_xor1), .fs_or0(arrdiv12_fs55_or0));
  fs fs_arrdiv12_fs56_out(.a(arrdiv12_mux2to140_xor0[0]), .b(b[8]), .bin(arrdiv12_fs55_or0[0]), .fs_xor1(arrdiv12_fs56_xor1), .fs_or0(arrdiv12_fs56_or0));
  fs fs_arrdiv12_fs57_out(.a(arrdiv12_mux2to141_xor0[0]), .b(b[9]), .bin(arrdiv12_fs56_or0[0]), .fs_xor1(arrdiv12_fs57_xor1), .fs_or0(arrdiv12_fs57_or0));
  fs fs_arrdiv12_fs58_out(.a(arrdiv12_mux2to142_xor0[0]), .b(b[10]), .bin(arrdiv12_fs57_or0[0]), .fs_xor1(arrdiv12_fs58_xor1), .fs_or0(arrdiv12_fs58_or0));
  fs fs_arrdiv12_fs59_out(.a(arrdiv12_mux2to143_xor0[0]), .b(b[11]), .bin(arrdiv12_fs58_or0[0]), .fs_xor1(arrdiv12_fs59_xor1), .fs_or0(arrdiv12_fs59_or0));
  mux2to1 mux2to1_arrdiv12_mux2to144_out(.d0(arrdiv12_fs48_xor0[0]), .d1(a[7]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to144_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to145_out(.d0(arrdiv12_fs49_xor1[0]), .d1(arrdiv12_mux2to133_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to145_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to146_out(.d0(arrdiv12_fs50_xor1[0]), .d1(arrdiv12_mux2to134_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to146_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to147_out(.d0(arrdiv12_fs51_xor1[0]), .d1(arrdiv12_mux2to135_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to147_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to148_out(.d0(arrdiv12_fs52_xor1[0]), .d1(arrdiv12_mux2to136_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to148_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to149_out(.d0(arrdiv12_fs53_xor1[0]), .d1(arrdiv12_mux2to137_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to149_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to150_out(.d0(arrdiv12_fs54_xor1[0]), .d1(arrdiv12_mux2to138_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to150_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to151_out(.d0(arrdiv12_fs55_xor1[0]), .d1(arrdiv12_mux2to139_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to151_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to152_out(.d0(arrdiv12_fs56_xor1[0]), .d1(arrdiv12_mux2to140_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to152_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to153_out(.d0(arrdiv12_fs57_xor1[0]), .d1(arrdiv12_mux2to141_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to153_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to154_out(.d0(arrdiv12_fs58_xor1[0]), .d1(arrdiv12_mux2to142_xor0[0]), .sel(arrdiv12_fs59_or0[0]), .mux2to1_xor0(arrdiv12_mux2to154_xor0));
  not_gate not_gate_arrdiv12_not4(.a(arrdiv12_fs59_or0[0]), .out(arrdiv12_not4));
  fs fs_arrdiv12_fs60_out(.a(a[6]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs60_xor0), .fs_or0(arrdiv12_fs60_and0));
  fs fs_arrdiv12_fs61_out(.a(arrdiv12_mux2to144_xor0[0]), .b(b[1]), .bin(arrdiv12_fs60_and0[0]), .fs_xor1(arrdiv12_fs61_xor1), .fs_or0(arrdiv12_fs61_or0));
  fs fs_arrdiv12_fs62_out(.a(arrdiv12_mux2to145_xor0[0]), .b(b[2]), .bin(arrdiv12_fs61_or0[0]), .fs_xor1(arrdiv12_fs62_xor1), .fs_or0(arrdiv12_fs62_or0));
  fs fs_arrdiv12_fs63_out(.a(arrdiv12_mux2to146_xor0[0]), .b(b[3]), .bin(arrdiv12_fs62_or0[0]), .fs_xor1(arrdiv12_fs63_xor1), .fs_or0(arrdiv12_fs63_or0));
  fs fs_arrdiv12_fs64_out(.a(arrdiv12_mux2to147_xor0[0]), .b(b[4]), .bin(arrdiv12_fs63_or0[0]), .fs_xor1(arrdiv12_fs64_xor1), .fs_or0(arrdiv12_fs64_or0));
  fs fs_arrdiv12_fs65_out(.a(arrdiv12_mux2to148_xor0[0]), .b(b[5]), .bin(arrdiv12_fs64_or0[0]), .fs_xor1(arrdiv12_fs65_xor1), .fs_or0(arrdiv12_fs65_or0));
  fs fs_arrdiv12_fs66_out(.a(arrdiv12_mux2to149_xor0[0]), .b(b[6]), .bin(arrdiv12_fs65_or0[0]), .fs_xor1(arrdiv12_fs66_xor1), .fs_or0(arrdiv12_fs66_or0));
  fs fs_arrdiv12_fs67_out(.a(arrdiv12_mux2to150_xor0[0]), .b(b[7]), .bin(arrdiv12_fs66_or0[0]), .fs_xor1(arrdiv12_fs67_xor1), .fs_or0(arrdiv12_fs67_or0));
  fs fs_arrdiv12_fs68_out(.a(arrdiv12_mux2to151_xor0[0]), .b(b[8]), .bin(arrdiv12_fs67_or0[0]), .fs_xor1(arrdiv12_fs68_xor1), .fs_or0(arrdiv12_fs68_or0));
  fs fs_arrdiv12_fs69_out(.a(arrdiv12_mux2to152_xor0[0]), .b(b[9]), .bin(arrdiv12_fs68_or0[0]), .fs_xor1(arrdiv12_fs69_xor1), .fs_or0(arrdiv12_fs69_or0));
  fs fs_arrdiv12_fs70_out(.a(arrdiv12_mux2to153_xor0[0]), .b(b[10]), .bin(arrdiv12_fs69_or0[0]), .fs_xor1(arrdiv12_fs70_xor1), .fs_or0(arrdiv12_fs70_or0));
  fs fs_arrdiv12_fs71_out(.a(arrdiv12_mux2to154_xor0[0]), .b(b[11]), .bin(arrdiv12_fs70_or0[0]), .fs_xor1(arrdiv12_fs71_xor1), .fs_or0(arrdiv12_fs71_or0));
  mux2to1 mux2to1_arrdiv12_mux2to155_out(.d0(arrdiv12_fs60_xor0[0]), .d1(a[6]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to155_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to156_out(.d0(arrdiv12_fs61_xor1[0]), .d1(arrdiv12_mux2to144_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to156_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to157_out(.d0(arrdiv12_fs62_xor1[0]), .d1(arrdiv12_mux2to145_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to157_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to158_out(.d0(arrdiv12_fs63_xor1[0]), .d1(arrdiv12_mux2to146_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to158_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to159_out(.d0(arrdiv12_fs64_xor1[0]), .d1(arrdiv12_mux2to147_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to159_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to160_out(.d0(arrdiv12_fs65_xor1[0]), .d1(arrdiv12_mux2to148_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to160_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to161_out(.d0(arrdiv12_fs66_xor1[0]), .d1(arrdiv12_mux2to149_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to161_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to162_out(.d0(arrdiv12_fs67_xor1[0]), .d1(arrdiv12_mux2to150_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to162_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to163_out(.d0(arrdiv12_fs68_xor1[0]), .d1(arrdiv12_mux2to151_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to163_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to164_out(.d0(arrdiv12_fs69_xor1[0]), .d1(arrdiv12_mux2to152_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to164_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to165_out(.d0(arrdiv12_fs70_xor1[0]), .d1(arrdiv12_mux2to153_xor0[0]), .sel(arrdiv12_fs71_or0[0]), .mux2to1_xor0(arrdiv12_mux2to165_xor0));
  not_gate not_gate_arrdiv12_not5(.a(arrdiv12_fs71_or0[0]), .out(arrdiv12_not5));
  fs fs_arrdiv12_fs72_out(.a(a[5]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs72_xor0), .fs_or0(arrdiv12_fs72_and0));
  fs fs_arrdiv12_fs73_out(.a(arrdiv12_mux2to155_xor0[0]), .b(b[1]), .bin(arrdiv12_fs72_and0[0]), .fs_xor1(arrdiv12_fs73_xor1), .fs_or0(arrdiv12_fs73_or0));
  fs fs_arrdiv12_fs74_out(.a(arrdiv12_mux2to156_xor0[0]), .b(b[2]), .bin(arrdiv12_fs73_or0[0]), .fs_xor1(arrdiv12_fs74_xor1), .fs_or0(arrdiv12_fs74_or0));
  fs fs_arrdiv12_fs75_out(.a(arrdiv12_mux2to157_xor0[0]), .b(b[3]), .bin(arrdiv12_fs74_or0[0]), .fs_xor1(arrdiv12_fs75_xor1), .fs_or0(arrdiv12_fs75_or0));
  fs fs_arrdiv12_fs76_out(.a(arrdiv12_mux2to158_xor0[0]), .b(b[4]), .bin(arrdiv12_fs75_or0[0]), .fs_xor1(arrdiv12_fs76_xor1), .fs_or0(arrdiv12_fs76_or0));
  fs fs_arrdiv12_fs77_out(.a(arrdiv12_mux2to159_xor0[0]), .b(b[5]), .bin(arrdiv12_fs76_or0[0]), .fs_xor1(arrdiv12_fs77_xor1), .fs_or0(arrdiv12_fs77_or0));
  fs fs_arrdiv12_fs78_out(.a(arrdiv12_mux2to160_xor0[0]), .b(b[6]), .bin(arrdiv12_fs77_or0[0]), .fs_xor1(arrdiv12_fs78_xor1), .fs_or0(arrdiv12_fs78_or0));
  fs fs_arrdiv12_fs79_out(.a(arrdiv12_mux2to161_xor0[0]), .b(b[7]), .bin(arrdiv12_fs78_or0[0]), .fs_xor1(arrdiv12_fs79_xor1), .fs_or0(arrdiv12_fs79_or0));
  fs fs_arrdiv12_fs80_out(.a(arrdiv12_mux2to162_xor0[0]), .b(b[8]), .bin(arrdiv12_fs79_or0[0]), .fs_xor1(arrdiv12_fs80_xor1), .fs_or0(arrdiv12_fs80_or0));
  fs fs_arrdiv12_fs81_out(.a(arrdiv12_mux2to163_xor0[0]), .b(b[9]), .bin(arrdiv12_fs80_or0[0]), .fs_xor1(arrdiv12_fs81_xor1), .fs_or0(arrdiv12_fs81_or0));
  fs fs_arrdiv12_fs82_out(.a(arrdiv12_mux2to164_xor0[0]), .b(b[10]), .bin(arrdiv12_fs81_or0[0]), .fs_xor1(arrdiv12_fs82_xor1), .fs_or0(arrdiv12_fs82_or0));
  fs fs_arrdiv12_fs83_out(.a(arrdiv12_mux2to165_xor0[0]), .b(b[11]), .bin(arrdiv12_fs82_or0[0]), .fs_xor1(arrdiv12_fs83_xor1), .fs_or0(arrdiv12_fs83_or0));
  mux2to1 mux2to1_arrdiv12_mux2to166_out(.d0(arrdiv12_fs72_xor0[0]), .d1(a[5]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to166_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to167_out(.d0(arrdiv12_fs73_xor1[0]), .d1(arrdiv12_mux2to155_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to167_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to168_out(.d0(arrdiv12_fs74_xor1[0]), .d1(arrdiv12_mux2to156_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to168_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to169_out(.d0(arrdiv12_fs75_xor1[0]), .d1(arrdiv12_mux2to157_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to169_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to170_out(.d0(arrdiv12_fs76_xor1[0]), .d1(arrdiv12_mux2to158_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to170_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to171_out(.d0(arrdiv12_fs77_xor1[0]), .d1(arrdiv12_mux2to159_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to171_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to172_out(.d0(arrdiv12_fs78_xor1[0]), .d1(arrdiv12_mux2to160_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to172_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to173_out(.d0(arrdiv12_fs79_xor1[0]), .d1(arrdiv12_mux2to161_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to173_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to174_out(.d0(arrdiv12_fs80_xor1[0]), .d1(arrdiv12_mux2to162_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to174_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to175_out(.d0(arrdiv12_fs81_xor1[0]), .d1(arrdiv12_mux2to163_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to175_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to176_out(.d0(arrdiv12_fs82_xor1[0]), .d1(arrdiv12_mux2to164_xor0[0]), .sel(arrdiv12_fs83_or0[0]), .mux2to1_xor0(arrdiv12_mux2to176_xor0));
  not_gate not_gate_arrdiv12_not6(.a(arrdiv12_fs83_or0[0]), .out(arrdiv12_not6));
  fs fs_arrdiv12_fs84_out(.a(a[4]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs84_xor0), .fs_or0(arrdiv12_fs84_and0));
  fs fs_arrdiv12_fs85_out(.a(arrdiv12_mux2to166_xor0[0]), .b(b[1]), .bin(arrdiv12_fs84_and0[0]), .fs_xor1(arrdiv12_fs85_xor1), .fs_or0(arrdiv12_fs85_or0));
  fs fs_arrdiv12_fs86_out(.a(arrdiv12_mux2to167_xor0[0]), .b(b[2]), .bin(arrdiv12_fs85_or0[0]), .fs_xor1(arrdiv12_fs86_xor1), .fs_or0(arrdiv12_fs86_or0));
  fs fs_arrdiv12_fs87_out(.a(arrdiv12_mux2to168_xor0[0]), .b(b[3]), .bin(arrdiv12_fs86_or0[0]), .fs_xor1(arrdiv12_fs87_xor1), .fs_or0(arrdiv12_fs87_or0));
  fs fs_arrdiv12_fs88_out(.a(arrdiv12_mux2to169_xor0[0]), .b(b[4]), .bin(arrdiv12_fs87_or0[0]), .fs_xor1(arrdiv12_fs88_xor1), .fs_or0(arrdiv12_fs88_or0));
  fs fs_arrdiv12_fs89_out(.a(arrdiv12_mux2to170_xor0[0]), .b(b[5]), .bin(arrdiv12_fs88_or0[0]), .fs_xor1(arrdiv12_fs89_xor1), .fs_or0(arrdiv12_fs89_or0));
  fs fs_arrdiv12_fs90_out(.a(arrdiv12_mux2to171_xor0[0]), .b(b[6]), .bin(arrdiv12_fs89_or0[0]), .fs_xor1(arrdiv12_fs90_xor1), .fs_or0(arrdiv12_fs90_or0));
  fs fs_arrdiv12_fs91_out(.a(arrdiv12_mux2to172_xor0[0]), .b(b[7]), .bin(arrdiv12_fs90_or0[0]), .fs_xor1(arrdiv12_fs91_xor1), .fs_or0(arrdiv12_fs91_or0));
  fs fs_arrdiv12_fs92_out(.a(arrdiv12_mux2to173_xor0[0]), .b(b[8]), .bin(arrdiv12_fs91_or0[0]), .fs_xor1(arrdiv12_fs92_xor1), .fs_or0(arrdiv12_fs92_or0));
  fs fs_arrdiv12_fs93_out(.a(arrdiv12_mux2to174_xor0[0]), .b(b[9]), .bin(arrdiv12_fs92_or0[0]), .fs_xor1(arrdiv12_fs93_xor1), .fs_or0(arrdiv12_fs93_or0));
  fs fs_arrdiv12_fs94_out(.a(arrdiv12_mux2to175_xor0[0]), .b(b[10]), .bin(arrdiv12_fs93_or0[0]), .fs_xor1(arrdiv12_fs94_xor1), .fs_or0(arrdiv12_fs94_or0));
  fs fs_arrdiv12_fs95_out(.a(arrdiv12_mux2to176_xor0[0]), .b(b[11]), .bin(arrdiv12_fs94_or0[0]), .fs_xor1(arrdiv12_fs95_xor1), .fs_or0(arrdiv12_fs95_or0));
  mux2to1 mux2to1_arrdiv12_mux2to177_out(.d0(arrdiv12_fs84_xor0[0]), .d1(a[4]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to177_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to178_out(.d0(arrdiv12_fs85_xor1[0]), .d1(arrdiv12_mux2to166_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to178_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to179_out(.d0(arrdiv12_fs86_xor1[0]), .d1(arrdiv12_mux2to167_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to179_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to180_out(.d0(arrdiv12_fs87_xor1[0]), .d1(arrdiv12_mux2to168_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to180_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to181_out(.d0(arrdiv12_fs88_xor1[0]), .d1(arrdiv12_mux2to169_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to181_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to182_out(.d0(arrdiv12_fs89_xor1[0]), .d1(arrdiv12_mux2to170_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to182_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to183_out(.d0(arrdiv12_fs90_xor1[0]), .d1(arrdiv12_mux2to171_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to183_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to184_out(.d0(arrdiv12_fs91_xor1[0]), .d1(arrdiv12_mux2to172_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to184_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to185_out(.d0(arrdiv12_fs92_xor1[0]), .d1(arrdiv12_mux2to173_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to185_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to186_out(.d0(arrdiv12_fs93_xor1[0]), .d1(arrdiv12_mux2to174_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to186_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to187_out(.d0(arrdiv12_fs94_xor1[0]), .d1(arrdiv12_mux2to175_xor0[0]), .sel(arrdiv12_fs95_or0[0]), .mux2to1_xor0(arrdiv12_mux2to187_xor0));
  not_gate not_gate_arrdiv12_not7(.a(arrdiv12_fs95_or0[0]), .out(arrdiv12_not7));
  fs fs_arrdiv12_fs96_out(.a(a[3]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs96_xor0), .fs_or0(arrdiv12_fs96_and0));
  fs fs_arrdiv12_fs97_out(.a(arrdiv12_mux2to177_xor0[0]), .b(b[1]), .bin(arrdiv12_fs96_and0[0]), .fs_xor1(arrdiv12_fs97_xor1), .fs_or0(arrdiv12_fs97_or0));
  fs fs_arrdiv12_fs98_out(.a(arrdiv12_mux2to178_xor0[0]), .b(b[2]), .bin(arrdiv12_fs97_or0[0]), .fs_xor1(arrdiv12_fs98_xor1), .fs_or0(arrdiv12_fs98_or0));
  fs fs_arrdiv12_fs99_out(.a(arrdiv12_mux2to179_xor0[0]), .b(b[3]), .bin(arrdiv12_fs98_or0[0]), .fs_xor1(arrdiv12_fs99_xor1), .fs_or0(arrdiv12_fs99_or0));
  fs fs_arrdiv12_fs100_out(.a(arrdiv12_mux2to180_xor0[0]), .b(b[4]), .bin(arrdiv12_fs99_or0[0]), .fs_xor1(arrdiv12_fs100_xor1), .fs_or0(arrdiv12_fs100_or0));
  fs fs_arrdiv12_fs101_out(.a(arrdiv12_mux2to181_xor0[0]), .b(b[5]), .bin(arrdiv12_fs100_or0[0]), .fs_xor1(arrdiv12_fs101_xor1), .fs_or0(arrdiv12_fs101_or0));
  fs fs_arrdiv12_fs102_out(.a(arrdiv12_mux2to182_xor0[0]), .b(b[6]), .bin(arrdiv12_fs101_or0[0]), .fs_xor1(arrdiv12_fs102_xor1), .fs_or0(arrdiv12_fs102_or0));
  fs fs_arrdiv12_fs103_out(.a(arrdiv12_mux2to183_xor0[0]), .b(b[7]), .bin(arrdiv12_fs102_or0[0]), .fs_xor1(arrdiv12_fs103_xor1), .fs_or0(arrdiv12_fs103_or0));
  fs fs_arrdiv12_fs104_out(.a(arrdiv12_mux2to184_xor0[0]), .b(b[8]), .bin(arrdiv12_fs103_or0[0]), .fs_xor1(arrdiv12_fs104_xor1), .fs_or0(arrdiv12_fs104_or0));
  fs fs_arrdiv12_fs105_out(.a(arrdiv12_mux2to185_xor0[0]), .b(b[9]), .bin(arrdiv12_fs104_or0[0]), .fs_xor1(arrdiv12_fs105_xor1), .fs_or0(arrdiv12_fs105_or0));
  fs fs_arrdiv12_fs106_out(.a(arrdiv12_mux2to186_xor0[0]), .b(b[10]), .bin(arrdiv12_fs105_or0[0]), .fs_xor1(arrdiv12_fs106_xor1), .fs_or0(arrdiv12_fs106_or0));
  fs fs_arrdiv12_fs107_out(.a(arrdiv12_mux2to187_xor0[0]), .b(b[11]), .bin(arrdiv12_fs106_or0[0]), .fs_xor1(arrdiv12_fs107_xor1), .fs_or0(arrdiv12_fs107_or0));
  mux2to1 mux2to1_arrdiv12_mux2to188_out(.d0(arrdiv12_fs96_xor0[0]), .d1(a[3]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to188_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to189_out(.d0(arrdiv12_fs97_xor1[0]), .d1(arrdiv12_mux2to177_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to189_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to190_out(.d0(arrdiv12_fs98_xor1[0]), .d1(arrdiv12_mux2to178_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to190_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to191_out(.d0(arrdiv12_fs99_xor1[0]), .d1(arrdiv12_mux2to179_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to191_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to192_out(.d0(arrdiv12_fs100_xor1[0]), .d1(arrdiv12_mux2to180_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to192_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to193_out(.d0(arrdiv12_fs101_xor1[0]), .d1(arrdiv12_mux2to181_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to193_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to194_out(.d0(arrdiv12_fs102_xor1[0]), .d1(arrdiv12_mux2to182_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to194_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to195_out(.d0(arrdiv12_fs103_xor1[0]), .d1(arrdiv12_mux2to183_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to195_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to196_out(.d0(arrdiv12_fs104_xor1[0]), .d1(arrdiv12_mux2to184_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to196_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to197_out(.d0(arrdiv12_fs105_xor1[0]), .d1(arrdiv12_mux2to185_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to197_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to198_out(.d0(arrdiv12_fs106_xor1[0]), .d1(arrdiv12_mux2to186_xor0[0]), .sel(arrdiv12_fs107_or0[0]), .mux2to1_xor0(arrdiv12_mux2to198_xor0));
  not_gate not_gate_arrdiv12_not8(.a(arrdiv12_fs107_or0[0]), .out(arrdiv12_not8));
  fs fs_arrdiv12_fs108_out(.a(a[2]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs108_xor0), .fs_or0(arrdiv12_fs108_and0));
  fs fs_arrdiv12_fs109_out(.a(arrdiv12_mux2to188_xor0[0]), .b(b[1]), .bin(arrdiv12_fs108_and0[0]), .fs_xor1(arrdiv12_fs109_xor1), .fs_or0(arrdiv12_fs109_or0));
  fs fs_arrdiv12_fs110_out(.a(arrdiv12_mux2to189_xor0[0]), .b(b[2]), .bin(arrdiv12_fs109_or0[0]), .fs_xor1(arrdiv12_fs110_xor1), .fs_or0(arrdiv12_fs110_or0));
  fs fs_arrdiv12_fs111_out(.a(arrdiv12_mux2to190_xor0[0]), .b(b[3]), .bin(arrdiv12_fs110_or0[0]), .fs_xor1(arrdiv12_fs111_xor1), .fs_or0(arrdiv12_fs111_or0));
  fs fs_arrdiv12_fs112_out(.a(arrdiv12_mux2to191_xor0[0]), .b(b[4]), .bin(arrdiv12_fs111_or0[0]), .fs_xor1(arrdiv12_fs112_xor1), .fs_or0(arrdiv12_fs112_or0));
  fs fs_arrdiv12_fs113_out(.a(arrdiv12_mux2to192_xor0[0]), .b(b[5]), .bin(arrdiv12_fs112_or0[0]), .fs_xor1(arrdiv12_fs113_xor1), .fs_or0(arrdiv12_fs113_or0));
  fs fs_arrdiv12_fs114_out(.a(arrdiv12_mux2to193_xor0[0]), .b(b[6]), .bin(arrdiv12_fs113_or0[0]), .fs_xor1(arrdiv12_fs114_xor1), .fs_or0(arrdiv12_fs114_or0));
  fs fs_arrdiv12_fs115_out(.a(arrdiv12_mux2to194_xor0[0]), .b(b[7]), .bin(arrdiv12_fs114_or0[0]), .fs_xor1(arrdiv12_fs115_xor1), .fs_or0(arrdiv12_fs115_or0));
  fs fs_arrdiv12_fs116_out(.a(arrdiv12_mux2to195_xor0[0]), .b(b[8]), .bin(arrdiv12_fs115_or0[0]), .fs_xor1(arrdiv12_fs116_xor1), .fs_or0(arrdiv12_fs116_or0));
  fs fs_arrdiv12_fs117_out(.a(arrdiv12_mux2to196_xor0[0]), .b(b[9]), .bin(arrdiv12_fs116_or0[0]), .fs_xor1(arrdiv12_fs117_xor1), .fs_or0(arrdiv12_fs117_or0));
  fs fs_arrdiv12_fs118_out(.a(arrdiv12_mux2to197_xor0[0]), .b(b[10]), .bin(arrdiv12_fs117_or0[0]), .fs_xor1(arrdiv12_fs118_xor1), .fs_or0(arrdiv12_fs118_or0));
  fs fs_arrdiv12_fs119_out(.a(arrdiv12_mux2to198_xor0[0]), .b(b[11]), .bin(arrdiv12_fs118_or0[0]), .fs_xor1(arrdiv12_fs119_xor1), .fs_or0(arrdiv12_fs119_or0));
  mux2to1 mux2to1_arrdiv12_mux2to199_out(.d0(arrdiv12_fs108_xor0[0]), .d1(a[2]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to199_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1100_out(.d0(arrdiv12_fs109_xor1[0]), .d1(arrdiv12_mux2to188_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1100_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1101_out(.d0(arrdiv12_fs110_xor1[0]), .d1(arrdiv12_mux2to189_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1101_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1102_out(.d0(arrdiv12_fs111_xor1[0]), .d1(arrdiv12_mux2to190_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1102_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1103_out(.d0(arrdiv12_fs112_xor1[0]), .d1(arrdiv12_mux2to191_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1103_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1104_out(.d0(arrdiv12_fs113_xor1[0]), .d1(arrdiv12_mux2to192_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1104_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1105_out(.d0(arrdiv12_fs114_xor1[0]), .d1(arrdiv12_mux2to193_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1105_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1106_out(.d0(arrdiv12_fs115_xor1[0]), .d1(arrdiv12_mux2to194_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1106_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1107_out(.d0(arrdiv12_fs116_xor1[0]), .d1(arrdiv12_mux2to195_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1107_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1108_out(.d0(arrdiv12_fs117_xor1[0]), .d1(arrdiv12_mux2to196_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1108_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1109_out(.d0(arrdiv12_fs118_xor1[0]), .d1(arrdiv12_mux2to197_xor0[0]), .sel(arrdiv12_fs119_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1109_xor0));
  not_gate not_gate_arrdiv12_not9(.a(arrdiv12_fs119_or0[0]), .out(arrdiv12_not9));
  fs fs_arrdiv12_fs120_out(.a(a[1]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs120_xor0), .fs_or0(arrdiv12_fs120_and0));
  fs fs_arrdiv12_fs121_out(.a(arrdiv12_mux2to199_xor0[0]), .b(b[1]), .bin(arrdiv12_fs120_and0[0]), .fs_xor1(arrdiv12_fs121_xor1), .fs_or0(arrdiv12_fs121_or0));
  fs fs_arrdiv12_fs122_out(.a(arrdiv12_mux2to1100_xor0[0]), .b(b[2]), .bin(arrdiv12_fs121_or0[0]), .fs_xor1(arrdiv12_fs122_xor1), .fs_or0(arrdiv12_fs122_or0));
  fs fs_arrdiv12_fs123_out(.a(arrdiv12_mux2to1101_xor0[0]), .b(b[3]), .bin(arrdiv12_fs122_or0[0]), .fs_xor1(arrdiv12_fs123_xor1), .fs_or0(arrdiv12_fs123_or0));
  fs fs_arrdiv12_fs124_out(.a(arrdiv12_mux2to1102_xor0[0]), .b(b[4]), .bin(arrdiv12_fs123_or0[0]), .fs_xor1(arrdiv12_fs124_xor1), .fs_or0(arrdiv12_fs124_or0));
  fs fs_arrdiv12_fs125_out(.a(arrdiv12_mux2to1103_xor0[0]), .b(b[5]), .bin(arrdiv12_fs124_or0[0]), .fs_xor1(arrdiv12_fs125_xor1), .fs_or0(arrdiv12_fs125_or0));
  fs fs_arrdiv12_fs126_out(.a(arrdiv12_mux2to1104_xor0[0]), .b(b[6]), .bin(arrdiv12_fs125_or0[0]), .fs_xor1(arrdiv12_fs126_xor1), .fs_or0(arrdiv12_fs126_or0));
  fs fs_arrdiv12_fs127_out(.a(arrdiv12_mux2to1105_xor0[0]), .b(b[7]), .bin(arrdiv12_fs126_or0[0]), .fs_xor1(arrdiv12_fs127_xor1), .fs_or0(arrdiv12_fs127_or0));
  fs fs_arrdiv12_fs128_out(.a(arrdiv12_mux2to1106_xor0[0]), .b(b[8]), .bin(arrdiv12_fs127_or0[0]), .fs_xor1(arrdiv12_fs128_xor1), .fs_or0(arrdiv12_fs128_or0));
  fs fs_arrdiv12_fs129_out(.a(arrdiv12_mux2to1107_xor0[0]), .b(b[9]), .bin(arrdiv12_fs128_or0[0]), .fs_xor1(arrdiv12_fs129_xor1), .fs_or0(arrdiv12_fs129_or0));
  fs fs_arrdiv12_fs130_out(.a(arrdiv12_mux2to1108_xor0[0]), .b(b[10]), .bin(arrdiv12_fs129_or0[0]), .fs_xor1(arrdiv12_fs130_xor1), .fs_or0(arrdiv12_fs130_or0));
  fs fs_arrdiv12_fs131_out(.a(arrdiv12_mux2to1109_xor0[0]), .b(b[11]), .bin(arrdiv12_fs130_or0[0]), .fs_xor1(arrdiv12_fs131_xor1), .fs_or0(arrdiv12_fs131_or0));
  mux2to1 mux2to1_arrdiv12_mux2to1110_out(.d0(arrdiv12_fs120_xor0[0]), .d1(a[1]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1110_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1111_out(.d0(arrdiv12_fs121_xor1[0]), .d1(arrdiv12_mux2to199_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1111_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1112_out(.d0(arrdiv12_fs122_xor1[0]), .d1(arrdiv12_mux2to1100_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1112_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1113_out(.d0(arrdiv12_fs123_xor1[0]), .d1(arrdiv12_mux2to1101_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1113_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1114_out(.d0(arrdiv12_fs124_xor1[0]), .d1(arrdiv12_mux2to1102_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1114_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1115_out(.d0(arrdiv12_fs125_xor1[0]), .d1(arrdiv12_mux2to1103_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1115_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1116_out(.d0(arrdiv12_fs126_xor1[0]), .d1(arrdiv12_mux2to1104_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1116_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1117_out(.d0(arrdiv12_fs127_xor1[0]), .d1(arrdiv12_mux2to1105_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1117_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1118_out(.d0(arrdiv12_fs128_xor1[0]), .d1(arrdiv12_mux2to1106_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1118_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1119_out(.d0(arrdiv12_fs129_xor1[0]), .d1(arrdiv12_mux2to1107_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1119_xor0));
  mux2to1 mux2to1_arrdiv12_mux2to1120_out(.d0(arrdiv12_fs130_xor1[0]), .d1(arrdiv12_mux2to1108_xor0[0]), .sel(arrdiv12_fs131_or0[0]), .mux2to1_xor0(arrdiv12_mux2to1120_xor0));
  not_gate not_gate_arrdiv12_not10(.a(arrdiv12_fs131_or0[0]), .out(arrdiv12_not10));
  fs fs_arrdiv12_fs132_out(.a(a[0]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv12_fs132_xor0), .fs_or0(arrdiv12_fs132_and0));
  fs fs_arrdiv12_fs133_out(.a(arrdiv12_mux2to1110_xor0[0]), .b(b[1]), .bin(arrdiv12_fs132_and0[0]), .fs_xor1(arrdiv12_fs133_xor1), .fs_or0(arrdiv12_fs133_or0));
  fs fs_arrdiv12_fs134_out(.a(arrdiv12_mux2to1111_xor0[0]), .b(b[2]), .bin(arrdiv12_fs133_or0[0]), .fs_xor1(arrdiv12_fs134_xor1), .fs_or0(arrdiv12_fs134_or0));
  fs fs_arrdiv12_fs135_out(.a(arrdiv12_mux2to1112_xor0[0]), .b(b[3]), .bin(arrdiv12_fs134_or0[0]), .fs_xor1(arrdiv12_fs135_xor1), .fs_or0(arrdiv12_fs135_or0));
  fs fs_arrdiv12_fs136_out(.a(arrdiv12_mux2to1113_xor0[0]), .b(b[4]), .bin(arrdiv12_fs135_or0[0]), .fs_xor1(arrdiv12_fs136_xor1), .fs_or0(arrdiv12_fs136_or0));
  fs fs_arrdiv12_fs137_out(.a(arrdiv12_mux2to1114_xor0[0]), .b(b[5]), .bin(arrdiv12_fs136_or0[0]), .fs_xor1(arrdiv12_fs137_xor1), .fs_or0(arrdiv12_fs137_or0));
  fs fs_arrdiv12_fs138_out(.a(arrdiv12_mux2to1115_xor0[0]), .b(b[6]), .bin(arrdiv12_fs137_or0[0]), .fs_xor1(arrdiv12_fs138_xor1), .fs_or0(arrdiv12_fs138_or0));
  fs fs_arrdiv12_fs139_out(.a(arrdiv12_mux2to1116_xor0[0]), .b(b[7]), .bin(arrdiv12_fs138_or0[0]), .fs_xor1(arrdiv12_fs139_xor1), .fs_or0(arrdiv12_fs139_or0));
  fs fs_arrdiv12_fs140_out(.a(arrdiv12_mux2to1117_xor0[0]), .b(b[8]), .bin(arrdiv12_fs139_or0[0]), .fs_xor1(arrdiv12_fs140_xor1), .fs_or0(arrdiv12_fs140_or0));
  fs fs_arrdiv12_fs141_out(.a(arrdiv12_mux2to1118_xor0[0]), .b(b[9]), .bin(arrdiv12_fs140_or0[0]), .fs_xor1(arrdiv12_fs141_xor1), .fs_or0(arrdiv12_fs141_or0));
  fs fs_arrdiv12_fs142_out(.a(arrdiv12_mux2to1119_xor0[0]), .b(b[10]), .bin(arrdiv12_fs141_or0[0]), .fs_xor1(arrdiv12_fs142_xor1), .fs_or0(arrdiv12_fs142_or0));
  fs fs_arrdiv12_fs143_out(.a(arrdiv12_mux2to1120_xor0[0]), .b(b[11]), .bin(arrdiv12_fs142_or0[0]), .fs_xor1(arrdiv12_fs143_xor1), .fs_or0(arrdiv12_fs143_or0));
  not_gate not_gate_arrdiv12_not11(.a(arrdiv12_fs143_or0[0]), .out(arrdiv12_not11));

  assign arrdiv12_out[0] = arrdiv12_not11[0];
  assign arrdiv12_out[1] = arrdiv12_not10[0];
  assign arrdiv12_out[2] = arrdiv12_not9[0];
  assign arrdiv12_out[3] = arrdiv12_not8[0];
  assign arrdiv12_out[4] = arrdiv12_not7[0];
  assign arrdiv12_out[5] = arrdiv12_not6[0];
  assign arrdiv12_out[6] = arrdiv12_not5[0];
  assign arrdiv12_out[7] = arrdiv12_not4[0];
  assign arrdiv12_out[8] = arrdiv12_not3[0];
  assign arrdiv12_out[9] = arrdiv12_not2[0];
  assign arrdiv12_out[10] = arrdiv12_not1[0];
  assign arrdiv12_out[11] = arrdiv12_not0[0];
endmodule