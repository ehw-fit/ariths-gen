module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(.a(a[0]), .b(b[0]), .out(pg_logic_or0));
  and_gate and_gate_pg_logic_and0(.a(a[0]), .b(b[0]), .out(pg_logic_and0));
  xor_gate xor_gate_pg_logic_xor0(.a(a[0]), .b(b[0]), .out(pg_logic_xor0));
endmodule

module u_cla14(input [13:0] a, input [13:0] b, output [14:0] u_cla14_out);
  wire [0:0] u_cla14_pg_logic0_or0;
  wire [0:0] u_cla14_pg_logic0_and0;
  wire [0:0] u_cla14_pg_logic0_xor0;
  wire [0:0] u_cla14_pg_logic1_or0;
  wire [0:0] u_cla14_pg_logic1_and0;
  wire [0:0] u_cla14_pg_logic1_xor0;
  wire [0:0] u_cla14_xor1;
  wire [0:0] u_cla14_and0;
  wire [0:0] u_cla14_or0;
  wire [0:0] u_cla14_pg_logic2_or0;
  wire [0:0] u_cla14_pg_logic2_and0;
  wire [0:0] u_cla14_pg_logic2_xor0;
  wire [0:0] u_cla14_xor2;
  wire [0:0] u_cla14_and1;
  wire [0:0] u_cla14_and2;
  wire [0:0] u_cla14_and3;
  wire [0:0] u_cla14_and4;
  wire [0:0] u_cla14_or1;
  wire [0:0] u_cla14_or2;
  wire [0:0] u_cla14_pg_logic3_or0;
  wire [0:0] u_cla14_pg_logic3_and0;
  wire [0:0] u_cla14_pg_logic3_xor0;
  wire [0:0] u_cla14_xor3;
  wire [0:0] u_cla14_and5;
  wire [0:0] u_cla14_and6;
  wire [0:0] u_cla14_and7;
  wire [0:0] u_cla14_and8;
  wire [0:0] u_cla14_and9;
  wire [0:0] u_cla14_and10;
  wire [0:0] u_cla14_and11;
  wire [0:0] u_cla14_or3;
  wire [0:0] u_cla14_or4;
  wire [0:0] u_cla14_or5;
  wire [0:0] u_cla14_pg_logic4_or0;
  wire [0:0] u_cla14_pg_logic4_and0;
  wire [0:0] u_cla14_pg_logic4_xor0;
  wire [0:0] u_cla14_xor4;
  wire [0:0] u_cla14_and12;
  wire [0:0] u_cla14_or6;
  wire [0:0] u_cla14_pg_logic5_or0;
  wire [0:0] u_cla14_pg_logic5_and0;
  wire [0:0] u_cla14_pg_logic5_xor0;
  wire [0:0] u_cla14_xor5;
  wire [0:0] u_cla14_and13;
  wire [0:0] u_cla14_and14;
  wire [0:0] u_cla14_and15;
  wire [0:0] u_cla14_or7;
  wire [0:0] u_cla14_or8;
  wire [0:0] u_cla14_pg_logic6_or0;
  wire [0:0] u_cla14_pg_logic6_and0;
  wire [0:0] u_cla14_pg_logic6_xor0;
  wire [0:0] u_cla14_xor6;
  wire [0:0] u_cla14_and16;
  wire [0:0] u_cla14_and17;
  wire [0:0] u_cla14_and18;
  wire [0:0] u_cla14_and19;
  wire [0:0] u_cla14_and20;
  wire [0:0] u_cla14_and21;
  wire [0:0] u_cla14_or9;
  wire [0:0] u_cla14_or10;
  wire [0:0] u_cla14_or11;
  wire [0:0] u_cla14_pg_logic7_or0;
  wire [0:0] u_cla14_pg_logic7_and0;
  wire [0:0] u_cla14_pg_logic7_xor0;
  wire [0:0] u_cla14_xor7;
  wire [0:0] u_cla14_and22;
  wire [0:0] u_cla14_and23;
  wire [0:0] u_cla14_and24;
  wire [0:0] u_cla14_and25;
  wire [0:0] u_cla14_and26;
  wire [0:0] u_cla14_and27;
  wire [0:0] u_cla14_and28;
  wire [0:0] u_cla14_and29;
  wire [0:0] u_cla14_and30;
  wire [0:0] u_cla14_and31;
  wire [0:0] u_cla14_or12;
  wire [0:0] u_cla14_or13;
  wire [0:0] u_cla14_or14;
  wire [0:0] u_cla14_or15;
  wire [0:0] u_cla14_pg_logic8_or0;
  wire [0:0] u_cla14_pg_logic8_and0;
  wire [0:0] u_cla14_pg_logic8_xor0;
  wire [0:0] u_cla14_xor8;
  wire [0:0] u_cla14_and32;
  wire [0:0] u_cla14_or16;
  wire [0:0] u_cla14_pg_logic9_or0;
  wire [0:0] u_cla14_pg_logic9_and0;
  wire [0:0] u_cla14_pg_logic9_xor0;
  wire [0:0] u_cla14_xor9;
  wire [0:0] u_cla14_and33;
  wire [0:0] u_cla14_and34;
  wire [0:0] u_cla14_and35;
  wire [0:0] u_cla14_or17;
  wire [0:0] u_cla14_or18;
  wire [0:0] u_cla14_pg_logic10_or0;
  wire [0:0] u_cla14_pg_logic10_and0;
  wire [0:0] u_cla14_pg_logic10_xor0;
  wire [0:0] u_cla14_xor10;
  wire [0:0] u_cla14_and36;
  wire [0:0] u_cla14_and37;
  wire [0:0] u_cla14_and38;
  wire [0:0] u_cla14_and39;
  wire [0:0] u_cla14_and40;
  wire [0:0] u_cla14_and41;
  wire [0:0] u_cla14_or19;
  wire [0:0] u_cla14_or20;
  wire [0:0] u_cla14_or21;
  wire [0:0] u_cla14_pg_logic11_or0;
  wire [0:0] u_cla14_pg_logic11_and0;
  wire [0:0] u_cla14_pg_logic11_xor0;
  wire [0:0] u_cla14_xor11;
  wire [0:0] u_cla14_and42;
  wire [0:0] u_cla14_and43;
  wire [0:0] u_cla14_and44;
  wire [0:0] u_cla14_and45;
  wire [0:0] u_cla14_and46;
  wire [0:0] u_cla14_and47;
  wire [0:0] u_cla14_and48;
  wire [0:0] u_cla14_and49;
  wire [0:0] u_cla14_and50;
  wire [0:0] u_cla14_and51;
  wire [0:0] u_cla14_or22;
  wire [0:0] u_cla14_or23;
  wire [0:0] u_cla14_or24;
  wire [0:0] u_cla14_or25;
  wire [0:0] u_cla14_pg_logic12_or0;
  wire [0:0] u_cla14_pg_logic12_and0;
  wire [0:0] u_cla14_pg_logic12_xor0;
  wire [0:0] u_cla14_xor12;
  wire [0:0] u_cla14_and52;
  wire [0:0] u_cla14_or26;
  wire [0:0] u_cla14_pg_logic13_or0;
  wire [0:0] u_cla14_pg_logic13_and0;
  wire [0:0] u_cla14_pg_logic13_xor0;
  wire [0:0] u_cla14_xor13;
  wire [0:0] u_cla14_and53;
  wire [0:0] u_cla14_and54;
  wire [0:0] u_cla14_and55;
  wire [0:0] u_cla14_or27;
  wire [0:0] u_cla14_or28;

  pg_logic pg_logic_u_cla14_pg_logic0_out(.a(a[0]), .b(b[0]), .pg_logic_or0(u_cla14_pg_logic0_or0), .pg_logic_and0(u_cla14_pg_logic0_and0), .pg_logic_xor0(u_cla14_pg_logic0_xor0));
  pg_logic pg_logic_u_cla14_pg_logic1_out(.a(a[1]), .b(b[1]), .pg_logic_or0(u_cla14_pg_logic1_or0), .pg_logic_and0(u_cla14_pg_logic1_and0), .pg_logic_xor0(u_cla14_pg_logic1_xor0));
  xor_gate xor_gate_u_cla14_xor1(.a(u_cla14_pg_logic1_xor0[0]), .b(u_cla14_pg_logic0_and0[0]), .out(u_cla14_xor1));
  and_gate and_gate_u_cla14_and0(.a(u_cla14_pg_logic0_and0[0]), .b(u_cla14_pg_logic1_or0[0]), .out(u_cla14_and0));
  or_gate or_gate_u_cla14_or0(.a(u_cla14_pg_logic1_and0[0]), .b(u_cla14_and0[0]), .out(u_cla14_or0));
  pg_logic pg_logic_u_cla14_pg_logic2_out(.a(a[2]), .b(b[2]), .pg_logic_or0(u_cla14_pg_logic2_or0), .pg_logic_and0(u_cla14_pg_logic2_and0), .pg_logic_xor0(u_cla14_pg_logic2_xor0));
  xor_gate xor_gate_u_cla14_xor2(.a(u_cla14_pg_logic2_xor0[0]), .b(u_cla14_or0[0]), .out(u_cla14_xor2));
  and_gate and_gate_u_cla14_and1(.a(u_cla14_pg_logic2_or0[0]), .b(u_cla14_pg_logic0_or0[0]), .out(u_cla14_and1));
  and_gate and_gate_u_cla14_and2(.a(u_cla14_pg_logic0_and0[0]), .b(u_cla14_pg_logic2_or0[0]), .out(u_cla14_and2));
  and_gate and_gate_u_cla14_and3(.a(u_cla14_and2[0]), .b(u_cla14_pg_logic1_or0[0]), .out(u_cla14_and3));
  and_gate and_gate_u_cla14_and4(.a(u_cla14_pg_logic1_and0[0]), .b(u_cla14_pg_logic2_or0[0]), .out(u_cla14_and4));
  or_gate or_gate_u_cla14_or1(.a(u_cla14_and3[0]), .b(u_cla14_and4[0]), .out(u_cla14_or1));
  or_gate or_gate_u_cla14_or2(.a(u_cla14_pg_logic2_and0[0]), .b(u_cla14_or1[0]), .out(u_cla14_or2));
  pg_logic pg_logic_u_cla14_pg_logic3_out(.a(a[3]), .b(b[3]), .pg_logic_or0(u_cla14_pg_logic3_or0), .pg_logic_and0(u_cla14_pg_logic3_and0), .pg_logic_xor0(u_cla14_pg_logic3_xor0));
  xor_gate xor_gate_u_cla14_xor3(.a(u_cla14_pg_logic3_xor0[0]), .b(u_cla14_or2[0]), .out(u_cla14_xor3));
  and_gate and_gate_u_cla14_and5(.a(u_cla14_pg_logic3_or0[0]), .b(u_cla14_pg_logic1_or0[0]), .out(u_cla14_and5));
  and_gate and_gate_u_cla14_and6(.a(u_cla14_pg_logic0_and0[0]), .b(u_cla14_pg_logic2_or0[0]), .out(u_cla14_and6));
  and_gate and_gate_u_cla14_and7(.a(u_cla14_pg_logic3_or0[0]), .b(u_cla14_pg_logic1_or0[0]), .out(u_cla14_and7));
  and_gate and_gate_u_cla14_and8(.a(u_cla14_and6[0]), .b(u_cla14_and7[0]), .out(u_cla14_and8));
  and_gate and_gate_u_cla14_and9(.a(u_cla14_pg_logic1_and0[0]), .b(u_cla14_pg_logic3_or0[0]), .out(u_cla14_and9));
  and_gate and_gate_u_cla14_and10(.a(u_cla14_and9[0]), .b(u_cla14_pg_logic2_or0[0]), .out(u_cla14_and10));
  and_gate and_gate_u_cla14_and11(.a(u_cla14_pg_logic2_and0[0]), .b(u_cla14_pg_logic3_or0[0]), .out(u_cla14_and11));
  or_gate or_gate_u_cla14_or3(.a(u_cla14_and8[0]), .b(u_cla14_and11[0]), .out(u_cla14_or3));
  or_gate or_gate_u_cla14_or4(.a(u_cla14_and10[0]), .b(u_cla14_or3[0]), .out(u_cla14_or4));
  or_gate or_gate_u_cla14_or5(.a(u_cla14_pg_logic3_and0[0]), .b(u_cla14_or4[0]), .out(u_cla14_or5));
  pg_logic pg_logic_u_cla14_pg_logic4_out(.a(a[4]), .b(b[4]), .pg_logic_or0(u_cla14_pg_logic4_or0), .pg_logic_and0(u_cla14_pg_logic4_and0), .pg_logic_xor0(u_cla14_pg_logic4_xor0));
  xor_gate xor_gate_u_cla14_xor4(.a(u_cla14_pg_logic4_xor0[0]), .b(u_cla14_or5[0]), .out(u_cla14_xor4));
  and_gate and_gate_u_cla14_and12(.a(u_cla14_or5[0]), .b(u_cla14_pg_logic4_or0[0]), .out(u_cla14_and12));
  or_gate or_gate_u_cla14_or6(.a(u_cla14_pg_logic4_and0[0]), .b(u_cla14_and12[0]), .out(u_cla14_or6));
  pg_logic pg_logic_u_cla14_pg_logic5_out(.a(a[5]), .b(b[5]), .pg_logic_or0(u_cla14_pg_logic5_or0), .pg_logic_and0(u_cla14_pg_logic5_and0), .pg_logic_xor0(u_cla14_pg_logic5_xor0));
  xor_gate xor_gate_u_cla14_xor5(.a(u_cla14_pg_logic5_xor0[0]), .b(u_cla14_or6[0]), .out(u_cla14_xor5));
  and_gate and_gate_u_cla14_and13(.a(u_cla14_or5[0]), .b(u_cla14_pg_logic5_or0[0]), .out(u_cla14_and13));
  and_gate and_gate_u_cla14_and14(.a(u_cla14_and13[0]), .b(u_cla14_pg_logic4_or0[0]), .out(u_cla14_and14));
  and_gate and_gate_u_cla14_and15(.a(u_cla14_pg_logic4_and0[0]), .b(u_cla14_pg_logic5_or0[0]), .out(u_cla14_and15));
  or_gate or_gate_u_cla14_or7(.a(u_cla14_and14[0]), .b(u_cla14_and15[0]), .out(u_cla14_or7));
  or_gate or_gate_u_cla14_or8(.a(u_cla14_pg_logic5_and0[0]), .b(u_cla14_or7[0]), .out(u_cla14_or8));
  pg_logic pg_logic_u_cla14_pg_logic6_out(.a(a[6]), .b(b[6]), .pg_logic_or0(u_cla14_pg_logic6_or0), .pg_logic_and0(u_cla14_pg_logic6_and0), .pg_logic_xor0(u_cla14_pg_logic6_xor0));
  xor_gate xor_gate_u_cla14_xor6(.a(u_cla14_pg_logic6_xor0[0]), .b(u_cla14_or8[0]), .out(u_cla14_xor6));
  and_gate and_gate_u_cla14_and16(.a(u_cla14_or5[0]), .b(u_cla14_pg_logic5_or0[0]), .out(u_cla14_and16));
  and_gate and_gate_u_cla14_and17(.a(u_cla14_pg_logic6_or0[0]), .b(u_cla14_pg_logic4_or0[0]), .out(u_cla14_and17));
  and_gate and_gate_u_cla14_and18(.a(u_cla14_and16[0]), .b(u_cla14_and17[0]), .out(u_cla14_and18));
  and_gate and_gate_u_cla14_and19(.a(u_cla14_pg_logic4_and0[0]), .b(u_cla14_pg_logic6_or0[0]), .out(u_cla14_and19));
  and_gate and_gate_u_cla14_and20(.a(u_cla14_and19[0]), .b(u_cla14_pg_logic5_or0[0]), .out(u_cla14_and20));
  and_gate and_gate_u_cla14_and21(.a(u_cla14_pg_logic5_and0[0]), .b(u_cla14_pg_logic6_or0[0]), .out(u_cla14_and21));
  or_gate or_gate_u_cla14_or9(.a(u_cla14_and18[0]), .b(u_cla14_and20[0]), .out(u_cla14_or9));
  or_gate or_gate_u_cla14_or10(.a(u_cla14_or9[0]), .b(u_cla14_and21[0]), .out(u_cla14_or10));
  or_gate or_gate_u_cla14_or11(.a(u_cla14_pg_logic6_and0[0]), .b(u_cla14_or10[0]), .out(u_cla14_or11));
  pg_logic pg_logic_u_cla14_pg_logic7_out(.a(a[7]), .b(b[7]), .pg_logic_or0(u_cla14_pg_logic7_or0), .pg_logic_and0(u_cla14_pg_logic7_and0), .pg_logic_xor0(u_cla14_pg_logic7_xor0));
  xor_gate xor_gate_u_cla14_xor7(.a(u_cla14_pg_logic7_xor0[0]), .b(u_cla14_or11[0]), .out(u_cla14_xor7));
  and_gate and_gate_u_cla14_and22(.a(u_cla14_or5[0]), .b(u_cla14_pg_logic6_or0[0]), .out(u_cla14_and22));
  and_gate and_gate_u_cla14_and23(.a(u_cla14_pg_logic7_or0[0]), .b(u_cla14_pg_logic5_or0[0]), .out(u_cla14_and23));
  and_gate and_gate_u_cla14_and24(.a(u_cla14_and22[0]), .b(u_cla14_and23[0]), .out(u_cla14_and24));
  and_gate and_gate_u_cla14_and25(.a(u_cla14_and24[0]), .b(u_cla14_pg_logic4_or0[0]), .out(u_cla14_and25));
  and_gate and_gate_u_cla14_and26(.a(u_cla14_pg_logic4_and0[0]), .b(u_cla14_pg_logic6_or0[0]), .out(u_cla14_and26));
  and_gate and_gate_u_cla14_and27(.a(u_cla14_pg_logic7_or0[0]), .b(u_cla14_pg_logic5_or0[0]), .out(u_cla14_and27));
  and_gate and_gate_u_cla14_and28(.a(u_cla14_and26[0]), .b(u_cla14_and27[0]), .out(u_cla14_and28));
  and_gate and_gate_u_cla14_and29(.a(u_cla14_pg_logic5_and0[0]), .b(u_cla14_pg_logic7_or0[0]), .out(u_cla14_and29));
  and_gate and_gate_u_cla14_and30(.a(u_cla14_and29[0]), .b(u_cla14_pg_logic6_or0[0]), .out(u_cla14_and30));
  and_gate and_gate_u_cla14_and31(.a(u_cla14_pg_logic6_and0[0]), .b(u_cla14_pg_logic7_or0[0]), .out(u_cla14_and31));
  or_gate or_gate_u_cla14_or12(.a(u_cla14_and25[0]), .b(u_cla14_and30[0]), .out(u_cla14_or12));
  or_gate or_gate_u_cla14_or13(.a(u_cla14_and28[0]), .b(u_cla14_and31[0]), .out(u_cla14_or13));
  or_gate or_gate_u_cla14_or14(.a(u_cla14_or12[0]), .b(u_cla14_or13[0]), .out(u_cla14_or14));
  or_gate or_gate_u_cla14_or15(.a(u_cla14_pg_logic7_and0[0]), .b(u_cla14_or14[0]), .out(u_cla14_or15));
  pg_logic pg_logic_u_cla14_pg_logic8_out(.a(a[8]), .b(b[8]), .pg_logic_or0(u_cla14_pg_logic8_or0), .pg_logic_and0(u_cla14_pg_logic8_and0), .pg_logic_xor0(u_cla14_pg_logic8_xor0));
  xor_gate xor_gate_u_cla14_xor8(.a(u_cla14_pg_logic8_xor0[0]), .b(u_cla14_or15[0]), .out(u_cla14_xor8));
  and_gate and_gate_u_cla14_and32(.a(u_cla14_or15[0]), .b(u_cla14_pg_logic8_or0[0]), .out(u_cla14_and32));
  or_gate or_gate_u_cla14_or16(.a(u_cla14_pg_logic8_and0[0]), .b(u_cla14_and32[0]), .out(u_cla14_or16));
  pg_logic pg_logic_u_cla14_pg_logic9_out(.a(a[9]), .b(b[9]), .pg_logic_or0(u_cla14_pg_logic9_or0), .pg_logic_and0(u_cla14_pg_logic9_and0), .pg_logic_xor0(u_cla14_pg_logic9_xor0));
  xor_gate xor_gate_u_cla14_xor9(.a(u_cla14_pg_logic9_xor0[0]), .b(u_cla14_or16[0]), .out(u_cla14_xor9));
  and_gate and_gate_u_cla14_and33(.a(u_cla14_or15[0]), .b(u_cla14_pg_logic9_or0[0]), .out(u_cla14_and33));
  and_gate and_gate_u_cla14_and34(.a(u_cla14_and33[0]), .b(u_cla14_pg_logic8_or0[0]), .out(u_cla14_and34));
  and_gate and_gate_u_cla14_and35(.a(u_cla14_pg_logic8_and0[0]), .b(u_cla14_pg_logic9_or0[0]), .out(u_cla14_and35));
  or_gate or_gate_u_cla14_or17(.a(u_cla14_and34[0]), .b(u_cla14_and35[0]), .out(u_cla14_or17));
  or_gate or_gate_u_cla14_or18(.a(u_cla14_pg_logic9_and0[0]), .b(u_cla14_or17[0]), .out(u_cla14_or18));
  pg_logic pg_logic_u_cla14_pg_logic10_out(.a(a[10]), .b(b[10]), .pg_logic_or0(u_cla14_pg_logic10_or0), .pg_logic_and0(u_cla14_pg_logic10_and0), .pg_logic_xor0(u_cla14_pg_logic10_xor0));
  xor_gate xor_gate_u_cla14_xor10(.a(u_cla14_pg_logic10_xor0[0]), .b(u_cla14_or18[0]), .out(u_cla14_xor10));
  and_gate and_gate_u_cla14_and36(.a(u_cla14_or15[0]), .b(u_cla14_pg_logic9_or0[0]), .out(u_cla14_and36));
  and_gate and_gate_u_cla14_and37(.a(u_cla14_pg_logic10_or0[0]), .b(u_cla14_pg_logic8_or0[0]), .out(u_cla14_and37));
  and_gate and_gate_u_cla14_and38(.a(u_cla14_and36[0]), .b(u_cla14_and37[0]), .out(u_cla14_and38));
  and_gate and_gate_u_cla14_and39(.a(u_cla14_pg_logic8_and0[0]), .b(u_cla14_pg_logic10_or0[0]), .out(u_cla14_and39));
  and_gate and_gate_u_cla14_and40(.a(u_cla14_and39[0]), .b(u_cla14_pg_logic9_or0[0]), .out(u_cla14_and40));
  and_gate and_gate_u_cla14_and41(.a(u_cla14_pg_logic9_and0[0]), .b(u_cla14_pg_logic10_or0[0]), .out(u_cla14_and41));
  or_gate or_gate_u_cla14_or19(.a(u_cla14_and38[0]), .b(u_cla14_and40[0]), .out(u_cla14_or19));
  or_gate or_gate_u_cla14_or20(.a(u_cla14_or19[0]), .b(u_cla14_and41[0]), .out(u_cla14_or20));
  or_gate or_gate_u_cla14_or21(.a(u_cla14_pg_logic10_and0[0]), .b(u_cla14_or20[0]), .out(u_cla14_or21));
  pg_logic pg_logic_u_cla14_pg_logic11_out(.a(a[11]), .b(b[11]), .pg_logic_or0(u_cla14_pg_logic11_or0), .pg_logic_and0(u_cla14_pg_logic11_and0), .pg_logic_xor0(u_cla14_pg_logic11_xor0));
  xor_gate xor_gate_u_cla14_xor11(.a(u_cla14_pg_logic11_xor0[0]), .b(u_cla14_or21[0]), .out(u_cla14_xor11));
  and_gate and_gate_u_cla14_and42(.a(u_cla14_or15[0]), .b(u_cla14_pg_logic10_or0[0]), .out(u_cla14_and42));
  and_gate and_gate_u_cla14_and43(.a(u_cla14_pg_logic11_or0[0]), .b(u_cla14_pg_logic9_or0[0]), .out(u_cla14_and43));
  and_gate and_gate_u_cla14_and44(.a(u_cla14_and42[0]), .b(u_cla14_and43[0]), .out(u_cla14_and44));
  and_gate and_gate_u_cla14_and45(.a(u_cla14_and44[0]), .b(u_cla14_pg_logic8_or0[0]), .out(u_cla14_and45));
  and_gate and_gate_u_cla14_and46(.a(u_cla14_pg_logic8_and0[0]), .b(u_cla14_pg_logic10_or0[0]), .out(u_cla14_and46));
  and_gate and_gate_u_cla14_and47(.a(u_cla14_pg_logic11_or0[0]), .b(u_cla14_pg_logic9_or0[0]), .out(u_cla14_and47));
  and_gate and_gate_u_cla14_and48(.a(u_cla14_and46[0]), .b(u_cla14_and47[0]), .out(u_cla14_and48));
  and_gate and_gate_u_cla14_and49(.a(u_cla14_pg_logic9_and0[0]), .b(u_cla14_pg_logic11_or0[0]), .out(u_cla14_and49));
  and_gate and_gate_u_cla14_and50(.a(u_cla14_and49[0]), .b(u_cla14_pg_logic10_or0[0]), .out(u_cla14_and50));
  and_gate and_gate_u_cla14_and51(.a(u_cla14_pg_logic10_and0[0]), .b(u_cla14_pg_logic11_or0[0]), .out(u_cla14_and51));
  or_gate or_gate_u_cla14_or22(.a(u_cla14_and45[0]), .b(u_cla14_and50[0]), .out(u_cla14_or22));
  or_gate or_gate_u_cla14_or23(.a(u_cla14_and48[0]), .b(u_cla14_and51[0]), .out(u_cla14_or23));
  or_gate or_gate_u_cla14_or24(.a(u_cla14_or22[0]), .b(u_cla14_or23[0]), .out(u_cla14_or24));
  or_gate or_gate_u_cla14_or25(.a(u_cla14_pg_logic11_and0[0]), .b(u_cla14_or24[0]), .out(u_cla14_or25));
  pg_logic pg_logic_u_cla14_pg_logic12_out(.a(a[12]), .b(b[12]), .pg_logic_or0(u_cla14_pg_logic12_or0), .pg_logic_and0(u_cla14_pg_logic12_and0), .pg_logic_xor0(u_cla14_pg_logic12_xor0));
  xor_gate xor_gate_u_cla14_xor12(.a(u_cla14_pg_logic12_xor0[0]), .b(u_cla14_or25[0]), .out(u_cla14_xor12));
  and_gate and_gate_u_cla14_and52(.a(u_cla14_or25[0]), .b(u_cla14_pg_logic12_or0[0]), .out(u_cla14_and52));
  or_gate or_gate_u_cla14_or26(.a(u_cla14_pg_logic12_and0[0]), .b(u_cla14_and52[0]), .out(u_cla14_or26));
  pg_logic pg_logic_u_cla14_pg_logic13_out(.a(a[13]), .b(b[13]), .pg_logic_or0(u_cla14_pg_logic13_or0), .pg_logic_and0(u_cla14_pg_logic13_and0), .pg_logic_xor0(u_cla14_pg_logic13_xor0));
  xor_gate xor_gate_u_cla14_xor13(.a(u_cla14_pg_logic13_xor0[0]), .b(u_cla14_or26[0]), .out(u_cla14_xor13));
  and_gate and_gate_u_cla14_and53(.a(u_cla14_or25[0]), .b(u_cla14_pg_logic13_or0[0]), .out(u_cla14_and53));
  and_gate and_gate_u_cla14_and54(.a(u_cla14_and53[0]), .b(u_cla14_pg_logic12_or0[0]), .out(u_cla14_and54));
  and_gate and_gate_u_cla14_and55(.a(u_cla14_pg_logic12_and0[0]), .b(u_cla14_pg_logic13_or0[0]), .out(u_cla14_and55));
  or_gate or_gate_u_cla14_or27(.a(u_cla14_and54[0]), .b(u_cla14_and55[0]), .out(u_cla14_or27));
  or_gate or_gate_u_cla14_or28(.a(u_cla14_pg_logic13_and0[0]), .b(u_cla14_or27[0]), .out(u_cla14_or28));

  assign u_cla14_out[0] = u_cla14_pg_logic0_xor0[0];
  assign u_cla14_out[1] = u_cla14_xor1[0];
  assign u_cla14_out[2] = u_cla14_xor2[0];
  assign u_cla14_out[3] = u_cla14_xor3[0];
  assign u_cla14_out[4] = u_cla14_xor4[0];
  assign u_cla14_out[5] = u_cla14_xor5[0];
  assign u_cla14_out[6] = u_cla14_xor6[0];
  assign u_cla14_out[7] = u_cla14_xor7[0];
  assign u_cla14_out[8] = u_cla14_xor8[0];
  assign u_cla14_out[9] = u_cla14_xor9[0];
  assign u_cla14_out[10] = u_cla14_xor10[0];
  assign u_cla14_out[11] = u_cla14_xor11[0];
  assign u_cla14_out[12] = u_cla14_xor12[0];
  assign u_cla14_out[13] = u_cla14_xor13[0];
  assign u_cla14_out[14] = u_cla14_or28[0];
endmodule

module u_dadda_cla8(input [7:0] a, input [7:0] b, output [15:0] u_dadda_cla8_out);
  wire [0:0] u_dadda_cla8_and_6_0;
  wire [0:0] u_dadda_cla8_and_5_1;
  wire [0:0] u_dadda_cla8_ha0_xor0;
  wire [0:0] u_dadda_cla8_ha0_and0;
  wire [0:0] u_dadda_cla8_and_7_0;
  wire [0:0] u_dadda_cla8_and_6_1;
  wire [0:0] u_dadda_cla8_fa0_xor1;
  wire [0:0] u_dadda_cla8_fa0_or0;
  wire [0:0] u_dadda_cla8_and_5_2;
  wire [0:0] u_dadda_cla8_and_4_3;
  wire [0:0] u_dadda_cla8_ha1_xor0;
  wire [0:0] u_dadda_cla8_ha1_and0;
  wire [0:0] u_dadda_cla8_and_7_1;
  wire [0:0] u_dadda_cla8_fa1_xor1;
  wire [0:0] u_dadda_cla8_fa1_or0;
  wire [0:0] u_dadda_cla8_and_6_2;
  wire [0:0] u_dadda_cla8_and_5_3;
  wire [0:0] u_dadda_cla8_ha2_xor0;
  wire [0:0] u_dadda_cla8_ha2_and0;
  wire [0:0] u_dadda_cla8_and_7_2;
  wire [0:0] u_dadda_cla8_fa2_xor1;
  wire [0:0] u_dadda_cla8_fa2_or0;
  wire [0:0] u_dadda_cla8_and_3_0;
  wire [0:0] u_dadda_cla8_and_2_1;
  wire [0:0] u_dadda_cla8_ha3_xor0;
  wire [0:0] u_dadda_cla8_ha3_and0;
  wire [0:0] u_dadda_cla8_and_4_0;
  wire [0:0] u_dadda_cla8_and_3_1;
  wire [0:0] u_dadda_cla8_fa3_xor1;
  wire [0:0] u_dadda_cla8_fa3_or0;
  wire [0:0] u_dadda_cla8_and_2_2;
  wire [0:0] u_dadda_cla8_and_1_3;
  wire [0:0] u_dadda_cla8_ha4_xor0;
  wire [0:0] u_dadda_cla8_ha4_and0;
  wire [0:0] u_dadda_cla8_and_5_0;
  wire [0:0] u_dadda_cla8_fa4_xor1;
  wire [0:0] u_dadda_cla8_fa4_or0;
  wire [0:0] u_dadda_cla8_and_4_1;
  wire [0:0] u_dadda_cla8_and_3_2;
  wire [0:0] u_dadda_cla8_and_2_3;
  wire [0:0] u_dadda_cla8_fa5_xor1;
  wire [0:0] u_dadda_cla8_fa5_or0;
  wire [0:0] u_dadda_cla8_and_1_4;
  wire [0:0] u_dadda_cla8_and_0_5;
  wire [0:0] u_dadda_cla8_ha5_xor0;
  wire [0:0] u_dadda_cla8_ha5_and0;
  wire [0:0] u_dadda_cla8_fa6_xor1;
  wire [0:0] u_dadda_cla8_fa6_or0;
  wire [0:0] u_dadda_cla8_and_4_2;
  wire [0:0] u_dadda_cla8_and_3_3;
  wire [0:0] u_dadda_cla8_and_2_4;
  wire [0:0] u_dadda_cla8_fa7_xor1;
  wire [0:0] u_dadda_cla8_fa7_or0;
  wire [0:0] u_dadda_cla8_and_1_5;
  wire [0:0] u_dadda_cla8_and_0_6;
  wire [0:0] u_dadda_cla8_fa8_xor1;
  wire [0:0] u_dadda_cla8_fa8_or0;
  wire [0:0] u_dadda_cla8_fa9_xor1;
  wire [0:0] u_dadda_cla8_fa9_or0;
  wire [0:0] u_dadda_cla8_and_3_4;
  wire [0:0] u_dadda_cla8_and_2_5;
  wire [0:0] u_dadda_cla8_and_1_6;
  wire [0:0] u_dadda_cla8_fa10_xor1;
  wire [0:0] u_dadda_cla8_fa10_or0;
  wire [0:0] u_dadda_cla8_and_0_7;
  wire [0:0] u_dadda_cla8_fa11_xor1;
  wire [0:0] u_dadda_cla8_fa11_or0;
  wire [0:0] u_dadda_cla8_fa12_xor1;
  wire [0:0] u_dadda_cla8_fa12_or0;
  wire [0:0] u_dadda_cla8_and_4_4;
  wire [0:0] u_dadda_cla8_and_3_5;
  wire [0:0] u_dadda_cla8_and_2_6;
  wire [0:0] u_dadda_cla8_fa13_xor1;
  wire [0:0] u_dadda_cla8_fa13_or0;
  wire [0:0] u_dadda_cla8_and_1_7;
  wire [0:0] u_dadda_cla8_fa14_xor1;
  wire [0:0] u_dadda_cla8_fa14_or0;
  wire [0:0] u_dadda_cla8_fa15_xor1;
  wire [0:0] u_dadda_cla8_fa15_or0;
  wire [0:0] u_dadda_cla8_and_6_3;
  wire [0:0] u_dadda_cla8_and_5_4;
  wire [0:0] u_dadda_cla8_and_4_5;
  wire [0:0] u_dadda_cla8_fa16_xor1;
  wire [0:0] u_dadda_cla8_fa16_or0;
  wire [0:0] u_dadda_cla8_and_3_6;
  wire [0:0] u_dadda_cla8_and_2_7;
  wire [0:0] u_dadda_cla8_fa17_xor1;
  wire [0:0] u_dadda_cla8_fa17_or0;
  wire [0:0] u_dadda_cla8_fa18_xor1;
  wire [0:0] u_dadda_cla8_fa18_or0;
  wire [0:0] u_dadda_cla8_and_7_3;
  wire [0:0] u_dadda_cla8_and_6_4;
  wire [0:0] u_dadda_cla8_fa19_xor1;
  wire [0:0] u_dadda_cla8_fa19_or0;
  wire [0:0] u_dadda_cla8_and_5_5;
  wire [0:0] u_dadda_cla8_and_4_6;
  wire [0:0] u_dadda_cla8_and_3_7;
  wire [0:0] u_dadda_cla8_fa20_xor1;
  wire [0:0] u_dadda_cla8_fa20_or0;
  wire [0:0] u_dadda_cla8_fa21_xor1;
  wire [0:0] u_dadda_cla8_fa21_or0;
  wire [0:0] u_dadda_cla8_and_7_4;
  wire [0:0] u_dadda_cla8_and_6_5;
  wire [0:0] u_dadda_cla8_and_5_6;
  wire [0:0] u_dadda_cla8_fa22_xor1;
  wire [0:0] u_dadda_cla8_fa22_or0;
  wire [0:0] u_dadda_cla8_and_7_5;
  wire [0:0] u_dadda_cla8_fa23_xor1;
  wire [0:0] u_dadda_cla8_fa23_or0;
  wire [0:0] u_dadda_cla8_and_2_0;
  wire [0:0] u_dadda_cla8_and_1_1;
  wire [0:0] u_dadda_cla8_ha6_xor0;
  wire [0:0] u_dadda_cla8_ha6_and0;
  wire [0:0] u_dadda_cla8_and_1_2;
  wire [0:0] u_dadda_cla8_and_0_3;
  wire [0:0] u_dadda_cla8_fa24_xor1;
  wire [0:0] u_dadda_cla8_fa24_or0;
  wire [0:0] u_dadda_cla8_and_0_4;
  wire [0:0] u_dadda_cla8_fa25_xor1;
  wire [0:0] u_dadda_cla8_fa25_or0;
  wire [0:0] u_dadda_cla8_fa26_xor1;
  wire [0:0] u_dadda_cla8_fa26_or0;
  wire [0:0] u_dadda_cla8_fa27_xor1;
  wire [0:0] u_dadda_cla8_fa27_or0;
  wire [0:0] u_dadda_cla8_fa28_xor1;
  wire [0:0] u_dadda_cla8_fa28_or0;
  wire [0:0] u_dadda_cla8_fa29_xor1;
  wire [0:0] u_dadda_cla8_fa29_or0;
  wire [0:0] u_dadda_cla8_fa30_xor1;
  wire [0:0] u_dadda_cla8_fa30_or0;
  wire [0:0] u_dadda_cla8_fa31_xor1;
  wire [0:0] u_dadda_cla8_fa31_or0;
  wire [0:0] u_dadda_cla8_and_4_7;
  wire [0:0] u_dadda_cla8_fa32_xor1;
  wire [0:0] u_dadda_cla8_fa32_or0;
  wire [0:0] u_dadda_cla8_and_6_6;
  wire [0:0] u_dadda_cla8_and_5_7;
  wire [0:0] u_dadda_cla8_fa33_xor1;
  wire [0:0] u_dadda_cla8_fa33_or0;
  wire [0:0] u_dadda_cla8_and_7_6;
  wire [0:0] u_dadda_cla8_fa34_xor1;
  wire [0:0] u_dadda_cla8_fa34_or0;
  wire [0:0] u_dadda_cla8_and_0_0;
  wire [0:0] u_dadda_cla8_and_1_0;
  wire [0:0] u_dadda_cla8_and_0_2;
  wire [0:0] u_dadda_cla8_and_6_7;
  wire [0:0] u_dadda_cla8_and_0_1;
  wire [0:0] u_dadda_cla8_and_7_7;
  wire [13:0] u_dadda_cla8_u_cla14_a;
  wire [13:0] u_dadda_cla8_u_cla14_b;
  wire [14:0] u_dadda_cla8_u_cla14_out;

  and_gate and_gate_u_dadda_cla8_and_6_0(.a(a[6]), .b(b[0]), .out(u_dadda_cla8_and_6_0));
  and_gate and_gate_u_dadda_cla8_and_5_1(.a(a[5]), .b(b[1]), .out(u_dadda_cla8_and_5_1));
  ha ha_u_dadda_cla8_ha0_out(.a(u_dadda_cla8_and_6_0[0]), .b(u_dadda_cla8_and_5_1[0]), .ha_xor0(u_dadda_cla8_ha0_xor0), .ha_and0(u_dadda_cla8_ha0_and0));
  and_gate and_gate_u_dadda_cla8_and_7_0(.a(a[7]), .b(b[0]), .out(u_dadda_cla8_and_7_0));
  and_gate and_gate_u_dadda_cla8_and_6_1(.a(a[6]), .b(b[1]), .out(u_dadda_cla8_and_6_1));
  fa fa_u_dadda_cla8_fa0_out(.a(u_dadda_cla8_ha0_and0[0]), .b(u_dadda_cla8_and_7_0[0]), .cin(u_dadda_cla8_and_6_1[0]), .fa_xor1(u_dadda_cla8_fa0_xor1), .fa_or0(u_dadda_cla8_fa0_or0));
  and_gate and_gate_u_dadda_cla8_and_5_2(.a(a[5]), .b(b[2]), .out(u_dadda_cla8_and_5_2));
  and_gate and_gate_u_dadda_cla8_and_4_3(.a(a[4]), .b(b[3]), .out(u_dadda_cla8_and_4_3));
  ha ha_u_dadda_cla8_ha1_out(.a(u_dadda_cla8_and_5_2[0]), .b(u_dadda_cla8_and_4_3[0]), .ha_xor0(u_dadda_cla8_ha1_xor0), .ha_and0(u_dadda_cla8_ha1_and0));
  and_gate and_gate_u_dadda_cla8_and_7_1(.a(a[7]), .b(b[1]), .out(u_dadda_cla8_and_7_1));
  fa fa_u_dadda_cla8_fa1_out(.a(u_dadda_cla8_ha1_and0[0]), .b(u_dadda_cla8_fa0_or0[0]), .cin(u_dadda_cla8_and_7_1[0]), .fa_xor1(u_dadda_cla8_fa1_xor1), .fa_or0(u_dadda_cla8_fa1_or0));
  and_gate and_gate_u_dadda_cla8_and_6_2(.a(a[6]), .b(b[2]), .out(u_dadda_cla8_and_6_2));
  and_gate and_gate_u_dadda_cla8_and_5_3(.a(a[5]), .b(b[3]), .out(u_dadda_cla8_and_5_3));
  ha ha_u_dadda_cla8_ha2_out(.a(u_dadda_cla8_and_6_2[0]), .b(u_dadda_cla8_and_5_3[0]), .ha_xor0(u_dadda_cla8_ha2_xor0), .ha_and0(u_dadda_cla8_ha2_and0));
  and_gate and_gate_u_dadda_cla8_and_7_2(.a(a[7]), .b(b[2]), .out(u_dadda_cla8_and_7_2));
  fa fa_u_dadda_cla8_fa2_out(.a(u_dadda_cla8_ha2_and0[0]), .b(u_dadda_cla8_fa1_or0[0]), .cin(u_dadda_cla8_and_7_2[0]), .fa_xor1(u_dadda_cla8_fa2_xor1), .fa_or0(u_dadda_cla8_fa2_or0));
  and_gate and_gate_u_dadda_cla8_and_3_0(.a(a[3]), .b(b[0]), .out(u_dadda_cla8_and_3_0));
  and_gate and_gate_u_dadda_cla8_and_2_1(.a(a[2]), .b(b[1]), .out(u_dadda_cla8_and_2_1));
  ha ha_u_dadda_cla8_ha3_out(.a(u_dadda_cla8_and_3_0[0]), .b(u_dadda_cla8_and_2_1[0]), .ha_xor0(u_dadda_cla8_ha3_xor0), .ha_and0(u_dadda_cla8_ha3_and0));
  and_gate and_gate_u_dadda_cla8_and_4_0(.a(a[4]), .b(b[0]), .out(u_dadda_cla8_and_4_0));
  and_gate and_gate_u_dadda_cla8_and_3_1(.a(a[3]), .b(b[1]), .out(u_dadda_cla8_and_3_1));
  fa fa_u_dadda_cla8_fa3_out(.a(u_dadda_cla8_ha3_and0[0]), .b(u_dadda_cla8_and_4_0[0]), .cin(u_dadda_cla8_and_3_1[0]), .fa_xor1(u_dadda_cla8_fa3_xor1), .fa_or0(u_dadda_cla8_fa3_or0));
  and_gate and_gate_u_dadda_cla8_and_2_2(.a(a[2]), .b(b[2]), .out(u_dadda_cla8_and_2_2));
  and_gate and_gate_u_dadda_cla8_and_1_3(.a(a[1]), .b(b[3]), .out(u_dadda_cla8_and_1_3));
  ha ha_u_dadda_cla8_ha4_out(.a(u_dadda_cla8_and_2_2[0]), .b(u_dadda_cla8_and_1_3[0]), .ha_xor0(u_dadda_cla8_ha4_xor0), .ha_and0(u_dadda_cla8_ha4_and0));
  and_gate and_gate_u_dadda_cla8_and_5_0(.a(a[5]), .b(b[0]), .out(u_dadda_cla8_and_5_0));
  fa fa_u_dadda_cla8_fa4_out(.a(u_dadda_cla8_ha4_and0[0]), .b(u_dadda_cla8_fa3_or0[0]), .cin(u_dadda_cla8_and_5_0[0]), .fa_xor1(u_dadda_cla8_fa4_xor1), .fa_or0(u_dadda_cla8_fa4_or0));
  and_gate and_gate_u_dadda_cla8_and_4_1(.a(a[4]), .b(b[1]), .out(u_dadda_cla8_and_4_1));
  and_gate and_gate_u_dadda_cla8_and_3_2(.a(a[3]), .b(b[2]), .out(u_dadda_cla8_and_3_2));
  and_gate and_gate_u_dadda_cla8_and_2_3(.a(a[2]), .b(b[3]), .out(u_dadda_cla8_and_2_3));
  fa fa_u_dadda_cla8_fa5_out(.a(u_dadda_cla8_and_4_1[0]), .b(u_dadda_cla8_and_3_2[0]), .cin(u_dadda_cla8_and_2_3[0]), .fa_xor1(u_dadda_cla8_fa5_xor1), .fa_or0(u_dadda_cla8_fa5_or0));
  and_gate and_gate_u_dadda_cla8_and_1_4(.a(a[1]), .b(b[4]), .out(u_dadda_cla8_and_1_4));
  and_gate and_gate_u_dadda_cla8_and_0_5(.a(a[0]), .b(b[5]), .out(u_dadda_cla8_and_0_5));
  ha ha_u_dadda_cla8_ha5_out(.a(u_dadda_cla8_and_1_4[0]), .b(u_dadda_cla8_and_0_5[0]), .ha_xor0(u_dadda_cla8_ha5_xor0), .ha_and0(u_dadda_cla8_ha5_and0));
  fa fa_u_dadda_cla8_fa6_out(.a(u_dadda_cla8_ha5_and0[0]), .b(u_dadda_cla8_fa5_or0[0]), .cin(u_dadda_cla8_fa4_or0[0]), .fa_xor1(u_dadda_cla8_fa6_xor1), .fa_or0(u_dadda_cla8_fa6_or0));
  and_gate and_gate_u_dadda_cla8_and_4_2(.a(a[4]), .b(b[2]), .out(u_dadda_cla8_and_4_2));
  and_gate and_gate_u_dadda_cla8_and_3_3(.a(a[3]), .b(b[3]), .out(u_dadda_cla8_and_3_3));
  and_gate and_gate_u_dadda_cla8_and_2_4(.a(a[2]), .b(b[4]), .out(u_dadda_cla8_and_2_4));
  fa fa_u_dadda_cla8_fa7_out(.a(u_dadda_cla8_and_4_2[0]), .b(u_dadda_cla8_and_3_3[0]), .cin(u_dadda_cla8_and_2_4[0]), .fa_xor1(u_dadda_cla8_fa7_xor1), .fa_or0(u_dadda_cla8_fa7_or0));
  and_gate and_gate_u_dadda_cla8_and_1_5(.a(a[1]), .b(b[5]), .out(u_dadda_cla8_and_1_5));
  and_gate and_gate_u_dadda_cla8_and_0_6(.a(a[0]), .b(b[6]), .out(u_dadda_cla8_and_0_6));
  fa fa_u_dadda_cla8_fa8_out(.a(u_dadda_cla8_and_1_5[0]), .b(u_dadda_cla8_and_0_6[0]), .cin(u_dadda_cla8_ha0_xor0[0]), .fa_xor1(u_dadda_cla8_fa8_xor1), .fa_or0(u_dadda_cla8_fa8_or0));
  fa fa_u_dadda_cla8_fa9_out(.a(u_dadda_cla8_fa8_or0[0]), .b(u_dadda_cla8_fa7_or0[0]), .cin(u_dadda_cla8_fa6_or0[0]), .fa_xor1(u_dadda_cla8_fa9_xor1), .fa_or0(u_dadda_cla8_fa9_or0));
  and_gate and_gate_u_dadda_cla8_and_3_4(.a(a[3]), .b(b[4]), .out(u_dadda_cla8_and_3_4));
  and_gate and_gate_u_dadda_cla8_and_2_5(.a(a[2]), .b(b[5]), .out(u_dadda_cla8_and_2_5));
  and_gate and_gate_u_dadda_cla8_and_1_6(.a(a[1]), .b(b[6]), .out(u_dadda_cla8_and_1_6));
  fa fa_u_dadda_cla8_fa10_out(.a(u_dadda_cla8_and_3_4[0]), .b(u_dadda_cla8_and_2_5[0]), .cin(u_dadda_cla8_and_1_6[0]), .fa_xor1(u_dadda_cla8_fa10_xor1), .fa_or0(u_dadda_cla8_fa10_or0));
  and_gate and_gate_u_dadda_cla8_and_0_7(.a(a[0]), .b(b[7]), .out(u_dadda_cla8_and_0_7));
  fa fa_u_dadda_cla8_fa11_out(.a(u_dadda_cla8_and_0_7[0]), .b(u_dadda_cla8_fa0_xor1[0]), .cin(u_dadda_cla8_ha1_xor0[0]), .fa_xor1(u_dadda_cla8_fa11_xor1), .fa_or0(u_dadda_cla8_fa11_or0));
  fa fa_u_dadda_cla8_fa12_out(.a(u_dadda_cla8_fa11_or0[0]), .b(u_dadda_cla8_fa10_or0[0]), .cin(u_dadda_cla8_fa9_or0[0]), .fa_xor1(u_dadda_cla8_fa12_xor1), .fa_or0(u_dadda_cla8_fa12_or0));
  and_gate and_gate_u_dadda_cla8_and_4_4(.a(a[4]), .b(b[4]), .out(u_dadda_cla8_and_4_4));
  and_gate and_gate_u_dadda_cla8_and_3_5(.a(a[3]), .b(b[5]), .out(u_dadda_cla8_and_3_5));
  and_gate and_gate_u_dadda_cla8_and_2_6(.a(a[2]), .b(b[6]), .out(u_dadda_cla8_and_2_6));
  fa fa_u_dadda_cla8_fa13_out(.a(u_dadda_cla8_and_4_4[0]), .b(u_dadda_cla8_and_3_5[0]), .cin(u_dadda_cla8_and_2_6[0]), .fa_xor1(u_dadda_cla8_fa13_xor1), .fa_or0(u_dadda_cla8_fa13_or0));
  and_gate and_gate_u_dadda_cla8_and_1_7(.a(a[1]), .b(b[7]), .out(u_dadda_cla8_and_1_7));
  fa fa_u_dadda_cla8_fa14_out(.a(u_dadda_cla8_and_1_7[0]), .b(u_dadda_cla8_fa1_xor1[0]), .cin(u_dadda_cla8_ha2_xor0[0]), .fa_xor1(u_dadda_cla8_fa14_xor1), .fa_or0(u_dadda_cla8_fa14_or0));
  fa fa_u_dadda_cla8_fa15_out(.a(u_dadda_cla8_fa14_or0[0]), .b(u_dadda_cla8_fa13_or0[0]), .cin(u_dadda_cla8_fa12_or0[0]), .fa_xor1(u_dadda_cla8_fa15_xor1), .fa_or0(u_dadda_cla8_fa15_or0));
  and_gate and_gate_u_dadda_cla8_and_6_3(.a(a[6]), .b(b[3]), .out(u_dadda_cla8_and_6_3));
  and_gate and_gate_u_dadda_cla8_and_5_4(.a(a[5]), .b(b[4]), .out(u_dadda_cla8_and_5_4));
  and_gate and_gate_u_dadda_cla8_and_4_5(.a(a[4]), .b(b[5]), .out(u_dadda_cla8_and_4_5));
  fa fa_u_dadda_cla8_fa16_out(.a(u_dadda_cla8_and_6_3[0]), .b(u_dadda_cla8_and_5_4[0]), .cin(u_dadda_cla8_and_4_5[0]), .fa_xor1(u_dadda_cla8_fa16_xor1), .fa_or0(u_dadda_cla8_fa16_or0));
  and_gate and_gate_u_dadda_cla8_and_3_6(.a(a[3]), .b(b[6]), .out(u_dadda_cla8_and_3_6));
  and_gate and_gate_u_dadda_cla8_and_2_7(.a(a[2]), .b(b[7]), .out(u_dadda_cla8_and_2_7));
  fa fa_u_dadda_cla8_fa17_out(.a(u_dadda_cla8_and_3_6[0]), .b(u_dadda_cla8_and_2_7[0]), .cin(u_dadda_cla8_fa2_xor1[0]), .fa_xor1(u_dadda_cla8_fa17_xor1), .fa_or0(u_dadda_cla8_fa17_or0));
  fa fa_u_dadda_cla8_fa18_out(.a(u_dadda_cla8_fa17_or0[0]), .b(u_dadda_cla8_fa16_or0[0]), .cin(u_dadda_cla8_fa15_or0[0]), .fa_xor1(u_dadda_cla8_fa18_xor1), .fa_or0(u_dadda_cla8_fa18_or0));
  and_gate and_gate_u_dadda_cla8_and_7_3(.a(a[7]), .b(b[3]), .out(u_dadda_cla8_and_7_3));
  and_gate and_gate_u_dadda_cla8_and_6_4(.a(a[6]), .b(b[4]), .out(u_dadda_cla8_and_6_4));
  fa fa_u_dadda_cla8_fa19_out(.a(u_dadda_cla8_fa2_or0[0]), .b(u_dadda_cla8_and_7_3[0]), .cin(u_dadda_cla8_and_6_4[0]), .fa_xor1(u_dadda_cla8_fa19_xor1), .fa_or0(u_dadda_cla8_fa19_or0));
  and_gate and_gate_u_dadda_cla8_and_5_5(.a(a[5]), .b(b[5]), .out(u_dadda_cla8_and_5_5));
  and_gate and_gate_u_dadda_cla8_and_4_6(.a(a[4]), .b(b[6]), .out(u_dadda_cla8_and_4_6));
  and_gate and_gate_u_dadda_cla8_and_3_7(.a(a[3]), .b(b[7]), .out(u_dadda_cla8_and_3_7));
  fa fa_u_dadda_cla8_fa20_out(.a(u_dadda_cla8_and_5_5[0]), .b(u_dadda_cla8_and_4_6[0]), .cin(u_dadda_cla8_and_3_7[0]), .fa_xor1(u_dadda_cla8_fa20_xor1), .fa_or0(u_dadda_cla8_fa20_or0));
  fa fa_u_dadda_cla8_fa21_out(.a(u_dadda_cla8_fa20_or0[0]), .b(u_dadda_cla8_fa19_or0[0]), .cin(u_dadda_cla8_fa18_or0[0]), .fa_xor1(u_dadda_cla8_fa21_xor1), .fa_or0(u_dadda_cla8_fa21_or0));
  and_gate and_gate_u_dadda_cla8_and_7_4(.a(a[7]), .b(b[4]), .out(u_dadda_cla8_and_7_4));
  and_gate and_gate_u_dadda_cla8_and_6_5(.a(a[6]), .b(b[5]), .out(u_dadda_cla8_and_6_5));
  and_gate and_gate_u_dadda_cla8_and_5_6(.a(a[5]), .b(b[6]), .out(u_dadda_cla8_and_5_6));
  fa fa_u_dadda_cla8_fa22_out(.a(u_dadda_cla8_and_7_4[0]), .b(u_dadda_cla8_and_6_5[0]), .cin(u_dadda_cla8_and_5_6[0]), .fa_xor1(u_dadda_cla8_fa22_xor1), .fa_or0(u_dadda_cla8_fa22_or0));
  and_gate and_gate_u_dadda_cla8_and_7_5(.a(a[7]), .b(b[5]), .out(u_dadda_cla8_and_7_5));
  fa fa_u_dadda_cla8_fa23_out(.a(u_dadda_cla8_fa22_or0[0]), .b(u_dadda_cla8_fa21_or0[0]), .cin(u_dadda_cla8_and_7_5[0]), .fa_xor1(u_dadda_cla8_fa23_xor1), .fa_or0(u_dadda_cla8_fa23_or0));
  and_gate and_gate_u_dadda_cla8_and_2_0(.a(a[2]), .b(b[0]), .out(u_dadda_cla8_and_2_0));
  and_gate and_gate_u_dadda_cla8_and_1_1(.a(a[1]), .b(b[1]), .out(u_dadda_cla8_and_1_1));
  ha ha_u_dadda_cla8_ha6_out(.a(u_dadda_cla8_and_2_0[0]), .b(u_dadda_cla8_and_1_1[0]), .ha_xor0(u_dadda_cla8_ha6_xor0), .ha_and0(u_dadda_cla8_ha6_and0));
  and_gate and_gate_u_dadda_cla8_and_1_2(.a(a[1]), .b(b[2]), .out(u_dadda_cla8_and_1_2));
  and_gate and_gate_u_dadda_cla8_and_0_3(.a(a[0]), .b(b[3]), .out(u_dadda_cla8_and_0_3));
  fa fa_u_dadda_cla8_fa24_out(.a(u_dadda_cla8_ha6_and0[0]), .b(u_dadda_cla8_and_1_2[0]), .cin(u_dadda_cla8_and_0_3[0]), .fa_xor1(u_dadda_cla8_fa24_xor1), .fa_or0(u_dadda_cla8_fa24_or0));
  and_gate and_gate_u_dadda_cla8_and_0_4(.a(a[0]), .b(b[4]), .out(u_dadda_cla8_and_0_4));
  fa fa_u_dadda_cla8_fa25_out(.a(u_dadda_cla8_fa24_or0[0]), .b(u_dadda_cla8_and_0_4[0]), .cin(u_dadda_cla8_fa3_xor1[0]), .fa_xor1(u_dadda_cla8_fa25_xor1), .fa_or0(u_dadda_cla8_fa25_or0));
  fa fa_u_dadda_cla8_fa26_out(.a(u_dadda_cla8_fa25_or0[0]), .b(u_dadda_cla8_fa4_xor1[0]), .cin(u_dadda_cla8_fa5_xor1[0]), .fa_xor1(u_dadda_cla8_fa26_xor1), .fa_or0(u_dadda_cla8_fa26_or0));
  fa fa_u_dadda_cla8_fa27_out(.a(u_dadda_cla8_fa26_or0[0]), .b(u_dadda_cla8_fa6_xor1[0]), .cin(u_dadda_cla8_fa7_xor1[0]), .fa_xor1(u_dadda_cla8_fa27_xor1), .fa_or0(u_dadda_cla8_fa27_or0));
  fa fa_u_dadda_cla8_fa28_out(.a(u_dadda_cla8_fa27_or0[0]), .b(u_dadda_cla8_fa9_xor1[0]), .cin(u_dadda_cla8_fa10_xor1[0]), .fa_xor1(u_dadda_cla8_fa28_xor1), .fa_or0(u_dadda_cla8_fa28_or0));
  fa fa_u_dadda_cla8_fa29_out(.a(u_dadda_cla8_fa28_or0[0]), .b(u_dadda_cla8_fa12_xor1[0]), .cin(u_dadda_cla8_fa13_xor1[0]), .fa_xor1(u_dadda_cla8_fa29_xor1), .fa_or0(u_dadda_cla8_fa29_or0));
  fa fa_u_dadda_cla8_fa30_out(.a(u_dadda_cla8_fa29_or0[0]), .b(u_dadda_cla8_fa15_xor1[0]), .cin(u_dadda_cla8_fa16_xor1[0]), .fa_xor1(u_dadda_cla8_fa30_xor1), .fa_or0(u_dadda_cla8_fa30_or0));
  fa fa_u_dadda_cla8_fa31_out(.a(u_dadda_cla8_fa30_or0[0]), .b(u_dadda_cla8_fa18_xor1[0]), .cin(u_dadda_cla8_fa19_xor1[0]), .fa_xor1(u_dadda_cla8_fa31_xor1), .fa_or0(u_dadda_cla8_fa31_or0));
  and_gate and_gate_u_dadda_cla8_and_4_7(.a(a[4]), .b(b[7]), .out(u_dadda_cla8_and_4_7));
  fa fa_u_dadda_cla8_fa32_out(.a(u_dadda_cla8_fa31_or0[0]), .b(u_dadda_cla8_and_4_7[0]), .cin(u_dadda_cla8_fa21_xor1[0]), .fa_xor1(u_dadda_cla8_fa32_xor1), .fa_or0(u_dadda_cla8_fa32_or0));
  and_gate and_gate_u_dadda_cla8_and_6_6(.a(a[6]), .b(b[6]), .out(u_dadda_cla8_and_6_6));
  and_gate and_gate_u_dadda_cla8_and_5_7(.a(a[5]), .b(b[7]), .out(u_dadda_cla8_and_5_7));
  fa fa_u_dadda_cla8_fa33_out(.a(u_dadda_cla8_fa32_or0[0]), .b(u_dadda_cla8_and_6_6[0]), .cin(u_dadda_cla8_and_5_7[0]), .fa_xor1(u_dadda_cla8_fa33_xor1), .fa_or0(u_dadda_cla8_fa33_or0));
  and_gate and_gate_u_dadda_cla8_and_7_6(.a(a[7]), .b(b[6]), .out(u_dadda_cla8_and_7_6));
  fa fa_u_dadda_cla8_fa34_out(.a(u_dadda_cla8_fa33_or0[0]), .b(u_dadda_cla8_fa23_or0[0]), .cin(u_dadda_cla8_and_7_6[0]), .fa_xor1(u_dadda_cla8_fa34_xor1), .fa_or0(u_dadda_cla8_fa34_or0));
  and_gate and_gate_u_dadda_cla8_and_0_0(.a(a[0]), .b(b[0]), .out(u_dadda_cla8_and_0_0));
  and_gate and_gate_u_dadda_cla8_and_1_0(.a(a[1]), .b(b[0]), .out(u_dadda_cla8_and_1_0));
  and_gate and_gate_u_dadda_cla8_and_0_2(.a(a[0]), .b(b[2]), .out(u_dadda_cla8_and_0_2));
  and_gate and_gate_u_dadda_cla8_and_6_7(.a(a[6]), .b(b[7]), .out(u_dadda_cla8_and_6_7));
  and_gate and_gate_u_dadda_cla8_and_0_1(.a(a[0]), .b(b[1]), .out(u_dadda_cla8_and_0_1));
  and_gate and_gate_u_dadda_cla8_and_7_7(.a(a[7]), .b(b[7]), .out(u_dadda_cla8_and_7_7));
  assign u_dadda_cla8_u_cla14_a[0] = u_dadda_cla8_and_1_0[0];
  assign u_dadda_cla8_u_cla14_a[1] = u_dadda_cla8_and_0_2[0];
  assign u_dadda_cla8_u_cla14_a[2] = u_dadda_cla8_ha3_xor0[0];
  assign u_dadda_cla8_u_cla14_a[3] = u_dadda_cla8_ha4_xor0[0];
  assign u_dadda_cla8_u_cla14_a[4] = u_dadda_cla8_ha5_xor0[0];
  assign u_dadda_cla8_u_cla14_a[5] = u_dadda_cla8_fa8_xor1[0];
  assign u_dadda_cla8_u_cla14_a[6] = u_dadda_cla8_fa11_xor1[0];
  assign u_dadda_cla8_u_cla14_a[7] = u_dadda_cla8_fa14_xor1[0];
  assign u_dadda_cla8_u_cla14_a[8] = u_dadda_cla8_fa17_xor1[0];
  assign u_dadda_cla8_u_cla14_a[9] = u_dadda_cla8_fa20_xor1[0];
  assign u_dadda_cla8_u_cla14_a[10] = u_dadda_cla8_fa22_xor1[0];
  assign u_dadda_cla8_u_cla14_a[11] = u_dadda_cla8_fa23_xor1[0];
  assign u_dadda_cla8_u_cla14_a[12] = u_dadda_cla8_and_6_7[0];
  assign u_dadda_cla8_u_cla14_a[13] = u_dadda_cla8_fa34_or0[0];
  assign u_dadda_cla8_u_cla14_b[0] = u_dadda_cla8_and_0_1[0];
  assign u_dadda_cla8_u_cla14_b[1] = u_dadda_cla8_ha6_xor0[0];
  assign u_dadda_cla8_u_cla14_b[2] = u_dadda_cla8_fa24_xor1[0];
  assign u_dadda_cla8_u_cla14_b[3] = u_dadda_cla8_fa25_xor1[0];
  assign u_dadda_cla8_u_cla14_b[4] = u_dadda_cla8_fa26_xor1[0];
  assign u_dadda_cla8_u_cla14_b[5] = u_dadda_cla8_fa27_xor1[0];
  assign u_dadda_cla8_u_cla14_b[6] = u_dadda_cla8_fa28_xor1[0];
  assign u_dadda_cla8_u_cla14_b[7] = u_dadda_cla8_fa29_xor1[0];
  assign u_dadda_cla8_u_cla14_b[8] = u_dadda_cla8_fa30_xor1[0];
  assign u_dadda_cla8_u_cla14_b[9] = u_dadda_cla8_fa31_xor1[0];
  assign u_dadda_cla8_u_cla14_b[10] = u_dadda_cla8_fa32_xor1[0];
  assign u_dadda_cla8_u_cla14_b[11] = u_dadda_cla8_fa33_xor1[0];
  assign u_dadda_cla8_u_cla14_b[12] = u_dadda_cla8_fa34_xor1[0];
  assign u_dadda_cla8_u_cla14_b[13] = u_dadda_cla8_and_7_7[0];
  u_cla14 u_cla14_u_dadda_cla8_u_cla14_out(.a(u_dadda_cla8_u_cla14_a), .b(u_dadda_cla8_u_cla14_b), .u_cla14_out(u_dadda_cla8_u_cla14_out));

  assign u_dadda_cla8_out[0] = u_dadda_cla8_and_0_0[0];
  assign u_dadda_cla8_out[1] = u_dadda_cla8_u_cla14_out[0];
  assign u_dadda_cla8_out[2] = u_dadda_cla8_u_cla14_out[1];
  assign u_dadda_cla8_out[3] = u_dadda_cla8_u_cla14_out[2];
  assign u_dadda_cla8_out[4] = u_dadda_cla8_u_cla14_out[3];
  assign u_dadda_cla8_out[5] = u_dadda_cla8_u_cla14_out[4];
  assign u_dadda_cla8_out[6] = u_dadda_cla8_u_cla14_out[5];
  assign u_dadda_cla8_out[7] = u_dadda_cla8_u_cla14_out[6];
  assign u_dadda_cla8_out[8] = u_dadda_cla8_u_cla14_out[7];
  assign u_dadda_cla8_out[9] = u_dadda_cla8_u_cla14_out[8];
  assign u_dadda_cla8_out[10] = u_dadda_cla8_u_cla14_out[9];
  assign u_dadda_cla8_out[11] = u_dadda_cla8_u_cla14_out[10];
  assign u_dadda_cla8_out[12] = u_dadda_cla8_u_cla14_out[11];
  assign u_dadda_cla8_out[13] = u_dadda_cla8_u_cla14_out[12];
  assign u_dadda_cla8_out[14] = u_dadda_cla8_u_cla14_out[13];
  assign u_dadda_cla8_out[15] = u_dadda_cla8_u_cla14_out[14];
endmodule