module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module nor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a | _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module constant_wire_value_0(input a, input b, output constant_wire_0);
  wire constant_wire_value_0_a;
  wire constant_wire_value_0_b;

  assign constant_wire_value_0_a = a;
  assign constant_wire_value_0_b = b;

  xor_gate xor_gate_constant_wire_value_0_y0(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y0);
  xnor_gate xnor_gate_constant_wire_value_0_y1(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y1);
  nor_gate nor_gate_constant_wire_0(constant_wire_value_0_y0, constant_wire_value_0_y1, constant_wire_0);
endmodule

module pg_logic(input a, input b, output pg_logic_y0, output pg_logic_y1, output pg_logic_y2);
  wire pg_logic_a;
  wire pg_logic_b;

  assign pg_logic_a = a;
  assign pg_logic_b = b;

  or_gate or_gate_pg_logic_y0(pg_logic_a, pg_logic_b, pg_logic_y0);
  and_gate and_gate_pg_logic_y1(pg_logic_a, pg_logic_b, pg_logic_y1);
  xor_gate xor_gate_pg_logic_y2(pg_logic_a, pg_logic_b, pg_logic_y2);
endmodule

module h_u_cla32(input [31:0] a, input [31:0] b, output [32:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire a_30;
  wire a_31;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire b_30;
  wire b_31;
  wire constant_wire_0;
  wire h_u_cla32_pg_logic0_y0;
  wire h_u_cla32_pg_logic0_y1;
  wire h_u_cla32_pg_logic0_y2;
  wire h_u_cla32_xor0_y0;
  wire h_u_cla32_and0_y0;
  wire h_u_cla32_or0_y0;
  wire h_u_cla32_pg_logic1_y0;
  wire h_u_cla32_pg_logic1_y1;
  wire h_u_cla32_pg_logic1_y2;
  wire h_u_cla32_xor1_y0;
  wire h_u_cla32_and1_y0;
  wire h_u_cla32_and2_y0;
  wire h_u_cla32_and3_y0;
  wire h_u_cla32_and4_y0;
  wire h_u_cla32_or1_y0;
  wire h_u_cla32_or2_y0;
  wire h_u_cla32_pg_logic2_y0;
  wire h_u_cla32_pg_logic2_y1;
  wire h_u_cla32_pg_logic2_y2;
  wire h_u_cla32_xor2_y0;
  wire h_u_cla32_and5_y0;
  wire h_u_cla32_and6_y0;
  wire h_u_cla32_and7_y0;
  wire h_u_cla32_and8_y0;
  wire h_u_cla32_and9_y0;
  wire h_u_cla32_and10_y0;
  wire h_u_cla32_and11_y0;
  wire h_u_cla32_and12_y0;
  wire h_u_cla32_and13_y0;
  wire h_u_cla32_or3_y0;
  wire h_u_cla32_or4_y0;
  wire h_u_cla32_or5_y0;
  wire h_u_cla32_pg_logic3_y0;
  wire h_u_cla32_pg_logic3_y1;
  wire h_u_cla32_pg_logic3_y2;
  wire h_u_cla32_xor3_y0;
  wire h_u_cla32_and14_y0;
  wire h_u_cla32_and15_y0;
  wire h_u_cla32_and16_y0;
  wire h_u_cla32_and17_y0;
  wire h_u_cla32_and18_y0;
  wire h_u_cla32_and19_y0;
  wire h_u_cla32_and20_y0;
  wire h_u_cla32_and21_y0;
  wire h_u_cla32_and22_y0;
  wire h_u_cla32_and23_y0;
  wire h_u_cla32_and24_y0;
  wire h_u_cla32_and25_y0;
  wire h_u_cla32_and26_y0;
  wire h_u_cla32_and27_y0;
  wire h_u_cla32_and28_y0;
  wire h_u_cla32_and29_y0;
  wire h_u_cla32_or6_y0;
  wire h_u_cla32_or7_y0;
  wire h_u_cla32_or8_y0;
  wire h_u_cla32_or9_y0;
  wire h_u_cla32_pg_logic4_y0;
  wire h_u_cla32_pg_logic4_y1;
  wire h_u_cla32_pg_logic4_y2;
  wire h_u_cla32_xor4_y0;
  wire h_u_cla32_and30_y0;
  wire h_u_cla32_and31_y0;
  wire h_u_cla32_and32_y0;
  wire h_u_cla32_and33_y0;
  wire h_u_cla32_and34_y0;
  wire h_u_cla32_and35_y0;
  wire h_u_cla32_and36_y0;
  wire h_u_cla32_and37_y0;
  wire h_u_cla32_and38_y0;
  wire h_u_cla32_and39_y0;
  wire h_u_cla32_and40_y0;
  wire h_u_cla32_and41_y0;
  wire h_u_cla32_and42_y0;
  wire h_u_cla32_and43_y0;
  wire h_u_cla32_and44_y0;
  wire h_u_cla32_and45_y0;
  wire h_u_cla32_and46_y0;
  wire h_u_cla32_and47_y0;
  wire h_u_cla32_and48_y0;
  wire h_u_cla32_and49_y0;
  wire h_u_cla32_and50_y0;
  wire h_u_cla32_and51_y0;
  wire h_u_cla32_and52_y0;
  wire h_u_cla32_and53_y0;
  wire h_u_cla32_and54_y0;
  wire h_u_cla32_or10_y0;
  wire h_u_cla32_or11_y0;
  wire h_u_cla32_or12_y0;
  wire h_u_cla32_or13_y0;
  wire h_u_cla32_or14_y0;
  wire h_u_cla32_pg_logic5_y0;
  wire h_u_cla32_pg_logic5_y1;
  wire h_u_cla32_pg_logic5_y2;
  wire h_u_cla32_xor5_y0;
  wire h_u_cla32_and55_y0;
  wire h_u_cla32_and56_y0;
  wire h_u_cla32_and57_y0;
  wire h_u_cla32_and58_y0;
  wire h_u_cla32_and59_y0;
  wire h_u_cla32_and60_y0;
  wire h_u_cla32_and61_y0;
  wire h_u_cla32_and62_y0;
  wire h_u_cla32_and63_y0;
  wire h_u_cla32_and64_y0;
  wire h_u_cla32_and65_y0;
  wire h_u_cla32_and66_y0;
  wire h_u_cla32_and67_y0;
  wire h_u_cla32_and68_y0;
  wire h_u_cla32_and69_y0;
  wire h_u_cla32_and70_y0;
  wire h_u_cla32_and71_y0;
  wire h_u_cla32_and72_y0;
  wire h_u_cla32_and73_y0;
  wire h_u_cla32_and74_y0;
  wire h_u_cla32_and75_y0;
  wire h_u_cla32_and76_y0;
  wire h_u_cla32_and77_y0;
  wire h_u_cla32_and78_y0;
  wire h_u_cla32_and79_y0;
  wire h_u_cla32_and80_y0;
  wire h_u_cla32_and81_y0;
  wire h_u_cla32_and82_y0;
  wire h_u_cla32_and83_y0;
  wire h_u_cla32_and84_y0;
  wire h_u_cla32_and85_y0;
  wire h_u_cla32_and86_y0;
  wire h_u_cla32_and87_y0;
  wire h_u_cla32_and88_y0;
  wire h_u_cla32_and89_y0;
  wire h_u_cla32_and90_y0;
  wire h_u_cla32_or15_y0;
  wire h_u_cla32_or16_y0;
  wire h_u_cla32_or17_y0;
  wire h_u_cla32_or18_y0;
  wire h_u_cla32_or19_y0;
  wire h_u_cla32_or20_y0;
  wire h_u_cla32_pg_logic6_y0;
  wire h_u_cla32_pg_logic6_y1;
  wire h_u_cla32_pg_logic6_y2;
  wire h_u_cla32_xor6_y0;
  wire h_u_cla32_and91_y0;
  wire h_u_cla32_and92_y0;
  wire h_u_cla32_and93_y0;
  wire h_u_cla32_and94_y0;
  wire h_u_cla32_and95_y0;
  wire h_u_cla32_and96_y0;
  wire h_u_cla32_and97_y0;
  wire h_u_cla32_and98_y0;
  wire h_u_cla32_and99_y0;
  wire h_u_cla32_and100_y0;
  wire h_u_cla32_and101_y0;
  wire h_u_cla32_and102_y0;
  wire h_u_cla32_and103_y0;
  wire h_u_cla32_and104_y0;
  wire h_u_cla32_and105_y0;
  wire h_u_cla32_and106_y0;
  wire h_u_cla32_and107_y0;
  wire h_u_cla32_and108_y0;
  wire h_u_cla32_and109_y0;
  wire h_u_cla32_and110_y0;
  wire h_u_cla32_and111_y0;
  wire h_u_cla32_and112_y0;
  wire h_u_cla32_and113_y0;
  wire h_u_cla32_and114_y0;
  wire h_u_cla32_and115_y0;
  wire h_u_cla32_and116_y0;
  wire h_u_cla32_and117_y0;
  wire h_u_cla32_and118_y0;
  wire h_u_cla32_and119_y0;
  wire h_u_cla32_and120_y0;
  wire h_u_cla32_and121_y0;
  wire h_u_cla32_and122_y0;
  wire h_u_cla32_and123_y0;
  wire h_u_cla32_and124_y0;
  wire h_u_cla32_and125_y0;
  wire h_u_cla32_and126_y0;
  wire h_u_cla32_and127_y0;
  wire h_u_cla32_and128_y0;
  wire h_u_cla32_and129_y0;
  wire h_u_cla32_and130_y0;
  wire h_u_cla32_and131_y0;
  wire h_u_cla32_and132_y0;
  wire h_u_cla32_and133_y0;
  wire h_u_cla32_and134_y0;
  wire h_u_cla32_and135_y0;
  wire h_u_cla32_and136_y0;
  wire h_u_cla32_and137_y0;
  wire h_u_cla32_and138_y0;
  wire h_u_cla32_and139_y0;
  wire h_u_cla32_or21_y0;
  wire h_u_cla32_or22_y0;
  wire h_u_cla32_or23_y0;
  wire h_u_cla32_or24_y0;
  wire h_u_cla32_or25_y0;
  wire h_u_cla32_or26_y0;
  wire h_u_cla32_or27_y0;
  wire h_u_cla32_pg_logic7_y0;
  wire h_u_cla32_pg_logic7_y1;
  wire h_u_cla32_pg_logic7_y2;
  wire h_u_cla32_xor7_y0;
  wire h_u_cla32_and140_y0;
  wire h_u_cla32_and141_y0;
  wire h_u_cla32_and142_y0;
  wire h_u_cla32_and143_y0;
  wire h_u_cla32_and144_y0;
  wire h_u_cla32_and145_y0;
  wire h_u_cla32_and146_y0;
  wire h_u_cla32_and147_y0;
  wire h_u_cla32_and148_y0;
  wire h_u_cla32_and149_y0;
  wire h_u_cla32_and150_y0;
  wire h_u_cla32_and151_y0;
  wire h_u_cla32_and152_y0;
  wire h_u_cla32_and153_y0;
  wire h_u_cla32_and154_y0;
  wire h_u_cla32_and155_y0;
  wire h_u_cla32_and156_y0;
  wire h_u_cla32_and157_y0;
  wire h_u_cla32_and158_y0;
  wire h_u_cla32_and159_y0;
  wire h_u_cla32_and160_y0;
  wire h_u_cla32_and161_y0;
  wire h_u_cla32_and162_y0;
  wire h_u_cla32_and163_y0;
  wire h_u_cla32_and164_y0;
  wire h_u_cla32_and165_y0;
  wire h_u_cla32_and166_y0;
  wire h_u_cla32_and167_y0;
  wire h_u_cla32_and168_y0;
  wire h_u_cla32_and169_y0;
  wire h_u_cla32_and170_y0;
  wire h_u_cla32_and171_y0;
  wire h_u_cla32_and172_y0;
  wire h_u_cla32_and173_y0;
  wire h_u_cla32_and174_y0;
  wire h_u_cla32_and175_y0;
  wire h_u_cla32_and176_y0;
  wire h_u_cla32_and177_y0;
  wire h_u_cla32_and178_y0;
  wire h_u_cla32_and179_y0;
  wire h_u_cla32_and180_y0;
  wire h_u_cla32_and181_y0;
  wire h_u_cla32_and182_y0;
  wire h_u_cla32_and183_y0;
  wire h_u_cla32_and184_y0;
  wire h_u_cla32_and185_y0;
  wire h_u_cla32_and186_y0;
  wire h_u_cla32_and187_y0;
  wire h_u_cla32_and188_y0;
  wire h_u_cla32_and189_y0;
  wire h_u_cla32_and190_y0;
  wire h_u_cla32_and191_y0;
  wire h_u_cla32_and192_y0;
  wire h_u_cla32_and193_y0;
  wire h_u_cla32_and194_y0;
  wire h_u_cla32_and195_y0;
  wire h_u_cla32_and196_y0;
  wire h_u_cla32_and197_y0;
  wire h_u_cla32_and198_y0;
  wire h_u_cla32_and199_y0;
  wire h_u_cla32_and200_y0;
  wire h_u_cla32_and201_y0;
  wire h_u_cla32_and202_y0;
  wire h_u_cla32_and203_y0;
  wire h_u_cla32_or28_y0;
  wire h_u_cla32_or29_y0;
  wire h_u_cla32_or30_y0;
  wire h_u_cla32_or31_y0;
  wire h_u_cla32_or32_y0;
  wire h_u_cla32_or33_y0;
  wire h_u_cla32_or34_y0;
  wire h_u_cla32_or35_y0;
  wire h_u_cla32_pg_logic8_y0;
  wire h_u_cla32_pg_logic8_y1;
  wire h_u_cla32_pg_logic8_y2;
  wire h_u_cla32_xor8_y0;
  wire h_u_cla32_and204_y0;
  wire h_u_cla32_and205_y0;
  wire h_u_cla32_and206_y0;
  wire h_u_cla32_and207_y0;
  wire h_u_cla32_and208_y0;
  wire h_u_cla32_and209_y0;
  wire h_u_cla32_and210_y0;
  wire h_u_cla32_and211_y0;
  wire h_u_cla32_and212_y0;
  wire h_u_cla32_and213_y0;
  wire h_u_cla32_and214_y0;
  wire h_u_cla32_and215_y0;
  wire h_u_cla32_and216_y0;
  wire h_u_cla32_and217_y0;
  wire h_u_cla32_and218_y0;
  wire h_u_cla32_and219_y0;
  wire h_u_cla32_and220_y0;
  wire h_u_cla32_and221_y0;
  wire h_u_cla32_and222_y0;
  wire h_u_cla32_and223_y0;
  wire h_u_cla32_and224_y0;
  wire h_u_cla32_and225_y0;
  wire h_u_cla32_and226_y0;
  wire h_u_cla32_and227_y0;
  wire h_u_cla32_and228_y0;
  wire h_u_cla32_and229_y0;
  wire h_u_cla32_and230_y0;
  wire h_u_cla32_and231_y0;
  wire h_u_cla32_and232_y0;
  wire h_u_cla32_and233_y0;
  wire h_u_cla32_and234_y0;
  wire h_u_cla32_and235_y0;
  wire h_u_cla32_and236_y0;
  wire h_u_cla32_and237_y0;
  wire h_u_cla32_and238_y0;
  wire h_u_cla32_and239_y0;
  wire h_u_cla32_and240_y0;
  wire h_u_cla32_and241_y0;
  wire h_u_cla32_and242_y0;
  wire h_u_cla32_and243_y0;
  wire h_u_cla32_and244_y0;
  wire h_u_cla32_and245_y0;
  wire h_u_cla32_and246_y0;
  wire h_u_cla32_and247_y0;
  wire h_u_cla32_and248_y0;
  wire h_u_cla32_and249_y0;
  wire h_u_cla32_and250_y0;
  wire h_u_cla32_and251_y0;
  wire h_u_cla32_and252_y0;
  wire h_u_cla32_and253_y0;
  wire h_u_cla32_and254_y0;
  wire h_u_cla32_and255_y0;
  wire h_u_cla32_and256_y0;
  wire h_u_cla32_and257_y0;
  wire h_u_cla32_and258_y0;
  wire h_u_cla32_and259_y0;
  wire h_u_cla32_and260_y0;
  wire h_u_cla32_and261_y0;
  wire h_u_cla32_and262_y0;
  wire h_u_cla32_and263_y0;
  wire h_u_cla32_and264_y0;
  wire h_u_cla32_and265_y0;
  wire h_u_cla32_and266_y0;
  wire h_u_cla32_and267_y0;
  wire h_u_cla32_and268_y0;
  wire h_u_cla32_and269_y0;
  wire h_u_cla32_and270_y0;
  wire h_u_cla32_and271_y0;
  wire h_u_cla32_and272_y0;
  wire h_u_cla32_and273_y0;
  wire h_u_cla32_and274_y0;
  wire h_u_cla32_and275_y0;
  wire h_u_cla32_and276_y0;
  wire h_u_cla32_and277_y0;
  wire h_u_cla32_and278_y0;
  wire h_u_cla32_and279_y0;
  wire h_u_cla32_and280_y0;
  wire h_u_cla32_and281_y0;
  wire h_u_cla32_and282_y0;
  wire h_u_cla32_and283_y0;
  wire h_u_cla32_and284_y0;
  wire h_u_cla32_or36_y0;
  wire h_u_cla32_or37_y0;
  wire h_u_cla32_or38_y0;
  wire h_u_cla32_or39_y0;
  wire h_u_cla32_or40_y0;
  wire h_u_cla32_or41_y0;
  wire h_u_cla32_or42_y0;
  wire h_u_cla32_or43_y0;
  wire h_u_cla32_or44_y0;
  wire h_u_cla32_pg_logic9_y0;
  wire h_u_cla32_pg_logic9_y1;
  wire h_u_cla32_pg_logic9_y2;
  wire h_u_cla32_xor9_y0;
  wire h_u_cla32_and285_y0;
  wire h_u_cla32_and286_y0;
  wire h_u_cla32_and287_y0;
  wire h_u_cla32_and288_y0;
  wire h_u_cla32_and289_y0;
  wire h_u_cla32_and290_y0;
  wire h_u_cla32_and291_y0;
  wire h_u_cla32_and292_y0;
  wire h_u_cla32_and293_y0;
  wire h_u_cla32_and294_y0;
  wire h_u_cla32_and295_y0;
  wire h_u_cla32_and296_y0;
  wire h_u_cla32_and297_y0;
  wire h_u_cla32_and298_y0;
  wire h_u_cla32_and299_y0;
  wire h_u_cla32_and300_y0;
  wire h_u_cla32_and301_y0;
  wire h_u_cla32_and302_y0;
  wire h_u_cla32_and303_y0;
  wire h_u_cla32_and304_y0;
  wire h_u_cla32_and305_y0;
  wire h_u_cla32_and306_y0;
  wire h_u_cla32_and307_y0;
  wire h_u_cla32_and308_y0;
  wire h_u_cla32_and309_y0;
  wire h_u_cla32_and310_y0;
  wire h_u_cla32_and311_y0;
  wire h_u_cla32_and312_y0;
  wire h_u_cla32_and313_y0;
  wire h_u_cla32_and314_y0;
  wire h_u_cla32_and315_y0;
  wire h_u_cla32_and316_y0;
  wire h_u_cla32_and317_y0;
  wire h_u_cla32_and318_y0;
  wire h_u_cla32_and319_y0;
  wire h_u_cla32_and320_y0;
  wire h_u_cla32_and321_y0;
  wire h_u_cla32_and322_y0;
  wire h_u_cla32_and323_y0;
  wire h_u_cla32_and324_y0;
  wire h_u_cla32_and325_y0;
  wire h_u_cla32_and326_y0;
  wire h_u_cla32_and327_y0;
  wire h_u_cla32_and328_y0;
  wire h_u_cla32_and329_y0;
  wire h_u_cla32_and330_y0;
  wire h_u_cla32_and331_y0;
  wire h_u_cla32_and332_y0;
  wire h_u_cla32_and333_y0;
  wire h_u_cla32_and334_y0;
  wire h_u_cla32_and335_y0;
  wire h_u_cla32_and336_y0;
  wire h_u_cla32_and337_y0;
  wire h_u_cla32_and338_y0;
  wire h_u_cla32_and339_y0;
  wire h_u_cla32_and340_y0;
  wire h_u_cla32_and341_y0;
  wire h_u_cla32_and342_y0;
  wire h_u_cla32_and343_y0;
  wire h_u_cla32_and344_y0;
  wire h_u_cla32_and345_y0;
  wire h_u_cla32_and346_y0;
  wire h_u_cla32_and347_y0;
  wire h_u_cla32_and348_y0;
  wire h_u_cla32_and349_y0;
  wire h_u_cla32_and350_y0;
  wire h_u_cla32_and351_y0;
  wire h_u_cla32_and352_y0;
  wire h_u_cla32_and353_y0;
  wire h_u_cla32_and354_y0;
  wire h_u_cla32_and355_y0;
  wire h_u_cla32_and356_y0;
  wire h_u_cla32_and357_y0;
  wire h_u_cla32_and358_y0;
  wire h_u_cla32_and359_y0;
  wire h_u_cla32_and360_y0;
  wire h_u_cla32_and361_y0;
  wire h_u_cla32_and362_y0;
  wire h_u_cla32_and363_y0;
  wire h_u_cla32_and364_y0;
  wire h_u_cla32_and365_y0;
  wire h_u_cla32_and366_y0;
  wire h_u_cla32_and367_y0;
  wire h_u_cla32_and368_y0;
  wire h_u_cla32_and369_y0;
  wire h_u_cla32_and370_y0;
  wire h_u_cla32_and371_y0;
  wire h_u_cla32_and372_y0;
  wire h_u_cla32_and373_y0;
  wire h_u_cla32_and374_y0;
  wire h_u_cla32_and375_y0;
  wire h_u_cla32_and376_y0;
  wire h_u_cla32_and377_y0;
  wire h_u_cla32_and378_y0;
  wire h_u_cla32_and379_y0;
  wire h_u_cla32_and380_y0;
  wire h_u_cla32_and381_y0;
  wire h_u_cla32_and382_y0;
  wire h_u_cla32_and383_y0;
  wire h_u_cla32_and384_y0;
  wire h_u_cla32_or45_y0;
  wire h_u_cla32_or46_y0;
  wire h_u_cla32_or47_y0;
  wire h_u_cla32_or48_y0;
  wire h_u_cla32_or49_y0;
  wire h_u_cla32_or50_y0;
  wire h_u_cla32_or51_y0;
  wire h_u_cla32_or52_y0;
  wire h_u_cla32_or53_y0;
  wire h_u_cla32_or54_y0;
  wire h_u_cla32_pg_logic10_y0;
  wire h_u_cla32_pg_logic10_y1;
  wire h_u_cla32_pg_logic10_y2;
  wire h_u_cla32_xor10_y0;
  wire h_u_cla32_and385_y0;
  wire h_u_cla32_and386_y0;
  wire h_u_cla32_and387_y0;
  wire h_u_cla32_and388_y0;
  wire h_u_cla32_and389_y0;
  wire h_u_cla32_and390_y0;
  wire h_u_cla32_and391_y0;
  wire h_u_cla32_and392_y0;
  wire h_u_cla32_and393_y0;
  wire h_u_cla32_and394_y0;
  wire h_u_cla32_and395_y0;
  wire h_u_cla32_and396_y0;
  wire h_u_cla32_and397_y0;
  wire h_u_cla32_and398_y0;
  wire h_u_cla32_and399_y0;
  wire h_u_cla32_and400_y0;
  wire h_u_cla32_and401_y0;
  wire h_u_cla32_and402_y0;
  wire h_u_cla32_and403_y0;
  wire h_u_cla32_and404_y0;
  wire h_u_cla32_and405_y0;
  wire h_u_cla32_and406_y0;
  wire h_u_cla32_and407_y0;
  wire h_u_cla32_and408_y0;
  wire h_u_cla32_and409_y0;
  wire h_u_cla32_and410_y0;
  wire h_u_cla32_and411_y0;
  wire h_u_cla32_and412_y0;
  wire h_u_cla32_and413_y0;
  wire h_u_cla32_and414_y0;
  wire h_u_cla32_and415_y0;
  wire h_u_cla32_and416_y0;
  wire h_u_cla32_and417_y0;
  wire h_u_cla32_and418_y0;
  wire h_u_cla32_and419_y0;
  wire h_u_cla32_and420_y0;
  wire h_u_cla32_and421_y0;
  wire h_u_cla32_and422_y0;
  wire h_u_cla32_and423_y0;
  wire h_u_cla32_and424_y0;
  wire h_u_cla32_and425_y0;
  wire h_u_cla32_and426_y0;
  wire h_u_cla32_and427_y0;
  wire h_u_cla32_and428_y0;
  wire h_u_cla32_and429_y0;
  wire h_u_cla32_and430_y0;
  wire h_u_cla32_and431_y0;
  wire h_u_cla32_and432_y0;
  wire h_u_cla32_and433_y0;
  wire h_u_cla32_and434_y0;
  wire h_u_cla32_and435_y0;
  wire h_u_cla32_and436_y0;
  wire h_u_cla32_and437_y0;
  wire h_u_cla32_and438_y0;
  wire h_u_cla32_and439_y0;
  wire h_u_cla32_and440_y0;
  wire h_u_cla32_and441_y0;
  wire h_u_cla32_and442_y0;
  wire h_u_cla32_and443_y0;
  wire h_u_cla32_and444_y0;
  wire h_u_cla32_and445_y0;
  wire h_u_cla32_and446_y0;
  wire h_u_cla32_and447_y0;
  wire h_u_cla32_and448_y0;
  wire h_u_cla32_and449_y0;
  wire h_u_cla32_and450_y0;
  wire h_u_cla32_and451_y0;
  wire h_u_cla32_and452_y0;
  wire h_u_cla32_and453_y0;
  wire h_u_cla32_and454_y0;
  wire h_u_cla32_and455_y0;
  wire h_u_cla32_and456_y0;
  wire h_u_cla32_and457_y0;
  wire h_u_cla32_and458_y0;
  wire h_u_cla32_and459_y0;
  wire h_u_cla32_and460_y0;
  wire h_u_cla32_and461_y0;
  wire h_u_cla32_and462_y0;
  wire h_u_cla32_and463_y0;
  wire h_u_cla32_and464_y0;
  wire h_u_cla32_and465_y0;
  wire h_u_cla32_and466_y0;
  wire h_u_cla32_and467_y0;
  wire h_u_cla32_and468_y0;
  wire h_u_cla32_and469_y0;
  wire h_u_cla32_and470_y0;
  wire h_u_cla32_and471_y0;
  wire h_u_cla32_and472_y0;
  wire h_u_cla32_and473_y0;
  wire h_u_cla32_and474_y0;
  wire h_u_cla32_and475_y0;
  wire h_u_cla32_and476_y0;
  wire h_u_cla32_and477_y0;
  wire h_u_cla32_and478_y0;
  wire h_u_cla32_and479_y0;
  wire h_u_cla32_and480_y0;
  wire h_u_cla32_and481_y0;
  wire h_u_cla32_and482_y0;
  wire h_u_cla32_and483_y0;
  wire h_u_cla32_and484_y0;
  wire h_u_cla32_and485_y0;
  wire h_u_cla32_and486_y0;
  wire h_u_cla32_and487_y0;
  wire h_u_cla32_and488_y0;
  wire h_u_cla32_and489_y0;
  wire h_u_cla32_and490_y0;
  wire h_u_cla32_and491_y0;
  wire h_u_cla32_and492_y0;
  wire h_u_cla32_and493_y0;
  wire h_u_cla32_and494_y0;
  wire h_u_cla32_and495_y0;
  wire h_u_cla32_and496_y0;
  wire h_u_cla32_and497_y0;
  wire h_u_cla32_and498_y0;
  wire h_u_cla32_and499_y0;
  wire h_u_cla32_and500_y0;
  wire h_u_cla32_and501_y0;
  wire h_u_cla32_and502_y0;
  wire h_u_cla32_and503_y0;
  wire h_u_cla32_and504_y0;
  wire h_u_cla32_and505_y0;
  wire h_u_cla32_or55_y0;
  wire h_u_cla32_or56_y0;
  wire h_u_cla32_or57_y0;
  wire h_u_cla32_or58_y0;
  wire h_u_cla32_or59_y0;
  wire h_u_cla32_or60_y0;
  wire h_u_cla32_or61_y0;
  wire h_u_cla32_or62_y0;
  wire h_u_cla32_or63_y0;
  wire h_u_cla32_or64_y0;
  wire h_u_cla32_or65_y0;
  wire h_u_cla32_pg_logic11_y0;
  wire h_u_cla32_pg_logic11_y1;
  wire h_u_cla32_pg_logic11_y2;
  wire h_u_cla32_xor11_y0;
  wire h_u_cla32_and506_y0;
  wire h_u_cla32_and507_y0;
  wire h_u_cla32_and508_y0;
  wire h_u_cla32_and509_y0;
  wire h_u_cla32_and510_y0;
  wire h_u_cla32_and511_y0;
  wire h_u_cla32_and512_y0;
  wire h_u_cla32_and513_y0;
  wire h_u_cla32_and514_y0;
  wire h_u_cla32_and515_y0;
  wire h_u_cla32_and516_y0;
  wire h_u_cla32_and517_y0;
  wire h_u_cla32_and518_y0;
  wire h_u_cla32_and519_y0;
  wire h_u_cla32_and520_y0;
  wire h_u_cla32_and521_y0;
  wire h_u_cla32_and522_y0;
  wire h_u_cla32_and523_y0;
  wire h_u_cla32_and524_y0;
  wire h_u_cla32_and525_y0;
  wire h_u_cla32_and526_y0;
  wire h_u_cla32_and527_y0;
  wire h_u_cla32_and528_y0;
  wire h_u_cla32_and529_y0;
  wire h_u_cla32_and530_y0;
  wire h_u_cla32_and531_y0;
  wire h_u_cla32_and532_y0;
  wire h_u_cla32_and533_y0;
  wire h_u_cla32_and534_y0;
  wire h_u_cla32_and535_y0;
  wire h_u_cla32_and536_y0;
  wire h_u_cla32_and537_y0;
  wire h_u_cla32_and538_y0;
  wire h_u_cla32_and539_y0;
  wire h_u_cla32_and540_y0;
  wire h_u_cla32_and541_y0;
  wire h_u_cla32_and542_y0;
  wire h_u_cla32_and543_y0;
  wire h_u_cla32_and544_y0;
  wire h_u_cla32_and545_y0;
  wire h_u_cla32_and546_y0;
  wire h_u_cla32_and547_y0;
  wire h_u_cla32_and548_y0;
  wire h_u_cla32_and549_y0;
  wire h_u_cla32_and550_y0;
  wire h_u_cla32_and551_y0;
  wire h_u_cla32_and552_y0;
  wire h_u_cla32_and553_y0;
  wire h_u_cla32_and554_y0;
  wire h_u_cla32_and555_y0;
  wire h_u_cla32_and556_y0;
  wire h_u_cla32_and557_y0;
  wire h_u_cla32_and558_y0;
  wire h_u_cla32_and559_y0;
  wire h_u_cla32_and560_y0;
  wire h_u_cla32_and561_y0;
  wire h_u_cla32_and562_y0;
  wire h_u_cla32_and563_y0;
  wire h_u_cla32_and564_y0;
  wire h_u_cla32_and565_y0;
  wire h_u_cla32_and566_y0;
  wire h_u_cla32_and567_y0;
  wire h_u_cla32_and568_y0;
  wire h_u_cla32_and569_y0;
  wire h_u_cla32_and570_y0;
  wire h_u_cla32_and571_y0;
  wire h_u_cla32_and572_y0;
  wire h_u_cla32_and573_y0;
  wire h_u_cla32_and574_y0;
  wire h_u_cla32_and575_y0;
  wire h_u_cla32_and576_y0;
  wire h_u_cla32_and577_y0;
  wire h_u_cla32_and578_y0;
  wire h_u_cla32_and579_y0;
  wire h_u_cla32_and580_y0;
  wire h_u_cla32_and581_y0;
  wire h_u_cla32_and582_y0;
  wire h_u_cla32_and583_y0;
  wire h_u_cla32_and584_y0;
  wire h_u_cla32_and585_y0;
  wire h_u_cla32_and586_y0;
  wire h_u_cla32_and587_y0;
  wire h_u_cla32_and588_y0;
  wire h_u_cla32_and589_y0;
  wire h_u_cla32_and590_y0;
  wire h_u_cla32_and591_y0;
  wire h_u_cla32_and592_y0;
  wire h_u_cla32_and593_y0;
  wire h_u_cla32_and594_y0;
  wire h_u_cla32_and595_y0;
  wire h_u_cla32_and596_y0;
  wire h_u_cla32_and597_y0;
  wire h_u_cla32_and598_y0;
  wire h_u_cla32_and599_y0;
  wire h_u_cla32_and600_y0;
  wire h_u_cla32_and601_y0;
  wire h_u_cla32_and602_y0;
  wire h_u_cla32_and603_y0;
  wire h_u_cla32_and604_y0;
  wire h_u_cla32_and605_y0;
  wire h_u_cla32_and606_y0;
  wire h_u_cla32_and607_y0;
  wire h_u_cla32_and608_y0;
  wire h_u_cla32_and609_y0;
  wire h_u_cla32_and610_y0;
  wire h_u_cla32_and611_y0;
  wire h_u_cla32_and612_y0;
  wire h_u_cla32_and613_y0;
  wire h_u_cla32_and614_y0;
  wire h_u_cla32_and615_y0;
  wire h_u_cla32_and616_y0;
  wire h_u_cla32_and617_y0;
  wire h_u_cla32_and618_y0;
  wire h_u_cla32_and619_y0;
  wire h_u_cla32_and620_y0;
  wire h_u_cla32_and621_y0;
  wire h_u_cla32_and622_y0;
  wire h_u_cla32_and623_y0;
  wire h_u_cla32_and624_y0;
  wire h_u_cla32_and625_y0;
  wire h_u_cla32_and626_y0;
  wire h_u_cla32_and627_y0;
  wire h_u_cla32_and628_y0;
  wire h_u_cla32_and629_y0;
  wire h_u_cla32_and630_y0;
  wire h_u_cla32_and631_y0;
  wire h_u_cla32_and632_y0;
  wire h_u_cla32_and633_y0;
  wire h_u_cla32_and634_y0;
  wire h_u_cla32_and635_y0;
  wire h_u_cla32_and636_y0;
  wire h_u_cla32_and637_y0;
  wire h_u_cla32_and638_y0;
  wire h_u_cla32_and639_y0;
  wire h_u_cla32_and640_y0;
  wire h_u_cla32_and641_y0;
  wire h_u_cla32_and642_y0;
  wire h_u_cla32_and643_y0;
  wire h_u_cla32_and644_y0;
  wire h_u_cla32_and645_y0;
  wire h_u_cla32_and646_y0;
  wire h_u_cla32_and647_y0;
  wire h_u_cla32_and648_y0;
  wire h_u_cla32_and649_y0;
  wire h_u_cla32_or66_y0;
  wire h_u_cla32_or67_y0;
  wire h_u_cla32_or68_y0;
  wire h_u_cla32_or69_y0;
  wire h_u_cla32_or70_y0;
  wire h_u_cla32_or71_y0;
  wire h_u_cla32_or72_y0;
  wire h_u_cla32_or73_y0;
  wire h_u_cla32_or74_y0;
  wire h_u_cla32_or75_y0;
  wire h_u_cla32_or76_y0;
  wire h_u_cla32_or77_y0;
  wire h_u_cla32_pg_logic12_y0;
  wire h_u_cla32_pg_logic12_y1;
  wire h_u_cla32_pg_logic12_y2;
  wire h_u_cla32_xor12_y0;
  wire h_u_cla32_and650_y0;
  wire h_u_cla32_and651_y0;
  wire h_u_cla32_and652_y0;
  wire h_u_cla32_and653_y0;
  wire h_u_cla32_and654_y0;
  wire h_u_cla32_and655_y0;
  wire h_u_cla32_and656_y0;
  wire h_u_cla32_and657_y0;
  wire h_u_cla32_and658_y0;
  wire h_u_cla32_and659_y0;
  wire h_u_cla32_and660_y0;
  wire h_u_cla32_and661_y0;
  wire h_u_cla32_and662_y0;
  wire h_u_cla32_and663_y0;
  wire h_u_cla32_and664_y0;
  wire h_u_cla32_and665_y0;
  wire h_u_cla32_and666_y0;
  wire h_u_cla32_and667_y0;
  wire h_u_cla32_and668_y0;
  wire h_u_cla32_and669_y0;
  wire h_u_cla32_and670_y0;
  wire h_u_cla32_and671_y0;
  wire h_u_cla32_and672_y0;
  wire h_u_cla32_and673_y0;
  wire h_u_cla32_and674_y0;
  wire h_u_cla32_and675_y0;
  wire h_u_cla32_and676_y0;
  wire h_u_cla32_and677_y0;
  wire h_u_cla32_and678_y0;
  wire h_u_cla32_and679_y0;
  wire h_u_cla32_and680_y0;
  wire h_u_cla32_and681_y0;
  wire h_u_cla32_and682_y0;
  wire h_u_cla32_and683_y0;
  wire h_u_cla32_and684_y0;
  wire h_u_cla32_and685_y0;
  wire h_u_cla32_and686_y0;
  wire h_u_cla32_and687_y0;
  wire h_u_cla32_and688_y0;
  wire h_u_cla32_and689_y0;
  wire h_u_cla32_and690_y0;
  wire h_u_cla32_and691_y0;
  wire h_u_cla32_and692_y0;
  wire h_u_cla32_and693_y0;
  wire h_u_cla32_and694_y0;
  wire h_u_cla32_and695_y0;
  wire h_u_cla32_and696_y0;
  wire h_u_cla32_and697_y0;
  wire h_u_cla32_and698_y0;
  wire h_u_cla32_and699_y0;
  wire h_u_cla32_and700_y0;
  wire h_u_cla32_and701_y0;
  wire h_u_cla32_and702_y0;
  wire h_u_cla32_and703_y0;
  wire h_u_cla32_and704_y0;
  wire h_u_cla32_and705_y0;
  wire h_u_cla32_and706_y0;
  wire h_u_cla32_and707_y0;
  wire h_u_cla32_and708_y0;
  wire h_u_cla32_and709_y0;
  wire h_u_cla32_and710_y0;
  wire h_u_cla32_and711_y0;
  wire h_u_cla32_and712_y0;
  wire h_u_cla32_and713_y0;
  wire h_u_cla32_and714_y0;
  wire h_u_cla32_and715_y0;
  wire h_u_cla32_and716_y0;
  wire h_u_cla32_and717_y0;
  wire h_u_cla32_and718_y0;
  wire h_u_cla32_and719_y0;
  wire h_u_cla32_and720_y0;
  wire h_u_cla32_and721_y0;
  wire h_u_cla32_and722_y0;
  wire h_u_cla32_and723_y0;
  wire h_u_cla32_and724_y0;
  wire h_u_cla32_and725_y0;
  wire h_u_cla32_and726_y0;
  wire h_u_cla32_and727_y0;
  wire h_u_cla32_and728_y0;
  wire h_u_cla32_and729_y0;
  wire h_u_cla32_and730_y0;
  wire h_u_cla32_and731_y0;
  wire h_u_cla32_and732_y0;
  wire h_u_cla32_and733_y0;
  wire h_u_cla32_and734_y0;
  wire h_u_cla32_and735_y0;
  wire h_u_cla32_and736_y0;
  wire h_u_cla32_and737_y0;
  wire h_u_cla32_and738_y0;
  wire h_u_cla32_and739_y0;
  wire h_u_cla32_and740_y0;
  wire h_u_cla32_and741_y0;
  wire h_u_cla32_and742_y0;
  wire h_u_cla32_and743_y0;
  wire h_u_cla32_and744_y0;
  wire h_u_cla32_and745_y0;
  wire h_u_cla32_and746_y0;
  wire h_u_cla32_and747_y0;
  wire h_u_cla32_and748_y0;
  wire h_u_cla32_and749_y0;
  wire h_u_cla32_and750_y0;
  wire h_u_cla32_and751_y0;
  wire h_u_cla32_and752_y0;
  wire h_u_cla32_and753_y0;
  wire h_u_cla32_and754_y0;
  wire h_u_cla32_and755_y0;
  wire h_u_cla32_and756_y0;
  wire h_u_cla32_and757_y0;
  wire h_u_cla32_and758_y0;
  wire h_u_cla32_and759_y0;
  wire h_u_cla32_and760_y0;
  wire h_u_cla32_and761_y0;
  wire h_u_cla32_and762_y0;
  wire h_u_cla32_and763_y0;
  wire h_u_cla32_and764_y0;
  wire h_u_cla32_and765_y0;
  wire h_u_cla32_and766_y0;
  wire h_u_cla32_and767_y0;
  wire h_u_cla32_and768_y0;
  wire h_u_cla32_and769_y0;
  wire h_u_cla32_and770_y0;
  wire h_u_cla32_and771_y0;
  wire h_u_cla32_and772_y0;
  wire h_u_cla32_and773_y0;
  wire h_u_cla32_and774_y0;
  wire h_u_cla32_and775_y0;
  wire h_u_cla32_and776_y0;
  wire h_u_cla32_and777_y0;
  wire h_u_cla32_and778_y0;
  wire h_u_cla32_and779_y0;
  wire h_u_cla32_and780_y0;
  wire h_u_cla32_and781_y0;
  wire h_u_cla32_and782_y0;
  wire h_u_cla32_and783_y0;
  wire h_u_cla32_and784_y0;
  wire h_u_cla32_and785_y0;
  wire h_u_cla32_and786_y0;
  wire h_u_cla32_and787_y0;
  wire h_u_cla32_and788_y0;
  wire h_u_cla32_and789_y0;
  wire h_u_cla32_and790_y0;
  wire h_u_cla32_and791_y0;
  wire h_u_cla32_and792_y0;
  wire h_u_cla32_and793_y0;
  wire h_u_cla32_and794_y0;
  wire h_u_cla32_and795_y0;
  wire h_u_cla32_and796_y0;
  wire h_u_cla32_and797_y0;
  wire h_u_cla32_and798_y0;
  wire h_u_cla32_and799_y0;
  wire h_u_cla32_and800_y0;
  wire h_u_cla32_and801_y0;
  wire h_u_cla32_and802_y0;
  wire h_u_cla32_and803_y0;
  wire h_u_cla32_and804_y0;
  wire h_u_cla32_and805_y0;
  wire h_u_cla32_and806_y0;
  wire h_u_cla32_and807_y0;
  wire h_u_cla32_and808_y0;
  wire h_u_cla32_and809_y0;
  wire h_u_cla32_and810_y0;
  wire h_u_cla32_and811_y0;
  wire h_u_cla32_and812_y0;
  wire h_u_cla32_and813_y0;
  wire h_u_cla32_and814_y0;
  wire h_u_cla32_and815_y0;
  wire h_u_cla32_and816_y0;
  wire h_u_cla32_and817_y0;
  wire h_u_cla32_and818_y0;
  wire h_u_cla32_or78_y0;
  wire h_u_cla32_or79_y0;
  wire h_u_cla32_or80_y0;
  wire h_u_cla32_or81_y0;
  wire h_u_cla32_or82_y0;
  wire h_u_cla32_or83_y0;
  wire h_u_cla32_or84_y0;
  wire h_u_cla32_or85_y0;
  wire h_u_cla32_or86_y0;
  wire h_u_cla32_or87_y0;
  wire h_u_cla32_or88_y0;
  wire h_u_cla32_or89_y0;
  wire h_u_cla32_or90_y0;
  wire h_u_cla32_pg_logic13_y0;
  wire h_u_cla32_pg_logic13_y1;
  wire h_u_cla32_pg_logic13_y2;
  wire h_u_cla32_xor13_y0;
  wire h_u_cla32_and819_y0;
  wire h_u_cla32_and820_y0;
  wire h_u_cla32_and821_y0;
  wire h_u_cla32_and822_y0;
  wire h_u_cla32_and823_y0;
  wire h_u_cla32_and824_y0;
  wire h_u_cla32_and825_y0;
  wire h_u_cla32_and826_y0;
  wire h_u_cla32_and827_y0;
  wire h_u_cla32_and828_y0;
  wire h_u_cla32_and829_y0;
  wire h_u_cla32_and830_y0;
  wire h_u_cla32_and831_y0;
  wire h_u_cla32_and832_y0;
  wire h_u_cla32_and833_y0;
  wire h_u_cla32_and834_y0;
  wire h_u_cla32_and835_y0;
  wire h_u_cla32_and836_y0;
  wire h_u_cla32_and837_y0;
  wire h_u_cla32_and838_y0;
  wire h_u_cla32_and839_y0;
  wire h_u_cla32_and840_y0;
  wire h_u_cla32_and841_y0;
  wire h_u_cla32_and842_y0;
  wire h_u_cla32_and843_y0;
  wire h_u_cla32_and844_y0;
  wire h_u_cla32_and845_y0;
  wire h_u_cla32_and846_y0;
  wire h_u_cla32_and847_y0;
  wire h_u_cla32_and848_y0;
  wire h_u_cla32_and849_y0;
  wire h_u_cla32_and850_y0;
  wire h_u_cla32_and851_y0;
  wire h_u_cla32_and852_y0;
  wire h_u_cla32_and853_y0;
  wire h_u_cla32_and854_y0;
  wire h_u_cla32_and855_y0;
  wire h_u_cla32_and856_y0;
  wire h_u_cla32_and857_y0;
  wire h_u_cla32_and858_y0;
  wire h_u_cla32_and859_y0;
  wire h_u_cla32_and860_y0;
  wire h_u_cla32_and861_y0;
  wire h_u_cla32_and862_y0;
  wire h_u_cla32_and863_y0;
  wire h_u_cla32_and864_y0;
  wire h_u_cla32_and865_y0;
  wire h_u_cla32_and866_y0;
  wire h_u_cla32_and867_y0;
  wire h_u_cla32_and868_y0;
  wire h_u_cla32_and869_y0;
  wire h_u_cla32_and870_y0;
  wire h_u_cla32_and871_y0;
  wire h_u_cla32_and872_y0;
  wire h_u_cla32_and873_y0;
  wire h_u_cla32_and874_y0;
  wire h_u_cla32_and875_y0;
  wire h_u_cla32_and876_y0;
  wire h_u_cla32_and877_y0;
  wire h_u_cla32_and878_y0;
  wire h_u_cla32_and879_y0;
  wire h_u_cla32_and880_y0;
  wire h_u_cla32_and881_y0;
  wire h_u_cla32_and882_y0;
  wire h_u_cla32_and883_y0;
  wire h_u_cla32_and884_y0;
  wire h_u_cla32_and885_y0;
  wire h_u_cla32_and886_y0;
  wire h_u_cla32_and887_y0;
  wire h_u_cla32_and888_y0;
  wire h_u_cla32_and889_y0;
  wire h_u_cla32_and890_y0;
  wire h_u_cla32_and891_y0;
  wire h_u_cla32_and892_y0;
  wire h_u_cla32_and893_y0;
  wire h_u_cla32_and894_y0;
  wire h_u_cla32_and895_y0;
  wire h_u_cla32_and896_y0;
  wire h_u_cla32_and897_y0;
  wire h_u_cla32_and898_y0;
  wire h_u_cla32_and899_y0;
  wire h_u_cla32_and900_y0;
  wire h_u_cla32_and901_y0;
  wire h_u_cla32_and902_y0;
  wire h_u_cla32_and903_y0;
  wire h_u_cla32_and904_y0;
  wire h_u_cla32_and905_y0;
  wire h_u_cla32_and906_y0;
  wire h_u_cla32_and907_y0;
  wire h_u_cla32_and908_y0;
  wire h_u_cla32_and909_y0;
  wire h_u_cla32_and910_y0;
  wire h_u_cla32_and911_y0;
  wire h_u_cla32_and912_y0;
  wire h_u_cla32_and913_y0;
  wire h_u_cla32_and914_y0;
  wire h_u_cla32_and915_y0;
  wire h_u_cla32_and916_y0;
  wire h_u_cla32_and917_y0;
  wire h_u_cla32_and918_y0;
  wire h_u_cla32_and919_y0;
  wire h_u_cla32_and920_y0;
  wire h_u_cla32_and921_y0;
  wire h_u_cla32_and922_y0;
  wire h_u_cla32_and923_y0;
  wire h_u_cla32_and924_y0;
  wire h_u_cla32_and925_y0;
  wire h_u_cla32_and926_y0;
  wire h_u_cla32_and927_y0;
  wire h_u_cla32_and928_y0;
  wire h_u_cla32_and929_y0;
  wire h_u_cla32_and930_y0;
  wire h_u_cla32_and931_y0;
  wire h_u_cla32_and932_y0;
  wire h_u_cla32_and933_y0;
  wire h_u_cla32_and934_y0;
  wire h_u_cla32_and935_y0;
  wire h_u_cla32_and936_y0;
  wire h_u_cla32_and937_y0;
  wire h_u_cla32_and938_y0;
  wire h_u_cla32_and939_y0;
  wire h_u_cla32_and940_y0;
  wire h_u_cla32_and941_y0;
  wire h_u_cla32_and942_y0;
  wire h_u_cla32_and943_y0;
  wire h_u_cla32_and944_y0;
  wire h_u_cla32_and945_y0;
  wire h_u_cla32_and946_y0;
  wire h_u_cla32_and947_y0;
  wire h_u_cla32_and948_y0;
  wire h_u_cla32_and949_y0;
  wire h_u_cla32_and950_y0;
  wire h_u_cla32_and951_y0;
  wire h_u_cla32_and952_y0;
  wire h_u_cla32_and953_y0;
  wire h_u_cla32_and954_y0;
  wire h_u_cla32_and955_y0;
  wire h_u_cla32_and956_y0;
  wire h_u_cla32_and957_y0;
  wire h_u_cla32_and958_y0;
  wire h_u_cla32_and959_y0;
  wire h_u_cla32_and960_y0;
  wire h_u_cla32_and961_y0;
  wire h_u_cla32_and962_y0;
  wire h_u_cla32_and963_y0;
  wire h_u_cla32_and964_y0;
  wire h_u_cla32_and965_y0;
  wire h_u_cla32_and966_y0;
  wire h_u_cla32_and967_y0;
  wire h_u_cla32_and968_y0;
  wire h_u_cla32_and969_y0;
  wire h_u_cla32_and970_y0;
  wire h_u_cla32_and971_y0;
  wire h_u_cla32_and972_y0;
  wire h_u_cla32_and973_y0;
  wire h_u_cla32_and974_y0;
  wire h_u_cla32_and975_y0;
  wire h_u_cla32_and976_y0;
  wire h_u_cla32_and977_y0;
  wire h_u_cla32_and978_y0;
  wire h_u_cla32_and979_y0;
  wire h_u_cla32_and980_y0;
  wire h_u_cla32_and981_y0;
  wire h_u_cla32_and982_y0;
  wire h_u_cla32_and983_y0;
  wire h_u_cla32_and984_y0;
  wire h_u_cla32_and985_y0;
  wire h_u_cla32_and986_y0;
  wire h_u_cla32_and987_y0;
  wire h_u_cla32_and988_y0;
  wire h_u_cla32_and989_y0;
  wire h_u_cla32_and990_y0;
  wire h_u_cla32_and991_y0;
  wire h_u_cla32_and992_y0;
  wire h_u_cla32_and993_y0;
  wire h_u_cla32_and994_y0;
  wire h_u_cla32_and995_y0;
  wire h_u_cla32_and996_y0;
  wire h_u_cla32_and997_y0;
  wire h_u_cla32_and998_y0;
  wire h_u_cla32_and999_y0;
  wire h_u_cla32_and1000_y0;
  wire h_u_cla32_and1001_y0;
  wire h_u_cla32_and1002_y0;
  wire h_u_cla32_and1003_y0;
  wire h_u_cla32_and1004_y0;
  wire h_u_cla32_and1005_y0;
  wire h_u_cla32_and1006_y0;
  wire h_u_cla32_and1007_y0;
  wire h_u_cla32_and1008_y0;
  wire h_u_cla32_and1009_y0;
  wire h_u_cla32_and1010_y0;
  wire h_u_cla32_and1011_y0;
  wire h_u_cla32_and1012_y0;
  wire h_u_cla32_and1013_y0;
  wire h_u_cla32_and1014_y0;
  wire h_u_cla32_or91_y0;
  wire h_u_cla32_or92_y0;
  wire h_u_cla32_or93_y0;
  wire h_u_cla32_or94_y0;
  wire h_u_cla32_or95_y0;
  wire h_u_cla32_or96_y0;
  wire h_u_cla32_or97_y0;
  wire h_u_cla32_or98_y0;
  wire h_u_cla32_or99_y0;
  wire h_u_cla32_or100_y0;
  wire h_u_cla32_or101_y0;
  wire h_u_cla32_or102_y0;
  wire h_u_cla32_or103_y0;
  wire h_u_cla32_or104_y0;
  wire h_u_cla32_pg_logic14_y0;
  wire h_u_cla32_pg_logic14_y1;
  wire h_u_cla32_pg_logic14_y2;
  wire h_u_cla32_xor14_y0;
  wire h_u_cla32_and1015_y0;
  wire h_u_cla32_and1016_y0;
  wire h_u_cla32_and1017_y0;
  wire h_u_cla32_and1018_y0;
  wire h_u_cla32_and1019_y0;
  wire h_u_cla32_and1020_y0;
  wire h_u_cla32_and1021_y0;
  wire h_u_cla32_and1022_y0;
  wire h_u_cla32_and1023_y0;
  wire h_u_cla32_and1024_y0;
  wire h_u_cla32_and1025_y0;
  wire h_u_cla32_and1026_y0;
  wire h_u_cla32_and1027_y0;
  wire h_u_cla32_and1028_y0;
  wire h_u_cla32_and1029_y0;
  wire h_u_cla32_and1030_y0;
  wire h_u_cla32_and1031_y0;
  wire h_u_cla32_and1032_y0;
  wire h_u_cla32_and1033_y0;
  wire h_u_cla32_and1034_y0;
  wire h_u_cla32_and1035_y0;
  wire h_u_cla32_and1036_y0;
  wire h_u_cla32_and1037_y0;
  wire h_u_cla32_and1038_y0;
  wire h_u_cla32_and1039_y0;
  wire h_u_cla32_and1040_y0;
  wire h_u_cla32_and1041_y0;
  wire h_u_cla32_and1042_y0;
  wire h_u_cla32_and1043_y0;
  wire h_u_cla32_and1044_y0;
  wire h_u_cla32_and1045_y0;
  wire h_u_cla32_and1046_y0;
  wire h_u_cla32_and1047_y0;
  wire h_u_cla32_and1048_y0;
  wire h_u_cla32_and1049_y0;
  wire h_u_cla32_and1050_y0;
  wire h_u_cla32_and1051_y0;
  wire h_u_cla32_and1052_y0;
  wire h_u_cla32_and1053_y0;
  wire h_u_cla32_and1054_y0;
  wire h_u_cla32_and1055_y0;
  wire h_u_cla32_and1056_y0;
  wire h_u_cla32_and1057_y0;
  wire h_u_cla32_and1058_y0;
  wire h_u_cla32_and1059_y0;
  wire h_u_cla32_and1060_y0;
  wire h_u_cla32_and1061_y0;
  wire h_u_cla32_and1062_y0;
  wire h_u_cla32_and1063_y0;
  wire h_u_cla32_and1064_y0;
  wire h_u_cla32_and1065_y0;
  wire h_u_cla32_and1066_y0;
  wire h_u_cla32_and1067_y0;
  wire h_u_cla32_and1068_y0;
  wire h_u_cla32_and1069_y0;
  wire h_u_cla32_and1070_y0;
  wire h_u_cla32_and1071_y0;
  wire h_u_cla32_and1072_y0;
  wire h_u_cla32_and1073_y0;
  wire h_u_cla32_and1074_y0;
  wire h_u_cla32_and1075_y0;
  wire h_u_cla32_and1076_y0;
  wire h_u_cla32_and1077_y0;
  wire h_u_cla32_and1078_y0;
  wire h_u_cla32_and1079_y0;
  wire h_u_cla32_and1080_y0;
  wire h_u_cla32_and1081_y0;
  wire h_u_cla32_and1082_y0;
  wire h_u_cla32_and1083_y0;
  wire h_u_cla32_and1084_y0;
  wire h_u_cla32_and1085_y0;
  wire h_u_cla32_and1086_y0;
  wire h_u_cla32_and1087_y0;
  wire h_u_cla32_and1088_y0;
  wire h_u_cla32_and1089_y0;
  wire h_u_cla32_and1090_y0;
  wire h_u_cla32_and1091_y0;
  wire h_u_cla32_and1092_y0;
  wire h_u_cla32_and1093_y0;
  wire h_u_cla32_and1094_y0;
  wire h_u_cla32_and1095_y0;
  wire h_u_cla32_and1096_y0;
  wire h_u_cla32_and1097_y0;
  wire h_u_cla32_and1098_y0;
  wire h_u_cla32_and1099_y0;
  wire h_u_cla32_and1100_y0;
  wire h_u_cla32_and1101_y0;
  wire h_u_cla32_and1102_y0;
  wire h_u_cla32_and1103_y0;
  wire h_u_cla32_and1104_y0;
  wire h_u_cla32_and1105_y0;
  wire h_u_cla32_and1106_y0;
  wire h_u_cla32_and1107_y0;
  wire h_u_cla32_and1108_y0;
  wire h_u_cla32_and1109_y0;
  wire h_u_cla32_and1110_y0;
  wire h_u_cla32_and1111_y0;
  wire h_u_cla32_and1112_y0;
  wire h_u_cla32_and1113_y0;
  wire h_u_cla32_and1114_y0;
  wire h_u_cla32_and1115_y0;
  wire h_u_cla32_and1116_y0;
  wire h_u_cla32_and1117_y0;
  wire h_u_cla32_and1118_y0;
  wire h_u_cla32_and1119_y0;
  wire h_u_cla32_and1120_y0;
  wire h_u_cla32_and1121_y0;
  wire h_u_cla32_and1122_y0;
  wire h_u_cla32_and1123_y0;
  wire h_u_cla32_and1124_y0;
  wire h_u_cla32_and1125_y0;
  wire h_u_cla32_and1126_y0;
  wire h_u_cla32_and1127_y0;
  wire h_u_cla32_and1128_y0;
  wire h_u_cla32_and1129_y0;
  wire h_u_cla32_and1130_y0;
  wire h_u_cla32_and1131_y0;
  wire h_u_cla32_and1132_y0;
  wire h_u_cla32_and1133_y0;
  wire h_u_cla32_and1134_y0;
  wire h_u_cla32_and1135_y0;
  wire h_u_cla32_and1136_y0;
  wire h_u_cla32_and1137_y0;
  wire h_u_cla32_and1138_y0;
  wire h_u_cla32_and1139_y0;
  wire h_u_cla32_and1140_y0;
  wire h_u_cla32_and1141_y0;
  wire h_u_cla32_and1142_y0;
  wire h_u_cla32_and1143_y0;
  wire h_u_cla32_and1144_y0;
  wire h_u_cla32_and1145_y0;
  wire h_u_cla32_and1146_y0;
  wire h_u_cla32_and1147_y0;
  wire h_u_cla32_and1148_y0;
  wire h_u_cla32_and1149_y0;
  wire h_u_cla32_and1150_y0;
  wire h_u_cla32_and1151_y0;
  wire h_u_cla32_and1152_y0;
  wire h_u_cla32_and1153_y0;
  wire h_u_cla32_and1154_y0;
  wire h_u_cla32_and1155_y0;
  wire h_u_cla32_and1156_y0;
  wire h_u_cla32_and1157_y0;
  wire h_u_cla32_and1158_y0;
  wire h_u_cla32_and1159_y0;
  wire h_u_cla32_and1160_y0;
  wire h_u_cla32_and1161_y0;
  wire h_u_cla32_and1162_y0;
  wire h_u_cla32_and1163_y0;
  wire h_u_cla32_and1164_y0;
  wire h_u_cla32_and1165_y0;
  wire h_u_cla32_and1166_y0;
  wire h_u_cla32_and1167_y0;
  wire h_u_cla32_and1168_y0;
  wire h_u_cla32_and1169_y0;
  wire h_u_cla32_and1170_y0;
  wire h_u_cla32_and1171_y0;
  wire h_u_cla32_and1172_y0;
  wire h_u_cla32_and1173_y0;
  wire h_u_cla32_and1174_y0;
  wire h_u_cla32_and1175_y0;
  wire h_u_cla32_and1176_y0;
  wire h_u_cla32_and1177_y0;
  wire h_u_cla32_and1178_y0;
  wire h_u_cla32_and1179_y0;
  wire h_u_cla32_and1180_y0;
  wire h_u_cla32_and1181_y0;
  wire h_u_cla32_and1182_y0;
  wire h_u_cla32_and1183_y0;
  wire h_u_cla32_and1184_y0;
  wire h_u_cla32_and1185_y0;
  wire h_u_cla32_and1186_y0;
  wire h_u_cla32_and1187_y0;
  wire h_u_cla32_and1188_y0;
  wire h_u_cla32_and1189_y0;
  wire h_u_cla32_and1190_y0;
  wire h_u_cla32_and1191_y0;
  wire h_u_cla32_and1192_y0;
  wire h_u_cla32_and1193_y0;
  wire h_u_cla32_and1194_y0;
  wire h_u_cla32_and1195_y0;
  wire h_u_cla32_and1196_y0;
  wire h_u_cla32_and1197_y0;
  wire h_u_cla32_and1198_y0;
  wire h_u_cla32_and1199_y0;
  wire h_u_cla32_and1200_y0;
  wire h_u_cla32_and1201_y0;
  wire h_u_cla32_and1202_y0;
  wire h_u_cla32_and1203_y0;
  wire h_u_cla32_and1204_y0;
  wire h_u_cla32_and1205_y0;
  wire h_u_cla32_and1206_y0;
  wire h_u_cla32_and1207_y0;
  wire h_u_cla32_and1208_y0;
  wire h_u_cla32_and1209_y0;
  wire h_u_cla32_and1210_y0;
  wire h_u_cla32_and1211_y0;
  wire h_u_cla32_and1212_y0;
  wire h_u_cla32_and1213_y0;
  wire h_u_cla32_and1214_y0;
  wire h_u_cla32_and1215_y0;
  wire h_u_cla32_and1216_y0;
  wire h_u_cla32_and1217_y0;
  wire h_u_cla32_and1218_y0;
  wire h_u_cla32_and1219_y0;
  wire h_u_cla32_and1220_y0;
  wire h_u_cla32_and1221_y0;
  wire h_u_cla32_and1222_y0;
  wire h_u_cla32_and1223_y0;
  wire h_u_cla32_and1224_y0;
  wire h_u_cla32_and1225_y0;
  wire h_u_cla32_and1226_y0;
  wire h_u_cla32_and1227_y0;
  wire h_u_cla32_and1228_y0;
  wire h_u_cla32_and1229_y0;
  wire h_u_cla32_and1230_y0;
  wire h_u_cla32_and1231_y0;
  wire h_u_cla32_and1232_y0;
  wire h_u_cla32_and1233_y0;
  wire h_u_cla32_and1234_y0;
  wire h_u_cla32_and1235_y0;
  wire h_u_cla32_and1236_y0;
  wire h_u_cla32_and1237_y0;
  wire h_u_cla32_and1238_y0;
  wire h_u_cla32_and1239_y0;
  wire h_u_cla32_or105_y0;
  wire h_u_cla32_or106_y0;
  wire h_u_cla32_or107_y0;
  wire h_u_cla32_or108_y0;
  wire h_u_cla32_or109_y0;
  wire h_u_cla32_or110_y0;
  wire h_u_cla32_or111_y0;
  wire h_u_cla32_or112_y0;
  wire h_u_cla32_or113_y0;
  wire h_u_cla32_or114_y0;
  wire h_u_cla32_or115_y0;
  wire h_u_cla32_or116_y0;
  wire h_u_cla32_or117_y0;
  wire h_u_cla32_or118_y0;
  wire h_u_cla32_or119_y0;
  wire h_u_cla32_pg_logic15_y0;
  wire h_u_cla32_pg_logic15_y1;
  wire h_u_cla32_pg_logic15_y2;
  wire h_u_cla32_xor15_y0;
  wire h_u_cla32_and1240_y0;
  wire h_u_cla32_and1241_y0;
  wire h_u_cla32_and1242_y0;
  wire h_u_cla32_and1243_y0;
  wire h_u_cla32_and1244_y0;
  wire h_u_cla32_and1245_y0;
  wire h_u_cla32_and1246_y0;
  wire h_u_cla32_and1247_y0;
  wire h_u_cla32_and1248_y0;
  wire h_u_cla32_and1249_y0;
  wire h_u_cla32_and1250_y0;
  wire h_u_cla32_and1251_y0;
  wire h_u_cla32_and1252_y0;
  wire h_u_cla32_and1253_y0;
  wire h_u_cla32_and1254_y0;
  wire h_u_cla32_and1255_y0;
  wire h_u_cla32_and1256_y0;
  wire h_u_cla32_and1257_y0;
  wire h_u_cla32_and1258_y0;
  wire h_u_cla32_and1259_y0;
  wire h_u_cla32_and1260_y0;
  wire h_u_cla32_and1261_y0;
  wire h_u_cla32_and1262_y0;
  wire h_u_cla32_and1263_y0;
  wire h_u_cla32_and1264_y0;
  wire h_u_cla32_and1265_y0;
  wire h_u_cla32_and1266_y0;
  wire h_u_cla32_and1267_y0;
  wire h_u_cla32_and1268_y0;
  wire h_u_cla32_and1269_y0;
  wire h_u_cla32_and1270_y0;
  wire h_u_cla32_and1271_y0;
  wire h_u_cla32_and1272_y0;
  wire h_u_cla32_and1273_y0;
  wire h_u_cla32_and1274_y0;
  wire h_u_cla32_and1275_y0;
  wire h_u_cla32_and1276_y0;
  wire h_u_cla32_and1277_y0;
  wire h_u_cla32_and1278_y0;
  wire h_u_cla32_and1279_y0;
  wire h_u_cla32_and1280_y0;
  wire h_u_cla32_and1281_y0;
  wire h_u_cla32_and1282_y0;
  wire h_u_cla32_and1283_y0;
  wire h_u_cla32_and1284_y0;
  wire h_u_cla32_and1285_y0;
  wire h_u_cla32_and1286_y0;
  wire h_u_cla32_and1287_y0;
  wire h_u_cla32_and1288_y0;
  wire h_u_cla32_and1289_y0;
  wire h_u_cla32_and1290_y0;
  wire h_u_cla32_and1291_y0;
  wire h_u_cla32_and1292_y0;
  wire h_u_cla32_and1293_y0;
  wire h_u_cla32_and1294_y0;
  wire h_u_cla32_and1295_y0;
  wire h_u_cla32_and1296_y0;
  wire h_u_cla32_and1297_y0;
  wire h_u_cla32_and1298_y0;
  wire h_u_cla32_and1299_y0;
  wire h_u_cla32_and1300_y0;
  wire h_u_cla32_and1301_y0;
  wire h_u_cla32_and1302_y0;
  wire h_u_cla32_and1303_y0;
  wire h_u_cla32_and1304_y0;
  wire h_u_cla32_and1305_y0;
  wire h_u_cla32_and1306_y0;
  wire h_u_cla32_and1307_y0;
  wire h_u_cla32_and1308_y0;
  wire h_u_cla32_and1309_y0;
  wire h_u_cla32_and1310_y0;
  wire h_u_cla32_and1311_y0;
  wire h_u_cla32_and1312_y0;
  wire h_u_cla32_and1313_y0;
  wire h_u_cla32_and1314_y0;
  wire h_u_cla32_and1315_y0;
  wire h_u_cla32_and1316_y0;
  wire h_u_cla32_and1317_y0;
  wire h_u_cla32_and1318_y0;
  wire h_u_cla32_and1319_y0;
  wire h_u_cla32_and1320_y0;
  wire h_u_cla32_and1321_y0;
  wire h_u_cla32_and1322_y0;
  wire h_u_cla32_and1323_y0;
  wire h_u_cla32_and1324_y0;
  wire h_u_cla32_and1325_y0;
  wire h_u_cla32_and1326_y0;
  wire h_u_cla32_and1327_y0;
  wire h_u_cla32_and1328_y0;
  wire h_u_cla32_and1329_y0;
  wire h_u_cla32_and1330_y0;
  wire h_u_cla32_and1331_y0;
  wire h_u_cla32_and1332_y0;
  wire h_u_cla32_and1333_y0;
  wire h_u_cla32_and1334_y0;
  wire h_u_cla32_and1335_y0;
  wire h_u_cla32_and1336_y0;
  wire h_u_cla32_and1337_y0;
  wire h_u_cla32_and1338_y0;
  wire h_u_cla32_and1339_y0;
  wire h_u_cla32_and1340_y0;
  wire h_u_cla32_and1341_y0;
  wire h_u_cla32_and1342_y0;
  wire h_u_cla32_and1343_y0;
  wire h_u_cla32_and1344_y0;
  wire h_u_cla32_and1345_y0;
  wire h_u_cla32_and1346_y0;
  wire h_u_cla32_and1347_y0;
  wire h_u_cla32_and1348_y0;
  wire h_u_cla32_and1349_y0;
  wire h_u_cla32_and1350_y0;
  wire h_u_cla32_and1351_y0;
  wire h_u_cla32_and1352_y0;
  wire h_u_cla32_and1353_y0;
  wire h_u_cla32_and1354_y0;
  wire h_u_cla32_and1355_y0;
  wire h_u_cla32_and1356_y0;
  wire h_u_cla32_and1357_y0;
  wire h_u_cla32_and1358_y0;
  wire h_u_cla32_and1359_y0;
  wire h_u_cla32_and1360_y0;
  wire h_u_cla32_and1361_y0;
  wire h_u_cla32_and1362_y0;
  wire h_u_cla32_and1363_y0;
  wire h_u_cla32_and1364_y0;
  wire h_u_cla32_and1365_y0;
  wire h_u_cla32_and1366_y0;
  wire h_u_cla32_and1367_y0;
  wire h_u_cla32_and1368_y0;
  wire h_u_cla32_and1369_y0;
  wire h_u_cla32_and1370_y0;
  wire h_u_cla32_and1371_y0;
  wire h_u_cla32_and1372_y0;
  wire h_u_cla32_and1373_y0;
  wire h_u_cla32_and1374_y0;
  wire h_u_cla32_and1375_y0;
  wire h_u_cla32_and1376_y0;
  wire h_u_cla32_and1377_y0;
  wire h_u_cla32_and1378_y0;
  wire h_u_cla32_and1379_y0;
  wire h_u_cla32_and1380_y0;
  wire h_u_cla32_and1381_y0;
  wire h_u_cla32_and1382_y0;
  wire h_u_cla32_and1383_y0;
  wire h_u_cla32_and1384_y0;
  wire h_u_cla32_and1385_y0;
  wire h_u_cla32_and1386_y0;
  wire h_u_cla32_and1387_y0;
  wire h_u_cla32_and1388_y0;
  wire h_u_cla32_and1389_y0;
  wire h_u_cla32_and1390_y0;
  wire h_u_cla32_and1391_y0;
  wire h_u_cla32_and1392_y0;
  wire h_u_cla32_and1393_y0;
  wire h_u_cla32_and1394_y0;
  wire h_u_cla32_and1395_y0;
  wire h_u_cla32_and1396_y0;
  wire h_u_cla32_and1397_y0;
  wire h_u_cla32_and1398_y0;
  wire h_u_cla32_and1399_y0;
  wire h_u_cla32_and1400_y0;
  wire h_u_cla32_and1401_y0;
  wire h_u_cla32_and1402_y0;
  wire h_u_cla32_and1403_y0;
  wire h_u_cla32_and1404_y0;
  wire h_u_cla32_and1405_y0;
  wire h_u_cla32_and1406_y0;
  wire h_u_cla32_and1407_y0;
  wire h_u_cla32_and1408_y0;
  wire h_u_cla32_and1409_y0;
  wire h_u_cla32_and1410_y0;
  wire h_u_cla32_and1411_y0;
  wire h_u_cla32_and1412_y0;
  wire h_u_cla32_and1413_y0;
  wire h_u_cla32_and1414_y0;
  wire h_u_cla32_and1415_y0;
  wire h_u_cla32_and1416_y0;
  wire h_u_cla32_and1417_y0;
  wire h_u_cla32_and1418_y0;
  wire h_u_cla32_and1419_y0;
  wire h_u_cla32_and1420_y0;
  wire h_u_cla32_and1421_y0;
  wire h_u_cla32_and1422_y0;
  wire h_u_cla32_and1423_y0;
  wire h_u_cla32_and1424_y0;
  wire h_u_cla32_and1425_y0;
  wire h_u_cla32_and1426_y0;
  wire h_u_cla32_and1427_y0;
  wire h_u_cla32_and1428_y0;
  wire h_u_cla32_and1429_y0;
  wire h_u_cla32_and1430_y0;
  wire h_u_cla32_and1431_y0;
  wire h_u_cla32_and1432_y0;
  wire h_u_cla32_and1433_y0;
  wire h_u_cla32_and1434_y0;
  wire h_u_cla32_and1435_y0;
  wire h_u_cla32_and1436_y0;
  wire h_u_cla32_and1437_y0;
  wire h_u_cla32_and1438_y0;
  wire h_u_cla32_and1439_y0;
  wire h_u_cla32_and1440_y0;
  wire h_u_cla32_and1441_y0;
  wire h_u_cla32_and1442_y0;
  wire h_u_cla32_and1443_y0;
  wire h_u_cla32_and1444_y0;
  wire h_u_cla32_and1445_y0;
  wire h_u_cla32_and1446_y0;
  wire h_u_cla32_and1447_y0;
  wire h_u_cla32_and1448_y0;
  wire h_u_cla32_and1449_y0;
  wire h_u_cla32_and1450_y0;
  wire h_u_cla32_and1451_y0;
  wire h_u_cla32_and1452_y0;
  wire h_u_cla32_and1453_y0;
  wire h_u_cla32_and1454_y0;
  wire h_u_cla32_and1455_y0;
  wire h_u_cla32_and1456_y0;
  wire h_u_cla32_and1457_y0;
  wire h_u_cla32_and1458_y0;
  wire h_u_cla32_and1459_y0;
  wire h_u_cla32_and1460_y0;
  wire h_u_cla32_and1461_y0;
  wire h_u_cla32_and1462_y0;
  wire h_u_cla32_and1463_y0;
  wire h_u_cla32_and1464_y0;
  wire h_u_cla32_and1465_y0;
  wire h_u_cla32_and1466_y0;
  wire h_u_cla32_and1467_y0;
  wire h_u_cla32_and1468_y0;
  wire h_u_cla32_and1469_y0;
  wire h_u_cla32_and1470_y0;
  wire h_u_cla32_and1471_y0;
  wire h_u_cla32_and1472_y0;
  wire h_u_cla32_and1473_y0;
  wire h_u_cla32_and1474_y0;
  wire h_u_cla32_and1475_y0;
  wire h_u_cla32_and1476_y0;
  wire h_u_cla32_and1477_y0;
  wire h_u_cla32_and1478_y0;
  wire h_u_cla32_and1479_y0;
  wire h_u_cla32_and1480_y0;
  wire h_u_cla32_and1481_y0;
  wire h_u_cla32_and1482_y0;
  wire h_u_cla32_and1483_y0;
  wire h_u_cla32_and1484_y0;
  wire h_u_cla32_and1485_y0;
  wire h_u_cla32_and1486_y0;
  wire h_u_cla32_and1487_y0;
  wire h_u_cla32_and1488_y0;
  wire h_u_cla32_and1489_y0;
  wire h_u_cla32_and1490_y0;
  wire h_u_cla32_and1491_y0;
  wire h_u_cla32_and1492_y0;
  wire h_u_cla32_and1493_y0;
  wire h_u_cla32_and1494_y0;
  wire h_u_cla32_and1495_y0;
  wire h_u_cla32_or120_y0;
  wire h_u_cla32_or121_y0;
  wire h_u_cla32_or122_y0;
  wire h_u_cla32_or123_y0;
  wire h_u_cla32_or124_y0;
  wire h_u_cla32_or125_y0;
  wire h_u_cla32_or126_y0;
  wire h_u_cla32_or127_y0;
  wire h_u_cla32_or128_y0;
  wire h_u_cla32_or129_y0;
  wire h_u_cla32_or130_y0;
  wire h_u_cla32_or131_y0;
  wire h_u_cla32_or132_y0;
  wire h_u_cla32_or133_y0;
  wire h_u_cla32_or134_y0;
  wire h_u_cla32_or135_y0;
  wire h_u_cla32_pg_logic16_y0;
  wire h_u_cla32_pg_logic16_y1;
  wire h_u_cla32_pg_logic16_y2;
  wire h_u_cla32_xor16_y0;
  wire h_u_cla32_and1496_y0;
  wire h_u_cla32_and1497_y0;
  wire h_u_cla32_and1498_y0;
  wire h_u_cla32_and1499_y0;
  wire h_u_cla32_and1500_y0;
  wire h_u_cla32_and1501_y0;
  wire h_u_cla32_and1502_y0;
  wire h_u_cla32_and1503_y0;
  wire h_u_cla32_and1504_y0;
  wire h_u_cla32_and1505_y0;
  wire h_u_cla32_and1506_y0;
  wire h_u_cla32_and1507_y0;
  wire h_u_cla32_and1508_y0;
  wire h_u_cla32_and1509_y0;
  wire h_u_cla32_and1510_y0;
  wire h_u_cla32_and1511_y0;
  wire h_u_cla32_and1512_y0;
  wire h_u_cla32_and1513_y0;
  wire h_u_cla32_and1514_y0;
  wire h_u_cla32_and1515_y0;
  wire h_u_cla32_and1516_y0;
  wire h_u_cla32_and1517_y0;
  wire h_u_cla32_and1518_y0;
  wire h_u_cla32_and1519_y0;
  wire h_u_cla32_and1520_y0;
  wire h_u_cla32_and1521_y0;
  wire h_u_cla32_and1522_y0;
  wire h_u_cla32_and1523_y0;
  wire h_u_cla32_and1524_y0;
  wire h_u_cla32_and1525_y0;
  wire h_u_cla32_and1526_y0;
  wire h_u_cla32_and1527_y0;
  wire h_u_cla32_and1528_y0;
  wire h_u_cla32_and1529_y0;
  wire h_u_cla32_and1530_y0;
  wire h_u_cla32_and1531_y0;
  wire h_u_cla32_and1532_y0;
  wire h_u_cla32_and1533_y0;
  wire h_u_cla32_and1534_y0;
  wire h_u_cla32_and1535_y0;
  wire h_u_cla32_and1536_y0;
  wire h_u_cla32_and1537_y0;
  wire h_u_cla32_and1538_y0;
  wire h_u_cla32_and1539_y0;
  wire h_u_cla32_and1540_y0;
  wire h_u_cla32_and1541_y0;
  wire h_u_cla32_and1542_y0;
  wire h_u_cla32_and1543_y0;
  wire h_u_cla32_and1544_y0;
  wire h_u_cla32_and1545_y0;
  wire h_u_cla32_and1546_y0;
  wire h_u_cla32_and1547_y0;
  wire h_u_cla32_and1548_y0;
  wire h_u_cla32_and1549_y0;
  wire h_u_cla32_and1550_y0;
  wire h_u_cla32_and1551_y0;
  wire h_u_cla32_and1552_y0;
  wire h_u_cla32_and1553_y0;
  wire h_u_cla32_and1554_y0;
  wire h_u_cla32_and1555_y0;
  wire h_u_cla32_and1556_y0;
  wire h_u_cla32_and1557_y0;
  wire h_u_cla32_and1558_y0;
  wire h_u_cla32_and1559_y0;
  wire h_u_cla32_and1560_y0;
  wire h_u_cla32_and1561_y0;
  wire h_u_cla32_and1562_y0;
  wire h_u_cla32_and1563_y0;
  wire h_u_cla32_and1564_y0;
  wire h_u_cla32_and1565_y0;
  wire h_u_cla32_and1566_y0;
  wire h_u_cla32_and1567_y0;
  wire h_u_cla32_and1568_y0;
  wire h_u_cla32_and1569_y0;
  wire h_u_cla32_and1570_y0;
  wire h_u_cla32_and1571_y0;
  wire h_u_cla32_and1572_y0;
  wire h_u_cla32_and1573_y0;
  wire h_u_cla32_and1574_y0;
  wire h_u_cla32_and1575_y0;
  wire h_u_cla32_and1576_y0;
  wire h_u_cla32_and1577_y0;
  wire h_u_cla32_and1578_y0;
  wire h_u_cla32_and1579_y0;
  wire h_u_cla32_and1580_y0;
  wire h_u_cla32_and1581_y0;
  wire h_u_cla32_and1582_y0;
  wire h_u_cla32_and1583_y0;
  wire h_u_cla32_and1584_y0;
  wire h_u_cla32_and1585_y0;
  wire h_u_cla32_and1586_y0;
  wire h_u_cla32_and1587_y0;
  wire h_u_cla32_and1588_y0;
  wire h_u_cla32_and1589_y0;
  wire h_u_cla32_and1590_y0;
  wire h_u_cla32_and1591_y0;
  wire h_u_cla32_and1592_y0;
  wire h_u_cla32_and1593_y0;
  wire h_u_cla32_and1594_y0;
  wire h_u_cla32_and1595_y0;
  wire h_u_cla32_and1596_y0;
  wire h_u_cla32_and1597_y0;
  wire h_u_cla32_and1598_y0;
  wire h_u_cla32_and1599_y0;
  wire h_u_cla32_and1600_y0;
  wire h_u_cla32_and1601_y0;
  wire h_u_cla32_and1602_y0;
  wire h_u_cla32_and1603_y0;
  wire h_u_cla32_and1604_y0;
  wire h_u_cla32_and1605_y0;
  wire h_u_cla32_and1606_y0;
  wire h_u_cla32_and1607_y0;
  wire h_u_cla32_and1608_y0;
  wire h_u_cla32_and1609_y0;
  wire h_u_cla32_and1610_y0;
  wire h_u_cla32_and1611_y0;
  wire h_u_cla32_and1612_y0;
  wire h_u_cla32_and1613_y0;
  wire h_u_cla32_and1614_y0;
  wire h_u_cla32_and1615_y0;
  wire h_u_cla32_and1616_y0;
  wire h_u_cla32_and1617_y0;
  wire h_u_cla32_and1618_y0;
  wire h_u_cla32_and1619_y0;
  wire h_u_cla32_and1620_y0;
  wire h_u_cla32_and1621_y0;
  wire h_u_cla32_and1622_y0;
  wire h_u_cla32_and1623_y0;
  wire h_u_cla32_and1624_y0;
  wire h_u_cla32_and1625_y0;
  wire h_u_cla32_and1626_y0;
  wire h_u_cla32_and1627_y0;
  wire h_u_cla32_and1628_y0;
  wire h_u_cla32_and1629_y0;
  wire h_u_cla32_and1630_y0;
  wire h_u_cla32_and1631_y0;
  wire h_u_cla32_and1632_y0;
  wire h_u_cla32_and1633_y0;
  wire h_u_cla32_and1634_y0;
  wire h_u_cla32_and1635_y0;
  wire h_u_cla32_and1636_y0;
  wire h_u_cla32_and1637_y0;
  wire h_u_cla32_and1638_y0;
  wire h_u_cla32_and1639_y0;
  wire h_u_cla32_and1640_y0;
  wire h_u_cla32_and1641_y0;
  wire h_u_cla32_and1642_y0;
  wire h_u_cla32_and1643_y0;
  wire h_u_cla32_and1644_y0;
  wire h_u_cla32_and1645_y0;
  wire h_u_cla32_and1646_y0;
  wire h_u_cla32_and1647_y0;
  wire h_u_cla32_and1648_y0;
  wire h_u_cla32_and1649_y0;
  wire h_u_cla32_and1650_y0;
  wire h_u_cla32_and1651_y0;
  wire h_u_cla32_and1652_y0;
  wire h_u_cla32_and1653_y0;
  wire h_u_cla32_and1654_y0;
  wire h_u_cla32_and1655_y0;
  wire h_u_cla32_and1656_y0;
  wire h_u_cla32_and1657_y0;
  wire h_u_cla32_and1658_y0;
  wire h_u_cla32_and1659_y0;
  wire h_u_cla32_and1660_y0;
  wire h_u_cla32_and1661_y0;
  wire h_u_cla32_and1662_y0;
  wire h_u_cla32_and1663_y0;
  wire h_u_cla32_and1664_y0;
  wire h_u_cla32_and1665_y0;
  wire h_u_cla32_and1666_y0;
  wire h_u_cla32_and1667_y0;
  wire h_u_cla32_and1668_y0;
  wire h_u_cla32_and1669_y0;
  wire h_u_cla32_and1670_y0;
  wire h_u_cla32_and1671_y0;
  wire h_u_cla32_and1672_y0;
  wire h_u_cla32_and1673_y0;
  wire h_u_cla32_and1674_y0;
  wire h_u_cla32_and1675_y0;
  wire h_u_cla32_and1676_y0;
  wire h_u_cla32_and1677_y0;
  wire h_u_cla32_and1678_y0;
  wire h_u_cla32_and1679_y0;
  wire h_u_cla32_and1680_y0;
  wire h_u_cla32_and1681_y0;
  wire h_u_cla32_and1682_y0;
  wire h_u_cla32_and1683_y0;
  wire h_u_cla32_and1684_y0;
  wire h_u_cla32_and1685_y0;
  wire h_u_cla32_and1686_y0;
  wire h_u_cla32_and1687_y0;
  wire h_u_cla32_and1688_y0;
  wire h_u_cla32_and1689_y0;
  wire h_u_cla32_and1690_y0;
  wire h_u_cla32_and1691_y0;
  wire h_u_cla32_and1692_y0;
  wire h_u_cla32_and1693_y0;
  wire h_u_cla32_and1694_y0;
  wire h_u_cla32_and1695_y0;
  wire h_u_cla32_and1696_y0;
  wire h_u_cla32_and1697_y0;
  wire h_u_cla32_and1698_y0;
  wire h_u_cla32_and1699_y0;
  wire h_u_cla32_and1700_y0;
  wire h_u_cla32_and1701_y0;
  wire h_u_cla32_and1702_y0;
  wire h_u_cla32_and1703_y0;
  wire h_u_cla32_and1704_y0;
  wire h_u_cla32_and1705_y0;
  wire h_u_cla32_and1706_y0;
  wire h_u_cla32_and1707_y0;
  wire h_u_cla32_and1708_y0;
  wire h_u_cla32_and1709_y0;
  wire h_u_cla32_and1710_y0;
  wire h_u_cla32_and1711_y0;
  wire h_u_cla32_and1712_y0;
  wire h_u_cla32_and1713_y0;
  wire h_u_cla32_and1714_y0;
  wire h_u_cla32_and1715_y0;
  wire h_u_cla32_and1716_y0;
  wire h_u_cla32_and1717_y0;
  wire h_u_cla32_and1718_y0;
  wire h_u_cla32_and1719_y0;
  wire h_u_cla32_and1720_y0;
  wire h_u_cla32_and1721_y0;
  wire h_u_cla32_and1722_y0;
  wire h_u_cla32_and1723_y0;
  wire h_u_cla32_and1724_y0;
  wire h_u_cla32_and1725_y0;
  wire h_u_cla32_and1726_y0;
  wire h_u_cla32_and1727_y0;
  wire h_u_cla32_and1728_y0;
  wire h_u_cla32_and1729_y0;
  wire h_u_cla32_and1730_y0;
  wire h_u_cla32_and1731_y0;
  wire h_u_cla32_and1732_y0;
  wire h_u_cla32_and1733_y0;
  wire h_u_cla32_and1734_y0;
  wire h_u_cla32_and1735_y0;
  wire h_u_cla32_and1736_y0;
  wire h_u_cla32_and1737_y0;
  wire h_u_cla32_and1738_y0;
  wire h_u_cla32_and1739_y0;
  wire h_u_cla32_and1740_y0;
  wire h_u_cla32_and1741_y0;
  wire h_u_cla32_and1742_y0;
  wire h_u_cla32_and1743_y0;
  wire h_u_cla32_and1744_y0;
  wire h_u_cla32_and1745_y0;
  wire h_u_cla32_and1746_y0;
  wire h_u_cla32_and1747_y0;
  wire h_u_cla32_and1748_y0;
  wire h_u_cla32_and1749_y0;
  wire h_u_cla32_and1750_y0;
  wire h_u_cla32_and1751_y0;
  wire h_u_cla32_and1752_y0;
  wire h_u_cla32_and1753_y0;
  wire h_u_cla32_and1754_y0;
  wire h_u_cla32_and1755_y0;
  wire h_u_cla32_and1756_y0;
  wire h_u_cla32_and1757_y0;
  wire h_u_cla32_and1758_y0;
  wire h_u_cla32_and1759_y0;
  wire h_u_cla32_and1760_y0;
  wire h_u_cla32_and1761_y0;
  wire h_u_cla32_and1762_y0;
  wire h_u_cla32_and1763_y0;
  wire h_u_cla32_and1764_y0;
  wire h_u_cla32_and1765_y0;
  wire h_u_cla32_and1766_y0;
  wire h_u_cla32_and1767_y0;
  wire h_u_cla32_and1768_y0;
  wire h_u_cla32_and1769_y0;
  wire h_u_cla32_and1770_y0;
  wire h_u_cla32_and1771_y0;
  wire h_u_cla32_and1772_y0;
  wire h_u_cla32_and1773_y0;
  wire h_u_cla32_and1774_y0;
  wire h_u_cla32_and1775_y0;
  wire h_u_cla32_and1776_y0;
  wire h_u_cla32_and1777_y0;
  wire h_u_cla32_and1778_y0;
  wire h_u_cla32_and1779_y0;
  wire h_u_cla32_and1780_y0;
  wire h_u_cla32_and1781_y0;
  wire h_u_cla32_and1782_y0;
  wire h_u_cla32_and1783_y0;
  wire h_u_cla32_and1784_y0;
  wire h_u_cla32_or136_y0;
  wire h_u_cla32_or137_y0;
  wire h_u_cla32_or138_y0;
  wire h_u_cla32_or139_y0;
  wire h_u_cla32_or140_y0;
  wire h_u_cla32_or141_y0;
  wire h_u_cla32_or142_y0;
  wire h_u_cla32_or143_y0;
  wire h_u_cla32_or144_y0;
  wire h_u_cla32_or145_y0;
  wire h_u_cla32_or146_y0;
  wire h_u_cla32_or147_y0;
  wire h_u_cla32_or148_y0;
  wire h_u_cla32_or149_y0;
  wire h_u_cla32_or150_y0;
  wire h_u_cla32_or151_y0;
  wire h_u_cla32_or152_y0;
  wire h_u_cla32_pg_logic17_y0;
  wire h_u_cla32_pg_logic17_y1;
  wire h_u_cla32_pg_logic17_y2;
  wire h_u_cla32_xor17_y0;
  wire h_u_cla32_and1785_y0;
  wire h_u_cla32_and1786_y0;
  wire h_u_cla32_and1787_y0;
  wire h_u_cla32_and1788_y0;
  wire h_u_cla32_and1789_y0;
  wire h_u_cla32_and1790_y0;
  wire h_u_cla32_and1791_y0;
  wire h_u_cla32_and1792_y0;
  wire h_u_cla32_and1793_y0;
  wire h_u_cla32_and1794_y0;
  wire h_u_cla32_and1795_y0;
  wire h_u_cla32_and1796_y0;
  wire h_u_cla32_and1797_y0;
  wire h_u_cla32_and1798_y0;
  wire h_u_cla32_and1799_y0;
  wire h_u_cla32_and1800_y0;
  wire h_u_cla32_and1801_y0;
  wire h_u_cla32_and1802_y0;
  wire h_u_cla32_and1803_y0;
  wire h_u_cla32_and1804_y0;
  wire h_u_cla32_and1805_y0;
  wire h_u_cla32_and1806_y0;
  wire h_u_cla32_and1807_y0;
  wire h_u_cla32_and1808_y0;
  wire h_u_cla32_and1809_y0;
  wire h_u_cla32_and1810_y0;
  wire h_u_cla32_and1811_y0;
  wire h_u_cla32_and1812_y0;
  wire h_u_cla32_and1813_y0;
  wire h_u_cla32_and1814_y0;
  wire h_u_cla32_and1815_y0;
  wire h_u_cla32_and1816_y0;
  wire h_u_cla32_and1817_y0;
  wire h_u_cla32_and1818_y0;
  wire h_u_cla32_and1819_y0;
  wire h_u_cla32_and1820_y0;
  wire h_u_cla32_and1821_y0;
  wire h_u_cla32_and1822_y0;
  wire h_u_cla32_and1823_y0;
  wire h_u_cla32_and1824_y0;
  wire h_u_cla32_and1825_y0;
  wire h_u_cla32_and1826_y0;
  wire h_u_cla32_and1827_y0;
  wire h_u_cla32_and1828_y0;
  wire h_u_cla32_and1829_y0;
  wire h_u_cla32_and1830_y0;
  wire h_u_cla32_and1831_y0;
  wire h_u_cla32_and1832_y0;
  wire h_u_cla32_and1833_y0;
  wire h_u_cla32_and1834_y0;
  wire h_u_cla32_and1835_y0;
  wire h_u_cla32_and1836_y0;
  wire h_u_cla32_and1837_y0;
  wire h_u_cla32_and1838_y0;
  wire h_u_cla32_and1839_y0;
  wire h_u_cla32_and1840_y0;
  wire h_u_cla32_and1841_y0;
  wire h_u_cla32_and1842_y0;
  wire h_u_cla32_and1843_y0;
  wire h_u_cla32_and1844_y0;
  wire h_u_cla32_and1845_y0;
  wire h_u_cla32_and1846_y0;
  wire h_u_cla32_and1847_y0;
  wire h_u_cla32_and1848_y0;
  wire h_u_cla32_and1849_y0;
  wire h_u_cla32_and1850_y0;
  wire h_u_cla32_and1851_y0;
  wire h_u_cla32_and1852_y0;
  wire h_u_cla32_and1853_y0;
  wire h_u_cla32_and1854_y0;
  wire h_u_cla32_and1855_y0;
  wire h_u_cla32_and1856_y0;
  wire h_u_cla32_and1857_y0;
  wire h_u_cla32_and1858_y0;
  wire h_u_cla32_and1859_y0;
  wire h_u_cla32_and1860_y0;
  wire h_u_cla32_and1861_y0;
  wire h_u_cla32_and1862_y0;
  wire h_u_cla32_and1863_y0;
  wire h_u_cla32_and1864_y0;
  wire h_u_cla32_and1865_y0;
  wire h_u_cla32_and1866_y0;
  wire h_u_cla32_and1867_y0;
  wire h_u_cla32_and1868_y0;
  wire h_u_cla32_and1869_y0;
  wire h_u_cla32_and1870_y0;
  wire h_u_cla32_and1871_y0;
  wire h_u_cla32_and1872_y0;
  wire h_u_cla32_and1873_y0;
  wire h_u_cla32_and1874_y0;
  wire h_u_cla32_and1875_y0;
  wire h_u_cla32_and1876_y0;
  wire h_u_cla32_and1877_y0;
  wire h_u_cla32_and1878_y0;
  wire h_u_cla32_and1879_y0;
  wire h_u_cla32_and1880_y0;
  wire h_u_cla32_and1881_y0;
  wire h_u_cla32_and1882_y0;
  wire h_u_cla32_and1883_y0;
  wire h_u_cla32_and1884_y0;
  wire h_u_cla32_and1885_y0;
  wire h_u_cla32_and1886_y0;
  wire h_u_cla32_and1887_y0;
  wire h_u_cla32_and1888_y0;
  wire h_u_cla32_and1889_y0;
  wire h_u_cla32_and1890_y0;
  wire h_u_cla32_and1891_y0;
  wire h_u_cla32_and1892_y0;
  wire h_u_cla32_and1893_y0;
  wire h_u_cla32_and1894_y0;
  wire h_u_cla32_and1895_y0;
  wire h_u_cla32_and1896_y0;
  wire h_u_cla32_and1897_y0;
  wire h_u_cla32_and1898_y0;
  wire h_u_cla32_and1899_y0;
  wire h_u_cla32_and1900_y0;
  wire h_u_cla32_and1901_y0;
  wire h_u_cla32_and1902_y0;
  wire h_u_cla32_and1903_y0;
  wire h_u_cla32_and1904_y0;
  wire h_u_cla32_and1905_y0;
  wire h_u_cla32_and1906_y0;
  wire h_u_cla32_and1907_y0;
  wire h_u_cla32_and1908_y0;
  wire h_u_cla32_and1909_y0;
  wire h_u_cla32_and1910_y0;
  wire h_u_cla32_and1911_y0;
  wire h_u_cla32_and1912_y0;
  wire h_u_cla32_and1913_y0;
  wire h_u_cla32_and1914_y0;
  wire h_u_cla32_and1915_y0;
  wire h_u_cla32_and1916_y0;
  wire h_u_cla32_and1917_y0;
  wire h_u_cla32_and1918_y0;
  wire h_u_cla32_and1919_y0;
  wire h_u_cla32_and1920_y0;
  wire h_u_cla32_and1921_y0;
  wire h_u_cla32_and1922_y0;
  wire h_u_cla32_and1923_y0;
  wire h_u_cla32_and1924_y0;
  wire h_u_cla32_and1925_y0;
  wire h_u_cla32_and1926_y0;
  wire h_u_cla32_and1927_y0;
  wire h_u_cla32_and1928_y0;
  wire h_u_cla32_and1929_y0;
  wire h_u_cla32_and1930_y0;
  wire h_u_cla32_and1931_y0;
  wire h_u_cla32_and1932_y0;
  wire h_u_cla32_and1933_y0;
  wire h_u_cla32_and1934_y0;
  wire h_u_cla32_and1935_y0;
  wire h_u_cla32_and1936_y0;
  wire h_u_cla32_and1937_y0;
  wire h_u_cla32_and1938_y0;
  wire h_u_cla32_and1939_y0;
  wire h_u_cla32_and1940_y0;
  wire h_u_cla32_and1941_y0;
  wire h_u_cla32_and1942_y0;
  wire h_u_cla32_and1943_y0;
  wire h_u_cla32_and1944_y0;
  wire h_u_cla32_and1945_y0;
  wire h_u_cla32_and1946_y0;
  wire h_u_cla32_and1947_y0;
  wire h_u_cla32_and1948_y0;
  wire h_u_cla32_and1949_y0;
  wire h_u_cla32_and1950_y0;
  wire h_u_cla32_and1951_y0;
  wire h_u_cla32_and1952_y0;
  wire h_u_cla32_and1953_y0;
  wire h_u_cla32_and1954_y0;
  wire h_u_cla32_and1955_y0;
  wire h_u_cla32_and1956_y0;
  wire h_u_cla32_and1957_y0;
  wire h_u_cla32_and1958_y0;
  wire h_u_cla32_and1959_y0;
  wire h_u_cla32_and1960_y0;
  wire h_u_cla32_and1961_y0;
  wire h_u_cla32_and1962_y0;
  wire h_u_cla32_and1963_y0;
  wire h_u_cla32_and1964_y0;
  wire h_u_cla32_and1965_y0;
  wire h_u_cla32_and1966_y0;
  wire h_u_cla32_and1967_y0;
  wire h_u_cla32_and1968_y0;
  wire h_u_cla32_and1969_y0;
  wire h_u_cla32_and1970_y0;
  wire h_u_cla32_and1971_y0;
  wire h_u_cla32_and1972_y0;
  wire h_u_cla32_and1973_y0;
  wire h_u_cla32_and1974_y0;
  wire h_u_cla32_and1975_y0;
  wire h_u_cla32_and1976_y0;
  wire h_u_cla32_and1977_y0;
  wire h_u_cla32_and1978_y0;
  wire h_u_cla32_and1979_y0;
  wire h_u_cla32_and1980_y0;
  wire h_u_cla32_and1981_y0;
  wire h_u_cla32_and1982_y0;
  wire h_u_cla32_and1983_y0;
  wire h_u_cla32_and1984_y0;
  wire h_u_cla32_and1985_y0;
  wire h_u_cla32_and1986_y0;
  wire h_u_cla32_and1987_y0;
  wire h_u_cla32_and1988_y0;
  wire h_u_cla32_and1989_y0;
  wire h_u_cla32_and1990_y0;
  wire h_u_cla32_and1991_y0;
  wire h_u_cla32_and1992_y0;
  wire h_u_cla32_and1993_y0;
  wire h_u_cla32_and1994_y0;
  wire h_u_cla32_and1995_y0;
  wire h_u_cla32_and1996_y0;
  wire h_u_cla32_and1997_y0;
  wire h_u_cla32_and1998_y0;
  wire h_u_cla32_and1999_y0;
  wire h_u_cla32_and2000_y0;
  wire h_u_cla32_and2001_y0;
  wire h_u_cla32_and2002_y0;
  wire h_u_cla32_and2003_y0;
  wire h_u_cla32_and2004_y0;
  wire h_u_cla32_and2005_y0;
  wire h_u_cla32_and2006_y0;
  wire h_u_cla32_and2007_y0;
  wire h_u_cla32_and2008_y0;
  wire h_u_cla32_and2009_y0;
  wire h_u_cla32_and2010_y0;
  wire h_u_cla32_and2011_y0;
  wire h_u_cla32_and2012_y0;
  wire h_u_cla32_and2013_y0;
  wire h_u_cla32_and2014_y0;
  wire h_u_cla32_and2015_y0;
  wire h_u_cla32_and2016_y0;
  wire h_u_cla32_and2017_y0;
  wire h_u_cla32_and2018_y0;
  wire h_u_cla32_and2019_y0;
  wire h_u_cla32_and2020_y0;
  wire h_u_cla32_and2021_y0;
  wire h_u_cla32_and2022_y0;
  wire h_u_cla32_and2023_y0;
  wire h_u_cla32_and2024_y0;
  wire h_u_cla32_and2025_y0;
  wire h_u_cla32_and2026_y0;
  wire h_u_cla32_and2027_y0;
  wire h_u_cla32_and2028_y0;
  wire h_u_cla32_and2029_y0;
  wire h_u_cla32_and2030_y0;
  wire h_u_cla32_and2031_y0;
  wire h_u_cla32_and2032_y0;
  wire h_u_cla32_and2033_y0;
  wire h_u_cla32_and2034_y0;
  wire h_u_cla32_and2035_y0;
  wire h_u_cla32_and2036_y0;
  wire h_u_cla32_and2037_y0;
  wire h_u_cla32_and2038_y0;
  wire h_u_cla32_and2039_y0;
  wire h_u_cla32_and2040_y0;
  wire h_u_cla32_and2041_y0;
  wire h_u_cla32_and2042_y0;
  wire h_u_cla32_and2043_y0;
  wire h_u_cla32_and2044_y0;
  wire h_u_cla32_and2045_y0;
  wire h_u_cla32_and2046_y0;
  wire h_u_cla32_and2047_y0;
  wire h_u_cla32_and2048_y0;
  wire h_u_cla32_and2049_y0;
  wire h_u_cla32_and2050_y0;
  wire h_u_cla32_and2051_y0;
  wire h_u_cla32_and2052_y0;
  wire h_u_cla32_and2053_y0;
  wire h_u_cla32_and2054_y0;
  wire h_u_cla32_and2055_y0;
  wire h_u_cla32_and2056_y0;
  wire h_u_cla32_and2057_y0;
  wire h_u_cla32_and2058_y0;
  wire h_u_cla32_and2059_y0;
  wire h_u_cla32_and2060_y0;
  wire h_u_cla32_and2061_y0;
  wire h_u_cla32_and2062_y0;
  wire h_u_cla32_and2063_y0;
  wire h_u_cla32_and2064_y0;
  wire h_u_cla32_and2065_y0;
  wire h_u_cla32_and2066_y0;
  wire h_u_cla32_and2067_y0;
  wire h_u_cla32_and2068_y0;
  wire h_u_cla32_and2069_y0;
  wire h_u_cla32_and2070_y0;
  wire h_u_cla32_and2071_y0;
  wire h_u_cla32_and2072_y0;
  wire h_u_cla32_and2073_y0;
  wire h_u_cla32_and2074_y0;
  wire h_u_cla32_and2075_y0;
  wire h_u_cla32_and2076_y0;
  wire h_u_cla32_and2077_y0;
  wire h_u_cla32_and2078_y0;
  wire h_u_cla32_and2079_y0;
  wire h_u_cla32_and2080_y0;
  wire h_u_cla32_and2081_y0;
  wire h_u_cla32_and2082_y0;
  wire h_u_cla32_and2083_y0;
  wire h_u_cla32_and2084_y0;
  wire h_u_cla32_and2085_y0;
  wire h_u_cla32_and2086_y0;
  wire h_u_cla32_and2087_y0;
  wire h_u_cla32_and2088_y0;
  wire h_u_cla32_and2089_y0;
  wire h_u_cla32_and2090_y0;
  wire h_u_cla32_and2091_y0;
  wire h_u_cla32_and2092_y0;
  wire h_u_cla32_and2093_y0;
  wire h_u_cla32_and2094_y0;
  wire h_u_cla32_and2095_y0;
  wire h_u_cla32_and2096_y0;
  wire h_u_cla32_and2097_y0;
  wire h_u_cla32_and2098_y0;
  wire h_u_cla32_and2099_y0;
  wire h_u_cla32_and2100_y0;
  wire h_u_cla32_and2101_y0;
  wire h_u_cla32_and2102_y0;
  wire h_u_cla32_and2103_y0;
  wire h_u_cla32_and2104_y0;
  wire h_u_cla32_and2105_y0;
  wire h_u_cla32_and2106_y0;
  wire h_u_cla32_and2107_y0;
  wire h_u_cla32_and2108_y0;
  wire h_u_cla32_or153_y0;
  wire h_u_cla32_or154_y0;
  wire h_u_cla32_or155_y0;
  wire h_u_cla32_or156_y0;
  wire h_u_cla32_or157_y0;
  wire h_u_cla32_or158_y0;
  wire h_u_cla32_or159_y0;
  wire h_u_cla32_or160_y0;
  wire h_u_cla32_or161_y0;
  wire h_u_cla32_or162_y0;
  wire h_u_cla32_or163_y0;
  wire h_u_cla32_or164_y0;
  wire h_u_cla32_or165_y0;
  wire h_u_cla32_or166_y0;
  wire h_u_cla32_or167_y0;
  wire h_u_cla32_or168_y0;
  wire h_u_cla32_or169_y0;
  wire h_u_cla32_or170_y0;
  wire h_u_cla32_pg_logic18_y0;
  wire h_u_cla32_pg_logic18_y1;
  wire h_u_cla32_pg_logic18_y2;
  wire h_u_cla32_xor18_y0;
  wire h_u_cla32_and2109_y0;
  wire h_u_cla32_and2110_y0;
  wire h_u_cla32_and2111_y0;
  wire h_u_cla32_and2112_y0;
  wire h_u_cla32_and2113_y0;
  wire h_u_cla32_and2114_y0;
  wire h_u_cla32_and2115_y0;
  wire h_u_cla32_and2116_y0;
  wire h_u_cla32_and2117_y0;
  wire h_u_cla32_and2118_y0;
  wire h_u_cla32_and2119_y0;
  wire h_u_cla32_and2120_y0;
  wire h_u_cla32_and2121_y0;
  wire h_u_cla32_and2122_y0;
  wire h_u_cla32_and2123_y0;
  wire h_u_cla32_and2124_y0;
  wire h_u_cla32_and2125_y0;
  wire h_u_cla32_and2126_y0;
  wire h_u_cla32_and2127_y0;
  wire h_u_cla32_and2128_y0;
  wire h_u_cla32_and2129_y0;
  wire h_u_cla32_and2130_y0;
  wire h_u_cla32_and2131_y0;
  wire h_u_cla32_and2132_y0;
  wire h_u_cla32_and2133_y0;
  wire h_u_cla32_and2134_y0;
  wire h_u_cla32_and2135_y0;
  wire h_u_cla32_and2136_y0;
  wire h_u_cla32_and2137_y0;
  wire h_u_cla32_and2138_y0;
  wire h_u_cla32_and2139_y0;
  wire h_u_cla32_and2140_y0;
  wire h_u_cla32_and2141_y0;
  wire h_u_cla32_and2142_y0;
  wire h_u_cla32_and2143_y0;
  wire h_u_cla32_and2144_y0;
  wire h_u_cla32_and2145_y0;
  wire h_u_cla32_and2146_y0;
  wire h_u_cla32_and2147_y0;
  wire h_u_cla32_and2148_y0;
  wire h_u_cla32_and2149_y0;
  wire h_u_cla32_and2150_y0;
  wire h_u_cla32_and2151_y0;
  wire h_u_cla32_and2152_y0;
  wire h_u_cla32_and2153_y0;
  wire h_u_cla32_and2154_y0;
  wire h_u_cla32_and2155_y0;
  wire h_u_cla32_and2156_y0;
  wire h_u_cla32_and2157_y0;
  wire h_u_cla32_and2158_y0;
  wire h_u_cla32_and2159_y0;
  wire h_u_cla32_and2160_y0;
  wire h_u_cla32_and2161_y0;
  wire h_u_cla32_and2162_y0;
  wire h_u_cla32_and2163_y0;
  wire h_u_cla32_and2164_y0;
  wire h_u_cla32_and2165_y0;
  wire h_u_cla32_and2166_y0;
  wire h_u_cla32_and2167_y0;
  wire h_u_cla32_and2168_y0;
  wire h_u_cla32_and2169_y0;
  wire h_u_cla32_and2170_y0;
  wire h_u_cla32_and2171_y0;
  wire h_u_cla32_and2172_y0;
  wire h_u_cla32_and2173_y0;
  wire h_u_cla32_and2174_y0;
  wire h_u_cla32_and2175_y0;
  wire h_u_cla32_and2176_y0;
  wire h_u_cla32_and2177_y0;
  wire h_u_cla32_and2178_y0;
  wire h_u_cla32_and2179_y0;
  wire h_u_cla32_and2180_y0;
  wire h_u_cla32_and2181_y0;
  wire h_u_cla32_and2182_y0;
  wire h_u_cla32_and2183_y0;
  wire h_u_cla32_and2184_y0;
  wire h_u_cla32_and2185_y0;
  wire h_u_cla32_and2186_y0;
  wire h_u_cla32_and2187_y0;
  wire h_u_cla32_and2188_y0;
  wire h_u_cla32_and2189_y0;
  wire h_u_cla32_and2190_y0;
  wire h_u_cla32_and2191_y0;
  wire h_u_cla32_and2192_y0;
  wire h_u_cla32_and2193_y0;
  wire h_u_cla32_and2194_y0;
  wire h_u_cla32_and2195_y0;
  wire h_u_cla32_and2196_y0;
  wire h_u_cla32_and2197_y0;
  wire h_u_cla32_and2198_y0;
  wire h_u_cla32_and2199_y0;
  wire h_u_cla32_and2200_y0;
  wire h_u_cla32_and2201_y0;
  wire h_u_cla32_and2202_y0;
  wire h_u_cla32_and2203_y0;
  wire h_u_cla32_and2204_y0;
  wire h_u_cla32_and2205_y0;
  wire h_u_cla32_and2206_y0;
  wire h_u_cla32_and2207_y0;
  wire h_u_cla32_and2208_y0;
  wire h_u_cla32_and2209_y0;
  wire h_u_cla32_and2210_y0;
  wire h_u_cla32_and2211_y0;
  wire h_u_cla32_and2212_y0;
  wire h_u_cla32_and2213_y0;
  wire h_u_cla32_and2214_y0;
  wire h_u_cla32_and2215_y0;
  wire h_u_cla32_and2216_y0;
  wire h_u_cla32_and2217_y0;
  wire h_u_cla32_and2218_y0;
  wire h_u_cla32_and2219_y0;
  wire h_u_cla32_and2220_y0;
  wire h_u_cla32_and2221_y0;
  wire h_u_cla32_and2222_y0;
  wire h_u_cla32_and2223_y0;
  wire h_u_cla32_and2224_y0;
  wire h_u_cla32_and2225_y0;
  wire h_u_cla32_and2226_y0;
  wire h_u_cla32_and2227_y0;
  wire h_u_cla32_and2228_y0;
  wire h_u_cla32_and2229_y0;
  wire h_u_cla32_and2230_y0;
  wire h_u_cla32_and2231_y0;
  wire h_u_cla32_and2232_y0;
  wire h_u_cla32_and2233_y0;
  wire h_u_cla32_and2234_y0;
  wire h_u_cla32_and2235_y0;
  wire h_u_cla32_and2236_y0;
  wire h_u_cla32_and2237_y0;
  wire h_u_cla32_and2238_y0;
  wire h_u_cla32_and2239_y0;
  wire h_u_cla32_and2240_y0;
  wire h_u_cla32_and2241_y0;
  wire h_u_cla32_and2242_y0;
  wire h_u_cla32_and2243_y0;
  wire h_u_cla32_and2244_y0;
  wire h_u_cla32_and2245_y0;
  wire h_u_cla32_and2246_y0;
  wire h_u_cla32_and2247_y0;
  wire h_u_cla32_and2248_y0;
  wire h_u_cla32_and2249_y0;
  wire h_u_cla32_and2250_y0;
  wire h_u_cla32_and2251_y0;
  wire h_u_cla32_and2252_y0;
  wire h_u_cla32_and2253_y0;
  wire h_u_cla32_and2254_y0;
  wire h_u_cla32_and2255_y0;
  wire h_u_cla32_and2256_y0;
  wire h_u_cla32_and2257_y0;
  wire h_u_cla32_and2258_y0;
  wire h_u_cla32_and2259_y0;
  wire h_u_cla32_and2260_y0;
  wire h_u_cla32_and2261_y0;
  wire h_u_cla32_and2262_y0;
  wire h_u_cla32_and2263_y0;
  wire h_u_cla32_and2264_y0;
  wire h_u_cla32_and2265_y0;
  wire h_u_cla32_and2266_y0;
  wire h_u_cla32_and2267_y0;
  wire h_u_cla32_and2268_y0;
  wire h_u_cla32_and2269_y0;
  wire h_u_cla32_and2270_y0;
  wire h_u_cla32_and2271_y0;
  wire h_u_cla32_and2272_y0;
  wire h_u_cla32_and2273_y0;
  wire h_u_cla32_and2274_y0;
  wire h_u_cla32_and2275_y0;
  wire h_u_cla32_and2276_y0;
  wire h_u_cla32_and2277_y0;
  wire h_u_cla32_and2278_y0;
  wire h_u_cla32_and2279_y0;
  wire h_u_cla32_and2280_y0;
  wire h_u_cla32_and2281_y0;
  wire h_u_cla32_and2282_y0;
  wire h_u_cla32_and2283_y0;
  wire h_u_cla32_and2284_y0;
  wire h_u_cla32_and2285_y0;
  wire h_u_cla32_and2286_y0;
  wire h_u_cla32_and2287_y0;
  wire h_u_cla32_and2288_y0;
  wire h_u_cla32_and2289_y0;
  wire h_u_cla32_and2290_y0;
  wire h_u_cla32_and2291_y0;
  wire h_u_cla32_and2292_y0;
  wire h_u_cla32_and2293_y0;
  wire h_u_cla32_and2294_y0;
  wire h_u_cla32_and2295_y0;
  wire h_u_cla32_and2296_y0;
  wire h_u_cla32_and2297_y0;
  wire h_u_cla32_and2298_y0;
  wire h_u_cla32_and2299_y0;
  wire h_u_cla32_and2300_y0;
  wire h_u_cla32_and2301_y0;
  wire h_u_cla32_and2302_y0;
  wire h_u_cla32_and2303_y0;
  wire h_u_cla32_and2304_y0;
  wire h_u_cla32_and2305_y0;
  wire h_u_cla32_and2306_y0;
  wire h_u_cla32_and2307_y0;
  wire h_u_cla32_and2308_y0;
  wire h_u_cla32_and2309_y0;
  wire h_u_cla32_and2310_y0;
  wire h_u_cla32_and2311_y0;
  wire h_u_cla32_and2312_y0;
  wire h_u_cla32_and2313_y0;
  wire h_u_cla32_and2314_y0;
  wire h_u_cla32_and2315_y0;
  wire h_u_cla32_and2316_y0;
  wire h_u_cla32_and2317_y0;
  wire h_u_cla32_and2318_y0;
  wire h_u_cla32_and2319_y0;
  wire h_u_cla32_and2320_y0;
  wire h_u_cla32_and2321_y0;
  wire h_u_cla32_and2322_y0;
  wire h_u_cla32_and2323_y0;
  wire h_u_cla32_and2324_y0;
  wire h_u_cla32_and2325_y0;
  wire h_u_cla32_and2326_y0;
  wire h_u_cla32_and2327_y0;
  wire h_u_cla32_and2328_y0;
  wire h_u_cla32_and2329_y0;
  wire h_u_cla32_and2330_y0;
  wire h_u_cla32_and2331_y0;
  wire h_u_cla32_and2332_y0;
  wire h_u_cla32_and2333_y0;
  wire h_u_cla32_and2334_y0;
  wire h_u_cla32_and2335_y0;
  wire h_u_cla32_and2336_y0;
  wire h_u_cla32_and2337_y0;
  wire h_u_cla32_and2338_y0;
  wire h_u_cla32_and2339_y0;
  wire h_u_cla32_and2340_y0;
  wire h_u_cla32_and2341_y0;
  wire h_u_cla32_and2342_y0;
  wire h_u_cla32_and2343_y0;
  wire h_u_cla32_and2344_y0;
  wire h_u_cla32_and2345_y0;
  wire h_u_cla32_and2346_y0;
  wire h_u_cla32_and2347_y0;
  wire h_u_cla32_and2348_y0;
  wire h_u_cla32_and2349_y0;
  wire h_u_cla32_and2350_y0;
  wire h_u_cla32_and2351_y0;
  wire h_u_cla32_and2352_y0;
  wire h_u_cla32_and2353_y0;
  wire h_u_cla32_and2354_y0;
  wire h_u_cla32_and2355_y0;
  wire h_u_cla32_and2356_y0;
  wire h_u_cla32_and2357_y0;
  wire h_u_cla32_and2358_y0;
  wire h_u_cla32_and2359_y0;
  wire h_u_cla32_and2360_y0;
  wire h_u_cla32_and2361_y0;
  wire h_u_cla32_and2362_y0;
  wire h_u_cla32_and2363_y0;
  wire h_u_cla32_and2364_y0;
  wire h_u_cla32_and2365_y0;
  wire h_u_cla32_and2366_y0;
  wire h_u_cla32_and2367_y0;
  wire h_u_cla32_and2368_y0;
  wire h_u_cla32_and2369_y0;
  wire h_u_cla32_and2370_y0;
  wire h_u_cla32_and2371_y0;
  wire h_u_cla32_and2372_y0;
  wire h_u_cla32_and2373_y0;
  wire h_u_cla32_and2374_y0;
  wire h_u_cla32_and2375_y0;
  wire h_u_cla32_and2376_y0;
  wire h_u_cla32_and2377_y0;
  wire h_u_cla32_and2378_y0;
  wire h_u_cla32_and2379_y0;
  wire h_u_cla32_and2380_y0;
  wire h_u_cla32_and2381_y0;
  wire h_u_cla32_and2382_y0;
  wire h_u_cla32_and2383_y0;
  wire h_u_cla32_and2384_y0;
  wire h_u_cla32_and2385_y0;
  wire h_u_cla32_and2386_y0;
  wire h_u_cla32_and2387_y0;
  wire h_u_cla32_and2388_y0;
  wire h_u_cla32_and2389_y0;
  wire h_u_cla32_and2390_y0;
  wire h_u_cla32_and2391_y0;
  wire h_u_cla32_and2392_y0;
  wire h_u_cla32_and2393_y0;
  wire h_u_cla32_and2394_y0;
  wire h_u_cla32_and2395_y0;
  wire h_u_cla32_and2396_y0;
  wire h_u_cla32_and2397_y0;
  wire h_u_cla32_and2398_y0;
  wire h_u_cla32_and2399_y0;
  wire h_u_cla32_and2400_y0;
  wire h_u_cla32_and2401_y0;
  wire h_u_cla32_and2402_y0;
  wire h_u_cla32_and2403_y0;
  wire h_u_cla32_and2404_y0;
  wire h_u_cla32_and2405_y0;
  wire h_u_cla32_and2406_y0;
  wire h_u_cla32_and2407_y0;
  wire h_u_cla32_and2408_y0;
  wire h_u_cla32_and2409_y0;
  wire h_u_cla32_and2410_y0;
  wire h_u_cla32_and2411_y0;
  wire h_u_cla32_and2412_y0;
  wire h_u_cla32_and2413_y0;
  wire h_u_cla32_and2414_y0;
  wire h_u_cla32_and2415_y0;
  wire h_u_cla32_and2416_y0;
  wire h_u_cla32_and2417_y0;
  wire h_u_cla32_and2418_y0;
  wire h_u_cla32_and2419_y0;
  wire h_u_cla32_and2420_y0;
  wire h_u_cla32_and2421_y0;
  wire h_u_cla32_and2422_y0;
  wire h_u_cla32_and2423_y0;
  wire h_u_cla32_and2424_y0;
  wire h_u_cla32_and2425_y0;
  wire h_u_cla32_and2426_y0;
  wire h_u_cla32_and2427_y0;
  wire h_u_cla32_and2428_y0;
  wire h_u_cla32_and2429_y0;
  wire h_u_cla32_and2430_y0;
  wire h_u_cla32_and2431_y0;
  wire h_u_cla32_and2432_y0;
  wire h_u_cla32_and2433_y0;
  wire h_u_cla32_and2434_y0;
  wire h_u_cla32_and2435_y0;
  wire h_u_cla32_and2436_y0;
  wire h_u_cla32_and2437_y0;
  wire h_u_cla32_and2438_y0;
  wire h_u_cla32_and2439_y0;
  wire h_u_cla32_and2440_y0;
  wire h_u_cla32_and2441_y0;
  wire h_u_cla32_and2442_y0;
  wire h_u_cla32_and2443_y0;
  wire h_u_cla32_and2444_y0;
  wire h_u_cla32_and2445_y0;
  wire h_u_cla32_and2446_y0;
  wire h_u_cla32_and2447_y0;
  wire h_u_cla32_and2448_y0;
  wire h_u_cla32_and2449_y0;
  wire h_u_cla32_and2450_y0;
  wire h_u_cla32_and2451_y0;
  wire h_u_cla32_and2452_y0;
  wire h_u_cla32_and2453_y0;
  wire h_u_cla32_and2454_y0;
  wire h_u_cla32_and2455_y0;
  wire h_u_cla32_and2456_y0;
  wire h_u_cla32_and2457_y0;
  wire h_u_cla32_and2458_y0;
  wire h_u_cla32_and2459_y0;
  wire h_u_cla32_and2460_y0;
  wire h_u_cla32_and2461_y0;
  wire h_u_cla32_and2462_y0;
  wire h_u_cla32_and2463_y0;
  wire h_u_cla32_and2464_y0;
  wire h_u_cla32_and2465_y0;
  wire h_u_cla32_and2466_y0;
  wire h_u_cla32_and2467_y0;
  wire h_u_cla32_and2468_y0;
  wire h_u_cla32_and2469_y0;
  wire h_u_cla32_or171_y0;
  wire h_u_cla32_or172_y0;
  wire h_u_cla32_or173_y0;
  wire h_u_cla32_or174_y0;
  wire h_u_cla32_or175_y0;
  wire h_u_cla32_or176_y0;
  wire h_u_cla32_or177_y0;
  wire h_u_cla32_or178_y0;
  wire h_u_cla32_or179_y0;
  wire h_u_cla32_or180_y0;
  wire h_u_cla32_or181_y0;
  wire h_u_cla32_or182_y0;
  wire h_u_cla32_or183_y0;
  wire h_u_cla32_or184_y0;
  wire h_u_cla32_or185_y0;
  wire h_u_cla32_or186_y0;
  wire h_u_cla32_or187_y0;
  wire h_u_cla32_or188_y0;
  wire h_u_cla32_or189_y0;
  wire h_u_cla32_pg_logic19_y0;
  wire h_u_cla32_pg_logic19_y1;
  wire h_u_cla32_pg_logic19_y2;
  wire h_u_cla32_xor19_y0;
  wire h_u_cla32_and2470_y0;
  wire h_u_cla32_and2471_y0;
  wire h_u_cla32_and2472_y0;
  wire h_u_cla32_and2473_y0;
  wire h_u_cla32_and2474_y0;
  wire h_u_cla32_and2475_y0;
  wire h_u_cla32_and2476_y0;
  wire h_u_cla32_and2477_y0;
  wire h_u_cla32_and2478_y0;
  wire h_u_cla32_and2479_y0;
  wire h_u_cla32_and2480_y0;
  wire h_u_cla32_and2481_y0;
  wire h_u_cla32_and2482_y0;
  wire h_u_cla32_and2483_y0;
  wire h_u_cla32_and2484_y0;
  wire h_u_cla32_and2485_y0;
  wire h_u_cla32_and2486_y0;
  wire h_u_cla32_and2487_y0;
  wire h_u_cla32_and2488_y0;
  wire h_u_cla32_and2489_y0;
  wire h_u_cla32_and2490_y0;
  wire h_u_cla32_and2491_y0;
  wire h_u_cla32_and2492_y0;
  wire h_u_cla32_and2493_y0;
  wire h_u_cla32_and2494_y0;
  wire h_u_cla32_and2495_y0;
  wire h_u_cla32_and2496_y0;
  wire h_u_cla32_and2497_y0;
  wire h_u_cla32_and2498_y0;
  wire h_u_cla32_and2499_y0;
  wire h_u_cla32_and2500_y0;
  wire h_u_cla32_and2501_y0;
  wire h_u_cla32_and2502_y0;
  wire h_u_cla32_and2503_y0;
  wire h_u_cla32_and2504_y0;
  wire h_u_cla32_and2505_y0;
  wire h_u_cla32_and2506_y0;
  wire h_u_cla32_and2507_y0;
  wire h_u_cla32_and2508_y0;
  wire h_u_cla32_and2509_y0;
  wire h_u_cla32_and2510_y0;
  wire h_u_cla32_and2511_y0;
  wire h_u_cla32_and2512_y0;
  wire h_u_cla32_and2513_y0;
  wire h_u_cla32_and2514_y0;
  wire h_u_cla32_and2515_y0;
  wire h_u_cla32_and2516_y0;
  wire h_u_cla32_and2517_y0;
  wire h_u_cla32_and2518_y0;
  wire h_u_cla32_and2519_y0;
  wire h_u_cla32_and2520_y0;
  wire h_u_cla32_and2521_y0;
  wire h_u_cla32_and2522_y0;
  wire h_u_cla32_and2523_y0;
  wire h_u_cla32_and2524_y0;
  wire h_u_cla32_and2525_y0;
  wire h_u_cla32_and2526_y0;
  wire h_u_cla32_and2527_y0;
  wire h_u_cla32_and2528_y0;
  wire h_u_cla32_and2529_y0;
  wire h_u_cla32_and2530_y0;
  wire h_u_cla32_and2531_y0;
  wire h_u_cla32_and2532_y0;
  wire h_u_cla32_and2533_y0;
  wire h_u_cla32_and2534_y0;
  wire h_u_cla32_and2535_y0;
  wire h_u_cla32_and2536_y0;
  wire h_u_cla32_and2537_y0;
  wire h_u_cla32_and2538_y0;
  wire h_u_cla32_and2539_y0;
  wire h_u_cla32_and2540_y0;
  wire h_u_cla32_and2541_y0;
  wire h_u_cla32_and2542_y0;
  wire h_u_cla32_and2543_y0;
  wire h_u_cla32_and2544_y0;
  wire h_u_cla32_and2545_y0;
  wire h_u_cla32_and2546_y0;
  wire h_u_cla32_and2547_y0;
  wire h_u_cla32_and2548_y0;
  wire h_u_cla32_and2549_y0;
  wire h_u_cla32_and2550_y0;
  wire h_u_cla32_and2551_y0;
  wire h_u_cla32_and2552_y0;
  wire h_u_cla32_and2553_y0;
  wire h_u_cla32_and2554_y0;
  wire h_u_cla32_and2555_y0;
  wire h_u_cla32_and2556_y0;
  wire h_u_cla32_and2557_y0;
  wire h_u_cla32_and2558_y0;
  wire h_u_cla32_and2559_y0;
  wire h_u_cla32_and2560_y0;
  wire h_u_cla32_and2561_y0;
  wire h_u_cla32_and2562_y0;
  wire h_u_cla32_and2563_y0;
  wire h_u_cla32_and2564_y0;
  wire h_u_cla32_and2565_y0;
  wire h_u_cla32_and2566_y0;
  wire h_u_cla32_and2567_y0;
  wire h_u_cla32_and2568_y0;
  wire h_u_cla32_and2569_y0;
  wire h_u_cla32_and2570_y0;
  wire h_u_cla32_and2571_y0;
  wire h_u_cla32_and2572_y0;
  wire h_u_cla32_and2573_y0;
  wire h_u_cla32_and2574_y0;
  wire h_u_cla32_and2575_y0;
  wire h_u_cla32_and2576_y0;
  wire h_u_cla32_and2577_y0;
  wire h_u_cla32_and2578_y0;
  wire h_u_cla32_and2579_y0;
  wire h_u_cla32_and2580_y0;
  wire h_u_cla32_and2581_y0;
  wire h_u_cla32_and2582_y0;
  wire h_u_cla32_and2583_y0;
  wire h_u_cla32_and2584_y0;
  wire h_u_cla32_and2585_y0;
  wire h_u_cla32_and2586_y0;
  wire h_u_cla32_and2587_y0;
  wire h_u_cla32_and2588_y0;
  wire h_u_cla32_and2589_y0;
  wire h_u_cla32_and2590_y0;
  wire h_u_cla32_and2591_y0;
  wire h_u_cla32_and2592_y0;
  wire h_u_cla32_and2593_y0;
  wire h_u_cla32_and2594_y0;
  wire h_u_cla32_and2595_y0;
  wire h_u_cla32_and2596_y0;
  wire h_u_cla32_and2597_y0;
  wire h_u_cla32_and2598_y0;
  wire h_u_cla32_and2599_y0;
  wire h_u_cla32_and2600_y0;
  wire h_u_cla32_and2601_y0;
  wire h_u_cla32_and2602_y0;
  wire h_u_cla32_and2603_y0;
  wire h_u_cla32_and2604_y0;
  wire h_u_cla32_and2605_y0;
  wire h_u_cla32_and2606_y0;
  wire h_u_cla32_and2607_y0;
  wire h_u_cla32_and2608_y0;
  wire h_u_cla32_and2609_y0;
  wire h_u_cla32_and2610_y0;
  wire h_u_cla32_and2611_y0;
  wire h_u_cla32_and2612_y0;
  wire h_u_cla32_and2613_y0;
  wire h_u_cla32_and2614_y0;
  wire h_u_cla32_and2615_y0;
  wire h_u_cla32_and2616_y0;
  wire h_u_cla32_and2617_y0;
  wire h_u_cla32_and2618_y0;
  wire h_u_cla32_and2619_y0;
  wire h_u_cla32_and2620_y0;
  wire h_u_cla32_and2621_y0;
  wire h_u_cla32_and2622_y0;
  wire h_u_cla32_and2623_y0;
  wire h_u_cla32_and2624_y0;
  wire h_u_cla32_and2625_y0;
  wire h_u_cla32_and2626_y0;
  wire h_u_cla32_and2627_y0;
  wire h_u_cla32_and2628_y0;
  wire h_u_cla32_and2629_y0;
  wire h_u_cla32_and2630_y0;
  wire h_u_cla32_and2631_y0;
  wire h_u_cla32_and2632_y0;
  wire h_u_cla32_and2633_y0;
  wire h_u_cla32_and2634_y0;
  wire h_u_cla32_and2635_y0;
  wire h_u_cla32_and2636_y0;
  wire h_u_cla32_and2637_y0;
  wire h_u_cla32_and2638_y0;
  wire h_u_cla32_and2639_y0;
  wire h_u_cla32_and2640_y0;
  wire h_u_cla32_and2641_y0;
  wire h_u_cla32_and2642_y0;
  wire h_u_cla32_and2643_y0;
  wire h_u_cla32_and2644_y0;
  wire h_u_cla32_and2645_y0;
  wire h_u_cla32_and2646_y0;
  wire h_u_cla32_and2647_y0;
  wire h_u_cla32_and2648_y0;
  wire h_u_cla32_and2649_y0;
  wire h_u_cla32_and2650_y0;
  wire h_u_cla32_and2651_y0;
  wire h_u_cla32_and2652_y0;
  wire h_u_cla32_and2653_y0;
  wire h_u_cla32_and2654_y0;
  wire h_u_cla32_and2655_y0;
  wire h_u_cla32_and2656_y0;
  wire h_u_cla32_and2657_y0;
  wire h_u_cla32_and2658_y0;
  wire h_u_cla32_and2659_y0;
  wire h_u_cla32_and2660_y0;
  wire h_u_cla32_and2661_y0;
  wire h_u_cla32_and2662_y0;
  wire h_u_cla32_and2663_y0;
  wire h_u_cla32_and2664_y0;
  wire h_u_cla32_and2665_y0;
  wire h_u_cla32_and2666_y0;
  wire h_u_cla32_and2667_y0;
  wire h_u_cla32_and2668_y0;
  wire h_u_cla32_and2669_y0;
  wire h_u_cla32_and2670_y0;
  wire h_u_cla32_and2671_y0;
  wire h_u_cla32_and2672_y0;
  wire h_u_cla32_and2673_y0;
  wire h_u_cla32_and2674_y0;
  wire h_u_cla32_and2675_y0;
  wire h_u_cla32_and2676_y0;
  wire h_u_cla32_and2677_y0;
  wire h_u_cla32_and2678_y0;
  wire h_u_cla32_and2679_y0;
  wire h_u_cla32_and2680_y0;
  wire h_u_cla32_and2681_y0;
  wire h_u_cla32_and2682_y0;
  wire h_u_cla32_and2683_y0;
  wire h_u_cla32_and2684_y0;
  wire h_u_cla32_and2685_y0;
  wire h_u_cla32_and2686_y0;
  wire h_u_cla32_and2687_y0;
  wire h_u_cla32_and2688_y0;
  wire h_u_cla32_and2689_y0;
  wire h_u_cla32_and2690_y0;
  wire h_u_cla32_and2691_y0;
  wire h_u_cla32_and2692_y0;
  wire h_u_cla32_and2693_y0;
  wire h_u_cla32_and2694_y0;
  wire h_u_cla32_and2695_y0;
  wire h_u_cla32_and2696_y0;
  wire h_u_cla32_and2697_y0;
  wire h_u_cla32_and2698_y0;
  wire h_u_cla32_and2699_y0;
  wire h_u_cla32_and2700_y0;
  wire h_u_cla32_and2701_y0;
  wire h_u_cla32_and2702_y0;
  wire h_u_cla32_and2703_y0;
  wire h_u_cla32_and2704_y0;
  wire h_u_cla32_and2705_y0;
  wire h_u_cla32_and2706_y0;
  wire h_u_cla32_and2707_y0;
  wire h_u_cla32_and2708_y0;
  wire h_u_cla32_and2709_y0;
  wire h_u_cla32_and2710_y0;
  wire h_u_cla32_and2711_y0;
  wire h_u_cla32_and2712_y0;
  wire h_u_cla32_and2713_y0;
  wire h_u_cla32_and2714_y0;
  wire h_u_cla32_and2715_y0;
  wire h_u_cla32_and2716_y0;
  wire h_u_cla32_and2717_y0;
  wire h_u_cla32_and2718_y0;
  wire h_u_cla32_and2719_y0;
  wire h_u_cla32_and2720_y0;
  wire h_u_cla32_and2721_y0;
  wire h_u_cla32_and2722_y0;
  wire h_u_cla32_and2723_y0;
  wire h_u_cla32_and2724_y0;
  wire h_u_cla32_and2725_y0;
  wire h_u_cla32_and2726_y0;
  wire h_u_cla32_and2727_y0;
  wire h_u_cla32_and2728_y0;
  wire h_u_cla32_and2729_y0;
  wire h_u_cla32_and2730_y0;
  wire h_u_cla32_and2731_y0;
  wire h_u_cla32_and2732_y0;
  wire h_u_cla32_and2733_y0;
  wire h_u_cla32_and2734_y0;
  wire h_u_cla32_and2735_y0;
  wire h_u_cla32_and2736_y0;
  wire h_u_cla32_and2737_y0;
  wire h_u_cla32_and2738_y0;
  wire h_u_cla32_and2739_y0;
  wire h_u_cla32_and2740_y0;
  wire h_u_cla32_and2741_y0;
  wire h_u_cla32_and2742_y0;
  wire h_u_cla32_and2743_y0;
  wire h_u_cla32_and2744_y0;
  wire h_u_cla32_and2745_y0;
  wire h_u_cla32_and2746_y0;
  wire h_u_cla32_and2747_y0;
  wire h_u_cla32_and2748_y0;
  wire h_u_cla32_and2749_y0;
  wire h_u_cla32_and2750_y0;
  wire h_u_cla32_and2751_y0;
  wire h_u_cla32_and2752_y0;
  wire h_u_cla32_and2753_y0;
  wire h_u_cla32_and2754_y0;
  wire h_u_cla32_and2755_y0;
  wire h_u_cla32_and2756_y0;
  wire h_u_cla32_and2757_y0;
  wire h_u_cla32_and2758_y0;
  wire h_u_cla32_and2759_y0;
  wire h_u_cla32_and2760_y0;
  wire h_u_cla32_and2761_y0;
  wire h_u_cla32_and2762_y0;
  wire h_u_cla32_and2763_y0;
  wire h_u_cla32_and2764_y0;
  wire h_u_cla32_and2765_y0;
  wire h_u_cla32_and2766_y0;
  wire h_u_cla32_and2767_y0;
  wire h_u_cla32_and2768_y0;
  wire h_u_cla32_and2769_y0;
  wire h_u_cla32_and2770_y0;
  wire h_u_cla32_and2771_y0;
  wire h_u_cla32_and2772_y0;
  wire h_u_cla32_and2773_y0;
  wire h_u_cla32_and2774_y0;
  wire h_u_cla32_and2775_y0;
  wire h_u_cla32_and2776_y0;
  wire h_u_cla32_and2777_y0;
  wire h_u_cla32_and2778_y0;
  wire h_u_cla32_and2779_y0;
  wire h_u_cla32_and2780_y0;
  wire h_u_cla32_and2781_y0;
  wire h_u_cla32_and2782_y0;
  wire h_u_cla32_and2783_y0;
  wire h_u_cla32_and2784_y0;
  wire h_u_cla32_and2785_y0;
  wire h_u_cla32_and2786_y0;
  wire h_u_cla32_and2787_y0;
  wire h_u_cla32_and2788_y0;
  wire h_u_cla32_and2789_y0;
  wire h_u_cla32_and2790_y0;
  wire h_u_cla32_and2791_y0;
  wire h_u_cla32_and2792_y0;
  wire h_u_cla32_and2793_y0;
  wire h_u_cla32_and2794_y0;
  wire h_u_cla32_and2795_y0;
  wire h_u_cla32_and2796_y0;
  wire h_u_cla32_and2797_y0;
  wire h_u_cla32_and2798_y0;
  wire h_u_cla32_and2799_y0;
  wire h_u_cla32_and2800_y0;
  wire h_u_cla32_and2801_y0;
  wire h_u_cla32_and2802_y0;
  wire h_u_cla32_and2803_y0;
  wire h_u_cla32_and2804_y0;
  wire h_u_cla32_and2805_y0;
  wire h_u_cla32_and2806_y0;
  wire h_u_cla32_and2807_y0;
  wire h_u_cla32_and2808_y0;
  wire h_u_cla32_and2809_y0;
  wire h_u_cla32_and2810_y0;
  wire h_u_cla32_and2811_y0;
  wire h_u_cla32_and2812_y0;
  wire h_u_cla32_and2813_y0;
  wire h_u_cla32_and2814_y0;
  wire h_u_cla32_and2815_y0;
  wire h_u_cla32_and2816_y0;
  wire h_u_cla32_and2817_y0;
  wire h_u_cla32_and2818_y0;
  wire h_u_cla32_and2819_y0;
  wire h_u_cla32_and2820_y0;
  wire h_u_cla32_and2821_y0;
  wire h_u_cla32_and2822_y0;
  wire h_u_cla32_and2823_y0;
  wire h_u_cla32_and2824_y0;
  wire h_u_cla32_and2825_y0;
  wire h_u_cla32_and2826_y0;
  wire h_u_cla32_and2827_y0;
  wire h_u_cla32_and2828_y0;
  wire h_u_cla32_and2829_y0;
  wire h_u_cla32_and2830_y0;
  wire h_u_cla32_and2831_y0;
  wire h_u_cla32_and2832_y0;
  wire h_u_cla32_and2833_y0;
  wire h_u_cla32_and2834_y0;
  wire h_u_cla32_and2835_y0;
  wire h_u_cla32_and2836_y0;
  wire h_u_cla32_and2837_y0;
  wire h_u_cla32_and2838_y0;
  wire h_u_cla32_and2839_y0;
  wire h_u_cla32_and2840_y0;
  wire h_u_cla32_and2841_y0;
  wire h_u_cla32_and2842_y0;
  wire h_u_cla32_and2843_y0;
  wire h_u_cla32_and2844_y0;
  wire h_u_cla32_and2845_y0;
  wire h_u_cla32_and2846_y0;
  wire h_u_cla32_and2847_y0;
  wire h_u_cla32_and2848_y0;
  wire h_u_cla32_and2849_y0;
  wire h_u_cla32_and2850_y0;
  wire h_u_cla32_and2851_y0;
  wire h_u_cla32_and2852_y0;
  wire h_u_cla32_and2853_y0;
  wire h_u_cla32_and2854_y0;
  wire h_u_cla32_and2855_y0;
  wire h_u_cla32_and2856_y0;
  wire h_u_cla32_and2857_y0;
  wire h_u_cla32_and2858_y0;
  wire h_u_cla32_and2859_y0;
  wire h_u_cla32_and2860_y0;
  wire h_u_cla32_and2861_y0;
  wire h_u_cla32_and2862_y0;
  wire h_u_cla32_and2863_y0;
  wire h_u_cla32_and2864_y0;
  wire h_u_cla32_and2865_y0;
  wire h_u_cla32_and2866_y0;
  wire h_u_cla32_and2867_y0;
  wire h_u_cla32_and2868_y0;
  wire h_u_cla32_and2869_y0;
  wire h_u_cla32_or190_y0;
  wire h_u_cla32_or191_y0;
  wire h_u_cla32_or192_y0;
  wire h_u_cla32_or193_y0;
  wire h_u_cla32_or194_y0;
  wire h_u_cla32_or195_y0;
  wire h_u_cla32_or196_y0;
  wire h_u_cla32_or197_y0;
  wire h_u_cla32_or198_y0;
  wire h_u_cla32_or199_y0;
  wire h_u_cla32_or200_y0;
  wire h_u_cla32_or201_y0;
  wire h_u_cla32_or202_y0;
  wire h_u_cla32_or203_y0;
  wire h_u_cla32_or204_y0;
  wire h_u_cla32_or205_y0;
  wire h_u_cla32_or206_y0;
  wire h_u_cla32_or207_y0;
  wire h_u_cla32_or208_y0;
  wire h_u_cla32_or209_y0;
  wire h_u_cla32_pg_logic20_y0;
  wire h_u_cla32_pg_logic20_y1;
  wire h_u_cla32_pg_logic20_y2;
  wire h_u_cla32_xor20_y0;
  wire h_u_cla32_and2870_y0;
  wire h_u_cla32_and2871_y0;
  wire h_u_cla32_and2872_y0;
  wire h_u_cla32_and2873_y0;
  wire h_u_cla32_and2874_y0;
  wire h_u_cla32_and2875_y0;
  wire h_u_cla32_and2876_y0;
  wire h_u_cla32_and2877_y0;
  wire h_u_cla32_and2878_y0;
  wire h_u_cla32_and2879_y0;
  wire h_u_cla32_and2880_y0;
  wire h_u_cla32_and2881_y0;
  wire h_u_cla32_and2882_y0;
  wire h_u_cla32_and2883_y0;
  wire h_u_cla32_and2884_y0;
  wire h_u_cla32_and2885_y0;
  wire h_u_cla32_and2886_y0;
  wire h_u_cla32_and2887_y0;
  wire h_u_cla32_and2888_y0;
  wire h_u_cla32_and2889_y0;
  wire h_u_cla32_and2890_y0;
  wire h_u_cla32_and2891_y0;
  wire h_u_cla32_and2892_y0;
  wire h_u_cla32_and2893_y0;
  wire h_u_cla32_and2894_y0;
  wire h_u_cla32_and2895_y0;
  wire h_u_cla32_and2896_y0;
  wire h_u_cla32_and2897_y0;
  wire h_u_cla32_and2898_y0;
  wire h_u_cla32_and2899_y0;
  wire h_u_cla32_and2900_y0;
  wire h_u_cla32_and2901_y0;
  wire h_u_cla32_and2902_y0;
  wire h_u_cla32_and2903_y0;
  wire h_u_cla32_and2904_y0;
  wire h_u_cla32_and2905_y0;
  wire h_u_cla32_and2906_y0;
  wire h_u_cla32_and2907_y0;
  wire h_u_cla32_and2908_y0;
  wire h_u_cla32_and2909_y0;
  wire h_u_cla32_and2910_y0;
  wire h_u_cla32_and2911_y0;
  wire h_u_cla32_and2912_y0;
  wire h_u_cla32_and2913_y0;
  wire h_u_cla32_and2914_y0;
  wire h_u_cla32_and2915_y0;
  wire h_u_cla32_and2916_y0;
  wire h_u_cla32_and2917_y0;
  wire h_u_cla32_and2918_y0;
  wire h_u_cla32_and2919_y0;
  wire h_u_cla32_and2920_y0;
  wire h_u_cla32_and2921_y0;
  wire h_u_cla32_and2922_y0;
  wire h_u_cla32_and2923_y0;
  wire h_u_cla32_and2924_y0;
  wire h_u_cla32_and2925_y0;
  wire h_u_cla32_and2926_y0;
  wire h_u_cla32_and2927_y0;
  wire h_u_cla32_and2928_y0;
  wire h_u_cla32_and2929_y0;
  wire h_u_cla32_and2930_y0;
  wire h_u_cla32_and2931_y0;
  wire h_u_cla32_and2932_y0;
  wire h_u_cla32_and2933_y0;
  wire h_u_cla32_and2934_y0;
  wire h_u_cla32_and2935_y0;
  wire h_u_cla32_and2936_y0;
  wire h_u_cla32_and2937_y0;
  wire h_u_cla32_and2938_y0;
  wire h_u_cla32_and2939_y0;
  wire h_u_cla32_and2940_y0;
  wire h_u_cla32_and2941_y0;
  wire h_u_cla32_and2942_y0;
  wire h_u_cla32_and2943_y0;
  wire h_u_cla32_and2944_y0;
  wire h_u_cla32_and2945_y0;
  wire h_u_cla32_and2946_y0;
  wire h_u_cla32_and2947_y0;
  wire h_u_cla32_and2948_y0;
  wire h_u_cla32_and2949_y0;
  wire h_u_cla32_and2950_y0;
  wire h_u_cla32_and2951_y0;
  wire h_u_cla32_and2952_y0;
  wire h_u_cla32_and2953_y0;
  wire h_u_cla32_and2954_y0;
  wire h_u_cla32_and2955_y0;
  wire h_u_cla32_and2956_y0;
  wire h_u_cla32_and2957_y0;
  wire h_u_cla32_and2958_y0;
  wire h_u_cla32_and2959_y0;
  wire h_u_cla32_and2960_y0;
  wire h_u_cla32_and2961_y0;
  wire h_u_cla32_and2962_y0;
  wire h_u_cla32_and2963_y0;
  wire h_u_cla32_and2964_y0;
  wire h_u_cla32_and2965_y0;
  wire h_u_cla32_and2966_y0;
  wire h_u_cla32_and2967_y0;
  wire h_u_cla32_and2968_y0;
  wire h_u_cla32_and2969_y0;
  wire h_u_cla32_and2970_y0;
  wire h_u_cla32_and2971_y0;
  wire h_u_cla32_and2972_y0;
  wire h_u_cla32_and2973_y0;
  wire h_u_cla32_and2974_y0;
  wire h_u_cla32_and2975_y0;
  wire h_u_cla32_and2976_y0;
  wire h_u_cla32_and2977_y0;
  wire h_u_cla32_and2978_y0;
  wire h_u_cla32_and2979_y0;
  wire h_u_cla32_and2980_y0;
  wire h_u_cla32_and2981_y0;
  wire h_u_cla32_and2982_y0;
  wire h_u_cla32_and2983_y0;
  wire h_u_cla32_and2984_y0;
  wire h_u_cla32_and2985_y0;
  wire h_u_cla32_and2986_y0;
  wire h_u_cla32_and2987_y0;
  wire h_u_cla32_and2988_y0;
  wire h_u_cla32_and2989_y0;
  wire h_u_cla32_and2990_y0;
  wire h_u_cla32_and2991_y0;
  wire h_u_cla32_and2992_y0;
  wire h_u_cla32_and2993_y0;
  wire h_u_cla32_and2994_y0;
  wire h_u_cla32_and2995_y0;
  wire h_u_cla32_and2996_y0;
  wire h_u_cla32_and2997_y0;
  wire h_u_cla32_and2998_y0;
  wire h_u_cla32_and2999_y0;
  wire h_u_cla32_and3000_y0;
  wire h_u_cla32_and3001_y0;
  wire h_u_cla32_and3002_y0;
  wire h_u_cla32_and3003_y0;
  wire h_u_cla32_and3004_y0;
  wire h_u_cla32_and3005_y0;
  wire h_u_cla32_and3006_y0;
  wire h_u_cla32_and3007_y0;
  wire h_u_cla32_and3008_y0;
  wire h_u_cla32_and3009_y0;
  wire h_u_cla32_and3010_y0;
  wire h_u_cla32_and3011_y0;
  wire h_u_cla32_and3012_y0;
  wire h_u_cla32_and3013_y0;
  wire h_u_cla32_and3014_y0;
  wire h_u_cla32_and3015_y0;
  wire h_u_cla32_and3016_y0;
  wire h_u_cla32_and3017_y0;
  wire h_u_cla32_and3018_y0;
  wire h_u_cla32_and3019_y0;
  wire h_u_cla32_and3020_y0;
  wire h_u_cla32_and3021_y0;
  wire h_u_cla32_and3022_y0;
  wire h_u_cla32_and3023_y0;
  wire h_u_cla32_and3024_y0;
  wire h_u_cla32_and3025_y0;
  wire h_u_cla32_and3026_y0;
  wire h_u_cla32_and3027_y0;
  wire h_u_cla32_and3028_y0;
  wire h_u_cla32_and3029_y0;
  wire h_u_cla32_and3030_y0;
  wire h_u_cla32_and3031_y0;
  wire h_u_cla32_and3032_y0;
  wire h_u_cla32_and3033_y0;
  wire h_u_cla32_and3034_y0;
  wire h_u_cla32_and3035_y0;
  wire h_u_cla32_and3036_y0;
  wire h_u_cla32_and3037_y0;
  wire h_u_cla32_and3038_y0;
  wire h_u_cla32_and3039_y0;
  wire h_u_cla32_and3040_y0;
  wire h_u_cla32_and3041_y0;
  wire h_u_cla32_and3042_y0;
  wire h_u_cla32_and3043_y0;
  wire h_u_cla32_and3044_y0;
  wire h_u_cla32_and3045_y0;
  wire h_u_cla32_and3046_y0;
  wire h_u_cla32_and3047_y0;
  wire h_u_cla32_and3048_y0;
  wire h_u_cla32_and3049_y0;
  wire h_u_cla32_and3050_y0;
  wire h_u_cla32_and3051_y0;
  wire h_u_cla32_and3052_y0;
  wire h_u_cla32_and3053_y0;
  wire h_u_cla32_and3054_y0;
  wire h_u_cla32_and3055_y0;
  wire h_u_cla32_and3056_y0;
  wire h_u_cla32_and3057_y0;
  wire h_u_cla32_and3058_y0;
  wire h_u_cla32_and3059_y0;
  wire h_u_cla32_and3060_y0;
  wire h_u_cla32_and3061_y0;
  wire h_u_cla32_and3062_y0;
  wire h_u_cla32_and3063_y0;
  wire h_u_cla32_and3064_y0;
  wire h_u_cla32_and3065_y0;
  wire h_u_cla32_and3066_y0;
  wire h_u_cla32_and3067_y0;
  wire h_u_cla32_and3068_y0;
  wire h_u_cla32_and3069_y0;
  wire h_u_cla32_and3070_y0;
  wire h_u_cla32_and3071_y0;
  wire h_u_cla32_and3072_y0;
  wire h_u_cla32_and3073_y0;
  wire h_u_cla32_and3074_y0;
  wire h_u_cla32_and3075_y0;
  wire h_u_cla32_and3076_y0;
  wire h_u_cla32_and3077_y0;
  wire h_u_cla32_and3078_y0;
  wire h_u_cla32_and3079_y0;
  wire h_u_cla32_and3080_y0;
  wire h_u_cla32_and3081_y0;
  wire h_u_cla32_and3082_y0;
  wire h_u_cla32_and3083_y0;
  wire h_u_cla32_and3084_y0;
  wire h_u_cla32_and3085_y0;
  wire h_u_cla32_and3086_y0;
  wire h_u_cla32_and3087_y0;
  wire h_u_cla32_and3088_y0;
  wire h_u_cla32_and3089_y0;
  wire h_u_cla32_and3090_y0;
  wire h_u_cla32_and3091_y0;
  wire h_u_cla32_and3092_y0;
  wire h_u_cla32_and3093_y0;
  wire h_u_cla32_and3094_y0;
  wire h_u_cla32_and3095_y0;
  wire h_u_cla32_and3096_y0;
  wire h_u_cla32_and3097_y0;
  wire h_u_cla32_and3098_y0;
  wire h_u_cla32_and3099_y0;
  wire h_u_cla32_and3100_y0;
  wire h_u_cla32_and3101_y0;
  wire h_u_cla32_and3102_y0;
  wire h_u_cla32_and3103_y0;
  wire h_u_cla32_and3104_y0;
  wire h_u_cla32_and3105_y0;
  wire h_u_cla32_and3106_y0;
  wire h_u_cla32_and3107_y0;
  wire h_u_cla32_and3108_y0;
  wire h_u_cla32_and3109_y0;
  wire h_u_cla32_and3110_y0;
  wire h_u_cla32_and3111_y0;
  wire h_u_cla32_and3112_y0;
  wire h_u_cla32_and3113_y0;
  wire h_u_cla32_and3114_y0;
  wire h_u_cla32_and3115_y0;
  wire h_u_cla32_and3116_y0;
  wire h_u_cla32_and3117_y0;
  wire h_u_cla32_and3118_y0;
  wire h_u_cla32_and3119_y0;
  wire h_u_cla32_and3120_y0;
  wire h_u_cla32_and3121_y0;
  wire h_u_cla32_and3122_y0;
  wire h_u_cla32_and3123_y0;
  wire h_u_cla32_and3124_y0;
  wire h_u_cla32_and3125_y0;
  wire h_u_cla32_and3126_y0;
  wire h_u_cla32_and3127_y0;
  wire h_u_cla32_and3128_y0;
  wire h_u_cla32_and3129_y0;
  wire h_u_cla32_and3130_y0;
  wire h_u_cla32_and3131_y0;
  wire h_u_cla32_and3132_y0;
  wire h_u_cla32_and3133_y0;
  wire h_u_cla32_and3134_y0;
  wire h_u_cla32_and3135_y0;
  wire h_u_cla32_and3136_y0;
  wire h_u_cla32_and3137_y0;
  wire h_u_cla32_and3138_y0;
  wire h_u_cla32_and3139_y0;
  wire h_u_cla32_and3140_y0;
  wire h_u_cla32_and3141_y0;
  wire h_u_cla32_and3142_y0;
  wire h_u_cla32_and3143_y0;
  wire h_u_cla32_and3144_y0;
  wire h_u_cla32_and3145_y0;
  wire h_u_cla32_and3146_y0;
  wire h_u_cla32_and3147_y0;
  wire h_u_cla32_and3148_y0;
  wire h_u_cla32_and3149_y0;
  wire h_u_cla32_and3150_y0;
  wire h_u_cla32_and3151_y0;
  wire h_u_cla32_and3152_y0;
  wire h_u_cla32_and3153_y0;
  wire h_u_cla32_and3154_y0;
  wire h_u_cla32_and3155_y0;
  wire h_u_cla32_and3156_y0;
  wire h_u_cla32_and3157_y0;
  wire h_u_cla32_and3158_y0;
  wire h_u_cla32_and3159_y0;
  wire h_u_cla32_and3160_y0;
  wire h_u_cla32_and3161_y0;
  wire h_u_cla32_and3162_y0;
  wire h_u_cla32_and3163_y0;
  wire h_u_cla32_and3164_y0;
  wire h_u_cla32_and3165_y0;
  wire h_u_cla32_and3166_y0;
  wire h_u_cla32_and3167_y0;
  wire h_u_cla32_and3168_y0;
  wire h_u_cla32_and3169_y0;
  wire h_u_cla32_and3170_y0;
  wire h_u_cla32_and3171_y0;
  wire h_u_cla32_and3172_y0;
  wire h_u_cla32_and3173_y0;
  wire h_u_cla32_and3174_y0;
  wire h_u_cla32_and3175_y0;
  wire h_u_cla32_and3176_y0;
  wire h_u_cla32_and3177_y0;
  wire h_u_cla32_and3178_y0;
  wire h_u_cla32_and3179_y0;
  wire h_u_cla32_and3180_y0;
  wire h_u_cla32_and3181_y0;
  wire h_u_cla32_and3182_y0;
  wire h_u_cla32_and3183_y0;
  wire h_u_cla32_and3184_y0;
  wire h_u_cla32_and3185_y0;
  wire h_u_cla32_and3186_y0;
  wire h_u_cla32_and3187_y0;
  wire h_u_cla32_and3188_y0;
  wire h_u_cla32_and3189_y0;
  wire h_u_cla32_and3190_y0;
  wire h_u_cla32_and3191_y0;
  wire h_u_cla32_and3192_y0;
  wire h_u_cla32_and3193_y0;
  wire h_u_cla32_and3194_y0;
  wire h_u_cla32_and3195_y0;
  wire h_u_cla32_and3196_y0;
  wire h_u_cla32_and3197_y0;
  wire h_u_cla32_and3198_y0;
  wire h_u_cla32_and3199_y0;
  wire h_u_cla32_and3200_y0;
  wire h_u_cla32_and3201_y0;
  wire h_u_cla32_and3202_y0;
  wire h_u_cla32_and3203_y0;
  wire h_u_cla32_and3204_y0;
  wire h_u_cla32_and3205_y0;
  wire h_u_cla32_and3206_y0;
  wire h_u_cla32_and3207_y0;
  wire h_u_cla32_and3208_y0;
  wire h_u_cla32_and3209_y0;
  wire h_u_cla32_and3210_y0;
  wire h_u_cla32_and3211_y0;
  wire h_u_cla32_and3212_y0;
  wire h_u_cla32_and3213_y0;
  wire h_u_cla32_and3214_y0;
  wire h_u_cla32_and3215_y0;
  wire h_u_cla32_and3216_y0;
  wire h_u_cla32_and3217_y0;
  wire h_u_cla32_and3218_y0;
  wire h_u_cla32_and3219_y0;
  wire h_u_cla32_and3220_y0;
  wire h_u_cla32_and3221_y0;
  wire h_u_cla32_and3222_y0;
  wire h_u_cla32_and3223_y0;
  wire h_u_cla32_and3224_y0;
  wire h_u_cla32_and3225_y0;
  wire h_u_cla32_and3226_y0;
  wire h_u_cla32_and3227_y0;
  wire h_u_cla32_and3228_y0;
  wire h_u_cla32_and3229_y0;
  wire h_u_cla32_and3230_y0;
  wire h_u_cla32_and3231_y0;
  wire h_u_cla32_and3232_y0;
  wire h_u_cla32_and3233_y0;
  wire h_u_cla32_and3234_y0;
  wire h_u_cla32_and3235_y0;
  wire h_u_cla32_and3236_y0;
  wire h_u_cla32_and3237_y0;
  wire h_u_cla32_and3238_y0;
  wire h_u_cla32_and3239_y0;
  wire h_u_cla32_and3240_y0;
  wire h_u_cla32_and3241_y0;
  wire h_u_cla32_and3242_y0;
  wire h_u_cla32_and3243_y0;
  wire h_u_cla32_and3244_y0;
  wire h_u_cla32_and3245_y0;
  wire h_u_cla32_and3246_y0;
  wire h_u_cla32_and3247_y0;
  wire h_u_cla32_and3248_y0;
  wire h_u_cla32_and3249_y0;
  wire h_u_cla32_and3250_y0;
  wire h_u_cla32_and3251_y0;
  wire h_u_cla32_and3252_y0;
  wire h_u_cla32_and3253_y0;
  wire h_u_cla32_and3254_y0;
  wire h_u_cla32_and3255_y0;
  wire h_u_cla32_and3256_y0;
  wire h_u_cla32_and3257_y0;
  wire h_u_cla32_and3258_y0;
  wire h_u_cla32_and3259_y0;
  wire h_u_cla32_and3260_y0;
  wire h_u_cla32_and3261_y0;
  wire h_u_cla32_and3262_y0;
  wire h_u_cla32_and3263_y0;
  wire h_u_cla32_and3264_y0;
  wire h_u_cla32_and3265_y0;
  wire h_u_cla32_and3266_y0;
  wire h_u_cla32_and3267_y0;
  wire h_u_cla32_and3268_y0;
  wire h_u_cla32_and3269_y0;
  wire h_u_cla32_and3270_y0;
  wire h_u_cla32_and3271_y0;
  wire h_u_cla32_and3272_y0;
  wire h_u_cla32_and3273_y0;
  wire h_u_cla32_and3274_y0;
  wire h_u_cla32_and3275_y0;
  wire h_u_cla32_and3276_y0;
  wire h_u_cla32_and3277_y0;
  wire h_u_cla32_and3278_y0;
  wire h_u_cla32_and3279_y0;
  wire h_u_cla32_and3280_y0;
  wire h_u_cla32_and3281_y0;
  wire h_u_cla32_and3282_y0;
  wire h_u_cla32_and3283_y0;
  wire h_u_cla32_and3284_y0;
  wire h_u_cla32_and3285_y0;
  wire h_u_cla32_and3286_y0;
  wire h_u_cla32_and3287_y0;
  wire h_u_cla32_and3288_y0;
  wire h_u_cla32_and3289_y0;
  wire h_u_cla32_and3290_y0;
  wire h_u_cla32_and3291_y0;
  wire h_u_cla32_and3292_y0;
  wire h_u_cla32_and3293_y0;
  wire h_u_cla32_and3294_y0;
  wire h_u_cla32_and3295_y0;
  wire h_u_cla32_and3296_y0;
  wire h_u_cla32_and3297_y0;
  wire h_u_cla32_and3298_y0;
  wire h_u_cla32_and3299_y0;
  wire h_u_cla32_and3300_y0;
  wire h_u_cla32_and3301_y0;
  wire h_u_cla32_and3302_y0;
  wire h_u_cla32_and3303_y0;
  wire h_u_cla32_and3304_y0;
  wire h_u_cla32_and3305_y0;
  wire h_u_cla32_and3306_y0;
  wire h_u_cla32_and3307_y0;
  wire h_u_cla32_and3308_y0;
  wire h_u_cla32_and3309_y0;
  wire h_u_cla32_and3310_y0;
  wire h_u_cla32_or210_y0;
  wire h_u_cla32_or211_y0;
  wire h_u_cla32_or212_y0;
  wire h_u_cla32_or213_y0;
  wire h_u_cla32_or214_y0;
  wire h_u_cla32_or215_y0;
  wire h_u_cla32_or216_y0;
  wire h_u_cla32_or217_y0;
  wire h_u_cla32_or218_y0;
  wire h_u_cla32_or219_y0;
  wire h_u_cla32_or220_y0;
  wire h_u_cla32_or221_y0;
  wire h_u_cla32_or222_y0;
  wire h_u_cla32_or223_y0;
  wire h_u_cla32_or224_y0;
  wire h_u_cla32_or225_y0;
  wire h_u_cla32_or226_y0;
  wire h_u_cla32_or227_y0;
  wire h_u_cla32_or228_y0;
  wire h_u_cla32_or229_y0;
  wire h_u_cla32_or230_y0;
  wire h_u_cla32_pg_logic21_y0;
  wire h_u_cla32_pg_logic21_y1;
  wire h_u_cla32_pg_logic21_y2;
  wire h_u_cla32_xor21_y0;
  wire h_u_cla32_and3311_y0;
  wire h_u_cla32_and3312_y0;
  wire h_u_cla32_and3313_y0;
  wire h_u_cla32_and3314_y0;
  wire h_u_cla32_and3315_y0;
  wire h_u_cla32_and3316_y0;
  wire h_u_cla32_and3317_y0;
  wire h_u_cla32_and3318_y0;
  wire h_u_cla32_and3319_y0;
  wire h_u_cla32_and3320_y0;
  wire h_u_cla32_and3321_y0;
  wire h_u_cla32_and3322_y0;
  wire h_u_cla32_and3323_y0;
  wire h_u_cla32_and3324_y0;
  wire h_u_cla32_and3325_y0;
  wire h_u_cla32_and3326_y0;
  wire h_u_cla32_and3327_y0;
  wire h_u_cla32_and3328_y0;
  wire h_u_cla32_and3329_y0;
  wire h_u_cla32_and3330_y0;
  wire h_u_cla32_and3331_y0;
  wire h_u_cla32_and3332_y0;
  wire h_u_cla32_and3333_y0;
  wire h_u_cla32_and3334_y0;
  wire h_u_cla32_and3335_y0;
  wire h_u_cla32_and3336_y0;
  wire h_u_cla32_and3337_y0;
  wire h_u_cla32_and3338_y0;
  wire h_u_cla32_and3339_y0;
  wire h_u_cla32_and3340_y0;
  wire h_u_cla32_and3341_y0;
  wire h_u_cla32_and3342_y0;
  wire h_u_cla32_and3343_y0;
  wire h_u_cla32_and3344_y0;
  wire h_u_cla32_and3345_y0;
  wire h_u_cla32_and3346_y0;
  wire h_u_cla32_and3347_y0;
  wire h_u_cla32_and3348_y0;
  wire h_u_cla32_and3349_y0;
  wire h_u_cla32_and3350_y0;
  wire h_u_cla32_and3351_y0;
  wire h_u_cla32_and3352_y0;
  wire h_u_cla32_and3353_y0;
  wire h_u_cla32_and3354_y0;
  wire h_u_cla32_and3355_y0;
  wire h_u_cla32_and3356_y0;
  wire h_u_cla32_and3357_y0;
  wire h_u_cla32_and3358_y0;
  wire h_u_cla32_and3359_y0;
  wire h_u_cla32_and3360_y0;
  wire h_u_cla32_and3361_y0;
  wire h_u_cla32_and3362_y0;
  wire h_u_cla32_and3363_y0;
  wire h_u_cla32_and3364_y0;
  wire h_u_cla32_and3365_y0;
  wire h_u_cla32_and3366_y0;
  wire h_u_cla32_and3367_y0;
  wire h_u_cla32_and3368_y0;
  wire h_u_cla32_and3369_y0;
  wire h_u_cla32_and3370_y0;
  wire h_u_cla32_and3371_y0;
  wire h_u_cla32_and3372_y0;
  wire h_u_cla32_and3373_y0;
  wire h_u_cla32_and3374_y0;
  wire h_u_cla32_and3375_y0;
  wire h_u_cla32_and3376_y0;
  wire h_u_cla32_and3377_y0;
  wire h_u_cla32_and3378_y0;
  wire h_u_cla32_and3379_y0;
  wire h_u_cla32_and3380_y0;
  wire h_u_cla32_and3381_y0;
  wire h_u_cla32_and3382_y0;
  wire h_u_cla32_and3383_y0;
  wire h_u_cla32_and3384_y0;
  wire h_u_cla32_and3385_y0;
  wire h_u_cla32_and3386_y0;
  wire h_u_cla32_and3387_y0;
  wire h_u_cla32_and3388_y0;
  wire h_u_cla32_and3389_y0;
  wire h_u_cla32_and3390_y0;
  wire h_u_cla32_and3391_y0;
  wire h_u_cla32_and3392_y0;
  wire h_u_cla32_and3393_y0;
  wire h_u_cla32_and3394_y0;
  wire h_u_cla32_and3395_y0;
  wire h_u_cla32_and3396_y0;
  wire h_u_cla32_and3397_y0;
  wire h_u_cla32_and3398_y0;
  wire h_u_cla32_and3399_y0;
  wire h_u_cla32_and3400_y0;
  wire h_u_cla32_and3401_y0;
  wire h_u_cla32_and3402_y0;
  wire h_u_cla32_and3403_y0;
  wire h_u_cla32_and3404_y0;
  wire h_u_cla32_and3405_y0;
  wire h_u_cla32_and3406_y0;
  wire h_u_cla32_and3407_y0;
  wire h_u_cla32_and3408_y0;
  wire h_u_cla32_and3409_y0;
  wire h_u_cla32_and3410_y0;
  wire h_u_cla32_and3411_y0;
  wire h_u_cla32_and3412_y0;
  wire h_u_cla32_and3413_y0;
  wire h_u_cla32_and3414_y0;
  wire h_u_cla32_and3415_y0;
  wire h_u_cla32_and3416_y0;
  wire h_u_cla32_and3417_y0;
  wire h_u_cla32_and3418_y0;
  wire h_u_cla32_and3419_y0;
  wire h_u_cla32_and3420_y0;
  wire h_u_cla32_and3421_y0;
  wire h_u_cla32_and3422_y0;
  wire h_u_cla32_and3423_y0;
  wire h_u_cla32_and3424_y0;
  wire h_u_cla32_and3425_y0;
  wire h_u_cla32_and3426_y0;
  wire h_u_cla32_and3427_y0;
  wire h_u_cla32_and3428_y0;
  wire h_u_cla32_and3429_y0;
  wire h_u_cla32_and3430_y0;
  wire h_u_cla32_and3431_y0;
  wire h_u_cla32_and3432_y0;
  wire h_u_cla32_and3433_y0;
  wire h_u_cla32_and3434_y0;
  wire h_u_cla32_and3435_y0;
  wire h_u_cla32_and3436_y0;
  wire h_u_cla32_and3437_y0;
  wire h_u_cla32_and3438_y0;
  wire h_u_cla32_and3439_y0;
  wire h_u_cla32_and3440_y0;
  wire h_u_cla32_and3441_y0;
  wire h_u_cla32_and3442_y0;
  wire h_u_cla32_and3443_y0;
  wire h_u_cla32_and3444_y0;
  wire h_u_cla32_and3445_y0;
  wire h_u_cla32_and3446_y0;
  wire h_u_cla32_and3447_y0;
  wire h_u_cla32_and3448_y0;
  wire h_u_cla32_and3449_y0;
  wire h_u_cla32_and3450_y0;
  wire h_u_cla32_and3451_y0;
  wire h_u_cla32_and3452_y0;
  wire h_u_cla32_and3453_y0;
  wire h_u_cla32_and3454_y0;
  wire h_u_cla32_and3455_y0;
  wire h_u_cla32_and3456_y0;
  wire h_u_cla32_and3457_y0;
  wire h_u_cla32_and3458_y0;
  wire h_u_cla32_and3459_y0;
  wire h_u_cla32_and3460_y0;
  wire h_u_cla32_and3461_y0;
  wire h_u_cla32_and3462_y0;
  wire h_u_cla32_and3463_y0;
  wire h_u_cla32_and3464_y0;
  wire h_u_cla32_and3465_y0;
  wire h_u_cla32_and3466_y0;
  wire h_u_cla32_and3467_y0;
  wire h_u_cla32_and3468_y0;
  wire h_u_cla32_and3469_y0;
  wire h_u_cla32_and3470_y0;
  wire h_u_cla32_and3471_y0;
  wire h_u_cla32_and3472_y0;
  wire h_u_cla32_and3473_y0;
  wire h_u_cla32_and3474_y0;
  wire h_u_cla32_and3475_y0;
  wire h_u_cla32_and3476_y0;
  wire h_u_cla32_and3477_y0;
  wire h_u_cla32_and3478_y0;
  wire h_u_cla32_and3479_y0;
  wire h_u_cla32_and3480_y0;
  wire h_u_cla32_and3481_y0;
  wire h_u_cla32_and3482_y0;
  wire h_u_cla32_and3483_y0;
  wire h_u_cla32_and3484_y0;
  wire h_u_cla32_and3485_y0;
  wire h_u_cla32_and3486_y0;
  wire h_u_cla32_and3487_y0;
  wire h_u_cla32_and3488_y0;
  wire h_u_cla32_and3489_y0;
  wire h_u_cla32_and3490_y0;
  wire h_u_cla32_and3491_y0;
  wire h_u_cla32_and3492_y0;
  wire h_u_cla32_and3493_y0;
  wire h_u_cla32_and3494_y0;
  wire h_u_cla32_and3495_y0;
  wire h_u_cla32_and3496_y0;
  wire h_u_cla32_and3497_y0;
  wire h_u_cla32_and3498_y0;
  wire h_u_cla32_and3499_y0;
  wire h_u_cla32_and3500_y0;
  wire h_u_cla32_and3501_y0;
  wire h_u_cla32_and3502_y0;
  wire h_u_cla32_and3503_y0;
  wire h_u_cla32_and3504_y0;
  wire h_u_cla32_and3505_y0;
  wire h_u_cla32_and3506_y0;
  wire h_u_cla32_and3507_y0;
  wire h_u_cla32_and3508_y0;
  wire h_u_cla32_and3509_y0;
  wire h_u_cla32_and3510_y0;
  wire h_u_cla32_and3511_y0;
  wire h_u_cla32_and3512_y0;
  wire h_u_cla32_and3513_y0;
  wire h_u_cla32_and3514_y0;
  wire h_u_cla32_and3515_y0;
  wire h_u_cla32_and3516_y0;
  wire h_u_cla32_and3517_y0;
  wire h_u_cla32_and3518_y0;
  wire h_u_cla32_and3519_y0;
  wire h_u_cla32_and3520_y0;
  wire h_u_cla32_and3521_y0;
  wire h_u_cla32_and3522_y0;
  wire h_u_cla32_and3523_y0;
  wire h_u_cla32_and3524_y0;
  wire h_u_cla32_and3525_y0;
  wire h_u_cla32_and3526_y0;
  wire h_u_cla32_and3527_y0;
  wire h_u_cla32_and3528_y0;
  wire h_u_cla32_and3529_y0;
  wire h_u_cla32_and3530_y0;
  wire h_u_cla32_and3531_y0;
  wire h_u_cla32_and3532_y0;
  wire h_u_cla32_and3533_y0;
  wire h_u_cla32_and3534_y0;
  wire h_u_cla32_and3535_y0;
  wire h_u_cla32_and3536_y0;
  wire h_u_cla32_and3537_y0;
  wire h_u_cla32_and3538_y0;
  wire h_u_cla32_and3539_y0;
  wire h_u_cla32_and3540_y0;
  wire h_u_cla32_and3541_y0;
  wire h_u_cla32_and3542_y0;
  wire h_u_cla32_and3543_y0;
  wire h_u_cla32_and3544_y0;
  wire h_u_cla32_and3545_y0;
  wire h_u_cla32_and3546_y0;
  wire h_u_cla32_and3547_y0;
  wire h_u_cla32_and3548_y0;
  wire h_u_cla32_and3549_y0;
  wire h_u_cla32_and3550_y0;
  wire h_u_cla32_and3551_y0;
  wire h_u_cla32_and3552_y0;
  wire h_u_cla32_and3553_y0;
  wire h_u_cla32_and3554_y0;
  wire h_u_cla32_and3555_y0;
  wire h_u_cla32_and3556_y0;
  wire h_u_cla32_and3557_y0;
  wire h_u_cla32_and3558_y0;
  wire h_u_cla32_and3559_y0;
  wire h_u_cla32_and3560_y0;
  wire h_u_cla32_and3561_y0;
  wire h_u_cla32_and3562_y0;
  wire h_u_cla32_and3563_y0;
  wire h_u_cla32_and3564_y0;
  wire h_u_cla32_and3565_y0;
  wire h_u_cla32_and3566_y0;
  wire h_u_cla32_and3567_y0;
  wire h_u_cla32_and3568_y0;
  wire h_u_cla32_and3569_y0;
  wire h_u_cla32_and3570_y0;
  wire h_u_cla32_and3571_y0;
  wire h_u_cla32_and3572_y0;
  wire h_u_cla32_and3573_y0;
  wire h_u_cla32_and3574_y0;
  wire h_u_cla32_and3575_y0;
  wire h_u_cla32_and3576_y0;
  wire h_u_cla32_and3577_y0;
  wire h_u_cla32_and3578_y0;
  wire h_u_cla32_and3579_y0;
  wire h_u_cla32_and3580_y0;
  wire h_u_cla32_and3581_y0;
  wire h_u_cla32_and3582_y0;
  wire h_u_cla32_and3583_y0;
  wire h_u_cla32_and3584_y0;
  wire h_u_cla32_and3585_y0;
  wire h_u_cla32_and3586_y0;
  wire h_u_cla32_and3587_y0;
  wire h_u_cla32_and3588_y0;
  wire h_u_cla32_and3589_y0;
  wire h_u_cla32_and3590_y0;
  wire h_u_cla32_and3591_y0;
  wire h_u_cla32_and3592_y0;
  wire h_u_cla32_and3593_y0;
  wire h_u_cla32_and3594_y0;
  wire h_u_cla32_and3595_y0;
  wire h_u_cla32_and3596_y0;
  wire h_u_cla32_and3597_y0;
  wire h_u_cla32_and3598_y0;
  wire h_u_cla32_and3599_y0;
  wire h_u_cla32_and3600_y0;
  wire h_u_cla32_and3601_y0;
  wire h_u_cla32_and3602_y0;
  wire h_u_cla32_and3603_y0;
  wire h_u_cla32_and3604_y0;
  wire h_u_cla32_and3605_y0;
  wire h_u_cla32_and3606_y0;
  wire h_u_cla32_and3607_y0;
  wire h_u_cla32_and3608_y0;
  wire h_u_cla32_and3609_y0;
  wire h_u_cla32_and3610_y0;
  wire h_u_cla32_and3611_y0;
  wire h_u_cla32_and3612_y0;
  wire h_u_cla32_and3613_y0;
  wire h_u_cla32_and3614_y0;
  wire h_u_cla32_and3615_y0;
  wire h_u_cla32_and3616_y0;
  wire h_u_cla32_and3617_y0;
  wire h_u_cla32_and3618_y0;
  wire h_u_cla32_and3619_y0;
  wire h_u_cla32_and3620_y0;
  wire h_u_cla32_and3621_y0;
  wire h_u_cla32_and3622_y0;
  wire h_u_cla32_and3623_y0;
  wire h_u_cla32_and3624_y0;
  wire h_u_cla32_and3625_y0;
  wire h_u_cla32_and3626_y0;
  wire h_u_cla32_and3627_y0;
  wire h_u_cla32_and3628_y0;
  wire h_u_cla32_and3629_y0;
  wire h_u_cla32_and3630_y0;
  wire h_u_cla32_and3631_y0;
  wire h_u_cla32_and3632_y0;
  wire h_u_cla32_and3633_y0;
  wire h_u_cla32_and3634_y0;
  wire h_u_cla32_and3635_y0;
  wire h_u_cla32_and3636_y0;
  wire h_u_cla32_and3637_y0;
  wire h_u_cla32_and3638_y0;
  wire h_u_cla32_and3639_y0;
  wire h_u_cla32_and3640_y0;
  wire h_u_cla32_and3641_y0;
  wire h_u_cla32_and3642_y0;
  wire h_u_cla32_and3643_y0;
  wire h_u_cla32_and3644_y0;
  wire h_u_cla32_and3645_y0;
  wire h_u_cla32_and3646_y0;
  wire h_u_cla32_and3647_y0;
  wire h_u_cla32_and3648_y0;
  wire h_u_cla32_and3649_y0;
  wire h_u_cla32_and3650_y0;
  wire h_u_cla32_and3651_y0;
  wire h_u_cla32_and3652_y0;
  wire h_u_cla32_and3653_y0;
  wire h_u_cla32_and3654_y0;
  wire h_u_cla32_and3655_y0;
  wire h_u_cla32_and3656_y0;
  wire h_u_cla32_and3657_y0;
  wire h_u_cla32_and3658_y0;
  wire h_u_cla32_and3659_y0;
  wire h_u_cla32_and3660_y0;
  wire h_u_cla32_and3661_y0;
  wire h_u_cla32_and3662_y0;
  wire h_u_cla32_and3663_y0;
  wire h_u_cla32_and3664_y0;
  wire h_u_cla32_and3665_y0;
  wire h_u_cla32_and3666_y0;
  wire h_u_cla32_and3667_y0;
  wire h_u_cla32_and3668_y0;
  wire h_u_cla32_and3669_y0;
  wire h_u_cla32_and3670_y0;
  wire h_u_cla32_and3671_y0;
  wire h_u_cla32_and3672_y0;
  wire h_u_cla32_and3673_y0;
  wire h_u_cla32_and3674_y0;
  wire h_u_cla32_and3675_y0;
  wire h_u_cla32_and3676_y0;
  wire h_u_cla32_and3677_y0;
  wire h_u_cla32_and3678_y0;
  wire h_u_cla32_and3679_y0;
  wire h_u_cla32_and3680_y0;
  wire h_u_cla32_and3681_y0;
  wire h_u_cla32_and3682_y0;
  wire h_u_cla32_and3683_y0;
  wire h_u_cla32_and3684_y0;
  wire h_u_cla32_and3685_y0;
  wire h_u_cla32_and3686_y0;
  wire h_u_cla32_and3687_y0;
  wire h_u_cla32_and3688_y0;
  wire h_u_cla32_and3689_y0;
  wire h_u_cla32_and3690_y0;
  wire h_u_cla32_and3691_y0;
  wire h_u_cla32_and3692_y0;
  wire h_u_cla32_and3693_y0;
  wire h_u_cla32_and3694_y0;
  wire h_u_cla32_and3695_y0;
  wire h_u_cla32_and3696_y0;
  wire h_u_cla32_and3697_y0;
  wire h_u_cla32_and3698_y0;
  wire h_u_cla32_and3699_y0;
  wire h_u_cla32_and3700_y0;
  wire h_u_cla32_and3701_y0;
  wire h_u_cla32_and3702_y0;
  wire h_u_cla32_and3703_y0;
  wire h_u_cla32_and3704_y0;
  wire h_u_cla32_and3705_y0;
  wire h_u_cla32_and3706_y0;
  wire h_u_cla32_and3707_y0;
  wire h_u_cla32_and3708_y0;
  wire h_u_cla32_and3709_y0;
  wire h_u_cla32_and3710_y0;
  wire h_u_cla32_and3711_y0;
  wire h_u_cla32_and3712_y0;
  wire h_u_cla32_and3713_y0;
  wire h_u_cla32_and3714_y0;
  wire h_u_cla32_and3715_y0;
  wire h_u_cla32_and3716_y0;
  wire h_u_cla32_and3717_y0;
  wire h_u_cla32_and3718_y0;
  wire h_u_cla32_and3719_y0;
  wire h_u_cla32_and3720_y0;
  wire h_u_cla32_and3721_y0;
  wire h_u_cla32_and3722_y0;
  wire h_u_cla32_and3723_y0;
  wire h_u_cla32_and3724_y0;
  wire h_u_cla32_and3725_y0;
  wire h_u_cla32_and3726_y0;
  wire h_u_cla32_and3727_y0;
  wire h_u_cla32_and3728_y0;
  wire h_u_cla32_and3729_y0;
  wire h_u_cla32_and3730_y0;
  wire h_u_cla32_and3731_y0;
  wire h_u_cla32_and3732_y0;
  wire h_u_cla32_and3733_y0;
  wire h_u_cla32_and3734_y0;
  wire h_u_cla32_and3735_y0;
  wire h_u_cla32_and3736_y0;
  wire h_u_cla32_and3737_y0;
  wire h_u_cla32_and3738_y0;
  wire h_u_cla32_and3739_y0;
  wire h_u_cla32_and3740_y0;
  wire h_u_cla32_and3741_y0;
  wire h_u_cla32_and3742_y0;
  wire h_u_cla32_and3743_y0;
  wire h_u_cla32_and3744_y0;
  wire h_u_cla32_and3745_y0;
  wire h_u_cla32_and3746_y0;
  wire h_u_cla32_and3747_y0;
  wire h_u_cla32_and3748_y0;
  wire h_u_cla32_and3749_y0;
  wire h_u_cla32_and3750_y0;
  wire h_u_cla32_and3751_y0;
  wire h_u_cla32_and3752_y0;
  wire h_u_cla32_and3753_y0;
  wire h_u_cla32_and3754_y0;
  wire h_u_cla32_and3755_y0;
  wire h_u_cla32_and3756_y0;
  wire h_u_cla32_and3757_y0;
  wire h_u_cla32_and3758_y0;
  wire h_u_cla32_and3759_y0;
  wire h_u_cla32_and3760_y0;
  wire h_u_cla32_and3761_y0;
  wire h_u_cla32_and3762_y0;
  wire h_u_cla32_and3763_y0;
  wire h_u_cla32_and3764_y0;
  wire h_u_cla32_and3765_y0;
  wire h_u_cla32_and3766_y0;
  wire h_u_cla32_and3767_y0;
  wire h_u_cla32_and3768_y0;
  wire h_u_cla32_and3769_y0;
  wire h_u_cla32_and3770_y0;
  wire h_u_cla32_and3771_y0;
  wire h_u_cla32_and3772_y0;
  wire h_u_cla32_and3773_y0;
  wire h_u_cla32_and3774_y0;
  wire h_u_cla32_and3775_y0;
  wire h_u_cla32_and3776_y0;
  wire h_u_cla32_and3777_y0;
  wire h_u_cla32_and3778_y0;
  wire h_u_cla32_and3779_y0;
  wire h_u_cla32_and3780_y0;
  wire h_u_cla32_and3781_y0;
  wire h_u_cla32_and3782_y0;
  wire h_u_cla32_and3783_y0;
  wire h_u_cla32_and3784_y0;
  wire h_u_cla32_and3785_y0;
  wire h_u_cla32_and3786_y0;
  wire h_u_cla32_and3787_y0;
  wire h_u_cla32_and3788_y0;
  wire h_u_cla32_and3789_y0;
  wire h_u_cla32_and3790_y0;
  wire h_u_cla32_and3791_y0;
  wire h_u_cla32_and3792_y0;
  wire h_u_cla32_and3793_y0;
  wire h_u_cla32_and3794_y0;
  wire h_u_cla32_or231_y0;
  wire h_u_cla32_or232_y0;
  wire h_u_cla32_or233_y0;
  wire h_u_cla32_or234_y0;
  wire h_u_cla32_or235_y0;
  wire h_u_cla32_or236_y0;
  wire h_u_cla32_or237_y0;
  wire h_u_cla32_or238_y0;
  wire h_u_cla32_or239_y0;
  wire h_u_cla32_or240_y0;
  wire h_u_cla32_or241_y0;
  wire h_u_cla32_or242_y0;
  wire h_u_cla32_or243_y0;
  wire h_u_cla32_or244_y0;
  wire h_u_cla32_or245_y0;
  wire h_u_cla32_or246_y0;
  wire h_u_cla32_or247_y0;
  wire h_u_cla32_or248_y0;
  wire h_u_cla32_or249_y0;
  wire h_u_cla32_or250_y0;
  wire h_u_cla32_or251_y0;
  wire h_u_cla32_or252_y0;
  wire h_u_cla32_pg_logic22_y0;
  wire h_u_cla32_pg_logic22_y1;
  wire h_u_cla32_pg_logic22_y2;
  wire h_u_cla32_xor22_y0;
  wire h_u_cla32_and3795_y0;
  wire h_u_cla32_and3796_y0;
  wire h_u_cla32_and3797_y0;
  wire h_u_cla32_and3798_y0;
  wire h_u_cla32_and3799_y0;
  wire h_u_cla32_and3800_y0;
  wire h_u_cla32_and3801_y0;
  wire h_u_cla32_and3802_y0;
  wire h_u_cla32_and3803_y0;
  wire h_u_cla32_and3804_y0;
  wire h_u_cla32_and3805_y0;
  wire h_u_cla32_and3806_y0;
  wire h_u_cla32_and3807_y0;
  wire h_u_cla32_and3808_y0;
  wire h_u_cla32_and3809_y0;
  wire h_u_cla32_and3810_y0;
  wire h_u_cla32_and3811_y0;
  wire h_u_cla32_and3812_y0;
  wire h_u_cla32_and3813_y0;
  wire h_u_cla32_and3814_y0;
  wire h_u_cla32_and3815_y0;
  wire h_u_cla32_and3816_y0;
  wire h_u_cla32_and3817_y0;
  wire h_u_cla32_and3818_y0;
  wire h_u_cla32_and3819_y0;
  wire h_u_cla32_and3820_y0;
  wire h_u_cla32_and3821_y0;
  wire h_u_cla32_and3822_y0;
  wire h_u_cla32_and3823_y0;
  wire h_u_cla32_and3824_y0;
  wire h_u_cla32_and3825_y0;
  wire h_u_cla32_and3826_y0;
  wire h_u_cla32_and3827_y0;
  wire h_u_cla32_and3828_y0;
  wire h_u_cla32_and3829_y0;
  wire h_u_cla32_and3830_y0;
  wire h_u_cla32_and3831_y0;
  wire h_u_cla32_and3832_y0;
  wire h_u_cla32_and3833_y0;
  wire h_u_cla32_and3834_y0;
  wire h_u_cla32_and3835_y0;
  wire h_u_cla32_and3836_y0;
  wire h_u_cla32_and3837_y0;
  wire h_u_cla32_and3838_y0;
  wire h_u_cla32_and3839_y0;
  wire h_u_cla32_and3840_y0;
  wire h_u_cla32_and3841_y0;
  wire h_u_cla32_and3842_y0;
  wire h_u_cla32_and3843_y0;
  wire h_u_cla32_and3844_y0;
  wire h_u_cla32_and3845_y0;
  wire h_u_cla32_and3846_y0;
  wire h_u_cla32_and3847_y0;
  wire h_u_cla32_and3848_y0;
  wire h_u_cla32_and3849_y0;
  wire h_u_cla32_and3850_y0;
  wire h_u_cla32_and3851_y0;
  wire h_u_cla32_and3852_y0;
  wire h_u_cla32_and3853_y0;
  wire h_u_cla32_and3854_y0;
  wire h_u_cla32_and3855_y0;
  wire h_u_cla32_and3856_y0;
  wire h_u_cla32_and3857_y0;
  wire h_u_cla32_and3858_y0;
  wire h_u_cla32_and3859_y0;
  wire h_u_cla32_and3860_y0;
  wire h_u_cla32_and3861_y0;
  wire h_u_cla32_and3862_y0;
  wire h_u_cla32_and3863_y0;
  wire h_u_cla32_and3864_y0;
  wire h_u_cla32_and3865_y0;
  wire h_u_cla32_and3866_y0;
  wire h_u_cla32_and3867_y0;
  wire h_u_cla32_and3868_y0;
  wire h_u_cla32_and3869_y0;
  wire h_u_cla32_and3870_y0;
  wire h_u_cla32_and3871_y0;
  wire h_u_cla32_and3872_y0;
  wire h_u_cla32_and3873_y0;
  wire h_u_cla32_and3874_y0;
  wire h_u_cla32_and3875_y0;
  wire h_u_cla32_and3876_y0;
  wire h_u_cla32_and3877_y0;
  wire h_u_cla32_and3878_y0;
  wire h_u_cla32_and3879_y0;
  wire h_u_cla32_and3880_y0;
  wire h_u_cla32_and3881_y0;
  wire h_u_cla32_and3882_y0;
  wire h_u_cla32_and3883_y0;
  wire h_u_cla32_and3884_y0;
  wire h_u_cla32_and3885_y0;
  wire h_u_cla32_and3886_y0;
  wire h_u_cla32_and3887_y0;
  wire h_u_cla32_and3888_y0;
  wire h_u_cla32_and3889_y0;
  wire h_u_cla32_and3890_y0;
  wire h_u_cla32_and3891_y0;
  wire h_u_cla32_and3892_y0;
  wire h_u_cla32_and3893_y0;
  wire h_u_cla32_and3894_y0;
  wire h_u_cla32_and3895_y0;
  wire h_u_cla32_and3896_y0;
  wire h_u_cla32_and3897_y0;
  wire h_u_cla32_and3898_y0;
  wire h_u_cla32_and3899_y0;
  wire h_u_cla32_and3900_y0;
  wire h_u_cla32_and3901_y0;
  wire h_u_cla32_and3902_y0;
  wire h_u_cla32_and3903_y0;
  wire h_u_cla32_and3904_y0;
  wire h_u_cla32_and3905_y0;
  wire h_u_cla32_and3906_y0;
  wire h_u_cla32_and3907_y0;
  wire h_u_cla32_and3908_y0;
  wire h_u_cla32_and3909_y0;
  wire h_u_cla32_and3910_y0;
  wire h_u_cla32_and3911_y0;
  wire h_u_cla32_and3912_y0;
  wire h_u_cla32_and3913_y0;
  wire h_u_cla32_and3914_y0;
  wire h_u_cla32_and3915_y0;
  wire h_u_cla32_and3916_y0;
  wire h_u_cla32_and3917_y0;
  wire h_u_cla32_and3918_y0;
  wire h_u_cla32_and3919_y0;
  wire h_u_cla32_and3920_y0;
  wire h_u_cla32_and3921_y0;
  wire h_u_cla32_and3922_y0;
  wire h_u_cla32_and3923_y0;
  wire h_u_cla32_and3924_y0;
  wire h_u_cla32_and3925_y0;
  wire h_u_cla32_and3926_y0;
  wire h_u_cla32_and3927_y0;
  wire h_u_cla32_and3928_y0;
  wire h_u_cla32_and3929_y0;
  wire h_u_cla32_and3930_y0;
  wire h_u_cla32_and3931_y0;
  wire h_u_cla32_and3932_y0;
  wire h_u_cla32_and3933_y0;
  wire h_u_cla32_and3934_y0;
  wire h_u_cla32_and3935_y0;
  wire h_u_cla32_and3936_y0;
  wire h_u_cla32_and3937_y0;
  wire h_u_cla32_and3938_y0;
  wire h_u_cla32_and3939_y0;
  wire h_u_cla32_and3940_y0;
  wire h_u_cla32_and3941_y0;
  wire h_u_cla32_and3942_y0;
  wire h_u_cla32_and3943_y0;
  wire h_u_cla32_and3944_y0;
  wire h_u_cla32_and3945_y0;
  wire h_u_cla32_and3946_y0;
  wire h_u_cla32_and3947_y0;
  wire h_u_cla32_and3948_y0;
  wire h_u_cla32_and3949_y0;
  wire h_u_cla32_and3950_y0;
  wire h_u_cla32_and3951_y0;
  wire h_u_cla32_and3952_y0;
  wire h_u_cla32_and3953_y0;
  wire h_u_cla32_and3954_y0;
  wire h_u_cla32_and3955_y0;
  wire h_u_cla32_and3956_y0;
  wire h_u_cla32_and3957_y0;
  wire h_u_cla32_and3958_y0;
  wire h_u_cla32_and3959_y0;
  wire h_u_cla32_and3960_y0;
  wire h_u_cla32_and3961_y0;
  wire h_u_cla32_and3962_y0;
  wire h_u_cla32_and3963_y0;
  wire h_u_cla32_and3964_y0;
  wire h_u_cla32_and3965_y0;
  wire h_u_cla32_and3966_y0;
  wire h_u_cla32_and3967_y0;
  wire h_u_cla32_and3968_y0;
  wire h_u_cla32_and3969_y0;
  wire h_u_cla32_and3970_y0;
  wire h_u_cla32_and3971_y0;
  wire h_u_cla32_and3972_y0;
  wire h_u_cla32_and3973_y0;
  wire h_u_cla32_and3974_y0;
  wire h_u_cla32_and3975_y0;
  wire h_u_cla32_and3976_y0;
  wire h_u_cla32_and3977_y0;
  wire h_u_cla32_and3978_y0;
  wire h_u_cla32_and3979_y0;
  wire h_u_cla32_and3980_y0;
  wire h_u_cla32_and3981_y0;
  wire h_u_cla32_and3982_y0;
  wire h_u_cla32_and3983_y0;
  wire h_u_cla32_and3984_y0;
  wire h_u_cla32_and3985_y0;
  wire h_u_cla32_and3986_y0;
  wire h_u_cla32_and3987_y0;
  wire h_u_cla32_and3988_y0;
  wire h_u_cla32_and3989_y0;
  wire h_u_cla32_and3990_y0;
  wire h_u_cla32_and3991_y0;
  wire h_u_cla32_and3992_y0;
  wire h_u_cla32_and3993_y0;
  wire h_u_cla32_and3994_y0;
  wire h_u_cla32_and3995_y0;
  wire h_u_cla32_and3996_y0;
  wire h_u_cla32_and3997_y0;
  wire h_u_cla32_and3998_y0;
  wire h_u_cla32_and3999_y0;
  wire h_u_cla32_and4000_y0;
  wire h_u_cla32_and4001_y0;
  wire h_u_cla32_and4002_y0;
  wire h_u_cla32_and4003_y0;
  wire h_u_cla32_and4004_y0;
  wire h_u_cla32_and4005_y0;
  wire h_u_cla32_and4006_y0;
  wire h_u_cla32_and4007_y0;
  wire h_u_cla32_and4008_y0;
  wire h_u_cla32_and4009_y0;
  wire h_u_cla32_and4010_y0;
  wire h_u_cla32_and4011_y0;
  wire h_u_cla32_and4012_y0;
  wire h_u_cla32_and4013_y0;
  wire h_u_cla32_and4014_y0;
  wire h_u_cla32_and4015_y0;
  wire h_u_cla32_and4016_y0;
  wire h_u_cla32_and4017_y0;
  wire h_u_cla32_and4018_y0;
  wire h_u_cla32_and4019_y0;
  wire h_u_cla32_and4020_y0;
  wire h_u_cla32_and4021_y0;
  wire h_u_cla32_and4022_y0;
  wire h_u_cla32_and4023_y0;
  wire h_u_cla32_and4024_y0;
  wire h_u_cla32_and4025_y0;
  wire h_u_cla32_and4026_y0;
  wire h_u_cla32_and4027_y0;
  wire h_u_cla32_and4028_y0;
  wire h_u_cla32_and4029_y0;
  wire h_u_cla32_and4030_y0;
  wire h_u_cla32_and4031_y0;
  wire h_u_cla32_and4032_y0;
  wire h_u_cla32_and4033_y0;
  wire h_u_cla32_and4034_y0;
  wire h_u_cla32_and4035_y0;
  wire h_u_cla32_and4036_y0;
  wire h_u_cla32_and4037_y0;
  wire h_u_cla32_and4038_y0;
  wire h_u_cla32_and4039_y0;
  wire h_u_cla32_and4040_y0;
  wire h_u_cla32_and4041_y0;
  wire h_u_cla32_and4042_y0;
  wire h_u_cla32_and4043_y0;
  wire h_u_cla32_and4044_y0;
  wire h_u_cla32_and4045_y0;
  wire h_u_cla32_and4046_y0;
  wire h_u_cla32_and4047_y0;
  wire h_u_cla32_and4048_y0;
  wire h_u_cla32_and4049_y0;
  wire h_u_cla32_and4050_y0;
  wire h_u_cla32_and4051_y0;
  wire h_u_cla32_and4052_y0;
  wire h_u_cla32_and4053_y0;
  wire h_u_cla32_and4054_y0;
  wire h_u_cla32_and4055_y0;
  wire h_u_cla32_and4056_y0;
  wire h_u_cla32_and4057_y0;
  wire h_u_cla32_and4058_y0;
  wire h_u_cla32_and4059_y0;
  wire h_u_cla32_and4060_y0;
  wire h_u_cla32_and4061_y0;
  wire h_u_cla32_and4062_y0;
  wire h_u_cla32_and4063_y0;
  wire h_u_cla32_and4064_y0;
  wire h_u_cla32_and4065_y0;
  wire h_u_cla32_and4066_y0;
  wire h_u_cla32_and4067_y0;
  wire h_u_cla32_and4068_y0;
  wire h_u_cla32_and4069_y0;
  wire h_u_cla32_and4070_y0;
  wire h_u_cla32_and4071_y0;
  wire h_u_cla32_and4072_y0;
  wire h_u_cla32_and4073_y0;
  wire h_u_cla32_and4074_y0;
  wire h_u_cla32_and4075_y0;
  wire h_u_cla32_and4076_y0;
  wire h_u_cla32_and4077_y0;
  wire h_u_cla32_and4078_y0;
  wire h_u_cla32_and4079_y0;
  wire h_u_cla32_and4080_y0;
  wire h_u_cla32_and4081_y0;
  wire h_u_cla32_and4082_y0;
  wire h_u_cla32_and4083_y0;
  wire h_u_cla32_and4084_y0;
  wire h_u_cla32_and4085_y0;
  wire h_u_cla32_and4086_y0;
  wire h_u_cla32_and4087_y0;
  wire h_u_cla32_and4088_y0;
  wire h_u_cla32_and4089_y0;
  wire h_u_cla32_and4090_y0;
  wire h_u_cla32_and4091_y0;
  wire h_u_cla32_and4092_y0;
  wire h_u_cla32_and4093_y0;
  wire h_u_cla32_and4094_y0;
  wire h_u_cla32_and4095_y0;
  wire h_u_cla32_and4096_y0;
  wire h_u_cla32_and4097_y0;
  wire h_u_cla32_and4098_y0;
  wire h_u_cla32_and4099_y0;
  wire h_u_cla32_and4100_y0;
  wire h_u_cla32_and4101_y0;
  wire h_u_cla32_and4102_y0;
  wire h_u_cla32_and4103_y0;
  wire h_u_cla32_and4104_y0;
  wire h_u_cla32_and4105_y0;
  wire h_u_cla32_and4106_y0;
  wire h_u_cla32_and4107_y0;
  wire h_u_cla32_and4108_y0;
  wire h_u_cla32_and4109_y0;
  wire h_u_cla32_and4110_y0;
  wire h_u_cla32_and4111_y0;
  wire h_u_cla32_and4112_y0;
  wire h_u_cla32_and4113_y0;
  wire h_u_cla32_and4114_y0;
  wire h_u_cla32_and4115_y0;
  wire h_u_cla32_and4116_y0;
  wire h_u_cla32_and4117_y0;
  wire h_u_cla32_and4118_y0;
  wire h_u_cla32_and4119_y0;
  wire h_u_cla32_and4120_y0;
  wire h_u_cla32_and4121_y0;
  wire h_u_cla32_and4122_y0;
  wire h_u_cla32_and4123_y0;
  wire h_u_cla32_and4124_y0;
  wire h_u_cla32_and4125_y0;
  wire h_u_cla32_and4126_y0;
  wire h_u_cla32_and4127_y0;
  wire h_u_cla32_and4128_y0;
  wire h_u_cla32_and4129_y0;
  wire h_u_cla32_and4130_y0;
  wire h_u_cla32_and4131_y0;
  wire h_u_cla32_and4132_y0;
  wire h_u_cla32_and4133_y0;
  wire h_u_cla32_and4134_y0;
  wire h_u_cla32_and4135_y0;
  wire h_u_cla32_and4136_y0;
  wire h_u_cla32_and4137_y0;
  wire h_u_cla32_and4138_y0;
  wire h_u_cla32_and4139_y0;
  wire h_u_cla32_and4140_y0;
  wire h_u_cla32_and4141_y0;
  wire h_u_cla32_and4142_y0;
  wire h_u_cla32_and4143_y0;
  wire h_u_cla32_and4144_y0;
  wire h_u_cla32_and4145_y0;
  wire h_u_cla32_and4146_y0;
  wire h_u_cla32_and4147_y0;
  wire h_u_cla32_and4148_y0;
  wire h_u_cla32_and4149_y0;
  wire h_u_cla32_and4150_y0;
  wire h_u_cla32_and4151_y0;
  wire h_u_cla32_and4152_y0;
  wire h_u_cla32_and4153_y0;
  wire h_u_cla32_and4154_y0;
  wire h_u_cla32_and4155_y0;
  wire h_u_cla32_and4156_y0;
  wire h_u_cla32_and4157_y0;
  wire h_u_cla32_and4158_y0;
  wire h_u_cla32_and4159_y0;
  wire h_u_cla32_and4160_y0;
  wire h_u_cla32_and4161_y0;
  wire h_u_cla32_and4162_y0;
  wire h_u_cla32_and4163_y0;
  wire h_u_cla32_and4164_y0;
  wire h_u_cla32_and4165_y0;
  wire h_u_cla32_and4166_y0;
  wire h_u_cla32_and4167_y0;
  wire h_u_cla32_and4168_y0;
  wire h_u_cla32_and4169_y0;
  wire h_u_cla32_and4170_y0;
  wire h_u_cla32_and4171_y0;
  wire h_u_cla32_and4172_y0;
  wire h_u_cla32_and4173_y0;
  wire h_u_cla32_and4174_y0;
  wire h_u_cla32_and4175_y0;
  wire h_u_cla32_and4176_y0;
  wire h_u_cla32_and4177_y0;
  wire h_u_cla32_and4178_y0;
  wire h_u_cla32_and4179_y0;
  wire h_u_cla32_and4180_y0;
  wire h_u_cla32_and4181_y0;
  wire h_u_cla32_and4182_y0;
  wire h_u_cla32_and4183_y0;
  wire h_u_cla32_and4184_y0;
  wire h_u_cla32_and4185_y0;
  wire h_u_cla32_and4186_y0;
  wire h_u_cla32_and4187_y0;
  wire h_u_cla32_and4188_y0;
  wire h_u_cla32_and4189_y0;
  wire h_u_cla32_and4190_y0;
  wire h_u_cla32_and4191_y0;
  wire h_u_cla32_and4192_y0;
  wire h_u_cla32_and4193_y0;
  wire h_u_cla32_and4194_y0;
  wire h_u_cla32_and4195_y0;
  wire h_u_cla32_and4196_y0;
  wire h_u_cla32_and4197_y0;
  wire h_u_cla32_and4198_y0;
  wire h_u_cla32_and4199_y0;
  wire h_u_cla32_and4200_y0;
  wire h_u_cla32_and4201_y0;
  wire h_u_cla32_and4202_y0;
  wire h_u_cla32_and4203_y0;
  wire h_u_cla32_and4204_y0;
  wire h_u_cla32_and4205_y0;
  wire h_u_cla32_and4206_y0;
  wire h_u_cla32_and4207_y0;
  wire h_u_cla32_and4208_y0;
  wire h_u_cla32_and4209_y0;
  wire h_u_cla32_and4210_y0;
  wire h_u_cla32_and4211_y0;
  wire h_u_cla32_and4212_y0;
  wire h_u_cla32_and4213_y0;
  wire h_u_cla32_and4214_y0;
  wire h_u_cla32_and4215_y0;
  wire h_u_cla32_and4216_y0;
  wire h_u_cla32_and4217_y0;
  wire h_u_cla32_and4218_y0;
  wire h_u_cla32_and4219_y0;
  wire h_u_cla32_and4220_y0;
  wire h_u_cla32_and4221_y0;
  wire h_u_cla32_and4222_y0;
  wire h_u_cla32_and4223_y0;
  wire h_u_cla32_and4224_y0;
  wire h_u_cla32_and4225_y0;
  wire h_u_cla32_and4226_y0;
  wire h_u_cla32_and4227_y0;
  wire h_u_cla32_and4228_y0;
  wire h_u_cla32_and4229_y0;
  wire h_u_cla32_and4230_y0;
  wire h_u_cla32_and4231_y0;
  wire h_u_cla32_and4232_y0;
  wire h_u_cla32_and4233_y0;
  wire h_u_cla32_and4234_y0;
  wire h_u_cla32_and4235_y0;
  wire h_u_cla32_and4236_y0;
  wire h_u_cla32_and4237_y0;
  wire h_u_cla32_and4238_y0;
  wire h_u_cla32_and4239_y0;
  wire h_u_cla32_and4240_y0;
  wire h_u_cla32_and4241_y0;
  wire h_u_cla32_and4242_y0;
  wire h_u_cla32_and4243_y0;
  wire h_u_cla32_and4244_y0;
  wire h_u_cla32_and4245_y0;
  wire h_u_cla32_and4246_y0;
  wire h_u_cla32_and4247_y0;
  wire h_u_cla32_and4248_y0;
  wire h_u_cla32_and4249_y0;
  wire h_u_cla32_and4250_y0;
  wire h_u_cla32_and4251_y0;
  wire h_u_cla32_and4252_y0;
  wire h_u_cla32_and4253_y0;
  wire h_u_cla32_and4254_y0;
  wire h_u_cla32_and4255_y0;
  wire h_u_cla32_and4256_y0;
  wire h_u_cla32_and4257_y0;
  wire h_u_cla32_and4258_y0;
  wire h_u_cla32_and4259_y0;
  wire h_u_cla32_and4260_y0;
  wire h_u_cla32_and4261_y0;
  wire h_u_cla32_and4262_y0;
  wire h_u_cla32_and4263_y0;
  wire h_u_cla32_and4264_y0;
  wire h_u_cla32_and4265_y0;
  wire h_u_cla32_and4266_y0;
  wire h_u_cla32_and4267_y0;
  wire h_u_cla32_and4268_y0;
  wire h_u_cla32_and4269_y0;
  wire h_u_cla32_and4270_y0;
  wire h_u_cla32_and4271_y0;
  wire h_u_cla32_and4272_y0;
  wire h_u_cla32_and4273_y0;
  wire h_u_cla32_and4274_y0;
  wire h_u_cla32_and4275_y0;
  wire h_u_cla32_and4276_y0;
  wire h_u_cla32_and4277_y0;
  wire h_u_cla32_and4278_y0;
  wire h_u_cla32_and4279_y0;
  wire h_u_cla32_and4280_y0;
  wire h_u_cla32_and4281_y0;
  wire h_u_cla32_and4282_y0;
  wire h_u_cla32_and4283_y0;
  wire h_u_cla32_and4284_y0;
  wire h_u_cla32_and4285_y0;
  wire h_u_cla32_and4286_y0;
  wire h_u_cla32_and4287_y0;
  wire h_u_cla32_and4288_y0;
  wire h_u_cla32_and4289_y0;
  wire h_u_cla32_and4290_y0;
  wire h_u_cla32_and4291_y0;
  wire h_u_cla32_and4292_y0;
  wire h_u_cla32_and4293_y0;
  wire h_u_cla32_and4294_y0;
  wire h_u_cla32_and4295_y0;
  wire h_u_cla32_and4296_y0;
  wire h_u_cla32_and4297_y0;
  wire h_u_cla32_and4298_y0;
  wire h_u_cla32_and4299_y0;
  wire h_u_cla32_and4300_y0;
  wire h_u_cla32_and4301_y0;
  wire h_u_cla32_and4302_y0;
  wire h_u_cla32_and4303_y0;
  wire h_u_cla32_and4304_y0;
  wire h_u_cla32_and4305_y0;
  wire h_u_cla32_and4306_y0;
  wire h_u_cla32_and4307_y0;
  wire h_u_cla32_and4308_y0;
  wire h_u_cla32_and4309_y0;
  wire h_u_cla32_and4310_y0;
  wire h_u_cla32_and4311_y0;
  wire h_u_cla32_and4312_y0;
  wire h_u_cla32_and4313_y0;
  wire h_u_cla32_and4314_y0;
  wire h_u_cla32_and4315_y0;
  wire h_u_cla32_and4316_y0;
  wire h_u_cla32_and4317_y0;
  wire h_u_cla32_and4318_y0;
  wire h_u_cla32_and4319_y0;
  wire h_u_cla32_and4320_y0;
  wire h_u_cla32_and4321_y0;
  wire h_u_cla32_and4322_y0;
  wire h_u_cla32_and4323_y0;
  wire h_u_cla32_or253_y0;
  wire h_u_cla32_or254_y0;
  wire h_u_cla32_or255_y0;
  wire h_u_cla32_or256_y0;
  wire h_u_cla32_or257_y0;
  wire h_u_cla32_or258_y0;
  wire h_u_cla32_or259_y0;
  wire h_u_cla32_or260_y0;
  wire h_u_cla32_or261_y0;
  wire h_u_cla32_or262_y0;
  wire h_u_cla32_or263_y0;
  wire h_u_cla32_or264_y0;
  wire h_u_cla32_or265_y0;
  wire h_u_cla32_or266_y0;
  wire h_u_cla32_or267_y0;
  wire h_u_cla32_or268_y0;
  wire h_u_cla32_or269_y0;
  wire h_u_cla32_or270_y0;
  wire h_u_cla32_or271_y0;
  wire h_u_cla32_or272_y0;
  wire h_u_cla32_or273_y0;
  wire h_u_cla32_or274_y0;
  wire h_u_cla32_or275_y0;
  wire h_u_cla32_pg_logic23_y0;
  wire h_u_cla32_pg_logic23_y1;
  wire h_u_cla32_pg_logic23_y2;
  wire h_u_cla32_xor23_y0;
  wire h_u_cla32_and4324_y0;
  wire h_u_cla32_and4325_y0;
  wire h_u_cla32_and4326_y0;
  wire h_u_cla32_and4327_y0;
  wire h_u_cla32_and4328_y0;
  wire h_u_cla32_and4329_y0;
  wire h_u_cla32_and4330_y0;
  wire h_u_cla32_and4331_y0;
  wire h_u_cla32_and4332_y0;
  wire h_u_cla32_and4333_y0;
  wire h_u_cla32_and4334_y0;
  wire h_u_cla32_and4335_y0;
  wire h_u_cla32_and4336_y0;
  wire h_u_cla32_and4337_y0;
  wire h_u_cla32_and4338_y0;
  wire h_u_cla32_and4339_y0;
  wire h_u_cla32_and4340_y0;
  wire h_u_cla32_and4341_y0;
  wire h_u_cla32_and4342_y0;
  wire h_u_cla32_and4343_y0;
  wire h_u_cla32_and4344_y0;
  wire h_u_cla32_and4345_y0;
  wire h_u_cla32_and4346_y0;
  wire h_u_cla32_and4347_y0;
  wire h_u_cla32_and4348_y0;
  wire h_u_cla32_and4349_y0;
  wire h_u_cla32_and4350_y0;
  wire h_u_cla32_and4351_y0;
  wire h_u_cla32_and4352_y0;
  wire h_u_cla32_and4353_y0;
  wire h_u_cla32_and4354_y0;
  wire h_u_cla32_and4355_y0;
  wire h_u_cla32_and4356_y0;
  wire h_u_cla32_and4357_y0;
  wire h_u_cla32_and4358_y0;
  wire h_u_cla32_and4359_y0;
  wire h_u_cla32_and4360_y0;
  wire h_u_cla32_and4361_y0;
  wire h_u_cla32_and4362_y0;
  wire h_u_cla32_and4363_y0;
  wire h_u_cla32_and4364_y0;
  wire h_u_cla32_and4365_y0;
  wire h_u_cla32_and4366_y0;
  wire h_u_cla32_and4367_y0;
  wire h_u_cla32_and4368_y0;
  wire h_u_cla32_and4369_y0;
  wire h_u_cla32_and4370_y0;
  wire h_u_cla32_and4371_y0;
  wire h_u_cla32_and4372_y0;
  wire h_u_cla32_and4373_y0;
  wire h_u_cla32_and4374_y0;
  wire h_u_cla32_and4375_y0;
  wire h_u_cla32_and4376_y0;
  wire h_u_cla32_and4377_y0;
  wire h_u_cla32_and4378_y0;
  wire h_u_cla32_and4379_y0;
  wire h_u_cla32_and4380_y0;
  wire h_u_cla32_and4381_y0;
  wire h_u_cla32_and4382_y0;
  wire h_u_cla32_and4383_y0;
  wire h_u_cla32_and4384_y0;
  wire h_u_cla32_and4385_y0;
  wire h_u_cla32_and4386_y0;
  wire h_u_cla32_and4387_y0;
  wire h_u_cla32_and4388_y0;
  wire h_u_cla32_and4389_y0;
  wire h_u_cla32_and4390_y0;
  wire h_u_cla32_and4391_y0;
  wire h_u_cla32_and4392_y0;
  wire h_u_cla32_and4393_y0;
  wire h_u_cla32_and4394_y0;
  wire h_u_cla32_and4395_y0;
  wire h_u_cla32_and4396_y0;
  wire h_u_cla32_and4397_y0;
  wire h_u_cla32_and4398_y0;
  wire h_u_cla32_and4399_y0;
  wire h_u_cla32_and4400_y0;
  wire h_u_cla32_and4401_y0;
  wire h_u_cla32_and4402_y0;
  wire h_u_cla32_and4403_y0;
  wire h_u_cla32_and4404_y0;
  wire h_u_cla32_and4405_y0;
  wire h_u_cla32_and4406_y0;
  wire h_u_cla32_and4407_y0;
  wire h_u_cla32_and4408_y0;
  wire h_u_cla32_and4409_y0;
  wire h_u_cla32_and4410_y0;
  wire h_u_cla32_and4411_y0;
  wire h_u_cla32_and4412_y0;
  wire h_u_cla32_and4413_y0;
  wire h_u_cla32_and4414_y0;
  wire h_u_cla32_and4415_y0;
  wire h_u_cla32_and4416_y0;
  wire h_u_cla32_and4417_y0;
  wire h_u_cla32_and4418_y0;
  wire h_u_cla32_and4419_y0;
  wire h_u_cla32_and4420_y0;
  wire h_u_cla32_and4421_y0;
  wire h_u_cla32_and4422_y0;
  wire h_u_cla32_and4423_y0;
  wire h_u_cla32_and4424_y0;
  wire h_u_cla32_and4425_y0;
  wire h_u_cla32_and4426_y0;
  wire h_u_cla32_and4427_y0;
  wire h_u_cla32_and4428_y0;
  wire h_u_cla32_and4429_y0;
  wire h_u_cla32_and4430_y0;
  wire h_u_cla32_and4431_y0;
  wire h_u_cla32_and4432_y0;
  wire h_u_cla32_and4433_y0;
  wire h_u_cla32_and4434_y0;
  wire h_u_cla32_and4435_y0;
  wire h_u_cla32_and4436_y0;
  wire h_u_cla32_and4437_y0;
  wire h_u_cla32_and4438_y0;
  wire h_u_cla32_and4439_y0;
  wire h_u_cla32_and4440_y0;
  wire h_u_cla32_and4441_y0;
  wire h_u_cla32_and4442_y0;
  wire h_u_cla32_and4443_y0;
  wire h_u_cla32_and4444_y0;
  wire h_u_cla32_and4445_y0;
  wire h_u_cla32_and4446_y0;
  wire h_u_cla32_and4447_y0;
  wire h_u_cla32_and4448_y0;
  wire h_u_cla32_and4449_y0;
  wire h_u_cla32_and4450_y0;
  wire h_u_cla32_and4451_y0;
  wire h_u_cla32_and4452_y0;
  wire h_u_cla32_and4453_y0;
  wire h_u_cla32_and4454_y0;
  wire h_u_cla32_and4455_y0;
  wire h_u_cla32_and4456_y0;
  wire h_u_cla32_and4457_y0;
  wire h_u_cla32_and4458_y0;
  wire h_u_cla32_and4459_y0;
  wire h_u_cla32_and4460_y0;
  wire h_u_cla32_and4461_y0;
  wire h_u_cla32_and4462_y0;
  wire h_u_cla32_and4463_y0;
  wire h_u_cla32_and4464_y0;
  wire h_u_cla32_and4465_y0;
  wire h_u_cla32_and4466_y0;
  wire h_u_cla32_and4467_y0;
  wire h_u_cla32_and4468_y0;
  wire h_u_cla32_and4469_y0;
  wire h_u_cla32_and4470_y0;
  wire h_u_cla32_and4471_y0;
  wire h_u_cla32_and4472_y0;
  wire h_u_cla32_and4473_y0;
  wire h_u_cla32_and4474_y0;
  wire h_u_cla32_and4475_y0;
  wire h_u_cla32_and4476_y0;
  wire h_u_cla32_and4477_y0;
  wire h_u_cla32_and4478_y0;
  wire h_u_cla32_and4479_y0;
  wire h_u_cla32_and4480_y0;
  wire h_u_cla32_and4481_y0;
  wire h_u_cla32_and4482_y0;
  wire h_u_cla32_and4483_y0;
  wire h_u_cla32_and4484_y0;
  wire h_u_cla32_and4485_y0;
  wire h_u_cla32_and4486_y0;
  wire h_u_cla32_and4487_y0;
  wire h_u_cla32_and4488_y0;
  wire h_u_cla32_and4489_y0;
  wire h_u_cla32_and4490_y0;
  wire h_u_cla32_and4491_y0;
  wire h_u_cla32_and4492_y0;
  wire h_u_cla32_and4493_y0;
  wire h_u_cla32_and4494_y0;
  wire h_u_cla32_and4495_y0;
  wire h_u_cla32_and4496_y0;
  wire h_u_cla32_and4497_y0;
  wire h_u_cla32_and4498_y0;
  wire h_u_cla32_and4499_y0;
  wire h_u_cla32_and4500_y0;
  wire h_u_cla32_and4501_y0;
  wire h_u_cla32_and4502_y0;
  wire h_u_cla32_and4503_y0;
  wire h_u_cla32_and4504_y0;
  wire h_u_cla32_and4505_y0;
  wire h_u_cla32_and4506_y0;
  wire h_u_cla32_and4507_y0;
  wire h_u_cla32_and4508_y0;
  wire h_u_cla32_and4509_y0;
  wire h_u_cla32_and4510_y0;
  wire h_u_cla32_and4511_y0;
  wire h_u_cla32_and4512_y0;
  wire h_u_cla32_and4513_y0;
  wire h_u_cla32_and4514_y0;
  wire h_u_cla32_and4515_y0;
  wire h_u_cla32_and4516_y0;
  wire h_u_cla32_and4517_y0;
  wire h_u_cla32_and4518_y0;
  wire h_u_cla32_and4519_y0;
  wire h_u_cla32_and4520_y0;
  wire h_u_cla32_and4521_y0;
  wire h_u_cla32_and4522_y0;
  wire h_u_cla32_and4523_y0;
  wire h_u_cla32_and4524_y0;
  wire h_u_cla32_and4525_y0;
  wire h_u_cla32_and4526_y0;
  wire h_u_cla32_and4527_y0;
  wire h_u_cla32_and4528_y0;
  wire h_u_cla32_and4529_y0;
  wire h_u_cla32_and4530_y0;
  wire h_u_cla32_and4531_y0;
  wire h_u_cla32_and4532_y0;
  wire h_u_cla32_and4533_y0;
  wire h_u_cla32_and4534_y0;
  wire h_u_cla32_and4535_y0;
  wire h_u_cla32_and4536_y0;
  wire h_u_cla32_and4537_y0;
  wire h_u_cla32_and4538_y0;
  wire h_u_cla32_and4539_y0;
  wire h_u_cla32_and4540_y0;
  wire h_u_cla32_and4541_y0;
  wire h_u_cla32_and4542_y0;
  wire h_u_cla32_and4543_y0;
  wire h_u_cla32_and4544_y0;
  wire h_u_cla32_and4545_y0;
  wire h_u_cla32_and4546_y0;
  wire h_u_cla32_and4547_y0;
  wire h_u_cla32_and4548_y0;
  wire h_u_cla32_and4549_y0;
  wire h_u_cla32_and4550_y0;
  wire h_u_cla32_and4551_y0;
  wire h_u_cla32_and4552_y0;
  wire h_u_cla32_and4553_y0;
  wire h_u_cla32_and4554_y0;
  wire h_u_cla32_and4555_y0;
  wire h_u_cla32_and4556_y0;
  wire h_u_cla32_and4557_y0;
  wire h_u_cla32_and4558_y0;
  wire h_u_cla32_and4559_y0;
  wire h_u_cla32_and4560_y0;
  wire h_u_cla32_and4561_y0;
  wire h_u_cla32_and4562_y0;
  wire h_u_cla32_and4563_y0;
  wire h_u_cla32_and4564_y0;
  wire h_u_cla32_and4565_y0;
  wire h_u_cla32_and4566_y0;
  wire h_u_cla32_and4567_y0;
  wire h_u_cla32_and4568_y0;
  wire h_u_cla32_and4569_y0;
  wire h_u_cla32_and4570_y0;
  wire h_u_cla32_and4571_y0;
  wire h_u_cla32_and4572_y0;
  wire h_u_cla32_and4573_y0;
  wire h_u_cla32_and4574_y0;
  wire h_u_cla32_and4575_y0;
  wire h_u_cla32_and4576_y0;
  wire h_u_cla32_and4577_y0;
  wire h_u_cla32_and4578_y0;
  wire h_u_cla32_and4579_y0;
  wire h_u_cla32_and4580_y0;
  wire h_u_cla32_and4581_y0;
  wire h_u_cla32_and4582_y0;
  wire h_u_cla32_and4583_y0;
  wire h_u_cla32_and4584_y0;
  wire h_u_cla32_and4585_y0;
  wire h_u_cla32_and4586_y0;
  wire h_u_cla32_and4587_y0;
  wire h_u_cla32_and4588_y0;
  wire h_u_cla32_and4589_y0;
  wire h_u_cla32_and4590_y0;
  wire h_u_cla32_and4591_y0;
  wire h_u_cla32_and4592_y0;
  wire h_u_cla32_and4593_y0;
  wire h_u_cla32_and4594_y0;
  wire h_u_cla32_and4595_y0;
  wire h_u_cla32_and4596_y0;
  wire h_u_cla32_and4597_y0;
  wire h_u_cla32_and4598_y0;
  wire h_u_cla32_and4599_y0;
  wire h_u_cla32_and4600_y0;
  wire h_u_cla32_and4601_y0;
  wire h_u_cla32_and4602_y0;
  wire h_u_cla32_and4603_y0;
  wire h_u_cla32_and4604_y0;
  wire h_u_cla32_and4605_y0;
  wire h_u_cla32_and4606_y0;
  wire h_u_cla32_and4607_y0;
  wire h_u_cla32_and4608_y0;
  wire h_u_cla32_and4609_y0;
  wire h_u_cla32_and4610_y0;
  wire h_u_cla32_and4611_y0;
  wire h_u_cla32_and4612_y0;
  wire h_u_cla32_and4613_y0;
  wire h_u_cla32_and4614_y0;
  wire h_u_cla32_and4615_y0;
  wire h_u_cla32_and4616_y0;
  wire h_u_cla32_and4617_y0;
  wire h_u_cla32_and4618_y0;
  wire h_u_cla32_and4619_y0;
  wire h_u_cla32_and4620_y0;
  wire h_u_cla32_and4621_y0;
  wire h_u_cla32_and4622_y0;
  wire h_u_cla32_and4623_y0;
  wire h_u_cla32_and4624_y0;
  wire h_u_cla32_and4625_y0;
  wire h_u_cla32_and4626_y0;
  wire h_u_cla32_and4627_y0;
  wire h_u_cla32_and4628_y0;
  wire h_u_cla32_and4629_y0;
  wire h_u_cla32_and4630_y0;
  wire h_u_cla32_and4631_y0;
  wire h_u_cla32_and4632_y0;
  wire h_u_cla32_and4633_y0;
  wire h_u_cla32_and4634_y0;
  wire h_u_cla32_and4635_y0;
  wire h_u_cla32_and4636_y0;
  wire h_u_cla32_and4637_y0;
  wire h_u_cla32_and4638_y0;
  wire h_u_cla32_and4639_y0;
  wire h_u_cla32_and4640_y0;
  wire h_u_cla32_and4641_y0;
  wire h_u_cla32_and4642_y0;
  wire h_u_cla32_and4643_y0;
  wire h_u_cla32_and4644_y0;
  wire h_u_cla32_and4645_y0;
  wire h_u_cla32_and4646_y0;
  wire h_u_cla32_and4647_y0;
  wire h_u_cla32_and4648_y0;
  wire h_u_cla32_and4649_y0;
  wire h_u_cla32_and4650_y0;
  wire h_u_cla32_and4651_y0;
  wire h_u_cla32_and4652_y0;
  wire h_u_cla32_and4653_y0;
  wire h_u_cla32_and4654_y0;
  wire h_u_cla32_and4655_y0;
  wire h_u_cla32_and4656_y0;
  wire h_u_cla32_and4657_y0;
  wire h_u_cla32_and4658_y0;
  wire h_u_cla32_and4659_y0;
  wire h_u_cla32_and4660_y0;
  wire h_u_cla32_and4661_y0;
  wire h_u_cla32_and4662_y0;
  wire h_u_cla32_and4663_y0;
  wire h_u_cla32_and4664_y0;
  wire h_u_cla32_and4665_y0;
  wire h_u_cla32_and4666_y0;
  wire h_u_cla32_and4667_y0;
  wire h_u_cla32_and4668_y0;
  wire h_u_cla32_and4669_y0;
  wire h_u_cla32_and4670_y0;
  wire h_u_cla32_and4671_y0;
  wire h_u_cla32_and4672_y0;
  wire h_u_cla32_and4673_y0;
  wire h_u_cla32_and4674_y0;
  wire h_u_cla32_and4675_y0;
  wire h_u_cla32_and4676_y0;
  wire h_u_cla32_and4677_y0;
  wire h_u_cla32_and4678_y0;
  wire h_u_cla32_and4679_y0;
  wire h_u_cla32_and4680_y0;
  wire h_u_cla32_and4681_y0;
  wire h_u_cla32_and4682_y0;
  wire h_u_cla32_and4683_y0;
  wire h_u_cla32_and4684_y0;
  wire h_u_cla32_and4685_y0;
  wire h_u_cla32_and4686_y0;
  wire h_u_cla32_and4687_y0;
  wire h_u_cla32_and4688_y0;
  wire h_u_cla32_and4689_y0;
  wire h_u_cla32_and4690_y0;
  wire h_u_cla32_and4691_y0;
  wire h_u_cla32_and4692_y0;
  wire h_u_cla32_and4693_y0;
  wire h_u_cla32_and4694_y0;
  wire h_u_cla32_and4695_y0;
  wire h_u_cla32_and4696_y0;
  wire h_u_cla32_and4697_y0;
  wire h_u_cla32_and4698_y0;
  wire h_u_cla32_and4699_y0;
  wire h_u_cla32_and4700_y0;
  wire h_u_cla32_and4701_y0;
  wire h_u_cla32_and4702_y0;
  wire h_u_cla32_and4703_y0;
  wire h_u_cla32_and4704_y0;
  wire h_u_cla32_and4705_y0;
  wire h_u_cla32_and4706_y0;
  wire h_u_cla32_and4707_y0;
  wire h_u_cla32_and4708_y0;
  wire h_u_cla32_and4709_y0;
  wire h_u_cla32_and4710_y0;
  wire h_u_cla32_and4711_y0;
  wire h_u_cla32_and4712_y0;
  wire h_u_cla32_and4713_y0;
  wire h_u_cla32_and4714_y0;
  wire h_u_cla32_and4715_y0;
  wire h_u_cla32_and4716_y0;
  wire h_u_cla32_and4717_y0;
  wire h_u_cla32_and4718_y0;
  wire h_u_cla32_and4719_y0;
  wire h_u_cla32_and4720_y0;
  wire h_u_cla32_and4721_y0;
  wire h_u_cla32_and4722_y0;
  wire h_u_cla32_and4723_y0;
  wire h_u_cla32_and4724_y0;
  wire h_u_cla32_and4725_y0;
  wire h_u_cla32_and4726_y0;
  wire h_u_cla32_and4727_y0;
  wire h_u_cla32_and4728_y0;
  wire h_u_cla32_and4729_y0;
  wire h_u_cla32_and4730_y0;
  wire h_u_cla32_and4731_y0;
  wire h_u_cla32_and4732_y0;
  wire h_u_cla32_and4733_y0;
  wire h_u_cla32_and4734_y0;
  wire h_u_cla32_and4735_y0;
  wire h_u_cla32_and4736_y0;
  wire h_u_cla32_and4737_y0;
  wire h_u_cla32_and4738_y0;
  wire h_u_cla32_and4739_y0;
  wire h_u_cla32_and4740_y0;
  wire h_u_cla32_and4741_y0;
  wire h_u_cla32_and4742_y0;
  wire h_u_cla32_and4743_y0;
  wire h_u_cla32_and4744_y0;
  wire h_u_cla32_and4745_y0;
  wire h_u_cla32_and4746_y0;
  wire h_u_cla32_and4747_y0;
  wire h_u_cla32_and4748_y0;
  wire h_u_cla32_and4749_y0;
  wire h_u_cla32_and4750_y0;
  wire h_u_cla32_and4751_y0;
  wire h_u_cla32_and4752_y0;
  wire h_u_cla32_and4753_y0;
  wire h_u_cla32_and4754_y0;
  wire h_u_cla32_and4755_y0;
  wire h_u_cla32_and4756_y0;
  wire h_u_cla32_and4757_y0;
  wire h_u_cla32_and4758_y0;
  wire h_u_cla32_and4759_y0;
  wire h_u_cla32_and4760_y0;
  wire h_u_cla32_and4761_y0;
  wire h_u_cla32_and4762_y0;
  wire h_u_cla32_and4763_y0;
  wire h_u_cla32_and4764_y0;
  wire h_u_cla32_and4765_y0;
  wire h_u_cla32_and4766_y0;
  wire h_u_cla32_and4767_y0;
  wire h_u_cla32_and4768_y0;
  wire h_u_cla32_and4769_y0;
  wire h_u_cla32_and4770_y0;
  wire h_u_cla32_and4771_y0;
  wire h_u_cla32_and4772_y0;
  wire h_u_cla32_and4773_y0;
  wire h_u_cla32_and4774_y0;
  wire h_u_cla32_and4775_y0;
  wire h_u_cla32_and4776_y0;
  wire h_u_cla32_and4777_y0;
  wire h_u_cla32_and4778_y0;
  wire h_u_cla32_and4779_y0;
  wire h_u_cla32_and4780_y0;
  wire h_u_cla32_and4781_y0;
  wire h_u_cla32_and4782_y0;
  wire h_u_cla32_and4783_y0;
  wire h_u_cla32_and4784_y0;
  wire h_u_cla32_and4785_y0;
  wire h_u_cla32_and4786_y0;
  wire h_u_cla32_and4787_y0;
  wire h_u_cla32_and4788_y0;
  wire h_u_cla32_and4789_y0;
  wire h_u_cla32_and4790_y0;
  wire h_u_cla32_and4791_y0;
  wire h_u_cla32_and4792_y0;
  wire h_u_cla32_and4793_y0;
  wire h_u_cla32_and4794_y0;
  wire h_u_cla32_and4795_y0;
  wire h_u_cla32_and4796_y0;
  wire h_u_cla32_and4797_y0;
  wire h_u_cla32_and4798_y0;
  wire h_u_cla32_and4799_y0;
  wire h_u_cla32_and4800_y0;
  wire h_u_cla32_and4801_y0;
  wire h_u_cla32_and4802_y0;
  wire h_u_cla32_and4803_y0;
  wire h_u_cla32_and4804_y0;
  wire h_u_cla32_and4805_y0;
  wire h_u_cla32_and4806_y0;
  wire h_u_cla32_and4807_y0;
  wire h_u_cla32_and4808_y0;
  wire h_u_cla32_and4809_y0;
  wire h_u_cla32_and4810_y0;
  wire h_u_cla32_and4811_y0;
  wire h_u_cla32_and4812_y0;
  wire h_u_cla32_and4813_y0;
  wire h_u_cla32_and4814_y0;
  wire h_u_cla32_and4815_y0;
  wire h_u_cla32_and4816_y0;
  wire h_u_cla32_and4817_y0;
  wire h_u_cla32_and4818_y0;
  wire h_u_cla32_and4819_y0;
  wire h_u_cla32_and4820_y0;
  wire h_u_cla32_and4821_y0;
  wire h_u_cla32_and4822_y0;
  wire h_u_cla32_and4823_y0;
  wire h_u_cla32_and4824_y0;
  wire h_u_cla32_and4825_y0;
  wire h_u_cla32_and4826_y0;
  wire h_u_cla32_and4827_y0;
  wire h_u_cla32_and4828_y0;
  wire h_u_cla32_and4829_y0;
  wire h_u_cla32_and4830_y0;
  wire h_u_cla32_and4831_y0;
  wire h_u_cla32_and4832_y0;
  wire h_u_cla32_and4833_y0;
  wire h_u_cla32_and4834_y0;
  wire h_u_cla32_and4835_y0;
  wire h_u_cla32_and4836_y0;
  wire h_u_cla32_and4837_y0;
  wire h_u_cla32_and4838_y0;
  wire h_u_cla32_and4839_y0;
  wire h_u_cla32_and4840_y0;
  wire h_u_cla32_and4841_y0;
  wire h_u_cla32_and4842_y0;
  wire h_u_cla32_and4843_y0;
  wire h_u_cla32_and4844_y0;
  wire h_u_cla32_and4845_y0;
  wire h_u_cla32_and4846_y0;
  wire h_u_cla32_and4847_y0;
  wire h_u_cla32_and4848_y0;
  wire h_u_cla32_and4849_y0;
  wire h_u_cla32_and4850_y0;
  wire h_u_cla32_and4851_y0;
  wire h_u_cla32_and4852_y0;
  wire h_u_cla32_and4853_y0;
  wire h_u_cla32_and4854_y0;
  wire h_u_cla32_and4855_y0;
  wire h_u_cla32_and4856_y0;
  wire h_u_cla32_and4857_y0;
  wire h_u_cla32_and4858_y0;
  wire h_u_cla32_and4859_y0;
  wire h_u_cla32_and4860_y0;
  wire h_u_cla32_and4861_y0;
  wire h_u_cla32_and4862_y0;
  wire h_u_cla32_and4863_y0;
  wire h_u_cla32_and4864_y0;
  wire h_u_cla32_and4865_y0;
  wire h_u_cla32_and4866_y0;
  wire h_u_cla32_and4867_y0;
  wire h_u_cla32_and4868_y0;
  wire h_u_cla32_and4869_y0;
  wire h_u_cla32_and4870_y0;
  wire h_u_cla32_and4871_y0;
  wire h_u_cla32_and4872_y0;
  wire h_u_cla32_and4873_y0;
  wire h_u_cla32_and4874_y0;
  wire h_u_cla32_and4875_y0;
  wire h_u_cla32_and4876_y0;
  wire h_u_cla32_and4877_y0;
  wire h_u_cla32_and4878_y0;
  wire h_u_cla32_and4879_y0;
  wire h_u_cla32_and4880_y0;
  wire h_u_cla32_and4881_y0;
  wire h_u_cla32_and4882_y0;
  wire h_u_cla32_and4883_y0;
  wire h_u_cla32_and4884_y0;
  wire h_u_cla32_and4885_y0;
  wire h_u_cla32_and4886_y0;
  wire h_u_cla32_and4887_y0;
  wire h_u_cla32_and4888_y0;
  wire h_u_cla32_and4889_y0;
  wire h_u_cla32_and4890_y0;
  wire h_u_cla32_and4891_y0;
  wire h_u_cla32_and4892_y0;
  wire h_u_cla32_and4893_y0;
  wire h_u_cla32_and4894_y0;
  wire h_u_cla32_and4895_y0;
  wire h_u_cla32_and4896_y0;
  wire h_u_cla32_and4897_y0;
  wire h_u_cla32_and4898_y0;
  wire h_u_cla32_and4899_y0;
  wire h_u_cla32_or276_y0;
  wire h_u_cla32_or277_y0;
  wire h_u_cla32_or278_y0;
  wire h_u_cla32_or279_y0;
  wire h_u_cla32_or280_y0;
  wire h_u_cla32_or281_y0;
  wire h_u_cla32_or282_y0;
  wire h_u_cla32_or283_y0;
  wire h_u_cla32_or284_y0;
  wire h_u_cla32_or285_y0;
  wire h_u_cla32_or286_y0;
  wire h_u_cla32_or287_y0;
  wire h_u_cla32_or288_y0;
  wire h_u_cla32_or289_y0;
  wire h_u_cla32_or290_y0;
  wire h_u_cla32_or291_y0;
  wire h_u_cla32_or292_y0;
  wire h_u_cla32_or293_y0;
  wire h_u_cla32_or294_y0;
  wire h_u_cla32_or295_y0;
  wire h_u_cla32_or296_y0;
  wire h_u_cla32_or297_y0;
  wire h_u_cla32_or298_y0;
  wire h_u_cla32_or299_y0;
  wire h_u_cla32_pg_logic24_y0;
  wire h_u_cla32_pg_logic24_y1;
  wire h_u_cla32_pg_logic24_y2;
  wire h_u_cla32_xor24_y0;
  wire h_u_cla32_and4900_y0;
  wire h_u_cla32_and4901_y0;
  wire h_u_cla32_and4902_y0;
  wire h_u_cla32_and4903_y0;
  wire h_u_cla32_and4904_y0;
  wire h_u_cla32_and4905_y0;
  wire h_u_cla32_and4906_y0;
  wire h_u_cla32_and4907_y0;
  wire h_u_cla32_and4908_y0;
  wire h_u_cla32_and4909_y0;
  wire h_u_cla32_and4910_y0;
  wire h_u_cla32_and4911_y0;
  wire h_u_cla32_and4912_y0;
  wire h_u_cla32_and4913_y0;
  wire h_u_cla32_and4914_y0;
  wire h_u_cla32_and4915_y0;
  wire h_u_cla32_and4916_y0;
  wire h_u_cla32_and4917_y0;
  wire h_u_cla32_and4918_y0;
  wire h_u_cla32_and4919_y0;
  wire h_u_cla32_and4920_y0;
  wire h_u_cla32_and4921_y0;
  wire h_u_cla32_and4922_y0;
  wire h_u_cla32_and4923_y0;
  wire h_u_cla32_and4924_y0;
  wire h_u_cla32_and4925_y0;
  wire h_u_cla32_and4926_y0;
  wire h_u_cla32_and4927_y0;
  wire h_u_cla32_and4928_y0;
  wire h_u_cla32_and4929_y0;
  wire h_u_cla32_and4930_y0;
  wire h_u_cla32_and4931_y0;
  wire h_u_cla32_and4932_y0;
  wire h_u_cla32_and4933_y0;
  wire h_u_cla32_and4934_y0;
  wire h_u_cla32_and4935_y0;
  wire h_u_cla32_and4936_y0;
  wire h_u_cla32_and4937_y0;
  wire h_u_cla32_and4938_y0;
  wire h_u_cla32_and4939_y0;
  wire h_u_cla32_and4940_y0;
  wire h_u_cla32_and4941_y0;
  wire h_u_cla32_and4942_y0;
  wire h_u_cla32_and4943_y0;
  wire h_u_cla32_and4944_y0;
  wire h_u_cla32_and4945_y0;
  wire h_u_cla32_and4946_y0;
  wire h_u_cla32_and4947_y0;
  wire h_u_cla32_and4948_y0;
  wire h_u_cla32_and4949_y0;
  wire h_u_cla32_and4950_y0;
  wire h_u_cla32_and4951_y0;
  wire h_u_cla32_and4952_y0;
  wire h_u_cla32_and4953_y0;
  wire h_u_cla32_and4954_y0;
  wire h_u_cla32_and4955_y0;
  wire h_u_cla32_and4956_y0;
  wire h_u_cla32_and4957_y0;
  wire h_u_cla32_and4958_y0;
  wire h_u_cla32_and4959_y0;
  wire h_u_cla32_and4960_y0;
  wire h_u_cla32_and4961_y0;
  wire h_u_cla32_and4962_y0;
  wire h_u_cla32_and4963_y0;
  wire h_u_cla32_and4964_y0;
  wire h_u_cla32_and4965_y0;
  wire h_u_cla32_and4966_y0;
  wire h_u_cla32_and4967_y0;
  wire h_u_cla32_and4968_y0;
  wire h_u_cla32_and4969_y0;
  wire h_u_cla32_and4970_y0;
  wire h_u_cla32_and4971_y0;
  wire h_u_cla32_and4972_y0;
  wire h_u_cla32_and4973_y0;
  wire h_u_cla32_and4974_y0;
  wire h_u_cla32_and4975_y0;
  wire h_u_cla32_and4976_y0;
  wire h_u_cla32_and4977_y0;
  wire h_u_cla32_and4978_y0;
  wire h_u_cla32_and4979_y0;
  wire h_u_cla32_and4980_y0;
  wire h_u_cla32_and4981_y0;
  wire h_u_cla32_and4982_y0;
  wire h_u_cla32_and4983_y0;
  wire h_u_cla32_and4984_y0;
  wire h_u_cla32_and4985_y0;
  wire h_u_cla32_and4986_y0;
  wire h_u_cla32_and4987_y0;
  wire h_u_cla32_and4988_y0;
  wire h_u_cla32_and4989_y0;
  wire h_u_cla32_and4990_y0;
  wire h_u_cla32_and4991_y0;
  wire h_u_cla32_and4992_y0;
  wire h_u_cla32_and4993_y0;
  wire h_u_cla32_and4994_y0;
  wire h_u_cla32_and4995_y0;
  wire h_u_cla32_and4996_y0;
  wire h_u_cla32_and4997_y0;
  wire h_u_cla32_and4998_y0;
  wire h_u_cla32_and4999_y0;
  wire h_u_cla32_and5000_y0;
  wire h_u_cla32_and5001_y0;
  wire h_u_cla32_and5002_y0;
  wire h_u_cla32_and5003_y0;
  wire h_u_cla32_and5004_y0;
  wire h_u_cla32_and5005_y0;
  wire h_u_cla32_and5006_y0;
  wire h_u_cla32_and5007_y0;
  wire h_u_cla32_and5008_y0;
  wire h_u_cla32_and5009_y0;
  wire h_u_cla32_and5010_y0;
  wire h_u_cla32_and5011_y0;
  wire h_u_cla32_and5012_y0;
  wire h_u_cla32_and5013_y0;
  wire h_u_cla32_and5014_y0;
  wire h_u_cla32_and5015_y0;
  wire h_u_cla32_and5016_y0;
  wire h_u_cla32_and5017_y0;
  wire h_u_cla32_and5018_y0;
  wire h_u_cla32_and5019_y0;
  wire h_u_cla32_and5020_y0;
  wire h_u_cla32_and5021_y0;
  wire h_u_cla32_and5022_y0;
  wire h_u_cla32_and5023_y0;
  wire h_u_cla32_and5024_y0;
  wire h_u_cla32_and5025_y0;
  wire h_u_cla32_and5026_y0;
  wire h_u_cla32_and5027_y0;
  wire h_u_cla32_and5028_y0;
  wire h_u_cla32_and5029_y0;
  wire h_u_cla32_and5030_y0;
  wire h_u_cla32_and5031_y0;
  wire h_u_cla32_and5032_y0;
  wire h_u_cla32_and5033_y0;
  wire h_u_cla32_and5034_y0;
  wire h_u_cla32_and5035_y0;
  wire h_u_cla32_and5036_y0;
  wire h_u_cla32_and5037_y0;
  wire h_u_cla32_and5038_y0;
  wire h_u_cla32_and5039_y0;
  wire h_u_cla32_and5040_y0;
  wire h_u_cla32_and5041_y0;
  wire h_u_cla32_and5042_y0;
  wire h_u_cla32_and5043_y0;
  wire h_u_cla32_and5044_y0;
  wire h_u_cla32_and5045_y0;
  wire h_u_cla32_and5046_y0;
  wire h_u_cla32_and5047_y0;
  wire h_u_cla32_and5048_y0;
  wire h_u_cla32_and5049_y0;
  wire h_u_cla32_and5050_y0;
  wire h_u_cla32_and5051_y0;
  wire h_u_cla32_and5052_y0;
  wire h_u_cla32_and5053_y0;
  wire h_u_cla32_and5054_y0;
  wire h_u_cla32_and5055_y0;
  wire h_u_cla32_and5056_y0;
  wire h_u_cla32_and5057_y0;
  wire h_u_cla32_and5058_y0;
  wire h_u_cla32_and5059_y0;
  wire h_u_cla32_and5060_y0;
  wire h_u_cla32_and5061_y0;
  wire h_u_cla32_and5062_y0;
  wire h_u_cla32_and5063_y0;
  wire h_u_cla32_and5064_y0;
  wire h_u_cla32_and5065_y0;
  wire h_u_cla32_and5066_y0;
  wire h_u_cla32_and5067_y0;
  wire h_u_cla32_and5068_y0;
  wire h_u_cla32_and5069_y0;
  wire h_u_cla32_and5070_y0;
  wire h_u_cla32_and5071_y0;
  wire h_u_cla32_and5072_y0;
  wire h_u_cla32_and5073_y0;
  wire h_u_cla32_and5074_y0;
  wire h_u_cla32_and5075_y0;
  wire h_u_cla32_and5076_y0;
  wire h_u_cla32_and5077_y0;
  wire h_u_cla32_and5078_y0;
  wire h_u_cla32_and5079_y0;
  wire h_u_cla32_and5080_y0;
  wire h_u_cla32_and5081_y0;
  wire h_u_cla32_and5082_y0;
  wire h_u_cla32_and5083_y0;
  wire h_u_cla32_and5084_y0;
  wire h_u_cla32_and5085_y0;
  wire h_u_cla32_and5086_y0;
  wire h_u_cla32_and5087_y0;
  wire h_u_cla32_and5088_y0;
  wire h_u_cla32_and5089_y0;
  wire h_u_cla32_and5090_y0;
  wire h_u_cla32_and5091_y0;
  wire h_u_cla32_and5092_y0;
  wire h_u_cla32_and5093_y0;
  wire h_u_cla32_and5094_y0;
  wire h_u_cla32_and5095_y0;
  wire h_u_cla32_and5096_y0;
  wire h_u_cla32_and5097_y0;
  wire h_u_cla32_and5098_y0;
  wire h_u_cla32_and5099_y0;
  wire h_u_cla32_and5100_y0;
  wire h_u_cla32_and5101_y0;
  wire h_u_cla32_and5102_y0;
  wire h_u_cla32_and5103_y0;
  wire h_u_cla32_and5104_y0;
  wire h_u_cla32_and5105_y0;
  wire h_u_cla32_and5106_y0;
  wire h_u_cla32_and5107_y0;
  wire h_u_cla32_and5108_y0;
  wire h_u_cla32_and5109_y0;
  wire h_u_cla32_and5110_y0;
  wire h_u_cla32_and5111_y0;
  wire h_u_cla32_and5112_y0;
  wire h_u_cla32_and5113_y0;
  wire h_u_cla32_and5114_y0;
  wire h_u_cla32_and5115_y0;
  wire h_u_cla32_and5116_y0;
  wire h_u_cla32_and5117_y0;
  wire h_u_cla32_and5118_y0;
  wire h_u_cla32_and5119_y0;
  wire h_u_cla32_and5120_y0;
  wire h_u_cla32_and5121_y0;
  wire h_u_cla32_and5122_y0;
  wire h_u_cla32_and5123_y0;
  wire h_u_cla32_and5124_y0;
  wire h_u_cla32_and5125_y0;
  wire h_u_cla32_and5126_y0;
  wire h_u_cla32_and5127_y0;
  wire h_u_cla32_and5128_y0;
  wire h_u_cla32_and5129_y0;
  wire h_u_cla32_and5130_y0;
  wire h_u_cla32_and5131_y0;
  wire h_u_cla32_and5132_y0;
  wire h_u_cla32_and5133_y0;
  wire h_u_cla32_and5134_y0;
  wire h_u_cla32_and5135_y0;
  wire h_u_cla32_and5136_y0;
  wire h_u_cla32_and5137_y0;
  wire h_u_cla32_and5138_y0;
  wire h_u_cla32_and5139_y0;
  wire h_u_cla32_and5140_y0;
  wire h_u_cla32_and5141_y0;
  wire h_u_cla32_and5142_y0;
  wire h_u_cla32_and5143_y0;
  wire h_u_cla32_and5144_y0;
  wire h_u_cla32_and5145_y0;
  wire h_u_cla32_and5146_y0;
  wire h_u_cla32_and5147_y0;
  wire h_u_cla32_and5148_y0;
  wire h_u_cla32_and5149_y0;
  wire h_u_cla32_and5150_y0;
  wire h_u_cla32_and5151_y0;
  wire h_u_cla32_and5152_y0;
  wire h_u_cla32_and5153_y0;
  wire h_u_cla32_and5154_y0;
  wire h_u_cla32_and5155_y0;
  wire h_u_cla32_and5156_y0;
  wire h_u_cla32_and5157_y0;
  wire h_u_cla32_and5158_y0;
  wire h_u_cla32_and5159_y0;
  wire h_u_cla32_and5160_y0;
  wire h_u_cla32_and5161_y0;
  wire h_u_cla32_and5162_y0;
  wire h_u_cla32_and5163_y0;
  wire h_u_cla32_and5164_y0;
  wire h_u_cla32_and5165_y0;
  wire h_u_cla32_and5166_y0;
  wire h_u_cla32_and5167_y0;
  wire h_u_cla32_and5168_y0;
  wire h_u_cla32_and5169_y0;
  wire h_u_cla32_and5170_y0;
  wire h_u_cla32_and5171_y0;
  wire h_u_cla32_and5172_y0;
  wire h_u_cla32_and5173_y0;
  wire h_u_cla32_and5174_y0;
  wire h_u_cla32_and5175_y0;
  wire h_u_cla32_and5176_y0;
  wire h_u_cla32_and5177_y0;
  wire h_u_cla32_and5178_y0;
  wire h_u_cla32_and5179_y0;
  wire h_u_cla32_and5180_y0;
  wire h_u_cla32_and5181_y0;
  wire h_u_cla32_and5182_y0;
  wire h_u_cla32_and5183_y0;
  wire h_u_cla32_and5184_y0;
  wire h_u_cla32_and5185_y0;
  wire h_u_cla32_and5186_y0;
  wire h_u_cla32_and5187_y0;
  wire h_u_cla32_and5188_y0;
  wire h_u_cla32_and5189_y0;
  wire h_u_cla32_and5190_y0;
  wire h_u_cla32_and5191_y0;
  wire h_u_cla32_and5192_y0;
  wire h_u_cla32_and5193_y0;
  wire h_u_cla32_and5194_y0;
  wire h_u_cla32_and5195_y0;
  wire h_u_cla32_and5196_y0;
  wire h_u_cla32_and5197_y0;
  wire h_u_cla32_and5198_y0;
  wire h_u_cla32_and5199_y0;
  wire h_u_cla32_and5200_y0;
  wire h_u_cla32_and5201_y0;
  wire h_u_cla32_and5202_y0;
  wire h_u_cla32_and5203_y0;
  wire h_u_cla32_and5204_y0;
  wire h_u_cla32_and5205_y0;
  wire h_u_cla32_and5206_y0;
  wire h_u_cla32_and5207_y0;
  wire h_u_cla32_and5208_y0;
  wire h_u_cla32_and5209_y0;
  wire h_u_cla32_and5210_y0;
  wire h_u_cla32_and5211_y0;
  wire h_u_cla32_and5212_y0;
  wire h_u_cla32_and5213_y0;
  wire h_u_cla32_and5214_y0;
  wire h_u_cla32_and5215_y0;
  wire h_u_cla32_and5216_y0;
  wire h_u_cla32_and5217_y0;
  wire h_u_cla32_and5218_y0;
  wire h_u_cla32_and5219_y0;
  wire h_u_cla32_and5220_y0;
  wire h_u_cla32_and5221_y0;
  wire h_u_cla32_and5222_y0;
  wire h_u_cla32_and5223_y0;
  wire h_u_cla32_and5224_y0;
  wire h_u_cla32_and5225_y0;
  wire h_u_cla32_and5226_y0;
  wire h_u_cla32_and5227_y0;
  wire h_u_cla32_and5228_y0;
  wire h_u_cla32_and5229_y0;
  wire h_u_cla32_and5230_y0;
  wire h_u_cla32_and5231_y0;
  wire h_u_cla32_and5232_y0;
  wire h_u_cla32_and5233_y0;
  wire h_u_cla32_and5234_y0;
  wire h_u_cla32_and5235_y0;
  wire h_u_cla32_and5236_y0;
  wire h_u_cla32_and5237_y0;
  wire h_u_cla32_and5238_y0;
  wire h_u_cla32_and5239_y0;
  wire h_u_cla32_and5240_y0;
  wire h_u_cla32_and5241_y0;
  wire h_u_cla32_and5242_y0;
  wire h_u_cla32_and5243_y0;
  wire h_u_cla32_and5244_y0;
  wire h_u_cla32_and5245_y0;
  wire h_u_cla32_and5246_y0;
  wire h_u_cla32_and5247_y0;
  wire h_u_cla32_and5248_y0;
  wire h_u_cla32_and5249_y0;
  wire h_u_cla32_and5250_y0;
  wire h_u_cla32_and5251_y0;
  wire h_u_cla32_and5252_y0;
  wire h_u_cla32_and5253_y0;
  wire h_u_cla32_and5254_y0;
  wire h_u_cla32_and5255_y0;
  wire h_u_cla32_and5256_y0;
  wire h_u_cla32_and5257_y0;
  wire h_u_cla32_and5258_y0;
  wire h_u_cla32_and5259_y0;
  wire h_u_cla32_and5260_y0;
  wire h_u_cla32_and5261_y0;
  wire h_u_cla32_and5262_y0;
  wire h_u_cla32_and5263_y0;
  wire h_u_cla32_and5264_y0;
  wire h_u_cla32_and5265_y0;
  wire h_u_cla32_and5266_y0;
  wire h_u_cla32_and5267_y0;
  wire h_u_cla32_and5268_y0;
  wire h_u_cla32_and5269_y0;
  wire h_u_cla32_and5270_y0;
  wire h_u_cla32_and5271_y0;
  wire h_u_cla32_and5272_y0;
  wire h_u_cla32_and5273_y0;
  wire h_u_cla32_and5274_y0;
  wire h_u_cla32_and5275_y0;
  wire h_u_cla32_and5276_y0;
  wire h_u_cla32_and5277_y0;
  wire h_u_cla32_and5278_y0;
  wire h_u_cla32_and5279_y0;
  wire h_u_cla32_and5280_y0;
  wire h_u_cla32_and5281_y0;
  wire h_u_cla32_and5282_y0;
  wire h_u_cla32_and5283_y0;
  wire h_u_cla32_and5284_y0;
  wire h_u_cla32_and5285_y0;
  wire h_u_cla32_and5286_y0;
  wire h_u_cla32_and5287_y0;
  wire h_u_cla32_and5288_y0;
  wire h_u_cla32_and5289_y0;
  wire h_u_cla32_and5290_y0;
  wire h_u_cla32_and5291_y0;
  wire h_u_cla32_and5292_y0;
  wire h_u_cla32_and5293_y0;
  wire h_u_cla32_and5294_y0;
  wire h_u_cla32_and5295_y0;
  wire h_u_cla32_and5296_y0;
  wire h_u_cla32_and5297_y0;
  wire h_u_cla32_and5298_y0;
  wire h_u_cla32_and5299_y0;
  wire h_u_cla32_and5300_y0;
  wire h_u_cla32_and5301_y0;
  wire h_u_cla32_and5302_y0;
  wire h_u_cla32_and5303_y0;
  wire h_u_cla32_and5304_y0;
  wire h_u_cla32_and5305_y0;
  wire h_u_cla32_and5306_y0;
  wire h_u_cla32_and5307_y0;
  wire h_u_cla32_and5308_y0;
  wire h_u_cla32_and5309_y0;
  wire h_u_cla32_and5310_y0;
  wire h_u_cla32_and5311_y0;
  wire h_u_cla32_and5312_y0;
  wire h_u_cla32_and5313_y0;
  wire h_u_cla32_and5314_y0;
  wire h_u_cla32_and5315_y0;
  wire h_u_cla32_and5316_y0;
  wire h_u_cla32_and5317_y0;
  wire h_u_cla32_and5318_y0;
  wire h_u_cla32_and5319_y0;
  wire h_u_cla32_and5320_y0;
  wire h_u_cla32_and5321_y0;
  wire h_u_cla32_and5322_y0;
  wire h_u_cla32_and5323_y0;
  wire h_u_cla32_and5324_y0;
  wire h_u_cla32_and5325_y0;
  wire h_u_cla32_and5326_y0;
  wire h_u_cla32_and5327_y0;
  wire h_u_cla32_and5328_y0;
  wire h_u_cla32_and5329_y0;
  wire h_u_cla32_and5330_y0;
  wire h_u_cla32_and5331_y0;
  wire h_u_cla32_and5332_y0;
  wire h_u_cla32_and5333_y0;
  wire h_u_cla32_and5334_y0;
  wire h_u_cla32_and5335_y0;
  wire h_u_cla32_and5336_y0;
  wire h_u_cla32_and5337_y0;
  wire h_u_cla32_and5338_y0;
  wire h_u_cla32_and5339_y0;
  wire h_u_cla32_and5340_y0;
  wire h_u_cla32_and5341_y0;
  wire h_u_cla32_and5342_y0;
  wire h_u_cla32_and5343_y0;
  wire h_u_cla32_and5344_y0;
  wire h_u_cla32_and5345_y0;
  wire h_u_cla32_and5346_y0;
  wire h_u_cla32_and5347_y0;
  wire h_u_cla32_and5348_y0;
  wire h_u_cla32_and5349_y0;
  wire h_u_cla32_and5350_y0;
  wire h_u_cla32_and5351_y0;
  wire h_u_cla32_and5352_y0;
  wire h_u_cla32_and5353_y0;
  wire h_u_cla32_and5354_y0;
  wire h_u_cla32_and5355_y0;
  wire h_u_cla32_and5356_y0;
  wire h_u_cla32_and5357_y0;
  wire h_u_cla32_and5358_y0;
  wire h_u_cla32_and5359_y0;
  wire h_u_cla32_and5360_y0;
  wire h_u_cla32_and5361_y0;
  wire h_u_cla32_and5362_y0;
  wire h_u_cla32_and5363_y0;
  wire h_u_cla32_and5364_y0;
  wire h_u_cla32_and5365_y0;
  wire h_u_cla32_and5366_y0;
  wire h_u_cla32_and5367_y0;
  wire h_u_cla32_and5368_y0;
  wire h_u_cla32_and5369_y0;
  wire h_u_cla32_and5370_y0;
  wire h_u_cla32_and5371_y0;
  wire h_u_cla32_and5372_y0;
  wire h_u_cla32_and5373_y0;
  wire h_u_cla32_and5374_y0;
  wire h_u_cla32_and5375_y0;
  wire h_u_cla32_and5376_y0;
  wire h_u_cla32_and5377_y0;
  wire h_u_cla32_and5378_y0;
  wire h_u_cla32_and5379_y0;
  wire h_u_cla32_and5380_y0;
  wire h_u_cla32_and5381_y0;
  wire h_u_cla32_and5382_y0;
  wire h_u_cla32_and5383_y0;
  wire h_u_cla32_and5384_y0;
  wire h_u_cla32_and5385_y0;
  wire h_u_cla32_and5386_y0;
  wire h_u_cla32_and5387_y0;
  wire h_u_cla32_and5388_y0;
  wire h_u_cla32_and5389_y0;
  wire h_u_cla32_and5390_y0;
  wire h_u_cla32_and5391_y0;
  wire h_u_cla32_and5392_y0;
  wire h_u_cla32_and5393_y0;
  wire h_u_cla32_and5394_y0;
  wire h_u_cla32_and5395_y0;
  wire h_u_cla32_and5396_y0;
  wire h_u_cla32_and5397_y0;
  wire h_u_cla32_and5398_y0;
  wire h_u_cla32_and5399_y0;
  wire h_u_cla32_and5400_y0;
  wire h_u_cla32_and5401_y0;
  wire h_u_cla32_and5402_y0;
  wire h_u_cla32_and5403_y0;
  wire h_u_cla32_and5404_y0;
  wire h_u_cla32_and5405_y0;
  wire h_u_cla32_and5406_y0;
  wire h_u_cla32_and5407_y0;
  wire h_u_cla32_and5408_y0;
  wire h_u_cla32_and5409_y0;
  wire h_u_cla32_and5410_y0;
  wire h_u_cla32_and5411_y0;
  wire h_u_cla32_and5412_y0;
  wire h_u_cla32_and5413_y0;
  wire h_u_cla32_and5414_y0;
  wire h_u_cla32_and5415_y0;
  wire h_u_cla32_and5416_y0;
  wire h_u_cla32_and5417_y0;
  wire h_u_cla32_and5418_y0;
  wire h_u_cla32_and5419_y0;
  wire h_u_cla32_and5420_y0;
  wire h_u_cla32_and5421_y0;
  wire h_u_cla32_and5422_y0;
  wire h_u_cla32_and5423_y0;
  wire h_u_cla32_and5424_y0;
  wire h_u_cla32_and5425_y0;
  wire h_u_cla32_and5426_y0;
  wire h_u_cla32_and5427_y0;
  wire h_u_cla32_and5428_y0;
  wire h_u_cla32_and5429_y0;
  wire h_u_cla32_and5430_y0;
  wire h_u_cla32_and5431_y0;
  wire h_u_cla32_and5432_y0;
  wire h_u_cla32_and5433_y0;
  wire h_u_cla32_and5434_y0;
  wire h_u_cla32_and5435_y0;
  wire h_u_cla32_and5436_y0;
  wire h_u_cla32_and5437_y0;
  wire h_u_cla32_and5438_y0;
  wire h_u_cla32_and5439_y0;
  wire h_u_cla32_and5440_y0;
  wire h_u_cla32_and5441_y0;
  wire h_u_cla32_and5442_y0;
  wire h_u_cla32_and5443_y0;
  wire h_u_cla32_and5444_y0;
  wire h_u_cla32_and5445_y0;
  wire h_u_cla32_and5446_y0;
  wire h_u_cla32_and5447_y0;
  wire h_u_cla32_and5448_y0;
  wire h_u_cla32_and5449_y0;
  wire h_u_cla32_and5450_y0;
  wire h_u_cla32_and5451_y0;
  wire h_u_cla32_and5452_y0;
  wire h_u_cla32_and5453_y0;
  wire h_u_cla32_and5454_y0;
  wire h_u_cla32_and5455_y0;
  wire h_u_cla32_and5456_y0;
  wire h_u_cla32_and5457_y0;
  wire h_u_cla32_and5458_y0;
  wire h_u_cla32_and5459_y0;
  wire h_u_cla32_and5460_y0;
  wire h_u_cla32_and5461_y0;
  wire h_u_cla32_and5462_y0;
  wire h_u_cla32_and5463_y0;
  wire h_u_cla32_and5464_y0;
  wire h_u_cla32_and5465_y0;
  wire h_u_cla32_and5466_y0;
  wire h_u_cla32_and5467_y0;
  wire h_u_cla32_and5468_y0;
  wire h_u_cla32_and5469_y0;
  wire h_u_cla32_and5470_y0;
  wire h_u_cla32_and5471_y0;
  wire h_u_cla32_and5472_y0;
  wire h_u_cla32_and5473_y0;
  wire h_u_cla32_and5474_y0;
  wire h_u_cla32_and5475_y0;
  wire h_u_cla32_and5476_y0;
  wire h_u_cla32_and5477_y0;
  wire h_u_cla32_and5478_y0;
  wire h_u_cla32_and5479_y0;
  wire h_u_cla32_and5480_y0;
  wire h_u_cla32_and5481_y0;
  wire h_u_cla32_and5482_y0;
  wire h_u_cla32_and5483_y0;
  wire h_u_cla32_and5484_y0;
  wire h_u_cla32_and5485_y0;
  wire h_u_cla32_and5486_y0;
  wire h_u_cla32_and5487_y0;
  wire h_u_cla32_and5488_y0;
  wire h_u_cla32_and5489_y0;
  wire h_u_cla32_and5490_y0;
  wire h_u_cla32_and5491_y0;
  wire h_u_cla32_and5492_y0;
  wire h_u_cla32_and5493_y0;
  wire h_u_cla32_and5494_y0;
  wire h_u_cla32_and5495_y0;
  wire h_u_cla32_and5496_y0;
  wire h_u_cla32_and5497_y0;
  wire h_u_cla32_and5498_y0;
  wire h_u_cla32_and5499_y0;
  wire h_u_cla32_and5500_y0;
  wire h_u_cla32_and5501_y0;
  wire h_u_cla32_and5502_y0;
  wire h_u_cla32_and5503_y0;
  wire h_u_cla32_and5504_y0;
  wire h_u_cla32_and5505_y0;
  wire h_u_cla32_and5506_y0;
  wire h_u_cla32_and5507_y0;
  wire h_u_cla32_and5508_y0;
  wire h_u_cla32_and5509_y0;
  wire h_u_cla32_and5510_y0;
  wire h_u_cla32_and5511_y0;
  wire h_u_cla32_and5512_y0;
  wire h_u_cla32_and5513_y0;
  wire h_u_cla32_and5514_y0;
  wire h_u_cla32_and5515_y0;
  wire h_u_cla32_and5516_y0;
  wire h_u_cla32_and5517_y0;
  wire h_u_cla32_and5518_y0;
  wire h_u_cla32_and5519_y0;
  wire h_u_cla32_and5520_y0;
  wire h_u_cla32_and5521_y0;
  wire h_u_cla32_and5522_y0;
  wire h_u_cla32_and5523_y0;
  wire h_u_cla32_and5524_y0;
  wire h_u_cla32_or300_y0;
  wire h_u_cla32_or301_y0;
  wire h_u_cla32_or302_y0;
  wire h_u_cla32_or303_y0;
  wire h_u_cla32_or304_y0;
  wire h_u_cla32_or305_y0;
  wire h_u_cla32_or306_y0;
  wire h_u_cla32_or307_y0;
  wire h_u_cla32_or308_y0;
  wire h_u_cla32_or309_y0;
  wire h_u_cla32_or310_y0;
  wire h_u_cla32_or311_y0;
  wire h_u_cla32_or312_y0;
  wire h_u_cla32_or313_y0;
  wire h_u_cla32_or314_y0;
  wire h_u_cla32_or315_y0;
  wire h_u_cla32_or316_y0;
  wire h_u_cla32_or317_y0;
  wire h_u_cla32_or318_y0;
  wire h_u_cla32_or319_y0;
  wire h_u_cla32_or320_y0;
  wire h_u_cla32_or321_y0;
  wire h_u_cla32_or322_y0;
  wire h_u_cla32_or323_y0;
  wire h_u_cla32_or324_y0;
  wire h_u_cla32_pg_logic25_y0;
  wire h_u_cla32_pg_logic25_y1;
  wire h_u_cla32_pg_logic25_y2;
  wire h_u_cla32_xor25_y0;
  wire h_u_cla32_and5525_y0;
  wire h_u_cla32_and5526_y0;
  wire h_u_cla32_and5527_y0;
  wire h_u_cla32_and5528_y0;
  wire h_u_cla32_and5529_y0;
  wire h_u_cla32_and5530_y0;
  wire h_u_cla32_and5531_y0;
  wire h_u_cla32_and5532_y0;
  wire h_u_cla32_and5533_y0;
  wire h_u_cla32_and5534_y0;
  wire h_u_cla32_and5535_y0;
  wire h_u_cla32_and5536_y0;
  wire h_u_cla32_and5537_y0;
  wire h_u_cla32_and5538_y0;
  wire h_u_cla32_and5539_y0;
  wire h_u_cla32_and5540_y0;
  wire h_u_cla32_and5541_y0;
  wire h_u_cla32_and5542_y0;
  wire h_u_cla32_and5543_y0;
  wire h_u_cla32_and5544_y0;
  wire h_u_cla32_and5545_y0;
  wire h_u_cla32_and5546_y0;
  wire h_u_cla32_and5547_y0;
  wire h_u_cla32_and5548_y0;
  wire h_u_cla32_and5549_y0;
  wire h_u_cla32_and5550_y0;
  wire h_u_cla32_and5551_y0;
  wire h_u_cla32_and5552_y0;
  wire h_u_cla32_and5553_y0;
  wire h_u_cla32_and5554_y0;
  wire h_u_cla32_and5555_y0;
  wire h_u_cla32_and5556_y0;
  wire h_u_cla32_and5557_y0;
  wire h_u_cla32_and5558_y0;
  wire h_u_cla32_and5559_y0;
  wire h_u_cla32_and5560_y0;
  wire h_u_cla32_and5561_y0;
  wire h_u_cla32_and5562_y0;
  wire h_u_cla32_and5563_y0;
  wire h_u_cla32_and5564_y0;
  wire h_u_cla32_and5565_y0;
  wire h_u_cla32_and5566_y0;
  wire h_u_cla32_and5567_y0;
  wire h_u_cla32_and5568_y0;
  wire h_u_cla32_and5569_y0;
  wire h_u_cla32_and5570_y0;
  wire h_u_cla32_and5571_y0;
  wire h_u_cla32_and5572_y0;
  wire h_u_cla32_and5573_y0;
  wire h_u_cla32_and5574_y0;
  wire h_u_cla32_and5575_y0;
  wire h_u_cla32_and5576_y0;
  wire h_u_cla32_and5577_y0;
  wire h_u_cla32_and5578_y0;
  wire h_u_cla32_and5579_y0;
  wire h_u_cla32_and5580_y0;
  wire h_u_cla32_and5581_y0;
  wire h_u_cla32_and5582_y0;
  wire h_u_cla32_and5583_y0;
  wire h_u_cla32_and5584_y0;
  wire h_u_cla32_and5585_y0;
  wire h_u_cla32_and5586_y0;
  wire h_u_cla32_and5587_y0;
  wire h_u_cla32_and5588_y0;
  wire h_u_cla32_and5589_y0;
  wire h_u_cla32_and5590_y0;
  wire h_u_cla32_and5591_y0;
  wire h_u_cla32_and5592_y0;
  wire h_u_cla32_and5593_y0;
  wire h_u_cla32_and5594_y0;
  wire h_u_cla32_and5595_y0;
  wire h_u_cla32_and5596_y0;
  wire h_u_cla32_and5597_y0;
  wire h_u_cla32_and5598_y0;
  wire h_u_cla32_and5599_y0;
  wire h_u_cla32_and5600_y0;
  wire h_u_cla32_and5601_y0;
  wire h_u_cla32_and5602_y0;
  wire h_u_cla32_and5603_y0;
  wire h_u_cla32_and5604_y0;
  wire h_u_cla32_and5605_y0;
  wire h_u_cla32_and5606_y0;
  wire h_u_cla32_and5607_y0;
  wire h_u_cla32_and5608_y0;
  wire h_u_cla32_and5609_y0;
  wire h_u_cla32_and5610_y0;
  wire h_u_cla32_and5611_y0;
  wire h_u_cla32_and5612_y0;
  wire h_u_cla32_and5613_y0;
  wire h_u_cla32_and5614_y0;
  wire h_u_cla32_and5615_y0;
  wire h_u_cla32_and5616_y0;
  wire h_u_cla32_and5617_y0;
  wire h_u_cla32_and5618_y0;
  wire h_u_cla32_and5619_y0;
  wire h_u_cla32_and5620_y0;
  wire h_u_cla32_and5621_y0;
  wire h_u_cla32_and5622_y0;
  wire h_u_cla32_and5623_y0;
  wire h_u_cla32_and5624_y0;
  wire h_u_cla32_and5625_y0;
  wire h_u_cla32_and5626_y0;
  wire h_u_cla32_and5627_y0;
  wire h_u_cla32_and5628_y0;
  wire h_u_cla32_and5629_y0;
  wire h_u_cla32_and5630_y0;
  wire h_u_cla32_and5631_y0;
  wire h_u_cla32_and5632_y0;
  wire h_u_cla32_and5633_y0;
  wire h_u_cla32_and5634_y0;
  wire h_u_cla32_and5635_y0;
  wire h_u_cla32_and5636_y0;
  wire h_u_cla32_and5637_y0;
  wire h_u_cla32_and5638_y0;
  wire h_u_cla32_and5639_y0;
  wire h_u_cla32_and5640_y0;
  wire h_u_cla32_and5641_y0;
  wire h_u_cla32_and5642_y0;
  wire h_u_cla32_and5643_y0;
  wire h_u_cla32_and5644_y0;
  wire h_u_cla32_and5645_y0;
  wire h_u_cla32_and5646_y0;
  wire h_u_cla32_and5647_y0;
  wire h_u_cla32_and5648_y0;
  wire h_u_cla32_and5649_y0;
  wire h_u_cla32_and5650_y0;
  wire h_u_cla32_and5651_y0;
  wire h_u_cla32_and5652_y0;
  wire h_u_cla32_and5653_y0;
  wire h_u_cla32_and5654_y0;
  wire h_u_cla32_and5655_y0;
  wire h_u_cla32_and5656_y0;
  wire h_u_cla32_and5657_y0;
  wire h_u_cla32_and5658_y0;
  wire h_u_cla32_and5659_y0;
  wire h_u_cla32_and5660_y0;
  wire h_u_cla32_and5661_y0;
  wire h_u_cla32_and5662_y0;
  wire h_u_cla32_and5663_y0;
  wire h_u_cla32_and5664_y0;
  wire h_u_cla32_and5665_y0;
  wire h_u_cla32_and5666_y0;
  wire h_u_cla32_and5667_y0;
  wire h_u_cla32_and5668_y0;
  wire h_u_cla32_and5669_y0;
  wire h_u_cla32_and5670_y0;
  wire h_u_cla32_and5671_y0;
  wire h_u_cla32_and5672_y0;
  wire h_u_cla32_and5673_y0;
  wire h_u_cla32_and5674_y0;
  wire h_u_cla32_and5675_y0;
  wire h_u_cla32_and5676_y0;
  wire h_u_cla32_and5677_y0;
  wire h_u_cla32_and5678_y0;
  wire h_u_cla32_and5679_y0;
  wire h_u_cla32_and5680_y0;
  wire h_u_cla32_and5681_y0;
  wire h_u_cla32_and5682_y0;
  wire h_u_cla32_and5683_y0;
  wire h_u_cla32_and5684_y0;
  wire h_u_cla32_and5685_y0;
  wire h_u_cla32_and5686_y0;
  wire h_u_cla32_and5687_y0;
  wire h_u_cla32_and5688_y0;
  wire h_u_cla32_and5689_y0;
  wire h_u_cla32_and5690_y0;
  wire h_u_cla32_and5691_y0;
  wire h_u_cla32_and5692_y0;
  wire h_u_cla32_and5693_y0;
  wire h_u_cla32_and5694_y0;
  wire h_u_cla32_and5695_y0;
  wire h_u_cla32_and5696_y0;
  wire h_u_cla32_and5697_y0;
  wire h_u_cla32_and5698_y0;
  wire h_u_cla32_and5699_y0;
  wire h_u_cla32_and5700_y0;
  wire h_u_cla32_and5701_y0;
  wire h_u_cla32_and5702_y0;
  wire h_u_cla32_and5703_y0;
  wire h_u_cla32_and5704_y0;
  wire h_u_cla32_and5705_y0;
  wire h_u_cla32_and5706_y0;
  wire h_u_cla32_and5707_y0;
  wire h_u_cla32_and5708_y0;
  wire h_u_cla32_and5709_y0;
  wire h_u_cla32_and5710_y0;
  wire h_u_cla32_and5711_y0;
  wire h_u_cla32_and5712_y0;
  wire h_u_cla32_and5713_y0;
  wire h_u_cla32_and5714_y0;
  wire h_u_cla32_and5715_y0;
  wire h_u_cla32_and5716_y0;
  wire h_u_cla32_and5717_y0;
  wire h_u_cla32_and5718_y0;
  wire h_u_cla32_and5719_y0;
  wire h_u_cla32_and5720_y0;
  wire h_u_cla32_and5721_y0;
  wire h_u_cla32_and5722_y0;
  wire h_u_cla32_and5723_y0;
  wire h_u_cla32_and5724_y0;
  wire h_u_cla32_and5725_y0;
  wire h_u_cla32_and5726_y0;
  wire h_u_cla32_and5727_y0;
  wire h_u_cla32_and5728_y0;
  wire h_u_cla32_and5729_y0;
  wire h_u_cla32_and5730_y0;
  wire h_u_cla32_and5731_y0;
  wire h_u_cla32_and5732_y0;
  wire h_u_cla32_and5733_y0;
  wire h_u_cla32_and5734_y0;
  wire h_u_cla32_and5735_y0;
  wire h_u_cla32_and5736_y0;
  wire h_u_cla32_and5737_y0;
  wire h_u_cla32_and5738_y0;
  wire h_u_cla32_and5739_y0;
  wire h_u_cla32_and5740_y0;
  wire h_u_cla32_and5741_y0;
  wire h_u_cla32_and5742_y0;
  wire h_u_cla32_and5743_y0;
  wire h_u_cla32_and5744_y0;
  wire h_u_cla32_and5745_y0;
  wire h_u_cla32_and5746_y0;
  wire h_u_cla32_and5747_y0;
  wire h_u_cla32_and5748_y0;
  wire h_u_cla32_and5749_y0;
  wire h_u_cla32_and5750_y0;
  wire h_u_cla32_and5751_y0;
  wire h_u_cla32_and5752_y0;
  wire h_u_cla32_and5753_y0;
  wire h_u_cla32_and5754_y0;
  wire h_u_cla32_and5755_y0;
  wire h_u_cla32_and5756_y0;
  wire h_u_cla32_and5757_y0;
  wire h_u_cla32_and5758_y0;
  wire h_u_cla32_and5759_y0;
  wire h_u_cla32_and5760_y0;
  wire h_u_cla32_and5761_y0;
  wire h_u_cla32_and5762_y0;
  wire h_u_cla32_and5763_y0;
  wire h_u_cla32_and5764_y0;
  wire h_u_cla32_and5765_y0;
  wire h_u_cla32_and5766_y0;
  wire h_u_cla32_and5767_y0;
  wire h_u_cla32_and5768_y0;
  wire h_u_cla32_and5769_y0;
  wire h_u_cla32_and5770_y0;
  wire h_u_cla32_and5771_y0;
  wire h_u_cla32_and5772_y0;
  wire h_u_cla32_and5773_y0;
  wire h_u_cla32_and5774_y0;
  wire h_u_cla32_and5775_y0;
  wire h_u_cla32_and5776_y0;
  wire h_u_cla32_and5777_y0;
  wire h_u_cla32_and5778_y0;
  wire h_u_cla32_and5779_y0;
  wire h_u_cla32_and5780_y0;
  wire h_u_cla32_and5781_y0;
  wire h_u_cla32_and5782_y0;
  wire h_u_cla32_and5783_y0;
  wire h_u_cla32_and5784_y0;
  wire h_u_cla32_and5785_y0;
  wire h_u_cla32_and5786_y0;
  wire h_u_cla32_and5787_y0;
  wire h_u_cla32_and5788_y0;
  wire h_u_cla32_and5789_y0;
  wire h_u_cla32_and5790_y0;
  wire h_u_cla32_and5791_y0;
  wire h_u_cla32_and5792_y0;
  wire h_u_cla32_and5793_y0;
  wire h_u_cla32_and5794_y0;
  wire h_u_cla32_and5795_y0;
  wire h_u_cla32_and5796_y0;
  wire h_u_cla32_and5797_y0;
  wire h_u_cla32_and5798_y0;
  wire h_u_cla32_and5799_y0;
  wire h_u_cla32_and5800_y0;
  wire h_u_cla32_and5801_y0;
  wire h_u_cla32_and5802_y0;
  wire h_u_cla32_and5803_y0;
  wire h_u_cla32_and5804_y0;
  wire h_u_cla32_and5805_y0;
  wire h_u_cla32_and5806_y0;
  wire h_u_cla32_and5807_y0;
  wire h_u_cla32_and5808_y0;
  wire h_u_cla32_and5809_y0;
  wire h_u_cla32_and5810_y0;
  wire h_u_cla32_and5811_y0;
  wire h_u_cla32_and5812_y0;
  wire h_u_cla32_and5813_y0;
  wire h_u_cla32_and5814_y0;
  wire h_u_cla32_and5815_y0;
  wire h_u_cla32_and5816_y0;
  wire h_u_cla32_and5817_y0;
  wire h_u_cla32_and5818_y0;
  wire h_u_cla32_and5819_y0;
  wire h_u_cla32_and5820_y0;
  wire h_u_cla32_and5821_y0;
  wire h_u_cla32_and5822_y0;
  wire h_u_cla32_and5823_y0;
  wire h_u_cla32_and5824_y0;
  wire h_u_cla32_and5825_y0;
  wire h_u_cla32_and5826_y0;
  wire h_u_cla32_and5827_y0;
  wire h_u_cla32_and5828_y0;
  wire h_u_cla32_and5829_y0;
  wire h_u_cla32_and5830_y0;
  wire h_u_cla32_and5831_y0;
  wire h_u_cla32_and5832_y0;
  wire h_u_cla32_and5833_y0;
  wire h_u_cla32_and5834_y0;
  wire h_u_cla32_and5835_y0;
  wire h_u_cla32_and5836_y0;
  wire h_u_cla32_and5837_y0;
  wire h_u_cla32_and5838_y0;
  wire h_u_cla32_and5839_y0;
  wire h_u_cla32_and5840_y0;
  wire h_u_cla32_and5841_y0;
  wire h_u_cla32_and5842_y0;
  wire h_u_cla32_and5843_y0;
  wire h_u_cla32_and5844_y0;
  wire h_u_cla32_and5845_y0;
  wire h_u_cla32_and5846_y0;
  wire h_u_cla32_and5847_y0;
  wire h_u_cla32_and5848_y0;
  wire h_u_cla32_and5849_y0;
  wire h_u_cla32_and5850_y0;
  wire h_u_cla32_and5851_y0;
  wire h_u_cla32_and5852_y0;
  wire h_u_cla32_and5853_y0;
  wire h_u_cla32_and5854_y0;
  wire h_u_cla32_and5855_y0;
  wire h_u_cla32_and5856_y0;
  wire h_u_cla32_and5857_y0;
  wire h_u_cla32_and5858_y0;
  wire h_u_cla32_and5859_y0;
  wire h_u_cla32_and5860_y0;
  wire h_u_cla32_and5861_y0;
  wire h_u_cla32_and5862_y0;
  wire h_u_cla32_and5863_y0;
  wire h_u_cla32_and5864_y0;
  wire h_u_cla32_and5865_y0;
  wire h_u_cla32_and5866_y0;
  wire h_u_cla32_and5867_y0;
  wire h_u_cla32_and5868_y0;
  wire h_u_cla32_and5869_y0;
  wire h_u_cla32_and5870_y0;
  wire h_u_cla32_and5871_y0;
  wire h_u_cla32_and5872_y0;
  wire h_u_cla32_and5873_y0;
  wire h_u_cla32_and5874_y0;
  wire h_u_cla32_and5875_y0;
  wire h_u_cla32_and5876_y0;
  wire h_u_cla32_and5877_y0;
  wire h_u_cla32_and5878_y0;
  wire h_u_cla32_and5879_y0;
  wire h_u_cla32_and5880_y0;
  wire h_u_cla32_and5881_y0;
  wire h_u_cla32_and5882_y0;
  wire h_u_cla32_and5883_y0;
  wire h_u_cla32_and5884_y0;
  wire h_u_cla32_and5885_y0;
  wire h_u_cla32_and5886_y0;
  wire h_u_cla32_and5887_y0;
  wire h_u_cla32_and5888_y0;
  wire h_u_cla32_and5889_y0;
  wire h_u_cla32_and5890_y0;
  wire h_u_cla32_and5891_y0;
  wire h_u_cla32_and5892_y0;
  wire h_u_cla32_and5893_y0;
  wire h_u_cla32_and5894_y0;
  wire h_u_cla32_and5895_y0;
  wire h_u_cla32_and5896_y0;
  wire h_u_cla32_and5897_y0;
  wire h_u_cla32_and5898_y0;
  wire h_u_cla32_and5899_y0;
  wire h_u_cla32_and5900_y0;
  wire h_u_cla32_and5901_y0;
  wire h_u_cla32_and5902_y0;
  wire h_u_cla32_and5903_y0;
  wire h_u_cla32_and5904_y0;
  wire h_u_cla32_and5905_y0;
  wire h_u_cla32_and5906_y0;
  wire h_u_cla32_and5907_y0;
  wire h_u_cla32_and5908_y0;
  wire h_u_cla32_and5909_y0;
  wire h_u_cla32_and5910_y0;
  wire h_u_cla32_and5911_y0;
  wire h_u_cla32_and5912_y0;
  wire h_u_cla32_and5913_y0;
  wire h_u_cla32_and5914_y0;
  wire h_u_cla32_and5915_y0;
  wire h_u_cla32_and5916_y0;
  wire h_u_cla32_and5917_y0;
  wire h_u_cla32_and5918_y0;
  wire h_u_cla32_and5919_y0;
  wire h_u_cla32_and5920_y0;
  wire h_u_cla32_and5921_y0;
  wire h_u_cla32_and5922_y0;
  wire h_u_cla32_and5923_y0;
  wire h_u_cla32_and5924_y0;
  wire h_u_cla32_and5925_y0;
  wire h_u_cla32_and5926_y0;
  wire h_u_cla32_and5927_y0;
  wire h_u_cla32_and5928_y0;
  wire h_u_cla32_and5929_y0;
  wire h_u_cla32_and5930_y0;
  wire h_u_cla32_and5931_y0;
  wire h_u_cla32_and5932_y0;
  wire h_u_cla32_and5933_y0;
  wire h_u_cla32_and5934_y0;
  wire h_u_cla32_and5935_y0;
  wire h_u_cla32_and5936_y0;
  wire h_u_cla32_and5937_y0;
  wire h_u_cla32_and5938_y0;
  wire h_u_cla32_and5939_y0;
  wire h_u_cla32_and5940_y0;
  wire h_u_cla32_and5941_y0;
  wire h_u_cla32_and5942_y0;
  wire h_u_cla32_and5943_y0;
  wire h_u_cla32_and5944_y0;
  wire h_u_cla32_and5945_y0;
  wire h_u_cla32_and5946_y0;
  wire h_u_cla32_and5947_y0;
  wire h_u_cla32_and5948_y0;
  wire h_u_cla32_and5949_y0;
  wire h_u_cla32_and5950_y0;
  wire h_u_cla32_and5951_y0;
  wire h_u_cla32_and5952_y0;
  wire h_u_cla32_and5953_y0;
  wire h_u_cla32_and5954_y0;
  wire h_u_cla32_and5955_y0;
  wire h_u_cla32_and5956_y0;
  wire h_u_cla32_and5957_y0;
  wire h_u_cla32_and5958_y0;
  wire h_u_cla32_and5959_y0;
  wire h_u_cla32_and5960_y0;
  wire h_u_cla32_and5961_y0;
  wire h_u_cla32_and5962_y0;
  wire h_u_cla32_and5963_y0;
  wire h_u_cla32_and5964_y0;
  wire h_u_cla32_and5965_y0;
  wire h_u_cla32_and5966_y0;
  wire h_u_cla32_and5967_y0;
  wire h_u_cla32_and5968_y0;
  wire h_u_cla32_and5969_y0;
  wire h_u_cla32_and5970_y0;
  wire h_u_cla32_and5971_y0;
  wire h_u_cla32_and5972_y0;
  wire h_u_cla32_and5973_y0;
  wire h_u_cla32_and5974_y0;
  wire h_u_cla32_and5975_y0;
  wire h_u_cla32_and5976_y0;
  wire h_u_cla32_and5977_y0;
  wire h_u_cla32_and5978_y0;
  wire h_u_cla32_and5979_y0;
  wire h_u_cla32_and5980_y0;
  wire h_u_cla32_and5981_y0;
  wire h_u_cla32_and5982_y0;
  wire h_u_cla32_and5983_y0;
  wire h_u_cla32_and5984_y0;
  wire h_u_cla32_and5985_y0;
  wire h_u_cla32_and5986_y0;
  wire h_u_cla32_and5987_y0;
  wire h_u_cla32_and5988_y0;
  wire h_u_cla32_and5989_y0;
  wire h_u_cla32_and5990_y0;
  wire h_u_cla32_and5991_y0;
  wire h_u_cla32_and5992_y0;
  wire h_u_cla32_and5993_y0;
  wire h_u_cla32_and5994_y0;
  wire h_u_cla32_and5995_y0;
  wire h_u_cla32_and5996_y0;
  wire h_u_cla32_and5997_y0;
  wire h_u_cla32_and5998_y0;
  wire h_u_cla32_and5999_y0;
  wire h_u_cla32_and6000_y0;
  wire h_u_cla32_and6001_y0;
  wire h_u_cla32_and6002_y0;
  wire h_u_cla32_and6003_y0;
  wire h_u_cla32_and6004_y0;
  wire h_u_cla32_and6005_y0;
  wire h_u_cla32_and6006_y0;
  wire h_u_cla32_and6007_y0;
  wire h_u_cla32_and6008_y0;
  wire h_u_cla32_and6009_y0;
  wire h_u_cla32_and6010_y0;
  wire h_u_cla32_and6011_y0;
  wire h_u_cla32_and6012_y0;
  wire h_u_cla32_and6013_y0;
  wire h_u_cla32_and6014_y0;
  wire h_u_cla32_and6015_y0;
  wire h_u_cla32_and6016_y0;
  wire h_u_cla32_and6017_y0;
  wire h_u_cla32_and6018_y0;
  wire h_u_cla32_and6019_y0;
  wire h_u_cla32_and6020_y0;
  wire h_u_cla32_and6021_y0;
  wire h_u_cla32_and6022_y0;
  wire h_u_cla32_and6023_y0;
  wire h_u_cla32_and6024_y0;
  wire h_u_cla32_and6025_y0;
  wire h_u_cla32_and6026_y0;
  wire h_u_cla32_and6027_y0;
  wire h_u_cla32_and6028_y0;
  wire h_u_cla32_and6029_y0;
  wire h_u_cla32_and6030_y0;
  wire h_u_cla32_and6031_y0;
  wire h_u_cla32_and6032_y0;
  wire h_u_cla32_and6033_y0;
  wire h_u_cla32_and6034_y0;
  wire h_u_cla32_and6035_y0;
  wire h_u_cla32_and6036_y0;
  wire h_u_cla32_and6037_y0;
  wire h_u_cla32_and6038_y0;
  wire h_u_cla32_and6039_y0;
  wire h_u_cla32_and6040_y0;
  wire h_u_cla32_and6041_y0;
  wire h_u_cla32_and6042_y0;
  wire h_u_cla32_and6043_y0;
  wire h_u_cla32_and6044_y0;
  wire h_u_cla32_and6045_y0;
  wire h_u_cla32_and6046_y0;
  wire h_u_cla32_and6047_y0;
  wire h_u_cla32_and6048_y0;
  wire h_u_cla32_and6049_y0;
  wire h_u_cla32_and6050_y0;
  wire h_u_cla32_and6051_y0;
  wire h_u_cla32_and6052_y0;
  wire h_u_cla32_and6053_y0;
  wire h_u_cla32_and6054_y0;
  wire h_u_cla32_and6055_y0;
  wire h_u_cla32_and6056_y0;
  wire h_u_cla32_and6057_y0;
  wire h_u_cla32_and6058_y0;
  wire h_u_cla32_and6059_y0;
  wire h_u_cla32_and6060_y0;
  wire h_u_cla32_and6061_y0;
  wire h_u_cla32_and6062_y0;
  wire h_u_cla32_and6063_y0;
  wire h_u_cla32_and6064_y0;
  wire h_u_cla32_and6065_y0;
  wire h_u_cla32_and6066_y0;
  wire h_u_cla32_and6067_y0;
  wire h_u_cla32_and6068_y0;
  wire h_u_cla32_and6069_y0;
  wire h_u_cla32_and6070_y0;
  wire h_u_cla32_and6071_y0;
  wire h_u_cla32_and6072_y0;
  wire h_u_cla32_and6073_y0;
  wire h_u_cla32_and6074_y0;
  wire h_u_cla32_and6075_y0;
  wire h_u_cla32_and6076_y0;
  wire h_u_cla32_and6077_y0;
  wire h_u_cla32_and6078_y0;
  wire h_u_cla32_and6079_y0;
  wire h_u_cla32_and6080_y0;
  wire h_u_cla32_and6081_y0;
  wire h_u_cla32_and6082_y0;
  wire h_u_cla32_and6083_y0;
  wire h_u_cla32_and6084_y0;
  wire h_u_cla32_and6085_y0;
  wire h_u_cla32_and6086_y0;
  wire h_u_cla32_and6087_y0;
  wire h_u_cla32_and6088_y0;
  wire h_u_cla32_and6089_y0;
  wire h_u_cla32_and6090_y0;
  wire h_u_cla32_and6091_y0;
  wire h_u_cla32_and6092_y0;
  wire h_u_cla32_and6093_y0;
  wire h_u_cla32_and6094_y0;
  wire h_u_cla32_and6095_y0;
  wire h_u_cla32_and6096_y0;
  wire h_u_cla32_and6097_y0;
  wire h_u_cla32_and6098_y0;
  wire h_u_cla32_and6099_y0;
  wire h_u_cla32_and6100_y0;
  wire h_u_cla32_and6101_y0;
  wire h_u_cla32_and6102_y0;
  wire h_u_cla32_and6103_y0;
  wire h_u_cla32_and6104_y0;
  wire h_u_cla32_and6105_y0;
  wire h_u_cla32_and6106_y0;
  wire h_u_cla32_and6107_y0;
  wire h_u_cla32_and6108_y0;
  wire h_u_cla32_and6109_y0;
  wire h_u_cla32_and6110_y0;
  wire h_u_cla32_and6111_y0;
  wire h_u_cla32_and6112_y0;
  wire h_u_cla32_and6113_y0;
  wire h_u_cla32_and6114_y0;
  wire h_u_cla32_and6115_y0;
  wire h_u_cla32_and6116_y0;
  wire h_u_cla32_and6117_y0;
  wire h_u_cla32_and6118_y0;
  wire h_u_cla32_and6119_y0;
  wire h_u_cla32_and6120_y0;
  wire h_u_cla32_and6121_y0;
  wire h_u_cla32_and6122_y0;
  wire h_u_cla32_and6123_y0;
  wire h_u_cla32_and6124_y0;
  wire h_u_cla32_and6125_y0;
  wire h_u_cla32_and6126_y0;
  wire h_u_cla32_and6127_y0;
  wire h_u_cla32_and6128_y0;
  wire h_u_cla32_and6129_y0;
  wire h_u_cla32_and6130_y0;
  wire h_u_cla32_and6131_y0;
  wire h_u_cla32_and6132_y0;
  wire h_u_cla32_and6133_y0;
  wire h_u_cla32_and6134_y0;
  wire h_u_cla32_and6135_y0;
  wire h_u_cla32_and6136_y0;
  wire h_u_cla32_and6137_y0;
  wire h_u_cla32_and6138_y0;
  wire h_u_cla32_and6139_y0;
  wire h_u_cla32_and6140_y0;
  wire h_u_cla32_and6141_y0;
  wire h_u_cla32_and6142_y0;
  wire h_u_cla32_and6143_y0;
  wire h_u_cla32_and6144_y0;
  wire h_u_cla32_and6145_y0;
  wire h_u_cla32_and6146_y0;
  wire h_u_cla32_and6147_y0;
  wire h_u_cla32_and6148_y0;
  wire h_u_cla32_and6149_y0;
  wire h_u_cla32_and6150_y0;
  wire h_u_cla32_and6151_y0;
  wire h_u_cla32_and6152_y0;
  wire h_u_cla32_and6153_y0;
  wire h_u_cla32_and6154_y0;
  wire h_u_cla32_and6155_y0;
  wire h_u_cla32_and6156_y0;
  wire h_u_cla32_and6157_y0;
  wire h_u_cla32_and6158_y0;
  wire h_u_cla32_and6159_y0;
  wire h_u_cla32_and6160_y0;
  wire h_u_cla32_and6161_y0;
  wire h_u_cla32_and6162_y0;
  wire h_u_cla32_and6163_y0;
  wire h_u_cla32_and6164_y0;
  wire h_u_cla32_and6165_y0;
  wire h_u_cla32_and6166_y0;
  wire h_u_cla32_and6167_y0;
  wire h_u_cla32_and6168_y0;
  wire h_u_cla32_and6169_y0;
  wire h_u_cla32_and6170_y0;
  wire h_u_cla32_and6171_y0;
  wire h_u_cla32_and6172_y0;
  wire h_u_cla32_and6173_y0;
  wire h_u_cla32_and6174_y0;
  wire h_u_cla32_and6175_y0;
  wire h_u_cla32_and6176_y0;
  wire h_u_cla32_and6177_y0;
  wire h_u_cla32_and6178_y0;
  wire h_u_cla32_and6179_y0;
  wire h_u_cla32_and6180_y0;
  wire h_u_cla32_and6181_y0;
  wire h_u_cla32_and6182_y0;
  wire h_u_cla32_and6183_y0;
  wire h_u_cla32_and6184_y0;
  wire h_u_cla32_and6185_y0;
  wire h_u_cla32_and6186_y0;
  wire h_u_cla32_and6187_y0;
  wire h_u_cla32_and6188_y0;
  wire h_u_cla32_and6189_y0;
  wire h_u_cla32_and6190_y0;
  wire h_u_cla32_and6191_y0;
  wire h_u_cla32_and6192_y0;
  wire h_u_cla32_and6193_y0;
  wire h_u_cla32_and6194_y0;
  wire h_u_cla32_and6195_y0;
  wire h_u_cla32_and6196_y0;
  wire h_u_cla32_and6197_y0;
  wire h_u_cla32_and6198_y0;
  wire h_u_cla32_and6199_y0;
  wire h_u_cla32_and6200_y0;
  wire h_u_cla32_or325_y0;
  wire h_u_cla32_or326_y0;
  wire h_u_cla32_or327_y0;
  wire h_u_cla32_or328_y0;
  wire h_u_cla32_or329_y0;
  wire h_u_cla32_or330_y0;
  wire h_u_cla32_or331_y0;
  wire h_u_cla32_or332_y0;
  wire h_u_cla32_or333_y0;
  wire h_u_cla32_or334_y0;
  wire h_u_cla32_or335_y0;
  wire h_u_cla32_or336_y0;
  wire h_u_cla32_or337_y0;
  wire h_u_cla32_or338_y0;
  wire h_u_cla32_or339_y0;
  wire h_u_cla32_or340_y0;
  wire h_u_cla32_or341_y0;
  wire h_u_cla32_or342_y0;
  wire h_u_cla32_or343_y0;
  wire h_u_cla32_or344_y0;
  wire h_u_cla32_or345_y0;
  wire h_u_cla32_or346_y0;
  wire h_u_cla32_or347_y0;
  wire h_u_cla32_or348_y0;
  wire h_u_cla32_or349_y0;
  wire h_u_cla32_or350_y0;
  wire h_u_cla32_pg_logic26_y0;
  wire h_u_cla32_pg_logic26_y1;
  wire h_u_cla32_pg_logic26_y2;
  wire h_u_cla32_xor26_y0;
  wire h_u_cla32_and6201_y0;
  wire h_u_cla32_and6202_y0;
  wire h_u_cla32_and6203_y0;
  wire h_u_cla32_and6204_y0;
  wire h_u_cla32_and6205_y0;
  wire h_u_cla32_and6206_y0;
  wire h_u_cla32_and6207_y0;
  wire h_u_cla32_and6208_y0;
  wire h_u_cla32_and6209_y0;
  wire h_u_cla32_and6210_y0;
  wire h_u_cla32_and6211_y0;
  wire h_u_cla32_and6212_y0;
  wire h_u_cla32_and6213_y0;
  wire h_u_cla32_and6214_y0;
  wire h_u_cla32_and6215_y0;
  wire h_u_cla32_and6216_y0;
  wire h_u_cla32_and6217_y0;
  wire h_u_cla32_and6218_y0;
  wire h_u_cla32_and6219_y0;
  wire h_u_cla32_and6220_y0;
  wire h_u_cla32_and6221_y0;
  wire h_u_cla32_and6222_y0;
  wire h_u_cla32_and6223_y0;
  wire h_u_cla32_and6224_y0;
  wire h_u_cla32_and6225_y0;
  wire h_u_cla32_and6226_y0;
  wire h_u_cla32_and6227_y0;
  wire h_u_cla32_and6228_y0;
  wire h_u_cla32_and6229_y0;
  wire h_u_cla32_and6230_y0;
  wire h_u_cla32_and6231_y0;
  wire h_u_cla32_and6232_y0;
  wire h_u_cla32_and6233_y0;
  wire h_u_cla32_and6234_y0;
  wire h_u_cla32_and6235_y0;
  wire h_u_cla32_and6236_y0;
  wire h_u_cla32_and6237_y0;
  wire h_u_cla32_and6238_y0;
  wire h_u_cla32_and6239_y0;
  wire h_u_cla32_and6240_y0;
  wire h_u_cla32_and6241_y0;
  wire h_u_cla32_and6242_y0;
  wire h_u_cla32_and6243_y0;
  wire h_u_cla32_and6244_y0;
  wire h_u_cla32_and6245_y0;
  wire h_u_cla32_and6246_y0;
  wire h_u_cla32_and6247_y0;
  wire h_u_cla32_and6248_y0;
  wire h_u_cla32_and6249_y0;
  wire h_u_cla32_and6250_y0;
  wire h_u_cla32_and6251_y0;
  wire h_u_cla32_and6252_y0;
  wire h_u_cla32_and6253_y0;
  wire h_u_cla32_and6254_y0;
  wire h_u_cla32_and6255_y0;
  wire h_u_cla32_and6256_y0;
  wire h_u_cla32_and6257_y0;
  wire h_u_cla32_and6258_y0;
  wire h_u_cla32_and6259_y0;
  wire h_u_cla32_and6260_y0;
  wire h_u_cla32_and6261_y0;
  wire h_u_cla32_and6262_y0;
  wire h_u_cla32_and6263_y0;
  wire h_u_cla32_and6264_y0;
  wire h_u_cla32_and6265_y0;
  wire h_u_cla32_and6266_y0;
  wire h_u_cla32_and6267_y0;
  wire h_u_cla32_and6268_y0;
  wire h_u_cla32_and6269_y0;
  wire h_u_cla32_and6270_y0;
  wire h_u_cla32_and6271_y0;
  wire h_u_cla32_and6272_y0;
  wire h_u_cla32_and6273_y0;
  wire h_u_cla32_and6274_y0;
  wire h_u_cla32_and6275_y0;
  wire h_u_cla32_and6276_y0;
  wire h_u_cla32_and6277_y0;
  wire h_u_cla32_and6278_y0;
  wire h_u_cla32_and6279_y0;
  wire h_u_cla32_and6280_y0;
  wire h_u_cla32_and6281_y0;
  wire h_u_cla32_and6282_y0;
  wire h_u_cla32_and6283_y0;
  wire h_u_cla32_and6284_y0;
  wire h_u_cla32_and6285_y0;
  wire h_u_cla32_and6286_y0;
  wire h_u_cla32_and6287_y0;
  wire h_u_cla32_and6288_y0;
  wire h_u_cla32_and6289_y0;
  wire h_u_cla32_and6290_y0;
  wire h_u_cla32_and6291_y0;
  wire h_u_cla32_and6292_y0;
  wire h_u_cla32_and6293_y0;
  wire h_u_cla32_and6294_y0;
  wire h_u_cla32_and6295_y0;
  wire h_u_cla32_and6296_y0;
  wire h_u_cla32_and6297_y0;
  wire h_u_cla32_and6298_y0;
  wire h_u_cla32_and6299_y0;
  wire h_u_cla32_and6300_y0;
  wire h_u_cla32_and6301_y0;
  wire h_u_cla32_and6302_y0;
  wire h_u_cla32_and6303_y0;
  wire h_u_cla32_and6304_y0;
  wire h_u_cla32_and6305_y0;
  wire h_u_cla32_and6306_y0;
  wire h_u_cla32_and6307_y0;
  wire h_u_cla32_and6308_y0;
  wire h_u_cla32_and6309_y0;
  wire h_u_cla32_and6310_y0;
  wire h_u_cla32_and6311_y0;
  wire h_u_cla32_and6312_y0;
  wire h_u_cla32_and6313_y0;
  wire h_u_cla32_and6314_y0;
  wire h_u_cla32_and6315_y0;
  wire h_u_cla32_and6316_y0;
  wire h_u_cla32_and6317_y0;
  wire h_u_cla32_and6318_y0;
  wire h_u_cla32_and6319_y0;
  wire h_u_cla32_and6320_y0;
  wire h_u_cla32_and6321_y0;
  wire h_u_cla32_and6322_y0;
  wire h_u_cla32_and6323_y0;
  wire h_u_cla32_and6324_y0;
  wire h_u_cla32_and6325_y0;
  wire h_u_cla32_and6326_y0;
  wire h_u_cla32_and6327_y0;
  wire h_u_cla32_and6328_y0;
  wire h_u_cla32_and6329_y0;
  wire h_u_cla32_and6330_y0;
  wire h_u_cla32_and6331_y0;
  wire h_u_cla32_and6332_y0;
  wire h_u_cla32_and6333_y0;
  wire h_u_cla32_and6334_y0;
  wire h_u_cla32_and6335_y0;
  wire h_u_cla32_and6336_y0;
  wire h_u_cla32_and6337_y0;
  wire h_u_cla32_and6338_y0;
  wire h_u_cla32_and6339_y0;
  wire h_u_cla32_and6340_y0;
  wire h_u_cla32_and6341_y0;
  wire h_u_cla32_and6342_y0;
  wire h_u_cla32_and6343_y0;
  wire h_u_cla32_and6344_y0;
  wire h_u_cla32_and6345_y0;
  wire h_u_cla32_and6346_y0;
  wire h_u_cla32_and6347_y0;
  wire h_u_cla32_and6348_y0;
  wire h_u_cla32_and6349_y0;
  wire h_u_cla32_and6350_y0;
  wire h_u_cla32_and6351_y0;
  wire h_u_cla32_and6352_y0;
  wire h_u_cla32_and6353_y0;
  wire h_u_cla32_and6354_y0;
  wire h_u_cla32_and6355_y0;
  wire h_u_cla32_and6356_y0;
  wire h_u_cla32_and6357_y0;
  wire h_u_cla32_and6358_y0;
  wire h_u_cla32_and6359_y0;
  wire h_u_cla32_and6360_y0;
  wire h_u_cla32_and6361_y0;
  wire h_u_cla32_and6362_y0;
  wire h_u_cla32_and6363_y0;
  wire h_u_cla32_and6364_y0;
  wire h_u_cla32_and6365_y0;
  wire h_u_cla32_and6366_y0;
  wire h_u_cla32_and6367_y0;
  wire h_u_cla32_and6368_y0;
  wire h_u_cla32_and6369_y0;
  wire h_u_cla32_and6370_y0;
  wire h_u_cla32_and6371_y0;
  wire h_u_cla32_and6372_y0;
  wire h_u_cla32_and6373_y0;
  wire h_u_cla32_and6374_y0;
  wire h_u_cla32_and6375_y0;
  wire h_u_cla32_and6376_y0;
  wire h_u_cla32_and6377_y0;
  wire h_u_cla32_and6378_y0;
  wire h_u_cla32_and6379_y0;
  wire h_u_cla32_and6380_y0;
  wire h_u_cla32_and6381_y0;
  wire h_u_cla32_and6382_y0;
  wire h_u_cla32_and6383_y0;
  wire h_u_cla32_and6384_y0;
  wire h_u_cla32_and6385_y0;
  wire h_u_cla32_and6386_y0;
  wire h_u_cla32_and6387_y0;
  wire h_u_cla32_and6388_y0;
  wire h_u_cla32_and6389_y0;
  wire h_u_cla32_and6390_y0;
  wire h_u_cla32_and6391_y0;
  wire h_u_cla32_and6392_y0;
  wire h_u_cla32_and6393_y0;
  wire h_u_cla32_and6394_y0;
  wire h_u_cla32_and6395_y0;
  wire h_u_cla32_and6396_y0;
  wire h_u_cla32_and6397_y0;
  wire h_u_cla32_and6398_y0;
  wire h_u_cla32_and6399_y0;
  wire h_u_cla32_and6400_y0;
  wire h_u_cla32_and6401_y0;
  wire h_u_cla32_and6402_y0;
  wire h_u_cla32_and6403_y0;
  wire h_u_cla32_and6404_y0;
  wire h_u_cla32_and6405_y0;
  wire h_u_cla32_and6406_y0;
  wire h_u_cla32_and6407_y0;
  wire h_u_cla32_and6408_y0;
  wire h_u_cla32_and6409_y0;
  wire h_u_cla32_and6410_y0;
  wire h_u_cla32_and6411_y0;
  wire h_u_cla32_and6412_y0;
  wire h_u_cla32_and6413_y0;
  wire h_u_cla32_and6414_y0;
  wire h_u_cla32_and6415_y0;
  wire h_u_cla32_and6416_y0;
  wire h_u_cla32_and6417_y0;
  wire h_u_cla32_and6418_y0;
  wire h_u_cla32_and6419_y0;
  wire h_u_cla32_and6420_y0;
  wire h_u_cla32_and6421_y0;
  wire h_u_cla32_and6422_y0;
  wire h_u_cla32_and6423_y0;
  wire h_u_cla32_and6424_y0;
  wire h_u_cla32_and6425_y0;
  wire h_u_cla32_and6426_y0;
  wire h_u_cla32_and6427_y0;
  wire h_u_cla32_and6428_y0;
  wire h_u_cla32_and6429_y0;
  wire h_u_cla32_and6430_y0;
  wire h_u_cla32_and6431_y0;
  wire h_u_cla32_and6432_y0;
  wire h_u_cla32_and6433_y0;
  wire h_u_cla32_and6434_y0;
  wire h_u_cla32_and6435_y0;
  wire h_u_cla32_and6436_y0;
  wire h_u_cla32_and6437_y0;
  wire h_u_cla32_and6438_y0;
  wire h_u_cla32_and6439_y0;
  wire h_u_cla32_and6440_y0;
  wire h_u_cla32_and6441_y0;
  wire h_u_cla32_and6442_y0;
  wire h_u_cla32_and6443_y0;
  wire h_u_cla32_and6444_y0;
  wire h_u_cla32_and6445_y0;
  wire h_u_cla32_and6446_y0;
  wire h_u_cla32_and6447_y0;
  wire h_u_cla32_and6448_y0;
  wire h_u_cla32_and6449_y0;
  wire h_u_cla32_and6450_y0;
  wire h_u_cla32_and6451_y0;
  wire h_u_cla32_and6452_y0;
  wire h_u_cla32_and6453_y0;
  wire h_u_cla32_and6454_y0;
  wire h_u_cla32_and6455_y0;
  wire h_u_cla32_and6456_y0;
  wire h_u_cla32_and6457_y0;
  wire h_u_cla32_and6458_y0;
  wire h_u_cla32_and6459_y0;
  wire h_u_cla32_and6460_y0;
  wire h_u_cla32_and6461_y0;
  wire h_u_cla32_and6462_y0;
  wire h_u_cla32_and6463_y0;
  wire h_u_cla32_and6464_y0;
  wire h_u_cla32_and6465_y0;
  wire h_u_cla32_and6466_y0;
  wire h_u_cla32_and6467_y0;
  wire h_u_cla32_and6468_y0;
  wire h_u_cla32_and6469_y0;
  wire h_u_cla32_and6470_y0;
  wire h_u_cla32_and6471_y0;
  wire h_u_cla32_and6472_y0;
  wire h_u_cla32_and6473_y0;
  wire h_u_cla32_and6474_y0;
  wire h_u_cla32_and6475_y0;
  wire h_u_cla32_and6476_y0;
  wire h_u_cla32_and6477_y0;
  wire h_u_cla32_and6478_y0;
  wire h_u_cla32_and6479_y0;
  wire h_u_cla32_and6480_y0;
  wire h_u_cla32_and6481_y0;
  wire h_u_cla32_and6482_y0;
  wire h_u_cla32_and6483_y0;
  wire h_u_cla32_and6484_y0;
  wire h_u_cla32_and6485_y0;
  wire h_u_cla32_and6486_y0;
  wire h_u_cla32_and6487_y0;
  wire h_u_cla32_and6488_y0;
  wire h_u_cla32_and6489_y0;
  wire h_u_cla32_and6490_y0;
  wire h_u_cla32_and6491_y0;
  wire h_u_cla32_and6492_y0;
  wire h_u_cla32_and6493_y0;
  wire h_u_cla32_and6494_y0;
  wire h_u_cla32_and6495_y0;
  wire h_u_cla32_and6496_y0;
  wire h_u_cla32_and6497_y0;
  wire h_u_cla32_and6498_y0;
  wire h_u_cla32_and6499_y0;
  wire h_u_cla32_and6500_y0;
  wire h_u_cla32_and6501_y0;
  wire h_u_cla32_and6502_y0;
  wire h_u_cla32_and6503_y0;
  wire h_u_cla32_and6504_y0;
  wire h_u_cla32_and6505_y0;
  wire h_u_cla32_and6506_y0;
  wire h_u_cla32_and6507_y0;
  wire h_u_cla32_and6508_y0;
  wire h_u_cla32_and6509_y0;
  wire h_u_cla32_and6510_y0;
  wire h_u_cla32_and6511_y0;
  wire h_u_cla32_and6512_y0;
  wire h_u_cla32_and6513_y0;
  wire h_u_cla32_and6514_y0;
  wire h_u_cla32_and6515_y0;
  wire h_u_cla32_and6516_y0;
  wire h_u_cla32_and6517_y0;
  wire h_u_cla32_and6518_y0;
  wire h_u_cla32_and6519_y0;
  wire h_u_cla32_and6520_y0;
  wire h_u_cla32_and6521_y0;
  wire h_u_cla32_and6522_y0;
  wire h_u_cla32_and6523_y0;
  wire h_u_cla32_and6524_y0;
  wire h_u_cla32_and6525_y0;
  wire h_u_cla32_and6526_y0;
  wire h_u_cla32_and6527_y0;
  wire h_u_cla32_and6528_y0;
  wire h_u_cla32_and6529_y0;
  wire h_u_cla32_and6530_y0;
  wire h_u_cla32_and6531_y0;
  wire h_u_cla32_and6532_y0;
  wire h_u_cla32_and6533_y0;
  wire h_u_cla32_and6534_y0;
  wire h_u_cla32_and6535_y0;
  wire h_u_cla32_and6536_y0;
  wire h_u_cla32_and6537_y0;
  wire h_u_cla32_and6538_y0;
  wire h_u_cla32_and6539_y0;
  wire h_u_cla32_and6540_y0;
  wire h_u_cla32_and6541_y0;
  wire h_u_cla32_and6542_y0;
  wire h_u_cla32_and6543_y0;
  wire h_u_cla32_and6544_y0;
  wire h_u_cla32_and6545_y0;
  wire h_u_cla32_and6546_y0;
  wire h_u_cla32_and6547_y0;
  wire h_u_cla32_and6548_y0;
  wire h_u_cla32_and6549_y0;
  wire h_u_cla32_and6550_y0;
  wire h_u_cla32_and6551_y0;
  wire h_u_cla32_and6552_y0;
  wire h_u_cla32_and6553_y0;
  wire h_u_cla32_and6554_y0;
  wire h_u_cla32_and6555_y0;
  wire h_u_cla32_and6556_y0;
  wire h_u_cla32_and6557_y0;
  wire h_u_cla32_and6558_y0;
  wire h_u_cla32_and6559_y0;
  wire h_u_cla32_and6560_y0;
  wire h_u_cla32_and6561_y0;
  wire h_u_cla32_and6562_y0;
  wire h_u_cla32_and6563_y0;
  wire h_u_cla32_and6564_y0;
  wire h_u_cla32_and6565_y0;
  wire h_u_cla32_and6566_y0;
  wire h_u_cla32_and6567_y0;
  wire h_u_cla32_and6568_y0;
  wire h_u_cla32_and6569_y0;
  wire h_u_cla32_and6570_y0;
  wire h_u_cla32_and6571_y0;
  wire h_u_cla32_and6572_y0;
  wire h_u_cla32_and6573_y0;
  wire h_u_cla32_and6574_y0;
  wire h_u_cla32_and6575_y0;
  wire h_u_cla32_and6576_y0;
  wire h_u_cla32_and6577_y0;
  wire h_u_cla32_and6578_y0;
  wire h_u_cla32_and6579_y0;
  wire h_u_cla32_and6580_y0;
  wire h_u_cla32_and6581_y0;
  wire h_u_cla32_and6582_y0;
  wire h_u_cla32_and6583_y0;
  wire h_u_cla32_and6584_y0;
  wire h_u_cla32_and6585_y0;
  wire h_u_cla32_and6586_y0;
  wire h_u_cla32_and6587_y0;
  wire h_u_cla32_and6588_y0;
  wire h_u_cla32_and6589_y0;
  wire h_u_cla32_and6590_y0;
  wire h_u_cla32_and6591_y0;
  wire h_u_cla32_and6592_y0;
  wire h_u_cla32_and6593_y0;
  wire h_u_cla32_and6594_y0;
  wire h_u_cla32_and6595_y0;
  wire h_u_cla32_and6596_y0;
  wire h_u_cla32_and6597_y0;
  wire h_u_cla32_and6598_y0;
  wire h_u_cla32_and6599_y0;
  wire h_u_cla32_and6600_y0;
  wire h_u_cla32_and6601_y0;
  wire h_u_cla32_and6602_y0;
  wire h_u_cla32_and6603_y0;
  wire h_u_cla32_and6604_y0;
  wire h_u_cla32_and6605_y0;
  wire h_u_cla32_and6606_y0;
  wire h_u_cla32_and6607_y0;
  wire h_u_cla32_and6608_y0;
  wire h_u_cla32_and6609_y0;
  wire h_u_cla32_and6610_y0;
  wire h_u_cla32_and6611_y0;
  wire h_u_cla32_and6612_y0;
  wire h_u_cla32_and6613_y0;
  wire h_u_cla32_and6614_y0;
  wire h_u_cla32_and6615_y0;
  wire h_u_cla32_and6616_y0;
  wire h_u_cla32_and6617_y0;
  wire h_u_cla32_and6618_y0;
  wire h_u_cla32_and6619_y0;
  wire h_u_cla32_and6620_y0;
  wire h_u_cla32_and6621_y0;
  wire h_u_cla32_and6622_y0;
  wire h_u_cla32_and6623_y0;
  wire h_u_cla32_and6624_y0;
  wire h_u_cla32_and6625_y0;
  wire h_u_cla32_and6626_y0;
  wire h_u_cla32_and6627_y0;
  wire h_u_cla32_and6628_y0;
  wire h_u_cla32_and6629_y0;
  wire h_u_cla32_and6630_y0;
  wire h_u_cla32_and6631_y0;
  wire h_u_cla32_and6632_y0;
  wire h_u_cla32_and6633_y0;
  wire h_u_cla32_and6634_y0;
  wire h_u_cla32_and6635_y0;
  wire h_u_cla32_and6636_y0;
  wire h_u_cla32_and6637_y0;
  wire h_u_cla32_and6638_y0;
  wire h_u_cla32_and6639_y0;
  wire h_u_cla32_and6640_y0;
  wire h_u_cla32_and6641_y0;
  wire h_u_cla32_and6642_y0;
  wire h_u_cla32_and6643_y0;
  wire h_u_cla32_and6644_y0;
  wire h_u_cla32_and6645_y0;
  wire h_u_cla32_and6646_y0;
  wire h_u_cla32_and6647_y0;
  wire h_u_cla32_and6648_y0;
  wire h_u_cla32_and6649_y0;
  wire h_u_cla32_and6650_y0;
  wire h_u_cla32_and6651_y0;
  wire h_u_cla32_and6652_y0;
  wire h_u_cla32_and6653_y0;
  wire h_u_cla32_and6654_y0;
  wire h_u_cla32_and6655_y0;
  wire h_u_cla32_and6656_y0;
  wire h_u_cla32_and6657_y0;
  wire h_u_cla32_and6658_y0;
  wire h_u_cla32_and6659_y0;
  wire h_u_cla32_and6660_y0;
  wire h_u_cla32_and6661_y0;
  wire h_u_cla32_and6662_y0;
  wire h_u_cla32_and6663_y0;
  wire h_u_cla32_and6664_y0;
  wire h_u_cla32_and6665_y0;
  wire h_u_cla32_and6666_y0;
  wire h_u_cla32_and6667_y0;
  wire h_u_cla32_and6668_y0;
  wire h_u_cla32_and6669_y0;
  wire h_u_cla32_and6670_y0;
  wire h_u_cla32_and6671_y0;
  wire h_u_cla32_and6672_y0;
  wire h_u_cla32_and6673_y0;
  wire h_u_cla32_and6674_y0;
  wire h_u_cla32_and6675_y0;
  wire h_u_cla32_and6676_y0;
  wire h_u_cla32_and6677_y0;
  wire h_u_cla32_and6678_y0;
  wire h_u_cla32_and6679_y0;
  wire h_u_cla32_and6680_y0;
  wire h_u_cla32_and6681_y0;
  wire h_u_cla32_and6682_y0;
  wire h_u_cla32_and6683_y0;
  wire h_u_cla32_and6684_y0;
  wire h_u_cla32_and6685_y0;
  wire h_u_cla32_and6686_y0;
  wire h_u_cla32_and6687_y0;
  wire h_u_cla32_and6688_y0;
  wire h_u_cla32_and6689_y0;
  wire h_u_cla32_and6690_y0;
  wire h_u_cla32_and6691_y0;
  wire h_u_cla32_and6692_y0;
  wire h_u_cla32_and6693_y0;
  wire h_u_cla32_and6694_y0;
  wire h_u_cla32_and6695_y0;
  wire h_u_cla32_and6696_y0;
  wire h_u_cla32_and6697_y0;
  wire h_u_cla32_and6698_y0;
  wire h_u_cla32_and6699_y0;
  wire h_u_cla32_and6700_y0;
  wire h_u_cla32_and6701_y0;
  wire h_u_cla32_and6702_y0;
  wire h_u_cla32_and6703_y0;
  wire h_u_cla32_and6704_y0;
  wire h_u_cla32_and6705_y0;
  wire h_u_cla32_and6706_y0;
  wire h_u_cla32_and6707_y0;
  wire h_u_cla32_and6708_y0;
  wire h_u_cla32_and6709_y0;
  wire h_u_cla32_and6710_y0;
  wire h_u_cla32_and6711_y0;
  wire h_u_cla32_and6712_y0;
  wire h_u_cla32_and6713_y0;
  wire h_u_cla32_and6714_y0;
  wire h_u_cla32_and6715_y0;
  wire h_u_cla32_and6716_y0;
  wire h_u_cla32_and6717_y0;
  wire h_u_cla32_and6718_y0;
  wire h_u_cla32_and6719_y0;
  wire h_u_cla32_and6720_y0;
  wire h_u_cla32_and6721_y0;
  wire h_u_cla32_and6722_y0;
  wire h_u_cla32_and6723_y0;
  wire h_u_cla32_and6724_y0;
  wire h_u_cla32_and6725_y0;
  wire h_u_cla32_and6726_y0;
  wire h_u_cla32_and6727_y0;
  wire h_u_cla32_and6728_y0;
  wire h_u_cla32_and6729_y0;
  wire h_u_cla32_and6730_y0;
  wire h_u_cla32_and6731_y0;
  wire h_u_cla32_and6732_y0;
  wire h_u_cla32_and6733_y0;
  wire h_u_cla32_and6734_y0;
  wire h_u_cla32_and6735_y0;
  wire h_u_cla32_and6736_y0;
  wire h_u_cla32_and6737_y0;
  wire h_u_cla32_and6738_y0;
  wire h_u_cla32_and6739_y0;
  wire h_u_cla32_and6740_y0;
  wire h_u_cla32_and6741_y0;
  wire h_u_cla32_and6742_y0;
  wire h_u_cla32_and6743_y0;
  wire h_u_cla32_and6744_y0;
  wire h_u_cla32_and6745_y0;
  wire h_u_cla32_and6746_y0;
  wire h_u_cla32_and6747_y0;
  wire h_u_cla32_and6748_y0;
  wire h_u_cla32_and6749_y0;
  wire h_u_cla32_and6750_y0;
  wire h_u_cla32_and6751_y0;
  wire h_u_cla32_and6752_y0;
  wire h_u_cla32_and6753_y0;
  wire h_u_cla32_and6754_y0;
  wire h_u_cla32_and6755_y0;
  wire h_u_cla32_and6756_y0;
  wire h_u_cla32_and6757_y0;
  wire h_u_cla32_and6758_y0;
  wire h_u_cla32_and6759_y0;
  wire h_u_cla32_and6760_y0;
  wire h_u_cla32_and6761_y0;
  wire h_u_cla32_and6762_y0;
  wire h_u_cla32_and6763_y0;
  wire h_u_cla32_and6764_y0;
  wire h_u_cla32_and6765_y0;
  wire h_u_cla32_and6766_y0;
  wire h_u_cla32_and6767_y0;
  wire h_u_cla32_and6768_y0;
  wire h_u_cla32_and6769_y0;
  wire h_u_cla32_and6770_y0;
  wire h_u_cla32_and6771_y0;
  wire h_u_cla32_and6772_y0;
  wire h_u_cla32_and6773_y0;
  wire h_u_cla32_and6774_y0;
  wire h_u_cla32_and6775_y0;
  wire h_u_cla32_and6776_y0;
  wire h_u_cla32_and6777_y0;
  wire h_u_cla32_and6778_y0;
  wire h_u_cla32_and6779_y0;
  wire h_u_cla32_and6780_y0;
  wire h_u_cla32_and6781_y0;
  wire h_u_cla32_and6782_y0;
  wire h_u_cla32_and6783_y0;
  wire h_u_cla32_and6784_y0;
  wire h_u_cla32_and6785_y0;
  wire h_u_cla32_and6786_y0;
  wire h_u_cla32_and6787_y0;
  wire h_u_cla32_and6788_y0;
  wire h_u_cla32_and6789_y0;
  wire h_u_cla32_and6790_y0;
  wire h_u_cla32_and6791_y0;
  wire h_u_cla32_and6792_y0;
  wire h_u_cla32_and6793_y0;
  wire h_u_cla32_and6794_y0;
  wire h_u_cla32_and6795_y0;
  wire h_u_cla32_and6796_y0;
  wire h_u_cla32_and6797_y0;
  wire h_u_cla32_and6798_y0;
  wire h_u_cla32_and6799_y0;
  wire h_u_cla32_and6800_y0;
  wire h_u_cla32_and6801_y0;
  wire h_u_cla32_and6802_y0;
  wire h_u_cla32_and6803_y0;
  wire h_u_cla32_and6804_y0;
  wire h_u_cla32_and6805_y0;
  wire h_u_cla32_and6806_y0;
  wire h_u_cla32_and6807_y0;
  wire h_u_cla32_and6808_y0;
  wire h_u_cla32_and6809_y0;
  wire h_u_cla32_and6810_y0;
  wire h_u_cla32_and6811_y0;
  wire h_u_cla32_and6812_y0;
  wire h_u_cla32_and6813_y0;
  wire h_u_cla32_and6814_y0;
  wire h_u_cla32_and6815_y0;
  wire h_u_cla32_and6816_y0;
  wire h_u_cla32_and6817_y0;
  wire h_u_cla32_and6818_y0;
  wire h_u_cla32_and6819_y0;
  wire h_u_cla32_and6820_y0;
  wire h_u_cla32_and6821_y0;
  wire h_u_cla32_and6822_y0;
  wire h_u_cla32_and6823_y0;
  wire h_u_cla32_and6824_y0;
  wire h_u_cla32_and6825_y0;
  wire h_u_cla32_and6826_y0;
  wire h_u_cla32_and6827_y0;
  wire h_u_cla32_and6828_y0;
  wire h_u_cla32_and6829_y0;
  wire h_u_cla32_and6830_y0;
  wire h_u_cla32_and6831_y0;
  wire h_u_cla32_and6832_y0;
  wire h_u_cla32_and6833_y0;
  wire h_u_cla32_and6834_y0;
  wire h_u_cla32_and6835_y0;
  wire h_u_cla32_and6836_y0;
  wire h_u_cla32_and6837_y0;
  wire h_u_cla32_and6838_y0;
  wire h_u_cla32_and6839_y0;
  wire h_u_cla32_and6840_y0;
  wire h_u_cla32_and6841_y0;
  wire h_u_cla32_and6842_y0;
  wire h_u_cla32_and6843_y0;
  wire h_u_cla32_and6844_y0;
  wire h_u_cla32_and6845_y0;
  wire h_u_cla32_and6846_y0;
  wire h_u_cla32_and6847_y0;
  wire h_u_cla32_and6848_y0;
  wire h_u_cla32_and6849_y0;
  wire h_u_cla32_and6850_y0;
  wire h_u_cla32_and6851_y0;
  wire h_u_cla32_and6852_y0;
  wire h_u_cla32_and6853_y0;
  wire h_u_cla32_and6854_y0;
  wire h_u_cla32_and6855_y0;
  wire h_u_cla32_and6856_y0;
  wire h_u_cla32_and6857_y0;
  wire h_u_cla32_and6858_y0;
  wire h_u_cla32_and6859_y0;
  wire h_u_cla32_and6860_y0;
  wire h_u_cla32_and6861_y0;
  wire h_u_cla32_and6862_y0;
  wire h_u_cla32_and6863_y0;
  wire h_u_cla32_and6864_y0;
  wire h_u_cla32_and6865_y0;
  wire h_u_cla32_and6866_y0;
  wire h_u_cla32_and6867_y0;
  wire h_u_cla32_and6868_y0;
  wire h_u_cla32_and6869_y0;
  wire h_u_cla32_and6870_y0;
  wire h_u_cla32_and6871_y0;
  wire h_u_cla32_and6872_y0;
  wire h_u_cla32_and6873_y0;
  wire h_u_cla32_and6874_y0;
  wire h_u_cla32_and6875_y0;
  wire h_u_cla32_and6876_y0;
  wire h_u_cla32_and6877_y0;
  wire h_u_cla32_and6878_y0;
  wire h_u_cla32_and6879_y0;
  wire h_u_cla32_and6880_y0;
  wire h_u_cla32_and6881_y0;
  wire h_u_cla32_and6882_y0;
  wire h_u_cla32_and6883_y0;
  wire h_u_cla32_and6884_y0;
  wire h_u_cla32_and6885_y0;
  wire h_u_cla32_and6886_y0;
  wire h_u_cla32_and6887_y0;
  wire h_u_cla32_and6888_y0;
  wire h_u_cla32_and6889_y0;
  wire h_u_cla32_and6890_y0;
  wire h_u_cla32_and6891_y0;
  wire h_u_cla32_and6892_y0;
  wire h_u_cla32_and6893_y0;
  wire h_u_cla32_and6894_y0;
  wire h_u_cla32_and6895_y0;
  wire h_u_cla32_and6896_y0;
  wire h_u_cla32_and6897_y0;
  wire h_u_cla32_and6898_y0;
  wire h_u_cla32_and6899_y0;
  wire h_u_cla32_and6900_y0;
  wire h_u_cla32_and6901_y0;
  wire h_u_cla32_and6902_y0;
  wire h_u_cla32_and6903_y0;
  wire h_u_cla32_and6904_y0;
  wire h_u_cla32_and6905_y0;
  wire h_u_cla32_and6906_y0;
  wire h_u_cla32_and6907_y0;
  wire h_u_cla32_and6908_y0;
  wire h_u_cla32_and6909_y0;
  wire h_u_cla32_and6910_y0;
  wire h_u_cla32_and6911_y0;
  wire h_u_cla32_and6912_y0;
  wire h_u_cla32_and6913_y0;
  wire h_u_cla32_and6914_y0;
  wire h_u_cla32_and6915_y0;
  wire h_u_cla32_and6916_y0;
  wire h_u_cla32_and6917_y0;
  wire h_u_cla32_and6918_y0;
  wire h_u_cla32_and6919_y0;
  wire h_u_cla32_and6920_y0;
  wire h_u_cla32_and6921_y0;
  wire h_u_cla32_and6922_y0;
  wire h_u_cla32_and6923_y0;
  wire h_u_cla32_and6924_y0;
  wire h_u_cla32_and6925_y0;
  wire h_u_cla32_and6926_y0;
  wire h_u_cla32_and6927_y0;
  wire h_u_cla32_and6928_y0;
  wire h_u_cla32_and6929_y0;
  wire h_u_cla32_or351_y0;
  wire h_u_cla32_or352_y0;
  wire h_u_cla32_or353_y0;
  wire h_u_cla32_or354_y0;
  wire h_u_cla32_or355_y0;
  wire h_u_cla32_or356_y0;
  wire h_u_cla32_or357_y0;
  wire h_u_cla32_or358_y0;
  wire h_u_cla32_or359_y0;
  wire h_u_cla32_or360_y0;
  wire h_u_cla32_or361_y0;
  wire h_u_cla32_or362_y0;
  wire h_u_cla32_or363_y0;
  wire h_u_cla32_or364_y0;
  wire h_u_cla32_or365_y0;
  wire h_u_cla32_or366_y0;
  wire h_u_cla32_or367_y0;
  wire h_u_cla32_or368_y0;
  wire h_u_cla32_or369_y0;
  wire h_u_cla32_or370_y0;
  wire h_u_cla32_or371_y0;
  wire h_u_cla32_or372_y0;
  wire h_u_cla32_or373_y0;
  wire h_u_cla32_or374_y0;
  wire h_u_cla32_or375_y0;
  wire h_u_cla32_or376_y0;
  wire h_u_cla32_or377_y0;
  wire h_u_cla32_pg_logic27_y0;
  wire h_u_cla32_pg_logic27_y1;
  wire h_u_cla32_pg_logic27_y2;
  wire h_u_cla32_xor27_y0;
  wire h_u_cla32_and6930_y0;
  wire h_u_cla32_and6931_y0;
  wire h_u_cla32_and6932_y0;
  wire h_u_cla32_and6933_y0;
  wire h_u_cla32_and6934_y0;
  wire h_u_cla32_and6935_y0;
  wire h_u_cla32_and6936_y0;
  wire h_u_cla32_and6937_y0;
  wire h_u_cla32_and6938_y0;
  wire h_u_cla32_and6939_y0;
  wire h_u_cla32_and6940_y0;
  wire h_u_cla32_and6941_y0;
  wire h_u_cla32_and6942_y0;
  wire h_u_cla32_and6943_y0;
  wire h_u_cla32_and6944_y0;
  wire h_u_cla32_and6945_y0;
  wire h_u_cla32_and6946_y0;
  wire h_u_cla32_and6947_y0;
  wire h_u_cla32_and6948_y0;
  wire h_u_cla32_and6949_y0;
  wire h_u_cla32_and6950_y0;
  wire h_u_cla32_and6951_y0;
  wire h_u_cla32_and6952_y0;
  wire h_u_cla32_and6953_y0;
  wire h_u_cla32_and6954_y0;
  wire h_u_cla32_and6955_y0;
  wire h_u_cla32_and6956_y0;
  wire h_u_cla32_and6957_y0;
  wire h_u_cla32_and6958_y0;
  wire h_u_cla32_and6959_y0;
  wire h_u_cla32_and6960_y0;
  wire h_u_cla32_and6961_y0;
  wire h_u_cla32_and6962_y0;
  wire h_u_cla32_and6963_y0;
  wire h_u_cla32_and6964_y0;
  wire h_u_cla32_and6965_y0;
  wire h_u_cla32_and6966_y0;
  wire h_u_cla32_and6967_y0;
  wire h_u_cla32_and6968_y0;
  wire h_u_cla32_and6969_y0;
  wire h_u_cla32_and6970_y0;
  wire h_u_cla32_and6971_y0;
  wire h_u_cla32_and6972_y0;
  wire h_u_cla32_and6973_y0;
  wire h_u_cla32_and6974_y0;
  wire h_u_cla32_and6975_y0;
  wire h_u_cla32_and6976_y0;
  wire h_u_cla32_and6977_y0;
  wire h_u_cla32_and6978_y0;
  wire h_u_cla32_and6979_y0;
  wire h_u_cla32_and6980_y0;
  wire h_u_cla32_and6981_y0;
  wire h_u_cla32_and6982_y0;
  wire h_u_cla32_and6983_y0;
  wire h_u_cla32_and6984_y0;
  wire h_u_cla32_and6985_y0;
  wire h_u_cla32_and6986_y0;
  wire h_u_cla32_and6987_y0;
  wire h_u_cla32_and6988_y0;
  wire h_u_cla32_and6989_y0;
  wire h_u_cla32_and6990_y0;
  wire h_u_cla32_and6991_y0;
  wire h_u_cla32_and6992_y0;
  wire h_u_cla32_and6993_y0;
  wire h_u_cla32_and6994_y0;
  wire h_u_cla32_and6995_y0;
  wire h_u_cla32_and6996_y0;
  wire h_u_cla32_and6997_y0;
  wire h_u_cla32_and6998_y0;
  wire h_u_cla32_and6999_y0;
  wire h_u_cla32_and7000_y0;
  wire h_u_cla32_and7001_y0;
  wire h_u_cla32_and7002_y0;
  wire h_u_cla32_and7003_y0;
  wire h_u_cla32_and7004_y0;
  wire h_u_cla32_and7005_y0;
  wire h_u_cla32_and7006_y0;
  wire h_u_cla32_and7007_y0;
  wire h_u_cla32_and7008_y0;
  wire h_u_cla32_and7009_y0;
  wire h_u_cla32_and7010_y0;
  wire h_u_cla32_and7011_y0;
  wire h_u_cla32_and7012_y0;
  wire h_u_cla32_and7013_y0;
  wire h_u_cla32_and7014_y0;
  wire h_u_cla32_and7015_y0;
  wire h_u_cla32_and7016_y0;
  wire h_u_cla32_and7017_y0;
  wire h_u_cla32_and7018_y0;
  wire h_u_cla32_and7019_y0;
  wire h_u_cla32_and7020_y0;
  wire h_u_cla32_and7021_y0;
  wire h_u_cla32_and7022_y0;
  wire h_u_cla32_and7023_y0;
  wire h_u_cla32_and7024_y0;
  wire h_u_cla32_and7025_y0;
  wire h_u_cla32_and7026_y0;
  wire h_u_cla32_and7027_y0;
  wire h_u_cla32_and7028_y0;
  wire h_u_cla32_and7029_y0;
  wire h_u_cla32_and7030_y0;
  wire h_u_cla32_and7031_y0;
  wire h_u_cla32_and7032_y0;
  wire h_u_cla32_and7033_y0;
  wire h_u_cla32_and7034_y0;
  wire h_u_cla32_and7035_y0;
  wire h_u_cla32_and7036_y0;
  wire h_u_cla32_and7037_y0;
  wire h_u_cla32_and7038_y0;
  wire h_u_cla32_and7039_y0;
  wire h_u_cla32_and7040_y0;
  wire h_u_cla32_and7041_y0;
  wire h_u_cla32_and7042_y0;
  wire h_u_cla32_and7043_y0;
  wire h_u_cla32_and7044_y0;
  wire h_u_cla32_and7045_y0;
  wire h_u_cla32_and7046_y0;
  wire h_u_cla32_and7047_y0;
  wire h_u_cla32_and7048_y0;
  wire h_u_cla32_and7049_y0;
  wire h_u_cla32_and7050_y0;
  wire h_u_cla32_and7051_y0;
  wire h_u_cla32_and7052_y0;
  wire h_u_cla32_and7053_y0;
  wire h_u_cla32_and7054_y0;
  wire h_u_cla32_and7055_y0;
  wire h_u_cla32_and7056_y0;
  wire h_u_cla32_and7057_y0;
  wire h_u_cla32_and7058_y0;
  wire h_u_cla32_and7059_y0;
  wire h_u_cla32_and7060_y0;
  wire h_u_cla32_and7061_y0;
  wire h_u_cla32_and7062_y0;
  wire h_u_cla32_and7063_y0;
  wire h_u_cla32_and7064_y0;
  wire h_u_cla32_and7065_y0;
  wire h_u_cla32_and7066_y0;
  wire h_u_cla32_and7067_y0;
  wire h_u_cla32_and7068_y0;
  wire h_u_cla32_and7069_y0;
  wire h_u_cla32_and7070_y0;
  wire h_u_cla32_and7071_y0;
  wire h_u_cla32_and7072_y0;
  wire h_u_cla32_and7073_y0;
  wire h_u_cla32_and7074_y0;
  wire h_u_cla32_and7075_y0;
  wire h_u_cla32_and7076_y0;
  wire h_u_cla32_and7077_y0;
  wire h_u_cla32_and7078_y0;
  wire h_u_cla32_and7079_y0;
  wire h_u_cla32_and7080_y0;
  wire h_u_cla32_and7081_y0;
  wire h_u_cla32_and7082_y0;
  wire h_u_cla32_and7083_y0;
  wire h_u_cla32_and7084_y0;
  wire h_u_cla32_and7085_y0;
  wire h_u_cla32_and7086_y0;
  wire h_u_cla32_and7087_y0;
  wire h_u_cla32_and7088_y0;
  wire h_u_cla32_and7089_y0;
  wire h_u_cla32_and7090_y0;
  wire h_u_cla32_and7091_y0;
  wire h_u_cla32_and7092_y0;
  wire h_u_cla32_and7093_y0;
  wire h_u_cla32_and7094_y0;
  wire h_u_cla32_and7095_y0;
  wire h_u_cla32_and7096_y0;
  wire h_u_cla32_and7097_y0;
  wire h_u_cla32_and7098_y0;
  wire h_u_cla32_and7099_y0;
  wire h_u_cla32_and7100_y0;
  wire h_u_cla32_and7101_y0;
  wire h_u_cla32_and7102_y0;
  wire h_u_cla32_and7103_y0;
  wire h_u_cla32_and7104_y0;
  wire h_u_cla32_and7105_y0;
  wire h_u_cla32_and7106_y0;
  wire h_u_cla32_and7107_y0;
  wire h_u_cla32_and7108_y0;
  wire h_u_cla32_and7109_y0;
  wire h_u_cla32_and7110_y0;
  wire h_u_cla32_and7111_y0;
  wire h_u_cla32_and7112_y0;
  wire h_u_cla32_and7113_y0;
  wire h_u_cla32_and7114_y0;
  wire h_u_cla32_and7115_y0;
  wire h_u_cla32_and7116_y0;
  wire h_u_cla32_and7117_y0;
  wire h_u_cla32_and7118_y0;
  wire h_u_cla32_and7119_y0;
  wire h_u_cla32_and7120_y0;
  wire h_u_cla32_and7121_y0;
  wire h_u_cla32_and7122_y0;
  wire h_u_cla32_and7123_y0;
  wire h_u_cla32_and7124_y0;
  wire h_u_cla32_and7125_y0;
  wire h_u_cla32_and7126_y0;
  wire h_u_cla32_and7127_y0;
  wire h_u_cla32_and7128_y0;
  wire h_u_cla32_and7129_y0;
  wire h_u_cla32_and7130_y0;
  wire h_u_cla32_and7131_y0;
  wire h_u_cla32_and7132_y0;
  wire h_u_cla32_and7133_y0;
  wire h_u_cla32_and7134_y0;
  wire h_u_cla32_and7135_y0;
  wire h_u_cla32_and7136_y0;
  wire h_u_cla32_and7137_y0;
  wire h_u_cla32_and7138_y0;
  wire h_u_cla32_and7139_y0;
  wire h_u_cla32_and7140_y0;
  wire h_u_cla32_and7141_y0;
  wire h_u_cla32_and7142_y0;
  wire h_u_cla32_and7143_y0;
  wire h_u_cla32_and7144_y0;
  wire h_u_cla32_and7145_y0;
  wire h_u_cla32_and7146_y0;
  wire h_u_cla32_and7147_y0;
  wire h_u_cla32_and7148_y0;
  wire h_u_cla32_and7149_y0;
  wire h_u_cla32_and7150_y0;
  wire h_u_cla32_and7151_y0;
  wire h_u_cla32_and7152_y0;
  wire h_u_cla32_and7153_y0;
  wire h_u_cla32_and7154_y0;
  wire h_u_cla32_and7155_y0;
  wire h_u_cla32_and7156_y0;
  wire h_u_cla32_and7157_y0;
  wire h_u_cla32_and7158_y0;
  wire h_u_cla32_and7159_y0;
  wire h_u_cla32_and7160_y0;
  wire h_u_cla32_and7161_y0;
  wire h_u_cla32_and7162_y0;
  wire h_u_cla32_and7163_y0;
  wire h_u_cla32_and7164_y0;
  wire h_u_cla32_and7165_y0;
  wire h_u_cla32_and7166_y0;
  wire h_u_cla32_and7167_y0;
  wire h_u_cla32_and7168_y0;
  wire h_u_cla32_and7169_y0;
  wire h_u_cla32_and7170_y0;
  wire h_u_cla32_and7171_y0;
  wire h_u_cla32_and7172_y0;
  wire h_u_cla32_and7173_y0;
  wire h_u_cla32_and7174_y0;
  wire h_u_cla32_and7175_y0;
  wire h_u_cla32_and7176_y0;
  wire h_u_cla32_and7177_y0;
  wire h_u_cla32_and7178_y0;
  wire h_u_cla32_and7179_y0;
  wire h_u_cla32_and7180_y0;
  wire h_u_cla32_and7181_y0;
  wire h_u_cla32_and7182_y0;
  wire h_u_cla32_and7183_y0;
  wire h_u_cla32_and7184_y0;
  wire h_u_cla32_and7185_y0;
  wire h_u_cla32_and7186_y0;
  wire h_u_cla32_and7187_y0;
  wire h_u_cla32_and7188_y0;
  wire h_u_cla32_and7189_y0;
  wire h_u_cla32_and7190_y0;
  wire h_u_cla32_and7191_y0;
  wire h_u_cla32_and7192_y0;
  wire h_u_cla32_and7193_y0;
  wire h_u_cla32_and7194_y0;
  wire h_u_cla32_and7195_y0;
  wire h_u_cla32_and7196_y0;
  wire h_u_cla32_and7197_y0;
  wire h_u_cla32_and7198_y0;
  wire h_u_cla32_and7199_y0;
  wire h_u_cla32_and7200_y0;
  wire h_u_cla32_and7201_y0;
  wire h_u_cla32_and7202_y0;
  wire h_u_cla32_and7203_y0;
  wire h_u_cla32_and7204_y0;
  wire h_u_cla32_and7205_y0;
  wire h_u_cla32_and7206_y0;
  wire h_u_cla32_and7207_y0;
  wire h_u_cla32_and7208_y0;
  wire h_u_cla32_and7209_y0;
  wire h_u_cla32_and7210_y0;
  wire h_u_cla32_and7211_y0;
  wire h_u_cla32_and7212_y0;
  wire h_u_cla32_and7213_y0;
  wire h_u_cla32_and7214_y0;
  wire h_u_cla32_and7215_y0;
  wire h_u_cla32_and7216_y0;
  wire h_u_cla32_and7217_y0;
  wire h_u_cla32_and7218_y0;
  wire h_u_cla32_and7219_y0;
  wire h_u_cla32_and7220_y0;
  wire h_u_cla32_and7221_y0;
  wire h_u_cla32_and7222_y0;
  wire h_u_cla32_and7223_y0;
  wire h_u_cla32_and7224_y0;
  wire h_u_cla32_and7225_y0;
  wire h_u_cla32_and7226_y0;
  wire h_u_cla32_and7227_y0;
  wire h_u_cla32_and7228_y0;
  wire h_u_cla32_and7229_y0;
  wire h_u_cla32_and7230_y0;
  wire h_u_cla32_and7231_y0;
  wire h_u_cla32_and7232_y0;
  wire h_u_cla32_and7233_y0;
  wire h_u_cla32_and7234_y0;
  wire h_u_cla32_and7235_y0;
  wire h_u_cla32_and7236_y0;
  wire h_u_cla32_and7237_y0;
  wire h_u_cla32_and7238_y0;
  wire h_u_cla32_and7239_y0;
  wire h_u_cla32_and7240_y0;
  wire h_u_cla32_and7241_y0;
  wire h_u_cla32_and7242_y0;
  wire h_u_cla32_and7243_y0;
  wire h_u_cla32_and7244_y0;
  wire h_u_cla32_and7245_y0;
  wire h_u_cla32_and7246_y0;
  wire h_u_cla32_and7247_y0;
  wire h_u_cla32_and7248_y0;
  wire h_u_cla32_and7249_y0;
  wire h_u_cla32_and7250_y0;
  wire h_u_cla32_and7251_y0;
  wire h_u_cla32_and7252_y0;
  wire h_u_cla32_and7253_y0;
  wire h_u_cla32_and7254_y0;
  wire h_u_cla32_and7255_y0;
  wire h_u_cla32_and7256_y0;
  wire h_u_cla32_and7257_y0;
  wire h_u_cla32_and7258_y0;
  wire h_u_cla32_and7259_y0;
  wire h_u_cla32_and7260_y0;
  wire h_u_cla32_and7261_y0;
  wire h_u_cla32_and7262_y0;
  wire h_u_cla32_and7263_y0;
  wire h_u_cla32_and7264_y0;
  wire h_u_cla32_and7265_y0;
  wire h_u_cla32_and7266_y0;
  wire h_u_cla32_and7267_y0;
  wire h_u_cla32_and7268_y0;
  wire h_u_cla32_and7269_y0;
  wire h_u_cla32_and7270_y0;
  wire h_u_cla32_and7271_y0;
  wire h_u_cla32_and7272_y0;
  wire h_u_cla32_and7273_y0;
  wire h_u_cla32_and7274_y0;
  wire h_u_cla32_and7275_y0;
  wire h_u_cla32_and7276_y0;
  wire h_u_cla32_and7277_y0;
  wire h_u_cla32_and7278_y0;
  wire h_u_cla32_and7279_y0;
  wire h_u_cla32_and7280_y0;
  wire h_u_cla32_and7281_y0;
  wire h_u_cla32_and7282_y0;
  wire h_u_cla32_and7283_y0;
  wire h_u_cla32_and7284_y0;
  wire h_u_cla32_and7285_y0;
  wire h_u_cla32_and7286_y0;
  wire h_u_cla32_and7287_y0;
  wire h_u_cla32_and7288_y0;
  wire h_u_cla32_and7289_y0;
  wire h_u_cla32_and7290_y0;
  wire h_u_cla32_and7291_y0;
  wire h_u_cla32_and7292_y0;
  wire h_u_cla32_and7293_y0;
  wire h_u_cla32_and7294_y0;
  wire h_u_cla32_and7295_y0;
  wire h_u_cla32_and7296_y0;
  wire h_u_cla32_and7297_y0;
  wire h_u_cla32_and7298_y0;
  wire h_u_cla32_and7299_y0;
  wire h_u_cla32_and7300_y0;
  wire h_u_cla32_and7301_y0;
  wire h_u_cla32_and7302_y0;
  wire h_u_cla32_and7303_y0;
  wire h_u_cla32_and7304_y0;
  wire h_u_cla32_and7305_y0;
  wire h_u_cla32_and7306_y0;
  wire h_u_cla32_and7307_y0;
  wire h_u_cla32_and7308_y0;
  wire h_u_cla32_and7309_y0;
  wire h_u_cla32_and7310_y0;
  wire h_u_cla32_and7311_y0;
  wire h_u_cla32_and7312_y0;
  wire h_u_cla32_and7313_y0;
  wire h_u_cla32_and7314_y0;
  wire h_u_cla32_and7315_y0;
  wire h_u_cla32_and7316_y0;
  wire h_u_cla32_and7317_y0;
  wire h_u_cla32_and7318_y0;
  wire h_u_cla32_and7319_y0;
  wire h_u_cla32_and7320_y0;
  wire h_u_cla32_and7321_y0;
  wire h_u_cla32_and7322_y0;
  wire h_u_cla32_and7323_y0;
  wire h_u_cla32_and7324_y0;
  wire h_u_cla32_and7325_y0;
  wire h_u_cla32_and7326_y0;
  wire h_u_cla32_and7327_y0;
  wire h_u_cla32_and7328_y0;
  wire h_u_cla32_and7329_y0;
  wire h_u_cla32_and7330_y0;
  wire h_u_cla32_and7331_y0;
  wire h_u_cla32_and7332_y0;
  wire h_u_cla32_and7333_y0;
  wire h_u_cla32_and7334_y0;
  wire h_u_cla32_and7335_y0;
  wire h_u_cla32_and7336_y0;
  wire h_u_cla32_and7337_y0;
  wire h_u_cla32_and7338_y0;
  wire h_u_cla32_and7339_y0;
  wire h_u_cla32_and7340_y0;
  wire h_u_cla32_and7341_y0;
  wire h_u_cla32_and7342_y0;
  wire h_u_cla32_and7343_y0;
  wire h_u_cla32_and7344_y0;
  wire h_u_cla32_and7345_y0;
  wire h_u_cla32_and7346_y0;
  wire h_u_cla32_and7347_y0;
  wire h_u_cla32_and7348_y0;
  wire h_u_cla32_and7349_y0;
  wire h_u_cla32_and7350_y0;
  wire h_u_cla32_and7351_y0;
  wire h_u_cla32_and7352_y0;
  wire h_u_cla32_and7353_y0;
  wire h_u_cla32_and7354_y0;
  wire h_u_cla32_and7355_y0;
  wire h_u_cla32_and7356_y0;
  wire h_u_cla32_and7357_y0;
  wire h_u_cla32_and7358_y0;
  wire h_u_cla32_and7359_y0;
  wire h_u_cla32_and7360_y0;
  wire h_u_cla32_and7361_y0;
  wire h_u_cla32_and7362_y0;
  wire h_u_cla32_and7363_y0;
  wire h_u_cla32_and7364_y0;
  wire h_u_cla32_and7365_y0;
  wire h_u_cla32_and7366_y0;
  wire h_u_cla32_and7367_y0;
  wire h_u_cla32_and7368_y0;
  wire h_u_cla32_and7369_y0;
  wire h_u_cla32_and7370_y0;
  wire h_u_cla32_and7371_y0;
  wire h_u_cla32_and7372_y0;
  wire h_u_cla32_and7373_y0;
  wire h_u_cla32_and7374_y0;
  wire h_u_cla32_and7375_y0;
  wire h_u_cla32_and7376_y0;
  wire h_u_cla32_and7377_y0;
  wire h_u_cla32_and7378_y0;
  wire h_u_cla32_and7379_y0;
  wire h_u_cla32_and7380_y0;
  wire h_u_cla32_and7381_y0;
  wire h_u_cla32_and7382_y0;
  wire h_u_cla32_and7383_y0;
  wire h_u_cla32_and7384_y0;
  wire h_u_cla32_and7385_y0;
  wire h_u_cla32_and7386_y0;
  wire h_u_cla32_and7387_y0;
  wire h_u_cla32_and7388_y0;
  wire h_u_cla32_and7389_y0;
  wire h_u_cla32_and7390_y0;
  wire h_u_cla32_and7391_y0;
  wire h_u_cla32_and7392_y0;
  wire h_u_cla32_and7393_y0;
  wire h_u_cla32_and7394_y0;
  wire h_u_cla32_and7395_y0;
  wire h_u_cla32_and7396_y0;
  wire h_u_cla32_and7397_y0;
  wire h_u_cla32_and7398_y0;
  wire h_u_cla32_and7399_y0;
  wire h_u_cla32_and7400_y0;
  wire h_u_cla32_and7401_y0;
  wire h_u_cla32_and7402_y0;
  wire h_u_cla32_and7403_y0;
  wire h_u_cla32_and7404_y0;
  wire h_u_cla32_and7405_y0;
  wire h_u_cla32_and7406_y0;
  wire h_u_cla32_and7407_y0;
  wire h_u_cla32_and7408_y0;
  wire h_u_cla32_and7409_y0;
  wire h_u_cla32_and7410_y0;
  wire h_u_cla32_and7411_y0;
  wire h_u_cla32_and7412_y0;
  wire h_u_cla32_and7413_y0;
  wire h_u_cla32_and7414_y0;
  wire h_u_cla32_and7415_y0;
  wire h_u_cla32_and7416_y0;
  wire h_u_cla32_and7417_y0;
  wire h_u_cla32_and7418_y0;
  wire h_u_cla32_and7419_y0;
  wire h_u_cla32_and7420_y0;
  wire h_u_cla32_and7421_y0;
  wire h_u_cla32_and7422_y0;
  wire h_u_cla32_and7423_y0;
  wire h_u_cla32_and7424_y0;
  wire h_u_cla32_and7425_y0;
  wire h_u_cla32_and7426_y0;
  wire h_u_cla32_and7427_y0;
  wire h_u_cla32_and7428_y0;
  wire h_u_cla32_and7429_y0;
  wire h_u_cla32_and7430_y0;
  wire h_u_cla32_and7431_y0;
  wire h_u_cla32_and7432_y0;
  wire h_u_cla32_and7433_y0;
  wire h_u_cla32_and7434_y0;
  wire h_u_cla32_and7435_y0;
  wire h_u_cla32_and7436_y0;
  wire h_u_cla32_and7437_y0;
  wire h_u_cla32_and7438_y0;
  wire h_u_cla32_and7439_y0;
  wire h_u_cla32_and7440_y0;
  wire h_u_cla32_and7441_y0;
  wire h_u_cla32_and7442_y0;
  wire h_u_cla32_and7443_y0;
  wire h_u_cla32_and7444_y0;
  wire h_u_cla32_and7445_y0;
  wire h_u_cla32_and7446_y0;
  wire h_u_cla32_and7447_y0;
  wire h_u_cla32_and7448_y0;
  wire h_u_cla32_and7449_y0;
  wire h_u_cla32_and7450_y0;
  wire h_u_cla32_and7451_y0;
  wire h_u_cla32_and7452_y0;
  wire h_u_cla32_and7453_y0;
  wire h_u_cla32_and7454_y0;
  wire h_u_cla32_and7455_y0;
  wire h_u_cla32_and7456_y0;
  wire h_u_cla32_and7457_y0;
  wire h_u_cla32_and7458_y0;
  wire h_u_cla32_and7459_y0;
  wire h_u_cla32_and7460_y0;
  wire h_u_cla32_and7461_y0;
  wire h_u_cla32_and7462_y0;
  wire h_u_cla32_and7463_y0;
  wire h_u_cla32_and7464_y0;
  wire h_u_cla32_and7465_y0;
  wire h_u_cla32_and7466_y0;
  wire h_u_cla32_and7467_y0;
  wire h_u_cla32_and7468_y0;
  wire h_u_cla32_and7469_y0;
  wire h_u_cla32_and7470_y0;
  wire h_u_cla32_and7471_y0;
  wire h_u_cla32_and7472_y0;
  wire h_u_cla32_and7473_y0;
  wire h_u_cla32_and7474_y0;
  wire h_u_cla32_and7475_y0;
  wire h_u_cla32_and7476_y0;
  wire h_u_cla32_and7477_y0;
  wire h_u_cla32_and7478_y0;
  wire h_u_cla32_and7479_y0;
  wire h_u_cla32_and7480_y0;
  wire h_u_cla32_and7481_y0;
  wire h_u_cla32_and7482_y0;
  wire h_u_cla32_and7483_y0;
  wire h_u_cla32_and7484_y0;
  wire h_u_cla32_and7485_y0;
  wire h_u_cla32_and7486_y0;
  wire h_u_cla32_and7487_y0;
  wire h_u_cla32_and7488_y0;
  wire h_u_cla32_and7489_y0;
  wire h_u_cla32_and7490_y0;
  wire h_u_cla32_and7491_y0;
  wire h_u_cla32_and7492_y0;
  wire h_u_cla32_and7493_y0;
  wire h_u_cla32_and7494_y0;
  wire h_u_cla32_and7495_y0;
  wire h_u_cla32_and7496_y0;
  wire h_u_cla32_and7497_y0;
  wire h_u_cla32_and7498_y0;
  wire h_u_cla32_and7499_y0;
  wire h_u_cla32_and7500_y0;
  wire h_u_cla32_and7501_y0;
  wire h_u_cla32_and7502_y0;
  wire h_u_cla32_and7503_y0;
  wire h_u_cla32_and7504_y0;
  wire h_u_cla32_and7505_y0;
  wire h_u_cla32_and7506_y0;
  wire h_u_cla32_and7507_y0;
  wire h_u_cla32_and7508_y0;
  wire h_u_cla32_and7509_y0;
  wire h_u_cla32_and7510_y0;
  wire h_u_cla32_and7511_y0;
  wire h_u_cla32_and7512_y0;
  wire h_u_cla32_and7513_y0;
  wire h_u_cla32_and7514_y0;
  wire h_u_cla32_and7515_y0;
  wire h_u_cla32_and7516_y0;
  wire h_u_cla32_and7517_y0;
  wire h_u_cla32_and7518_y0;
  wire h_u_cla32_and7519_y0;
  wire h_u_cla32_and7520_y0;
  wire h_u_cla32_and7521_y0;
  wire h_u_cla32_and7522_y0;
  wire h_u_cla32_and7523_y0;
  wire h_u_cla32_and7524_y0;
  wire h_u_cla32_and7525_y0;
  wire h_u_cla32_and7526_y0;
  wire h_u_cla32_and7527_y0;
  wire h_u_cla32_and7528_y0;
  wire h_u_cla32_and7529_y0;
  wire h_u_cla32_and7530_y0;
  wire h_u_cla32_and7531_y0;
  wire h_u_cla32_and7532_y0;
  wire h_u_cla32_and7533_y0;
  wire h_u_cla32_and7534_y0;
  wire h_u_cla32_and7535_y0;
  wire h_u_cla32_and7536_y0;
  wire h_u_cla32_and7537_y0;
  wire h_u_cla32_and7538_y0;
  wire h_u_cla32_and7539_y0;
  wire h_u_cla32_and7540_y0;
  wire h_u_cla32_and7541_y0;
  wire h_u_cla32_and7542_y0;
  wire h_u_cla32_and7543_y0;
  wire h_u_cla32_and7544_y0;
  wire h_u_cla32_and7545_y0;
  wire h_u_cla32_and7546_y0;
  wire h_u_cla32_and7547_y0;
  wire h_u_cla32_and7548_y0;
  wire h_u_cla32_and7549_y0;
  wire h_u_cla32_and7550_y0;
  wire h_u_cla32_and7551_y0;
  wire h_u_cla32_and7552_y0;
  wire h_u_cla32_and7553_y0;
  wire h_u_cla32_and7554_y0;
  wire h_u_cla32_and7555_y0;
  wire h_u_cla32_and7556_y0;
  wire h_u_cla32_and7557_y0;
  wire h_u_cla32_and7558_y0;
  wire h_u_cla32_and7559_y0;
  wire h_u_cla32_and7560_y0;
  wire h_u_cla32_and7561_y0;
  wire h_u_cla32_and7562_y0;
  wire h_u_cla32_and7563_y0;
  wire h_u_cla32_and7564_y0;
  wire h_u_cla32_and7565_y0;
  wire h_u_cla32_and7566_y0;
  wire h_u_cla32_and7567_y0;
  wire h_u_cla32_and7568_y0;
  wire h_u_cla32_and7569_y0;
  wire h_u_cla32_and7570_y0;
  wire h_u_cla32_and7571_y0;
  wire h_u_cla32_and7572_y0;
  wire h_u_cla32_and7573_y0;
  wire h_u_cla32_and7574_y0;
  wire h_u_cla32_and7575_y0;
  wire h_u_cla32_and7576_y0;
  wire h_u_cla32_and7577_y0;
  wire h_u_cla32_and7578_y0;
  wire h_u_cla32_and7579_y0;
  wire h_u_cla32_and7580_y0;
  wire h_u_cla32_and7581_y0;
  wire h_u_cla32_and7582_y0;
  wire h_u_cla32_and7583_y0;
  wire h_u_cla32_and7584_y0;
  wire h_u_cla32_and7585_y0;
  wire h_u_cla32_and7586_y0;
  wire h_u_cla32_and7587_y0;
  wire h_u_cla32_and7588_y0;
  wire h_u_cla32_and7589_y0;
  wire h_u_cla32_and7590_y0;
  wire h_u_cla32_and7591_y0;
  wire h_u_cla32_and7592_y0;
  wire h_u_cla32_and7593_y0;
  wire h_u_cla32_and7594_y0;
  wire h_u_cla32_and7595_y0;
  wire h_u_cla32_and7596_y0;
  wire h_u_cla32_and7597_y0;
  wire h_u_cla32_and7598_y0;
  wire h_u_cla32_and7599_y0;
  wire h_u_cla32_and7600_y0;
  wire h_u_cla32_and7601_y0;
  wire h_u_cla32_and7602_y0;
  wire h_u_cla32_and7603_y0;
  wire h_u_cla32_and7604_y0;
  wire h_u_cla32_and7605_y0;
  wire h_u_cla32_and7606_y0;
  wire h_u_cla32_and7607_y0;
  wire h_u_cla32_and7608_y0;
  wire h_u_cla32_and7609_y0;
  wire h_u_cla32_and7610_y0;
  wire h_u_cla32_and7611_y0;
  wire h_u_cla32_and7612_y0;
  wire h_u_cla32_and7613_y0;
  wire h_u_cla32_and7614_y0;
  wire h_u_cla32_and7615_y0;
  wire h_u_cla32_and7616_y0;
  wire h_u_cla32_and7617_y0;
  wire h_u_cla32_and7618_y0;
  wire h_u_cla32_and7619_y0;
  wire h_u_cla32_and7620_y0;
  wire h_u_cla32_and7621_y0;
  wire h_u_cla32_and7622_y0;
  wire h_u_cla32_and7623_y0;
  wire h_u_cla32_and7624_y0;
  wire h_u_cla32_and7625_y0;
  wire h_u_cla32_and7626_y0;
  wire h_u_cla32_and7627_y0;
  wire h_u_cla32_and7628_y0;
  wire h_u_cla32_and7629_y0;
  wire h_u_cla32_and7630_y0;
  wire h_u_cla32_and7631_y0;
  wire h_u_cla32_and7632_y0;
  wire h_u_cla32_and7633_y0;
  wire h_u_cla32_and7634_y0;
  wire h_u_cla32_and7635_y0;
  wire h_u_cla32_and7636_y0;
  wire h_u_cla32_and7637_y0;
  wire h_u_cla32_and7638_y0;
  wire h_u_cla32_and7639_y0;
  wire h_u_cla32_and7640_y0;
  wire h_u_cla32_and7641_y0;
  wire h_u_cla32_and7642_y0;
  wire h_u_cla32_and7643_y0;
  wire h_u_cla32_and7644_y0;
  wire h_u_cla32_and7645_y0;
  wire h_u_cla32_and7646_y0;
  wire h_u_cla32_and7647_y0;
  wire h_u_cla32_and7648_y0;
  wire h_u_cla32_and7649_y0;
  wire h_u_cla32_and7650_y0;
  wire h_u_cla32_and7651_y0;
  wire h_u_cla32_and7652_y0;
  wire h_u_cla32_and7653_y0;
  wire h_u_cla32_and7654_y0;
  wire h_u_cla32_and7655_y0;
  wire h_u_cla32_and7656_y0;
  wire h_u_cla32_and7657_y0;
  wire h_u_cla32_and7658_y0;
  wire h_u_cla32_and7659_y0;
  wire h_u_cla32_and7660_y0;
  wire h_u_cla32_and7661_y0;
  wire h_u_cla32_and7662_y0;
  wire h_u_cla32_and7663_y0;
  wire h_u_cla32_and7664_y0;
  wire h_u_cla32_and7665_y0;
  wire h_u_cla32_and7666_y0;
  wire h_u_cla32_and7667_y0;
  wire h_u_cla32_and7668_y0;
  wire h_u_cla32_and7669_y0;
  wire h_u_cla32_and7670_y0;
  wire h_u_cla32_and7671_y0;
  wire h_u_cla32_and7672_y0;
  wire h_u_cla32_and7673_y0;
  wire h_u_cla32_and7674_y0;
  wire h_u_cla32_and7675_y0;
  wire h_u_cla32_and7676_y0;
  wire h_u_cla32_and7677_y0;
  wire h_u_cla32_and7678_y0;
  wire h_u_cla32_and7679_y0;
  wire h_u_cla32_and7680_y0;
  wire h_u_cla32_and7681_y0;
  wire h_u_cla32_and7682_y0;
  wire h_u_cla32_and7683_y0;
  wire h_u_cla32_and7684_y0;
  wire h_u_cla32_and7685_y0;
  wire h_u_cla32_and7686_y0;
  wire h_u_cla32_and7687_y0;
  wire h_u_cla32_and7688_y0;
  wire h_u_cla32_and7689_y0;
  wire h_u_cla32_and7690_y0;
  wire h_u_cla32_and7691_y0;
  wire h_u_cla32_and7692_y0;
  wire h_u_cla32_and7693_y0;
  wire h_u_cla32_and7694_y0;
  wire h_u_cla32_and7695_y0;
  wire h_u_cla32_and7696_y0;
  wire h_u_cla32_and7697_y0;
  wire h_u_cla32_and7698_y0;
  wire h_u_cla32_and7699_y0;
  wire h_u_cla32_and7700_y0;
  wire h_u_cla32_and7701_y0;
  wire h_u_cla32_and7702_y0;
  wire h_u_cla32_and7703_y0;
  wire h_u_cla32_and7704_y0;
  wire h_u_cla32_and7705_y0;
  wire h_u_cla32_and7706_y0;
  wire h_u_cla32_and7707_y0;
  wire h_u_cla32_and7708_y0;
  wire h_u_cla32_and7709_y0;
  wire h_u_cla32_and7710_y0;
  wire h_u_cla32_and7711_y0;
  wire h_u_cla32_and7712_y0;
  wire h_u_cla32_and7713_y0;
  wire h_u_cla32_or378_y0;
  wire h_u_cla32_or379_y0;
  wire h_u_cla32_or380_y0;
  wire h_u_cla32_or381_y0;
  wire h_u_cla32_or382_y0;
  wire h_u_cla32_or383_y0;
  wire h_u_cla32_or384_y0;
  wire h_u_cla32_or385_y0;
  wire h_u_cla32_or386_y0;
  wire h_u_cla32_or387_y0;
  wire h_u_cla32_or388_y0;
  wire h_u_cla32_or389_y0;
  wire h_u_cla32_or390_y0;
  wire h_u_cla32_or391_y0;
  wire h_u_cla32_or392_y0;
  wire h_u_cla32_or393_y0;
  wire h_u_cla32_or394_y0;
  wire h_u_cla32_or395_y0;
  wire h_u_cla32_or396_y0;
  wire h_u_cla32_or397_y0;
  wire h_u_cla32_or398_y0;
  wire h_u_cla32_or399_y0;
  wire h_u_cla32_or400_y0;
  wire h_u_cla32_or401_y0;
  wire h_u_cla32_or402_y0;
  wire h_u_cla32_or403_y0;
  wire h_u_cla32_or404_y0;
  wire h_u_cla32_or405_y0;
  wire h_u_cla32_pg_logic28_y0;
  wire h_u_cla32_pg_logic28_y1;
  wire h_u_cla32_pg_logic28_y2;
  wire h_u_cla32_xor28_y0;
  wire h_u_cla32_and7714_y0;
  wire h_u_cla32_and7715_y0;
  wire h_u_cla32_and7716_y0;
  wire h_u_cla32_and7717_y0;
  wire h_u_cla32_and7718_y0;
  wire h_u_cla32_and7719_y0;
  wire h_u_cla32_and7720_y0;
  wire h_u_cla32_and7721_y0;
  wire h_u_cla32_and7722_y0;
  wire h_u_cla32_and7723_y0;
  wire h_u_cla32_and7724_y0;
  wire h_u_cla32_and7725_y0;
  wire h_u_cla32_and7726_y0;
  wire h_u_cla32_and7727_y0;
  wire h_u_cla32_and7728_y0;
  wire h_u_cla32_and7729_y0;
  wire h_u_cla32_and7730_y0;
  wire h_u_cla32_and7731_y0;
  wire h_u_cla32_and7732_y0;
  wire h_u_cla32_and7733_y0;
  wire h_u_cla32_and7734_y0;
  wire h_u_cla32_and7735_y0;
  wire h_u_cla32_and7736_y0;
  wire h_u_cla32_and7737_y0;
  wire h_u_cla32_and7738_y0;
  wire h_u_cla32_and7739_y0;
  wire h_u_cla32_and7740_y0;
  wire h_u_cla32_and7741_y0;
  wire h_u_cla32_and7742_y0;
  wire h_u_cla32_and7743_y0;
  wire h_u_cla32_and7744_y0;
  wire h_u_cla32_and7745_y0;
  wire h_u_cla32_and7746_y0;
  wire h_u_cla32_and7747_y0;
  wire h_u_cla32_and7748_y0;
  wire h_u_cla32_and7749_y0;
  wire h_u_cla32_and7750_y0;
  wire h_u_cla32_and7751_y0;
  wire h_u_cla32_and7752_y0;
  wire h_u_cla32_and7753_y0;
  wire h_u_cla32_and7754_y0;
  wire h_u_cla32_and7755_y0;
  wire h_u_cla32_and7756_y0;
  wire h_u_cla32_and7757_y0;
  wire h_u_cla32_and7758_y0;
  wire h_u_cla32_and7759_y0;
  wire h_u_cla32_and7760_y0;
  wire h_u_cla32_and7761_y0;
  wire h_u_cla32_and7762_y0;
  wire h_u_cla32_and7763_y0;
  wire h_u_cla32_and7764_y0;
  wire h_u_cla32_and7765_y0;
  wire h_u_cla32_and7766_y0;
  wire h_u_cla32_and7767_y0;
  wire h_u_cla32_and7768_y0;
  wire h_u_cla32_and7769_y0;
  wire h_u_cla32_and7770_y0;
  wire h_u_cla32_and7771_y0;
  wire h_u_cla32_and7772_y0;
  wire h_u_cla32_and7773_y0;
  wire h_u_cla32_and7774_y0;
  wire h_u_cla32_and7775_y0;
  wire h_u_cla32_and7776_y0;
  wire h_u_cla32_and7777_y0;
  wire h_u_cla32_and7778_y0;
  wire h_u_cla32_and7779_y0;
  wire h_u_cla32_and7780_y0;
  wire h_u_cla32_and7781_y0;
  wire h_u_cla32_and7782_y0;
  wire h_u_cla32_and7783_y0;
  wire h_u_cla32_and7784_y0;
  wire h_u_cla32_and7785_y0;
  wire h_u_cla32_and7786_y0;
  wire h_u_cla32_and7787_y0;
  wire h_u_cla32_and7788_y0;
  wire h_u_cla32_and7789_y0;
  wire h_u_cla32_and7790_y0;
  wire h_u_cla32_and7791_y0;
  wire h_u_cla32_and7792_y0;
  wire h_u_cla32_and7793_y0;
  wire h_u_cla32_and7794_y0;
  wire h_u_cla32_and7795_y0;
  wire h_u_cla32_and7796_y0;
  wire h_u_cla32_and7797_y0;
  wire h_u_cla32_and7798_y0;
  wire h_u_cla32_and7799_y0;
  wire h_u_cla32_and7800_y0;
  wire h_u_cla32_and7801_y0;
  wire h_u_cla32_and7802_y0;
  wire h_u_cla32_and7803_y0;
  wire h_u_cla32_and7804_y0;
  wire h_u_cla32_and7805_y0;
  wire h_u_cla32_and7806_y0;
  wire h_u_cla32_and7807_y0;
  wire h_u_cla32_and7808_y0;
  wire h_u_cla32_and7809_y0;
  wire h_u_cla32_and7810_y0;
  wire h_u_cla32_and7811_y0;
  wire h_u_cla32_and7812_y0;
  wire h_u_cla32_and7813_y0;
  wire h_u_cla32_and7814_y0;
  wire h_u_cla32_and7815_y0;
  wire h_u_cla32_and7816_y0;
  wire h_u_cla32_and7817_y0;
  wire h_u_cla32_and7818_y0;
  wire h_u_cla32_and7819_y0;
  wire h_u_cla32_and7820_y0;
  wire h_u_cla32_and7821_y0;
  wire h_u_cla32_and7822_y0;
  wire h_u_cla32_and7823_y0;
  wire h_u_cla32_and7824_y0;
  wire h_u_cla32_and7825_y0;
  wire h_u_cla32_and7826_y0;
  wire h_u_cla32_and7827_y0;
  wire h_u_cla32_and7828_y0;
  wire h_u_cla32_and7829_y0;
  wire h_u_cla32_and7830_y0;
  wire h_u_cla32_and7831_y0;
  wire h_u_cla32_and7832_y0;
  wire h_u_cla32_and7833_y0;
  wire h_u_cla32_and7834_y0;
  wire h_u_cla32_and7835_y0;
  wire h_u_cla32_and7836_y0;
  wire h_u_cla32_and7837_y0;
  wire h_u_cla32_and7838_y0;
  wire h_u_cla32_and7839_y0;
  wire h_u_cla32_and7840_y0;
  wire h_u_cla32_and7841_y0;
  wire h_u_cla32_and7842_y0;
  wire h_u_cla32_and7843_y0;
  wire h_u_cla32_and7844_y0;
  wire h_u_cla32_and7845_y0;
  wire h_u_cla32_and7846_y0;
  wire h_u_cla32_and7847_y0;
  wire h_u_cla32_and7848_y0;
  wire h_u_cla32_and7849_y0;
  wire h_u_cla32_and7850_y0;
  wire h_u_cla32_and7851_y0;
  wire h_u_cla32_and7852_y0;
  wire h_u_cla32_and7853_y0;
  wire h_u_cla32_and7854_y0;
  wire h_u_cla32_and7855_y0;
  wire h_u_cla32_and7856_y0;
  wire h_u_cla32_and7857_y0;
  wire h_u_cla32_and7858_y0;
  wire h_u_cla32_and7859_y0;
  wire h_u_cla32_and7860_y0;
  wire h_u_cla32_and7861_y0;
  wire h_u_cla32_and7862_y0;
  wire h_u_cla32_and7863_y0;
  wire h_u_cla32_and7864_y0;
  wire h_u_cla32_and7865_y0;
  wire h_u_cla32_and7866_y0;
  wire h_u_cla32_and7867_y0;
  wire h_u_cla32_and7868_y0;
  wire h_u_cla32_and7869_y0;
  wire h_u_cla32_and7870_y0;
  wire h_u_cla32_and7871_y0;
  wire h_u_cla32_and7872_y0;
  wire h_u_cla32_and7873_y0;
  wire h_u_cla32_and7874_y0;
  wire h_u_cla32_and7875_y0;
  wire h_u_cla32_and7876_y0;
  wire h_u_cla32_and7877_y0;
  wire h_u_cla32_and7878_y0;
  wire h_u_cla32_and7879_y0;
  wire h_u_cla32_and7880_y0;
  wire h_u_cla32_and7881_y0;
  wire h_u_cla32_and7882_y0;
  wire h_u_cla32_and7883_y0;
  wire h_u_cla32_and7884_y0;
  wire h_u_cla32_and7885_y0;
  wire h_u_cla32_and7886_y0;
  wire h_u_cla32_and7887_y0;
  wire h_u_cla32_and7888_y0;
  wire h_u_cla32_and7889_y0;
  wire h_u_cla32_and7890_y0;
  wire h_u_cla32_and7891_y0;
  wire h_u_cla32_and7892_y0;
  wire h_u_cla32_and7893_y0;
  wire h_u_cla32_and7894_y0;
  wire h_u_cla32_and7895_y0;
  wire h_u_cla32_and7896_y0;
  wire h_u_cla32_and7897_y0;
  wire h_u_cla32_and7898_y0;
  wire h_u_cla32_and7899_y0;
  wire h_u_cla32_and7900_y0;
  wire h_u_cla32_and7901_y0;
  wire h_u_cla32_and7902_y0;
  wire h_u_cla32_and7903_y0;
  wire h_u_cla32_and7904_y0;
  wire h_u_cla32_and7905_y0;
  wire h_u_cla32_and7906_y0;
  wire h_u_cla32_and7907_y0;
  wire h_u_cla32_and7908_y0;
  wire h_u_cla32_and7909_y0;
  wire h_u_cla32_and7910_y0;
  wire h_u_cla32_and7911_y0;
  wire h_u_cla32_and7912_y0;
  wire h_u_cla32_and7913_y0;
  wire h_u_cla32_and7914_y0;
  wire h_u_cla32_and7915_y0;
  wire h_u_cla32_and7916_y0;
  wire h_u_cla32_and7917_y0;
  wire h_u_cla32_and7918_y0;
  wire h_u_cla32_and7919_y0;
  wire h_u_cla32_and7920_y0;
  wire h_u_cla32_and7921_y0;
  wire h_u_cla32_and7922_y0;
  wire h_u_cla32_and7923_y0;
  wire h_u_cla32_and7924_y0;
  wire h_u_cla32_and7925_y0;
  wire h_u_cla32_and7926_y0;
  wire h_u_cla32_and7927_y0;
  wire h_u_cla32_and7928_y0;
  wire h_u_cla32_and7929_y0;
  wire h_u_cla32_and7930_y0;
  wire h_u_cla32_and7931_y0;
  wire h_u_cla32_and7932_y0;
  wire h_u_cla32_and7933_y0;
  wire h_u_cla32_and7934_y0;
  wire h_u_cla32_and7935_y0;
  wire h_u_cla32_and7936_y0;
  wire h_u_cla32_and7937_y0;
  wire h_u_cla32_and7938_y0;
  wire h_u_cla32_and7939_y0;
  wire h_u_cla32_and7940_y0;
  wire h_u_cla32_and7941_y0;
  wire h_u_cla32_and7942_y0;
  wire h_u_cla32_and7943_y0;
  wire h_u_cla32_and7944_y0;
  wire h_u_cla32_and7945_y0;
  wire h_u_cla32_and7946_y0;
  wire h_u_cla32_and7947_y0;
  wire h_u_cla32_and7948_y0;
  wire h_u_cla32_and7949_y0;
  wire h_u_cla32_and7950_y0;
  wire h_u_cla32_and7951_y0;
  wire h_u_cla32_and7952_y0;
  wire h_u_cla32_and7953_y0;
  wire h_u_cla32_and7954_y0;
  wire h_u_cla32_and7955_y0;
  wire h_u_cla32_and7956_y0;
  wire h_u_cla32_and7957_y0;
  wire h_u_cla32_and7958_y0;
  wire h_u_cla32_and7959_y0;
  wire h_u_cla32_and7960_y0;
  wire h_u_cla32_and7961_y0;
  wire h_u_cla32_and7962_y0;
  wire h_u_cla32_and7963_y0;
  wire h_u_cla32_and7964_y0;
  wire h_u_cla32_and7965_y0;
  wire h_u_cla32_and7966_y0;
  wire h_u_cla32_and7967_y0;
  wire h_u_cla32_and7968_y0;
  wire h_u_cla32_and7969_y0;
  wire h_u_cla32_and7970_y0;
  wire h_u_cla32_and7971_y0;
  wire h_u_cla32_and7972_y0;
  wire h_u_cla32_and7973_y0;
  wire h_u_cla32_and7974_y0;
  wire h_u_cla32_and7975_y0;
  wire h_u_cla32_and7976_y0;
  wire h_u_cla32_and7977_y0;
  wire h_u_cla32_and7978_y0;
  wire h_u_cla32_and7979_y0;
  wire h_u_cla32_and7980_y0;
  wire h_u_cla32_and7981_y0;
  wire h_u_cla32_and7982_y0;
  wire h_u_cla32_and7983_y0;
  wire h_u_cla32_and7984_y0;
  wire h_u_cla32_and7985_y0;
  wire h_u_cla32_and7986_y0;
  wire h_u_cla32_and7987_y0;
  wire h_u_cla32_and7988_y0;
  wire h_u_cla32_and7989_y0;
  wire h_u_cla32_and7990_y0;
  wire h_u_cla32_and7991_y0;
  wire h_u_cla32_and7992_y0;
  wire h_u_cla32_and7993_y0;
  wire h_u_cla32_and7994_y0;
  wire h_u_cla32_and7995_y0;
  wire h_u_cla32_and7996_y0;
  wire h_u_cla32_and7997_y0;
  wire h_u_cla32_and7998_y0;
  wire h_u_cla32_and7999_y0;
  wire h_u_cla32_and8000_y0;
  wire h_u_cla32_and8001_y0;
  wire h_u_cla32_and8002_y0;
  wire h_u_cla32_and8003_y0;
  wire h_u_cla32_and8004_y0;
  wire h_u_cla32_and8005_y0;
  wire h_u_cla32_and8006_y0;
  wire h_u_cla32_and8007_y0;
  wire h_u_cla32_and8008_y0;
  wire h_u_cla32_and8009_y0;
  wire h_u_cla32_and8010_y0;
  wire h_u_cla32_and8011_y0;
  wire h_u_cla32_and8012_y0;
  wire h_u_cla32_and8013_y0;
  wire h_u_cla32_and8014_y0;
  wire h_u_cla32_and8015_y0;
  wire h_u_cla32_and8016_y0;
  wire h_u_cla32_and8017_y0;
  wire h_u_cla32_and8018_y0;
  wire h_u_cla32_and8019_y0;
  wire h_u_cla32_and8020_y0;
  wire h_u_cla32_and8021_y0;
  wire h_u_cla32_and8022_y0;
  wire h_u_cla32_and8023_y0;
  wire h_u_cla32_and8024_y0;
  wire h_u_cla32_and8025_y0;
  wire h_u_cla32_and8026_y0;
  wire h_u_cla32_and8027_y0;
  wire h_u_cla32_and8028_y0;
  wire h_u_cla32_and8029_y0;
  wire h_u_cla32_and8030_y0;
  wire h_u_cla32_and8031_y0;
  wire h_u_cla32_and8032_y0;
  wire h_u_cla32_and8033_y0;
  wire h_u_cla32_and8034_y0;
  wire h_u_cla32_and8035_y0;
  wire h_u_cla32_and8036_y0;
  wire h_u_cla32_and8037_y0;
  wire h_u_cla32_and8038_y0;
  wire h_u_cla32_and8039_y0;
  wire h_u_cla32_and8040_y0;
  wire h_u_cla32_and8041_y0;
  wire h_u_cla32_and8042_y0;
  wire h_u_cla32_and8043_y0;
  wire h_u_cla32_and8044_y0;
  wire h_u_cla32_and8045_y0;
  wire h_u_cla32_and8046_y0;
  wire h_u_cla32_and8047_y0;
  wire h_u_cla32_and8048_y0;
  wire h_u_cla32_and8049_y0;
  wire h_u_cla32_and8050_y0;
  wire h_u_cla32_and8051_y0;
  wire h_u_cla32_and8052_y0;
  wire h_u_cla32_and8053_y0;
  wire h_u_cla32_and8054_y0;
  wire h_u_cla32_and8055_y0;
  wire h_u_cla32_and8056_y0;
  wire h_u_cla32_and8057_y0;
  wire h_u_cla32_and8058_y0;
  wire h_u_cla32_and8059_y0;
  wire h_u_cla32_and8060_y0;
  wire h_u_cla32_and8061_y0;
  wire h_u_cla32_and8062_y0;
  wire h_u_cla32_and8063_y0;
  wire h_u_cla32_and8064_y0;
  wire h_u_cla32_and8065_y0;
  wire h_u_cla32_and8066_y0;
  wire h_u_cla32_and8067_y0;
  wire h_u_cla32_and8068_y0;
  wire h_u_cla32_and8069_y0;
  wire h_u_cla32_and8070_y0;
  wire h_u_cla32_and8071_y0;
  wire h_u_cla32_and8072_y0;
  wire h_u_cla32_and8073_y0;
  wire h_u_cla32_and8074_y0;
  wire h_u_cla32_and8075_y0;
  wire h_u_cla32_and8076_y0;
  wire h_u_cla32_and8077_y0;
  wire h_u_cla32_and8078_y0;
  wire h_u_cla32_and8079_y0;
  wire h_u_cla32_and8080_y0;
  wire h_u_cla32_and8081_y0;
  wire h_u_cla32_and8082_y0;
  wire h_u_cla32_and8083_y0;
  wire h_u_cla32_and8084_y0;
  wire h_u_cla32_and8085_y0;
  wire h_u_cla32_and8086_y0;
  wire h_u_cla32_and8087_y0;
  wire h_u_cla32_and8088_y0;
  wire h_u_cla32_and8089_y0;
  wire h_u_cla32_and8090_y0;
  wire h_u_cla32_and8091_y0;
  wire h_u_cla32_and8092_y0;
  wire h_u_cla32_and8093_y0;
  wire h_u_cla32_and8094_y0;
  wire h_u_cla32_and8095_y0;
  wire h_u_cla32_and8096_y0;
  wire h_u_cla32_and8097_y0;
  wire h_u_cla32_and8098_y0;
  wire h_u_cla32_and8099_y0;
  wire h_u_cla32_and8100_y0;
  wire h_u_cla32_and8101_y0;
  wire h_u_cla32_and8102_y0;
  wire h_u_cla32_and8103_y0;
  wire h_u_cla32_and8104_y0;
  wire h_u_cla32_and8105_y0;
  wire h_u_cla32_and8106_y0;
  wire h_u_cla32_and8107_y0;
  wire h_u_cla32_and8108_y0;
  wire h_u_cla32_and8109_y0;
  wire h_u_cla32_and8110_y0;
  wire h_u_cla32_and8111_y0;
  wire h_u_cla32_and8112_y0;
  wire h_u_cla32_and8113_y0;
  wire h_u_cla32_and8114_y0;
  wire h_u_cla32_and8115_y0;
  wire h_u_cla32_and8116_y0;
  wire h_u_cla32_and8117_y0;
  wire h_u_cla32_and8118_y0;
  wire h_u_cla32_and8119_y0;
  wire h_u_cla32_and8120_y0;
  wire h_u_cla32_and8121_y0;
  wire h_u_cla32_and8122_y0;
  wire h_u_cla32_and8123_y0;
  wire h_u_cla32_and8124_y0;
  wire h_u_cla32_and8125_y0;
  wire h_u_cla32_and8126_y0;
  wire h_u_cla32_and8127_y0;
  wire h_u_cla32_and8128_y0;
  wire h_u_cla32_and8129_y0;
  wire h_u_cla32_and8130_y0;
  wire h_u_cla32_and8131_y0;
  wire h_u_cla32_and8132_y0;
  wire h_u_cla32_and8133_y0;
  wire h_u_cla32_and8134_y0;
  wire h_u_cla32_and8135_y0;
  wire h_u_cla32_and8136_y0;
  wire h_u_cla32_and8137_y0;
  wire h_u_cla32_and8138_y0;
  wire h_u_cla32_and8139_y0;
  wire h_u_cla32_and8140_y0;
  wire h_u_cla32_and8141_y0;
  wire h_u_cla32_and8142_y0;
  wire h_u_cla32_and8143_y0;
  wire h_u_cla32_and8144_y0;
  wire h_u_cla32_and8145_y0;
  wire h_u_cla32_and8146_y0;
  wire h_u_cla32_and8147_y0;
  wire h_u_cla32_and8148_y0;
  wire h_u_cla32_and8149_y0;
  wire h_u_cla32_and8150_y0;
  wire h_u_cla32_and8151_y0;
  wire h_u_cla32_and8152_y0;
  wire h_u_cla32_and8153_y0;
  wire h_u_cla32_and8154_y0;
  wire h_u_cla32_and8155_y0;
  wire h_u_cla32_and8156_y0;
  wire h_u_cla32_and8157_y0;
  wire h_u_cla32_and8158_y0;
  wire h_u_cla32_and8159_y0;
  wire h_u_cla32_and8160_y0;
  wire h_u_cla32_and8161_y0;
  wire h_u_cla32_and8162_y0;
  wire h_u_cla32_and8163_y0;
  wire h_u_cla32_and8164_y0;
  wire h_u_cla32_and8165_y0;
  wire h_u_cla32_and8166_y0;
  wire h_u_cla32_and8167_y0;
  wire h_u_cla32_and8168_y0;
  wire h_u_cla32_and8169_y0;
  wire h_u_cla32_and8170_y0;
  wire h_u_cla32_and8171_y0;
  wire h_u_cla32_and8172_y0;
  wire h_u_cla32_and8173_y0;
  wire h_u_cla32_and8174_y0;
  wire h_u_cla32_and8175_y0;
  wire h_u_cla32_and8176_y0;
  wire h_u_cla32_and8177_y0;
  wire h_u_cla32_and8178_y0;
  wire h_u_cla32_and8179_y0;
  wire h_u_cla32_and8180_y0;
  wire h_u_cla32_and8181_y0;
  wire h_u_cla32_and8182_y0;
  wire h_u_cla32_and8183_y0;
  wire h_u_cla32_and8184_y0;
  wire h_u_cla32_and8185_y0;
  wire h_u_cla32_and8186_y0;
  wire h_u_cla32_and8187_y0;
  wire h_u_cla32_and8188_y0;
  wire h_u_cla32_and8189_y0;
  wire h_u_cla32_and8190_y0;
  wire h_u_cla32_and8191_y0;
  wire h_u_cla32_and8192_y0;
  wire h_u_cla32_and8193_y0;
  wire h_u_cla32_and8194_y0;
  wire h_u_cla32_and8195_y0;
  wire h_u_cla32_and8196_y0;
  wire h_u_cla32_and8197_y0;
  wire h_u_cla32_and8198_y0;
  wire h_u_cla32_and8199_y0;
  wire h_u_cla32_and8200_y0;
  wire h_u_cla32_and8201_y0;
  wire h_u_cla32_and8202_y0;
  wire h_u_cla32_and8203_y0;
  wire h_u_cla32_and8204_y0;
  wire h_u_cla32_and8205_y0;
  wire h_u_cla32_and8206_y0;
  wire h_u_cla32_and8207_y0;
  wire h_u_cla32_and8208_y0;
  wire h_u_cla32_and8209_y0;
  wire h_u_cla32_and8210_y0;
  wire h_u_cla32_and8211_y0;
  wire h_u_cla32_and8212_y0;
  wire h_u_cla32_and8213_y0;
  wire h_u_cla32_and8214_y0;
  wire h_u_cla32_and8215_y0;
  wire h_u_cla32_and8216_y0;
  wire h_u_cla32_and8217_y0;
  wire h_u_cla32_and8218_y0;
  wire h_u_cla32_and8219_y0;
  wire h_u_cla32_and8220_y0;
  wire h_u_cla32_and8221_y0;
  wire h_u_cla32_and8222_y0;
  wire h_u_cla32_and8223_y0;
  wire h_u_cla32_and8224_y0;
  wire h_u_cla32_and8225_y0;
  wire h_u_cla32_and8226_y0;
  wire h_u_cla32_and8227_y0;
  wire h_u_cla32_and8228_y0;
  wire h_u_cla32_and8229_y0;
  wire h_u_cla32_and8230_y0;
  wire h_u_cla32_and8231_y0;
  wire h_u_cla32_and8232_y0;
  wire h_u_cla32_and8233_y0;
  wire h_u_cla32_and8234_y0;
  wire h_u_cla32_and8235_y0;
  wire h_u_cla32_and8236_y0;
  wire h_u_cla32_and8237_y0;
  wire h_u_cla32_and8238_y0;
  wire h_u_cla32_and8239_y0;
  wire h_u_cla32_and8240_y0;
  wire h_u_cla32_and8241_y0;
  wire h_u_cla32_and8242_y0;
  wire h_u_cla32_and8243_y0;
  wire h_u_cla32_and8244_y0;
  wire h_u_cla32_and8245_y0;
  wire h_u_cla32_and8246_y0;
  wire h_u_cla32_and8247_y0;
  wire h_u_cla32_and8248_y0;
  wire h_u_cla32_and8249_y0;
  wire h_u_cla32_and8250_y0;
  wire h_u_cla32_and8251_y0;
  wire h_u_cla32_and8252_y0;
  wire h_u_cla32_and8253_y0;
  wire h_u_cla32_and8254_y0;
  wire h_u_cla32_and8255_y0;
  wire h_u_cla32_and8256_y0;
  wire h_u_cla32_and8257_y0;
  wire h_u_cla32_and8258_y0;
  wire h_u_cla32_and8259_y0;
  wire h_u_cla32_and8260_y0;
  wire h_u_cla32_and8261_y0;
  wire h_u_cla32_and8262_y0;
  wire h_u_cla32_and8263_y0;
  wire h_u_cla32_and8264_y0;
  wire h_u_cla32_and8265_y0;
  wire h_u_cla32_and8266_y0;
  wire h_u_cla32_and8267_y0;
  wire h_u_cla32_and8268_y0;
  wire h_u_cla32_and8269_y0;
  wire h_u_cla32_and8270_y0;
  wire h_u_cla32_and8271_y0;
  wire h_u_cla32_and8272_y0;
  wire h_u_cla32_and8273_y0;
  wire h_u_cla32_and8274_y0;
  wire h_u_cla32_and8275_y0;
  wire h_u_cla32_and8276_y0;
  wire h_u_cla32_and8277_y0;
  wire h_u_cla32_and8278_y0;
  wire h_u_cla32_and8279_y0;
  wire h_u_cla32_and8280_y0;
  wire h_u_cla32_and8281_y0;
  wire h_u_cla32_and8282_y0;
  wire h_u_cla32_and8283_y0;
  wire h_u_cla32_and8284_y0;
  wire h_u_cla32_and8285_y0;
  wire h_u_cla32_and8286_y0;
  wire h_u_cla32_and8287_y0;
  wire h_u_cla32_and8288_y0;
  wire h_u_cla32_and8289_y0;
  wire h_u_cla32_and8290_y0;
  wire h_u_cla32_and8291_y0;
  wire h_u_cla32_and8292_y0;
  wire h_u_cla32_and8293_y0;
  wire h_u_cla32_and8294_y0;
  wire h_u_cla32_and8295_y0;
  wire h_u_cla32_and8296_y0;
  wire h_u_cla32_and8297_y0;
  wire h_u_cla32_and8298_y0;
  wire h_u_cla32_and8299_y0;
  wire h_u_cla32_and8300_y0;
  wire h_u_cla32_and8301_y0;
  wire h_u_cla32_and8302_y0;
  wire h_u_cla32_and8303_y0;
  wire h_u_cla32_and8304_y0;
  wire h_u_cla32_and8305_y0;
  wire h_u_cla32_and8306_y0;
  wire h_u_cla32_and8307_y0;
  wire h_u_cla32_and8308_y0;
  wire h_u_cla32_and8309_y0;
  wire h_u_cla32_and8310_y0;
  wire h_u_cla32_and8311_y0;
  wire h_u_cla32_and8312_y0;
  wire h_u_cla32_and8313_y0;
  wire h_u_cla32_and8314_y0;
  wire h_u_cla32_and8315_y0;
  wire h_u_cla32_and8316_y0;
  wire h_u_cla32_and8317_y0;
  wire h_u_cla32_and8318_y0;
  wire h_u_cla32_and8319_y0;
  wire h_u_cla32_and8320_y0;
  wire h_u_cla32_and8321_y0;
  wire h_u_cla32_and8322_y0;
  wire h_u_cla32_and8323_y0;
  wire h_u_cla32_and8324_y0;
  wire h_u_cla32_and8325_y0;
  wire h_u_cla32_and8326_y0;
  wire h_u_cla32_and8327_y0;
  wire h_u_cla32_and8328_y0;
  wire h_u_cla32_and8329_y0;
  wire h_u_cla32_and8330_y0;
  wire h_u_cla32_and8331_y0;
  wire h_u_cla32_and8332_y0;
  wire h_u_cla32_and8333_y0;
  wire h_u_cla32_and8334_y0;
  wire h_u_cla32_and8335_y0;
  wire h_u_cla32_and8336_y0;
  wire h_u_cla32_and8337_y0;
  wire h_u_cla32_and8338_y0;
  wire h_u_cla32_and8339_y0;
  wire h_u_cla32_and8340_y0;
  wire h_u_cla32_and8341_y0;
  wire h_u_cla32_and8342_y0;
  wire h_u_cla32_and8343_y0;
  wire h_u_cla32_and8344_y0;
  wire h_u_cla32_and8345_y0;
  wire h_u_cla32_and8346_y0;
  wire h_u_cla32_and8347_y0;
  wire h_u_cla32_and8348_y0;
  wire h_u_cla32_and8349_y0;
  wire h_u_cla32_and8350_y0;
  wire h_u_cla32_and8351_y0;
  wire h_u_cla32_and8352_y0;
  wire h_u_cla32_and8353_y0;
  wire h_u_cla32_and8354_y0;
  wire h_u_cla32_and8355_y0;
  wire h_u_cla32_and8356_y0;
  wire h_u_cla32_and8357_y0;
  wire h_u_cla32_and8358_y0;
  wire h_u_cla32_and8359_y0;
  wire h_u_cla32_and8360_y0;
  wire h_u_cla32_and8361_y0;
  wire h_u_cla32_and8362_y0;
  wire h_u_cla32_and8363_y0;
  wire h_u_cla32_and8364_y0;
  wire h_u_cla32_and8365_y0;
  wire h_u_cla32_and8366_y0;
  wire h_u_cla32_and8367_y0;
  wire h_u_cla32_and8368_y0;
  wire h_u_cla32_and8369_y0;
  wire h_u_cla32_and8370_y0;
  wire h_u_cla32_and8371_y0;
  wire h_u_cla32_and8372_y0;
  wire h_u_cla32_and8373_y0;
  wire h_u_cla32_and8374_y0;
  wire h_u_cla32_and8375_y0;
  wire h_u_cla32_and8376_y0;
  wire h_u_cla32_and8377_y0;
  wire h_u_cla32_and8378_y0;
  wire h_u_cla32_and8379_y0;
  wire h_u_cla32_and8380_y0;
  wire h_u_cla32_and8381_y0;
  wire h_u_cla32_and8382_y0;
  wire h_u_cla32_and8383_y0;
  wire h_u_cla32_and8384_y0;
  wire h_u_cla32_and8385_y0;
  wire h_u_cla32_and8386_y0;
  wire h_u_cla32_and8387_y0;
  wire h_u_cla32_and8388_y0;
  wire h_u_cla32_and8389_y0;
  wire h_u_cla32_and8390_y0;
  wire h_u_cla32_and8391_y0;
  wire h_u_cla32_and8392_y0;
  wire h_u_cla32_and8393_y0;
  wire h_u_cla32_and8394_y0;
  wire h_u_cla32_and8395_y0;
  wire h_u_cla32_and8396_y0;
  wire h_u_cla32_and8397_y0;
  wire h_u_cla32_and8398_y0;
  wire h_u_cla32_and8399_y0;
  wire h_u_cla32_and8400_y0;
  wire h_u_cla32_and8401_y0;
  wire h_u_cla32_and8402_y0;
  wire h_u_cla32_and8403_y0;
  wire h_u_cla32_and8404_y0;
  wire h_u_cla32_and8405_y0;
  wire h_u_cla32_and8406_y0;
  wire h_u_cla32_and8407_y0;
  wire h_u_cla32_and8408_y0;
  wire h_u_cla32_and8409_y0;
  wire h_u_cla32_and8410_y0;
  wire h_u_cla32_and8411_y0;
  wire h_u_cla32_and8412_y0;
  wire h_u_cla32_and8413_y0;
  wire h_u_cla32_and8414_y0;
  wire h_u_cla32_and8415_y0;
  wire h_u_cla32_and8416_y0;
  wire h_u_cla32_and8417_y0;
  wire h_u_cla32_and8418_y0;
  wire h_u_cla32_and8419_y0;
  wire h_u_cla32_and8420_y0;
  wire h_u_cla32_and8421_y0;
  wire h_u_cla32_and8422_y0;
  wire h_u_cla32_and8423_y0;
  wire h_u_cla32_and8424_y0;
  wire h_u_cla32_and8425_y0;
  wire h_u_cla32_and8426_y0;
  wire h_u_cla32_and8427_y0;
  wire h_u_cla32_and8428_y0;
  wire h_u_cla32_and8429_y0;
  wire h_u_cla32_and8430_y0;
  wire h_u_cla32_and8431_y0;
  wire h_u_cla32_and8432_y0;
  wire h_u_cla32_and8433_y0;
  wire h_u_cla32_and8434_y0;
  wire h_u_cla32_and8435_y0;
  wire h_u_cla32_and8436_y0;
  wire h_u_cla32_and8437_y0;
  wire h_u_cla32_and8438_y0;
  wire h_u_cla32_and8439_y0;
  wire h_u_cla32_and8440_y0;
  wire h_u_cla32_and8441_y0;
  wire h_u_cla32_and8442_y0;
  wire h_u_cla32_and8443_y0;
  wire h_u_cla32_and8444_y0;
  wire h_u_cla32_and8445_y0;
  wire h_u_cla32_and8446_y0;
  wire h_u_cla32_and8447_y0;
  wire h_u_cla32_and8448_y0;
  wire h_u_cla32_and8449_y0;
  wire h_u_cla32_and8450_y0;
  wire h_u_cla32_and8451_y0;
  wire h_u_cla32_and8452_y0;
  wire h_u_cla32_and8453_y0;
  wire h_u_cla32_and8454_y0;
  wire h_u_cla32_and8455_y0;
  wire h_u_cla32_and8456_y0;
  wire h_u_cla32_and8457_y0;
  wire h_u_cla32_and8458_y0;
  wire h_u_cla32_and8459_y0;
  wire h_u_cla32_and8460_y0;
  wire h_u_cla32_and8461_y0;
  wire h_u_cla32_and8462_y0;
  wire h_u_cla32_and8463_y0;
  wire h_u_cla32_and8464_y0;
  wire h_u_cla32_and8465_y0;
  wire h_u_cla32_and8466_y0;
  wire h_u_cla32_and8467_y0;
  wire h_u_cla32_and8468_y0;
  wire h_u_cla32_and8469_y0;
  wire h_u_cla32_and8470_y0;
  wire h_u_cla32_and8471_y0;
  wire h_u_cla32_and8472_y0;
  wire h_u_cla32_and8473_y0;
  wire h_u_cla32_and8474_y0;
  wire h_u_cla32_and8475_y0;
  wire h_u_cla32_and8476_y0;
  wire h_u_cla32_and8477_y0;
  wire h_u_cla32_and8478_y0;
  wire h_u_cla32_and8479_y0;
  wire h_u_cla32_and8480_y0;
  wire h_u_cla32_and8481_y0;
  wire h_u_cla32_and8482_y0;
  wire h_u_cla32_and8483_y0;
  wire h_u_cla32_and8484_y0;
  wire h_u_cla32_and8485_y0;
  wire h_u_cla32_and8486_y0;
  wire h_u_cla32_and8487_y0;
  wire h_u_cla32_and8488_y0;
  wire h_u_cla32_and8489_y0;
  wire h_u_cla32_and8490_y0;
  wire h_u_cla32_and8491_y0;
  wire h_u_cla32_and8492_y0;
  wire h_u_cla32_and8493_y0;
  wire h_u_cla32_and8494_y0;
  wire h_u_cla32_and8495_y0;
  wire h_u_cla32_and8496_y0;
  wire h_u_cla32_and8497_y0;
  wire h_u_cla32_and8498_y0;
  wire h_u_cla32_and8499_y0;
  wire h_u_cla32_and8500_y0;
  wire h_u_cla32_and8501_y0;
  wire h_u_cla32_and8502_y0;
  wire h_u_cla32_and8503_y0;
  wire h_u_cla32_and8504_y0;
  wire h_u_cla32_and8505_y0;
  wire h_u_cla32_and8506_y0;
  wire h_u_cla32_and8507_y0;
  wire h_u_cla32_and8508_y0;
  wire h_u_cla32_and8509_y0;
  wire h_u_cla32_and8510_y0;
  wire h_u_cla32_and8511_y0;
  wire h_u_cla32_and8512_y0;
  wire h_u_cla32_and8513_y0;
  wire h_u_cla32_and8514_y0;
  wire h_u_cla32_and8515_y0;
  wire h_u_cla32_and8516_y0;
  wire h_u_cla32_and8517_y0;
  wire h_u_cla32_and8518_y0;
  wire h_u_cla32_and8519_y0;
  wire h_u_cla32_and8520_y0;
  wire h_u_cla32_and8521_y0;
  wire h_u_cla32_and8522_y0;
  wire h_u_cla32_and8523_y0;
  wire h_u_cla32_and8524_y0;
  wire h_u_cla32_and8525_y0;
  wire h_u_cla32_and8526_y0;
  wire h_u_cla32_and8527_y0;
  wire h_u_cla32_and8528_y0;
  wire h_u_cla32_and8529_y0;
  wire h_u_cla32_and8530_y0;
  wire h_u_cla32_and8531_y0;
  wire h_u_cla32_and8532_y0;
  wire h_u_cla32_and8533_y0;
  wire h_u_cla32_and8534_y0;
  wire h_u_cla32_and8535_y0;
  wire h_u_cla32_and8536_y0;
  wire h_u_cla32_and8537_y0;
  wire h_u_cla32_and8538_y0;
  wire h_u_cla32_and8539_y0;
  wire h_u_cla32_and8540_y0;
  wire h_u_cla32_and8541_y0;
  wire h_u_cla32_and8542_y0;
  wire h_u_cla32_and8543_y0;
  wire h_u_cla32_and8544_y0;
  wire h_u_cla32_and8545_y0;
  wire h_u_cla32_and8546_y0;
  wire h_u_cla32_and8547_y0;
  wire h_u_cla32_and8548_y0;
  wire h_u_cla32_and8549_y0;
  wire h_u_cla32_and8550_y0;
  wire h_u_cla32_and8551_y0;
  wire h_u_cla32_and8552_y0;
  wire h_u_cla32_and8553_y0;
  wire h_u_cla32_and8554_y0;
  wire h_u_cla32_or406_y0;
  wire h_u_cla32_or407_y0;
  wire h_u_cla32_or408_y0;
  wire h_u_cla32_or409_y0;
  wire h_u_cla32_or410_y0;
  wire h_u_cla32_or411_y0;
  wire h_u_cla32_or412_y0;
  wire h_u_cla32_or413_y0;
  wire h_u_cla32_or414_y0;
  wire h_u_cla32_or415_y0;
  wire h_u_cla32_or416_y0;
  wire h_u_cla32_or417_y0;
  wire h_u_cla32_or418_y0;
  wire h_u_cla32_or419_y0;
  wire h_u_cla32_or420_y0;
  wire h_u_cla32_or421_y0;
  wire h_u_cla32_or422_y0;
  wire h_u_cla32_or423_y0;
  wire h_u_cla32_or424_y0;
  wire h_u_cla32_or425_y0;
  wire h_u_cla32_or426_y0;
  wire h_u_cla32_or427_y0;
  wire h_u_cla32_or428_y0;
  wire h_u_cla32_or429_y0;
  wire h_u_cla32_or430_y0;
  wire h_u_cla32_or431_y0;
  wire h_u_cla32_or432_y0;
  wire h_u_cla32_or433_y0;
  wire h_u_cla32_or434_y0;
  wire h_u_cla32_pg_logic29_y0;
  wire h_u_cla32_pg_logic29_y1;
  wire h_u_cla32_pg_logic29_y2;
  wire h_u_cla32_xor29_y0;
  wire h_u_cla32_and8555_y0;
  wire h_u_cla32_and8556_y0;
  wire h_u_cla32_and8557_y0;
  wire h_u_cla32_and8558_y0;
  wire h_u_cla32_and8559_y0;
  wire h_u_cla32_and8560_y0;
  wire h_u_cla32_and8561_y0;
  wire h_u_cla32_and8562_y0;
  wire h_u_cla32_and8563_y0;
  wire h_u_cla32_and8564_y0;
  wire h_u_cla32_and8565_y0;
  wire h_u_cla32_and8566_y0;
  wire h_u_cla32_and8567_y0;
  wire h_u_cla32_and8568_y0;
  wire h_u_cla32_and8569_y0;
  wire h_u_cla32_and8570_y0;
  wire h_u_cla32_and8571_y0;
  wire h_u_cla32_and8572_y0;
  wire h_u_cla32_and8573_y0;
  wire h_u_cla32_and8574_y0;
  wire h_u_cla32_and8575_y0;
  wire h_u_cla32_and8576_y0;
  wire h_u_cla32_and8577_y0;
  wire h_u_cla32_and8578_y0;
  wire h_u_cla32_and8579_y0;
  wire h_u_cla32_and8580_y0;
  wire h_u_cla32_and8581_y0;
  wire h_u_cla32_and8582_y0;
  wire h_u_cla32_and8583_y0;
  wire h_u_cla32_and8584_y0;
  wire h_u_cla32_and8585_y0;
  wire h_u_cla32_and8586_y0;
  wire h_u_cla32_and8587_y0;
  wire h_u_cla32_and8588_y0;
  wire h_u_cla32_and8589_y0;
  wire h_u_cla32_and8590_y0;
  wire h_u_cla32_and8591_y0;
  wire h_u_cla32_and8592_y0;
  wire h_u_cla32_and8593_y0;
  wire h_u_cla32_and8594_y0;
  wire h_u_cla32_and8595_y0;
  wire h_u_cla32_and8596_y0;
  wire h_u_cla32_and8597_y0;
  wire h_u_cla32_and8598_y0;
  wire h_u_cla32_and8599_y0;
  wire h_u_cla32_and8600_y0;
  wire h_u_cla32_and8601_y0;
  wire h_u_cla32_and8602_y0;
  wire h_u_cla32_and8603_y0;
  wire h_u_cla32_and8604_y0;
  wire h_u_cla32_and8605_y0;
  wire h_u_cla32_and8606_y0;
  wire h_u_cla32_and8607_y0;
  wire h_u_cla32_and8608_y0;
  wire h_u_cla32_and8609_y0;
  wire h_u_cla32_and8610_y0;
  wire h_u_cla32_and8611_y0;
  wire h_u_cla32_and8612_y0;
  wire h_u_cla32_and8613_y0;
  wire h_u_cla32_and8614_y0;
  wire h_u_cla32_and8615_y0;
  wire h_u_cla32_and8616_y0;
  wire h_u_cla32_and8617_y0;
  wire h_u_cla32_and8618_y0;
  wire h_u_cla32_and8619_y0;
  wire h_u_cla32_and8620_y0;
  wire h_u_cla32_and8621_y0;
  wire h_u_cla32_and8622_y0;
  wire h_u_cla32_and8623_y0;
  wire h_u_cla32_and8624_y0;
  wire h_u_cla32_and8625_y0;
  wire h_u_cla32_and8626_y0;
  wire h_u_cla32_and8627_y0;
  wire h_u_cla32_and8628_y0;
  wire h_u_cla32_and8629_y0;
  wire h_u_cla32_and8630_y0;
  wire h_u_cla32_and8631_y0;
  wire h_u_cla32_and8632_y0;
  wire h_u_cla32_and8633_y0;
  wire h_u_cla32_and8634_y0;
  wire h_u_cla32_and8635_y0;
  wire h_u_cla32_and8636_y0;
  wire h_u_cla32_and8637_y0;
  wire h_u_cla32_and8638_y0;
  wire h_u_cla32_and8639_y0;
  wire h_u_cla32_and8640_y0;
  wire h_u_cla32_and8641_y0;
  wire h_u_cla32_and8642_y0;
  wire h_u_cla32_and8643_y0;
  wire h_u_cla32_and8644_y0;
  wire h_u_cla32_and8645_y0;
  wire h_u_cla32_and8646_y0;
  wire h_u_cla32_and8647_y0;
  wire h_u_cla32_and8648_y0;
  wire h_u_cla32_and8649_y0;
  wire h_u_cla32_and8650_y0;
  wire h_u_cla32_and8651_y0;
  wire h_u_cla32_and8652_y0;
  wire h_u_cla32_and8653_y0;
  wire h_u_cla32_and8654_y0;
  wire h_u_cla32_and8655_y0;
  wire h_u_cla32_and8656_y0;
  wire h_u_cla32_and8657_y0;
  wire h_u_cla32_and8658_y0;
  wire h_u_cla32_and8659_y0;
  wire h_u_cla32_and8660_y0;
  wire h_u_cla32_and8661_y0;
  wire h_u_cla32_and8662_y0;
  wire h_u_cla32_and8663_y0;
  wire h_u_cla32_and8664_y0;
  wire h_u_cla32_and8665_y0;
  wire h_u_cla32_and8666_y0;
  wire h_u_cla32_and8667_y0;
  wire h_u_cla32_and8668_y0;
  wire h_u_cla32_and8669_y0;
  wire h_u_cla32_and8670_y0;
  wire h_u_cla32_and8671_y0;
  wire h_u_cla32_and8672_y0;
  wire h_u_cla32_and8673_y0;
  wire h_u_cla32_and8674_y0;
  wire h_u_cla32_and8675_y0;
  wire h_u_cla32_and8676_y0;
  wire h_u_cla32_and8677_y0;
  wire h_u_cla32_and8678_y0;
  wire h_u_cla32_and8679_y0;
  wire h_u_cla32_and8680_y0;
  wire h_u_cla32_and8681_y0;
  wire h_u_cla32_and8682_y0;
  wire h_u_cla32_and8683_y0;
  wire h_u_cla32_and8684_y0;
  wire h_u_cla32_and8685_y0;
  wire h_u_cla32_and8686_y0;
  wire h_u_cla32_and8687_y0;
  wire h_u_cla32_and8688_y0;
  wire h_u_cla32_and8689_y0;
  wire h_u_cla32_and8690_y0;
  wire h_u_cla32_and8691_y0;
  wire h_u_cla32_and8692_y0;
  wire h_u_cla32_and8693_y0;
  wire h_u_cla32_and8694_y0;
  wire h_u_cla32_and8695_y0;
  wire h_u_cla32_and8696_y0;
  wire h_u_cla32_and8697_y0;
  wire h_u_cla32_and8698_y0;
  wire h_u_cla32_and8699_y0;
  wire h_u_cla32_and8700_y0;
  wire h_u_cla32_and8701_y0;
  wire h_u_cla32_and8702_y0;
  wire h_u_cla32_and8703_y0;
  wire h_u_cla32_and8704_y0;
  wire h_u_cla32_and8705_y0;
  wire h_u_cla32_and8706_y0;
  wire h_u_cla32_and8707_y0;
  wire h_u_cla32_and8708_y0;
  wire h_u_cla32_and8709_y0;
  wire h_u_cla32_and8710_y0;
  wire h_u_cla32_and8711_y0;
  wire h_u_cla32_and8712_y0;
  wire h_u_cla32_and8713_y0;
  wire h_u_cla32_and8714_y0;
  wire h_u_cla32_and8715_y0;
  wire h_u_cla32_and8716_y0;
  wire h_u_cla32_and8717_y0;
  wire h_u_cla32_and8718_y0;
  wire h_u_cla32_and8719_y0;
  wire h_u_cla32_and8720_y0;
  wire h_u_cla32_and8721_y0;
  wire h_u_cla32_and8722_y0;
  wire h_u_cla32_and8723_y0;
  wire h_u_cla32_and8724_y0;
  wire h_u_cla32_and8725_y0;
  wire h_u_cla32_and8726_y0;
  wire h_u_cla32_and8727_y0;
  wire h_u_cla32_and8728_y0;
  wire h_u_cla32_and8729_y0;
  wire h_u_cla32_and8730_y0;
  wire h_u_cla32_and8731_y0;
  wire h_u_cla32_and8732_y0;
  wire h_u_cla32_and8733_y0;
  wire h_u_cla32_and8734_y0;
  wire h_u_cla32_and8735_y0;
  wire h_u_cla32_and8736_y0;
  wire h_u_cla32_and8737_y0;
  wire h_u_cla32_and8738_y0;
  wire h_u_cla32_and8739_y0;
  wire h_u_cla32_and8740_y0;
  wire h_u_cla32_and8741_y0;
  wire h_u_cla32_and8742_y0;
  wire h_u_cla32_and8743_y0;
  wire h_u_cla32_and8744_y0;
  wire h_u_cla32_and8745_y0;
  wire h_u_cla32_and8746_y0;
  wire h_u_cla32_and8747_y0;
  wire h_u_cla32_and8748_y0;
  wire h_u_cla32_and8749_y0;
  wire h_u_cla32_and8750_y0;
  wire h_u_cla32_and8751_y0;
  wire h_u_cla32_and8752_y0;
  wire h_u_cla32_and8753_y0;
  wire h_u_cla32_and8754_y0;
  wire h_u_cla32_and8755_y0;
  wire h_u_cla32_and8756_y0;
  wire h_u_cla32_and8757_y0;
  wire h_u_cla32_and8758_y0;
  wire h_u_cla32_and8759_y0;
  wire h_u_cla32_and8760_y0;
  wire h_u_cla32_and8761_y0;
  wire h_u_cla32_and8762_y0;
  wire h_u_cla32_and8763_y0;
  wire h_u_cla32_and8764_y0;
  wire h_u_cla32_and8765_y0;
  wire h_u_cla32_and8766_y0;
  wire h_u_cla32_and8767_y0;
  wire h_u_cla32_and8768_y0;
  wire h_u_cla32_and8769_y0;
  wire h_u_cla32_and8770_y0;
  wire h_u_cla32_and8771_y0;
  wire h_u_cla32_and8772_y0;
  wire h_u_cla32_and8773_y0;
  wire h_u_cla32_and8774_y0;
  wire h_u_cla32_and8775_y0;
  wire h_u_cla32_and8776_y0;
  wire h_u_cla32_and8777_y0;
  wire h_u_cla32_and8778_y0;
  wire h_u_cla32_and8779_y0;
  wire h_u_cla32_and8780_y0;
  wire h_u_cla32_and8781_y0;
  wire h_u_cla32_and8782_y0;
  wire h_u_cla32_and8783_y0;
  wire h_u_cla32_and8784_y0;
  wire h_u_cla32_and8785_y0;
  wire h_u_cla32_and8786_y0;
  wire h_u_cla32_and8787_y0;
  wire h_u_cla32_and8788_y0;
  wire h_u_cla32_and8789_y0;
  wire h_u_cla32_and8790_y0;
  wire h_u_cla32_and8791_y0;
  wire h_u_cla32_and8792_y0;
  wire h_u_cla32_and8793_y0;
  wire h_u_cla32_and8794_y0;
  wire h_u_cla32_and8795_y0;
  wire h_u_cla32_and8796_y0;
  wire h_u_cla32_and8797_y0;
  wire h_u_cla32_and8798_y0;
  wire h_u_cla32_and8799_y0;
  wire h_u_cla32_and8800_y0;
  wire h_u_cla32_and8801_y0;
  wire h_u_cla32_and8802_y0;
  wire h_u_cla32_and8803_y0;
  wire h_u_cla32_and8804_y0;
  wire h_u_cla32_and8805_y0;
  wire h_u_cla32_and8806_y0;
  wire h_u_cla32_and8807_y0;
  wire h_u_cla32_and8808_y0;
  wire h_u_cla32_and8809_y0;
  wire h_u_cla32_and8810_y0;
  wire h_u_cla32_and8811_y0;
  wire h_u_cla32_and8812_y0;
  wire h_u_cla32_and8813_y0;
  wire h_u_cla32_and8814_y0;
  wire h_u_cla32_and8815_y0;
  wire h_u_cla32_and8816_y0;
  wire h_u_cla32_and8817_y0;
  wire h_u_cla32_and8818_y0;
  wire h_u_cla32_and8819_y0;
  wire h_u_cla32_and8820_y0;
  wire h_u_cla32_and8821_y0;
  wire h_u_cla32_and8822_y0;
  wire h_u_cla32_and8823_y0;
  wire h_u_cla32_and8824_y0;
  wire h_u_cla32_and8825_y0;
  wire h_u_cla32_and8826_y0;
  wire h_u_cla32_and8827_y0;
  wire h_u_cla32_and8828_y0;
  wire h_u_cla32_and8829_y0;
  wire h_u_cla32_and8830_y0;
  wire h_u_cla32_and8831_y0;
  wire h_u_cla32_and8832_y0;
  wire h_u_cla32_and8833_y0;
  wire h_u_cla32_and8834_y0;
  wire h_u_cla32_and8835_y0;
  wire h_u_cla32_and8836_y0;
  wire h_u_cla32_and8837_y0;
  wire h_u_cla32_and8838_y0;
  wire h_u_cla32_and8839_y0;
  wire h_u_cla32_and8840_y0;
  wire h_u_cla32_and8841_y0;
  wire h_u_cla32_and8842_y0;
  wire h_u_cla32_and8843_y0;
  wire h_u_cla32_and8844_y0;
  wire h_u_cla32_and8845_y0;
  wire h_u_cla32_and8846_y0;
  wire h_u_cla32_and8847_y0;
  wire h_u_cla32_and8848_y0;
  wire h_u_cla32_and8849_y0;
  wire h_u_cla32_and8850_y0;
  wire h_u_cla32_and8851_y0;
  wire h_u_cla32_and8852_y0;
  wire h_u_cla32_and8853_y0;
  wire h_u_cla32_and8854_y0;
  wire h_u_cla32_and8855_y0;
  wire h_u_cla32_and8856_y0;
  wire h_u_cla32_and8857_y0;
  wire h_u_cla32_and8858_y0;
  wire h_u_cla32_and8859_y0;
  wire h_u_cla32_and8860_y0;
  wire h_u_cla32_and8861_y0;
  wire h_u_cla32_and8862_y0;
  wire h_u_cla32_and8863_y0;
  wire h_u_cla32_and8864_y0;
  wire h_u_cla32_and8865_y0;
  wire h_u_cla32_and8866_y0;
  wire h_u_cla32_and8867_y0;
  wire h_u_cla32_and8868_y0;
  wire h_u_cla32_and8869_y0;
  wire h_u_cla32_and8870_y0;
  wire h_u_cla32_and8871_y0;
  wire h_u_cla32_and8872_y0;
  wire h_u_cla32_and8873_y0;
  wire h_u_cla32_and8874_y0;
  wire h_u_cla32_and8875_y0;
  wire h_u_cla32_and8876_y0;
  wire h_u_cla32_and8877_y0;
  wire h_u_cla32_and8878_y0;
  wire h_u_cla32_and8879_y0;
  wire h_u_cla32_and8880_y0;
  wire h_u_cla32_and8881_y0;
  wire h_u_cla32_and8882_y0;
  wire h_u_cla32_and8883_y0;
  wire h_u_cla32_and8884_y0;
  wire h_u_cla32_and8885_y0;
  wire h_u_cla32_and8886_y0;
  wire h_u_cla32_and8887_y0;
  wire h_u_cla32_and8888_y0;
  wire h_u_cla32_and8889_y0;
  wire h_u_cla32_and8890_y0;
  wire h_u_cla32_and8891_y0;
  wire h_u_cla32_and8892_y0;
  wire h_u_cla32_and8893_y0;
  wire h_u_cla32_and8894_y0;
  wire h_u_cla32_and8895_y0;
  wire h_u_cla32_and8896_y0;
  wire h_u_cla32_and8897_y0;
  wire h_u_cla32_and8898_y0;
  wire h_u_cla32_and8899_y0;
  wire h_u_cla32_and8900_y0;
  wire h_u_cla32_and8901_y0;
  wire h_u_cla32_and8902_y0;
  wire h_u_cla32_and8903_y0;
  wire h_u_cla32_and8904_y0;
  wire h_u_cla32_and8905_y0;
  wire h_u_cla32_and8906_y0;
  wire h_u_cla32_and8907_y0;
  wire h_u_cla32_and8908_y0;
  wire h_u_cla32_and8909_y0;
  wire h_u_cla32_and8910_y0;
  wire h_u_cla32_and8911_y0;
  wire h_u_cla32_and8912_y0;
  wire h_u_cla32_and8913_y0;
  wire h_u_cla32_and8914_y0;
  wire h_u_cla32_and8915_y0;
  wire h_u_cla32_and8916_y0;
  wire h_u_cla32_and8917_y0;
  wire h_u_cla32_and8918_y0;
  wire h_u_cla32_and8919_y0;
  wire h_u_cla32_and8920_y0;
  wire h_u_cla32_and8921_y0;
  wire h_u_cla32_and8922_y0;
  wire h_u_cla32_and8923_y0;
  wire h_u_cla32_and8924_y0;
  wire h_u_cla32_and8925_y0;
  wire h_u_cla32_and8926_y0;
  wire h_u_cla32_and8927_y0;
  wire h_u_cla32_and8928_y0;
  wire h_u_cla32_and8929_y0;
  wire h_u_cla32_and8930_y0;
  wire h_u_cla32_and8931_y0;
  wire h_u_cla32_and8932_y0;
  wire h_u_cla32_and8933_y0;
  wire h_u_cla32_and8934_y0;
  wire h_u_cla32_and8935_y0;
  wire h_u_cla32_and8936_y0;
  wire h_u_cla32_and8937_y0;
  wire h_u_cla32_and8938_y0;
  wire h_u_cla32_and8939_y0;
  wire h_u_cla32_and8940_y0;
  wire h_u_cla32_and8941_y0;
  wire h_u_cla32_and8942_y0;
  wire h_u_cla32_and8943_y0;
  wire h_u_cla32_and8944_y0;
  wire h_u_cla32_and8945_y0;
  wire h_u_cla32_and8946_y0;
  wire h_u_cla32_and8947_y0;
  wire h_u_cla32_and8948_y0;
  wire h_u_cla32_and8949_y0;
  wire h_u_cla32_and8950_y0;
  wire h_u_cla32_and8951_y0;
  wire h_u_cla32_and8952_y0;
  wire h_u_cla32_and8953_y0;
  wire h_u_cla32_and8954_y0;
  wire h_u_cla32_and8955_y0;
  wire h_u_cla32_and8956_y0;
  wire h_u_cla32_and8957_y0;
  wire h_u_cla32_and8958_y0;
  wire h_u_cla32_and8959_y0;
  wire h_u_cla32_and8960_y0;
  wire h_u_cla32_and8961_y0;
  wire h_u_cla32_and8962_y0;
  wire h_u_cla32_and8963_y0;
  wire h_u_cla32_and8964_y0;
  wire h_u_cla32_and8965_y0;
  wire h_u_cla32_and8966_y0;
  wire h_u_cla32_and8967_y0;
  wire h_u_cla32_and8968_y0;
  wire h_u_cla32_and8969_y0;
  wire h_u_cla32_and8970_y0;
  wire h_u_cla32_and8971_y0;
  wire h_u_cla32_and8972_y0;
  wire h_u_cla32_and8973_y0;
  wire h_u_cla32_and8974_y0;
  wire h_u_cla32_and8975_y0;
  wire h_u_cla32_and8976_y0;
  wire h_u_cla32_and8977_y0;
  wire h_u_cla32_and8978_y0;
  wire h_u_cla32_and8979_y0;
  wire h_u_cla32_and8980_y0;
  wire h_u_cla32_and8981_y0;
  wire h_u_cla32_and8982_y0;
  wire h_u_cla32_and8983_y0;
  wire h_u_cla32_and8984_y0;
  wire h_u_cla32_and8985_y0;
  wire h_u_cla32_and8986_y0;
  wire h_u_cla32_and8987_y0;
  wire h_u_cla32_and8988_y0;
  wire h_u_cla32_and8989_y0;
  wire h_u_cla32_and8990_y0;
  wire h_u_cla32_and8991_y0;
  wire h_u_cla32_and8992_y0;
  wire h_u_cla32_and8993_y0;
  wire h_u_cla32_and8994_y0;
  wire h_u_cla32_and8995_y0;
  wire h_u_cla32_and8996_y0;
  wire h_u_cla32_and8997_y0;
  wire h_u_cla32_and8998_y0;
  wire h_u_cla32_and8999_y0;
  wire h_u_cla32_and9000_y0;
  wire h_u_cla32_and9001_y0;
  wire h_u_cla32_and9002_y0;
  wire h_u_cla32_and9003_y0;
  wire h_u_cla32_and9004_y0;
  wire h_u_cla32_and9005_y0;
  wire h_u_cla32_and9006_y0;
  wire h_u_cla32_and9007_y0;
  wire h_u_cla32_and9008_y0;
  wire h_u_cla32_and9009_y0;
  wire h_u_cla32_and9010_y0;
  wire h_u_cla32_and9011_y0;
  wire h_u_cla32_and9012_y0;
  wire h_u_cla32_and9013_y0;
  wire h_u_cla32_and9014_y0;
  wire h_u_cla32_and9015_y0;
  wire h_u_cla32_and9016_y0;
  wire h_u_cla32_and9017_y0;
  wire h_u_cla32_and9018_y0;
  wire h_u_cla32_and9019_y0;
  wire h_u_cla32_and9020_y0;
  wire h_u_cla32_and9021_y0;
  wire h_u_cla32_and9022_y0;
  wire h_u_cla32_and9023_y0;
  wire h_u_cla32_and9024_y0;
  wire h_u_cla32_and9025_y0;
  wire h_u_cla32_and9026_y0;
  wire h_u_cla32_and9027_y0;
  wire h_u_cla32_and9028_y0;
  wire h_u_cla32_and9029_y0;
  wire h_u_cla32_and9030_y0;
  wire h_u_cla32_and9031_y0;
  wire h_u_cla32_and9032_y0;
  wire h_u_cla32_and9033_y0;
  wire h_u_cla32_and9034_y0;
  wire h_u_cla32_and9035_y0;
  wire h_u_cla32_and9036_y0;
  wire h_u_cla32_and9037_y0;
  wire h_u_cla32_and9038_y0;
  wire h_u_cla32_and9039_y0;
  wire h_u_cla32_and9040_y0;
  wire h_u_cla32_and9041_y0;
  wire h_u_cla32_and9042_y0;
  wire h_u_cla32_and9043_y0;
  wire h_u_cla32_and9044_y0;
  wire h_u_cla32_and9045_y0;
  wire h_u_cla32_and9046_y0;
  wire h_u_cla32_and9047_y0;
  wire h_u_cla32_and9048_y0;
  wire h_u_cla32_and9049_y0;
  wire h_u_cla32_and9050_y0;
  wire h_u_cla32_and9051_y0;
  wire h_u_cla32_and9052_y0;
  wire h_u_cla32_and9053_y0;
  wire h_u_cla32_and9054_y0;
  wire h_u_cla32_and9055_y0;
  wire h_u_cla32_and9056_y0;
  wire h_u_cla32_and9057_y0;
  wire h_u_cla32_and9058_y0;
  wire h_u_cla32_and9059_y0;
  wire h_u_cla32_and9060_y0;
  wire h_u_cla32_and9061_y0;
  wire h_u_cla32_and9062_y0;
  wire h_u_cla32_and9063_y0;
  wire h_u_cla32_and9064_y0;
  wire h_u_cla32_and9065_y0;
  wire h_u_cla32_and9066_y0;
  wire h_u_cla32_and9067_y0;
  wire h_u_cla32_and9068_y0;
  wire h_u_cla32_and9069_y0;
  wire h_u_cla32_and9070_y0;
  wire h_u_cla32_and9071_y0;
  wire h_u_cla32_and9072_y0;
  wire h_u_cla32_and9073_y0;
  wire h_u_cla32_and9074_y0;
  wire h_u_cla32_and9075_y0;
  wire h_u_cla32_and9076_y0;
  wire h_u_cla32_and9077_y0;
  wire h_u_cla32_and9078_y0;
  wire h_u_cla32_and9079_y0;
  wire h_u_cla32_and9080_y0;
  wire h_u_cla32_and9081_y0;
  wire h_u_cla32_and9082_y0;
  wire h_u_cla32_and9083_y0;
  wire h_u_cla32_and9084_y0;
  wire h_u_cla32_and9085_y0;
  wire h_u_cla32_and9086_y0;
  wire h_u_cla32_and9087_y0;
  wire h_u_cla32_and9088_y0;
  wire h_u_cla32_and9089_y0;
  wire h_u_cla32_and9090_y0;
  wire h_u_cla32_and9091_y0;
  wire h_u_cla32_and9092_y0;
  wire h_u_cla32_and9093_y0;
  wire h_u_cla32_and9094_y0;
  wire h_u_cla32_and9095_y0;
  wire h_u_cla32_and9096_y0;
  wire h_u_cla32_and9097_y0;
  wire h_u_cla32_and9098_y0;
  wire h_u_cla32_and9099_y0;
  wire h_u_cla32_and9100_y0;
  wire h_u_cla32_and9101_y0;
  wire h_u_cla32_and9102_y0;
  wire h_u_cla32_and9103_y0;
  wire h_u_cla32_and9104_y0;
  wire h_u_cla32_and9105_y0;
  wire h_u_cla32_and9106_y0;
  wire h_u_cla32_and9107_y0;
  wire h_u_cla32_and9108_y0;
  wire h_u_cla32_and9109_y0;
  wire h_u_cla32_and9110_y0;
  wire h_u_cla32_and9111_y0;
  wire h_u_cla32_and9112_y0;
  wire h_u_cla32_and9113_y0;
  wire h_u_cla32_and9114_y0;
  wire h_u_cla32_and9115_y0;
  wire h_u_cla32_and9116_y0;
  wire h_u_cla32_and9117_y0;
  wire h_u_cla32_and9118_y0;
  wire h_u_cla32_and9119_y0;
  wire h_u_cla32_and9120_y0;
  wire h_u_cla32_and9121_y0;
  wire h_u_cla32_and9122_y0;
  wire h_u_cla32_and9123_y0;
  wire h_u_cla32_and9124_y0;
  wire h_u_cla32_and9125_y0;
  wire h_u_cla32_and9126_y0;
  wire h_u_cla32_and9127_y0;
  wire h_u_cla32_and9128_y0;
  wire h_u_cla32_and9129_y0;
  wire h_u_cla32_and9130_y0;
  wire h_u_cla32_and9131_y0;
  wire h_u_cla32_and9132_y0;
  wire h_u_cla32_and9133_y0;
  wire h_u_cla32_and9134_y0;
  wire h_u_cla32_and9135_y0;
  wire h_u_cla32_and9136_y0;
  wire h_u_cla32_and9137_y0;
  wire h_u_cla32_and9138_y0;
  wire h_u_cla32_and9139_y0;
  wire h_u_cla32_and9140_y0;
  wire h_u_cla32_and9141_y0;
  wire h_u_cla32_and9142_y0;
  wire h_u_cla32_and9143_y0;
  wire h_u_cla32_and9144_y0;
  wire h_u_cla32_and9145_y0;
  wire h_u_cla32_and9146_y0;
  wire h_u_cla32_and9147_y0;
  wire h_u_cla32_and9148_y0;
  wire h_u_cla32_and9149_y0;
  wire h_u_cla32_and9150_y0;
  wire h_u_cla32_and9151_y0;
  wire h_u_cla32_and9152_y0;
  wire h_u_cla32_and9153_y0;
  wire h_u_cla32_and9154_y0;
  wire h_u_cla32_and9155_y0;
  wire h_u_cla32_and9156_y0;
  wire h_u_cla32_and9157_y0;
  wire h_u_cla32_and9158_y0;
  wire h_u_cla32_and9159_y0;
  wire h_u_cla32_and9160_y0;
  wire h_u_cla32_and9161_y0;
  wire h_u_cla32_and9162_y0;
  wire h_u_cla32_and9163_y0;
  wire h_u_cla32_and9164_y0;
  wire h_u_cla32_and9165_y0;
  wire h_u_cla32_and9166_y0;
  wire h_u_cla32_and9167_y0;
  wire h_u_cla32_and9168_y0;
  wire h_u_cla32_and9169_y0;
  wire h_u_cla32_and9170_y0;
  wire h_u_cla32_and9171_y0;
  wire h_u_cla32_and9172_y0;
  wire h_u_cla32_and9173_y0;
  wire h_u_cla32_and9174_y0;
  wire h_u_cla32_and9175_y0;
  wire h_u_cla32_and9176_y0;
  wire h_u_cla32_and9177_y0;
  wire h_u_cla32_and9178_y0;
  wire h_u_cla32_and9179_y0;
  wire h_u_cla32_and9180_y0;
  wire h_u_cla32_and9181_y0;
  wire h_u_cla32_and9182_y0;
  wire h_u_cla32_and9183_y0;
  wire h_u_cla32_and9184_y0;
  wire h_u_cla32_and9185_y0;
  wire h_u_cla32_and9186_y0;
  wire h_u_cla32_and9187_y0;
  wire h_u_cla32_and9188_y0;
  wire h_u_cla32_and9189_y0;
  wire h_u_cla32_and9190_y0;
  wire h_u_cla32_and9191_y0;
  wire h_u_cla32_and9192_y0;
  wire h_u_cla32_and9193_y0;
  wire h_u_cla32_and9194_y0;
  wire h_u_cla32_and9195_y0;
  wire h_u_cla32_and9196_y0;
  wire h_u_cla32_and9197_y0;
  wire h_u_cla32_and9198_y0;
  wire h_u_cla32_and9199_y0;
  wire h_u_cla32_and9200_y0;
  wire h_u_cla32_and9201_y0;
  wire h_u_cla32_and9202_y0;
  wire h_u_cla32_and9203_y0;
  wire h_u_cla32_and9204_y0;
  wire h_u_cla32_and9205_y0;
  wire h_u_cla32_and9206_y0;
  wire h_u_cla32_and9207_y0;
  wire h_u_cla32_and9208_y0;
  wire h_u_cla32_and9209_y0;
  wire h_u_cla32_and9210_y0;
  wire h_u_cla32_and9211_y0;
  wire h_u_cla32_and9212_y0;
  wire h_u_cla32_and9213_y0;
  wire h_u_cla32_and9214_y0;
  wire h_u_cla32_and9215_y0;
  wire h_u_cla32_and9216_y0;
  wire h_u_cla32_and9217_y0;
  wire h_u_cla32_and9218_y0;
  wire h_u_cla32_and9219_y0;
  wire h_u_cla32_and9220_y0;
  wire h_u_cla32_and9221_y0;
  wire h_u_cla32_and9222_y0;
  wire h_u_cla32_and9223_y0;
  wire h_u_cla32_and9224_y0;
  wire h_u_cla32_and9225_y0;
  wire h_u_cla32_and9226_y0;
  wire h_u_cla32_and9227_y0;
  wire h_u_cla32_and9228_y0;
  wire h_u_cla32_and9229_y0;
  wire h_u_cla32_and9230_y0;
  wire h_u_cla32_and9231_y0;
  wire h_u_cla32_and9232_y0;
  wire h_u_cla32_and9233_y0;
  wire h_u_cla32_and9234_y0;
  wire h_u_cla32_and9235_y0;
  wire h_u_cla32_and9236_y0;
  wire h_u_cla32_and9237_y0;
  wire h_u_cla32_and9238_y0;
  wire h_u_cla32_and9239_y0;
  wire h_u_cla32_and9240_y0;
  wire h_u_cla32_and9241_y0;
  wire h_u_cla32_and9242_y0;
  wire h_u_cla32_and9243_y0;
  wire h_u_cla32_and9244_y0;
  wire h_u_cla32_and9245_y0;
  wire h_u_cla32_and9246_y0;
  wire h_u_cla32_and9247_y0;
  wire h_u_cla32_and9248_y0;
  wire h_u_cla32_and9249_y0;
  wire h_u_cla32_and9250_y0;
  wire h_u_cla32_and9251_y0;
  wire h_u_cla32_and9252_y0;
  wire h_u_cla32_and9253_y0;
  wire h_u_cla32_and9254_y0;
  wire h_u_cla32_and9255_y0;
  wire h_u_cla32_and9256_y0;
  wire h_u_cla32_and9257_y0;
  wire h_u_cla32_and9258_y0;
  wire h_u_cla32_and9259_y0;
  wire h_u_cla32_and9260_y0;
  wire h_u_cla32_and9261_y0;
  wire h_u_cla32_and9262_y0;
  wire h_u_cla32_and9263_y0;
  wire h_u_cla32_and9264_y0;
  wire h_u_cla32_and9265_y0;
  wire h_u_cla32_and9266_y0;
  wire h_u_cla32_and9267_y0;
  wire h_u_cla32_and9268_y0;
  wire h_u_cla32_and9269_y0;
  wire h_u_cla32_and9270_y0;
  wire h_u_cla32_and9271_y0;
  wire h_u_cla32_and9272_y0;
  wire h_u_cla32_and9273_y0;
  wire h_u_cla32_and9274_y0;
  wire h_u_cla32_and9275_y0;
  wire h_u_cla32_and9276_y0;
  wire h_u_cla32_and9277_y0;
  wire h_u_cla32_and9278_y0;
  wire h_u_cla32_and9279_y0;
  wire h_u_cla32_and9280_y0;
  wire h_u_cla32_and9281_y0;
  wire h_u_cla32_and9282_y0;
  wire h_u_cla32_and9283_y0;
  wire h_u_cla32_and9284_y0;
  wire h_u_cla32_and9285_y0;
  wire h_u_cla32_and9286_y0;
  wire h_u_cla32_and9287_y0;
  wire h_u_cla32_and9288_y0;
  wire h_u_cla32_and9289_y0;
  wire h_u_cla32_and9290_y0;
  wire h_u_cla32_and9291_y0;
  wire h_u_cla32_and9292_y0;
  wire h_u_cla32_and9293_y0;
  wire h_u_cla32_and9294_y0;
  wire h_u_cla32_and9295_y0;
  wire h_u_cla32_and9296_y0;
  wire h_u_cla32_and9297_y0;
  wire h_u_cla32_and9298_y0;
  wire h_u_cla32_and9299_y0;
  wire h_u_cla32_and9300_y0;
  wire h_u_cla32_and9301_y0;
  wire h_u_cla32_and9302_y0;
  wire h_u_cla32_and9303_y0;
  wire h_u_cla32_and9304_y0;
  wire h_u_cla32_and9305_y0;
  wire h_u_cla32_and9306_y0;
  wire h_u_cla32_and9307_y0;
  wire h_u_cla32_and9308_y0;
  wire h_u_cla32_and9309_y0;
  wire h_u_cla32_and9310_y0;
  wire h_u_cla32_and9311_y0;
  wire h_u_cla32_and9312_y0;
  wire h_u_cla32_and9313_y0;
  wire h_u_cla32_and9314_y0;
  wire h_u_cla32_and9315_y0;
  wire h_u_cla32_and9316_y0;
  wire h_u_cla32_and9317_y0;
  wire h_u_cla32_and9318_y0;
  wire h_u_cla32_and9319_y0;
  wire h_u_cla32_and9320_y0;
  wire h_u_cla32_and9321_y0;
  wire h_u_cla32_and9322_y0;
  wire h_u_cla32_and9323_y0;
  wire h_u_cla32_and9324_y0;
  wire h_u_cla32_and9325_y0;
  wire h_u_cla32_and9326_y0;
  wire h_u_cla32_and9327_y0;
  wire h_u_cla32_and9328_y0;
  wire h_u_cla32_and9329_y0;
  wire h_u_cla32_and9330_y0;
  wire h_u_cla32_and9331_y0;
  wire h_u_cla32_and9332_y0;
  wire h_u_cla32_and9333_y0;
  wire h_u_cla32_and9334_y0;
  wire h_u_cla32_and9335_y0;
  wire h_u_cla32_and9336_y0;
  wire h_u_cla32_and9337_y0;
  wire h_u_cla32_and9338_y0;
  wire h_u_cla32_and9339_y0;
  wire h_u_cla32_and9340_y0;
  wire h_u_cla32_and9341_y0;
  wire h_u_cla32_and9342_y0;
  wire h_u_cla32_and9343_y0;
  wire h_u_cla32_and9344_y0;
  wire h_u_cla32_and9345_y0;
  wire h_u_cla32_and9346_y0;
  wire h_u_cla32_and9347_y0;
  wire h_u_cla32_and9348_y0;
  wire h_u_cla32_and9349_y0;
  wire h_u_cla32_and9350_y0;
  wire h_u_cla32_and9351_y0;
  wire h_u_cla32_and9352_y0;
  wire h_u_cla32_and9353_y0;
  wire h_u_cla32_and9354_y0;
  wire h_u_cla32_and9355_y0;
  wire h_u_cla32_and9356_y0;
  wire h_u_cla32_and9357_y0;
  wire h_u_cla32_and9358_y0;
  wire h_u_cla32_and9359_y0;
  wire h_u_cla32_and9360_y0;
  wire h_u_cla32_and9361_y0;
  wire h_u_cla32_and9362_y0;
  wire h_u_cla32_and9363_y0;
  wire h_u_cla32_and9364_y0;
  wire h_u_cla32_and9365_y0;
  wire h_u_cla32_and9366_y0;
  wire h_u_cla32_and9367_y0;
  wire h_u_cla32_and9368_y0;
  wire h_u_cla32_and9369_y0;
  wire h_u_cla32_and9370_y0;
  wire h_u_cla32_and9371_y0;
  wire h_u_cla32_and9372_y0;
  wire h_u_cla32_and9373_y0;
  wire h_u_cla32_and9374_y0;
  wire h_u_cla32_and9375_y0;
  wire h_u_cla32_and9376_y0;
  wire h_u_cla32_and9377_y0;
  wire h_u_cla32_and9378_y0;
  wire h_u_cla32_and9379_y0;
  wire h_u_cla32_and9380_y0;
  wire h_u_cla32_and9381_y0;
  wire h_u_cla32_and9382_y0;
  wire h_u_cla32_and9383_y0;
  wire h_u_cla32_and9384_y0;
  wire h_u_cla32_and9385_y0;
  wire h_u_cla32_and9386_y0;
  wire h_u_cla32_and9387_y0;
  wire h_u_cla32_and9388_y0;
  wire h_u_cla32_and9389_y0;
  wire h_u_cla32_and9390_y0;
  wire h_u_cla32_and9391_y0;
  wire h_u_cla32_and9392_y0;
  wire h_u_cla32_and9393_y0;
  wire h_u_cla32_and9394_y0;
  wire h_u_cla32_and9395_y0;
  wire h_u_cla32_and9396_y0;
  wire h_u_cla32_and9397_y0;
  wire h_u_cla32_and9398_y0;
  wire h_u_cla32_and9399_y0;
  wire h_u_cla32_and9400_y0;
  wire h_u_cla32_and9401_y0;
  wire h_u_cla32_and9402_y0;
  wire h_u_cla32_and9403_y0;
  wire h_u_cla32_and9404_y0;
  wire h_u_cla32_and9405_y0;
  wire h_u_cla32_and9406_y0;
  wire h_u_cla32_and9407_y0;
  wire h_u_cla32_and9408_y0;
  wire h_u_cla32_and9409_y0;
  wire h_u_cla32_and9410_y0;
  wire h_u_cla32_and9411_y0;
  wire h_u_cla32_and9412_y0;
  wire h_u_cla32_and9413_y0;
  wire h_u_cla32_and9414_y0;
  wire h_u_cla32_and9415_y0;
  wire h_u_cla32_and9416_y0;
  wire h_u_cla32_and9417_y0;
  wire h_u_cla32_and9418_y0;
  wire h_u_cla32_and9419_y0;
  wire h_u_cla32_and9420_y0;
  wire h_u_cla32_and9421_y0;
  wire h_u_cla32_and9422_y0;
  wire h_u_cla32_and9423_y0;
  wire h_u_cla32_and9424_y0;
  wire h_u_cla32_and9425_y0;
  wire h_u_cla32_and9426_y0;
  wire h_u_cla32_and9427_y0;
  wire h_u_cla32_and9428_y0;
  wire h_u_cla32_and9429_y0;
  wire h_u_cla32_and9430_y0;
  wire h_u_cla32_and9431_y0;
  wire h_u_cla32_and9432_y0;
  wire h_u_cla32_and9433_y0;
  wire h_u_cla32_and9434_y0;
  wire h_u_cla32_and9435_y0;
  wire h_u_cla32_and9436_y0;
  wire h_u_cla32_and9437_y0;
  wire h_u_cla32_and9438_y0;
  wire h_u_cla32_and9439_y0;
  wire h_u_cla32_and9440_y0;
  wire h_u_cla32_and9441_y0;
  wire h_u_cla32_and9442_y0;
  wire h_u_cla32_and9443_y0;
  wire h_u_cla32_and9444_y0;
  wire h_u_cla32_and9445_y0;
  wire h_u_cla32_and9446_y0;
  wire h_u_cla32_and9447_y0;
  wire h_u_cla32_and9448_y0;
  wire h_u_cla32_and9449_y0;
  wire h_u_cla32_and9450_y0;
  wire h_u_cla32_and9451_y0;
  wire h_u_cla32_and9452_y0;
  wire h_u_cla32_and9453_y0;
  wire h_u_cla32_and9454_y0;
  wire h_u_cla32_or435_y0;
  wire h_u_cla32_or436_y0;
  wire h_u_cla32_or437_y0;
  wire h_u_cla32_or438_y0;
  wire h_u_cla32_or439_y0;
  wire h_u_cla32_or440_y0;
  wire h_u_cla32_or441_y0;
  wire h_u_cla32_or442_y0;
  wire h_u_cla32_or443_y0;
  wire h_u_cla32_or444_y0;
  wire h_u_cla32_or445_y0;
  wire h_u_cla32_or446_y0;
  wire h_u_cla32_or447_y0;
  wire h_u_cla32_or448_y0;
  wire h_u_cla32_or449_y0;
  wire h_u_cla32_or450_y0;
  wire h_u_cla32_or451_y0;
  wire h_u_cla32_or452_y0;
  wire h_u_cla32_or453_y0;
  wire h_u_cla32_or454_y0;
  wire h_u_cla32_or455_y0;
  wire h_u_cla32_or456_y0;
  wire h_u_cla32_or457_y0;
  wire h_u_cla32_or458_y0;
  wire h_u_cla32_or459_y0;
  wire h_u_cla32_or460_y0;
  wire h_u_cla32_or461_y0;
  wire h_u_cla32_or462_y0;
  wire h_u_cla32_or463_y0;
  wire h_u_cla32_or464_y0;
  wire h_u_cla32_pg_logic30_y0;
  wire h_u_cla32_pg_logic30_y1;
  wire h_u_cla32_pg_logic30_y2;
  wire h_u_cla32_xor30_y0;
  wire h_u_cla32_and9455_y0;
  wire h_u_cla32_and9456_y0;
  wire h_u_cla32_and9457_y0;
  wire h_u_cla32_and9458_y0;
  wire h_u_cla32_and9459_y0;
  wire h_u_cla32_and9460_y0;
  wire h_u_cla32_and9461_y0;
  wire h_u_cla32_and9462_y0;
  wire h_u_cla32_and9463_y0;
  wire h_u_cla32_and9464_y0;
  wire h_u_cla32_and9465_y0;
  wire h_u_cla32_and9466_y0;
  wire h_u_cla32_and9467_y0;
  wire h_u_cla32_and9468_y0;
  wire h_u_cla32_and9469_y0;
  wire h_u_cla32_and9470_y0;
  wire h_u_cla32_and9471_y0;
  wire h_u_cla32_and9472_y0;
  wire h_u_cla32_and9473_y0;
  wire h_u_cla32_and9474_y0;
  wire h_u_cla32_and9475_y0;
  wire h_u_cla32_and9476_y0;
  wire h_u_cla32_and9477_y0;
  wire h_u_cla32_and9478_y0;
  wire h_u_cla32_and9479_y0;
  wire h_u_cla32_and9480_y0;
  wire h_u_cla32_and9481_y0;
  wire h_u_cla32_and9482_y0;
  wire h_u_cla32_and9483_y0;
  wire h_u_cla32_and9484_y0;
  wire h_u_cla32_and9485_y0;
  wire h_u_cla32_and9486_y0;
  wire h_u_cla32_and9487_y0;
  wire h_u_cla32_and9488_y0;
  wire h_u_cla32_and9489_y0;
  wire h_u_cla32_and9490_y0;
  wire h_u_cla32_and9491_y0;
  wire h_u_cla32_and9492_y0;
  wire h_u_cla32_and9493_y0;
  wire h_u_cla32_and9494_y0;
  wire h_u_cla32_and9495_y0;
  wire h_u_cla32_and9496_y0;
  wire h_u_cla32_and9497_y0;
  wire h_u_cla32_and9498_y0;
  wire h_u_cla32_and9499_y0;
  wire h_u_cla32_and9500_y0;
  wire h_u_cla32_and9501_y0;
  wire h_u_cla32_and9502_y0;
  wire h_u_cla32_and9503_y0;
  wire h_u_cla32_and9504_y0;
  wire h_u_cla32_and9505_y0;
  wire h_u_cla32_and9506_y0;
  wire h_u_cla32_and9507_y0;
  wire h_u_cla32_and9508_y0;
  wire h_u_cla32_and9509_y0;
  wire h_u_cla32_and9510_y0;
  wire h_u_cla32_and9511_y0;
  wire h_u_cla32_and9512_y0;
  wire h_u_cla32_and9513_y0;
  wire h_u_cla32_and9514_y0;
  wire h_u_cla32_and9515_y0;
  wire h_u_cla32_and9516_y0;
  wire h_u_cla32_and9517_y0;
  wire h_u_cla32_and9518_y0;
  wire h_u_cla32_and9519_y0;
  wire h_u_cla32_and9520_y0;
  wire h_u_cla32_and9521_y0;
  wire h_u_cla32_and9522_y0;
  wire h_u_cla32_and9523_y0;
  wire h_u_cla32_and9524_y0;
  wire h_u_cla32_and9525_y0;
  wire h_u_cla32_and9526_y0;
  wire h_u_cla32_and9527_y0;
  wire h_u_cla32_and9528_y0;
  wire h_u_cla32_and9529_y0;
  wire h_u_cla32_and9530_y0;
  wire h_u_cla32_and9531_y0;
  wire h_u_cla32_and9532_y0;
  wire h_u_cla32_and9533_y0;
  wire h_u_cla32_and9534_y0;
  wire h_u_cla32_and9535_y0;
  wire h_u_cla32_and9536_y0;
  wire h_u_cla32_and9537_y0;
  wire h_u_cla32_and9538_y0;
  wire h_u_cla32_and9539_y0;
  wire h_u_cla32_and9540_y0;
  wire h_u_cla32_and9541_y0;
  wire h_u_cla32_and9542_y0;
  wire h_u_cla32_and9543_y0;
  wire h_u_cla32_and9544_y0;
  wire h_u_cla32_and9545_y0;
  wire h_u_cla32_and9546_y0;
  wire h_u_cla32_and9547_y0;
  wire h_u_cla32_and9548_y0;
  wire h_u_cla32_and9549_y0;
  wire h_u_cla32_and9550_y0;
  wire h_u_cla32_and9551_y0;
  wire h_u_cla32_and9552_y0;
  wire h_u_cla32_and9553_y0;
  wire h_u_cla32_and9554_y0;
  wire h_u_cla32_and9555_y0;
  wire h_u_cla32_and9556_y0;
  wire h_u_cla32_and9557_y0;
  wire h_u_cla32_and9558_y0;
  wire h_u_cla32_and9559_y0;
  wire h_u_cla32_and9560_y0;
  wire h_u_cla32_and9561_y0;
  wire h_u_cla32_and9562_y0;
  wire h_u_cla32_and9563_y0;
  wire h_u_cla32_and9564_y0;
  wire h_u_cla32_and9565_y0;
  wire h_u_cla32_and9566_y0;
  wire h_u_cla32_and9567_y0;
  wire h_u_cla32_and9568_y0;
  wire h_u_cla32_and9569_y0;
  wire h_u_cla32_and9570_y0;
  wire h_u_cla32_and9571_y0;
  wire h_u_cla32_and9572_y0;
  wire h_u_cla32_and9573_y0;
  wire h_u_cla32_and9574_y0;
  wire h_u_cla32_and9575_y0;
  wire h_u_cla32_and9576_y0;
  wire h_u_cla32_and9577_y0;
  wire h_u_cla32_and9578_y0;
  wire h_u_cla32_and9579_y0;
  wire h_u_cla32_and9580_y0;
  wire h_u_cla32_and9581_y0;
  wire h_u_cla32_and9582_y0;
  wire h_u_cla32_and9583_y0;
  wire h_u_cla32_and9584_y0;
  wire h_u_cla32_and9585_y0;
  wire h_u_cla32_and9586_y0;
  wire h_u_cla32_and9587_y0;
  wire h_u_cla32_and9588_y0;
  wire h_u_cla32_and9589_y0;
  wire h_u_cla32_and9590_y0;
  wire h_u_cla32_and9591_y0;
  wire h_u_cla32_and9592_y0;
  wire h_u_cla32_and9593_y0;
  wire h_u_cla32_and9594_y0;
  wire h_u_cla32_and9595_y0;
  wire h_u_cla32_and9596_y0;
  wire h_u_cla32_and9597_y0;
  wire h_u_cla32_and9598_y0;
  wire h_u_cla32_and9599_y0;
  wire h_u_cla32_and9600_y0;
  wire h_u_cla32_and9601_y0;
  wire h_u_cla32_and9602_y0;
  wire h_u_cla32_and9603_y0;
  wire h_u_cla32_and9604_y0;
  wire h_u_cla32_and9605_y0;
  wire h_u_cla32_and9606_y0;
  wire h_u_cla32_and9607_y0;
  wire h_u_cla32_and9608_y0;
  wire h_u_cla32_and9609_y0;
  wire h_u_cla32_and9610_y0;
  wire h_u_cla32_and9611_y0;
  wire h_u_cla32_and9612_y0;
  wire h_u_cla32_and9613_y0;
  wire h_u_cla32_and9614_y0;
  wire h_u_cla32_and9615_y0;
  wire h_u_cla32_and9616_y0;
  wire h_u_cla32_and9617_y0;
  wire h_u_cla32_and9618_y0;
  wire h_u_cla32_and9619_y0;
  wire h_u_cla32_and9620_y0;
  wire h_u_cla32_and9621_y0;
  wire h_u_cla32_and9622_y0;
  wire h_u_cla32_and9623_y0;
  wire h_u_cla32_and9624_y0;
  wire h_u_cla32_and9625_y0;
  wire h_u_cla32_and9626_y0;
  wire h_u_cla32_and9627_y0;
  wire h_u_cla32_and9628_y0;
  wire h_u_cla32_and9629_y0;
  wire h_u_cla32_and9630_y0;
  wire h_u_cla32_and9631_y0;
  wire h_u_cla32_and9632_y0;
  wire h_u_cla32_and9633_y0;
  wire h_u_cla32_and9634_y0;
  wire h_u_cla32_and9635_y0;
  wire h_u_cla32_and9636_y0;
  wire h_u_cla32_and9637_y0;
  wire h_u_cla32_and9638_y0;
  wire h_u_cla32_and9639_y0;
  wire h_u_cla32_and9640_y0;
  wire h_u_cla32_and9641_y0;
  wire h_u_cla32_and9642_y0;
  wire h_u_cla32_and9643_y0;
  wire h_u_cla32_and9644_y0;
  wire h_u_cla32_and9645_y0;
  wire h_u_cla32_and9646_y0;
  wire h_u_cla32_and9647_y0;
  wire h_u_cla32_and9648_y0;
  wire h_u_cla32_and9649_y0;
  wire h_u_cla32_and9650_y0;
  wire h_u_cla32_and9651_y0;
  wire h_u_cla32_and9652_y0;
  wire h_u_cla32_and9653_y0;
  wire h_u_cla32_and9654_y0;
  wire h_u_cla32_and9655_y0;
  wire h_u_cla32_and9656_y0;
  wire h_u_cla32_and9657_y0;
  wire h_u_cla32_and9658_y0;
  wire h_u_cla32_and9659_y0;
  wire h_u_cla32_and9660_y0;
  wire h_u_cla32_and9661_y0;
  wire h_u_cla32_and9662_y0;
  wire h_u_cla32_and9663_y0;
  wire h_u_cla32_and9664_y0;
  wire h_u_cla32_and9665_y0;
  wire h_u_cla32_and9666_y0;
  wire h_u_cla32_and9667_y0;
  wire h_u_cla32_and9668_y0;
  wire h_u_cla32_and9669_y0;
  wire h_u_cla32_and9670_y0;
  wire h_u_cla32_and9671_y0;
  wire h_u_cla32_and9672_y0;
  wire h_u_cla32_and9673_y0;
  wire h_u_cla32_and9674_y0;
  wire h_u_cla32_and9675_y0;
  wire h_u_cla32_and9676_y0;
  wire h_u_cla32_and9677_y0;
  wire h_u_cla32_and9678_y0;
  wire h_u_cla32_and9679_y0;
  wire h_u_cla32_and9680_y0;
  wire h_u_cla32_and9681_y0;
  wire h_u_cla32_and9682_y0;
  wire h_u_cla32_and9683_y0;
  wire h_u_cla32_and9684_y0;
  wire h_u_cla32_and9685_y0;
  wire h_u_cla32_and9686_y0;
  wire h_u_cla32_and9687_y0;
  wire h_u_cla32_and9688_y0;
  wire h_u_cla32_and9689_y0;
  wire h_u_cla32_and9690_y0;
  wire h_u_cla32_and9691_y0;
  wire h_u_cla32_and9692_y0;
  wire h_u_cla32_and9693_y0;
  wire h_u_cla32_and9694_y0;
  wire h_u_cla32_and9695_y0;
  wire h_u_cla32_and9696_y0;
  wire h_u_cla32_and9697_y0;
  wire h_u_cla32_and9698_y0;
  wire h_u_cla32_and9699_y0;
  wire h_u_cla32_and9700_y0;
  wire h_u_cla32_and9701_y0;
  wire h_u_cla32_and9702_y0;
  wire h_u_cla32_and9703_y0;
  wire h_u_cla32_and9704_y0;
  wire h_u_cla32_and9705_y0;
  wire h_u_cla32_and9706_y0;
  wire h_u_cla32_and9707_y0;
  wire h_u_cla32_and9708_y0;
  wire h_u_cla32_and9709_y0;
  wire h_u_cla32_and9710_y0;
  wire h_u_cla32_and9711_y0;
  wire h_u_cla32_and9712_y0;
  wire h_u_cla32_and9713_y0;
  wire h_u_cla32_and9714_y0;
  wire h_u_cla32_and9715_y0;
  wire h_u_cla32_and9716_y0;
  wire h_u_cla32_and9717_y0;
  wire h_u_cla32_and9718_y0;
  wire h_u_cla32_and9719_y0;
  wire h_u_cla32_and9720_y0;
  wire h_u_cla32_and9721_y0;
  wire h_u_cla32_and9722_y0;
  wire h_u_cla32_and9723_y0;
  wire h_u_cla32_and9724_y0;
  wire h_u_cla32_and9725_y0;
  wire h_u_cla32_and9726_y0;
  wire h_u_cla32_and9727_y0;
  wire h_u_cla32_and9728_y0;
  wire h_u_cla32_and9729_y0;
  wire h_u_cla32_and9730_y0;
  wire h_u_cla32_and9731_y0;
  wire h_u_cla32_and9732_y0;
  wire h_u_cla32_and9733_y0;
  wire h_u_cla32_and9734_y0;
  wire h_u_cla32_and9735_y0;
  wire h_u_cla32_and9736_y0;
  wire h_u_cla32_and9737_y0;
  wire h_u_cla32_and9738_y0;
  wire h_u_cla32_and9739_y0;
  wire h_u_cla32_and9740_y0;
  wire h_u_cla32_and9741_y0;
  wire h_u_cla32_and9742_y0;
  wire h_u_cla32_and9743_y0;
  wire h_u_cla32_and9744_y0;
  wire h_u_cla32_and9745_y0;
  wire h_u_cla32_and9746_y0;
  wire h_u_cla32_and9747_y0;
  wire h_u_cla32_and9748_y0;
  wire h_u_cla32_and9749_y0;
  wire h_u_cla32_and9750_y0;
  wire h_u_cla32_and9751_y0;
  wire h_u_cla32_and9752_y0;
  wire h_u_cla32_and9753_y0;
  wire h_u_cla32_and9754_y0;
  wire h_u_cla32_and9755_y0;
  wire h_u_cla32_and9756_y0;
  wire h_u_cla32_and9757_y0;
  wire h_u_cla32_and9758_y0;
  wire h_u_cla32_and9759_y0;
  wire h_u_cla32_and9760_y0;
  wire h_u_cla32_and9761_y0;
  wire h_u_cla32_and9762_y0;
  wire h_u_cla32_and9763_y0;
  wire h_u_cla32_and9764_y0;
  wire h_u_cla32_and9765_y0;
  wire h_u_cla32_and9766_y0;
  wire h_u_cla32_and9767_y0;
  wire h_u_cla32_and9768_y0;
  wire h_u_cla32_and9769_y0;
  wire h_u_cla32_and9770_y0;
  wire h_u_cla32_and9771_y0;
  wire h_u_cla32_and9772_y0;
  wire h_u_cla32_and9773_y0;
  wire h_u_cla32_and9774_y0;
  wire h_u_cla32_and9775_y0;
  wire h_u_cla32_and9776_y0;
  wire h_u_cla32_and9777_y0;
  wire h_u_cla32_and9778_y0;
  wire h_u_cla32_and9779_y0;
  wire h_u_cla32_and9780_y0;
  wire h_u_cla32_and9781_y0;
  wire h_u_cla32_and9782_y0;
  wire h_u_cla32_and9783_y0;
  wire h_u_cla32_and9784_y0;
  wire h_u_cla32_and9785_y0;
  wire h_u_cla32_and9786_y0;
  wire h_u_cla32_and9787_y0;
  wire h_u_cla32_and9788_y0;
  wire h_u_cla32_and9789_y0;
  wire h_u_cla32_and9790_y0;
  wire h_u_cla32_and9791_y0;
  wire h_u_cla32_and9792_y0;
  wire h_u_cla32_and9793_y0;
  wire h_u_cla32_and9794_y0;
  wire h_u_cla32_and9795_y0;
  wire h_u_cla32_and9796_y0;
  wire h_u_cla32_and9797_y0;
  wire h_u_cla32_and9798_y0;
  wire h_u_cla32_and9799_y0;
  wire h_u_cla32_and9800_y0;
  wire h_u_cla32_and9801_y0;
  wire h_u_cla32_and9802_y0;
  wire h_u_cla32_and9803_y0;
  wire h_u_cla32_and9804_y0;
  wire h_u_cla32_and9805_y0;
  wire h_u_cla32_and9806_y0;
  wire h_u_cla32_and9807_y0;
  wire h_u_cla32_and9808_y0;
  wire h_u_cla32_and9809_y0;
  wire h_u_cla32_and9810_y0;
  wire h_u_cla32_and9811_y0;
  wire h_u_cla32_and9812_y0;
  wire h_u_cla32_and9813_y0;
  wire h_u_cla32_and9814_y0;
  wire h_u_cla32_and9815_y0;
  wire h_u_cla32_and9816_y0;
  wire h_u_cla32_and9817_y0;
  wire h_u_cla32_and9818_y0;
  wire h_u_cla32_and9819_y0;
  wire h_u_cla32_and9820_y0;
  wire h_u_cla32_and9821_y0;
  wire h_u_cla32_and9822_y0;
  wire h_u_cla32_and9823_y0;
  wire h_u_cla32_and9824_y0;
  wire h_u_cla32_and9825_y0;
  wire h_u_cla32_and9826_y0;
  wire h_u_cla32_and9827_y0;
  wire h_u_cla32_and9828_y0;
  wire h_u_cla32_and9829_y0;
  wire h_u_cla32_and9830_y0;
  wire h_u_cla32_and9831_y0;
  wire h_u_cla32_and9832_y0;
  wire h_u_cla32_and9833_y0;
  wire h_u_cla32_and9834_y0;
  wire h_u_cla32_and9835_y0;
  wire h_u_cla32_and9836_y0;
  wire h_u_cla32_and9837_y0;
  wire h_u_cla32_and9838_y0;
  wire h_u_cla32_and9839_y0;
  wire h_u_cla32_and9840_y0;
  wire h_u_cla32_and9841_y0;
  wire h_u_cla32_and9842_y0;
  wire h_u_cla32_and9843_y0;
  wire h_u_cla32_and9844_y0;
  wire h_u_cla32_and9845_y0;
  wire h_u_cla32_and9846_y0;
  wire h_u_cla32_and9847_y0;
  wire h_u_cla32_and9848_y0;
  wire h_u_cla32_and9849_y0;
  wire h_u_cla32_and9850_y0;
  wire h_u_cla32_and9851_y0;
  wire h_u_cla32_and9852_y0;
  wire h_u_cla32_and9853_y0;
  wire h_u_cla32_and9854_y0;
  wire h_u_cla32_and9855_y0;
  wire h_u_cla32_and9856_y0;
  wire h_u_cla32_and9857_y0;
  wire h_u_cla32_and9858_y0;
  wire h_u_cla32_and9859_y0;
  wire h_u_cla32_and9860_y0;
  wire h_u_cla32_and9861_y0;
  wire h_u_cla32_and9862_y0;
  wire h_u_cla32_and9863_y0;
  wire h_u_cla32_and9864_y0;
  wire h_u_cla32_and9865_y0;
  wire h_u_cla32_and9866_y0;
  wire h_u_cla32_and9867_y0;
  wire h_u_cla32_and9868_y0;
  wire h_u_cla32_and9869_y0;
  wire h_u_cla32_and9870_y0;
  wire h_u_cla32_and9871_y0;
  wire h_u_cla32_and9872_y0;
  wire h_u_cla32_and9873_y0;
  wire h_u_cla32_and9874_y0;
  wire h_u_cla32_and9875_y0;
  wire h_u_cla32_and9876_y0;
  wire h_u_cla32_and9877_y0;
  wire h_u_cla32_and9878_y0;
  wire h_u_cla32_and9879_y0;
  wire h_u_cla32_and9880_y0;
  wire h_u_cla32_and9881_y0;
  wire h_u_cla32_and9882_y0;
  wire h_u_cla32_and9883_y0;
  wire h_u_cla32_and9884_y0;
  wire h_u_cla32_and9885_y0;
  wire h_u_cla32_and9886_y0;
  wire h_u_cla32_and9887_y0;
  wire h_u_cla32_and9888_y0;
  wire h_u_cla32_and9889_y0;
  wire h_u_cla32_and9890_y0;
  wire h_u_cla32_and9891_y0;
  wire h_u_cla32_and9892_y0;
  wire h_u_cla32_and9893_y0;
  wire h_u_cla32_and9894_y0;
  wire h_u_cla32_and9895_y0;
  wire h_u_cla32_and9896_y0;
  wire h_u_cla32_and9897_y0;
  wire h_u_cla32_and9898_y0;
  wire h_u_cla32_and9899_y0;
  wire h_u_cla32_and9900_y0;
  wire h_u_cla32_and9901_y0;
  wire h_u_cla32_and9902_y0;
  wire h_u_cla32_and9903_y0;
  wire h_u_cla32_and9904_y0;
  wire h_u_cla32_and9905_y0;
  wire h_u_cla32_and9906_y0;
  wire h_u_cla32_and9907_y0;
  wire h_u_cla32_and9908_y0;
  wire h_u_cla32_and9909_y0;
  wire h_u_cla32_and9910_y0;
  wire h_u_cla32_and9911_y0;
  wire h_u_cla32_and9912_y0;
  wire h_u_cla32_and9913_y0;
  wire h_u_cla32_and9914_y0;
  wire h_u_cla32_and9915_y0;
  wire h_u_cla32_and9916_y0;
  wire h_u_cla32_and9917_y0;
  wire h_u_cla32_and9918_y0;
  wire h_u_cla32_and9919_y0;
  wire h_u_cla32_and9920_y0;
  wire h_u_cla32_and9921_y0;
  wire h_u_cla32_and9922_y0;
  wire h_u_cla32_and9923_y0;
  wire h_u_cla32_and9924_y0;
  wire h_u_cla32_and9925_y0;
  wire h_u_cla32_and9926_y0;
  wire h_u_cla32_and9927_y0;
  wire h_u_cla32_and9928_y0;
  wire h_u_cla32_and9929_y0;
  wire h_u_cla32_and9930_y0;
  wire h_u_cla32_and9931_y0;
  wire h_u_cla32_and9932_y0;
  wire h_u_cla32_and9933_y0;
  wire h_u_cla32_and9934_y0;
  wire h_u_cla32_and9935_y0;
  wire h_u_cla32_and9936_y0;
  wire h_u_cla32_and9937_y0;
  wire h_u_cla32_and9938_y0;
  wire h_u_cla32_and9939_y0;
  wire h_u_cla32_and9940_y0;
  wire h_u_cla32_and9941_y0;
  wire h_u_cla32_and9942_y0;
  wire h_u_cla32_and9943_y0;
  wire h_u_cla32_and9944_y0;
  wire h_u_cla32_and9945_y0;
  wire h_u_cla32_and9946_y0;
  wire h_u_cla32_and9947_y0;
  wire h_u_cla32_and9948_y0;
  wire h_u_cla32_and9949_y0;
  wire h_u_cla32_and9950_y0;
  wire h_u_cla32_and9951_y0;
  wire h_u_cla32_and9952_y0;
  wire h_u_cla32_and9953_y0;
  wire h_u_cla32_and9954_y0;
  wire h_u_cla32_and9955_y0;
  wire h_u_cla32_and9956_y0;
  wire h_u_cla32_and9957_y0;
  wire h_u_cla32_and9958_y0;
  wire h_u_cla32_and9959_y0;
  wire h_u_cla32_and9960_y0;
  wire h_u_cla32_and9961_y0;
  wire h_u_cla32_and9962_y0;
  wire h_u_cla32_and9963_y0;
  wire h_u_cla32_and9964_y0;
  wire h_u_cla32_and9965_y0;
  wire h_u_cla32_and9966_y0;
  wire h_u_cla32_and9967_y0;
  wire h_u_cla32_and9968_y0;
  wire h_u_cla32_and9969_y0;
  wire h_u_cla32_and9970_y0;
  wire h_u_cla32_and9971_y0;
  wire h_u_cla32_and9972_y0;
  wire h_u_cla32_and9973_y0;
  wire h_u_cla32_and9974_y0;
  wire h_u_cla32_and9975_y0;
  wire h_u_cla32_and9976_y0;
  wire h_u_cla32_and9977_y0;
  wire h_u_cla32_and9978_y0;
  wire h_u_cla32_and9979_y0;
  wire h_u_cla32_and9980_y0;
  wire h_u_cla32_and9981_y0;
  wire h_u_cla32_and9982_y0;
  wire h_u_cla32_and9983_y0;
  wire h_u_cla32_and9984_y0;
  wire h_u_cla32_and9985_y0;
  wire h_u_cla32_and9986_y0;
  wire h_u_cla32_and9987_y0;
  wire h_u_cla32_and9988_y0;
  wire h_u_cla32_and9989_y0;
  wire h_u_cla32_and9990_y0;
  wire h_u_cla32_and9991_y0;
  wire h_u_cla32_and9992_y0;
  wire h_u_cla32_and9993_y0;
  wire h_u_cla32_and9994_y0;
  wire h_u_cla32_and9995_y0;
  wire h_u_cla32_and9996_y0;
  wire h_u_cla32_and9997_y0;
  wire h_u_cla32_and9998_y0;
  wire h_u_cla32_and9999_y0;
  wire h_u_cla32_and10000_y0;
  wire h_u_cla32_and10001_y0;
  wire h_u_cla32_and10002_y0;
  wire h_u_cla32_and10003_y0;
  wire h_u_cla32_and10004_y0;
  wire h_u_cla32_and10005_y0;
  wire h_u_cla32_and10006_y0;
  wire h_u_cla32_and10007_y0;
  wire h_u_cla32_and10008_y0;
  wire h_u_cla32_and10009_y0;
  wire h_u_cla32_and10010_y0;
  wire h_u_cla32_and10011_y0;
  wire h_u_cla32_and10012_y0;
  wire h_u_cla32_and10013_y0;
  wire h_u_cla32_and10014_y0;
  wire h_u_cla32_and10015_y0;
  wire h_u_cla32_and10016_y0;
  wire h_u_cla32_and10017_y0;
  wire h_u_cla32_and10018_y0;
  wire h_u_cla32_and10019_y0;
  wire h_u_cla32_and10020_y0;
  wire h_u_cla32_and10021_y0;
  wire h_u_cla32_and10022_y0;
  wire h_u_cla32_and10023_y0;
  wire h_u_cla32_and10024_y0;
  wire h_u_cla32_and10025_y0;
  wire h_u_cla32_and10026_y0;
  wire h_u_cla32_and10027_y0;
  wire h_u_cla32_and10028_y0;
  wire h_u_cla32_and10029_y0;
  wire h_u_cla32_and10030_y0;
  wire h_u_cla32_and10031_y0;
  wire h_u_cla32_and10032_y0;
  wire h_u_cla32_and10033_y0;
  wire h_u_cla32_and10034_y0;
  wire h_u_cla32_and10035_y0;
  wire h_u_cla32_and10036_y0;
  wire h_u_cla32_and10037_y0;
  wire h_u_cla32_and10038_y0;
  wire h_u_cla32_and10039_y0;
  wire h_u_cla32_and10040_y0;
  wire h_u_cla32_and10041_y0;
  wire h_u_cla32_and10042_y0;
  wire h_u_cla32_and10043_y0;
  wire h_u_cla32_and10044_y0;
  wire h_u_cla32_and10045_y0;
  wire h_u_cla32_and10046_y0;
  wire h_u_cla32_and10047_y0;
  wire h_u_cla32_and10048_y0;
  wire h_u_cla32_and10049_y0;
  wire h_u_cla32_and10050_y0;
  wire h_u_cla32_and10051_y0;
  wire h_u_cla32_and10052_y0;
  wire h_u_cla32_and10053_y0;
  wire h_u_cla32_and10054_y0;
  wire h_u_cla32_and10055_y0;
  wire h_u_cla32_and10056_y0;
  wire h_u_cla32_and10057_y0;
  wire h_u_cla32_and10058_y0;
  wire h_u_cla32_and10059_y0;
  wire h_u_cla32_and10060_y0;
  wire h_u_cla32_and10061_y0;
  wire h_u_cla32_and10062_y0;
  wire h_u_cla32_and10063_y0;
  wire h_u_cla32_and10064_y0;
  wire h_u_cla32_and10065_y0;
  wire h_u_cla32_and10066_y0;
  wire h_u_cla32_and10067_y0;
  wire h_u_cla32_and10068_y0;
  wire h_u_cla32_and10069_y0;
  wire h_u_cla32_and10070_y0;
  wire h_u_cla32_and10071_y0;
  wire h_u_cla32_and10072_y0;
  wire h_u_cla32_and10073_y0;
  wire h_u_cla32_and10074_y0;
  wire h_u_cla32_and10075_y0;
  wire h_u_cla32_and10076_y0;
  wire h_u_cla32_and10077_y0;
  wire h_u_cla32_and10078_y0;
  wire h_u_cla32_and10079_y0;
  wire h_u_cla32_and10080_y0;
  wire h_u_cla32_and10081_y0;
  wire h_u_cla32_and10082_y0;
  wire h_u_cla32_and10083_y0;
  wire h_u_cla32_and10084_y0;
  wire h_u_cla32_and10085_y0;
  wire h_u_cla32_and10086_y0;
  wire h_u_cla32_and10087_y0;
  wire h_u_cla32_and10088_y0;
  wire h_u_cla32_and10089_y0;
  wire h_u_cla32_and10090_y0;
  wire h_u_cla32_and10091_y0;
  wire h_u_cla32_and10092_y0;
  wire h_u_cla32_and10093_y0;
  wire h_u_cla32_and10094_y0;
  wire h_u_cla32_and10095_y0;
  wire h_u_cla32_and10096_y0;
  wire h_u_cla32_and10097_y0;
  wire h_u_cla32_and10098_y0;
  wire h_u_cla32_and10099_y0;
  wire h_u_cla32_and10100_y0;
  wire h_u_cla32_and10101_y0;
  wire h_u_cla32_and10102_y0;
  wire h_u_cla32_and10103_y0;
  wire h_u_cla32_and10104_y0;
  wire h_u_cla32_and10105_y0;
  wire h_u_cla32_and10106_y0;
  wire h_u_cla32_and10107_y0;
  wire h_u_cla32_and10108_y0;
  wire h_u_cla32_and10109_y0;
  wire h_u_cla32_and10110_y0;
  wire h_u_cla32_and10111_y0;
  wire h_u_cla32_and10112_y0;
  wire h_u_cla32_and10113_y0;
  wire h_u_cla32_and10114_y0;
  wire h_u_cla32_and10115_y0;
  wire h_u_cla32_and10116_y0;
  wire h_u_cla32_and10117_y0;
  wire h_u_cla32_and10118_y0;
  wire h_u_cla32_and10119_y0;
  wire h_u_cla32_and10120_y0;
  wire h_u_cla32_and10121_y0;
  wire h_u_cla32_and10122_y0;
  wire h_u_cla32_and10123_y0;
  wire h_u_cla32_and10124_y0;
  wire h_u_cla32_and10125_y0;
  wire h_u_cla32_and10126_y0;
  wire h_u_cla32_and10127_y0;
  wire h_u_cla32_and10128_y0;
  wire h_u_cla32_and10129_y0;
  wire h_u_cla32_and10130_y0;
  wire h_u_cla32_and10131_y0;
  wire h_u_cla32_and10132_y0;
  wire h_u_cla32_and10133_y0;
  wire h_u_cla32_and10134_y0;
  wire h_u_cla32_and10135_y0;
  wire h_u_cla32_and10136_y0;
  wire h_u_cla32_and10137_y0;
  wire h_u_cla32_and10138_y0;
  wire h_u_cla32_and10139_y0;
  wire h_u_cla32_and10140_y0;
  wire h_u_cla32_and10141_y0;
  wire h_u_cla32_and10142_y0;
  wire h_u_cla32_and10143_y0;
  wire h_u_cla32_and10144_y0;
  wire h_u_cla32_and10145_y0;
  wire h_u_cla32_and10146_y0;
  wire h_u_cla32_and10147_y0;
  wire h_u_cla32_and10148_y0;
  wire h_u_cla32_and10149_y0;
  wire h_u_cla32_and10150_y0;
  wire h_u_cla32_and10151_y0;
  wire h_u_cla32_and10152_y0;
  wire h_u_cla32_and10153_y0;
  wire h_u_cla32_and10154_y0;
  wire h_u_cla32_and10155_y0;
  wire h_u_cla32_and10156_y0;
  wire h_u_cla32_and10157_y0;
  wire h_u_cla32_and10158_y0;
  wire h_u_cla32_and10159_y0;
  wire h_u_cla32_and10160_y0;
  wire h_u_cla32_and10161_y0;
  wire h_u_cla32_and10162_y0;
  wire h_u_cla32_and10163_y0;
  wire h_u_cla32_and10164_y0;
  wire h_u_cla32_and10165_y0;
  wire h_u_cla32_and10166_y0;
  wire h_u_cla32_and10167_y0;
  wire h_u_cla32_and10168_y0;
  wire h_u_cla32_and10169_y0;
  wire h_u_cla32_and10170_y0;
  wire h_u_cla32_and10171_y0;
  wire h_u_cla32_and10172_y0;
  wire h_u_cla32_and10173_y0;
  wire h_u_cla32_and10174_y0;
  wire h_u_cla32_and10175_y0;
  wire h_u_cla32_and10176_y0;
  wire h_u_cla32_and10177_y0;
  wire h_u_cla32_and10178_y0;
  wire h_u_cla32_and10179_y0;
  wire h_u_cla32_and10180_y0;
  wire h_u_cla32_and10181_y0;
  wire h_u_cla32_and10182_y0;
  wire h_u_cla32_and10183_y0;
  wire h_u_cla32_and10184_y0;
  wire h_u_cla32_and10185_y0;
  wire h_u_cla32_and10186_y0;
  wire h_u_cla32_and10187_y0;
  wire h_u_cla32_and10188_y0;
  wire h_u_cla32_and10189_y0;
  wire h_u_cla32_and10190_y0;
  wire h_u_cla32_and10191_y0;
  wire h_u_cla32_and10192_y0;
  wire h_u_cla32_and10193_y0;
  wire h_u_cla32_and10194_y0;
  wire h_u_cla32_and10195_y0;
  wire h_u_cla32_and10196_y0;
  wire h_u_cla32_and10197_y0;
  wire h_u_cla32_and10198_y0;
  wire h_u_cla32_and10199_y0;
  wire h_u_cla32_and10200_y0;
  wire h_u_cla32_and10201_y0;
  wire h_u_cla32_and10202_y0;
  wire h_u_cla32_and10203_y0;
  wire h_u_cla32_and10204_y0;
  wire h_u_cla32_and10205_y0;
  wire h_u_cla32_and10206_y0;
  wire h_u_cla32_and10207_y0;
  wire h_u_cla32_and10208_y0;
  wire h_u_cla32_and10209_y0;
  wire h_u_cla32_and10210_y0;
  wire h_u_cla32_and10211_y0;
  wire h_u_cla32_and10212_y0;
  wire h_u_cla32_and10213_y0;
  wire h_u_cla32_and10214_y0;
  wire h_u_cla32_and10215_y0;
  wire h_u_cla32_and10216_y0;
  wire h_u_cla32_and10217_y0;
  wire h_u_cla32_and10218_y0;
  wire h_u_cla32_and10219_y0;
  wire h_u_cla32_and10220_y0;
  wire h_u_cla32_and10221_y0;
  wire h_u_cla32_and10222_y0;
  wire h_u_cla32_and10223_y0;
  wire h_u_cla32_and10224_y0;
  wire h_u_cla32_and10225_y0;
  wire h_u_cla32_and10226_y0;
  wire h_u_cla32_and10227_y0;
  wire h_u_cla32_and10228_y0;
  wire h_u_cla32_and10229_y0;
  wire h_u_cla32_and10230_y0;
  wire h_u_cla32_and10231_y0;
  wire h_u_cla32_and10232_y0;
  wire h_u_cla32_and10233_y0;
  wire h_u_cla32_and10234_y0;
  wire h_u_cla32_and10235_y0;
  wire h_u_cla32_and10236_y0;
  wire h_u_cla32_and10237_y0;
  wire h_u_cla32_and10238_y0;
  wire h_u_cla32_and10239_y0;
  wire h_u_cla32_and10240_y0;
  wire h_u_cla32_and10241_y0;
  wire h_u_cla32_and10242_y0;
  wire h_u_cla32_and10243_y0;
  wire h_u_cla32_and10244_y0;
  wire h_u_cla32_and10245_y0;
  wire h_u_cla32_and10246_y0;
  wire h_u_cla32_and10247_y0;
  wire h_u_cla32_and10248_y0;
  wire h_u_cla32_and10249_y0;
  wire h_u_cla32_and10250_y0;
  wire h_u_cla32_and10251_y0;
  wire h_u_cla32_and10252_y0;
  wire h_u_cla32_and10253_y0;
  wire h_u_cla32_and10254_y0;
  wire h_u_cla32_and10255_y0;
  wire h_u_cla32_and10256_y0;
  wire h_u_cla32_and10257_y0;
  wire h_u_cla32_and10258_y0;
  wire h_u_cla32_and10259_y0;
  wire h_u_cla32_and10260_y0;
  wire h_u_cla32_and10261_y0;
  wire h_u_cla32_and10262_y0;
  wire h_u_cla32_and10263_y0;
  wire h_u_cla32_and10264_y0;
  wire h_u_cla32_and10265_y0;
  wire h_u_cla32_and10266_y0;
  wire h_u_cla32_and10267_y0;
  wire h_u_cla32_and10268_y0;
  wire h_u_cla32_and10269_y0;
  wire h_u_cla32_and10270_y0;
  wire h_u_cla32_and10271_y0;
  wire h_u_cla32_and10272_y0;
  wire h_u_cla32_and10273_y0;
  wire h_u_cla32_and10274_y0;
  wire h_u_cla32_and10275_y0;
  wire h_u_cla32_and10276_y0;
  wire h_u_cla32_and10277_y0;
  wire h_u_cla32_and10278_y0;
  wire h_u_cla32_and10279_y0;
  wire h_u_cla32_and10280_y0;
  wire h_u_cla32_and10281_y0;
  wire h_u_cla32_and10282_y0;
  wire h_u_cla32_and10283_y0;
  wire h_u_cla32_and10284_y0;
  wire h_u_cla32_and10285_y0;
  wire h_u_cla32_and10286_y0;
  wire h_u_cla32_and10287_y0;
  wire h_u_cla32_and10288_y0;
  wire h_u_cla32_and10289_y0;
  wire h_u_cla32_and10290_y0;
  wire h_u_cla32_and10291_y0;
  wire h_u_cla32_and10292_y0;
  wire h_u_cla32_and10293_y0;
  wire h_u_cla32_and10294_y0;
  wire h_u_cla32_and10295_y0;
  wire h_u_cla32_and10296_y0;
  wire h_u_cla32_and10297_y0;
  wire h_u_cla32_and10298_y0;
  wire h_u_cla32_and10299_y0;
  wire h_u_cla32_and10300_y0;
  wire h_u_cla32_and10301_y0;
  wire h_u_cla32_and10302_y0;
  wire h_u_cla32_and10303_y0;
  wire h_u_cla32_and10304_y0;
  wire h_u_cla32_and10305_y0;
  wire h_u_cla32_and10306_y0;
  wire h_u_cla32_and10307_y0;
  wire h_u_cla32_and10308_y0;
  wire h_u_cla32_and10309_y0;
  wire h_u_cla32_and10310_y0;
  wire h_u_cla32_and10311_y0;
  wire h_u_cla32_and10312_y0;
  wire h_u_cla32_and10313_y0;
  wire h_u_cla32_and10314_y0;
  wire h_u_cla32_and10315_y0;
  wire h_u_cla32_and10316_y0;
  wire h_u_cla32_and10317_y0;
  wire h_u_cla32_and10318_y0;
  wire h_u_cla32_and10319_y0;
  wire h_u_cla32_and10320_y0;
  wire h_u_cla32_and10321_y0;
  wire h_u_cla32_and10322_y0;
  wire h_u_cla32_and10323_y0;
  wire h_u_cla32_and10324_y0;
  wire h_u_cla32_and10325_y0;
  wire h_u_cla32_and10326_y0;
  wire h_u_cla32_and10327_y0;
  wire h_u_cla32_and10328_y0;
  wire h_u_cla32_and10329_y0;
  wire h_u_cla32_and10330_y0;
  wire h_u_cla32_and10331_y0;
  wire h_u_cla32_and10332_y0;
  wire h_u_cla32_and10333_y0;
  wire h_u_cla32_and10334_y0;
  wire h_u_cla32_and10335_y0;
  wire h_u_cla32_and10336_y0;
  wire h_u_cla32_and10337_y0;
  wire h_u_cla32_and10338_y0;
  wire h_u_cla32_and10339_y0;
  wire h_u_cla32_and10340_y0;
  wire h_u_cla32_and10341_y0;
  wire h_u_cla32_and10342_y0;
  wire h_u_cla32_and10343_y0;
  wire h_u_cla32_and10344_y0;
  wire h_u_cla32_and10345_y0;
  wire h_u_cla32_and10346_y0;
  wire h_u_cla32_and10347_y0;
  wire h_u_cla32_and10348_y0;
  wire h_u_cla32_and10349_y0;
  wire h_u_cla32_and10350_y0;
  wire h_u_cla32_and10351_y0;
  wire h_u_cla32_and10352_y0;
  wire h_u_cla32_and10353_y0;
  wire h_u_cla32_and10354_y0;
  wire h_u_cla32_and10355_y0;
  wire h_u_cla32_and10356_y0;
  wire h_u_cla32_and10357_y0;
  wire h_u_cla32_and10358_y0;
  wire h_u_cla32_and10359_y0;
  wire h_u_cla32_and10360_y0;
  wire h_u_cla32_and10361_y0;
  wire h_u_cla32_and10362_y0;
  wire h_u_cla32_and10363_y0;
  wire h_u_cla32_and10364_y0;
  wire h_u_cla32_and10365_y0;
  wire h_u_cla32_and10366_y0;
  wire h_u_cla32_and10367_y0;
  wire h_u_cla32_and10368_y0;
  wire h_u_cla32_and10369_y0;
  wire h_u_cla32_and10370_y0;
  wire h_u_cla32_and10371_y0;
  wire h_u_cla32_and10372_y0;
  wire h_u_cla32_and10373_y0;
  wire h_u_cla32_and10374_y0;
  wire h_u_cla32_and10375_y0;
  wire h_u_cla32_and10376_y0;
  wire h_u_cla32_and10377_y0;
  wire h_u_cla32_and10378_y0;
  wire h_u_cla32_and10379_y0;
  wire h_u_cla32_and10380_y0;
  wire h_u_cla32_and10381_y0;
  wire h_u_cla32_and10382_y0;
  wire h_u_cla32_and10383_y0;
  wire h_u_cla32_and10384_y0;
  wire h_u_cla32_and10385_y0;
  wire h_u_cla32_and10386_y0;
  wire h_u_cla32_and10387_y0;
  wire h_u_cla32_and10388_y0;
  wire h_u_cla32_and10389_y0;
  wire h_u_cla32_and10390_y0;
  wire h_u_cla32_and10391_y0;
  wire h_u_cla32_and10392_y0;
  wire h_u_cla32_and10393_y0;
  wire h_u_cla32_and10394_y0;
  wire h_u_cla32_and10395_y0;
  wire h_u_cla32_and10396_y0;
  wire h_u_cla32_and10397_y0;
  wire h_u_cla32_and10398_y0;
  wire h_u_cla32_and10399_y0;
  wire h_u_cla32_and10400_y0;
  wire h_u_cla32_and10401_y0;
  wire h_u_cla32_and10402_y0;
  wire h_u_cla32_and10403_y0;
  wire h_u_cla32_and10404_y0;
  wire h_u_cla32_and10405_y0;
  wire h_u_cla32_and10406_y0;
  wire h_u_cla32_and10407_y0;
  wire h_u_cla32_and10408_y0;
  wire h_u_cla32_and10409_y0;
  wire h_u_cla32_and10410_y0;
  wire h_u_cla32_and10411_y0;
  wire h_u_cla32_and10412_y0;
  wire h_u_cla32_and10413_y0;
  wire h_u_cla32_and10414_y0;
  wire h_u_cla32_and10415_y0;
  wire h_u_cla32_or465_y0;
  wire h_u_cla32_or466_y0;
  wire h_u_cla32_or467_y0;
  wire h_u_cla32_or468_y0;
  wire h_u_cla32_or469_y0;
  wire h_u_cla32_or470_y0;
  wire h_u_cla32_or471_y0;
  wire h_u_cla32_or472_y0;
  wire h_u_cla32_or473_y0;
  wire h_u_cla32_or474_y0;
  wire h_u_cla32_or475_y0;
  wire h_u_cla32_or476_y0;
  wire h_u_cla32_or477_y0;
  wire h_u_cla32_or478_y0;
  wire h_u_cla32_or479_y0;
  wire h_u_cla32_or480_y0;
  wire h_u_cla32_or481_y0;
  wire h_u_cla32_or482_y0;
  wire h_u_cla32_or483_y0;
  wire h_u_cla32_or484_y0;
  wire h_u_cla32_or485_y0;
  wire h_u_cla32_or486_y0;
  wire h_u_cla32_or487_y0;
  wire h_u_cla32_or488_y0;
  wire h_u_cla32_or489_y0;
  wire h_u_cla32_or490_y0;
  wire h_u_cla32_or491_y0;
  wire h_u_cla32_or492_y0;
  wire h_u_cla32_or493_y0;
  wire h_u_cla32_or494_y0;
  wire h_u_cla32_or495_y0;
  wire h_u_cla32_pg_logic31_y0;
  wire h_u_cla32_pg_logic31_y1;
  wire h_u_cla32_pg_logic31_y2;
  wire h_u_cla32_xor31_y0;
  wire h_u_cla32_and10416_y0;
  wire h_u_cla32_and10417_y0;
  wire h_u_cla32_and10418_y0;
  wire h_u_cla32_and10419_y0;
  wire h_u_cla32_and10420_y0;
  wire h_u_cla32_and10421_y0;
  wire h_u_cla32_and10422_y0;
  wire h_u_cla32_and10423_y0;
  wire h_u_cla32_and10424_y0;
  wire h_u_cla32_and10425_y0;
  wire h_u_cla32_and10426_y0;
  wire h_u_cla32_and10427_y0;
  wire h_u_cla32_and10428_y0;
  wire h_u_cla32_and10429_y0;
  wire h_u_cla32_and10430_y0;
  wire h_u_cla32_and10431_y0;
  wire h_u_cla32_and10432_y0;
  wire h_u_cla32_and10433_y0;
  wire h_u_cla32_and10434_y0;
  wire h_u_cla32_and10435_y0;
  wire h_u_cla32_and10436_y0;
  wire h_u_cla32_and10437_y0;
  wire h_u_cla32_and10438_y0;
  wire h_u_cla32_and10439_y0;
  wire h_u_cla32_and10440_y0;
  wire h_u_cla32_and10441_y0;
  wire h_u_cla32_and10442_y0;
  wire h_u_cla32_and10443_y0;
  wire h_u_cla32_and10444_y0;
  wire h_u_cla32_and10445_y0;
  wire h_u_cla32_and10446_y0;
  wire h_u_cla32_and10447_y0;
  wire h_u_cla32_and10448_y0;
  wire h_u_cla32_and10449_y0;
  wire h_u_cla32_and10450_y0;
  wire h_u_cla32_and10451_y0;
  wire h_u_cla32_and10452_y0;
  wire h_u_cla32_and10453_y0;
  wire h_u_cla32_and10454_y0;
  wire h_u_cla32_and10455_y0;
  wire h_u_cla32_and10456_y0;
  wire h_u_cla32_and10457_y0;
  wire h_u_cla32_and10458_y0;
  wire h_u_cla32_and10459_y0;
  wire h_u_cla32_and10460_y0;
  wire h_u_cla32_and10461_y0;
  wire h_u_cla32_and10462_y0;
  wire h_u_cla32_and10463_y0;
  wire h_u_cla32_and10464_y0;
  wire h_u_cla32_and10465_y0;
  wire h_u_cla32_and10466_y0;
  wire h_u_cla32_and10467_y0;
  wire h_u_cla32_and10468_y0;
  wire h_u_cla32_and10469_y0;
  wire h_u_cla32_and10470_y0;
  wire h_u_cla32_and10471_y0;
  wire h_u_cla32_and10472_y0;
  wire h_u_cla32_and10473_y0;
  wire h_u_cla32_and10474_y0;
  wire h_u_cla32_and10475_y0;
  wire h_u_cla32_and10476_y0;
  wire h_u_cla32_and10477_y0;
  wire h_u_cla32_and10478_y0;
  wire h_u_cla32_and10479_y0;
  wire h_u_cla32_and10480_y0;
  wire h_u_cla32_and10481_y0;
  wire h_u_cla32_and10482_y0;
  wire h_u_cla32_and10483_y0;
  wire h_u_cla32_and10484_y0;
  wire h_u_cla32_and10485_y0;
  wire h_u_cla32_and10486_y0;
  wire h_u_cla32_and10487_y0;
  wire h_u_cla32_and10488_y0;
  wire h_u_cla32_and10489_y0;
  wire h_u_cla32_and10490_y0;
  wire h_u_cla32_and10491_y0;
  wire h_u_cla32_and10492_y0;
  wire h_u_cla32_and10493_y0;
  wire h_u_cla32_and10494_y0;
  wire h_u_cla32_and10495_y0;
  wire h_u_cla32_and10496_y0;
  wire h_u_cla32_and10497_y0;
  wire h_u_cla32_and10498_y0;
  wire h_u_cla32_and10499_y0;
  wire h_u_cla32_and10500_y0;
  wire h_u_cla32_and10501_y0;
  wire h_u_cla32_and10502_y0;
  wire h_u_cla32_and10503_y0;
  wire h_u_cla32_and10504_y0;
  wire h_u_cla32_and10505_y0;
  wire h_u_cla32_and10506_y0;
  wire h_u_cla32_and10507_y0;
  wire h_u_cla32_and10508_y0;
  wire h_u_cla32_and10509_y0;
  wire h_u_cla32_and10510_y0;
  wire h_u_cla32_and10511_y0;
  wire h_u_cla32_and10512_y0;
  wire h_u_cla32_and10513_y0;
  wire h_u_cla32_and10514_y0;
  wire h_u_cla32_and10515_y0;
  wire h_u_cla32_and10516_y0;
  wire h_u_cla32_and10517_y0;
  wire h_u_cla32_and10518_y0;
  wire h_u_cla32_and10519_y0;
  wire h_u_cla32_and10520_y0;
  wire h_u_cla32_and10521_y0;
  wire h_u_cla32_and10522_y0;
  wire h_u_cla32_and10523_y0;
  wire h_u_cla32_and10524_y0;
  wire h_u_cla32_and10525_y0;
  wire h_u_cla32_and10526_y0;
  wire h_u_cla32_and10527_y0;
  wire h_u_cla32_and10528_y0;
  wire h_u_cla32_and10529_y0;
  wire h_u_cla32_and10530_y0;
  wire h_u_cla32_and10531_y0;
  wire h_u_cla32_and10532_y0;
  wire h_u_cla32_and10533_y0;
  wire h_u_cla32_and10534_y0;
  wire h_u_cla32_and10535_y0;
  wire h_u_cla32_and10536_y0;
  wire h_u_cla32_and10537_y0;
  wire h_u_cla32_and10538_y0;
  wire h_u_cla32_and10539_y0;
  wire h_u_cla32_and10540_y0;
  wire h_u_cla32_and10541_y0;
  wire h_u_cla32_and10542_y0;
  wire h_u_cla32_and10543_y0;
  wire h_u_cla32_and10544_y0;
  wire h_u_cla32_and10545_y0;
  wire h_u_cla32_and10546_y0;
  wire h_u_cla32_and10547_y0;
  wire h_u_cla32_and10548_y0;
  wire h_u_cla32_and10549_y0;
  wire h_u_cla32_and10550_y0;
  wire h_u_cla32_and10551_y0;
  wire h_u_cla32_and10552_y0;
  wire h_u_cla32_and10553_y0;
  wire h_u_cla32_and10554_y0;
  wire h_u_cla32_and10555_y0;
  wire h_u_cla32_and10556_y0;
  wire h_u_cla32_and10557_y0;
  wire h_u_cla32_and10558_y0;
  wire h_u_cla32_and10559_y0;
  wire h_u_cla32_and10560_y0;
  wire h_u_cla32_and10561_y0;
  wire h_u_cla32_and10562_y0;
  wire h_u_cla32_and10563_y0;
  wire h_u_cla32_and10564_y0;
  wire h_u_cla32_and10565_y0;
  wire h_u_cla32_and10566_y0;
  wire h_u_cla32_and10567_y0;
  wire h_u_cla32_and10568_y0;
  wire h_u_cla32_and10569_y0;
  wire h_u_cla32_and10570_y0;
  wire h_u_cla32_and10571_y0;
  wire h_u_cla32_and10572_y0;
  wire h_u_cla32_and10573_y0;
  wire h_u_cla32_and10574_y0;
  wire h_u_cla32_and10575_y0;
  wire h_u_cla32_and10576_y0;
  wire h_u_cla32_and10577_y0;
  wire h_u_cla32_and10578_y0;
  wire h_u_cla32_and10579_y0;
  wire h_u_cla32_and10580_y0;
  wire h_u_cla32_and10581_y0;
  wire h_u_cla32_and10582_y0;
  wire h_u_cla32_and10583_y0;
  wire h_u_cla32_and10584_y0;
  wire h_u_cla32_and10585_y0;
  wire h_u_cla32_and10586_y0;
  wire h_u_cla32_and10587_y0;
  wire h_u_cla32_and10588_y0;
  wire h_u_cla32_and10589_y0;
  wire h_u_cla32_and10590_y0;
  wire h_u_cla32_and10591_y0;
  wire h_u_cla32_and10592_y0;
  wire h_u_cla32_and10593_y0;
  wire h_u_cla32_and10594_y0;
  wire h_u_cla32_and10595_y0;
  wire h_u_cla32_and10596_y0;
  wire h_u_cla32_and10597_y0;
  wire h_u_cla32_and10598_y0;
  wire h_u_cla32_and10599_y0;
  wire h_u_cla32_and10600_y0;
  wire h_u_cla32_and10601_y0;
  wire h_u_cla32_and10602_y0;
  wire h_u_cla32_and10603_y0;
  wire h_u_cla32_and10604_y0;
  wire h_u_cla32_and10605_y0;
  wire h_u_cla32_and10606_y0;
  wire h_u_cla32_and10607_y0;
  wire h_u_cla32_and10608_y0;
  wire h_u_cla32_and10609_y0;
  wire h_u_cla32_and10610_y0;
  wire h_u_cla32_and10611_y0;
  wire h_u_cla32_and10612_y0;
  wire h_u_cla32_and10613_y0;
  wire h_u_cla32_and10614_y0;
  wire h_u_cla32_and10615_y0;
  wire h_u_cla32_and10616_y0;
  wire h_u_cla32_and10617_y0;
  wire h_u_cla32_and10618_y0;
  wire h_u_cla32_and10619_y0;
  wire h_u_cla32_and10620_y0;
  wire h_u_cla32_and10621_y0;
  wire h_u_cla32_and10622_y0;
  wire h_u_cla32_and10623_y0;
  wire h_u_cla32_and10624_y0;
  wire h_u_cla32_and10625_y0;
  wire h_u_cla32_and10626_y0;
  wire h_u_cla32_and10627_y0;
  wire h_u_cla32_and10628_y0;
  wire h_u_cla32_and10629_y0;
  wire h_u_cla32_and10630_y0;
  wire h_u_cla32_and10631_y0;
  wire h_u_cla32_and10632_y0;
  wire h_u_cla32_and10633_y0;
  wire h_u_cla32_and10634_y0;
  wire h_u_cla32_and10635_y0;
  wire h_u_cla32_and10636_y0;
  wire h_u_cla32_and10637_y0;
  wire h_u_cla32_and10638_y0;
  wire h_u_cla32_and10639_y0;
  wire h_u_cla32_and10640_y0;
  wire h_u_cla32_and10641_y0;
  wire h_u_cla32_and10642_y0;
  wire h_u_cla32_and10643_y0;
  wire h_u_cla32_and10644_y0;
  wire h_u_cla32_and10645_y0;
  wire h_u_cla32_and10646_y0;
  wire h_u_cla32_and10647_y0;
  wire h_u_cla32_and10648_y0;
  wire h_u_cla32_and10649_y0;
  wire h_u_cla32_and10650_y0;
  wire h_u_cla32_and10651_y0;
  wire h_u_cla32_and10652_y0;
  wire h_u_cla32_and10653_y0;
  wire h_u_cla32_and10654_y0;
  wire h_u_cla32_and10655_y0;
  wire h_u_cla32_and10656_y0;
  wire h_u_cla32_and10657_y0;
  wire h_u_cla32_and10658_y0;
  wire h_u_cla32_and10659_y0;
  wire h_u_cla32_and10660_y0;
  wire h_u_cla32_and10661_y0;
  wire h_u_cla32_and10662_y0;
  wire h_u_cla32_and10663_y0;
  wire h_u_cla32_and10664_y0;
  wire h_u_cla32_and10665_y0;
  wire h_u_cla32_and10666_y0;
  wire h_u_cla32_and10667_y0;
  wire h_u_cla32_and10668_y0;
  wire h_u_cla32_and10669_y0;
  wire h_u_cla32_and10670_y0;
  wire h_u_cla32_and10671_y0;
  wire h_u_cla32_and10672_y0;
  wire h_u_cla32_and10673_y0;
  wire h_u_cla32_and10674_y0;
  wire h_u_cla32_and10675_y0;
  wire h_u_cla32_and10676_y0;
  wire h_u_cla32_and10677_y0;
  wire h_u_cla32_and10678_y0;
  wire h_u_cla32_and10679_y0;
  wire h_u_cla32_and10680_y0;
  wire h_u_cla32_and10681_y0;
  wire h_u_cla32_and10682_y0;
  wire h_u_cla32_and10683_y0;
  wire h_u_cla32_and10684_y0;
  wire h_u_cla32_and10685_y0;
  wire h_u_cla32_and10686_y0;
  wire h_u_cla32_and10687_y0;
  wire h_u_cla32_and10688_y0;
  wire h_u_cla32_and10689_y0;
  wire h_u_cla32_and10690_y0;
  wire h_u_cla32_and10691_y0;
  wire h_u_cla32_and10692_y0;
  wire h_u_cla32_and10693_y0;
  wire h_u_cla32_and10694_y0;
  wire h_u_cla32_and10695_y0;
  wire h_u_cla32_and10696_y0;
  wire h_u_cla32_and10697_y0;
  wire h_u_cla32_and10698_y0;
  wire h_u_cla32_and10699_y0;
  wire h_u_cla32_and10700_y0;
  wire h_u_cla32_and10701_y0;
  wire h_u_cla32_and10702_y0;
  wire h_u_cla32_and10703_y0;
  wire h_u_cla32_and10704_y0;
  wire h_u_cla32_and10705_y0;
  wire h_u_cla32_and10706_y0;
  wire h_u_cla32_and10707_y0;
  wire h_u_cla32_and10708_y0;
  wire h_u_cla32_and10709_y0;
  wire h_u_cla32_and10710_y0;
  wire h_u_cla32_and10711_y0;
  wire h_u_cla32_and10712_y0;
  wire h_u_cla32_and10713_y0;
  wire h_u_cla32_and10714_y0;
  wire h_u_cla32_and10715_y0;
  wire h_u_cla32_and10716_y0;
  wire h_u_cla32_and10717_y0;
  wire h_u_cla32_and10718_y0;
  wire h_u_cla32_and10719_y0;
  wire h_u_cla32_and10720_y0;
  wire h_u_cla32_and10721_y0;
  wire h_u_cla32_and10722_y0;
  wire h_u_cla32_and10723_y0;
  wire h_u_cla32_and10724_y0;
  wire h_u_cla32_and10725_y0;
  wire h_u_cla32_and10726_y0;
  wire h_u_cla32_and10727_y0;
  wire h_u_cla32_and10728_y0;
  wire h_u_cla32_and10729_y0;
  wire h_u_cla32_and10730_y0;
  wire h_u_cla32_and10731_y0;
  wire h_u_cla32_and10732_y0;
  wire h_u_cla32_and10733_y0;
  wire h_u_cla32_and10734_y0;
  wire h_u_cla32_and10735_y0;
  wire h_u_cla32_and10736_y0;
  wire h_u_cla32_and10737_y0;
  wire h_u_cla32_and10738_y0;
  wire h_u_cla32_and10739_y0;
  wire h_u_cla32_and10740_y0;
  wire h_u_cla32_and10741_y0;
  wire h_u_cla32_and10742_y0;
  wire h_u_cla32_and10743_y0;
  wire h_u_cla32_and10744_y0;
  wire h_u_cla32_and10745_y0;
  wire h_u_cla32_and10746_y0;
  wire h_u_cla32_and10747_y0;
  wire h_u_cla32_and10748_y0;
  wire h_u_cla32_and10749_y0;
  wire h_u_cla32_and10750_y0;
  wire h_u_cla32_and10751_y0;
  wire h_u_cla32_and10752_y0;
  wire h_u_cla32_and10753_y0;
  wire h_u_cla32_and10754_y0;
  wire h_u_cla32_and10755_y0;
  wire h_u_cla32_and10756_y0;
  wire h_u_cla32_and10757_y0;
  wire h_u_cla32_and10758_y0;
  wire h_u_cla32_and10759_y0;
  wire h_u_cla32_and10760_y0;
  wire h_u_cla32_and10761_y0;
  wire h_u_cla32_and10762_y0;
  wire h_u_cla32_and10763_y0;
  wire h_u_cla32_and10764_y0;
  wire h_u_cla32_and10765_y0;
  wire h_u_cla32_and10766_y0;
  wire h_u_cla32_and10767_y0;
  wire h_u_cla32_and10768_y0;
  wire h_u_cla32_and10769_y0;
  wire h_u_cla32_and10770_y0;
  wire h_u_cla32_and10771_y0;
  wire h_u_cla32_and10772_y0;
  wire h_u_cla32_and10773_y0;
  wire h_u_cla32_and10774_y0;
  wire h_u_cla32_and10775_y0;
  wire h_u_cla32_and10776_y0;
  wire h_u_cla32_and10777_y0;
  wire h_u_cla32_and10778_y0;
  wire h_u_cla32_and10779_y0;
  wire h_u_cla32_and10780_y0;
  wire h_u_cla32_and10781_y0;
  wire h_u_cla32_and10782_y0;
  wire h_u_cla32_and10783_y0;
  wire h_u_cla32_and10784_y0;
  wire h_u_cla32_and10785_y0;
  wire h_u_cla32_and10786_y0;
  wire h_u_cla32_and10787_y0;
  wire h_u_cla32_and10788_y0;
  wire h_u_cla32_and10789_y0;
  wire h_u_cla32_and10790_y0;
  wire h_u_cla32_and10791_y0;
  wire h_u_cla32_and10792_y0;
  wire h_u_cla32_and10793_y0;
  wire h_u_cla32_and10794_y0;
  wire h_u_cla32_and10795_y0;
  wire h_u_cla32_and10796_y0;
  wire h_u_cla32_and10797_y0;
  wire h_u_cla32_and10798_y0;
  wire h_u_cla32_and10799_y0;
  wire h_u_cla32_and10800_y0;
  wire h_u_cla32_and10801_y0;
  wire h_u_cla32_and10802_y0;
  wire h_u_cla32_and10803_y0;
  wire h_u_cla32_and10804_y0;
  wire h_u_cla32_and10805_y0;
  wire h_u_cla32_and10806_y0;
  wire h_u_cla32_and10807_y0;
  wire h_u_cla32_and10808_y0;
  wire h_u_cla32_and10809_y0;
  wire h_u_cla32_and10810_y0;
  wire h_u_cla32_and10811_y0;
  wire h_u_cla32_and10812_y0;
  wire h_u_cla32_and10813_y0;
  wire h_u_cla32_and10814_y0;
  wire h_u_cla32_and10815_y0;
  wire h_u_cla32_and10816_y0;
  wire h_u_cla32_and10817_y0;
  wire h_u_cla32_and10818_y0;
  wire h_u_cla32_and10819_y0;
  wire h_u_cla32_and10820_y0;
  wire h_u_cla32_and10821_y0;
  wire h_u_cla32_and10822_y0;
  wire h_u_cla32_and10823_y0;
  wire h_u_cla32_and10824_y0;
  wire h_u_cla32_and10825_y0;
  wire h_u_cla32_and10826_y0;
  wire h_u_cla32_and10827_y0;
  wire h_u_cla32_and10828_y0;
  wire h_u_cla32_and10829_y0;
  wire h_u_cla32_and10830_y0;
  wire h_u_cla32_and10831_y0;
  wire h_u_cla32_and10832_y0;
  wire h_u_cla32_and10833_y0;
  wire h_u_cla32_and10834_y0;
  wire h_u_cla32_and10835_y0;
  wire h_u_cla32_and10836_y0;
  wire h_u_cla32_and10837_y0;
  wire h_u_cla32_and10838_y0;
  wire h_u_cla32_and10839_y0;
  wire h_u_cla32_and10840_y0;
  wire h_u_cla32_and10841_y0;
  wire h_u_cla32_and10842_y0;
  wire h_u_cla32_and10843_y0;
  wire h_u_cla32_and10844_y0;
  wire h_u_cla32_and10845_y0;
  wire h_u_cla32_and10846_y0;
  wire h_u_cla32_and10847_y0;
  wire h_u_cla32_and10848_y0;
  wire h_u_cla32_and10849_y0;
  wire h_u_cla32_and10850_y0;
  wire h_u_cla32_and10851_y0;
  wire h_u_cla32_and10852_y0;
  wire h_u_cla32_and10853_y0;
  wire h_u_cla32_and10854_y0;
  wire h_u_cla32_and10855_y0;
  wire h_u_cla32_and10856_y0;
  wire h_u_cla32_and10857_y0;
  wire h_u_cla32_and10858_y0;
  wire h_u_cla32_and10859_y0;
  wire h_u_cla32_and10860_y0;
  wire h_u_cla32_and10861_y0;
  wire h_u_cla32_and10862_y0;
  wire h_u_cla32_and10863_y0;
  wire h_u_cla32_and10864_y0;
  wire h_u_cla32_and10865_y0;
  wire h_u_cla32_and10866_y0;
  wire h_u_cla32_and10867_y0;
  wire h_u_cla32_and10868_y0;
  wire h_u_cla32_and10869_y0;
  wire h_u_cla32_and10870_y0;
  wire h_u_cla32_and10871_y0;
  wire h_u_cla32_and10872_y0;
  wire h_u_cla32_and10873_y0;
  wire h_u_cla32_and10874_y0;
  wire h_u_cla32_and10875_y0;
  wire h_u_cla32_and10876_y0;
  wire h_u_cla32_and10877_y0;
  wire h_u_cla32_and10878_y0;
  wire h_u_cla32_and10879_y0;
  wire h_u_cla32_and10880_y0;
  wire h_u_cla32_and10881_y0;
  wire h_u_cla32_and10882_y0;
  wire h_u_cla32_and10883_y0;
  wire h_u_cla32_and10884_y0;
  wire h_u_cla32_and10885_y0;
  wire h_u_cla32_and10886_y0;
  wire h_u_cla32_and10887_y0;
  wire h_u_cla32_and10888_y0;
  wire h_u_cla32_and10889_y0;
  wire h_u_cla32_and10890_y0;
  wire h_u_cla32_and10891_y0;
  wire h_u_cla32_and10892_y0;
  wire h_u_cla32_and10893_y0;
  wire h_u_cla32_and10894_y0;
  wire h_u_cla32_and10895_y0;
  wire h_u_cla32_and10896_y0;
  wire h_u_cla32_and10897_y0;
  wire h_u_cla32_and10898_y0;
  wire h_u_cla32_and10899_y0;
  wire h_u_cla32_and10900_y0;
  wire h_u_cla32_and10901_y0;
  wire h_u_cla32_and10902_y0;
  wire h_u_cla32_and10903_y0;
  wire h_u_cla32_and10904_y0;
  wire h_u_cla32_and10905_y0;
  wire h_u_cla32_and10906_y0;
  wire h_u_cla32_and10907_y0;
  wire h_u_cla32_and10908_y0;
  wire h_u_cla32_and10909_y0;
  wire h_u_cla32_and10910_y0;
  wire h_u_cla32_and10911_y0;
  wire h_u_cla32_and10912_y0;
  wire h_u_cla32_and10913_y0;
  wire h_u_cla32_and10914_y0;
  wire h_u_cla32_and10915_y0;
  wire h_u_cla32_and10916_y0;
  wire h_u_cla32_and10917_y0;
  wire h_u_cla32_and10918_y0;
  wire h_u_cla32_and10919_y0;
  wire h_u_cla32_and10920_y0;
  wire h_u_cla32_and10921_y0;
  wire h_u_cla32_and10922_y0;
  wire h_u_cla32_and10923_y0;
  wire h_u_cla32_and10924_y0;
  wire h_u_cla32_and10925_y0;
  wire h_u_cla32_and10926_y0;
  wire h_u_cla32_and10927_y0;
  wire h_u_cla32_and10928_y0;
  wire h_u_cla32_and10929_y0;
  wire h_u_cla32_and10930_y0;
  wire h_u_cla32_and10931_y0;
  wire h_u_cla32_and10932_y0;
  wire h_u_cla32_and10933_y0;
  wire h_u_cla32_and10934_y0;
  wire h_u_cla32_and10935_y0;
  wire h_u_cla32_and10936_y0;
  wire h_u_cla32_and10937_y0;
  wire h_u_cla32_and10938_y0;
  wire h_u_cla32_and10939_y0;
  wire h_u_cla32_and10940_y0;
  wire h_u_cla32_and10941_y0;
  wire h_u_cla32_and10942_y0;
  wire h_u_cla32_and10943_y0;
  wire h_u_cla32_and10944_y0;
  wire h_u_cla32_and10945_y0;
  wire h_u_cla32_and10946_y0;
  wire h_u_cla32_and10947_y0;
  wire h_u_cla32_and10948_y0;
  wire h_u_cla32_and10949_y0;
  wire h_u_cla32_and10950_y0;
  wire h_u_cla32_and10951_y0;
  wire h_u_cla32_and10952_y0;
  wire h_u_cla32_and10953_y0;
  wire h_u_cla32_and10954_y0;
  wire h_u_cla32_and10955_y0;
  wire h_u_cla32_and10956_y0;
  wire h_u_cla32_and10957_y0;
  wire h_u_cla32_and10958_y0;
  wire h_u_cla32_and10959_y0;
  wire h_u_cla32_and10960_y0;
  wire h_u_cla32_and10961_y0;
  wire h_u_cla32_and10962_y0;
  wire h_u_cla32_and10963_y0;
  wire h_u_cla32_and10964_y0;
  wire h_u_cla32_and10965_y0;
  wire h_u_cla32_and10966_y0;
  wire h_u_cla32_and10967_y0;
  wire h_u_cla32_and10968_y0;
  wire h_u_cla32_and10969_y0;
  wire h_u_cla32_and10970_y0;
  wire h_u_cla32_and10971_y0;
  wire h_u_cla32_and10972_y0;
  wire h_u_cla32_and10973_y0;
  wire h_u_cla32_and10974_y0;
  wire h_u_cla32_and10975_y0;
  wire h_u_cla32_and10976_y0;
  wire h_u_cla32_and10977_y0;
  wire h_u_cla32_and10978_y0;
  wire h_u_cla32_and10979_y0;
  wire h_u_cla32_and10980_y0;
  wire h_u_cla32_and10981_y0;
  wire h_u_cla32_and10982_y0;
  wire h_u_cla32_and10983_y0;
  wire h_u_cla32_and10984_y0;
  wire h_u_cla32_and10985_y0;
  wire h_u_cla32_and10986_y0;
  wire h_u_cla32_and10987_y0;
  wire h_u_cla32_and10988_y0;
  wire h_u_cla32_and10989_y0;
  wire h_u_cla32_and10990_y0;
  wire h_u_cla32_and10991_y0;
  wire h_u_cla32_and10992_y0;
  wire h_u_cla32_and10993_y0;
  wire h_u_cla32_and10994_y0;
  wire h_u_cla32_and10995_y0;
  wire h_u_cla32_and10996_y0;
  wire h_u_cla32_and10997_y0;
  wire h_u_cla32_and10998_y0;
  wire h_u_cla32_and10999_y0;
  wire h_u_cla32_and11000_y0;
  wire h_u_cla32_and11001_y0;
  wire h_u_cla32_and11002_y0;
  wire h_u_cla32_and11003_y0;
  wire h_u_cla32_and11004_y0;
  wire h_u_cla32_and11005_y0;
  wire h_u_cla32_and11006_y0;
  wire h_u_cla32_and11007_y0;
  wire h_u_cla32_and11008_y0;
  wire h_u_cla32_and11009_y0;
  wire h_u_cla32_and11010_y0;
  wire h_u_cla32_and11011_y0;
  wire h_u_cla32_and11012_y0;
  wire h_u_cla32_and11013_y0;
  wire h_u_cla32_and11014_y0;
  wire h_u_cla32_and11015_y0;
  wire h_u_cla32_and11016_y0;
  wire h_u_cla32_and11017_y0;
  wire h_u_cla32_and11018_y0;
  wire h_u_cla32_and11019_y0;
  wire h_u_cla32_and11020_y0;
  wire h_u_cla32_and11021_y0;
  wire h_u_cla32_and11022_y0;
  wire h_u_cla32_and11023_y0;
  wire h_u_cla32_and11024_y0;
  wire h_u_cla32_and11025_y0;
  wire h_u_cla32_and11026_y0;
  wire h_u_cla32_and11027_y0;
  wire h_u_cla32_and11028_y0;
  wire h_u_cla32_and11029_y0;
  wire h_u_cla32_and11030_y0;
  wire h_u_cla32_and11031_y0;
  wire h_u_cla32_and11032_y0;
  wire h_u_cla32_and11033_y0;
  wire h_u_cla32_and11034_y0;
  wire h_u_cla32_and11035_y0;
  wire h_u_cla32_and11036_y0;
  wire h_u_cla32_and11037_y0;
  wire h_u_cla32_and11038_y0;
  wire h_u_cla32_and11039_y0;
  wire h_u_cla32_and11040_y0;
  wire h_u_cla32_and11041_y0;
  wire h_u_cla32_and11042_y0;
  wire h_u_cla32_and11043_y0;
  wire h_u_cla32_and11044_y0;
  wire h_u_cla32_and11045_y0;
  wire h_u_cla32_and11046_y0;
  wire h_u_cla32_and11047_y0;
  wire h_u_cla32_and11048_y0;
  wire h_u_cla32_and11049_y0;
  wire h_u_cla32_and11050_y0;
  wire h_u_cla32_and11051_y0;
  wire h_u_cla32_and11052_y0;
  wire h_u_cla32_and11053_y0;
  wire h_u_cla32_and11054_y0;
  wire h_u_cla32_and11055_y0;
  wire h_u_cla32_and11056_y0;
  wire h_u_cla32_and11057_y0;
  wire h_u_cla32_and11058_y0;
  wire h_u_cla32_and11059_y0;
  wire h_u_cla32_and11060_y0;
  wire h_u_cla32_and11061_y0;
  wire h_u_cla32_and11062_y0;
  wire h_u_cla32_and11063_y0;
  wire h_u_cla32_and11064_y0;
  wire h_u_cla32_and11065_y0;
  wire h_u_cla32_and11066_y0;
  wire h_u_cla32_and11067_y0;
  wire h_u_cla32_and11068_y0;
  wire h_u_cla32_and11069_y0;
  wire h_u_cla32_and11070_y0;
  wire h_u_cla32_and11071_y0;
  wire h_u_cla32_and11072_y0;
  wire h_u_cla32_and11073_y0;
  wire h_u_cla32_and11074_y0;
  wire h_u_cla32_and11075_y0;
  wire h_u_cla32_and11076_y0;
  wire h_u_cla32_and11077_y0;
  wire h_u_cla32_and11078_y0;
  wire h_u_cla32_and11079_y0;
  wire h_u_cla32_and11080_y0;
  wire h_u_cla32_and11081_y0;
  wire h_u_cla32_and11082_y0;
  wire h_u_cla32_and11083_y0;
  wire h_u_cla32_and11084_y0;
  wire h_u_cla32_and11085_y0;
  wire h_u_cla32_and11086_y0;
  wire h_u_cla32_and11087_y0;
  wire h_u_cla32_and11088_y0;
  wire h_u_cla32_and11089_y0;
  wire h_u_cla32_and11090_y0;
  wire h_u_cla32_and11091_y0;
  wire h_u_cla32_and11092_y0;
  wire h_u_cla32_and11093_y0;
  wire h_u_cla32_and11094_y0;
  wire h_u_cla32_and11095_y0;
  wire h_u_cla32_and11096_y0;
  wire h_u_cla32_and11097_y0;
  wire h_u_cla32_and11098_y0;
  wire h_u_cla32_and11099_y0;
  wire h_u_cla32_and11100_y0;
  wire h_u_cla32_and11101_y0;
  wire h_u_cla32_and11102_y0;
  wire h_u_cla32_and11103_y0;
  wire h_u_cla32_and11104_y0;
  wire h_u_cla32_and11105_y0;
  wire h_u_cla32_and11106_y0;
  wire h_u_cla32_and11107_y0;
  wire h_u_cla32_and11108_y0;
  wire h_u_cla32_and11109_y0;
  wire h_u_cla32_and11110_y0;
  wire h_u_cla32_and11111_y0;
  wire h_u_cla32_and11112_y0;
  wire h_u_cla32_and11113_y0;
  wire h_u_cla32_and11114_y0;
  wire h_u_cla32_and11115_y0;
  wire h_u_cla32_and11116_y0;
  wire h_u_cla32_and11117_y0;
  wire h_u_cla32_and11118_y0;
  wire h_u_cla32_and11119_y0;
  wire h_u_cla32_and11120_y0;
  wire h_u_cla32_and11121_y0;
  wire h_u_cla32_and11122_y0;
  wire h_u_cla32_and11123_y0;
  wire h_u_cla32_and11124_y0;
  wire h_u_cla32_and11125_y0;
  wire h_u_cla32_and11126_y0;
  wire h_u_cla32_and11127_y0;
  wire h_u_cla32_and11128_y0;
  wire h_u_cla32_and11129_y0;
  wire h_u_cla32_and11130_y0;
  wire h_u_cla32_and11131_y0;
  wire h_u_cla32_and11132_y0;
  wire h_u_cla32_and11133_y0;
  wire h_u_cla32_and11134_y0;
  wire h_u_cla32_and11135_y0;
  wire h_u_cla32_and11136_y0;
  wire h_u_cla32_and11137_y0;
  wire h_u_cla32_and11138_y0;
  wire h_u_cla32_and11139_y0;
  wire h_u_cla32_and11140_y0;
  wire h_u_cla32_and11141_y0;
  wire h_u_cla32_and11142_y0;
  wire h_u_cla32_and11143_y0;
  wire h_u_cla32_and11144_y0;
  wire h_u_cla32_and11145_y0;
  wire h_u_cla32_and11146_y0;
  wire h_u_cla32_and11147_y0;
  wire h_u_cla32_and11148_y0;
  wire h_u_cla32_and11149_y0;
  wire h_u_cla32_and11150_y0;
  wire h_u_cla32_and11151_y0;
  wire h_u_cla32_and11152_y0;
  wire h_u_cla32_and11153_y0;
  wire h_u_cla32_and11154_y0;
  wire h_u_cla32_and11155_y0;
  wire h_u_cla32_and11156_y0;
  wire h_u_cla32_and11157_y0;
  wire h_u_cla32_and11158_y0;
  wire h_u_cla32_and11159_y0;
  wire h_u_cla32_and11160_y0;
  wire h_u_cla32_and11161_y0;
  wire h_u_cla32_and11162_y0;
  wire h_u_cla32_and11163_y0;
  wire h_u_cla32_and11164_y0;
  wire h_u_cla32_and11165_y0;
  wire h_u_cla32_and11166_y0;
  wire h_u_cla32_and11167_y0;
  wire h_u_cla32_and11168_y0;
  wire h_u_cla32_and11169_y0;
  wire h_u_cla32_and11170_y0;
  wire h_u_cla32_and11171_y0;
  wire h_u_cla32_and11172_y0;
  wire h_u_cla32_and11173_y0;
  wire h_u_cla32_and11174_y0;
  wire h_u_cla32_and11175_y0;
  wire h_u_cla32_and11176_y0;
  wire h_u_cla32_and11177_y0;
  wire h_u_cla32_and11178_y0;
  wire h_u_cla32_and11179_y0;
  wire h_u_cla32_and11180_y0;
  wire h_u_cla32_and11181_y0;
  wire h_u_cla32_and11182_y0;
  wire h_u_cla32_and11183_y0;
  wire h_u_cla32_and11184_y0;
  wire h_u_cla32_and11185_y0;
  wire h_u_cla32_and11186_y0;
  wire h_u_cla32_and11187_y0;
  wire h_u_cla32_and11188_y0;
  wire h_u_cla32_and11189_y0;
  wire h_u_cla32_and11190_y0;
  wire h_u_cla32_and11191_y0;
  wire h_u_cla32_and11192_y0;
  wire h_u_cla32_and11193_y0;
  wire h_u_cla32_and11194_y0;
  wire h_u_cla32_and11195_y0;
  wire h_u_cla32_and11196_y0;
  wire h_u_cla32_and11197_y0;
  wire h_u_cla32_and11198_y0;
  wire h_u_cla32_and11199_y0;
  wire h_u_cla32_and11200_y0;
  wire h_u_cla32_and11201_y0;
  wire h_u_cla32_and11202_y0;
  wire h_u_cla32_and11203_y0;
  wire h_u_cla32_and11204_y0;
  wire h_u_cla32_and11205_y0;
  wire h_u_cla32_and11206_y0;
  wire h_u_cla32_and11207_y0;
  wire h_u_cla32_and11208_y0;
  wire h_u_cla32_and11209_y0;
  wire h_u_cla32_and11210_y0;
  wire h_u_cla32_and11211_y0;
  wire h_u_cla32_and11212_y0;
  wire h_u_cla32_and11213_y0;
  wire h_u_cla32_and11214_y0;
  wire h_u_cla32_and11215_y0;
  wire h_u_cla32_and11216_y0;
  wire h_u_cla32_and11217_y0;
  wire h_u_cla32_and11218_y0;
  wire h_u_cla32_and11219_y0;
  wire h_u_cla32_and11220_y0;
  wire h_u_cla32_and11221_y0;
  wire h_u_cla32_and11222_y0;
  wire h_u_cla32_and11223_y0;
  wire h_u_cla32_and11224_y0;
  wire h_u_cla32_and11225_y0;
  wire h_u_cla32_and11226_y0;
  wire h_u_cla32_and11227_y0;
  wire h_u_cla32_and11228_y0;
  wire h_u_cla32_and11229_y0;
  wire h_u_cla32_and11230_y0;
  wire h_u_cla32_and11231_y0;
  wire h_u_cla32_and11232_y0;
  wire h_u_cla32_and11233_y0;
  wire h_u_cla32_and11234_y0;
  wire h_u_cla32_and11235_y0;
  wire h_u_cla32_and11236_y0;
  wire h_u_cla32_and11237_y0;
  wire h_u_cla32_and11238_y0;
  wire h_u_cla32_and11239_y0;
  wire h_u_cla32_and11240_y0;
  wire h_u_cla32_and11241_y0;
  wire h_u_cla32_and11242_y0;
  wire h_u_cla32_and11243_y0;
  wire h_u_cla32_and11244_y0;
  wire h_u_cla32_and11245_y0;
  wire h_u_cla32_and11246_y0;
  wire h_u_cla32_and11247_y0;
  wire h_u_cla32_and11248_y0;
  wire h_u_cla32_and11249_y0;
  wire h_u_cla32_and11250_y0;
  wire h_u_cla32_and11251_y0;
  wire h_u_cla32_and11252_y0;
  wire h_u_cla32_and11253_y0;
  wire h_u_cla32_and11254_y0;
  wire h_u_cla32_and11255_y0;
  wire h_u_cla32_and11256_y0;
  wire h_u_cla32_and11257_y0;
  wire h_u_cla32_and11258_y0;
  wire h_u_cla32_and11259_y0;
  wire h_u_cla32_and11260_y0;
  wire h_u_cla32_and11261_y0;
  wire h_u_cla32_and11262_y0;
  wire h_u_cla32_and11263_y0;
  wire h_u_cla32_and11264_y0;
  wire h_u_cla32_and11265_y0;
  wire h_u_cla32_and11266_y0;
  wire h_u_cla32_and11267_y0;
  wire h_u_cla32_and11268_y0;
  wire h_u_cla32_and11269_y0;
  wire h_u_cla32_and11270_y0;
  wire h_u_cla32_and11271_y0;
  wire h_u_cla32_and11272_y0;
  wire h_u_cla32_and11273_y0;
  wire h_u_cla32_and11274_y0;
  wire h_u_cla32_and11275_y0;
  wire h_u_cla32_and11276_y0;
  wire h_u_cla32_and11277_y0;
  wire h_u_cla32_and11278_y0;
  wire h_u_cla32_and11279_y0;
  wire h_u_cla32_and11280_y0;
  wire h_u_cla32_and11281_y0;
  wire h_u_cla32_and11282_y0;
  wire h_u_cla32_and11283_y0;
  wire h_u_cla32_and11284_y0;
  wire h_u_cla32_and11285_y0;
  wire h_u_cla32_and11286_y0;
  wire h_u_cla32_and11287_y0;
  wire h_u_cla32_and11288_y0;
  wire h_u_cla32_and11289_y0;
  wire h_u_cla32_and11290_y0;
  wire h_u_cla32_and11291_y0;
  wire h_u_cla32_and11292_y0;
  wire h_u_cla32_and11293_y0;
  wire h_u_cla32_and11294_y0;
  wire h_u_cla32_and11295_y0;
  wire h_u_cla32_and11296_y0;
  wire h_u_cla32_and11297_y0;
  wire h_u_cla32_and11298_y0;
  wire h_u_cla32_and11299_y0;
  wire h_u_cla32_and11300_y0;
  wire h_u_cla32_and11301_y0;
  wire h_u_cla32_and11302_y0;
  wire h_u_cla32_and11303_y0;
  wire h_u_cla32_and11304_y0;
  wire h_u_cla32_and11305_y0;
  wire h_u_cla32_and11306_y0;
  wire h_u_cla32_and11307_y0;
  wire h_u_cla32_and11308_y0;
  wire h_u_cla32_and11309_y0;
  wire h_u_cla32_and11310_y0;
  wire h_u_cla32_and11311_y0;
  wire h_u_cla32_and11312_y0;
  wire h_u_cla32_and11313_y0;
  wire h_u_cla32_and11314_y0;
  wire h_u_cla32_and11315_y0;
  wire h_u_cla32_and11316_y0;
  wire h_u_cla32_and11317_y0;
  wire h_u_cla32_and11318_y0;
  wire h_u_cla32_and11319_y0;
  wire h_u_cla32_and11320_y0;
  wire h_u_cla32_and11321_y0;
  wire h_u_cla32_and11322_y0;
  wire h_u_cla32_and11323_y0;
  wire h_u_cla32_and11324_y0;
  wire h_u_cla32_and11325_y0;
  wire h_u_cla32_and11326_y0;
  wire h_u_cla32_and11327_y0;
  wire h_u_cla32_and11328_y0;
  wire h_u_cla32_and11329_y0;
  wire h_u_cla32_and11330_y0;
  wire h_u_cla32_and11331_y0;
  wire h_u_cla32_and11332_y0;
  wire h_u_cla32_and11333_y0;
  wire h_u_cla32_and11334_y0;
  wire h_u_cla32_and11335_y0;
  wire h_u_cla32_and11336_y0;
  wire h_u_cla32_and11337_y0;
  wire h_u_cla32_and11338_y0;
  wire h_u_cla32_and11339_y0;
  wire h_u_cla32_and11340_y0;
  wire h_u_cla32_and11341_y0;
  wire h_u_cla32_and11342_y0;
  wire h_u_cla32_and11343_y0;
  wire h_u_cla32_and11344_y0;
  wire h_u_cla32_and11345_y0;
  wire h_u_cla32_and11346_y0;
  wire h_u_cla32_and11347_y0;
  wire h_u_cla32_and11348_y0;
  wire h_u_cla32_and11349_y0;
  wire h_u_cla32_and11350_y0;
  wire h_u_cla32_and11351_y0;
  wire h_u_cla32_and11352_y0;
  wire h_u_cla32_and11353_y0;
  wire h_u_cla32_and11354_y0;
  wire h_u_cla32_and11355_y0;
  wire h_u_cla32_and11356_y0;
  wire h_u_cla32_and11357_y0;
  wire h_u_cla32_and11358_y0;
  wire h_u_cla32_and11359_y0;
  wire h_u_cla32_and11360_y0;
  wire h_u_cla32_and11361_y0;
  wire h_u_cla32_and11362_y0;
  wire h_u_cla32_and11363_y0;
  wire h_u_cla32_and11364_y0;
  wire h_u_cla32_and11365_y0;
  wire h_u_cla32_and11366_y0;
  wire h_u_cla32_and11367_y0;
  wire h_u_cla32_and11368_y0;
  wire h_u_cla32_and11369_y0;
  wire h_u_cla32_and11370_y0;
  wire h_u_cla32_and11371_y0;
  wire h_u_cla32_and11372_y0;
  wire h_u_cla32_and11373_y0;
  wire h_u_cla32_and11374_y0;
  wire h_u_cla32_and11375_y0;
  wire h_u_cla32_and11376_y0;
  wire h_u_cla32_and11377_y0;
  wire h_u_cla32_and11378_y0;
  wire h_u_cla32_and11379_y0;
  wire h_u_cla32_and11380_y0;
  wire h_u_cla32_and11381_y0;
  wire h_u_cla32_and11382_y0;
  wire h_u_cla32_and11383_y0;
  wire h_u_cla32_and11384_y0;
  wire h_u_cla32_and11385_y0;
  wire h_u_cla32_and11386_y0;
  wire h_u_cla32_and11387_y0;
  wire h_u_cla32_and11388_y0;
  wire h_u_cla32_and11389_y0;
  wire h_u_cla32_and11390_y0;
  wire h_u_cla32_and11391_y0;
  wire h_u_cla32_and11392_y0;
  wire h_u_cla32_and11393_y0;
  wire h_u_cla32_and11394_y0;
  wire h_u_cla32_and11395_y0;
  wire h_u_cla32_and11396_y0;
  wire h_u_cla32_and11397_y0;
  wire h_u_cla32_and11398_y0;
  wire h_u_cla32_and11399_y0;
  wire h_u_cla32_and11400_y0;
  wire h_u_cla32_and11401_y0;
  wire h_u_cla32_and11402_y0;
  wire h_u_cla32_and11403_y0;
  wire h_u_cla32_and11404_y0;
  wire h_u_cla32_and11405_y0;
  wire h_u_cla32_and11406_y0;
  wire h_u_cla32_and11407_y0;
  wire h_u_cla32_and11408_y0;
  wire h_u_cla32_and11409_y0;
  wire h_u_cla32_and11410_y0;
  wire h_u_cla32_and11411_y0;
  wire h_u_cla32_and11412_y0;
  wire h_u_cla32_and11413_y0;
  wire h_u_cla32_and11414_y0;
  wire h_u_cla32_and11415_y0;
  wire h_u_cla32_and11416_y0;
  wire h_u_cla32_and11417_y0;
  wire h_u_cla32_and11418_y0;
  wire h_u_cla32_and11419_y0;
  wire h_u_cla32_and11420_y0;
  wire h_u_cla32_and11421_y0;
  wire h_u_cla32_and11422_y0;
  wire h_u_cla32_and11423_y0;
  wire h_u_cla32_and11424_y0;
  wire h_u_cla32_and11425_y0;
  wire h_u_cla32_and11426_y0;
  wire h_u_cla32_and11427_y0;
  wire h_u_cla32_and11428_y0;
  wire h_u_cla32_and11429_y0;
  wire h_u_cla32_and11430_y0;
  wire h_u_cla32_and11431_y0;
  wire h_u_cla32_and11432_y0;
  wire h_u_cla32_and11433_y0;
  wire h_u_cla32_and11434_y0;
  wire h_u_cla32_and11435_y0;
  wire h_u_cla32_and11436_y0;
  wire h_u_cla32_and11437_y0;
  wire h_u_cla32_and11438_y0;
  wire h_u_cla32_and11439_y0;
  wire h_u_cla32_or496_y0;
  wire h_u_cla32_or497_y0;
  wire h_u_cla32_or498_y0;
  wire h_u_cla32_or499_y0;
  wire h_u_cla32_or500_y0;
  wire h_u_cla32_or501_y0;
  wire h_u_cla32_or502_y0;
  wire h_u_cla32_or503_y0;
  wire h_u_cla32_or504_y0;
  wire h_u_cla32_or505_y0;
  wire h_u_cla32_or506_y0;
  wire h_u_cla32_or507_y0;
  wire h_u_cla32_or508_y0;
  wire h_u_cla32_or509_y0;
  wire h_u_cla32_or510_y0;
  wire h_u_cla32_or511_y0;
  wire h_u_cla32_or512_y0;
  wire h_u_cla32_or513_y0;
  wire h_u_cla32_or514_y0;
  wire h_u_cla32_or515_y0;
  wire h_u_cla32_or516_y0;
  wire h_u_cla32_or517_y0;
  wire h_u_cla32_or518_y0;
  wire h_u_cla32_or519_y0;
  wire h_u_cla32_or520_y0;
  wire h_u_cla32_or521_y0;
  wire h_u_cla32_or522_y0;
  wire h_u_cla32_or523_y0;
  wire h_u_cla32_or524_y0;
  wire h_u_cla32_or525_y0;
  wire h_u_cla32_or526_y0;
  wire h_u_cla32_or527_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign a_30 = a[30];
  assign a_31 = a[31];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  assign b_30 = b[30];
  assign b_31 = b[31];
  constant_wire_value_0 constant_wire_value_0_constant_wire_0(a_0, b_0, constant_wire_0);
  pg_logic pg_logic_h_u_cla32_pg_logic0_y0(a_0, b_0, h_u_cla32_pg_logic0_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_pg_logic0_y2);
  xor_gate xor_gate_h_u_cla32_xor0_y0(h_u_cla32_pg_logic0_y2, constant_wire_0, h_u_cla32_xor0_y0);
  and_gate and_gate_h_u_cla32_and0_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and0_y0);
  or_gate or_gate_h_u_cla32_or0_y0(h_u_cla32_pg_logic0_y1, h_u_cla32_and0_y0, h_u_cla32_or0_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic1_y0(a_1, b_1, h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_pg_logic1_y2);
  xor_gate xor_gate_h_u_cla32_xor1_y0(h_u_cla32_pg_logic1_y2, h_u_cla32_or0_y0, h_u_cla32_xor1_y0);
  and_gate and_gate_h_u_cla32_and1_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and1_y0);
  and_gate and_gate_h_u_cla32_and2_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and2_y0);
  and_gate and_gate_h_u_cla32_and3_y0(h_u_cla32_and2_y0, h_u_cla32_and1_y0, h_u_cla32_and3_y0);
  and_gate and_gate_h_u_cla32_and4_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4_y0);
  or_gate or_gate_h_u_cla32_or1_y0(h_u_cla32_and4_y0, h_u_cla32_and3_y0, h_u_cla32_or1_y0);
  or_gate or_gate_h_u_cla32_or2_y0(h_u_cla32_pg_logic1_y1, h_u_cla32_or1_y0, h_u_cla32_or2_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic2_y0(a_2, b_2, h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_pg_logic2_y2);
  xor_gate xor_gate_h_u_cla32_xor2_y0(h_u_cla32_pg_logic2_y2, h_u_cla32_or2_y0, h_u_cla32_xor2_y0);
  and_gate and_gate_h_u_cla32_and5_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and5_y0);
  and_gate and_gate_h_u_cla32_and6_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and6_y0);
  and_gate and_gate_h_u_cla32_and7_y0(h_u_cla32_and6_y0, h_u_cla32_and5_y0, h_u_cla32_and7_y0);
  and_gate and_gate_h_u_cla32_and8_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and8_y0);
  and_gate and_gate_h_u_cla32_and9_y0(h_u_cla32_and8_y0, h_u_cla32_and7_y0, h_u_cla32_and9_y0);
  and_gate and_gate_h_u_cla32_and10_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10_y0);
  and_gate and_gate_h_u_cla32_and11_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and11_y0);
  and_gate and_gate_h_u_cla32_and12_y0(h_u_cla32_and11_y0, h_u_cla32_and10_y0, h_u_cla32_and12_y0);
  and_gate and_gate_h_u_cla32_and13_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and13_y0);
  or_gate or_gate_h_u_cla32_or3_y0(h_u_cla32_and13_y0, h_u_cla32_and9_y0, h_u_cla32_or3_y0);
  or_gate or_gate_h_u_cla32_or4_y0(h_u_cla32_or3_y0, h_u_cla32_and12_y0, h_u_cla32_or4_y0);
  or_gate or_gate_h_u_cla32_or5_y0(h_u_cla32_pg_logic2_y1, h_u_cla32_or4_y0, h_u_cla32_or5_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic3_y0(a_3, b_3, h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_pg_logic3_y2);
  xor_gate xor_gate_h_u_cla32_xor3_y0(h_u_cla32_pg_logic3_y2, h_u_cla32_or5_y0, h_u_cla32_xor3_y0);
  and_gate and_gate_h_u_cla32_and14_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and14_y0);
  and_gate and_gate_h_u_cla32_and15_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and15_y0);
  and_gate and_gate_h_u_cla32_and16_y0(h_u_cla32_and15_y0, h_u_cla32_and14_y0, h_u_cla32_and16_y0);
  and_gate and_gate_h_u_cla32_and17_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and17_y0);
  and_gate and_gate_h_u_cla32_and18_y0(h_u_cla32_and17_y0, h_u_cla32_and16_y0, h_u_cla32_and18_y0);
  and_gate and_gate_h_u_cla32_and19_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and19_y0);
  and_gate and_gate_h_u_cla32_and20_y0(h_u_cla32_and19_y0, h_u_cla32_and18_y0, h_u_cla32_and20_y0);
  and_gate and_gate_h_u_cla32_and21_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and21_y0);
  and_gate and_gate_h_u_cla32_and22_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and22_y0);
  and_gate and_gate_h_u_cla32_and23_y0(h_u_cla32_and22_y0, h_u_cla32_and21_y0, h_u_cla32_and23_y0);
  and_gate and_gate_h_u_cla32_and24_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and24_y0);
  and_gate and_gate_h_u_cla32_and25_y0(h_u_cla32_and24_y0, h_u_cla32_and23_y0, h_u_cla32_and25_y0);
  and_gate and_gate_h_u_cla32_and26_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and26_y0);
  and_gate and_gate_h_u_cla32_and27_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and27_y0);
  and_gate and_gate_h_u_cla32_and28_y0(h_u_cla32_and27_y0, h_u_cla32_and26_y0, h_u_cla32_and28_y0);
  and_gate and_gate_h_u_cla32_and29_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and29_y0);
  or_gate or_gate_h_u_cla32_or6_y0(h_u_cla32_and29_y0, h_u_cla32_and20_y0, h_u_cla32_or6_y0);
  or_gate or_gate_h_u_cla32_or7_y0(h_u_cla32_or6_y0, h_u_cla32_and25_y0, h_u_cla32_or7_y0);
  or_gate or_gate_h_u_cla32_or8_y0(h_u_cla32_or7_y0, h_u_cla32_and28_y0, h_u_cla32_or8_y0);
  or_gate or_gate_h_u_cla32_or9_y0(h_u_cla32_pg_logic3_y1, h_u_cla32_or8_y0, h_u_cla32_or9_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic4_y0(a_4, b_4, h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_pg_logic4_y2);
  xor_gate xor_gate_h_u_cla32_xor4_y0(h_u_cla32_pg_logic4_y2, h_u_cla32_or9_y0, h_u_cla32_xor4_y0);
  and_gate and_gate_h_u_cla32_and30_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and30_y0);
  and_gate and_gate_h_u_cla32_and31_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and31_y0);
  and_gate and_gate_h_u_cla32_and32_y0(h_u_cla32_and31_y0, h_u_cla32_and30_y0, h_u_cla32_and32_y0);
  and_gate and_gate_h_u_cla32_and33_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and33_y0);
  and_gate and_gate_h_u_cla32_and34_y0(h_u_cla32_and33_y0, h_u_cla32_and32_y0, h_u_cla32_and34_y0);
  and_gate and_gate_h_u_cla32_and35_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and35_y0);
  and_gate and_gate_h_u_cla32_and36_y0(h_u_cla32_and35_y0, h_u_cla32_and34_y0, h_u_cla32_and36_y0);
  and_gate and_gate_h_u_cla32_and37_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and37_y0);
  and_gate and_gate_h_u_cla32_and38_y0(h_u_cla32_and37_y0, h_u_cla32_and36_y0, h_u_cla32_and38_y0);
  and_gate and_gate_h_u_cla32_and39_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and39_y0);
  and_gate and_gate_h_u_cla32_and40_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and40_y0);
  and_gate and_gate_h_u_cla32_and41_y0(h_u_cla32_and40_y0, h_u_cla32_and39_y0, h_u_cla32_and41_y0);
  and_gate and_gate_h_u_cla32_and42_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and42_y0);
  and_gate and_gate_h_u_cla32_and43_y0(h_u_cla32_and42_y0, h_u_cla32_and41_y0, h_u_cla32_and43_y0);
  and_gate and_gate_h_u_cla32_and44_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and44_y0);
  and_gate and_gate_h_u_cla32_and45_y0(h_u_cla32_and44_y0, h_u_cla32_and43_y0, h_u_cla32_and45_y0);
  and_gate and_gate_h_u_cla32_and46_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and46_y0);
  and_gate and_gate_h_u_cla32_and47_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and47_y0);
  and_gate and_gate_h_u_cla32_and48_y0(h_u_cla32_and47_y0, h_u_cla32_and46_y0, h_u_cla32_and48_y0);
  and_gate and_gate_h_u_cla32_and49_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and49_y0);
  and_gate and_gate_h_u_cla32_and50_y0(h_u_cla32_and49_y0, h_u_cla32_and48_y0, h_u_cla32_and50_y0);
  and_gate and_gate_h_u_cla32_and51_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and51_y0);
  and_gate and_gate_h_u_cla32_and52_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and52_y0);
  and_gate and_gate_h_u_cla32_and53_y0(h_u_cla32_and52_y0, h_u_cla32_and51_y0, h_u_cla32_and53_y0);
  and_gate and_gate_h_u_cla32_and54_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and54_y0);
  or_gate or_gate_h_u_cla32_or10_y0(h_u_cla32_and54_y0, h_u_cla32_and38_y0, h_u_cla32_or10_y0);
  or_gate or_gate_h_u_cla32_or11_y0(h_u_cla32_or10_y0, h_u_cla32_and45_y0, h_u_cla32_or11_y0);
  or_gate or_gate_h_u_cla32_or12_y0(h_u_cla32_or11_y0, h_u_cla32_and50_y0, h_u_cla32_or12_y0);
  or_gate or_gate_h_u_cla32_or13_y0(h_u_cla32_or12_y0, h_u_cla32_and53_y0, h_u_cla32_or13_y0);
  or_gate or_gate_h_u_cla32_or14_y0(h_u_cla32_pg_logic4_y1, h_u_cla32_or13_y0, h_u_cla32_or14_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic5_y0(a_5, b_5, h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_pg_logic5_y2);
  xor_gate xor_gate_h_u_cla32_xor5_y0(h_u_cla32_pg_logic5_y2, h_u_cla32_or14_y0, h_u_cla32_xor5_y0);
  and_gate and_gate_h_u_cla32_and55_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and55_y0);
  and_gate and_gate_h_u_cla32_and56_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and56_y0);
  and_gate and_gate_h_u_cla32_and57_y0(h_u_cla32_and56_y0, h_u_cla32_and55_y0, h_u_cla32_and57_y0);
  and_gate and_gate_h_u_cla32_and58_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and58_y0);
  and_gate and_gate_h_u_cla32_and59_y0(h_u_cla32_and58_y0, h_u_cla32_and57_y0, h_u_cla32_and59_y0);
  and_gate and_gate_h_u_cla32_and60_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and60_y0);
  and_gate and_gate_h_u_cla32_and61_y0(h_u_cla32_and60_y0, h_u_cla32_and59_y0, h_u_cla32_and61_y0);
  and_gate and_gate_h_u_cla32_and62_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and62_y0);
  and_gate and_gate_h_u_cla32_and63_y0(h_u_cla32_and62_y0, h_u_cla32_and61_y0, h_u_cla32_and63_y0);
  and_gate and_gate_h_u_cla32_and64_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and64_y0);
  and_gate and_gate_h_u_cla32_and65_y0(h_u_cla32_and64_y0, h_u_cla32_and63_y0, h_u_cla32_and65_y0);
  and_gate and_gate_h_u_cla32_and66_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and66_y0);
  and_gate and_gate_h_u_cla32_and67_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and67_y0);
  and_gate and_gate_h_u_cla32_and68_y0(h_u_cla32_and67_y0, h_u_cla32_and66_y0, h_u_cla32_and68_y0);
  and_gate and_gate_h_u_cla32_and69_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and69_y0);
  and_gate and_gate_h_u_cla32_and70_y0(h_u_cla32_and69_y0, h_u_cla32_and68_y0, h_u_cla32_and70_y0);
  and_gate and_gate_h_u_cla32_and71_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and71_y0);
  and_gate and_gate_h_u_cla32_and72_y0(h_u_cla32_and71_y0, h_u_cla32_and70_y0, h_u_cla32_and72_y0);
  and_gate and_gate_h_u_cla32_and73_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and73_y0);
  and_gate and_gate_h_u_cla32_and74_y0(h_u_cla32_and73_y0, h_u_cla32_and72_y0, h_u_cla32_and74_y0);
  and_gate and_gate_h_u_cla32_and75_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and75_y0);
  and_gate and_gate_h_u_cla32_and76_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and76_y0);
  and_gate and_gate_h_u_cla32_and77_y0(h_u_cla32_and76_y0, h_u_cla32_and75_y0, h_u_cla32_and77_y0);
  and_gate and_gate_h_u_cla32_and78_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and78_y0);
  and_gate and_gate_h_u_cla32_and79_y0(h_u_cla32_and78_y0, h_u_cla32_and77_y0, h_u_cla32_and79_y0);
  and_gate and_gate_h_u_cla32_and80_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and80_y0);
  and_gate and_gate_h_u_cla32_and81_y0(h_u_cla32_and80_y0, h_u_cla32_and79_y0, h_u_cla32_and81_y0);
  and_gate and_gate_h_u_cla32_and82_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and82_y0);
  and_gate and_gate_h_u_cla32_and83_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and83_y0);
  and_gate and_gate_h_u_cla32_and84_y0(h_u_cla32_and83_y0, h_u_cla32_and82_y0, h_u_cla32_and84_y0);
  and_gate and_gate_h_u_cla32_and85_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and85_y0);
  and_gate and_gate_h_u_cla32_and86_y0(h_u_cla32_and85_y0, h_u_cla32_and84_y0, h_u_cla32_and86_y0);
  and_gate and_gate_h_u_cla32_and87_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and87_y0);
  and_gate and_gate_h_u_cla32_and88_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and88_y0);
  and_gate and_gate_h_u_cla32_and89_y0(h_u_cla32_and88_y0, h_u_cla32_and87_y0, h_u_cla32_and89_y0);
  and_gate and_gate_h_u_cla32_and90_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and90_y0);
  or_gate or_gate_h_u_cla32_or15_y0(h_u_cla32_and90_y0, h_u_cla32_and65_y0, h_u_cla32_or15_y0);
  or_gate or_gate_h_u_cla32_or16_y0(h_u_cla32_or15_y0, h_u_cla32_and74_y0, h_u_cla32_or16_y0);
  or_gate or_gate_h_u_cla32_or17_y0(h_u_cla32_or16_y0, h_u_cla32_and81_y0, h_u_cla32_or17_y0);
  or_gate or_gate_h_u_cla32_or18_y0(h_u_cla32_or17_y0, h_u_cla32_and86_y0, h_u_cla32_or18_y0);
  or_gate or_gate_h_u_cla32_or19_y0(h_u_cla32_or18_y0, h_u_cla32_and89_y0, h_u_cla32_or19_y0);
  or_gate or_gate_h_u_cla32_or20_y0(h_u_cla32_pg_logic5_y1, h_u_cla32_or19_y0, h_u_cla32_or20_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic6_y0(a_6, b_6, h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_pg_logic6_y2);
  xor_gate xor_gate_h_u_cla32_xor6_y0(h_u_cla32_pg_logic6_y2, h_u_cla32_or20_y0, h_u_cla32_xor6_y0);
  and_gate and_gate_h_u_cla32_and91_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and91_y0);
  and_gate and_gate_h_u_cla32_and92_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and92_y0);
  and_gate and_gate_h_u_cla32_and93_y0(h_u_cla32_and92_y0, h_u_cla32_and91_y0, h_u_cla32_and93_y0);
  and_gate and_gate_h_u_cla32_and94_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and94_y0);
  and_gate and_gate_h_u_cla32_and95_y0(h_u_cla32_and94_y0, h_u_cla32_and93_y0, h_u_cla32_and95_y0);
  and_gate and_gate_h_u_cla32_and96_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and96_y0);
  and_gate and_gate_h_u_cla32_and97_y0(h_u_cla32_and96_y0, h_u_cla32_and95_y0, h_u_cla32_and97_y0);
  and_gate and_gate_h_u_cla32_and98_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and98_y0);
  and_gate and_gate_h_u_cla32_and99_y0(h_u_cla32_and98_y0, h_u_cla32_and97_y0, h_u_cla32_and99_y0);
  and_gate and_gate_h_u_cla32_and100_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and100_y0);
  and_gate and_gate_h_u_cla32_and101_y0(h_u_cla32_and100_y0, h_u_cla32_and99_y0, h_u_cla32_and101_y0);
  and_gate and_gate_h_u_cla32_and102_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and102_y0);
  and_gate and_gate_h_u_cla32_and103_y0(h_u_cla32_and102_y0, h_u_cla32_and101_y0, h_u_cla32_and103_y0);
  and_gate and_gate_h_u_cla32_and104_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and104_y0);
  and_gate and_gate_h_u_cla32_and105_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and105_y0);
  and_gate and_gate_h_u_cla32_and106_y0(h_u_cla32_and105_y0, h_u_cla32_and104_y0, h_u_cla32_and106_y0);
  and_gate and_gate_h_u_cla32_and107_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and107_y0);
  and_gate and_gate_h_u_cla32_and108_y0(h_u_cla32_and107_y0, h_u_cla32_and106_y0, h_u_cla32_and108_y0);
  and_gate and_gate_h_u_cla32_and109_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and109_y0);
  and_gate and_gate_h_u_cla32_and110_y0(h_u_cla32_and109_y0, h_u_cla32_and108_y0, h_u_cla32_and110_y0);
  and_gate and_gate_h_u_cla32_and111_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and111_y0);
  and_gate and_gate_h_u_cla32_and112_y0(h_u_cla32_and111_y0, h_u_cla32_and110_y0, h_u_cla32_and112_y0);
  and_gate and_gate_h_u_cla32_and113_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and113_y0);
  and_gate and_gate_h_u_cla32_and114_y0(h_u_cla32_and113_y0, h_u_cla32_and112_y0, h_u_cla32_and114_y0);
  and_gate and_gate_h_u_cla32_and115_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and115_y0);
  and_gate and_gate_h_u_cla32_and116_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and116_y0);
  and_gate and_gate_h_u_cla32_and117_y0(h_u_cla32_and116_y0, h_u_cla32_and115_y0, h_u_cla32_and117_y0);
  and_gate and_gate_h_u_cla32_and118_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and118_y0);
  and_gate and_gate_h_u_cla32_and119_y0(h_u_cla32_and118_y0, h_u_cla32_and117_y0, h_u_cla32_and119_y0);
  and_gate and_gate_h_u_cla32_and120_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and120_y0);
  and_gate and_gate_h_u_cla32_and121_y0(h_u_cla32_and120_y0, h_u_cla32_and119_y0, h_u_cla32_and121_y0);
  and_gate and_gate_h_u_cla32_and122_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and122_y0);
  and_gate and_gate_h_u_cla32_and123_y0(h_u_cla32_and122_y0, h_u_cla32_and121_y0, h_u_cla32_and123_y0);
  and_gate and_gate_h_u_cla32_and124_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and124_y0);
  and_gate and_gate_h_u_cla32_and125_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and125_y0);
  and_gate and_gate_h_u_cla32_and126_y0(h_u_cla32_and125_y0, h_u_cla32_and124_y0, h_u_cla32_and126_y0);
  and_gate and_gate_h_u_cla32_and127_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and127_y0);
  and_gate and_gate_h_u_cla32_and128_y0(h_u_cla32_and127_y0, h_u_cla32_and126_y0, h_u_cla32_and128_y0);
  and_gate and_gate_h_u_cla32_and129_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and129_y0);
  and_gate and_gate_h_u_cla32_and130_y0(h_u_cla32_and129_y0, h_u_cla32_and128_y0, h_u_cla32_and130_y0);
  and_gate and_gate_h_u_cla32_and131_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and131_y0);
  and_gate and_gate_h_u_cla32_and132_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and132_y0);
  and_gate and_gate_h_u_cla32_and133_y0(h_u_cla32_and132_y0, h_u_cla32_and131_y0, h_u_cla32_and133_y0);
  and_gate and_gate_h_u_cla32_and134_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and134_y0);
  and_gate and_gate_h_u_cla32_and135_y0(h_u_cla32_and134_y0, h_u_cla32_and133_y0, h_u_cla32_and135_y0);
  and_gate and_gate_h_u_cla32_and136_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and136_y0);
  and_gate and_gate_h_u_cla32_and137_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and137_y0);
  and_gate and_gate_h_u_cla32_and138_y0(h_u_cla32_and137_y0, h_u_cla32_and136_y0, h_u_cla32_and138_y0);
  and_gate and_gate_h_u_cla32_and139_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and139_y0);
  or_gate or_gate_h_u_cla32_or21_y0(h_u_cla32_and139_y0, h_u_cla32_and103_y0, h_u_cla32_or21_y0);
  or_gate or_gate_h_u_cla32_or22_y0(h_u_cla32_or21_y0, h_u_cla32_and114_y0, h_u_cla32_or22_y0);
  or_gate or_gate_h_u_cla32_or23_y0(h_u_cla32_or22_y0, h_u_cla32_and123_y0, h_u_cla32_or23_y0);
  or_gate or_gate_h_u_cla32_or24_y0(h_u_cla32_or23_y0, h_u_cla32_and130_y0, h_u_cla32_or24_y0);
  or_gate or_gate_h_u_cla32_or25_y0(h_u_cla32_or24_y0, h_u_cla32_and135_y0, h_u_cla32_or25_y0);
  or_gate or_gate_h_u_cla32_or26_y0(h_u_cla32_or25_y0, h_u_cla32_and138_y0, h_u_cla32_or26_y0);
  or_gate or_gate_h_u_cla32_or27_y0(h_u_cla32_pg_logic6_y1, h_u_cla32_or26_y0, h_u_cla32_or27_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic7_y0(a_7, b_7, h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_pg_logic7_y2);
  xor_gate xor_gate_h_u_cla32_xor7_y0(h_u_cla32_pg_logic7_y2, h_u_cla32_or27_y0, h_u_cla32_xor7_y0);
  and_gate and_gate_h_u_cla32_and140_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and140_y0);
  and_gate and_gate_h_u_cla32_and141_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and141_y0);
  and_gate and_gate_h_u_cla32_and142_y0(h_u_cla32_and141_y0, h_u_cla32_and140_y0, h_u_cla32_and142_y0);
  and_gate and_gate_h_u_cla32_and143_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and143_y0);
  and_gate and_gate_h_u_cla32_and144_y0(h_u_cla32_and143_y0, h_u_cla32_and142_y0, h_u_cla32_and144_y0);
  and_gate and_gate_h_u_cla32_and145_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and145_y0);
  and_gate and_gate_h_u_cla32_and146_y0(h_u_cla32_and145_y0, h_u_cla32_and144_y0, h_u_cla32_and146_y0);
  and_gate and_gate_h_u_cla32_and147_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and147_y0);
  and_gate and_gate_h_u_cla32_and148_y0(h_u_cla32_and147_y0, h_u_cla32_and146_y0, h_u_cla32_and148_y0);
  and_gate and_gate_h_u_cla32_and149_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and149_y0);
  and_gate and_gate_h_u_cla32_and150_y0(h_u_cla32_and149_y0, h_u_cla32_and148_y0, h_u_cla32_and150_y0);
  and_gate and_gate_h_u_cla32_and151_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and151_y0);
  and_gate and_gate_h_u_cla32_and152_y0(h_u_cla32_and151_y0, h_u_cla32_and150_y0, h_u_cla32_and152_y0);
  and_gate and_gate_h_u_cla32_and153_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and153_y0);
  and_gate and_gate_h_u_cla32_and154_y0(h_u_cla32_and153_y0, h_u_cla32_and152_y0, h_u_cla32_and154_y0);
  and_gate and_gate_h_u_cla32_and155_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and155_y0);
  and_gate and_gate_h_u_cla32_and156_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and156_y0);
  and_gate and_gate_h_u_cla32_and157_y0(h_u_cla32_and156_y0, h_u_cla32_and155_y0, h_u_cla32_and157_y0);
  and_gate and_gate_h_u_cla32_and158_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and158_y0);
  and_gate and_gate_h_u_cla32_and159_y0(h_u_cla32_and158_y0, h_u_cla32_and157_y0, h_u_cla32_and159_y0);
  and_gate and_gate_h_u_cla32_and160_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and160_y0);
  and_gate and_gate_h_u_cla32_and161_y0(h_u_cla32_and160_y0, h_u_cla32_and159_y0, h_u_cla32_and161_y0);
  and_gate and_gate_h_u_cla32_and162_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and162_y0);
  and_gate and_gate_h_u_cla32_and163_y0(h_u_cla32_and162_y0, h_u_cla32_and161_y0, h_u_cla32_and163_y0);
  and_gate and_gate_h_u_cla32_and164_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and164_y0);
  and_gate and_gate_h_u_cla32_and165_y0(h_u_cla32_and164_y0, h_u_cla32_and163_y0, h_u_cla32_and165_y0);
  and_gate and_gate_h_u_cla32_and166_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and166_y0);
  and_gate and_gate_h_u_cla32_and167_y0(h_u_cla32_and166_y0, h_u_cla32_and165_y0, h_u_cla32_and167_y0);
  and_gate and_gate_h_u_cla32_and168_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and168_y0);
  and_gate and_gate_h_u_cla32_and169_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and169_y0);
  and_gate and_gate_h_u_cla32_and170_y0(h_u_cla32_and169_y0, h_u_cla32_and168_y0, h_u_cla32_and170_y0);
  and_gate and_gate_h_u_cla32_and171_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and171_y0);
  and_gate and_gate_h_u_cla32_and172_y0(h_u_cla32_and171_y0, h_u_cla32_and170_y0, h_u_cla32_and172_y0);
  and_gate and_gate_h_u_cla32_and173_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and173_y0);
  and_gate and_gate_h_u_cla32_and174_y0(h_u_cla32_and173_y0, h_u_cla32_and172_y0, h_u_cla32_and174_y0);
  and_gate and_gate_h_u_cla32_and175_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and175_y0);
  and_gate and_gate_h_u_cla32_and176_y0(h_u_cla32_and175_y0, h_u_cla32_and174_y0, h_u_cla32_and176_y0);
  and_gate and_gate_h_u_cla32_and177_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and177_y0);
  and_gate and_gate_h_u_cla32_and178_y0(h_u_cla32_and177_y0, h_u_cla32_and176_y0, h_u_cla32_and178_y0);
  and_gate and_gate_h_u_cla32_and179_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and179_y0);
  and_gate and_gate_h_u_cla32_and180_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and180_y0);
  and_gate and_gate_h_u_cla32_and181_y0(h_u_cla32_and180_y0, h_u_cla32_and179_y0, h_u_cla32_and181_y0);
  and_gate and_gate_h_u_cla32_and182_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and182_y0);
  and_gate and_gate_h_u_cla32_and183_y0(h_u_cla32_and182_y0, h_u_cla32_and181_y0, h_u_cla32_and183_y0);
  and_gate and_gate_h_u_cla32_and184_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and184_y0);
  and_gate and_gate_h_u_cla32_and185_y0(h_u_cla32_and184_y0, h_u_cla32_and183_y0, h_u_cla32_and185_y0);
  and_gate and_gate_h_u_cla32_and186_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and186_y0);
  and_gate and_gate_h_u_cla32_and187_y0(h_u_cla32_and186_y0, h_u_cla32_and185_y0, h_u_cla32_and187_y0);
  and_gate and_gate_h_u_cla32_and188_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and188_y0);
  and_gate and_gate_h_u_cla32_and189_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and189_y0);
  and_gate and_gate_h_u_cla32_and190_y0(h_u_cla32_and189_y0, h_u_cla32_and188_y0, h_u_cla32_and190_y0);
  and_gate and_gate_h_u_cla32_and191_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and191_y0);
  and_gate and_gate_h_u_cla32_and192_y0(h_u_cla32_and191_y0, h_u_cla32_and190_y0, h_u_cla32_and192_y0);
  and_gate and_gate_h_u_cla32_and193_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and193_y0);
  and_gate and_gate_h_u_cla32_and194_y0(h_u_cla32_and193_y0, h_u_cla32_and192_y0, h_u_cla32_and194_y0);
  and_gate and_gate_h_u_cla32_and195_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and195_y0);
  and_gate and_gate_h_u_cla32_and196_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and196_y0);
  and_gate and_gate_h_u_cla32_and197_y0(h_u_cla32_and196_y0, h_u_cla32_and195_y0, h_u_cla32_and197_y0);
  and_gate and_gate_h_u_cla32_and198_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and198_y0);
  and_gate and_gate_h_u_cla32_and199_y0(h_u_cla32_and198_y0, h_u_cla32_and197_y0, h_u_cla32_and199_y0);
  and_gate and_gate_h_u_cla32_and200_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and200_y0);
  and_gate and_gate_h_u_cla32_and201_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and201_y0);
  and_gate and_gate_h_u_cla32_and202_y0(h_u_cla32_and201_y0, h_u_cla32_and200_y0, h_u_cla32_and202_y0);
  and_gate and_gate_h_u_cla32_and203_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and203_y0);
  or_gate or_gate_h_u_cla32_or28_y0(h_u_cla32_and203_y0, h_u_cla32_and154_y0, h_u_cla32_or28_y0);
  or_gate or_gate_h_u_cla32_or29_y0(h_u_cla32_or28_y0, h_u_cla32_and167_y0, h_u_cla32_or29_y0);
  or_gate or_gate_h_u_cla32_or30_y0(h_u_cla32_or29_y0, h_u_cla32_and178_y0, h_u_cla32_or30_y0);
  or_gate or_gate_h_u_cla32_or31_y0(h_u_cla32_or30_y0, h_u_cla32_and187_y0, h_u_cla32_or31_y0);
  or_gate or_gate_h_u_cla32_or32_y0(h_u_cla32_or31_y0, h_u_cla32_and194_y0, h_u_cla32_or32_y0);
  or_gate or_gate_h_u_cla32_or33_y0(h_u_cla32_or32_y0, h_u_cla32_and199_y0, h_u_cla32_or33_y0);
  or_gate or_gate_h_u_cla32_or34_y0(h_u_cla32_or33_y0, h_u_cla32_and202_y0, h_u_cla32_or34_y0);
  or_gate or_gate_h_u_cla32_or35_y0(h_u_cla32_pg_logic7_y1, h_u_cla32_or34_y0, h_u_cla32_or35_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic8_y0(a_8, b_8, h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_pg_logic8_y2);
  xor_gate xor_gate_h_u_cla32_xor8_y0(h_u_cla32_pg_logic8_y2, h_u_cla32_or35_y0, h_u_cla32_xor8_y0);
  and_gate and_gate_h_u_cla32_and204_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and204_y0);
  and_gate and_gate_h_u_cla32_and205_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and205_y0);
  and_gate and_gate_h_u_cla32_and206_y0(h_u_cla32_and205_y0, h_u_cla32_and204_y0, h_u_cla32_and206_y0);
  and_gate and_gate_h_u_cla32_and207_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and207_y0);
  and_gate and_gate_h_u_cla32_and208_y0(h_u_cla32_and207_y0, h_u_cla32_and206_y0, h_u_cla32_and208_y0);
  and_gate and_gate_h_u_cla32_and209_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and209_y0);
  and_gate and_gate_h_u_cla32_and210_y0(h_u_cla32_and209_y0, h_u_cla32_and208_y0, h_u_cla32_and210_y0);
  and_gate and_gate_h_u_cla32_and211_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and211_y0);
  and_gate and_gate_h_u_cla32_and212_y0(h_u_cla32_and211_y0, h_u_cla32_and210_y0, h_u_cla32_and212_y0);
  and_gate and_gate_h_u_cla32_and213_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and213_y0);
  and_gate and_gate_h_u_cla32_and214_y0(h_u_cla32_and213_y0, h_u_cla32_and212_y0, h_u_cla32_and214_y0);
  and_gate and_gate_h_u_cla32_and215_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and215_y0);
  and_gate and_gate_h_u_cla32_and216_y0(h_u_cla32_and215_y0, h_u_cla32_and214_y0, h_u_cla32_and216_y0);
  and_gate and_gate_h_u_cla32_and217_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and217_y0);
  and_gate and_gate_h_u_cla32_and218_y0(h_u_cla32_and217_y0, h_u_cla32_and216_y0, h_u_cla32_and218_y0);
  and_gate and_gate_h_u_cla32_and219_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and219_y0);
  and_gate and_gate_h_u_cla32_and220_y0(h_u_cla32_and219_y0, h_u_cla32_and218_y0, h_u_cla32_and220_y0);
  and_gate and_gate_h_u_cla32_and221_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and221_y0);
  and_gate and_gate_h_u_cla32_and222_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and222_y0);
  and_gate and_gate_h_u_cla32_and223_y0(h_u_cla32_and222_y0, h_u_cla32_and221_y0, h_u_cla32_and223_y0);
  and_gate and_gate_h_u_cla32_and224_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and224_y0);
  and_gate and_gate_h_u_cla32_and225_y0(h_u_cla32_and224_y0, h_u_cla32_and223_y0, h_u_cla32_and225_y0);
  and_gate and_gate_h_u_cla32_and226_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and226_y0);
  and_gate and_gate_h_u_cla32_and227_y0(h_u_cla32_and226_y0, h_u_cla32_and225_y0, h_u_cla32_and227_y0);
  and_gate and_gate_h_u_cla32_and228_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and228_y0);
  and_gate and_gate_h_u_cla32_and229_y0(h_u_cla32_and228_y0, h_u_cla32_and227_y0, h_u_cla32_and229_y0);
  and_gate and_gate_h_u_cla32_and230_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and230_y0);
  and_gate and_gate_h_u_cla32_and231_y0(h_u_cla32_and230_y0, h_u_cla32_and229_y0, h_u_cla32_and231_y0);
  and_gate and_gate_h_u_cla32_and232_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and232_y0);
  and_gate and_gate_h_u_cla32_and233_y0(h_u_cla32_and232_y0, h_u_cla32_and231_y0, h_u_cla32_and233_y0);
  and_gate and_gate_h_u_cla32_and234_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and234_y0);
  and_gate and_gate_h_u_cla32_and235_y0(h_u_cla32_and234_y0, h_u_cla32_and233_y0, h_u_cla32_and235_y0);
  and_gate and_gate_h_u_cla32_and236_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and236_y0);
  and_gate and_gate_h_u_cla32_and237_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and237_y0);
  and_gate and_gate_h_u_cla32_and238_y0(h_u_cla32_and237_y0, h_u_cla32_and236_y0, h_u_cla32_and238_y0);
  and_gate and_gate_h_u_cla32_and239_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and239_y0);
  and_gate and_gate_h_u_cla32_and240_y0(h_u_cla32_and239_y0, h_u_cla32_and238_y0, h_u_cla32_and240_y0);
  and_gate and_gate_h_u_cla32_and241_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and241_y0);
  and_gate and_gate_h_u_cla32_and242_y0(h_u_cla32_and241_y0, h_u_cla32_and240_y0, h_u_cla32_and242_y0);
  and_gate and_gate_h_u_cla32_and243_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and243_y0);
  and_gate and_gate_h_u_cla32_and244_y0(h_u_cla32_and243_y0, h_u_cla32_and242_y0, h_u_cla32_and244_y0);
  and_gate and_gate_h_u_cla32_and245_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and245_y0);
  and_gate and_gate_h_u_cla32_and246_y0(h_u_cla32_and245_y0, h_u_cla32_and244_y0, h_u_cla32_and246_y0);
  and_gate and_gate_h_u_cla32_and247_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and247_y0);
  and_gate and_gate_h_u_cla32_and248_y0(h_u_cla32_and247_y0, h_u_cla32_and246_y0, h_u_cla32_and248_y0);
  and_gate and_gate_h_u_cla32_and249_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and249_y0);
  and_gate and_gate_h_u_cla32_and250_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and250_y0);
  and_gate and_gate_h_u_cla32_and251_y0(h_u_cla32_and250_y0, h_u_cla32_and249_y0, h_u_cla32_and251_y0);
  and_gate and_gate_h_u_cla32_and252_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and252_y0);
  and_gate and_gate_h_u_cla32_and253_y0(h_u_cla32_and252_y0, h_u_cla32_and251_y0, h_u_cla32_and253_y0);
  and_gate and_gate_h_u_cla32_and254_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and254_y0);
  and_gate and_gate_h_u_cla32_and255_y0(h_u_cla32_and254_y0, h_u_cla32_and253_y0, h_u_cla32_and255_y0);
  and_gate and_gate_h_u_cla32_and256_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and256_y0);
  and_gate and_gate_h_u_cla32_and257_y0(h_u_cla32_and256_y0, h_u_cla32_and255_y0, h_u_cla32_and257_y0);
  and_gate and_gate_h_u_cla32_and258_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and258_y0);
  and_gate and_gate_h_u_cla32_and259_y0(h_u_cla32_and258_y0, h_u_cla32_and257_y0, h_u_cla32_and259_y0);
  and_gate and_gate_h_u_cla32_and260_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and260_y0);
  and_gate and_gate_h_u_cla32_and261_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and261_y0);
  and_gate and_gate_h_u_cla32_and262_y0(h_u_cla32_and261_y0, h_u_cla32_and260_y0, h_u_cla32_and262_y0);
  and_gate and_gate_h_u_cla32_and263_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and263_y0);
  and_gate and_gate_h_u_cla32_and264_y0(h_u_cla32_and263_y0, h_u_cla32_and262_y0, h_u_cla32_and264_y0);
  and_gate and_gate_h_u_cla32_and265_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and265_y0);
  and_gate and_gate_h_u_cla32_and266_y0(h_u_cla32_and265_y0, h_u_cla32_and264_y0, h_u_cla32_and266_y0);
  and_gate and_gate_h_u_cla32_and267_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and267_y0);
  and_gate and_gate_h_u_cla32_and268_y0(h_u_cla32_and267_y0, h_u_cla32_and266_y0, h_u_cla32_and268_y0);
  and_gate and_gate_h_u_cla32_and269_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and269_y0);
  and_gate and_gate_h_u_cla32_and270_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and270_y0);
  and_gate and_gate_h_u_cla32_and271_y0(h_u_cla32_and270_y0, h_u_cla32_and269_y0, h_u_cla32_and271_y0);
  and_gate and_gate_h_u_cla32_and272_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and272_y0);
  and_gate and_gate_h_u_cla32_and273_y0(h_u_cla32_and272_y0, h_u_cla32_and271_y0, h_u_cla32_and273_y0);
  and_gate and_gate_h_u_cla32_and274_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and274_y0);
  and_gate and_gate_h_u_cla32_and275_y0(h_u_cla32_and274_y0, h_u_cla32_and273_y0, h_u_cla32_and275_y0);
  and_gate and_gate_h_u_cla32_and276_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and276_y0);
  and_gate and_gate_h_u_cla32_and277_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and277_y0);
  and_gate and_gate_h_u_cla32_and278_y0(h_u_cla32_and277_y0, h_u_cla32_and276_y0, h_u_cla32_and278_y0);
  and_gate and_gate_h_u_cla32_and279_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and279_y0);
  and_gate and_gate_h_u_cla32_and280_y0(h_u_cla32_and279_y0, h_u_cla32_and278_y0, h_u_cla32_and280_y0);
  and_gate and_gate_h_u_cla32_and281_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and281_y0);
  and_gate and_gate_h_u_cla32_and282_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and282_y0);
  and_gate and_gate_h_u_cla32_and283_y0(h_u_cla32_and282_y0, h_u_cla32_and281_y0, h_u_cla32_and283_y0);
  and_gate and_gate_h_u_cla32_and284_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and284_y0);
  or_gate or_gate_h_u_cla32_or36_y0(h_u_cla32_and284_y0, h_u_cla32_and220_y0, h_u_cla32_or36_y0);
  or_gate or_gate_h_u_cla32_or37_y0(h_u_cla32_or36_y0, h_u_cla32_and235_y0, h_u_cla32_or37_y0);
  or_gate or_gate_h_u_cla32_or38_y0(h_u_cla32_or37_y0, h_u_cla32_and248_y0, h_u_cla32_or38_y0);
  or_gate or_gate_h_u_cla32_or39_y0(h_u_cla32_or38_y0, h_u_cla32_and259_y0, h_u_cla32_or39_y0);
  or_gate or_gate_h_u_cla32_or40_y0(h_u_cla32_or39_y0, h_u_cla32_and268_y0, h_u_cla32_or40_y0);
  or_gate or_gate_h_u_cla32_or41_y0(h_u_cla32_or40_y0, h_u_cla32_and275_y0, h_u_cla32_or41_y0);
  or_gate or_gate_h_u_cla32_or42_y0(h_u_cla32_or41_y0, h_u_cla32_and280_y0, h_u_cla32_or42_y0);
  or_gate or_gate_h_u_cla32_or43_y0(h_u_cla32_or42_y0, h_u_cla32_and283_y0, h_u_cla32_or43_y0);
  or_gate or_gate_h_u_cla32_or44_y0(h_u_cla32_pg_logic8_y1, h_u_cla32_or43_y0, h_u_cla32_or44_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic9_y0(a_9, b_9, h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_pg_logic9_y2);
  xor_gate xor_gate_h_u_cla32_xor9_y0(h_u_cla32_pg_logic9_y2, h_u_cla32_or44_y0, h_u_cla32_xor9_y0);
  and_gate and_gate_h_u_cla32_and285_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and285_y0);
  and_gate and_gate_h_u_cla32_and286_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and286_y0);
  and_gate and_gate_h_u_cla32_and287_y0(h_u_cla32_and286_y0, h_u_cla32_and285_y0, h_u_cla32_and287_y0);
  and_gate and_gate_h_u_cla32_and288_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and288_y0);
  and_gate and_gate_h_u_cla32_and289_y0(h_u_cla32_and288_y0, h_u_cla32_and287_y0, h_u_cla32_and289_y0);
  and_gate and_gate_h_u_cla32_and290_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and290_y0);
  and_gate and_gate_h_u_cla32_and291_y0(h_u_cla32_and290_y0, h_u_cla32_and289_y0, h_u_cla32_and291_y0);
  and_gate and_gate_h_u_cla32_and292_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and292_y0);
  and_gate and_gate_h_u_cla32_and293_y0(h_u_cla32_and292_y0, h_u_cla32_and291_y0, h_u_cla32_and293_y0);
  and_gate and_gate_h_u_cla32_and294_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and294_y0);
  and_gate and_gate_h_u_cla32_and295_y0(h_u_cla32_and294_y0, h_u_cla32_and293_y0, h_u_cla32_and295_y0);
  and_gate and_gate_h_u_cla32_and296_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and296_y0);
  and_gate and_gate_h_u_cla32_and297_y0(h_u_cla32_and296_y0, h_u_cla32_and295_y0, h_u_cla32_and297_y0);
  and_gate and_gate_h_u_cla32_and298_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and298_y0);
  and_gate and_gate_h_u_cla32_and299_y0(h_u_cla32_and298_y0, h_u_cla32_and297_y0, h_u_cla32_and299_y0);
  and_gate and_gate_h_u_cla32_and300_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and300_y0);
  and_gate and_gate_h_u_cla32_and301_y0(h_u_cla32_and300_y0, h_u_cla32_and299_y0, h_u_cla32_and301_y0);
  and_gate and_gate_h_u_cla32_and302_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and302_y0);
  and_gate and_gate_h_u_cla32_and303_y0(h_u_cla32_and302_y0, h_u_cla32_and301_y0, h_u_cla32_and303_y0);
  and_gate and_gate_h_u_cla32_and304_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and304_y0);
  and_gate and_gate_h_u_cla32_and305_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and305_y0);
  and_gate and_gate_h_u_cla32_and306_y0(h_u_cla32_and305_y0, h_u_cla32_and304_y0, h_u_cla32_and306_y0);
  and_gate and_gate_h_u_cla32_and307_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and307_y0);
  and_gate and_gate_h_u_cla32_and308_y0(h_u_cla32_and307_y0, h_u_cla32_and306_y0, h_u_cla32_and308_y0);
  and_gate and_gate_h_u_cla32_and309_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and309_y0);
  and_gate and_gate_h_u_cla32_and310_y0(h_u_cla32_and309_y0, h_u_cla32_and308_y0, h_u_cla32_and310_y0);
  and_gate and_gate_h_u_cla32_and311_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and311_y0);
  and_gate and_gate_h_u_cla32_and312_y0(h_u_cla32_and311_y0, h_u_cla32_and310_y0, h_u_cla32_and312_y0);
  and_gate and_gate_h_u_cla32_and313_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and313_y0);
  and_gate and_gate_h_u_cla32_and314_y0(h_u_cla32_and313_y0, h_u_cla32_and312_y0, h_u_cla32_and314_y0);
  and_gate and_gate_h_u_cla32_and315_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and315_y0);
  and_gate and_gate_h_u_cla32_and316_y0(h_u_cla32_and315_y0, h_u_cla32_and314_y0, h_u_cla32_and316_y0);
  and_gate and_gate_h_u_cla32_and317_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and317_y0);
  and_gate and_gate_h_u_cla32_and318_y0(h_u_cla32_and317_y0, h_u_cla32_and316_y0, h_u_cla32_and318_y0);
  and_gate and_gate_h_u_cla32_and319_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and319_y0);
  and_gate and_gate_h_u_cla32_and320_y0(h_u_cla32_and319_y0, h_u_cla32_and318_y0, h_u_cla32_and320_y0);
  and_gate and_gate_h_u_cla32_and321_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and321_y0);
  and_gate and_gate_h_u_cla32_and322_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and322_y0);
  and_gate and_gate_h_u_cla32_and323_y0(h_u_cla32_and322_y0, h_u_cla32_and321_y0, h_u_cla32_and323_y0);
  and_gate and_gate_h_u_cla32_and324_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and324_y0);
  and_gate and_gate_h_u_cla32_and325_y0(h_u_cla32_and324_y0, h_u_cla32_and323_y0, h_u_cla32_and325_y0);
  and_gate and_gate_h_u_cla32_and326_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and326_y0);
  and_gate and_gate_h_u_cla32_and327_y0(h_u_cla32_and326_y0, h_u_cla32_and325_y0, h_u_cla32_and327_y0);
  and_gate and_gate_h_u_cla32_and328_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and328_y0);
  and_gate and_gate_h_u_cla32_and329_y0(h_u_cla32_and328_y0, h_u_cla32_and327_y0, h_u_cla32_and329_y0);
  and_gate and_gate_h_u_cla32_and330_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and330_y0);
  and_gate and_gate_h_u_cla32_and331_y0(h_u_cla32_and330_y0, h_u_cla32_and329_y0, h_u_cla32_and331_y0);
  and_gate and_gate_h_u_cla32_and332_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and332_y0);
  and_gate and_gate_h_u_cla32_and333_y0(h_u_cla32_and332_y0, h_u_cla32_and331_y0, h_u_cla32_and333_y0);
  and_gate and_gate_h_u_cla32_and334_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and334_y0);
  and_gate and_gate_h_u_cla32_and335_y0(h_u_cla32_and334_y0, h_u_cla32_and333_y0, h_u_cla32_and335_y0);
  and_gate and_gate_h_u_cla32_and336_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and336_y0);
  and_gate and_gate_h_u_cla32_and337_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and337_y0);
  and_gate and_gate_h_u_cla32_and338_y0(h_u_cla32_and337_y0, h_u_cla32_and336_y0, h_u_cla32_and338_y0);
  and_gate and_gate_h_u_cla32_and339_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and339_y0);
  and_gate and_gate_h_u_cla32_and340_y0(h_u_cla32_and339_y0, h_u_cla32_and338_y0, h_u_cla32_and340_y0);
  and_gate and_gate_h_u_cla32_and341_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and341_y0);
  and_gate and_gate_h_u_cla32_and342_y0(h_u_cla32_and341_y0, h_u_cla32_and340_y0, h_u_cla32_and342_y0);
  and_gate and_gate_h_u_cla32_and343_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and343_y0);
  and_gate and_gate_h_u_cla32_and344_y0(h_u_cla32_and343_y0, h_u_cla32_and342_y0, h_u_cla32_and344_y0);
  and_gate and_gate_h_u_cla32_and345_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and345_y0);
  and_gate and_gate_h_u_cla32_and346_y0(h_u_cla32_and345_y0, h_u_cla32_and344_y0, h_u_cla32_and346_y0);
  and_gate and_gate_h_u_cla32_and347_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and347_y0);
  and_gate and_gate_h_u_cla32_and348_y0(h_u_cla32_and347_y0, h_u_cla32_and346_y0, h_u_cla32_and348_y0);
  and_gate and_gate_h_u_cla32_and349_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and349_y0);
  and_gate and_gate_h_u_cla32_and350_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and350_y0);
  and_gate and_gate_h_u_cla32_and351_y0(h_u_cla32_and350_y0, h_u_cla32_and349_y0, h_u_cla32_and351_y0);
  and_gate and_gate_h_u_cla32_and352_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and352_y0);
  and_gate and_gate_h_u_cla32_and353_y0(h_u_cla32_and352_y0, h_u_cla32_and351_y0, h_u_cla32_and353_y0);
  and_gate and_gate_h_u_cla32_and354_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and354_y0);
  and_gate and_gate_h_u_cla32_and355_y0(h_u_cla32_and354_y0, h_u_cla32_and353_y0, h_u_cla32_and355_y0);
  and_gate and_gate_h_u_cla32_and356_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and356_y0);
  and_gate and_gate_h_u_cla32_and357_y0(h_u_cla32_and356_y0, h_u_cla32_and355_y0, h_u_cla32_and357_y0);
  and_gate and_gate_h_u_cla32_and358_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and358_y0);
  and_gate and_gate_h_u_cla32_and359_y0(h_u_cla32_and358_y0, h_u_cla32_and357_y0, h_u_cla32_and359_y0);
  and_gate and_gate_h_u_cla32_and360_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and360_y0);
  and_gate and_gate_h_u_cla32_and361_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and361_y0);
  and_gate and_gate_h_u_cla32_and362_y0(h_u_cla32_and361_y0, h_u_cla32_and360_y0, h_u_cla32_and362_y0);
  and_gate and_gate_h_u_cla32_and363_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and363_y0);
  and_gate and_gate_h_u_cla32_and364_y0(h_u_cla32_and363_y0, h_u_cla32_and362_y0, h_u_cla32_and364_y0);
  and_gate and_gate_h_u_cla32_and365_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and365_y0);
  and_gate and_gate_h_u_cla32_and366_y0(h_u_cla32_and365_y0, h_u_cla32_and364_y0, h_u_cla32_and366_y0);
  and_gate and_gate_h_u_cla32_and367_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and367_y0);
  and_gate and_gate_h_u_cla32_and368_y0(h_u_cla32_and367_y0, h_u_cla32_and366_y0, h_u_cla32_and368_y0);
  and_gate and_gate_h_u_cla32_and369_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and369_y0);
  and_gate and_gate_h_u_cla32_and370_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and370_y0);
  and_gate and_gate_h_u_cla32_and371_y0(h_u_cla32_and370_y0, h_u_cla32_and369_y0, h_u_cla32_and371_y0);
  and_gate and_gate_h_u_cla32_and372_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and372_y0);
  and_gate and_gate_h_u_cla32_and373_y0(h_u_cla32_and372_y0, h_u_cla32_and371_y0, h_u_cla32_and373_y0);
  and_gate and_gate_h_u_cla32_and374_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and374_y0);
  and_gate and_gate_h_u_cla32_and375_y0(h_u_cla32_and374_y0, h_u_cla32_and373_y0, h_u_cla32_and375_y0);
  and_gate and_gate_h_u_cla32_and376_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and376_y0);
  and_gate and_gate_h_u_cla32_and377_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and377_y0);
  and_gate and_gate_h_u_cla32_and378_y0(h_u_cla32_and377_y0, h_u_cla32_and376_y0, h_u_cla32_and378_y0);
  and_gate and_gate_h_u_cla32_and379_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and379_y0);
  and_gate and_gate_h_u_cla32_and380_y0(h_u_cla32_and379_y0, h_u_cla32_and378_y0, h_u_cla32_and380_y0);
  and_gate and_gate_h_u_cla32_and381_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and381_y0);
  and_gate and_gate_h_u_cla32_and382_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and382_y0);
  and_gate and_gate_h_u_cla32_and383_y0(h_u_cla32_and382_y0, h_u_cla32_and381_y0, h_u_cla32_and383_y0);
  and_gate and_gate_h_u_cla32_and384_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and384_y0);
  or_gate or_gate_h_u_cla32_or45_y0(h_u_cla32_and384_y0, h_u_cla32_and303_y0, h_u_cla32_or45_y0);
  or_gate or_gate_h_u_cla32_or46_y0(h_u_cla32_or45_y0, h_u_cla32_and320_y0, h_u_cla32_or46_y0);
  or_gate or_gate_h_u_cla32_or47_y0(h_u_cla32_or46_y0, h_u_cla32_and335_y0, h_u_cla32_or47_y0);
  or_gate or_gate_h_u_cla32_or48_y0(h_u_cla32_or47_y0, h_u_cla32_and348_y0, h_u_cla32_or48_y0);
  or_gate or_gate_h_u_cla32_or49_y0(h_u_cla32_or48_y0, h_u_cla32_and359_y0, h_u_cla32_or49_y0);
  or_gate or_gate_h_u_cla32_or50_y0(h_u_cla32_or49_y0, h_u_cla32_and368_y0, h_u_cla32_or50_y0);
  or_gate or_gate_h_u_cla32_or51_y0(h_u_cla32_or50_y0, h_u_cla32_and375_y0, h_u_cla32_or51_y0);
  or_gate or_gate_h_u_cla32_or52_y0(h_u_cla32_or51_y0, h_u_cla32_and380_y0, h_u_cla32_or52_y0);
  or_gate or_gate_h_u_cla32_or53_y0(h_u_cla32_or52_y0, h_u_cla32_and383_y0, h_u_cla32_or53_y0);
  or_gate or_gate_h_u_cla32_or54_y0(h_u_cla32_pg_logic9_y1, h_u_cla32_or53_y0, h_u_cla32_or54_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic10_y0(a_10, b_10, h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_pg_logic10_y2);
  xor_gate xor_gate_h_u_cla32_xor10_y0(h_u_cla32_pg_logic10_y2, h_u_cla32_or54_y0, h_u_cla32_xor10_y0);
  and_gate and_gate_h_u_cla32_and385_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and385_y0);
  and_gate and_gate_h_u_cla32_and386_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and386_y0);
  and_gate and_gate_h_u_cla32_and387_y0(h_u_cla32_and386_y0, h_u_cla32_and385_y0, h_u_cla32_and387_y0);
  and_gate and_gate_h_u_cla32_and388_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and388_y0);
  and_gate and_gate_h_u_cla32_and389_y0(h_u_cla32_and388_y0, h_u_cla32_and387_y0, h_u_cla32_and389_y0);
  and_gate and_gate_h_u_cla32_and390_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and390_y0);
  and_gate and_gate_h_u_cla32_and391_y0(h_u_cla32_and390_y0, h_u_cla32_and389_y0, h_u_cla32_and391_y0);
  and_gate and_gate_h_u_cla32_and392_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and392_y0);
  and_gate and_gate_h_u_cla32_and393_y0(h_u_cla32_and392_y0, h_u_cla32_and391_y0, h_u_cla32_and393_y0);
  and_gate and_gate_h_u_cla32_and394_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and394_y0);
  and_gate and_gate_h_u_cla32_and395_y0(h_u_cla32_and394_y0, h_u_cla32_and393_y0, h_u_cla32_and395_y0);
  and_gate and_gate_h_u_cla32_and396_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and396_y0);
  and_gate and_gate_h_u_cla32_and397_y0(h_u_cla32_and396_y0, h_u_cla32_and395_y0, h_u_cla32_and397_y0);
  and_gate and_gate_h_u_cla32_and398_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and398_y0);
  and_gate and_gate_h_u_cla32_and399_y0(h_u_cla32_and398_y0, h_u_cla32_and397_y0, h_u_cla32_and399_y0);
  and_gate and_gate_h_u_cla32_and400_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and400_y0);
  and_gate and_gate_h_u_cla32_and401_y0(h_u_cla32_and400_y0, h_u_cla32_and399_y0, h_u_cla32_and401_y0);
  and_gate and_gate_h_u_cla32_and402_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and402_y0);
  and_gate and_gate_h_u_cla32_and403_y0(h_u_cla32_and402_y0, h_u_cla32_and401_y0, h_u_cla32_and403_y0);
  and_gate and_gate_h_u_cla32_and404_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and404_y0);
  and_gate and_gate_h_u_cla32_and405_y0(h_u_cla32_and404_y0, h_u_cla32_and403_y0, h_u_cla32_and405_y0);
  and_gate and_gate_h_u_cla32_and406_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and406_y0);
  and_gate and_gate_h_u_cla32_and407_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and407_y0);
  and_gate and_gate_h_u_cla32_and408_y0(h_u_cla32_and407_y0, h_u_cla32_and406_y0, h_u_cla32_and408_y0);
  and_gate and_gate_h_u_cla32_and409_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and409_y0);
  and_gate and_gate_h_u_cla32_and410_y0(h_u_cla32_and409_y0, h_u_cla32_and408_y0, h_u_cla32_and410_y0);
  and_gate and_gate_h_u_cla32_and411_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and411_y0);
  and_gate and_gate_h_u_cla32_and412_y0(h_u_cla32_and411_y0, h_u_cla32_and410_y0, h_u_cla32_and412_y0);
  and_gate and_gate_h_u_cla32_and413_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and413_y0);
  and_gate and_gate_h_u_cla32_and414_y0(h_u_cla32_and413_y0, h_u_cla32_and412_y0, h_u_cla32_and414_y0);
  and_gate and_gate_h_u_cla32_and415_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and415_y0);
  and_gate and_gate_h_u_cla32_and416_y0(h_u_cla32_and415_y0, h_u_cla32_and414_y0, h_u_cla32_and416_y0);
  and_gate and_gate_h_u_cla32_and417_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and417_y0);
  and_gate and_gate_h_u_cla32_and418_y0(h_u_cla32_and417_y0, h_u_cla32_and416_y0, h_u_cla32_and418_y0);
  and_gate and_gate_h_u_cla32_and419_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and419_y0);
  and_gate and_gate_h_u_cla32_and420_y0(h_u_cla32_and419_y0, h_u_cla32_and418_y0, h_u_cla32_and420_y0);
  and_gate and_gate_h_u_cla32_and421_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and421_y0);
  and_gate and_gate_h_u_cla32_and422_y0(h_u_cla32_and421_y0, h_u_cla32_and420_y0, h_u_cla32_and422_y0);
  and_gate and_gate_h_u_cla32_and423_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and423_y0);
  and_gate and_gate_h_u_cla32_and424_y0(h_u_cla32_and423_y0, h_u_cla32_and422_y0, h_u_cla32_and424_y0);
  and_gate and_gate_h_u_cla32_and425_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and425_y0);
  and_gate and_gate_h_u_cla32_and426_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and426_y0);
  and_gate and_gate_h_u_cla32_and427_y0(h_u_cla32_and426_y0, h_u_cla32_and425_y0, h_u_cla32_and427_y0);
  and_gate and_gate_h_u_cla32_and428_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and428_y0);
  and_gate and_gate_h_u_cla32_and429_y0(h_u_cla32_and428_y0, h_u_cla32_and427_y0, h_u_cla32_and429_y0);
  and_gate and_gate_h_u_cla32_and430_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and430_y0);
  and_gate and_gate_h_u_cla32_and431_y0(h_u_cla32_and430_y0, h_u_cla32_and429_y0, h_u_cla32_and431_y0);
  and_gate and_gate_h_u_cla32_and432_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and432_y0);
  and_gate and_gate_h_u_cla32_and433_y0(h_u_cla32_and432_y0, h_u_cla32_and431_y0, h_u_cla32_and433_y0);
  and_gate and_gate_h_u_cla32_and434_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and434_y0);
  and_gate and_gate_h_u_cla32_and435_y0(h_u_cla32_and434_y0, h_u_cla32_and433_y0, h_u_cla32_and435_y0);
  and_gate and_gate_h_u_cla32_and436_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and436_y0);
  and_gate and_gate_h_u_cla32_and437_y0(h_u_cla32_and436_y0, h_u_cla32_and435_y0, h_u_cla32_and437_y0);
  and_gate and_gate_h_u_cla32_and438_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and438_y0);
  and_gate and_gate_h_u_cla32_and439_y0(h_u_cla32_and438_y0, h_u_cla32_and437_y0, h_u_cla32_and439_y0);
  and_gate and_gate_h_u_cla32_and440_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and440_y0);
  and_gate and_gate_h_u_cla32_and441_y0(h_u_cla32_and440_y0, h_u_cla32_and439_y0, h_u_cla32_and441_y0);
  and_gate and_gate_h_u_cla32_and442_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and442_y0);
  and_gate and_gate_h_u_cla32_and443_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and443_y0);
  and_gate and_gate_h_u_cla32_and444_y0(h_u_cla32_and443_y0, h_u_cla32_and442_y0, h_u_cla32_and444_y0);
  and_gate and_gate_h_u_cla32_and445_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and445_y0);
  and_gate and_gate_h_u_cla32_and446_y0(h_u_cla32_and445_y0, h_u_cla32_and444_y0, h_u_cla32_and446_y0);
  and_gate and_gate_h_u_cla32_and447_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and447_y0);
  and_gate and_gate_h_u_cla32_and448_y0(h_u_cla32_and447_y0, h_u_cla32_and446_y0, h_u_cla32_and448_y0);
  and_gate and_gate_h_u_cla32_and449_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and449_y0);
  and_gate and_gate_h_u_cla32_and450_y0(h_u_cla32_and449_y0, h_u_cla32_and448_y0, h_u_cla32_and450_y0);
  and_gate and_gate_h_u_cla32_and451_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and451_y0);
  and_gate and_gate_h_u_cla32_and452_y0(h_u_cla32_and451_y0, h_u_cla32_and450_y0, h_u_cla32_and452_y0);
  and_gate and_gate_h_u_cla32_and453_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and453_y0);
  and_gate and_gate_h_u_cla32_and454_y0(h_u_cla32_and453_y0, h_u_cla32_and452_y0, h_u_cla32_and454_y0);
  and_gate and_gate_h_u_cla32_and455_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and455_y0);
  and_gate and_gate_h_u_cla32_and456_y0(h_u_cla32_and455_y0, h_u_cla32_and454_y0, h_u_cla32_and456_y0);
  and_gate and_gate_h_u_cla32_and457_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and457_y0);
  and_gate and_gate_h_u_cla32_and458_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and458_y0);
  and_gate and_gate_h_u_cla32_and459_y0(h_u_cla32_and458_y0, h_u_cla32_and457_y0, h_u_cla32_and459_y0);
  and_gate and_gate_h_u_cla32_and460_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and460_y0);
  and_gate and_gate_h_u_cla32_and461_y0(h_u_cla32_and460_y0, h_u_cla32_and459_y0, h_u_cla32_and461_y0);
  and_gate and_gate_h_u_cla32_and462_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and462_y0);
  and_gate and_gate_h_u_cla32_and463_y0(h_u_cla32_and462_y0, h_u_cla32_and461_y0, h_u_cla32_and463_y0);
  and_gate and_gate_h_u_cla32_and464_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and464_y0);
  and_gate and_gate_h_u_cla32_and465_y0(h_u_cla32_and464_y0, h_u_cla32_and463_y0, h_u_cla32_and465_y0);
  and_gate and_gate_h_u_cla32_and466_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and466_y0);
  and_gate and_gate_h_u_cla32_and467_y0(h_u_cla32_and466_y0, h_u_cla32_and465_y0, h_u_cla32_and467_y0);
  and_gate and_gate_h_u_cla32_and468_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and468_y0);
  and_gate and_gate_h_u_cla32_and469_y0(h_u_cla32_and468_y0, h_u_cla32_and467_y0, h_u_cla32_and469_y0);
  and_gate and_gate_h_u_cla32_and470_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and470_y0);
  and_gate and_gate_h_u_cla32_and471_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and471_y0);
  and_gate and_gate_h_u_cla32_and472_y0(h_u_cla32_and471_y0, h_u_cla32_and470_y0, h_u_cla32_and472_y0);
  and_gate and_gate_h_u_cla32_and473_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and473_y0);
  and_gate and_gate_h_u_cla32_and474_y0(h_u_cla32_and473_y0, h_u_cla32_and472_y0, h_u_cla32_and474_y0);
  and_gate and_gate_h_u_cla32_and475_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and475_y0);
  and_gate and_gate_h_u_cla32_and476_y0(h_u_cla32_and475_y0, h_u_cla32_and474_y0, h_u_cla32_and476_y0);
  and_gate and_gate_h_u_cla32_and477_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and477_y0);
  and_gate and_gate_h_u_cla32_and478_y0(h_u_cla32_and477_y0, h_u_cla32_and476_y0, h_u_cla32_and478_y0);
  and_gate and_gate_h_u_cla32_and479_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and479_y0);
  and_gate and_gate_h_u_cla32_and480_y0(h_u_cla32_and479_y0, h_u_cla32_and478_y0, h_u_cla32_and480_y0);
  and_gate and_gate_h_u_cla32_and481_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and481_y0);
  and_gate and_gate_h_u_cla32_and482_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and482_y0);
  and_gate and_gate_h_u_cla32_and483_y0(h_u_cla32_and482_y0, h_u_cla32_and481_y0, h_u_cla32_and483_y0);
  and_gate and_gate_h_u_cla32_and484_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and484_y0);
  and_gate and_gate_h_u_cla32_and485_y0(h_u_cla32_and484_y0, h_u_cla32_and483_y0, h_u_cla32_and485_y0);
  and_gate and_gate_h_u_cla32_and486_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and486_y0);
  and_gate and_gate_h_u_cla32_and487_y0(h_u_cla32_and486_y0, h_u_cla32_and485_y0, h_u_cla32_and487_y0);
  and_gate and_gate_h_u_cla32_and488_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and488_y0);
  and_gate and_gate_h_u_cla32_and489_y0(h_u_cla32_and488_y0, h_u_cla32_and487_y0, h_u_cla32_and489_y0);
  and_gate and_gate_h_u_cla32_and490_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and490_y0);
  and_gate and_gate_h_u_cla32_and491_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and491_y0);
  and_gate and_gate_h_u_cla32_and492_y0(h_u_cla32_and491_y0, h_u_cla32_and490_y0, h_u_cla32_and492_y0);
  and_gate and_gate_h_u_cla32_and493_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and493_y0);
  and_gate and_gate_h_u_cla32_and494_y0(h_u_cla32_and493_y0, h_u_cla32_and492_y0, h_u_cla32_and494_y0);
  and_gate and_gate_h_u_cla32_and495_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and495_y0);
  and_gate and_gate_h_u_cla32_and496_y0(h_u_cla32_and495_y0, h_u_cla32_and494_y0, h_u_cla32_and496_y0);
  and_gate and_gate_h_u_cla32_and497_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and497_y0);
  and_gate and_gate_h_u_cla32_and498_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and498_y0);
  and_gate and_gate_h_u_cla32_and499_y0(h_u_cla32_and498_y0, h_u_cla32_and497_y0, h_u_cla32_and499_y0);
  and_gate and_gate_h_u_cla32_and500_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and500_y0);
  and_gate and_gate_h_u_cla32_and501_y0(h_u_cla32_and500_y0, h_u_cla32_and499_y0, h_u_cla32_and501_y0);
  and_gate and_gate_h_u_cla32_and502_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and502_y0);
  and_gate and_gate_h_u_cla32_and503_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and503_y0);
  and_gate and_gate_h_u_cla32_and504_y0(h_u_cla32_and503_y0, h_u_cla32_and502_y0, h_u_cla32_and504_y0);
  and_gate and_gate_h_u_cla32_and505_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and505_y0);
  or_gate or_gate_h_u_cla32_or55_y0(h_u_cla32_and505_y0, h_u_cla32_and405_y0, h_u_cla32_or55_y0);
  or_gate or_gate_h_u_cla32_or56_y0(h_u_cla32_or55_y0, h_u_cla32_and424_y0, h_u_cla32_or56_y0);
  or_gate or_gate_h_u_cla32_or57_y0(h_u_cla32_or56_y0, h_u_cla32_and441_y0, h_u_cla32_or57_y0);
  or_gate or_gate_h_u_cla32_or58_y0(h_u_cla32_or57_y0, h_u_cla32_and456_y0, h_u_cla32_or58_y0);
  or_gate or_gate_h_u_cla32_or59_y0(h_u_cla32_or58_y0, h_u_cla32_and469_y0, h_u_cla32_or59_y0);
  or_gate or_gate_h_u_cla32_or60_y0(h_u_cla32_or59_y0, h_u_cla32_and480_y0, h_u_cla32_or60_y0);
  or_gate or_gate_h_u_cla32_or61_y0(h_u_cla32_or60_y0, h_u_cla32_and489_y0, h_u_cla32_or61_y0);
  or_gate or_gate_h_u_cla32_or62_y0(h_u_cla32_or61_y0, h_u_cla32_and496_y0, h_u_cla32_or62_y0);
  or_gate or_gate_h_u_cla32_or63_y0(h_u_cla32_or62_y0, h_u_cla32_and501_y0, h_u_cla32_or63_y0);
  or_gate or_gate_h_u_cla32_or64_y0(h_u_cla32_or63_y0, h_u_cla32_and504_y0, h_u_cla32_or64_y0);
  or_gate or_gate_h_u_cla32_or65_y0(h_u_cla32_pg_logic10_y1, h_u_cla32_or64_y0, h_u_cla32_or65_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic11_y0(a_11, b_11, h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_pg_logic11_y2);
  xor_gate xor_gate_h_u_cla32_xor11_y0(h_u_cla32_pg_logic11_y2, h_u_cla32_or65_y0, h_u_cla32_xor11_y0);
  and_gate and_gate_h_u_cla32_and506_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and506_y0);
  and_gate and_gate_h_u_cla32_and507_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and507_y0);
  and_gate and_gate_h_u_cla32_and508_y0(h_u_cla32_and507_y0, h_u_cla32_and506_y0, h_u_cla32_and508_y0);
  and_gate and_gate_h_u_cla32_and509_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and509_y0);
  and_gate and_gate_h_u_cla32_and510_y0(h_u_cla32_and509_y0, h_u_cla32_and508_y0, h_u_cla32_and510_y0);
  and_gate and_gate_h_u_cla32_and511_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and511_y0);
  and_gate and_gate_h_u_cla32_and512_y0(h_u_cla32_and511_y0, h_u_cla32_and510_y0, h_u_cla32_and512_y0);
  and_gate and_gate_h_u_cla32_and513_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and513_y0);
  and_gate and_gate_h_u_cla32_and514_y0(h_u_cla32_and513_y0, h_u_cla32_and512_y0, h_u_cla32_and514_y0);
  and_gate and_gate_h_u_cla32_and515_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and515_y0);
  and_gate and_gate_h_u_cla32_and516_y0(h_u_cla32_and515_y0, h_u_cla32_and514_y0, h_u_cla32_and516_y0);
  and_gate and_gate_h_u_cla32_and517_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and517_y0);
  and_gate and_gate_h_u_cla32_and518_y0(h_u_cla32_and517_y0, h_u_cla32_and516_y0, h_u_cla32_and518_y0);
  and_gate and_gate_h_u_cla32_and519_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and519_y0);
  and_gate and_gate_h_u_cla32_and520_y0(h_u_cla32_and519_y0, h_u_cla32_and518_y0, h_u_cla32_and520_y0);
  and_gate and_gate_h_u_cla32_and521_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and521_y0);
  and_gate and_gate_h_u_cla32_and522_y0(h_u_cla32_and521_y0, h_u_cla32_and520_y0, h_u_cla32_and522_y0);
  and_gate and_gate_h_u_cla32_and523_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and523_y0);
  and_gate and_gate_h_u_cla32_and524_y0(h_u_cla32_and523_y0, h_u_cla32_and522_y0, h_u_cla32_and524_y0);
  and_gate and_gate_h_u_cla32_and525_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and525_y0);
  and_gate and_gate_h_u_cla32_and526_y0(h_u_cla32_and525_y0, h_u_cla32_and524_y0, h_u_cla32_and526_y0);
  and_gate and_gate_h_u_cla32_and527_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and527_y0);
  and_gate and_gate_h_u_cla32_and528_y0(h_u_cla32_and527_y0, h_u_cla32_and526_y0, h_u_cla32_and528_y0);
  and_gate and_gate_h_u_cla32_and529_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and529_y0);
  and_gate and_gate_h_u_cla32_and530_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and530_y0);
  and_gate and_gate_h_u_cla32_and531_y0(h_u_cla32_and530_y0, h_u_cla32_and529_y0, h_u_cla32_and531_y0);
  and_gate and_gate_h_u_cla32_and532_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and532_y0);
  and_gate and_gate_h_u_cla32_and533_y0(h_u_cla32_and532_y0, h_u_cla32_and531_y0, h_u_cla32_and533_y0);
  and_gate and_gate_h_u_cla32_and534_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and534_y0);
  and_gate and_gate_h_u_cla32_and535_y0(h_u_cla32_and534_y0, h_u_cla32_and533_y0, h_u_cla32_and535_y0);
  and_gate and_gate_h_u_cla32_and536_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and536_y0);
  and_gate and_gate_h_u_cla32_and537_y0(h_u_cla32_and536_y0, h_u_cla32_and535_y0, h_u_cla32_and537_y0);
  and_gate and_gate_h_u_cla32_and538_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and538_y0);
  and_gate and_gate_h_u_cla32_and539_y0(h_u_cla32_and538_y0, h_u_cla32_and537_y0, h_u_cla32_and539_y0);
  and_gate and_gate_h_u_cla32_and540_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and540_y0);
  and_gate and_gate_h_u_cla32_and541_y0(h_u_cla32_and540_y0, h_u_cla32_and539_y0, h_u_cla32_and541_y0);
  and_gate and_gate_h_u_cla32_and542_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and542_y0);
  and_gate and_gate_h_u_cla32_and543_y0(h_u_cla32_and542_y0, h_u_cla32_and541_y0, h_u_cla32_and543_y0);
  and_gate and_gate_h_u_cla32_and544_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and544_y0);
  and_gate and_gate_h_u_cla32_and545_y0(h_u_cla32_and544_y0, h_u_cla32_and543_y0, h_u_cla32_and545_y0);
  and_gate and_gate_h_u_cla32_and546_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and546_y0);
  and_gate and_gate_h_u_cla32_and547_y0(h_u_cla32_and546_y0, h_u_cla32_and545_y0, h_u_cla32_and547_y0);
  and_gate and_gate_h_u_cla32_and548_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and548_y0);
  and_gate and_gate_h_u_cla32_and549_y0(h_u_cla32_and548_y0, h_u_cla32_and547_y0, h_u_cla32_and549_y0);
  and_gate and_gate_h_u_cla32_and550_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and550_y0);
  and_gate and_gate_h_u_cla32_and551_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and551_y0);
  and_gate and_gate_h_u_cla32_and552_y0(h_u_cla32_and551_y0, h_u_cla32_and550_y0, h_u_cla32_and552_y0);
  and_gate and_gate_h_u_cla32_and553_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and553_y0);
  and_gate and_gate_h_u_cla32_and554_y0(h_u_cla32_and553_y0, h_u_cla32_and552_y0, h_u_cla32_and554_y0);
  and_gate and_gate_h_u_cla32_and555_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and555_y0);
  and_gate and_gate_h_u_cla32_and556_y0(h_u_cla32_and555_y0, h_u_cla32_and554_y0, h_u_cla32_and556_y0);
  and_gate and_gate_h_u_cla32_and557_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and557_y0);
  and_gate and_gate_h_u_cla32_and558_y0(h_u_cla32_and557_y0, h_u_cla32_and556_y0, h_u_cla32_and558_y0);
  and_gate and_gate_h_u_cla32_and559_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and559_y0);
  and_gate and_gate_h_u_cla32_and560_y0(h_u_cla32_and559_y0, h_u_cla32_and558_y0, h_u_cla32_and560_y0);
  and_gate and_gate_h_u_cla32_and561_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and561_y0);
  and_gate and_gate_h_u_cla32_and562_y0(h_u_cla32_and561_y0, h_u_cla32_and560_y0, h_u_cla32_and562_y0);
  and_gate and_gate_h_u_cla32_and563_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and563_y0);
  and_gate and_gate_h_u_cla32_and564_y0(h_u_cla32_and563_y0, h_u_cla32_and562_y0, h_u_cla32_and564_y0);
  and_gate and_gate_h_u_cla32_and565_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and565_y0);
  and_gate and_gate_h_u_cla32_and566_y0(h_u_cla32_and565_y0, h_u_cla32_and564_y0, h_u_cla32_and566_y0);
  and_gate and_gate_h_u_cla32_and567_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and567_y0);
  and_gate and_gate_h_u_cla32_and568_y0(h_u_cla32_and567_y0, h_u_cla32_and566_y0, h_u_cla32_and568_y0);
  and_gate and_gate_h_u_cla32_and569_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and569_y0);
  and_gate and_gate_h_u_cla32_and570_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and570_y0);
  and_gate and_gate_h_u_cla32_and571_y0(h_u_cla32_and570_y0, h_u_cla32_and569_y0, h_u_cla32_and571_y0);
  and_gate and_gate_h_u_cla32_and572_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and572_y0);
  and_gate and_gate_h_u_cla32_and573_y0(h_u_cla32_and572_y0, h_u_cla32_and571_y0, h_u_cla32_and573_y0);
  and_gate and_gate_h_u_cla32_and574_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and574_y0);
  and_gate and_gate_h_u_cla32_and575_y0(h_u_cla32_and574_y0, h_u_cla32_and573_y0, h_u_cla32_and575_y0);
  and_gate and_gate_h_u_cla32_and576_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and576_y0);
  and_gate and_gate_h_u_cla32_and577_y0(h_u_cla32_and576_y0, h_u_cla32_and575_y0, h_u_cla32_and577_y0);
  and_gate and_gate_h_u_cla32_and578_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and578_y0);
  and_gate and_gate_h_u_cla32_and579_y0(h_u_cla32_and578_y0, h_u_cla32_and577_y0, h_u_cla32_and579_y0);
  and_gate and_gate_h_u_cla32_and580_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and580_y0);
  and_gate and_gate_h_u_cla32_and581_y0(h_u_cla32_and580_y0, h_u_cla32_and579_y0, h_u_cla32_and581_y0);
  and_gate and_gate_h_u_cla32_and582_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and582_y0);
  and_gate and_gate_h_u_cla32_and583_y0(h_u_cla32_and582_y0, h_u_cla32_and581_y0, h_u_cla32_and583_y0);
  and_gate and_gate_h_u_cla32_and584_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and584_y0);
  and_gate and_gate_h_u_cla32_and585_y0(h_u_cla32_and584_y0, h_u_cla32_and583_y0, h_u_cla32_and585_y0);
  and_gate and_gate_h_u_cla32_and586_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and586_y0);
  and_gate and_gate_h_u_cla32_and587_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and587_y0);
  and_gate and_gate_h_u_cla32_and588_y0(h_u_cla32_and587_y0, h_u_cla32_and586_y0, h_u_cla32_and588_y0);
  and_gate and_gate_h_u_cla32_and589_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and589_y0);
  and_gate and_gate_h_u_cla32_and590_y0(h_u_cla32_and589_y0, h_u_cla32_and588_y0, h_u_cla32_and590_y0);
  and_gate and_gate_h_u_cla32_and591_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and591_y0);
  and_gate and_gate_h_u_cla32_and592_y0(h_u_cla32_and591_y0, h_u_cla32_and590_y0, h_u_cla32_and592_y0);
  and_gate and_gate_h_u_cla32_and593_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and593_y0);
  and_gate and_gate_h_u_cla32_and594_y0(h_u_cla32_and593_y0, h_u_cla32_and592_y0, h_u_cla32_and594_y0);
  and_gate and_gate_h_u_cla32_and595_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and595_y0);
  and_gate and_gate_h_u_cla32_and596_y0(h_u_cla32_and595_y0, h_u_cla32_and594_y0, h_u_cla32_and596_y0);
  and_gate and_gate_h_u_cla32_and597_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and597_y0);
  and_gate and_gate_h_u_cla32_and598_y0(h_u_cla32_and597_y0, h_u_cla32_and596_y0, h_u_cla32_and598_y0);
  and_gate and_gate_h_u_cla32_and599_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and599_y0);
  and_gate and_gate_h_u_cla32_and600_y0(h_u_cla32_and599_y0, h_u_cla32_and598_y0, h_u_cla32_and600_y0);
  and_gate and_gate_h_u_cla32_and601_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and601_y0);
  and_gate and_gate_h_u_cla32_and602_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and602_y0);
  and_gate and_gate_h_u_cla32_and603_y0(h_u_cla32_and602_y0, h_u_cla32_and601_y0, h_u_cla32_and603_y0);
  and_gate and_gate_h_u_cla32_and604_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and604_y0);
  and_gate and_gate_h_u_cla32_and605_y0(h_u_cla32_and604_y0, h_u_cla32_and603_y0, h_u_cla32_and605_y0);
  and_gate and_gate_h_u_cla32_and606_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and606_y0);
  and_gate and_gate_h_u_cla32_and607_y0(h_u_cla32_and606_y0, h_u_cla32_and605_y0, h_u_cla32_and607_y0);
  and_gate and_gate_h_u_cla32_and608_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and608_y0);
  and_gate and_gate_h_u_cla32_and609_y0(h_u_cla32_and608_y0, h_u_cla32_and607_y0, h_u_cla32_and609_y0);
  and_gate and_gate_h_u_cla32_and610_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and610_y0);
  and_gate and_gate_h_u_cla32_and611_y0(h_u_cla32_and610_y0, h_u_cla32_and609_y0, h_u_cla32_and611_y0);
  and_gate and_gate_h_u_cla32_and612_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and612_y0);
  and_gate and_gate_h_u_cla32_and613_y0(h_u_cla32_and612_y0, h_u_cla32_and611_y0, h_u_cla32_and613_y0);
  and_gate and_gate_h_u_cla32_and614_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and614_y0);
  and_gate and_gate_h_u_cla32_and615_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and615_y0);
  and_gate and_gate_h_u_cla32_and616_y0(h_u_cla32_and615_y0, h_u_cla32_and614_y0, h_u_cla32_and616_y0);
  and_gate and_gate_h_u_cla32_and617_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and617_y0);
  and_gate and_gate_h_u_cla32_and618_y0(h_u_cla32_and617_y0, h_u_cla32_and616_y0, h_u_cla32_and618_y0);
  and_gate and_gate_h_u_cla32_and619_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and619_y0);
  and_gate and_gate_h_u_cla32_and620_y0(h_u_cla32_and619_y0, h_u_cla32_and618_y0, h_u_cla32_and620_y0);
  and_gate and_gate_h_u_cla32_and621_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and621_y0);
  and_gate and_gate_h_u_cla32_and622_y0(h_u_cla32_and621_y0, h_u_cla32_and620_y0, h_u_cla32_and622_y0);
  and_gate and_gate_h_u_cla32_and623_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and623_y0);
  and_gate and_gate_h_u_cla32_and624_y0(h_u_cla32_and623_y0, h_u_cla32_and622_y0, h_u_cla32_and624_y0);
  and_gate and_gate_h_u_cla32_and625_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and625_y0);
  and_gate and_gate_h_u_cla32_and626_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and626_y0);
  and_gate and_gate_h_u_cla32_and627_y0(h_u_cla32_and626_y0, h_u_cla32_and625_y0, h_u_cla32_and627_y0);
  and_gate and_gate_h_u_cla32_and628_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and628_y0);
  and_gate and_gate_h_u_cla32_and629_y0(h_u_cla32_and628_y0, h_u_cla32_and627_y0, h_u_cla32_and629_y0);
  and_gate and_gate_h_u_cla32_and630_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and630_y0);
  and_gate and_gate_h_u_cla32_and631_y0(h_u_cla32_and630_y0, h_u_cla32_and629_y0, h_u_cla32_and631_y0);
  and_gate and_gate_h_u_cla32_and632_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and632_y0);
  and_gate and_gate_h_u_cla32_and633_y0(h_u_cla32_and632_y0, h_u_cla32_and631_y0, h_u_cla32_and633_y0);
  and_gate and_gate_h_u_cla32_and634_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and634_y0);
  and_gate and_gate_h_u_cla32_and635_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and635_y0);
  and_gate and_gate_h_u_cla32_and636_y0(h_u_cla32_and635_y0, h_u_cla32_and634_y0, h_u_cla32_and636_y0);
  and_gate and_gate_h_u_cla32_and637_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and637_y0);
  and_gate and_gate_h_u_cla32_and638_y0(h_u_cla32_and637_y0, h_u_cla32_and636_y0, h_u_cla32_and638_y0);
  and_gate and_gate_h_u_cla32_and639_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and639_y0);
  and_gate and_gate_h_u_cla32_and640_y0(h_u_cla32_and639_y0, h_u_cla32_and638_y0, h_u_cla32_and640_y0);
  and_gate and_gate_h_u_cla32_and641_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and641_y0);
  and_gate and_gate_h_u_cla32_and642_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and642_y0);
  and_gate and_gate_h_u_cla32_and643_y0(h_u_cla32_and642_y0, h_u_cla32_and641_y0, h_u_cla32_and643_y0);
  and_gate and_gate_h_u_cla32_and644_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and644_y0);
  and_gate and_gate_h_u_cla32_and645_y0(h_u_cla32_and644_y0, h_u_cla32_and643_y0, h_u_cla32_and645_y0);
  and_gate and_gate_h_u_cla32_and646_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and646_y0);
  and_gate and_gate_h_u_cla32_and647_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and647_y0);
  and_gate and_gate_h_u_cla32_and648_y0(h_u_cla32_and647_y0, h_u_cla32_and646_y0, h_u_cla32_and648_y0);
  and_gate and_gate_h_u_cla32_and649_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and649_y0);
  or_gate or_gate_h_u_cla32_or66_y0(h_u_cla32_and649_y0, h_u_cla32_and528_y0, h_u_cla32_or66_y0);
  or_gate or_gate_h_u_cla32_or67_y0(h_u_cla32_or66_y0, h_u_cla32_and549_y0, h_u_cla32_or67_y0);
  or_gate or_gate_h_u_cla32_or68_y0(h_u_cla32_or67_y0, h_u_cla32_and568_y0, h_u_cla32_or68_y0);
  or_gate or_gate_h_u_cla32_or69_y0(h_u_cla32_or68_y0, h_u_cla32_and585_y0, h_u_cla32_or69_y0);
  or_gate or_gate_h_u_cla32_or70_y0(h_u_cla32_or69_y0, h_u_cla32_and600_y0, h_u_cla32_or70_y0);
  or_gate or_gate_h_u_cla32_or71_y0(h_u_cla32_or70_y0, h_u_cla32_and613_y0, h_u_cla32_or71_y0);
  or_gate or_gate_h_u_cla32_or72_y0(h_u_cla32_or71_y0, h_u_cla32_and624_y0, h_u_cla32_or72_y0);
  or_gate or_gate_h_u_cla32_or73_y0(h_u_cla32_or72_y0, h_u_cla32_and633_y0, h_u_cla32_or73_y0);
  or_gate or_gate_h_u_cla32_or74_y0(h_u_cla32_or73_y0, h_u_cla32_and640_y0, h_u_cla32_or74_y0);
  or_gate or_gate_h_u_cla32_or75_y0(h_u_cla32_or74_y0, h_u_cla32_and645_y0, h_u_cla32_or75_y0);
  or_gate or_gate_h_u_cla32_or76_y0(h_u_cla32_or75_y0, h_u_cla32_and648_y0, h_u_cla32_or76_y0);
  or_gate or_gate_h_u_cla32_or77_y0(h_u_cla32_pg_logic11_y1, h_u_cla32_or76_y0, h_u_cla32_or77_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic12_y0(a_12, b_12, h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_pg_logic12_y2);
  xor_gate xor_gate_h_u_cla32_xor12_y0(h_u_cla32_pg_logic12_y2, h_u_cla32_or77_y0, h_u_cla32_xor12_y0);
  and_gate and_gate_h_u_cla32_and650_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and650_y0);
  and_gate and_gate_h_u_cla32_and651_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and651_y0);
  and_gate and_gate_h_u_cla32_and652_y0(h_u_cla32_and651_y0, h_u_cla32_and650_y0, h_u_cla32_and652_y0);
  and_gate and_gate_h_u_cla32_and653_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and653_y0);
  and_gate and_gate_h_u_cla32_and654_y0(h_u_cla32_and653_y0, h_u_cla32_and652_y0, h_u_cla32_and654_y0);
  and_gate and_gate_h_u_cla32_and655_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and655_y0);
  and_gate and_gate_h_u_cla32_and656_y0(h_u_cla32_and655_y0, h_u_cla32_and654_y0, h_u_cla32_and656_y0);
  and_gate and_gate_h_u_cla32_and657_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and657_y0);
  and_gate and_gate_h_u_cla32_and658_y0(h_u_cla32_and657_y0, h_u_cla32_and656_y0, h_u_cla32_and658_y0);
  and_gate and_gate_h_u_cla32_and659_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and659_y0);
  and_gate and_gate_h_u_cla32_and660_y0(h_u_cla32_and659_y0, h_u_cla32_and658_y0, h_u_cla32_and660_y0);
  and_gate and_gate_h_u_cla32_and661_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and661_y0);
  and_gate and_gate_h_u_cla32_and662_y0(h_u_cla32_and661_y0, h_u_cla32_and660_y0, h_u_cla32_and662_y0);
  and_gate and_gate_h_u_cla32_and663_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and663_y0);
  and_gate and_gate_h_u_cla32_and664_y0(h_u_cla32_and663_y0, h_u_cla32_and662_y0, h_u_cla32_and664_y0);
  and_gate and_gate_h_u_cla32_and665_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and665_y0);
  and_gate and_gate_h_u_cla32_and666_y0(h_u_cla32_and665_y0, h_u_cla32_and664_y0, h_u_cla32_and666_y0);
  and_gate and_gate_h_u_cla32_and667_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and667_y0);
  and_gate and_gate_h_u_cla32_and668_y0(h_u_cla32_and667_y0, h_u_cla32_and666_y0, h_u_cla32_and668_y0);
  and_gate and_gate_h_u_cla32_and669_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and669_y0);
  and_gate and_gate_h_u_cla32_and670_y0(h_u_cla32_and669_y0, h_u_cla32_and668_y0, h_u_cla32_and670_y0);
  and_gate and_gate_h_u_cla32_and671_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and671_y0);
  and_gate and_gate_h_u_cla32_and672_y0(h_u_cla32_and671_y0, h_u_cla32_and670_y0, h_u_cla32_and672_y0);
  and_gate and_gate_h_u_cla32_and673_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and673_y0);
  and_gate and_gate_h_u_cla32_and674_y0(h_u_cla32_and673_y0, h_u_cla32_and672_y0, h_u_cla32_and674_y0);
  and_gate and_gate_h_u_cla32_and675_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and675_y0);
  and_gate and_gate_h_u_cla32_and676_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and676_y0);
  and_gate and_gate_h_u_cla32_and677_y0(h_u_cla32_and676_y0, h_u_cla32_and675_y0, h_u_cla32_and677_y0);
  and_gate and_gate_h_u_cla32_and678_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and678_y0);
  and_gate and_gate_h_u_cla32_and679_y0(h_u_cla32_and678_y0, h_u_cla32_and677_y0, h_u_cla32_and679_y0);
  and_gate and_gate_h_u_cla32_and680_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and680_y0);
  and_gate and_gate_h_u_cla32_and681_y0(h_u_cla32_and680_y0, h_u_cla32_and679_y0, h_u_cla32_and681_y0);
  and_gate and_gate_h_u_cla32_and682_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and682_y0);
  and_gate and_gate_h_u_cla32_and683_y0(h_u_cla32_and682_y0, h_u_cla32_and681_y0, h_u_cla32_and683_y0);
  and_gate and_gate_h_u_cla32_and684_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and684_y0);
  and_gate and_gate_h_u_cla32_and685_y0(h_u_cla32_and684_y0, h_u_cla32_and683_y0, h_u_cla32_and685_y0);
  and_gate and_gate_h_u_cla32_and686_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and686_y0);
  and_gate and_gate_h_u_cla32_and687_y0(h_u_cla32_and686_y0, h_u_cla32_and685_y0, h_u_cla32_and687_y0);
  and_gate and_gate_h_u_cla32_and688_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and688_y0);
  and_gate and_gate_h_u_cla32_and689_y0(h_u_cla32_and688_y0, h_u_cla32_and687_y0, h_u_cla32_and689_y0);
  and_gate and_gate_h_u_cla32_and690_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and690_y0);
  and_gate and_gate_h_u_cla32_and691_y0(h_u_cla32_and690_y0, h_u_cla32_and689_y0, h_u_cla32_and691_y0);
  and_gate and_gate_h_u_cla32_and692_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and692_y0);
  and_gate and_gate_h_u_cla32_and693_y0(h_u_cla32_and692_y0, h_u_cla32_and691_y0, h_u_cla32_and693_y0);
  and_gate and_gate_h_u_cla32_and694_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and694_y0);
  and_gate and_gate_h_u_cla32_and695_y0(h_u_cla32_and694_y0, h_u_cla32_and693_y0, h_u_cla32_and695_y0);
  and_gate and_gate_h_u_cla32_and696_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and696_y0);
  and_gate and_gate_h_u_cla32_and697_y0(h_u_cla32_and696_y0, h_u_cla32_and695_y0, h_u_cla32_and697_y0);
  and_gate and_gate_h_u_cla32_and698_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and698_y0);
  and_gate and_gate_h_u_cla32_and699_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and699_y0);
  and_gate and_gate_h_u_cla32_and700_y0(h_u_cla32_and699_y0, h_u_cla32_and698_y0, h_u_cla32_and700_y0);
  and_gate and_gate_h_u_cla32_and701_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and701_y0);
  and_gate and_gate_h_u_cla32_and702_y0(h_u_cla32_and701_y0, h_u_cla32_and700_y0, h_u_cla32_and702_y0);
  and_gate and_gate_h_u_cla32_and703_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and703_y0);
  and_gate and_gate_h_u_cla32_and704_y0(h_u_cla32_and703_y0, h_u_cla32_and702_y0, h_u_cla32_and704_y0);
  and_gate and_gate_h_u_cla32_and705_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and705_y0);
  and_gate and_gate_h_u_cla32_and706_y0(h_u_cla32_and705_y0, h_u_cla32_and704_y0, h_u_cla32_and706_y0);
  and_gate and_gate_h_u_cla32_and707_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and707_y0);
  and_gate and_gate_h_u_cla32_and708_y0(h_u_cla32_and707_y0, h_u_cla32_and706_y0, h_u_cla32_and708_y0);
  and_gate and_gate_h_u_cla32_and709_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and709_y0);
  and_gate and_gate_h_u_cla32_and710_y0(h_u_cla32_and709_y0, h_u_cla32_and708_y0, h_u_cla32_and710_y0);
  and_gate and_gate_h_u_cla32_and711_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and711_y0);
  and_gate and_gate_h_u_cla32_and712_y0(h_u_cla32_and711_y0, h_u_cla32_and710_y0, h_u_cla32_and712_y0);
  and_gate and_gate_h_u_cla32_and713_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and713_y0);
  and_gate and_gate_h_u_cla32_and714_y0(h_u_cla32_and713_y0, h_u_cla32_and712_y0, h_u_cla32_and714_y0);
  and_gate and_gate_h_u_cla32_and715_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and715_y0);
  and_gate and_gate_h_u_cla32_and716_y0(h_u_cla32_and715_y0, h_u_cla32_and714_y0, h_u_cla32_and716_y0);
  and_gate and_gate_h_u_cla32_and717_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and717_y0);
  and_gate and_gate_h_u_cla32_and718_y0(h_u_cla32_and717_y0, h_u_cla32_and716_y0, h_u_cla32_and718_y0);
  and_gate and_gate_h_u_cla32_and719_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and719_y0);
  and_gate and_gate_h_u_cla32_and720_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and720_y0);
  and_gate and_gate_h_u_cla32_and721_y0(h_u_cla32_and720_y0, h_u_cla32_and719_y0, h_u_cla32_and721_y0);
  and_gate and_gate_h_u_cla32_and722_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and722_y0);
  and_gate and_gate_h_u_cla32_and723_y0(h_u_cla32_and722_y0, h_u_cla32_and721_y0, h_u_cla32_and723_y0);
  and_gate and_gate_h_u_cla32_and724_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and724_y0);
  and_gate and_gate_h_u_cla32_and725_y0(h_u_cla32_and724_y0, h_u_cla32_and723_y0, h_u_cla32_and725_y0);
  and_gate and_gate_h_u_cla32_and726_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and726_y0);
  and_gate and_gate_h_u_cla32_and727_y0(h_u_cla32_and726_y0, h_u_cla32_and725_y0, h_u_cla32_and727_y0);
  and_gate and_gate_h_u_cla32_and728_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and728_y0);
  and_gate and_gate_h_u_cla32_and729_y0(h_u_cla32_and728_y0, h_u_cla32_and727_y0, h_u_cla32_and729_y0);
  and_gate and_gate_h_u_cla32_and730_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and730_y0);
  and_gate and_gate_h_u_cla32_and731_y0(h_u_cla32_and730_y0, h_u_cla32_and729_y0, h_u_cla32_and731_y0);
  and_gate and_gate_h_u_cla32_and732_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and732_y0);
  and_gate and_gate_h_u_cla32_and733_y0(h_u_cla32_and732_y0, h_u_cla32_and731_y0, h_u_cla32_and733_y0);
  and_gate and_gate_h_u_cla32_and734_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and734_y0);
  and_gate and_gate_h_u_cla32_and735_y0(h_u_cla32_and734_y0, h_u_cla32_and733_y0, h_u_cla32_and735_y0);
  and_gate and_gate_h_u_cla32_and736_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and736_y0);
  and_gate and_gate_h_u_cla32_and737_y0(h_u_cla32_and736_y0, h_u_cla32_and735_y0, h_u_cla32_and737_y0);
  and_gate and_gate_h_u_cla32_and738_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and738_y0);
  and_gate and_gate_h_u_cla32_and739_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and739_y0);
  and_gate and_gate_h_u_cla32_and740_y0(h_u_cla32_and739_y0, h_u_cla32_and738_y0, h_u_cla32_and740_y0);
  and_gate and_gate_h_u_cla32_and741_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and741_y0);
  and_gate and_gate_h_u_cla32_and742_y0(h_u_cla32_and741_y0, h_u_cla32_and740_y0, h_u_cla32_and742_y0);
  and_gate and_gate_h_u_cla32_and743_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and743_y0);
  and_gate and_gate_h_u_cla32_and744_y0(h_u_cla32_and743_y0, h_u_cla32_and742_y0, h_u_cla32_and744_y0);
  and_gate and_gate_h_u_cla32_and745_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and745_y0);
  and_gate and_gate_h_u_cla32_and746_y0(h_u_cla32_and745_y0, h_u_cla32_and744_y0, h_u_cla32_and746_y0);
  and_gate and_gate_h_u_cla32_and747_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and747_y0);
  and_gate and_gate_h_u_cla32_and748_y0(h_u_cla32_and747_y0, h_u_cla32_and746_y0, h_u_cla32_and748_y0);
  and_gate and_gate_h_u_cla32_and749_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and749_y0);
  and_gate and_gate_h_u_cla32_and750_y0(h_u_cla32_and749_y0, h_u_cla32_and748_y0, h_u_cla32_and750_y0);
  and_gate and_gate_h_u_cla32_and751_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and751_y0);
  and_gate and_gate_h_u_cla32_and752_y0(h_u_cla32_and751_y0, h_u_cla32_and750_y0, h_u_cla32_and752_y0);
  and_gate and_gate_h_u_cla32_and753_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and753_y0);
  and_gate and_gate_h_u_cla32_and754_y0(h_u_cla32_and753_y0, h_u_cla32_and752_y0, h_u_cla32_and754_y0);
  and_gate and_gate_h_u_cla32_and755_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and755_y0);
  and_gate and_gate_h_u_cla32_and756_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and756_y0);
  and_gate and_gate_h_u_cla32_and757_y0(h_u_cla32_and756_y0, h_u_cla32_and755_y0, h_u_cla32_and757_y0);
  and_gate and_gate_h_u_cla32_and758_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and758_y0);
  and_gate and_gate_h_u_cla32_and759_y0(h_u_cla32_and758_y0, h_u_cla32_and757_y0, h_u_cla32_and759_y0);
  and_gate and_gate_h_u_cla32_and760_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and760_y0);
  and_gate and_gate_h_u_cla32_and761_y0(h_u_cla32_and760_y0, h_u_cla32_and759_y0, h_u_cla32_and761_y0);
  and_gate and_gate_h_u_cla32_and762_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and762_y0);
  and_gate and_gate_h_u_cla32_and763_y0(h_u_cla32_and762_y0, h_u_cla32_and761_y0, h_u_cla32_and763_y0);
  and_gate and_gate_h_u_cla32_and764_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and764_y0);
  and_gate and_gate_h_u_cla32_and765_y0(h_u_cla32_and764_y0, h_u_cla32_and763_y0, h_u_cla32_and765_y0);
  and_gate and_gate_h_u_cla32_and766_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and766_y0);
  and_gate and_gate_h_u_cla32_and767_y0(h_u_cla32_and766_y0, h_u_cla32_and765_y0, h_u_cla32_and767_y0);
  and_gate and_gate_h_u_cla32_and768_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and768_y0);
  and_gate and_gate_h_u_cla32_and769_y0(h_u_cla32_and768_y0, h_u_cla32_and767_y0, h_u_cla32_and769_y0);
  and_gate and_gate_h_u_cla32_and770_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and770_y0);
  and_gate and_gate_h_u_cla32_and771_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and771_y0);
  and_gate and_gate_h_u_cla32_and772_y0(h_u_cla32_and771_y0, h_u_cla32_and770_y0, h_u_cla32_and772_y0);
  and_gate and_gate_h_u_cla32_and773_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and773_y0);
  and_gate and_gate_h_u_cla32_and774_y0(h_u_cla32_and773_y0, h_u_cla32_and772_y0, h_u_cla32_and774_y0);
  and_gate and_gate_h_u_cla32_and775_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and775_y0);
  and_gate and_gate_h_u_cla32_and776_y0(h_u_cla32_and775_y0, h_u_cla32_and774_y0, h_u_cla32_and776_y0);
  and_gate and_gate_h_u_cla32_and777_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and777_y0);
  and_gate and_gate_h_u_cla32_and778_y0(h_u_cla32_and777_y0, h_u_cla32_and776_y0, h_u_cla32_and778_y0);
  and_gate and_gate_h_u_cla32_and779_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and779_y0);
  and_gate and_gate_h_u_cla32_and780_y0(h_u_cla32_and779_y0, h_u_cla32_and778_y0, h_u_cla32_and780_y0);
  and_gate and_gate_h_u_cla32_and781_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and781_y0);
  and_gate and_gate_h_u_cla32_and782_y0(h_u_cla32_and781_y0, h_u_cla32_and780_y0, h_u_cla32_and782_y0);
  and_gate and_gate_h_u_cla32_and783_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and783_y0);
  and_gate and_gate_h_u_cla32_and784_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and784_y0);
  and_gate and_gate_h_u_cla32_and785_y0(h_u_cla32_and784_y0, h_u_cla32_and783_y0, h_u_cla32_and785_y0);
  and_gate and_gate_h_u_cla32_and786_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and786_y0);
  and_gate and_gate_h_u_cla32_and787_y0(h_u_cla32_and786_y0, h_u_cla32_and785_y0, h_u_cla32_and787_y0);
  and_gate and_gate_h_u_cla32_and788_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and788_y0);
  and_gate and_gate_h_u_cla32_and789_y0(h_u_cla32_and788_y0, h_u_cla32_and787_y0, h_u_cla32_and789_y0);
  and_gate and_gate_h_u_cla32_and790_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and790_y0);
  and_gate and_gate_h_u_cla32_and791_y0(h_u_cla32_and790_y0, h_u_cla32_and789_y0, h_u_cla32_and791_y0);
  and_gate and_gate_h_u_cla32_and792_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and792_y0);
  and_gate and_gate_h_u_cla32_and793_y0(h_u_cla32_and792_y0, h_u_cla32_and791_y0, h_u_cla32_and793_y0);
  and_gate and_gate_h_u_cla32_and794_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and794_y0);
  and_gate and_gate_h_u_cla32_and795_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and795_y0);
  and_gate and_gate_h_u_cla32_and796_y0(h_u_cla32_and795_y0, h_u_cla32_and794_y0, h_u_cla32_and796_y0);
  and_gate and_gate_h_u_cla32_and797_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and797_y0);
  and_gate and_gate_h_u_cla32_and798_y0(h_u_cla32_and797_y0, h_u_cla32_and796_y0, h_u_cla32_and798_y0);
  and_gate and_gate_h_u_cla32_and799_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and799_y0);
  and_gate and_gate_h_u_cla32_and800_y0(h_u_cla32_and799_y0, h_u_cla32_and798_y0, h_u_cla32_and800_y0);
  and_gate and_gate_h_u_cla32_and801_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and801_y0);
  and_gate and_gate_h_u_cla32_and802_y0(h_u_cla32_and801_y0, h_u_cla32_and800_y0, h_u_cla32_and802_y0);
  and_gate and_gate_h_u_cla32_and803_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and803_y0);
  and_gate and_gate_h_u_cla32_and804_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and804_y0);
  and_gate and_gate_h_u_cla32_and805_y0(h_u_cla32_and804_y0, h_u_cla32_and803_y0, h_u_cla32_and805_y0);
  and_gate and_gate_h_u_cla32_and806_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and806_y0);
  and_gate and_gate_h_u_cla32_and807_y0(h_u_cla32_and806_y0, h_u_cla32_and805_y0, h_u_cla32_and807_y0);
  and_gate and_gate_h_u_cla32_and808_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and808_y0);
  and_gate and_gate_h_u_cla32_and809_y0(h_u_cla32_and808_y0, h_u_cla32_and807_y0, h_u_cla32_and809_y0);
  and_gate and_gate_h_u_cla32_and810_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and810_y0);
  and_gate and_gate_h_u_cla32_and811_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and811_y0);
  and_gate and_gate_h_u_cla32_and812_y0(h_u_cla32_and811_y0, h_u_cla32_and810_y0, h_u_cla32_and812_y0);
  and_gate and_gate_h_u_cla32_and813_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and813_y0);
  and_gate and_gate_h_u_cla32_and814_y0(h_u_cla32_and813_y0, h_u_cla32_and812_y0, h_u_cla32_and814_y0);
  and_gate and_gate_h_u_cla32_and815_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and815_y0);
  and_gate and_gate_h_u_cla32_and816_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and816_y0);
  and_gate and_gate_h_u_cla32_and817_y0(h_u_cla32_and816_y0, h_u_cla32_and815_y0, h_u_cla32_and817_y0);
  and_gate and_gate_h_u_cla32_and818_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and818_y0);
  or_gate or_gate_h_u_cla32_or78_y0(h_u_cla32_and818_y0, h_u_cla32_and674_y0, h_u_cla32_or78_y0);
  or_gate or_gate_h_u_cla32_or79_y0(h_u_cla32_or78_y0, h_u_cla32_and697_y0, h_u_cla32_or79_y0);
  or_gate or_gate_h_u_cla32_or80_y0(h_u_cla32_or79_y0, h_u_cla32_and718_y0, h_u_cla32_or80_y0);
  or_gate or_gate_h_u_cla32_or81_y0(h_u_cla32_or80_y0, h_u_cla32_and737_y0, h_u_cla32_or81_y0);
  or_gate or_gate_h_u_cla32_or82_y0(h_u_cla32_or81_y0, h_u_cla32_and754_y0, h_u_cla32_or82_y0);
  or_gate or_gate_h_u_cla32_or83_y0(h_u_cla32_or82_y0, h_u_cla32_and769_y0, h_u_cla32_or83_y0);
  or_gate or_gate_h_u_cla32_or84_y0(h_u_cla32_or83_y0, h_u_cla32_and782_y0, h_u_cla32_or84_y0);
  or_gate or_gate_h_u_cla32_or85_y0(h_u_cla32_or84_y0, h_u_cla32_and793_y0, h_u_cla32_or85_y0);
  or_gate or_gate_h_u_cla32_or86_y0(h_u_cla32_or85_y0, h_u_cla32_and802_y0, h_u_cla32_or86_y0);
  or_gate or_gate_h_u_cla32_or87_y0(h_u_cla32_or86_y0, h_u_cla32_and809_y0, h_u_cla32_or87_y0);
  or_gate or_gate_h_u_cla32_or88_y0(h_u_cla32_or87_y0, h_u_cla32_and814_y0, h_u_cla32_or88_y0);
  or_gate or_gate_h_u_cla32_or89_y0(h_u_cla32_or88_y0, h_u_cla32_and817_y0, h_u_cla32_or89_y0);
  or_gate or_gate_h_u_cla32_or90_y0(h_u_cla32_pg_logic12_y1, h_u_cla32_or89_y0, h_u_cla32_or90_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic13_y0(a_13, b_13, h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_pg_logic13_y2);
  xor_gate xor_gate_h_u_cla32_xor13_y0(h_u_cla32_pg_logic13_y2, h_u_cla32_or90_y0, h_u_cla32_xor13_y0);
  and_gate and_gate_h_u_cla32_and819_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and819_y0);
  and_gate and_gate_h_u_cla32_and820_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and820_y0);
  and_gate and_gate_h_u_cla32_and821_y0(h_u_cla32_and820_y0, h_u_cla32_and819_y0, h_u_cla32_and821_y0);
  and_gate and_gate_h_u_cla32_and822_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and822_y0);
  and_gate and_gate_h_u_cla32_and823_y0(h_u_cla32_and822_y0, h_u_cla32_and821_y0, h_u_cla32_and823_y0);
  and_gate and_gate_h_u_cla32_and824_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and824_y0);
  and_gate and_gate_h_u_cla32_and825_y0(h_u_cla32_and824_y0, h_u_cla32_and823_y0, h_u_cla32_and825_y0);
  and_gate and_gate_h_u_cla32_and826_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and826_y0);
  and_gate and_gate_h_u_cla32_and827_y0(h_u_cla32_and826_y0, h_u_cla32_and825_y0, h_u_cla32_and827_y0);
  and_gate and_gate_h_u_cla32_and828_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and828_y0);
  and_gate and_gate_h_u_cla32_and829_y0(h_u_cla32_and828_y0, h_u_cla32_and827_y0, h_u_cla32_and829_y0);
  and_gate and_gate_h_u_cla32_and830_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and830_y0);
  and_gate and_gate_h_u_cla32_and831_y0(h_u_cla32_and830_y0, h_u_cla32_and829_y0, h_u_cla32_and831_y0);
  and_gate and_gate_h_u_cla32_and832_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and832_y0);
  and_gate and_gate_h_u_cla32_and833_y0(h_u_cla32_and832_y0, h_u_cla32_and831_y0, h_u_cla32_and833_y0);
  and_gate and_gate_h_u_cla32_and834_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and834_y0);
  and_gate and_gate_h_u_cla32_and835_y0(h_u_cla32_and834_y0, h_u_cla32_and833_y0, h_u_cla32_and835_y0);
  and_gate and_gate_h_u_cla32_and836_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and836_y0);
  and_gate and_gate_h_u_cla32_and837_y0(h_u_cla32_and836_y0, h_u_cla32_and835_y0, h_u_cla32_and837_y0);
  and_gate and_gate_h_u_cla32_and838_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and838_y0);
  and_gate and_gate_h_u_cla32_and839_y0(h_u_cla32_and838_y0, h_u_cla32_and837_y0, h_u_cla32_and839_y0);
  and_gate and_gate_h_u_cla32_and840_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and840_y0);
  and_gate and_gate_h_u_cla32_and841_y0(h_u_cla32_and840_y0, h_u_cla32_and839_y0, h_u_cla32_and841_y0);
  and_gate and_gate_h_u_cla32_and842_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and842_y0);
  and_gate and_gate_h_u_cla32_and843_y0(h_u_cla32_and842_y0, h_u_cla32_and841_y0, h_u_cla32_and843_y0);
  and_gate and_gate_h_u_cla32_and844_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and844_y0);
  and_gate and_gate_h_u_cla32_and845_y0(h_u_cla32_and844_y0, h_u_cla32_and843_y0, h_u_cla32_and845_y0);
  and_gate and_gate_h_u_cla32_and846_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and846_y0);
  and_gate and_gate_h_u_cla32_and847_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and847_y0);
  and_gate and_gate_h_u_cla32_and848_y0(h_u_cla32_and847_y0, h_u_cla32_and846_y0, h_u_cla32_and848_y0);
  and_gate and_gate_h_u_cla32_and849_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and849_y0);
  and_gate and_gate_h_u_cla32_and850_y0(h_u_cla32_and849_y0, h_u_cla32_and848_y0, h_u_cla32_and850_y0);
  and_gate and_gate_h_u_cla32_and851_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and851_y0);
  and_gate and_gate_h_u_cla32_and852_y0(h_u_cla32_and851_y0, h_u_cla32_and850_y0, h_u_cla32_and852_y0);
  and_gate and_gate_h_u_cla32_and853_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and853_y0);
  and_gate and_gate_h_u_cla32_and854_y0(h_u_cla32_and853_y0, h_u_cla32_and852_y0, h_u_cla32_and854_y0);
  and_gate and_gate_h_u_cla32_and855_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and855_y0);
  and_gate and_gate_h_u_cla32_and856_y0(h_u_cla32_and855_y0, h_u_cla32_and854_y0, h_u_cla32_and856_y0);
  and_gate and_gate_h_u_cla32_and857_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and857_y0);
  and_gate and_gate_h_u_cla32_and858_y0(h_u_cla32_and857_y0, h_u_cla32_and856_y0, h_u_cla32_and858_y0);
  and_gate and_gate_h_u_cla32_and859_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and859_y0);
  and_gate and_gate_h_u_cla32_and860_y0(h_u_cla32_and859_y0, h_u_cla32_and858_y0, h_u_cla32_and860_y0);
  and_gate and_gate_h_u_cla32_and861_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and861_y0);
  and_gate and_gate_h_u_cla32_and862_y0(h_u_cla32_and861_y0, h_u_cla32_and860_y0, h_u_cla32_and862_y0);
  and_gate and_gate_h_u_cla32_and863_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and863_y0);
  and_gate and_gate_h_u_cla32_and864_y0(h_u_cla32_and863_y0, h_u_cla32_and862_y0, h_u_cla32_and864_y0);
  and_gate and_gate_h_u_cla32_and865_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and865_y0);
  and_gate and_gate_h_u_cla32_and866_y0(h_u_cla32_and865_y0, h_u_cla32_and864_y0, h_u_cla32_and866_y0);
  and_gate and_gate_h_u_cla32_and867_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and867_y0);
  and_gate and_gate_h_u_cla32_and868_y0(h_u_cla32_and867_y0, h_u_cla32_and866_y0, h_u_cla32_and868_y0);
  and_gate and_gate_h_u_cla32_and869_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and869_y0);
  and_gate and_gate_h_u_cla32_and870_y0(h_u_cla32_and869_y0, h_u_cla32_and868_y0, h_u_cla32_and870_y0);
  and_gate and_gate_h_u_cla32_and871_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and871_y0);
  and_gate and_gate_h_u_cla32_and872_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and872_y0);
  and_gate and_gate_h_u_cla32_and873_y0(h_u_cla32_and872_y0, h_u_cla32_and871_y0, h_u_cla32_and873_y0);
  and_gate and_gate_h_u_cla32_and874_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and874_y0);
  and_gate and_gate_h_u_cla32_and875_y0(h_u_cla32_and874_y0, h_u_cla32_and873_y0, h_u_cla32_and875_y0);
  and_gate and_gate_h_u_cla32_and876_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and876_y0);
  and_gate and_gate_h_u_cla32_and877_y0(h_u_cla32_and876_y0, h_u_cla32_and875_y0, h_u_cla32_and877_y0);
  and_gate and_gate_h_u_cla32_and878_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and878_y0);
  and_gate and_gate_h_u_cla32_and879_y0(h_u_cla32_and878_y0, h_u_cla32_and877_y0, h_u_cla32_and879_y0);
  and_gate and_gate_h_u_cla32_and880_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and880_y0);
  and_gate and_gate_h_u_cla32_and881_y0(h_u_cla32_and880_y0, h_u_cla32_and879_y0, h_u_cla32_and881_y0);
  and_gate and_gate_h_u_cla32_and882_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and882_y0);
  and_gate and_gate_h_u_cla32_and883_y0(h_u_cla32_and882_y0, h_u_cla32_and881_y0, h_u_cla32_and883_y0);
  and_gate and_gate_h_u_cla32_and884_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and884_y0);
  and_gate and_gate_h_u_cla32_and885_y0(h_u_cla32_and884_y0, h_u_cla32_and883_y0, h_u_cla32_and885_y0);
  and_gate and_gate_h_u_cla32_and886_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and886_y0);
  and_gate and_gate_h_u_cla32_and887_y0(h_u_cla32_and886_y0, h_u_cla32_and885_y0, h_u_cla32_and887_y0);
  and_gate and_gate_h_u_cla32_and888_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and888_y0);
  and_gate and_gate_h_u_cla32_and889_y0(h_u_cla32_and888_y0, h_u_cla32_and887_y0, h_u_cla32_and889_y0);
  and_gate and_gate_h_u_cla32_and890_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and890_y0);
  and_gate and_gate_h_u_cla32_and891_y0(h_u_cla32_and890_y0, h_u_cla32_and889_y0, h_u_cla32_and891_y0);
  and_gate and_gate_h_u_cla32_and892_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and892_y0);
  and_gate and_gate_h_u_cla32_and893_y0(h_u_cla32_and892_y0, h_u_cla32_and891_y0, h_u_cla32_and893_y0);
  and_gate and_gate_h_u_cla32_and894_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and894_y0);
  and_gate and_gate_h_u_cla32_and895_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and895_y0);
  and_gate and_gate_h_u_cla32_and896_y0(h_u_cla32_and895_y0, h_u_cla32_and894_y0, h_u_cla32_and896_y0);
  and_gate and_gate_h_u_cla32_and897_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and897_y0);
  and_gate and_gate_h_u_cla32_and898_y0(h_u_cla32_and897_y0, h_u_cla32_and896_y0, h_u_cla32_and898_y0);
  and_gate and_gate_h_u_cla32_and899_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and899_y0);
  and_gate and_gate_h_u_cla32_and900_y0(h_u_cla32_and899_y0, h_u_cla32_and898_y0, h_u_cla32_and900_y0);
  and_gate and_gate_h_u_cla32_and901_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and901_y0);
  and_gate and_gate_h_u_cla32_and902_y0(h_u_cla32_and901_y0, h_u_cla32_and900_y0, h_u_cla32_and902_y0);
  and_gate and_gate_h_u_cla32_and903_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and903_y0);
  and_gate and_gate_h_u_cla32_and904_y0(h_u_cla32_and903_y0, h_u_cla32_and902_y0, h_u_cla32_and904_y0);
  and_gate and_gate_h_u_cla32_and905_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and905_y0);
  and_gate and_gate_h_u_cla32_and906_y0(h_u_cla32_and905_y0, h_u_cla32_and904_y0, h_u_cla32_and906_y0);
  and_gate and_gate_h_u_cla32_and907_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and907_y0);
  and_gate and_gate_h_u_cla32_and908_y0(h_u_cla32_and907_y0, h_u_cla32_and906_y0, h_u_cla32_and908_y0);
  and_gate and_gate_h_u_cla32_and909_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and909_y0);
  and_gate and_gate_h_u_cla32_and910_y0(h_u_cla32_and909_y0, h_u_cla32_and908_y0, h_u_cla32_and910_y0);
  and_gate and_gate_h_u_cla32_and911_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and911_y0);
  and_gate and_gate_h_u_cla32_and912_y0(h_u_cla32_and911_y0, h_u_cla32_and910_y0, h_u_cla32_and912_y0);
  and_gate and_gate_h_u_cla32_and913_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and913_y0);
  and_gate and_gate_h_u_cla32_and914_y0(h_u_cla32_and913_y0, h_u_cla32_and912_y0, h_u_cla32_and914_y0);
  and_gate and_gate_h_u_cla32_and915_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and915_y0);
  and_gate and_gate_h_u_cla32_and916_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and916_y0);
  and_gate and_gate_h_u_cla32_and917_y0(h_u_cla32_and916_y0, h_u_cla32_and915_y0, h_u_cla32_and917_y0);
  and_gate and_gate_h_u_cla32_and918_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and918_y0);
  and_gate and_gate_h_u_cla32_and919_y0(h_u_cla32_and918_y0, h_u_cla32_and917_y0, h_u_cla32_and919_y0);
  and_gate and_gate_h_u_cla32_and920_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and920_y0);
  and_gate and_gate_h_u_cla32_and921_y0(h_u_cla32_and920_y0, h_u_cla32_and919_y0, h_u_cla32_and921_y0);
  and_gate and_gate_h_u_cla32_and922_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and922_y0);
  and_gate and_gate_h_u_cla32_and923_y0(h_u_cla32_and922_y0, h_u_cla32_and921_y0, h_u_cla32_and923_y0);
  and_gate and_gate_h_u_cla32_and924_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and924_y0);
  and_gate and_gate_h_u_cla32_and925_y0(h_u_cla32_and924_y0, h_u_cla32_and923_y0, h_u_cla32_and925_y0);
  and_gate and_gate_h_u_cla32_and926_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and926_y0);
  and_gate and_gate_h_u_cla32_and927_y0(h_u_cla32_and926_y0, h_u_cla32_and925_y0, h_u_cla32_and927_y0);
  and_gate and_gate_h_u_cla32_and928_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and928_y0);
  and_gate and_gate_h_u_cla32_and929_y0(h_u_cla32_and928_y0, h_u_cla32_and927_y0, h_u_cla32_and929_y0);
  and_gate and_gate_h_u_cla32_and930_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and930_y0);
  and_gate and_gate_h_u_cla32_and931_y0(h_u_cla32_and930_y0, h_u_cla32_and929_y0, h_u_cla32_and931_y0);
  and_gate and_gate_h_u_cla32_and932_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and932_y0);
  and_gate and_gate_h_u_cla32_and933_y0(h_u_cla32_and932_y0, h_u_cla32_and931_y0, h_u_cla32_and933_y0);
  and_gate and_gate_h_u_cla32_and934_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and934_y0);
  and_gate and_gate_h_u_cla32_and935_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and935_y0);
  and_gate and_gate_h_u_cla32_and936_y0(h_u_cla32_and935_y0, h_u_cla32_and934_y0, h_u_cla32_and936_y0);
  and_gate and_gate_h_u_cla32_and937_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and937_y0);
  and_gate and_gate_h_u_cla32_and938_y0(h_u_cla32_and937_y0, h_u_cla32_and936_y0, h_u_cla32_and938_y0);
  and_gate and_gate_h_u_cla32_and939_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and939_y0);
  and_gate and_gate_h_u_cla32_and940_y0(h_u_cla32_and939_y0, h_u_cla32_and938_y0, h_u_cla32_and940_y0);
  and_gate and_gate_h_u_cla32_and941_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and941_y0);
  and_gate and_gate_h_u_cla32_and942_y0(h_u_cla32_and941_y0, h_u_cla32_and940_y0, h_u_cla32_and942_y0);
  and_gate and_gate_h_u_cla32_and943_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and943_y0);
  and_gate and_gate_h_u_cla32_and944_y0(h_u_cla32_and943_y0, h_u_cla32_and942_y0, h_u_cla32_and944_y0);
  and_gate and_gate_h_u_cla32_and945_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and945_y0);
  and_gate and_gate_h_u_cla32_and946_y0(h_u_cla32_and945_y0, h_u_cla32_and944_y0, h_u_cla32_and946_y0);
  and_gate and_gate_h_u_cla32_and947_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and947_y0);
  and_gate and_gate_h_u_cla32_and948_y0(h_u_cla32_and947_y0, h_u_cla32_and946_y0, h_u_cla32_and948_y0);
  and_gate and_gate_h_u_cla32_and949_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and949_y0);
  and_gate and_gate_h_u_cla32_and950_y0(h_u_cla32_and949_y0, h_u_cla32_and948_y0, h_u_cla32_and950_y0);
  and_gate and_gate_h_u_cla32_and951_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and951_y0);
  and_gate and_gate_h_u_cla32_and952_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and952_y0);
  and_gate and_gate_h_u_cla32_and953_y0(h_u_cla32_and952_y0, h_u_cla32_and951_y0, h_u_cla32_and953_y0);
  and_gate and_gate_h_u_cla32_and954_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and954_y0);
  and_gate and_gate_h_u_cla32_and955_y0(h_u_cla32_and954_y0, h_u_cla32_and953_y0, h_u_cla32_and955_y0);
  and_gate and_gate_h_u_cla32_and956_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and956_y0);
  and_gate and_gate_h_u_cla32_and957_y0(h_u_cla32_and956_y0, h_u_cla32_and955_y0, h_u_cla32_and957_y0);
  and_gate and_gate_h_u_cla32_and958_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and958_y0);
  and_gate and_gate_h_u_cla32_and959_y0(h_u_cla32_and958_y0, h_u_cla32_and957_y0, h_u_cla32_and959_y0);
  and_gate and_gate_h_u_cla32_and960_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and960_y0);
  and_gate and_gate_h_u_cla32_and961_y0(h_u_cla32_and960_y0, h_u_cla32_and959_y0, h_u_cla32_and961_y0);
  and_gate and_gate_h_u_cla32_and962_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and962_y0);
  and_gate and_gate_h_u_cla32_and963_y0(h_u_cla32_and962_y0, h_u_cla32_and961_y0, h_u_cla32_and963_y0);
  and_gate and_gate_h_u_cla32_and964_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and964_y0);
  and_gate and_gate_h_u_cla32_and965_y0(h_u_cla32_and964_y0, h_u_cla32_and963_y0, h_u_cla32_and965_y0);
  and_gate and_gate_h_u_cla32_and966_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and966_y0);
  and_gate and_gate_h_u_cla32_and967_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and967_y0);
  and_gate and_gate_h_u_cla32_and968_y0(h_u_cla32_and967_y0, h_u_cla32_and966_y0, h_u_cla32_and968_y0);
  and_gate and_gate_h_u_cla32_and969_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and969_y0);
  and_gate and_gate_h_u_cla32_and970_y0(h_u_cla32_and969_y0, h_u_cla32_and968_y0, h_u_cla32_and970_y0);
  and_gate and_gate_h_u_cla32_and971_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and971_y0);
  and_gate and_gate_h_u_cla32_and972_y0(h_u_cla32_and971_y0, h_u_cla32_and970_y0, h_u_cla32_and972_y0);
  and_gate and_gate_h_u_cla32_and973_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and973_y0);
  and_gate and_gate_h_u_cla32_and974_y0(h_u_cla32_and973_y0, h_u_cla32_and972_y0, h_u_cla32_and974_y0);
  and_gate and_gate_h_u_cla32_and975_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and975_y0);
  and_gate and_gate_h_u_cla32_and976_y0(h_u_cla32_and975_y0, h_u_cla32_and974_y0, h_u_cla32_and976_y0);
  and_gate and_gate_h_u_cla32_and977_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and977_y0);
  and_gate and_gate_h_u_cla32_and978_y0(h_u_cla32_and977_y0, h_u_cla32_and976_y0, h_u_cla32_and978_y0);
  and_gate and_gate_h_u_cla32_and979_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and979_y0);
  and_gate and_gate_h_u_cla32_and980_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and980_y0);
  and_gate and_gate_h_u_cla32_and981_y0(h_u_cla32_and980_y0, h_u_cla32_and979_y0, h_u_cla32_and981_y0);
  and_gate and_gate_h_u_cla32_and982_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and982_y0);
  and_gate and_gate_h_u_cla32_and983_y0(h_u_cla32_and982_y0, h_u_cla32_and981_y0, h_u_cla32_and983_y0);
  and_gate and_gate_h_u_cla32_and984_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and984_y0);
  and_gate and_gate_h_u_cla32_and985_y0(h_u_cla32_and984_y0, h_u_cla32_and983_y0, h_u_cla32_and985_y0);
  and_gate and_gate_h_u_cla32_and986_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and986_y0);
  and_gate and_gate_h_u_cla32_and987_y0(h_u_cla32_and986_y0, h_u_cla32_and985_y0, h_u_cla32_and987_y0);
  and_gate and_gate_h_u_cla32_and988_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and988_y0);
  and_gate and_gate_h_u_cla32_and989_y0(h_u_cla32_and988_y0, h_u_cla32_and987_y0, h_u_cla32_and989_y0);
  and_gate and_gate_h_u_cla32_and990_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and990_y0);
  and_gate and_gate_h_u_cla32_and991_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and991_y0);
  and_gate and_gate_h_u_cla32_and992_y0(h_u_cla32_and991_y0, h_u_cla32_and990_y0, h_u_cla32_and992_y0);
  and_gate and_gate_h_u_cla32_and993_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and993_y0);
  and_gate and_gate_h_u_cla32_and994_y0(h_u_cla32_and993_y0, h_u_cla32_and992_y0, h_u_cla32_and994_y0);
  and_gate and_gate_h_u_cla32_and995_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and995_y0);
  and_gate and_gate_h_u_cla32_and996_y0(h_u_cla32_and995_y0, h_u_cla32_and994_y0, h_u_cla32_and996_y0);
  and_gate and_gate_h_u_cla32_and997_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and997_y0);
  and_gate and_gate_h_u_cla32_and998_y0(h_u_cla32_and997_y0, h_u_cla32_and996_y0, h_u_cla32_and998_y0);
  and_gate and_gate_h_u_cla32_and999_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and999_y0);
  and_gate and_gate_h_u_cla32_and1000_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1000_y0);
  and_gate and_gate_h_u_cla32_and1001_y0(h_u_cla32_and1000_y0, h_u_cla32_and999_y0, h_u_cla32_and1001_y0);
  and_gate and_gate_h_u_cla32_and1002_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1002_y0);
  and_gate and_gate_h_u_cla32_and1003_y0(h_u_cla32_and1002_y0, h_u_cla32_and1001_y0, h_u_cla32_and1003_y0);
  and_gate and_gate_h_u_cla32_and1004_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1004_y0);
  and_gate and_gate_h_u_cla32_and1005_y0(h_u_cla32_and1004_y0, h_u_cla32_and1003_y0, h_u_cla32_and1005_y0);
  and_gate and_gate_h_u_cla32_and1006_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1006_y0);
  and_gate and_gate_h_u_cla32_and1007_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1007_y0);
  and_gate and_gate_h_u_cla32_and1008_y0(h_u_cla32_and1007_y0, h_u_cla32_and1006_y0, h_u_cla32_and1008_y0);
  and_gate and_gate_h_u_cla32_and1009_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1009_y0);
  and_gate and_gate_h_u_cla32_and1010_y0(h_u_cla32_and1009_y0, h_u_cla32_and1008_y0, h_u_cla32_and1010_y0);
  and_gate and_gate_h_u_cla32_and1011_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1011_y0);
  and_gate and_gate_h_u_cla32_and1012_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1012_y0);
  and_gate and_gate_h_u_cla32_and1013_y0(h_u_cla32_and1012_y0, h_u_cla32_and1011_y0, h_u_cla32_and1013_y0);
  and_gate and_gate_h_u_cla32_and1014_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1014_y0);
  or_gate or_gate_h_u_cla32_or91_y0(h_u_cla32_and1014_y0, h_u_cla32_and845_y0, h_u_cla32_or91_y0);
  or_gate or_gate_h_u_cla32_or92_y0(h_u_cla32_or91_y0, h_u_cla32_and870_y0, h_u_cla32_or92_y0);
  or_gate or_gate_h_u_cla32_or93_y0(h_u_cla32_or92_y0, h_u_cla32_and893_y0, h_u_cla32_or93_y0);
  or_gate or_gate_h_u_cla32_or94_y0(h_u_cla32_or93_y0, h_u_cla32_and914_y0, h_u_cla32_or94_y0);
  or_gate or_gate_h_u_cla32_or95_y0(h_u_cla32_or94_y0, h_u_cla32_and933_y0, h_u_cla32_or95_y0);
  or_gate or_gate_h_u_cla32_or96_y0(h_u_cla32_or95_y0, h_u_cla32_and950_y0, h_u_cla32_or96_y0);
  or_gate or_gate_h_u_cla32_or97_y0(h_u_cla32_or96_y0, h_u_cla32_and965_y0, h_u_cla32_or97_y0);
  or_gate or_gate_h_u_cla32_or98_y0(h_u_cla32_or97_y0, h_u_cla32_and978_y0, h_u_cla32_or98_y0);
  or_gate or_gate_h_u_cla32_or99_y0(h_u_cla32_or98_y0, h_u_cla32_and989_y0, h_u_cla32_or99_y0);
  or_gate or_gate_h_u_cla32_or100_y0(h_u_cla32_or99_y0, h_u_cla32_and998_y0, h_u_cla32_or100_y0);
  or_gate or_gate_h_u_cla32_or101_y0(h_u_cla32_or100_y0, h_u_cla32_and1005_y0, h_u_cla32_or101_y0);
  or_gate or_gate_h_u_cla32_or102_y0(h_u_cla32_or101_y0, h_u_cla32_and1010_y0, h_u_cla32_or102_y0);
  or_gate or_gate_h_u_cla32_or103_y0(h_u_cla32_or102_y0, h_u_cla32_and1013_y0, h_u_cla32_or103_y0);
  or_gate or_gate_h_u_cla32_or104_y0(h_u_cla32_pg_logic13_y1, h_u_cla32_or103_y0, h_u_cla32_or104_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic14_y0(a_14, b_14, h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_pg_logic14_y2);
  xor_gate xor_gate_h_u_cla32_xor14_y0(h_u_cla32_pg_logic14_y2, h_u_cla32_or104_y0, h_u_cla32_xor14_y0);
  and_gate and_gate_h_u_cla32_and1015_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and1015_y0);
  and_gate and_gate_h_u_cla32_and1016_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and1016_y0);
  and_gate and_gate_h_u_cla32_and1017_y0(h_u_cla32_and1016_y0, h_u_cla32_and1015_y0, h_u_cla32_and1017_y0);
  and_gate and_gate_h_u_cla32_and1018_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and1018_y0);
  and_gate and_gate_h_u_cla32_and1019_y0(h_u_cla32_and1018_y0, h_u_cla32_and1017_y0, h_u_cla32_and1019_y0);
  and_gate and_gate_h_u_cla32_and1020_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and1020_y0);
  and_gate and_gate_h_u_cla32_and1021_y0(h_u_cla32_and1020_y0, h_u_cla32_and1019_y0, h_u_cla32_and1021_y0);
  and_gate and_gate_h_u_cla32_and1022_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and1022_y0);
  and_gate and_gate_h_u_cla32_and1023_y0(h_u_cla32_and1022_y0, h_u_cla32_and1021_y0, h_u_cla32_and1023_y0);
  and_gate and_gate_h_u_cla32_and1024_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and1024_y0);
  and_gate and_gate_h_u_cla32_and1025_y0(h_u_cla32_and1024_y0, h_u_cla32_and1023_y0, h_u_cla32_and1025_y0);
  and_gate and_gate_h_u_cla32_and1026_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and1026_y0);
  and_gate and_gate_h_u_cla32_and1027_y0(h_u_cla32_and1026_y0, h_u_cla32_and1025_y0, h_u_cla32_and1027_y0);
  and_gate and_gate_h_u_cla32_and1028_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and1028_y0);
  and_gate and_gate_h_u_cla32_and1029_y0(h_u_cla32_and1028_y0, h_u_cla32_and1027_y0, h_u_cla32_and1029_y0);
  and_gate and_gate_h_u_cla32_and1030_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and1030_y0);
  and_gate and_gate_h_u_cla32_and1031_y0(h_u_cla32_and1030_y0, h_u_cla32_and1029_y0, h_u_cla32_and1031_y0);
  and_gate and_gate_h_u_cla32_and1032_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and1032_y0);
  and_gate and_gate_h_u_cla32_and1033_y0(h_u_cla32_and1032_y0, h_u_cla32_and1031_y0, h_u_cla32_and1033_y0);
  and_gate and_gate_h_u_cla32_and1034_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and1034_y0);
  and_gate and_gate_h_u_cla32_and1035_y0(h_u_cla32_and1034_y0, h_u_cla32_and1033_y0, h_u_cla32_and1035_y0);
  and_gate and_gate_h_u_cla32_and1036_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and1036_y0);
  and_gate and_gate_h_u_cla32_and1037_y0(h_u_cla32_and1036_y0, h_u_cla32_and1035_y0, h_u_cla32_and1037_y0);
  and_gate and_gate_h_u_cla32_and1038_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and1038_y0);
  and_gate and_gate_h_u_cla32_and1039_y0(h_u_cla32_and1038_y0, h_u_cla32_and1037_y0, h_u_cla32_and1039_y0);
  and_gate and_gate_h_u_cla32_and1040_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and1040_y0);
  and_gate and_gate_h_u_cla32_and1041_y0(h_u_cla32_and1040_y0, h_u_cla32_and1039_y0, h_u_cla32_and1041_y0);
  and_gate and_gate_h_u_cla32_and1042_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and1042_y0);
  and_gate and_gate_h_u_cla32_and1043_y0(h_u_cla32_and1042_y0, h_u_cla32_and1041_y0, h_u_cla32_and1043_y0);
  and_gate and_gate_h_u_cla32_and1044_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1044_y0);
  and_gate and_gate_h_u_cla32_and1045_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1045_y0);
  and_gate and_gate_h_u_cla32_and1046_y0(h_u_cla32_and1045_y0, h_u_cla32_and1044_y0, h_u_cla32_and1046_y0);
  and_gate and_gate_h_u_cla32_and1047_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1047_y0);
  and_gate and_gate_h_u_cla32_and1048_y0(h_u_cla32_and1047_y0, h_u_cla32_and1046_y0, h_u_cla32_and1048_y0);
  and_gate and_gate_h_u_cla32_and1049_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1049_y0);
  and_gate and_gate_h_u_cla32_and1050_y0(h_u_cla32_and1049_y0, h_u_cla32_and1048_y0, h_u_cla32_and1050_y0);
  and_gate and_gate_h_u_cla32_and1051_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1051_y0);
  and_gate and_gate_h_u_cla32_and1052_y0(h_u_cla32_and1051_y0, h_u_cla32_and1050_y0, h_u_cla32_and1052_y0);
  and_gate and_gate_h_u_cla32_and1053_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1053_y0);
  and_gate and_gate_h_u_cla32_and1054_y0(h_u_cla32_and1053_y0, h_u_cla32_and1052_y0, h_u_cla32_and1054_y0);
  and_gate and_gate_h_u_cla32_and1055_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1055_y0);
  and_gate and_gate_h_u_cla32_and1056_y0(h_u_cla32_and1055_y0, h_u_cla32_and1054_y0, h_u_cla32_and1056_y0);
  and_gate and_gate_h_u_cla32_and1057_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1057_y0);
  and_gate and_gate_h_u_cla32_and1058_y0(h_u_cla32_and1057_y0, h_u_cla32_and1056_y0, h_u_cla32_and1058_y0);
  and_gate and_gate_h_u_cla32_and1059_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1059_y0);
  and_gate and_gate_h_u_cla32_and1060_y0(h_u_cla32_and1059_y0, h_u_cla32_and1058_y0, h_u_cla32_and1060_y0);
  and_gate and_gate_h_u_cla32_and1061_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1061_y0);
  and_gate and_gate_h_u_cla32_and1062_y0(h_u_cla32_and1061_y0, h_u_cla32_and1060_y0, h_u_cla32_and1062_y0);
  and_gate and_gate_h_u_cla32_and1063_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1063_y0);
  and_gate and_gate_h_u_cla32_and1064_y0(h_u_cla32_and1063_y0, h_u_cla32_and1062_y0, h_u_cla32_and1064_y0);
  and_gate and_gate_h_u_cla32_and1065_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1065_y0);
  and_gate and_gate_h_u_cla32_and1066_y0(h_u_cla32_and1065_y0, h_u_cla32_and1064_y0, h_u_cla32_and1066_y0);
  and_gate and_gate_h_u_cla32_and1067_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1067_y0);
  and_gate and_gate_h_u_cla32_and1068_y0(h_u_cla32_and1067_y0, h_u_cla32_and1066_y0, h_u_cla32_and1068_y0);
  and_gate and_gate_h_u_cla32_and1069_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1069_y0);
  and_gate and_gate_h_u_cla32_and1070_y0(h_u_cla32_and1069_y0, h_u_cla32_and1068_y0, h_u_cla32_and1070_y0);
  and_gate and_gate_h_u_cla32_and1071_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1071_y0);
  and_gate and_gate_h_u_cla32_and1072_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1072_y0);
  and_gate and_gate_h_u_cla32_and1073_y0(h_u_cla32_and1072_y0, h_u_cla32_and1071_y0, h_u_cla32_and1073_y0);
  and_gate and_gate_h_u_cla32_and1074_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1074_y0);
  and_gate and_gate_h_u_cla32_and1075_y0(h_u_cla32_and1074_y0, h_u_cla32_and1073_y0, h_u_cla32_and1075_y0);
  and_gate and_gate_h_u_cla32_and1076_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1076_y0);
  and_gate and_gate_h_u_cla32_and1077_y0(h_u_cla32_and1076_y0, h_u_cla32_and1075_y0, h_u_cla32_and1077_y0);
  and_gate and_gate_h_u_cla32_and1078_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1078_y0);
  and_gate and_gate_h_u_cla32_and1079_y0(h_u_cla32_and1078_y0, h_u_cla32_and1077_y0, h_u_cla32_and1079_y0);
  and_gate and_gate_h_u_cla32_and1080_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1080_y0);
  and_gate and_gate_h_u_cla32_and1081_y0(h_u_cla32_and1080_y0, h_u_cla32_and1079_y0, h_u_cla32_and1081_y0);
  and_gate and_gate_h_u_cla32_and1082_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1082_y0);
  and_gate and_gate_h_u_cla32_and1083_y0(h_u_cla32_and1082_y0, h_u_cla32_and1081_y0, h_u_cla32_and1083_y0);
  and_gate and_gate_h_u_cla32_and1084_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1084_y0);
  and_gate and_gate_h_u_cla32_and1085_y0(h_u_cla32_and1084_y0, h_u_cla32_and1083_y0, h_u_cla32_and1085_y0);
  and_gate and_gate_h_u_cla32_and1086_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1086_y0);
  and_gate and_gate_h_u_cla32_and1087_y0(h_u_cla32_and1086_y0, h_u_cla32_and1085_y0, h_u_cla32_and1087_y0);
  and_gate and_gate_h_u_cla32_and1088_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1088_y0);
  and_gate and_gate_h_u_cla32_and1089_y0(h_u_cla32_and1088_y0, h_u_cla32_and1087_y0, h_u_cla32_and1089_y0);
  and_gate and_gate_h_u_cla32_and1090_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1090_y0);
  and_gate and_gate_h_u_cla32_and1091_y0(h_u_cla32_and1090_y0, h_u_cla32_and1089_y0, h_u_cla32_and1091_y0);
  and_gate and_gate_h_u_cla32_and1092_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1092_y0);
  and_gate and_gate_h_u_cla32_and1093_y0(h_u_cla32_and1092_y0, h_u_cla32_and1091_y0, h_u_cla32_and1093_y0);
  and_gate and_gate_h_u_cla32_and1094_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1094_y0);
  and_gate and_gate_h_u_cla32_and1095_y0(h_u_cla32_and1094_y0, h_u_cla32_and1093_y0, h_u_cla32_and1095_y0);
  and_gate and_gate_h_u_cla32_and1096_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1096_y0);
  and_gate and_gate_h_u_cla32_and1097_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1097_y0);
  and_gate and_gate_h_u_cla32_and1098_y0(h_u_cla32_and1097_y0, h_u_cla32_and1096_y0, h_u_cla32_and1098_y0);
  and_gate and_gate_h_u_cla32_and1099_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1099_y0);
  and_gate and_gate_h_u_cla32_and1100_y0(h_u_cla32_and1099_y0, h_u_cla32_and1098_y0, h_u_cla32_and1100_y0);
  and_gate and_gate_h_u_cla32_and1101_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1101_y0);
  and_gate and_gate_h_u_cla32_and1102_y0(h_u_cla32_and1101_y0, h_u_cla32_and1100_y0, h_u_cla32_and1102_y0);
  and_gate and_gate_h_u_cla32_and1103_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1103_y0);
  and_gate and_gate_h_u_cla32_and1104_y0(h_u_cla32_and1103_y0, h_u_cla32_and1102_y0, h_u_cla32_and1104_y0);
  and_gate and_gate_h_u_cla32_and1105_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1105_y0);
  and_gate and_gate_h_u_cla32_and1106_y0(h_u_cla32_and1105_y0, h_u_cla32_and1104_y0, h_u_cla32_and1106_y0);
  and_gate and_gate_h_u_cla32_and1107_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1107_y0);
  and_gate and_gate_h_u_cla32_and1108_y0(h_u_cla32_and1107_y0, h_u_cla32_and1106_y0, h_u_cla32_and1108_y0);
  and_gate and_gate_h_u_cla32_and1109_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1109_y0);
  and_gate and_gate_h_u_cla32_and1110_y0(h_u_cla32_and1109_y0, h_u_cla32_and1108_y0, h_u_cla32_and1110_y0);
  and_gate and_gate_h_u_cla32_and1111_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1111_y0);
  and_gate and_gate_h_u_cla32_and1112_y0(h_u_cla32_and1111_y0, h_u_cla32_and1110_y0, h_u_cla32_and1112_y0);
  and_gate and_gate_h_u_cla32_and1113_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1113_y0);
  and_gate and_gate_h_u_cla32_and1114_y0(h_u_cla32_and1113_y0, h_u_cla32_and1112_y0, h_u_cla32_and1114_y0);
  and_gate and_gate_h_u_cla32_and1115_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1115_y0);
  and_gate and_gate_h_u_cla32_and1116_y0(h_u_cla32_and1115_y0, h_u_cla32_and1114_y0, h_u_cla32_and1116_y0);
  and_gate and_gate_h_u_cla32_and1117_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1117_y0);
  and_gate and_gate_h_u_cla32_and1118_y0(h_u_cla32_and1117_y0, h_u_cla32_and1116_y0, h_u_cla32_and1118_y0);
  and_gate and_gate_h_u_cla32_and1119_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1119_y0);
  and_gate and_gate_h_u_cla32_and1120_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1120_y0);
  and_gate and_gate_h_u_cla32_and1121_y0(h_u_cla32_and1120_y0, h_u_cla32_and1119_y0, h_u_cla32_and1121_y0);
  and_gate and_gate_h_u_cla32_and1122_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1122_y0);
  and_gate and_gate_h_u_cla32_and1123_y0(h_u_cla32_and1122_y0, h_u_cla32_and1121_y0, h_u_cla32_and1123_y0);
  and_gate and_gate_h_u_cla32_and1124_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1124_y0);
  and_gate and_gate_h_u_cla32_and1125_y0(h_u_cla32_and1124_y0, h_u_cla32_and1123_y0, h_u_cla32_and1125_y0);
  and_gate and_gate_h_u_cla32_and1126_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1126_y0);
  and_gate and_gate_h_u_cla32_and1127_y0(h_u_cla32_and1126_y0, h_u_cla32_and1125_y0, h_u_cla32_and1127_y0);
  and_gate and_gate_h_u_cla32_and1128_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1128_y0);
  and_gate and_gate_h_u_cla32_and1129_y0(h_u_cla32_and1128_y0, h_u_cla32_and1127_y0, h_u_cla32_and1129_y0);
  and_gate and_gate_h_u_cla32_and1130_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1130_y0);
  and_gate and_gate_h_u_cla32_and1131_y0(h_u_cla32_and1130_y0, h_u_cla32_and1129_y0, h_u_cla32_and1131_y0);
  and_gate and_gate_h_u_cla32_and1132_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1132_y0);
  and_gate and_gate_h_u_cla32_and1133_y0(h_u_cla32_and1132_y0, h_u_cla32_and1131_y0, h_u_cla32_and1133_y0);
  and_gate and_gate_h_u_cla32_and1134_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1134_y0);
  and_gate and_gate_h_u_cla32_and1135_y0(h_u_cla32_and1134_y0, h_u_cla32_and1133_y0, h_u_cla32_and1135_y0);
  and_gate and_gate_h_u_cla32_and1136_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1136_y0);
  and_gate and_gate_h_u_cla32_and1137_y0(h_u_cla32_and1136_y0, h_u_cla32_and1135_y0, h_u_cla32_and1137_y0);
  and_gate and_gate_h_u_cla32_and1138_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1138_y0);
  and_gate and_gate_h_u_cla32_and1139_y0(h_u_cla32_and1138_y0, h_u_cla32_and1137_y0, h_u_cla32_and1139_y0);
  and_gate and_gate_h_u_cla32_and1140_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1140_y0);
  and_gate and_gate_h_u_cla32_and1141_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1141_y0);
  and_gate and_gate_h_u_cla32_and1142_y0(h_u_cla32_and1141_y0, h_u_cla32_and1140_y0, h_u_cla32_and1142_y0);
  and_gate and_gate_h_u_cla32_and1143_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1143_y0);
  and_gate and_gate_h_u_cla32_and1144_y0(h_u_cla32_and1143_y0, h_u_cla32_and1142_y0, h_u_cla32_and1144_y0);
  and_gate and_gate_h_u_cla32_and1145_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1145_y0);
  and_gate and_gate_h_u_cla32_and1146_y0(h_u_cla32_and1145_y0, h_u_cla32_and1144_y0, h_u_cla32_and1146_y0);
  and_gate and_gate_h_u_cla32_and1147_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1147_y0);
  and_gate and_gate_h_u_cla32_and1148_y0(h_u_cla32_and1147_y0, h_u_cla32_and1146_y0, h_u_cla32_and1148_y0);
  and_gate and_gate_h_u_cla32_and1149_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1149_y0);
  and_gate and_gate_h_u_cla32_and1150_y0(h_u_cla32_and1149_y0, h_u_cla32_and1148_y0, h_u_cla32_and1150_y0);
  and_gate and_gate_h_u_cla32_and1151_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1151_y0);
  and_gate and_gate_h_u_cla32_and1152_y0(h_u_cla32_and1151_y0, h_u_cla32_and1150_y0, h_u_cla32_and1152_y0);
  and_gate and_gate_h_u_cla32_and1153_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1153_y0);
  and_gate and_gate_h_u_cla32_and1154_y0(h_u_cla32_and1153_y0, h_u_cla32_and1152_y0, h_u_cla32_and1154_y0);
  and_gate and_gate_h_u_cla32_and1155_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1155_y0);
  and_gate and_gate_h_u_cla32_and1156_y0(h_u_cla32_and1155_y0, h_u_cla32_and1154_y0, h_u_cla32_and1156_y0);
  and_gate and_gate_h_u_cla32_and1157_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1157_y0);
  and_gate and_gate_h_u_cla32_and1158_y0(h_u_cla32_and1157_y0, h_u_cla32_and1156_y0, h_u_cla32_and1158_y0);
  and_gate and_gate_h_u_cla32_and1159_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1159_y0);
  and_gate and_gate_h_u_cla32_and1160_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1160_y0);
  and_gate and_gate_h_u_cla32_and1161_y0(h_u_cla32_and1160_y0, h_u_cla32_and1159_y0, h_u_cla32_and1161_y0);
  and_gate and_gate_h_u_cla32_and1162_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1162_y0);
  and_gate and_gate_h_u_cla32_and1163_y0(h_u_cla32_and1162_y0, h_u_cla32_and1161_y0, h_u_cla32_and1163_y0);
  and_gate and_gate_h_u_cla32_and1164_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1164_y0);
  and_gate and_gate_h_u_cla32_and1165_y0(h_u_cla32_and1164_y0, h_u_cla32_and1163_y0, h_u_cla32_and1165_y0);
  and_gate and_gate_h_u_cla32_and1166_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1166_y0);
  and_gate and_gate_h_u_cla32_and1167_y0(h_u_cla32_and1166_y0, h_u_cla32_and1165_y0, h_u_cla32_and1167_y0);
  and_gate and_gate_h_u_cla32_and1168_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1168_y0);
  and_gate and_gate_h_u_cla32_and1169_y0(h_u_cla32_and1168_y0, h_u_cla32_and1167_y0, h_u_cla32_and1169_y0);
  and_gate and_gate_h_u_cla32_and1170_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1170_y0);
  and_gate and_gate_h_u_cla32_and1171_y0(h_u_cla32_and1170_y0, h_u_cla32_and1169_y0, h_u_cla32_and1171_y0);
  and_gate and_gate_h_u_cla32_and1172_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1172_y0);
  and_gate and_gate_h_u_cla32_and1173_y0(h_u_cla32_and1172_y0, h_u_cla32_and1171_y0, h_u_cla32_and1173_y0);
  and_gate and_gate_h_u_cla32_and1174_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1174_y0);
  and_gate and_gate_h_u_cla32_and1175_y0(h_u_cla32_and1174_y0, h_u_cla32_and1173_y0, h_u_cla32_and1175_y0);
  and_gate and_gate_h_u_cla32_and1176_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1176_y0);
  and_gate and_gate_h_u_cla32_and1177_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1177_y0);
  and_gate and_gate_h_u_cla32_and1178_y0(h_u_cla32_and1177_y0, h_u_cla32_and1176_y0, h_u_cla32_and1178_y0);
  and_gate and_gate_h_u_cla32_and1179_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1179_y0);
  and_gate and_gate_h_u_cla32_and1180_y0(h_u_cla32_and1179_y0, h_u_cla32_and1178_y0, h_u_cla32_and1180_y0);
  and_gate and_gate_h_u_cla32_and1181_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1181_y0);
  and_gate and_gate_h_u_cla32_and1182_y0(h_u_cla32_and1181_y0, h_u_cla32_and1180_y0, h_u_cla32_and1182_y0);
  and_gate and_gate_h_u_cla32_and1183_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1183_y0);
  and_gate and_gate_h_u_cla32_and1184_y0(h_u_cla32_and1183_y0, h_u_cla32_and1182_y0, h_u_cla32_and1184_y0);
  and_gate and_gate_h_u_cla32_and1185_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1185_y0);
  and_gate and_gate_h_u_cla32_and1186_y0(h_u_cla32_and1185_y0, h_u_cla32_and1184_y0, h_u_cla32_and1186_y0);
  and_gate and_gate_h_u_cla32_and1187_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1187_y0);
  and_gate and_gate_h_u_cla32_and1188_y0(h_u_cla32_and1187_y0, h_u_cla32_and1186_y0, h_u_cla32_and1188_y0);
  and_gate and_gate_h_u_cla32_and1189_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1189_y0);
  and_gate and_gate_h_u_cla32_and1190_y0(h_u_cla32_and1189_y0, h_u_cla32_and1188_y0, h_u_cla32_and1190_y0);
  and_gate and_gate_h_u_cla32_and1191_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1191_y0);
  and_gate and_gate_h_u_cla32_and1192_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1192_y0);
  and_gate and_gate_h_u_cla32_and1193_y0(h_u_cla32_and1192_y0, h_u_cla32_and1191_y0, h_u_cla32_and1193_y0);
  and_gate and_gate_h_u_cla32_and1194_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1194_y0);
  and_gate and_gate_h_u_cla32_and1195_y0(h_u_cla32_and1194_y0, h_u_cla32_and1193_y0, h_u_cla32_and1195_y0);
  and_gate and_gate_h_u_cla32_and1196_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1196_y0);
  and_gate and_gate_h_u_cla32_and1197_y0(h_u_cla32_and1196_y0, h_u_cla32_and1195_y0, h_u_cla32_and1197_y0);
  and_gate and_gate_h_u_cla32_and1198_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1198_y0);
  and_gate and_gate_h_u_cla32_and1199_y0(h_u_cla32_and1198_y0, h_u_cla32_and1197_y0, h_u_cla32_and1199_y0);
  and_gate and_gate_h_u_cla32_and1200_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1200_y0);
  and_gate and_gate_h_u_cla32_and1201_y0(h_u_cla32_and1200_y0, h_u_cla32_and1199_y0, h_u_cla32_and1201_y0);
  and_gate and_gate_h_u_cla32_and1202_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1202_y0);
  and_gate and_gate_h_u_cla32_and1203_y0(h_u_cla32_and1202_y0, h_u_cla32_and1201_y0, h_u_cla32_and1203_y0);
  and_gate and_gate_h_u_cla32_and1204_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1204_y0);
  and_gate and_gate_h_u_cla32_and1205_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1205_y0);
  and_gate and_gate_h_u_cla32_and1206_y0(h_u_cla32_and1205_y0, h_u_cla32_and1204_y0, h_u_cla32_and1206_y0);
  and_gate and_gate_h_u_cla32_and1207_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1207_y0);
  and_gate and_gate_h_u_cla32_and1208_y0(h_u_cla32_and1207_y0, h_u_cla32_and1206_y0, h_u_cla32_and1208_y0);
  and_gate and_gate_h_u_cla32_and1209_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1209_y0);
  and_gate and_gate_h_u_cla32_and1210_y0(h_u_cla32_and1209_y0, h_u_cla32_and1208_y0, h_u_cla32_and1210_y0);
  and_gate and_gate_h_u_cla32_and1211_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1211_y0);
  and_gate and_gate_h_u_cla32_and1212_y0(h_u_cla32_and1211_y0, h_u_cla32_and1210_y0, h_u_cla32_and1212_y0);
  and_gate and_gate_h_u_cla32_and1213_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1213_y0);
  and_gate and_gate_h_u_cla32_and1214_y0(h_u_cla32_and1213_y0, h_u_cla32_and1212_y0, h_u_cla32_and1214_y0);
  and_gate and_gate_h_u_cla32_and1215_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1215_y0);
  and_gate and_gate_h_u_cla32_and1216_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1216_y0);
  and_gate and_gate_h_u_cla32_and1217_y0(h_u_cla32_and1216_y0, h_u_cla32_and1215_y0, h_u_cla32_and1217_y0);
  and_gate and_gate_h_u_cla32_and1218_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1218_y0);
  and_gate and_gate_h_u_cla32_and1219_y0(h_u_cla32_and1218_y0, h_u_cla32_and1217_y0, h_u_cla32_and1219_y0);
  and_gate and_gate_h_u_cla32_and1220_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1220_y0);
  and_gate and_gate_h_u_cla32_and1221_y0(h_u_cla32_and1220_y0, h_u_cla32_and1219_y0, h_u_cla32_and1221_y0);
  and_gate and_gate_h_u_cla32_and1222_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1222_y0);
  and_gate and_gate_h_u_cla32_and1223_y0(h_u_cla32_and1222_y0, h_u_cla32_and1221_y0, h_u_cla32_and1223_y0);
  and_gate and_gate_h_u_cla32_and1224_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1224_y0);
  and_gate and_gate_h_u_cla32_and1225_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1225_y0);
  and_gate and_gate_h_u_cla32_and1226_y0(h_u_cla32_and1225_y0, h_u_cla32_and1224_y0, h_u_cla32_and1226_y0);
  and_gate and_gate_h_u_cla32_and1227_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1227_y0);
  and_gate and_gate_h_u_cla32_and1228_y0(h_u_cla32_and1227_y0, h_u_cla32_and1226_y0, h_u_cla32_and1228_y0);
  and_gate and_gate_h_u_cla32_and1229_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1229_y0);
  and_gate and_gate_h_u_cla32_and1230_y0(h_u_cla32_and1229_y0, h_u_cla32_and1228_y0, h_u_cla32_and1230_y0);
  and_gate and_gate_h_u_cla32_and1231_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1231_y0);
  and_gate and_gate_h_u_cla32_and1232_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1232_y0);
  and_gate and_gate_h_u_cla32_and1233_y0(h_u_cla32_and1232_y0, h_u_cla32_and1231_y0, h_u_cla32_and1233_y0);
  and_gate and_gate_h_u_cla32_and1234_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1234_y0);
  and_gate and_gate_h_u_cla32_and1235_y0(h_u_cla32_and1234_y0, h_u_cla32_and1233_y0, h_u_cla32_and1235_y0);
  and_gate and_gate_h_u_cla32_and1236_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1236_y0);
  and_gate and_gate_h_u_cla32_and1237_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1237_y0);
  and_gate and_gate_h_u_cla32_and1238_y0(h_u_cla32_and1237_y0, h_u_cla32_and1236_y0, h_u_cla32_and1238_y0);
  and_gate and_gate_h_u_cla32_and1239_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and1239_y0);
  or_gate or_gate_h_u_cla32_or105_y0(h_u_cla32_and1239_y0, h_u_cla32_and1043_y0, h_u_cla32_or105_y0);
  or_gate or_gate_h_u_cla32_or106_y0(h_u_cla32_or105_y0, h_u_cla32_and1070_y0, h_u_cla32_or106_y0);
  or_gate or_gate_h_u_cla32_or107_y0(h_u_cla32_or106_y0, h_u_cla32_and1095_y0, h_u_cla32_or107_y0);
  or_gate or_gate_h_u_cla32_or108_y0(h_u_cla32_or107_y0, h_u_cla32_and1118_y0, h_u_cla32_or108_y0);
  or_gate or_gate_h_u_cla32_or109_y0(h_u_cla32_or108_y0, h_u_cla32_and1139_y0, h_u_cla32_or109_y0);
  or_gate or_gate_h_u_cla32_or110_y0(h_u_cla32_or109_y0, h_u_cla32_and1158_y0, h_u_cla32_or110_y0);
  or_gate or_gate_h_u_cla32_or111_y0(h_u_cla32_or110_y0, h_u_cla32_and1175_y0, h_u_cla32_or111_y0);
  or_gate or_gate_h_u_cla32_or112_y0(h_u_cla32_or111_y0, h_u_cla32_and1190_y0, h_u_cla32_or112_y0);
  or_gate or_gate_h_u_cla32_or113_y0(h_u_cla32_or112_y0, h_u_cla32_and1203_y0, h_u_cla32_or113_y0);
  or_gate or_gate_h_u_cla32_or114_y0(h_u_cla32_or113_y0, h_u_cla32_and1214_y0, h_u_cla32_or114_y0);
  or_gate or_gate_h_u_cla32_or115_y0(h_u_cla32_or114_y0, h_u_cla32_and1223_y0, h_u_cla32_or115_y0);
  or_gate or_gate_h_u_cla32_or116_y0(h_u_cla32_or115_y0, h_u_cla32_and1230_y0, h_u_cla32_or116_y0);
  or_gate or_gate_h_u_cla32_or117_y0(h_u_cla32_or116_y0, h_u_cla32_and1235_y0, h_u_cla32_or117_y0);
  or_gate or_gate_h_u_cla32_or118_y0(h_u_cla32_or117_y0, h_u_cla32_and1238_y0, h_u_cla32_or118_y0);
  or_gate or_gate_h_u_cla32_or119_y0(h_u_cla32_pg_logic14_y1, h_u_cla32_or118_y0, h_u_cla32_or119_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic15_y0(a_15, b_15, h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_pg_logic15_y2);
  xor_gate xor_gate_h_u_cla32_xor15_y0(h_u_cla32_pg_logic15_y2, h_u_cla32_or119_y0, h_u_cla32_xor15_y0);
  and_gate and_gate_h_u_cla32_and1240_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and1240_y0);
  and_gate and_gate_h_u_cla32_and1241_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and1241_y0);
  and_gate and_gate_h_u_cla32_and1242_y0(h_u_cla32_and1241_y0, h_u_cla32_and1240_y0, h_u_cla32_and1242_y0);
  and_gate and_gate_h_u_cla32_and1243_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and1243_y0);
  and_gate and_gate_h_u_cla32_and1244_y0(h_u_cla32_and1243_y0, h_u_cla32_and1242_y0, h_u_cla32_and1244_y0);
  and_gate and_gate_h_u_cla32_and1245_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and1245_y0);
  and_gate and_gate_h_u_cla32_and1246_y0(h_u_cla32_and1245_y0, h_u_cla32_and1244_y0, h_u_cla32_and1246_y0);
  and_gate and_gate_h_u_cla32_and1247_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and1247_y0);
  and_gate and_gate_h_u_cla32_and1248_y0(h_u_cla32_and1247_y0, h_u_cla32_and1246_y0, h_u_cla32_and1248_y0);
  and_gate and_gate_h_u_cla32_and1249_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and1249_y0);
  and_gate and_gate_h_u_cla32_and1250_y0(h_u_cla32_and1249_y0, h_u_cla32_and1248_y0, h_u_cla32_and1250_y0);
  and_gate and_gate_h_u_cla32_and1251_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and1251_y0);
  and_gate and_gate_h_u_cla32_and1252_y0(h_u_cla32_and1251_y0, h_u_cla32_and1250_y0, h_u_cla32_and1252_y0);
  and_gate and_gate_h_u_cla32_and1253_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and1253_y0);
  and_gate and_gate_h_u_cla32_and1254_y0(h_u_cla32_and1253_y0, h_u_cla32_and1252_y0, h_u_cla32_and1254_y0);
  and_gate and_gate_h_u_cla32_and1255_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and1255_y0);
  and_gate and_gate_h_u_cla32_and1256_y0(h_u_cla32_and1255_y0, h_u_cla32_and1254_y0, h_u_cla32_and1256_y0);
  and_gate and_gate_h_u_cla32_and1257_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and1257_y0);
  and_gate and_gate_h_u_cla32_and1258_y0(h_u_cla32_and1257_y0, h_u_cla32_and1256_y0, h_u_cla32_and1258_y0);
  and_gate and_gate_h_u_cla32_and1259_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and1259_y0);
  and_gate and_gate_h_u_cla32_and1260_y0(h_u_cla32_and1259_y0, h_u_cla32_and1258_y0, h_u_cla32_and1260_y0);
  and_gate and_gate_h_u_cla32_and1261_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and1261_y0);
  and_gate and_gate_h_u_cla32_and1262_y0(h_u_cla32_and1261_y0, h_u_cla32_and1260_y0, h_u_cla32_and1262_y0);
  and_gate and_gate_h_u_cla32_and1263_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and1263_y0);
  and_gate and_gate_h_u_cla32_and1264_y0(h_u_cla32_and1263_y0, h_u_cla32_and1262_y0, h_u_cla32_and1264_y0);
  and_gate and_gate_h_u_cla32_and1265_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and1265_y0);
  and_gate and_gate_h_u_cla32_and1266_y0(h_u_cla32_and1265_y0, h_u_cla32_and1264_y0, h_u_cla32_and1266_y0);
  and_gate and_gate_h_u_cla32_and1267_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and1267_y0);
  and_gate and_gate_h_u_cla32_and1268_y0(h_u_cla32_and1267_y0, h_u_cla32_and1266_y0, h_u_cla32_and1268_y0);
  and_gate and_gate_h_u_cla32_and1269_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and1269_y0);
  and_gate and_gate_h_u_cla32_and1270_y0(h_u_cla32_and1269_y0, h_u_cla32_and1268_y0, h_u_cla32_and1270_y0);
  and_gate and_gate_h_u_cla32_and1271_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1271_y0);
  and_gate and_gate_h_u_cla32_and1272_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1272_y0);
  and_gate and_gate_h_u_cla32_and1273_y0(h_u_cla32_and1272_y0, h_u_cla32_and1271_y0, h_u_cla32_and1273_y0);
  and_gate and_gate_h_u_cla32_and1274_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1274_y0);
  and_gate and_gate_h_u_cla32_and1275_y0(h_u_cla32_and1274_y0, h_u_cla32_and1273_y0, h_u_cla32_and1275_y0);
  and_gate and_gate_h_u_cla32_and1276_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1276_y0);
  and_gate and_gate_h_u_cla32_and1277_y0(h_u_cla32_and1276_y0, h_u_cla32_and1275_y0, h_u_cla32_and1277_y0);
  and_gate and_gate_h_u_cla32_and1278_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1278_y0);
  and_gate and_gate_h_u_cla32_and1279_y0(h_u_cla32_and1278_y0, h_u_cla32_and1277_y0, h_u_cla32_and1279_y0);
  and_gate and_gate_h_u_cla32_and1280_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1280_y0);
  and_gate and_gate_h_u_cla32_and1281_y0(h_u_cla32_and1280_y0, h_u_cla32_and1279_y0, h_u_cla32_and1281_y0);
  and_gate and_gate_h_u_cla32_and1282_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1282_y0);
  and_gate and_gate_h_u_cla32_and1283_y0(h_u_cla32_and1282_y0, h_u_cla32_and1281_y0, h_u_cla32_and1283_y0);
  and_gate and_gate_h_u_cla32_and1284_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1284_y0);
  and_gate and_gate_h_u_cla32_and1285_y0(h_u_cla32_and1284_y0, h_u_cla32_and1283_y0, h_u_cla32_and1285_y0);
  and_gate and_gate_h_u_cla32_and1286_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1286_y0);
  and_gate and_gate_h_u_cla32_and1287_y0(h_u_cla32_and1286_y0, h_u_cla32_and1285_y0, h_u_cla32_and1287_y0);
  and_gate and_gate_h_u_cla32_and1288_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1288_y0);
  and_gate and_gate_h_u_cla32_and1289_y0(h_u_cla32_and1288_y0, h_u_cla32_and1287_y0, h_u_cla32_and1289_y0);
  and_gate and_gate_h_u_cla32_and1290_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1290_y0);
  and_gate and_gate_h_u_cla32_and1291_y0(h_u_cla32_and1290_y0, h_u_cla32_and1289_y0, h_u_cla32_and1291_y0);
  and_gate and_gate_h_u_cla32_and1292_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1292_y0);
  and_gate and_gate_h_u_cla32_and1293_y0(h_u_cla32_and1292_y0, h_u_cla32_and1291_y0, h_u_cla32_and1293_y0);
  and_gate and_gate_h_u_cla32_and1294_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1294_y0);
  and_gate and_gate_h_u_cla32_and1295_y0(h_u_cla32_and1294_y0, h_u_cla32_and1293_y0, h_u_cla32_and1295_y0);
  and_gate and_gate_h_u_cla32_and1296_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1296_y0);
  and_gate and_gate_h_u_cla32_and1297_y0(h_u_cla32_and1296_y0, h_u_cla32_and1295_y0, h_u_cla32_and1297_y0);
  and_gate and_gate_h_u_cla32_and1298_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1298_y0);
  and_gate and_gate_h_u_cla32_and1299_y0(h_u_cla32_and1298_y0, h_u_cla32_and1297_y0, h_u_cla32_and1299_y0);
  and_gate and_gate_h_u_cla32_and1300_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1300_y0);
  and_gate and_gate_h_u_cla32_and1301_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1301_y0);
  and_gate and_gate_h_u_cla32_and1302_y0(h_u_cla32_and1301_y0, h_u_cla32_and1300_y0, h_u_cla32_and1302_y0);
  and_gate and_gate_h_u_cla32_and1303_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1303_y0);
  and_gate and_gate_h_u_cla32_and1304_y0(h_u_cla32_and1303_y0, h_u_cla32_and1302_y0, h_u_cla32_and1304_y0);
  and_gate and_gate_h_u_cla32_and1305_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1305_y0);
  and_gate and_gate_h_u_cla32_and1306_y0(h_u_cla32_and1305_y0, h_u_cla32_and1304_y0, h_u_cla32_and1306_y0);
  and_gate and_gate_h_u_cla32_and1307_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1307_y0);
  and_gate and_gate_h_u_cla32_and1308_y0(h_u_cla32_and1307_y0, h_u_cla32_and1306_y0, h_u_cla32_and1308_y0);
  and_gate and_gate_h_u_cla32_and1309_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1309_y0);
  and_gate and_gate_h_u_cla32_and1310_y0(h_u_cla32_and1309_y0, h_u_cla32_and1308_y0, h_u_cla32_and1310_y0);
  and_gate and_gate_h_u_cla32_and1311_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1311_y0);
  and_gate and_gate_h_u_cla32_and1312_y0(h_u_cla32_and1311_y0, h_u_cla32_and1310_y0, h_u_cla32_and1312_y0);
  and_gate and_gate_h_u_cla32_and1313_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1313_y0);
  and_gate and_gate_h_u_cla32_and1314_y0(h_u_cla32_and1313_y0, h_u_cla32_and1312_y0, h_u_cla32_and1314_y0);
  and_gate and_gate_h_u_cla32_and1315_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1315_y0);
  and_gate and_gate_h_u_cla32_and1316_y0(h_u_cla32_and1315_y0, h_u_cla32_and1314_y0, h_u_cla32_and1316_y0);
  and_gate and_gate_h_u_cla32_and1317_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1317_y0);
  and_gate and_gate_h_u_cla32_and1318_y0(h_u_cla32_and1317_y0, h_u_cla32_and1316_y0, h_u_cla32_and1318_y0);
  and_gate and_gate_h_u_cla32_and1319_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1319_y0);
  and_gate and_gate_h_u_cla32_and1320_y0(h_u_cla32_and1319_y0, h_u_cla32_and1318_y0, h_u_cla32_and1320_y0);
  and_gate and_gate_h_u_cla32_and1321_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1321_y0);
  and_gate and_gate_h_u_cla32_and1322_y0(h_u_cla32_and1321_y0, h_u_cla32_and1320_y0, h_u_cla32_and1322_y0);
  and_gate and_gate_h_u_cla32_and1323_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1323_y0);
  and_gate and_gate_h_u_cla32_and1324_y0(h_u_cla32_and1323_y0, h_u_cla32_and1322_y0, h_u_cla32_and1324_y0);
  and_gate and_gate_h_u_cla32_and1325_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1325_y0);
  and_gate and_gate_h_u_cla32_and1326_y0(h_u_cla32_and1325_y0, h_u_cla32_and1324_y0, h_u_cla32_and1326_y0);
  and_gate and_gate_h_u_cla32_and1327_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1327_y0);
  and_gate and_gate_h_u_cla32_and1328_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1328_y0);
  and_gate and_gate_h_u_cla32_and1329_y0(h_u_cla32_and1328_y0, h_u_cla32_and1327_y0, h_u_cla32_and1329_y0);
  and_gate and_gate_h_u_cla32_and1330_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1330_y0);
  and_gate and_gate_h_u_cla32_and1331_y0(h_u_cla32_and1330_y0, h_u_cla32_and1329_y0, h_u_cla32_and1331_y0);
  and_gate and_gate_h_u_cla32_and1332_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1332_y0);
  and_gate and_gate_h_u_cla32_and1333_y0(h_u_cla32_and1332_y0, h_u_cla32_and1331_y0, h_u_cla32_and1333_y0);
  and_gate and_gate_h_u_cla32_and1334_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1334_y0);
  and_gate and_gate_h_u_cla32_and1335_y0(h_u_cla32_and1334_y0, h_u_cla32_and1333_y0, h_u_cla32_and1335_y0);
  and_gate and_gate_h_u_cla32_and1336_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1336_y0);
  and_gate and_gate_h_u_cla32_and1337_y0(h_u_cla32_and1336_y0, h_u_cla32_and1335_y0, h_u_cla32_and1337_y0);
  and_gate and_gate_h_u_cla32_and1338_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1338_y0);
  and_gate and_gate_h_u_cla32_and1339_y0(h_u_cla32_and1338_y0, h_u_cla32_and1337_y0, h_u_cla32_and1339_y0);
  and_gate and_gate_h_u_cla32_and1340_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1340_y0);
  and_gate and_gate_h_u_cla32_and1341_y0(h_u_cla32_and1340_y0, h_u_cla32_and1339_y0, h_u_cla32_and1341_y0);
  and_gate and_gate_h_u_cla32_and1342_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1342_y0);
  and_gate and_gate_h_u_cla32_and1343_y0(h_u_cla32_and1342_y0, h_u_cla32_and1341_y0, h_u_cla32_and1343_y0);
  and_gate and_gate_h_u_cla32_and1344_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1344_y0);
  and_gate and_gate_h_u_cla32_and1345_y0(h_u_cla32_and1344_y0, h_u_cla32_and1343_y0, h_u_cla32_and1345_y0);
  and_gate and_gate_h_u_cla32_and1346_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1346_y0);
  and_gate and_gate_h_u_cla32_and1347_y0(h_u_cla32_and1346_y0, h_u_cla32_and1345_y0, h_u_cla32_and1347_y0);
  and_gate and_gate_h_u_cla32_and1348_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1348_y0);
  and_gate and_gate_h_u_cla32_and1349_y0(h_u_cla32_and1348_y0, h_u_cla32_and1347_y0, h_u_cla32_and1349_y0);
  and_gate and_gate_h_u_cla32_and1350_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1350_y0);
  and_gate and_gate_h_u_cla32_and1351_y0(h_u_cla32_and1350_y0, h_u_cla32_and1349_y0, h_u_cla32_and1351_y0);
  and_gate and_gate_h_u_cla32_and1352_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1352_y0);
  and_gate and_gate_h_u_cla32_and1353_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1353_y0);
  and_gate and_gate_h_u_cla32_and1354_y0(h_u_cla32_and1353_y0, h_u_cla32_and1352_y0, h_u_cla32_and1354_y0);
  and_gate and_gate_h_u_cla32_and1355_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1355_y0);
  and_gate and_gate_h_u_cla32_and1356_y0(h_u_cla32_and1355_y0, h_u_cla32_and1354_y0, h_u_cla32_and1356_y0);
  and_gate and_gate_h_u_cla32_and1357_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1357_y0);
  and_gate and_gate_h_u_cla32_and1358_y0(h_u_cla32_and1357_y0, h_u_cla32_and1356_y0, h_u_cla32_and1358_y0);
  and_gate and_gate_h_u_cla32_and1359_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1359_y0);
  and_gate and_gate_h_u_cla32_and1360_y0(h_u_cla32_and1359_y0, h_u_cla32_and1358_y0, h_u_cla32_and1360_y0);
  and_gate and_gate_h_u_cla32_and1361_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1361_y0);
  and_gate and_gate_h_u_cla32_and1362_y0(h_u_cla32_and1361_y0, h_u_cla32_and1360_y0, h_u_cla32_and1362_y0);
  and_gate and_gate_h_u_cla32_and1363_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1363_y0);
  and_gate and_gate_h_u_cla32_and1364_y0(h_u_cla32_and1363_y0, h_u_cla32_and1362_y0, h_u_cla32_and1364_y0);
  and_gate and_gate_h_u_cla32_and1365_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1365_y0);
  and_gate and_gate_h_u_cla32_and1366_y0(h_u_cla32_and1365_y0, h_u_cla32_and1364_y0, h_u_cla32_and1366_y0);
  and_gate and_gate_h_u_cla32_and1367_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1367_y0);
  and_gate and_gate_h_u_cla32_and1368_y0(h_u_cla32_and1367_y0, h_u_cla32_and1366_y0, h_u_cla32_and1368_y0);
  and_gate and_gate_h_u_cla32_and1369_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1369_y0);
  and_gate and_gate_h_u_cla32_and1370_y0(h_u_cla32_and1369_y0, h_u_cla32_and1368_y0, h_u_cla32_and1370_y0);
  and_gate and_gate_h_u_cla32_and1371_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1371_y0);
  and_gate and_gate_h_u_cla32_and1372_y0(h_u_cla32_and1371_y0, h_u_cla32_and1370_y0, h_u_cla32_and1372_y0);
  and_gate and_gate_h_u_cla32_and1373_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1373_y0);
  and_gate and_gate_h_u_cla32_and1374_y0(h_u_cla32_and1373_y0, h_u_cla32_and1372_y0, h_u_cla32_and1374_y0);
  and_gate and_gate_h_u_cla32_and1375_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1375_y0);
  and_gate and_gate_h_u_cla32_and1376_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1376_y0);
  and_gate and_gate_h_u_cla32_and1377_y0(h_u_cla32_and1376_y0, h_u_cla32_and1375_y0, h_u_cla32_and1377_y0);
  and_gate and_gate_h_u_cla32_and1378_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1378_y0);
  and_gate and_gate_h_u_cla32_and1379_y0(h_u_cla32_and1378_y0, h_u_cla32_and1377_y0, h_u_cla32_and1379_y0);
  and_gate and_gate_h_u_cla32_and1380_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1380_y0);
  and_gate and_gate_h_u_cla32_and1381_y0(h_u_cla32_and1380_y0, h_u_cla32_and1379_y0, h_u_cla32_and1381_y0);
  and_gate and_gate_h_u_cla32_and1382_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1382_y0);
  and_gate and_gate_h_u_cla32_and1383_y0(h_u_cla32_and1382_y0, h_u_cla32_and1381_y0, h_u_cla32_and1383_y0);
  and_gate and_gate_h_u_cla32_and1384_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1384_y0);
  and_gate and_gate_h_u_cla32_and1385_y0(h_u_cla32_and1384_y0, h_u_cla32_and1383_y0, h_u_cla32_and1385_y0);
  and_gate and_gate_h_u_cla32_and1386_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1386_y0);
  and_gate and_gate_h_u_cla32_and1387_y0(h_u_cla32_and1386_y0, h_u_cla32_and1385_y0, h_u_cla32_and1387_y0);
  and_gate and_gate_h_u_cla32_and1388_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1388_y0);
  and_gate and_gate_h_u_cla32_and1389_y0(h_u_cla32_and1388_y0, h_u_cla32_and1387_y0, h_u_cla32_and1389_y0);
  and_gate and_gate_h_u_cla32_and1390_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1390_y0);
  and_gate and_gate_h_u_cla32_and1391_y0(h_u_cla32_and1390_y0, h_u_cla32_and1389_y0, h_u_cla32_and1391_y0);
  and_gate and_gate_h_u_cla32_and1392_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1392_y0);
  and_gate and_gate_h_u_cla32_and1393_y0(h_u_cla32_and1392_y0, h_u_cla32_and1391_y0, h_u_cla32_and1393_y0);
  and_gate and_gate_h_u_cla32_and1394_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1394_y0);
  and_gate and_gate_h_u_cla32_and1395_y0(h_u_cla32_and1394_y0, h_u_cla32_and1393_y0, h_u_cla32_and1395_y0);
  and_gate and_gate_h_u_cla32_and1396_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1396_y0);
  and_gate and_gate_h_u_cla32_and1397_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1397_y0);
  and_gate and_gate_h_u_cla32_and1398_y0(h_u_cla32_and1397_y0, h_u_cla32_and1396_y0, h_u_cla32_and1398_y0);
  and_gate and_gate_h_u_cla32_and1399_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1399_y0);
  and_gate and_gate_h_u_cla32_and1400_y0(h_u_cla32_and1399_y0, h_u_cla32_and1398_y0, h_u_cla32_and1400_y0);
  and_gate and_gate_h_u_cla32_and1401_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1401_y0);
  and_gate and_gate_h_u_cla32_and1402_y0(h_u_cla32_and1401_y0, h_u_cla32_and1400_y0, h_u_cla32_and1402_y0);
  and_gate and_gate_h_u_cla32_and1403_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1403_y0);
  and_gate and_gate_h_u_cla32_and1404_y0(h_u_cla32_and1403_y0, h_u_cla32_and1402_y0, h_u_cla32_and1404_y0);
  and_gate and_gate_h_u_cla32_and1405_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1405_y0);
  and_gate and_gate_h_u_cla32_and1406_y0(h_u_cla32_and1405_y0, h_u_cla32_and1404_y0, h_u_cla32_and1406_y0);
  and_gate and_gate_h_u_cla32_and1407_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1407_y0);
  and_gate and_gate_h_u_cla32_and1408_y0(h_u_cla32_and1407_y0, h_u_cla32_and1406_y0, h_u_cla32_and1408_y0);
  and_gate and_gate_h_u_cla32_and1409_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1409_y0);
  and_gate and_gate_h_u_cla32_and1410_y0(h_u_cla32_and1409_y0, h_u_cla32_and1408_y0, h_u_cla32_and1410_y0);
  and_gate and_gate_h_u_cla32_and1411_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1411_y0);
  and_gate and_gate_h_u_cla32_and1412_y0(h_u_cla32_and1411_y0, h_u_cla32_and1410_y0, h_u_cla32_and1412_y0);
  and_gate and_gate_h_u_cla32_and1413_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1413_y0);
  and_gate and_gate_h_u_cla32_and1414_y0(h_u_cla32_and1413_y0, h_u_cla32_and1412_y0, h_u_cla32_and1414_y0);
  and_gate and_gate_h_u_cla32_and1415_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1415_y0);
  and_gate and_gate_h_u_cla32_and1416_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1416_y0);
  and_gate and_gate_h_u_cla32_and1417_y0(h_u_cla32_and1416_y0, h_u_cla32_and1415_y0, h_u_cla32_and1417_y0);
  and_gate and_gate_h_u_cla32_and1418_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1418_y0);
  and_gate and_gate_h_u_cla32_and1419_y0(h_u_cla32_and1418_y0, h_u_cla32_and1417_y0, h_u_cla32_and1419_y0);
  and_gate and_gate_h_u_cla32_and1420_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1420_y0);
  and_gate and_gate_h_u_cla32_and1421_y0(h_u_cla32_and1420_y0, h_u_cla32_and1419_y0, h_u_cla32_and1421_y0);
  and_gate and_gate_h_u_cla32_and1422_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1422_y0);
  and_gate and_gate_h_u_cla32_and1423_y0(h_u_cla32_and1422_y0, h_u_cla32_and1421_y0, h_u_cla32_and1423_y0);
  and_gate and_gate_h_u_cla32_and1424_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1424_y0);
  and_gate and_gate_h_u_cla32_and1425_y0(h_u_cla32_and1424_y0, h_u_cla32_and1423_y0, h_u_cla32_and1425_y0);
  and_gate and_gate_h_u_cla32_and1426_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1426_y0);
  and_gate and_gate_h_u_cla32_and1427_y0(h_u_cla32_and1426_y0, h_u_cla32_and1425_y0, h_u_cla32_and1427_y0);
  and_gate and_gate_h_u_cla32_and1428_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1428_y0);
  and_gate and_gate_h_u_cla32_and1429_y0(h_u_cla32_and1428_y0, h_u_cla32_and1427_y0, h_u_cla32_and1429_y0);
  and_gate and_gate_h_u_cla32_and1430_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1430_y0);
  and_gate and_gate_h_u_cla32_and1431_y0(h_u_cla32_and1430_y0, h_u_cla32_and1429_y0, h_u_cla32_and1431_y0);
  and_gate and_gate_h_u_cla32_and1432_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1432_y0);
  and_gate and_gate_h_u_cla32_and1433_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1433_y0);
  and_gate and_gate_h_u_cla32_and1434_y0(h_u_cla32_and1433_y0, h_u_cla32_and1432_y0, h_u_cla32_and1434_y0);
  and_gate and_gate_h_u_cla32_and1435_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1435_y0);
  and_gate and_gate_h_u_cla32_and1436_y0(h_u_cla32_and1435_y0, h_u_cla32_and1434_y0, h_u_cla32_and1436_y0);
  and_gate and_gate_h_u_cla32_and1437_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1437_y0);
  and_gate and_gate_h_u_cla32_and1438_y0(h_u_cla32_and1437_y0, h_u_cla32_and1436_y0, h_u_cla32_and1438_y0);
  and_gate and_gate_h_u_cla32_and1439_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1439_y0);
  and_gate and_gate_h_u_cla32_and1440_y0(h_u_cla32_and1439_y0, h_u_cla32_and1438_y0, h_u_cla32_and1440_y0);
  and_gate and_gate_h_u_cla32_and1441_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1441_y0);
  and_gate and_gate_h_u_cla32_and1442_y0(h_u_cla32_and1441_y0, h_u_cla32_and1440_y0, h_u_cla32_and1442_y0);
  and_gate and_gate_h_u_cla32_and1443_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1443_y0);
  and_gate and_gate_h_u_cla32_and1444_y0(h_u_cla32_and1443_y0, h_u_cla32_and1442_y0, h_u_cla32_and1444_y0);
  and_gate and_gate_h_u_cla32_and1445_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1445_y0);
  and_gate and_gate_h_u_cla32_and1446_y0(h_u_cla32_and1445_y0, h_u_cla32_and1444_y0, h_u_cla32_and1446_y0);
  and_gate and_gate_h_u_cla32_and1447_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1447_y0);
  and_gate and_gate_h_u_cla32_and1448_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1448_y0);
  and_gate and_gate_h_u_cla32_and1449_y0(h_u_cla32_and1448_y0, h_u_cla32_and1447_y0, h_u_cla32_and1449_y0);
  and_gate and_gate_h_u_cla32_and1450_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1450_y0);
  and_gate and_gate_h_u_cla32_and1451_y0(h_u_cla32_and1450_y0, h_u_cla32_and1449_y0, h_u_cla32_and1451_y0);
  and_gate and_gate_h_u_cla32_and1452_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1452_y0);
  and_gate and_gate_h_u_cla32_and1453_y0(h_u_cla32_and1452_y0, h_u_cla32_and1451_y0, h_u_cla32_and1453_y0);
  and_gate and_gate_h_u_cla32_and1454_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1454_y0);
  and_gate and_gate_h_u_cla32_and1455_y0(h_u_cla32_and1454_y0, h_u_cla32_and1453_y0, h_u_cla32_and1455_y0);
  and_gate and_gate_h_u_cla32_and1456_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1456_y0);
  and_gate and_gate_h_u_cla32_and1457_y0(h_u_cla32_and1456_y0, h_u_cla32_and1455_y0, h_u_cla32_and1457_y0);
  and_gate and_gate_h_u_cla32_and1458_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1458_y0);
  and_gate and_gate_h_u_cla32_and1459_y0(h_u_cla32_and1458_y0, h_u_cla32_and1457_y0, h_u_cla32_and1459_y0);
  and_gate and_gate_h_u_cla32_and1460_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1460_y0);
  and_gate and_gate_h_u_cla32_and1461_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1461_y0);
  and_gate and_gate_h_u_cla32_and1462_y0(h_u_cla32_and1461_y0, h_u_cla32_and1460_y0, h_u_cla32_and1462_y0);
  and_gate and_gate_h_u_cla32_and1463_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1463_y0);
  and_gate and_gate_h_u_cla32_and1464_y0(h_u_cla32_and1463_y0, h_u_cla32_and1462_y0, h_u_cla32_and1464_y0);
  and_gate and_gate_h_u_cla32_and1465_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1465_y0);
  and_gate and_gate_h_u_cla32_and1466_y0(h_u_cla32_and1465_y0, h_u_cla32_and1464_y0, h_u_cla32_and1466_y0);
  and_gate and_gate_h_u_cla32_and1467_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1467_y0);
  and_gate and_gate_h_u_cla32_and1468_y0(h_u_cla32_and1467_y0, h_u_cla32_and1466_y0, h_u_cla32_and1468_y0);
  and_gate and_gate_h_u_cla32_and1469_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1469_y0);
  and_gate and_gate_h_u_cla32_and1470_y0(h_u_cla32_and1469_y0, h_u_cla32_and1468_y0, h_u_cla32_and1470_y0);
  and_gate and_gate_h_u_cla32_and1471_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1471_y0);
  and_gate and_gate_h_u_cla32_and1472_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1472_y0);
  and_gate and_gate_h_u_cla32_and1473_y0(h_u_cla32_and1472_y0, h_u_cla32_and1471_y0, h_u_cla32_and1473_y0);
  and_gate and_gate_h_u_cla32_and1474_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1474_y0);
  and_gate and_gate_h_u_cla32_and1475_y0(h_u_cla32_and1474_y0, h_u_cla32_and1473_y0, h_u_cla32_and1475_y0);
  and_gate and_gate_h_u_cla32_and1476_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1476_y0);
  and_gate and_gate_h_u_cla32_and1477_y0(h_u_cla32_and1476_y0, h_u_cla32_and1475_y0, h_u_cla32_and1477_y0);
  and_gate and_gate_h_u_cla32_and1478_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1478_y0);
  and_gate and_gate_h_u_cla32_and1479_y0(h_u_cla32_and1478_y0, h_u_cla32_and1477_y0, h_u_cla32_and1479_y0);
  and_gate and_gate_h_u_cla32_and1480_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1480_y0);
  and_gate and_gate_h_u_cla32_and1481_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1481_y0);
  and_gate and_gate_h_u_cla32_and1482_y0(h_u_cla32_and1481_y0, h_u_cla32_and1480_y0, h_u_cla32_and1482_y0);
  and_gate and_gate_h_u_cla32_and1483_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1483_y0);
  and_gate and_gate_h_u_cla32_and1484_y0(h_u_cla32_and1483_y0, h_u_cla32_and1482_y0, h_u_cla32_and1484_y0);
  and_gate and_gate_h_u_cla32_and1485_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1485_y0);
  and_gate and_gate_h_u_cla32_and1486_y0(h_u_cla32_and1485_y0, h_u_cla32_and1484_y0, h_u_cla32_and1486_y0);
  and_gate and_gate_h_u_cla32_and1487_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1487_y0);
  and_gate and_gate_h_u_cla32_and1488_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1488_y0);
  and_gate and_gate_h_u_cla32_and1489_y0(h_u_cla32_and1488_y0, h_u_cla32_and1487_y0, h_u_cla32_and1489_y0);
  and_gate and_gate_h_u_cla32_and1490_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1490_y0);
  and_gate and_gate_h_u_cla32_and1491_y0(h_u_cla32_and1490_y0, h_u_cla32_and1489_y0, h_u_cla32_and1491_y0);
  and_gate and_gate_h_u_cla32_and1492_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and1492_y0);
  and_gate and_gate_h_u_cla32_and1493_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and1493_y0);
  and_gate and_gate_h_u_cla32_and1494_y0(h_u_cla32_and1493_y0, h_u_cla32_and1492_y0, h_u_cla32_and1494_y0);
  and_gate and_gate_h_u_cla32_and1495_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and1495_y0);
  or_gate or_gate_h_u_cla32_or120_y0(h_u_cla32_and1495_y0, h_u_cla32_and1270_y0, h_u_cla32_or120_y0);
  or_gate or_gate_h_u_cla32_or121_y0(h_u_cla32_or120_y0, h_u_cla32_and1299_y0, h_u_cla32_or121_y0);
  or_gate or_gate_h_u_cla32_or122_y0(h_u_cla32_or121_y0, h_u_cla32_and1326_y0, h_u_cla32_or122_y0);
  or_gate or_gate_h_u_cla32_or123_y0(h_u_cla32_or122_y0, h_u_cla32_and1351_y0, h_u_cla32_or123_y0);
  or_gate or_gate_h_u_cla32_or124_y0(h_u_cla32_or123_y0, h_u_cla32_and1374_y0, h_u_cla32_or124_y0);
  or_gate or_gate_h_u_cla32_or125_y0(h_u_cla32_or124_y0, h_u_cla32_and1395_y0, h_u_cla32_or125_y0);
  or_gate or_gate_h_u_cla32_or126_y0(h_u_cla32_or125_y0, h_u_cla32_and1414_y0, h_u_cla32_or126_y0);
  or_gate or_gate_h_u_cla32_or127_y0(h_u_cla32_or126_y0, h_u_cla32_and1431_y0, h_u_cla32_or127_y0);
  or_gate or_gate_h_u_cla32_or128_y0(h_u_cla32_or127_y0, h_u_cla32_and1446_y0, h_u_cla32_or128_y0);
  or_gate or_gate_h_u_cla32_or129_y0(h_u_cla32_or128_y0, h_u_cla32_and1459_y0, h_u_cla32_or129_y0);
  or_gate or_gate_h_u_cla32_or130_y0(h_u_cla32_or129_y0, h_u_cla32_and1470_y0, h_u_cla32_or130_y0);
  or_gate or_gate_h_u_cla32_or131_y0(h_u_cla32_or130_y0, h_u_cla32_and1479_y0, h_u_cla32_or131_y0);
  or_gate or_gate_h_u_cla32_or132_y0(h_u_cla32_or131_y0, h_u_cla32_and1486_y0, h_u_cla32_or132_y0);
  or_gate or_gate_h_u_cla32_or133_y0(h_u_cla32_or132_y0, h_u_cla32_and1491_y0, h_u_cla32_or133_y0);
  or_gate or_gate_h_u_cla32_or134_y0(h_u_cla32_or133_y0, h_u_cla32_and1494_y0, h_u_cla32_or134_y0);
  or_gate or_gate_h_u_cla32_or135_y0(h_u_cla32_pg_logic15_y1, h_u_cla32_or134_y0, h_u_cla32_or135_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic16_y0(a_16, b_16, h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_pg_logic16_y2);
  xor_gate xor_gate_h_u_cla32_xor16_y0(h_u_cla32_pg_logic16_y2, h_u_cla32_or135_y0, h_u_cla32_xor16_y0);
  and_gate and_gate_h_u_cla32_and1496_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and1496_y0);
  and_gate and_gate_h_u_cla32_and1497_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and1497_y0);
  and_gate and_gate_h_u_cla32_and1498_y0(h_u_cla32_and1497_y0, h_u_cla32_and1496_y0, h_u_cla32_and1498_y0);
  and_gate and_gate_h_u_cla32_and1499_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and1499_y0);
  and_gate and_gate_h_u_cla32_and1500_y0(h_u_cla32_and1499_y0, h_u_cla32_and1498_y0, h_u_cla32_and1500_y0);
  and_gate and_gate_h_u_cla32_and1501_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and1501_y0);
  and_gate and_gate_h_u_cla32_and1502_y0(h_u_cla32_and1501_y0, h_u_cla32_and1500_y0, h_u_cla32_and1502_y0);
  and_gate and_gate_h_u_cla32_and1503_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and1503_y0);
  and_gate and_gate_h_u_cla32_and1504_y0(h_u_cla32_and1503_y0, h_u_cla32_and1502_y0, h_u_cla32_and1504_y0);
  and_gate and_gate_h_u_cla32_and1505_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and1505_y0);
  and_gate and_gate_h_u_cla32_and1506_y0(h_u_cla32_and1505_y0, h_u_cla32_and1504_y0, h_u_cla32_and1506_y0);
  and_gate and_gate_h_u_cla32_and1507_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and1507_y0);
  and_gate and_gate_h_u_cla32_and1508_y0(h_u_cla32_and1507_y0, h_u_cla32_and1506_y0, h_u_cla32_and1508_y0);
  and_gate and_gate_h_u_cla32_and1509_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and1509_y0);
  and_gate and_gate_h_u_cla32_and1510_y0(h_u_cla32_and1509_y0, h_u_cla32_and1508_y0, h_u_cla32_and1510_y0);
  and_gate and_gate_h_u_cla32_and1511_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and1511_y0);
  and_gate and_gate_h_u_cla32_and1512_y0(h_u_cla32_and1511_y0, h_u_cla32_and1510_y0, h_u_cla32_and1512_y0);
  and_gate and_gate_h_u_cla32_and1513_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and1513_y0);
  and_gate and_gate_h_u_cla32_and1514_y0(h_u_cla32_and1513_y0, h_u_cla32_and1512_y0, h_u_cla32_and1514_y0);
  and_gate and_gate_h_u_cla32_and1515_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and1515_y0);
  and_gate and_gate_h_u_cla32_and1516_y0(h_u_cla32_and1515_y0, h_u_cla32_and1514_y0, h_u_cla32_and1516_y0);
  and_gate and_gate_h_u_cla32_and1517_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and1517_y0);
  and_gate and_gate_h_u_cla32_and1518_y0(h_u_cla32_and1517_y0, h_u_cla32_and1516_y0, h_u_cla32_and1518_y0);
  and_gate and_gate_h_u_cla32_and1519_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and1519_y0);
  and_gate and_gate_h_u_cla32_and1520_y0(h_u_cla32_and1519_y0, h_u_cla32_and1518_y0, h_u_cla32_and1520_y0);
  and_gate and_gate_h_u_cla32_and1521_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and1521_y0);
  and_gate and_gate_h_u_cla32_and1522_y0(h_u_cla32_and1521_y0, h_u_cla32_and1520_y0, h_u_cla32_and1522_y0);
  and_gate and_gate_h_u_cla32_and1523_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and1523_y0);
  and_gate and_gate_h_u_cla32_and1524_y0(h_u_cla32_and1523_y0, h_u_cla32_and1522_y0, h_u_cla32_and1524_y0);
  and_gate and_gate_h_u_cla32_and1525_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and1525_y0);
  and_gate and_gate_h_u_cla32_and1526_y0(h_u_cla32_and1525_y0, h_u_cla32_and1524_y0, h_u_cla32_and1526_y0);
  and_gate and_gate_h_u_cla32_and1527_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and1527_y0);
  and_gate and_gate_h_u_cla32_and1528_y0(h_u_cla32_and1527_y0, h_u_cla32_and1526_y0, h_u_cla32_and1528_y0);
  and_gate and_gate_h_u_cla32_and1529_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1529_y0);
  and_gate and_gate_h_u_cla32_and1530_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1530_y0);
  and_gate and_gate_h_u_cla32_and1531_y0(h_u_cla32_and1530_y0, h_u_cla32_and1529_y0, h_u_cla32_and1531_y0);
  and_gate and_gate_h_u_cla32_and1532_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1532_y0);
  and_gate and_gate_h_u_cla32_and1533_y0(h_u_cla32_and1532_y0, h_u_cla32_and1531_y0, h_u_cla32_and1533_y0);
  and_gate and_gate_h_u_cla32_and1534_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1534_y0);
  and_gate and_gate_h_u_cla32_and1535_y0(h_u_cla32_and1534_y0, h_u_cla32_and1533_y0, h_u_cla32_and1535_y0);
  and_gate and_gate_h_u_cla32_and1536_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1536_y0);
  and_gate and_gate_h_u_cla32_and1537_y0(h_u_cla32_and1536_y0, h_u_cla32_and1535_y0, h_u_cla32_and1537_y0);
  and_gate and_gate_h_u_cla32_and1538_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1538_y0);
  and_gate and_gate_h_u_cla32_and1539_y0(h_u_cla32_and1538_y0, h_u_cla32_and1537_y0, h_u_cla32_and1539_y0);
  and_gate and_gate_h_u_cla32_and1540_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1540_y0);
  and_gate and_gate_h_u_cla32_and1541_y0(h_u_cla32_and1540_y0, h_u_cla32_and1539_y0, h_u_cla32_and1541_y0);
  and_gate and_gate_h_u_cla32_and1542_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1542_y0);
  and_gate and_gate_h_u_cla32_and1543_y0(h_u_cla32_and1542_y0, h_u_cla32_and1541_y0, h_u_cla32_and1543_y0);
  and_gate and_gate_h_u_cla32_and1544_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1544_y0);
  and_gate and_gate_h_u_cla32_and1545_y0(h_u_cla32_and1544_y0, h_u_cla32_and1543_y0, h_u_cla32_and1545_y0);
  and_gate and_gate_h_u_cla32_and1546_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1546_y0);
  and_gate and_gate_h_u_cla32_and1547_y0(h_u_cla32_and1546_y0, h_u_cla32_and1545_y0, h_u_cla32_and1547_y0);
  and_gate and_gate_h_u_cla32_and1548_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1548_y0);
  and_gate and_gate_h_u_cla32_and1549_y0(h_u_cla32_and1548_y0, h_u_cla32_and1547_y0, h_u_cla32_and1549_y0);
  and_gate and_gate_h_u_cla32_and1550_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1550_y0);
  and_gate and_gate_h_u_cla32_and1551_y0(h_u_cla32_and1550_y0, h_u_cla32_and1549_y0, h_u_cla32_and1551_y0);
  and_gate and_gate_h_u_cla32_and1552_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1552_y0);
  and_gate and_gate_h_u_cla32_and1553_y0(h_u_cla32_and1552_y0, h_u_cla32_and1551_y0, h_u_cla32_and1553_y0);
  and_gate and_gate_h_u_cla32_and1554_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1554_y0);
  and_gate and_gate_h_u_cla32_and1555_y0(h_u_cla32_and1554_y0, h_u_cla32_and1553_y0, h_u_cla32_and1555_y0);
  and_gate and_gate_h_u_cla32_and1556_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1556_y0);
  and_gate and_gate_h_u_cla32_and1557_y0(h_u_cla32_and1556_y0, h_u_cla32_and1555_y0, h_u_cla32_and1557_y0);
  and_gate and_gate_h_u_cla32_and1558_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1558_y0);
  and_gate and_gate_h_u_cla32_and1559_y0(h_u_cla32_and1558_y0, h_u_cla32_and1557_y0, h_u_cla32_and1559_y0);
  and_gate and_gate_h_u_cla32_and1560_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1560_y0);
  and_gate and_gate_h_u_cla32_and1561_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1561_y0);
  and_gate and_gate_h_u_cla32_and1562_y0(h_u_cla32_and1561_y0, h_u_cla32_and1560_y0, h_u_cla32_and1562_y0);
  and_gate and_gate_h_u_cla32_and1563_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1563_y0);
  and_gate and_gate_h_u_cla32_and1564_y0(h_u_cla32_and1563_y0, h_u_cla32_and1562_y0, h_u_cla32_and1564_y0);
  and_gate and_gate_h_u_cla32_and1565_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1565_y0);
  and_gate and_gate_h_u_cla32_and1566_y0(h_u_cla32_and1565_y0, h_u_cla32_and1564_y0, h_u_cla32_and1566_y0);
  and_gate and_gate_h_u_cla32_and1567_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1567_y0);
  and_gate and_gate_h_u_cla32_and1568_y0(h_u_cla32_and1567_y0, h_u_cla32_and1566_y0, h_u_cla32_and1568_y0);
  and_gate and_gate_h_u_cla32_and1569_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1569_y0);
  and_gate and_gate_h_u_cla32_and1570_y0(h_u_cla32_and1569_y0, h_u_cla32_and1568_y0, h_u_cla32_and1570_y0);
  and_gate and_gate_h_u_cla32_and1571_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1571_y0);
  and_gate and_gate_h_u_cla32_and1572_y0(h_u_cla32_and1571_y0, h_u_cla32_and1570_y0, h_u_cla32_and1572_y0);
  and_gate and_gate_h_u_cla32_and1573_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1573_y0);
  and_gate and_gate_h_u_cla32_and1574_y0(h_u_cla32_and1573_y0, h_u_cla32_and1572_y0, h_u_cla32_and1574_y0);
  and_gate and_gate_h_u_cla32_and1575_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1575_y0);
  and_gate and_gate_h_u_cla32_and1576_y0(h_u_cla32_and1575_y0, h_u_cla32_and1574_y0, h_u_cla32_and1576_y0);
  and_gate and_gate_h_u_cla32_and1577_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1577_y0);
  and_gate and_gate_h_u_cla32_and1578_y0(h_u_cla32_and1577_y0, h_u_cla32_and1576_y0, h_u_cla32_and1578_y0);
  and_gate and_gate_h_u_cla32_and1579_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1579_y0);
  and_gate and_gate_h_u_cla32_and1580_y0(h_u_cla32_and1579_y0, h_u_cla32_and1578_y0, h_u_cla32_and1580_y0);
  and_gate and_gate_h_u_cla32_and1581_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1581_y0);
  and_gate and_gate_h_u_cla32_and1582_y0(h_u_cla32_and1581_y0, h_u_cla32_and1580_y0, h_u_cla32_and1582_y0);
  and_gate and_gate_h_u_cla32_and1583_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1583_y0);
  and_gate and_gate_h_u_cla32_and1584_y0(h_u_cla32_and1583_y0, h_u_cla32_and1582_y0, h_u_cla32_and1584_y0);
  and_gate and_gate_h_u_cla32_and1585_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1585_y0);
  and_gate and_gate_h_u_cla32_and1586_y0(h_u_cla32_and1585_y0, h_u_cla32_and1584_y0, h_u_cla32_and1586_y0);
  and_gate and_gate_h_u_cla32_and1587_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1587_y0);
  and_gate and_gate_h_u_cla32_and1588_y0(h_u_cla32_and1587_y0, h_u_cla32_and1586_y0, h_u_cla32_and1588_y0);
  and_gate and_gate_h_u_cla32_and1589_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1589_y0);
  and_gate and_gate_h_u_cla32_and1590_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1590_y0);
  and_gate and_gate_h_u_cla32_and1591_y0(h_u_cla32_and1590_y0, h_u_cla32_and1589_y0, h_u_cla32_and1591_y0);
  and_gate and_gate_h_u_cla32_and1592_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1592_y0);
  and_gate and_gate_h_u_cla32_and1593_y0(h_u_cla32_and1592_y0, h_u_cla32_and1591_y0, h_u_cla32_and1593_y0);
  and_gate and_gate_h_u_cla32_and1594_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1594_y0);
  and_gate and_gate_h_u_cla32_and1595_y0(h_u_cla32_and1594_y0, h_u_cla32_and1593_y0, h_u_cla32_and1595_y0);
  and_gate and_gate_h_u_cla32_and1596_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1596_y0);
  and_gate and_gate_h_u_cla32_and1597_y0(h_u_cla32_and1596_y0, h_u_cla32_and1595_y0, h_u_cla32_and1597_y0);
  and_gate and_gate_h_u_cla32_and1598_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1598_y0);
  and_gate and_gate_h_u_cla32_and1599_y0(h_u_cla32_and1598_y0, h_u_cla32_and1597_y0, h_u_cla32_and1599_y0);
  and_gate and_gate_h_u_cla32_and1600_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1600_y0);
  and_gate and_gate_h_u_cla32_and1601_y0(h_u_cla32_and1600_y0, h_u_cla32_and1599_y0, h_u_cla32_and1601_y0);
  and_gate and_gate_h_u_cla32_and1602_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1602_y0);
  and_gate and_gate_h_u_cla32_and1603_y0(h_u_cla32_and1602_y0, h_u_cla32_and1601_y0, h_u_cla32_and1603_y0);
  and_gate and_gate_h_u_cla32_and1604_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1604_y0);
  and_gate and_gate_h_u_cla32_and1605_y0(h_u_cla32_and1604_y0, h_u_cla32_and1603_y0, h_u_cla32_and1605_y0);
  and_gate and_gate_h_u_cla32_and1606_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1606_y0);
  and_gate and_gate_h_u_cla32_and1607_y0(h_u_cla32_and1606_y0, h_u_cla32_and1605_y0, h_u_cla32_and1607_y0);
  and_gate and_gate_h_u_cla32_and1608_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1608_y0);
  and_gate and_gate_h_u_cla32_and1609_y0(h_u_cla32_and1608_y0, h_u_cla32_and1607_y0, h_u_cla32_and1609_y0);
  and_gate and_gate_h_u_cla32_and1610_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1610_y0);
  and_gate and_gate_h_u_cla32_and1611_y0(h_u_cla32_and1610_y0, h_u_cla32_and1609_y0, h_u_cla32_and1611_y0);
  and_gate and_gate_h_u_cla32_and1612_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1612_y0);
  and_gate and_gate_h_u_cla32_and1613_y0(h_u_cla32_and1612_y0, h_u_cla32_and1611_y0, h_u_cla32_and1613_y0);
  and_gate and_gate_h_u_cla32_and1614_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1614_y0);
  and_gate and_gate_h_u_cla32_and1615_y0(h_u_cla32_and1614_y0, h_u_cla32_and1613_y0, h_u_cla32_and1615_y0);
  and_gate and_gate_h_u_cla32_and1616_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1616_y0);
  and_gate and_gate_h_u_cla32_and1617_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1617_y0);
  and_gate and_gate_h_u_cla32_and1618_y0(h_u_cla32_and1617_y0, h_u_cla32_and1616_y0, h_u_cla32_and1618_y0);
  and_gate and_gate_h_u_cla32_and1619_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1619_y0);
  and_gate and_gate_h_u_cla32_and1620_y0(h_u_cla32_and1619_y0, h_u_cla32_and1618_y0, h_u_cla32_and1620_y0);
  and_gate and_gate_h_u_cla32_and1621_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1621_y0);
  and_gate and_gate_h_u_cla32_and1622_y0(h_u_cla32_and1621_y0, h_u_cla32_and1620_y0, h_u_cla32_and1622_y0);
  and_gate and_gate_h_u_cla32_and1623_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1623_y0);
  and_gate and_gate_h_u_cla32_and1624_y0(h_u_cla32_and1623_y0, h_u_cla32_and1622_y0, h_u_cla32_and1624_y0);
  and_gate and_gate_h_u_cla32_and1625_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1625_y0);
  and_gate and_gate_h_u_cla32_and1626_y0(h_u_cla32_and1625_y0, h_u_cla32_and1624_y0, h_u_cla32_and1626_y0);
  and_gate and_gate_h_u_cla32_and1627_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1627_y0);
  and_gate and_gate_h_u_cla32_and1628_y0(h_u_cla32_and1627_y0, h_u_cla32_and1626_y0, h_u_cla32_and1628_y0);
  and_gate and_gate_h_u_cla32_and1629_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1629_y0);
  and_gate and_gate_h_u_cla32_and1630_y0(h_u_cla32_and1629_y0, h_u_cla32_and1628_y0, h_u_cla32_and1630_y0);
  and_gate and_gate_h_u_cla32_and1631_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1631_y0);
  and_gate and_gate_h_u_cla32_and1632_y0(h_u_cla32_and1631_y0, h_u_cla32_and1630_y0, h_u_cla32_and1632_y0);
  and_gate and_gate_h_u_cla32_and1633_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1633_y0);
  and_gate and_gate_h_u_cla32_and1634_y0(h_u_cla32_and1633_y0, h_u_cla32_and1632_y0, h_u_cla32_and1634_y0);
  and_gate and_gate_h_u_cla32_and1635_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1635_y0);
  and_gate and_gate_h_u_cla32_and1636_y0(h_u_cla32_and1635_y0, h_u_cla32_and1634_y0, h_u_cla32_and1636_y0);
  and_gate and_gate_h_u_cla32_and1637_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1637_y0);
  and_gate and_gate_h_u_cla32_and1638_y0(h_u_cla32_and1637_y0, h_u_cla32_and1636_y0, h_u_cla32_and1638_y0);
  and_gate and_gate_h_u_cla32_and1639_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1639_y0);
  and_gate and_gate_h_u_cla32_and1640_y0(h_u_cla32_and1639_y0, h_u_cla32_and1638_y0, h_u_cla32_and1640_y0);
  and_gate and_gate_h_u_cla32_and1641_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1641_y0);
  and_gate and_gate_h_u_cla32_and1642_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1642_y0);
  and_gate and_gate_h_u_cla32_and1643_y0(h_u_cla32_and1642_y0, h_u_cla32_and1641_y0, h_u_cla32_and1643_y0);
  and_gate and_gate_h_u_cla32_and1644_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1644_y0);
  and_gate and_gate_h_u_cla32_and1645_y0(h_u_cla32_and1644_y0, h_u_cla32_and1643_y0, h_u_cla32_and1645_y0);
  and_gate and_gate_h_u_cla32_and1646_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1646_y0);
  and_gate and_gate_h_u_cla32_and1647_y0(h_u_cla32_and1646_y0, h_u_cla32_and1645_y0, h_u_cla32_and1647_y0);
  and_gate and_gate_h_u_cla32_and1648_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1648_y0);
  and_gate and_gate_h_u_cla32_and1649_y0(h_u_cla32_and1648_y0, h_u_cla32_and1647_y0, h_u_cla32_and1649_y0);
  and_gate and_gate_h_u_cla32_and1650_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1650_y0);
  and_gate and_gate_h_u_cla32_and1651_y0(h_u_cla32_and1650_y0, h_u_cla32_and1649_y0, h_u_cla32_and1651_y0);
  and_gate and_gate_h_u_cla32_and1652_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1652_y0);
  and_gate and_gate_h_u_cla32_and1653_y0(h_u_cla32_and1652_y0, h_u_cla32_and1651_y0, h_u_cla32_and1653_y0);
  and_gate and_gate_h_u_cla32_and1654_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1654_y0);
  and_gate and_gate_h_u_cla32_and1655_y0(h_u_cla32_and1654_y0, h_u_cla32_and1653_y0, h_u_cla32_and1655_y0);
  and_gate and_gate_h_u_cla32_and1656_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1656_y0);
  and_gate and_gate_h_u_cla32_and1657_y0(h_u_cla32_and1656_y0, h_u_cla32_and1655_y0, h_u_cla32_and1657_y0);
  and_gate and_gate_h_u_cla32_and1658_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1658_y0);
  and_gate and_gate_h_u_cla32_and1659_y0(h_u_cla32_and1658_y0, h_u_cla32_and1657_y0, h_u_cla32_and1659_y0);
  and_gate and_gate_h_u_cla32_and1660_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1660_y0);
  and_gate and_gate_h_u_cla32_and1661_y0(h_u_cla32_and1660_y0, h_u_cla32_and1659_y0, h_u_cla32_and1661_y0);
  and_gate and_gate_h_u_cla32_and1662_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1662_y0);
  and_gate and_gate_h_u_cla32_and1663_y0(h_u_cla32_and1662_y0, h_u_cla32_and1661_y0, h_u_cla32_and1663_y0);
  and_gate and_gate_h_u_cla32_and1664_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1664_y0);
  and_gate and_gate_h_u_cla32_and1665_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1665_y0);
  and_gate and_gate_h_u_cla32_and1666_y0(h_u_cla32_and1665_y0, h_u_cla32_and1664_y0, h_u_cla32_and1666_y0);
  and_gate and_gate_h_u_cla32_and1667_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1667_y0);
  and_gate and_gate_h_u_cla32_and1668_y0(h_u_cla32_and1667_y0, h_u_cla32_and1666_y0, h_u_cla32_and1668_y0);
  and_gate and_gate_h_u_cla32_and1669_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1669_y0);
  and_gate and_gate_h_u_cla32_and1670_y0(h_u_cla32_and1669_y0, h_u_cla32_and1668_y0, h_u_cla32_and1670_y0);
  and_gate and_gate_h_u_cla32_and1671_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1671_y0);
  and_gate and_gate_h_u_cla32_and1672_y0(h_u_cla32_and1671_y0, h_u_cla32_and1670_y0, h_u_cla32_and1672_y0);
  and_gate and_gate_h_u_cla32_and1673_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1673_y0);
  and_gate and_gate_h_u_cla32_and1674_y0(h_u_cla32_and1673_y0, h_u_cla32_and1672_y0, h_u_cla32_and1674_y0);
  and_gate and_gate_h_u_cla32_and1675_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1675_y0);
  and_gate and_gate_h_u_cla32_and1676_y0(h_u_cla32_and1675_y0, h_u_cla32_and1674_y0, h_u_cla32_and1676_y0);
  and_gate and_gate_h_u_cla32_and1677_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1677_y0);
  and_gate and_gate_h_u_cla32_and1678_y0(h_u_cla32_and1677_y0, h_u_cla32_and1676_y0, h_u_cla32_and1678_y0);
  and_gate and_gate_h_u_cla32_and1679_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1679_y0);
  and_gate and_gate_h_u_cla32_and1680_y0(h_u_cla32_and1679_y0, h_u_cla32_and1678_y0, h_u_cla32_and1680_y0);
  and_gate and_gate_h_u_cla32_and1681_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1681_y0);
  and_gate and_gate_h_u_cla32_and1682_y0(h_u_cla32_and1681_y0, h_u_cla32_and1680_y0, h_u_cla32_and1682_y0);
  and_gate and_gate_h_u_cla32_and1683_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1683_y0);
  and_gate and_gate_h_u_cla32_and1684_y0(h_u_cla32_and1683_y0, h_u_cla32_and1682_y0, h_u_cla32_and1684_y0);
  and_gate and_gate_h_u_cla32_and1685_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1685_y0);
  and_gate and_gate_h_u_cla32_and1686_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1686_y0);
  and_gate and_gate_h_u_cla32_and1687_y0(h_u_cla32_and1686_y0, h_u_cla32_and1685_y0, h_u_cla32_and1687_y0);
  and_gate and_gate_h_u_cla32_and1688_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1688_y0);
  and_gate and_gate_h_u_cla32_and1689_y0(h_u_cla32_and1688_y0, h_u_cla32_and1687_y0, h_u_cla32_and1689_y0);
  and_gate and_gate_h_u_cla32_and1690_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1690_y0);
  and_gate and_gate_h_u_cla32_and1691_y0(h_u_cla32_and1690_y0, h_u_cla32_and1689_y0, h_u_cla32_and1691_y0);
  and_gate and_gate_h_u_cla32_and1692_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1692_y0);
  and_gate and_gate_h_u_cla32_and1693_y0(h_u_cla32_and1692_y0, h_u_cla32_and1691_y0, h_u_cla32_and1693_y0);
  and_gate and_gate_h_u_cla32_and1694_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1694_y0);
  and_gate and_gate_h_u_cla32_and1695_y0(h_u_cla32_and1694_y0, h_u_cla32_and1693_y0, h_u_cla32_and1695_y0);
  and_gate and_gate_h_u_cla32_and1696_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1696_y0);
  and_gate and_gate_h_u_cla32_and1697_y0(h_u_cla32_and1696_y0, h_u_cla32_and1695_y0, h_u_cla32_and1697_y0);
  and_gate and_gate_h_u_cla32_and1698_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1698_y0);
  and_gate and_gate_h_u_cla32_and1699_y0(h_u_cla32_and1698_y0, h_u_cla32_and1697_y0, h_u_cla32_and1699_y0);
  and_gate and_gate_h_u_cla32_and1700_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1700_y0);
  and_gate and_gate_h_u_cla32_and1701_y0(h_u_cla32_and1700_y0, h_u_cla32_and1699_y0, h_u_cla32_and1701_y0);
  and_gate and_gate_h_u_cla32_and1702_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1702_y0);
  and_gate and_gate_h_u_cla32_and1703_y0(h_u_cla32_and1702_y0, h_u_cla32_and1701_y0, h_u_cla32_and1703_y0);
  and_gate and_gate_h_u_cla32_and1704_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1704_y0);
  and_gate and_gate_h_u_cla32_and1705_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1705_y0);
  and_gate and_gate_h_u_cla32_and1706_y0(h_u_cla32_and1705_y0, h_u_cla32_and1704_y0, h_u_cla32_and1706_y0);
  and_gate and_gate_h_u_cla32_and1707_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1707_y0);
  and_gate and_gate_h_u_cla32_and1708_y0(h_u_cla32_and1707_y0, h_u_cla32_and1706_y0, h_u_cla32_and1708_y0);
  and_gate and_gate_h_u_cla32_and1709_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1709_y0);
  and_gate and_gate_h_u_cla32_and1710_y0(h_u_cla32_and1709_y0, h_u_cla32_and1708_y0, h_u_cla32_and1710_y0);
  and_gate and_gate_h_u_cla32_and1711_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1711_y0);
  and_gate and_gate_h_u_cla32_and1712_y0(h_u_cla32_and1711_y0, h_u_cla32_and1710_y0, h_u_cla32_and1712_y0);
  and_gate and_gate_h_u_cla32_and1713_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1713_y0);
  and_gate and_gate_h_u_cla32_and1714_y0(h_u_cla32_and1713_y0, h_u_cla32_and1712_y0, h_u_cla32_and1714_y0);
  and_gate and_gate_h_u_cla32_and1715_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1715_y0);
  and_gate and_gate_h_u_cla32_and1716_y0(h_u_cla32_and1715_y0, h_u_cla32_and1714_y0, h_u_cla32_and1716_y0);
  and_gate and_gate_h_u_cla32_and1717_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1717_y0);
  and_gate and_gate_h_u_cla32_and1718_y0(h_u_cla32_and1717_y0, h_u_cla32_and1716_y0, h_u_cla32_and1718_y0);
  and_gate and_gate_h_u_cla32_and1719_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and1719_y0);
  and_gate and_gate_h_u_cla32_and1720_y0(h_u_cla32_and1719_y0, h_u_cla32_and1718_y0, h_u_cla32_and1720_y0);
  and_gate and_gate_h_u_cla32_and1721_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1721_y0);
  and_gate and_gate_h_u_cla32_and1722_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1722_y0);
  and_gate and_gate_h_u_cla32_and1723_y0(h_u_cla32_and1722_y0, h_u_cla32_and1721_y0, h_u_cla32_and1723_y0);
  and_gate and_gate_h_u_cla32_and1724_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1724_y0);
  and_gate and_gate_h_u_cla32_and1725_y0(h_u_cla32_and1724_y0, h_u_cla32_and1723_y0, h_u_cla32_and1725_y0);
  and_gate and_gate_h_u_cla32_and1726_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1726_y0);
  and_gate and_gate_h_u_cla32_and1727_y0(h_u_cla32_and1726_y0, h_u_cla32_and1725_y0, h_u_cla32_and1727_y0);
  and_gate and_gate_h_u_cla32_and1728_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1728_y0);
  and_gate and_gate_h_u_cla32_and1729_y0(h_u_cla32_and1728_y0, h_u_cla32_and1727_y0, h_u_cla32_and1729_y0);
  and_gate and_gate_h_u_cla32_and1730_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1730_y0);
  and_gate and_gate_h_u_cla32_and1731_y0(h_u_cla32_and1730_y0, h_u_cla32_and1729_y0, h_u_cla32_and1731_y0);
  and_gate and_gate_h_u_cla32_and1732_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1732_y0);
  and_gate and_gate_h_u_cla32_and1733_y0(h_u_cla32_and1732_y0, h_u_cla32_and1731_y0, h_u_cla32_and1733_y0);
  and_gate and_gate_h_u_cla32_and1734_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and1734_y0);
  and_gate and_gate_h_u_cla32_and1735_y0(h_u_cla32_and1734_y0, h_u_cla32_and1733_y0, h_u_cla32_and1735_y0);
  and_gate and_gate_h_u_cla32_and1736_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1736_y0);
  and_gate and_gate_h_u_cla32_and1737_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1737_y0);
  and_gate and_gate_h_u_cla32_and1738_y0(h_u_cla32_and1737_y0, h_u_cla32_and1736_y0, h_u_cla32_and1738_y0);
  and_gate and_gate_h_u_cla32_and1739_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1739_y0);
  and_gate and_gate_h_u_cla32_and1740_y0(h_u_cla32_and1739_y0, h_u_cla32_and1738_y0, h_u_cla32_and1740_y0);
  and_gate and_gate_h_u_cla32_and1741_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1741_y0);
  and_gate and_gate_h_u_cla32_and1742_y0(h_u_cla32_and1741_y0, h_u_cla32_and1740_y0, h_u_cla32_and1742_y0);
  and_gate and_gate_h_u_cla32_and1743_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1743_y0);
  and_gate and_gate_h_u_cla32_and1744_y0(h_u_cla32_and1743_y0, h_u_cla32_and1742_y0, h_u_cla32_and1744_y0);
  and_gate and_gate_h_u_cla32_and1745_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1745_y0);
  and_gate and_gate_h_u_cla32_and1746_y0(h_u_cla32_and1745_y0, h_u_cla32_and1744_y0, h_u_cla32_and1746_y0);
  and_gate and_gate_h_u_cla32_and1747_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and1747_y0);
  and_gate and_gate_h_u_cla32_and1748_y0(h_u_cla32_and1747_y0, h_u_cla32_and1746_y0, h_u_cla32_and1748_y0);
  and_gate and_gate_h_u_cla32_and1749_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1749_y0);
  and_gate and_gate_h_u_cla32_and1750_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1750_y0);
  and_gate and_gate_h_u_cla32_and1751_y0(h_u_cla32_and1750_y0, h_u_cla32_and1749_y0, h_u_cla32_and1751_y0);
  and_gate and_gate_h_u_cla32_and1752_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1752_y0);
  and_gate and_gate_h_u_cla32_and1753_y0(h_u_cla32_and1752_y0, h_u_cla32_and1751_y0, h_u_cla32_and1753_y0);
  and_gate and_gate_h_u_cla32_and1754_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1754_y0);
  and_gate and_gate_h_u_cla32_and1755_y0(h_u_cla32_and1754_y0, h_u_cla32_and1753_y0, h_u_cla32_and1755_y0);
  and_gate and_gate_h_u_cla32_and1756_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1756_y0);
  and_gate and_gate_h_u_cla32_and1757_y0(h_u_cla32_and1756_y0, h_u_cla32_and1755_y0, h_u_cla32_and1757_y0);
  and_gate and_gate_h_u_cla32_and1758_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and1758_y0);
  and_gate and_gate_h_u_cla32_and1759_y0(h_u_cla32_and1758_y0, h_u_cla32_and1757_y0, h_u_cla32_and1759_y0);
  and_gate and_gate_h_u_cla32_and1760_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1760_y0);
  and_gate and_gate_h_u_cla32_and1761_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1761_y0);
  and_gate and_gate_h_u_cla32_and1762_y0(h_u_cla32_and1761_y0, h_u_cla32_and1760_y0, h_u_cla32_and1762_y0);
  and_gate and_gate_h_u_cla32_and1763_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1763_y0);
  and_gate and_gate_h_u_cla32_and1764_y0(h_u_cla32_and1763_y0, h_u_cla32_and1762_y0, h_u_cla32_and1764_y0);
  and_gate and_gate_h_u_cla32_and1765_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1765_y0);
  and_gate and_gate_h_u_cla32_and1766_y0(h_u_cla32_and1765_y0, h_u_cla32_and1764_y0, h_u_cla32_and1766_y0);
  and_gate and_gate_h_u_cla32_and1767_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and1767_y0);
  and_gate and_gate_h_u_cla32_and1768_y0(h_u_cla32_and1767_y0, h_u_cla32_and1766_y0, h_u_cla32_and1768_y0);
  and_gate and_gate_h_u_cla32_and1769_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1769_y0);
  and_gate and_gate_h_u_cla32_and1770_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1770_y0);
  and_gate and_gate_h_u_cla32_and1771_y0(h_u_cla32_and1770_y0, h_u_cla32_and1769_y0, h_u_cla32_and1771_y0);
  and_gate and_gate_h_u_cla32_and1772_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1772_y0);
  and_gate and_gate_h_u_cla32_and1773_y0(h_u_cla32_and1772_y0, h_u_cla32_and1771_y0, h_u_cla32_and1773_y0);
  and_gate and_gate_h_u_cla32_and1774_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and1774_y0);
  and_gate and_gate_h_u_cla32_and1775_y0(h_u_cla32_and1774_y0, h_u_cla32_and1773_y0, h_u_cla32_and1775_y0);
  and_gate and_gate_h_u_cla32_and1776_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and1776_y0);
  and_gate and_gate_h_u_cla32_and1777_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and1777_y0);
  and_gate and_gate_h_u_cla32_and1778_y0(h_u_cla32_and1777_y0, h_u_cla32_and1776_y0, h_u_cla32_and1778_y0);
  and_gate and_gate_h_u_cla32_and1779_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and1779_y0);
  and_gate and_gate_h_u_cla32_and1780_y0(h_u_cla32_and1779_y0, h_u_cla32_and1778_y0, h_u_cla32_and1780_y0);
  and_gate and_gate_h_u_cla32_and1781_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and1781_y0);
  and_gate and_gate_h_u_cla32_and1782_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and1782_y0);
  and_gate and_gate_h_u_cla32_and1783_y0(h_u_cla32_and1782_y0, h_u_cla32_and1781_y0, h_u_cla32_and1783_y0);
  and_gate and_gate_h_u_cla32_and1784_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and1784_y0);
  or_gate or_gate_h_u_cla32_or136_y0(h_u_cla32_and1784_y0, h_u_cla32_and1528_y0, h_u_cla32_or136_y0);
  or_gate or_gate_h_u_cla32_or137_y0(h_u_cla32_or136_y0, h_u_cla32_and1559_y0, h_u_cla32_or137_y0);
  or_gate or_gate_h_u_cla32_or138_y0(h_u_cla32_or137_y0, h_u_cla32_and1588_y0, h_u_cla32_or138_y0);
  or_gate or_gate_h_u_cla32_or139_y0(h_u_cla32_or138_y0, h_u_cla32_and1615_y0, h_u_cla32_or139_y0);
  or_gate or_gate_h_u_cla32_or140_y0(h_u_cla32_or139_y0, h_u_cla32_and1640_y0, h_u_cla32_or140_y0);
  or_gate or_gate_h_u_cla32_or141_y0(h_u_cla32_or140_y0, h_u_cla32_and1663_y0, h_u_cla32_or141_y0);
  or_gate or_gate_h_u_cla32_or142_y0(h_u_cla32_or141_y0, h_u_cla32_and1684_y0, h_u_cla32_or142_y0);
  or_gate or_gate_h_u_cla32_or143_y0(h_u_cla32_or142_y0, h_u_cla32_and1703_y0, h_u_cla32_or143_y0);
  or_gate or_gate_h_u_cla32_or144_y0(h_u_cla32_or143_y0, h_u_cla32_and1720_y0, h_u_cla32_or144_y0);
  or_gate or_gate_h_u_cla32_or145_y0(h_u_cla32_or144_y0, h_u_cla32_and1735_y0, h_u_cla32_or145_y0);
  or_gate or_gate_h_u_cla32_or146_y0(h_u_cla32_or145_y0, h_u_cla32_and1748_y0, h_u_cla32_or146_y0);
  or_gate or_gate_h_u_cla32_or147_y0(h_u_cla32_or146_y0, h_u_cla32_and1759_y0, h_u_cla32_or147_y0);
  or_gate or_gate_h_u_cla32_or148_y0(h_u_cla32_or147_y0, h_u_cla32_and1768_y0, h_u_cla32_or148_y0);
  or_gate or_gate_h_u_cla32_or149_y0(h_u_cla32_or148_y0, h_u_cla32_and1775_y0, h_u_cla32_or149_y0);
  or_gate or_gate_h_u_cla32_or150_y0(h_u_cla32_or149_y0, h_u_cla32_and1780_y0, h_u_cla32_or150_y0);
  or_gate or_gate_h_u_cla32_or151_y0(h_u_cla32_or150_y0, h_u_cla32_and1783_y0, h_u_cla32_or151_y0);
  or_gate or_gate_h_u_cla32_or152_y0(h_u_cla32_pg_logic16_y1, h_u_cla32_or151_y0, h_u_cla32_or152_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic17_y0(a_17, b_17, h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_pg_logic17_y2);
  xor_gate xor_gate_h_u_cla32_xor17_y0(h_u_cla32_pg_logic17_y2, h_u_cla32_or152_y0, h_u_cla32_xor17_y0);
  and_gate and_gate_h_u_cla32_and1785_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and1785_y0);
  and_gate and_gate_h_u_cla32_and1786_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and1786_y0);
  and_gate and_gate_h_u_cla32_and1787_y0(h_u_cla32_and1786_y0, h_u_cla32_and1785_y0, h_u_cla32_and1787_y0);
  and_gate and_gate_h_u_cla32_and1788_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and1788_y0);
  and_gate and_gate_h_u_cla32_and1789_y0(h_u_cla32_and1788_y0, h_u_cla32_and1787_y0, h_u_cla32_and1789_y0);
  and_gate and_gate_h_u_cla32_and1790_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and1790_y0);
  and_gate and_gate_h_u_cla32_and1791_y0(h_u_cla32_and1790_y0, h_u_cla32_and1789_y0, h_u_cla32_and1791_y0);
  and_gate and_gate_h_u_cla32_and1792_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and1792_y0);
  and_gate and_gate_h_u_cla32_and1793_y0(h_u_cla32_and1792_y0, h_u_cla32_and1791_y0, h_u_cla32_and1793_y0);
  and_gate and_gate_h_u_cla32_and1794_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and1794_y0);
  and_gate and_gate_h_u_cla32_and1795_y0(h_u_cla32_and1794_y0, h_u_cla32_and1793_y0, h_u_cla32_and1795_y0);
  and_gate and_gate_h_u_cla32_and1796_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and1796_y0);
  and_gate and_gate_h_u_cla32_and1797_y0(h_u_cla32_and1796_y0, h_u_cla32_and1795_y0, h_u_cla32_and1797_y0);
  and_gate and_gate_h_u_cla32_and1798_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and1798_y0);
  and_gate and_gate_h_u_cla32_and1799_y0(h_u_cla32_and1798_y0, h_u_cla32_and1797_y0, h_u_cla32_and1799_y0);
  and_gate and_gate_h_u_cla32_and1800_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and1800_y0);
  and_gate and_gate_h_u_cla32_and1801_y0(h_u_cla32_and1800_y0, h_u_cla32_and1799_y0, h_u_cla32_and1801_y0);
  and_gate and_gate_h_u_cla32_and1802_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and1802_y0);
  and_gate and_gate_h_u_cla32_and1803_y0(h_u_cla32_and1802_y0, h_u_cla32_and1801_y0, h_u_cla32_and1803_y0);
  and_gate and_gate_h_u_cla32_and1804_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and1804_y0);
  and_gate and_gate_h_u_cla32_and1805_y0(h_u_cla32_and1804_y0, h_u_cla32_and1803_y0, h_u_cla32_and1805_y0);
  and_gate and_gate_h_u_cla32_and1806_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and1806_y0);
  and_gate and_gate_h_u_cla32_and1807_y0(h_u_cla32_and1806_y0, h_u_cla32_and1805_y0, h_u_cla32_and1807_y0);
  and_gate and_gate_h_u_cla32_and1808_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and1808_y0);
  and_gate and_gate_h_u_cla32_and1809_y0(h_u_cla32_and1808_y0, h_u_cla32_and1807_y0, h_u_cla32_and1809_y0);
  and_gate and_gate_h_u_cla32_and1810_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and1810_y0);
  and_gate and_gate_h_u_cla32_and1811_y0(h_u_cla32_and1810_y0, h_u_cla32_and1809_y0, h_u_cla32_and1811_y0);
  and_gate and_gate_h_u_cla32_and1812_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and1812_y0);
  and_gate and_gate_h_u_cla32_and1813_y0(h_u_cla32_and1812_y0, h_u_cla32_and1811_y0, h_u_cla32_and1813_y0);
  and_gate and_gate_h_u_cla32_and1814_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and1814_y0);
  and_gate and_gate_h_u_cla32_and1815_y0(h_u_cla32_and1814_y0, h_u_cla32_and1813_y0, h_u_cla32_and1815_y0);
  and_gate and_gate_h_u_cla32_and1816_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and1816_y0);
  and_gate and_gate_h_u_cla32_and1817_y0(h_u_cla32_and1816_y0, h_u_cla32_and1815_y0, h_u_cla32_and1817_y0);
  and_gate and_gate_h_u_cla32_and1818_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and1818_y0);
  and_gate and_gate_h_u_cla32_and1819_y0(h_u_cla32_and1818_y0, h_u_cla32_and1817_y0, h_u_cla32_and1819_y0);
  and_gate and_gate_h_u_cla32_and1820_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1820_y0);
  and_gate and_gate_h_u_cla32_and1821_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1821_y0);
  and_gate and_gate_h_u_cla32_and1822_y0(h_u_cla32_and1821_y0, h_u_cla32_and1820_y0, h_u_cla32_and1822_y0);
  and_gate and_gate_h_u_cla32_and1823_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1823_y0);
  and_gate and_gate_h_u_cla32_and1824_y0(h_u_cla32_and1823_y0, h_u_cla32_and1822_y0, h_u_cla32_and1824_y0);
  and_gate and_gate_h_u_cla32_and1825_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1825_y0);
  and_gate and_gate_h_u_cla32_and1826_y0(h_u_cla32_and1825_y0, h_u_cla32_and1824_y0, h_u_cla32_and1826_y0);
  and_gate and_gate_h_u_cla32_and1827_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1827_y0);
  and_gate and_gate_h_u_cla32_and1828_y0(h_u_cla32_and1827_y0, h_u_cla32_and1826_y0, h_u_cla32_and1828_y0);
  and_gate and_gate_h_u_cla32_and1829_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1829_y0);
  and_gate and_gate_h_u_cla32_and1830_y0(h_u_cla32_and1829_y0, h_u_cla32_and1828_y0, h_u_cla32_and1830_y0);
  and_gate and_gate_h_u_cla32_and1831_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1831_y0);
  and_gate and_gate_h_u_cla32_and1832_y0(h_u_cla32_and1831_y0, h_u_cla32_and1830_y0, h_u_cla32_and1832_y0);
  and_gate and_gate_h_u_cla32_and1833_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1833_y0);
  and_gate and_gate_h_u_cla32_and1834_y0(h_u_cla32_and1833_y0, h_u_cla32_and1832_y0, h_u_cla32_and1834_y0);
  and_gate and_gate_h_u_cla32_and1835_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1835_y0);
  and_gate and_gate_h_u_cla32_and1836_y0(h_u_cla32_and1835_y0, h_u_cla32_and1834_y0, h_u_cla32_and1836_y0);
  and_gate and_gate_h_u_cla32_and1837_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1837_y0);
  and_gate and_gate_h_u_cla32_and1838_y0(h_u_cla32_and1837_y0, h_u_cla32_and1836_y0, h_u_cla32_and1838_y0);
  and_gate and_gate_h_u_cla32_and1839_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1839_y0);
  and_gate and_gate_h_u_cla32_and1840_y0(h_u_cla32_and1839_y0, h_u_cla32_and1838_y0, h_u_cla32_and1840_y0);
  and_gate and_gate_h_u_cla32_and1841_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1841_y0);
  and_gate and_gate_h_u_cla32_and1842_y0(h_u_cla32_and1841_y0, h_u_cla32_and1840_y0, h_u_cla32_and1842_y0);
  and_gate and_gate_h_u_cla32_and1843_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1843_y0);
  and_gate and_gate_h_u_cla32_and1844_y0(h_u_cla32_and1843_y0, h_u_cla32_and1842_y0, h_u_cla32_and1844_y0);
  and_gate and_gate_h_u_cla32_and1845_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1845_y0);
  and_gate and_gate_h_u_cla32_and1846_y0(h_u_cla32_and1845_y0, h_u_cla32_and1844_y0, h_u_cla32_and1846_y0);
  and_gate and_gate_h_u_cla32_and1847_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1847_y0);
  and_gate and_gate_h_u_cla32_and1848_y0(h_u_cla32_and1847_y0, h_u_cla32_and1846_y0, h_u_cla32_and1848_y0);
  and_gate and_gate_h_u_cla32_and1849_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1849_y0);
  and_gate and_gate_h_u_cla32_and1850_y0(h_u_cla32_and1849_y0, h_u_cla32_and1848_y0, h_u_cla32_and1850_y0);
  and_gate and_gate_h_u_cla32_and1851_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and1851_y0);
  and_gate and_gate_h_u_cla32_and1852_y0(h_u_cla32_and1851_y0, h_u_cla32_and1850_y0, h_u_cla32_and1852_y0);
  and_gate and_gate_h_u_cla32_and1853_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1853_y0);
  and_gate and_gate_h_u_cla32_and1854_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1854_y0);
  and_gate and_gate_h_u_cla32_and1855_y0(h_u_cla32_and1854_y0, h_u_cla32_and1853_y0, h_u_cla32_and1855_y0);
  and_gate and_gate_h_u_cla32_and1856_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1856_y0);
  and_gate and_gate_h_u_cla32_and1857_y0(h_u_cla32_and1856_y0, h_u_cla32_and1855_y0, h_u_cla32_and1857_y0);
  and_gate and_gate_h_u_cla32_and1858_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1858_y0);
  and_gate and_gate_h_u_cla32_and1859_y0(h_u_cla32_and1858_y0, h_u_cla32_and1857_y0, h_u_cla32_and1859_y0);
  and_gate and_gate_h_u_cla32_and1860_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1860_y0);
  and_gate and_gate_h_u_cla32_and1861_y0(h_u_cla32_and1860_y0, h_u_cla32_and1859_y0, h_u_cla32_and1861_y0);
  and_gate and_gate_h_u_cla32_and1862_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1862_y0);
  and_gate and_gate_h_u_cla32_and1863_y0(h_u_cla32_and1862_y0, h_u_cla32_and1861_y0, h_u_cla32_and1863_y0);
  and_gate and_gate_h_u_cla32_and1864_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1864_y0);
  and_gate and_gate_h_u_cla32_and1865_y0(h_u_cla32_and1864_y0, h_u_cla32_and1863_y0, h_u_cla32_and1865_y0);
  and_gate and_gate_h_u_cla32_and1866_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1866_y0);
  and_gate and_gate_h_u_cla32_and1867_y0(h_u_cla32_and1866_y0, h_u_cla32_and1865_y0, h_u_cla32_and1867_y0);
  and_gate and_gate_h_u_cla32_and1868_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1868_y0);
  and_gate and_gate_h_u_cla32_and1869_y0(h_u_cla32_and1868_y0, h_u_cla32_and1867_y0, h_u_cla32_and1869_y0);
  and_gate and_gate_h_u_cla32_and1870_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1870_y0);
  and_gate and_gate_h_u_cla32_and1871_y0(h_u_cla32_and1870_y0, h_u_cla32_and1869_y0, h_u_cla32_and1871_y0);
  and_gate and_gate_h_u_cla32_and1872_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1872_y0);
  and_gate and_gate_h_u_cla32_and1873_y0(h_u_cla32_and1872_y0, h_u_cla32_and1871_y0, h_u_cla32_and1873_y0);
  and_gate and_gate_h_u_cla32_and1874_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1874_y0);
  and_gate and_gate_h_u_cla32_and1875_y0(h_u_cla32_and1874_y0, h_u_cla32_and1873_y0, h_u_cla32_and1875_y0);
  and_gate and_gate_h_u_cla32_and1876_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1876_y0);
  and_gate and_gate_h_u_cla32_and1877_y0(h_u_cla32_and1876_y0, h_u_cla32_and1875_y0, h_u_cla32_and1877_y0);
  and_gate and_gate_h_u_cla32_and1878_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1878_y0);
  and_gate and_gate_h_u_cla32_and1879_y0(h_u_cla32_and1878_y0, h_u_cla32_and1877_y0, h_u_cla32_and1879_y0);
  and_gate and_gate_h_u_cla32_and1880_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1880_y0);
  and_gate and_gate_h_u_cla32_and1881_y0(h_u_cla32_and1880_y0, h_u_cla32_and1879_y0, h_u_cla32_and1881_y0);
  and_gate and_gate_h_u_cla32_and1882_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and1882_y0);
  and_gate and_gate_h_u_cla32_and1883_y0(h_u_cla32_and1882_y0, h_u_cla32_and1881_y0, h_u_cla32_and1883_y0);
  and_gate and_gate_h_u_cla32_and1884_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1884_y0);
  and_gate and_gate_h_u_cla32_and1885_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1885_y0);
  and_gate and_gate_h_u_cla32_and1886_y0(h_u_cla32_and1885_y0, h_u_cla32_and1884_y0, h_u_cla32_and1886_y0);
  and_gate and_gate_h_u_cla32_and1887_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1887_y0);
  and_gate and_gate_h_u_cla32_and1888_y0(h_u_cla32_and1887_y0, h_u_cla32_and1886_y0, h_u_cla32_and1888_y0);
  and_gate and_gate_h_u_cla32_and1889_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1889_y0);
  and_gate and_gate_h_u_cla32_and1890_y0(h_u_cla32_and1889_y0, h_u_cla32_and1888_y0, h_u_cla32_and1890_y0);
  and_gate and_gate_h_u_cla32_and1891_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1891_y0);
  and_gate and_gate_h_u_cla32_and1892_y0(h_u_cla32_and1891_y0, h_u_cla32_and1890_y0, h_u_cla32_and1892_y0);
  and_gate and_gate_h_u_cla32_and1893_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1893_y0);
  and_gate and_gate_h_u_cla32_and1894_y0(h_u_cla32_and1893_y0, h_u_cla32_and1892_y0, h_u_cla32_and1894_y0);
  and_gate and_gate_h_u_cla32_and1895_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1895_y0);
  and_gate and_gate_h_u_cla32_and1896_y0(h_u_cla32_and1895_y0, h_u_cla32_and1894_y0, h_u_cla32_and1896_y0);
  and_gate and_gate_h_u_cla32_and1897_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1897_y0);
  and_gate and_gate_h_u_cla32_and1898_y0(h_u_cla32_and1897_y0, h_u_cla32_and1896_y0, h_u_cla32_and1898_y0);
  and_gate and_gate_h_u_cla32_and1899_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1899_y0);
  and_gate and_gate_h_u_cla32_and1900_y0(h_u_cla32_and1899_y0, h_u_cla32_and1898_y0, h_u_cla32_and1900_y0);
  and_gate and_gate_h_u_cla32_and1901_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1901_y0);
  and_gate and_gate_h_u_cla32_and1902_y0(h_u_cla32_and1901_y0, h_u_cla32_and1900_y0, h_u_cla32_and1902_y0);
  and_gate and_gate_h_u_cla32_and1903_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1903_y0);
  and_gate and_gate_h_u_cla32_and1904_y0(h_u_cla32_and1903_y0, h_u_cla32_and1902_y0, h_u_cla32_and1904_y0);
  and_gate and_gate_h_u_cla32_and1905_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1905_y0);
  and_gate and_gate_h_u_cla32_and1906_y0(h_u_cla32_and1905_y0, h_u_cla32_and1904_y0, h_u_cla32_and1906_y0);
  and_gate and_gate_h_u_cla32_and1907_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1907_y0);
  and_gate and_gate_h_u_cla32_and1908_y0(h_u_cla32_and1907_y0, h_u_cla32_and1906_y0, h_u_cla32_and1908_y0);
  and_gate and_gate_h_u_cla32_and1909_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1909_y0);
  and_gate and_gate_h_u_cla32_and1910_y0(h_u_cla32_and1909_y0, h_u_cla32_and1908_y0, h_u_cla32_and1910_y0);
  and_gate and_gate_h_u_cla32_and1911_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and1911_y0);
  and_gate and_gate_h_u_cla32_and1912_y0(h_u_cla32_and1911_y0, h_u_cla32_and1910_y0, h_u_cla32_and1912_y0);
  and_gate and_gate_h_u_cla32_and1913_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1913_y0);
  and_gate and_gate_h_u_cla32_and1914_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1914_y0);
  and_gate and_gate_h_u_cla32_and1915_y0(h_u_cla32_and1914_y0, h_u_cla32_and1913_y0, h_u_cla32_and1915_y0);
  and_gate and_gate_h_u_cla32_and1916_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1916_y0);
  and_gate and_gate_h_u_cla32_and1917_y0(h_u_cla32_and1916_y0, h_u_cla32_and1915_y0, h_u_cla32_and1917_y0);
  and_gate and_gate_h_u_cla32_and1918_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1918_y0);
  and_gate and_gate_h_u_cla32_and1919_y0(h_u_cla32_and1918_y0, h_u_cla32_and1917_y0, h_u_cla32_and1919_y0);
  and_gate and_gate_h_u_cla32_and1920_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1920_y0);
  and_gate and_gate_h_u_cla32_and1921_y0(h_u_cla32_and1920_y0, h_u_cla32_and1919_y0, h_u_cla32_and1921_y0);
  and_gate and_gate_h_u_cla32_and1922_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1922_y0);
  and_gate and_gate_h_u_cla32_and1923_y0(h_u_cla32_and1922_y0, h_u_cla32_and1921_y0, h_u_cla32_and1923_y0);
  and_gate and_gate_h_u_cla32_and1924_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1924_y0);
  and_gate and_gate_h_u_cla32_and1925_y0(h_u_cla32_and1924_y0, h_u_cla32_and1923_y0, h_u_cla32_and1925_y0);
  and_gate and_gate_h_u_cla32_and1926_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1926_y0);
  and_gate and_gate_h_u_cla32_and1927_y0(h_u_cla32_and1926_y0, h_u_cla32_and1925_y0, h_u_cla32_and1927_y0);
  and_gate and_gate_h_u_cla32_and1928_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1928_y0);
  and_gate and_gate_h_u_cla32_and1929_y0(h_u_cla32_and1928_y0, h_u_cla32_and1927_y0, h_u_cla32_and1929_y0);
  and_gate and_gate_h_u_cla32_and1930_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1930_y0);
  and_gate and_gate_h_u_cla32_and1931_y0(h_u_cla32_and1930_y0, h_u_cla32_and1929_y0, h_u_cla32_and1931_y0);
  and_gate and_gate_h_u_cla32_and1932_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1932_y0);
  and_gate and_gate_h_u_cla32_and1933_y0(h_u_cla32_and1932_y0, h_u_cla32_and1931_y0, h_u_cla32_and1933_y0);
  and_gate and_gate_h_u_cla32_and1934_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1934_y0);
  and_gate and_gate_h_u_cla32_and1935_y0(h_u_cla32_and1934_y0, h_u_cla32_and1933_y0, h_u_cla32_and1935_y0);
  and_gate and_gate_h_u_cla32_and1936_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1936_y0);
  and_gate and_gate_h_u_cla32_and1937_y0(h_u_cla32_and1936_y0, h_u_cla32_and1935_y0, h_u_cla32_and1937_y0);
  and_gate and_gate_h_u_cla32_and1938_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and1938_y0);
  and_gate and_gate_h_u_cla32_and1939_y0(h_u_cla32_and1938_y0, h_u_cla32_and1937_y0, h_u_cla32_and1939_y0);
  and_gate and_gate_h_u_cla32_and1940_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1940_y0);
  and_gate and_gate_h_u_cla32_and1941_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1941_y0);
  and_gate and_gate_h_u_cla32_and1942_y0(h_u_cla32_and1941_y0, h_u_cla32_and1940_y0, h_u_cla32_and1942_y0);
  and_gate and_gate_h_u_cla32_and1943_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1943_y0);
  and_gate and_gate_h_u_cla32_and1944_y0(h_u_cla32_and1943_y0, h_u_cla32_and1942_y0, h_u_cla32_and1944_y0);
  and_gate and_gate_h_u_cla32_and1945_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1945_y0);
  and_gate and_gate_h_u_cla32_and1946_y0(h_u_cla32_and1945_y0, h_u_cla32_and1944_y0, h_u_cla32_and1946_y0);
  and_gate and_gate_h_u_cla32_and1947_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1947_y0);
  and_gate and_gate_h_u_cla32_and1948_y0(h_u_cla32_and1947_y0, h_u_cla32_and1946_y0, h_u_cla32_and1948_y0);
  and_gate and_gate_h_u_cla32_and1949_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1949_y0);
  and_gate and_gate_h_u_cla32_and1950_y0(h_u_cla32_and1949_y0, h_u_cla32_and1948_y0, h_u_cla32_and1950_y0);
  and_gate and_gate_h_u_cla32_and1951_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1951_y0);
  and_gate and_gate_h_u_cla32_and1952_y0(h_u_cla32_and1951_y0, h_u_cla32_and1950_y0, h_u_cla32_and1952_y0);
  and_gate and_gate_h_u_cla32_and1953_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1953_y0);
  and_gate and_gate_h_u_cla32_and1954_y0(h_u_cla32_and1953_y0, h_u_cla32_and1952_y0, h_u_cla32_and1954_y0);
  and_gate and_gate_h_u_cla32_and1955_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1955_y0);
  and_gate and_gate_h_u_cla32_and1956_y0(h_u_cla32_and1955_y0, h_u_cla32_and1954_y0, h_u_cla32_and1956_y0);
  and_gate and_gate_h_u_cla32_and1957_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1957_y0);
  and_gate and_gate_h_u_cla32_and1958_y0(h_u_cla32_and1957_y0, h_u_cla32_and1956_y0, h_u_cla32_and1958_y0);
  and_gate and_gate_h_u_cla32_and1959_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1959_y0);
  and_gate and_gate_h_u_cla32_and1960_y0(h_u_cla32_and1959_y0, h_u_cla32_and1958_y0, h_u_cla32_and1960_y0);
  and_gate and_gate_h_u_cla32_and1961_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1961_y0);
  and_gate and_gate_h_u_cla32_and1962_y0(h_u_cla32_and1961_y0, h_u_cla32_and1960_y0, h_u_cla32_and1962_y0);
  and_gate and_gate_h_u_cla32_and1963_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and1963_y0);
  and_gate and_gate_h_u_cla32_and1964_y0(h_u_cla32_and1963_y0, h_u_cla32_and1962_y0, h_u_cla32_and1964_y0);
  and_gate and_gate_h_u_cla32_and1965_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1965_y0);
  and_gate and_gate_h_u_cla32_and1966_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1966_y0);
  and_gate and_gate_h_u_cla32_and1967_y0(h_u_cla32_and1966_y0, h_u_cla32_and1965_y0, h_u_cla32_and1967_y0);
  and_gate and_gate_h_u_cla32_and1968_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1968_y0);
  and_gate and_gate_h_u_cla32_and1969_y0(h_u_cla32_and1968_y0, h_u_cla32_and1967_y0, h_u_cla32_and1969_y0);
  and_gate and_gate_h_u_cla32_and1970_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1970_y0);
  and_gate and_gate_h_u_cla32_and1971_y0(h_u_cla32_and1970_y0, h_u_cla32_and1969_y0, h_u_cla32_and1971_y0);
  and_gate and_gate_h_u_cla32_and1972_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1972_y0);
  and_gate and_gate_h_u_cla32_and1973_y0(h_u_cla32_and1972_y0, h_u_cla32_and1971_y0, h_u_cla32_and1973_y0);
  and_gate and_gate_h_u_cla32_and1974_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1974_y0);
  and_gate and_gate_h_u_cla32_and1975_y0(h_u_cla32_and1974_y0, h_u_cla32_and1973_y0, h_u_cla32_and1975_y0);
  and_gate and_gate_h_u_cla32_and1976_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1976_y0);
  and_gate and_gate_h_u_cla32_and1977_y0(h_u_cla32_and1976_y0, h_u_cla32_and1975_y0, h_u_cla32_and1977_y0);
  and_gate and_gate_h_u_cla32_and1978_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1978_y0);
  and_gate and_gate_h_u_cla32_and1979_y0(h_u_cla32_and1978_y0, h_u_cla32_and1977_y0, h_u_cla32_and1979_y0);
  and_gate and_gate_h_u_cla32_and1980_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1980_y0);
  and_gate and_gate_h_u_cla32_and1981_y0(h_u_cla32_and1980_y0, h_u_cla32_and1979_y0, h_u_cla32_and1981_y0);
  and_gate and_gate_h_u_cla32_and1982_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1982_y0);
  and_gate and_gate_h_u_cla32_and1983_y0(h_u_cla32_and1982_y0, h_u_cla32_and1981_y0, h_u_cla32_and1983_y0);
  and_gate and_gate_h_u_cla32_and1984_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1984_y0);
  and_gate and_gate_h_u_cla32_and1985_y0(h_u_cla32_and1984_y0, h_u_cla32_and1983_y0, h_u_cla32_and1985_y0);
  and_gate and_gate_h_u_cla32_and1986_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and1986_y0);
  and_gate and_gate_h_u_cla32_and1987_y0(h_u_cla32_and1986_y0, h_u_cla32_and1985_y0, h_u_cla32_and1987_y0);
  and_gate and_gate_h_u_cla32_and1988_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1988_y0);
  and_gate and_gate_h_u_cla32_and1989_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1989_y0);
  and_gate and_gate_h_u_cla32_and1990_y0(h_u_cla32_and1989_y0, h_u_cla32_and1988_y0, h_u_cla32_and1990_y0);
  and_gate and_gate_h_u_cla32_and1991_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1991_y0);
  and_gate and_gate_h_u_cla32_and1992_y0(h_u_cla32_and1991_y0, h_u_cla32_and1990_y0, h_u_cla32_and1992_y0);
  and_gate and_gate_h_u_cla32_and1993_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1993_y0);
  and_gate and_gate_h_u_cla32_and1994_y0(h_u_cla32_and1993_y0, h_u_cla32_and1992_y0, h_u_cla32_and1994_y0);
  and_gate and_gate_h_u_cla32_and1995_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1995_y0);
  and_gate and_gate_h_u_cla32_and1996_y0(h_u_cla32_and1995_y0, h_u_cla32_and1994_y0, h_u_cla32_and1996_y0);
  and_gate and_gate_h_u_cla32_and1997_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1997_y0);
  and_gate and_gate_h_u_cla32_and1998_y0(h_u_cla32_and1997_y0, h_u_cla32_and1996_y0, h_u_cla32_and1998_y0);
  and_gate and_gate_h_u_cla32_and1999_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and1999_y0);
  and_gate and_gate_h_u_cla32_and2000_y0(h_u_cla32_and1999_y0, h_u_cla32_and1998_y0, h_u_cla32_and2000_y0);
  and_gate and_gate_h_u_cla32_and2001_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2001_y0);
  and_gate and_gate_h_u_cla32_and2002_y0(h_u_cla32_and2001_y0, h_u_cla32_and2000_y0, h_u_cla32_and2002_y0);
  and_gate and_gate_h_u_cla32_and2003_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2003_y0);
  and_gate and_gate_h_u_cla32_and2004_y0(h_u_cla32_and2003_y0, h_u_cla32_and2002_y0, h_u_cla32_and2004_y0);
  and_gate and_gate_h_u_cla32_and2005_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2005_y0);
  and_gate and_gate_h_u_cla32_and2006_y0(h_u_cla32_and2005_y0, h_u_cla32_and2004_y0, h_u_cla32_and2006_y0);
  and_gate and_gate_h_u_cla32_and2007_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2007_y0);
  and_gate and_gate_h_u_cla32_and2008_y0(h_u_cla32_and2007_y0, h_u_cla32_and2006_y0, h_u_cla32_and2008_y0);
  and_gate and_gate_h_u_cla32_and2009_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2009_y0);
  and_gate and_gate_h_u_cla32_and2010_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2010_y0);
  and_gate and_gate_h_u_cla32_and2011_y0(h_u_cla32_and2010_y0, h_u_cla32_and2009_y0, h_u_cla32_and2011_y0);
  and_gate and_gate_h_u_cla32_and2012_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2012_y0);
  and_gate and_gate_h_u_cla32_and2013_y0(h_u_cla32_and2012_y0, h_u_cla32_and2011_y0, h_u_cla32_and2013_y0);
  and_gate and_gate_h_u_cla32_and2014_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2014_y0);
  and_gate and_gate_h_u_cla32_and2015_y0(h_u_cla32_and2014_y0, h_u_cla32_and2013_y0, h_u_cla32_and2015_y0);
  and_gate and_gate_h_u_cla32_and2016_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2016_y0);
  and_gate and_gate_h_u_cla32_and2017_y0(h_u_cla32_and2016_y0, h_u_cla32_and2015_y0, h_u_cla32_and2017_y0);
  and_gate and_gate_h_u_cla32_and2018_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2018_y0);
  and_gate and_gate_h_u_cla32_and2019_y0(h_u_cla32_and2018_y0, h_u_cla32_and2017_y0, h_u_cla32_and2019_y0);
  and_gate and_gate_h_u_cla32_and2020_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2020_y0);
  and_gate and_gate_h_u_cla32_and2021_y0(h_u_cla32_and2020_y0, h_u_cla32_and2019_y0, h_u_cla32_and2021_y0);
  and_gate and_gate_h_u_cla32_and2022_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2022_y0);
  and_gate and_gate_h_u_cla32_and2023_y0(h_u_cla32_and2022_y0, h_u_cla32_and2021_y0, h_u_cla32_and2023_y0);
  and_gate and_gate_h_u_cla32_and2024_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2024_y0);
  and_gate and_gate_h_u_cla32_and2025_y0(h_u_cla32_and2024_y0, h_u_cla32_and2023_y0, h_u_cla32_and2025_y0);
  and_gate and_gate_h_u_cla32_and2026_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2026_y0);
  and_gate and_gate_h_u_cla32_and2027_y0(h_u_cla32_and2026_y0, h_u_cla32_and2025_y0, h_u_cla32_and2027_y0);
  and_gate and_gate_h_u_cla32_and2028_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2028_y0);
  and_gate and_gate_h_u_cla32_and2029_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2029_y0);
  and_gate and_gate_h_u_cla32_and2030_y0(h_u_cla32_and2029_y0, h_u_cla32_and2028_y0, h_u_cla32_and2030_y0);
  and_gate and_gate_h_u_cla32_and2031_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2031_y0);
  and_gate and_gate_h_u_cla32_and2032_y0(h_u_cla32_and2031_y0, h_u_cla32_and2030_y0, h_u_cla32_and2032_y0);
  and_gate and_gate_h_u_cla32_and2033_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2033_y0);
  and_gate and_gate_h_u_cla32_and2034_y0(h_u_cla32_and2033_y0, h_u_cla32_and2032_y0, h_u_cla32_and2034_y0);
  and_gate and_gate_h_u_cla32_and2035_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2035_y0);
  and_gate and_gate_h_u_cla32_and2036_y0(h_u_cla32_and2035_y0, h_u_cla32_and2034_y0, h_u_cla32_and2036_y0);
  and_gate and_gate_h_u_cla32_and2037_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2037_y0);
  and_gate and_gate_h_u_cla32_and2038_y0(h_u_cla32_and2037_y0, h_u_cla32_and2036_y0, h_u_cla32_and2038_y0);
  and_gate and_gate_h_u_cla32_and2039_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2039_y0);
  and_gate and_gate_h_u_cla32_and2040_y0(h_u_cla32_and2039_y0, h_u_cla32_and2038_y0, h_u_cla32_and2040_y0);
  and_gate and_gate_h_u_cla32_and2041_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2041_y0);
  and_gate and_gate_h_u_cla32_and2042_y0(h_u_cla32_and2041_y0, h_u_cla32_and2040_y0, h_u_cla32_and2042_y0);
  and_gate and_gate_h_u_cla32_and2043_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2043_y0);
  and_gate and_gate_h_u_cla32_and2044_y0(h_u_cla32_and2043_y0, h_u_cla32_and2042_y0, h_u_cla32_and2044_y0);
  and_gate and_gate_h_u_cla32_and2045_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2045_y0);
  and_gate and_gate_h_u_cla32_and2046_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2046_y0);
  and_gate and_gate_h_u_cla32_and2047_y0(h_u_cla32_and2046_y0, h_u_cla32_and2045_y0, h_u_cla32_and2047_y0);
  and_gate and_gate_h_u_cla32_and2048_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2048_y0);
  and_gate and_gate_h_u_cla32_and2049_y0(h_u_cla32_and2048_y0, h_u_cla32_and2047_y0, h_u_cla32_and2049_y0);
  and_gate and_gate_h_u_cla32_and2050_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2050_y0);
  and_gate and_gate_h_u_cla32_and2051_y0(h_u_cla32_and2050_y0, h_u_cla32_and2049_y0, h_u_cla32_and2051_y0);
  and_gate and_gate_h_u_cla32_and2052_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2052_y0);
  and_gate and_gate_h_u_cla32_and2053_y0(h_u_cla32_and2052_y0, h_u_cla32_and2051_y0, h_u_cla32_and2053_y0);
  and_gate and_gate_h_u_cla32_and2054_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2054_y0);
  and_gate and_gate_h_u_cla32_and2055_y0(h_u_cla32_and2054_y0, h_u_cla32_and2053_y0, h_u_cla32_and2055_y0);
  and_gate and_gate_h_u_cla32_and2056_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2056_y0);
  and_gate and_gate_h_u_cla32_and2057_y0(h_u_cla32_and2056_y0, h_u_cla32_and2055_y0, h_u_cla32_and2057_y0);
  and_gate and_gate_h_u_cla32_and2058_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2058_y0);
  and_gate and_gate_h_u_cla32_and2059_y0(h_u_cla32_and2058_y0, h_u_cla32_and2057_y0, h_u_cla32_and2059_y0);
  and_gate and_gate_h_u_cla32_and2060_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2060_y0);
  and_gate and_gate_h_u_cla32_and2061_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2061_y0);
  and_gate and_gate_h_u_cla32_and2062_y0(h_u_cla32_and2061_y0, h_u_cla32_and2060_y0, h_u_cla32_and2062_y0);
  and_gate and_gate_h_u_cla32_and2063_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2063_y0);
  and_gate and_gate_h_u_cla32_and2064_y0(h_u_cla32_and2063_y0, h_u_cla32_and2062_y0, h_u_cla32_and2064_y0);
  and_gate and_gate_h_u_cla32_and2065_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2065_y0);
  and_gate and_gate_h_u_cla32_and2066_y0(h_u_cla32_and2065_y0, h_u_cla32_and2064_y0, h_u_cla32_and2066_y0);
  and_gate and_gate_h_u_cla32_and2067_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2067_y0);
  and_gate and_gate_h_u_cla32_and2068_y0(h_u_cla32_and2067_y0, h_u_cla32_and2066_y0, h_u_cla32_and2068_y0);
  and_gate and_gate_h_u_cla32_and2069_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2069_y0);
  and_gate and_gate_h_u_cla32_and2070_y0(h_u_cla32_and2069_y0, h_u_cla32_and2068_y0, h_u_cla32_and2070_y0);
  and_gate and_gate_h_u_cla32_and2071_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2071_y0);
  and_gate and_gate_h_u_cla32_and2072_y0(h_u_cla32_and2071_y0, h_u_cla32_and2070_y0, h_u_cla32_and2072_y0);
  and_gate and_gate_h_u_cla32_and2073_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2073_y0);
  and_gate and_gate_h_u_cla32_and2074_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2074_y0);
  and_gate and_gate_h_u_cla32_and2075_y0(h_u_cla32_and2074_y0, h_u_cla32_and2073_y0, h_u_cla32_and2075_y0);
  and_gate and_gate_h_u_cla32_and2076_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2076_y0);
  and_gate and_gate_h_u_cla32_and2077_y0(h_u_cla32_and2076_y0, h_u_cla32_and2075_y0, h_u_cla32_and2077_y0);
  and_gate and_gate_h_u_cla32_and2078_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2078_y0);
  and_gate and_gate_h_u_cla32_and2079_y0(h_u_cla32_and2078_y0, h_u_cla32_and2077_y0, h_u_cla32_and2079_y0);
  and_gate and_gate_h_u_cla32_and2080_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2080_y0);
  and_gate and_gate_h_u_cla32_and2081_y0(h_u_cla32_and2080_y0, h_u_cla32_and2079_y0, h_u_cla32_and2081_y0);
  and_gate and_gate_h_u_cla32_and2082_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2082_y0);
  and_gate and_gate_h_u_cla32_and2083_y0(h_u_cla32_and2082_y0, h_u_cla32_and2081_y0, h_u_cla32_and2083_y0);
  and_gate and_gate_h_u_cla32_and2084_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2084_y0);
  and_gate and_gate_h_u_cla32_and2085_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2085_y0);
  and_gate and_gate_h_u_cla32_and2086_y0(h_u_cla32_and2085_y0, h_u_cla32_and2084_y0, h_u_cla32_and2086_y0);
  and_gate and_gate_h_u_cla32_and2087_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2087_y0);
  and_gate and_gate_h_u_cla32_and2088_y0(h_u_cla32_and2087_y0, h_u_cla32_and2086_y0, h_u_cla32_and2088_y0);
  and_gate and_gate_h_u_cla32_and2089_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2089_y0);
  and_gate and_gate_h_u_cla32_and2090_y0(h_u_cla32_and2089_y0, h_u_cla32_and2088_y0, h_u_cla32_and2090_y0);
  and_gate and_gate_h_u_cla32_and2091_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2091_y0);
  and_gate and_gate_h_u_cla32_and2092_y0(h_u_cla32_and2091_y0, h_u_cla32_and2090_y0, h_u_cla32_and2092_y0);
  and_gate and_gate_h_u_cla32_and2093_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2093_y0);
  and_gate and_gate_h_u_cla32_and2094_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2094_y0);
  and_gate and_gate_h_u_cla32_and2095_y0(h_u_cla32_and2094_y0, h_u_cla32_and2093_y0, h_u_cla32_and2095_y0);
  and_gate and_gate_h_u_cla32_and2096_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2096_y0);
  and_gate and_gate_h_u_cla32_and2097_y0(h_u_cla32_and2096_y0, h_u_cla32_and2095_y0, h_u_cla32_and2097_y0);
  and_gate and_gate_h_u_cla32_and2098_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2098_y0);
  and_gate and_gate_h_u_cla32_and2099_y0(h_u_cla32_and2098_y0, h_u_cla32_and2097_y0, h_u_cla32_and2099_y0);
  and_gate and_gate_h_u_cla32_and2100_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2100_y0);
  and_gate and_gate_h_u_cla32_and2101_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2101_y0);
  and_gate and_gate_h_u_cla32_and2102_y0(h_u_cla32_and2101_y0, h_u_cla32_and2100_y0, h_u_cla32_and2102_y0);
  and_gate and_gate_h_u_cla32_and2103_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2103_y0);
  and_gate and_gate_h_u_cla32_and2104_y0(h_u_cla32_and2103_y0, h_u_cla32_and2102_y0, h_u_cla32_and2104_y0);
  and_gate and_gate_h_u_cla32_and2105_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2105_y0);
  and_gate and_gate_h_u_cla32_and2106_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2106_y0);
  and_gate and_gate_h_u_cla32_and2107_y0(h_u_cla32_and2106_y0, h_u_cla32_and2105_y0, h_u_cla32_and2107_y0);
  and_gate and_gate_h_u_cla32_and2108_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and2108_y0);
  or_gate or_gate_h_u_cla32_or153_y0(h_u_cla32_and2108_y0, h_u_cla32_and1819_y0, h_u_cla32_or153_y0);
  or_gate or_gate_h_u_cla32_or154_y0(h_u_cla32_or153_y0, h_u_cla32_and1852_y0, h_u_cla32_or154_y0);
  or_gate or_gate_h_u_cla32_or155_y0(h_u_cla32_or154_y0, h_u_cla32_and1883_y0, h_u_cla32_or155_y0);
  or_gate or_gate_h_u_cla32_or156_y0(h_u_cla32_or155_y0, h_u_cla32_and1912_y0, h_u_cla32_or156_y0);
  or_gate or_gate_h_u_cla32_or157_y0(h_u_cla32_or156_y0, h_u_cla32_and1939_y0, h_u_cla32_or157_y0);
  or_gate or_gate_h_u_cla32_or158_y0(h_u_cla32_or157_y0, h_u_cla32_and1964_y0, h_u_cla32_or158_y0);
  or_gate or_gate_h_u_cla32_or159_y0(h_u_cla32_or158_y0, h_u_cla32_and1987_y0, h_u_cla32_or159_y0);
  or_gate or_gate_h_u_cla32_or160_y0(h_u_cla32_or159_y0, h_u_cla32_and2008_y0, h_u_cla32_or160_y0);
  or_gate or_gate_h_u_cla32_or161_y0(h_u_cla32_or160_y0, h_u_cla32_and2027_y0, h_u_cla32_or161_y0);
  or_gate or_gate_h_u_cla32_or162_y0(h_u_cla32_or161_y0, h_u_cla32_and2044_y0, h_u_cla32_or162_y0);
  or_gate or_gate_h_u_cla32_or163_y0(h_u_cla32_or162_y0, h_u_cla32_and2059_y0, h_u_cla32_or163_y0);
  or_gate or_gate_h_u_cla32_or164_y0(h_u_cla32_or163_y0, h_u_cla32_and2072_y0, h_u_cla32_or164_y0);
  or_gate or_gate_h_u_cla32_or165_y0(h_u_cla32_or164_y0, h_u_cla32_and2083_y0, h_u_cla32_or165_y0);
  or_gate or_gate_h_u_cla32_or166_y0(h_u_cla32_or165_y0, h_u_cla32_and2092_y0, h_u_cla32_or166_y0);
  or_gate or_gate_h_u_cla32_or167_y0(h_u_cla32_or166_y0, h_u_cla32_and2099_y0, h_u_cla32_or167_y0);
  or_gate or_gate_h_u_cla32_or168_y0(h_u_cla32_or167_y0, h_u_cla32_and2104_y0, h_u_cla32_or168_y0);
  or_gate or_gate_h_u_cla32_or169_y0(h_u_cla32_or168_y0, h_u_cla32_and2107_y0, h_u_cla32_or169_y0);
  or_gate or_gate_h_u_cla32_or170_y0(h_u_cla32_pg_logic17_y1, h_u_cla32_or169_y0, h_u_cla32_or170_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic18_y0(a_18, b_18, h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_pg_logic18_y2);
  xor_gate xor_gate_h_u_cla32_xor18_y0(h_u_cla32_pg_logic18_y2, h_u_cla32_or170_y0, h_u_cla32_xor18_y0);
  and_gate and_gate_h_u_cla32_and2109_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and2109_y0);
  and_gate and_gate_h_u_cla32_and2110_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and2110_y0);
  and_gate and_gate_h_u_cla32_and2111_y0(h_u_cla32_and2110_y0, h_u_cla32_and2109_y0, h_u_cla32_and2111_y0);
  and_gate and_gate_h_u_cla32_and2112_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and2112_y0);
  and_gate and_gate_h_u_cla32_and2113_y0(h_u_cla32_and2112_y0, h_u_cla32_and2111_y0, h_u_cla32_and2113_y0);
  and_gate and_gate_h_u_cla32_and2114_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and2114_y0);
  and_gate and_gate_h_u_cla32_and2115_y0(h_u_cla32_and2114_y0, h_u_cla32_and2113_y0, h_u_cla32_and2115_y0);
  and_gate and_gate_h_u_cla32_and2116_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and2116_y0);
  and_gate and_gate_h_u_cla32_and2117_y0(h_u_cla32_and2116_y0, h_u_cla32_and2115_y0, h_u_cla32_and2117_y0);
  and_gate and_gate_h_u_cla32_and2118_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and2118_y0);
  and_gate and_gate_h_u_cla32_and2119_y0(h_u_cla32_and2118_y0, h_u_cla32_and2117_y0, h_u_cla32_and2119_y0);
  and_gate and_gate_h_u_cla32_and2120_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and2120_y0);
  and_gate and_gate_h_u_cla32_and2121_y0(h_u_cla32_and2120_y0, h_u_cla32_and2119_y0, h_u_cla32_and2121_y0);
  and_gate and_gate_h_u_cla32_and2122_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and2122_y0);
  and_gate and_gate_h_u_cla32_and2123_y0(h_u_cla32_and2122_y0, h_u_cla32_and2121_y0, h_u_cla32_and2123_y0);
  and_gate and_gate_h_u_cla32_and2124_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and2124_y0);
  and_gate and_gate_h_u_cla32_and2125_y0(h_u_cla32_and2124_y0, h_u_cla32_and2123_y0, h_u_cla32_and2125_y0);
  and_gate and_gate_h_u_cla32_and2126_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and2126_y0);
  and_gate and_gate_h_u_cla32_and2127_y0(h_u_cla32_and2126_y0, h_u_cla32_and2125_y0, h_u_cla32_and2127_y0);
  and_gate and_gate_h_u_cla32_and2128_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and2128_y0);
  and_gate and_gate_h_u_cla32_and2129_y0(h_u_cla32_and2128_y0, h_u_cla32_and2127_y0, h_u_cla32_and2129_y0);
  and_gate and_gate_h_u_cla32_and2130_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and2130_y0);
  and_gate and_gate_h_u_cla32_and2131_y0(h_u_cla32_and2130_y0, h_u_cla32_and2129_y0, h_u_cla32_and2131_y0);
  and_gate and_gate_h_u_cla32_and2132_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and2132_y0);
  and_gate and_gate_h_u_cla32_and2133_y0(h_u_cla32_and2132_y0, h_u_cla32_and2131_y0, h_u_cla32_and2133_y0);
  and_gate and_gate_h_u_cla32_and2134_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and2134_y0);
  and_gate and_gate_h_u_cla32_and2135_y0(h_u_cla32_and2134_y0, h_u_cla32_and2133_y0, h_u_cla32_and2135_y0);
  and_gate and_gate_h_u_cla32_and2136_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and2136_y0);
  and_gate and_gate_h_u_cla32_and2137_y0(h_u_cla32_and2136_y0, h_u_cla32_and2135_y0, h_u_cla32_and2137_y0);
  and_gate and_gate_h_u_cla32_and2138_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and2138_y0);
  and_gate and_gate_h_u_cla32_and2139_y0(h_u_cla32_and2138_y0, h_u_cla32_and2137_y0, h_u_cla32_and2139_y0);
  and_gate and_gate_h_u_cla32_and2140_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and2140_y0);
  and_gate and_gate_h_u_cla32_and2141_y0(h_u_cla32_and2140_y0, h_u_cla32_and2139_y0, h_u_cla32_and2141_y0);
  and_gate and_gate_h_u_cla32_and2142_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and2142_y0);
  and_gate and_gate_h_u_cla32_and2143_y0(h_u_cla32_and2142_y0, h_u_cla32_and2141_y0, h_u_cla32_and2143_y0);
  and_gate and_gate_h_u_cla32_and2144_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and2144_y0);
  and_gate and_gate_h_u_cla32_and2145_y0(h_u_cla32_and2144_y0, h_u_cla32_and2143_y0, h_u_cla32_and2145_y0);
  and_gate and_gate_h_u_cla32_and2146_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2146_y0);
  and_gate and_gate_h_u_cla32_and2147_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2147_y0);
  and_gate and_gate_h_u_cla32_and2148_y0(h_u_cla32_and2147_y0, h_u_cla32_and2146_y0, h_u_cla32_and2148_y0);
  and_gate and_gate_h_u_cla32_and2149_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2149_y0);
  and_gate and_gate_h_u_cla32_and2150_y0(h_u_cla32_and2149_y0, h_u_cla32_and2148_y0, h_u_cla32_and2150_y0);
  and_gate and_gate_h_u_cla32_and2151_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2151_y0);
  and_gate and_gate_h_u_cla32_and2152_y0(h_u_cla32_and2151_y0, h_u_cla32_and2150_y0, h_u_cla32_and2152_y0);
  and_gate and_gate_h_u_cla32_and2153_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2153_y0);
  and_gate and_gate_h_u_cla32_and2154_y0(h_u_cla32_and2153_y0, h_u_cla32_and2152_y0, h_u_cla32_and2154_y0);
  and_gate and_gate_h_u_cla32_and2155_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2155_y0);
  and_gate and_gate_h_u_cla32_and2156_y0(h_u_cla32_and2155_y0, h_u_cla32_and2154_y0, h_u_cla32_and2156_y0);
  and_gate and_gate_h_u_cla32_and2157_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2157_y0);
  and_gate and_gate_h_u_cla32_and2158_y0(h_u_cla32_and2157_y0, h_u_cla32_and2156_y0, h_u_cla32_and2158_y0);
  and_gate and_gate_h_u_cla32_and2159_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2159_y0);
  and_gate and_gate_h_u_cla32_and2160_y0(h_u_cla32_and2159_y0, h_u_cla32_and2158_y0, h_u_cla32_and2160_y0);
  and_gate and_gate_h_u_cla32_and2161_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2161_y0);
  and_gate and_gate_h_u_cla32_and2162_y0(h_u_cla32_and2161_y0, h_u_cla32_and2160_y0, h_u_cla32_and2162_y0);
  and_gate and_gate_h_u_cla32_and2163_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2163_y0);
  and_gate and_gate_h_u_cla32_and2164_y0(h_u_cla32_and2163_y0, h_u_cla32_and2162_y0, h_u_cla32_and2164_y0);
  and_gate and_gate_h_u_cla32_and2165_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2165_y0);
  and_gate and_gate_h_u_cla32_and2166_y0(h_u_cla32_and2165_y0, h_u_cla32_and2164_y0, h_u_cla32_and2166_y0);
  and_gate and_gate_h_u_cla32_and2167_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2167_y0);
  and_gate and_gate_h_u_cla32_and2168_y0(h_u_cla32_and2167_y0, h_u_cla32_and2166_y0, h_u_cla32_and2168_y0);
  and_gate and_gate_h_u_cla32_and2169_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2169_y0);
  and_gate and_gate_h_u_cla32_and2170_y0(h_u_cla32_and2169_y0, h_u_cla32_and2168_y0, h_u_cla32_and2170_y0);
  and_gate and_gate_h_u_cla32_and2171_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2171_y0);
  and_gate and_gate_h_u_cla32_and2172_y0(h_u_cla32_and2171_y0, h_u_cla32_and2170_y0, h_u_cla32_and2172_y0);
  and_gate and_gate_h_u_cla32_and2173_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2173_y0);
  and_gate and_gate_h_u_cla32_and2174_y0(h_u_cla32_and2173_y0, h_u_cla32_and2172_y0, h_u_cla32_and2174_y0);
  and_gate and_gate_h_u_cla32_and2175_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2175_y0);
  and_gate and_gate_h_u_cla32_and2176_y0(h_u_cla32_and2175_y0, h_u_cla32_and2174_y0, h_u_cla32_and2176_y0);
  and_gate and_gate_h_u_cla32_and2177_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2177_y0);
  and_gate and_gate_h_u_cla32_and2178_y0(h_u_cla32_and2177_y0, h_u_cla32_and2176_y0, h_u_cla32_and2178_y0);
  and_gate and_gate_h_u_cla32_and2179_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2179_y0);
  and_gate and_gate_h_u_cla32_and2180_y0(h_u_cla32_and2179_y0, h_u_cla32_and2178_y0, h_u_cla32_and2180_y0);
  and_gate and_gate_h_u_cla32_and2181_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2181_y0);
  and_gate and_gate_h_u_cla32_and2182_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2182_y0);
  and_gate and_gate_h_u_cla32_and2183_y0(h_u_cla32_and2182_y0, h_u_cla32_and2181_y0, h_u_cla32_and2183_y0);
  and_gate and_gate_h_u_cla32_and2184_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2184_y0);
  and_gate and_gate_h_u_cla32_and2185_y0(h_u_cla32_and2184_y0, h_u_cla32_and2183_y0, h_u_cla32_and2185_y0);
  and_gate and_gate_h_u_cla32_and2186_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2186_y0);
  and_gate and_gate_h_u_cla32_and2187_y0(h_u_cla32_and2186_y0, h_u_cla32_and2185_y0, h_u_cla32_and2187_y0);
  and_gate and_gate_h_u_cla32_and2188_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2188_y0);
  and_gate and_gate_h_u_cla32_and2189_y0(h_u_cla32_and2188_y0, h_u_cla32_and2187_y0, h_u_cla32_and2189_y0);
  and_gate and_gate_h_u_cla32_and2190_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2190_y0);
  and_gate and_gate_h_u_cla32_and2191_y0(h_u_cla32_and2190_y0, h_u_cla32_and2189_y0, h_u_cla32_and2191_y0);
  and_gate and_gate_h_u_cla32_and2192_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2192_y0);
  and_gate and_gate_h_u_cla32_and2193_y0(h_u_cla32_and2192_y0, h_u_cla32_and2191_y0, h_u_cla32_and2193_y0);
  and_gate and_gate_h_u_cla32_and2194_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2194_y0);
  and_gate and_gate_h_u_cla32_and2195_y0(h_u_cla32_and2194_y0, h_u_cla32_and2193_y0, h_u_cla32_and2195_y0);
  and_gate and_gate_h_u_cla32_and2196_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2196_y0);
  and_gate and_gate_h_u_cla32_and2197_y0(h_u_cla32_and2196_y0, h_u_cla32_and2195_y0, h_u_cla32_and2197_y0);
  and_gate and_gate_h_u_cla32_and2198_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2198_y0);
  and_gate and_gate_h_u_cla32_and2199_y0(h_u_cla32_and2198_y0, h_u_cla32_and2197_y0, h_u_cla32_and2199_y0);
  and_gate and_gate_h_u_cla32_and2200_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2200_y0);
  and_gate and_gate_h_u_cla32_and2201_y0(h_u_cla32_and2200_y0, h_u_cla32_and2199_y0, h_u_cla32_and2201_y0);
  and_gate and_gate_h_u_cla32_and2202_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2202_y0);
  and_gate and_gate_h_u_cla32_and2203_y0(h_u_cla32_and2202_y0, h_u_cla32_and2201_y0, h_u_cla32_and2203_y0);
  and_gate and_gate_h_u_cla32_and2204_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2204_y0);
  and_gate and_gate_h_u_cla32_and2205_y0(h_u_cla32_and2204_y0, h_u_cla32_and2203_y0, h_u_cla32_and2205_y0);
  and_gate and_gate_h_u_cla32_and2206_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2206_y0);
  and_gate and_gate_h_u_cla32_and2207_y0(h_u_cla32_and2206_y0, h_u_cla32_and2205_y0, h_u_cla32_and2207_y0);
  and_gate and_gate_h_u_cla32_and2208_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2208_y0);
  and_gate and_gate_h_u_cla32_and2209_y0(h_u_cla32_and2208_y0, h_u_cla32_and2207_y0, h_u_cla32_and2209_y0);
  and_gate and_gate_h_u_cla32_and2210_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2210_y0);
  and_gate and_gate_h_u_cla32_and2211_y0(h_u_cla32_and2210_y0, h_u_cla32_and2209_y0, h_u_cla32_and2211_y0);
  and_gate and_gate_h_u_cla32_and2212_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2212_y0);
  and_gate and_gate_h_u_cla32_and2213_y0(h_u_cla32_and2212_y0, h_u_cla32_and2211_y0, h_u_cla32_and2213_y0);
  and_gate and_gate_h_u_cla32_and2214_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2214_y0);
  and_gate and_gate_h_u_cla32_and2215_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2215_y0);
  and_gate and_gate_h_u_cla32_and2216_y0(h_u_cla32_and2215_y0, h_u_cla32_and2214_y0, h_u_cla32_and2216_y0);
  and_gate and_gate_h_u_cla32_and2217_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2217_y0);
  and_gate and_gate_h_u_cla32_and2218_y0(h_u_cla32_and2217_y0, h_u_cla32_and2216_y0, h_u_cla32_and2218_y0);
  and_gate and_gate_h_u_cla32_and2219_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2219_y0);
  and_gate and_gate_h_u_cla32_and2220_y0(h_u_cla32_and2219_y0, h_u_cla32_and2218_y0, h_u_cla32_and2220_y0);
  and_gate and_gate_h_u_cla32_and2221_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2221_y0);
  and_gate and_gate_h_u_cla32_and2222_y0(h_u_cla32_and2221_y0, h_u_cla32_and2220_y0, h_u_cla32_and2222_y0);
  and_gate and_gate_h_u_cla32_and2223_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2223_y0);
  and_gate and_gate_h_u_cla32_and2224_y0(h_u_cla32_and2223_y0, h_u_cla32_and2222_y0, h_u_cla32_and2224_y0);
  and_gate and_gate_h_u_cla32_and2225_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2225_y0);
  and_gate and_gate_h_u_cla32_and2226_y0(h_u_cla32_and2225_y0, h_u_cla32_and2224_y0, h_u_cla32_and2226_y0);
  and_gate and_gate_h_u_cla32_and2227_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2227_y0);
  and_gate and_gate_h_u_cla32_and2228_y0(h_u_cla32_and2227_y0, h_u_cla32_and2226_y0, h_u_cla32_and2228_y0);
  and_gate and_gate_h_u_cla32_and2229_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2229_y0);
  and_gate and_gate_h_u_cla32_and2230_y0(h_u_cla32_and2229_y0, h_u_cla32_and2228_y0, h_u_cla32_and2230_y0);
  and_gate and_gate_h_u_cla32_and2231_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2231_y0);
  and_gate and_gate_h_u_cla32_and2232_y0(h_u_cla32_and2231_y0, h_u_cla32_and2230_y0, h_u_cla32_and2232_y0);
  and_gate and_gate_h_u_cla32_and2233_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2233_y0);
  and_gate and_gate_h_u_cla32_and2234_y0(h_u_cla32_and2233_y0, h_u_cla32_and2232_y0, h_u_cla32_and2234_y0);
  and_gate and_gate_h_u_cla32_and2235_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2235_y0);
  and_gate and_gate_h_u_cla32_and2236_y0(h_u_cla32_and2235_y0, h_u_cla32_and2234_y0, h_u_cla32_and2236_y0);
  and_gate and_gate_h_u_cla32_and2237_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2237_y0);
  and_gate and_gate_h_u_cla32_and2238_y0(h_u_cla32_and2237_y0, h_u_cla32_and2236_y0, h_u_cla32_and2238_y0);
  and_gate and_gate_h_u_cla32_and2239_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2239_y0);
  and_gate and_gate_h_u_cla32_and2240_y0(h_u_cla32_and2239_y0, h_u_cla32_and2238_y0, h_u_cla32_and2240_y0);
  and_gate and_gate_h_u_cla32_and2241_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2241_y0);
  and_gate and_gate_h_u_cla32_and2242_y0(h_u_cla32_and2241_y0, h_u_cla32_and2240_y0, h_u_cla32_and2242_y0);
  and_gate and_gate_h_u_cla32_and2243_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2243_y0);
  and_gate and_gate_h_u_cla32_and2244_y0(h_u_cla32_and2243_y0, h_u_cla32_and2242_y0, h_u_cla32_and2244_y0);
  and_gate and_gate_h_u_cla32_and2245_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2245_y0);
  and_gate and_gate_h_u_cla32_and2246_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2246_y0);
  and_gate and_gate_h_u_cla32_and2247_y0(h_u_cla32_and2246_y0, h_u_cla32_and2245_y0, h_u_cla32_and2247_y0);
  and_gate and_gate_h_u_cla32_and2248_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2248_y0);
  and_gate and_gate_h_u_cla32_and2249_y0(h_u_cla32_and2248_y0, h_u_cla32_and2247_y0, h_u_cla32_and2249_y0);
  and_gate and_gate_h_u_cla32_and2250_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2250_y0);
  and_gate and_gate_h_u_cla32_and2251_y0(h_u_cla32_and2250_y0, h_u_cla32_and2249_y0, h_u_cla32_and2251_y0);
  and_gate and_gate_h_u_cla32_and2252_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2252_y0);
  and_gate and_gate_h_u_cla32_and2253_y0(h_u_cla32_and2252_y0, h_u_cla32_and2251_y0, h_u_cla32_and2253_y0);
  and_gate and_gate_h_u_cla32_and2254_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2254_y0);
  and_gate and_gate_h_u_cla32_and2255_y0(h_u_cla32_and2254_y0, h_u_cla32_and2253_y0, h_u_cla32_and2255_y0);
  and_gate and_gate_h_u_cla32_and2256_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2256_y0);
  and_gate and_gate_h_u_cla32_and2257_y0(h_u_cla32_and2256_y0, h_u_cla32_and2255_y0, h_u_cla32_and2257_y0);
  and_gate and_gate_h_u_cla32_and2258_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2258_y0);
  and_gate and_gate_h_u_cla32_and2259_y0(h_u_cla32_and2258_y0, h_u_cla32_and2257_y0, h_u_cla32_and2259_y0);
  and_gate and_gate_h_u_cla32_and2260_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2260_y0);
  and_gate and_gate_h_u_cla32_and2261_y0(h_u_cla32_and2260_y0, h_u_cla32_and2259_y0, h_u_cla32_and2261_y0);
  and_gate and_gate_h_u_cla32_and2262_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2262_y0);
  and_gate and_gate_h_u_cla32_and2263_y0(h_u_cla32_and2262_y0, h_u_cla32_and2261_y0, h_u_cla32_and2263_y0);
  and_gate and_gate_h_u_cla32_and2264_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2264_y0);
  and_gate and_gate_h_u_cla32_and2265_y0(h_u_cla32_and2264_y0, h_u_cla32_and2263_y0, h_u_cla32_and2265_y0);
  and_gate and_gate_h_u_cla32_and2266_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2266_y0);
  and_gate and_gate_h_u_cla32_and2267_y0(h_u_cla32_and2266_y0, h_u_cla32_and2265_y0, h_u_cla32_and2267_y0);
  and_gate and_gate_h_u_cla32_and2268_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2268_y0);
  and_gate and_gate_h_u_cla32_and2269_y0(h_u_cla32_and2268_y0, h_u_cla32_and2267_y0, h_u_cla32_and2269_y0);
  and_gate and_gate_h_u_cla32_and2270_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2270_y0);
  and_gate and_gate_h_u_cla32_and2271_y0(h_u_cla32_and2270_y0, h_u_cla32_and2269_y0, h_u_cla32_and2271_y0);
  and_gate and_gate_h_u_cla32_and2272_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2272_y0);
  and_gate and_gate_h_u_cla32_and2273_y0(h_u_cla32_and2272_y0, h_u_cla32_and2271_y0, h_u_cla32_and2273_y0);
  and_gate and_gate_h_u_cla32_and2274_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2274_y0);
  and_gate and_gate_h_u_cla32_and2275_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2275_y0);
  and_gate and_gate_h_u_cla32_and2276_y0(h_u_cla32_and2275_y0, h_u_cla32_and2274_y0, h_u_cla32_and2276_y0);
  and_gate and_gate_h_u_cla32_and2277_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2277_y0);
  and_gate and_gate_h_u_cla32_and2278_y0(h_u_cla32_and2277_y0, h_u_cla32_and2276_y0, h_u_cla32_and2278_y0);
  and_gate and_gate_h_u_cla32_and2279_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2279_y0);
  and_gate and_gate_h_u_cla32_and2280_y0(h_u_cla32_and2279_y0, h_u_cla32_and2278_y0, h_u_cla32_and2280_y0);
  and_gate and_gate_h_u_cla32_and2281_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2281_y0);
  and_gate and_gate_h_u_cla32_and2282_y0(h_u_cla32_and2281_y0, h_u_cla32_and2280_y0, h_u_cla32_and2282_y0);
  and_gate and_gate_h_u_cla32_and2283_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2283_y0);
  and_gate and_gate_h_u_cla32_and2284_y0(h_u_cla32_and2283_y0, h_u_cla32_and2282_y0, h_u_cla32_and2284_y0);
  and_gate and_gate_h_u_cla32_and2285_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2285_y0);
  and_gate and_gate_h_u_cla32_and2286_y0(h_u_cla32_and2285_y0, h_u_cla32_and2284_y0, h_u_cla32_and2286_y0);
  and_gate and_gate_h_u_cla32_and2287_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2287_y0);
  and_gate and_gate_h_u_cla32_and2288_y0(h_u_cla32_and2287_y0, h_u_cla32_and2286_y0, h_u_cla32_and2288_y0);
  and_gate and_gate_h_u_cla32_and2289_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2289_y0);
  and_gate and_gate_h_u_cla32_and2290_y0(h_u_cla32_and2289_y0, h_u_cla32_and2288_y0, h_u_cla32_and2290_y0);
  and_gate and_gate_h_u_cla32_and2291_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2291_y0);
  and_gate and_gate_h_u_cla32_and2292_y0(h_u_cla32_and2291_y0, h_u_cla32_and2290_y0, h_u_cla32_and2292_y0);
  and_gate and_gate_h_u_cla32_and2293_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2293_y0);
  and_gate and_gate_h_u_cla32_and2294_y0(h_u_cla32_and2293_y0, h_u_cla32_and2292_y0, h_u_cla32_and2294_y0);
  and_gate and_gate_h_u_cla32_and2295_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2295_y0);
  and_gate and_gate_h_u_cla32_and2296_y0(h_u_cla32_and2295_y0, h_u_cla32_and2294_y0, h_u_cla32_and2296_y0);
  and_gate and_gate_h_u_cla32_and2297_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2297_y0);
  and_gate and_gate_h_u_cla32_and2298_y0(h_u_cla32_and2297_y0, h_u_cla32_and2296_y0, h_u_cla32_and2298_y0);
  and_gate and_gate_h_u_cla32_and2299_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2299_y0);
  and_gate and_gate_h_u_cla32_and2300_y0(h_u_cla32_and2299_y0, h_u_cla32_and2298_y0, h_u_cla32_and2300_y0);
  and_gate and_gate_h_u_cla32_and2301_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2301_y0);
  and_gate and_gate_h_u_cla32_and2302_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2302_y0);
  and_gate and_gate_h_u_cla32_and2303_y0(h_u_cla32_and2302_y0, h_u_cla32_and2301_y0, h_u_cla32_and2303_y0);
  and_gate and_gate_h_u_cla32_and2304_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2304_y0);
  and_gate and_gate_h_u_cla32_and2305_y0(h_u_cla32_and2304_y0, h_u_cla32_and2303_y0, h_u_cla32_and2305_y0);
  and_gate and_gate_h_u_cla32_and2306_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2306_y0);
  and_gate and_gate_h_u_cla32_and2307_y0(h_u_cla32_and2306_y0, h_u_cla32_and2305_y0, h_u_cla32_and2307_y0);
  and_gate and_gate_h_u_cla32_and2308_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2308_y0);
  and_gate and_gate_h_u_cla32_and2309_y0(h_u_cla32_and2308_y0, h_u_cla32_and2307_y0, h_u_cla32_and2309_y0);
  and_gate and_gate_h_u_cla32_and2310_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2310_y0);
  and_gate and_gate_h_u_cla32_and2311_y0(h_u_cla32_and2310_y0, h_u_cla32_and2309_y0, h_u_cla32_and2311_y0);
  and_gate and_gate_h_u_cla32_and2312_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2312_y0);
  and_gate and_gate_h_u_cla32_and2313_y0(h_u_cla32_and2312_y0, h_u_cla32_and2311_y0, h_u_cla32_and2313_y0);
  and_gate and_gate_h_u_cla32_and2314_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2314_y0);
  and_gate and_gate_h_u_cla32_and2315_y0(h_u_cla32_and2314_y0, h_u_cla32_and2313_y0, h_u_cla32_and2315_y0);
  and_gate and_gate_h_u_cla32_and2316_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2316_y0);
  and_gate and_gate_h_u_cla32_and2317_y0(h_u_cla32_and2316_y0, h_u_cla32_and2315_y0, h_u_cla32_and2317_y0);
  and_gate and_gate_h_u_cla32_and2318_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2318_y0);
  and_gate and_gate_h_u_cla32_and2319_y0(h_u_cla32_and2318_y0, h_u_cla32_and2317_y0, h_u_cla32_and2319_y0);
  and_gate and_gate_h_u_cla32_and2320_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2320_y0);
  and_gate and_gate_h_u_cla32_and2321_y0(h_u_cla32_and2320_y0, h_u_cla32_and2319_y0, h_u_cla32_and2321_y0);
  and_gate and_gate_h_u_cla32_and2322_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2322_y0);
  and_gate and_gate_h_u_cla32_and2323_y0(h_u_cla32_and2322_y0, h_u_cla32_and2321_y0, h_u_cla32_and2323_y0);
  and_gate and_gate_h_u_cla32_and2324_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2324_y0);
  and_gate and_gate_h_u_cla32_and2325_y0(h_u_cla32_and2324_y0, h_u_cla32_and2323_y0, h_u_cla32_and2325_y0);
  and_gate and_gate_h_u_cla32_and2326_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2326_y0);
  and_gate and_gate_h_u_cla32_and2327_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2327_y0);
  and_gate and_gate_h_u_cla32_and2328_y0(h_u_cla32_and2327_y0, h_u_cla32_and2326_y0, h_u_cla32_and2328_y0);
  and_gate and_gate_h_u_cla32_and2329_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2329_y0);
  and_gate and_gate_h_u_cla32_and2330_y0(h_u_cla32_and2329_y0, h_u_cla32_and2328_y0, h_u_cla32_and2330_y0);
  and_gate and_gate_h_u_cla32_and2331_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2331_y0);
  and_gate and_gate_h_u_cla32_and2332_y0(h_u_cla32_and2331_y0, h_u_cla32_and2330_y0, h_u_cla32_and2332_y0);
  and_gate and_gate_h_u_cla32_and2333_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2333_y0);
  and_gate and_gate_h_u_cla32_and2334_y0(h_u_cla32_and2333_y0, h_u_cla32_and2332_y0, h_u_cla32_and2334_y0);
  and_gate and_gate_h_u_cla32_and2335_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2335_y0);
  and_gate and_gate_h_u_cla32_and2336_y0(h_u_cla32_and2335_y0, h_u_cla32_and2334_y0, h_u_cla32_and2336_y0);
  and_gate and_gate_h_u_cla32_and2337_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2337_y0);
  and_gate and_gate_h_u_cla32_and2338_y0(h_u_cla32_and2337_y0, h_u_cla32_and2336_y0, h_u_cla32_and2338_y0);
  and_gate and_gate_h_u_cla32_and2339_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2339_y0);
  and_gate and_gate_h_u_cla32_and2340_y0(h_u_cla32_and2339_y0, h_u_cla32_and2338_y0, h_u_cla32_and2340_y0);
  and_gate and_gate_h_u_cla32_and2341_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2341_y0);
  and_gate and_gate_h_u_cla32_and2342_y0(h_u_cla32_and2341_y0, h_u_cla32_and2340_y0, h_u_cla32_and2342_y0);
  and_gate and_gate_h_u_cla32_and2343_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2343_y0);
  and_gate and_gate_h_u_cla32_and2344_y0(h_u_cla32_and2343_y0, h_u_cla32_and2342_y0, h_u_cla32_and2344_y0);
  and_gate and_gate_h_u_cla32_and2345_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2345_y0);
  and_gate and_gate_h_u_cla32_and2346_y0(h_u_cla32_and2345_y0, h_u_cla32_and2344_y0, h_u_cla32_and2346_y0);
  and_gate and_gate_h_u_cla32_and2347_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2347_y0);
  and_gate and_gate_h_u_cla32_and2348_y0(h_u_cla32_and2347_y0, h_u_cla32_and2346_y0, h_u_cla32_and2348_y0);
  and_gate and_gate_h_u_cla32_and2349_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2349_y0);
  and_gate and_gate_h_u_cla32_and2350_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2350_y0);
  and_gate and_gate_h_u_cla32_and2351_y0(h_u_cla32_and2350_y0, h_u_cla32_and2349_y0, h_u_cla32_and2351_y0);
  and_gate and_gate_h_u_cla32_and2352_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2352_y0);
  and_gate and_gate_h_u_cla32_and2353_y0(h_u_cla32_and2352_y0, h_u_cla32_and2351_y0, h_u_cla32_and2353_y0);
  and_gate and_gate_h_u_cla32_and2354_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2354_y0);
  and_gate and_gate_h_u_cla32_and2355_y0(h_u_cla32_and2354_y0, h_u_cla32_and2353_y0, h_u_cla32_and2355_y0);
  and_gate and_gate_h_u_cla32_and2356_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2356_y0);
  and_gate and_gate_h_u_cla32_and2357_y0(h_u_cla32_and2356_y0, h_u_cla32_and2355_y0, h_u_cla32_and2357_y0);
  and_gate and_gate_h_u_cla32_and2358_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2358_y0);
  and_gate and_gate_h_u_cla32_and2359_y0(h_u_cla32_and2358_y0, h_u_cla32_and2357_y0, h_u_cla32_and2359_y0);
  and_gate and_gate_h_u_cla32_and2360_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2360_y0);
  and_gate and_gate_h_u_cla32_and2361_y0(h_u_cla32_and2360_y0, h_u_cla32_and2359_y0, h_u_cla32_and2361_y0);
  and_gate and_gate_h_u_cla32_and2362_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2362_y0);
  and_gate and_gate_h_u_cla32_and2363_y0(h_u_cla32_and2362_y0, h_u_cla32_and2361_y0, h_u_cla32_and2363_y0);
  and_gate and_gate_h_u_cla32_and2364_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2364_y0);
  and_gate and_gate_h_u_cla32_and2365_y0(h_u_cla32_and2364_y0, h_u_cla32_and2363_y0, h_u_cla32_and2365_y0);
  and_gate and_gate_h_u_cla32_and2366_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2366_y0);
  and_gate and_gate_h_u_cla32_and2367_y0(h_u_cla32_and2366_y0, h_u_cla32_and2365_y0, h_u_cla32_and2367_y0);
  and_gate and_gate_h_u_cla32_and2368_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2368_y0);
  and_gate and_gate_h_u_cla32_and2369_y0(h_u_cla32_and2368_y0, h_u_cla32_and2367_y0, h_u_cla32_and2369_y0);
  and_gate and_gate_h_u_cla32_and2370_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2370_y0);
  and_gate and_gate_h_u_cla32_and2371_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2371_y0);
  and_gate and_gate_h_u_cla32_and2372_y0(h_u_cla32_and2371_y0, h_u_cla32_and2370_y0, h_u_cla32_and2372_y0);
  and_gate and_gate_h_u_cla32_and2373_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2373_y0);
  and_gate and_gate_h_u_cla32_and2374_y0(h_u_cla32_and2373_y0, h_u_cla32_and2372_y0, h_u_cla32_and2374_y0);
  and_gate and_gate_h_u_cla32_and2375_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2375_y0);
  and_gate and_gate_h_u_cla32_and2376_y0(h_u_cla32_and2375_y0, h_u_cla32_and2374_y0, h_u_cla32_and2376_y0);
  and_gate and_gate_h_u_cla32_and2377_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2377_y0);
  and_gate and_gate_h_u_cla32_and2378_y0(h_u_cla32_and2377_y0, h_u_cla32_and2376_y0, h_u_cla32_and2378_y0);
  and_gate and_gate_h_u_cla32_and2379_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2379_y0);
  and_gate and_gate_h_u_cla32_and2380_y0(h_u_cla32_and2379_y0, h_u_cla32_and2378_y0, h_u_cla32_and2380_y0);
  and_gate and_gate_h_u_cla32_and2381_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2381_y0);
  and_gate and_gate_h_u_cla32_and2382_y0(h_u_cla32_and2381_y0, h_u_cla32_and2380_y0, h_u_cla32_and2382_y0);
  and_gate and_gate_h_u_cla32_and2383_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2383_y0);
  and_gate and_gate_h_u_cla32_and2384_y0(h_u_cla32_and2383_y0, h_u_cla32_and2382_y0, h_u_cla32_and2384_y0);
  and_gate and_gate_h_u_cla32_and2385_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2385_y0);
  and_gate and_gate_h_u_cla32_and2386_y0(h_u_cla32_and2385_y0, h_u_cla32_and2384_y0, h_u_cla32_and2386_y0);
  and_gate and_gate_h_u_cla32_and2387_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2387_y0);
  and_gate and_gate_h_u_cla32_and2388_y0(h_u_cla32_and2387_y0, h_u_cla32_and2386_y0, h_u_cla32_and2388_y0);
  and_gate and_gate_h_u_cla32_and2389_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2389_y0);
  and_gate and_gate_h_u_cla32_and2390_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2390_y0);
  and_gate and_gate_h_u_cla32_and2391_y0(h_u_cla32_and2390_y0, h_u_cla32_and2389_y0, h_u_cla32_and2391_y0);
  and_gate and_gate_h_u_cla32_and2392_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2392_y0);
  and_gate and_gate_h_u_cla32_and2393_y0(h_u_cla32_and2392_y0, h_u_cla32_and2391_y0, h_u_cla32_and2393_y0);
  and_gate and_gate_h_u_cla32_and2394_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2394_y0);
  and_gate and_gate_h_u_cla32_and2395_y0(h_u_cla32_and2394_y0, h_u_cla32_and2393_y0, h_u_cla32_and2395_y0);
  and_gate and_gate_h_u_cla32_and2396_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2396_y0);
  and_gate and_gate_h_u_cla32_and2397_y0(h_u_cla32_and2396_y0, h_u_cla32_and2395_y0, h_u_cla32_and2397_y0);
  and_gate and_gate_h_u_cla32_and2398_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2398_y0);
  and_gate and_gate_h_u_cla32_and2399_y0(h_u_cla32_and2398_y0, h_u_cla32_and2397_y0, h_u_cla32_and2399_y0);
  and_gate and_gate_h_u_cla32_and2400_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2400_y0);
  and_gate and_gate_h_u_cla32_and2401_y0(h_u_cla32_and2400_y0, h_u_cla32_and2399_y0, h_u_cla32_and2401_y0);
  and_gate and_gate_h_u_cla32_and2402_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2402_y0);
  and_gate and_gate_h_u_cla32_and2403_y0(h_u_cla32_and2402_y0, h_u_cla32_and2401_y0, h_u_cla32_and2403_y0);
  and_gate and_gate_h_u_cla32_and2404_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2404_y0);
  and_gate and_gate_h_u_cla32_and2405_y0(h_u_cla32_and2404_y0, h_u_cla32_and2403_y0, h_u_cla32_and2405_y0);
  and_gate and_gate_h_u_cla32_and2406_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2406_y0);
  and_gate and_gate_h_u_cla32_and2407_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2407_y0);
  and_gate and_gate_h_u_cla32_and2408_y0(h_u_cla32_and2407_y0, h_u_cla32_and2406_y0, h_u_cla32_and2408_y0);
  and_gate and_gate_h_u_cla32_and2409_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2409_y0);
  and_gate and_gate_h_u_cla32_and2410_y0(h_u_cla32_and2409_y0, h_u_cla32_and2408_y0, h_u_cla32_and2410_y0);
  and_gate and_gate_h_u_cla32_and2411_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2411_y0);
  and_gate and_gate_h_u_cla32_and2412_y0(h_u_cla32_and2411_y0, h_u_cla32_and2410_y0, h_u_cla32_and2412_y0);
  and_gate and_gate_h_u_cla32_and2413_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2413_y0);
  and_gate and_gate_h_u_cla32_and2414_y0(h_u_cla32_and2413_y0, h_u_cla32_and2412_y0, h_u_cla32_and2414_y0);
  and_gate and_gate_h_u_cla32_and2415_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2415_y0);
  and_gate and_gate_h_u_cla32_and2416_y0(h_u_cla32_and2415_y0, h_u_cla32_and2414_y0, h_u_cla32_and2416_y0);
  and_gate and_gate_h_u_cla32_and2417_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2417_y0);
  and_gate and_gate_h_u_cla32_and2418_y0(h_u_cla32_and2417_y0, h_u_cla32_and2416_y0, h_u_cla32_and2418_y0);
  and_gate and_gate_h_u_cla32_and2419_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2419_y0);
  and_gate and_gate_h_u_cla32_and2420_y0(h_u_cla32_and2419_y0, h_u_cla32_and2418_y0, h_u_cla32_and2420_y0);
  and_gate and_gate_h_u_cla32_and2421_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2421_y0);
  and_gate and_gate_h_u_cla32_and2422_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2422_y0);
  and_gate and_gate_h_u_cla32_and2423_y0(h_u_cla32_and2422_y0, h_u_cla32_and2421_y0, h_u_cla32_and2423_y0);
  and_gate and_gate_h_u_cla32_and2424_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2424_y0);
  and_gate and_gate_h_u_cla32_and2425_y0(h_u_cla32_and2424_y0, h_u_cla32_and2423_y0, h_u_cla32_and2425_y0);
  and_gate and_gate_h_u_cla32_and2426_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2426_y0);
  and_gate and_gate_h_u_cla32_and2427_y0(h_u_cla32_and2426_y0, h_u_cla32_and2425_y0, h_u_cla32_and2427_y0);
  and_gate and_gate_h_u_cla32_and2428_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2428_y0);
  and_gate and_gate_h_u_cla32_and2429_y0(h_u_cla32_and2428_y0, h_u_cla32_and2427_y0, h_u_cla32_and2429_y0);
  and_gate and_gate_h_u_cla32_and2430_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2430_y0);
  and_gate and_gate_h_u_cla32_and2431_y0(h_u_cla32_and2430_y0, h_u_cla32_and2429_y0, h_u_cla32_and2431_y0);
  and_gate and_gate_h_u_cla32_and2432_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2432_y0);
  and_gate and_gate_h_u_cla32_and2433_y0(h_u_cla32_and2432_y0, h_u_cla32_and2431_y0, h_u_cla32_and2433_y0);
  and_gate and_gate_h_u_cla32_and2434_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2434_y0);
  and_gate and_gate_h_u_cla32_and2435_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2435_y0);
  and_gate and_gate_h_u_cla32_and2436_y0(h_u_cla32_and2435_y0, h_u_cla32_and2434_y0, h_u_cla32_and2436_y0);
  and_gate and_gate_h_u_cla32_and2437_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2437_y0);
  and_gate and_gate_h_u_cla32_and2438_y0(h_u_cla32_and2437_y0, h_u_cla32_and2436_y0, h_u_cla32_and2438_y0);
  and_gate and_gate_h_u_cla32_and2439_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2439_y0);
  and_gate and_gate_h_u_cla32_and2440_y0(h_u_cla32_and2439_y0, h_u_cla32_and2438_y0, h_u_cla32_and2440_y0);
  and_gate and_gate_h_u_cla32_and2441_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2441_y0);
  and_gate and_gate_h_u_cla32_and2442_y0(h_u_cla32_and2441_y0, h_u_cla32_and2440_y0, h_u_cla32_and2442_y0);
  and_gate and_gate_h_u_cla32_and2443_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2443_y0);
  and_gate and_gate_h_u_cla32_and2444_y0(h_u_cla32_and2443_y0, h_u_cla32_and2442_y0, h_u_cla32_and2444_y0);
  and_gate and_gate_h_u_cla32_and2445_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2445_y0);
  and_gate and_gate_h_u_cla32_and2446_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2446_y0);
  and_gate and_gate_h_u_cla32_and2447_y0(h_u_cla32_and2446_y0, h_u_cla32_and2445_y0, h_u_cla32_and2447_y0);
  and_gate and_gate_h_u_cla32_and2448_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2448_y0);
  and_gate and_gate_h_u_cla32_and2449_y0(h_u_cla32_and2448_y0, h_u_cla32_and2447_y0, h_u_cla32_and2449_y0);
  and_gate and_gate_h_u_cla32_and2450_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2450_y0);
  and_gate and_gate_h_u_cla32_and2451_y0(h_u_cla32_and2450_y0, h_u_cla32_and2449_y0, h_u_cla32_and2451_y0);
  and_gate and_gate_h_u_cla32_and2452_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2452_y0);
  and_gate and_gate_h_u_cla32_and2453_y0(h_u_cla32_and2452_y0, h_u_cla32_and2451_y0, h_u_cla32_and2453_y0);
  and_gate and_gate_h_u_cla32_and2454_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2454_y0);
  and_gate and_gate_h_u_cla32_and2455_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2455_y0);
  and_gate and_gate_h_u_cla32_and2456_y0(h_u_cla32_and2455_y0, h_u_cla32_and2454_y0, h_u_cla32_and2456_y0);
  and_gate and_gate_h_u_cla32_and2457_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2457_y0);
  and_gate and_gate_h_u_cla32_and2458_y0(h_u_cla32_and2457_y0, h_u_cla32_and2456_y0, h_u_cla32_and2458_y0);
  and_gate and_gate_h_u_cla32_and2459_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2459_y0);
  and_gate and_gate_h_u_cla32_and2460_y0(h_u_cla32_and2459_y0, h_u_cla32_and2458_y0, h_u_cla32_and2460_y0);
  and_gate and_gate_h_u_cla32_and2461_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2461_y0);
  and_gate and_gate_h_u_cla32_and2462_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2462_y0);
  and_gate and_gate_h_u_cla32_and2463_y0(h_u_cla32_and2462_y0, h_u_cla32_and2461_y0, h_u_cla32_and2463_y0);
  and_gate and_gate_h_u_cla32_and2464_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2464_y0);
  and_gate and_gate_h_u_cla32_and2465_y0(h_u_cla32_and2464_y0, h_u_cla32_and2463_y0, h_u_cla32_and2465_y0);
  and_gate and_gate_h_u_cla32_and2466_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and2466_y0);
  and_gate and_gate_h_u_cla32_and2467_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and2467_y0);
  and_gate and_gate_h_u_cla32_and2468_y0(h_u_cla32_and2467_y0, h_u_cla32_and2466_y0, h_u_cla32_and2468_y0);
  and_gate and_gate_h_u_cla32_and2469_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and2469_y0);
  or_gate or_gate_h_u_cla32_or171_y0(h_u_cla32_and2469_y0, h_u_cla32_and2145_y0, h_u_cla32_or171_y0);
  or_gate or_gate_h_u_cla32_or172_y0(h_u_cla32_or171_y0, h_u_cla32_and2180_y0, h_u_cla32_or172_y0);
  or_gate or_gate_h_u_cla32_or173_y0(h_u_cla32_or172_y0, h_u_cla32_and2213_y0, h_u_cla32_or173_y0);
  or_gate or_gate_h_u_cla32_or174_y0(h_u_cla32_or173_y0, h_u_cla32_and2244_y0, h_u_cla32_or174_y0);
  or_gate or_gate_h_u_cla32_or175_y0(h_u_cla32_or174_y0, h_u_cla32_and2273_y0, h_u_cla32_or175_y0);
  or_gate or_gate_h_u_cla32_or176_y0(h_u_cla32_or175_y0, h_u_cla32_and2300_y0, h_u_cla32_or176_y0);
  or_gate or_gate_h_u_cla32_or177_y0(h_u_cla32_or176_y0, h_u_cla32_and2325_y0, h_u_cla32_or177_y0);
  or_gate or_gate_h_u_cla32_or178_y0(h_u_cla32_or177_y0, h_u_cla32_and2348_y0, h_u_cla32_or178_y0);
  or_gate or_gate_h_u_cla32_or179_y0(h_u_cla32_or178_y0, h_u_cla32_and2369_y0, h_u_cla32_or179_y0);
  or_gate or_gate_h_u_cla32_or180_y0(h_u_cla32_or179_y0, h_u_cla32_and2388_y0, h_u_cla32_or180_y0);
  or_gate or_gate_h_u_cla32_or181_y0(h_u_cla32_or180_y0, h_u_cla32_and2405_y0, h_u_cla32_or181_y0);
  or_gate or_gate_h_u_cla32_or182_y0(h_u_cla32_or181_y0, h_u_cla32_and2420_y0, h_u_cla32_or182_y0);
  or_gate or_gate_h_u_cla32_or183_y0(h_u_cla32_or182_y0, h_u_cla32_and2433_y0, h_u_cla32_or183_y0);
  or_gate or_gate_h_u_cla32_or184_y0(h_u_cla32_or183_y0, h_u_cla32_and2444_y0, h_u_cla32_or184_y0);
  or_gate or_gate_h_u_cla32_or185_y0(h_u_cla32_or184_y0, h_u_cla32_and2453_y0, h_u_cla32_or185_y0);
  or_gate or_gate_h_u_cla32_or186_y0(h_u_cla32_or185_y0, h_u_cla32_and2460_y0, h_u_cla32_or186_y0);
  or_gate or_gate_h_u_cla32_or187_y0(h_u_cla32_or186_y0, h_u_cla32_and2465_y0, h_u_cla32_or187_y0);
  or_gate or_gate_h_u_cla32_or188_y0(h_u_cla32_or187_y0, h_u_cla32_and2468_y0, h_u_cla32_or188_y0);
  or_gate or_gate_h_u_cla32_or189_y0(h_u_cla32_pg_logic18_y1, h_u_cla32_or188_y0, h_u_cla32_or189_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic19_y0(a_19, b_19, h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_pg_logic19_y2);
  xor_gate xor_gate_h_u_cla32_xor19_y0(h_u_cla32_pg_logic19_y2, h_u_cla32_or189_y0, h_u_cla32_xor19_y0);
  and_gate and_gate_h_u_cla32_and2470_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and2470_y0);
  and_gate and_gate_h_u_cla32_and2471_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and2471_y0);
  and_gate and_gate_h_u_cla32_and2472_y0(h_u_cla32_and2471_y0, h_u_cla32_and2470_y0, h_u_cla32_and2472_y0);
  and_gate and_gate_h_u_cla32_and2473_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and2473_y0);
  and_gate and_gate_h_u_cla32_and2474_y0(h_u_cla32_and2473_y0, h_u_cla32_and2472_y0, h_u_cla32_and2474_y0);
  and_gate and_gate_h_u_cla32_and2475_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and2475_y0);
  and_gate and_gate_h_u_cla32_and2476_y0(h_u_cla32_and2475_y0, h_u_cla32_and2474_y0, h_u_cla32_and2476_y0);
  and_gate and_gate_h_u_cla32_and2477_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and2477_y0);
  and_gate and_gate_h_u_cla32_and2478_y0(h_u_cla32_and2477_y0, h_u_cla32_and2476_y0, h_u_cla32_and2478_y0);
  and_gate and_gate_h_u_cla32_and2479_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and2479_y0);
  and_gate and_gate_h_u_cla32_and2480_y0(h_u_cla32_and2479_y0, h_u_cla32_and2478_y0, h_u_cla32_and2480_y0);
  and_gate and_gate_h_u_cla32_and2481_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and2481_y0);
  and_gate and_gate_h_u_cla32_and2482_y0(h_u_cla32_and2481_y0, h_u_cla32_and2480_y0, h_u_cla32_and2482_y0);
  and_gate and_gate_h_u_cla32_and2483_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and2483_y0);
  and_gate and_gate_h_u_cla32_and2484_y0(h_u_cla32_and2483_y0, h_u_cla32_and2482_y0, h_u_cla32_and2484_y0);
  and_gate and_gate_h_u_cla32_and2485_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and2485_y0);
  and_gate and_gate_h_u_cla32_and2486_y0(h_u_cla32_and2485_y0, h_u_cla32_and2484_y0, h_u_cla32_and2486_y0);
  and_gate and_gate_h_u_cla32_and2487_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and2487_y0);
  and_gate and_gate_h_u_cla32_and2488_y0(h_u_cla32_and2487_y0, h_u_cla32_and2486_y0, h_u_cla32_and2488_y0);
  and_gate and_gate_h_u_cla32_and2489_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and2489_y0);
  and_gate and_gate_h_u_cla32_and2490_y0(h_u_cla32_and2489_y0, h_u_cla32_and2488_y0, h_u_cla32_and2490_y0);
  and_gate and_gate_h_u_cla32_and2491_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and2491_y0);
  and_gate and_gate_h_u_cla32_and2492_y0(h_u_cla32_and2491_y0, h_u_cla32_and2490_y0, h_u_cla32_and2492_y0);
  and_gate and_gate_h_u_cla32_and2493_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and2493_y0);
  and_gate and_gate_h_u_cla32_and2494_y0(h_u_cla32_and2493_y0, h_u_cla32_and2492_y0, h_u_cla32_and2494_y0);
  and_gate and_gate_h_u_cla32_and2495_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and2495_y0);
  and_gate and_gate_h_u_cla32_and2496_y0(h_u_cla32_and2495_y0, h_u_cla32_and2494_y0, h_u_cla32_and2496_y0);
  and_gate and_gate_h_u_cla32_and2497_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and2497_y0);
  and_gate and_gate_h_u_cla32_and2498_y0(h_u_cla32_and2497_y0, h_u_cla32_and2496_y0, h_u_cla32_and2498_y0);
  and_gate and_gate_h_u_cla32_and2499_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and2499_y0);
  and_gate and_gate_h_u_cla32_and2500_y0(h_u_cla32_and2499_y0, h_u_cla32_and2498_y0, h_u_cla32_and2500_y0);
  and_gate and_gate_h_u_cla32_and2501_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and2501_y0);
  and_gate and_gate_h_u_cla32_and2502_y0(h_u_cla32_and2501_y0, h_u_cla32_and2500_y0, h_u_cla32_and2502_y0);
  and_gate and_gate_h_u_cla32_and2503_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and2503_y0);
  and_gate and_gate_h_u_cla32_and2504_y0(h_u_cla32_and2503_y0, h_u_cla32_and2502_y0, h_u_cla32_and2504_y0);
  and_gate and_gate_h_u_cla32_and2505_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and2505_y0);
  and_gate and_gate_h_u_cla32_and2506_y0(h_u_cla32_and2505_y0, h_u_cla32_and2504_y0, h_u_cla32_and2506_y0);
  and_gate and_gate_h_u_cla32_and2507_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and2507_y0);
  and_gate and_gate_h_u_cla32_and2508_y0(h_u_cla32_and2507_y0, h_u_cla32_and2506_y0, h_u_cla32_and2508_y0);
  and_gate and_gate_h_u_cla32_and2509_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2509_y0);
  and_gate and_gate_h_u_cla32_and2510_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2510_y0);
  and_gate and_gate_h_u_cla32_and2511_y0(h_u_cla32_and2510_y0, h_u_cla32_and2509_y0, h_u_cla32_and2511_y0);
  and_gate and_gate_h_u_cla32_and2512_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2512_y0);
  and_gate and_gate_h_u_cla32_and2513_y0(h_u_cla32_and2512_y0, h_u_cla32_and2511_y0, h_u_cla32_and2513_y0);
  and_gate and_gate_h_u_cla32_and2514_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2514_y0);
  and_gate and_gate_h_u_cla32_and2515_y0(h_u_cla32_and2514_y0, h_u_cla32_and2513_y0, h_u_cla32_and2515_y0);
  and_gate and_gate_h_u_cla32_and2516_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2516_y0);
  and_gate and_gate_h_u_cla32_and2517_y0(h_u_cla32_and2516_y0, h_u_cla32_and2515_y0, h_u_cla32_and2517_y0);
  and_gate and_gate_h_u_cla32_and2518_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2518_y0);
  and_gate and_gate_h_u_cla32_and2519_y0(h_u_cla32_and2518_y0, h_u_cla32_and2517_y0, h_u_cla32_and2519_y0);
  and_gate and_gate_h_u_cla32_and2520_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2520_y0);
  and_gate and_gate_h_u_cla32_and2521_y0(h_u_cla32_and2520_y0, h_u_cla32_and2519_y0, h_u_cla32_and2521_y0);
  and_gate and_gate_h_u_cla32_and2522_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2522_y0);
  and_gate and_gate_h_u_cla32_and2523_y0(h_u_cla32_and2522_y0, h_u_cla32_and2521_y0, h_u_cla32_and2523_y0);
  and_gate and_gate_h_u_cla32_and2524_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2524_y0);
  and_gate and_gate_h_u_cla32_and2525_y0(h_u_cla32_and2524_y0, h_u_cla32_and2523_y0, h_u_cla32_and2525_y0);
  and_gate and_gate_h_u_cla32_and2526_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2526_y0);
  and_gate and_gate_h_u_cla32_and2527_y0(h_u_cla32_and2526_y0, h_u_cla32_and2525_y0, h_u_cla32_and2527_y0);
  and_gate and_gate_h_u_cla32_and2528_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2528_y0);
  and_gate and_gate_h_u_cla32_and2529_y0(h_u_cla32_and2528_y0, h_u_cla32_and2527_y0, h_u_cla32_and2529_y0);
  and_gate and_gate_h_u_cla32_and2530_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2530_y0);
  and_gate and_gate_h_u_cla32_and2531_y0(h_u_cla32_and2530_y0, h_u_cla32_and2529_y0, h_u_cla32_and2531_y0);
  and_gate and_gate_h_u_cla32_and2532_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2532_y0);
  and_gate and_gate_h_u_cla32_and2533_y0(h_u_cla32_and2532_y0, h_u_cla32_and2531_y0, h_u_cla32_and2533_y0);
  and_gate and_gate_h_u_cla32_and2534_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2534_y0);
  and_gate and_gate_h_u_cla32_and2535_y0(h_u_cla32_and2534_y0, h_u_cla32_and2533_y0, h_u_cla32_and2535_y0);
  and_gate and_gate_h_u_cla32_and2536_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2536_y0);
  and_gate and_gate_h_u_cla32_and2537_y0(h_u_cla32_and2536_y0, h_u_cla32_and2535_y0, h_u_cla32_and2537_y0);
  and_gate and_gate_h_u_cla32_and2538_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2538_y0);
  and_gate and_gate_h_u_cla32_and2539_y0(h_u_cla32_and2538_y0, h_u_cla32_and2537_y0, h_u_cla32_and2539_y0);
  and_gate and_gate_h_u_cla32_and2540_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2540_y0);
  and_gate and_gate_h_u_cla32_and2541_y0(h_u_cla32_and2540_y0, h_u_cla32_and2539_y0, h_u_cla32_and2541_y0);
  and_gate and_gate_h_u_cla32_and2542_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2542_y0);
  and_gate and_gate_h_u_cla32_and2543_y0(h_u_cla32_and2542_y0, h_u_cla32_and2541_y0, h_u_cla32_and2543_y0);
  and_gate and_gate_h_u_cla32_and2544_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2544_y0);
  and_gate and_gate_h_u_cla32_and2545_y0(h_u_cla32_and2544_y0, h_u_cla32_and2543_y0, h_u_cla32_and2545_y0);
  and_gate and_gate_h_u_cla32_and2546_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2546_y0);
  and_gate and_gate_h_u_cla32_and2547_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2547_y0);
  and_gate and_gate_h_u_cla32_and2548_y0(h_u_cla32_and2547_y0, h_u_cla32_and2546_y0, h_u_cla32_and2548_y0);
  and_gate and_gate_h_u_cla32_and2549_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2549_y0);
  and_gate and_gate_h_u_cla32_and2550_y0(h_u_cla32_and2549_y0, h_u_cla32_and2548_y0, h_u_cla32_and2550_y0);
  and_gate and_gate_h_u_cla32_and2551_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2551_y0);
  and_gate and_gate_h_u_cla32_and2552_y0(h_u_cla32_and2551_y0, h_u_cla32_and2550_y0, h_u_cla32_and2552_y0);
  and_gate and_gate_h_u_cla32_and2553_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2553_y0);
  and_gate and_gate_h_u_cla32_and2554_y0(h_u_cla32_and2553_y0, h_u_cla32_and2552_y0, h_u_cla32_and2554_y0);
  and_gate and_gate_h_u_cla32_and2555_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2555_y0);
  and_gate and_gate_h_u_cla32_and2556_y0(h_u_cla32_and2555_y0, h_u_cla32_and2554_y0, h_u_cla32_and2556_y0);
  and_gate and_gate_h_u_cla32_and2557_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2557_y0);
  and_gate and_gate_h_u_cla32_and2558_y0(h_u_cla32_and2557_y0, h_u_cla32_and2556_y0, h_u_cla32_and2558_y0);
  and_gate and_gate_h_u_cla32_and2559_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2559_y0);
  and_gate and_gate_h_u_cla32_and2560_y0(h_u_cla32_and2559_y0, h_u_cla32_and2558_y0, h_u_cla32_and2560_y0);
  and_gate and_gate_h_u_cla32_and2561_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2561_y0);
  and_gate and_gate_h_u_cla32_and2562_y0(h_u_cla32_and2561_y0, h_u_cla32_and2560_y0, h_u_cla32_and2562_y0);
  and_gate and_gate_h_u_cla32_and2563_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2563_y0);
  and_gate and_gate_h_u_cla32_and2564_y0(h_u_cla32_and2563_y0, h_u_cla32_and2562_y0, h_u_cla32_and2564_y0);
  and_gate and_gate_h_u_cla32_and2565_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2565_y0);
  and_gate and_gate_h_u_cla32_and2566_y0(h_u_cla32_and2565_y0, h_u_cla32_and2564_y0, h_u_cla32_and2566_y0);
  and_gate and_gate_h_u_cla32_and2567_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2567_y0);
  and_gate and_gate_h_u_cla32_and2568_y0(h_u_cla32_and2567_y0, h_u_cla32_and2566_y0, h_u_cla32_and2568_y0);
  and_gate and_gate_h_u_cla32_and2569_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2569_y0);
  and_gate and_gate_h_u_cla32_and2570_y0(h_u_cla32_and2569_y0, h_u_cla32_and2568_y0, h_u_cla32_and2570_y0);
  and_gate and_gate_h_u_cla32_and2571_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2571_y0);
  and_gate and_gate_h_u_cla32_and2572_y0(h_u_cla32_and2571_y0, h_u_cla32_and2570_y0, h_u_cla32_and2572_y0);
  and_gate and_gate_h_u_cla32_and2573_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2573_y0);
  and_gate and_gate_h_u_cla32_and2574_y0(h_u_cla32_and2573_y0, h_u_cla32_and2572_y0, h_u_cla32_and2574_y0);
  and_gate and_gate_h_u_cla32_and2575_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2575_y0);
  and_gate and_gate_h_u_cla32_and2576_y0(h_u_cla32_and2575_y0, h_u_cla32_and2574_y0, h_u_cla32_and2576_y0);
  and_gate and_gate_h_u_cla32_and2577_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2577_y0);
  and_gate and_gate_h_u_cla32_and2578_y0(h_u_cla32_and2577_y0, h_u_cla32_and2576_y0, h_u_cla32_and2578_y0);
  and_gate and_gate_h_u_cla32_and2579_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2579_y0);
  and_gate and_gate_h_u_cla32_and2580_y0(h_u_cla32_and2579_y0, h_u_cla32_and2578_y0, h_u_cla32_and2580_y0);
  and_gate and_gate_h_u_cla32_and2581_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2581_y0);
  and_gate and_gate_h_u_cla32_and2582_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2582_y0);
  and_gate and_gate_h_u_cla32_and2583_y0(h_u_cla32_and2582_y0, h_u_cla32_and2581_y0, h_u_cla32_and2583_y0);
  and_gate and_gate_h_u_cla32_and2584_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2584_y0);
  and_gate and_gate_h_u_cla32_and2585_y0(h_u_cla32_and2584_y0, h_u_cla32_and2583_y0, h_u_cla32_and2585_y0);
  and_gate and_gate_h_u_cla32_and2586_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2586_y0);
  and_gate and_gate_h_u_cla32_and2587_y0(h_u_cla32_and2586_y0, h_u_cla32_and2585_y0, h_u_cla32_and2587_y0);
  and_gate and_gate_h_u_cla32_and2588_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2588_y0);
  and_gate and_gate_h_u_cla32_and2589_y0(h_u_cla32_and2588_y0, h_u_cla32_and2587_y0, h_u_cla32_and2589_y0);
  and_gate and_gate_h_u_cla32_and2590_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2590_y0);
  and_gate and_gate_h_u_cla32_and2591_y0(h_u_cla32_and2590_y0, h_u_cla32_and2589_y0, h_u_cla32_and2591_y0);
  and_gate and_gate_h_u_cla32_and2592_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2592_y0);
  and_gate and_gate_h_u_cla32_and2593_y0(h_u_cla32_and2592_y0, h_u_cla32_and2591_y0, h_u_cla32_and2593_y0);
  and_gate and_gate_h_u_cla32_and2594_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2594_y0);
  and_gate and_gate_h_u_cla32_and2595_y0(h_u_cla32_and2594_y0, h_u_cla32_and2593_y0, h_u_cla32_and2595_y0);
  and_gate and_gate_h_u_cla32_and2596_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2596_y0);
  and_gate and_gate_h_u_cla32_and2597_y0(h_u_cla32_and2596_y0, h_u_cla32_and2595_y0, h_u_cla32_and2597_y0);
  and_gate and_gate_h_u_cla32_and2598_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2598_y0);
  and_gate and_gate_h_u_cla32_and2599_y0(h_u_cla32_and2598_y0, h_u_cla32_and2597_y0, h_u_cla32_and2599_y0);
  and_gate and_gate_h_u_cla32_and2600_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2600_y0);
  and_gate and_gate_h_u_cla32_and2601_y0(h_u_cla32_and2600_y0, h_u_cla32_and2599_y0, h_u_cla32_and2601_y0);
  and_gate and_gate_h_u_cla32_and2602_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2602_y0);
  and_gate and_gate_h_u_cla32_and2603_y0(h_u_cla32_and2602_y0, h_u_cla32_and2601_y0, h_u_cla32_and2603_y0);
  and_gate and_gate_h_u_cla32_and2604_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2604_y0);
  and_gate and_gate_h_u_cla32_and2605_y0(h_u_cla32_and2604_y0, h_u_cla32_and2603_y0, h_u_cla32_and2605_y0);
  and_gate and_gate_h_u_cla32_and2606_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2606_y0);
  and_gate and_gate_h_u_cla32_and2607_y0(h_u_cla32_and2606_y0, h_u_cla32_and2605_y0, h_u_cla32_and2607_y0);
  and_gate and_gate_h_u_cla32_and2608_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2608_y0);
  and_gate and_gate_h_u_cla32_and2609_y0(h_u_cla32_and2608_y0, h_u_cla32_and2607_y0, h_u_cla32_and2609_y0);
  and_gate and_gate_h_u_cla32_and2610_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2610_y0);
  and_gate and_gate_h_u_cla32_and2611_y0(h_u_cla32_and2610_y0, h_u_cla32_and2609_y0, h_u_cla32_and2611_y0);
  and_gate and_gate_h_u_cla32_and2612_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2612_y0);
  and_gate and_gate_h_u_cla32_and2613_y0(h_u_cla32_and2612_y0, h_u_cla32_and2611_y0, h_u_cla32_and2613_y0);
  and_gate and_gate_h_u_cla32_and2614_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2614_y0);
  and_gate and_gate_h_u_cla32_and2615_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2615_y0);
  and_gate and_gate_h_u_cla32_and2616_y0(h_u_cla32_and2615_y0, h_u_cla32_and2614_y0, h_u_cla32_and2616_y0);
  and_gate and_gate_h_u_cla32_and2617_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2617_y0);
  and_gate and_gate_h_u_cla32_and2618_y0(h_u_cla32_and2617_y0, h_u_cla32_and2616_y0, h_u_cla32_and2618_y0);
  and_gate and_gate_h_u_cla32_and2619_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2619_y0);
  and_gate and_gate_h_u_cla32_and2620_y0(h_u_cla32_and2619_y0, h_u_cla32_and2618_y0, h_u_cla32_and2620_y0);
  and_gate and_gate_h_u_cla32_and2621_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2621_y0);
  and_gate and_gate_h_u_cla32_and2622_y0(h_u_cla32_and2621_y0, h_u_cla32_and2620_y0, h_u_cla32_and2622_y0);
  and_gate and_gate_h_u_cla32_and2623_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2623_y0);
  and_gate and_gate_h_u_cla32_and2624_y0(h_u_cla32_and2623_y0, h_u_cla32_and2622_y0, h_u_cla32_and2624_y0);
  and_gate and_gate_h_u_cla32_and2625_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2625_y0);
  and_gate and_gate_h_u_cla32_and2626_y0(h_u_cla32_and2625_y0, h_u_cla32_and2624_y0, h_u_cla32_and2626_y0);
  and_gate and_gate_h_u_cla32_and2627_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2627_y0);
  and_gate and_gate_h_u_cla32_and2628_y0(h_u_cla32_and2627_y0, h_u_cla32_and2626_y0, h_u_cla32_and2628_y0);
  and_gate and_gate_h_u_cla32_and2629_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2629_y0);
  and_gate and_gate_h_u_cla32_and2630_y0(h_u_cla32_and2629_y0, h_u_cla32_and2628_y0, h_u_cla32_and2630_y0);
  and_gate and_gate_h_u_cla32_and2631_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2631_y0);
  and_gate and_gate_h_u_cla32_and2632_y0(h_u_cla32_and2631_y0, h_u_cla32_and2630_y0, h_u_cla32_and2632_y0);
  and_gate and_gate_h_u_cla32_and2633_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2633_y0);
  and_gate and_gate_h_u_cla32_and2634_y0(h_u_cla32_and2633_y0, h_u_cla32_and2632_y0, h_u_cla32_and2634_y0);
  and_gate and_gate_h_u_cla32_and2635_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2635_y0);
  and_gate and_gate_h_u_cla32_and2636_y0(h_u_cla32_and2635_y0, h_u_cla32_and2634_y0, h_u_cla32_and2636_y0);
  and_gate and_gate_h_u_cla32_and2637_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2637_y0);
  and_gate and_gate_h_u_cla32_and2638_y0(h_u_cla32_and2637_y0, h_u_cla32_and2636_y0, h_u_cla32_and2638_y0);
  and_gate and_gate_h_u_cla32_and2639_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2639_y0);
  and_gate and_gate_h_u_cla32_and2640_y0(h_u_cla32_and2639_y0, h_u_cla32_and2638_y0, h_u_cla32_and2640_y0);
  and_gate and_gate_h_u_cla32_and2641_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2641_y0);
  and_gate and_gate_h_u_cla32_and2642_y0(h_u_cla32_and2641_y0, h_u_cla32_and2640_y0, h_u_cla32_and2642_y0);
  and_gate and_gate_h_u_cla32_and2643_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and2643_y0);
  and_gate and_gate_h_u_cla32_and2644_y0(h_u_cla32_and2643_y0, h_u_cla32_and2642_y0, h_u_cla32_and2644_y0);
  and_gate and_gate_h_u_cla32_and2645_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2645_y0);
  and_gate and_gate_h_u_cla32_and2646_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2646_y0);
  and_gate and_gate_h_u_cla32_and2647_y0(h_u_cla32_and2646_y0, h_u_cla32_and2645_y0, h_u_cla32_and2647_y0);
  and_gate and_gate_h_u_cla32_and2648_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2648_y0);
  and_gate and_gate_h_u_cla32_and2649_y0(h_u_cla32_and2648_y0, h_u_cla32_and2647_y0, h_u_cla32_and2649_y0);
  and_gate and_gate_h_u_cla32_and2650_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2650_y0);
  and_gate and_gate_h_u_cla32_and2651_y0(h_u_cla32_and2650_y0, h_u_cla32_and2649_y0, h_u_cla32_and2651_y0);
  and_gate and_gate_h_u_cla32_and2652_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2652_y0);
  and_gate and_gate_h_u_cla32_and2653_y0(h_u_cla32_and2652_y0, h_u_cla32_and2651_y0, h_u_cla32_and2653_y0);
  and_gate and_gate_h_u_cla32_and2654_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2654_y0);
  and_gate and_gate_h_u_cla32_and2655_y0(h_u_cla32_and2654_y0, h_u_cla32_and2653_y0, h_u_cla32_and2655_y0);
  and_gate and_gate_h_u_cla32_and2656_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2656_y0);
  and_gate and_gate_h_u_cla32_and2657_y0(h_u_cla32_and2656_y0, h_u_cla32_and2655_y0, h_u_cla32_and2657_y0);
  and_gate and_gate_h_u_cla32_and2658_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2658_y0);
  and_gate and_gate_h_u_cla32_and2659_y0(h_u_cla32_and2658_y0, h_u_cla32_and2657_y0, h_u_cla32_and2659_y0);
  and_gate and_gate_h_u_cla32_and2660_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2660_y0);
  and_gate and_gate_h_u_cla32_and2661_y0(h_u_cla32_and2660_y0, h_u_cla32_and2659_y0, h_u_cla32_and2661_y0);
  and_gate and_gate_h_u_cla32_and2662_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2662_y0);
  and_gate and_gate_h_u_cla32_and2663_y0(h_u_cla32_and2662_y0, h_u_cla32_and2661_y0, h_u_cla32_and2663_y0);
  and_gate and_gate_h_u_cla32_and2664_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2664_y0);
  and_gate and_gate_h_u_cla32_and2665_y0(h_u_cla32_and2664_y0, h_u_cla32_and2663_y0, h_u_cla32_and2665_y0);
  and_gate and_gate_h_u_cla32_and2666_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2666_y0);
  and_gate and_gate_h_u_cla32_and2667_y0(h_u_cla32_and2666_y0, h_u_cla32_and2665_y0, h_u_cla32_and2667_y0);
  and_gate and_gate_h_u_cla32_and2668_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2668_y0);
  and_gate and_gate_h_u_cla32_and2669_y0(h_u_cla32_and2668_y0, h_u_cla32_and2667_y0, h_u_cla32_and2669_y0);
  and_gate and_gate_h_u_cla32_and2670_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2670_y0);
  and_gate and_gate_h_u_cla32_and2671_y0(h_u_cla32_and2670_y0, h_u_cla32_and2669_y0, h_u_cla32_and2671_y0);
  and_gate and_gate_h_u_cla32_and2672_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and2672_y0);
  and_gate and_gate_h_u_cla32_and2673_y0(h_u_cla32_and2672_y0, h_u_cla32_and2671_y0, h_u_cla32_and2673_y0);
  and_gate and_gate_h_u_cla32_and2674_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2674_y0);
  and_gate and_gate_h_u_cla32_and2675_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2675_y0);
  and_gate and_gate_h_u_cla32_and2676_y0(h_u_cla32_and2675_y0, h_u_cla32_and2674_y0, h_u_cla32_and2676_y0);
  and_gate and_gate_h_u_cla32_and2677_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2677_y0);
  and_gate and_gate_h_u_cla32_and2678_y0(h_u_cla32_and2677_y0, h_u_cla32_and2676_y0, h_u_cla32_and2678_y0);
  and_gate and_gate_h_u_cla32_and2679_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2679_y0);
  and_gate and_gate_h_u_cla32_and2680_y0(h_u_cla32_and2679_y0, h_u_cla32_and2678_y0, h_u_cla32_and2680_y0);
  and_gate and_gate_h_u_cla32_and2681_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2681_y0);
  and_gate and_gate_h_u_cla32_and2682_y0(h_u_cla32_and2681_y0, h_u_cla32_and2680_y0, h_u_cla32_and2682_y0);
  and_gate and_gate_h_u_cla32_and2683_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2683_y0);
  and_gate and_gate_h_u_cla32_and2684_y0(h_u_cla32_and2683_y0, h_u_cla32_and2682_y0, h_u_cla32_and2684_y0);
  and_gate and_gate_h_u_cla32_and2685_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2685_y0);
  and_gate and_gate_h_u_cla32_and2686_y0(h_u_cla32_and2685_y0, h_u_cla32_and2684_y0, h_u_cla32_and2686_y0);
  and_gate and_gate_h_u_cla32_and2687_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2687_y0);
  and_gate and_gate_h_u_cla32_and2688_y0(h_u_cla32_and2687_y0, h_u_cla32_and2686_y0, h_u_cla32_and2688_y0);
  and_gate and_gate_h_u_cla32_and2689_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2689_y0);
  and_gate and_gate_h_u_cla32_and2690_y0(h_u_cla32_and2689_y0, h_u_cla32_and2688_y0, h_u_cla32_and2690_y0);
  and_gate and_gate_h_u_cla32_and2691_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2691_y0);
  and_gate and_gate_h_u_cla32_and2692_y0(h_u_cla32_and2691_y0, h_u_cla32_and2690_y0, h_u_cla32_and2692_y0);
  and_gate and_gate_h_u_cla32_and2693_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2693_y0);
  and_gate and_gate_h_u_cla32_and2694_y0(h_u_cla32_and2693_y0, h_u_cla32_and2692_y0, h_u_cla32_and2694_y0);
  and_gate and_gate_h_u_cla32_and2695_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2695_y0);
  and_gate and_gate_h_u_cla32_and2696_y0(h_u_cla32_and2695_y0, h_u_cla32_and2694_y0, h_u_cla32_and2696_y0);
  and_gate and_gate_h_u_cla32_and2697_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2697_y0);
  and_gate and_gate_h_u_cla32_and2698_y0(h_u_cla32_and2697_y0, h_u_cla32_and2696_y0, h_u_cla32_and2698_y0);
  and_gate and_gate_h_u_cla32_and2699_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and2699_y0);
  and_gate and_gate_h_u_cla32_and2700_y0(h_u_cla32_and2699_y0, h_u_cla32_and2698_y0, h_u_cla32_and2700_y0);
  and_gate and_gate_h_u_cla32_and2701_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2701_y0);
  and_gate and_gate_h_u_cla32_and2702_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2702_y0);
  and_gate and_gate_h_u_cla32_and2703_y0(h_u_cla32_and2702_y0, h_u_cla32_and2701_y0, h_u_cla32_and2703_y0);
  and_gate and_gate_h_u_cla32_and2704_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2704_y0);
  and_gate and_gate_h_u_cla32_and2705_y0(h_u_cla32_and2704_y0, h_u_cla32_and2703_y0, h_u_cla32_and2705_y0);
  and_gate and_gate_h_u_cla32_and2706_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2706_y0);
  and_gate and_gate_h_u_cla32_and2707_y0(h_u_cla32_and2706_y0, h_u_cla32_and2705_y0, h_u_cla32_and2707_y0);
  and_gate and_gate_h_u_cla32_and2708_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2708_y0);
  and_gate and_gate_h_u_cla32_and2709_y0(h_u_cla32_and2708_y0, h_u_cla32_and2707_y0, h_u_cla32_and2709_y0);
  and_gate and_gate_h_u_cla32_and2710_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2710_y0);
  and_gate and_gate_h_u_cla32_and2711_y0(h_u_cla32_and2710_y0, h_u_cla32_and2709_y0, h_u_cla32_and2711_y0);
  and_gate and_gate_h_u_cla32_and2712_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2712_y0);
  and_gate and_gate_h_u_cla32_and2713_y0(h_u_cla32_and2712_y0, h_u_cla32_and2711_y0, h_u_cla32_and2713_y0);
  and_gate and_gate_h_u_cla32_and2714_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2714_y0);
  and_gate and_gate_h_u_cla32_and2715_y0(h_u_cla32_and2714_y0, h_u_cla32_and2713_y0, h_u_cla32_and2715_y0);
  and_gate and_gate_h_u_cla32_and2716_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2716_y0);
  and_gate and_gate_h_u_cla32_and2717_y0(h_u_cla32_and2716_y0, h_u_cla32_and2715_y0, h_u_cla32_and2717_y0);
  and_gate and_gate_h_u_cla32_and2718_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2718_y0);
  and_gate and_gate_h_u_cla32_and2719_y0(h_u_cla32_and2718_y0, h_u_cla32_and2717_y0, h_u_cla32_and2719_y0);
  and_gate and_gate_h_u_cla32_and2720_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2720_y0);
  and_gate and_gate_h_u_cla32_and2721_y0(h_u_cla32_and2720_y0, h_u_cla32_and2719_y0, h_u_cla32_and2721_y0);
  and_gate and_gate_h_u_cla32_and2722_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2722_y0);
  and_gate and_gate_h_u_cla32_and2723_y0(h_u_cla32_and2722_y0, h_u_cla32_and2721_y0, h_u_cla32_and2723_y0);
  and_gate and_gate_h_u_cla32_and2724_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and2724_y0);
  and_gate and_gate_h_u_cla32_and2725_y0(h_u_cla32_and2724_y0, h_u_cla32_and2723_y0, h_u_cla32_and2725_y0);
  and_gate and_gate_h_u_cla32_and2726_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2726_y0);
  and_gate and_gate_h_u_cla32_and2727_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2727_y0);
  and_gate and_gate_h_u_cla32_and2728_y0(h_u_cla32_and2727_y0, h_u_cla32_and2726_y0, h_u_cla32_and2728_y0);
  and_gate and_gate_h_u_cla32_and2729_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2729_y0);
  and_gate and_gate_h_u_cla32_and2730_y0(h_u_cla32_and2729_y0, h_u_cla32_and2728_y0, h_u_cla32_and2730_y0);
  and_gate and_gate_h_u_cla32_and2731_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2731_y0);
  and_gate and_gate_h_u_cla32_and2732_y0(h_u_cla32_and2731_y0, h_u_cla32_and2730_y0, h_u_cla32_and2732_y0);
  and_gate and_gate_h_u_cla32_and2733_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2733_y0);
  and_gate and_gate_h_u_cla32_and2734_y0(h_u_cla32_and2733_y0, h_u_cla32_and2732_y0, h_u_cla32_and2734_y0);
  and_gate and_gate_h_u_cla32_and2735_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2735_y0);
  and_gate and_gate_h_u_cla32_and2736_y0(h_u_cla32_and2735_y0, h_u_cla32_and2734_y0, h_u_cla32_and2736_y0);
  and_gate and_gate_h_u_cla32_and2737_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2737_y0);
  and_gate and_gate_h_u_cla32_and2738_y0(h_u_cla32_and2737_y0, h_u_cla32_and2736_y0, h_u_cla32_and2738_y0);
  and_gate and_gate_h_u_cla32_and2739_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2739_y0);
  and_gate and_gate_h_u_cla32_and2740_y0(h_u_cla32_and2739_y0, h_u_cla32_and2738_y0, h_u_cla32_and2740_y0);
  and_gate and_gate_h_u_cla32_and2741_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2741_y0);
  and_gate and_gate_h_u_cla32_and2742_y0(h_u_cla32_and2741_y0, h_u_cla32_and2740_y0, h_u_cla32_and2742_y0);
  and_gate and_gate_h_u_cla32_and2743_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2743_y0);
  and_gate and_gate_h_u_cla32_and2744_y0(h_u_cla32_and2743_y0, h_u_cla32_and2742_y0, h_u_cla32_and2744_y0);
  and_gate and_gate_h_u_cla32_and2745_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2745_y0);
  and_gate and_gate_h_u_cla32_and2746_y0(h_u_cla32_and2745_y0, h_u_cla32_and2744_y0, h_u_cla32_and2746_y0);
  and_gate and_gate_h_u_cla32_and2747_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and2747_y0);
  and_gate and_gate_h_u_cla32_and2748_y0(h_u_cla32_and2747_y0, h_u_cla32_and2746_y0, h_u_cla32_and2748_y0);
  and_gate and_gate_h_u_cla32_and2749_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2749_y0);
  and_gate and_gate_h_u_cla32_and2750_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2750_y0);
  and_gate and_gate_h_u_cla32_and2751_y0(h_u_cla32_and2750_y0, h_u_cla32_and2749_y0, h_u_cla32_and2751_y0);
  and_gate and_gate_h_u_cla32_and2752_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2752_y0);
  and_gate and_gate_h_u_cla32_and2753_y0(h_u_cla32_and2752_y0, h_u_cla32_and2751_y0, h_u_cla32_and2753_y0);
  and_gate and_gate_h_u_cla32_and2754_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2754_y0);
  and_gate and_gate_h_u_cla32_and2755_y0(h_u_cla32_and2754_y0, h_u_cla32_and2753_y0, h_u_cla32_and2755_y0);
  and_gate and_gate_h_u_cla32_and2756_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2756_y0);
  and_gate and_gate_h_u_cla32_and2757_y0(h_u_cla32_and2756_y0, h_u_cla32_and2755_y0, h_u_cla32_and2757_y0);
  and_gate and_gate_h_u_cla32_and2758_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2758_y0);
  and_gate and_gate_h_u_cla32_and2759_y0(h_u_cla32_and2758_y0, h_u_cla32_and2757_y0, h_u_cla32_and2759_y0);
  and_gate and_gate_h_u_cla32_and2760_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2760_y0);
  and_gate and_gate_h_u_cla32_and2761_y0(h_u_cla32_and2760_y0, h_u_cla32_and2759_y0, h_u_cla32_and2761_y0);
  and_gate and_gate_h_u_cla32_and2762_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2762_y0);
  and_gate and_gate_h_u_cla32_and2763_y0(h_u_cla32_and2762_y0, h_u_cla32_and2761_y0, h_u_cla32_and2763_y0);
  and_gate and_gate_h_u_cla32_and2764_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2764_y0);
  and_gate and_gate_h_u_cla32_and2765_y0(h_u_cla32_and2764_y0, h_u_cla32_and2763_y0, h_u_cla32_and2765_y0);
  and_gate and_gate_h_u_cla32_and2766_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2766_y0);
  and_gate and_gate_h_u_cla32_and2767_y0(h_u_cla32_and2766_y0, h_u_cla32_and2765_y0, h_u_cla32_and2767_y0);
  and_gate and_gate_h_u_cla32_and2768_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and2768_y0);
  and_gate and_gate_h_u_cla32_and2769_y0(h_u_cla32_and2768_y0, h_u_cla32_and2767_y0, h_u_cla32_and2769_y0);
  and_gate and_gate_h_u_cla32_and2770_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2770_y0);
  and_gate and_gate_h_u_cla32_and2771_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2771_y0);
  and_gate and_gate_h_u_cla32_and2772_y0(h_u_cla32_and2771_y0, h_u_cla32_and2770_y0, h_u_cla32_and2772_y0);
  and_gate and_gate_h_u_cla32_and2773_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2773_y0);
  and_gate and_gate_h_u_cla32_and2774_y0(h_u_cla32_and2773_y0, h_u_cla32_and2772_y0, h_u_cla32_and2774_y0);
  and_gate and_gate_h_u_cla32_and2775_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2775_y0);
  and_gate and_gate_h_u_cla32_and2776_y0(h_u_cla32_and2775_y0, h_u_cla32_and2774_y0, h_u_cla32_and2776_y0);
  and_gate and_gate_h_u_cla32_and2777_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2777_y0);
  and_gate and_gate_h_u_cla32_and2778_y0(h_u_cla32_and2777_y0, h_u_cla32_and2776_y0, h_u_cla32_and2778_y0);
  and_gate and_gate_h_u_cla32_and2779_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2779_y0);
  and_gate and_gate_h_u_cla32_and2780_y0(h_u_cla32_and2779_y0, h_u_cla32_and2778_y0, h_u_cla32_and2780_y0);
  and_gate and_gate_h_u_cla32_and2781_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2781_y0);
  and_gate and_gate_h_u_cla32_and2782_y0(h_u_cla32_and2781_y0, h_u_cla32_and2780_y0, h_u_cla32_and2782_y0);
  and_gate and_gate_h_u_cla32_and2783_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2783_y0);
  and_gate and_gate_h_u_cla32_and2784_y0(h_u_cla32_and2783_y0, h_u_cla32_and2782_y0, h_u_cla32_and2784_y0);
  and_gate and_gate_h_u_cla32_and2785_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2785_y0);
  and_gate and_gate_h_u_cla32_and2786_y0(h_u_cla32_and2785_y0, h_u_cla32_and2784_y0, h_u_cla32_and2786_y0);
  and_gate and_gate_h_u_cla32_and2787_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and2787_y0);
  and_gate and_gate_h_u_cla32_and2788_y0(h_u_cla32_and2787_y0, h_u_cla32_and2786_y0, h_u_cla32_and2788_y0);
  and_gate and_gate_h_u_cla32_and2789_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2789_y0);
  and_gate and_gate_h_u_cla32_and2790_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2790_y0);
  and_gate and_gate_h_u_cla32_and2791_y0(h_u_cla32_and2790_y0, h_u_cla32_and2789_y0, h_u_cla32_and2791_y0);
  and_gate and_gate_h_u_cla32_and2792_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2792_y0);
  and_gate and_gate_h_u_cla32_and2793_y0(h_u_cla32_and2792_y0, h_u_cla32_and2791_y0, h_u_cla32_and2793_y0);
  and_gate and_gate_h_u_cla32_and2794_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2794_y0);
  and_gate and_gate_h_u_cla32_and2795_y0(h_u_cla32_and2794_y0, h_u_cla32_and2793_y0, h_u_cla32_and2795_y0);
  and_gate and_gate_h_u_cla32_and2796_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2796_y0);
  and_gate and_gate_h_u_cla32_and2797_y0(h_u_cla32_and2796_y0, h_u_cla32_and2795_y0, h_u_cla32_and2797_y0);
  and_gate and_gate_h_u_cla32_and2798_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2798_y0);
  and_gate and_gate_h_u_cla32_and2799_y0(h_u_cla32_and2798_y0, h_u_cla32_and2797_y0, h_u_cla32_and2799_y0);
  and_gate and_gate_h_u_cla32_and2800_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2800_y0);
  and_gate and_gate_h_u_cla32_and2801_y0(h_u_cla32_and2800_y0, h_u_cla32_and2799_y0, h_u_cla32_and2801_y0);
  and_gate and_gate_h_u_cla32_and2802_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2802_y0);
  and_gate and_gate_h_u_cla32_and2803_y0(h_u_cla32_and2802_y0, h_u_cla32_and2801_y0, h_u_cla32_and2803_y0);
  and_gate and_gate_h_u_cla32_and2804_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and2804_y0);
  and_gate and_gate_h_u_cla32_and2805_y0(h_u_cla32_and2804_y0, h_u_cla32_and2803_y0, h_u_cla32_and2805_y0);
  and_gate and_gate_h_u_cla32_and2806_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2806_y0);
  and_gate and_gate_h_u_cla32_and2807_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2807_y0);
  and_gate and_gate_h_u_cla32_and2808_y0(h_u_cla32_and2807_y0, h_u_cla32_and2806_y0, h_u_cla32_and2808_y0);
  and_gate and_gate_h_u_cla32_and2809_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2809_y0);
  and_gate and_gate_h_u_cla32_and2810_y0(h_u_cla32_and2809_y0, h_u_cla32_and2808_y0, h_u_cla32_and2810_y0);
  and_gate and_gate_h_u_cla32_and2811_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2811_y0);
  and_gate and_gate_h_u_cla32_and2812_y0(h_u_cla32_and2811_y0, h_u_cla32_and2810_y0, h_u_cla32_and2812_y0);
  and_gate and_gate_h_u_cla32_and2813_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2813_y0);
  and_gate and_gate_h_u_cla32_and2814_y0(h_u_cla32_and2813_y0, h_u_cla32_and2812_y0, h_u_cla32_and2814_y0);
  and_gate and_gate_h_u_cla32_and2815_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2815_y0);
  and_gate and_gate_h_u_cla32_and2816_y0(h_u_cla32_and2815_y0, h_u_cla32_and2814_y0, h_u_cla32_and2816_y0);
  and_gate and_gate_h_u_cla32_and2817_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2817_y0);
  and_gate and_gate_h_u_cla32_and2818_y0(h_u_cla32_and2817_y0, h_u_cla32_and2816_y0, h_u_cla32_and2818_y0);
  and_gate and_gate_h_u_cla32_and2819_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and2819_y0);
  and_gate and_gate_h_u_cla32_and2820_y0(h_u_cla32_and2819_y0, h_u_cla32_and2818_y0, h_u_cla32_and2820_y0);
  and_gate and_gate_h_u_cla32_and2821_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2821_y0);
  and_gate and_gate_h_u_cla32_and2822_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2822_y0);
  and_gate and_gate_h_u_cla32_and2823_y0(h_u_cla32_and2822_y0, h_u_cla32_and2821_y0, h_u_cla32_and2823_y0);
  and_gate and_gate_h_u_cla32_and2824_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2824_y0);
  and_gate and_gate_h_u_cla32_and2825_y0(h_u_cla32_and2824_y0, h_u_cla32_and2823_y0, h_u_cla32_and2825_y0);
  and_gate and_gate_h_u_cla32_and2826_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2826_y0);
  and_gate and_gate_h_u_cla32_and2827_y0(h_u_cla32_and2826_y0, h_u_cla32_and2825_y0, h_u_cla32_and2827_y0);
  and_gate and_gate_h_u_cla32_and2828_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2828_y0);
  and_gate and_gate_h_u_cla32_and2829_y0(h_u_cla32_and2828_y0, h_u_cla32_and2827_y0, h_u_cla32_and2829_y0);
  and_gate and_gate_h_u_cla32_and2830_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2830_y0);
  and_gate and_gate_h_u_cla32_and2831_y0(h_u_cla32_and2830_y0, h_u_cla32_and2829_y0, h_u_cla32_and2831_y0);
  and_gate and_gate_h_u_cla32_and2832_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and2832_y0);
  and_gate and_gate_h_u_cla32_and2833_y0(h_u_cla32_and2832_y0, h_u_cla32_and2831_y0, h_u_cla32_and2833_y0);
  and_gate and_gate_h_u_cla32_and2834_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2834_y0);
  and_gate and_gate_h_u_cla32_and2835_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2835_y0);
  and_gate and_gate_h_u_cla32_and2836_y0(h_u_cla32_and2835_y0, h_u_cla32_and2834_y0, h_u_cla32_and2836_y0);
  and_gate and_gate_h_u_cla32_and2837_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2837_y0);
  and_gate and_gate_h_u_cla32_and2838_y0(h_u_cla32_and2837_y0, h_u_cla32_and2836_y0, h_u_cla32_and2838_y0);
  and_gate and_gate_h_u_cla32_and2839_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2839_y0);
  and_gate and_gate_h_u_cla32_and2840_y0(h_u_cla32_and2839_y0, h_u_cla32_and2838_y0, h_u_cla32_and2840_y0);
  and_gate and_gate_h_u_cla32_and2841_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2841_y0);
  and_gate and_gate_h_u_cla32_and2842_y0(h_u_cla32_and2841_y0, h_u_cla32_and2840_y0, h_u_cla32_and2842_y0);
  and_gate and_gate_h_u_cla32_and2843_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and2843_y0);
  and_gate and_gate_h_u_cla32_and2844_y0(h_u_cla32_and2843_y0, h_u_cla32_and2842_y0, h_u_cla32_and2844_y0);
  and_gate and_gate_h_u_cla32_and2845_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2845_y0);
  and_gate and_gate_h_u_cla32_and2846_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2846_y0);
  and_gate and_gate_h_u_cla32_and2847_y0(h_u_cla32_and2846_y0, h_u_cla32_and2845_y0, h_u_cla32_and2847_y0);
  and_gate and_gate_h_u_cla32_and2848_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2848_y0);
  and_gate and_gate_h_u_cla32_and2849_y0(h_u_cla32_and2848_y0, h_u_cla32_and2847_y0, h_u_cla32_and2849_y0);
  and_gate and_gate_h_u_cla32_and2850_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2850_y0);
  and_gate and_gate_h_u_cla32_and2851_y0(h_u_cla32_and2850_y0, h_u_cla32_and2849_y0, h_u_cla32_and2851_y0);
  and_gate and_gate_h_u_cla32_and2852_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and2852_y0);
  and_gate and_gate_h_u_cla32_and2853_y0(h_u_cla32_and2852_y0, h_u_cla32_and2851_y0, h_u_cla32_and2853_y0);
  and_gate and_gate_h_u_cla32_and2854_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2854_y0);
  and_gate and_gate_h_u_cla32_and2855_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2855_y0);
  and_gate and_gate_h_u_cla32_and2856_y0(h_u_cla32_and2855_y0, h_u_cla32_and2854_y0, h_u_cla32_and2856_y0);
  and_gate and_gate_h_u_cla32_and2857_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2857_y0);
  and_gate and_gate_h_u_cla32_and2858_y0(h_u_cla32_and2857_y0, h_u_cla32_and2856_y0, h_u_cla32_and2858_y0);
  and_gate and_gate_h_u_cla32_and2859_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and2859_y0);
  and_gate and_gate_h_u_cla32_and2860_y0(h_u_cla32_and2859_y0, h_u_cla32_and2858_y0, h_u_cla32_and2860_y0);
  and_gate and_gate_h_u_cla32_and2861_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and2861_y0);
  and_gate and_gate_h_u_cla32_and2862_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and2862_y0);
  and_gate and_gate_h_u_cla32_and2863_y0(h_u_cla32_and2862_y0, h_u_cla32_and2861_y0, h_u_cla32_and2863_y0);
  and_gate and_gate_h_u_cla32_and2864_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and2864_y0);
  and_gate and_gate_h_u_cla32_and2865_y0(h_u_cla32_and2864_y0, h_u_cla32_and2863_y0, h_u_cla32_and2865_y0);
  and_gate and_gate_h_u_cla32_and2866_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and2866_y0);
  and_gate and_gate_h_u_cla32_and2867_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and2867_y0);
  and_gate and_gate_h_u_cla32_and2868_y0(h_u_cla32_and2867_y0, h_u_cla32_and2866_y0, h_u_cla32_and2868_y0);
  and_gate and_gate_h_u_cla32_and2869_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and2869_y0);
  or_gate or_gate_h_u_cla32_or190_y0(h_u_cla32_and2869_y0, h_u_cla32_and2508_y0, h_u_cla32_or190_y0);
  or_gate or_gate_h_u_cla32_or191_y0(h_u_cla32_or190_y0, h_u_cla32_and2545_y0, h_u_cla32_or191_y0);
  or_gate or_gate_h_u_cla32_or192_y0(h_u_cla32_or191_y0, h_u_cla32_and2580_y0, h_u_cla32_or192_y0);
  or_gate or_gate_h_u_cla32_or193_y0(h_u_cla32_or192_y0, h_u_cla32_and2613_y0, h_u_cla32_or193_y0);
  or_gate or_gate_h_u_cla32_or194_y0(h_u_cla32_or193_y0, h_u_cla32_and2644_y0, h_u_cla32_or194_y0);
  or_gate or_gate_h_u_cla32_or195_y0(h_u_cla32_or194_y0, h_u_cla32_and2673_y0, h_u_cla32_or195_y0);
  or_gate or_gate_h_u_cla32_or196_y0(h_u_cla32_or195_y0, h_u_cla32_and2700_y0, h_u_cla32_or196_y0);
  or_gate or_gate_h_u_cla32_or197_y0(h_u_cla32_or196_y0, h_u_cla32_and2725_y0, h_u_cla32_or197_y0);
  or_gate or_gate_h_u_cla32_or198_y0(h_u_cla32_or197_y0, h_u_cla32_and2748_y0, h_u_cla32_or198_y0);
  or_gate or_gate_h_u_cla32_or199_y0(h_u_cla32_or198_y0, h_u_cla32_and2769_y0, h_u_cla32_or199_y0);
  or_gate or_gate_h_u_cla32_or200_y0(h_u_cla32_or199_y0, h_u_cla32_and2788_y0, h_u_cla32_or200_y0);
  or_gate or_gate_h_u_cla32_or201_y0(h_u_cla32_or200_y0, h_u_cla32_and2805_y0, h_u_cla32_or201_y0);
  or_gate or_gate_h_u_cla32_or202_y0(h_u_cla32_or201_y0, h_u_cla32_and2820_y0, h_u_cla32_or202_y0);
  or_gate or_gate_h_u_cla32_or203_y0(h_u_cla32_or202_y0, h_u_cla32_and2833_y0, h_u_cla32_or203_y0);
  or_gate or_gate_h_u_cla32_or204_y0(h_u_cla32_or203_y0, h_u_cla32_and2844_y0, h_u_cla32_or204_y0);
  or_gate or_gate_h_u_cla32_or205_y0(h_u_cla32_or204_y0, h_u_cla32_and2853_y0, h_u_cla32_or205_y0);
  or_gate or_gate_h_u_cla32_or206_y0(h_u_cla32_or205_y0, h_u_cla32_and2860_y0, h_u_cla32_or206_y0);
  or_gate or_gate_h_u_cla32_or207_y0(h_u_cla32_or206_y0, h_u_cla32_and2865_y0, h_u_cla32_or207_y0);
  or_gate or_gate_h_u_cla32_or208_y0(h_u_cla32_or207_y0, h_u_cla32_and2868_y0, h_u_cla32_or208_y0);
  or_gate or_gate_h_u_cla32_or209_y0(h_u_cla32_pg_logic19_y1, h_u_cla32_or208_y0, h_u_cla32_or209_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic20_y0(a_20, b_20, h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_pg_logic20_y2);
  xor_gate xor_gate_h_u_cla32_xor20_y0(h_u_cla32_pg_logic20_y2, h_u_cla32_or209_y0, h_u_cla32_xor20_y0);
  and_gate and_gate_h_u_cla32_and2870_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and2870_y0);
  and_gate and_gate_h_u_cla32_and2871_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and2871_y0);
  and_gate and_gate_h_u_cla32_and2872_y0(h_u_cla32_and2871_y0, h_u_cla32_and2870_y0, h_u_cla32_and2872_y0);
  and_gate and_gate_h_u_cla32_and2873_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and2873_y0);
  and_gate and_gate_h_u_cla32_and2874_y0(h_u_cla32_and2873_y0, h_u_cla32_and2872_y0, h_u_cla32_and2874_y0);
  and_gate and_gate_h_u_cla32_and2875_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and2875_y0);
  and_gate and_gate_h_u_cla32_and2876_y0(h_u_cla32_and2875_y0, h_u_cla32_and2874_y0, h_u_cla32_and2876_y0);
  and_gate and_gate_h_u_cla32_and2877_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and2877_y0);
  and_gate and_gate_h_u_cla32_and2878_y0(h_u_cla32_and2877_y0, h_u_cla32_and2876_y0, h_u_cla32_and2878_y0);
  and_gate and_gate_h_u_cla32_and2879_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and2879_y0);
  and_gate and_gate_h_u_cla32_and2880_y0(h_u_cla32_and2879_y0, h_u_cla32_and2878_y0, h_u_cla32_and2880_y0);
  and_gate and_gate_h_u_cla32_and2881_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and2881_y0);
  and_gate and_gate_h_u_cla32_and2882_y0(h_u_cla32_and2881_y0, h_u_cla32_and2880_y0, h_u_cla32_and2882_y0);
  and_gate and_gate_h_u_cla32_and2883_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and2883_y0);
  and_gate and_gate_h_u_cla32_and2884_y0(h_u_cla32_and2883_y0, h_u_cla32_and2882_y0, h_u_cla32_and2884_y0);
  and_gate and_gate_h_u_cla32_and2885_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and2885_y0);
  and_gate and_gate_h_u_cla32_and2886_y0(h_u_cla32_and2885_y0, h_u_cla32_and2884_y0, h_u_cla32_and2886_y0);
  and_gate and_gate_h_u_cla32_and2887_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and2887_y0);
  and_gate and_gate_h_u_cla32_and2888_y0(h_u_cla32_and2887_y0, h_u_cla32_and2886_y0, h_u_cla32_and2888_y0);
  and_gate and_gate_h_u_cla32_and2889_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and2889_y0);
  and_gate and_gate_h_u_cla32_and2890_y0(h_u_cla32_and2889_y0, h_u_cla32_and2888_y0, h_u_cla32_and2890_y0);
  and_gate and_gate_h_u_cla32_and2891_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and2891_y0);
  and_gate and_gate_h_u_cla32_and2892_y0(h_u_cla32_and2891_y0, h_u_cla32_and2890_y0, h_u_cla32_and2892_y0);
  and_gate and_gate_h_u_cla32_and2893_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and2893_y0);
  and_gate and_gate_h_u_cla32_and2894_y0(h_u_cla32_and2893_y0, h_u_cla32_and2892_y0, h_u_cla32_and2894_y0);
  and_gate and_gate_h_u_cla32_and2895_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and2895_y0);
  and_gate and_gate_h_u_cla32_and2896_y0(h_u_cla32_and2895_y0, h_u_cla32_and2894_y0, h_u_cla32_and2896_y0);
  and_gate and_gate_h_u_cla32_and2897_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and2897_y0);
  and_gate and_gate_h_u_cla32_and2898_y0(h_u_cla32_and2897_y0, h_u_cla32_and2896_y0, h_u_cla32_and2898_y0);
  and_gate and_gate_h_u_cla32_and2899_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and2899_y0);
  and_gate and_gate_h_u_cla32_and2900_y0(h_u_cla32_and2899_y0, h_u_cla32_and2898_y0, h_u_cla32_and2900_y0);
  and_gate and_gate_h_u_cla32_and2901_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and2901_y0);
  and_gate and_gate_h_u_cla32_and2902_y0(h_u_cla32_and2901_y0, h_u_cla32_and2900_y0, h_u_cla32_and2902_y0);
  and_gate and_gate_h_u_cla32_and2903_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and2903_y0);
  and_gate and_gate_h_u_cla32_and2904_y0(h_u_cla32_and2903_y0, h_u_cla32_and2902_y0, h_u_cla32_and2904_y0);
  and_gate and_gate_h_u_cla32_and2905_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and2905_y0);
  and_gate and_gate_h_u_cla32_and2906_y0(h_u_cla32_and2905_y0, h_u_cla32_and2904_y0, h_u_cla32_and2906_y0);
  and_gate and_gate_h_u_cla32_and2907_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and2907_y0);
  and_gate and_gate_h_u_cla32_and2908_y0(h_u_cla32_and2907_y0, h_u_cla32_and2906_y0, h_u_cla32_and2908_y0);
  and_gate and_gate_h_u_cla32_and2909_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and2909_y0);
  and_gate and_gate_h_u_cla32_and2910_y0(h_u_cla32_and2909_y0, h_u_cla32_and2908_y0, h_u_cla32_and2910_y0);
  and_gate and_gate_h_u_cla32_and2911_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2911_y0);
  and_gate and_gate_h_u_cla32_and2912_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2912_y0);
  and_gate and_gate_h_u_cla32_and2913_y0(h_u_cla32_and2912_y0, h_u_cla32_and2911_y0, h_u_cla32_and2913_y0);
  and_gate and_gate_h_u_cla32_and2914_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2914_y0);
  and_gate and_gate_h_u_cla32_and2915_y0(h_u_cla32_and2914_y0, h_u_cla32_and2913_y0, h_u_cla32_and2915_y0);
  and_gate and_gate_h_u_cla32_and2916_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2916_y0);
  and_gate and_gate_h_u_cla32_and2917_y0(h_u_cla32_and2916_y0, h_u_cla32_and2915_y0, h_u_cla32_and2917_y0);
  and_gate and_gate_h_u_cla32_and2918_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2918_y0);
  and_gate and_gate_h_u_cla32_and2919_y0(h_u_cla32_and2918_y0, h_u_cla32_and2917_y0, h_u_cla32_and2919_y0);
  and_gate and_gate_h_u_cla32_and2920_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2920_y0);
  and_gate and_gate_h_u_cla32_and2921_y0(h_u_cla32_and2920_y0, h_u_cla32_and2919_y0, h_u_cla32_and2921_y0);
  and_gate and_gate_h_u_cla32_and2922_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2922_y0);
  and_gate and_gate_h_u_cla32_and2923_y0(h_u_cla32_and2922_y0, h_u_cla32_and2921_y0, h_u_cla32_and2923_y0);
  and_gate and_gate_h_u_cla32_and2924_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2924_y0);
  and_gate and_gate_h_u_cla32_and2925_y0(h_u_cla32_and2924_y0, h_u_cla32_and2923_y0, h_u_cla32_and2925_y0);
  and_gate and_gate_h_u_cla32_and2926_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2926_y0);
  and_gate and_gate_h_u_cla32_and2927_y0(h_u_cla32_and2926_y0, h_u_cla32_and2925_y0, h_u_cla32_and2927_y0);
  and_gate and_gate_h_u_cla32_and2928_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2928_y0);
  and_gate and_gate_h_u_cla32_and2929_y0(h_u_cla32_and2928_y0, h_u_cla32_and2927_y0, h_u_cla32_and2929_y0);
  and_gate and_gate_h_u_cla32_and2930_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2930_y0);
  and_gate and_gate_h_u_cla32_and2931_y0(h_u_cla32_and2930_y0, h_u_cla32_and2929_y0, h_u_cla32_and2931_y0);
  and_gate and_gate_h_u_cla32_and2932_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2932_y0);
  and_gate and_gate_h_u_cla32_and2933_y0(h_u_cla32_and2932_y0, h_u_cla32_and2931_y0, h_u_cla32_and2933_y0);
  and_gate and_gate_h_u_cla32_and2934_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2934_y0);
  and_gate and_gate_h_u_cla32_and2935_y0(h_u_cla32_and2934_y0, h_u_cla32_and2933_y0, h_u_cla32_and2935_y0);
  and_gate and_gate_h_u_cla32_and2936_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2936_y0);
  and_gate and_gate_h_u_cla32_and2937_y0(h_u_cla32_and2936_y0, h_u_cla32_and2935_y0, h_u_cla32_and2937_y0);
  and_gate and_gate_h_u_cla32_and2938_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2938_y0);
  and_gate and_gate_h_u_cla32_and2939_y0(h_u_cla32_and2938_y0, h_u_cla32_and2937_y0, h_u_cla32_and2939_y0);
  and_gate and_gate_h_u_cla32_and2940_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2940_y0);
  and_gate and_gate_h_u_cla32_and2941_y0(h_u_cla32_and2940_y0, h_u_cla32_and2939_y0, h_u_cla32_and2941_y0);
  and_gate and_gate_h_u_cla32_and2942_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2942_y0);
  and_gate and_gate_h_u_cla32_and2943_y0(h_u_cla32_and2942_y0, h_u_cla32_and2941_y0, h_u_cla32_and2943_y0);
  and_gate and_gate_h_u_cla32_and2944_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2944_y0);
  and_gate and_gate_h_u_cla32_and2945_y0(h_u_cla32_and2944_y0, h_u_cla32_and2943_y0, h_u_cla32_and2945_y0);
  and_gate and_gate_h_u_cla32_and2946_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2946_y0);
  and_gate and_gate_h_u_cla32_and2947_y0(h_u_cla32_and2946_y0, h_u_cla32_and2945_y0, h_u_cla32_and2947_y0);
  and_gate and_gate_h_u_cla32_and2948_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and2948_y0);
  and_gate and_gate_h_u_cla32_and2949_y0(h_u_cla32_and2948_y0, h_u_cla32_and2947_y0, h_u_cla32_and2949_y0);
  and_gate and_gate_h_u_cla32_and2950_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2950_y0);
  and_gate and_gate_h_u_cla32_and2951_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2951_y0);
  and_gate and_gate_h_u_cla32_and2952_y0(h_u_cla32_and2951_y0, h_u_cla32_and2950_y0, h_u_cla32_and2952_y0);
  and_gate and_gate_h_u_cla32_and2953_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2953_y0);
  and_gate and_gate_h_u_cla32_and2954_y0(h_u_cla32_and2953_y0, h_u_cla32_and2952_y0, h_u_cla32_and2954_y0);
  and_gate and_gate_h_u_cla32_and2955_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2955_y0);
  and_gate and_gate_h_u_cla32_and2956_y0(h_u_cla32_and2955_y0, h_u_cla32_and2954_y0, h_u_cla32_and2956_y0);
  and_gate and_gate_h_u_cla32_and2957_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2957_y0);
  and_gate and_gate_h_u_cla32_and2958_y0(h_u_cla32_and2957_y0, h_u_cla32_and2956_y0, h_u_cla32_and2958_y0);
  and_gate and_gate_h_u_cla32_and2959_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2959_y0);
  and_gate and_gate_h_u_cla32_and2960_y0(h_u_cla32_and2959_y0, h_u_cla32_and2958_y0, h_u_cla32_and2960_y0);
  and_gate and_gate_h_u_cla32_and2961_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2961_y0);
  and_gate and_gate_h_u_cla32_and2962_y0(h_u_cla32_and2961_y0, h_u_cla32_and2960_y0, h_u_cla32_and2962_y0);
  and_gate and_gate_h_u_cla32_and2963_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2963_y0);
  and_gate and_gate_h_u_cla32_and2964_y0(h_u_cla32_and2963_y0, h_u_cla32_and2962_y0, h_u_cla32_and2964_y0);
  and_gate and_gate_h_u_cla32_and2965_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2965_y0);
  and_gate and_gate_h_u_cla32_and2966_y0(h_u_cla32_and2965_y0, h_u_cla32_and2964_y0, h_u_cla32_and2966_y0);
  and_gate and_gate_h_u_cla32_and2967_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2967_y0);
  and_gate and_gate_h_u_cla32_and2968_y0(h_u_cla32_and2967_y0, h_u_cla32_and2966_y0, h_u_cla32_and2968_y0);
  and_gate and_gate_h_u_cla32_and2969_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2969_y0);
  and_gate and_gate_h_u_cla32_and2970_y0(h_u_cla32_and2969_y0, h_u_cla32_and2968_y0, h_u_cla32_and2970_y0);
  and_gate and_gate_h_u_cla32_and2971_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2971_y0);
  and_gate and_gate_h_u_cla32_and2972_y0(h_u_cla32_and2971_y0, h_u_cla32_and2970_y0, h_u_cla32_and2972_y0);
  and_gate and_gate_h_u_cla32_and2973_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2973_y0);
  and_gate and_gate_h_u_cla32_and2974_y0(h_u_cla32_and2973_y0, h_u_cla32_and2972_y0, h_u_cla32_and2974_y0);
  and_gate and_gate_h_u_cla32_and2975_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2975_y0);
  and_gate and_gate_h_u_cla32_and2976_y0(h_u_cla32_and2975_y0, h_u_cla32_and2974_y0, h_u_cla32_and2976_y0);
  and_gate and_gate_h_u_cla32_and2977_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2977_y0);
  and_gate and_gate_h_u_cla32_and2978_y0(h_u_cla32_and2977_y0, h_u_cla32_and2976_y0, h_u_cla32_and2978_y0);
  and_gate and_gate_h_u_cla32_and2979_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2979_y0);
  and_gate and_gate_h_u_cla32_and2980_y0(h_u_cla32_and2979_y0, h_u_cla32_and2978_y0, h_u_cla32_and2980_y0);
  and_gate and_gate_h_u_cla32_and2981_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2981_y0);
  and_gate and_gate_h_u_cla32_and2982_y0(h_u_cla32_and2981_y0, h_u_cla32_and2980_y0, h_u_cla32_and2982_y0);
  and_gate and_gate_h_u_cla32_and2983_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2983_y0);
  and_gate and_gate_h_u_cla32_and2984_y0(h_u_cla32_and2983_y0, h_u_cla32_and2982_y0, h_u_cla32_and2984_y0);
  and_gate and_gate_h_u_cla32_and2985_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and2985_y0);
  and_gate and_gate_h_u_cla32_and2986_y0(h_u_cla32_and2985_y0, h_u_cla32_and2984_y0, h_u_cla32_and2986_y0);
  and_gate and_gate_h_u_cla32_and2987_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2987_y0);
  and_gate and_gate_h_u_cla32_and2988_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2988_y0);
  and_gate and_gate_h_u_cla32_and2989_y0(h_u_cla32_and2988_y0, h_u_cla32_and2987_y0, h_u_cla32_and2989_y0);
  and_gate and_gate_h_u_cla32_and2990_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2990_y0);
  and_gate and_gate_h_u_cla32_and2991_y0(h_u_cla32_and2990_y0, h_u_cla32_and2989_y0, h_u_cla32_and2991_y0);
  and_gate and_gate_h_u_cla32_and2992_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2992_y0);
  and_gate and_gate_h_u_cla32_and2993_y0(h_u_cla32_and2992_y0, h_u_cla32_and2991_y0, h_u_cla32_and2993_y0);
  and_gate and_gate_h_u_cla32_and2994_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2994_y0);
  and_gate and_gate_h_u_cla32_and2995_y0(h_u_cla32_and2994_y0, h_u_cla32_and2993_y0, h_u_cla32_and2995_y0);
  and_gate and_gate_h_u_cla32_and2996_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2996_y0);
  and_gate and_gate_h_u_cla32_and2997_y0(h_u_cla32_and2996_y0, h_u_cla32_and2995_y0, h_u_cla32_and2997_y0);
  and_gate and_gate_h_u_cla32_and2998_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and2998_y0);
  and_gate and_gate_h_u_cla32_and2999_y0(h_u_cla32_and2998_y0, h_u_cla32_and2997_y0, h_u_cla32_and2999_y0);
  and_gate and_gate_h_u_cla32_and3000_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3000_y0);
  and_gate and_gate_h_u_cla32_and3001_y0(h_u_cla32_and3000_y0, h_u_cla32_and2999_y0, h_u_cla32_and3001_y0);
  and_gate and_gate_h_u_cla32_and3002_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3002_y0);
  and_gate and_gate_h_u_cla32_and3003_y0(h_u_cla32_and3002_y0, h_u_cla32_and3001_y0, h_u_cla32_and3003_y0);
  and_gate and_gate_h_u_cla32_and3004_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3004_y0);
  and_gate and_gate_h_u_cla32_and3005_y0(h_u_cla32_and3004_y0, h_u_cla32_and3003_y0, h_u_cla32_and3005_y0);
  and_gate and_gate_h_u_cla32_and3006_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3006_y0);
  and_gate and_gate_h_u_cla32_and3007_y0(h_u_cla32_and3006_y0, h_u_cla32_and3005_y0, h_u_cla32_and3007_y0);
  and_gate and_gate_h_u_cla32_and3008_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3008_y0);
  and_gate and_gate_h_u_cla32_and3009_y0(h_u_cla32_and3008_y0, h_u_cla32_and3007_y0, h_u_cla32_and3009_y0);
  and_gate and_gate_h_u_cla32_and3010_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3010_y0);
  and_gate and_gate_h_u_cla32_and3011_y0(h_u_cla32_and3010_y0, h_u_cla32_and3009_y0, h_u_cla32_and3011_y0);
  and_gate and_gate_h_u_cla32_and3012_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3012_y0);
  and_gate and_gate_h_u_cla32_and3013_y0(h_u_cla32_and3012_y0, h_u_cla32_and3011_y0, h_u_cla32_and3013_y0);
  and_gate and_gate_h_u_cla32_and3014_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3014_y0);
  and_gate and_gate_h_u_cla32_and3015_y0(h_u_cla32_and3014_y0, h_u_cla32_and3013_y0, h_u_cla32_and3015_y0);
  and_gate and_gate_h_u_cla32_and3016_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3016_y0);
  and_gate and_gate_h_u_cla32_and3017_y0(h_u_cla32_and3016_y0, h_u_cla32_and3015_y0, h_u_cla32_and3017_y0);
  and_gate and_gate_h_u_cla32_and3018_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3018_y0);
  and_gate and_gate_h_u_cla32_and3019_y0(h_u_cla32_and3018_y0, h_u_cla32_and3017_y0, h_u_cla32_and3019_y0);
  and_gate and_gate_h_u_cla32_and3020_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3020_y0);
  and_gate and_gate_h_u_cla32_and3021_y0(h_u_cla32_and3020_y0, h_u_cla32_and3019_y0, h_u_cla32_and3021_y0);
  and_gate and_gate_h_u_cla32_and3022_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3022_y0);
  and_gate and_gate_h_u_cla32_and3023_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3023_y0);
  and_gate and_gate_h_u_cla32_and3024_y0(h_u_cla32_and3023_y0, h_u_cla32_and3022_y0, h_u_cla32_and3024_y0);
  and_gate and_gate_h_u_cla32_and3025_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3025_y0);
  and_gate and_gate_h_u_cla32_and3026_y0(h_u_cla32_and3025_y0, h_u_cla32_and3024_y0, h_u_cla32_and3026_y0);
  and_gate and_gate_h_u_cla32_and3027_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3027_y0);
  and_gate and_gate_h_u_cla32_and3028_y0(h_u_cla32_and3027_y0, h_u_cla32_and3026_y0, h_u_cla32_and3028_y0);
  and_gate and_gate_h_u_cla32_and3029_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3029_y0);
  and_gate and_gate_h_u_cla32_and3030_y0(h_u_cla32_and3029_y0, h_u_cla32_and3028_y0, h_u_cla32_and3030_y0);
  and_gate and_gate_h_u_cla32_and3031_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3031_y0);
  and_gate and_gate_h_u_cla32_and3032_y0(h_u_cla32_and3031_y0, h_u_cla32_and3030_y0, h_u_cla32_and3032_y0);
  and_gate and_gate_h_u_cla32_and3033_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3033_y0);
  and_gate and_gate_h_u_cla32_and3034_y0(h_u_cla32_and3033_y0, h_u_cla32_and3032_y0, h_u_cla32_and3034_y0);
  and_gate and_gate_h_u_cla32_and3035_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3035_y0);
  and_gate and_gate_h_u_cla32_and3036_y0(h_u_cla32_and3035_y0, h_u_cla32_and3034_y0, h_u_cla32_and3036_y0);
  and_gate and_gate_h_u_cla32_and3037_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3037_y0);
  and_gate and_gate_h_u_cla32_and3038_y0(h_u_cla32_and3037_y0, h_u_cla32_and3036_y0, h_u_cla32_and3038_y0);
  and_gate and_gate_h_u_cla32_and3039_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3039_y0);
  and_gate and_gate_h_u_cla32_and3040_y0(h_u_cla32_and3039_y0, h_u_cla32_and3038_y0, h_u_cla32_and3040_y0);
  and_gate and_gate_h_u_cla32_and3041_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3041_y0);
  and_gate and_gate_h_u_cla32_and3042_y0(h_u_cla32_and3041_y0, h_u_cla32_and3040_y0, h_u_cla32_and3042_y0);
  and_gate and_gate_h_u_cla32_and3043_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3043_y0);
  and_gate and_gate_h_u_cla32_and3044_y0(h_u_cla32_and3043_y0, h_u_cla32_and3042_y0, h_u_cla32_and3044_y0);
  and_gate and_gate_h_u_cla32_and3045_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3045_y0);
  and_gate and_gate_h_u_cla32_and3046_y0(h_u_cla32_and3045_y0, h_u_cla32_and3044_y0, h_u_cla32_and3046_y0);
  and_gate and_gate_h_u_cla32_and3047_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3047_y0);
  and_gate and_gate_h_u_cla32_and3048_y0(h_u_cla32_and3047_y0, h_u_cla32_and3046_y0, h_u_cla32_and3048_y0);
  and_gate and_gate_h_u_cla32_and3049_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3049_y0);
  and_gate and_gate_h_u_cla32_and3050_y0(h_u_cla32_and3049_y0, h_u_cla32_and3048_y0, h_u_cla32_and3050_y0);
  and_gate and_gate_h_u_cla32_and3051_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3051_y0);
  and_gate and_gate_h_u_cla32_and3052_y0(h_u_cla32_and3051_y0, h_u_cla32_and3050_y0, h_u_cla32_and3052_y0);
  and_gate and_gate_h_u_cla32_and3053_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3053_y0);
  and_gate and_gate_h_u_cla32_and3054_y0(h_u_cla32_and3053_y0, h_u_cla32_and3052_y0, h_u_cla32_and3054_y0);
  and_gate and_gate_h_u_cla32_and3055_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3055_y0);
  and_gate and_gate_h_u_cla32_and3056_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3056_y0);
  and_gate and_gate_h_u_cla32_and3057_y0(h_u_cla32_and3056_y0, h_u_cla32_and3055_y0, h_u_cla32_and3057_y0);
  and_gate and_gate_h_u_cla32_and3058_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3058_y0);
  and_gate and_gate_h_u_cla32_and3059_y0(h_u_cla32_and3058_y0, h_u_cla32_and3057_y0, h_u_cla32_and3059_y0);
  and_gate and_gate_h_u_cla32_and3060_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3060_y0);
  and_gate and_gate_h_u_cla32_and3061_y0(h_u_cla32_and3060_y0, h_u_cla32_and3059_y0, h_u_cla32_and3061_y0);
  and_gate and_gate_h_u_cla32_and3062_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3062_y0);
  and_gate and_gate_h_u_cla32_and3063_y0(h_u_cla32_and3062_y0, h_u_cla32_and3061_y0, h_u_cla32_and3063_y0);
  and_gate and_gate_h_u_cla32_and3064_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3064_y0);
  and_gate and_gate_h_u_cla32_and3065_y0(h_u_cla32_and3064_y0, h_u_cla32_and3063_y0, h_u_cla32_and3065_y0);
  and_gate and_gate_h_u_cla32_and3066_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3066_y0);
  and_gate and_gate_h_u_cla32_and3067_y0(h_u_cla32_and3066_y0, h_u_cla32_and3065_y0, h_u_cla32_and3067_y0);
  and_gate and_gate_h_u_cla32_and3068_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3068_y0);
  and_gate and_gate_h_u_cla32_and3069_y0(h_u_cla32_and3068_y0, h_u_cla32_and3067_y0, h_u_cla32_and3069_y0);
  and_gate and_gate_h_u_cla32_and3070_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3070_y0);
  and_gate and_gate_h_u_cla32_and3071_y0(h_u_cla32_and3070_y0, h_u_cla32_and3069_y0, h_u_cla32_and3071_y0);
  and_gate and_gate_h_u_cla32_and3072_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3072_y0);
  and_gate and_gate_h_u_cla32_and3073_y0(h_u_cla32_and3072_y0, h_u_cla32_and3071_y0, h_u_cla32_and3073_y0);
  and_gate and_gate_h_u_cla32_and3074_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3074_y0);
  and_gate and_gate_h_u_cla32_and3075_y0(h_u_cla32_and3074_y0, h_u_cla32_and3073_y0, h_u_cla32_and3075_y0);
  and_gate and_gate_h_u_cla32_and3076_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3076_y0);
  and_gate and_gate_h_u_cla32_and3077_y0(h_u_cla32_and3076_y0, h_u_cla32_and3075_y0, h_u_cla32_and3077_y0);
  and_gate and_gate_h_u_cla32_and3078_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3078_y0);
  and_gate and_gate_h_u_cla32_and3079_y0(h_u_cla32_and3078_y0, h_u_cla32_and3077_y0, h_u_cla32_and3079_y0);
  and_gate and_gate_h_u_cla32_and3080_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3080_y0);
  and_gate and_gate_h_u_cla32_and3081_y0(h_u_cla32_and3080_y0, h_u_cla32_and3079_y0, h_u_cla32_and3081_y0);
  and_gate and_gate_h_u_cla32_and3082_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3082_y0);
  and_gate and_gate_h_u_cla32_and3083_y0(h_u_cla32_and3082_y0, h_u_cla32_and3081_y0, h_u_cla32_and3083_y0);
  and_gate and_gate_h_u_cla32_and3084_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3084_y0);
  and_gate and_gate_h_u_cla32_and3085_y0(h_u_cla32_and3084_y0, h_u_cla32_and3083_y0, h_u_cla32_and3085_y0);
  and_gate and_gate_h_u_cla32_and3086_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3086_y0);
  and_gate and_gate_h_u_cla32_and3087_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3087_y0);
  and_gate and_gate_h_u_cla32_and3088_y0(h_u_cla32_and3087_y0, h_u_cla32_and3086_y0, h_u_cla32_and3088_y0);
  and_gate and_gate_h_u_cla32_and3089_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3089_y0);
  and_gate and_gate_h_u_cla32_and3090_y0(h_u_cla32_and3089_y0, h_u_cla32_and3088_y0, h_u_cla32_and3090_y0);
  and_gate and_gate_h_u_cla32_and3091_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3091_y0);
  and_gate and_gate_h_u_cla32_and3092_y0(h_u_cla32_and3091_y0, h_u_cla32_and3090_y0, h_u_cla32_and3092_y0);
  and_gate and_gate_h_u_cla32_and3093_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3093_y0);
  and_gate and_gate_h_u_cla32_and3094_y0(h_u_cla32_and3093_y0, h_u_cla32_and3092_y0, h_u_cla32_and3094_y0);
  and_gate and_gate_h_u_cla32_and3095_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3095_y0);
  and_gate and_gate_h_u_cla32_and3096_y0(h_u_cla32_and3095_y0, h_u_cla32_and3094_y0, h_u_cla32_and3096_y0);
  and_gate and_gate_h_u_cla32_and3097_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3097_y0);
  and_gate and_gate_h_u_cla32_and3098_y0(h_u_cla32_and3097_y0, h_u_cla32_and3096_y0, h_u_cla32_and3098_y0);
  and_gate and_gate_h_u_cla32_and3099_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3099_y0);
  and_gate and_gate_h_u_cla32_and3100_y0(h_u_cla32_and3099_y0, h_u_cla32_and3098_y0, h_u_cla32_and3100_y0);
  and_gate and_gate_h_u_cla32_and3101_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3101_y0);
  and_gate and_gate_h_u_cla32_and3102_y0(h_u_cla32_and3101_y0, h_u_cla32_and3100_y0, h_u_cla32_and3102_y0);
  and_gate and_gate_h_u_cla32_and3103_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3103_y0);
  and_gate and_gate_h_u_cla32_and3104_y0(h_u_cla32_and3103_y0, h_u_cla32_and3102_y0, h_u_cla32_and3104_y0);
  and_gate and_gate_h_u_cla32_and3105_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3105_y0);
  and_gate and_gate_h_u_cla32_and3106_y0(h_u_cla32_and3105_y0, h_u_cla32_and3104_y0, h_u_cla32_and3106_y0);
  and_gate and_gate_h_u_cla32_and3107_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3107_y0);
  and_gate and_gate_h_u_cla32_and3108_y0(h_u_cla32_and3107_y0, h_u_cla32_and3106_y0, h_u_cla32_and3108_y0);
  and_gate and_gate_h_u_cla32_and3109_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3109_y0);
  and_gate and_gate_h_u_cla32_and3110_y0(h_u_cla32_and3109_y0, h_u_cla32_and3108_y0, h_u_cla32_and3110_y0);
  and_gate and_gate_h_u_cla32_and3111_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3111_y0);
  and_gate and_gate_h_u_cla32_and3112_y0(h_u_cla32_and3111_y0, h_u_cla32_and3110_y0, h_u_cla32_and3112_y0);
  and_gate and_gate_h_u_cla32_and3113_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3113_y0);
  and_gate and_gate_h_u_cla32_and3114_y0(h_u_cla32_and3113_y0, h_u_cla32_and3112_y0, h_u_cla32_and3114_y0);
  and_gate and_gate_h_u_cla32_and3115_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3115_y0);
  and_gate and_gate_h_u_cla32_and3116_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3116_y0);
  and_gate and_gate_h_u_cla32_and3117_y0(h_u_cla32_and3116_y0, h_u_cla32_and3115_y0, h_u_cla32_and3117_y0);
  and_gate and_gate_h_u_cla32_and3118_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3118_y0);
  and_gate and_gate_h_u_cla32_and3119_y0(h_u_cla32_and3118_y0, h_u_cla32_and3117_y0, h_u_cla32_and3119_y0);
  and_gate and_gate_h_u_cla32_and3120_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3120_y0);
  and_gate and_gate_h_u_cla32_and3121_y0(h_u_cla32_and3120_y0, h_u_cla32_and3119_y0, h_u_cla32_and3121_y0);
  and_gate and_gate_h_u_cla32_and3122_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3122_y0);
  and_gate and_gate_h_u_cla32_and3123_y0(h_u_cla32_and3122_y0, h_u_cla32_and3121_y0, h_u_cla32_and3123_y0);
  and_gate and_gate_h_u_cla32_and3124_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3124_y0);
  and_gate and_gate_h_u_cla32_and3125_y0(h_u_cla32_and3124_y0, h_u_cla32_and3123_y0, h_u_cla32_and3125_y0);
  and_gate and_gate_h_u_cla32_and3126_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3126_y0);
  and_gate and_gate_h_u_cla32_and3127_y0(h_u_cla32_and3126_y0, h_u_cla32_and3125_y0, h_u_cla32_and3127_y0);
  and_gate and_gate_h_u_cla32_and3128_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3128_y0);
  and_gate and_gate_h_u_cla32_and3129_y0(h_u_cla32_and3128_y0, h_u_cla32_and3127_y0, h_u_cla32_and3129_y0);
  and_gate and_gate_h_u_cla32_and3130_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3130_y0);
  and_gate and_gate_h_u_cla32_and3131_y0(h_u_cla32_and3130_y0, h_u_cla32_and3129_y0, h_u_cla32_and3131_y0);
  and_gate and_gate_h_u_cla32_and3132_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3132_y0);
  and_gate and_gate_h_u_cla32_and3133_y0(h_u_cla32_and3132_y0, h_u_cla32_and3131_y0, h_u_cla32_and3133_y0);
  and_gate and_gate_h_u_cla32_and3134_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3134_y0);
  and_gate and_gate_h_u_cla32_and3135_y0(h_u_cla32_and3134_y0, h_u_cla32_and3133_y0, h_u_cla32_and3135_y0);
  and_gate and_gate_h_u_cla32_and3136_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3136_y0);
  and_gate and_gate_h_u_cla32_and3137_y0(h_u_cla32_and3136_y0, h_u_cla32_and3135_y0, h_u_cla32_and3137_y0);
  and_gate and_gate_h_u_cla32_and3138_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3138_y0);
  and_gate and_gate_h_u_cla32_and3139_y0(h_u_cla32_and3138_y0, h_u_cla32_and3137_y0, h_u_cla32_and3139_y0);
  and_gate and_gate_h_u_cla32_and3140_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3140_y0);
  and_gate and_gate_h_u_cla32_and3141_y0(h_u_cla32_and3140_y0, h_u_cla32_and3139_y0, h_u_cla32_and3141_y0);
  and_gate and_gate_h_u_cla32_and3142_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3142_y0);
  and_gate and_gate_h_u_cla32_and3143_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3143_y0);
  and_gate and_gate_h_u_cla32_and3144_y0(h_u_cla32_and3143_y0, h_u_cla32_and3142_y0, h_u_cla32_and3144_y0);
  and_gate and_gate_h_u_cla32_and3145_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3145_y0);
  and_gate and_gate_h_u_cla32_and3146_y0(h_u_cla32_and3145_y0, h_u_cla32_and3144_y0, h_u_cla32_and3146_y0);
  and_gate and_gate_h_u_cla32_and3147_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3147_y0);
  and_gate and_gate_h_u_cla32_and3148_y0(h_u_cla32_and3147_y0, h_u_cla32_and3146_y0, h_u_cla32_and3148_y0);
  and_gate and_gate_h_u_cla32_and3149_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3149_y0);
  and_gate and_gate_h_u_cla32_and3150_y0(h_u_cla32_and3149_y0, h_u_cla32_and3148_y0, h_u_cla32_and3150_y0);
  and_gate and_gate_h_u_cla32_and3151_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3151_y0);
  and_gate and_gate_h_u_cla32_and3152_y0(h_u_cla32_and3151_y0, h_u_cla32_and3150_y0, h_u_cla32_and3152_y0);
  and_gate and_gate_h_u_cla32_and3153_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3153_y0);
  and_gate and_gate_h_u_cla32_and3154_y0(h_u_cla32_and3153_y0, h_u_cla32_and3152_y0, h_u_cla32_and3154_y0);
  and_gate and_gate_h_u_cla32_and3155_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3155_y0);
  and_gate and_gate_h_u_cla32_and3156_y0(h_u_cla32_and3155_y0, h_u_cla32_and3154_y0, h_u_cla32_and3156_y0);
  and_gate and_gate_h_u_cla32_and3157_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3157_y0);
  and_gate and_gate_h_u_cla32_and3158_y0(h_u_cla32_and3157_y0, h_u_cla32_and3156_y0, h_u_cla32_and3158_y0);
  and_gate and_gate_h_u_cla32_and3159_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3159_y0);
  and_gate and_gate_h_u_cla32_and3160_y0(h_u_cla32_and3159_y0, h_u_cla32_and3158_y0, h_u_cla32_and3160_y0);
  and_gate and_gate_h_u_cla32_and3161_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3161_y0);
  and_gate and_gate_h_u_cla32_and3162_y0(h_u_cla32_and3161_y0, h_u_cla32_and3160_y0, h_u_cla32_and3162_y0);
  and_gate and_gate_h_u_cla32_and3163_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3163_y0);
  and_gate and_gate_h_u_cla32_and3164_y0(h_u_cla32_and3163_y0, h_u_cla32_and3162_y0, h_u_cla32_and3164_y0);
  and_gate and_gate_h_u_cla32_and3165_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3165_y0);
  and_gate and_gate_h_u_cla32_and3166_y0(h_u_cla32_and3165_y0, h_u_cla32_and3164_y0, h_u_cla32_and3166_y0);
  and_gate and_gate_h_u_cla32_and3167_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3167_y0);
  and_gate and_gate_h_u_cla32_and3168_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3168_y0);
  and_gate and_gate_h_u_cla32_and3169_y0(h_u_cla32_and3168_y0, h_u_cla32_and3167_y0, h_u_cla32_and3169_y0);
  and_gate and_gate_h_u_cla32_and3170_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3170_y0);
  and_gate and_gate_h_u_cla32_and3171_y0(h_u_cla32_and3170_y0, h_u_cla32_and3169_y0, h_u_cla32_and3171_y0);
  and_gate and_gate_h_u_cla32_and3172_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3172_y0);
  and_gate and_gate_h_u_cla32_and3173_y0(h_u_cla32_and3172_y0, h_u_cla32_and3171_y0, h_u_cla32_and3173_y0);
  and_gate and_gate_h_u_cla32_and3174_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3174_y0);
  and_gate and_gate_h_u_cla32_and3175_y0(h_u_cla32_and3174_y0, h_u_cla32_and3173_y0, h_u_cla32_and3175_y0);
  and_gate and_gate_h_u_cla32_and3176_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3176_y0);
  and_gate and_gate_h_u_cla32_and3177_y0(h_u_cla32_and3176_y0, h_u_cla32_and3175_y0, h_u_cla32_and3177_y0);
  and_gate and_gate_h_u_cla32_and3178_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3178_y0);
  and_gate and_gate_h_u_cla32_and3179_y0(h_u_cla32_and3178_y0, h_u_cla32_and3177_y0, h_u_cla32_and3179_y0);
  and_gate and_gate_h_u_cla32_and3180_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3180_y0);
  and_gate and_gate_h_u_cla32_and3181_y0(h_u_cla32_and3180_y0, h_u_cla32_and3179_y0, h_u_cla32_and3181_y0);
  and_gate and_gate_h_u_cla32_and3182_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3182_y0);
  and_gate and_gate_h_u_cla32_and3183_y0(h_u_cla32_and3182_y0, h_u_cla32_and3181_y0, h_u_cla32_and3183_y0);
  and_gate and_gate_h_u_cla32_and3184_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3184_y0);
  and_gate and_gate_h_u_cla32_and3185_y0(h_u_cla32_and3184_y0, h_u_cla32_and3183_y0, h_u_cla32_and3185_y0);
  and_gate and_gate_h_u_cla32_and3186_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3186_y0);
  and_gate and_gate_h_u_cla32_and3187_y0(h_u_cla32_and3186_y0, h_u_cla32_and3185_y0, h_u_cla32_and3187_y0);
  and_gate and_gate_h_u_cla32_and3188_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3188_y0);
  and_gate and_gate_h_u_cla32_and3189_y0(h_u_cla32_and3188_y0, h_u_cla32_and3187_y0, h_u_cla32_and3189_y0);
  and_gate and_gate_h_u_cla32_and3190_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3190_y0);
  and_gate and_gate_h_u_cla32_and3191_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3191_y0);
  and_gate and_gate_h_u_cla32_and3192_y0(h_u_cla32_and3191_y0, h_u_cla32_and3190_y0, h_u_cla32_and3192_y0);
  and_gate and_gate_h_u_cla32_and3193_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3193_y0);
  and_gate and_gate_h_u_cla32_and3194_y0(h_u_cla32_and3193_y0, h_u_cla32_and3192_y0, h_u_cla32_and3194_y0);
  and_gate and_gate_h_u_cla32_and3195_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3195_y0);
  and_gate and_gate_h_u_cla32_and3196_y0(h_u_cla32_and3195_y0, h_u_cla32_and3194_y0, h_u_cla32_and3196_y0);
  and_gate and_gate_h_u_cla32_and3197_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3197_y0);
  and_gate and_gate_h_u_cla32_and3198_y0(h_u_cla32_and3197_y0, h_u_cla32_and3196_y0, h_u_cla32_and3198_y0);
  and_gate and_gate_h_u_cla32_and3199_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3199_y0);
  and_gate and_gate_h_u_cla32_and3200_y0(h_u_cla32_and3199_y0, h_u_cla32_and3198_y0, h_u_cla32_and3200_y0);
  and_gate and_gate_h_u_cla32_and3201_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3201_y0);
  and_gate and_gate_h_u_cla32_and3202_y0(h_u_cla32_and3201_y0, h_u_cla32_and3200_y0, h_u_cla32_and3202_y0);
  and_gate and_gate_h_u_cla32_and3203_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3203_y0);
  and_gate and_gate_h_u_cla32_and3204_y0(h_u_cla32_and3203_y0, h_u_cla32_and3202_y0, h_u_cla32_and3204_y0);
  and_gate and_gate_h_u_cla32_and3205_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3205_y0);
  and_gate and_gate_h_u_cla32_and3206_y0(h_u_cla32_and3205_y0, h_u_cla32_and3204_y0, h_u_cla32_and3206_y0);
  and_gate and_gate_h_u_cla32_and3207_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3207_y0);
  and_gate and_gate_h_u_cla32_and3208_y0(h_u_cla32_and3207_y0, h_u_cla32_and3206_y0, h_u_cla32_and3208_y0);
  and_gate and_gate_h_u_cla32_and3209_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3209_y0);
  and_gate and_gate_h_u_cla32_and3210_y0(h_u_cla32_and3209_y0, h_u_cla32_and3208_y0, h_u_cla32_and3210_y0);
  and_gate and_gate_h_u_cla32_and3211_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3211_y0);
  and_gate and_gate_h_u_cla32_and3212_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3212_y0);
  and_gate and_gate_h_u_cla32_and3213_y0(h_u_cla32_and3212_y0, h_u_cla32_and3211_y0, h_u_cla32_and3213_y0);
  and_gate and_gate_h_u_cla32_and3214_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3214_y0);
  and_gate and_gate_h_u_cla32_and3215_y0(h_u_cla32_and3214_y0, h_u_cla32_and3213_y0, h_u_cla32_and3215_y0);
  and_gate and_gate_h_u_cla32_and3216_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3216_y0);
  and_gate and_gate_h_u_cla32_and3217_y0(h_u_cla32_and3216_y0, h_u_cla32_and3215_y0, h_u_cla32_and3217_y0);
  and_gate and_gate_h_u_cla32_and3218_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3218_y0);
  and_gate and_gate_h_u_cla32_and3219_y0(h_u_cla32_and3218_y0, h_u_cla32_and3217_y0, h_u_cla32_and3219_y0);
  and_gate and_gate_h_u_cla32_and3220_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3220_y0);
  and_gate and_gate_h_u_cla32_and3221_y0(h_u_cla32_and3220_y0, h_u_cla32_and3219_y0, h_u_cla32_and3221_y0);
  and_gate and_gate_h_u_cla32_and3222_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3222_y0);
  and_gate and_gate_h_u_cla32_and3223_y0(h_u_cla32_and3222_y0, h_u_cla32_and3221_y0, h_u_cla32_and3223_y0);
  and_gate and_gate_h_u_cla32_and3224_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3224_y0);
  and_gate and_gate_h_u_cla32_and3225_y0(h_u_cla32_and3224_y0, h_u_cla32_and3223_y0, h_u_cla32_and3225_y0);
  and_gate and_gate_h_u_cla32_and3226_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3226_y0);
  and_gate and_gate_h_u_cla32_and3227_y0(h_u_cla32_and3226_y0, h_u_cla32_and3225_y0, h_u_cla32_and3227_y0);
  and_gate and_gate_h_u_cla32_and3228_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3228_y0);
  and_gate and_gate_h_u_cla32_and3229_y0(h_u_cla32_and3228_y0, h_u_cla32_and3227_y0, h_u_cla32_and3229_y0);
  and_gate and_gate_h_u_cla32_and3230_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3230_y0);
  and_gate and_gate_h_u_cla32_and3231_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3231_y0);
  and_gate and_gate_h_u_cla32_and3232_y0(h_u_cla32_and3231_y0, h_u_cla32_and3230_y0, h_u_cla32_and3232_y0);
  and_gate and_gate_h_u_cla32_and3233_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3233_y0);
  and_gate and_gate_h_u_cla32_and3234_y0(h_u_cla32_and3233_y0, h_u_cla32_and3232_y0, h_u_cla32_and3234_y0);
  and_gate and_gate_h_u_cla32_and3235_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3235_y0);
  and_gate and_gate_h_u_cla32_and3236_y0(h_u_cla32_and3235_y0, h_u_cla32_and3234_y0, h_u_cla32_and3236_y0);
  and_gate and_gate_h_u_cla32_and3237_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3237_y0);
  and_gate and_gate_h_u_cla32_and3238_y0(h_u_cla32_and3237_y0, h_u_cla32_and3236_y0, h_u_cla32_and3238_y0);
  and_gate and_gate_h_u_cla32_and3239_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3239_y0);
  and_gate and_gate_h_u_cla32_and3240_y0(h_u_cla32_and3239_y0, h_u_cla32_and3238_y0, h_u_cla32_and3240_y0);
  and_gate and_gate_h_u_cla32_and3241_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3241_y0);
  and_gate and_gate_h_u_cla32_and3242_y0(h_u_cla32_and3241_y0, h_u_cla32_and3240_y0, h_u_cla32_and3242_y0);
  and_gate and_gate_h_u_cla32_and3243_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3243_y0);
  and_gate and_gate_h_u_cla32_and3244_y0(h_u_cla32_and3243_y0, h_u_cla32_and3242_y0, h_u_cla32_and3244_y0);
  and_gate and_gate_h_u_cla32_and3245_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3245_y0);
  and_gate and_gate_h_u_cla32_and3246_y0(h_u_cla32_and3245_y0, h_u_cla32_and3244_y0, h_u_cla32_and3246_y0);
  and_gate and_gate_h_u_cla32_and3247_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3247_y0);
  and_gate and_gate_h_u_cla32_and3248_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3248_y0);
  and_gate and_gate_h_u_cla32_and3249_y0(h_u_cla32_and3248_y0, h_u_cla32_and3247_y0, h_u_cla32_and3249_y0);
  and_gate and_gate_h_u_cla32_and3250_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3250_y0);
  and_gate and_gate_h_u_cla32_and3251_y0(h_u_cla32_and3250_y0, h_u_cla32_and3249_y0, h_u_cla32_and3251_y0);
  and_gate and_gate_h_u_cla32_and3252_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3252_y0);
  and_gate and_gate_h_u_cla32_and3253_y0(h_u_cla32_and3252_y0, h_u_cla32_and3251_y0, h_u_cla32_and3253_y0);
  and_gate and_gate_h_u_cla32_and3254_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3254_y0);
  and_gate and_gate_h_u_cla32_and3255_y0(h_u_cla32_and3254_y0, h_u_cla32_and3253_y0, h_u_cla32_and3255_y0);
  and_gate and_gate_h_u_cla32_and3256_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3256_y0);
  and_gate and_gate_h_u_cla32_and3257_y0(h_u_cla32_and3256_y0, h_u_cla32_and3255_y0, h_u_cla32_and3257_y0);
  and_gate and_gate_h_u_cla32_and3258_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3258_y0);
  and_gate and_gate_h_u_cla32_and3259_y0(h_u_cla32_and3258_y0, h_u_cla32_and3257_y0, h_u_cla32_and3259_y0);
  and_gate and_gate_h_u_cla32_and3260_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3260_y0);
  and_gate and_gate_h_u_cla32_and3261_y0(h_u_cla32_and3260_y0, h_u_cla32_and3259_y0, h_u_cla32_and3261_y0);
  and_gate and_gate_h_u_cla32_and3262_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3262_y0);
  and_gate and_gate_h_u_cla32_and3263_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3263_y0);
  and_gate and_gate_h_u_cla32_and3264_y0(h_u_cla32_and3263_y0, h_u_cla32_and3262_y0, h_u_cla32_and3264_y0);
  and_gate and_gate_h_u_cla32_and3265_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3265_y0);
  and_gate and_gate_h_u_cla32_and3266_y0(h_u_cla32_and3265_y0, h_u_cla32_and3264_y0, h_u_cla32_and3266_y0);
  and_gate and_gate_h_u_cla32_and3267_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3267_y0);
  and_gate and_gate_h_u_cla32_and3268_y0(h_u_cla32_and3267_y0, h_u_cla32_and3266_y0, h_u_cla32_and3268_y0);
  and_gate and_gate_h_u_cla32_and3269_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3269_y0);
  and_gate and_gate_h_u_cla32_and3270_y0(h_u_cla32_and3269_y0, h_u_cla32_and3268_y0, h_u_cla32_and3270_y0);
  and_gate and_gate_h_u_cla32_and3271_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3271_y0);
  and_gate and_gate_h_u_cla32_and3272_y0(h_u_cla32_and3271_y0, h_u_cla32_and3270_y0, h_u_cla32_and3272_y0);
  and_gate and_gate_h_u_cla32_and3273_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3273_y0);
  and_gate and_gate_h_u_cla32_and3274_y0(h_u_cla32_and3273_y0, h_u_cla32_and3272_y0, h_u_cla32_and3274_y0);
  and_gate and_gate_h_u_cla32_and3275_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3275_y0);
  and_gate and_gate_h_u_cla32_and3276_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3276_y0);
  and_gate and_gate_h_u_cla32_and3277_y0(h_u_cla32_and3276_y0, h_u_cla32_and3275_y0, h_u_cla32_and3277_y0);
  and_gate and_gate_h_u_cla32_and3278_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3278_y0);
  and_gate and_gate_h_u_cla32_and3279_y0(h_u_cla32_and3278_y0, h_u_cla32_and3277_y0, h_u_cla32_and3279_y0);
  and_gate and_gate_h_u_cla32_and3280_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3280_y0);
  and_gate and_gate_h_u_cla32_and3281_y0(h_u_cla32_and3280_y0, h_u_cla32_and3279_y0, h_u_cla32_and3281_y0);
  and_gate and_gate_h_u_cla32_and3282_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3282_y0);
  and_gate and_gate_h_u_cla32_and3283_y0(h_u_cla32_and3282_y0, h_u_cla32_and3281_y0, h_u_cla32_and3283_y0);
  and_gate and_gate_h_u_cla32_and3284_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3284_y0);
  and_gate and_gate_h_u_cla32_and3285_y0(h_u_cla32_and3284_y0, h_u_cla32_and3283_y0, h_u_cla32_and3285_y0);
  and_gate and_gate_h_u_cla32_and3286_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3286_y0);
  and_gate and_gate_h_u_cla32_and3287_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3287_y0);
  and_gate and_gate_h_u_cla32_and3288_y0(h_u_cla32_and3287_y0, h_u_cla32_and3286_y0, h_u_cla32_and3288_y0);
  and_gate and_gate_h_u_cla32_and3289_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3289_y0);
  and_gate and_gate_h_u_cla32_and3290_y0(h_u_cla32_and3289_y0, h_u_cla32_and3288_y0, h_u_cla32_and3290_y0);
  and_gate and_gate_h_u_cla32_and3291_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3291_y0);
  and_gate and_gate_h_u_cla32_and3292_y0(h_u_cla32_and3291_y0, h_u_cla32_and3290_y0, h_u_cla32_and3292_y0);
  and_gate and_gate_h_u_cla32_and3293_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3293_y0);
  and_gate and_gate_h_u_cla32_and3294_y0(h_u_cla32_and3293_y0, h_u_cla32_and3292_y0, h_u_cla32_and3294_y0);
  and_gate and_gate_h_u_cla32_and3295_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3295_y0);
  and_gate and_gate_h_u_cla32_and3296_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3296_y0);
  and_gate and_gate_h_u_cla32_and3297_y0(h_u_cla32_and3296_y0, h_u_cla32_and3295_y0, h_u_cla32_and3297_y0);
  and_gate and_gate_h_u_cla32_and3298_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3298_y0);
  and_gate and_gate_h_u_cla32_and3299_y0(h_u_cla32_and3298_y0, h_u_cla32_and3297_y0, h_u_cla32_and3299_y0);
  and_gate and_gate_h_u_cla32_and3300_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3300_y0);
  and_gate and_gate_h_u_cla32_and3301_y0(h_u_cla32_and3300_y0, h_u_cla32_and3299_y0, h_u_cla32_and3301_y0);
  and_gate and_gate_h_u_cla32_and3302_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3302_y0);
  and_gate and_gate_h_u_cla32_and3303_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3303_y0);
  and_gate and_gate_h_u_cla32_and3304_y0(h_u_cla32_and3303_y0, h_u_cla32_and3302_y0, h_u_cla32_and3304_y0);
  and_gate and_gate_h_u_cla32_and3305_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3305_y0);
  and_gate and_gate_h_u_cla32_and3306_y0(h_u_cla32_and3305_y0, h_u_cla32_and3304_y0, h_u_cla32_and3306_y0);
  and_gate and_gate_h_u_cla32_and3307_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and3307_y0);
  and_gate and_gate_h_u_cla32_and3308_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and3308_y0);
  and_gate and_gate_h_u_cla32_and3309_y0(h_u_cla32_and3308_y0, h_u_cla32_and3307_y0, h_u_cla32_and3309_y0);
  and_gate and_gate_h_u_cla32_and3310_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and3310_y0);
  or_gate or_gate_h_u_cla32_or210_y0(h_u_cla32_and3310_y0, h_u_cla32_and2910_y0, h_u_cla32_or210_y0);
  or_gate or_gate_h_u_cla32_or211_y0(h_u_cla32_or210_y0, h_u_cla32_and2949_y0, h_u_cla32_or211_y0);
  or_gate or_gate_h_u_cla32_or212_y0(h_u_cla32_or211_y0, h_u_cla32_and2986_y0, h_u_cla32_or212_y0);
  or_gate or_gate_h_u_cla32_or213_y0(h_u_cla32_or212_y0, h_u_cla32_and3021_y0, h_u_cla32_or213_y0);
  or_gate or_gate_h_u_cla32_or214_y0(h_u_cla32_or213_y0, h_u_cla32_and3054_y0, h_u_cla32_or214_y0);
  or_gate or_gate_h_u_cla32_or215_y0(h_u_cla32_or214_y0, h_u_cla32_and3085_y0, h_u_cla32_or215_y0);
  or_gate or_gate_h_u_cla32_or216_y0(h_u_cla32_or215_y0, h_u_cla32_and3114_y0, h_u_cla32_or216_y0);
  or_gate or_gate_h_u_cla32_or217_y0(h_u_cla32_or216_y0, h_u_cla32_and3141_y0, h_u_cla32_or217_y0);
  or_gate or_gate_h_u_cla32_or218_y0(h_u_cla32_or217_y0, h_u_cla32_and3166_y0, h_u_cla32_or218_y0);
  or_gate or_gate_h_u_cla32_or219_y0(h_u_cla32_or218_y0, h_u_cla32_and3189_y0, h_u_cla32_or219_y0);
  or_gate or_gate_h_u_cla32_or220_y0(h_u_cla32_or219_y0, h_u_cla32_and3210_y0, h_u_cla32_or220_y0);
  or_gate or_gate_h_u_cla32_or221_y0(h_u_cla32_or220_y0, h_u_cla32_and3229_y0, h_u_cla32_or221_y0);
  or_gate or_gate_h_u_cla32_or222_y0(h_u_cla32_or221_y0, h_u_cla32_and3246_y0, h_u_cla32_or222_y0);
  or_gate or_gate_h_u_cla32_or223_y0(h_u_cla32_or222_y0, h_u_cla32_and3261_y0, h_u_cla32_or223_y0);
  or_gate or_gate_h_u_cla32_or224_y0(h_u_cla32_or223_y0, h_u_cla32_and3274_y0, h_u_cla32_or224_y0);
  or_gate or_gate_h_u_cla32_or225_y0(h_u_cla32_or224_y0, h_u_cla32_and3285_y0, h_u_cla32_or225_y0);
  or_gate or_gate_h_u_cla32_or226_y0(h_u_cla32_or225_y0, h_u_cla32_and3294_y0, h_u_cla32_or226_y0);
  or_gate or_gate_h_u_cla32_or227_y0(h_u_cla32_or226_y0, h_u_cla32_and3301_y0, h_u_cla32_or227_y0);
  or_gate or_gate_h_u_cla32_or228_y0(h_u_cla32_or227_y0, h_u_cla32_and3306_y0, h_u_cla32_or228_y0);
  or_gate or_gate_h_u_cla32_or229_y0(h_u_cla32_or228_y0, h_u_cla32_and3309_y0, h_u_cla32_or229_y0);
  or_gate or_gate_h_u_cla32_or230_y0(h_u_cla32_pg_logic20_y1, h_u_cla32_or229_y0, h_u_cla32_or230_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic21_y0(a_21, b_21, h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_pg_logic21_y2);
  xor_gate xor_gate_h_u_cla32_xor21_y0(h_u_cla32_pg_logic21_y2, h_u_cla32_or230_y0, h_u_cla32_xor21_y0);
  and_gate and_gate_h_u_cla32_and3311_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and3311_y0);
  and_gate and_gate_h_u_cla32_and3312_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and3312_y0);
  and_gate and_gate_h_u_cla32_and3313_y0(h_u_cla32_and3312_y0, h_u_cla32_and3311_y0, h_u_cla32_and3313_y0);
  and_gate and_gate_h_u_cla32_and3314_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and3314_y0);
  and_gate and_gate_h_u_cla32_and3315_y0(h_u_cla32_and3314_y0, h_u_cla32_and3313_y0, h_u_cla32_and3315_y0);
  and_gate and_gate_h_u_cla32_and3316_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and3316_y0);
  and_gate and_gate_h_u_cla32_and3317_y0(h_u_cla32_and3316_y0, h_u_cla32_and3315_y0, h_u_cla32_and3317_y0);
  and_gate and_gate_h_u_cla32_and3318_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and3318_y0);
  and_gate and_gate_h_u_cla32_and3319_y0(h_u_cla32_and3318_y0, h_u_cla32_and3317_y0, h_u_cla32_and3319_y0);
  and_gate and_gate_h_u_cla32_and3320_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and3320_y0);
  and_gate and_gate_h_u_cla32_and3321_y0(h_u_cla32_and3320_y0, h_u_cla32_and3319_y0, h_u_cla32_and3321_y0);
  and_gate and_gate_h_u_cla32_and3322_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and3322_y0);
  and_gate and_gate_h_u_cla32_and3323_y0(h_u_cla32_and3322_y0, h_u_cla32_and3321_y0, h_u_cla32_and3323_y0);
  and_gate and_gate_h_u_cla32_and3324_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and3324_y0);
  and_gate and_gate_h_u_cla32_and3325_y0(h_u_cla32_and3324_y0, h_u_cla32_and3323_y0, h_u_cla32_and3325_y0);
  and_gate and_gate_h_u_cla32_and3326_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and3326_y0);
  and_gate and_gate_h_u_cla32_and3327_y0(h_u_cla32_and3326_y0, h_u_cla32_and3325_y0, h_u_cla32_and3327_y0);
  and_gate and_gate_h_u_cla32_and3328_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and3328_y0);
  and_gate and_gate_h_u_cla32_and3329_y0(h_u_cla32_and3328_y0, h_u_cla32_and3327_y0, h_u_cla32_and3329_y0);
  and_gate and_gate_h_u_cla32_and3330_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and3330_y0);
  and_gate and_gate_h_u_cla32_and3331_y0(h_u_cla32_and3330_y0, h_u_cla32_and3329_y0, h_u_cla32_and3331_y0);
  and_gate and_gate_h_u_cla32_and3332_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and3332_y0);
  and_gate and_gate_h_u_cla32_and3333_y0(h_u_cla32_and3332_y0, h_u_cla32_and3331_y0, h_u_cla32_and3333_y0);
  and_gate and_gate_h_u_cla32_and3334_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and3334_y0);
  and_gate and_gate_h_u_cla32_and3335_y0(h_u_cla32_and3334_y0, h_u_cla32_and3333_y0, h_u_cla32_and3335_y0);
  and_gate and_gate_h_u_cla32_and3336_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and3336_y0);
  and_gate and_gate_h_u_cla32_and3337_y0(h_u_cla32_and3336_y0, h_u_cla32_and3335_y0, h_u_cla32_and3337_y0);
  and_gate and_gate_h_u_cla32_and3338_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and3338_y0);
  and_gate and_gate_h_u_cla32_and3339_y0(h_u_cla32_and3338_y0, h_u_cla32_and3337_y0, h_u_cla32_and3339_y0);
  and_gate and_gate_h_u_cla32_and3340_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and3340_y0);
  and_gate and_gate_h_u_cla32_and3341_y0(h_u_cla32_and3340_y0, h_u_cla32_and3339_y0, h_u_cla32_and3341_y0);
  and_gate and_gate_h_u_cla32_and3342_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and3342_y0);
  and_gate and_gate_h_u_cla32_and3343_y0(h_u_cla32_and3342_y0, h_u_cla32_and3341_y0, h_u_cla32_and3343_y0);
  and_gate and_gate_h_u_cla32_and3344_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and3344_y0);
  and_gate and_gate_h_u_cla32_and3345_y0(h_u_cla32_and3344_y0, h_u_cla32_and3343_y0, h_u_cla32_and3345_y0);
  and_gate and_gate_h_u_cla32_and3346_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and3346_y0);
  and_gate and_gate_h_u_cla32_and3347_y0(h_u_cla32_and3346_y0, h_u_cla32_and3345_y0, h_u_cla32_and3347_y0);
  and_gate and_gate_h_u_cla32_and3348_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and3348_y0);
  and_gate and_gate_h_u_cla32_and3349_y0(h_u_cla32_and3348_y0, h_u_cla32_and3347_y0, h_u_cla32_and3349_y0);
  and_gate and_gate_h_u_cla32_and3350_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and3350_y0);
  and_gate and_gate_h_u_cla32_and3351_y0(h_u_cla32_and3350_y0, h_u_cla32_and3349_y0, h_u_cla32_and3351_y0);
  and_gate and_gate_h_u_cla32_and3352_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and3352_y0);
  and_gate and_gate_h_u_cla32_and3353_y0(h_u_cla32_and3352_y0, h_u_cla32_and3351_y0, h_u_cla32_and3353_y0);
  and_gate and_gate_h_u_cla32_and3354_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3354_y0);
  and_gate and_gate_h_u_cla32_and3355_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3355_y0);
  and_gate and_gate_h_u_cla32_and3356_y0(h_u_cla32_and3355_y0, h_u_cla32_and3354_y0, h_u_cla32_and3356_y0);
  and_gate and_gate_h_u_cla32_and3357_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3357_y0);
  and_gate and_gate_h_u_cla32_and3358_y0(h_u_cla32_and3357_y0, h_u_cla32_and3356_y0, h_u_cla32_and3358_y0);
  and_gate and_gate_h_u_cla32_and3359_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3359_y0);
  and_gate and_gate_h_u_cla32_and3360_y0(h_u_cla32_and3359_y0, h_u_cla32_and3358_y0, h_u_cla32_and3360_y0);
  and_gate and_gate_h_u_cla32_and3361_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3361_y0);
  and_gate and_gate_h_u_cla32_and3362_y0(h_u_cla32_and3361_y0, h_u_cla32_and3360_y0, h_u_cla32_and3362_y0);
  and_gate and_gate_h_u_cla32_and3363_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3363_y0);
  and_gate and_gate_h_u_cla32_and3364_y0(h_u_cla32_and3363_y0, h_u_cla32_and3362_y0, h_u_cla32_and3364_y0);
  and_gate and_gate_h_u_cla32_and3365_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3365_y0);
  and_gate and_gate_h_u_cla32_and3366_y0(h_u_cla32_and3365_y0, h_u_cla32_and3364_y0, h_u_cla32_and3366_y0);
  and_gate and_gate_h_u_cla32_and3367_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3367_y0);
  and_gate and_gate_h_u_cla32_and3368_y0(h_u_cla32_and3367_y0, h_u_cla32_and3366_y0, h_u_cla32_and3368_y0);
  and_gate and_gate_h_u_cla32_and3369_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3369_y0);
  and_gate and_gate_h_u_cla32_and3370_y0(h_u_cla32_and3369_y0, h_u_cla32_and3368_y0, h_u_cla32_and3370_y0);
  and_gate and_gate_h_u_cla32_and3371_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3371_y0);
  and_gate and_gate_h_u_cla32_and3372_y0(h_u_cla32_and3371_y0, h_u_cla32_and3370_y0, h_u_cla32_and3372_y0);
  and_gate and_gate_h_u_cla32_and3373_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3373_y0);
  and_gate and_gate_h_u_cla32_and3374_y0(h_u_cla32_and3373_y0, h_u_cla32_and3372_y0, h_u_cla32_and3374_y0);
  and_gate and_gate_h_u_cla32_and3375_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3375_y0);
  and_gate and_gate_h_u_cla32_and3376_y0(h_u_cla32_and3375_y0, h_u_cla32_and3374_y0, h_u_cla32_and3376_y0);
  and_gate and_gate_h_u_cla32_and3377_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3377_y0);
  and_gate and_gate_h_u_cla32_and3378_y0(h_u_cla32_and3377_y0, h_u_cla32_and3376_y0, h_u_cla32_and3378_y0);
  and_gate and_gate_h_u_cla32_and3379_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3379_y0);
  and_gate and_gate_h_u_cla32_and3380_y0(h_u_cla32_and3379_y0, h_u_cla32_and3378_y0, h_u_cla32_and3380_y0);
  and_gate and_gate_h_u_cla32_and3381_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3381_y0);
  and_gate and_gate_h_u_cla32_and3382_y0(h_u_cla32_and3381_y0, h_u_cla32_and3380_y0, h_u_cla32_and3382_y0);
  and_gate and_gate_h_u_cla32_and3383_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3383_y0);
  and_gate and_gate_h_u_cla32_and3384_y0(h_u_cla32_and3383_y0, h_u_cla32_and3382_y0, h_u_cla32_and3384_y0);
  and_gate and_gate_h_u_cla32_and3385_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3385_y0);
  and_gate and_gate_h_u_cla32_and3386_y0(h_u_cla32_and3385_y0, h_u_cla32_and3384_y0, h_u_cla32_and3386_y0);
  and_gate and_gate_h_u_cla32_and3387_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3387_y0);
  and_gate and_gate_h_u_cla32_and3388_y0(h_u_cla32_and3387_y0, h_u_cla32_and3386_y0, h_u_cla32_and3388_y0);
  and_gate and_gate_h_u_cla32_and3389_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3389_y0);
  and_gate and_gate_h_u_cla32_and3390_y0(h_u_cla32_and3389_y0, h_u_cla32_and3388_y0, h_u_cla32_and3390_y0);
  and_gate and_gate_h_u_cla32_and3391_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3391_y0);
  and_gate and_gate_h_u_cla32_and3392_y0(h_u_cla32_and3391_y0, h_u_cla32_and3390_y0, h_u_cla32_and3392_y0);
  and_gate and_gate_h_u_cla32_and3393_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3393_y0);
  and_gate and_gate_h_u_cla32_and3394_y0(h_u_cla32_and3393_y0, h_u_cla32_and3392_y0, h_u_cla32_and3394_y0);
  and_gate and_gate_h_u_cla32_and3395_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3395_y0);
  and_gate and_gate_h_u_cla32_and3396_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3396_y0);
  and_gate and_gate_h_u_cla32_and3397_y0(h_u_cla32_and3396_y0, h_u_cla32_and3395_y0, h_u_cla32_and3397_y0);
  and_gate and_gate_h_u_cla32_and3398_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3398_y0);
  and_gate and_gate_h_u_cla32_and3399_y0(h_u_cla32_and3398_y0, h_u_cla32_and3397_y0, h_u_cla32_and3399_y0);
  and_gate and_gate_h_u_cla32_and3400_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3400_y0);
  and_gate and_gate_h_u_cla32_and3401_y0(h_u_cla32_and3400_y0, h_u_cla32_and3399_y0, h_u_cla32_and3401_y0);
  and_gate and_gate_h_u_cla32_and3402_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3402_y0);
  and_gate and_gate_h_u_cla32_and3403_y0(h_u_cla32_and3402_y0, h_u_cla32_and3401_y0, h_u_cla32_and3403_y0);
  and_gate and_gate_h_u_cla32_and3404_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3404_y0);
  and_gate and_gate_h_u_cla32_and3405_y0(h_u_cla32_and3404_y0, h_u_cla32_and3403_y0, h_u_cla32_and3405_y0);
  and_gate and_gate_h_u_cla32_and3406_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3406_y0);
  and_gate and_gate_h_u_cla32_and3407_y0(h_u_cla32_and3406_y0, h_u_cla32_and3405_y0, h_u_cla32_and3407_y0);
  and_gate and_gate_h_u_cla32_and3408_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3408_y0);
  and_gate and_gate_h_u_cla32_and3409_y0(h_u_cla32_and3408_y0, h_u_cla32_and3407_y0, h_u_cla32_and3409_y0);
  and_gate and_gate_h_u_cla32_and3410_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3410_y0);
  and_gate and_gate_h_u_cla32_and3411_y0(h_u_cla32_and3410_y0, h_u_cla32_and3409_y0, h_u_cla32_and3411_y0);
  and_gate and_gate_h_u_cla32_and3412_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3412_y0);
  and_gate and_gate_h_u_cla32_and3413_y0(h_u_cla32_and3412_y0, h_u_cla32_and3411_y0, h_u_cla32_and3413_y0);
  and_gate and_gate_h_u_cla32_and3414_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3414_y0);
  and_gate and_gate_h_u_cla32_and3415_y0(h_u_cla32_and3414_y0, h_u_cla32_and3413_y0, h_u_cla32_and3415_y0);
  and_gate and_gate_h_u_cla32_and3416_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3416_y0);
  and_gate and_gate_h_u_cla32_and3417_y0(h_u_cla32_and3416_y0, h_u_cla32_and3415_y0, h_u_cla32_and3417_y0);
  and_gate and_gate_h_u_cla32_and3418_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3418_y0);
  and_gate and_gate_h_u_cla32_and3419_y0(h_u_cla32_and3418_y0, h_u_cla32_and3417_y0, h_u_cla32_and3419_y0);
  and_gate and_gate_h_u_cla32_and3420_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3420_y0);
  and_gate and_gate_h_u_cla32_and3421_y0(h_u_cla32_and3420_y0, h_u_cla32_and3419_y0, h_u_cla32_and3421_y0);
  and_gate and_gate_h_u_cla32_and3422_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3422_y0);
  and_gate and_gate_h_u_cla32_and3423_y0(h_u_cla32_and3422_y0, h_u_cla32_and3421_y0, h_u_cla32_and3423_y0);
  and_gate and_gate_h_u_cla32_and3424_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3424_y0);
  and_gate and_gate_h_u_cla32_and3425_y0(h_u_cla32_and3424_y0, h_u_cla32_and3423_y0, h_u_cla32_and3425_y0);
  and_gate and_gate_h_u_cla32_and3426_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3426_y0);
  and_gate and_gate_h_u_cla32_and3427_y0(h_u_cla32_and3426_y0, h_u_cla32_and3425_y0, h_u_cla32_and3427_y0);
  and_gate and_gate_h_u_cla32_and3428_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3428_y0);
  and_gate and_gate_h_u_cla32_and3429_y0(h_u_cla32_and3428_y0, h_u_cla32_and3427_y0, h_u_cla32_and3429_y0);
  and_gate and_gate_h_u_cla32_and3430_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3430_y0);
  and_gate and_gate_h_u_cla32_and3431_y0(h_u_cla32_and3430_y0, h_u_cla32_and3429_y0, h_u_cla32_and3431_y0);
  and_gate and_gate_h_u_cla32_and3432_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3432_y0);
  and_gate and_gate_h_u_cla32_and3433_y0(h_u_cla32_and3432_y0, h_u_cla32_and3431_y0, h_u_cla32_and3433_y0);
  and_gate and_gate_h_u_cla32_and3434_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3434_y0);
  and_gate and_gate_h_u_cla32_and3435_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3435_y0);
  and_gate and_gate_h_u_cla32_and3436_y0(h_u_cla32_and3435_y0, h_u_cla32_and3434_y0, h_u_cla32_and3436_y0);
  and_gate and_gate_h_u_cla32_and3437_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3437_y0);
  and_gate and_gate_h_u_cla32_and3438_y0(h_u_cla32_and3437_y0, h_u_cla32_and3436_y0, h_u_cla32_and3438_y0);
  and_gate and_gate_h_u_cla32_and3439_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3439_y0);
  and_gate and_gate_h_u_cla32_and3440_y0(h_u_cla32_and3439_y0, h_u_cla32_and3438_y0, h_u_cla32_and3440_y0);
  and_gate and_gate_h_u_cla32_and3441_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3441_y0);
  and_gate and_gate_h_u_cla32_and3442_y0(h_u_cla32_and3441_y0, h_u_cla32_and3440_y0, h_u_cla32_and3442_y0);
  and_gate and_gate_h_u_cla32_and3443_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3443_y0);
  and_gate and_gate_h_u_cla32_and3444_y0(h_u_cla32_and3443_y0, h_u_cla32_and3442_y0, h_u_cla32_and3444_y0);
  and_gate and_gate_h_u_cla32_and3445_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3445_y0);
  and_gate and_gate_h_u_cla32_and3446_y0(h_u_cla32_and3445_y0, h_u_cla32_and3444_y0, h_u_cla32_and3446_y0);
  and_gate and_gate_h_u_cla32_and3447_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3447_y0);
  and_gate and_gate_h_u_cla32_and3448_y0(h_u_cla32_and3447_y0, h_u_cla32_and3446_y0, h_u_cla32_and3448_y0);
  and_gate and_gate_h_u_cla32_and3449_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3449_y0);
  and_gate and_gate_h_u_cla32_and3450_y0(h_u_cla32_and3449_y0, h_u_cla32_and3448_y0, h_u_cla32_and3450_y0);
  and_gate and_gate_h_u_cla32_and3451_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3451_y0);
  and_gate and_gate_h_u_cla32_and3452_y0(h_u_cla32_and3451_y0, h_u_cla32_and3450_y0, h_u_cla32_and3452_y0);
  and_gate and_gate_h_u_cla32_and3453_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3453_y0);
  and_gate and_gate_h_u_cla32_and3454_y0(h_u_cla32_and3453_y0, h_u_cla32_and3452_y0, h_u_cla32_and3454_y0);
  and_gate and_gate_h_u_cla32_and3455_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3455_y0);
  and_gate and_gate_h_u_cla32_and3456_y0(h_u_cla32_and3455_y0, h_u_cla32_and3454_y0, h_u_cla32_and3456_y0);
  and_gate and_gate_h_u_cla32_and3457_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3457_y0);
  and_gate and_gate_h_u_cla32_and3458_y0(h_u_cla32_and3457_y0, h_u_cla32_and3456_y0, h_u_cla32_and3458_y0);
  and_gate and_gate_h_u_cla32_and3459_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3459_y0);
  and_gate and_gate_h_u_cla32_and3460_y0(h_u_cla32_and3459_y0, h_u_cla32_and3458_y0, h_u_cla32_and3460_y0);
  and_gate and_gate_h_u_cla32_and3461_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3461_y0);
  and_gate and_gate_h_u_cla32_and3462_y0(h_u_cla32_and3461_y0, h_u_cla32_and3460_y0, h_u_cla32_and3462_y0);
  and_gate and_gate_h_u_cla32_and3463_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3463_y0);
  and_gate and_gate_h_u_cla32_and3464_y0(h_u_cla32_and3463_y0, h_u_cla32_and3462_y0, h_u_cla32_and3464_y0);
  and_gate and_gate_h_u_cla32_and3465_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3465_y0);
  and_gate and_gate_h_u_cla32_and3466_y0(h_u_cla32_and3465_y0, h_u_cla32_and3464_y0, h_u_cla32_and3466_y0);
  and_gate and_gate_h_u_cla32_and3467_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3467_y0);
  and_gate and_gate_h_u_cla32_and3468_y0(h_u_cla32_and3467_y0, h_u_cla32_and3466_y0, h_u_cla32_and3468_y0);
  and_gate and_gate_h_u_cla32_and3469_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3469_y0);
  and_gate and_gate_h_u_cla32_and3470_y0(h_u_cla32_and3469_y0, h_u_cla32_and3468_y0, h_u_cla32_and3470_y0);
  and_gate and_gate_h_u_cla32_and3471_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3471_y0);
  and_gate and_gate_h_u_cla32_and3472_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3472_y0);
  and_gate and_gate_h_u_cla32_and3473_y0(h_u_cla32_and3472_y0, h_u_cla32_and3471_y0, h_u_cla32_and3473_y0);
  and_gate and_gate_h_u_cla32_and3474_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3474_y0);
  and_gate and_gate_h_u_cla32_and3475_y0(h_u_cla32_and3474_y0, h_u_cla32_and3473_y0, h_u_cla32_and3475_y0);
  and_gate and_gate_h_u_cla32_and3476_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3476_y0);
  and_gate and_gate_h_u_cla32_and3477_y0(h_u_cla32_and3476_y0, h_u_cla32_and3475_y0, h_u_cla32_and3477_y0);
  and_gate and_gate_h_u_cla32_and3478_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3478_y0);
  and_gate and_gate_h_u_cla32_and3479_y0(h_u_cla32_and3478_y0, h_u_cla32_and3477_y0, h_u_cla32_and3479_y0);
  and_gate and_gate_h_u_cla32_and3480_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3480_y0);
  and_gate and_gate_h_u_cla32_and3481_y0(h_u_cla32_and3480_y0, h_u_cla32_and3479_y0, h_u_cla32_and3481_y0);
  and_gate and_gate_h_u_cla32_and3482_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3482_y0);
  and_gate and_gate_h_u_cla32_and3483_y0(h_u_cla32_and3482_y0, h_u_cla32_and3481_y0, h_u_cla32_and3483_y0);
  and_gate and_gate_h_u_cla32_and3484_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3484_y0);
  and_gate and_gate_h_u_cla32_and3485_y0(h_u_cla32_and3484_y0, h_u_cla32_and3483_y0, h_u_cla32_and3485_y0);
  and_gate and_gate_h_u_cla32_and3486_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3486_y0);
  and_gate and_gate_h_u_cla32_and3487_y0(h_u_cla32_and3486_y0, h_u_cla32_and3485_y0, h_u_cla32_and3487_y0);
  and_gate and_gate_h_u_cla32_and3488_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3488_y0);
  and_gate and_gate_h_u_cla32_and3489_y0(h_u_cla32_and3488_y0, h_u_cla32_and3487_y0, h_u_cla32_and3489_y0);
  and_gate and_gate_h_u_cla32_and3490_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3490_y0);
  and_gate and_gate_h_u_cla32_and3491_y0(h_u_cla32_and3490_y0, h_u_cla32_and3489_y0, h_u_cla32_and3491_y0);
  and_gate and_gate_h_u_cla32_and3492_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3492_y0);
  and_gate and_gate_h_u_cla32_and3493_y0(h_u_cla32_and3492_y0, h_u_cla32_and3491_y0, h_u_cla32_and3493_y0);
  and_gate and_gate_h_u_cla32_and3494_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3494_y0);
  and_gate and_gate_h_u_cla32_and3495_y0(h_u_cla32_and3494_y0, h_u_cla32_and3493_y0, h_u_cla32_and3495_y0);
  and_gate and_gate_h_u_cla32_and3496_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3496_y0);
  and_gate and_gate_h_u_cla32_and3497_y0(h_u_cla32_and3496_y0, h_u_cla32_and3495_y0, h_u_cla32_and3497_y0);
  and_gate and_gate_h_u_cla32_and3498_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3498_y0);
  and_gate and_gate_h_u_cla32_and3499_y0(h_u_cla32_and3498_y0, h_u_cla32_and3497_y0, h_u_cla32_and3499_y0);
  and_gate and_gate_h_u_cla32_and3500_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3500_y0);
  and_gate and_gate_h_u_cla32_and3501_y0(h_u_cla32_and3500_y0, h_u_cla32_and3499_y0, h_u_cla32_and3501_y0);
  and_gate and_gate_h_u_cla32_and3502_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3502_y0);
  and_gate and_gate_h_u_cla32_and3503_y0(h_u_cla32_and3502_y0, h_u_cla32_and3501_y0, h_u_cla32_and3503_y0);
  and_gate and_gate_h_u_cla32_and3504_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3504_y0);
  and_gate and_gate_h_u_cla32_and3505_y0(h_u_cla32_and3504_y0, h_u_cla32_and3503_y0, h_u_cla32_and3505_y0);
  and_gate and_gate_h_u_cla32_and3506_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3506_y0);
  and_gate and_gate_h_u_cla32_and3507_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3507_y0);
  and_gate and_gate_h_u_cla32_and3508_y0(h_u_cla32_and3507_y0, h_u_cla32_and3506_y0, h_u_cla32_and3508_y0);
  and_gate and_gate_h_u_cla32_and3509_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3509_y0);
  and_gate and_gate_h_u_cla32_and3510_y0(h_u_cla32_and3509_y0, h_u_cla32_and3508_y0, h_u_cla32_and3510_y0);
  and_gate and_gate_h_u_cla32_and3511_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3511_y0);
  and_gate and_gate_h_u_cla32_and3512_y0(h_u_cla32_and3511_y0, h_u_cla32_and3510_y0, h_u_cla32_and3512_y0);
  and_gate and_gate_h_u_cla32_and3513_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3513_y0);
  and_gate and_gate_h_u_cla32_and3514_y0(h_u_cla32_and3513_y0, h_u_cla32_and3512_y0, h_u_cla32_and3514_y0);
  and_gate and_gate_h_u_cla32_and3515_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3515_y0);
  and_gate and_gate_h_u_cla32_and3516_y0(h_u_cla32_and3515_y0, h_u_cla32_and3514_y0, h_u_cla32_and3516_y0);
  and_gate and_gate_h_u_cla32_and3517_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3517_y0);
  and_gate and_gate_h_u_cla32_and3518_y0(h_u_cla32_and3517_y0, h_u_cla32_and3516_y0, h_u_cla32_and3518_y0);
  and_gate and_gate_h_u_cla32_and3519_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3519_y0);
  and_gate and_gate_h_u_cla32_and3520_y0(h_u_cla32_and3519_y0, h_u_cla32_and3518_y0, h_u_cla32_and3520_y0);
  and_gate and_gate_h_u_cla32_and3521_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3521_y0);
  and_gate and_gate_h_u_cla32_and3522_y0(h_u_cla32_and3521_y0, h_u_cla32_and3520_y0, h_u_cla32_and3522_y0);
  and_gate and_gate_h_u_cla32_and3523_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3523_y0);
  and_gate and_gate_h_u_cla32_and3524_y0(h_u_cla32_and3523_y0, h_u_cla32_and3522_y0, h_u_cla32_and3524_y0);
  and_gate and_gate_h_u_cla32_and3525_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3525_y0);
  and_gate and_gate_h_u_cla32_and3526_y0(h_u_cla32_and3525_y0, h_u_cla32_and3524_y0, h_u_cla32_and3526_y0);
  and_gate and_gate_h_u_cla32_and3527_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3527_y0);
  and_gate and_gate_h_u_cla32_and3528_y0(h_u_cla32_and3527_y0, h_u_cla32_and3526_y0, h_u_cla32_and3528_y0);
  and_gate and_gate_h_u_cla32_and3529_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3529_y0);
  and_gate and_gate_h_u_cla32_and3530_y0(h_u_cla32_and3529_y0, h_u_cla32_and3528_y0, h_u_cla32_and3530_y0);
  and_gate and_gate_h_u_cla32_and3531_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3531_y0);
  and_gate and_gate_h_u_cla32_and3532_y0(h_u_cla32_and3531_y0, h_u_cla32_and3530_y0, h_u_cla32_and3532_y0);
  and_gate and_gate_h_u_cla32_and3533_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3533_y0);
  and_gate and_gate_h_u_cla32_and3534_y0(h_u_cla32_and3533_y0, h_u_cla32_and3532_y0, h_u_cla32_and3534_y0);
  and_gate and_gate_h_u_cla32_and3535_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3535_y0);
  and_gate and_gate_h_u_cla32_and3536_y0(h_u_cla32_and3535_y0, h_u_cla32_and3534_y0, h_u_cla32_and3536_y0);
  and_gate and_gate_h_u_cla32_and3537_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and3537_y0);
  and_gate and_gate_h_u_cla32_and3538_y0(h_u_cla32_and3537_y0, h_u_cla32_and3536_y0, h_u_cla32_and3538_y0);
  and_gate and_gate_h_u_cla32_and3539_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3539_y0);
  and_gate and_gate_h_u_cla32_and3540_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3540_y0);
  and_gate and_gate_h_u_cla32_and3541_y0(h_u_cla32_and3540_y0, h_u_cla32_and3539_y0, h_u_cla32_and3541_y0);
  and_gate and_gate_h_u_cla32_and3542_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3542_y0);
  and_gate and_gate_h_u_cla32_and3543_y0(h_u_cla32_and3542_y0, h_u_cla32_and3541_y0, h_u_cla32_and3543_y0);
  and_gate and_gate_h_u_cla32_and3544_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3544_y0);
  and_gate and_gate_h_u_cla32_and3545_y0(h_u_cla32_and3544_y0, h_u_cla32_and3543_y0, h_u_cla32_and3545_y0);
  and_gate and_gate_h_u_cla32_and3546_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3546_y0);
  and_gate and_gate_h_u_cla32_and3547_y0(h_u_cla32_and3546_y0, h_u_cla32_and3545_y0, h_u_cla32_and3547_y0);
  and_gate and_gate_h_u_cla32_and3548_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3548_y0);
  and_gate and_gate_h_u_cla32_and3549_y0(h_u_cla32_and3548_y0, h_u_cla32_and3547_y0, h_u_cla32_and3549_y0);
  and_gate and_gate_h_u_cla32_and3550_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3550_y0);
  and_gate and_gate_h_u_cla32_and3551_y0(h_u_cla32_and3550_y0, h_u_cla32_and3549_y0, h_u_cla32_and3551_y0);
  and_gate and_gate_h_u_cla32_and3552_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3552_y0);
  and_gate and_gate_h_u_cla32_and3553_y0(h_u_cla32_and3552_y0, h_u_cla32_and3551_y0, h_u_cla32_and3553_y0);
  and_gate and_gate_h_u_cla32_and3554_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3554_y0);
  and_gate and_gate_h_u_cla32_and3555_y0(h_u_cla32_and3554_y0, h_u_cla32_and3553_y0, h_u_cla32_and3555_y0);
  and_gate and_gate_h_u_cla32_and3556_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3556_y0);
  and_gate and_gate_h_u_cla32_and3557_y0(h_u_cla32_and3556_y0, h_u_cla32_and3555_y0, h_u_cla32_and3557_y0);
  and_gate and_gate_h_u_cla32_and3558_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3558_y0);
  and_gate and_gate_h_u_cla32_and3559_y0(h_u_cla32_and3558_y0, h_u_cla32_and3557_y0, h_u_cla32_and3559_y0);
  and_gate and_gate_h_u_cla32_and3560_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3560_y0);
  and_gate and_gate_h_u_cla32_and3561_y0(h_u_cla32_and3560_y0, h_u_cla32_and3559_y0, h_u_cla32_and3561_y0);
  and_gate and_gate_h_u_cla32_and3562_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3562_y0);
  and_gate and_gate_h_u_cla32_and3563_y0(h_u_cla32_and3562_y0, h_u_cla32_and3561_y0, h_u_cla32_and3563_y0);
  and_gate and_gate_h_u_cla32_and3564_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3564_y0);
  and_gate and_gate_h_u_cla32_and3565_y0(h_u_cla32_and3564_y0, h_u_cla32_and3563_y0, h_u_cla32_and3565_y0);
  and_gate and_gate_h_u_cla32_and3566_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3566_y0);
  and_gate and_gate_h_u_cla32_and3567_y0(h_u_cla32_and3566_y0, h_u_cla32_and3565_y0, h_u_cla32_and3567_y0);
  and_gate and_gate_h_u_cla32_and3568_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and3568_y0);
  and_gate and_gate_h_u_cla32_and3569_y0(h_u_cla32_and3568_y0, h_u_cla32_and3567_y0, h_u_cla32_and3569_y0);
  and_gate and_gate_h_u_cla32_and3570_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3570_y0);
  and_gate and_gate_h_u_cla32_and3571_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3571_y0);
  and_gate and_gate_h_u_cla32_and3572_y0(h_u_cla32_and3571_y0, h_u_cla32_and3570_y0, h_u_cla32_and3572_y0);
  and_gate and_gate_h_u_cla32_and3573_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3573_y0);
  and_gate and_gate_h_u_cla32_and3574_y0(h_u_cla32_and3573_y0, h_u_cla32_and3572_y0, h_u_cla32_and3574_y0);
  and_gate and_gate_h_u_cla32_and3575_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3575_y0);
  and_gate and_gate_h_u_cla32_and3576_y0(h_u_cla32_and3575_y0, h_u_cla32_and3574_y0, h_u_cla32_and3576_y0);
  and_gate and_gate_h_u_cla32_and3577_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3577_y0);
  and_gate and_gate_h_u_cla32_and3578_y0(h_u_cla32_and3577_y0, h_u_cla32_and3576_y0, h_u_cla32_and3578_y0);
  and_gate and_gate_h_u_cla32_and3579_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3579_y0);
  and_gate and_gate_h_u_cla32_and3580_y0(h_u_cla32_and3579_y0, h_u_cla32_and3578_y0, h_u_cla32_and3580_y0);
  and_gate and_gate_h_u_cla32_and3581_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3581_y0);
  and_gate and_gate_h_u_cla32_and3582_y0(h_u_cla32_and3581_y0, h_u_cla32_and3580_y0, h_u_cla32_and3582_y0);
  and_gate and_gate_h_u_cla32_and3583_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3583_y0);
  and_gate and_gate_h_u_cla32_and3584_y0(h_u_cla32_and3583_y0, h_u_cla32_and3582_y0, h_u_cla32_and3584_y0);
  and_gate and_gate_h_u_cla32_and3585_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3585_y0);
  and_gate and_gate_h_u_cla32_and3586_y0(h_u_cla32_and3585_y0, h_u_cla32_and3584_y0, h_u_cla32_and3586_y0);
  and_gate and_gate_h_u_cla32_and3587_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3587_y0);
  and_gate and_gate_h_u_cla32_and3588_y0(h_u_cla32_and3587_y0, h_u_cla32_and3586_y0, h_u_cla32_and3588_y0);
  and_gate and_gate_h_u_cla32_and3589_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3589_y0);
  and_gate and_gate_h_u_cla32_and3590_y0(h_u_cla32_and3589_y0, h_u_cla32_and3588_y0, h_u_cla32_and3590_y0);
  and_gate and_gate_h_u_cla32_and3591_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3591_y0);
  and_gate and_gate_h_u_cla32_and3592_y0(h_u_cla32_and3591_y0, h_u_cla32_and3590_y0, h_u_cla32_and3592_y0);
  and_gate and_gate_h_u_cla32_and3593_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3593_y0);
  and_gate and_gate_h_u_cla32_and3594_y0(h_u_cla32_and3593_y0, h_u_cla32_and3592_y0, h_u_cla32_and3594_y0);
  and_gate and_gate_h_u_cla32_and3595_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3595_y0);
  and_gate and_gate_h_u_cla32_and3596_y0(h_u_cla32_and3595_y0, h_u_cla32_and3594_y0, h_u_cla32_and3596_y0);
  and_gate and_gate_h_u_cla32_and3597_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and3597_y0);
  and_gate and_gate_h_u_cla32_and3598_y0(h_u_cla32_and3597_y0, h_u_cla32_and3596_y0, h_u_cla32_and3598_y0);
  and_gate and_gate_h_u_cla32_and3599_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3599_y0);
  and_gate and_gate_h_u_cla32_and3600_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3600_y0);
  and_gate and_gate_h_u_cla32_and3601_y0(h_u_cla32_and3600_y0, h_u_cla32_and3599_y0, h_u_cla32_and3601_y0);
  and_gate and_gate_h_u_cla32_and3602_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3602_y0);
  and_gate and_gate_h_u_cla32_and3603_y0(h_u_cla32_and3602_y0, h_u_cla32_and3601_y0, h_u_cla32_and3603_y0);
  and_gate and_gate_h_u_cla32_and3604_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3604_y0);
  and_gate and_gate_h_u_cla32_and3605_y0(h_u_cla32_and3604_y0, h_u_cla32_and3603_y0, h_u_cla32_and3605_y0);
  and_gate and_gate_h_u_cla32_and3606_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3606_y0);
  and_gate and_gate_h_u_cla32_and3607_y0(h_u_cla32_and3606_y0, h_u_cla32_and3605_y0, h_u_cla32_and3607_y0);
  and_gate and_gate_h_u_cla32_and3608_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3608_y0);
  and_gate and_gate_h_u_cla32_and3609_y0(h_u_cla32_and3608_y0, h_u_cla32_and3607_y0, h_u_cla32_and3609_y0);
  and_gate and_gate_h_u_cla32_and3610_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3610_y0);
  and_gate and_gate_h_u_cla32_and3611_y0(h_u_cla32_and3610_y0, h_u_cla32_and3609_y0, h_u_cla32_and3611_y0);
  and_gate and_gate_h_u_cla32_and3612_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3612_y0);
  and_gate and_gate_h_u_cla32_and3613_y0(h_u_cla32_and3612_y0, h_u_cla32_and3611_y0, h_u_cla32_and3613_y0);
  and_gate and_gate_h_u_cla32_and3614_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3614_y0);
  and_gate and_gate_h_u_cla32_and3615_y0(h_u_cla32_and3614_y0, h_u_cla32_and3613_y0, h_u_cla32_and3615_y0);
  and_gate and_gate_h_u_cla32_and3616_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3616_y0);
  and_gate and_gate_h_u_cla32_and3617_y0(h_u_cla32_and3616_y0, h_u_cla32_and3615_y0, h_u_cla32_and3617_y0);
  and_gate and_gate_h_u_cla32_and3618_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3618_y0);
  and_gate and_gate_h_u_cla32_and3619_y0(h_u_cla32_and3618_y0, h_u_cla32_and3617_y0, h_u_cla32_and3619_y0);
  and_gate and_gate_h_u_cla32_and3620_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3620_y0);
  and_gate and_gate_h_u_cla32_and3621_y0(h_u_cla32_and3620_y0, h_u_cla32_and3619_y0, h_u_cla32_and3621_y0);
  and_gate and_gate_h_u_cla32_and3622_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3622_y0);
  and_gate and_gate_h_u_cla32_and3623_y0(h_u_cla32_and3622_y0, h_u_cla32_and3621_y0, h_u_cla32_and3623_y0);
  and_gate and_gate_h_u_cla32_and3624_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and3624_y0);
  and_gate and_gate_h_u_cla32_and3625_y0(h_u_cla32_and3624_y0, h_u_cla32_and3623_y0, h_u_cla32_and3625_y0);
  and_gate and_gate_h_u_cla32_and3626_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3626_y0);
  and_gate and_gate_h_u_cla32_and3627_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3627_y0);
  and_gate and_gate_h_u_cla32_and3628_y0(h_u_cla32_and3627_y0, h_u_cla32_and3626_y0, h_u_cla32_and3628_y0);
  and_gate and_gate_h_u_cla32_and3629_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3629_y0);
  and_gate and_gate_h_u_cla32_and3630_y0(h_u_cla32_and3629_y0, h_u_cla32_and3628_y0, h_u_cla32_and3630_y0);
  and_gate and_gate_h_u_cla32_and3631_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3631_y0);
  and_gate and_gate_h_u_cla32_and3632_y0(h_u_cla32_and3631_y0, h_u_cla32_and3630_y0, h_u_cla32_and3632_y0);
  and_gate and_gate_h_u_cla32_and3633_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3633_y0);
  and_gate and_gate_h_u_cla32_and3634_y0(h_u_cla32_and3633_y0, h_u_cla32_and3632_y0, h_u_cla32_and3634_y0);
  and_gate and_gate_h_u_cla32_and3635_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3635_y0);
  and_gate and_gate_h_u_cla32_and3636_y0(h_u_cla32_and3635_y0, h_u_cla32_and3634_y0, h_u_cla32_and3636_y0);
  and_gate and_gate_h_u_cla32_and3637_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3637_y0);
  and_gate and_gate_h_u_cla32_and3638_y0(h_u_cla32_and3637_y0, h_u_cla32_and3636_y0, h_u_cla32_and3638_y0);
  and_gate and_gate_h_u_cla32_and3639_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3639_y0);
  and_gate and_gate_h_u_cla32_and3640_y0(h_u_cla32_and3639_y0, h_u_cla32_and3638_y0, h_u_cla32_and3640_y0);
  and_gate and_gate_h_u_cla32_and3641_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3641_y0);
  and_gate and_gate_h_u_cla32_and3642_y0(h_u_cla32_and3641_y0, h_u_cla32_and3640_y0, h_u_cla32_and3642_y0);
  and_gate and_gate_h_u_cla32_and3643_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3643_y0);
  and_gate and_gate_h_u_cla32_and3644_y0(h_u_cla32_and3643_y0, h_u_cla32_and3642_y0, h_u_cla32_and3644_y0);
  and_gate and_gate_h_u_cla32_and3645_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3645_y0);
  and_gate and_gate_h_u_cla32_and3646_y0(h_u_cla32_and3645_y0, h_u_cla32_and3644_y0, h_u_cla32_and3646_y0);
  and_gate and_gate_h_u_cla32_and3647_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3647_y0);
  and_gate and_gate_h_u_cla32_and3648_y0(h_u_cla32_and3647_y0, h_u_cla32_and3646_y0, h_u_cla32_and3648_y0);
  and_gate and_gate_h_u_cla32_and3649_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and3649_y0);
  and_gate and_gate_h_u_cla32_and3650_y0(h_u_cla32_and3649_y0, h_u_cla32_and3648_y0, h_u_cla32_and3650_y0);
  and_gate and_gate_h_u_cla32_and3651_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3651_y0);
  and_gate and_gate_h_u_cla32_and3652_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3652_y0);
  and_gate and_gate_h_u_cla32_and3653_y0(h_u_cla32_and3652_y0, h_u_cla32_and3651_y0, h_u_cla32_and3653_y0);
  and_gate and_gate_h_u_cla32_and3654_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3654_y0);
  and_gate and_gate_h_u_cla32_and3655_y0(h_u_cla32_and3654_y0, h_u_cla32_and3653_y0, h_u_cla32_and3655_y0);
  and_gate and_gate_h_u_cla32_and3656_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3656_y0);
  and_gate and_gate_h_u_cla32_and3657_y0(h_u_cla32_and3656_y0, h_u_cla32_and3655_y0, h_u_cla32_and3657_y0);
  and_gate and_gate_h_u_cla32_and3658_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3658_y0);
  and_gate and_gate_h_u_cla32_and3659_y0(h_u_cla32_and3658_y0, h_u_cla32_and3657_y0, h_u_cla32_and3659_y0);
  and_gate and_gate_h_u_cla32_and3660_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3660_y0);
  and_gate and_gate_h_u_cla32_and3661_y0(h_u_cla32_and3660_y0, h_u_cla32_and3659_y0, h_u_cla32_and3661_y0);
  and_gate and_gate_h_u_cla32_and3662_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3662_y0);
  and_gate and_gate_h_u_cla32_and3663_y0(h_u_cla32_and3662_y0, h_u_cla32_and3661_y0, h_u_cla32_and3663_y0);
  and_gate and_gate_h_u_cla32_and3664_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3664_y0);
  and_gate and_gate_h_u_cla32_and3665_y0(h_u_cla32_and3664_y0, h_u_cla32_and3663_y0, h_u_cla32_and3665_y0);
  and_gate and_gate_h_u_cla32_and3666_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3666_y0);
  and_gate and_gate_h_u_cla32_and3667_y0(h_u_cla32_and3666_y0, h_u_cla32_and3665_y0, h_u_cla32_and3667_y0);
  and_gate and_gate_h_u_cla32_and3668_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3668_y0);
  and_gate and_gate_h_u_cla32_and3669_y0(h_u_cla32_and3668_y0, h_u_cla32_and3667_y0, h_u_cla32_and3669_y0);
  and_gate and_gate_h_u_cla32_and3670_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3670_y0);
  and_gate and_gate_h_u_cla32_and3671_y0(h_u_cla32_and3670_y0, h_u_cla32_and3669_y0, h_u_cla32_and3671_y0);
  and_gate and_gate_h_u_cla32_and3672_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and3672_y0);
  and_gate and_gate_h_u_cla32_and3673_y0(h_u_cla32_and3672_y0, h_u_cla32_and3671_y0, h_u_cla32_and3673_y0);
  and_gate and_gate_h_u_cla32_and3674_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3674_y0);
  and_gate and_gate_h_u_cla32_and3675_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3675_y0);
  and_gate and_gate_h_u_cla32_and3676_y0(h_u_cla32_and3675_y0, h_u_cla32_and3674_y0, h_u_cla32_and3676_y0);
  and_gate and_gate_h_u_cla32_and3677_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3677_y0);
  and_gate and_gate_h_u_cla32_and3678_y0(h_u_cla32_and3677_y0, h_u_cla32_and3676_y0, h_u_cla32_and3678_y0);
  and_gate and_gate_h_u_cla32_and3679_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3679_y0);
  and_gate and_gate_h_u_cla32_and3680_y0(h_u_cla32_and3679_y0, h_u_cla32_and3678_y0, h_u_cla32_and3680_y0);
  and_gate and_gate_h_u_cla32_and3681_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3681_y0);
  and_gate and_gate_h_u_cla32_and3682_y0(h_u_cla32_and3681_y0, h_u_cla32_and3680_y0, h_u_cla32_and3682_y0);
  and_gate and_gate_h_u_cla32_and3683_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3683_y0);
  and_gate and_gate_h_u_cla32_and3684_y0(h_u_cla32_and3683_y0, h_u_cla32_and3682_y0, h_u_cla32_and3684_y0);
  and_gate and_gate_h_u_cla32_and3685_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3685_y0);
  and_gate and_gate_h_u_cla32_and3686_y0(h_u_cla32_and3685_y0, h_u_cla32_and3684_y0, h_u_cla32_and3686_y0);
  and_gate and_gate_h_u_cla32_and3687_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3687_y0);
  and_gate and_gate_h_u_cla32_and3688_y0(h_u_cla32_and3687_y0, h_u_cla32_and3686_y0, h_u_cla32_and3688_y0);
  and_gate and_gate_h_u_cla32_and3689_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3689_y0);
  and_gate and_gate_h_u_cla32_and3690_y0(h_u_cla32_and3689_y0, h_u_cla32_and3688_y0, h_u_cla32_and3690_y0);
  and_gate and_gate_h_u_cla32_and3691_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3691_y0);
  and_gate and_gate_h_u_cla32_and3692_y0(h_u_cla32_and3691_y0, h_u_cla32_and3690_y0, h_u_cla32_and3692_y0);
  and_gate and_gate_h_u_cla32_and3693_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and3693_y0);
  and_gate and_gate_h_u_cla32_and3694_y0(h_u_cla32_and3693_y0, h_u_cla32_and3692_y0, h_u_cla32_and3694_y0);
  and_gate and_gate_h_u_cla32_and3695_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3695_y0);
  and_gate and_gate_h_u_cla32_and3696_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3696_y0);
  and_gate and_gate_h_u_cla32_and3697_y0(h_u_cla32_and3696_y0, h_u_cla32_and3695_y0, h_u_cla32_and3697_y0);
  and_gate and_gate_h_u_cla32_and3698_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3698_y0);
  and_gate and_gate_h_u_cla32_and3699_y0(h_u_cla32_and3698_y0, h_u_cla32_and3697_y0, h_u_cla32_and3699_y0);
  and_gate and_gate_h_u_cla32_and3700_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3700_y0);
  and_gate and_gate_h_u_cla32_and3701_y0(h_u_cla32_and3700_y0, h_u_cla32_and3699_y0, h_u_cla32_and3701_y0);
  and_gate and_gate_h_u_cla32_and3702_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3702_y0);
  and_gate and_gate_h_u_cla32_and3703_y0(h_u_cla32_and3702_y0, h_u_cla32_and3701_y0, h_u_cla32_and3703_y0);
  and_gate and_gate_h_u_cla32_and3704_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3704_y0);
  and_gate and_gate_h_u_cla32_and3705_y0(h_u_cla32_and3704_y0, h_u_cla32_and3703_y0, h_u_cla32_and3705_y0);
  and_gate and_gate_h_u_cla32_and3706_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3706_y0);
  and_gate and_gate_h_u_cla32_and3707_y0(h_u_cla32_and3706_y0, h_u_cla32_and3705_y0, h_u_cla32_and3707_y0);
  and_gate and_gate_h_u_cla32_and3708_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3708_y0);
  and_gate and_gate_h_u_cla32_and3709_y0(h_u_cla32_and3708_y0, h_u_cla32_and3707_y0, h_u_cla32_and3709_y0);
  and_gate and_gate_h_u_cla32_and3710_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3710_y0);
  and_gate and_gate_h_u_cla32_and3711_y0(h_u_cla32_and3710_y0, h_u_cla32_and3709_y0, h_u_cla32_and3711_y0);
  and_gate and_gate_h_u_cla32_and3712_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and3712_y0);
  and_gate and_gate_h_u_cla32_and3713_y0(h_u_cla32_and3712_y0, h_u_cla32_and3711_y0, h_u_cla32_and3713_y0);
  and_gate and_gate_h_u_cla32_and3714_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3714_y0);
  and_gate and_gate_h_u_cla32_and3715_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3715_y0);
  and_gate and_gate_h_u_cla32_and3716_y0(h_u_cla32_and3715_y0, h_u_cla32_and3714_y0, h_u_cla32_and3716_y0);
  and_gate and_gate_h_u_cla32_and3717_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3717_y0);
  and_gate and_gate_h_u_cla32_and3718_y0(h_u_cla32_and3717_y0, h_u_cla32_and3716_y0, h_u_cla32_and3718_y0);
  and_gate and_gate_h_u_cla32_and3719_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3719_y0);
  and_gate and_gate_h_u_cla32_and3720_y0(h_u_cla32_and3719_y0, h_u_cla32_and3718_y0, h_u_cla32_and3720_y0);
  and_gate and_gate_h_u_cla32_and3721_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3721_y0);
  and_gate and_gate_h_u_cla32_and3722_y0(h_u_cla32_and3721_y0, h_u_cla32_and3720_y0, h_u_cla32_and3722_y0);
  and_gate and_gate_h_u_cla32_and3723_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3723_y0);
  and_gate and_gate_h_u_cla32_and3724_y0(h_u_cla32_and3723_y0, h_u_cla32_and3722_y0, h_u_cla32_and3724_y0);
  and_gate and_gate_h_u_cla32_and3725_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3725_y0);
  and_gate and_gate_h_u_cla32_and3726_y0(h_u_cla32_and3725_y0, h_u_cla32_and3724_y0, h_u_cla32_and3726_y0);
  and_gate and_gate_h_u_cla32_and3727_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3727_y0);
  and_gate and_gate_h_u_cla32_and3728_y0(h_u_cla32_and3727_y0, h_u_cla32_and3726_y0, h_u_cla32_and3728_y0);
  and_gate and_gate_h_u_cla32_and3729_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and3729_y0);
  and_gate and_gate_h_u_cla32_and3730_y0(h_u_cla32_and3729_y0, h_u_cla32_and3728_y0, h_u_cla32_and3730_y0);
  and_gate and_gate_h_u_cla32_and3731_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3731_y0);
  and_gate and_gate_h_u_cla32_and3732_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3732_y0);
  and_gate and_gate_h_u_cla32_and3733_y0(h_u_cla32_and3732_y0, h_u_cla32_and3731_y0, h_u_cla32_and3733_y0);
  and_gate and_gate_h_u_cla32_and3734_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3734_y0);
  and_gate and_gate_h_u_cla32_and3735_y0(h_u_cla32_and3734_y0, h_u_cla32_and3733_y0, h_u_cla32_and3735_y0);
  and_gate and_gate_h_u_cla32_and3736_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3736_y0);
  and_gate and_gate_h_u_cla32_and3737_y0(h_u_cla32_and3736_y0, h_u_cla32_and3735_y0, h_u_cla32_and3737_y0);
  and_gate and_gate_h_u_cla32_and3738_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3738_y0);
  and_gate and_gate_h_u_cla32_and3739_y0(h_u_cla32_and3738_y0, h_u_cla32_and3737_y0, h_u_cla32_and3739_y0);
  and_gate and_gate_h_u_cla32_and3740_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3740_y0);
  and_gate and_gate_h_u_cla32_and3741_y0(h_u_cla32_and3740_y0, h_u_cla32_and3739_y0, h_u_cla32_and3741_y0);
  and_gate and_gate_h_u_cla32_and3742_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3742_y0);
  and_gate and_gate_h_u_cla32_and3743_y0(h_u_cla32_and3742_y0, h_u_cla32_and3741_y0, h_u_cla32_and3743_y0);
  and_gate and_gate_h_u_cla32_and3744_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and3744_y0);
  and_gate and_gate_h_u_cla32_and3745_y0(h_u_cla32_and3744_y0, h_u_cla32_and3743_y0, h_u_cla32_and3745_y0);
  and_gate and_gate_h_u_cla32_and3746_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3746_y0);
  and_gate and_gate_h_u_cla32_and3747_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3747_y0);
  and_gate and_gate_h_u_cla32_and3748_y0(h_u_cla32_and3747_y0, h_u_cla32_and3746_y0, h_u_cla32_and3748_y0);
  and_gate and_gate_h_u_cla32_and3749_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3749_y0);
  and_gate and_gate_h_u_cla32_and3750_y0(h_u_cla32_and3749_y0, h_u_cla32_and3748_y0, h_u_cla32_and3750_y0);
  and_gate and_gate_h_u_cla32_and3751_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3751_y0);
  and_gate and_gate_h_u_cla32_and3752_y0(h_u_cla32_and3751_y0, h_u_cla32_and3750_y0, h_u_cla32_and3752_y0);
  and_gate and_gate_h_u_cla32_and3753_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3753_y0);
  and_gate and_gate_h_u_cla32_and3754_y0(h_u_cla32_and3753_y0, h_u_cla32_and3752_y0, h_u_cla32_and3754_y0);
  and_gate and_gate_h_u_cla32_and3755_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3755_y0);
  and_gate and_gate_h_u_cla32_and3756_y0(h_u_cla32_and3755_y0, h_u_cla32_and3754_y0, h_u_cla32_and3756_y0);
  and_gate and_gate_h_u_cla32_and3757_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and3757_y0);
  and_gate and_gate_h_u_cla32_and3758_y0(h_u_cla32_and3757_y0, h_u_cla32_and3756_y0, h_u_cla32_and3758_y0);
  and_gate and_gate_h_u_cla32_and3759_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3759_y0);
  and_gate and_gate_h_u_cla32_and3760_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3760_y0);
  and_gate and_gate_h_u_cla32_and3761_y0(h_u_cla32_and3760_y0, h_u_cla32_and3759_y0, h_u_cla32_and3761_y0);
  and_gate and_gate_h_u_cla32_and3762_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3762_y0);
  and_gate and_gate_h_u_cla32_and3763_y0(h_u_cla32_and3762_y0, h_u_cla32_and3761_y0, h_u_cla32_and3763_y0);
  and_gate and_gate_h_u_cla32_and3764_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3764_y0);
  and_gate and_gate_h_u_cla32_and3765_y0(h_u_cla32_and3764_y0, h_u_cla32_and3763_y0, h_u_cla32_and3765_y0);
  and_gate and_gate_h_u_cla32_and3766_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3766_y0);
  and_gate and_gate_h_u_cla32_and3767_y0(h_u_cla32_and3766_y0, h_u_cla32_and3765_y0, h_u_cla32_and3767_y0);
  and_gate and_gate_h_u_cla32_and3768_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and3768_y0);
  and_gate and_gate_h_u_cla32_and3769_y0(h_u_cla32_and3768_y0, h_u_cla32_and3767_y0, h_u_cla32_and3769_y0);
  and_gate and_gate_h_u_cla32_and3770_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3770_y0);
  and_gate and_gate_h_u_cla32_and3771_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3771_y0);
  and_gate and_gate_h_u_cla32_and3772_y0(h_u_cla32_and3771_y0, h_u_cla32_and3770_y0, h_u_cla32_and3772_y0);
  and_gate and_gate_h_u_cla32_and3773_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3773_y0);
  and_gate and_gate_h_u_cla32_and3774_y0(h_u_cla32_and3773_y0, h_u_cla32_and3772_y0, h_u_cla32_and3774_y0);
  and_gate and_gate_h_u_cla32_and3775_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3775_y0);
  and_gate and_gate_h_u_cla32_and3776_y0(h_u_cla32_and3775_y0, h_u_cla32_and3774_y0, h_u_cla32_and3776_y0);
  and_gate and_gate_h_u_cla32_and3777_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and3777_y0);
  and_gate and_gate_h_u_cla32_and3778_y0(h_u_cla32_and3777_y0, h_u_cla32_and3776_y0, h_u_cla32_and3778_y0);
  and_gate and_gate_h_u_cla32_and3779_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3779_y0);
  and_gate and_gate_h_u_cla32_and3780_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3780_y0);
  and_gate and_gate_h_u_cla32_and3781_y0(h_u_cla32_and3780_y0, h_u_cla32_and3779_y0, h_u_cla32_and3781_y0);
  and_gate and_gate_h_u_cla32_and3782_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3782_y0);
  and_gate and_gate_h_u_cla32_and3783_y0(h_u_cla32_and3782_y0, h_u_cla32_and3781_y0, h_u_cla32_and3783_y0);
  and_gate and_gate_h_u_cla32_and3784_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and3784_y0);
  and_gate and_gate_h_u_cla32_and3785_y0(h_u_cla32_and3784_y0, h_u_cla32_and3783_y0, h_u_cla32_and3785_y0);
  and_gate and_gate_h_u_cla32_and3786_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and3786_y0);
  and_gate and_gate_h_u_cla32_and3787_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and3787_y0);
  and_gate and_gate_h_u_cla32_and3788_y0(h_u_cla32_and3787_y0, h_u_cla32_and3786_y0, h_u_cla32_and3788_y0);
  and_gate and_gate_h_u_cla32_and3789_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and3789_y0);
  and_gate and_gate_h_u_cla32_and3790_y0(h_u_cla32_and3789_y0, h_u_cla32_and3788_y0, h_u_cla32_and3790_y0);
  and_gate and_gate_h_u_cla32_and3791_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and3791_y0);
  and_gate and_gate_h_u_cla32_and3792_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and3792_y0);
  and_gate and_gate_h_u_cla32_and3793_y0(h_u_cla32_and3792_y0, h_u_cla32_and3791_y0, h_u_cla32_and3793_y0);
  and_gate and_gate_h_u_cla32_and3794_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and3794_y0);
  or_gate or_gate_h_u_cla32_or231_y0(h_u_cla32_and3794_y0, h_u_cla32_and3353_y0, h_u_cla32_or231_y0);
  or_gate or_gate_h_u_cla32_or232_y0(h_u_cla32_or231_y0, h_u_cla32_and3394_y0, h_u_cla32_or232_y0);
  or_gate or_gate_h_u_cla32_or233_y0(h_u_cla32_or232_y0, h_u_cla32_and3433_y0, h_u_cla32_or233_y0);
  or_gate or_gate_h_u_cla32_or234_y0(h_u_cla32_or233_y0, h_u_cla32_and3470_y0, h_u_cla32_or234_y0);
  or_gate or_gate_h_u_cla32_or235_y0(h_u_cla32_or234_y0, h_u_cla32_and3505_y0, h_u_cla32_or235_y0);
  or_gate or_gate_h_u_cla32_or236_y0(h_u_cla32_or235_y0, h_u_cla32_and3538_y0, h_u_cla32_or236_y0);
  or_gate or_gate_h_u_cla32_or237_y0(h_u_cla32_or236_y0, h_u_cla32_and3569_y0, h_u_cla32_or237_y0);
  or_gate or_gate_h_u_cla32_or238_y0(h_u_cla32_or237_y0, h_u_cla32_and3598_y0, h_u_cla32_or238_y0);
  or_gate or_gate_h_u_cla32_or239_y0(h_u_cla32_or238_y0, h_u_cla32_and3625_y0, h_u_cla32_or239_y0);
  or_gate or_gate_h_u_cla32_or240_y0(h_u_cla32_or239_y0, h_u_cla32_and3650_y0, h_u_cla32_or240_y0);
  or_gate or_gate_h_u_cla32_or241_y0(h_u_cla32_or240_y0, h_u_cla32_and3673_y0, h_u_cla32_or241_y0);
  or_gate or_gate_h_u_cla32_or242_y0(h_u_cla32_or241_y0, h_u_cla32_and3694_y0, h_u_cla32_or242_y0);
  or_gate or_gate_h_u_cla32_or243_y0(h_u_cla32_or242_y0, h_u_cla32_and3713_y0, h_u_cla32_or243_y0);
  or_gate or_gate_h_u_cla32_or244_y0(h_u_cla32_or243_y0, h_u_cla32_and3730_y0, h_u_cla32_or244_y0);
  or_gate or_gate_h_u_cla32_or245_y0(h_u_cla32_or244_y0, h_u_cla32_and3745_y0, h_u_cla32_or245_y0);
  or_gate or_gate_h_u_cla32_or246_y0(h_u_cla32_or245_y0, h_u_cla32_and3758_y0, h_u_cla32_or246_y0);
  or_gate or_gate_h_u_cla32_or247_y0(h_u_cla32_or246_y0, h_u_cla32_and3769_y0, h_u_cla32_or247_y0);
  or_gate or_gate_h_u_cla32_or248_y0(h_u_cla32_or247_y0, h_u_cla32_and3778_y0, h_u_cla32_or248_y0);
  or_gate or_gate_h_u_cla32_or249_y0(h_u_cla32_or248_y0, h_u_cla32_and3785_y0, h_u_cla32_or249_y0);
  or_gate or_gate_h_u_cla32_or250_y0(h_u_cla32_or249_y0, h_u_cla32_and3790_y0, h_u_cla32_or250_y0);
  or_gate or_gate_h_u_cla32_or251_y0(h_u_cla32_or250_y0, h_u_cla32_and3793_y0, h_u_cla32_or251_y0);
  or_gate or_gate_h_u_cla32_or252_y0(h_u_cla32_pg_logic21_y1, h_u_cla32_or251_y0, h_u_cla32_or252_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic22_y0(a_22, b_22, h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_pg_logic22_y2);
  xor_gate xor_gate_h_u_cla32_xor22_y0(h_u_cla32_pg_logic22_y2, h_u_cla32_or252_y0, h_u_cla32_xor22_y0);
  and_gate and_gate_h_u_cla32_and3795_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and3795_y0);
  and_gate and_gate_h_u_cla32_and3796_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and3796_y0);
  and_gate and_gate_h_u_cla32_and3797_y0(h_u_cla32_and3796_y0, h_u_cla32_and3795_y0, h_u_cla32_and3797_y0);
  and_gate and_gate_h_u_cla32_and3798_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and3798_y0);
  and_gate and_gate_h_u_cla32_and3799_y0(h_u_cla32_and3798_y0, h_u_cla32_and3797_y0, h_u_cla32_and3799_y0);
  and_gate and_gate_h_u_cla32_and3800_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and3800_y0);
  and_gate and_gate_h_u_cla32_and3801_y0(h_u_cla32_and3800_y0, h_u_cla32_and3799_y0, h_u_cla32_and3801_y0);
  and_gate and_gate_h_u_cla32_and3802_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and3802_y0);
  and_gate and_gate_h_u_cla32_and3803_y0(h_u_cla32_and3802_y0, h_u_cla32_and3801_y0, h_u_cla32_and3803_y0);
  and_gate and_gate_h_u_cla32_and3804_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and3804_y0);
  and_gate and_gate_h_u_cla32_and3805_y0(h_u_cla32_and3804_y0, h_u_cla32_and3803_y0, h_u_cla32_and3805_y0);
  and_gate and_gate_h_u_cla32_and3806_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and3806_y0);
  and_gate and_gate_h_u_cla32_and3807_y0(h_u_cla32_and3806_y0, h_u_cla32_and3805_y0, h_u_cla32_and3807_y0);
  and_gate and_gate_h_u_cla32_and3808_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and3808_y0);
  and_gate and_gate_h_u_cla32_and3809_y0(h_u_cla32_and3808_y0, h_u_cla32_and3807_y0, h_u_cla32_and3809_y0);
  and_gate and_gate_h_u_cla32_and3810_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and3810_y0);
  and_gate and_gate_h_u_cla32_and3811_y0(h_u_cla32_and3810_y0, h_u_cla32_and3809_y0, h_u_cla32_and3811_y0);
  and_gate and_gate_h_u_cla32_and3812_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and3812_y0);
  and_gate and_gate_h_u_cla32_and3813_y0(h_u_cla32_and3812_y0, h_u_cla32_and3811_y0, h_u_cla32_and3813_y0);
  and_gate and_gate_h_u_cla32_and3814_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and3814_y0);
  and_gate and_gate_h_u_cla32_and3815_y0(h_u_cla32_and3814_y0, h_u_cla32_and3813_y0, h_u_cla32_and3815_y0);
  and_gate and_gate_h_u_cla32_and3816_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and3816_y0);
  and_gate and_gate_h_u_cla32_and3817_y0(h_u_cla32_and3816_y0, h_u_cla32_and3815_y0, h_u_cla32_and3817_y0);
  and_gate and_gate_h_u_cla32_and3818_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and3818_y0);
  and_gate and_gate_h_u_cla32_and3819_y0(h_u_cla32_and3818_y0, h_u_cla32_and3817_y0, h_u_cla32_and3819_y0);
  and_gate and_gate_h_u_cla32_and3820_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and3820_y0);
  and_gate and_gate_h_u_cla32_and3821_y0(h_u_cla32_and3820_y0, h_u_cla32_and3819_y0, h_u_cla32_and3821_y0);
  and_gate and_gate_h_u_cla32_and3822_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and3822_y0);
  and_gate and_gate_h_u_cla32_and3823_y0(h_u_cla32_and3822_y0, h_u_cla32_and3821_y0, h_u_cla32_and3823_y0);
  and_gate and_gate_h_u_cla32_and3824_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and3824_y0);
  and_gate and_gate_h_u_cla32_and3825_y0(h_u_cla32_and3824_y0, h_u_cla32_and3823_y0, h_u_cla32_and3825_y0);
  and_gate and_gate_h_u_cla32_and3826_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and3826_y0);
  and_gate and_gate_h_u_cla32_and3827_y0(h_u_cla32_and3826_y0, h_u_cla32_and3825_y0, h_u_cla32_and3827_y0);
  and_gate and_gate_h_u_cla32_and3828_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and3828_y0);
  and_gate and_gate_h_u_cla32_and3829_y0(h_u_cla32_and3828_y0, h_u_cla32_and3827_y0, h_u_cla32_and3829_y0);
  and_gate and_gate_h_u_cla32_and3830_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and3830_y0);
  and_gate and_gate_h_u_cla32_and3831_y0(h_u_cla32_and3830_y0, h_u_cla32_and3829_y0, h_u_cla32_and3831_y0);
  and_gate and_gate_h_u_cla32_and3832_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and3832_y0);
  and_gate and_gate_h_u_cla32_and3833_y0(h_u_cla32_and3832_y0, h_u_cla32_and3831_y0, h_u_cla32_and3833_y0);
  and_gate and_gate_h_u_cla32_and3834_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and3834_y0);
  and_gate and_gate_h_u_cla32_and3835_y0(h_u_cla32_and3834_y0, h_u_cla32_and3833_y0, h_u_cla32_and3835_y0);
  and_gate and_gate_h_u_cla32_and3836_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and3836_y0);
  and_gate and_gate_h_u_cla32_and3837_y0(h_u_cla32_and3836_y0, h_u_cla32_and3835_y0, h_u_cla32_and3837_y0);
  and_gate and_gate_h_u_cla32_and3838_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and3838_y0);
  and_gate and_gate_h_u_cla32_and3839_y0(h_u_cla32_and3838_y0, h_u_cla32_and3837_y0, h_u_cla32_and3839_y0);
  and_gate and_gate_h_u_cla32_and3840_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3840_y0);
  and_gate and_gate_h_u_cla32_and3841_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3841_y0);
  and_gate and_gate_h_u_cla32_and3842_y0(h_u_cla32_and3841_y0, h_u_cla32_and3840_y0, h_u_cla32_and3842_y0);
  and_gate and_gate_h_u_cla32_and3843_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3843_y0);
  and_gate and_gate_h_u_cla32_and3844_y0(h_u_cla32_and3843_y0, h_u_cla32_and3842_y0, h_u_cla32_and3844_y0);
  and_gate and_gate_h_u_cla32_and3845_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3845_y0);
  and_gate and_gate_h_u_cla32_and3846_y0(h_u_cla32_and3845_y0, h_u_cla32_and3844_y0, h_u_cla32_and3846_y0);
  and_gate and_gate_h_u_cla32_and3847_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3847_y0);
  and_gate and_gate_h_u_cla32_and3848_y0(h_u_cla32_and3847_y0, h_u_cla32_and3846_y0, h_u_cla32_and3848_y0);
  and_gate and_gate_h_u_cla32_and3849_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3849_y0);
  and_gate and_gate_h_u_cla32_and3850_y0(h_u_cla32_and3849_y0, h_u_cla32_and3848_y0, h_u_cla32_and3850_y0);
  and_gate and_gate_h_u_cla32_and3851_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3851_y0);
  and_gate and_gate_h_u_cla32_and3852_y0(h_u_cla32_and3851_y0, h_u_cla32_and3850_y0, h_u_cla32_and3852_y0);
  and_gate and_gate_h_u_cla32_and3853_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3853_y0);
  and_gate and_gate_h_u_cla32_and3854_y0(h_u_cla32_and3853_y0, h_u_cla32_and3852_y0, h_u_cla32_and3854_y0);
  and_gate and_gate_h_u_cla32_and3855_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3855_y0);
  and_gate and_gate_h_u_cla32_and3856_y0(h_u_cla32_and3855_y0, h_u_cla32_and3854_y0, h_u_cla32_and3856_y0);
  and_gate and_gate_h_u_cla32_and3857_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3857_y0);
  and_gate and_gate_h_u_cla32_and3858_y0(h_u_cla32_and3857_y0, h_u_cla32_and3856_y0, h_u_cla32_and3858_y0);
  and_gate and_gate_h_u_cla32_and3859_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3859_y0);
  and_gate and_gate_h_u_cla32_and3860_y0(h_u_cla32_and3859_y0, h_u_cla32_and3858_y0, h_u_cla32_and3860_y0);
  and_gate and_gate_h_u_cla32_and3861_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3861_y0);
  and_gate and_gate_h_u_cla32_and3862_y0(h_u_cla32_and3861_y0, h_u_cla32_and3860_y0, h_u_cla32_and3862_y0);
  and_gate and_gate_h_u_cla32_and3863_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3863_y0);
  and_gate and_gate_h_u_cla32_and3864_y0(h_u_cla32_and3863_y0, h_u_cla32_and3862_y0, h_u_cla32_and3864_y0);
  and_gate and_gate_h_u_cla32_and3865_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3865_y0);
  and_gate and_gate_h_u_cla32_and3866_y0(h_u_cla32_and3865_y0, h_u_cla32_and3864_y0, h_u_cla32_and3866_y0);
  and_gate and_gate_h_u_cla32_and3867_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3867_y0);
  and_gate and_gate_h_u_cla32_and3868_y0(h_u_cla32_and3867_y0, h_u_cla32_and3866_y0, h_u_cla32_and3868_y0);
  and_gate and_gate_h_u_cla32_and3869_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3869_y0);
  and_gate and_gate_h_u_cla32_and3870_y0(h_u_cla32_and3869_y0, h_u_cla32_and3868_y0, h_u_cla32_and3870_y0);
  and_gate and_gate_h_u_cla32_and3871_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3871_y0);
  and_gate and_gate_h_u_cla32_and3872_y0(h_u_cla32_and3871_y0, h_u_cla32_and3870_y0, h_u_cla32_and3872_y0);
  and_gate and_gate_h_u_cla32_and3873_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3873_y0);
  and_gate and_gate_h_u_cla32_and3874_y0(h_u_cla32_and3873_y0, h_u_cla32_and3872_y0, h_u_cla32_and3874_y0);
  and_gate and_gate_h_u_cla32_and3875_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3875_y0);
  and_gate and_gate_h_u_cla32_and3876_y0(h_u_cla32_and3875_y0, h_u_cla32_and3874_y0, h_u_cla32_and3876_y0);
  and_gate and_gate_h_u_cla32_and3877_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3877_y0);
  and_gate and_gate_h_u_cla32_and3878_y0(h_u_cla32_and3877_y0, h_u_cla32_and3876_y0, h_u_cla32_and3878_y0);
  and_gate and_gate_h_u_cla32_and3879_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3879_y0);
  and_gate and_gate_h_u_cla32_and3880_y0(h_u_cla32_and3879_y0, h_u_cla32_and3878_y0, h_u_cla32_and3880_y0);
  and_gate and_gate_h_u_cla32_and3881_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and3881_y0);
  and_gate and_gate_h_u_cla32_and3882_y0(h_u_cla32_and3881_y0, h_u_cla32_and3880_y0, h_u_cla32_and3882_y0);
  and_gate and_gate_h_u_cla32_and3883_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3883_y0);
  and_gate and_gate_h_u_cla32_and3884_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3884_y0);
  and_gate and_gate_h_u_cla32_and3885_y0(h_u_cla32_and3884_y0, h_u_cla32_and3883_y0, h_u_cla32_and3885_y0);
  and_gate and_gate_h_u_cla32_and3886_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3886_y0);
  and_gate and_gate_h_u_cla32_and3887_y0(h_u_cla32_and3886_y0, h_u_cla32_and3885_y0, h_u_cla32_and3887_y0);
  and_gate and_gate_h_u_cla32_and3888_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3888_y0);
  and_gate and_gate_h_u_cla32_and3889_y0(h_u_cla32_and3888_y0, h_u_cla32_and3887_y0, h_u_cla32_and3889_y0);
  and_gate and_gate_h_u_cla32_and3890_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3890_y0);
  and_gate and_gate_h_u_cla32_and3891_y0(h_u_cla32_and3890_y0, h_u_cla32_and3889_y0, h_u_cla32_and3891_y0);
  and_gate and_gate_h_u_cla32_and3892_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3892_y0);
  and_gate and_gate_h_u_cla32_and3893_y0(h_u_cla32_and3892_y0, h_u_cla32_and3891_y0, h_u_cla32_and3893_y0);
  and_gate and_gate_h_u_cla32_and3894_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3894_y0);
  and_gate and_gate_h_u_cla32_and3895_y0(h_u_cla32_and3894_y0, h_u_cla32_and3893_y0, h_u_cla32_and3895_y0);
  and_gate and_gate_h_u_cla32_and3896_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3896_y0);
  and_gate and_gate_h_u_cla32_and3897_y0(h_u_cla32_and3896_y0, h_u_cla32_and3895_y0, h_u_cla32_and3897_y0);
  and_gate and_gate_h_u_cla32_and3898_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3898_y0);
  and_gate and_gate_h_u_cla32_and3899_y0(h_u_cla32_and3898_y0, h_u_cla32_and3897_y0, h_u_cla32_and3899_y0);
  and_gate and_gate_h_u_cla32_and3900_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3900_y0);
  and_gate and_gate_h_u_cla32_and3901_y0(h_u_cla32_and3900_y0, h_u_cla32_and3899_y0, h_u_cla32_and3901_y0);
  and_gate and_gate_h_u_cla32_and3902_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3902_y0);
  and_gate and_gate_h_u_cla32_and3903_y0(h_u_cla32_and3902_y0, h_u_cla32_and3901_y0, h_u_cla32_and3903_y0);
  and_gate and_gate_h_u_cla32_and3904_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3904_y0);
  and_gate and_gate_h_u_cla32_and3905_y0(h_u_cla32_and3904_y0, h_u_cla32_and3903_y0, h_u_cla32_and3905_y0);
  and_gate and_gate_h_u_cla32_and3906_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3906_y0);
  and_gate and_gate_h_u_cla32_and3907_y0(h_u_cla32_and3906_y0, h_u_cla32_and3905_y0, h_u_cla32_and3907_y0);
  and_gate and_gate_h_u_cla32_and3908_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3908_y0);
  and_gate and_gate_h_u_cla32_and3909_y0(h_u_cla32_and3908_y0, h_u_cla32_and3907_y0, h_u_cla32_and3909_y0);
  and_gate and_gate_h_u_cla32_and3910_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3910_y0);
  and_gate and_gate_h_u_cla32_and3911_y0(h_u_cla32_and3910_y0, h_u_cla32_and3909_y0, h_u_cla32_and3911_y0);
  and_gate and_gate_h_u_cla32_and3912_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3912_y0);
  and_gate and_gate_h_u_cla32_and3913_y0(h_u_cla32_and3912_y0, h_u_cla32_and3911_y0, h_u_cla32_and3913_y0);
  and_gate and_gate_h_u_cla32_and3914_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3914_y0);
  and_gate and_gate_h_u_cla32_and3915_y0(h_u_cla32_and3914_y0, h_u_cla32_and3913_y0, h_u_cla32_and3915_y0);
  and_gate and_gate_h_u_cla32_and3916_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3916_y0);
  and_gate and_gate_h_u_cla32_and3917_y0(h_u_cla32_and3916_y0, h_u_cla32_and3915_y0, h_u_cla32_and3917_y0);
  and_gate and_gate_h_u_cla32_and3918_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3918_y0);
  and_gate and_gate_h_u_cla32_and3919_y0(h_u_cla32_and3918_y0, h_u_cla32_and3917_y0, h_u_cla32_and3919_y0);
  and_gate and_gate_h_u_cla32_and3920_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3920_y0);
  and_gate and_gate_h_u_cla32_and3921_y0(h_u_cla32_and3920_y0, h_u_cla32_and3919_y0, h_u_cla32_and3921_y0);
  and_gate and_gate_h_u_cla32_and3922_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and3922_y0);
  and_gate and_gate_h_u_cla32_and3923_y0(h_u_cla32_and3922_y0, h_u_cla32_and3921_y0, h_u_cla32_and3923_y0);
  and_gate and_gate_h_u_cla32_and3924_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3924_y0);
  and_gate and_gate_h_u_cla32_and3925_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3925_y0);
  and_gate and_gate_h_u_cla32_and3926_y0(h_u_cla32_and3925_y0, h_u_cla32_and3924_y0, h_u_cla32_and3926_y0);
  and_gate and_gate_h_u_cla32_and3927_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3927_y0);
  and_gate and_gate_h_u_cla32_and3928_y0(h_u_cla32_and3927_y0, h_u_cla32_and3926_y0, h_u_cla32_and3928_y0);
  and_gate and_gate_h_u_cla32_and3929_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3929_y0);
  and_gate and_gate_h_u_cla32_and3930_y0(h_u_cla32_and3929_y0, h_u_cla32_and3928_y0, h_u_cla32_and3930_y0);
  and_gate and_gate_h_u_cla32_and3931_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3931_y0);
  and_gate and_gate_h_u_cla32_and3932_y0(h_u_cla32_and3931_y0, h_u_cla32_and3930_y0, h_u_cla32_and3932_y0);
  and_gate and_gate_h_u_cla32_and3933_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3933_y0);
  and_gate and_gate_h_u_cla32_and3934_y0(h_u_cla32_and3933_y0, h_u_cla32_and3932_y0, h_u_cla32_and3934_y0);
  and_gate and_gate_h_u_cla32_and3935_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3935_y0);
  and_gate and_gate_h_u_cla32_and3936_y0(h_u_cla32_and3935_y0, h_u_cla32_and3934_y0, h_u_cla32_and3936_y0);
  and_gate and_gate_h_u_cla32_and3937_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3937_y0);
  and_gate and_gate_h_u_cla32_and3938_y0(h_u_cla32_and3937_y0, h_u_cla32_and3936_y0, h_u_cla32_and3938_y0);
  and_gate and_gate_h_u_cla32_and3939_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3939_y0);
  and_gate and_gate_h_u_cla32_and3940_y0(h_u_cla32_and3939_y0, h_u_cla32_and3938_y0, h_u_cla32_and3940_y0);
  and_gate and_gate_h_u_cla32_and3941_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3941_y0);
  and_gate and_gate_h_u_cla32_and3942_y0(h_u_cla32_and3941_y0, h_u_cla32_and3940_y0, h_u_cla32_and3942_y0);
  and_gate and_gate_h_u_cla32_and3943_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3943_y0);
  and_gate and_gate_h_u_cla32_and3944_y0(h_u_cla32_and3943_y0, h_u_cla32_and3942_y0, h_u_cla32_and3944_y0);
  and_gate and_gate_h_u_cla32_and3945_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3945_y0);
  and_gate and_gate_h_u_cla32_and3946_y0(h_u_cla32_and3945_y0, h_u_cla32_and3944_y0, h_u_cla32_and3946_y0);
  and_gate and_gate_h_u_cla32_and3947_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3947_y0);
  and_gate and_gate_h_u_cla32_and3948_y0(h_u_cla32_and3947_y0, h_u_cla32_and3946_y0, h_u_cla32_and3948_y0);
  and_gate and_gate_h_u_cla32_and3949_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3949_y0);
  and_gate and_gate_h_u_cla32_and3950_y0(h_u_cla32_and3949_y0, h_u_cla32_and3948_y0, h_u_cla32_and3950_y0);
  and_gate and_gate_h_u_cla32_and3951_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3951_y0);
  and_gate and_gate_h_u_cla32_and3952_y0(h_u_cla32_and3951_y0, h_u_cla32_and3950_y0, h_u_cla32_and3952_y0);
  and_gate and_gate_h_u_cla32_and3953_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3953_y0);
  and_gate and_gate_h_u_cla32_and3954_y0(h_u_cla32_and3953_y0, h_u_cla32_and3952_y0, h_u_cla32_and3954_y0);
  and_gate and_gate_h_u_cla32_and3955_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3955_y0);
  and_gate and_gate_h_u_cla32_and3956_y0(h_u_cla32_and3955_y0, h_u_cla32_and3954_y0, h_u_cla32_and3956_y0);
  and_gate and_gate_h_u_cla32_and3957_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3957_y0);
  and_gate and_gate_h_u_cla32_and3958_y0(h_u_cla32_and3957_y0, h_u_cla32_and3956_y0, h_u_cla32_and3958_y0);
  and_gate and_gate_h_u_cla32_and3959_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3959_y0);
  and_gate and_gate_h_u_cla32_and3960_y0(h_u_cla32_and3959_y0, h_u_cla32_and3958_y0, h_u_cla32_and3960_y0);
  and_gate and_gate_h_u_cla32_and3961_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and3961_y0);
  and_gate and_gate_h_u_cla32_and3962_y0(h_u_cla32_and3961_y0, h_u_cla32_and3960_y0, h_u_cla32_and3962_y0);
  and_gate and_gate_h_u_cla32_and3963_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3963_y0);
  and_gate and_gate_h_u_cla32_and3964_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3964_y0);
  and_gate and_gate_h_u_cla32_and3965_y0(h_u_cla32_and3964_y0, h_u_cla32_and3963_y0, h_u_cla32_and3965_y0);
  and_gate and_gate_h_u_cla32_and3966_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3966_y0);
  and_gate and_gate_h_u_cla32_and3967_y0(h_u_cla32_and3966_y0, h_u_cla32_and3965_y0, h_u_cla32_and3967_y0);
  and_gate and_gate_h_u_cla32_and3968_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3968_y0);
  and_gate and_gate_h_u_cla32_and3969_y0(h_u_cla32_and3968_y0, h_u_cla32_and3967_y0, h_u_cla32_and3969_y0);
  and_gate and_gate_h_u_cla32_and3970_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3970_y0);
  and_gate and_gate_h_u_cla32_and3971_y0(h_u_cla32_and3970_y0, h_u_cla32_and3969_y0, h_u_cla32_and3971_y0);
  and_gate and_gate_h_u_cla32_and3972_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3972_y0);
  and_gate and_gate_h_u_cla32_and3973_y0(h_u_cla32_and3972_y0, h_u_cla32_and3971_y0, h_u_cla32_and3973_y0);
  and_gate and_gate_h_u_cla32_and3974_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3974_y0);
  and_gate and_gate_h_u_cla32_and3975_y0(h_u_cla32_and3974_y0, h_u_cla32_and3973_y0, h_u_cla32_and3975_y0);
  and_gate and_gate_h_u_cla32_and3976_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3976_y0);
  and_gate and_gate_h_u_cla32_and3977_y0(h_u_cla32_and3976_y0, h_u_cla32_and3975_y0, h_u_cla32_and3977_y0);
  and_gate and_gate_h_u_cla32_and3978_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3978_y0);
  and_gate and_gate_h_u_cla32_and3979_y0(h_u_cla32_and3978_y0, h_u_cla32_and3977_y0, h_u_cla32_and3979_y0);
  and_gate and_gate_h_u_cla32_and3980_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3980_y0);
  and_gate and_gate_h_u_cla32_and3981_y0(h_u_cla32_and3980_y0, h_u_cla32_and3979_y0, h_u_cla32_and3981_y0);
  and_gate and_gate_h_u_cla32_and3982_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3982_y0);
  and_gate and_gate_h_u_cla32_and3983_y0(h_u_cla32_and3982_y0, h_u_cla32_and3981_y0, h_u_cla32_and3983_y0);
  and_gate and_gate_h_u_cla32_and3984_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3984_y0);
  and_gate and_gate_h_u_cla32_and3985_y0(h_u_cla32_and3984_y0, h_u_cla32_and3983_y0, h_u_cla32_and3985_y0);
  and_gate and_gate_h_u_cla32_and3986_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3986_y0);
  and_gate and_gate_h_u_cla32_and3987_y0(h_u_cla32_and3986_y0, h_u_cla32_and3985_y0, h_u_cla32_and3987_y0);
  and_gate and_gate_h_u_cla32_and3988_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3988_y0);
  and_gate and_gate_h_u_cla32_and3989_y0(h_u_cla32_and3988_y0, h_u_cla32_and3987_y0, h_u_cla32_and3989_y0);
  and_gate and_gate_h_u_cla32_and3990_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3990_y0);
  and_gate and_gate_h_u_cla32_and3991_y0(h_u_cla32_and3990_y0, h_u_cla32_and3989_y0, h_u_cla32_and3991_y0);
  and_gate and_gate_h_u_cla32_and3992_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3992_y0);
  and_gate and_gate_h_u_cla32_and3993_y0(h_u_cla32_and3992_y0, h_u_cla32_and3991_y0, h_u_cla32_and3993_y0);
  and_gate and_gate_h_u_cla32_and3994_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3994_y0);
  and_gate and_gate_h_u_cla32_and3995_y0(h_u_cla32_and3994_y0, h_u_cla32_and3993_y0, h_u_cla32_and3995_y0);
  and_gate and_gate_h_u_cla32_and3996_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3996_y0);
  and_gate and_gate_h_u_cla32_and3997_y0(h_u_cla32_and3996_y0, h_u_cla32_and3995_y0, h_u_cla32_and3997_y0);
  and_gate and_gate_h_u_cla32_and3998_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and3998_y0);
  and_gate and_gate_h_u_cla32_and3999_y0(h_u_cla32_and3998_y0, h_u_cla32_and3997_y0, h_u_cla32_and3999_y0);
  and_gate and_gate_h_u_cla32_and4000_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4000_y0);
  and_gate and_gate_h_u_cla32_and4001_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4001_y0);
  and_gate and_gate_h_u_cla32_and4002_y0(h_u_cla32_and4001_y0, h_u_cla32_and4000_y0, h_u_cla32_and4002_y0);
  and_gate and_gate_h_u_cla32_and4003_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4003_y0);
  and_gate and_gate_h_u_cla32_and4004_y0(h_u_cla32_and4003_y0, h_u_cla32_and4002_y0, h_u_cla32_and4004_y0);
  and_gate and_gate_h_u_cla32_and4005_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4005_y0);
  and_gate and_gate_h_u_cla32_and4006_y0(h_u_cla32_and4005_y0, h_u_cla32_and4004_y0, h_u_cla32_and4006_y0);
  and_gate and_gate_h_u_cla32_and4007_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4007_y0);
  and_gate and_gate_h_u_cla32_and4008_y0(h_u_cla32_and4007_y0, h_u_cla32_and4006_y0, h_u_cla32_and4008_y0);
  and_gate and_gate_h_u_cla32_and4009_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4009_y0);
  and_gate and_gate_h_u_cla32_and4010_y0(h_u_cla32_and4009_y0, h_u_cla32_and4008_y0, h_u_cla32_and4010_y0);
  and_gate and_gate_h_u_cla32_and4011_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4011_y0);
  and_gate and_gate_h_u_cla32_and4012_y0(h_u_cla32_and4011_y0, h_u_cla32_and4010_y0, h_u_cla32_and4012_y0);
  and_gate and_gate_h_u_cla32_and4013_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4013_y0);
  and_gate and_gate_h_u_cla32_and4014_y0(h_u_cla32_and4013_y0, h_u_cla32_and4012_y0, h_u_cla32_and4014_y0);
  and_gate and_gate_h_u_cla32_and4015_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4015_y0);
  and_gate and_gate_h_u_cla32_and4016_y0(h_u_cla32_and4015_y0, h_u_cla32_and4014_y0, h_u_cla32_and4016_y0);
  and_gate and_gate_h_u_cla32_and4017_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4017_y0);
  and_gate and_gate_h_u_cla32_and4018_y0(h_u_cla32_and4017_y0, h_u_cla32_and4016_y0, h_u_cla32_and4018_y0);
  and_gate and_gate_h_u_cla32_and4019_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4019_y0);
  and_gate and_gate_h_u_cla32_and4020_y0(h_u_cla32_and4019_y0, h_u_cla32_and4018_y0, h_u_cla32_and4020_y0);
  and_gate and_gate_h_u_cla32_and4021_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4021_y0);
  and_gate and_gate_h_u_cla32_and4022_y0(h_u_cla32_and4021_y0, h_u_cla32_and4020_y0, h_u_cla32_and4022_y0);
  and_gate and_gate_h_u_cla32_and4023_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4023_y0);
  and_gate and_gate_h_u_cla32_and4024_y0(h_u_cla32_and4023_y0, h_u_cla32_and4022_y0, h_u_cla32_and4024_y0);
  and_gate and_gate_h_u_cla32_and4025_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4025_y0);
  and_gate and_gate_h_u_cla32_and4026_y0(h_u_cla32_and4025_y0, h_u_cla32_and4024_y0, h_u_cla32_and4026_y0);
  and_gate and_gate_h_u_cla32_and4027_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4027_y0);
  and_gate and_gate_h_u_cla32_and4028_y0(h_u_cla32_and4027_y0, h_u_cla32_and4026_y0, h_u_cla32_and4028_y0);
  and_gate and_gate_h_u_cla32_and4029_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4029_y0);
  and_gate and_gate_h_u_cla32_and4030_y0(h_u_cla32_and4029_y0, h_u_cla32_and4028_y0, h_u_cla32_and4030_y0);
  and_gate and_gate_h_u_cla32_and4031_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4031_y0);
  and_gate and_gate_h_u_cla32_and4032_y0(h_u_cla32_and4031_y0, h_u_cla32_and4030_y0, h_u_cla32_and4032_y0);
  and_gate and_gate_h_u_cla32_and4033_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4033_y0);
  and_gate and_gate_h_u_cla32_and4034_y0(h_u_cla32_and4033_y0, h_u_cla32_and4032_y0, h_u_cla32_and4034_y0);
  and_gate and_gate_h_u_cla32_and4035_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4035_y0);
  and_gate and_gate_h_u_cla32_and4036_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4036_y0);
  and_gate and_gate_h_u_cla32_and4037_y0(h_u_cla32_and4036_y0, h_u_cla32_and4035_y0, h_u_cla32_and4037_y0);
  and_gate and_gate_h_u_cla32_and4038_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4038_y0);
  and_gate and_gate_h_u_cla32_and4039_y0(h_u_cla32_and4038_y0, h_u_cla32_and4037_y0, h_u_cla32_and4039_y0);
  and_gate and_gate_h_u_cla32_and4040_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4040_y0);
  and_gate and_gate_h_u_cla32_and4041_y0(h_u_cla32_and4040_y0, h_u_cla32_and4039_y0, h_u_cla32_and4041_y0);
  and_gate and_gate_h_u_cla32_and4042_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4042_y0);
  and_gate and_gate_h_u_cla32_and4043_y0(h_u_cla32_and4042_y0, h_u_cla32_and4041_y0, h_u_cla32_and4043_y0);
  and_gate and_gate_h_u_cla32_and4044_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4044_y0);
  and_gate and_gate_h_u_cla32_and4045_y0(h_u_cla32_and4044_y0, h_u_cla32_and4043_y0, h_u_cla32_and4045_y0);
  and_gate and_gate_h_u_cla32_and4046_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4046_y0);
  and_gate and_gate_h_u_cla32_and4047_y0(h_u_cla32_and4046_y0, h_u_cla32_and4045_y0, h_u_cla32_and4047_y0);
  and_gate and_gate_h_u_cla32_and4048_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4048_y0);
  and_gate and_gate_h_u_cla32_and4049_y0(h_u_cla32_and4048_y0, h_u_cla32_and4047_y0, h_u_cla32_and4049_y0);
  and_gate and_gate_h_u_cla32_and4050_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4050_y0);
  and_gate and_gate_h_u_cla32_and4051_y0(h_u_cla32_and4050_y0, h_u_cla32_and4049_y0, h_u_cla32_and4051_y0);
  and_gate and_gate_h_u_cla32_and4052_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4052_y0);
  and_gate and_gate_h_u_cla32_and4053_y0(h_u_cla32_and4052_y0, h_u_cla32_and4051_y0, h_u_cla32_and4053_y0);
  and_gate and_gate_h_u_cla32_and4054_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4054_y0);
  and_gate and_gate_h_u_cla32_and4055_y0(h_u_cla32_and4054_y0, h_u_cla32_and4053_y0, h_u_cla32_and4055_y0);
  and_gate and_gate_h_u_cla32_and4056_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4056_y0);
  and_gate and_gate_h_u_cla32_and4057_y0(h_u_cla32_and4056_y0, h_u_cla32_and4055_y0, h_u_cla32_and4057_y0);
  and_gate and_gate_h_u_cla32_and4058_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4058_y0);
  and_gate and_gate_h_u_cla32_and4059_y0(h_u_cla32_and4058_y0, h_u_cla32_and4057_y0, h_u_cla32_and4059_y0);
  and_gate and_gate_h_u_cla32_and4060_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4060_y0);
  and_gate and_gate_h_u_cla32_and4061_y0(h_u_cla32_and4060_y0, h_u_cla32_and4059_y0, h_u_cla32_and4061_y0);
  and_gate and_gate_h_u_cla32_and4062_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4062_y0);
  and_gate and_gate_h_u_cla32_and4063_y0(h_u_cla32_and4062_y0, h_u_cla32_and4061_y0, h_u_cla32_and4063_y0);
  and_gate and_gate_h_u_cla32_and4064_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4064_y0);
  and_gate and_gate_h_u_cla32_and4065_y0(h_u_cla32_and4064_y0, h_u_cla32_and4063_y0, h_u_cla32_and4065_y0);
  and_gate and_gate_h_u_cla32_and4066_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4066_y0);
  and_gate and_gate_h_u_cla32_and4067_y0(h_u_cla32_and4066_y0, h_u_cla32_and4065_y0, h_u_cla32_and4067_y0);
  and_gate and_gate_h_u_cla32_and4068_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4068_y0);
  and_gate and_gate_h_u_cla32_and4069_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4069_y0);
  and_gate and_gate_h_u_cla32_and4070_y0(h_u_cla32_and4069_y0, h_u_cla32_and4068_y0, h_u_cla32_and4070_y0);
  and_gate and_gate_h_u_cla32_and4071_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4071_y0);
  and_gate and_gate_h_u_cla32_and4072_y0(h_u_cla32_and4071_y0, h_u_cla32_and4070_y0, h_u_cla32_and4072_y0);
  and_gate and_gate_h_u_cla32_and4073_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4073_y0);
  and_gate and_gate_h_u_cla32_and4074_y0(h_u_cla32_and4073_y0, h_u_cla32_and4072_y0, h_u_cla32_and4074_y0);
  and_gate and_gate_h_u_cla32_and4075_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4075_y0);
  and_gate and_gate_h_u_cla32_and4076_y0(h_u_cla32_and4075_y0, h_u_cla32_and4074_y0, h_u_cla32_and4076_y0);
  and_gate and_gate_h_u_cla32_and4077_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4077_y0);
  and_gate and_gate_h_u_cla32_and4078_y0(h_u_cla32_and4077_y0, h_u_cla32_and4076_y0, h_u_cla32_and4078_y0);
  and_gate and_gate_h_u_cla32_and4079_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4079_y0);
  and_gate and_gate_h_u_cla32_and4080_y0(h_u_cla32_and4079_y0, h_u_cla32_and4078_y0, h_u_cla32_and4080_y0);
  and_gate and_gate_h_u_cla32_and4081_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4081_y0);
  and_gate and_gate_h_u_cla32_and4082_y0(h_u_cla32_and4081_y0, h_u_cla32_and4080_y0, h_u_cla32_and4082_y0);
  and_gate and_gate_h_u_cla32_and4083_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4083_y0);
  and_gate and_gate_h_u_cla32_and4084_y0(h_u_cla32_and4083_y0, h_u_cla32_and4082_y0, h_u_cla32_and4084_y0);
  and_gate and_gate_h_u_cla32_and4085_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4085_y0);
  and_gate and_gate_h_u_cla32_and4086_y0(h_u_cla32_and4085_y0, h_u_cla32_and4084_y0, h_u_cla32_and4086_y0);
  and_gate and_gate_h_u_cla32_and4087_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4087_y0);
  and_gate and_gate_h_u_cla32_and4088_y0(h_u_cla32_and4087_y0, h_u_cla32_and4086_y0, h_u_cla32_and4088_y0);
  and_gate and_gate_h_u_cla32_and4089_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4089_y0);
  and_gate and_gate_h_u_cla32_and4090_y0(h_u_cla32_and4089_y0, h_u_cla32_and4088_y0, h_u_cla32_and4090_y0);
  and_gate and_gate_h_u_cla32_and4091_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4091_y0);
  and_gate and_gate_h_u_cla32_and4092_y0(h_u_cla32_and4091_y0, h_u_cla32_and4090_y0, h_u_cla32_and4092_y0);
  and_gate and_gate_h_u_cla32_and4093_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4093_y0);
  and_gate and_gate_h_u_cla32_and4094_y0(h_u_cla32_and4093_y0, h_u_cla32_and4092_y0, h_u_cla32_and4094_y0);
  and_gate and_gate_h_u_cla32_and4095_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4095_y0);
  and_gate and_gate_h_u_cla32_and4096_y0(h_u_cla32_and4095_y0, h_u_cla32_and4094_y0, h_u_cla32_and4096_y0);
  and_gate and_gate_h_u_cla32_and4097_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4097_y0);
  and_gate and_gate_h_u_cla32_and4098_y0(h_u_cla32_and4097_y0, h_u_cla32_and4096_y0, h_u_cla32_and4098_y0);
  and_gate and_gate_h_u_cla32_and4099_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4099_y0);
  and_gate and_gate_h_u_cla32_and4100_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4100_y0);
  and_gate and_gate_h_u_cla32_and4101_y0(h_u_cla32_and4100_y0, h_u_cla32_and4099_y0, h_u_cla32_and4101_y0);
  and_gate and_gate_h_u_cla32_and4102_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4102_y0);
  and_gate and_gate_h_u_cla32_and4103_y0(h_u_cla32_and4102_y0, h_u_cla32_and4101_y0, h_u_cla32_and4103_y0);
  and_gate and_gate_h_u_cla32_and4104_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4104_y0);
  and_gate and_gate_h_u_cla32_and4105_y0(h_u_cla32_and4104_y0, h_u_cla32_and4103_y0, h_u_cla32_and4105_y0);
  and_gate and_gate_h_u_cla32_and4106_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4106_y0);
  and_gate and_gate_h_u_cla32_and4107_y0(h_u_cla32_and4106_y0, h_u_cla32_and4105_y0, h_u_cla32_and4107_y0);
  and_gate and_gate_h_u_cla32_and4108_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4108_y0);
  and_gate and_gate_h_u_cla32_and4109_y0(h_u_cla32_and4108_y0, h_u_cla32_and4107_y0, h_u_cla32_and4109_y0);
  and_gate and_gate_h_u_cla32_and4110_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4110_y0);
  and_gate and_gate_h_u_cla32_and4111_y0(h_u_cla32_and4110_y0, h_u_cla32_and4109_y0, h_u_cla32_and4111_y0);
  and_gate and_gate_h_u_cla32_and4112_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4112_y0);
  and_gate and_gate_h_u_cla32_and4113_y0(h_u_cla32_and4112_y0, h_u_cla32_and4111_y0, h_u_cla32_and4113_y0);
  and_gate and_gate_h_u_cla32_and4114_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4114_y0);
  and_gate and_gate_h_u_cla32_and4115_y0(h_u_cla32_and4114_y0, h_u_cla32_and4113_y0, h_u_cla32_and4115_y0);
  and_gate and_gate_h_u_cla32_and4116_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4116_y0);
  and_gate and_gate_h_u_cla32_and4117_y0(h_u_cla32_and4116_y0, h_u_cla32_and4115_y0, h_u_cla32_and4117_y0);
  and_gate and_gate_h_u_cla32_and4118_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4118_y0);
  and_gate and_gate_h_u_cla32_and4119_y0(h_u_cla32_and4118_y0, h_u_cla32_and4117_y0, h_u_cla32_and4119_y0);
  and_gate and_gate_h_u_cla32_and4120_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4120_y0);
  and_gate and_gate_h_u_cla32_and4121_y0(h_u_cla32_and4120_y0, h_u_cla32_and4119_y0, h_u_cla32_and4121_y0);
  and_gate and_gate_h_u_cla32_and4122_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4122_y0);
  and_gate and_gate_h_u_cla32_and4123_y0(h_u_cla32_and4122_y0, h_u_cla32_and4121_y0, h_u_cla32_and4123_y0);
  and_gate and_gate_h_u_cla32_and4124_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4124_y0);
  and_gate and_gate_h_u_cla32_and4125_y0(h_u_cla32_and4124_y0, h_u_cla32_and4123_y0, h_u_cla32_and4125_y0);
  and_gate and_gate_h_u_cla32_and4126_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4126_y0);
  and_gate and_gate_h_u_cla32_and4127_y0(h_u_cla32_and4126_y0, h_u_cla32_and4125_y0, h_u_cla32_and4127_y0);
  and_gate and_gate_h_u_cla32_and4128_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4128_y0);
  and_gate and_gate_h_u_cla32_and4129_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4129_y0);
  and_gate and_gate_h_u_cla32_and4130_y0(h_u_cla32_and4129_y0, h_u_cla32_and4128_y0, h_u_cla32_and4130_y0);
  and_gate and_gate_h_u_cla32_and4131_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4131_y0);
  and_gate and_gate_h_u_cla32_and4132_y0(h_u_cla32_and4131_y0, h_u_cla32_and4130_y0, h_u_cla32_and4132_y0);
  and_gate and_gate_h_u_cla32_and4133_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4133_y0);
  and_gate and_gate_h_u_cla32_and4134_y0(h_u_cla32_and4133_y0, h_u_cla32_and4132_y0, h_u_cla32_and4134_y0);
  and_gate and_gate_h_u_cla32_and4135_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4135_y0);
  and_gate and_gate_h_u_cla32_and4136_y0(h_u_cla32_and4135_y0, h_u_cla32_and4134_y0, h_u_cla32_and4136_y0);
  and_gate and_gate_h_u_cla32_and4137_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4137_y0);
  and_gate and_gate_h_u_cla32_and4138_y0(h_u_cla32_and4137_y0, h_u_cla32_and4136_y0, h_u_cla32_and4138_y0);
  and_gate and_gate_h_u_cla32_and4139_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4139_y0);
  and_gate and_gate_h_u_cla32_and4140_y0(h_u_cla32_and4139_y0, h_u_cla32_and4138_y0, h_u_cla32_and4140_y0);
  and_gate and_gate_h_u_cla32_and4141_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4141_y0);
  and_gate and_gate_h_u_cla32_and4142_y0(h_u_cla32_and4141_y0, h_u_cla32_and4140_y0, h_u_cla32_and4142_y0);
  and_gate and_gate_h_u_cla32_and4143_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4143_y0);
  and_gate and_gate_h_u_cla32_and4144_y0(h_u_cla32_and4143_y0, h_u_cla32_and4142_y0, h_u_cla32_and4144_y0);
  and_gate and_gate_h_u_cla32_and4145_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4145_y0);
  and_gate and_gate_h_u_cla32_and4146_y0(h_u_cla32_and4145_y0, h_u_cla32_and4144_y0, h_u_cla32_and4146_y0);
  and_gate and_gate_h_u_cla32_and4147_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4147_y0);
  and_gate and_gate_h_u_cla32_and4148_y0(h_u_cla32_and4147_y0, h_u_cla32_and4146_y0, h_u_cla32_and4148_y0);
  and_gate and_gate_h_u_cla32_and4149_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4149_y0);
  and_gate and_gate_h_u_cla32_and4150_y0(h_u_cla32_and4149_y0, h_u_cla32_and4148_y0, h_u_cla32_and4150_y0);
  and_gate and_gate_h_u_cla32_and4151_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4151_y0);
  and_gate and_gate_h_u_cla32_and4152_y0(h_u_cla32_and4151_y0, h_u_cla32_and4150_y0, h_u_cla32_and4152_y0);
  and_gate and_gate_h_u_cla32_and4153_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4153_y0);
  and_gate and_gate_h_u_cla32_and4154_y0(h_u_cla32_and4153_y0, h_u_cla32_and4152_y0, h_u_cla32_and4154_y0);
  and_gate and_gate_h_u_cla32_and4155_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4155_y0);
  and_gate and_gate_h_u_cla32_and4156_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4156_y0);
  and_gate and_gate_h_u_cla32_and4157_y0(h_u_cla32_and4156_y0, h_u_cla32_and4155_y0, h_u_cla32_and4157_y0);
  and_gate and_gate_h_u_cla32_and4158_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4158_y0);
  and_gate and_gate_h_u_cla32_and4159_y0(h_u_cla32_and4158_y0, h_u_cla32_and4157_y0, h_u_cla32_and4159_y0);
  and_gate and_gate_h_u_cla32_and4160_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4160_y0);
  and_gate and_gate_h_u_cla32_and4161_y0(h_u_cla32_and4160_y0, h_u_cla32_and4159_y0, h_u_cla32_and4161_y0);
  and_gate and_gate_h_u_cla32_and4162_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4162_y0);
  and_gate and_gate_h_u_cla32_and4163_y0(h_u_cla32_and4162_y0, h_u_cla32_and4161_y0, h_u_cla32_and4163_y0);
  and_gate and_gate_h_u_cla32_and4164_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4164_y0);
  and_gate and_gate_h_u_cla32_and4165_y0(h_u_cla32_and4164_y0, h_u_cla32_and4163_y0, h_u_cla32_and4165_y0);
  and_gate and_gate_h_u_cla32_and4166_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4166_y0);
  and_gate and_gate_h_u_cla32_and4167_y0(h_u_cla32_and4166_y0, h_u_cla32_and4165_y0, h_u_cla32_and4167_y0);
  and_gate and_gate_h_u_cla32_and4168_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4168_y0);
  and_gate and_gate_h_u_cla32_and4169_y0(h_u_cla32_and4168_y0, h_u_cla32_and4167_y0, h_u_cla32_and4169_y0);
  and_gate and_gate_h_u_cla32_and4170_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4170_y0);
  and_gate and_gate_h_u_cla32_and4171_y0(h_u_cla32_and4170_y0, h_u_cla32_and4169_y0, h_u_cla32_and4171_y0);
  and_gate and_gate_h_u_cla32_and4172_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4172_y0);
  and_gate and_gate_h_u_cla32_and4173_y0(h_u_cla32_and4172_y0, h_u_cla32_and4171_y0, h_u_cla32_and4173_y0);
  and_gate and_gate_h_u_cla32_and4174_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4174_y0);
  and_gate and_gate_h_u_cla32_and4175_y0(h_u_cla32_and4174_y0, h_u_cla32_and4173_y0, h_u_cla32_and4175_y0);
  and_gate and_gate_h_u_cla32_and4176_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4176_y0);
  and_gate and_gate_h_u_cla32_and4177_y0(h_u_cla32_and4176_y0, h_u_cla32_and4175_y0, h_u_cla32_and4177_y0);
  and_gate and_gate_h_u_cla32_and4178_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4178_y0);
  and_gate and_gate_h_u_cla32_and4179_y0(h_u_cla32_and4178_y0, h_u_cla32_and4177_y0, h_u_cla32_and4179_y0);
  and_gate and_gate_h_u_cla32_and4180_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4180_y0);
  and_gate and_gate_h_u_cla32_and4181_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4181_y0);
  and_gate and_gate_h_u_cla32_and4182_y0(h_u_cla32_and4181_y0, h_u_cla32_and4180_y0, h_u_cla32_and4182_y0);
  and_gate and_gate_h_u_cla32_and4183_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4183_y0);
  and_gate and_gate_h_u_cla32_and4184_y0(h_u_cla32_and4183_y0, h_u_cla32_and4182_y0, h_u_cla32_and4184_y0);
  and_gate and_gate_h_u_cla32_and4185_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4185_y0);
  and_gate and_gate_h_u_cla32_and4186_y0(h_u_cla32_and4185_y0, h_u_cla32_and4184_y0, h_u_cla32_and4186_y0);
  and_gate and_gate_h_u_cla32_and4187_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4187_y0);
  and_gate and_gate_h_u_cla32_and4188_y0(h_u_cla32_and4187_y0, h_u_cla32_and4186_y0, h_u_cla32_and4188_y0);
  and_gate and_gate_h_u_cla32_and4189_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4189_y0);
  and_gate and_gate_h_u_cla32_and4190_y0(h_u_cla32_and4189_y0, h_u_cla32_and4188_y0, h_u_cla32_and4190_y0);
  and_gate and_gate_h_u_cla32_and4191_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4191_y0);
  and_gate and_gate_h_u_cla32_and4192_y0(h_u_cla32_and4191_y0, h_u_cla32_and4190_y0, h_u_cla32_and4192_y0);
  and_gate and_gate_h_u_cla32_and4193_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4193_y0);
  and_gate and_gate_h_u_cla32_and4194_y0(h_u_cla32_and4193_y0, h_u_cla32_and4192_y0, h_u_cla32_and4194_y0);
  and_gate and_gate_h_u_cla32_and4195_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4195_y0);
  and_gate and_gate_h_u_cla32_and4196_y0(h_u_cla32_and4195_y0, h_u_cla32_and4194_y0, h_u_cla32_and4196_y0);
  and_gate and_gate_h_u_cla32_and4197_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4197_y0);
  and_gate and_gate_h_u_cla32_and4198_y0(h_u_cla32_and4197_y0, h_u_cla32_and4196_y0, h_u_cla32_and4198_y0);
  and_gate and_gate_h_u_cla32_and4199_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4199_y0);
  and_gate and_gate_h_u_cla32_and4200_y0(h_u_cla32_and4199_y0, h_u_cla32_and4198_y0, h_u_cla32_and4200_y0);
  and_gate and_gate_h_u_cla32_and4201_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4201_y0);
  and_gate and_gate_h_u_cla32_and4202_y0(h_u_cla32_and4201_y0, h_u_cla32_and4200_y0, h_u_cla32_and4202_y0);
  and_gate and_gate_h_u_cla32_and4203_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4203_y0);
  and_gate and_gate_h_u_cla32_and4204_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4204_y0);
  and_gate and_gate_h_u_cla32_and4205_y0(h_u_cla32_and4204_y0, h_u_cla32_and4203_y0, h_u_cla32_and4205_y0);
  and_gate and_gate_h_u_cla32_and4206_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4206_y0);
  and_gate and_gate_h_u_cla32_and4207_y0(h_u_cla32_and4206_y0, h_u_cla32_and4205_y0, h_u_cla32_and4207_y0);
  and_gate and_gate_h_u_cla32_and4208_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4208_y0);
  and_gate and_gate_h_u_cla32_and4209_y0(h_u_cla32_and4208_y0, h_u_cla32_and4207_y0, h_u_cla32_and4209_y0);
  and_gate and_gate_h_u_cla32_and4210_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4210_y0);
  and_gate and_gate_h_u_cla32_and4211_y0(h_u_cla32_and4210_y0, h_u_cla32_and4209_y0, h_u_cla32_and4211_y0);
  and_gate and_gate_h_u_cla32_and4212_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4212_y0);
  and_gate and_gate_h_u_cla32_and4213_y0(h_u_cla32_and4212_y0, h_u_cla32_and4211_y0, h_u_cla32_and4213_y0);
  and_gate and_gate_h_u_cla32_and4214_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4214_y0);
  and_gate and_gate_h_u_cla32_and4215_y0(h_u_cla32_and4214_y0, h_u_cla32_and4213_y0, h_u_cla32_and4215_y0);
  and_gate and_gate_h_u_cla32_and4216_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4216_y0);
  and_gate and_gate_h_u_cla32_and4217_y0(h_u_cla32_and4216_y0, h_u_cla32_and4215_y0, h_u_cla32_and4217_y0);
  and_gate and_gate_h_u_cla32_and4218_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4218_y0);
  and_gate and_gate_h_u_cla32_and4219_y0(h_u_cla32_and4218_y0, h_u_cla32_and4217_y0, h_u_cla32_and4219_y0);
  and_gate and_gate_h_u_cla32_and4220_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4220_y0);
  and_gate and_gate_h_u_cla32_and4221_y0(h_u_cla32_and4220_y0, h_u_cla32_and4219_y0, h_u_cla32_and4221_y0);
  and_gate and_gate_h_u_cla32_and4222_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4222_y0);
  and_gate and_gate_h_u_cla32_and4223_y0(h_u_cla32_and4222_y0, h_u_cla32_and4221_y0, h_u_cla32_and4223_y0);
  and_gate and_gate_h_u_cla32_and4224_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4224_y0);
  and_gate and_gate_h_u_cla32_and4225_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4225_y0);
  and_gate and_gate_h_u_cla32_and4226_y0(h_u_cla32_and4225_y0, h_u_cla32_and4224_y0, h_u_cla32_and4226_y0);
  and_gate and_gate_h_u_cla32_and4227_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4227_y0);
  and_gate and_gate_h_u_cla32_and4228_y0(h_u_cla32_and4227_y0, h_u_cla32_and4226_y0, h_u_cla32_and4228_y0);
  and_gate and_gate_h_u_cla32_and4229_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4229_y0);
  and_gate and_gate_h_u_cla32_and4230_y0(h_u_cla32_and4229_y0, h_u_cla32_and4228_y0, h_u_cla32_and4230_y0);
  and_gate and_gate_h_u_cla32_and4231_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4231_y0);
  and_gate and_gate_h_u_cla32_and4232_y0(h_u_cla32_and4231_y0, h_u_cla32_and4230_y0, h_u_cla32_and4232_y0);
  and_gate and_gate_h_u_cla32_and4233_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4233_y0);
  and_gate and_gate_h_u_cla32_and4234_y0(h_u_cla32_and4233_y0, h_u_cla32_and4232_y0, h_u_cla32_and4234_y0);
  and_gate and_gate_h_u_cla32_and4235_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4235_y0);
  and_gate and_gate_h_u_cla32_and4236_y0(h_u_cla32_and4235_y0, h_u_cla32_and4234_y0, h_u_cla32_and4236_y0);
  and_gate and_gate_h_u_cla32_and4237_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4237_y0);
  and_gate and_gate_h_u_cla32_and4238_y0(h_u_cla32_and4237_y0, h_u_cla32_and4236_y0, h_u_cla32_and4238_y0);
  and_gate and_gate_h_u_cla32_and4239_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4239_y0);
  and_gate and_gate_h_u_cla32_and4240_y0(h_u_cla32_and4239_y0, h_u_cla32_and4238_y0, h_u_cla32_and4240_y0);
  and_gate and_gate_h_u_cla32_and4241_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4241_y0);
  and_gate and_gate_h_u_cla32_and4242_y0(h_u_cla32_and4241_y0, h_u_cla32_and4240_y0, h_u_cla32_and4242_y0);
  and_gate and_gate_h_u_cla32_and4243_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4243_y0);
  and_gate and_gate_h_u_cla32_and4244_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4244_y0);
  and_gate and_gate_h_u_cla32_and4245_y0(h_u_cla32_and4244_y0, h_u_cla32_and4243_y0, h_u_cla32_and4245_y0);
  and_gate and_gate_h_u_cla32_and4246_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4246_y0);
  and_gate and_gate_h_u_cla32_and4247_y0(h_u_cla32_and4246_y0, h_u_cla32_and4245_y0, h_u_cla32_and4247_y0);
  and_gate and_gate_h_u_cla32_and4248_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4248_y0);
  and_gate and_gate_h_u_cla32_and4249_y0(h_u_cla32_and4248_y0, h_u_cla32_and4247_y0, h_u_cla32_and4249_y0);
  and_gate and_gate_h_u_cla32_and4250_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4250_y0);
  and_gate and_gate_h_u_cla32_and4251_y0(h_u_cla32_and4250_y0, h_u_cla32_and4249_y0, h_u_cla32_and4251_y0);
  and_gate and_gate_h_u_cla32_and4252_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4252_y0);
  and_gate and_gate_h_u_cla32_and4253_y0(h_u_cla32_and4252_y0, h_u_cla32_and4251_y0, h_u_cla32_and4253_y0);
  and_gate and_gate_h_u_cla32_and4254_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4254_y0);
  and_gate and_gate_h_u_cla32_and4255_y0(h_u_cla32_and4254_y0, h_u_cla32_and4253_y0, h_u_cla32_and4255_y0);
  and_gate and_gate_h_u_cla32_and4256_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4256_y0);
  and_gate and_gate_h_u_cla32_and4257_y0(h_u_cla32_and4256_y0, h_u_cla32_and4255_y0, h_u_cla32_and4257_y0);
  and_gate and_gate_h_u_cla32_and4258_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4258_y0);
  and_gate and_gate_h_u_cla32_and4259_y0(h_u_cla32_and4258_y0, h_u_cla32_and4257_y0, h_u_cla32_and4259_y0);
  and_gate and_gate_h_u_cla32_and4260_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4260_y0);
  and_gate and_gate_h_u_cla32_and4261_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4261_y0);
  and_gate and_gate_h_u_cla32_and4262_y0(h_u_cla32_and4261_y0, h_u_cla32_and4260_y0, h_u_cla32_and4262_y0);
  and_gate and_gate_h_u_cla32_and4263_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4263_y0);
  and_gate and_gate_h_u_cla32_and4264_y0(h_u_cla32_and4263_y0, h_u_cla32_and4262_y0, h_u_cla32_and4264_y0);
  and_gate and_gate_h_u_cla32_and4265_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4265_y0);
  and_gate and_gate_h_u_cla32_and4266_y0(h_u_cla32_and4265_y0, h_u_cla32_and4264_y0, h_u_cla32_and4266_y0);
  and_gate and_gate_h_u_cla32_and4267_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4267_y0);
  and_gate and_gate_h_u_cla32_and4268_y0(h_u_cla32_and4267_y0, h_u_cla32_and4266_y0, h_u_cla32_and4268_y0);
  and_gate and_gate_h_u_cla32_and4269_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4269_y0);
  and_gate and_gate_h_u_cla32_and4270_y0(h_u_cla32_and4269_y0, h_u_cla32_and4268_y0, h_u_cla32_and4270_y0);
  and_gate and_gate_h_u_cla32_and4271_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4271_y0);
  and_gate and_gate_h_u_cla32_and4272_y0(h_u_cla32_and4271_y0, h_u_cla32_and4270_y0, h_u_cla32_and4272_y0);
  and_gate and_gate_h_u_cla32_and4273_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4273_y0);
  and_gate and_gate_h_u_cla32_and4274_y0(h_u_cla32_and4273_y0, h_u_cla32_and4272_y0, h_u_cla32_and4274_y0);
  and_gate and_gate_h_u_cla32_and4275_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4275_y0);
  and_gate and_gate_h_u_cla32_and4276_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4276_y0);
  and_gate and_gate_h_u_cla32_and4277_y0(h_u_cla32_and4276_y0, h_u_cla32_and4275_y0, h_u_cla32_and4277_y0);
  and_gate and_gate_h_u_cla32_and4278_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4278_y0);
  and_gate and_gate_h_u_cla32_and4279_y0(h_u_cla32_and4278_y0, h_u_cla32_and4277_y0, h_u_cla32_and4279_y0);
  and_gate and_gate_h_u_cla32_and4280_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4280_y0);
  and_gate and_gate_h_u_cla32_and4281_y0(h_u_cla32_and4280_y0, h_u_cla32_and4279_y0, h_u_cla32_and4281_y0);
  and_gate and_gate_h_u_cla32_and4282_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4282_y0);
  and_gate and_gate_h_u_cla32_and4283_y0(h_u_cla32_and4282_y0, h_u_cla32_and4281_y0, h_u_cla32_and4283_y0);
  and_gate and_gate_h_u_cla32_and4284_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4284_y0);
  and_gate and_gate_h_u_cla32_and4285_y0(h_u_cla32_and4284_y0, h_u_cla32_and4283_y0, h_u_cla32_and4285_y0);
  and_gate and_gate_h_u_cla32_and4286_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4286_y0);
  and_gate and_gate_h_u_cla32_and4287_y0(h_u_cla32_and4286_y0, h_u_cla32_and4285_y0, h_u_cla32_and4287_y0);
  and_gate and_gate_h_u_cla32_and4288_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4288_y0);
  and_gate and_gate_h_u_cla32_and4289_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4289_y0);
  and_gate and_gate_h_u_cla32_and4290_y0(h_u_cla32_and4289_y0, h_u_cla32_and4288_y0, h_u_cla32_and4290_y0);
  and_gate and_gate_h_u_cla32_and4291_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4291_y0);
  and_gate and_gate_h_u_cla32_and4292_y0(h_u_cla32_and4291_y0, h_u_cla32_and4290_y0, h_u_cla32_and4292_y0);
  and_gate and_gate_h_u_cla32_and4293_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4293_y0);
  and_gate and_gate_h_u_cla32_and4294_y0(h_u_cla32_and4293_y0, h_u_cla32_and4292_y0, h_u_cla32_and4294_y0);
  and_gate and_gate_h_u_cla32_and4295_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4295_y0);
  and_gate and_gate_h_u_cla32_and4296_y0(h_u_cla32_and4295_y0, h_u_cla32_and4294_y0, h_u_cla32_and4296_y0);
  and_gate and_gate_h_u_cla32_and4297_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4297_y0);
  and_gate and_gate_h_u_cla32_and4298_y0(h_u_cla32_and4297_y0, h_u_cla32_and4296_y0, h_u_cla32_and4298_y0);
  and_gate and_gate_h_u_cla32_and4299_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4299_y0);
  and_gate and_gate_h_u_cla32_and4300_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4300_y0);
  and_gate and_gate_h_u_cla32_and4301_y0(h_u_cla32_and4300_y0, h_u_cla32_and4299_y0, h_u_cla32_and4301_y0);
  and_gate and_gate_h_u_cla32_and4302_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4302_y0);
  and_gate and_gate_h_u_cla32_and4303_y0(h_u_cla32_and4302_y0, h_u_cla32_and4301_y0, h_u_cla32_and4303_y0);
  and_gate and_gate_h_u_cla32_and4304_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4304_y0);
  and_gate and_gate_h_u_cla32_and4305_y0(h_u_cla32_and4304_y0, h_u_cla32_and4303_y0, h_u_cla32_and4305_y0);
  and_gate and_gate_h_u_cla32_and4306_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4306_y0);
  and_gate and_gate_h_u_cla32_and4307_y0(h_u_cla32_and4306_y0, h_u_cla32_and4305_y0, h_u_cla32_and4307_y0);
  and_gate and_gate_h_u_cla32_and4308_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4308_y0);
  and_gate and_gate_h_u_cla32_and4309_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4309_y0);
  and_gate and_gate_h_u_cla32_and4310_y0(h_u_cla32_and4309_y0, h_u_cla32_and4308_y0, h_u_cla32_and4310_y0);
  and_gate and_gate_h_u_cla32_and4311_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4311_y0);
  and_gate and_gate_h_u_cla32_and4312_y0(h_u_cla32_and4311_y0, h_u_cla32_and4310_y0, h_u_cla32_and4312_y0);
  and_gate and_gate_h_u_cla32_and4313_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4313_y0);
  and_gate and_gate_h_u_cla32_and4314_y0(h_u_cla32_and4313_y0, h_u_cla32_and4312_y0, h_u_cla32_and4314_y0);
  and_gate and_gate_h_u_cla32_and4315_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4315_y0);
  and_gate and_gate_h_u_cla32_and4316_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4316_y0);
  and_gate and_gate_h_u_cla32_and4317_y0(h_u_cla32_and4316_y0, h_u_cla32_and4315_y0, h_u_cla32_and4317_y0);
  and_gate and_gate_h_u_cla32_and4318_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4318_y0);
  and_gate and_gate_h_u_cla32_and4319_y0(h_u_cla32_and4318_y0, h_u_cla32_and4317_y0, h_u_cla32_and4319_y0);
  and_gate and_gate_h_u_cla32_and4320_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and4320_y0);
  and_gate and_gate_h_u_cla32_and4321_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and4321_y0);
  and_gate and_gate_h_u_cla32_and4322_y0(h_u_cla32_and4321_y0, h_u_cla32_and4320_y0, h_u_cla32_and4322_y0);
  and_gate and_gate_h_u_cla32_and4323_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and4323_y0);
  or_gate or_gate_h_u_cla32_or253_y0(h_u_cla32_and4323_y0, h_u_cla32_and3839_y0, h_u_cla32_or253_y0);
  or_gate or_gate_h_u_cla32_or254_y0(h_u_cla32_or253_y0, h_u_cla32_and3882_y0, h_u_cla32_or254_y0);
  or_gate or_gate_h_u_cla32_or255_y0(h_u_cla32_or254_y0, h_u_cla32_and3923_y0, h_u_cla32_or255_y0);
  or_gate or_gate_h_u_cla32_or256_y0(h_u_cla32_or255_y0, h_u_cla32_and3962_y0, h_u_cla32_or256_y0);
  or_gate or_gate_h_u_cla32_or257_y0(h_u_cla32_or256_y0, h_u_cla32_and3999_y0, h_u_cla32_or257_y0);
  or_gate or_gate_h_u_cla32_or258_y0(h_u_cla32_or257_y0, h_u_cla32_and4034_y0, h_u_cla32_or258_y0);
  or_gate or_gate_h_u_cla32_or259_y0(h_u_cla32_or258_y0, h_u_cla32_and4067_y0, h_u_cla32_or259_y0);
  or_gate or_gate_h_u_cla32_or260_y0(h_u_cla32_or259_y0, h_u_cla32_and4098_y0, h_u_cla32_or260_y0);
  or_gate or_gate_h_u_cla32_or261_y0(h_u_cla32_or260_y0, h_u_cla32_and4127_y0, h_u_cla32_or261_y0);
  or_gate or_gate_h_u_cla32_or262_y0(h_u_cla32_or261_y0, h_u_cla32_and4154_y0, h_u_cla32_or262_y0);
  or_gate or_gate_h_u_cla32_or263_y0(h_u_cla32_or262_y0, h_u_cla32_and4179_y0, h_u_cla32_or263_y0);
  or_gate or_gate_h_u_cla32_or264_y0(h_u_cla32_or263_y0, h_u_cla32_and4202_y0, h_u_cla32_or264_y0);
  or_gate or_gate_h_u_cla32_or265_y0(h_u_cla32_or264_y0, h_u_cla32_and4223_y0, h_u_cla32_or265_y0);
  or_gate or_gate_h_u_cla32_or266_y0(h_u_cla32_or265_y0, h_u_cla32_and4242_y0, h_u_cla32_or266_y0);
  or_gate or_gate_h_u_cla32_or267_y0(h_u_cla32_or266_y0, h_u_cla32_and4259_y0, h_u_cla32_or267_y0);
  or_gate or_gate_h_u_cla32_or268_y0(h_u_cla32_or267_y0, h_u_cla32_and4274_y0, h_u_cla32_or268_y0);
  or_gate or_gate_h_u_cla32_or269_y0(h_u_cla32_or268_y0, h_u_cla32_and4287_y0, h_u_cla32_or269_y0);
  or_gate or_gate_h_u_cla32_or270_y0(h_u_cla32_or269_y0, h_u_cla32_and4298_y0, h_u_cla32_or270_y0);
  or_gate or_gate_h_u_cla32_or271_y0(h_u_cla32_or270_y0, h_u_cla32_and4307_y0, h_u_cla32_or271_y0);
  or_gate or_gate_h_u_cla32_or272_y0(h_u_cla32_or271_y0, h_u_cla32_and4314_y0, h_u_cla32_or272_y0);
  or_gate or_gate_h_u_cla32_or273_y0(h_u_cla32_or272_y0, h_u_cla32_and4319_y0, h_u_cla32_or273_y0);
  or_gate or_gate_h_u_cla32_or274_y0(h_u_cla32_or273_y0, h_u_cla32_and4322_y0, h_u_cla32_or274_y0);
  or_gate or_gate_h_u_cla32_or275_y0(h_u_cla32_pg_logic22_y1, h_u_cla32_or274_y0, h_u_cla32_or275_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic23_y0(a_23, b_23, h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_pg_logic23_y2);
  xor_gate xor_gate_h_u_cla32_xor23_y0(h_u_cla32_pg_logic23_y2, h_u_cla32_or275_y0, h_u_cla32_xor23_y0);
  and_gate and_gate_h_u_cla32_and4324_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and4324_y0);
  and_gate and_gate_h_u_cla32_and4325_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and4325_y0);
  and_gate and_gate_h_u_cla32_and4326_y0(h_u_cla32_and4325_y0, h_u_cla32_and4324_y0, h_u_cla32_and4326_y0);
  and_gate and_gate_h_u_cla32_and4327_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and4327_y0);
  and_gate and_gate_h_u_cla32_and4328_y0(h_u_cla32_and4327_y0, h_u_cla32_and4326_y0, h_u_cla32_and4328_y0);
  and_gate and_gate_h_u_cla32_and4329_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and4329_y0);
  and_gate and_gate_h_u_cla32_and4330_y0(h_u_cla32_and4329_y0, h_u_cla32_and4328_y0, h_u_cla32_and4330_y0);
  and_gate and_gate_h_u_cla32_and4331_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and4331_y0);
  and_gate and_gate_h_u_cla32_and4332_y0(h_u_cla32_and4331_y0, h_u_cla32_and4330_y0, h_u_cla32_and4332_y0);
  and_gate and_gate_h_u_cla32_and4333_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and4333_y0);
  and_gate and_gate_h_u_cla32_and4334_y0(h_u_cla32_and4333_y0, h_u_cla32_and4332_y0, h_u_cla32_and4334_y0);
  and_gate and_gate_h_u_cla32_and4335_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and4335_y0);
  and_gate and_gate_h_u_cla32_and4336_y0(h_u_cla32_and4335_y0, h_u_cla32_and4334_y0, h_u_cla32_and4336_y0);
  and_gate and_gate_h_u_cla32_and4337_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and4337_y0);
  and_gate and_gate_h_u_cla32_and4338_y0(h_u_cla32_and4337_y0, h_u_cla32_and4336_y0, h_u_cla32_and4338_y0);
  and_gate and_gate_h_u_cla32_and4339_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and4339_y0);
  and_gate and_gate_h_u_cla32_and4340_y0(h_u_cla32_and4339_y0, h_u_cla32_and4338_y0, h_u_cla32_and4340_y0);
  and_gate and_gate_h_u_cla32_and4341_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and4341_y0);
  and_gate and_gate_h_u_cla32_and4342_y0(h_u_cla32_and4341_y0, h_u_cla32_and4340_y0, h_u_cla32_and4342_y0);
  and_gate and_gate_h_u_cla32_and4343_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and4343_y0);
  and_gate and_gate_h_u_cla32_and4344_y0(h_u_cla32_and4343_y0, h_u_cla32_and4342_y0, h_u_cla32_and4344_y0);
  and_gate and_gate_h_u_cla32_and4345_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and4345_y0);
  and_gate and_gate_h_u_cla32_and4346_y0(h_u_cla32_and4345_y0, h_u_cla32_and4344_y0, h_u_cla32_and4346_y0);
  and_gate and_gate_h_u_cla32_and4347_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and4347_y0);
  and_gate and_gate_h_u_cla32_and4348_y0(h_u_cla32_and4347_y0, h_u_cla32_and4346_y0, h_u_cla32_and4348_y0);
  and_gate and_gate_h_u_cla32_and4349_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and4349_y0);
  and_gate and_gate_h_u_cla32_and4350_y0(h_u_cla32_and4349_y0, h_u_cla32_and4348_y0, h_u_cla32_and4350_y0);
  and_gate and_gate_h_u_cla32_and4351_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and4351_y0);
  and_gate and_gate_h_u_cla32_and4352_y0(h_u_cla32_and4351_y0, h_u_cla32_and4350_y0, h_u_cla32_and4352_y0);
  and_gate and_gate_h_u_cla32_and4353_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and4353_y0);
  and_gate and_gate_h_u_cla32_and4354_y0(h_u_cla32_and4353_y0, h_u_cla32_and4352_y0, h_u_cla32_and4354_y0);
  and_gate and_gate_h_u_cla32_and4355_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and4355_y0);
  and_gate and_gate_h_u_cla32_and4356_y0(h_u_cla32_and4355_y0, h_u_cla32_and4354_y0, h_u_cla32_and4356_y0);
  and_gate and_gate_h_u_cla32_and4357_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and4357_y0);
  and_gate and_gate_h_u_cla32_and4358_y0(h_u_cla32_and4357_y0, h_u_cla32_and4356_y0, h_u_cla32_and4358_y0);
  and_gate and_gate_h_u_cla32_and4359_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and4359_y0);
  and_gate and_gate_h_u_cla32_and4360_y0(h_u_cla32_and4359_y0, h_u_cla32_and4358_y0, h_u_cla32_and4360_y0);
  and_gate and_gate_h_u_cla32_and4361_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and4361_y0);
  and_gate and_gate_h_u_cla32_and4362_y0(h_u_cla32_and4361_y0, h_u_cla32_and4360_y0, h_u_cla32_and4362_y0);
  and_gate and_gate_h_u_cla32_and4363_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and4363_y0);
  and_gate and_gate_h_u_cla32_and4364_y0(h_u_cla32_and4363_y0, h_u_cla32_and4362_y0, h_u_cla32_and4364_y0);
  and_gate and_gate_h_u_cla32_and4365_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and4365_y0);
  and_gate and_gate_h_u_cla32_and4366_y0(h_u_cla32_and4365_y0, h_u_cla32_and4364_y0, h_u_cla32_and4366_y0);
  and_gate and_gate_h_u_cla32_and4367_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and4367_y0);
  and_gate and_gate_h_u_cla32_and4368_y0(h_u_cla32_and4367_y0, h_u_cla32_and4366_y0, h_u_cla32_and4368_y0);
  and_gate and_gate_h_u_cla32_and4369_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and4369_y0);
  and_gate and_gate_h_u_cla32_and4370_y0(h_u_cla32_and4369_y0, h_u_cla32_and4368_y0, h_u_cla32_and4370_y0);
  and_gate and_gate_h_u_cla32_and4371_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4371_y0);
  and_gate and_gate_h_u_cla32_and4372_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4372_y0);
  and_gate and_gate_h_u_cla32_and4373_y0(h_u_cla32_and4372_y0, h_u_cla32_and4371_y0, h_u_cla32_and4373_y0);
  and_gate and_gate_h_u_cla32_and4374_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4374_y0);
  and_gate and_gate_h_u_cla32_and4375_y0(h_u_cla32_and4374_y0, h_u_cla32_and4373_y0, h_u_cla32_and4375_y0);
  and_gate and_gate_h_u_cla32_and4376_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4376_y0);
  and_gate and_gate_h_u_cla32_and4377_y0(h_u_cla32_and4376_y0, h_u_cla32_and4375_y0, h_u_cla32_and4377_y0);
  and_gate and_gate_h_u_cla32_and4378_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4378_y0);
  and_gate and_gate_h_u_cla32_and4379_y0(h_u_cla32_and4378_y0, h_u_cla32_and4377_y0, h_u_cla32_and4379_y0);
  and_gate and_gate_h_u_cla32_and4380_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4380_y0);
  and_gate and_gate_h_u_cla32_and4381_y0(h_u_cla32_and4380_y0, h_u_cla32_and4379_y0, h_u_cla32_and4381_y0);
  and_gate and_gate_h_u_cla32_and4382_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4382_y0);
  and_gate and_gate_h_u_cla32_and4383_y0(h_u_cla32_and4382_y0, h_u_cla32_and4381_y0, h_u_cla32_and4383_y0);
  and_gate and_gate_h_u_cla32_and4384_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4384_y0);
  and_gate and_gate_h_u_cla32_and4385_y0(h_u_cla32_and4384_y0, h_u_cla32_and4383_y0, h_u_cla32_and4385_y0);
  and_gate and_gate_h_u_cla32_and4386_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4386_y0);
  and_gate and_gate_h_u_cla32_and4387_y0(h_u_cla32_and4386_y0, h_u_cla32_and4385_y0, h_u_cla32_and4387_y0);
  and_gate and_gate_h_u_cla32_and4388_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4388_y0);
  and_gate and_gate_h_u_cla32_and4389_y0(h_u_cla32_and4388_y0, h_u_cla32_and4387_y0, h_u_cla32_and4389_y0);
  and_gate and_gate_h_u_cla32_and4390_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4390_y0);
  and_gate and_gate_h_u_cla32_and4391_y0(h_u_cla32_and4390_y0, h_u_cla32_and4389_y0, h_u_cla32_and4391_y0);
  and_gate and_gate_h_u_cla32_and4392_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4392_y0);
  and_gate and_gate_h_u_cla32_and4393_y0(h_u_cla32_and4392_y0, h_u_cla32_and4391_y0, h_u_cla32_and4393_y0);
  and_gate and_gate_h_u_cla32_and4394_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4394_y0);
  and_gate and_gate_h_u_cla32_and4395_y0(h_u_cla32_and4394_y0, h_u_cla32_and4393_y0, h_u_cla32_and4395_y0);
  and_gate and_gate_h_u_cla32_and4396_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4396_y0);
  and_gate and_gate_h_u_cla32_and4397_y0(h_u_cla32_and4396_y0, h_u_cla32_and4395_y0, h_u_cla32_and4397_y0);
  and_gate and_gate_h_u_cla32_and4398_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4398_y0);
  and_gate and_gate_h_u_cla32_and4399_y0(h_u_cla32_and4398_y0, h_u_cla32_and4397_y0, h_u_cla32_and4399_y0);
  and_gate and_gate_h_u_cla32_and4400_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4400_y0);
  and_gate and_gate_h_u_cla32_and4401_y0(h_u_cla32_and4400_y0, h_u_cla32_and4399_y0, h_u_cla32_and4401_y0);
  and_gate and_gate_h_u_cla32_and4402_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4402_y0);
  and_gate and_gate_h_u_cla32_and4403_y0(h_u_cla32_and4402_y0, h_u_cla32_and4401_y0, h_u_cla32_and4403_y0);
  and_gate and_gate_h_u_cla32_and4404_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4404_y0);
  and_gate and_gate_h_u_cla32_and4405_y0(h_u_cla32_and4404_y0, h_u_cla32_and4403_y0, h_u_cla32_and4405_y0);
  and_gate and_gate_h_u_cla32_and4406_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4406_y0);
  and_gate and_gate_h_u_cla32_and4407_y0(h_u_cla32_and4406_y0, h_u_cla32_and4405_y0, h_u_cla32_and4407_y0);
  and_gate and_gate_h_u_cla32_and4408_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4408_y0);
  and_gate and_gate_h_u_cla32_and4409_y0(h_u_cla32_and4408_y0, h_u_cla32_and4407_y0, h_u_cla32_and4409_y0);
  and_gate and_gate_h_u_cla32_and4410_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4410_y0);
  and_gate and_gate_h_u_cla32_and4411_y0(h_u_cla32_and4410_y0, h_u_cla32_and4409_y0, h_u_cla32_and4411_y0);
  and_gate and_gate_h_u_cla32_and4412_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4412_y0);
  and_gate and_gate_h_u_cla32_and4413_y0(h_u_cla32_and4412_y0, h_u_cla32_and4411_y0, h_u_cla32_and4413_y0);
  and_gate and_gate_h_u_cla32_and4414_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4414_y0);
  and_gate and_gate_h_u_cla32_and4415_y0(h_u_cla32_and4414_y0, h_u_cla32_and4413_y0, h_u_cla32_and4415_y0);
  and_gate and_gate_h_u_cla32_and4416_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4416_y0);
  and_gate and_gate_h_u_cla32_and4417_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4417_y0);
  and_gate and_gate_h_u_cla32_and4418_y0(h_u_cla32_and4417_y0, h_u_cla32_and4416_y0, h_u_cla32_and4418_y0);
  and_gate and_gate_h_u_cla32_and4419_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4419_y0);
  and_gate and_gate_h_u_cla32_and4420_y0(h_u_cla32_and4419_y0, h_u_cla32_and4418_y0, h_u_cla32_and4420_y0);
  and_gate and_gate_h_u_cla32_and4421_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4421_y0);
  and_gate and_gate_h_u_cla32_and4422_y0(h_u_cla32_and4421_y0, h_u_cla32_and4420_y0, h_u_cla32_and4422_y0);
  and_gate and_gate_h_u_cla32_and4423_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4423_y0);
  and_gate and_gate_h_u_cla32_and4424_y0(h_u_cla32_and4423_y0, h_u_cla32_and4422_y0, h_u_cla32_and4424_y0);
  and_gate and_gate_h_u_cla32_and4425_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4425_y0);
  and_gate and_gate_h_u_cla32_and4426_y0(h_u_cla32_and4425_y0, h_u_cla32_and4424_y0, h_u_cla32_and4426_y0);
  and_gate and_gate_h_u_cla32_and4427_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4427_y0);
  and_gate and_gate_h_u_cla32_and4428_y0(h_u_cla32_and4427_y0, h_u_cla32_and4426_y0, h_u_cla32_and4428_y0);
  and_gate and_gate_h_u_cla32_and4429_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4429_y0);
  and_gate and_gate_h_u_cla32_and4430_y0(h_u_cla32_and4429_y0, h_u_cla32_and4428_y0, h_u_cla32_and4430_y0);
  and_gate and_gate_h_u_cla32_and4431_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4431_y0);
  and_gate and_gate_h_u_cla32_and4432_y0(h_u_cla32_and4431_y0, h_u_cla32_and4430_y0, h_u_cla32_and4432_y0);
  and_gate and_gate_h_u_cla32_and4433_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4433_y0);
  and_gate and_gate_h_u_cla32_and4434_y0(h_u_cla32_and4433_y0, h_u_cla32_and4432_y0, h_u_cla32_and4434_y0);
  and_gate and_gate_h_u_cla32_and4435_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4435_y0);
  and_gate and_gate_h_u_cla32_and4436_y0(h_u_cla32_and4435_y0, h_u_cla32_and4434_y0, h_u_cla32_and4436_y0);
  and_gate and_gate_h_u_cla32_and4437_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4437_y0);
  and_gate and_gate_h_u_cla32_and4438_y0(h_u_cla32_and4437_y0, h_u_cla32_and4436_y0, h_u_cla32_and4438_y0);
  and_gate and_gate_h_u_cla32_and4439_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4439_y0);
  and_gate and_gate_h_u_cla32_and4440_y0(h_u_cla32_and4439_y0, h_u_cla32_and4438_y0, h_u_cla32_and4440_y0);
  and_gate and_gate_h_u_cla32_and4441_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4441_y0);
  and_gate and_gate_h_u_cla32_and4442_y0(h_u_cla32_and4441_y0, h_u_cla32_and4440_y0, h_u_cla32_and4442_y0);
  and_gate and_gate_h_u_cla32_and4443_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4443_y0);
  and_gate and_gate_h_u_cla32_and4444_y0(h_u_cla32_and4443_y0, h_u_cla32_and4442_y0, h_u_cla32_and4444_y0);
  and_gate and_gate_h_u_cla32_and4445_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4445_y0);
  and_gate and_gate_h_u_cla32_and4446_y0(h_u_cla32_and4445_y0, h_u_cla32_and4444_y0, h_u_cla32_and4446_y0);
  and_gate and_gate_h_u_cla32_and4447_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4447_y0);
  and_gate and_gate_h_u_cla32_and4448_y0(h_u_cla32_and4447_y0, h_u_cla32_and4446_y0, h_u_cla32_and4448_y0);
  and_gate and_gate_h_u_cla32_and4449_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4449_y0);
  and_gate and_gate_h_u_cla32_and4450_y0(h_u_cla32_and4449_y0, h_u_cla32_and4448_y0, h_u_cla32_and4450_y0);
  and_gate and_gate_h_u_cla32_and4451_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4451_y0);
  and_gate and_gate_h_u_cla32_and4452_y0(h_u_cla32_and4451_y0, h_u_cla32_and4450_y0, h_u_cla32_and4452_y0);
  and_gate and_gate_h_u_cla32_and4453_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4453_y0);
  and_gate and_gate_h_u_cla32_and4454_y0(h_u_cla32_and4453_y0, h_u_cla32_and4452_y0, h_u_cla32_and4454_y0);
  and_gate and_gate_h_u_cla32_and4455_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4455_y0);
  and_gate and_gate_h_u_cla32_and4456_y0(h_u_cla32_and4455_y0, h_u_cla32_and4454_y0, h_u_cla32_and4456_y0);
  and_gate and_gate_h_u_cla32_and4457_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4457_y0);
  and_gate and_gate_h_u_cla32_and4458_y0(h_u_cla32_and4457_y0, h_u_cla32_and4456_y0, h_u_cla32_and4458_y0);
  and_gate and_gate_h_u_cla32_and4459_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4459_y0);
  and_gate and_gate_h_u_cla32_and4460_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4460_y0);
  and_gate and_gate_h_u_cla32_and4461_y0(h_u_cla32_and4460_y0, h_u_cla32_and4459_y0, h_u_cla32_and4461_y0);
  and_gate and_gate_h_u_cla32_and4462_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4462_y0);
  and_gate and_gate_h_u_cla32_and4463_y0(h_u_cla32_and4462_y0, h_u_cla32_and4461_y0, h_u_cla32_and4463_y0);
  and_gate and_gate_h_u_cla32_and4464_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4464_y0);
  and_gate and_gate_h_u_cla32_and4465_y0(h_u_cla32_and4464_y0, h_u_cla32_and4463_y0, h_u_cla32_and4465_y0);
  and_gate and_gate_h_u_cla32_and4466_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4466_y0);
  and_gate and_gate_h_u_cla32_and4467_y0(h_u_cla32_and4466_y0, h_u_cla32_and4465_y0, h_u_cla32_and4467_y0);
  and_gate and_gate_h_u_cla32_and4468_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4468_y0);
  and_gate and_gate_h_u_cla32_and4469_y0(h_u_cla32_and4468_y0, h_u_cla32_and4467_y0, h_u_cla32_and4469_y0);
  and_gate and_gate_h_u_cla32_and4470_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4470_y0);
  and_gate and_gate_h_u_cla32_and4471_y0(h_u_cla32_and4470_y0, h_u_cla32_and4469_y0, h_u_cla32_and4471_y0);
  and_gate and_gate_h_u_cla32_and4472_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4472_y0);
  and_gate and_gate_h_u_cla32_and4473_y0(h_u_cla32_and4472_y0, h_u_cla32_and4471_y0, h_u_cla32_and4473_y0);
  and_gate and_gate_h_u_cla32_and4474_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4474_y0);
  and_gate and_gate_h_u_cla32_and4475_y0(h_u_cla32_and4474_y0, h_u_cla32_and4473_y0, h_u_cla32_and4475_y0);
  and_gate and_gate_h_u_cla32_and4476_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4476_y0);
  and_gate and_gate_h_u_cla32_and4477_y0(h_u_cla32_and4476_y0, h_u_cla32_and4475_y0, h_u_cla32_and4477_y0);
  and_gate and_gate_h_u_cla32_and4478_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4478_y0);
  and_gate and_gate_h_u_cla32_and4479_y0(h_u_cla32_and4478_y0, h_u_cla32_and4477_y0, h_u_cla32_and4479_y0);
  and_gate and_gate_h_u_cla32_and4480_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4480_y0);
  and_gate and_gate_h_u_cla32_and4481_y0(h_u_cla32_and4480_y0, h_u_cla32_and4479_y0, h_u_cla32_and4481_y0);
  and_gate and_gate_h_u_cla32_and4482_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4482_y0);
  and_gate and_gate_h_u_cla32_and4483_y0(h_u_cla32_and4482_y0, h_u_cla32_and4481_y0, h_u_cla32_and4483_y0);
  and_gate and_gate_h_u_cla32_and4484_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4484_y0);
  and_gate and_gate_h_u_cla32_and4485_y0(h_u_cla32_and4484_y0, h_u_cla32_and4483_y0, h_u_cla32_and4485_y0);
  and_gate and_gate_h_u_cla32_and4486_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4486_y0);
  and_gate and_gate_h_u_cla32_and4487_y0(h_u_cla32_and4486_y0, h_u_cla32_and4485_y0, h_u_cla32_and4487_y0);
  and_gate and_gate_h_u_cla32_and4488_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4488_y0);
  and_gate and_gate_h_u_cla32_and4489_y0(h_u_cla32_and4488_y0, h_u_cla32_and4487_y0, h_u_cla32_and4489_y0);
  and_gate and_gate_h_u_cla32_and4490_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4490_y0);
  and_gate and_gate_h_u_cla32_and4491_y0(h_u_cla32_and4490_y0, h_u_cla32_and4489_y0, h_u_cla32_and4491_y0);
  and_gate and_gate_h_u_cla32_and4492_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4492_y0);
  and_gate and_gate_h_u_cla32_and4493_y0(h_u_cla32_and4492_y0, h_u_cla32_and4491_y0, h_u_cla32_and4493_y0);
  and_gate and_gate_h_u_cla32_and4494_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4494_y0);
  and_gate and_gate_h_u_cla32_and4495_y0(h_u_cla32_and4494_y0, h_u_cla32_and4493_y0, h_u_cla32_and4495_y0);
  and_gate and_gate_h_u_cla32_and4496_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4496_y0);
  and_gate and_gate_h_u_cla32_and4497_y0(h_u_cla32_and4496_y0, h_u_cla32_and4495_y0, h_u_cla32_and4497_y0);
  and_gate and_gate_h_u_cla32_and4498_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and4498_y0);
  and_gate and_gate_h_u_cla32_and4499_y0(h_u_cla32_and4498_y0, h_u_cla32_and4497_y0, h_u_cla32_and4499_y0);
  and_gate and_gate_h_u_cla32_and4500_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4500_y0);
  and_gate and_gate_h_u_cla32_and4501_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4501_y0);
  and_gate and_gate_h_u_cla32_and4502_y0(h_u_cla32_and4501_y0, h_u_cla32_and4500_y0, h_u_cla32_and4502_y0);
  and_gate and_gate_h_u_cla32_and4503_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4503_y0);
  and_gate and_gate_h_u_cla32_and4504_y0(h_u_cla32_and4503_y0, h_u_cla32_and4502_y0, h_u_cla32_and4504_y0);
  and_gate and_gate_h_u_cla32_and4505_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4505_y0);
  and_gate and_gate_h_u_cla32_and4506_y0(h_u_cla32_and4505_y0, h_u_cla32_and4504_y0, h_u_cla32_and4506_y0);
  and_gate and_gate_h_u_cla32_and4507_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4507_y0);
  and_gate and_gate_h_u_cla32_and4508_y0(h_u_cla32_and4507_y0, h_u_cla32_and4506_y0, h_u_cla32_and4508_y0);
  and_gate and_gate_h_u_cla32_and4509_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4509_y0);
  and_gate and_gate_h_u_cla32_and4510_y0(h_u_cla32_and4509_y0, h_u_cla32_and4508_y0, h_u_cla32_and4510_y0);
  and_gate and_gate_h_u_cla32_and4511_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4511_y0);
  and_gate and_gate_h_u_cla32_and4512_y0(h_u_cla32_and4511_y0, h_u_cla32_and4510_y0, h_u_cla32_and4512_y0);
  and_gate and_gate_h_u_cla32_and4513_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4513_y0);
  and_gate and_gate_h_u_cla32_and4514_y0(h_u_cla32_and4513_y0, h_u_cla32_and4512_y0, h_u_cla32_and4514_y0);
  and_gate and_gate_h_u_cla32_and4515_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4515_y0);
  and_gate and_gate_h_u_cla32_and4516_y0(h_u_cla32_and4515_y0, h_u_cla32_and4514_y0, h_u_cla32_and4516_y0);
  and_gate and_gate_h_u_cla32_and4517_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4517_y0);
  and_gate and_gate_h_u_cla32_and4518_y0(h_u_cla32_and4517_y0, h_u_cla32_and4516_y0, h_u_cla32_and4518_y0);
  and_gate and_gate_h_u_cla32_and4519_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4519_y0);
  and_gate and_gate_h_u_cla32_and4520_y0(h_u_cla32_and4519_y0, h_u_cla32_and4518_y0, h_u_cla32_and4520_y0);
  and_gate and_gate_h_u_cla32_and4521_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4521_y0);
  and_gate and_gate_h_u_cla32_and4522_y0(h_u_cla32_and4521_y0, h_u_cla32_and4520_y0, h_u_cla32_and4522_y0);
  and_gate and_gate_h_u_cla32_and4523_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4523_y0);
  and_gate and_gate_h_u_cla32_and4524_y0(h_u_cla32_and4523_y0, h_u_cla32_and4522_y0, h_u_cla32_and4524_y0);
  and_gate and_gate_h_u_cla32_and4525_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4525_y0);
  and_gate and_gate_h_u_cla32_and4526_y0(h_u_cla32_and4525_y0, h_u_cla32_and4524_y0, h_u_cla32_and4526_y0);
  and_gate and_gate_h_u_cla32_and4527_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4527_y0);
  and_gate and_gate_h_u_cla32_and4528_y0(h_u_cla32_and4527_y0, h_u_cla32_and4526_y0, h_u_cla32_and4528_y0);
  and_gate and_gate_h_u_cla32_and4529_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4529_y0);
  and_gate and_gate_h_u_cla32_and4530_y0(h_u_cla32_and4529_y0, h_u_cla32_and4528_y0, h_u_cla32_and4530_y0);
  and_gate and_gate_h_u_cla32_and4531_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4531_y0);
  and_gate and_gate_h_u_cla32_and4532_y0(h_u_cla32_and4531_y0, h_u_cla32_and4530_y0, h_u_cla32_and4532_y0);
  and_gate and_gate_h_u_cla32_and4533_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4533_y0);
  and_gate and_gate_h_u_cla32_and4534_y0(h_u_cla32_and4533_y0, h_u_cla32_and4532_y0, h_u_cla32_and4534_y0);
  and_gate and_gate_h_u_cla32_and4535_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4535_y0);
  and_gate and_gate_h_u_cla32_and4536_y0(h_u_cla32_and4535_y0, h_u_cla32_and4534_y0, h_u_cla32_and4536_y0);
  and_gate and_gate_h_u_cla32_and4537_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and4537_y0);
  and_gate and_gate_h_u_cla32_and4538_y0(h_u_cla32_and4537_y0, h_u_cla32_and4536_y0, h_u_cla32_and4538_y0);
  and_gate and_gate_h_u_cla32_and4539_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4539_y0);
  and_gate and_gate_h_u_cla32_and4540_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4540_y0);
  and_gate and_gate_h_u_cla32_and4541_y0(h_u_cla32_and4540_y0, h_u_cla32_and4539_y0, h_u_cla32_and4541_y0);
  and_gate and_gate_h_u_cla32_and4542_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4542_y0);
  and_gate and_gate_h_u_cla32_and4543_y0(h_u_cla32_and4542_y0, h_u_cla32_and4541_y0, h_u_cla32_and4543_y0);
  and_gate and_gate_h_u_cla32_and4544_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4544_y0);
  and_gate and_gate_h_u_cla32_and4545_y0(h_u_cla32_and4544_y0, h_u_cla32_and4543_y0, h_u_cla32_and4545_y0);
  and_gate and_gate_h_u_cla32_and4546_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4546_y0);
  and_gate and_gate_h_u_cla32_and4547_y0(h_u_cla32_and4546_y0, h_u_cla32_and4545_y0, h_u_cla32_and4547_y0);
  and_gate and_gate_h_u_cla32_and4548_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4548_y0);
  and_gate and_gate_h_u_cla32_and4549_y0(h_u_cla32_and4548_y0, h_u_cla32_and4547_y0, h_u_cla32_and4549_y0);
  and_gate and_gate_h_u_cla32_and4550_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4550_y0);
  and_gate and_gate_h_u_cla32_and4551_y0(h_u_cla32_and4550_y0, h_u_cla32_and4549_y0, h_u_cla32_and4551_y0);
  and_gate and_gate_h_u_cla32_and4552_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4552_y0);
  and_gate and_gate_h_u_cla32_and4553_y0(h_u_cla32_and4552_y0, h_u_cla32_and4551_y0, h_u_cla32_and4553_y0);
  and_gate and_gate_h_u_cla32_and4554_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4554_y0);
  and_gate and_gate_h_u_cla32_and4555_y0(h_u_cla32_and4554_y0, h_u_cla32_and4553_y0, h_u_cla32_and4555_y0);
  and_gate and_gate_h_u_cla32_and4556_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4556_y0);
  and_gate and_gate_h_u_cla32_and4557_y0(h_u_cla32_and4556_y0, h_u_cla32_and4555_y0, h_u_cla32_and4557_y0);
  and_gate and_gate_h_u_cla32_and4558_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4558_y0);
  and_gate and_gate_h_u_cla32_and4559_y0(h_u_cla32_and4558_y0, h_u_cla32_and4557_y0, h_u_cla32_and4559_y0);
  and_gate and_gate_h_u_cla32_and4560_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4560_y0);
  and_gate and_gate_h_u_cla32_and4561_y0(h_u_cla32_and4560_y0, h_u_cla32_and4559_y0, h_u_cla32_and4561_y0);
  and_gate and_gate_h_u_cla32_and4562_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4562_y0);
  and_gate and_gate_h_u_cla32_and4563_y0(h_u_cla32_and4562_y0, h_u_cla32_and4561_y0, h_u_cla32_and4563_y0);
  and_gate and_gate_h_u_cla32_and4564_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4564_y0);
  and_gate and_gate_h_u_cla32_and4565_y0(h_u_cla32_and4564_y0, h_u_cla32_and4563_y0, h_u_cla32_and4565_y0);
  and_gate and_gate_h_u_cla32_and4566_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4566_y0);
  and_gate and_gate_h_u_cla32_and4567_y0(h_u_cla32_and4566_y0, h_u_cla32_and4565_y0, h_u_cla32_and4567_y0);
  and_gate and_gate_h_u_cla32_and4568_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4568_y0);
  and_gate and_gate_h_u_cla32_and4569_y0(h_u_cla32_and4568_y0, h_u_cla32_and4567_y0, h_u_cla32_and4569_y0);
  and_gate and_gate_h_u_cla32_and4570_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4570_y0);
  and_gate and_gate_h_u_cla32_and4571_y0(h_u_cla32_and4570_y0, h_u_cla32_and4569_y0, h_u_cla32_and4571_y0);
  and_gate and_gate_h_u_cla32_and4572_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4572_y0);
  and_gate and_gate_h_u_cla32_and4573_y0(h_u_cla32_and4572_y0, h_u_cla32_and4571_y0, h_u_cla32_and4573_y0);
  and_gate and_gate_h_u_cla32_and4574_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and4574_y0);
  and_gate and_gate_h_u_cla32_and4575_y0(h_u_cla32_and4574_y0, h_u_cla32_and4573_y0, h_u_cla32_and4575_y0);
  and_gate and_gate_h_u_cla32_and4576_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4576_y0);
  and_gate and_gate_h_u_cla32_and4577_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4577_y0);
  and_gate and_gate_h_u_cla32_and4578_y0(h_u_cla32_and4577_y0, h_u_cla32_and4576_y0, h_u_cla32_and4578_y0);
  and_gate and_gate_h_u_cla32_and4579_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4579_y0);
  and_gate and_gate_h_u_cla32_and4580_y0(h_u_cla32_and4579_y0, h_u_cla32_and4578_y0, h_u_cla32_and4580_y0);
  and_gate and_gate_h_u_cla32_and4581_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4581_y0);
  and_gate and_gate_h_u_cla32_and4582_y0(h_u_cla32_and4581_y0, h_u_cla32_and4580_y0, h_u_cla32_and4582_y0);
  and_gate and_gate_h_u_cla32_and4583_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4583_y0);
  and_gate and_gate_h_u_cla32_and4584_y0(h_u_cla32_and4583_y0, h_u_cla32_and4582_y0, h_u_cla32_and4584_y0);
  and_gate and_gate_h_u_cla32_and4585_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4585_y0);
  and_gate and_gate_h_u_cla32_and4586_y0(h_u_cla32_and4585_y0, h_u_cla32_and4584_y0, h_u_cla32_and4586_y0);
  and_gate and_gate_h_u_cla32_and4587_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4587_y0);
  and_gate and_gate_h_u_cla32_and4588_y0(h_u_cla32_and4587_y0, h_u_cla32_and4586_y0, h_u_cla32_and4588_y0);
  and_gate and_gate_h_u_cla32_and4589_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4589_y0);
  and_gate and_gate_h_u_cla32_and4590_y0(h_u_cla32_and4589_y0, h_u_cla32_and4588_y0, h_u_cla32_and4590_y0);
  and_gate and_gate_h_u_cla32_and4591_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4591_y0);
  and_gate and_gate_h_u_cla32_and4592_y0(h_u_cla32_and4591_y0, h_u_cla32_and4590_y0, h_u_cla32_and4592_y0);
  and_gate and_gate_h_u_cla32_and4593_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4593_y0);
  and_gate and_gate_h_u_cla32_and4594_y0(h_u_cla32_and4593_y0, h_u_cla32_and4592_y0, h_u_cla32_and4594_y0);
  and_gate and_gate_h_u_cla32_and4595_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4595_y0);
  and_gate and_gate_h_u_cla32_and4596_y0(h_u_cla32_and4595_y0, h_u_cla32_and4594_y0, h_u_cla32_and4596_y0);
  and_gate and_gate_h_u_cla32_and4597_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4597_y0);
  and_gate and_gate_h_u_cla32_and4598_y0(h_u_cla32_and4597_y0, h_u_cla32_and4596_y0, h_u_cla32_and4598_y0);
  and_gate and_gate_h_u_cla32_and4599_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4599_y0);
  and_gate and_gate_h_u_cla32_and4600_y0(h_u_cla32_and4599_y0, h_u_cla32_and4598_y0, h_u_cla32_and4600_y0);
  and_gate and_gate_h_u_cla32_and4601_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4601_y0);
  and_gate and_gate_h_u_cla32_and4602_y0(h_u_cla32_and4601_y0, h_u_cla32_and4600_y0, h_u_cla32_and4602_y0);
  and_gate and_gate_h_u_cla32_and4603_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4603_y0);
  and_gate and_gate_h_u_cla32_and4604_y0(h_u_cla32_and4603_y0, h_u_cla32_and4602_y0, h_u_cla32_and4604_y0);
  and_gate and_gate_h_u_cla32_and4605_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4605_y0);
  and_gate and_gate_h_u_cla32_and4606_y0(h_u_cla32_and4605_y0, h_u_cla32_and4604_y0, h_u_cla32_and4606_y0);
  and_gate and_gate_h_u_cla32_and4607_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4607_y0);
  and_gate and_gate_h_u_cla32_and4608_y0(h_u_cla32_and4607_y0, h_u_cla32_and4606_y0, h_u_cla32_and4608_y0);
  and_gate and_gate_h_u_cla32_and4609_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and4609_y0);
  and_gate and_gate_h_u_cla32_and4610_y0(h_u_cla32_and4609_y0, h_u_cla32_and4608_y0, h_u_cla32_and4610_y0);
  and_gate and_gate_h_u_cla32_and4611_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4611_y0);
  and_gate and_gate_h_u_cla32_and4612_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4612_y0);
  and_gate and_gate_h_u_cla32_and4613_y0(h_u_cla32_and4612_y0, h_u_cla32_and4611_y0, h_u_cla32_and4613_y0);
  and_gate and_gate_h_u_cla32_and4614_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4614_y0);
  and_gate and_gate_h_u_cla32_and4615_y0(h_u_cla32_and4614_y0, h_u_cla32_and4613_y0, h_u_cla32_and4615_y0);
  and_gate and_gate_h_u_cla32_and4616_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4616_y0);
  and_gate and_gate_h_u_cla32_and4617_y0(h_u_cla32_and4616_y0, h_u_cla32_and4615_y0, h_u_cla32_and4617_y0);
  and_gate and_gate_h_u_cla32_and4618_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4618_y0);
  and_gate and_gate_h_u_cla32_and4619_y0(h_u_cla32_and4618_y0, h_u_cla32_and4617_y0, h_u_cla32_and4619_y0);
  and_gate and_gate_h_u_cla32_and4620_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4620_y0);
  and_gate and_gate_h_u_cla32_and4621_y0(h_u_cla32_and4620_y0, h_u_cla32_and4619_y0, h_u_cla32_and4621_y0);
  and_gate and_gate_h_u_cla32_and4622_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4622_y0);
  and_gate and_gate_h_u_cla32_and4623_y0(h_u_cla32_and4622_y0, h_u_cla32_and4621_y0, h_u_cla32_and4623_y0);
  and_gate and_gate_h_u_cla32_and4624_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4624_y0);
  and_gate and_gate_h_u_cla32_and4625_y0(h_u_cla32_and4624_y0, h_u_cla32_and4623_y0, h_u_cla32_and4625_y0);
  and_gate and_gate_h_u_cla32_and4626_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4626_y0);
  and_gate and_gate_h_u_cla32_and4627_y0(h_u_cla32_and4626_y0, h_u_cla32_and4625_y0, h_u_cla32_and4627_y0);
  and_gate and_gate_h_u_cla32_and4628_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4628_y0);
  and_gate and_gate_h_u_cla32_and4629_y0(h_u_cla32_and4628_y0, h_u_cla32_and4627_y0, h_u_cla32_and4629_y0);
  and_gate and_gate_h_u_cla32_and4630_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4630_y0);
  and_gate and_gate_h_u_cla32_and4631_y0(h_u_cla32_and4630_y0, h_u_cla32_and4629_y0, h_u_cla32_and4631_y0);
  and_gate and_gate_h_u_cla32_and4632_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4632_y0);
  and_gate and_gate_h_u_cla32_and4633_y0(h_u_cla32_and4632_y0, h_u_cla32_and4631_y0, h_u_cla32_and4633_y0);
  and_gate and_gate_h_u_cla32_and4634_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4634_y0);
  and_gate and_gate_h_u_cla32_and4635_y0(h_u_cla32_and4634_y0, h_u_cla32_and4633_y0, h_u_cla32_and4635_y0);
  and_gate and_gate_h_u_cla32_and4636_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4636_y0);
  and_gate and_gate_h_u_cla32_and4637_y0(h_u_cla32_and4636_y0, h_u_cla32_and4635_y0, h_u_cla32_and4637_y0);
  and_gate and_gate_h_u_cla32_and4638_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4638_y0);
  and_gate and_gate_h_u_cla32_and4639_y0(h_u_cla32_and4638_y0, h_u_cla32_and4637_y0, h_u_cla32_and4639_y0);
  and_gate and_gate_h_u_cla32_and4640_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4640_y0);
  and_gate and_gate_h_u_cla32_and4641_y0(h_u_cla32_and4640_y0, h_u_cla32_and4639_y0, h_u_cla32_and4641_y0);
  and_gate and_gate_h_u_cla32_and4642_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and4642_y0);
  and_gate and_gate_h_u_cla32_and4643_y0(h_u_cla32_and4642_y0, h_u_cla32_and4641_y0, h_u_cla32_and4643_y0);
  and_gate and_gate_h_u_cla32_and4644_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4644_y0);
  and_gate and_gate_h_u_cla32_and4645_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4645_y0);
  and_gate and_gate_h_u_cla32_and4646_y0(h_u_cla32_and4645_y0, h_u_cla32_and4644_y0, h_u_cla32_and4646_y0);
  and_gate and_gate_h_u_cla32_and4647_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4647_y0);
  and_gate and_gate_h_u_cla32_and4648_y0(h_u_cla32_and4647_y0, h_u_cla32_and4646_y0, h_u_cla32_and4648_y0);
  and_gate and_gate_h_u_cla32_and4649_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4649_y0);
  and_gate and_gate_h_u_cla32_and4650_y0(h_u_cla32_and4649_y0, h_u_cla32_and4648_y0, h_u_cla32_and4650_y0);
  and_gate and_gate_h_u_cla32_and4651_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4651_y0);
  and_gate and_gate_h_u_cla32_and4652_y0(h_u_cla32_and4651_y0, h_u_cla32_and4650_y0, h_u_cla32_and4652_y0);
  and_gate and_gate_h_u_cla32_and4653_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4653_y0);
  and_gate and_gate_h_u_cla32_and4654_y0(h_u_cla32_and4653_y0, h_u_cla32_and4652_y0, h_u_cla32_and4654_y0);
  and_gate and_gate_h_u_cla32_and4655_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4655_y0);
  and_gate and_gate_h_u_cla32_and4656_y0(h_u_cla32_and4655_y0, h_u_cla32_and4654_y0, h_u_cla32_and4656_y0);
  and_gate and_gate_h_u_cla32_and4657_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4657_y0);
  and_gate and_gate_h_u_cla32_and4658_y0(h_u_cla32_and4657_y0, h_u_cla32_and4656_y0, h_u_cla32_and4658_y0);
  and_gate and_gate_h_u_cla32_and4659_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4659_y0);
  and_gate and_gate_h_u_cla32_and4660_y0(h_u_cla32_and4659_y0, h_u_cla32_and4658_y0, h_u_cla32_and4660_y0);
  and_gate and_gate_h_u_cla32_and4661_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4661_y0);
  and_gate and_gate_h_u_cla32_and4662_y0(h_u_cla32_and4661_y0, h_u_cla32_and4660_y0, h_u_cla32_and4662_y0);
  and_gate and_gate_h_u_cla32_and4663_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4663_y0);
  and_gate and_gate_h_u_cla32_and4664_y0(h_u_cla32_and4663_y0, h_u_cla32_and4662_y0, h_u_cla32_and4664_y0);
  and_gate and_gate_h_u_cla32_and4665_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4665_y0);
  and_gate and_gate_h_u_cla32_and4666_y0(h_u_cla32_and4665_y0, h_u_cla32_and4664_y0, h_u_cla32_and4666_y0);
  and_gate and_gate_h_u_cla32_and4667_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4667_y0);
  and_gate and_gate_h_u_cla32_and4668_y0(h_u_cla32_and4667_y0, h_u_cla32_and4666_y0, h_u_cla32_and4668_y0);
  and_gate and_gate_h_u_cla32_and4669_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4669_y0);
  and_gate and_gate_h_u_cla32_and4670_y0(h_u_cla32_and4669_y0, h_u_cla32_and4668_y0, h_u_cla32_and4670_y0);
  and_gate and_gate_h_u_cla32_and4671_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4671_y0);
  and_gate and_gate_h_u_cla32_and4672_y0(h_u_cla32_and4671_y0, h_u_cla32_and4670_y0, h_u_cla32_and4672_y0);
  and_gate and_gate_h_u_cla32_and4673_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and4673_y0);
  and_gate and_gate_h_u_cla32_and4674_y0(h_u_cla32_and4673_y0, h_u_cla32_and4672_y0, h_u_cla32_and4674_y0);
  and_gate and_gate_h_u_cla32_and4675_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4675_y0);
  and_gate and_gate_h_u_cla32_and4676_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4676_y0);
  and_gate and_gate_h_u_cla32_and4677_y0(h_u_cla32_and4676_y0, h_u_cla32_and4675_y0, h_u_cla32_and4677_y0);
  and_gate and_gate_h_u_cla32_and4678_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4678_y0);
  and_gate and_gate_h_u_cla32_and4679_y0(h_u_cla32_and4678_y0, h_u_cla32_and4677_y0, h_u_cla32_and4679_y0);
  and_gate and_gate_h_u_cla32_and4680_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4680_y0);
  and_gate and_gate_h_u_cla32_and4681_y0(h_u_cla32_and4680_y0, h_u_cla32_and4679_y0, h_u_cla32_and4681_y0);
  and_gate and_gate_h_u_cla32_and4682_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4682_y0);
  and_gate and_gate_h_u_cla32_and4683_y0(h_u_cla32_and4682_y0, h_u_cla32_and4681_y0, h_u_cla32_and4683_y0);
  and_gate and_gate_h_u_cla32_and4684_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4684_y0);
  and_gate and_gate_h_u_cla32_and4685_y0(h_u_cla32_and4684_y0, h_u_cla32_and4683_y0, h_u_cla32_and4685_y0);
  and_gate and_gate_h_u_cla32_and4686_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4686_y0);
  and_gate and_gate_h_u_cla32_and4687_y0(h_u_cla32_and4686_y0, h_u_cla32_and4685_y0, h_u_cla32_and4687_y0);
  and_gate and_gate_h_u_cla32_and4688_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4688_y0);
  and_gate and_gate_h_u_cla32_and4689_y0(h_u_cla32_and4688_y0, h_u_cla32_and4687_y0, h_u_cla32_and4689_y0);
  and_gate and_gate_h_u_cla32_and4690_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4690_y0);
  and_gate and_gate_h_u_cla32_and4691_y0(h_u_cla32_and4690_y0, h_u_cla32_and4689_y0, h_u_cla32_and4691_y0);
  and_gate and_gate_h_u_cla32_and4692_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4692_y0);
  and_gate and_gate_h_u_cla32_and4693_y0(h_u_cla32_and4692_y0, h_u_cla32_and4691_y0, h_u_cla32_and4693_y0);
  and_gate and_gate_h_u_cla32_and4694_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4694_y0);
  and_gate and_gate_h_u_cla32_and4695_y0(h_u_cla32_and4694_y0, h_u_cla32_and4693_y0, h_u_cla32_and4695_y0);
  and_gate and_gate_h_u_cla32_and4696_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4696_y0);
  and_gate and_gate_h_u_cla32_and4697_y0(h_u_cla32_and4696_y0, h_u_cla32_and4695_y0, h_u_cla32_and4697_y0);
  and_gate and_gate_h_u_cla32_and4698_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4698_y0);
  and_gate and_gate_h_u_cla32_and4699_y0(h_u_cla32_and4698_y0, h_u_cla32_and4697_y0, h_u_cla32_and4699_y0);
  and_gate and_gate_h_u_cla32_and4700_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4700_y0);
  and_gate and_gate_h_u_cla32_and4701_y0(h_u_cla32_and4700_y0, h_u_cla32_and4699_y0, h_u_cla32_and4701_y0);
  and_gate and_gate_h_u_cla32_and4702_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and4702_y0);
  and_gate and_gate_h_u_cla32_and4703_y0(h_u_cla32_and4702_y0, h_u_cla32_and4701_y0, h_u_cla32_and4703_y0);
  and_gate and_gate_h_u_cla32_and4704_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4704_y0);
  and_gate and_gate_h_u_cla32_and4705_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4705_y0);
  and_gate and_gate_h_u_cla32_and4706_y0(h_u_cla32_and4705_y0, h_u_cla32_and4704_y0, h_u_cla32_and4706_y0);
  and_gate and_gate_h_u_cla32_and4707_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4707_y0);
  and_gate and_gate_h_u_cla32_and4708_y0(h_u_cla32_and4707_y0, h_u_cla32_and4706_y0, h_u_cla32_and4708_y0);
  and_gate and_gate_h_u_cla32_and4709_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4709_y0);
  and_gate and_gate_h_u_cla32_and4710_y0(h_u_cla32_and4709_y0, h_u_cla32_and4708_y0, h_u_cla32_and4710_y0);
  and_gate and_gate_h_u_cla32_and4711_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4711_y0);
  and_gate and_gate_h_u_cla32_and4712_y0(h_u_cla32_and4711_y0, h_u_cla32_and4710_y0, h_u_cla32_and4712_y0);
  and_gate and_gate_h_u_cla32_and4713_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4713_y0);
  and_gate and_gate_h_u_cla32_and4714_y0(h_u_cla32_and4713_y0, h_u_cla32_and4712_y0, h_u_cla32_and4714_y0);
  and_gate and_gate_h_u_cla32_and4715_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4715_y0);
  and_gate and_gate_h_u_cla32_and4716_y0(h_u_cla32_and4715_y0, h_u_cla32_and4714_y0, h_u_cla32_and4716_y0);
  and_gate and_gate_h_u_cla32_and4717_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4717_y0);
  and_gate and_gate_h_u_cla32_and4718_y0(h_u_cla32_and4717_y0, h_u_cla32_and4716_y0, h_u_cla32_and4718_y0);
  and_gate and_gate_h_u_cla32_and4719_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4719_y0);
  and_gate and_gate_h_u_cla32_and4720_y0(h_u_cla32_and4719_y0, h_u_cla32_and4718_y0, h_u_cla32_and4720_y0);
  and_gate and_gate_h_u_cla32_and4721_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4721_y0);
  and_gate and_gate_h_u_cla32_and4722_y0(h_u_cla32_and4721_y0, h_u_cla32_and4720_y0, h_u_cla32_and4722_y0);
  and_gate and_gate_h_u_cla32_and4723_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4723_y0);
  and_gate and_gate_h_u_cla32_and4724_y0(h_u_cla32_and4723_y0, h_u_cla32_and4722_y0, h_u_cla32_and4724_y0);
  and_gate and_gate_h_u_cla32_and4725_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4725_y0);
  and_gate and_gate_h_u_cla32_and4726_y0(h_u_cla32_and4725_y0, h_u_cla32_and4724_y0, h_u_cla32_and4726_y0);
  and_gate and_gate_h_u_cla32_and4727_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4727_y0);
  and_gate and_gate_h_u_cla32_and4728_y0(h_u_cla32_and4727_y0, h_u_cla32_and4726_y0, h_u_cla32_and4728_y0);
  and_gate and_gate_h_u_cla32_and4729_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and4729_y0);
  and_gate and_gate_h_u_cla32_and4730_y0(h_u_cla32_and4729_y0, h_u_cla32_and4728_y0, h_u_cla32_and4730_y0);
  and_gate and_gate_h_u_cla32_and4731_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4731_y0);
  and_gate and_gate_h_u_cla32_and4732_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4732_y0);
  and_gate and_gate_h_u_cla32_and4733_y0(h_u_cla32_and4732_y0, h_u_cla32_and4731_y0, h_u_cla32_and4733_y0);
  and_gate and_gate_h_u_cla32_and4734_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4734_y0);
  and_gate and_gate_h_u_cla32_and4735_y0(h_u_cla32_and4734_y0, h_u_cla32_and4733_y0, h_u_cla32_and4735_y0);
  and_gate and_gate_h_u_cla32_and4736_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4736_y0);
  and_gate and_gate_h_u_cla32_and4737_y0(h_u_cla32_and4736_y0, h_u_cla32_and4735_y0, h_u_cla32_and4737_y0);
  and_gate and_gate_h_u_cla32_and4738_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4738_y0);
  and_gate and_gate_h_u_cla32_and4739_y0(h_u_cla32_and4738_y0, h_u_cla32_and4737_y0, h_u_cla32_and4739_y0);
  and_gate and_gate_h_u_cla32_and4740_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4740_y0);
  and_gate and_gate_h_u_cla32_and4741_y0(h_u_cla32_and4740_y0, h_u_cla32_and4739_y0, h_u_cla32_and4741_y0);
  and_gate and_gate_h_u_cla32_and4742_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4742_y0);
  and_gate and_gate_h_u_cla32_and4743_y0(h_u_cla32_and4742_y0, h_u_cla32_and4741_y0, h_u_cla32_and4743_y0);
  and_gate and_gate_h_u_cla32_and4744_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4744_y0);
  and_gate and_gate_h_u_cla32_and4745_y0(h_u_cla32_and4744_y0, h_u_cla32_and4743_y0, h_u_cla32_and4745_y0);
  and_gate and_gate_h_u_cla32_and4746_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4746_y0);
  and_gate and_gate_h_u_cla32_and4747_y0(h_u_cla32_and4746_y0, h_u_cla32_and4745_y0, h_u_cla32_and4747_y0);
  and_gate and_gate_h_u_cla32_and4748_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4748_y0);
  and_gate and_gate_h_u_cla32_and4749_y0(h_u_cla32_and4748_y0, h_u_cla32_and4747_y0, h_u_cla32_and4749_y0);
  and_gate and_gate_h_u_cla32_and4750_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4750_y0);
  and_gate and_gate_h_u_cla32_and4751_y0(h_u_cla32_and4750_y0, h_u_cla32_and4749_y0, h_u_cla32_and4751_y0);
  and_gate and_gate_h_u_cla32_and4752_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4752_y0);
  and_gate and_gate_h_u_cla32_and4753_y0(h_u_cla32_and4752_y0, h_u_cla32_and4751_y0, h_u_cla32_and4753_y0);
  and_gate and_gate_h_u_cla32_and4754_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and4754_y0);
  and_gate and_gate_h_u_cla32_and4755_y0(h_u_cla32_and4754_y0, h_u_cla32_and4753_y0, h_u_cla32_and4755_y0);
  and_gate and_gate_h_u_cla32_and4756_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4756_y0);
  and_gate and_gate_h_u_cla32_and4757_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4757_y0);
  and_gate and_gate_h_u_cla32_and4758_y0(h_u_cla32_and4757_y0, h_u_cla32_and4756_y0, h_u_cla32_and4758_y0);
  and_gate and_gate_h_u_cla32_and4759_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4759_y0);
  and_gate and_gate_h_u_cla32_and4760_y0(h_u_cla32_and4759_y0, h_u_cla32_and4758_y0, h_u_cla32_and4760_y0);
  and_gate and_gate_h_u_cla32_and4761_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4761_y0);
  and_gate and_gate_h_u_cla32_and4762_y0(h_u_cla32_and4761_y0, h_u_cla32_and4760_y0, h_u_cla32_and4762_y0);
  and_gate and_gate_h_u_cla32_and4763_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4763_y0);
  and_gate and_gate_h_u_cla32_and4764_y0(h_u_cla32_and4763_y0, h_u_cla32_and4762_y0, h_u_cla32_and4764_y0);
  and_gate and_gate_h_u_cla32_and4765_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4765_y0);
  and_gate and_gate_h_u_cla32_and4766_y0(h_u_cla32_and4765_y0, h_u_cla32_and4764_y0, h_u_cla32_and4766_y0);
  and_gate and_gate_h_u_cla32_and4767_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4767_y0);
  and_gate and_gate_h_u_cla32_and4768_y0(h_u_cla32_and4767_y0, h_u_cla32_and4766_y0, h_u_cla32_and4768_y0);
  and_gate and_gate_h_u_cla32_and4769_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4769_y0);
  and_gate and_gate_h_u_cla32_and4770_y0(h_u_cla32_and4769_y0, h_u_cla32_and4768_y0, h_u_cla32_and4770_y0);
  and_gate and_gate_h_u_cla32_and4771_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4771_y0);
  and_gate and_gate_h_u_cla32_and4772_y0(h_u_cla32_and4771_y0, h_u_cla32_and4770_y0, h_u_cla32_and4772_y0);
  and_gate and_gate_h_u_cla32_and4773_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4773_y0);
  and_gate and_gate_h_u_cla32_and4774_y0(h_u_cla32_and4773_y0, h_u_cla32_and4772_y0, h_u_cla32_and4774_y0);
  and_gate and_gate_h_u_cla32_and4775_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4775_y0);
  and_gate and_gate_h_u_cla32_and4776_y0(h_u_cla32_and4775_y0, h_u_cla32_and4774_y0, h_u_cla32_and4776_y0);
  and_gate and_gate_h_u_cla32_and4777_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and4777_y0);
  and_gate and_gate_h_u_cla32_and4778_y0(h_u_cla32_and4777_y0, h_u_cla32_and4776_y0, h_u_cla32_and4778_y0);
  and_gate and_gate_h_u_cla32_and4779_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4779_y0);
  and_gate and_gate_h_u_cla32_and4780_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4780_y0);
  and_gate and_gate_h_u_cla32_and4781_y0(h_u_cla32_and4780_y0, h_u_cla32_and4779_y0, h_u_cla32_and4781_y0);
  and_gate and_gate_h_u_cla32_and4782_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4782_y0);
  and_gate and_gate_h_u_cla32_and4783_y0(h_u_cla32_and4782_y0, h_u_cla32_and4781_y0, h_u_cla32_and4783_y0);
  and_gate and_gate_h_u_cla32_and4784_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4784_y0);
  and_gate and_gate_h_u_cla32_and4785_y0(h_u_cla32_and4784_y0, h_u_cla32_and4783_y0, h_u_cla32_and4785_y0);
  and_gate and_gate_h_u_cla32_and4786_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4786_y0);
  and_gate and_gate_h_u_cla32_and4787_y0(h_u_cla32_and4786_y0, h_u_cla32_and4785_y0, h_u_cla32_and4787_y0);
  and_gate and_gate_h_u_cla32_and4788_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4788_y0);
  and_gate and_gate_h_u_cla32_and4789_y0(h_u_cla32_and4788_y0, h_u_cla32_and4787_y0, h_u_cla32_and4789_y0);
  and_gate and_gate_h_u_cla32_and4790_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4790_y0);
  and_gate and_gate_h_u_cla32_and4791_y0(h_u_cla32_and4790_y0, h_u_cla32_and4789_y0, h_u_cla32_and4791_y0);
  and_gate and_gate_h_u_cla32_and4792_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4792_y0);
  and_gate and_gate_h_u_cla32_and4793_y0(h_u_cla32_and4792_y0, h_u_cla32_and4791_y0, h_u_cla32_and4793_y0);
  and_gate and_gate_h_u_cla32_and4794_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4794_y0);
  and_gate and_gate_h_u_cla32_and4795_y0(h_u_cla32_and4794_y0, h_u_cla32_and4793_y0, h_u_cla32_and4795_y0);
  and_gate and_gate_h_u_cla32_and4796_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4796_y0);
  and_gate and_gate_h_u_cla32_and4797_y0(h_u_cla32_and4796_y0, h_u_cla32_and4795_y0, h_u_cla32_and4797_y0);
  and_gate and_gate_h_u_cla32_and4798_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and4798_y0);
  and_gate and_gate_h_u_cla32_and4799_y0(h_u_cla32_and4798_y0, h_u_cla32_and4797_y0, h_u_cla32_and4799_y0);
  and_gate and_gate_h_u_cla32_and4800_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4800_y0);
  and_gate and_gate_h_u_cla32_and4801_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4801_y0);
  and_gate and_gate_h_u_cla32_and4802_y0(h_u_cla32_and4801_y0, h_u_cla32_and4800_y0, h_u_cla32_and4802_y0);
  and_gate and_gate_h_u_cla32_and4803_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4803_y0);
  and_gate and_gate_h_u_cla32_and4804_y0(h_u_cla32_and4803_y0, h_u_cla32_and4802_y0, h_u_cla32_and4804_y0);
  and_gate and_gate_h_u_cla32_and4805_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4805_y0);
  and_gate and_gate_h_u_cla32_and4806_y0(h_u_cla32_and4805_y0, h_u_cla32_and4804_y0, h_u_cla32_and4806_y0);
  and_gate and_gate_h_u_cla32_and4807_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4807_y0);
  and_gate and_gate_h_u_cla32_and4808_y0(h_u_cla32_and4807_y0, h_u_cla32_and4806_y0, h_u_cla32_and4808_y0);
  and_gate and_gate_h_u_cla32_and4809_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4809_y0);
  and_gate and_gate_h_u_cla32_and4810_y0(h_u_cla32_and4809_y0, h_u_cla32_and4808_y0, h_u_cla32_and4810_y0);
  and_gate and_gate_h_u_cla32_and4811_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4811_y0);
  and_gate and_gate_h_u_cla32_and4812_y0(h_u_cla32_and4811_y0, h_u_cla32_and4810_y0, h_u_cla32_and4812_y0);
  and_gate and_gate_h_u_cla32_and4813_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4813_y0);
  and_gate and_gate_h_u_cla32_and4814_y0(h_u_cla32_and4813_y0, h_u_cla32_and4812_y0, h_u_cla32_and4814_y0);
  and_gate and_gate_h_u_cla32_and4815_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4815_y0);
  and_gate and_gate_h_u_cla32_and4816_y0(h_u_cla32_and4815_y0, h_u_cla32_and4814_y0, h_u_cla32_and4816_y0);
  and_gate and_gate_h_u_cla32_and4817_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and4817_y0);
  and_gate and_gate_h_u_cla32_and4818_y0(h_u_cla32_and4817_y0, h_u_cla32_and4816_y0, h_u_cla32_and4818_y0);
  and_gate and_gate_h_u_cla32_and4819_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4819_y0);
  and_gate and_gate_h_u_cla32_and4820_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4820_y0);
  and_gate and_gate_h_u_cla32_and4821_y0(h_u_cla32_and4820_y0, h_u_cla32_and4819_y0, h_u_cla32_and4821_y0);
  and_gate and_gate_h_u_cla32_and4822_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4822_y0);
  and_gate and_gate_h_u_cla32_and4823_y0(h_u_cla32_and4822_y0, h_u_cla32_and4821_y0, h_u_cla32_and4823_y0);
  and_gate and_gate_h_u_cla32_and4824_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4824_y0);
  and_gate and_gate_h_u_cla32_and4825_y0(h_u_cla32_and4824_y0, h_u_cla32_and4823_y0, h_u_cla32_and4825_y0);
  and_gate and_gate_h_u_cla32_and4826_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4826_y0);
  and_gate and_gate_h_u_cla32_and4827_y0(h_u_cla32_and4826_y0, h_u_cla32_and4825_y0, h_u_cla32_and4827_y0);
  and_gate and_gate_h_u_cla32_and4828_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4828_y0);
  and_gate and_gate_h_u_cla32_and4829_y0(h_u_cla32_and4828_y0, h_u_cla32_and4827_y0, h_u_cla32_and4829_y0);
  and_gate and_gate_h_u_cla32_and4830_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4830_y0);
  and_gate and_gate_h_u_cla32_and4831_y0(h_u_cla32_and4830_y0, h_u_cla32_and4829_y0, h_u_cla32_and4831_y0);
  and_gate and_gate_h_u_cla32_and4832_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4832_y0);
  and_gate and_gate_h_u_cla32_and4833_y0(h_u_cla32_and4832_y0, h_u_cla32_and4831_y0, h_u_cla32_and4833_y0);
  and_gate and_gate_h_u_cla32_and4834_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and4834_y0);
  and_gate and_gate_h_u_cla32_and4835_y0(h_u_cla32_and4834_y0, h_u_cla32_and4833_y0, h_u_cla32_and4835_y0);
  and_gate and_gate_h_u_cla32_and4836_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4836_y0);
  and_gate and_gate_h_u_cla32_and4837_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4837_y0);
  and_gate and_gate_h_u_cla32_and4838_y0(h_u_cla32_and4837_y0, h_u_cla32_and4836_y0, h_u_cla32_and4838_y0);
  and_gate and_gate_h_u_cla32_and4839_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4839_y0);
  and_gate and_gate_h_u_cla32_and4840_y0(h_u_cla32_and4839_y0, h_u_cla32_and4838_y0, h_u_cla32_and4840_y0);
  and_gate and_gate_h_u_cla32_and4841_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4841_y0);
  and_gate and_gate_h_u_cla32_and4842_y0(h_u_cla32_and4841_y0, h_u_cla32_and4840_y0, h_u_cla32_and4842_y0);
  and_gate and_gate_h_u_cla32_and4843_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4843_y0);
  and_gate and_gate_h_u_cla32_and4844_y0(h_u_cla32_and4843_y0, h_u_cla32_and4842_y0, h_u_cla32_and4844_y0);
  and_gate and_gate_h_u_cla32_and4845_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4845_y0);
  and_gate and_gate_h_u_cla32_and4846_y0(h_u_cla32_and4845_y0, h_u_cla32_and4844_y0, h_u_cla32_and4846_y0);
  and_gate and_gate_h_u_cla32_and4847_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4847_y0);
  and_gate and_gate_h_u_cla32_and4848_y0(h_u_cla32_and4847_y0, h_u_cla32_and4846_y0, h_u_cla32_and4848_y0);
  and_gate and_gate_h_u_cla32_and4849_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and4849_y0);
  and_gate and_gate_h_u_cla32_and4850_y0(h_u_cla32_and4849_y0, h_u_cla32_and4848_y0, h_u_cla32_and4850_y0);
  and_gate and_gate_h_u_cla32_and4851_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4851_y0);
  and_gate and_gate_h_u_cla32_and4852_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4852_y0);
  and_gate and_gate_h_u_cla32_and4853_y0(h_u_cla32_and4852_y0, h_u_cla32_and4851_y0, h_u_cla32_and4853_y0);
  and_gate and_gate_h_u_cla32_and4854_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4854_y0);
  and_gate and_gate_h_u_cla32_and4855_y0(h_u_cla32_and4854_y0, h_u_cla32_and4853_y0, h_u_cla32_and4855_y0);
  and_gate and_gate_h_u_cla32_and4856_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4856_y0);
  and_gate and_gate_h_u_cla32_and4857_y0(h_u_cla32_and4856_y0, h_u_cla32_and4855_y0, h_u_cla32_and4857_y0);
  and_gate and_gate_h_u_cla32_and4858_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4858_y0);
  and_gate and_gate_h_u_cla32_and4859_y0(h_u_cla32_and4858_y0, h_u_cla32_and4857_y0, h_u_cla32_and4859_y0);
  and_gate and_gate_h_u_cla32_and4860_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4860_y0);
  and_gate and_gate_h_u_cla32_and4861_y0(h_u_cla32_and4860_y0, h_u_cla32_and4859_y0, h_u_cla32_and4861_y0);
  and_gate and_gate_h_u_cla32_and4862_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and4862_y0);
  and_gate and_gate_h_u_cla32_and4863_y0(h_u_cla32_and4862_y0, h_u_cla32_and4861_y0, h_u_cla32_and4863_y0);
  and_gate and_gate_h_u_cla32_and4864_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4864_y0);
  and_gate and_gate_h_u_cla32_and4865_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4865_y0);
  and_gate and_gate_h_u_cla32_and4866_y0(h_u_cla32_and4865_y0, h_u_cla32_and4864_y0, h_u_cla32_and4866_y0);
  and_gate and_gate_h_u_cla32_and4867_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4867_y0);
  and_gate and_gate_h_u_cla32_and4868_y0(h_u_cla32_and4867_y0, h_u_cla32_and4866_y0, h_u_cla32_and4868_y0);
  and_gate and_gate_h_u_cla32_and4869_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4869_y0);
  and_gate and_gate_h_u_cla32_and4870_y0(h_u_cla32_and4869_y0, h_u_cla32_and4868_y0, h_u_cla32_and4870_y0);
  and_gate and_gate_h_u_cla32_and4871_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4871_y0);
  and_gate and_gate_h_u_cla32_and4872_y0(h_u_cla32_and4871_y0, h_u_cla32_and4870_y0, h_u_cla32_and4872_y0);
  and_gate and_gate_h_u_cla32_and4873_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and4873_y0);
  and_gate and_gate_h_u_cla32_and4874_y0(h_u_cla32_and4873_y0, h_u_cla32_and4872_y0, h_u_cla32_and4874_y0);
  and_gate and_gate_h_u_cla32_and4875_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4875_y0);
  and_gate and_gate_h_u_cla32_and4876_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4876_y0);
  and_gate and_gate_h_u_cla32_and4877_y0(h_u_cla32_and4876_y0, h_u_cla32_and4875_y0, h_u_cla32_and4877_y0);
  and_gate and_gate_h_u_cla32_and4878_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4878_y0);
  and_gate and_gate_h_u_cla32_and4879_y0(h_u_cla32_and4878_y0, h_u_cla32_and4877_y0, h_u_cla32_and4879_y0);
  and_gate and_gate_h_u_cla32_and4880_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4880_y0);
  and_gate and_gate_h_u_cla32_and4881_y0(h_u_cla32_and4880_y0, h_u_cla32_and4879_y0, h_u_cla32_and4881_y0);
  and_gate and_gate_h_u_cla32_and4882_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and4882_y0);
  and_gate and_gate_h_u_cla32_and4883_y0(h_u_cla32_and4882_y0, h_u_cla32_and4881_y0, h_u_cla32_and4883_y0);
  and_gate and_gate_h_u_cla32_and4884_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4884_y0);
  and_gate and_gate_h_u_cla32_and4885_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4885_y0);
  and_gate and_gate_h_u_cla32_and4886_y0(h_u_cla32_and4885_y0, h_u_cla32_and4884_y0, h_u_cla32_and4886_y0);
  and_gate and_gate_h_u_cla32_and4887_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4887_y0);
  and_gate and_gate_h_u_cla32_and4888_y0(h_u_cla32_and4887_y0, h_u_cla32_and4886_y0, h_u_cla32_and4888_y0);
  and_gate and_gate_h_u_cla32_and4889_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and4889_y0);
  and_gate and_gate_h_u_cla32_and4890_y0(h_u_cla32_and4889_y0, h_u_cla32_and4888_y0, h_u_cla32_and4890_y0);
  and_gate and_gate_h_u_cla32_and4891_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and4891_y0);
  and_gate and_gate_h_u_cla32_and4892_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and4892_y0);
  and_gate and_gate_h_u_cla32_and4893_y0(h_u_cla32_and4892_y0, h_u_cla32_and4891_y0, h_u_cla32_and4893_y0);
  and_gate and_gate_h_u_cla32_and4894_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and4894_y0);
  and_gate and_gate_h_u_cla32_and4895_y0(h_u_cla32_and4894_y0, h_u_cla32_and4893_y0, h_u_cla32_and4895_y0);
  and_gate and_gate_h_u_cla32_and4896_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and4896_y0);
  and_gate and_gate_h_u_cla32_and4897_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and4897_y0);
  and_gate and_gate_h_u_cla32_and4898_y0(h_u_cla32_and4897_y0, h_u_cla32_and4896_y0, h_u_cla32_and4898_y0);
  and_gate and_gate_h_u_cla32_and4899_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and4899_y0);
  or_gate or_gate_h_u_cla32_or276_y0(h_u_cla32_and4899_y0, h_u_cla32_and4370_y0, h_u_cla32_or276_y0);
  or_gate or_gate_h_u_cla32_or277_y0(h_u_cla32_or276_y0, h_u_cla32_and4415_y0, h_u_cla32_or277_y0);
  or_gate or_gate_h_u_cla32_or278_y0(h_u_cla32_or277_y0, h_u_cla32_and4458_y0, h_u_cla32_or278_y0);
  or_gate or_gate_h_u_cla32_or279_y0(h_u_cla32_or278_y0, h_u_cla32_and4499_y0, h_u_cla32_or279_y0);
  or_gate or_gate_h_u_cla32_or280_y0(h_u_cla32_or279_y0, h_u_cla32_and4538_y0, h_u_cla32_or280_y0);
  or_gate or_gate_h_u_cla32_or281_y0(h_u_cla32_or280_y0, h_u_cla32_and4575_y0, h_u_cla32_or281_y0);
  or_gate or_gate_h_u_cla32_or282_y0(h_u_cla32_or281_y0, h_u_cla32_and4610_y0, h_u_cla32_or282_y0);
  or_gate or_gate_h_u_cla32_or283_y0(h_u_cla32_or282_y0, h_u_cla32_and4643_y0, h_u_cla32_or283_y0);
  or_gate or_gate_h_u_cla32_or284_y0(h_u_cla32_or283_y0, h_u_cla32_and4674_y0, h_u_cla32_or284_y0);
  or_gate or_gate_h_u_cla32_or285_y0(h_u_cla32_or284_y0, h_u_cla32_and4703_y0, h_u_cla32_or285_y0);
  or_gate or_gate_h_u_cla32_or286_y0(h_u_cla32_or285_y0, h_u_cla32_and4730_y0, h_u_cla32_or286_y0);
  or_gate or_gate_h_u_cla32_or287_y0(h_u_cla32_or286_y0, h_u_cla32_and4755_y0, h_u_cla32_or287_y0);
  or_gate or_gate_h_u_cla32_or288_y0(h_u_cla32_or287_y0, h_u_cla32_and4778_y0, h_u_cla32_or288_y0);
  or_gate or_gate_h_u_cla32_or289_y0(h_u_cla32_or288_y0, h_u_cla32_and4799_y0, h_u_cla32_or289_y0);
  or_gate or_gate_h_u_cla32_or290_y0(h_u_cla32_or289_y0, h_u_cla32_and4818_y0, h_u_cla32_or290_y0);
  or_gate or_gate_h_u_cla32_or291_y0(h_u_cla32_or290_y0, h_u_cla32_and4835_y0, h_u_cla32_or291_y0);
  or_gate or_gate_h_u_cla32_or292_y0(h_u_cla32_or291_y0, h_u_cla32_and4850_y0, h_u_cla32_or292_y0);
  or_gate or_gate_h_u_cla32_or293_y0(h_u_cla32_or292_y0, h_u_cla32_and4863_y0, h_u_cla32_or293_y0);
  or_gate or_gate_h_u_cla32_or294_y0(h_u_cla32_or293_y0, h_u_cla32_and4874_y0, h_u_cla32_or294_y0);
  or_gate or_gate_h_u_cla32_or295_y0(h_u_cla32_or294_y0, h_u_cla32_and4883_y0, h_u_cla32_or295_y0);
  or_gate or_gate_h_u_cla32_or296_y0(h_u_cla32_or295_y0, h_u_cla32_and4890_y0, h_u_cla32_or296_y0);
  or_gate or_gate_h_u_cla32_or297_y0(h_u_cla32_or296_y0, h_u_cla32_and4895_y0, h_u_cla32_or297_y0);
  or_gate or_gate_h_u_cla32_or298_y0(h_u_cla32_or297_y0, h_u_cla32_and4898_y0, h_u_cla32_or298_y0);
  or_gate or_gate_h_u_cla32_or299_y0(h_u_cla32_pg_logic23_y1, h_u_cla32_or298_y0, h_u_cla32_or299_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic24_y0(a_24, b_24, h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_pg_logic24_y2);
  xor_gate xor_gate_h_u_cla32_xor24_y0(h_u_cla32_pg_logic24_y2, h_u_cla32_or299_y0, h_u_cla32_xor24_y0);
  and_gate and_gate_h_u_cla32_and4900_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and4900_y0);
  and_gate and_gate_h_u_cla32_and4901_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and4901_y0);
  and_gate and_gate_h_u_cla32_and4902_y0(h_u_cla32_and4901_y0, h_u_cla32_and4900_y0, h_u_cla32_and4902_y0);
  and_gate and_gate_h_u_cla32_and4903_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and4903_y0);
  and_gate and_gate_h_u_cla32_and4904_y0(h_u_cla32_and4903_y0, h_u_cla32_and4902_y0, h_u_cla32_and4904_y0);
  and_gate and_gate_h_u_cla32_and4905_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and4905_y0);
  and_gate and_gate_h_u_cla32_and4906_y0(h_u_cla32_and4905_y0, h_u_cla32_and4904_y0, h_u_cla32_and4906_y0);
  and_gate and_gate_h_u_cla32_and4907_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and4907_y0);
  and_gate and_gate_h_u_cla32_and4908_y0(h_u_cla32_and4907_y0, h_u_cla32_and4906_y0, h_u_cla32_and4908_y0);
  and_gate and_gate_h_u_cla32_and4909_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and4909_y0);
  and_gate and_gate_h_u_cla32_and4910_y0(h_u_cla32_and4909_y0, h_u_cla32_and4908_y0, h_u_cla32_and4910_y0);
  and_gate and_gate_h_u_cla32_and4911_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and4911_y0);
  and_gate and_gate_h_u_cla32_and4912_y0(h_u_cla32_and4911_y0, h_u_cla32_and4910_y0, h_u_cla32_and4912_y0);
  and_gate and_gate_h_u_cla32_and4913_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and4913_y0);
  and_gate and_gate_h_u_cla32_and4914_y0(h_u_cla32_and4913_y0, h_u_cla32_and4912_y0, h_u_cla32_and4914_y0);
  and_gate and_gate_h_u_cla32_and4915_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and4915_y0);
  and_gate and_gate_h_u_cla32_and4916_y0(h_u_cla32_and4915_y0, h_u_cla32_and4914_y0, h_u_cla32_and4916_y0);
  and_gate and_gate_h_u_cla32_and4917_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and4917_y0);
  and_gate and_gate_h_u_cla32_and4918_y0(h_u_cla32_and4917_y0, h_u_cla32_and4916_y0, h_u_cla32_and4918_y0);
  and_gate and_gate_h_u_cla32_and4919_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and4919_y0);
  and_gate and_gate_h_u_cla32_and4920_y0(h_u_cla32_and4919_y0, h_u_cla32_and4918_y0, h_u_cla32_and4920_y0);
  and_gate and_gate_h_u_cla32_and4921_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and4921_y0);
  and_gate and_gate_h_u_cla32_and4922_y0(h_u_cla32_and4921_y0, h_u_cla32_and4920_y0, h_u_cla32_and4922_y0);
  and_gate and_gate_h_u_cla32_and4923_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and4923_y0);
  and_gate and_gate_h_u_cla32_and4924_y0(h_u_cla32_and4923_y0, h_u_cla32_and4922_y0, h_u_cla32_and4924_y0);
  and_gate and_gate_h_u_cla32_and4925_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and4925_y0);
  and_gate and_gate_h_u_cla32_and4926_y0(h_u_cla32_and4925_y0, h_u_cla32_and4924_y0, h_u_cla32_and4926_y0);
  and_gate and_gate_h_u_cla32_and4927_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and4927_y0);
  and_gate and_gate_h_u_cla32_and4928_y0(h_u_cla32_and4927_y0, h_u_cla32_and4926_y0, h_u_cla32_and4928_y0);
  and_gate and_gate_h_u_cla32_and4929_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and4929_y0);
  and_gate and_gate_h_u_cla32_and4930_y0(h_u_cla32_and4929_y0, h_u_cla32_and4928_y0, h_u_cla32_and4930_y0);
  and_gate and_gate_h_u_cla32_and4931_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and4931_y0);
  and_gate and_gate_h_u_cla32_and4932_y0(h_u_cla32_and4931_y0, h_u_cla32_and4930_y0, h_u_cla32_and4932_y0);
  and_gate and_gate_h_u_cla32_and4933_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and4933_y0);
  and_gate and_gate_h_u_cla32_and4934_y0(h_u_cla32_and4933_y0, h_u_cla32_and4932_y0, h_u_cla32_and4934_y0);
  and_gate and_gate_h_u_cla32_and4935_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and4935_y0);
  and_gate and_gate_h_u_cla32_and4936_y0(h_u_cla32_and4935_y0, h_u_cla32_and4934_y0, h_u_cla32_and4936_y0);
  and_gate and_gate_h_u_cla32_and4937_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and4937_y0);
  and_gate and_gate_h_u_cla32_and4938_y0(h_u_cla32_and4937_y0, h_u_cla32_and4936_y0, h_u_cla32_and4938_y0);
  and_gate and_gate_h_u_cla32_and4939_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and4939_y0);
  and_gate and_gate_h_u_cla32_and4940_y0(h_u_cla32_and4939_y0, h_u_cla32_and4938_y0, h_u_cla32_and4940_y0);
  and_gate and_gate_h_u_cla32_and4941_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and4941_y0);
  and_gate and_gate_h_u_cla32_and4942_y0(h_u_cla32_and4941_y0, h_u_cla32_and4940_y0, h_u_cla32_and4942_y0);
  and_gate and_gate_h_u_cla32_and4943_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and4943_y0);
  and_gate and_gate_h_u_cla32_and4944_y0(h_u_cla32_and4943_y0, h_u_cla32_and4942_y0, h_u_cla32_and4944_y0);
  and_gate and_gate_h_u_cla32_and4945_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and4945_y0);
  and_gate and_gate_h_u_cla32_and4946_y0(h_u_cla32_and4945_y0, h_u_cla32_and4944_y0, h_u_cla32_and4946_y0);
  and_gate and_gate_h_u_cla32_and4947_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and4947_y0);
  and_gate and_gate_h_u_cla32_and4948_y0(h_u_cla32_and4947_y0, h_u_cla32_and4946_y0, h_u_cla32_and4948_y0);
  and_gate and_gate_h_u_cla32_and4949_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4949_y0);
  and_gate and_gate_h_u_cla32_and4950_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4950_y0);
  and_gate and_gate_h_u_cla32_and4951_y0(h_u_cla32_and4950_y0, h_u_cla32_and4949_y0, h_u_cla32_and4951_y0);
  and_gate and_gate_h_u_cla32_and4952_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4952_y0);
  and_gate and_gate_h_u_cla32_and4953_y0(h_u_cla32_and4952_y0, h_u_cla32_and4951_y0, h_u_cla32_and4953_y0);
  and_gate and_gate_h_u_cla32_and4954_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4954_y0);
  and_gate and_gate_h_u_cla32_and4955_y0(h_u_cla32_and4954_y0, h_u_cla32_and4953_y0, h_u_cla32_and4955_y0);
  and_gate and_gate_h_u_cla32_and4956_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4956_y0);
  and_gate and_gate_h_u_cla32_and4957_y0(h_u_cla32_and4956_y0, h_u_cla32_and4955_y0, h_u_cla32_and4957_y0);
  and_gate and_gate_h_u_cla32_and4958_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4958_y0);
  and_gate and_gate_h_u_cla32_and4959_y0(h_u_cla32_and4958_y0, h_u_cla32_and4957_y0, h_u_cla32_and4959_y0);
  and_gate and_gate_h_u_cla32_and4960_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4960_y0);
  and_gate and_gate_h_u_cla32_and4961_y0(h_u_cla32_and4960_y0, h_u_cla32_and4959_y0, h_u_cla32_and4961_y0);
  and_gate and_gate_h_u_cla32_and4962_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4962_y0);
  and_gate and_gate_h_u_cla32_and4963_y0(h_u_cla32_and4962_y0, h_u_cla32_and4961_y0, h_u_cla32_and4963_y0);
  and_gate and_gate_h_u_cla32_and4964_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4964_y0);
  and_gate and_gate_h_u_cla32_and4965_y0(h_u_cla32_and4964_y0, h_u_cla32_and4963_y0, h_u_cla32_and4965_y0);
  and_gate and_gate_h_u_cla32_and4966_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4966_y0);
  and_gate and_gate_h_u_cla32_and4967_y0(h_u_cla32_and4966_y0, h_u_cla32_and4965_y0, h_u_cla32_and4967_y0);
  and_gate and_gate_h_u_cla32_and4968_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4968_y0);
  and_gate and_gate_h_u_cla32_and4969_y0(h_u_cla32_and4968_y0, h_u_cla32_and4967_y0, h_u_cla32_and4969_y0);
  and_gate and_gate_h_u_cla32_and4970_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4970_y0);
  and_gate and_gate_h_u_cla32_and4971_y0(h_u_cla32_and4970_y0, h_u_cla32_and4969_y0, h_u_cla32_and4971_y0);
  and_gate and_gate_h_u_cla32_and4972_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4972_y0);
  and_gate and_gate_h_u_cla32_and4973_y0(h_u_cla32_and4972_y0, h_u_cla32_and4971_y0, h_u_cla32_and4973_y0);
  and_gate and_gate_h_u_cla32_and4974_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4974_y0);
  and_gate and_gate_h_u_cla32_and4975_y0(h_u_cla32_and4974_y0, h_u_cla32_and4973_y0, h_u_cla32_and4975_y0);
  and_gate and_gate_h_u_cla32_and4976_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4976_y0);
  and_gate and_gate_h_u_cla32_and4977_y0(h_u_cla32_and4976_y0, h_u_cla32_and4975_y0, h_u_cla32_and4977_y0);
  and_gate and_gate_h_u_cla32_and4978_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4978_y0);
  and_gate and_gate_h_u_cla32_and4979_y0(h_u_cla32_and4978_y0, h_u_cla32_and4977_y0, h_u_cla32_and4979_y0);
  and_gate and_gate_h_u_cla32_and4980_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4980_y0);
  and_gate and_gate_h_u_cla32_and4981_y0(h_u_cla32_and4980_y0, h_u_cla32_and4979_y0, h_u_cla32_and4981_y0);
  and_gate and_gate_h_u_cla32_and4982_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4982_y0);
  and_gate and_gate_h_u_cla32_and4983_y0(h_u_cla32_and4982_y0, h_u_cla32_and4981_y0, h_u_cla32_and4983_y0);
  and_gate and_gate_h_u_cla32_and4984_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4984_y0);
  and_gate and_gate_h_u_cla32_and4985_y0(h_u_cla32_and4984_y0, h_u_cla32_and4983_y0, h_u_cla32_and4985_y0);
  and_gate and_gate_h_u_cla32_and4986_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4986_y0);
  and_gate and_gate_h_u_cla32_and4987_y0(h_u_cla32_and4986_y0, h_u_cla32_and4985_y0, h_u_cla32_and4987_y0);
  and_gate and_gate_h_u_cla32_and4988_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4988_y0);
  and_gate and_gate_h_u_cla32_and4989_y0(h_u_cla32_and4988_y0, h_u_cla32_and4987_y0, h_u_cla32_and4989_y0);
  and_gate and_gate_h_u_cla32_and4990_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4990_y0);
  and_gate and_gate_h_u_cla32_and4991_y0(h_u_cla32_and4990_y0, h_u_cla32_and4989_y0, h_u_cla32_and4991_y0);
  and_gate and_gate_h_u_cla32_and4992_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4992_y0);
  and_gate and_gate_h_u_cla32_and4993_y0(h_u_cla32_and4992_y0, h_u_cla32_and4991_y0, h_u_cla32_and4993_y0);
  and_gate and_gate_h_u_cla32_and4994_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and4994_y0);
  and_gate and_gate_h_u_cla32_and4995_y0(h_u_cla32_and4994_y0, h_u_cla32_and4993_y0, h_u_cla32_and4995_y0);
  and_gate and_gate_h_u_cla32_and4996_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4996_y0);
  and_gate and_gate_h_u_cla32_and4997_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4997_y0);
  and_gate and_gate_h_u_cla32_and4998_y0(h_u_cla32_and4997_y0, h_u_cla32_and4996_y0, h_u_cla32_and4998_y0);
  and_gate and_gate_h_u_cla32_and4999_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and4999_y0);
  and_gate and_gate_h_u_cla32_and5000_y0(h_u_cla32_and4999_y0, h_u_cla32_and4998_y0, h_u_cla32_and5000_y0);
  and_gate and_gate_h_u_cla32_and5001_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5001_y0);
  and_gate and_gate_h_u_cla32_and5002_y0(h_u_cla32_and5001_y0, h_u_cla32_and5000_y0, h_u_cla32_and5002_y0);
  and_gate and_gate_h_u_cla32_and5003_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5003_y0);
  and_gate and_gate_h_u_cla32_and5004_y0(h_u_cla32_and5003_y0, h_u_cla32_and5002_y0, h_u_cla32_and5004_y0);
  and_gate and_gate_h_u_cla32_and5005_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5005_y0);
  and_gate and_gate_h_u_cla32_and5006_y0(h_u_cla32_and5005_y0, h_u_cla32_and5004_y0, h_u_cla32_and5006_y0);
  and_gate and_gate_h_u_cla32_and5007_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5007_y0);
  and_gate and_gate_h_u_cla32_and5008_y0(h_u_cla32_and5007_y0, h_u_cla32_and5006_y0, h_u_cla32_and5008_y0);
  and_gate and_gate_h_u_cla32_and5009_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5009_y0);
  and_gate and_gate_h_u_cla32_and5010_y0(h_u_cla32_and5009_y0, h_u_cla32_and5008_y0, h_u_cla32_and5010_y0);
  and_gate and_gate_h_u_cla32_and5011_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5011_y0);
  and_gate and_gate_h_u_cla32_and5012_y0(h_u_cla32_and5011_y0, h_u_cla32_and5010_y0, h_u_cla32_and5012_y0);
  and_gate and_gate_h_u_cla32_and5013_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5013_y0);
  and_gate and_gate_h_u_cla32_and5014_y0(h_u_cla32_and5013_y0, h_u_cla32_and5012_y0, h_u_cla32_and5014_y0);
  and_gate and_gate_h_u_cla32_and5015_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5015_y0);
  and_gate and_gate_h_u_cla32_and5016_y0(h_u_cla32_and5015_y0, h_u_cla32_and5014_y0, h_u_cla32_and5016_y0);
  and_gate and_gate_h_u_cla32_and5017_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5017_y0);
  and_gate and_gate_h_u_cla32_and5018_y0(h_u_cla32_and5017_y0, h_u_cla32_and5016_y0, h_u_cla32_and5018_y0);
  and_gate and_gate_h_u_cla32_and5019_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5019_y0);
  and_gate and_gate_h_u_cla32_and5020_y0(h_u_cla32_and5019_y0, h_u_cla32_and5018_y0, h_u_cla32_and5020_y0);
  and_gate and_gate_h_u_cla32_and5021_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5021_y0);
  and_gate and_gate_h_u_cla32_and5022_y0(h_u_cla32_and5021_y0, h_u_cla32_and5020_y0, h_u_cla32_and5022_y0);
  and_gate and_gate_h_u_cla32_and5023_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5023_y0);
  and_gate and_gate_h_u_cla32_and5024_y0(h_u_cla32_and5023_y0, h_u_cla32_and5022_y0, h_u_cla32_and5024_y0);
  and_gate and_gate_h_u_cla32_and5025_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5025_y0);
  and_gate and_gate_h_u_cla32_and5026_y0(h_u_cla32_and5025_y0, h_u_cla32_and5024_y0, h_u_cla32_and5026_y0);
  and_gate and_gate_h_u_cla32_and5027_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5027_y0);
  and_gate and_gate_h_u_cla32_and5028_y0(h_u_cla32_and5027_y0, h_u_cla32_and5026_y0, h_u_cla32_and5028_y0);
  and_gate and_gate_h_u_cla32_and5029_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5029_y0);
  and_gate and_gate_h_u_cla32_and5030_y0(h_u_cla32_and5029_y0, h_u_cla32_and5028_y0, h_u_cla32_and5030_y0);
  and_gate and_gate_h_u_cla32_and5031_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5031_y0);
  and_gate and_gate_h_u_cla32_and5032_y0(h_u_cla32_and5031_y0, h_u_cla32_and5030_y0, h_u_cla32_and5032_y0);
  and_gate and_gate_h_u_cla32_and5033_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5033_y0);
  and_gate and_gate_h_u_cla32_and5034_y0(h_u_cla32_and5033_y0, h_u_cla32_and5032_y0, h_u_cla32_and5034_y0);
  and_gate and_gate_h_u_cla32_and5035_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5035_y0);
  and_gate and_gate_h_u_cla32_and5036_y0(h_u_cla32_and5035_y0, h_u_cla32_and5034_y0, h_u_cla32_and5036_y0);
  and_gate and_gate_h_u_cla32_and5037_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5037_y0);
  and_gate and_gate_h_u_cla32_and5038_y0(h_u_cla32_and5037_y0, h_u_cla32_and5036_y0, h_u_cla32_and5038_y0);
  and_gate and_gate_h_u_cla32_and5039_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5039_y0);
  and_gate and_gate_h_u_cla32_and5040_y0(h_u_cla32_and5039_y0, h_u_cla32_and5038_y0, h_u_cla32_and5040_y0);
  and_gate and_gate_h_u_cla32_and5041_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5041_y0);
  and_gate and_gate_h_u_cla32_and5042_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5042_y0);
  and_gate and_gate_h_u_cla32_and5043_y0(h_u_cla32_and5042_y0, h_u_cla32_and5041_y0, h_u_cla32_and5043_y0);
  and_gate and_gate_h_u_cla32_and5044_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5044_y0);
  and_gate and_gate_h_u_cla32_and5045_y0(h_u_cla32_and5044_y0, h_u_cla32_and5043_y0, h_u_cla32_and5045_y0);
  and_gate and_gate_h_u_cla32_and5046_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5046_y0);
  and_gate and_gate_h_u_cla32_and5047_y0(h_u_cla32_and5046_y0, h_u_cla32_and5045_y0, h_u_cla32_and5047_y0);
  and_gate and_gate_h_u_cla32_and5048_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5048_y0);
  and_gate and_gate_h_u_cla32_and5049_y0(h_u_cla32_and5048_y0, h_u_cla32_and5047_y0, h_u_cla32_and5049_y0);
  and_gate and_gate_h_u_cla32_and5050_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5050_y0);
  and_gate and_gate_h_u_cla32_and5051_y0(h_u_cla32_and5050_y0, h_u_cla32_and5049_y0, h_u_cla32_and5051_y0);
  and_gate and_gate_h_u_cla32_and5052_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5052_y0);
  and_gate and_gate_h_u_cla32_and5053_y0(h_u_cla32_and5052_y0, h_u_cla32_and5051_y0, h_u_cla32_and5053_y0);
  and_gate and_gate_h_u_cla32_and5054_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5054_y0);
  and_gate and_gate_h_u_cla32_and5055_y0(h_u_cla32_and5054_y0, h_u_cla32_and5053_y0, h_u_cla32_and5055_y0);
  and_gate and_gate_h_u_cla32_and5056_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5056_y0);
  and_gate and_gate_h_u_cla32_and5057_y0(h_u_cla32_and5056_y0, h_u_cla32_and5055_y0, h_u_cla32_and5057_y0);
  and_gate and_gate_h_u_cla32_and5058_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5058_y0);
  and_gate and_gate_h_u_cla32_and5059_y0(h_u_cla32_and5058_y0, h_u_cla32_and5057_y0, h_u_cla32_and5059_y0);
  and_gate and_gate_h_u_cla32_and5060_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5060_y0);
  and_gate and_gate_h_u_cla32_and5061_y0(h_u_cla32_and5060_y0, h_u_cla32_and5059_y0, h_u_cla32_and5061_y0);
  and_gate and_gate_h_u_cla32_and5062_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5062_y0);
  and_gate and_gate_h_u_cla32_and5063_y0(h_u_cla32_and5062_y0, h_u_cla32_and5061_y0, h_u_cla32_and5063_y0);
  and_gate and_gate_h_u_cla32_and5064_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5064_y0);
  and_gate and_gate_h_u_cla32_and5065_y0(h_u_cla32_and5064_y0, h_u_cla32_and5063_y0, h_u_cla32_and5065_y0);
  and_gate and_gate_h_u_cla32_and5066_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5066_y0);
  and_gate and_gate_h_u_cla32_and5067_y0(h_u_cla32_and5066_y0, h_u_cla32_and5065_y0, h_u_cla32_and5067_y0);
  and_gate and_gate_h_u_cla32_and5068_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5068_y0);
  and_gate and_gate_h_u_cla32_and5069_y0(h_u_cla32_and5068_y0, h_u_cla32_and5067_y0, h_u_cla32_and5069_y0);
  and_gate and_gate_h_u_cla32_and5070_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5070_y0);
  and_gate and_gate_h_u_cla32_and5071_y0(h_u_cla32_and5070_y0, h_u_cla32_and5069_y0, h_u_cla32_and5071_y0);
  and_gate and_gate_h_u_cla32_and5072_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5072_y0);
  and_gate and_gate_h_u_cla32_and5073_y0(h_u_cla32_and5072_y0, h_u_cla32_and5071_y0, h_u_cla32_and5073_y0);
  and_gate and_gate_h_u_cla32_and5074_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5074_y0);
  and_gate and_gate_h_u_cla32_and5075_y0(h_u_cla32_and5074_y0, h_u_cla32_and5073_y0, h_u_cla32_and5075_y0);
  and_gate and_gate_h_u_cla32_and5076_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5076_y0);
  and_gate and_gate_h_u_cla32_and5077_y0(h_u_cla32_and5076_y0, h_u_cla32_and5075_y0, h_u_cla32_and5077_y0);
  and_gate and_gate_h_u_cla32_and5078_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5078_y0);
  and_gate and_gate_h_u_cla32_and5079_y0(h_u_cla32_and5078_y0, h_u_cla32_and5077_y0, h_u_cla32_and5079_y0);
  and_gate and_gate_h_u_cla32_and5080_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5080_y0);
  and_gate and_gate_h_u_cla32_and5081_y0(h_u_cla32_and5080_y0, h_u_cla32_and5079_y0, h_u_cla32_and5081_y0);
  and_gate and_gate_h_u_cla32_and5082_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5082_y0);
  and_gate and_gate_h_u_cla32_and5083_y0(h_u_cla32_and5082_y0, h_u_cla32_and5081_y0, h_u_cla32_and5083_y0);
  and_gate and_gate_h_u_cla32_and5084_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5084_y0);
  and_gate and_gate_h_u_cla32_and5085_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5085_y0);
  and_gate and_gate_h_u_cla32_and5086_y0(h_u_cla32_and5085_y0, h_u_cla32_and5084_y0, h_u_cla32_and5086_y0);
  and_gate and_gate_h_u_cla32_and5087_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5087_y0);
  and_gate and_gate_h_u_cla32_and5088_y0(h_u_cla32_and5087_y0, h_u_cla32_and5086_y0, h_u_cla32_and5088_y0);
  and_gate and_gate_h_u_cla32_and5089_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5089_y0);
  and_gate and_gate_h_u_cla32_and5090_y0(h_u_cla32_and5089_y0, h_u_cla32_and5088_y0, h_u_cla32_and5090_y0);
  and_gate and_gate_h_u_cla32_and5091_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5091_y0);
  and_gate and_gate_h_u_cla32_and5092_y0(h_u_cla32_and5091_y0, h_u_cla32_and5090_y0, h_u_cla32_and5092_y0);
  and_gate and_gate_h_u_cla32_and5093_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5093_y0);
  and_gate and_gate_h_u_cla32_and5094_y0(h_u_cla32_and5093_y0, h_u_cla32_and5092_y0, h_u_cla32_and5094_y0);
  and_gate and_gate_h_u_cla32_and5095_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5095_y0);
  and_gate and_gate_h_u_cla32_and5096_y0(h_u_cla32_and5095_y0, h_u_cla32_and5094_y0, h_u_cla32_and5096_y0);
  and_gate and_gate_h_u_cla32_and5097_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5097_y0);
  and_gate and_gate_h_u_cla32_and5098_y0(h_u_cla32_and5097_y0, h_u_cla32_and5096_y0, h_u_cla32_and5098_y0);
  and_gate and_gate_h_u_cla32_and5099_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5099_y0);
  and_gate and_gate_h_u_cla32_and5100_y0(h_u_cla32_and5099_y0, h_u_cla32_and5098_y0, h_u_cla32_and5100_y0);
  and_gate and_gate_h_u_cla32_and5101_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5101_y0);
  and_gate and_gate_h_u_cla32_and5102_y0(h_u_cla32_and5101_y0, h_u_cla32_and5100_y0, h_u_cla32_and5102_y0);
  and_gate and_gate_h_u_cla32_and5103_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5103_y0);
  and_gate and_gate_h_u_cla32_and5104_y0(h_u_cla32_and5103_y0, h_u_cla32_and5102_y0, h_u_cla32_and5104_y0);
  and_gate and_gate_h_u_cla32_and5105_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5105_y0);
  and_gate and_gate_h_u_cla32_and5106_y0(h_u_cla32_and5105_y0, h_u_cla32_and5104_y0, h_u_cla32_and5106_y0);
  and_gate and_gate_h_u_cla32_and5107_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5107_y0);
  and_gate and_gate_h_u_cla32_and5108_y0(h_u_cla32_and5107_y0, h_u_cla32_and5106_y0, h_u_cla32_and5108_y0);
  and_gate and_gate_h_u_cla32_and5109_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5109_y0);
  and_gate and_gate_h_u_cla32_and5110_y0(h_u_cla32_and5109_y0, h_u_cla32_and5108_y0, h_u_cla32_and5110_y0);
  and_gate and_gate_h_u_cla32_and5111_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5111_y0);
  and_gate and_gate_h_u_cla32_and5112_y0(h_u_cla32_and5111_y0, h_u_cla32_and5110_y0, h_u_cla32_and5112_y0);
  and_gate and_gate_h_u_cla32_and5113_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5113_y0);
  and_gate and_gate_h_u_cla32_and5114_y0(h_u_cla32_and5113_y0, h_u_cla32_and5112_y0, h_u_cla32_and5114_y0);
  and_gate and_gate_h_u_cla32_and5115_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5115_y0);
  and_gate and_gate_h_u_cla32_and5116_y0(h_u_cla32_and5115_y0, h_u_cla32_and5114_y0, h_u_cla32_and5116_y0);
  and_gate and_gate_h_u_cla32_and5117_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5117_y0);
  and_gate and_gate_h_u_cla32_and5118_y0(h_u_cla32_and5117_y0, h_u_cla32_and5116_y0, h_u_cla32_and5118_y0);
  and_gate and_gate_h_u_cla32_and5119_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5119_y0);
  and_gate and_gate_h_u_cla32_and5120_y0(h_u_cla32_and5119_y0, h_u_cla32_and5118_y0, h_u_cla32_and5120_y0);
  and_gate and_gate_h_u_cla32_and5121_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5121_y0);
  and_gate and_gate_h_u_cla32_and5122_y0(h_u_cla32_and5121_y0, h_u_cla32_and5120_y0, h_u_cla32_and5122_y0);
  and_gate and_gate_h_u_cla32_and5123_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5123_y0);
  and_gate and_gate_h_u_cla32_and5124_y0(h_u_cla32_and5123_y0, h_u_cla32_and5122_y0, h_u_cla32_and5124_y0);
  and_gate and_gate_h_u_cla32_and5125_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5125_y0);
  and_gate and_gate_h_u_cla32_and5126_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5126_y0);
  and_gate and_gate_h_u_cla32_and5127_y0(h_u_cla32_and5126_y0, h_u_cla32_and5125_y0, h_u_cla32_and5127_y0);
  and_gate and_gate_h_u_cla32_and5128_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5128_y0);
  and_gate and_gate_h_u_cla32_and5129_y0(h_u_cla32_and5128_y0, h_u_cla32_and5127_y0, h_u_cla32_and5129_y0);
  and_gate and_gate_h_u_cla32_and5130_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5130_y0);
  and_gate and_gate_h_u_cla32_and5131_y0(h_u_cla32_and5130_y0, h_u_cla32_and5129_y0, h_u_cla32_and5131_y0);
  and_gate and_gate_h_u_cla32_and5132_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5132_y0);
  and_gate and_gate_h_u_cla32_and5133_y0(h_u_cla32_and5132_y0, h_u_cla32_and5131_y0, h_u_cla32_and5133_y0);
  and_gate and_gate_h_u_cla32_and5134_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5134_y0);
  and_gate and_gate_h_u_cla32_and5135_y0(h_u_cla32_and5134_y0, h_u_cla32_and5133_y0, h_u_cla32_and5135_y0);
  and_gate and_gate_h_u_cla32_and5136_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5136_y0);
  and_gate and_gate_h_u_cla32_and5137_y0(h_u_cla32_and5136_y0, h_u_cla32_and5135_y0, h_u_cla32_and5137_y0);
  and_gate and_gate_h_u_cla32_and5138_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5138_y0);
  and_gate and_gate_h_u_cla32_and5139_y0(h_u_cla32_and5138_y0, h_u_cla32_and5137_y0, h_u_cla32_and5139_y0);
  and_gate and_gate_h_u_cla32_and5140_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5140_y0);
  and_gate and_gate_h_u_cla32_and5141_y0(h_u_cla32_and5140_y0, h_u_cla32_and5139_y0, h_u_cla32_and5141_y0);
  and_gate and_gate_h_u_cla32_and5142_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5142_y0);
  and_gate and_gate_h_u_cla32_and5143_y0(h_u_cla32_and5142_y0, h_u_cla32_and5141_y0, h_u_cla32_and5143_y0);
  and_gate and_gate_h_u_cla32_and5144_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5144_y0);
  and_gate and_gate_h_u_cla32_and5145_y0(h_u_cla32_and5144_y0, h_u_cla32_and5143_y0, h_u_cla32_and5145_y0);
  and_gate and_gate_h_u_cla32_and5146_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5146_y0);
  and_gate and_gate_h_u_cla32_and5147_y0(h_u_cla32_and5146_y0, h_u_cla32_and5145_y0, h_u_cla32_and5147_y0);
  and_gate and_gate_h_u_cla32_and5148_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5148_y0);
  and_gate and_gate_h_u_cla32_and5149_y0(h_u_cla32_and5148_y0, h_u_cla32_and5147_y0, h_u_cla32_and5149_y0);
  and_gate and_gate_h_u_cla32_and5150_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5150_y0);
  and_gate and_gate_h_u_cla32_and5151_y0(h_u_cla32_and5150_y0, h_u_cla32_and5149_y0, h_u_cla32_and5151_y0);
  and_gate and_gate_h_u_cla32_and5152_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5152_y0);
  and_gate and_gate_h_u_cla32_and5153_y0(h_u_cla32_and5152_y0, h_u_cla32_and5151_y0, h_u_cla32_and5153_y0);
  and_gate and_gate_h_u_cla32_and5154_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5154_y0);
  and_gate and_gate_h_u_cla32_and5155_y0(h_u_cla32_and5154_y0, h_u_cla32_and5153_y0, h_u_cla32_and5155_y0);
  and_gate and_gate_h_u_cla32_and5156_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5156_y0);
  and_gate and_gate_h_u_cla32_and5157_y0(h_u_cla32_and5156_y0, h_u_cla32_and5155_y0, h_u_cla32_and5157_y0);
  and_gate and_gate_h_u_cla32_and5158_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5158_y0);
  and_gate and_gate_h_u_cla32_and5159_y0(h_u_cla32_and5158_y0, h_u_cla32_and5157_y0, h_u_cla32_and5159_y0);
  and_gate and_gate_h_u_cla32_and5160_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5160_y0);
  and_gate and_gate_h_u_cla32_and5161_y0(h_u_cla32_and5160_y0, h_u_cla32_and5159_y0, h_u_cla32_and5161_y0);
  and_gate and_gate_h_u_cla32_and5162_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5162_y0);
  and_gate and_gate_h_u_cla32_and5163_y0(h_u_cla32_and5162_y0, h_u_cla32_and5161_y0, h_u_cla32_and5163_y0);
  and_gate and_gate_h_u_cla32_and5164_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5164_y0);
  and_gate and_gate_h_u_cla32_and5165_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5165_y0);
  and_gate and_gate_h_u_cla32_and5166_y0(h_u_cla32_and5165_y0, h_u_cla32_and5164_y0, h_u_cla32_and5166_y0);
  and_gate and_gate_h_u_cla32_and5167_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5167_y0);
  and_gate and_gate_h_u_cla32_and5168_y0(h_u_cla32_and5167_y0, h_u_cla32_and5166_y0, h_u_cla32_and5168_y0);
  and_gate and_gate_h_u_cla32_and5169_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5169_y0);
  and_gate and_gate_h_u_cla32_and5170_y0(h_u_cla32_and5169_y0, h_u_cla32_and5168_y0, h_u_cla32_and5170_y0);
  and_gate and_gate_h_u_cla32_and5171_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5171_y0);
  and_gate and_gate_h_u_cla32_and5172_y0(h_u_cla32_and5171_y0, h_u_cla32_and5170_y0, h_u_cla32_and5172_y0);
  and_gate and_gate_h_u_cla32_and5173_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5173_y0);
  and_gate and_gate_h_u_cla32_and5174_y0(h_u_cla32_and5173_y0, h_u_cla32_and5172_y0, h_u_cla32_and5174_y0);
  and_gate and_gate_h_u_cla32_and5175_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5175_y0);
  and_gate and_gate_h_u_cla32_and5176_y0(h_u_cla32_and5175_y0, h_u_cla32_and5174_y0, h_u_cla32_and5176_y0);
  and_gate and_gate_h_u_cla32_and5177_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5177_y0);
  and_gate and_gate_h_u_cla32_and5178_y0(h_u_cla32_and5177_y0, h_u_cla32_and5176_y0, h_u_cla32_and5178_y0);
  and_gate and_gate_h_u_cla32_and5179_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5179_y0);
  and_gate and_gate_h_u_cla32_and5180_y0(h_u_cla32_and5179_y0, h_u_cla32_and5178_y0, h_u_cla32_and5180_y0);
  and_gate and_gate_h_u_cla32_and5181_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5181_y0);
  and_gate and_gate_h_u_cla32_and5182_y0(h_u_cla32_and5181_y0, h_u_cla32_and5180_y0, h_u_cla32_and5182_y0);
  and_gate and_gate_h_u_cla32_and5183_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5183_y0);
  and_gate and_gate_h_u_cla32_and5184_y0(h_u_cla32_and5183_y0, h_u_cla32_and5182_y0, h_u_cla32_and5184_y0);
  and_gate and_gate_h_u_cla32_and5185_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5185_y0);
  and_gate and_gate_h_u_cla32_and5186_y0(h_u_cla32_and5185_y0, h_u_cla32_and5184_y0, h_u_cla32_and5186_y0);
  and_gate and_gate_h_u_cla32_and5187_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5187_y0);
  and_gate and_gate_h_u_cla32_and5188_y0(h_u_cla32_and5187_y0, h_u_cla32_and5186_y0, h_u_cla32_and5188_y0);
  and_gate and_gate_h_u_cla32_and5189_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5189_y0);
  and_gate and_gate_h_u_cla32_and5190_y0(h_u_cla32_and5189_y0, h_u_cla32_and5188_y0, h_u_cla32_and5190_y0);
  and_gate and_gate_h_u_cla32_and5191_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5191_y0);
  and_gate and_gate_h_u_cla32_and5192_y0(h_u_cla32_and5191_y0, h_u_cla32_and5190_y0, h_u_cla32_and5192_y0);
  and_gate and_gate_h_u_cla32_and5193_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5193_y0);
  and_gate and_gate_h_u_cla32_and5194_y0(h_u_cla32_and5193_y0, h_u_cla32_and5192_y0, h_u_cla32_and5194_y0);
  and_gate and_gate_h_u_cla32_and5195_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5195_y0);
  and_gate and_gate_h_u_cla32_and5196_y0(h_u_cla32_and5195_y0, h_u_cla32_and5194_y0, h_u_cla32_and5196_y0);
  and_gate and_gate_h_u_cla32_and5197_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5197_y0);
  and_gate and_gate_h_u_cla32_and5198_y0(h_u_cla32_and5197_y0, h_u_cla32_and5196_y0, h_u_cla32_and5198_y0);
  and_gate and_gate_h_u_cla32_and5199_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5199_y0);
  and_gate and_gate_h_u_cla32_and5200_y0(h_u_cla32_and5199_y0, h_u_cla32_and5198_y0, h_u_cla32_and5200_y0);
  and_gate and_gate_h_u_cla32_and5201_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5201_y0);
  and_gate and_gate_h_u_cla32_and5202_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5202_y0);
  and_gate and_gate_h_u_cla32_and5203_y0(h_u_cla32_and5202_y0, h_u_cla32_and5201_y0, h_u_cla32_and5203_y0);
  and_gate and_gate_h_u_cla32_and5204_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5204_y0);
  and_gate and_gate_h_u_cla32_and5205_y0(h_u_cla32_and5204_y0, h_u_cla32_and5203_y0, h_u_cla32_and5205_y0);
  and_gate and_gate_h_u_cla32_and5206_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5206_y0);
  and_gate and_gate_h_u_cla32_and5207_y0(h_u_cla32_and5206_y0, h_u_cla32_and5205_y0, h_u_cla32_and5207_y0);
  and_gate and_gate_h_u_cla32_and5208_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5208_y0);
  and_gate and_gate_h_u_cla32_and5209_y0(h_u_cla32_and5208_y0, h_u_cla32_and5207_y0, h_u_cla32_and5209_y0);
  and_gate and_gate_h_u_cla32_and5210_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5210_y0);
  and_gate and_gate_h_u_cla32_and5211_y0(h_u_cla32_and5210_y0, h_u_cla32_and5209_y0, h_u_cla32_and5211_y0);
  and_gate and_gate_h_u_cla32_and5212_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5212_y0);
  and_gate and_gate_h_u_cla32_and5213_y0(h_u_cla32_and5212_y0, h_u_cla32_and5211_y0, h_u_cla32_and5213_y0);
  and_gate and_gate_h_u_cla32_and5214_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5214_y0);
  and_gate and_gate_h_u_cla32_and5215_y0(h_u_cla32_and5214_y0, h_u_cla32_and5213_y0, h_u_cla32_and5215_y0);
  and_gate and_gate_h_u_cla32_and5216_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5216_y0);
  and_gate and_gate_h_u_cla32_and5217_y0(h_u_cla32_and5216_y0, h_u_cla32_and5215_y0, h_u_cla32_and5217_y0);
  and_gate and_gate_h_u_cla32_and5218_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5218_y0);
  and_gate and_gate_h_u_cla32_and5219_y0(h_u_cla32_and5218_y0, h_u_cla32_and5217_y0, h_u_cla32_and5219_y0);
  and_gate and_gate_h_u_cla32_and5220_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5220_y0);
  and_gate and_gate_h_u_cla32_and5221_y0(h_u_cla32_and5220_y0, h_u_cla32_and5219_y0, h_u_cla32_and5221_y0);
  and_gate and_gate_h_u_cla32_and5222_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5222_y0);
  and_gate and_gate_h_u_cla32_and5223_y0(h_u_cla32_and5222_y0, h_u_cla32_and5221_y0, h_u_cla32_and5223_y0);
  and_gate and_gate_h_u_cla32_and5224_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5224_y0);
  and_gate and_gate_h_u_cla32_and5225_y0(h_u_cla32_and5224_y0, h_u_cla32_and5223_y0, h_u_cla32_and5225_y0);
  and_gate and_gate_h_u_cla32_and5226_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5226_y0);
  and_gate and_gate_h_u_cla32_and5227_y0(h_u_cla32_and5226_y0, h_u_cla32_and5225_y0, h_u_cla32_and5227_y0);
  and_gate and_gate_h_u_cla32_and5228_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5228_y0);
  and_gate and_gate_h_u_cla32_and5229_y0(h_u_cla32_and5228_y0, h_u_cla32_and5227_y0, h_u_cla32_and5229_y0);
  and_gate and_gate_h_u_cla32_and5230_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5230_y0);
  and_gate and_gate_h_u_cla32_and5231_y0(h_u_cla32_and5230_y0, h_u_cla32_and5229_y0, h_u_cla32_and5231_y0);
  and_gate and_gate_h_u_cla32_and5232_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5232_y0);
  and_gate and_gate_h_u_cla32_and5233_y0(h_u_cla32_and5232_y0, h_u_cla32_and5231_y0, h_u_cla32_and5233_y0);
  and_gate and_gate_h_u_cla32_and5234_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5234_y0);
  and_gate and_gate_h_u_cla32_and5235_y0(h_u_cla32_and5234_y0, h_u_cla32_and5233_y0, h_u_cla32_and5235_y0);
  and_gate and_gate_h_u_cla32_and5236_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5236_y0);
  and_gate and_gate_h_u_cla32_and5237_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5237_y0);
  and_gate and_gate_h_u_cla32_and5238_y0(h_u_cla32_and5237_y0, h_u_cla32_and5236_y0, h_u_cla32_and5238_y0);
  and_gate and_gate_h_u_cla32_and5239_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5239_y0);
  and_gate and_gate_h_u_cla32_and5240_y0(h_u_cla32_and5239_y0, h_u_cla32_and5238_y0, h_u_cla32_and5240_y0);
  and_gate and_gate_h_u_cla32_and5241_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5241_y0);
  and_gate and_gate_h_u_cla32_and5242_y0(h_u_cla32_and5241_y0, h_u_cla32_and5240_y0, h_u_cla32_and5242_y0);
  and_gate and_gate_h_u_cla32_and5243_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5243_y0);
  and_gate and_gate_h_u_cla32_and5244_y0(h_u_cla32_and5243_y0, h_u_cla32_and5242_y0, h_u_cla32_and5244_y0);
  and_gate and_gate_h_u_cla32_and5245_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5245_y0);
  and_gate and_gate_h_u_cla32_and5246_y0(h_u_cla32_and5245_y0, h_u_cla32_and5244_y0, h_u_cla32_and5246_y0);
  and_gate and_gate_h_u_cla32_and5247_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5247_y0);
  and_gate and_gate_h_u_cla32_and5248_y0(h_u_cla32_and5247_y0, h_u_cla32_and5246_y0, h_u_cla32_and5248_y0);
  and_gate and_gate_h_u_cla32_and5249_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5249_y0);
  and_gate and_gate_h_u_cla32_and5250_y0(h_u_cla32_and5249_y0, h_u_cla32_and5248_y0, h_u_cla32_and5250_y0);
  and_gate and_gate_h_u_cla32_and5251_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5251_y0);
  and_gate and_gate_h_u_cla32_and5252_y0(h_u_cla32_and5251_y0, h_u_cla32_and5250_y0, h_u_cla32_and5252_y0);
  and_gate and_gate_h_u_cla32_and5253_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5253_y0);
  and_gate and_gate_h_u_cla32_and5254_y0(h_u_cla32_and5253_y0, h_u_cla32_and5252_y0, h_u_cla32_and5254_y0);
  and_gate and_gate_h_u_cla32_and5255_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5255_y0);
  and_gate and_gate_h_u_cla32_and5256_y0(h_u_cla32_and5255_y0, h_u_cla32_and5254_y0, h_u_cla32_and5256_y0);
  and_gate and_gate_h_u_cla32_and5257_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5257_y0);
  and_gate and_gate_h_u_cla32_and5258_y0(h_u_cla32_and5257_y0, h_u_cla32_and5256_y0, h_u_cla32_and5258_y0);
  and_gate and_gate_h_u_cla32_and5259_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5259_y0);
  and_gate and_gate_h_u_cla32_and5260_y0(h_u_cla32_and5259_y0, h_u_cla32_and5258_y0, h_u_cla32_and5260_y0);
  and_gate and_gate_h_u_cla32_and5261_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5261_y0);
  and_gate and_gate_h_u_cla32_and5262_y0(h_u_cla32_and5261_y0, h_u_cla32_and5260_y0, h_u_cla32_and5262_y0);
  and_gate and_gate_h_u_cla32_and5263_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5263_y0);
  and_gate and_gate_h_u_cla32_and5264_y0(h_u_cla32_and5263_y0, h_u_cla32_and5262_y0, h_u_cla32_and5264_y0);
  and_gate and_gate_h_u_cla32_and5265_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5265_y0);
  and_gate and_gate_h_u_cla32_and5266_y0(h_u_cla32_and5265_y0, h_u_cla32_and5264_y0, h_u_cla32_and5266_y0);
  and_gate and_gate_h_u_cla32_and5267_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5267_y0);
  and_gate and_gate_h_u_cla32_and5268_y0(h_u_cla32_and5267_y0, h_u_cla32_and5266_y0, h_u_cla32_and5268_y0);
  and_gate and_gate_h_u_cla32_and5269_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5269_y0);
  and_gate and_gate_h_u_cla32_and5270_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5270_y0);
  and_gate and_gate_h_u_cla32_and5271_y0(h_u_cla32_and5270_y0, h_u_cla32_and5269_y0, h_u_cla32_and5271_y0);
  and_gate and_gate_h_u_cla32_and5272_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5272_y0);
  and_gate and_gate_h_u_cla32_and5273_y0(h_u_cla32_and5272_y0, h_u_cla32_and5271_y0, h_u_cla32_and5273_y0);
  and_gate and_gate_h_u_cla32_and5274_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5274_y0);
  and_gate and_gate_h_u_cla32_and5275_y0(h_u_cla32_and5274_y0, h_u_cla32_and5273_y0, h_u_cla32_and5275_y0);
  and_gate and_gate_h_u_cla32_and5276_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5276_y0);
  and_gate and_gate_h_u_cla32_and5277_y0(h_u_cla32_and5276_y0, h_u_cla32_and5275_y0, h_u_cla32_and5277_y0);
  and_gate and_gate_h_u_cla32_and5278_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5278_y0);
  and_gate and_gate_h_u_cla32_and5279_y0(h_u_cla32_and5278_y0, h_u_cla32_and5277_y0, h_u_cla32_and5279_y0);
  and_gate and_gate_h_u_cla32_and5280_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5280_y0);
  and_gate and_gate_h_u_cla32_and5281_y0(h_u_cla32_and5280_y0, h_u_cla32_and5279_y0, h_u_cla32_and5281_y0);
  and_gate and_gate_h_u_cla32_and5282_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5282_y0);
  and_gate and_gate_h_u_cla32_and5283_y0(h_u_cla32_and5282_y0, h_u_cla32_and5281_y0, h_u_cla32_and5283_y0);
  and_gate and_gate_h_u_cla32_and5284_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5284_y0);
  and_gate and_gate_h_u_cla32_and5285_y0(h_u_cla32_and5284_y0, h_u_cla32_and5283_y0, h_u_cla32_and5285_y0);
  and_gate and_gate_h_u_cla32_and5286_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5286_y0);
  and_gate and_gate_h_u_cla32_and5287_y0(h_u_cla32_and5286_y0, h_u_cla32_and5285_y0, h_u_cla32_and5287_y0);
  and_gate and_gate_h_u_cla32_and5288_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5288_y0);
  and_gate and_gate_h_u_cla32_and5289_y0(h_u_cla32_and5288_y0, h_u_cla32_and5287_y0, h_u_cla32_and5289_y0);
  and_gate and_gate_h_u_cla32_and5290_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5290_y0);
  and_gate and_gate_h_u_cla32_and5291_y0(h_u_cla32_and5290_y0, h_u_cla32_and5289_y0, h_u_cla32_and5291_y0);
  and_gate and_gate_h_u_cla32_and5292_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5292_y0);
  and_gate and_gate_h_u_cla32_and5293_y0(h_u_cla32_and5292_y0, h_u_cla32_and5291_y0, h_u_cla32_and5293_y0);
  and_gate and_gate_h_u_cla32_and5294_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5294_y0);
  and_gate and_gate_h_u_cla32_and5295_y0(h_u_cla32_and5294_y0, h_u_cla32_and5293_y0, h_u_cla32_and5295_y0);
  and_gate and_gate_h_u_cla32_and5296_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5296_y0);
  and_gate and_gate_h_u_cla32_and5297_y0(h_u_cla32_and5296_y0, h_u_cla32_and5295_y0, h_u_cla32_and5297_y0);
  and_gate and_gate_h_u_cla32_and5298_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5298_y0);
  and_gate and_gate_h_u_cla32_and5299_y0(h_u_cla32_and5298_y0, h_u_cla32_and5297_y0, h_u_cla32_and5299_y0);
  and_gate and_gate_h_u_cla32_and5300_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5300_y0);
  and_gate and_gate_h_u_cla32_and5301_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5301_y0);
  and_gate and_gate_h_u_cla32_and5302_y0(h_u_cla32_and5301_y0, h_u_cla32_and5300_y0, h_u_cla32_and5302_y0);
  and_gate and_gate_h_u_cla32_and5303_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5303_y0);
  and_gate and_gate_h_u_cla32_and5304_y0(h_u_cla32_and5303_y0, h_u_cla32_and5302_y0, h_u_cla32_and5304_y0);
  and_gate and_gate_h_u_cla32_and5305_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5305_y0);
  and_gate and_gate_h_u_cla32_and5306_y0(h_u_cla32_and5305_y0, h_u_cla32_and5304_y0, h_u_cla32_and5306_y0);
  and_gate and_gate_h_u_cla32_and5307_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5307_y0);
  and_gate and_gate_h_u_cla32_and5308_y0(h_u_cla32_and5307_y0, h_u_cla32_and5306_y0, h_u_cla32_and5308_y0);
  and_gate and_gate_h_u_cla32_and5309_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5309_y0);
  and_gate and_gate_h_u_cla32_and5310_y0(h_u_cla32_and5309_y0, h_u_cla32_and5308_y0, h_u_cla32_and5310_y0);
  and_gate and_gate_h_u_cla32_and5311_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5311_y0);
  and_gate and_gate_h_u_cla32_and5312_y0(h_u_cla32_and5311_y0, h_u_cla32_and5310_y0, h_u_cla32_and5312_y0);
  and_gate and_gate_h_u_cla32_and5313_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5313_y0);
  and_gate and_gate_h_u_cla32_and5314_y0(h_u_cla32_and5313_y0, h_u_cla32_and5312_y0, h_u_cla32_and5314_y0);
  and_gate and_gate_h_u_cla32_and5315_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5315_y0);
  and_gate and_gate_h_u_cla32_and5316_y0(h_u_cla32_and5315_y0, h_u_cla32_and5314_y0, h_u_cla32_and5316_y0);
  and_gate and_gate_h_u_cla32_and5317_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5317_y0);
  and_gate and_gate_h_u_cla32_and5318_y0(h_u_cla32_and5317_y0, h_u_cla32_and5316_y0, h_u_cla32_and5318_y0);
  and_gate and_gate_h_u_cla32_and5319_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5319_y0);
  and_gate and_gate_h_u_cla32_and5320_y0(h_u_cla32_and5319_y0, h_u_cla32_and5318_y0, h_u_cla32_and5320_y0);
  and_gate and_gate_h_u_cla32_and5321_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5321_y0);
  and_gate and_gate_h_u_cla32_and5322_y0(h_u_cla32_and5321_y0, h_u_cla32_and5320_y0, h_u_cla32_and5322_y0);
  and_gate and_gate_h_u_cla32_and5323_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5323_y0);
  and_gate and_gate_h_u_cla32_and5324_y0(h_u_cla32_and5323_y0, h_u_cla32_and5322_y0, h_u_cla32_and5324_y0);
  and_gate and_gate_h_u_cla32_and5325_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5325_y0);
  and_gate and_gate_h_u_cla32_and5326_y0(h_u_cla32_and5325_y0, h_u_cla32_and5324_y0, h_u_cla32_and5326_y0);
  and_gate and_gate_h_u_cla32_and5327_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5327_y0);
  and_gate and_gate_h_u_cla32_and5328_y0(h_u_cla32_and5327_y0, h_u_cla32_and5326_y0, h_u_cla32_and5328_y0);
  and_gate and_gate_h_u_cla32_and5329_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5329_y0);
  and_gate and_gate_h_u_cla32_and5330_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5330_y0);
  and_gate and_gate_h_u_cla32_and5331_y0(h_u_cla32_and5330_y0, h_u_cla32_and5329_y0, h_u_cla32_and5331_y0);
  and_gate and_gate_h_u_cla32_and5332_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5332_y0);
  and_gate and_gate_h_u_cla32_and5333_y0(h_u_cla32_and5332_y0, h_u_cla32_and5331_y0, h_u_cla32_and5333_y0);
  and_gate and_gate_h_u_cla32_and5334_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5334_y0);
  and_gate and_gate_h_u_cla32_and5335_y0(h_u_cla32_and5334_y0, h_u_cla32_and5333_y0, h_u_cla32_and5335_y0);
  and_gate and_gate_h_u_cla32_and5336_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5336_y0);
  and_gate and_gate_h_u_cla32_and5337_y0(h_u_cla32_and5336_y0, h_u_cla32_and5335_y0, h_u_cla32_and5337_y0);
  and_gate and_gate_h_u_cla32_and5338_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5338_y0);
  and_gate and_gate_h_u_cla32_and5339_y0(h_u_cla32_and5338_y0, h_u_cla32_and5337_y0, h_u_cla32_and5339_y0);
  and_gate and_gate_h_u_cla32_and5340_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5340_y0);
  and_gate and_gate_h_u_cla32_and5341_y0(h_u_cla32_and5340_y0, h_u_cla32_and5339_y0, h_u_cla32_and5341_y0);
  and_gate and_gate_h_u_cla32_and5342_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5342_y0);
  and_gate and_gate_h_u_cla32_and5343_y0(h_u_cla32_and5342_y0, h_u_cla32_and5341_y0, h_u_cla32_and5343_y0);
  and_gate and_gate_h_u_cla32_and5344_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5344_y0);
  and_gate and_gate_h_u_cla32_and5345_y0(h_u_cla32_and5344_y0, h_u_cla32_and5343_y0, h_u_cla32_and5345_y0);
  and_gate and_gate_h_u_cla32_and5346_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5346_y0);
  and_gate and_gate_h_u_cla32_and5347_y0(h_u_cla32_and5346_y0, h_u_cla32_and5345_y0, h_u_cla32_and5347_y0);
  and_gate and_gate_h_u_cla32_and5348_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5348_y0);
  and_gate and_gate_h_u_cla32_and5349_y0(h_u_cla32_and5348_y0, h_u_cla32_and5347_y0, h_u_cla32_and5349_y0);
  and_gate and_gate_h_u_cla32_and5350_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5350_y0);
  and_gate and_gate_h_u_cla32_and5351_y0(h_u_cla32_and5350_y0, h_u_cla32_and5349_y0, h_u_cla32_and5351_y0);
  and_gate and_gate_h_u_cla32_and5352_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5352_y0);
  and_gate and_gate_h_u_cla32_and5353_y0(h_u_cla32_and5352_y0, h_u_cla32_and5351_y0, h_u_cla32_and5353_y0);
  and_gate and_gate_h_u_cla32_and5354_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5354_y0);
  and_gate and_gate_h_u_cla32_and5355_y0(h_u_cla32_and5354_y0, h_u_cla32_and5353_y0, h_u_cla32_and5355_y0);
  and_gate and_gate_h_u_cla32_and5356_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5356_y0);
  and_gate and_gate_h_u_cla32_and5357_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5357_y0);
  and_gate and_gate_h_u_cla32_and5358_y0(h_u_cla32_and5357_y0, h_u_cla32_and5356_y0, h_u_cla32_and5358_y0);
  and_gate and_gate_h_u_cla32_and5359_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5359_y0);
  and_gate and_gate_h_u_cla32_and5360_y0(h_u_cla32_and5359_y0, h_u_cla32_and5358_y0, h_u_cla32_and5360_y0);
  and_gate and_gate_h_u_cla32_and5361_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5361_y0);
  and_gate and_gate_h_u_cla32_and5362_y0(h_u_cla32_and5361_y0, h_u_cla32_and5360_y0, h_u_cla32_and5362_y0);
  and_gate and_gate_h_u_cla32_and5363_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5363_y0);
  and_gate and_gate_h_u_cla32_and5364_y0(h_u_cla32_and5363_y0, h_u_cla32_and5362_y0, h_u_cla32_and5364_y0);
  and_gate and_gate_h_u_cla32_and5365_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5365_y0);
  and_gate and_gate_h_u_cla32_and5366_y0(h_u_cla32_and5365_y0, h_u_cla32_and5364_y0, h_u_cla32_and5366_y0);
  and_gate and_gate_h_u_cla32_and5367_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5367_y0);
  and_gate and_gate_h_u_cla32_and5368_y0(h_u_cla32_and5367_y0, h_u_cla32_and5366_y0, h_u_cla32_and5368_y0);
  and_gate and_gate_h_u_cla32_and5369_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5369_y0);
  and_gate and_gate_h_u_cla32_and5370_y0(h_u_cla32_and5369_y0, h_u_cla32_and5368_y0, h_u_cla32_and5370_y0);
  and_gate and_gate_h_u_cla32_and5371_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5371_y0);
  and_gate and_gate_h_u_cla32_and5372_y0(h_u_cla32_and5371_y0, h_u_cla32_and5370_y0, h_u_cla32_and5372_y0);
  and_gate and_gate_h_u_cla32_and5373_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5373_y0);
  and_gate and_gate_h_u_cla32_and5374_y0(h_u_cla32_and5373_y0, h_u_cla32_and5372_y0, h_u_cla32_and5374_y0);
  and_gate and_gate_h_u_cla32_and5375_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5375_y0);
  and_gate and_gate_h_u_cla32_and5376_y0(h_u_cla32_and5375_y0, h_u_cla32_and5374_y0, h_u_cla32_and5376_y0);
  and_gate and_gate_h_u_cla32_and5377_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5377_y0);
  and_gate and_gate_h_u_cla32_and5378_y0(h_u_cla32_and5377_y0, h_u_cla32_and5376_y0, h_u_cla32_and5378_y0);
  and_gate and_gate_h_u_cla32_and5379_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and5379_y0);
  and_gate and_gate_h_u_cla32_and5380_y0(h_u_cla32_and5379_y0, h_u_cla32_and5378_y0, h_u_cla32_and5380_y0);
  and_gate and_gate_h_u_cla32_and5381_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5381_y0);
  and_gate and_gate_h_u_cla32_and5382_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5382_y0);
  and_gate and_gate_h_u_cla32_and5383_y0(h_u_cla32_and5382_y0, h_u_cla32_and5381_y0, h_u_cla32_and5383_y0);
  and_gate and_gate_h_u_cla32_and5384_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5384_y0);
  and_gate and_gate_h_u_cla32_and5385_y0(h_u_cla32_and5384_y0, h_u_cla32_and5383_y0, h_u_cla32_and5385_y0);
  and_gate and_gate_h_u_cla32_and5386_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5386_y0);
  and_gate and_gate_h_u_cla32_and5387_y0(h_u_cla32_and5386_y0, h_u_cla32_and5385_y0, h_u_cla32_and5387_y0);
  and_gate and_gate_h_u_cla32_and5388_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5388_y0);
  and_gate and_gate_h_u_cla32_and5389_y0(h_u_cla32_and5388_y0, h_u_cla32_and5387_y0, h_u_cla32_and5389_y0);
  and_gate and_gate_h_u_cla32_and5390_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5390_y0);
  and_gate and_gate_h_u_cla32_and5391_y0(h_u_cla32_and5390_y0, h_u_cla32_and5389_y0, h_u_cla32_and5391_y0);
  and_gate and_gate_h_u_cla32_and5392_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5392_y0);
  and_gate and_gate_h_u_cla32_and5393_y0(h_u_cla32_and5392_y0, h_u_cla32_and5391_y0, h_u_cla32_and5393_y0);
  and_gate and_gate_h_u_cla32_and5394_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5394_y0);
  and_gate and_gate_h_u_cla32_and5395_y0(h_u_cla32_and5394_y0, h_u_cla32_and5393_y0, h_u_cla32_and5395_y0);
  and_gate and_gate_h_u_cla32_and5396_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5396_y0);
  and_gate and_gate_h_u_cla32_and5397_y0(h_u_cla32_and5396_y0, h_u_cla32_and5395_y0, h_u_cla32_and5397_y0);
  and_gate and_gate_h_u_cla32_and5398_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5398_y0);
  and_gate and_gate_h_u_cla32_and5399_y0(h_u_cla32_and5398_y0, h_u_cla32_and5397_y0, h_u_cla32_and5399_y0);
  and_gate and_gate_h_u_cla32_and5400_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5400_y0);
  and_gate and_gate_h_u_cla32_and5401_y0(h_u_cla32_and5400_y0, h_u_cla32_and5399_y0, h_u_cla32_and5401_y0);
  and_gate and_gate_h_u_cla32_and5402_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and5402_y0);
  and_gate and_gate_h_u_cla32_and5403_y0(h_u_cla32_and5402_y0, h_u_cla32_and5401_y0, h_u_cla32_and5403_y0);
  and_gate and_gate_h_u_cla32_and5404_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5404_y0);
  and_gate and_gate_h_u_cla32_and5405_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5405_y0);
  and_gate and_gate_h_u_cla32_and5406_y0(h_u_cla32_and5405_y0, h_u_cla32_and5404_y0, h_u_cla32_and5406_y0);
  and_gate and_gate_h_u_cla32_and5407_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5407_y0);
  and_gate and_gate_h_u_cla32_and5408_y0(h_u_cla32_and5407_y0, h_u_cla32_and5406_y0, h_u_cla32_and5408_y0);
  and_gate and_gate_h_u_cla32_and5409_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5409_y0);
  and_gate and_gate_h_u_cla32_and5410_y0(h_u_cla32_and5409_y0, h_u_cla32_and5408_y0, h_u_cla32_and5410_y0);
  and_gate and_gate_h_u_cla32_and5411_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5411_y0);
  and_gate and_gate_h_u_cla32_and5412_y0(h_u_cla32_and5411_y0, h_u_cla32_and5410_y0, h_u_cla32_and5412_y0);
  and_gate and_gate_h_u_cla32_and5413_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5413_y0);
  and_gate and_gate_h_u_cla32_and5414_y0(h_u_cla32_and5413_y0, h_u_cla32_and5412_y0, h_u_cla32_and5414_y0);
  and_gate and_gate_h_u_cla32_and5415_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5415_y0);
  and_gate and_gate_h_u_cla32_and5416_y0(h_u_cla32_and5415_y0, h_u_cla32_and5414_y0, h_u_cla32_and5416_y0);
  and_gate and_gate_h_u_cla32_and5417_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5417_y0);
  and_gate and_gate_h_u_cla32_and5418_y0(h_u_cla32_and5417_y0, h_u_cla32_and5416_y0, h_u_cla32_and5418_y0);
  and_gate and_gate_h_u_cla32_and5419_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5419_y0);
  and_gate and_gate_h_u_cla32_and5420_y0(h_u_cla32_and5419_y0, h_u_cla32_and5418_y0, h_u_cla32_and5420_y0);
  and_gate and_gate_h_u_cla32_and5421_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5421_y0);
  and_gate and_gate_h_u_cla32_and5422_y0(h_u_cla32_and5421_y0, h_u_cla32_and5420_y0, h_u_cla32_and5422_y0);
  and_gate and_gate_h_u_cla32_and5423_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and5423_y0);
  and_gate and_gate_h_u_cla32_and5424_y0(h_u_cla32_and5423_y0, h_u_cla32_and5422_y0, h_u_cla32_and5424_y0);
  and_gate and_gate_h_u_cla32_and5425_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5425_y0);
  and_gate and_gate_h_u_cla32_and5426_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5426_y0);
  and_gate and_gate_h_u_cla32_and5427_y0(h_u_cla32_and5426_y0, h_u_cla32_and5425_y0, h_u_cla32_and5427_y0);
  and_gate and_gate_h_u_cla32_and5428_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5428_y0);
  and_gate and_gate_h_u_cla32_and5429_y0(h_u_cla32_and5428_y0, h_u_cla32_and5427_y0, h_u_cla32_and5429_y0);
  and_gate and_gate_h_u_cla32_and5430_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5430_y0);
  and_gate and_gate_h_u_cla32_and5431_y0(h_u_cla32_and5430_y0, h_u_cla32_and5429_y0, h_u_cla32_and5431_y0);
  and_gate and_gate_h_u_cla32_and5432_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5432_y0);
  and_gate and_gate_h_u_cla32_and5433_y0(h_u_cla32_and5432_y0, h_u_cla32_and5431_y0, h_u_cla32_and5433_y0);
  and_gate and_gate_h_u_cla32_and5434_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5434_y0);
  and_gate and_gate_h_u_cla32_and5435_y0(h_u_cla32_and5434_y0, h_u_cla32_and5433_y0, h_u_cla32_and5435_y0);
  and_gate and_gate_h_u_cla32_and5436_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5436_y0);
  and_gate and_gate_h_u_cla32_and5437_y0(h_u_cla32_and5436_y0, h_u_cla32_and5435_y0, h_u_cla32_and5437_y0);
  and_gate and_gate_h_u_cla32_and5438_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5438_y0);
  and_gate and_gate_h_u_cla32_and5439_y0(h_u_cla32_and5438_y0, h_u_cla32_and5437_y0, h_u_cla32_and5439_y0);
  and_gate and_gate_h_u_cla32_and5440_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5440_y0);
  and_gate and_gate_h_u_cla32_and5441_y0(h_u_cla32_and5440_y0, h_u_cla32_and5439_y0, h_u_cla32_and5441_y0);
  and_gate and_gate_h_u_cla32_and5442_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and5442_y0);
  and_gate and_gate_h_u_cla32_and5443_y0(h_u_cla32_and5442_y0, h_u_cla32_and5441_y0, h_u_cla32_and5443_y0);
  and_gate and_gate_h_u_cla32_and5444_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5444_y0);
  and_gate and_gate_h_u_cla32_and5445_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5445_y0);
  and_gate and_gate_h_u_cla32_and5446_y0(h_u_cla32_and5445_y0, h_u_cla32_and5444_y0, h_u_cla32_and5446_y0);
  and_gate and_gate_h_u_cla32_and5447_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5447_y0);
  and_gate and_gate_h_u_cla32_and5448_y0(h_u_cla32_and5447_y0, h_u_cla32_and5446_y0, h_u_cla32_and5448_y0);
  and_gate and_gate_h_u_cla32_and5449_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5449_y0);
  and_gate and_gate_h_u_cla32_and5450_y0(h_u_cla32_and5449_y0, h_u_cla32_and5448_y0, h_u_cla32_and5450_y0);
  and_gate and_gate_h_u_cla32_and5451_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5451_y0);
  and_gate and_gate_h_u_cla32_and5452_y0(h_u_cla32_and5451_y0, h_u_cla32_and5450_y0, h_u_cla32_and5452_y0);
  and_gate and_gate_h_u_cla32_and5453_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5453_y0);
  and_gate and_gate_h_u_cla32_and5454_y0(h_u_cla32_and5453_y0, h_u_cla32_and5452_y0, h_u_cla32_and5454_y0);
  and_gate and_gate_h_u_cla32_and5455_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5455_y0);
  and_gate and_gate_h_u_cla32_and5456_y0(h_u_cla32_and5455_y0, h_u_cla32_and5454_y0, h_u_cla32_and5456_y0);
  and_gate and_gate_h_u_cla32_and5457_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5457_y0);
  and_gate and_gate_h_u_cla32_and5458_y0(h_u_cla32_and5457_y0, h_u_cla32_and5456_y0, h_u_cla32_and5458_y0);
  and_gate and_gate_h_u_cla32_and5459_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and5459_y0);
  and_gate and_gate_h_u_cla32_and5460_y0(h_u_cla32_and5459_y0, h_u_cla32_and5458_y0, h_u_cla32_and5460_y0);
  and_gate and_gate_h_u_cla32_and5461_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5461_y0);
  and_gate and_gate_h_u_cla32_and5462_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5462_y0);
  and_gate and_gate_h_u_cla32_and5463_y0(h_u_cla32_and5462_y0, h_u_cla32_and5461_y0, h_u_cla32_and5463_y0);
  and_gate and_gate_h_u_cla32_and5464_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5464_y0);
  and_gate and_gate_h_u_cla32_and5465_y0(h_u_cla32_and5464_y0, h_u_cla32_and5463_y0, h_u_cla32_and5465_y0);
  and_gate and_gate_h_u_cla32_and5466_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5466_y0);
  and_gate and_gate_h_u_cla32_and5467_y0(h_u_cla32_and5466_y0, h_u_cla32_and5465_y0, h_u_cla32_and5467_y0);
  and_gate and_gate_h_u_cla32_and5468_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5468_y0);
  and_gate and_gate_h_u_cla32_and5469_y0(h_u_cla32_and5468_y0, h_u_cla32_and5467_y0, h_u_cla32_and5469_y0);
  and_gate and_gate_h_u_cla32_and5470_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5470_y0);
  and_gate and_gate_h_u_cla32_and5471_y0(h_u_cla32_and5470_y0, h_u_cla32_and5469_y0, h_u_cla32_and5471_y0);
  and_gate and_gate_h_u_cla32_and5472_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5472_y0);
  and_gate and_gate_h_u_cla32_and5473_y0(h_u_cla32_and5472_y0, h_u_cla32_and5471_y0, h_u_cla32_and5473_y0);
  and_gate and_gate_h_u_cla32_and5474_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and5474_y0);
  and_gate and_gate_h_u_cla32_and5475_y0(h_u_cla32_and5474_y0, h_u_cla32_and5473_y0, h_u_cla32_and5475_y0);
  and_gate and_gate_h_u_cla32_and5476_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5476_y0);
  and_gate and_gate_h_u_cla32_and5477_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5477_y0);
  and_gate and_gate_h_u_cla32_and5478_y0(h_u_cla32_and5477_y0, h_u_cla32_and5476_y0, h_u_cla32_and5478_y0);
  and_gate and_gate_h_u_cla32_and5479_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5479_y0);
  and_gate and_gate_h_u_cla32_and5480_y0(h_u_cla32_and5479_y0, h_u_cla32_and5478_y0, h_u_cla32_and5480_y0);
  and_gate and_gate_h_u_cla32_and5481_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5481_y0);
  and_gate and_gate_h_u_cla32_and5482_y0(h_u_cla32_and5481_y0, h_u_cla32_and5480_y0, h_u_cla32_and5482_y0);
  and_gate and_gate_h_u_cla32_and5483_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5483_y0);
  and_gate and_gate_h_u_cla32_and5484_y0(h_u_cla32_and5483_y0, h_u_cla32_and5482_y0, h_u_cla32_and5484_y0);
  and_gate and_gate_h_u_cla32_and5485_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5485_y0);
  and_gate and_gate_h_u_cla32_and5486_y0(h_u_cla32_and5485_y0, h_u_cla32_and5484_y0, h_u_cla32_and5486_y0);
  and_gate and_gate_h_u_cla32_and5487_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and5487_y0);
  and_gate and_gate_h_u_cla32_and5488_y0(h_u_cla32_and5487_y0, h_u_cla32_and5486_y0, h_u_cla32_and5488_y0);
  and_gate and_gate_h_u_cla32_and5489_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and5489_y0);
  and_gate and_gate_h_u_cla32_and5490_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and5490_y0);
  and_gate and_gate_h_u_cla32_and5491_y0(h_u_cla32_and5490_y0, h_u_cla32_and5489_y0, h_u_cla32_and5491_y0);
  and_gate and_gate_h_u_cla32_and5492_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and5492_y0);
  and_gate and_gate_h_u_cla32_and5493_y0(h_u_cla32_and5492_y0, h_u_cla32_and5491_y0, h_u_cla32_and5493_y0);
  and_gate and_gate_h_u_cla32_and5494_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and5494_y0);
  and_gate and_gate_h_u_cla32_and5495_y0(h_u_cla32_and5494_y0, h_u_cla32_and5493_y0, h_u_cla32_and5495_y0);
  and_gate and_gate_h_u_cla32_and5496_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and5496_y0);
  and_gate and_gate_h_u_cla32_and5497_y0(h_u_cla32_and5496_y0, h_u_cla32_and5495_y0, h_u_cla32_and5497_y0);
  and_gate and_gate_h_u_cla32_and5498_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and5498_y0);
  and_gate and_gate_h_u_cla32_and5499_y0(h_u_cla32_and5498_y0, h_u_cla32_and5497_y0, h_u_cla32_and5499_y0);
  and_gate and_gate_h_u_cla32_and5500_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and5500_y0);
  and_gate and_gate_h_u_cla32_and5501_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and5501_y0);
  and_gate and_gate_h_u_cla32_and5502_y0(h_u_cla32_and5501_y0, h_u_cla32_and5500_y0, h_u_cla32_and5502_y0);
  and_gate and_gate_h_u_cla32_and5503_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and5503_y0);
  and_gate and_gate_h_u_cla32_and5504_y0(h_u_cla32_and5503_y0, h_u_cla32_and5502_y0, h_u_cla32_and5504_y0);
  and_gate and_gate_h_u_cla32_and5505_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and5505_y0);
  and_gate and_gate_h_u_cla32_and5506_y0(h_u_cla32_and5505_y0, h_u_cla32_and5504_y0, h_u_cla32_and5506_y0);
  and_gate and_gate_h_u_cla32_and5507_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and5507_y0);
  and_gate and_gate_h_u_cla32_and5508_y0(h_u_cla32_and5507_y0, h_u_cla32_and5506_y0, h_u_cla32_and5508_y0);
  and_gate and_gate_h_u_cla32_and5509_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and5509_y0);
  and_gate and_gate_h_u_cla32_and5510_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and5510_y0);
  and_gate and_gate_h_u_cla32_and5511_y0(h_u_cla32_and5510_y0, h_u_cla32_and5509_y0, h_u_cla32_and5511_y0);
  and_gate and_gate_h_u_cla32_and5512_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and5512_y0);
  and_gate and_gate_h_u_cla32_and5513_y0(h_u_cla32_and5512_y0, h_u_cla32_and5511_y0, h_u_cla32_and5513_y0);
  and_gate and_gate_h_u_cla32_and5514_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and5514_y0);
  and_gate and_gate_h_u_cla32_and5515_y0(h_u_cla32_and5514_y0, h_u_cla32_and5513_y0, h_u_cla32_and5515_y0);
  and_gate and_gate_h_u_cla32_and5516_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and5516_y0);
  and_gate and_gate_h_u_cla32_and5517_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and5517_y0);
  and_gate and_gate_h_u_cla32_and5518_y0(h_u_cla32_and5517_y0, h_u_cla32_and5516_y0, h_u_cla32_and5518_y0);
  and_gate and_gate_h_u_cla32_and5519_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and5519_y0);
  and_gate and_gate_h_u_cla32_and5520_y0(h_u_cla32_and5519_y0, h_u_cla32_and5518_y0, h_u_cla32_and5520_y0);
  and_gate and_gate_h_u_cla32_and5521_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and5521_y0);
  and_gate and_gate_h_u_cla32_and5522_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and5522_y0);
  and_gate and_gate_h_u_cla32_and5523_y0(h_u_cla32_and5522_y0, h_u_cla32_and5521_y0, h_u_cla32_and5523_y0);
  and_gate and_gate_h_u_cla32_and5524_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and5524_y0);
  or_gate or_gate_h_u_cla32_or300_y0(h_u_cla32_and5524_y0, h_u_cla32_and4948_y0, h_u_cla32_or300_y0);
  or_gate or_gate_h_u_cla32_or301_y0(h_u_cla32_or300_y0, h_u_cla32_and4995_y0, h_u_cla32_or301_y0);
  or_gate or_gate_h_u_cla32_or302_y0(h_u_cla32_or301_y0, h_u_cla32_and5040_y0, h_u_cla32_or302_y0);
  or_gate or_gate_h_u_cla32_or303_y0(h_u_cla32_or302_y0, h_u_cla32_and5083_y0, h_u_cla32_or303_y0);
  or_gate or_gate_h_u_cla32_or304_y0(h_u_cla32_or303_y0, h_u_cla32_and5124_y0, h_u_cla32_or304_y0);
  or_gate or_gate_h_u_cla32_or305_y0(h_u_cla32_or304_y0, h_u_cla32_and5163_y0, h_u_cla32_or305_y0);
  or_gate or_gate_h_u_cla32_or306_y0(h_u_cla32_or305_y0, h_u_cla32_and5200_y0, h_u_cla32_or306_y0);
  or_gate or_gate_h_u_cla32_or307_y0(h_u_cla32_or306_y0, h_u_cla32_and5235_y0, h_u_cla32_or307_y0);
  or_gate or_gate_h_u_cla32_or308_y0(h_u_cla32_or307_y0, h_u_cla32_and5268_y0, h_u_cla32_or308_y0);
  or_gate or_gate_h_u_cla32_or309_y0(h_u_cla32_or308_y0, h_u_cla32_and5299_y0, h_u_cla32_or309_y0);
  or_gate or_gate_h_u_cla32_or310_y0(h_u_cla32_or309_y0, h_u_cla32_and5328_y0, h_u_cla32_or310_y0);
  or_gate or_gate_h_u_cla32_or311_y0(h_u_cla32_or310_y0, h_u_cla32_and5355_y0, h_u_cla32_or311_y0);
  or_gate or_gate_h_u_cla32_or312_y0(h_u_cla32_or311_y0, h_u_cla32_and5380_y0, h_u_cla32_or312_y0);
  or_gate or_gate_h_u_cla32_or313_y0(h_u_cla32_or312_y0, h_u_cla32_and5403_y0, h_u_cla32_or313_y0);
  or_gate or_gate_h_u_cla32_or314_y0(h_u_cla32_or313_y0, h_u_cla32_and5424_y0, h_u_cla32_or314_y0);
  or_gate or_gate_h_u_cla32_or315_y0(h_u_cla32_or314_y0, h_u_cla32_and5443_y0, h_u_cla32_or315_y0);
  or_gate or_gate_h_u_cla32_or316_y0(h_u_cla32_or315_y0, h_u_cla32_and5460_y0, h_u_cla32_or316_y0);
  or_gate or_gate_h_u_cla32_or317_y0(h_u_cla32_or316_y0, h_u_cla32_and5475_y0, h_u_cla32_or317_y0);
  or_gate or_gate_h_u_cla32_or318_y0(h_u_cla32_or317_y0, h_u_cla32_and5488_y0, h_u_cla32_or318_y0);
  or_gate or_gate_h_u_cla32_or319_y0(h_u_cla32_or318_y0, h_u_cla32_and5499_y0, h_u_cla32_or319_y0);
  or_gate or_gate_h_u_cla32_or320_y0(h_u_cla32_or319_y0, h_u_cla32_and5508_y0, h_u_cla32_or320_y0);
  or_gate or_gate_h_u_cla32_or321_y0(h_u_cla32_or320_y0, h_u_cla32_and5515_y0, h_u_cla32_or321_y0);
  or_gate or_gate_h_u_cla32_or322_y0(h_u_cla32_or321_y0, h_u_cla32_and5520_y0, h_u_cla32_or322_y0);
  or_gate or_gate_h_u_cla32_or323_y0(h_u_cla32_or322_y0, h_u_cla32_and5523_y0, h_u_cla32_or323_y0);
  or_gate or_gate_h_u_cla32_or324_y0(h_u_cla32_pg_logic24_y1, h_u_cla32_or323_y0, h_u_cla32_or324_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic25_y0(a_25, b_25, h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_pg_logic25_y2);
  xor_gate xor_gate_h_u_cla32_xor25_y0(h_u_cla32_pg_logic25_y2, h_u_cla32_or324_y0, h_u_cla32_xor25_y0);
  and_gate and_gate_h_u_cla32_and5525_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and5525_y0);
  and_gate and_gate_h_u_cla32_and5526_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and5526_y0);
  and_gate and_gate_h_u_cla32_and5527_y0(h_u_cla32_and5526_y0, h_u_cla32_and5525_y0, h_u_cla32_and5527_y0);
  and_gate and_gate_h_u_cla32_and5528_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and5528_y0);
  and_gate and_gate_h_u_cla32_and5529_y0(h_u_cla32_and5528_y0, h_u_cla32_and5527_y0, h_u_cla32_and5529_y0);
  and_gate and_gate_h_u_cla32_and5530_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and5530_y0);
  and_gate and_gate_h_u_cla32_and5531_y0(h_u_cla32_and5530_y0, h_u_cla32_and5529_y0, h_u_cla32_and5531_y0);
  and_gate and_gate_h_u_cla32_and5532_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and5532_y0);
  and_gate and_gate_h_u_cla32_and5533_y0(h_u_cla32_and5532_y0, h_u_cla32_and5531_y0, h_u_cla32_and5533_y0);
  and_gate and_gate_h_u_cla32_and5534_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and5534_y0);
  and_gate and_gate_h_u_cla32_and5535_y0(h_u_cla32_and5534_y0, h_u_cla32_and5533_y0, h_u_cla32_and5535_y0);
  and_gate and_gate_h_u_cla32_and5536_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and5536_y0);
  and_gate and_gate_h_u_cla32_and5537_y0(h_u_cla32_and5536_y0, h_u_cla32_and5535_y0, h_u_cla32_and5537_y0);
  and_gate and_gate_h_u_cla32_and5538_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and5538_y0);
  and_gate and_gate_h_u_cla32_and5539_y0(h_u_cla32_and5538_y0, h_u_cla32_and5537_y0, h_u_cla32_and5539_y0);
  and_gate and_gate_h_u_cla32_and5540_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and5540_y0);
  and_gate and_gate_h_u_cla32_and5541_y0(h_u_cla32_and5540_y0, h_u_cla32_and5539_y0, h_u_cla32_and5541_y0);
  and_gate and_gate_h_u_cla32_and5542_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and5542_y0);
  and_gate and_gate_h_u_cla32_and5543_y0(h_u_cla32_and5542_y0, h_u_cla32_and5541_y0, h_u_cla32_and5543_y0);
  and_gate and_gate_h_u_cla32_and5544_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and5544_y0);
  and_gate and_gate_h_u_cla32_and5545_y0(h_u_cla32_and5544_y0, h_u_cla32_and5543_y0, h_u_cla32_and5545_y0);
  and_gate and_gate_h_u_cla32_and5546_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and5546_y0);
  and_gate and_gate_h_u_cla32_and5547_y0(h_u_cla32_and5546_y0, h_u_cla32_and5545_y0, h_u_cla32_and5547_y0);
  and_gate and_gate_h_u_cla32_and5548_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and5548_y0);
  and_gate and_gate_h_u_cla32_and5549_y0(h_u_cla32_and5548_y0, h_u_cla32_and5547_y0, h_u_cla32_and5549_y0);
  and_gate and_gate_h_u_cla32_and5550_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and5550_y0);
  and_gate and_gate_h_u_cla32_and5551_y0(h_u_cla32_and5550_y0, h_u_cla32_and5549_y0, h_u_cla32_and5551_y0);
  and_gate and_gate_h_u_cla32_and5552_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and5552_y0);
  and_gate and_gate_h_u_cla32_and5553_y0(h_u_cla32_and5552_y0, h_u_cla32_and5551_y0, h_u_cla32_and5553_y0);
  and_gate and_gate_h_u_cla32_and5554_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and5554_y0);
  and_gate and_gate_h_u_cla32_and5555_y0(h_u_cla32_and5554_y0, h_u_cla32_and5553_y0, h_u_cla32_and5555_y0);
  and_gate and_gate_h_u_cla32_and5556_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and5556_y0);
  and_gate and_gate_h_u_cla32_and5557_y0(h_u_cla32_and5556_y0, h_u_cla32_and5555_y0, h_u_cla32_and5557_y0);
  and_gate and_gate_h_u_cla32_and5558_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and5558_y0);
  and_gate and_gate_h_u_cla32_and5559_y0(h_u_cla32_and5558_y0, h_u_cla32_and5557_y0, h_u_cla32_and5559_y0);
  and_gate and_gate_h_u_cla32_and5560_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and5560_y0);
  and_gate and_gate_h_u_cla32_and5561_y0(h_u_cla32_and5560_y0, h_u_cla32_and5559_y0, h_u_cla32_and5561_y0);
  and_gate and_gate_h_u_cla32_and5562_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and5562_y0);
  and_gate and_gate_h_u_cla32_and5563_y0(h_u_cla32_and5562_y0, h_u_cla32_and5561_y0, h_u_cla32_and5563_y0);
  and_gate and_gate_h_u_cla32_and5564_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and5564_y0);
  and_gate and_gate_h_u_cla32_and5565_y0(h_u_cla32_and5564_y0, h_u_cla32_and5563_y0, h_u_cla32_and5565_y0);
  and_gate and_gate_h_u_cla32_and5566_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and5566_y0);
  and_gate and_gate_h_u_cla32_and5567_y0(h_u_cla32_and5566_y0, h_u_cla32_and5565_y0, h_u_cla32_and5567_y0);
  and_gate and_gate_h_u_cla32_and5568_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and5568_y0);
  and_gate and_gate_h_u_cla32_and5569_y0(h_u_cla32_and5568_y0, h_u_cla32_and5567_y0, h_u_cla32_and5569_y0);
  and_gate and_gate_h_u_cla32_and5570_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and5570_y0);
  and_gate and_gate_h_u_cla32_and5571_y0(h_u_cla32_and5570_y0, h_u_cla32_and5569_y0, h_u_cla32_and5571_y0);
  and_gate and_gate_h_u_cla32_and5572_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and5572_y0);
  and_gate and_gate_h_u_cla32_and5573_y0(h_u_cla32_and5572_y0, h_u_cla32_and5571_y0, h_u_cla32_and5573_y0);
  and_gate and_gate_h_u_cla32_and5574_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and5574_y0);
  and_gate and_gate_h_u_cla32_and5575_y0(h_u_cla32_and5574_y0, h_u_cla32_and5573_y0, h_u_cla32_and5575_y0);
  and_gate and_gate_h_u_cla32_and5576_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5576_y0);
  and_gate and_gate_h_u_cla32_and5577_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5577_y0);
  and_gate and_gate_h_u_cla32_and5578_y0(h_u_cla32_and5577_y0, h_u_cla32_and5576_y0, h_u_cla32_and5578_y0);
  and_gate and_gate_h_u_cla32_and5579_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5579_y0);
  and_gate and_gate_h_u_cla32_and5580_y0(h_u_cla32_and5579_y0, h_u_cla32_and5578_y0, h_u_cla32_and5580_y0);
  and_gate and_gate_h_u_cla32_and5581_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5581_y0);
  and_gate and_gate_h_u_cla32_and5582_y0(h_u_cla32_and5581_y0, h_u_cla32_and5580_y0, h_u_cla32_and5582_y0);
  and_gate and_gate_h_u_cla32_and5583_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5583_y0);
  and_gate and_gate_h_u_cla32_and5584_y0(h_u_cla32_and5583_y0, h_u_cla32_and5582_y0, h_u_cla32_and5584_y0);
  and_gate and_gate_h_u_cla32_and5585_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5585_y0);
  and_gate and_gate_h_u_cla32_and5586_y0(h_u_cla32_and5585_y0, h_u_cla32_and5584_y0, h_u_cla32_and5586_y0);
  and_gate and_gate_h_u_cla32_and5587_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5587_y0);
  and_gate and_gate_h_u_cla32_and5588_y0(h_u_cla32_and5587_y0, h_u_cla32_and5586_y0, h_u_cla32_and5588_y0);
  and_gate and_gate_h_u_cla32_and5589_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5589_y0);
  and_gate and_gate_h_u_cla32_and5590_y0(h_u_cla32_and5589_y0, h_u_cla32_and5588_y0, h_u_cla32_and5590_y0);
  and_gate and_gate_h_u_cla32_and5591_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5591_y0);
  and_gate and_gate_h_u_cla32_and5592_y0(h_u_cla32_and5591_y0, h_u_cla32_and5590_y0, h_u_cla32_and5592_y0);
  and_gate and_gate_h_u_cla32_and5593_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5593_y0);
  and_gate and_gate_h_u_cla32_and5594_y0(h_u_cla32_and5593_y0, h_u_cla32_and5592_y0, h_u_cla32_and5594_y0);
  and_gate and_gate_h_u_cla32_and5595_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5595_y0);
  and_gate and_gate_h_u_cla32_and5596_y0(h_u_cla32_and5595_y0, h_u_cla32_and5594_y0, h_u_cla32_and5596_y0);
  and_gate and_gate_h_u_cla32_and5597_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5597_y0);
  and_gate and_gate_h_u_cla32_and5598_y0(h_u_cla32_and5597_y0, h_u_cla32_and5596_y0, h_u_cla32_and5598_y0);
  and_gate and_gate_h_u_cla32_and5599_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5599_y0);
  and_gate and_gate_h_u_cla32_and5600_y0(h_u_cla32_and5599_y0, h_u_cla32_and5598_y0, h_u_cla32_and5600_y0);
  and_gate and_gate_h_u_cla32_and5601_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5601_y0);
  and_gate and_gate_h_u_cla32_and5602_y0(h_u_cla32_and5601_y0, h_u_cla32_and5600_y0, h_u_cla32_and5602_y0);
  and_gate and_gate_h_u_cla32_and5603_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5603_y0);
  and_gate and_gate_h_u_cla32_and5604_y0(h_u_cla32_and5603_y0, h_u_cla32_and5602_y0, h_u_cla32_and5604_y0);
  and_gate and_gate_h_u_cla32_and5605_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5605_y0);
  and_gate and_gate_h_u_cla32_and5606_y0(h_u_cla32_and5605_y0, h_u_cla32_and5604_y0, h_u_cla32_and5606_y0);
  and_gate and_gate_h_u_cla32_and5607_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5607_y0);
  and_gate and_gate_h_u_cla32_and5608_y0(h_u_cla32_and5607_y0, h_u_cla32_and5606_y0, h_u_cla32_and5608_y0);
  and_gate and_gate_h_u_cla32_and5609_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5609_y0);
  and_gate and_gate_h_u_cla32_and5610_y0(h_u_cla32_and5609_y0, h_u_cla32_and5608_y0, h_u_cla32_and5610_y0);
  and_gate and_gate_h_u_cla32_and5611_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5611_y0);
  and_gate and_gate_h_u_cla32_and5612_y0(h_u_cla32_and5611_y0, h_u_cla32_and5610_y0, h_u_cla32_and5612_y0);
  and_gate and_gate_h_u_cla32_and5613_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5613_y0);
  and_gate and_gate_h_u_cla32_and5614_y0(h_u_cla32_and5613_y0, h_u_cla32_and5612_y0, h_u_cla32_and5614_y0);
  and_gate and_gate_h_u_cla32_and5615_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5615_y0);
  and_gate and_gate_h_u_cla32_and5616_y0(h_u_cla32_and5615_y0, h_u_cla32_and5614_y0, h_u_cla32_and5616_y0);
  and_gate and_gate_h_u_cla32_and5617_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5617_y0);
  and_gate and_gate_h_u_cla32_and5618_y0(h_u_cla32_and5617_y0, h_u_cla32_and5616_y0, h_u_cla32_and5618_y0);
  and_gate and_gate_h_u_cla32_and5619_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5619_y0);
  and_gate and_gate_h_u_cla32_and5620_y0(h_u_cla32_and5619_y0, h_u_cla32_and5618_y0, h_u_cla32_and5620_y0);
  and_gate and_gate_h_u_cla32_and5621_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5621_y0);
  and_gate and_gate_h_u_cla32_and5622_y0(h_u_cla32_and5621_y0, h_u_cla32_and5620_y0, h_u_cla32_and5622_y0);
  and_gate and_gate_h_u_cla32_and5623_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and5623_y0);
  and_gate and_gate_h_u_cla32_and5624_y0(h_u_cla32_and5623_y0, h_u_cla32_and5622_y0, h_u_cla32_and5624_y0);
  and_gate and_gate_h_u_cla32_and5625_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5625_y0);
  and_gate and_gate_h_u_cla32_and5626_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5626_y0);
  and_gate and_gate_h_u_cla32_and5627_y0(h_u_cla32_and5626_y0, h_u_cla32_and5625_y0, h_u_cla32_and5627_y0);
  and_gate and_gate_h_u_cla32_and5628_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5628_y0);
  and_gate and_gate_h_u_cla32_and5629_y0(h_u_cla32_and5628_y0, h_u_cla32_and5627_y0, h_u_cla32_and5629_y0);
  and_gate and_gate_h_u_cla32_and5630_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5630_y0);
  and_gate and_gate_h_u_cla32_and5631_y0(h_u_cla32_and5630_y0, h_u_cla32_and5629_y0, h_u_cla32_and5631_y0);
  and_gate and_gate_h_u_cla32_and5632_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5632_y0);
  and_gate and_gate_h_u_cla32_and5633_y0(h_u_cla32_and5632_y0, h_u_cla32_and5631_y0, h_u_cla32_and5633_y0);
  and_gate and_gate_h_u_cla32_and5634_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5634_y0);
  and_gate and_gate_h_u_cla32_and5635_y0(h_u_cla32_and5634_y0, h_u_cla32_and5633_y0, h_u_cla32_and5635_y0);
  and_gate and_gate_h_u_cla32_and5636_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5636_y0);
  and_gate and_gate_h_u_cla32_and5637_y0(h_u_cla32_and5636_y0, h_u_cla32_and5635_y0, h_u_cla32_and5637_y0);
  and_gate and_gate_h_u_cla32_and5638_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5638_y0);
  and_gate and_gate_h_u_cla32_and5639_y0(h_u_cla32_and5638_y0, h_u_cla32_and5637_y0, h_u_cla32_and5639_y0);
  and_gate and_gate_h_u_cla32_and5640_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5640_y0);
  and_gate and_gate_h_u_cla32_and5641_y0(h_u_cla32_and5640_y0, h_u_cla32_and5639_y0, h_u_cla32_and5641_y0);
  and_gate and_gate_h_u_cla32_and5642_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5642_y0);
  and_gate and_gate_h_u_cla32_and5643_y0(h_u_cla32_and5642_y0, h_u_cla32_and5641_y0, h_u_cla32_and5643_y0);
  and_gate and_gate_h_u_cla32_and5644_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5644_y0);
  and_gate and_gate_h_u_cla32_and5645_y0(h_u_cla32_and5644_y0, h_u_cla32_and5643_y0, h_u_cla32_and5645_y0);
  and_gate and_gate_h_u_cla32_and5646_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5646_y0);
  and_gate and_gate_h_u_cla32_and5647_y0(h_u_cla32_and5646_y0, h_u_cla32_and5645_y0, h_u_cla32_and5647_y0);
  and_gate and_gate_h_u_cla32_and5648_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5648_y0);
  and_gate and_gate_h_u_cla32_and5649_y0(h_u_cla32_and5648_y0, h_u_cla32_and5647_y0, h_u_cla32_and5649_y0);
  and_gate and_gate_h_u_cla32_and5650_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5650_y0);
  and_gate and_gate_h_u_cla32_and5651_y0(h_u_cla32_and5650_y0, h_u_cla32_and5649_y0, h_u_cla32_and5651_y0);
  and_gate and_gate_h_u_cla32_and5652_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5652_y0);
  and_gate and_gate_h_u_cla32_and5653_y0(h_u_cla32_and5652_y0, h_u_cla32_and5651_y0, h_u_cla32_and5653_y0);
  and_gate and_gate_h_u_cla32_and5654_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5654_y0);
  and_gate and_gate_h_u_cla32_and5655_y0(h_u_cla32_and5654_y0, h_u_cla32_and5653_y0, h_u_cla32_and5655_y0);
  and_gate and_gate_h_u_cla32_and5656_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5656_y0);
  and_gate and_gate_h_u_cla32_and5657_y0(h_u_cla32_and5656_y0, h_u_cla32_and5655_y0, h_u_cla32_and5657_y0);
  and_gate and_gate_h_u_cla32_and5658_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5658_y0);
  and_gate and_gate_h_u_cla32_and5659_y0(h_u_cla32_and5658_y0, h_u_cla32_and5657_y0, h_u_cla32_and5659_y0);
  and_gate and_gate_h_u_cla32_and5660_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5660_y0);
  and_gate and_gate_h_u_cla32_and5661_y0(h_u_cla32_and5660_y0, h_u_cla32_and5659_y0, h_u_cla32_and5661_y0);
  and_gate and_gate_h_u_cla32_and5662_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5662_y0);
  and_gate and_gate_h_u_cla32_and5663_y0(h_u_cla32_and5662_y0, h_u_cla32_and5661_y0, h_u_cla32_and5663_y0);
  and_gate and_gate_h_u_cla32_and5664_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5664_y0);
  and_gate and_gate_h_u_cla32_and5665_y0(h_u_cla32_and5664_y0, h_u_cla32_and5663_y0, h_u_cla32_and5665_y0);
  and_gate and_gate_h_u_cla32_and5666_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5666_y0);
  and_gate and_gate_h_u_cla32_and5667_y0(h_u_cla32_and5666_y0, h_u_cla32_and5665_y0, h_u_cla32_and5667_y0);
  and_gate and_gate_h_u_cla32_and5668_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5668_y0);
  and_gate and_gate_h_u_cla32_and5669_y0(h_u_cla32_and5668_y0, h_u_cla32_and5667_y0, h_u_cla32_and5669_y0);
  and_gate and_gate_h_u_cla32_and5670_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and5670_y0);
  and_gate and_gate_h_u_cla32_and5671_y0(h_u_cla32_and5670_y0, h_u_cla32_and5669_y0, h_u_cla32_and5671_y0);
  and_gate and_gate_h_u_cla32_and5672_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5672_y0);
  and_gate and_gate_h_u_cla32_and5673_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5673_y0);
  and_gate and_gate_h_u_cla32_and5674_y0(h_u_cla32_and5673_y0, h_u_cla32_and5672_y0, h_u_cla32_and5674_y0);
  and_gate and_gate_h_u_cla32_and5675_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5675_y0);
  and_gate and_gate_h_u_cla32_and5676_y0(h_u_cla32_and5675_y0, h_u_cla32_and5674_y0, h_u_cla32_and5676_y0);
  and_gate and_gate_h_u_cla32_and5677_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5677_y0);
  and_gate and_gate_h_u_cla32_and5678_y0(h_u_cla32_and5677_y0, h_u_cla32_and5676_y0, h_u_cla32_and5678_y0);
  and_gate and_gate_h_u_cla32_and5679_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5679_y0);
  and_gate and_gate_h_u_cla32_and5680_y0(h_u_cla32_and5679_y0, h_u_cla32_and5678_y0, h_u_cla32_and5680_y0);
  and_gate and_gate_h_u_cla32_and5681_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5681_y0);
  and_gate and_gate_h_u_cla32_and5682_y0(h_u_cla32_and5681_y0, h_u_cla32_and5680_y0, h_u_cla32_and5682_y0);
  and_gate and_gate_h_u_cla32_and5683_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5683_y0);
  and_gate and_gate_h_u_cla32_and5684_y0(h_u_cla32_and5683_y0, h_u_cla32_and5682_y0, h_u_cla32_and5684_y0);
  and_gate and_gate_h_u_cla32_and5685_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5685_y0);
  and_gate and_gate_h_u_cla32_and5686_y0(h_u_cla32_and5685_y0, h_u_cla32_and5684_y0, h_u_cla32_and5686_y0);
  and_gate and_gate_h_u_cla32_and5687_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5687_y0);
  and_gate and_gate_h_u_cla32_and5688_y0(h_u_cla32_and5687_y0, h_u_cla32_and5686_y0, h_u_cla32_and5688_y0);
  and_gate and_gate_h_u_cla32_and5689_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5689_y0);
  and_gate and_gate_h_u_cla32_and5690_y0(h_u_cla32_and5689_y0, h_u_cla32_and5688_y0, h_u_cla32_and5690_y0);
  and_gate and_gate_h_u_cla32_and5691_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5691_y0);
  and_gate and_gate_h_u_cla32_and5692_y0(h_u_cla32_and5691_y0, h_u_cla32_and5690_y0, h_u_cla32_and5692_y0);
  and_gate and_gate_h_u_cla32_and5693_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5693_y0);
  and_gate and_gate_h_u_cla32_and5694_y0(h_u_cla32_and5693_y0, h_u_cla32_and5692_y0, h_u_cla32_and5694_y0);
  and_gate and_gate_h_u_cla32_and5695_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5695_y0);
  and_gate and_gate_h_u_cla32_and5696_y0(h_u_cla32_and5695_y0, h_u_cla32_and5694_y0, h_u_cla32_and5696_y0);
  and_gate and_gate_h_u_cla32_and5697_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5697_y0);
  and_gate and_gate_h_u_cla32_and5698_y0(h_u_cla32_and5697_y0, h_u_cla32_and5696_y0, h_u_cla32_and5698_y0);
  and_gate and_gate_h_u_cla32_and5699_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5699_y0);
  and_gate and_gate_h_u_cla32_and5700_y0(h_u_cla32_and5699_y0, h_u_cla32_and5698_y0, h_u_cla32_and5700_y0);
  and_gate and_gate_h_u_cla32_and5701_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5701_y0);
  and_gate and_gate_h_u_cla32_and5702_y0(h_u_cla32_and5701_y0, h_u_cla32_and5700_y0, h_u_cla32_and5702_y0);
  and_gate and_gate_h_u_cla32_and5703_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5703_y0);
  and_gate and_gate_h_u_cla32_and5704_y0(h_u_cla32_and5703_y0, h_u_cla32_and5702_y0, h_u_cla32_and5704_y0);
  and_gate and_gate_h_u_cla32_and5705_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5705_y0);
  and_gate and_gate_h_u_cla32_and5706_y0(h_u_cla32_and5705_y0, h_u_cla32_and5704_y0, h_u_cla32_and5706_y0);
  and_gate and_gate_h_u_cla32_and5707_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5707_y0);
  and_gate and_gate_h_u_cla32_and5708_y0(h_u_cla32_and5707_y0, h_u_cla32_and5706_y0, h_u_cla32_and5708_y0);
  and_gate and_gate_h_u_cla32_and5709_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5709_y0);
  and_gate and_gate_h_u_cla32_and5710_y0(h_u_cla32_and5709_y0, h_u_cla32_and5708_y0, h_u_cla32_and5710_y0);
  and_gate and_gate_h_u_cla32_and5711_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5711_y0);
  and_gate and_gate_h_u_cla32_and5712_y0(h_u_cla32_and5711_y0, h_u_cla32_and5710_y0, h_u_cla32_and5712_y0);
  and_gate and_gate_h_u_cla32_and5713_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5713_y0);
  and_gate and_gate_h_u_cla32_and5714_y0(h_u_cla32_and5713_y0, h_u_cla32_and5712_y0, h_u_cla32_and5714_y0);
  and_gate and_gate_h_u_cla32_and5715_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and5715_y0);
  and_gate and_gate_h_u_cla32_and5716_y0(h_u_cla32_and5715_y0, h_u_cla32_and5714_y0, h_u_cla32_and5716_y0);
  and_gate and_gate_h_u_cla32_and5717_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5717_y0);
  and_gate and_gate_h_u_cla32_and5718_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5718_y0);
  and_gate and_gate_h_u_cla32_and5719_y0(h_u_cla32_and5718_y0, h_u_cla32_and5717_y0, h_u_cla32_and5719_y0);
  and_gate and_gate_h_u_cla32_and5720_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5720_y0);
  and_gate and_gate_h_u_cla32_and5721_y0(h_u_cla32_and5720_y0, h_u_cla32_and5719_y0, h_u_cla32_and5721_y0);
  and_gate and_gate_h_u_cla32_and5722_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5722_y0);
  and_gate and_gate_h_u_cla32_and5723_y0(h_u_cla32_and5722_y0, h_u_cla32_and5721_y0, h_u_cla32_and5723_y0);
  and_gate and_gate_h_u_cla32_and5724_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5724_y0);
  and_gate and_gate_h_u_cla32_and5725_y0(h_u_cla32_and5724_y0, h_u_cla32_and5723_y0, h_u_cla32_and5725_y0);
  and_gate and_gate_h_u_cla32_and5726_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5726_y0);
  and_gate and_gate_h_u_cla32_and5727_y0(h_u_cla32_and5726_y0, h_u_cla32_and5725_y0, h_u_cla32_and5727_y0);
  and_gate and_gate_h_u_cla32_and5728_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5728_y0);
  and_gate and_gate_h_u_cla32_and5729_y0(h_u_cla32_and5728_y0, h_u_cla32_and5727_y0, h_u_cla32_and5729_y0);
  and_gate and_gate_h_u_cla32_and5730_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5730_y0);
  and_gate and_gate_h_u_cla32_and5731_y0(h_u_cla32_and5730_y0, h_u_cla32_and5729_y0, h_u_cla32_and5731_y0);
  and_gate and_gate_h_u_cla32_and5732_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5732_y0);
  and_gate and_gate_h_u_cla32_and5733_y0(h_u_cla32_and5732_y0, h_u_cla32_and5731_y0, h_u_cla32_and5733_y0);
  and_gate and_gate_h_u_cla32_and5734_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5734_y0);
  and_gate and_gate_h_u_cla32_and5735_y0(h_u_cla32_and5734_y0, h_u_cla32_and5733_y0, h_u_cla32_and5735_y0);
  and_gate and_gate_h_u_cla32_and5736_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5736_y0);
  and_gate and_gate_h_u_cla32_and5737_y0(h_u_cla32_and5736_y0, h_u_cla32_and5735_y0, h_u_cla32_and5737_y0);
  and_gate and_gate_h_u_cla32_and5738_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5738_y0);
  and_gate and_gate_h_u_cla32_and5739_y0(h_u_cla32_and5738_y0, h_u_cla32_and5737_y0, h_u_cla32_and5739_y0);
  and_gate and_gate_h_u_cla32_and5740_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5740_y0);
  and_gate and_gate_h_u_cla32_and5741_y0(h_u_cla32_and5740_y0, h_u_cla32_and5739_y0, h_u_cla32_and5741_y0);
  and_gate and_gate_h_u_cla32_and5742_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5742_y0);
  and_gate and_gate_h_u_cla32_and5743_y0(h_u_cla32_and5742_y0, h_u_cla32_and5741_y0, h_u_cla32_and5743_y0);
  and_gate and_gate_h_u_cla32_and5744_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5744_y0);
  and_gate and_gate_h_u_cla32_and5745_y0(h_u_cla32_and5744_y0, h_u_cla32_and5743_y0, h_u_cla32_and5745_y0);
  and_gate and_gate_h_u_cla32_and5746_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5746_y0);
  and_gate and_gate_h_u_cla32_and5747_y0(h_u_cla32_and5746_y0, h_u_cla32_and5745_y0, h_u_cla32_and5747_y0);
  and_gate and_gate_h_u_cla32_and5748_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5748_y0);
  and_gate and_gate_h_u_cla32_and5749_y0(h_u_cla32_and5748_y0, h_u_cla32_and5747_y0, h_u_cla32_and5749_y0);
  and_gate and_gate_h_u_cla32_and5750_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5750_y0);
  and_gate and_gate_h_u_cla32_and5751_y0(h_u_cla32_and5750_y0, h_u_cla32_and5749_y0, h_u_cla32_and5751_y0);
  and_gate and_gate_h_u_cla32_and5752_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5752_y0);
  and_gate and_gate_h_u_cla32_and5753_y0(h_u_cla32_and5752_y0, h_u_cla32_and5751_y0, h_u_cla32_and5753_y0);
  and_gate and_gate_h_u_cla32_and5754_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5754_y0);
  and_gate and_gate_h_u_cla32_and5755_y0(h_u_cla32_and5754_y0, h_u_cla32_and5753_y0, h_u_cla32_and5755_y0);
  and_gate and_gate_h_u_cla32_and5756_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5756_y0);
  and_gate and_gate_h_u_cla32_and5757_y0(h_u_cla32_and5756_y0, h_u_cla32_and5755_y0, h_u_cla32_and5757_y0);
  and_gate and_gate_h_u_cla32_and5758_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and5758_y0);
  and_gate and_gate_h_u_cla32_and5759_y0(h_u_cla32_and5758_y0, h_u_cla32_and5757_y0, h_u_cla32_and5759_y0);
  and_gate and_gate_h_u_cla32_and5760_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5760_y0);
  and_gate and_gate_h_u_cla32_and5761_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5761_y0);
  and_gate and_gate_h_u_cla32_and5762_y0(h_u_cla32_and5761_y0, h_u_cla32_and5760_y0, h_u_cla32_and5762_y0);
  and_gate and_gate_h_u_cla32_and5763_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5763_y0);
  and_gate and_gate_h_u_cla32_and5764_y0(h_u_cla32_and5763_y0, h_u_cla32_and5762_y0, h_u_cla32_and5764_y0);
  and_gate and_gate_h_u_cla32_and5765_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5765_y0);
  and_gate and_gate_h_u_cla32_and5766_y0(h_u_cla32_and5765_y0, h_u_cla32_and5764_y0, h_u_cla32_and5766_y0);
  and_gate and_gate_h_u_cla32_and5767_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5767_y0);
  and_gate and_gate_h_u_cla32_and5768_y0(h_u_cla32_and5767_y0, h_u_cla32_and5766_y0, h_u_cla32_and5768_y0);
  and_gate and_gate_h_u_cla32_and5769_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5769_y0);
  and_gate and_gate_h_u_cla32_and5770_y0(h_u_cla32_and5769_y0, h_u_cla32_and5768_y0, h_u_cla32_and5770_y0);
  and_gate and_gate_h_u_cla32_and5771_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5771_y0);
  and_gate and_gate_h_u_cla32_and5772_y0(h_u_cla32_and5771_y0, h_u_cla32_and5770_y0, h_u_cla32_and5772_y0);
  and_gate and_gate_h_u_cla32_and5773_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5773_y0);
  and_gate and_gate_h_u_cla32_and5774_y0(h_u_cla32_and5773_y0, h_u_cla32_and5772_y0, h_u_cla32_and5774_y0);
  and_gate and_gate_h_u_cla32_and5775_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5775_y0);
  and_gate and_gate_h_u_cla32_and5776_y0(h_u_cla32_and5775_y0, h_u_cla32_and5774_y0, h_u_cla32_and5776_y0);
  and_gate and_gate_h_u_cla32_and5777_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5777_y0);
  and_gate and_gate_h_u_cla32_and5778_y0(h_u_cla32_and5777_y0, h_u_cla32_and5776_y0, h_u_cla32_and5778_y0);
  and_gate and_gate_h_u_cla32_and5779_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5779_y0);
  and_gate and_gate_h_u_cla32_and5780_y0(h_u_cla32_and5779_y0, h_u_cla32_and5778_y0, h_u_cla32_and5780_y0);
  and_gate and_gate_h_u_cla32_and5781_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5781_y0);
  and_gate and_gate_h_u_cla32_and5782_y0(h_u_cla32_and5781_y0, h_u_cla32_and5780_y0, h_u_cla32_and5782_y0);
  and_gate and_gate_h_u_cla32_and5783_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5783_y0);
  and_gate and_gate_h_u_cla32_and5784_y0(h_u_cla32_and5783_y0, h_u_cla32_and5782_y0, h_u_cla32_and5784_y0);
  and_gate and_gate_h_u_cla32_and5785_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5785_y0);
  and_gate and_gate_h_u_cla32_and5786_y0(h_u_cla32_and5785_y0, h_u_cla32_and5784_y0, h_u_cla32_and5786_y0);
  and_gate and_gate_h_u_cla32_and5787_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5787_y0);
  and_gate and_gate_h_u_cla32_and5788_y0(h_u_cla32_and5787_y0, h_u_cla32_and5786_y0, h_u_cla32_and5788_y0);
  and_gate and_gate_h_u_cla32_and5789_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5789_y0);
  and_gate and_gate_h_u_cla32_and5790_y0(h_u_cla32_and5789_y0, h_u_cla32_and5788_y0, h_u_cla32_and5790_y0);
  and_gate and_gate_h_u_cla32_and5791_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5791_y0);
  and_gate and_gate_h_u_cla32_and5792_y0(h_u_cla32_and5791_y0, h_u_cla32_and5790_y0, h_u_cla32_and5792_y0);
  and_gate and_gate_h_u_cla32_and5793_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5793_y0);
  and_gate and_gate_h_u_cla32_and5794_y0(h_u_cla32_and5793_y0, h_u_cla32_and5792_y0, h_u_cla32_and5794_y0);
  and_gate and_gate_h_u_cla32_and5795_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5795_y0);
  and_gate and_gate_h_u_cla32_and5796_y0(h_u_cla32_and5795_y0, h_u_cla32_and5794_y0, h_u_cla32_and5796_y0);
  and_gate and_gate_h_u_cla32_and5797_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5797_y0);
  and_gate and_gate_h_u_cla32_and5798_y0(h_u_cla32_and5797_y0, h_u_cla32_and5796_y0, h_u_cla32_and5798_y0);
  and_gate and_gate_h_u_cla32_and5799_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and5799_y0);
  and_gate and_gate_h_u_cla32_and5800_y0(h_u_cla32_and5799_y0, h_u_cla32_and5798_y0, h_u_cla32_and5800_y0);
  and_gate and_gate_h_u_cla32_and5801_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5801_y0);
  and_gate and_gate_h_u_cla32_and5802_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5802_y0);
  and_gate and_gate_h_u_cla32_and5803_y0(h_u_cla32_and5802_y0, h_u_cla32_and5801_y0, h_u_cla32_and5803_y0);
  and_gate and_gate_h_u_cla32_and5804_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5804_y0);
  and_gate and_gate_h_u_cla32_and5805_y0(h_u_cla32_and5804_y0, h_u_cla32_and5803_y0, h_u_cla32_and5805_y0);
  and_gate and_gate_h_u_cla32_and5806_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5806_y0);
  and_gate and_gate_h_u_cla32_and5807_y0(h_u_cla32_and5806_y0, h_u_cla32_and5805_y0, h_u_cla32_and5807_y0);
  and_gate and_gate_h_u_cla32_and5808_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5808_y0);
  and_gate and_gate_h_u_cla32_and5809_y0(h_u_cla32_and5808_y0, h_u_cla32_and5807_y0, h_u_cla32_and5809_y0);
  and_gate and_gate_h_u_cla32_and5810_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5810_y0);
  and_gate and_gate_h_u_cla32_and5811_y0(h_u_cla32_and5810_y0, h_u_cla32_and5809_y0, h_u_cla32_and5811_y0);
  and_gate and_gate_h_u_cla32_and5812_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5812_y0);
  and_gate and_gate_h_u_cla32_and5813_y0(h_u_cla32_and5812_y0, h_u_cla32_and5811_y0, h_u_cla32_and5813_y0);
  and_gate and_gate_h_u_cla32_and5814_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5814_y0);
  and_gate and_gate_h_u_cla32_and5815_y0(h_u_cla32_and5814_y0, h_u_cla32_and5813_y0, h_u_cla32_and5815_y0);
  and_gate and_gate_h_u_cla32_and5816_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5816_y0);
  and_gate and_gate_h_u_cla32_and5817_y0(h_u_cla32_and5816_y0, h_u_cla32_and5815_y0, h_u_cla32_and5817_y0);
  and_gate and_gate_h_u_cla32_and5818_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5818_y0);
  and_gate and_gate_h_u_cla32_and5819_y0(h_u_cla32_and5818_y0, h_u_cla32_and5817_y0, h_u_cla32_and5819_y0);
  and_gate and_gate_h_u_cla32_and5820_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5820_y0);
  and_gate and_gate_h_u_cla32_and5821_y0(h_u_cla32_and5820_y0, h_u_cla32_and5819_y0, h_u_cla32_and5821_y0);
  and_gate and_gate_h_u_cla32_and5822_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5822_y0);
  and_gate and_gate_h_u_cla32_and5823_y0(h_u_cla32_and5822_y0, h_u_cla32_and5821_y0, h_u_cla32_and5823_y0);
  and_gate and_gate_h_u_cla32_and5824_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5824_y0);
  and_gate and_gate_h_u_cla32_and5825_y0(h_u_cla32_and5824_y0, h_u_cla32_and5823_y0, h_u_cla32_and5825_y0);
  and_gate and_gate_h_u_cla32_and5826_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5826_y0);
  and_gate and_gate_h_u_cla32_and5827_y0(h_u_cla32_and5826_y0, h_u_cla32_and5825_y0, h_u_cla32_and5827_y0);
  and_gate and_gate_h_u_cla32_and5828_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5828_y0);
  and_gate and_gate_h_u_cla32_and5829_y0(h_u_cla32_and5828_y0, h_u_cla32_and5827_y0, h_u_cla32_and5829_y0);
  and_gate and_gate_h_u_cla32_and5830_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5830_y0);
  and_gate and_gate_h_u_cla32_and5831_y0(h_u_cla32_and5830_y0, h_u_cla32_and5829_y0, h_u_cla32_and5831_y0);
  and_gate and_gate_h_u_cla32_and5832_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5832_y0);
  and_gate and_gate_h_u_cla32_and5833_y0(h_u_cla32_and5832_y0, h_u_cla32_and5831_y0, h_u_cla32_and5833_y0);
  and_gate and_gate_h_u_cla32_and5834_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5834_y0);
  and_gate and_gate_h_u_cla32_and5835_y0(h_u_cla32_and5834_y0, h_u_cla32_and5833_y0, h_u_cla32_and5835_y0);
  and_gate and_gate_h_u_cla32_and5836_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5836_y0);
  and_gate and_gate_h_u_cla32_and5837_y0(h_u_cla32_and5836_y0, h_u_cla32_and5835_y0, h_u_cla32_and5837_y0);
  and_gate and_gate_h_u_cla32_and5838_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and5838_y0);
  and_gate and_gate_h_u_cla32_and5839_y0(h_u_cla32_and5838_y0, h_u_cla32_and5837_y0, h_u_cla32_and5839_y0);
  and_gate and_gate_h_u_cla32_and5840_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5840_y0);
  and_gate and_gate_h_u_cla32_and5841_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5841_y0);
  and_gate and_gate_h_u_cla32_and5842_y0(h_u_cla32_and5841_y0, h_u_cla32_and5840_y0, h_u_cla32_and5842_y0);
  and_gate and_gate_h_u_cla32_and5843_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5843_y0);
  and_gate and_gate_h_u_cla32_and5844_y0(h_u_cla32_and5843_y0, h_u_cla32_and5842_y0, h_u_cla32_and5844_y0);
  and_gate and_gate_h_u_cla32_and5845_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5845_y0);
  and_gate and_gate_h_u_cla32_and5846_y0(h_u_cla32_and5845_y0, h_u_cla32_and5844_y0, h_u_cla32_and5846_y0);
  and_gate and_gate_h_u_cla32_and5847_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5847_y0);
  and_gate and_gate_h_u_cla32_and5848_y0(h_u_cla32_and5847_y0, h_u_cla32_and5846_y0, h_u_cla32_and5848_y0);
  and_gate and_gate_h_u_cla32_and5849_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5849_y0);
  and_gate and_gate_h_u_cla32_and5850_y0(h_u_cla32_and5849_y0, h_u_cla32_and5848_y0, h_u_cla32_and5850_y0);
  and_gate and_gate_h_u_cla32_and5851_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5851_y0);
  and_gate and_gate_h_u_cla32_and5852_y0(h_u_cla32_and5851_y0, h_u_cla32_and5850_y0, h_u_cla32_and5852_y0);
  and_gate and_gate_h_u_cla32_and5853_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5853_y0);
  and_gate and_gate_h_u_cla32_and5854_y0(h_u_cla32_and5853_y0, h_u_cla32_and5852_y0, h_u_cla32_and5854_y0);
  and_gate and_gate_h_u_cla32_and5855_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5855_y0);
  and_gate and_gate_h_u_cla32_and5856_y0(h_u_cla32_and5855_y0, h_u_cla32_and5854_y0, h_u_cla32_and5856_y0);
  and_gate and_gate_h_u_cla32_and5857_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5857_y0);
  and_gate and_gate_h_u_cla32_and5858_y0(h_u_cla32_and5857_y0, h_u_cla32_and5856_y0, h_u_cla32_and5858_y0);
  and_gate and_gate_h_u_cla32_and5859_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5859_y0);
  and_gate and_gate_h_u_cla32_and5860_y0(h_u_cla32_and5859_y0, h_u_cla32_and5858_y0, h_u_cla32_and5860_y0);
  and_gate and_gate_h_u_cla32_and5861_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5861_y0);
  and_gate and_gate_h_u_cla32_and5862_y0(h_u_cla32_and5861_y0, h_u_cla32_and5860_y0, h_u_cla32_and5862_y0);
  and_gate and_gate_h_u_cla32_and5863_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5863_y0);
  and_gate and_gate_h_u_cla32_and5864_y0(h_u_cla32_and5863_y0, h_u_cla32_and5862_y0, h_u_cla32_and5864_y0);
  and_gate and_gate_h_u_cla32_and5865_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5865_y0);
  and_gate and_gate_h_u_cla32_and5866_y0(h_u_cla32_and5865_y0, h_u_cla32_and5864_y0, h_u_cla32_and5866_y0);
  and_gate and_gate_h_u_cla32_and5867_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5867_y0);
  and_gate and_gate_h_u_cla32_and5868_y0(h_u_cla32_and5867_y0, h_u_cla32_and5866_y0, h_u_cla32_and5868_y0);
  and_gate and_gate_h_u_cla32_and5869_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5869_y0);
  and_gate and_gate_h_u_cla32_and5870_y0(h_u_cla32_and5869_y0, h_u_cla32_and5868_y0, h_u_cla32_and5870_y0);
  and_gate and_gate_h_u_cla32_and5871_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5871_y0);
  and_gate and_gate_h_u_cla32_and5872_y0(h_u_cla32_and5871_y0, h_u_cla32_and5870_y0, h_u_cla32_and5872_y0);
  and_gate and_gate_h_u_cla32_and5873_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5873_y0);
  and_gate and_gate_h_u_cla32_and5874_y0(h_u_cla32_and5873_y0, h_u_cla32_and5872_y0, h_u_cla32_and5874_y0);
  and_gate and_gate_h_u_cla32_and5875_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and5875_y0);
  and_gate and_gate_h_u_cla32_and5876_y0(h_u_cla32_and5875_y0, h_u_cla32_and5874_y0, h_u_cla32_and5876_y0);
  and_gate and_gate_h_u_cla32_and5877_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5877_y0);
  and_gate and_gate_h_u_cla32_and5878_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5878_y0);
  and_gate and_gate_h_u_cla32_and5879_y0(h_u_cla32_and5878_y0, h_u_cla32_and5877_y0, h_u_cla32_and5879_y0);
  and_gate and_gate_h_u_cla32_and5880_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5880_y0);
  and_gate and_gate_h_u_cla32_and5881_y0(h_u_cla32_and5880_y0, h_u_cla32_and5879_y0, h_u_cla32_and5881_y0);
  and_gate and_gate_h_u_cla32_and5882_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5882_y0);
  and_gate and_gate_h_u_cla32_and5883_y0(h_u_cla32_and5882_y0, h_u_cla32_and5881_y0, h_u_cla32_and5883_y0);
  and_gate and_gate_h_u_cla32_and5884_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5884_y0);
  and_gate and_gate_h_u_cla32_and5885_y0(h_u_cla32_and5884_y0, h_u_cla32_and5883_y0, h_u_cla32_and5885_y0);
  and_gate and_gate_h_u_cla32_and5886_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5886_y0);
  and_gate and_gate_h_u_cla32_and5887_y0(h_u_cla32_and5886_y0, h_u_cla32_and5885_y0, h_u_cla32_and5887_y0);
  and_gate and_gate_h_u_cla32_and5888_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5888_y0);
  and_gate and_gate_h_u_cla32_and5889_y0(h_u_cla32_and5888_y0, h_u_cla32_and5887_y0, h_u_cla32_and5889_y0);
  and_gate and_gate_h_u_cla32_and5890_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5890_y0);
  and_gate and_gate_h_u_cla32_and5891_y0(h_u_cla32_and5890_y0, h_u_cla32_and5889_y0, h_u_cla32_and5891_y0);
  and_gate and_gate_h_u_cla32_and5892_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5892_y0);
  and_gate and_gate_h_u_cla32_and5893_y0(h_u_cla32_and5892_y0, h_u_cla32_and5891_y0, h_u_cla32_and5893_y0);
  and_gate and_gate_h_u_cla32_and5894_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5894_y0);
  and_gate and_gate_h_u_cla32_and5895_y0(h_u_cla32_and5894_y0, h_u_cla32_and5893_y0, h_u_cla32_and5895_y0);
  and_gate and_gate_h_u_cla32_and5896_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5896_y0);
  and_gate and_gate_h_u_cla32_and5897_y0(h_u_cla32_and5896_y0, h_u_cla32_and5895_y0, h_u_cla32_and5897_y0);
  and_gate and_gate_h_u_cla32_and5898_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5898_y0);
  and_gate and_gate_h_u_cla32_and5899_y0(h_u_cla32_and5898_y0, h_u_cla32_and5897_y0, h_u_cla32_and5899_y0);
  and_gate and_gate_h_u_cla32_and5900_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5900_y0);
  and_gate and_gate_h_u_cla32_and5901_y0(h_u_cla32_and5900_y0, h_u_cla32_and5899_y0, h_u_cla32_and5901_y0);
  and_gate and_gate_h_u_cla32_and5902_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5902_y0);
  and_gate and_gate_h_u_cla32_and5903_y0(h_u_cla32_and5902_y0, h_u_cla32_and5901_y0, h_u_cla32_and5903_y0);
  and_gate and_gate_h_u_cla32_and5904_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5904_y0);
  and_gate and_gate_h_u_cla32_and5905_y0(h_u_cla32_and5904_y0, h_u_cla32_and5903_y0, h_u_cla32_and5905_y0);
  and_gate and_gate_h_u_cla32_and5906_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5906_y0);
  and_gate and_gate_h_u_cla32_and5907_y0(h_u_cla32_and5906_y0, h_u_cla32_and5905_y0, h_u_cla32_and5907_y0);
  and_gate and_gate_h_u_cla32_and5908_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5908_y0);
  and_gate and_gate_h_u_cla32_and5909_y0(h_u_cla32_and5908_y0, h_u_cla32_and5907_y0, h_u_cla32_and5909_y0);
  and_gate and_gate_h_u_cla32_and5910_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and5910_y0);
  and_gate and_gate_h_u_cla32_and5911_y0(h_u_cla32_and5910_y0, h_u_cla32_and5909_y0, h_u_cla32_and5911_y0);
  and_gate and_gate_h_u_cla32_and5912_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5912_y0);
  and_gate and_gate_h_u_cla32_and5913_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5913_y0);
  and_gate and_gate_h_u_cla32_and5914_y0(h_u_cla32_and5913_y0, h_u_cla32_and5912_y0, h_u_cla32_and5914_y0);
  and_gate and_gate_h_u_cla32_and5915_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5915_y0);
  and_gate and_gate_h_u_cla32_and5916_y0(h_u_cla32_and5915_y0, h_u_cla32_and5914_y0, h_u_cla32_and5916_y0);
  and_gate and_gate_h_u_cla32_and5917_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5917_y0);
  and_gate and_gate_h_u_cla32_and5918_y0(h_u_cla32_and5917_y0, h_u_cla32_and5916_y0, h_u_cla32_and5918_y0);
  and_gate and_gate_h_u_cla32_and5919_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5919_y0);
  and_gate and_gate_h_u_cla32_and5920_y0(h_u_cla32_and5919_y0, h_u_cla32_and5918_y0, h_u_cla32_and5920_y0);
  and_gate and_gate_h_u_cla32_and5921_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5921_y0);
  and_gate and_gate_h_u_cla32_and5922_y0(h_u_cla32_and5921_y0, h_u_cla32_and5920_y0, h_u_cla32_and5922_y0);
  and_gate and_gate_h_u_cla32_and5923_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5923_y0);
  and_gate and_gate_h_u_cla32_and5924_y0(h_u_cla32_and5923_y0, h_u_cla32_and5922_y0, h_u_cla32_and5924_y0);
  and_gate and_gate_h_u_cla32_and5925_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5925_y0);
  and_gate and_gate_h_u_cla32_and5926_y0(h_u_cla32_and5925_y0, h_u_cla32_and5924_y0, h_u_cla32_and5926_y0);
  and_gate and_gate_h_u_cla32_and5927_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5927_y0);
  and_gate and_gate_h_u_cla32_and5928_y0(h_u_cla32_and5927_y0, h_u_cla32_and5926_y0, h_u_cla32_and5928_y0);
  and_gate and_gate_h_u_cla32_and5929_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5929_y0);
  and_gate and_gate_h_u_cla32_and5930_y0(h_u_cla32_and5929_y0, h_u_cla32_and5928_y0, h_u_cla32_and5930_y0);
  and_gate and_gate_h_u_cla32_and5931_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5931_y0);
  and_gate and_gate_h_u_cla32_and5932_y0(h_u_cla32_and5931_y0, h_u_cla32_and5930_y0, h_u_cla32_and5932_y0);
  and_gate and_gate_h_u_cla32_and5933_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5933_y0);
  and_gate and_gate_h_u_cla32_and5934_y0(h_u_cla32_and5933_y0, h_u_cla32_and5932_y0, h_u_cla32_and5934_y0);
  and_gate and_gate_h_u_cla32_and5935_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5935_y0);
  and_gate and_gate_h_u_cla32_and5936_y0(h_u_cla32_and5935_y0, h_u_cla32_and5934_y0, h_u_cla32_and5936_y0);
  and_gate and_gate_h_u_cla32_and5937_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5937_y0);
  and_gate and_gate_h_u_cla32_and5938_y0(h_u_cla32_and5937_y0, h_u_cla32_and5936_y0, h_u_cla32_and5938_y0);
  and_gate and_gate_h_u_cla32_and5939_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5939_y0);
  and_gate and_gate_h_u_cla32_and5940_y0(h_u_cla32_and5939_y0, h_u_cla32_and5938_y0, h_u_cla32_and5940_y0);
  and_gate and_gate_h_u_cla32_and5941_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5941_y0);
  and_gate and_gate_h_u_cla32_and5942_y0(h_u_cla32_and5941_y0, h_u_cla32_and5940_y0, h_u_cla32_and5942_y0);
  and_gate and_gate_h_u_cla32_and5943_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and5943_y0);
  and_gate and_gate_h_u_cla32_and5944_y0(h_u_cla32_and5943_y0, h_u_cla32_and5942_y0, h_u_cla32_and5944_y0);
  and_gate and_gate_h_u_cla32_and5945_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5945_y0);
  and_gate and_gate_h_u_cla32_and5946_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5946_y0);
  and_gate and_gate_h_u_cla32_and5947_y0(h_u_cla32_and5946_y0, h_u_cla32_and5945_y0, h_u_cla32_and5947_y0);
  and_gate and_gate_h_u_cla32_and5948_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5948_y0);
  and_gate and_gate_h_u_cla32_and5949_y0(h_u_cla32_and5948_y0, h_u_cla32_and5947_y0, h_u_cla32_and5949_y0);
  and_gate and_gate_h_u_cla32_and5950_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5950_y0);
  and_gate and_gate_h_u_cla32_and5951_y0(h_u_cla32_and5950_y0, h_u_cla32_and5949_y0, h_u_cla32_and5951_y0);
  and_gate and_gate_h_u_cla32_and5952_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5952_y0);
  and_gate and_gate_h_u_cla32_and5953_y0(h_u_cla32_and5952_y0, h_u_cla32_and5951_y0, h_u_cla32_and5953_y0);
  and_gate and_gate_h_u_cla32_and5954_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5954_y0);
  and_gate and_gate_h_u_cla32_and5955_y0(h_u_cla32_and5954_y0, h_u_cla32_and5953_y0, h_u_cla32_and5955_y0);
  and_gate and_gate_h_u_cla32_and5956_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5956_y0);
  and_gate and_gate_h_u_cla32_and5957_y0(h_u_cla32_and5956_y0, h_u_cla32_and5955_y0, h_u_cla32_and5957_y0);
  and_gate and_gate_h_u_cla32_and5958_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5958_y0);
  and_gate and_gate_h_u_cla32_and5959_y0(h_u_cla32_and5958_y0, h_u_cla32_and5957_y0, h_u_cla32_and5959_y0);
  and_gate and_gate_h_u_cla32_and5960_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5960_y0);
  and_gate and_gate_h_u_cla32_and5961_y0(h_u_cla32_and5960_y0, h_u_cla32_and5959_y0, h_u_cla32_and5961_y0);
  and_gate and_gate_h_u_cla32_and5962_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5962_y0);
  and_gate and_gate_h_u_cla32_and5963_y0(h_u_cla32_and5962_y0, h_u_cla32_and5961_y0, h_u_cla32_and5963_y0);
  and_gate and_gate_h_u_cla32_and5964_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5964_y0);
  and_gate and_gate_h_u_cla32_and5965_y0(h_u_cla32_and5964_y0, h_u_cla32_and5963_y0, h_u_cla32_and5965_y0);
  and_gate and_gate_h_u_cla32_and5966_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5966_y0);
  and_gate and_gate_h_u_cla32_and5967_y0(h_u_cla32_and5966_y0, h_u_cla32_and5965_y0, h_u_cla32_and5967_y0);
  and_gate and_gate_h_u_cla32_and5968_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5968_y0);
  and_gate and_gate_h_u_cla32_and5969_y0(h_u_cla32_and5968_y0, h_u_cla32_and5967_y0, h_u_cla32_and5969_y0);
  and_gate and_gate_h_u_cla32_and5970_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5970_y0);
  and_gate and_gate_h_u_cla32_and5971_y0(h_u_cla32_and5970_y0, h_u_cla32_and5969_y0, h_u_cla32_and5971_y0);
  and_gate and_gate_h_u_cla32_and5972_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5972_y0);
  and_gate and_gate_h_u_cla32_and5973_y0(h_u_cla32_and5972_y0, h_u_cla32_and5971_y0, h_u_cla32_and5973_y0);
  and_gate and_gate_h_u_cla32_and5974_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and5974_y0);
  and_gate and_gate_h_u_cla32_and5975_y0(h_u_cla32_and5974_y0, h_u_cla32_and5973_y0, h_u_cla32_and5975_y0);
  and_gate and_gate_h_u_cla32_and5976_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5976_y0);
  and_gate and_gate_h_u_cla32_and5977_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5977_y0);
  and_gate and_gate_h_u_cla32_and5978_y0(h_u_cla32_and5977_y0, h_u_cla32_and5976_y0, h_u_cla32_and5978_y0);
  and_gate and_gate_h_u_cla32_and5979_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5979_y0);
  and_gate and_gate_h_u_cla32_and5980_y0(h_u_cla32_and5979_y0, h_u_cla32_and5978_y0, h_u_cla32_and5980_y0);
  and_gate and_gate_h_u_cla32_and5981_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5981_y0);
  and_gate and_gate_h_u_cla32_and5982_y0(h_u_cla32_and5981_y0, h_u_cla32_and5980_y0, h_u_cla32_and5982_y0);
  and_gate and_gate_h_u_cla32_and5983_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5983_y0);
  and_gate and_gate_h_u_cla32_and5984_y0(h_u_cla32_and5983_y0, h_u_cla32_and5982_y0, h_u_cla32_and5984_y0);
  and_gate and_gate_h_u_cla32_and5985_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5985_y0);
  and_gate and_gate_h_u_cla32_and5986_y0(h_u_cla32_and5985_y0, h_u_cla32_and5984_y0, h_u_cla32_and5986_y0);
  and_gate and_gate_h_u_cla32_and5987_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5987_y0);
  and_gate and_gate_h_u_cla32_and5988_y0(h_u_cla32_and5987_y0, h_u_cla32_and5986_y0, h_u_cla32_and5988_y0);
  and_gate and_gate_h_u_cla32_and5989_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5989_y0);
  and_gate and_gate_h_u_cla32_and5990_y0(h_u_cla32_and5989_y0, h_u_cla32_and5988_y0, h_u_cla32_and5990_y0);
  and_gate and_gate_h_u_cla32_and5991_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5991_y0);
  and_gate and_gate_h_u_cla32_and5992_y0(h_u_cla32_and5991_y0, h_u_cla32_and5990_y0, h_u_cla32_and5992_y0);
  and_gate and_gate_h_u_cla32_and5993_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5993_y0);
  and_gate and_gate_h_u_cla32_and5994_y0(h_u_cla32_and5993_y0, h_u_cla32_and5992_y0, h_u_cla32_and5994_y0);
  and_gate and_gate_h_u_cla32_and5995_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5995_y0);
  and_gate and_gate_h_u_cla32_and5996_y0(h_u_cla32_and5995_y0, h_u_cla32_and5994_y0, h_u_cla32_and5996_y0);
  and_gate and_gate_h_u_cla32_and5997_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5997_y0);
  and_gate and_gate_h_u_cla32_and5998_y0(h_u_cla32_and5997_y0, h_u_cla32_and5996_y0, h_u_cla32_and5998_y0);
  and_gate and_gate_h_u_cla32_and5999_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and5999_y0);
  and_gate and_gate_h_u_cla32_and6000_y0(h_u_cla32_and5999_y0, h_u_cla32_and5998_y0, h_u_cla32_and6000_y0);
  and_gate and_gate_h_u_cla32_and6001_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6001_y0);
  and_gate and_gate_h_u_cla32_and6002_y0(h_u_cla32_and6001_y0, h_u_cla32_and6000_y0, h_u_cla32_and6002_y0);
  and_gate and_gate_h_u_cla32_and6003_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6003_y0);
  and_gate and_gate_h_u_cla32_and6004_y0(h_u_cla32_and6003_y0, h_u_cla32_and6002_y0, h_u_cla32_and6004_y0);
  and_gate and_gate_h_u_cla32_and6005_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6005_y0);
  and_gate and_gate_h_u_cla32_and6006_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6006_y0);
  and_gate and_gate_h_u_cla32_and6007_y0(h_u_cla32_and6006_y0, h_u_cla32_and6005_y0, h_u_cla32_and6007_y0);
  and_gate and_gate_h_u_cla32_and6008_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6008_y0);
  and_gate and_gate_h_u_cla32_and6009_y0(h_u_cla32_and6008_y0, h_u_cla32_and6007_y0, h_u_cla32_and6009_y0);
  and_gate and_gate_h_u_cla32_and6010_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6010_y0);
  and_gate and_gate_h_u_cla32_and6011_y0(h_u_cla32_and6010_y0, h_u_cla32_and6009_y0, h_u_cla32_and6011_y0);
  and_gate and_gate_h_u_cla32_and6012_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6012_y0);
  and_gate and_gate_h_u_cla32_and6013_y0(h_u_cla32_and6012_y0, h_u_cla32_and6011_y0, h_u_cla32_and6013_y0);
  and_gate and_gate_h_u_cla32_and6014_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6014_y0);
  and_gate and_gate_h_u_cla32_and6015_y0(h_u_cla32_and6014_y0, h_u_cla32_and6013_y0, h_u_cla32_and6015_y0);
  and_gate and_gate_h_u_cla32_and6016_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6016_y0);
  and_gate and_gate_h_u_cla32_and6017_y0(h_u_cla32_and6016_y0, h_u_cla32_and6015_y0, h_u_cla32_and6017_y0);
  and_gate and_gate_h_u_cla32_and6018_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6018_y0);
  and_gate and_gate_h_u_cla32_and6019_y0(h_u_cla32_and6018_y0, h_u_cla32_and6017_y0, h_u_cla32_and6019_y0);
  and_gate and_gate_h_u_cla32_and6020_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6020_y0);
  and_gate and_gate_h_u_cla32_and6021_y0(h_u_cla32_and6020_y0, h_u_cla32_and6019_y0, h_u_cla32_and6021_y0);
  and_gate and_gate_h_u_cla32_and6022_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6022_y0);
  and_gate and_gate_h_u_cla32_and6023_y0(h_u_cla32_and6022_y0, h_u_cla32_and6021_y0, h_u_cla32_and6023_y0);
  and_gate and_gate_h_u_cla32_and6024_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6024_y0);
  and_gate and_gate_h_u_cla32_and6025_y0(h_u_cla32_and6024_y0, h_u_cla32_and6023_y0, h_u_cla32_and6025_y0);
  and_gate and_gate_h_u_cla32_and6026_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6026_y0);
  and_gate and_gate_h_u_cla32_and6027_y0(h_u_cla32_and6026_y0, h_u_cla32_and6025_y0, h_u_cla32_and6027_y0);
  and_gate and_gate_h_u_cla32_and6028_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6028_y0);
  and_gate and_gate_h_u_cla32_and6029_y0(h_u_cla32_and6028_y0, h_u_cla32_and6027_y0, h_u_cla32_and6029_y0);
  and_gate and_gate_h_u_cla32_and6030_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6030_y0);
  and_gate and_gate_h_u_cla32_and6031_y0(h_u_cla32_and6030_y0, h_u_cla32_and6029_y0, h_u_cla32_and6031_y0);
  and_gate and_gate_h_u_cla32_and6032_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6032_y0);
  and_gate and_gate_h_u_cla32_and6033_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6033_y0);
  and_gate and_gate_h_u_cla32_and6034_y0(h_u_cla32_and6033_y0, h_u_cla32_and6032_y0, h_u_cla32_and6034_y0);
  and_gate and_gate_h_u_cla32_and6035_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6035_y0);
  and_gate and_gate_h_u_cla32_and6036_y0(h_u_cla32_and6035_y0, h_u_cla32_and6034_y0, h_u_cla32_and6036_y0);
  and_gate and_gate_h_u_cla32_and6037_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6037_y0);
  and_gate and_gate_h_u_cla32_and6038_y0(h_u_cla32_and6037_y0, h_u_cla32_and6036_y0, h_u_cla32_and6038_y0);
  and_gate and_gate_h_u_cla32_and6039_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6039_y0);
  and_gate and_gate_h_u_cla32_and6040_y0(h_u_cla32_and6039_y0, h_u_cla32_and6038_y0, h_u_cla32_and6040_y0);
  and_gate and_gate_h_u_cla32_and6041_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6041_y0);
  and_gate and_gate_h_u_cla32_and6042_y0(h_u_cla32_and6041_y0, h_u_cla32_and6040_y0, h_u_cla32_and6042_y0);
  and_gate and_gate_h_u_cla32_and6043_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6043_y0);
  and_gate and_gate_h_u_cla32_and6044_y0(h_u_cla32_and6043_y0, h_u_cla32_and6042_y0, h_u_cla32_and6044_y0);
  and_gate and_gate_h_u_cla32_and6045_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6045_y0);
  and_gate and_gate_h_u_cla32_and6046_y0(h_u_cla32_and6045_y0, h_u_cla32_and6044_y0, h_u_cla32_and6046_y0);
  and_gate and_gate_h_u_cla32_and6047_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6047_y0);
  and_gate and_gate_h_u_cla32_and6048_y0(h_u_cla32_and6047_y0, h_u_cla32_and6046_y0, h_u_cla32_and6048_y0);
  and_gate and_gate_h_u_cla32_and6049_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6049_y0);
  and_gate and_gate_h_u_cla32_and6050_y0(h_u_cla32_and6049_y0, h_u_cla32_and6048_y0, h_u_cla32_and6050_y0);
  and_gate and_gate_h_u_cla32_and6051_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6051_y0);
  and_gate and_gate_h_u_cla32_and6052_y0(h_u_cla32_and6051_y0, h_u_cla32_and6050_y0, h_u_cla32_and6052_y0);
  and_gate and_gate_h_u_cla32_and6053_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6053_y0);
  and_gate and_gate_h_u_cla32_and6054_y0(h_u_cla32_and6053_y0, h_u_cla32_and6052_y0, h_u_cla32_and6054_y0);
  and_gate and_gate_h_u_cla32_and6055_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6055_y0);
  and_gate and_gate_h_u_cla32_and6056_y0(h_u_cla32_and6055_y0, h_u_cla32_and6054_y0, h_u_cla32_and6056_y0);
  and_gate and_gate_h_u_cla32_and6057_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6057_y0);
  and_gate and_gate_h_u_cla32_and6058_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6058_y0);
  and_gate and_gate_h_u_cla32_and6059_y0(h_u_cla32_and6058_y0, h_u_cla32_and6057_y0, h_u_cla32_and6059_y0);
  and_gate and_gate_h_u_cla32_and6060_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6060_y0);
  and_gate and_gate_h_u_cla32_and6061_y0(h_u_cla32_and6060_y0, h_u_cla32_and6059_y0, h_u_cla32_and6061_y0);
  and_gate and_gate_h_u_cla32_and6062_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6062_y0);
  and_gate and_gate_h_u_cla32_and6063_y0(h_u_cla32_and6062_y0, h_u_cla32_and6061_y0, h_u_cla32_and6063_y0);
  and_gate and_gate_h_u_cla32_and6064_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6064_y0);
  and_gate and_gate_h_u_cla32_and6065_y0(h_u_cla32_and6064_y0, h_u_cla32_and6063_y0, h_u_cla32_and6065_y0);
  and_gate and_gate_h_u_cla32_and6066_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6066_y0);
  and_gate and_gate_h_u_cla32_and6067_y0(h_u_cla32_and6066_y0, h_u_cla32_and6065_y0, h_u_cla32_and6067_y0);
  and_gate and_gate_h_u_cla32_and6068_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6068_y0);
  and_gate and_gate_h_u_cla32_and6069_y0(h_u_cla32_and6068_y0, h_u_cla32_and6067_y0, h_u_cla32_and6069_y0);
  and_gate and_gate_h_u_cla32_and6070_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6070_y0);
  and_gate and_gate_h_u_cla32_and6071_y0(h_u_cla32_and6070_y0, h_u_cla32_and6069_y0, h_u_cla32_and6071_y0);
  and_gate and_gate_h_u_cla32_and6072_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6072_y0);
  and_gate and_gate_h_u_cla32_and6073_y0(h_u_cla32_and6072_y0, h_u_cla32_and6071_y0, h_u_cla32_and6073_y0);
  and_gate and_gate_h_u_cla32_and6074_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6074_y0);
  and_gate and_gate_h_u_cla32_and6075_y0(h_u_cla32_and6074_y0, h_u_cla32_and6073_y0, h_u_cla32_and6075_y0);
  and_gate and_gate_h_u_cla32_and6076_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6076_y0);
  and_gate and_gate_h_u_cla32_and6077_y0(h_u_cla32_and6076_y0, h_u_cla32_and6075_y0, h_u_cla32_and6077_y0);
  and_gate and_gate_h_u_cla32_and6078_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6078_y0);
  and_gate and_gate_h_u_cla32_and6079_y0(h_u_cla32_and6078_y0, h_u_cla32_and6077_y0, h_u_cla32_and6079_y0);
  and_gate and_gate_h_u_cla32_and6080_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6080_y0);
  and_gate and_gate_h_u_cla32_and6081_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6081_y0);
  and_gate and_gate_h_u_cla32_and6082_y0(h_u_cla32_and6081_y0, h_u_cla32_and6080_y0, h_u_cla32_and6082_y0);
  and_gate and_gate_h_u_cla32_and6083_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6083_y0);
  and_gate and_gate_h_u_cla32_and6084_y0(h_u_cla32_and6083_y0, h_u_cla32_and6082_y0, h_u_cla32_and6084_y0);
  and_gate and_gate_h_u_cla32_and6085_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6085_y0);
  and_gate and_gate_h_u_cla32_and6086_y0(h_u_cla32_and6085_y0, h_u_cla32_and6084_y0, h_u_cla32_and6086_y0);
  and_gate and_gate_h_u_cla32_and6087_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6087_y0);
  and_gate and_gate_h_u_cla32_and6088_y0(h_u_cla32_and6087_y0, h_u_cla32_and6086_y0, h_u_cla32_and6088_y0);
  and_gate and_gate_h_u_cla32_and6089_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6089_y0);
  and_gate and_gate_h_u_cla32_and6090_y0(h_u_cla32_and6089_y0, h_u_cla32_and6088_y0, h_u_cla32_and6090_y0);
  and_gate and_gate_h_u_cla32_and6091_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6091_y0);
  and_gate and_gate_h_u_cla32_and6092_y0(h_u_cla32_and6091_y0, h_u_cla32_and6090_y0, h_u_cla32_and6092_y0);
  and_gate and_gate_h_u_cla32_and6093_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6093_y0);
  and_gate and_gate_h_u_cla32_and6094_y0(h_u_cla32_and6093_y0, h_u_cla32_and6092_y0, h_u_cla32_and6094_y0);
  and_gate and_gate_h_u_cla32_and6095_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6095_y0);
  and_gate and_gate_h_u_cla32_and6096_y0(h_u_cla32_and6095_y0, h_u_cla32_and6094_y0, h_u_cla32_and6096_y0);
  and_gate and_gate_h_u_cla32_and6097_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6097_y0);
  and_gate and_gate_h_u_cla32_and6098_y0(h_u_cla32_and6097_y0, h_u_cla32_and6096_y0, h_u_cla32_and6098_y0);
  and_gate and_gate_h_u_cla32_and6099_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6099_y0);
  and_gate and_gate_h_u_cla32_and6100_y0(h_u_cla32_and6099_y0, h_u_cla32_and6098_y0, h_u_cla32_and6100_y0);
  and_gate and_gate_h_u_cla32_and6101_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6101_y0);
  and_gate and_gate_h_u_cla32_and6102_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6102_y0);
  and_gate and_gate_h_u_cla32_and6103_y0(h_u_cla32_and6102_y0, h_u_cla32_and6101_y0, h_u_cla32_and6103_y0);
  and_gate and_gate_h_u_cla32_and6104_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6104_y0);
  and_gate and_gate_h_u_cla32_and6105_y0(h_u_cla32_and6104_y0, h_u_cla32_and6103_y0, h_u_cla32_and6105_y0);
  and_gate and_gate_h_u_cla32_and6106_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6106_y0);
  and_gate and_gate_h_u_cla32_and6107_y0(h_u_cla32_and6106_y0, h_u_cla32_and6105_y0, h_u_cla32_and6107_y0);
  and_gate and_gate_h_u_cla32_and6108_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6108_y0);
  and_gate and_gate_h_u_cla32_and6109_y0(h_u_cla32_and6108_y0, h_u_cla32_and6107_y0, h_u_cla32_and6109_y0);
  and_gate and_gate_h_u_cla32_and6110_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6110_y0);
  and_gate and_gate_h_u_cla32_and6111_y0(h_u_cla32_and6110_y0, h_u_cla32_and6109_y0, h_u_cla32_and6111_y0);
  and_gate and_gate_h_u_cla32_and6112_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6112_y0);
  and_gate and_gate_h_u_cla32_and6113_y0(h_u_cla32_and6112_y0, h_u_cla32_and6111_y0, h_u_cla32_and6113_y0);
  and_gate and_gate_h_u_cla32_and6114_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6114_y0);
  and_gate and_gate_h_u_cla32_and6115_y0(h_u_cla32_and6114_y0, h_u_cla32_and6113_y0, h_u_cla32_and6115_y0);
  and_gate and_gate_h_u_cla32_and6116_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6116_y0);
  and_gate and_gate_h_u_cla32_and6117_y0(h_u_cla32_and6116_y0, h_u_cla32_and6115_y0, h_u_cla32_and6117_y0);
  and_gate and_gate_h_u_cla32_and6118_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6118_y0);
  and_gate and_gate_h_u_cla32_and6119_y0(h_u_cla32_and6118_y0, h_u_cla32_and6117_y0, h_u_cla32_and6119_y0);
  and_gate and_gate_h_u_cla32_and6120_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6120_y0);
  and_gate and_gate_h_u_cla32_and6121_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6121_y0);
  and_gate and_gate_h_u_cla32_and6122_y0(h_u_cla32_and6121_y0, h_u_cla32_and6120_y0, h_u_cla32_and6122_y0);
  and_gate and_gate_h_u_cla32_and6123_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6123_y0);
  and_gate and_gate_h_u_cla32_and6124_y0(h_u_cla32_and6123_y0, h_u_cla32_and6122_y0, h_u_cla32_and6124_y0);
  and_gate and_gate_h_u_cla32_and6125_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6125_y0);
  and_gate and_gate_h_u_cla32_and6126_y0(h_u_cla32_and6125_y0, h_u_cla32_and6124_y0, h_u_cla32_and6126_y0);
  and_gate and_gate_h_u_cla32_and6127_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6127_y0);
  and_gate and_gate_h_u_cla32_and6128_y0(h_u_cla32_and6127_y0, h_u_cla32_and6126_y0, h_u_cla32_and6128_y0);
  and_gate and_gate_h_u_cla32_and6129_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6129_y0);
  and_gate and_gate_h_u_cla32_and6130_y0(h_u_cla32_and6129_y0, h_u_cla32_and6128_y0, h_u_cla32_and6130_y0);
  and_gate and_gate_h_u_cla32_and6131_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6131_y0);
  and_gate and_gate_h_u_cla32_and6132_y0(h_u_cla32_and6131_y0, h_u_cla32_and6130_y0, h_u_cla32_and6132_y0);
  and_gate and_gate_h_u_cla32_and6133_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6133_y0);
  and_gate and_gate_h_u_cla32_and6134_y0(h_u_cla32_and6133_y0, h_u_cla32_and6132_y0, h_u_cla32_and6134_y0);
  and_gate and_gate_h_u_cla32_and6135_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6135_y0);
  and_gate and_gate_h_u_cla32_and6136_y0(h_u_cla32_and6135_y0, h_u_cla32_and6134_y0, h_u_cla32_and6136_y0);
  and_gate and_gate_h_u_cla32_and6137_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6137_y0);
  and_gate and_gate_h_u_cla32_and6138_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6138_y0);
  and_gate and_gate_h_u_cla32_and6139_y0(h_u_cla32_and6138_y0, h_u_cla32_and6137_y0, h_u_cla32_and6139_y0);
  and_gate and_gate_h_u_cla32_and6140_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6140_y0);
  and_gate and_gate_h_u_cla32_and6141_y0(h_u_cla32_and6140_y0, h_u_cla32_and6139_y0, h_u_cla32_and6141_y0);
  and_gate and_gate_h_u_cla32_and6142_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6142_y0);
  and_gate and_gate_h_u_cla32_and6143_y0(h_u_cla32_and6142_y0, h_u_cla32_and6141_y0, h_u_cla32_and6143_y0);
  and_gate and_gate_h_u_cla32_and6144_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6144_y0);
  and_gate and_gate_h_u_cla32_and6145_y0(h_u_cla32_and6144_y0, h_u_cla32_and6143_y0, h_u_cla32_and6145_y0);
  and_gate and_gate_h_u_cla32_and6146_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6146_y0);
  and_gate and_gate_h_u_cla32_and6147_y0(h_u_cla32_and6146_y0, h_u_cla32_and6145_y0, h_u_cla32_and6147_y0);
  and_gate and_gate_h_u_cla32_and6148_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6148_y0);
  and_gate and_gate_h_u_cla32_and6149_y0(h_u_cla32_and6148_y0, h_u_cla32_and6147_y0, h_u_cla32_and6149_y0);
  and_gate and_gate_h_u_cla32_and6150_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6150_y0);
  and_gate and_gate_h_u_cla32_and6151_y0(h_u_cla32_and6150_y0, h_u_cla32_and6149_y0, h_u_cla32_and6151_y0);
  and_gate and_gate_h_u_cla32_and6152_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6152_y0);
  and_gate and_gate_h_u_cla32_and6153_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6153_y0);
  and_gate and_gate_h_u_cla32_and6154_y0(h_u_cla32_and6153_y0, h_u_cla32_and6152_y0, h_u_cla32_and6154_y0);
  and_gate and_gate_h_u_cla32_and6155_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6155_y0);
  and_gate and_gate_h_u_cla32_and6156_y0(h_u_cla32_and6155_y0, h_u_cla32_and6154_y0, h_u_cla32_and6156_y0);
  and_gate and_gate_h_u_cla32_and6157_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6157_y0);
  and_gate and_gate_h_u_cla32_and6158_y0(h_u_cla32_and6157_y0, h_u_cla32_and6156_y0, h_u_cla32_and6158_y0);
  and_gate and_gate_h_u_cla32_and6159_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6159_y0);
  and_gate and_gate_h_u_cla32_and6160_y0(h_u_cla32_and6159_y0, h_u_cla32_and6158_y0, h_u_cla32_and6160_y0);
  and_gate and_gate_h_u_cla32_and6161_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6161_y0);
  and_gate and_gate_h_u_cla32_and6162_y0(h_u_cla32_and6161_y0, h_u_cla32_and6160_y0, h_u_cla32_and6162_y0);
  and_gate and_gate_h_u_cla32_and6163_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6163_y0);
  and_gate and_gate_h_u_cla32_and6164_y0(h_u_cla32_and6163_y0, h_u_cla32_and6162_y0, h_u_cla32_and6164_y0);
  and_gate and_gate_h_u_cla32_and6165_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6165_y0);
  and_gate and_gate_h_u_cla32_and6166_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6166_y0);
  and_gate and_gate_h_u_cla32_and6167_y0(h_u_cla32_and6166_y0, h_u_cla32_and6165_y0, h_u_cla32_and6167_y0);
  and_gate and_gate_h_u_cla32_and6168_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6168_y0);
  and_gate and_gate_h_u_cla32_and6169_y0(h_u_cla32_and6168_y0, h_u_cla32_and6167_y0, h_u_cla32_and6169_y0);
  and_gate and_gate_h_u_cla32_and6170_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6170_y0);
  and_gate and_gate_h_u_cla32_and6171_y0(h_u_cla32_and6170_y0, h_u_cla32_and6169_y0, h_u_cla32_and6171_y0);
  and_gate and_gate_h_u_cla32_and6172_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6172_y0);
  and_gate and_gate_h_u_cla32_and6173_y0(h_u_cla32_and6172_y0, h_u_cla32_and6171_y0, h_u_cla32_and6173_y0);
  and_gate and_gate_h_u_cla32_and6174_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6174_y0);
  and_gate and_gate_h_u_cla32_and6175_y0(h_u_cla32_and6174_y0, h_u_cla32_and6173_y0, h_u_cla32_and6175_y0);
  and_gate and_gate_h_u_cla32_and6176_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6176_y0);
  and_gate and_gate_h_u_cla32_and6177_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6177_y0);
  and_gate and_gate_h_u_cla32_and6178_y0(h_u_cla32_and6177_y0, h_u_cla32_and6176_y0, h_u_cla32_and6178_y0);
  and_gate and_gate_h_u_cla32_and6179_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6179_y0);
  and_gate and_gate_h_u_cla32_and6180_y0(h_u_cla32_and6179_y0, h_u_cla32_and6178_y0, h_u_cla32_and6180_y0);
  and_gate and_gate_h_u_cla32_and6181_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6181_y0);
  and_gate and_gate_h_u_cla32_and6182_y0(h_u_cla32_and6181_y0, h_u_cla32_and6180_y0, h_u_cla32_and6182_y0);
  and_gate and_gate_h_u_cla32_and6183_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6183_y0);
  and_gate and_gate_h_u_cla32_and6184_y0(h_u_cla32_and6183_y0, h_u_cla32_and6182_y0, h_u_cla32_and6184_y0);
  and_gate and_gate_h_u_cla32_and6185_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6185_y0);
  and_gate and_gate_h_u_cla32_and6186_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6186_y0);
  and_gate and_gate_h_u_cla32_and6187_y0(h_u_cla32_and6186_y0, h_u_cla32_and6185_y0, h_u_cla32_and6187_y0);
  and_gate and_gate_h_u_cla32_and6188_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6188_y0);
  and_gate and_gate_h_u_cla32_and6189_y0(h_u_cla32_and6188_y0, h_u_cla32_and6187_y0, h_u_cla32_and6189_y0);
  and_gate and_gate_h_u_cla32_and6190_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6190_y0);
  and_gate and_gate_h_u_cla32_and6191_y0(h_u_cla32_and6190_y0, h_u_cla32_and6189_y0, h_u_cla32_and6191_y0);
  and_gate and_gate_h_u_cla32_and6192_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6192_y0);
  and_gate and_gate_h_u_cla32_and6193_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6193_y0);
  and_gate and_gate_h_u_cla32_and6194_y0(h_u_cla32_and6193_y0, h_u_cla32_and6192_y0, h_u_cla32_and6194_y0);
  and_gate and_gate_h_u_cla32_and6195_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6195_y0);
  and_gate and_gate_h_u_cla32_and6196_y0(h_u_cla32_and6195_y0, h_u_cla32_and6194_y0, h_u_cla32_and6196_y0);
  and_gate and_gate_h_u_cla32_and6197_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and6197_y0);
  and_gate and_gate_h_u_cla32_and6198_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and6198_y0);
  and_gate and_gate_h_u_cla32_and6199_y0(h_u_cla32_and6198_y0, h_u_cla32_and6197_y0, h_u_cla32_and6199_y0);
  and_gate and_gate_h_u_cla32_and6200_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and6200_y0);
  or_gate or_gate_h_u_cla32_or325_y0(h_u_cla32_and6200_y0, h_u_cla32_and5575_y0, h_u_cla32_or325_y0);
  or_gate or_gate_h_u_cla32_or326_y0(h_u_cla32_or325_y0, h_u_cla32_and5624_y0, h_u_cla32_or326_y0);
  or_gate or_gate_h_u_cla32_or327_y0(h_u_cla32_or326_y0, h_u_cla32_and5671_y0, h_u_cla32_or327_y0);
  or_gate or_gate_h_u_cla32_or328_y0(h_u_cla32_or327_y0, h_u_cla32_and5716_y0, h_u_cla32_or328_y0);
  or_gate or_gate_h_u_cla32_or329_y0(h_u_cla32_or328_y0, h_u_cla32_and5759_y0, h_u_cla32_or329_y0);
  or_gate or_gate_h_u_cla32_or330_y0(h_u_cla32_or329_y0, h_u_cla32_and5800_y0, h_u_cla32_or330_y0);
  or_gate or_gate_h_u_cla32_or331_y0(h_u_cla32_or330_y0, h_u_cla32_and5839_y0, h_u_cla32_or331_y0);
  or_gate or_gate_h_u_cla32_or332_y0(h_u_cla32_or331_y0, h_u_cla32_and5876_y0, h_u_cla32_or332_y0);
  or_gate or_gate_h_u_cla32_or333_y0(h_u_cla32_or332_y0, h_u_cla32_and5911_y0, h_u_cla32_or333_y0);
  or_gate or_gate_h_u_cla32_or334_y0(h_u_cla32_or333_y0, h_u_cla32_and5944_y0, h_u_cla32_or334_y0);
  or_gate or_gate_h_u_cla32_or335_y0(h_u_cla32_or334_y0, h_u_cla32_and5975_y0, h_u_cla32_or335_y0);
  or_gate or_gate_h_u_cla32_or336_y0(h_u_cla32_or335_y0, h_u_cla32_and6004_y0, h_u_cla32_or336_y0);
  or_gate or_gate_h_u_cla32_or337_y0(h_u_cla32_or336_y0, h_u_cla32_and6031_y0, h_u_cla32_or337_y0);
  or_gate or_gate_h_u_cla32_or338_y0(h_u_cla32_or337_y0, h_u_cla32_and6056_y0, h_u_cla32_or338_y0);
  or_gate or_gate_h_u_cla32_or339_y0(h_u_cla32_or338_y0, h_u_cla32_and6079_y0, h_u_cla32_or339_y0);
  or_gate or_gate_h_u_cla32_or340_y0(h_u_cla32_or339_y0, h_u_cla32_and6100_y0, h_u_cla32_or340_y0);
  or_gate or_gate_h_u_cla32_or341_y0(h_u_cla32_or340_y0, h_u_cla32_and6119_y0, h_u_cla32_or341_y0);
  or_gate or_gate_h_u_cla32_or342_y0(h_u_cla32_or341_y0, h_u_cla32_and6136_y0, h_u_cla32_or342_y0);
  or_gate or_gate_h_u_cla32_or343_y0(h_u_cla32_or342_y0, h_u_cla32_and6151_y0, h_u_cla32_or343_y0);
  or_gate or_gate_h_u_cla32_or344_y0(h_u_cla32_or343_y0, h_u_cla32_and6164_y0, h_u_cla32_or344_y0);
  or_gate or_gate_h_u_cla32_or345_y0(h_u_cla32_or344_y0, h_u_cla32_and6175_y0, h_u_cla32_or345_y0);
  or_gate or_gate_h_u_cla32_or346_y0(h_u_cla32_or345_y0, h_u_cla32_and6184_y0, h_u_cla32_or346_y0);
  or_gate or_gate_h_u_cla32_or347_y0(h_u_cla32_or346_y0, h_u_cla32_and6191_y0, h_u_cla32_or347_y0);
  or_gate or_gate_h_u_cla32_or348_y0(h_u_cla32_or347_y0, h_u_cla32_and6196_y0, h_u_cla32_or348_y0);
  or_gate or_gate_h_u_cla32_or349_y0(h_u_cla32_or348_y0, h_u_cla32_and6199_y0, h_u_cla32_or349_y0);
  or_gate or_gate_h_u_cla32_or350_y0(h_u_cla32_pg_logic25_y1, h_u_cla32_or349_y0, h_u_cla32_or350_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic26_y0(a_26, b_26, h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_pg_logic26_y2);
  xor_gate xor_gate_h_u_cla32_xor26_y0(h_u_cla32_pg_logic26_y2, h_u_cla32_or350_y0, h_u_cla32_xor26_y0);
  and_gate and_gate_h_u_cla32_and6201_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and6201_y0);
  and_gate and_gate_h_u_cla32_and6202_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and6202_y0);
  and_gate and_gate_h_u_cla32_and6203_y0(h_u_cla32_and6202_y0, h_u_cla32_and6201_y0, h_u_cla32_and6203_y0);
  and_gate and_gate_h_u_cla32_and6204_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and6204_y0);
  and_gate and_gate_h_u_cla32_and6205_y0(h_u_cla32_and6204_y0, h_u_cla32_and6203_y0, h_u_cla32_and6205_y0);
  and_gate and_gate_h_u_cla32_and6206_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and6206_y0);
  and_gate and_gate_h_u_cla32_and6207_y0(h_u_cla32_and6206_y0, h_u_cla32_and6205_y0, h_u_cla32_and6207_y0);
  and_gate and_gate_h_u_cla32_and6208_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and6208_y0);
  and_gate and_gate_h_u_cla32_and6209_y0(h_u_cla32_and6208_y0, h_u_cla32_and6207_y0, h_u_cla32_and6209_y0);
  and_gate and_gate_h_u_cla32_and6210_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and6210_y0);
  and_gate and_gate_h_u_cla32_and6211_y0(h_u_cla32_and6210_y0, h_u_cla32_and6209_y0, h_u_cla32_and6211_y0);
  and_gate and_gate_h_u_cla32_and6212_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and6212_y0);
  and_gate and_gate_h_u_cla32_and6213_y0(h_u_cla32_and6212_y0, h_u_cla32_and6211_y0, h_u_cla32_and6213_y0);
  and_gate and_gate_h_u_cla32_and6214_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and6214_y0);
  and_gate and_gate_h_u_cla32_and6215_y0(h_u_cla32_and6214_y0, h_u_cla32_and6213_y0, h_u_cla32_and6215_y0);
  and_gate and_gate_h_u_cla32_and6216_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and6216_y0);
  and_gate and_gate_h_u_cla32_and6217_y0(h_u_cla32_and6216_y0, h_u_cla32_and6215_y0, h_u_cla32_and6217_y0);
  and_gate and_gate_h_u_cla32_and6218_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and6218_y0);
  and_gate and_gate_h_u_cla32_and6219_y0(h_u_cla32_and6218_y0, h_u_cla32_and6217_y0, h_u_cla32_and6219_y0);
  and_gate and_gate_h_u_cla32_and6220_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and6220_y0);
  and_gate and_gate_h_u_cla32_and6221_y0(h_u_cla32_and6220_y0, h_u_cla32_and6219_y0, h_u_cla32_and6221_y0);
  and_gate and_gate_h_u_cla32_and6222_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and6222_y0);
  and_gate and_gate_h_u_cla32_and6223_y0(h_u_cla32_and6222_y0, h_u_cla32_and6221_y0, h_u_cla32_and6223_y0);
  and_gate and_gate_h_u_cla32_and6224_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and6224_y0);
  and_gate and_gate_h_u_cla32_and6225_y0(h_u_cla32_and6224_y0, h_u_cla32_and6223_y0, h_u_cla32_and6225_y0);
  and_gate and_gate_h_u_cla32_and6226_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and6226_y0);
  and_gate and_gate_h_u_cla32_and6227_y0(h_u_cla32_and6226_y0, h_u_cla32_and6225_y0, h_u_cla32_and6227_y0);
  and_gate and_gate_h_u_cla32_and6228_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and6228_y0);
  and_gate and_gate_h_u_cla32_and6229_y0(h_u_cla32_and6228_y0, h_u_cla32_and6227_y0, h_u_cla32_and6229_y0);
  and_gate and_gate_h_u_cla32_and6230_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and6230_y0);
  and_gate and_gate_h_u_cla32_and6231_y0(h_u_cla32_and6230_y0, h_u_cla32_and6229_y0, h_u_cla32_and6231_y0);
  and_gate and_gate_h_u_cla32_and6232_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and6232_y0);
  and_gate and_gate_h_u_cla32_and6233_y0(h_u_cla32_and6232_y0, h_u_cla32_and6231_y0, h_u_cla32_and6233_y0);
  and_gate and_gate_h_u_cla32_and6234_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and6234_y0);
  and_gate and_gate_h_u_cla32_and6235_y0(h_u_cla32_and6234_y0, h_u_cla32_and6233_y0, h_u_cla32_and6235_y0);
  and_gate and_gate_h_u_cla32_and6236_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and6236_y0);
  and_gate and_gate_h_u_cla32_and6237_y0(h_u_cla32_and6236_y0, h_u_cla32_and6235_y0, h_u_cla32_and6237_y0);
  and_gate and_gate_h_u_cla32_and6238_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and6238_y0);
  and_gate and_gate_h_u_cla32_and6239_y0(h_u_cla32_and6238_y0, h_u_cla32_and6237_y0, h_u_cla32_and6239_y0);
  and_gate and_gate_h_u_cla32_and6240_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and6240_y0);
  and_gate and_gate_h_u_cla32_and6241_y0(h_u_cla32_and6240_y0, h_u_cla32_and6239_y0, h_u_cla32_and6241_y0);
  and_gate and_gate_h_u_cla32_and6242_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and6242_y0);
  and_gate and_gate_h_u_cla32_and6243_y0(h_u_cla32_and6242_y0, h_u_cla32_and6241_y0, h_u_cla32_and6243_y0);
  and_gate and_gate_h_u_cla32_and6244_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and6244_y0);
  and_gate and_gate_h_u_cla32_and6245_y0(h_u_cla32_and6244_y0, h_u_cla32_and6243_y0, h_u_cla32_and6245_y0);
  and_gate and_gate_h_u_cla32_and6246_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and6246_y0);
  and_gate and_gate_h_u_cla32_and6247_y0(h_u_cla32_and6246_y0, h_u_cla32_and6245_y0, h_u_cla32_and6247_y0);
  and_gate and_gate_h_u_cla32_and6248_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and6248_y0);
  and_gate and_gate_h_u_cla32_and6249_y0(h_u_cla32_and6248_y0, h_u_cla32_and6247_y0, h_u_cla32_and6249_y0);
  and_gate and_gate_h_u_cla32_and6250_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and6250_y0);
  and_gate and_gate_h_u_cla32_and6251_y0(h_u_cla32_and6250_y0, h_u_cla32_and6249_y0, h_u_cla32_and6251_y0);
  and_gate and_gate_h_u_cla32_and6252_y0(h_u_cla32_pg_logic26_y0, constant_wire_0, h_u_cla32_and6252_y0);
  and_gate and_gate_h_u_cla32_and6253_y0(h_u_cla32_and6252_y0, h_u_cla32_and6251_y0, h_u_cla32_and6253_y0);
  and_gate and_gate_h_u_cla32_and6254_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6254_y0);
  and_gate and_gate_h_u_cla32_and6255_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6255_y0);
  and_gate and_gate_h_u_cla32_and6256_y0(h_u_cla32_and6255_y0, h_u_cla32_and6254_y0, h_u_cla32_and6256_y0);
  and_gate and_gate_h_u_cla32_and6257_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6257_y0);
  and_gate and_gate_h_u_cla32_and6258_y0(h_u_cla32_and6257_y0, h_u_cla32_and6256_y0, h_u_cla32_and6258_y0);
  and_gate and_gate_h_u_cla32_and6259_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6259_y0);
  and_gate and_gate_h_u_cla32_and6260_y0(h_u_cla32_and6259_y0, h_u_cla32_and6258_y0, h_u_cla32_and6260_y0);
  and_gate and_gate_h_u_cla32_and6261_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6261_y0);
  and_gate and_gate_h_u_cla32_and6262_y0(h_u_cla32_and6261_y0, h_u_cla32_and6260_y0, h_u_cla32_and6262_y0);
  and_gate and_gate_h_u_cla32_and6263_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6263_y0);
  and_gate and_gate_h_u_cla32_and6264_y0(h_u_cla32_and6263_y0, h_u_cla32_and6262_y0, h_u_cla32_and6264_y0);
  and_gate and_gate_h_u_cla32_and6265_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6265_y0);
  and_gate and_gate_h_u_cla32_and6266_y0(h_u_cla32_and6265_y0, h_u_cla32_and6264_y0, h_u_cla32_and6266_y0);
  and_gate and_gate_h_u_cla32_and6267_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6267_y0);
  and_gate and_gate_h_u_cla32_and6268_y0(h_u_cla32_and6267_y0, h_u_cla32_and6266_y0, h_u_cla32_and6268_y0);
  and_gate and_gate_h_u_cla32_and6269_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6269_y0);
  and_gate and_gate_h_u_cla32_and6270_y0(h_u_cla32_and6269_y0, h_u_cla32_and6268_y0, h_u_cla32_and6270_y0);
  and_gate and_gate_h_u_cla32_and6271_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6271_y0);
  and_gate and_gate_h_u_cla32_and6272_y0(h_u_cla32_and6271_y0, h_u_cla32_and6270_y0, h_u_cla32_and6272_y0);
  and_gate and_gate_h_u_cla32_and6273_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6273_y0);
  and_gate and_gate_h_u_cla32_and6274_y0(h_u_cla32_and6273_y0, h_u_cla32_and6272_y0, h_u_cla32_and6274_y0);
  and_gate and_gate_h_u_cla32_and6275_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6275_y0);
  and_gate and_gate_h_u_cla32_and6276_y0(h_u_cla32_and6275_y0, h_u_cla32_and6274_y0, h_u_cla32_and6276_y0);
  and_gate and_gate_h_u_cla32_and6277_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6277_y0);
  and_gate and_gate_h_u_cla32_and6278_y0(h_u_cla32_and6277_y0, h_u_cla32_and6276_y0, h_u_cla32_and6278_y0);
  and_gate and_gate_h_u_cla32_and6279_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6279_y0);
  and_gate and_gate_h_u_cla32_and6280_y0(h_u_cla32_and6279_y0, h_u_cla32_and6278_y0, h_u_cla32_and6280_y0);
  and_gate and_gate_h_u_cla32_and6281_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6281_y0);
  and_gate and_gate_h_u_cla32_and6282_y0(h_u_cla32_and6281_y0, h_u_cla32_and6280_y0, h_u_cla32_and6282_y0);
  and_gate and_gate_h_u_cla32_and6283_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6283_y0);
  and_gate and_gate_h_u_cla32_and6284_y0(h_u_cla32_and6283_y0, h_u_cla32_and6282_y0, h_u_cla32_and6284_y0);
  and_gate and_gate_h_u_cla32_and6285_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6285_y0);
  and_gate and_gate_h_u_cla32_and6286_y0(h_u_cla32_and6285_y0, h_u_cla32_and6284_y0, h_u_cla32_and6286_y0);
  and_gate and_gate_h_u_cla32_and6287_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6287_y0);
  and_gate and_gate_h_u_cla32_and6288_y0(h_u_cla32_and6287_y0, h_u_cla32_and6286_y0, h_u_cla32_and6288_y0);
  and_gate and_gate_h_u_cla32_and6289_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6289_y0);
  and_gate and_gate_h_u_cla32_and6290_y0(h_u_cla32_and6289_y0, h_u_cla32_and6288_y0, h_u_cla32_and6290_y0);
  and_gate and_gate_h_u_cla32_and6291_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6291_y0);
  and_gate and_gate_h_u_cla32_and6292_y0(h_u_cla32_and6291_y0, h_u_cla32_and6290_y0, h_u_cla32_and6292_y0);
  and_gate and_gate_h_u_cla32_and6293_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6293_y0);
  and_gate and_gate_h_u_cla32_and6294_y0(h_u_cla32_and6293_y0, h_u_cla32_and6292_y0, h_u_cla32_and6294_y0);
  and_gate and_gate_h_u_cla32_and6295_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6295_y0);
  and_gate and_gate_h_u_cla32_and6296_y0(h_u_cla32_and6295_y0, h_u_cla32_and6294_y0, h_u_cla32_and6296_y0);
  and_gate and_gate_h_u_cla32_and6297_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6297_y0);
  and_gate and_gate_h_u_cla32_and6298_y0(h_u_cla32_and6297_y0, h_u_cla32_and6296_y0, h_u_cla32_and6298_y0);
  and_gate and_gate_h_u_cla32_and6299_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6299_y0);
  and_gate and_gate_h_u_cla32_and6300_y0(h_u_cla32_and6299_y0, h_u_cla32_and6298_y0, h_u_cla32_and6300_y0);
  and_gate and_gate_h_u_cla32_and6301_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6301_y0);
  and_gate and_gate_h_u_cla32_and6302_y0(h_u_cla32_and6301_y0, h_u_cla32_and6300_y0, h_u_cla32_and6302_y0);
  and_gate and_gate_h_u_cla32_and6303_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6303_y0);
  and_gate and_gate_h_u_cla32_and6304_y0(h_u_cla32_and6303_y0, h_u_cla32_and6302_y0, h_u_cla32_and6304_y0);
  and_gate and_gate_h_u_cla32_and6305_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6305_y0);
  and_gate and_gate_h_u_cla32_and6306_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6306_y0);
  and_gate and_gate_h_u_cla32_and6307_y0(h_u_cla32_and6306_y0, h_u_cla32_and6305_y0, h_u_cla32_and6307_y0);
  and_gate and_gate_h_u_cla32_and6308_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6308_y0);
  and_gate and_gate_h_u_cla32_and6309_y0(h_u_cla32_and6308_y0, h_u_cla32_and6307_y0, h_u_cla32_and6309_y0);
  and_gate and_gate_h_u_cla32_and6310_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6310_y0);
  and_gate and_gate_h_u_cla32_and6311_y0(h_u_cla32_and6310_y0, h_u_cla32_and6309_y0, h_u_cla32_and6311_y0);
  and_gate and_gate_h_u_cla32_and6312_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6312_y0);
  and_gate and_gate_h_u_cla32_and6313_y0(h_u_cla32_and6312_y0, h_u_cla32_and6311_y0, h_u_cla32_and6313_y0);
  and_gate and_gate_h_u_cla32_and6314_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6314_y0);
  and_gate and_gate_h_u_cla32_and6315_y0(h_u_cla32_and6314_y0, h_u_cla32_and6313_y0, h_u_cla32_and6315_y0);
  and_gate and_gate_h_u_cla32_and6316_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6316_y0);
  and_gate and_gate_h_u_cla32_and6317_y0(h_u_cla32_and6316_y0, h_u_cla32_and6315_y0, h_u_cla32_and6317_y0);
  and_gate and_gate_h_u_cla32_and6318_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6318_y0);
  and_gate and_gate_h_u_cla32_and6319_y0(h_u_cla32_and6318_y0, h_u_cla32_and6317_y0, h_u_cla32_and6319_y0);
  and_gate and_gate_h_u_cla32_and6320_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6320_y0);
  and_gate and_gate_h_u_cla32_and6321_y0(h_u_cla32_and6320_y0, h_u_cla32_and6319_y0, h_u_cla32_and6321_y0);
  and_gate and_gate_h_u_cla32_and6322_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6322_y0);
  and_gate and_gate_h_u_cla32_and6323_y0(h_u_cla32_and6322_y0, h_u_cla32_and6321_y0, h_u_cla32_and6323_y0);
  and_gate and_gate_h_u_cla32_and6324_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6324_y0);
  and_gate and_gate_h_u_cla32_and6325_y0(h_u_cla32_and6324_y0, h_u_cla32_and6323_y0, h_u_cla32_and6325_y0);
  and_gate and_gate_h_u_cla32_and6326_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6326_y0);
  and_gate and_gate_h_u_cla32_and6327_y0(h_u_cla32_and6326_y0, h_u_cla32_and6325_y0, h_u_cla32_and6327_y0);
  and_gate and_gate_h_u_cla32_and6328_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6328_y0);
  and_gate and_gate_h_u_cla32_and6329_y0(h_u_cla32_and6328_y0, h_u_cla32_and6327_y0, h_u_cla32_and6329_y0);
  and_gate and_gate_h_u_cla32_and6330_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6330_y0);
  and_gate and_gate_h_u_cla32_and6331_y0(h_u_cla32_and6330_y0, h_u_cla32_and6329_y0, h_u_cla32_and6331_y0);
  and_gate and_gate_h_u_cla32_and6332_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6332_y0);
  and_gate and_gate_h_u_cla32_and6333_y0(h_u_cla32_and6332_y0, h_u_cla32_and6331_y0, h_u_cla32_and6333_y0);
  and_gate and_gate_h_u_cla32_and6334_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6334_y0);
  and_gate and_gate_h_u_cla32_and6335_y0(h_u_cla32_and6334_y0, h_u_cla32_and6333_y0, h_u_cla32_and6335_y0);
  and_gate and_gate_h_u_cla32_and6336_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6336_y0);
  and_gate and_gate_h_u_cla32_and6337_y0(h_u_cla32_and6336_y0, h_u_cla32_and6335_y0, h_u_cla32_and6337_y0);
  and_gate and_gate_h_u_cla32_and6338_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6338_y0);
  and_gate and_gate_h_u_cla32_and6339_y0(h_u_cla32_and6338_y0, h_u_cla32_and6337_y0, h_u_cla32_and6339_y0);
  and_gate and_gate_h_u_cla32_and6340_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6340_y0);
  and_gate and_gate_h_u_cla32_and6341_y0(h_u_cla32_and6340_y0, h_u_cla32_and6339_y0, h_u_cla32_and6341_y0);
  and_gate and_gate_h_u_cla32_and6342_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6342_y0);
  and_gate and_gate_h_u_cla32_and6343_y0(h_u_cla32_and6342_y0, h_u_cla32_and6341_y0, h_u_cla32_and6343_y0);
  and_gate and_gate_h_u_cla32_and6344_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6344_y0);
  and_gate and_gate_h_u_cla32_and6345_y0(h_u_cla32_and6344_y0, h_u_cla32_and6343_y0, h_u_cla32_and6345_y0);
  and_gate and_gate_h_u_cla32_and6346_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6346_y0);
  and_gate and_gate_h_u_cla32_and6347_y0(h_u_cla32_and6346_y0, h_u_cla32_and6345_y0, h_u_cla32_and6347_y0);
  and_gate and_gate_h_u_cla32_and6348_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6348_y0);
  and_gate and_gate_h_u_cla32_and6349_y0(h_u_cla32_and6348_y0, h_u_cla32_and6347_y0, h_u_cla32_and6349_y0);
  and_gate and_gate_h_u_cla32_and6350_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6350_y0);
  and_gate and_gate_h_u_cla32_and6351_y0(h_u_cla32_and6350_y0, h_u_cla32_and6349_y0, h_u_cla32_and6351_y0);
  and_gate and_gate_h_u_cla32_and6352_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and6352_y0);
  and_gate and_gate_h_u_cla32_and6353_y0(h_u_cla32_and6352_y0, h_u_cla32_and6351_y0, h_u_cla32_and6353_y0);
  and_gate and_gate_h_u_cla32_and6354_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6354_y0);
  and_gate and_gate_h_u_cla32_and6355_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6355_y0);
  and_gate and_gate_h_u_cla32_and6356_y0(h_u_cla32_and6355_y0, h_u_cla32_and6354_y0, h_u_cla32_and6356_y0);
  and_gate and_gate_h_u_cla32_and6357_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6357_y0);
  and_gate and_gate_h_u_cla32_and6358_y0(h_u_cla32_and6357_y0, h_u_cla32_and6356_y0, h_u_cla32_and6358_y0);
  and_gate and_gate_h_u_cla32_and6359_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6359_y0);
  and_gate and_gate_h_u_cla32_and6360_y0(h_u_cla32_and6359_y0, h_u_cla32_and6358_y0, h_u_cla32_and6360_y0);
  and_gate and_gate_h_u_cla32_and6361_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6361_y0);
  and_gate and_gate_h_u_cla32_and6362_y0(h_u_cla32_and6361_y0, h_u_cla32_and6360_y0, h_u_cla32_and6362_y0);
  and_gate and_gate_h_u_cla32_and6363_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6363_y0);
  and_gate and_gate_h_u_cla32_and6364_y0(h_u_cla32_and6363_y0, h_u_cla32_and6362_y0, h_u_cla32_and6364_y0);
  and_gate and_gate_h_u_cla32_and6365_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6365_y0);
  and_gate and_gate_h_u_cla32_and6366_y0(h_u_cla32_and6365_y0, h_u_cla32_and6364_y0, h_u_cla32_and6366_y0);
  and_gate and_gate_h_u_cla32_and6367_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6367_y0);
  and_gate and_gate_h_u_cla32_and6368_y0(h_u_cla32_and6367_y0, h_u_cla32_and6366_y0, h_u_cla32_and6368_y0);
  and_gate and_gate_h_u_cla32_and6369_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6369_y0);
  and_gate and_gate_h_u_cla32_and6370_y0(h_u_cla32_and6369_y0, h_u_cla32_and6368_y0, h_u_cla32_and6370_y0);
  and_gate and_gate_h_u_cla32_and6371_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6371_y0);
  and_gate and_gate_h_u_cla32_and6372_y0(h_u_cla32_and6371_y0, h_u_cla32_and6370_y0, h_u_cla32_and6372_y0);
  and_gate and_gate_h_u_cla32_and6373_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6373_y0);
  and_gate and_gate_h_u_cla32_and6374_y0(h_u_cla32_and6373_y0, h_u_cla32_and6372_y0, h_u_cla32_and6374_y0);
  and_gate and_gate_h_u_cla32_and6375_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6375_y0);
  and_gate and_gate_h_u_cla32_and6376_y0(h_u_cla32_and6375_y0, h_u_cla32_and6374_y0, h_u_cla32_and6376_y0);
  and_gate and_gate_h_u_cla32_and6377_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6377_y0);
  and_gate and_gate_h_u_cla32_and6378_y0(h_u_cla32_and6377_y0, h_u_cla32_and6376_y0, h_u_cla32_and6378_y0);
  and_gate and_gate_h_u_cla32_and6379_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6379_y0);
  and_gate and_gate_h_u_cla32_and6380_y0(h_u_cla32_and6379_y0, h_u_cla32_and6378_y0, h_u_cla32_and6380_y0);
  and_gate and_gate_h_u_cla32_and6381_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6381_y0);
  and_gate and_gate_h_u_cla32_and6382_y0(h_u_cla32_and6381_y0, h_u_cla32_and6380_y0, h_u_cla32_and6382_y0);
  and_gate and_gate_h_u_cla32_and6383_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6383_y0);
  and_gate and_gate_h_u_cla32_and6384_y0(h_u_cla32_and6383_y0, h_u_cla32_and6382_y0, h_u_cla32_and6384_y0);
  and_gate and_gate_h_u_cla32_and6385_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6385_y0);
  and_gate and_gate_h_u_cla32_and6386_y0(h_u_cla32_and6385_y0, h_u_cla32_and6384_y0, h_u_cla32_and6386_y0);
  and_gate and_gate_h_u_cla32_and6387_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6387_y0);
  and_gate and_gate_h_u_cla32_and6388_y0(h_u_cla32_and6387_y0, h_u_cla32_and6386_y0, h_u_cla32_and6388_y0);
  and_gate and_gate_h_u_cla32_and6389_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6389_y0);
  and_gate and_gate_h_u_cla32_and6390_y0(h_u_cla32_and6389_y0, h_u_cla32_and6388_y0, h_u_cla32_and6390_y0);
  and_gate and_gate_h_u_cla32_and6391_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6391_y0);
  and_gate and_gate_h_u_cla32_and6392_y0(h_u_cla32_and6391_y0, h_u_cla32_and6390_y0, h_u_cla32_and6392_y0);
  and_gate and_gate_h_u_cla32_and6393_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6393_y0);
  and_gate and_gate_h_u_cla32_and6394_y0(h_u_cla32_and6393_y0, h_u_cla32_and6392_y0, h_u_cla32_and6394_y0);
  and_gate and_gate_h_u_cla32_and6395_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6395_y0);
  and_gate and_gate_h_u_cla32_and6396_y0(h_u_cla32_and6395_y0, h_u_cla32_and6394_y0, h_u_cla32_and6396_y0);
  and_gate and_gate_h_u_cla32_and6397_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6397_y0);
  and_gate and_gate_h_u_cla32_and6398_y0(h_u_cla32_and6397_y0, h_u_cla32_and6396_y0, h_u_cla32_and6398_y0);
  and_gate and_gate_h_u_cla32_and6399_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and6399_y0);
  and_gate and_gate_h_u_cla32_and6400_y0(h_u_cla32_and6399_y0, h_u_cla32_and6398_y0, h_u_cla32_and6400_y0);
  and_gate and_gate_h_u_cla32_and6401_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6401_y0);
  and_gate and_gate_h_u_cla32_and6402_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6402_y0);
  and_gate and_gate_h_u_cla32_and6403_y0(h_u_cla32_and6402_y0, h_u_cla32_and6401_y0, h_u_cla32_and6403_y0);
  and_gate and_gate_h_u_cla32_and6404_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6404_y0);
  and_gate and_gate_h_u_cla32_and6405_y0(h_u_cla32_and6404_y0, h_u_cla32_and6403_y0, h_u_cla32_and6405_y0);
  and_gate and_gate_h_u_cla32_and6406_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6406_y0);
  and_gate and_gate_h_u_cla32_and6407_y0(h_u_cla32_and6406_y0, h_u_cla32_and6405_y0, h_u_cla32_and6407_y0);
  and_gate and_gate_h_u_cla32_and6408_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6408_y0);
  and_gate and_gate_h_u_cla32_and6409_y0(h_u_cla32_and6408_y0, h_u_cla32_and6407_y0, h_u_cla32_and6409_y0);
  and_gate and_gate_h_u_cla32_and6410_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6410_y0);
  and_gate and_gate_h_u_cla32_and6411_y0(h_u_cla32_and6410_y0, h_u_cla32_and6409_y0, h_u_cla32_and6411_y0);
  and_gate and_gate_h_u_cla32_and6412_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6412_y0);
  and_gate and_gate_h_u_cla32_and6413_y0(h_u_cla32_and6412_y0, h_u_cla32_and6411_y0, h_u_cla32_and6413_y0);
  and_gate and_gate_h_u_cla32_and6414_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6414_y0);
  and_gate and_gate_h_u_cla32_and6415_y0(h_u_cla32_and6414_y0, h_u_cla32_and6413_y0, h_u_cla32_and6415_y0);
  and_gate and_gate_h_u_cla32_and6416_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6416_y0);
  and_gate and_gate_h_u_cla32_and6417_y0(h_u_cla32_and6416_y0, h_u_cla32_and6415_y0, h_u_cla32_and6417_y0);
  and_gate and_gate_h_u_cla32_and6418_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6418_y0);
  and_gate and_gate_h_u_cla32_and6419_y0(h_u_cla32_and6418_y0, h_u_cla32_and6417_y0, h_u_cla32_and6419_y0);
  and_gate and_gate_h_u_cla32_and6420_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6420_y0);
  and_gate and_gate_h_u_cla32_and6421_y0(h_u_cla32_and6420_y0, h_u_cla32_and6419_y0, h_u_cla32_and6421_y0);
  and_gate and_gate_h_u_cla32_and6422_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6422_y0);
  and_gate and_gate_h_u_cla32_and6423_y0(h_u_cla32_and6422_y0, h_u_cla32_and6421_y0, h_u_cla32_and6423_y0);
  and_gate and_gate_h_u_cla32_and6424_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6424_y0);
  and_gate and_gate_h_u_cla32_and6425_y0(h_u_cla32_and6424_y0, h_u_cla32_and6423_y0, h_u_cla32_and6425_y0);
  and_gate and_gate_h_u_cla32_and6426_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6426_y0);
  and_gate and_gate_h_u_cla32_and6427_y0(h_u_cla32_and6426_y0, h_u_cla32_and6425_y0, h_u_cla32_and6427_y0);
  and_gate and_gate_h_u_cla32_and6428_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6428_y0);
  and_gate and_gate_h_u_cla32_and6429_y0(h_u_cla32_and6428_y0, h_u_cla32_and6427_y0, h_u_cla32_and6429_y0);
  and_gate and_gate_h_u_cla32_and6430_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6430_y0);
  and_gate and_gate_h_u_cla32_and6431_y0(h_u_cla32_and6430_y0, h_u_cla32_and6429_y0, h_u_cla32_and6431_y0);
  and_gate and_gate_h_u_cla32_and6432_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6432_y0);
  and_gate and_gate_h_u_cla32_and6433_y0(h_u_cla32_and6432_y0, h_u_cla32_and6431_y0, h_u_cla32_and6433_y0);
  and_gate and_gate_h_u_cla32_and6434_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6434_y0);
  and_gate and_gate_h_u_cla32_and6435_y0(h_u_cla32_and6434_y0, h_u_cla32_and6433_y0, h_u_cla32_and6435_y0);
  and_gate and_gate_h_u_cla32_and6436_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6436_y0);
  and_gate and_gate_h_u_cla32_and6437_y0(h_u_cla32_and6436_y0, h_u_cla32_and6435_y0, h_u_cla32_and6437_y0);
  and_gate and_gate_h_u_cla32_and6438_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6438_y0);
  and_gate and_gate_h_u_cla32_and6439_y0(h_u_cla32_and6438_y0, h_u_cla32_and6437_y0, h_u_cla32_and6439_y0);
  and_gate and_gate_h_u_cla32_and6440_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6440_y0);
  and_gate and_gate_h_u_cla32_and6441_y0(h_u_cla32_and6440_y0, h_u_cla32_and6439_y0, h_u_cla32_and6441_y0);
  and_gate and_gate_h_u_cla32_and6442_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6442_y0);
  and_gate and_gate_h_u_cla32_and6443_y0(h_u_cla32_and6442_y0, h_u_cla32_and6441_y0, h_u_cla32_and6443_y0);
  and_gate and_gate_h_u_cla32_and6444_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and6444_y0);
  and_gate and_gate_h_u_cla32_and6445_y0(h_u_cla32_and6444_y0, h_u_cla32_and6443_y0, h_u_cla32_and6445_y0);
  and_gate and_gate_h_u_cla32_and6446_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6446_y0);
  and_gate and_gate_h_u_cla32_and6447_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6447_y0);
  and_gate and_gate_h_u_cla32_and6448_y0(h_u_cla32_and6447_y0, h_u_cla32_and6446_y0, h_u_cla32_and6448_y0);
  and_gate and_gate_h_u_cla32_and6449_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6449_y0);
  and_gate and_gate_h_u_cla32_and6450_y0(h_u_cla32_and6449_y0, h_u_cla32_and6448_y0, h_u_cla32_and6450_y0);
  and_gate and_gate_h_u_cla32_and6451_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6451_y0);
  and_gate and_gate_h_u_cla32_and6452_y0(h_u_cla32_and6451_y0, h_u_cla32_and6450_y0, h_u_cla32_and6452_y0);
  and_gate and_gate_h_u_cla32_and6453_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6453_y0);
  and_gate and_gate_h_u_cla32_and6454_y0(h_u_cla32_and6453_y0, h_u_cla32_and6452_y0, h_u_cla32_and6454_y0);
  and_gate and_gate_h_u_cla32_and6455_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6455_y0);
  and_gate and_gate_h_u_cla32_and6456_y0(h_u_cla32_and6455_y0, h_u_cla32_and6454_y0, h_u_cla32_and6456_y0);
  and_gate and_gate_h_u_cla32_and6457_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6457_y0);
  and_gate and_gate_h_u_cla32_and6458_y0(h_u_cla32_and6457_y0, h_u_cla32_and6456_y0, h_u_cla32_and6458_y0);
  and_gate and_gate_h_u_cla32_and6459_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6459_y0);
  and_gate and_gate_h_u_cla32_and6460_y0(h_u_cla32_and6459_y0, h_u_cla32_and6458_y0, h_u_cla32_and6460_y0);
  and_gate and_gate_h_u_cla32_and6461_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6461_y0);
  and_gate and_gate_h_u_cla32_and6462_y0(h_u_cla32_and6461_y0, h_u_cla32_and6460_y0, h_u_cla32_and6462_y0);
  and_gate and_gate_h_u_cla32_and6463_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6463_y0);
  and_gate and_gate_h_u_cla32_and6464_y0(h_u_cla32_and6463_y0, h_u_cla32_and6462_y0, h_u_cla32_and6464_y0);
  and_gate and_gate_h_u_cla32_and6465_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6465_y0);
  and_gate and_gate_h_u_cla32_and6466_y0(h_u_cla32_and6465_y0, h_u_cla32_and6464_y0, h_u_cla32_and6466_y0);
  and_gate and_gate_h_u_cla32_and6467_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6467_y0);
  and_gate and_gate_h_u_cla32_and6468_y0(h_u_cla32_and6467_y0, h_u_cla32_and6466_y0, h_u_cla32_and6468_y0);
  and_gate and_gate_h_u_cla32_and6469_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6469_y0);
  and_gate and_gate_h_u_cla32_and6470_y0(h_u_cla32_and6469_y0, h_u_cla32_and6468_y0, h_u_cla32_and6470_y0);
  and_gate and_gate_h_u_cla32_and6471_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6471_y0);
  and_gate and_gate_h_u_cla32_and6472_y0(h_u_cla32_and6471_y0, h_u_cla32_and6470_y0, h_u_cla32_and6472_y0);
  and_gate and_gate_h_u_cla32_and6473_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6473_y0);
  and_gate and_gate_h_u_cla32_and6474_y0(h_u_cla32_and6473_y0, h_u_cla32_and6472_y0, h_u_cla32_and6474_y0);
  and_gate and_gate_h_u_cla32_and6475_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6475_y0);
  and_gate and_gate_h_u_cla32_and6476_y0(h_u_cla32_and6475_y0, h_u_cla32_and6474_y0, h_u_cla32_and6476_y0);
  and_gate and_gate_h_u_cla32_and6477_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6477_y0);
  and_gate and_gate_h_u_cla32_and6478_y0(h_u_cla32_and6477_y0, h_u_cla32_and6476_y0, h_u_cla32_and6478_y0);
  and_gate and_gate_h_u_cla32_and6479_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6479_y0);
  and_gate and_gate_h_u_cla32_and6480_y0(h_u_cla32_and6479_y0, h_u_cla32_and6478_y0, h_u_cla32_and6480_y0);
  and_gate and_gate_h_u_cla32_and6481_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6481_y0);
  and_gate and_gate_h_u_cla32_and6482_y0(h_u_cla32_and6481_y0, h_u_cla32_and6480_y0, h_u_cla32_and6482_y0);
  and_gate and_gate_h_u_cla32_and6483_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6483_y0);
  and_gate and_gate_h_u_cla32_and6484_y0(h_u_cla32_and6483_y0, h_u_cla32_and6482_y0, h_u_cla32_and6484_y0);
  and_gate and_gate_h_u_cla32_and6485_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6485_y0);
  and_gate and_gate_h_u_cla32_and6486_y0(h_u_cla32_and6485_y0, h_u_cla32_and6484_y0, h_u_cla32_and6486_y0);
  and_gate and_gate_h_u_cla32_and6487_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and6487_y0);
  and_gate and_gate_h_u_cla32_and6488_y0(h_u_cla32_and6487_y0, h_u_cla32_and6486_y0, h_u_cla32_and6488_y0);
  and_gate and_gate_h_u_cla32_and6489_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6489_y0);
  and_gate and_gate_h_u_cla32_and6490_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6490_y0);
  and_gate and_gate_h_u_cla32_and6491_y0(h_u_cla32_and6490_y0, h_u_cla32_and6489_y0, h_u_cla32_and6491_y0);
  and_gate and_gate_h_u_cla32_and6492_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6492_y0);
  and_gate and_gate_h_u_cla32_and6493_y0(h_u_cla32_and6492_y0, h_u_cla32_and6491_y0, h_u_cla32_and6493_y0);
  and_gate and_gate_h_u_cla32_and6494_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6494_y0);
  and_gate and_gate_h_u_cla32_and6495_y0(h_u_cla32_and6494_y0, h_u_cla32_and6493_y0, h_u_cla32_and6495_y0);
  and_gate and_gate_h_u_cla32_and6496_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6496_y0);
  and_gate and_gate_h_u_cla32_and6497_y0(h_u_cla32_and6496_y0, h_u_cla32_and6495_y0, h_u_cla32_and6497_y0);
  and_gate and_gate_h_u_cla32_and6498_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6498_y0);
  and_gate and_gate_h_u_cla32_and6499_y0(h_u_cla32_and6498_y0, h_u_cla32_and6497_y0, h_u_cla32_and6499_y0);
  and_gate and_gate_h_u_cla32_and6500_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6500_y0);
  and_gate and_gate_h_u_cla32_and6501_y0(h_u_cla32_and6500_y0, h_u_cla32_and6499_y0, h_u_cla32_and6501_y0);
  and_gate and_gate_h_u_cla32_and6502_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6502_y0);
  and_gate and_gate_h_u_cla32_and6503_y0(h_u_cla32_and6502_y0, h_u_cla32_and6501_y0, h_u_cla32_and6503_y0);
  and_gate and_gate_h_u_cla32_and6504_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6504_y0);
  and_gate and_gate_h_u_cla32_and6505_y0(h_u_cla32_and6504_y0, h_u_cla32_and6503_y0, h_u_cla32_and6505_y0);
  and_gate and_gate_h_u_cla32_and6506_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6506_y0);
  and_gate and_gate_h_u_cla32_and6507_y0(h_u_cla32_and6506_y0, h_u_cla32_and6505_y0, h_u_cla32_and6507_y0);
  and_gate and_gate_h_u_cla32_and6508_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6508_y0);
  and_gate and_gate_h_u_cla32_and6509_y0(h_u_cla32_and6508_y0, h_u_cla32_and6507_y0, h_u_cla32_and6509_y0);
  and_gate and_gate_h_u_cla32_and6510_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6510_y0);
  and_gate and_gate_h_u_cla32_and6511_y0(h_u_cla32_and6510_y0, h_u_cla32_and6509_y0, h_u_cla32_and6511_y0);
  and_gate and_gate_h_u_cla32_and6512_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6512_y0);
  and_gate and_gate_h_u_cla32_and6513_y0(h_u_cla32_and6512_y0, h_u_cla32_and6511_y0, h_u_cla32_and6513_y0);
  and_gate and_gate_h_u_cla32_and6514_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6514_y0);
  and_gate and_gate_h_u_cla32_and6515_y0(h_u_cla32_and6514_y0, h_u_cla32_and6513_y0, h_u_cla32_and6515_y0);
  and_gate and_gate_h_u_cla32_and6516_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6516_y0);
  and_gate and_gate_h_u_cla32_and6517_y0(h_u_cla32_and6516_y0, h_u_cla32_and6515_y0, h_u_cla32_and6517_y0);
  and_gate and_gate_h_u_cla32_and6518_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6518_y0);
  and_gate and_gate_h_u_cla32_and6519_y0(h_u_cla32_and6518_y0, h_u_cla32_and6517_y0, h_u_cla32_and6519_y0);
  and_gate and_gate_h_u_cla32_and6520_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6520_y0);
  and_gate and_gate_h_u_cla32_and6521_y0(h_u_cla32_and6520_y0, h_u_cla32_and6519_y0, h_u_cla32_and6521_y0);
  and_gate and_gate_h_u_cla32_and6522_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6522_y0);
  and_gate and_gate_h_u_cla32_and6523_y0(h_u_cla32_and6522_y0, h_u_cla32_and6521_y0, h_u_cla32_and6523_y0);
  and_gate and_gate_h_u_cla32_and6524_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6524_y0);
  and_gate and_gate_h_u_cla32_and6525_y0(h_u_cla32_and6524_y0, h_u_cla32_and6523_y0, h_u_cla32_and6525_y0);
  and_gate and_gate_h_u_cla32_and6526_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6526_y0);
  and_gate and_gate_h_u_cla32_and6527_y0(h_u_cla32_and6526_y0, h_u_cla32_and6525_y0, h_u_cla32_and6527_y0);
  and_gate and_gate_h_u_cla32_and6528_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and6528_y0);
  and_gate and_gate_h_u_cla32_and6529_y0(h_u_cla32_and6528_y0, h_u_cla32_and6527_y0, h_u_cla32_and6529_y0);
  and_gate and_gate_h_u_cla32_and6530_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6530_y0);
  and_gate and_gate_h_u_cla32_and6531_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6531_y0);
  and_gate and_gate_h_u_cla32_and6532_y0(h_u_cla32_and6531_y0, h_u_cla32_and6530_y0, h_u_cla32_and6532_y0);
  and_gate and_gate_h_u_cla32_and6533_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6533_y0);
  and_gate and_gate_h_u_cla32_and6534_y0(h_u_cla32_and6533_y0, h_u_cla32_and6532_y0, h_u_cla32_and6534_y0);
  and_gate and_gate_h_u_cla32_and6535_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6535_y0);
  and_gate and_gate_h_u_cla32_and6536_y0(h_u_cla32_and6535_y0, h_u_cla32_and6534_y0, h_u_cla32_and6536_y0);
  and_gate and_gate_h_u_cla32_and6537_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6537_y0);
  and_gate and_gate_h_u_cla32_and6538_y0(h_u_cla32_and6537_y0, h_u_cla32_and6536_y0, h_u_cla32_and6538_y0);
  and_gate and_gate_h_u_cla32_and6539_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6539_y0);
  and_gate and_gate_h_u_cla32_and6540_y0(h_u_cla32_and6539_y0, h_u_cla32_and6538_y0, h_u_cla32_and6540_y0);
  and_gate and_gate_h_u_cla32_and6541_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6541_y0);
  and_gate and_gate_h_u_cla32_and6542_y0(h_u_cla32_and6541_y0, h_u_cla32_and6540_y0, h_u_cla32_and6542_y0);
  and_gate and_gate_h_u_cla32_and6543_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6543_y0);
  and_gate and_gate_h_u_cla32_and6544_y0(h_u_cla32_and6543_y0, h_u_cla32_and6542_y0, h_u_cla32_and6544_y0);
  and_gate and_gate_h_u_cla32_and6545_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6545_y0);
  and_gate and_gate_h_u_cla32_and6546_y0(h_u_cla32_and6545_y0, h_u_cla32_and6544_y0, h_u_cla32_and6546_y0);
  and_gate and_gate_h_u_cla32_and6547_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6547_y0);
  and_gate and_gate_h_u_cla32_and6548_y0(h_u_cla32_and6547_y0, h_u_cla32_and6546_y0, h_u_cla32_and6548_y0);
  and_gate and_gate_h_u_cla32_and6549_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6549_y0);
  and_gate and_gate_h_u_cla32_and6550_y0(h_u_cla32_and6549_y0, h_u_cla32_and6548_y0, h_u_cla32_and6550_y0);
  and_gate and_gate_h_u_cla32_and6551_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6551_y0);
  and_gate and_gate_h_u_cla32_and6552_y0(h_u_cla32_and6551_y0, h_u_cla32_and6550_y0, h_u_cla32_and6552_y0);
  and_gate and_gate_h_u_cla32_and6553_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6553_y0);
  and_gate and_gate_h_u_cla32_and6554_y0(h_u_cla32_and6553_y0, h_u_cla32_and6552_y0, h_u_cla32_and6554_y0);
  and_gate and_gate_h_u_cla32_and6555_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6555_y0);
  and_gate and_gate_h_u_cla32_and6556_y0(h_u_cla32_and6555_y0, h_u_cla32_and6554_y0, h_u_cla32_and6556_y0);
  and_gate and_gate_h_u_cla32_and6557_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6557_y0);
  and_gate and_gate_h_u_cla32_and6558_y0(h_u_cla32_and6557_y0, h_u_cla32_and6556_y0, h_u_cla32_and6558_y0);
  and_gate and_gate_h_u_cla32_and6559_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6559_y0);
  and_gate and_gate_h_u_cla32_and6560_y0(h_u_cla32_and6559_y0, h_u_cla32_and6558_y0, h_u_cla32_and6560_y0);
  and_gate and_gate_h_u_cla32_and6561_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6561_y0);
  and_gate and_gate_h_u_cla32_and6562_y0(h_u_cla32_and6561_y0, h_u_cla32_and6560_y0, h_u_cla32_and6562_y0);
  and_gate and_gate_h_u_cla32_and6563_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6563_y0);
  and_gate and_gate_h_u_cla32_and6564_y0(h_u_cla32_and6563_y0, h_u_cla32_and6562_y0, h_u_cla32_and6564_y0);
  and_gate and_gate_h_u_cla32_and6565_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6565_y0);
  and_gate and_gate_h_u_cla32_and6566_y0(h_u_cla32_and6565_y0, h_u_cla32_and6564_y0, h_u_cla32_and6566_y0);
  and_gate and_gate_h_u_cla32_and6567_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and6567_y0);
  and_gate and_gate_h_u_cla32_and6568_y0(h_u_cla32_and6567_y0, h_u_cla32_and6566_y0, h_u_cla32_and6568_y0);
  and_gate and_gate_h_u_cla32_and6569_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6569_y0);
  and_gate and_gate_h_u_cla32_and6570_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6570_y0);
  and_gate and_gate_h_u_cla32_and6571_y0(h_u_cla32_and6570_y0, h_u_cla32_and6569_y0, h_u_cla32_and6571_y0);
  and_gate and_gate_h_u_cla32_and6572_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6572_y0);
  and_gate and_gate_h_u_cla32_and6573_y0(h_u_cla32_and6572_y0, h_u_cla32_and6571_y0, h_u_cla32_and6573_y0);
  and_gate and_gate_h_u_cla32_and6574_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6574_y0);
  and_gate and_gate_h_u_cla32_and6575_y0(h_u_cla32_and6574_y0, h_u_cla32_and6573_y0, h_u_cla32_and6575_y0);
  and_gate and_gate_h_u_cla32_and6576_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6576_y0);
  and_gate and_gate_h_u_cla32_and6577_y0(h_u_cla32_and6576_y0, h_u_cla32_and6575_y0, h_u_cla32_and6577_y0);
  and_gate and_gate_h_u_cla32_and6578_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6578_y0);
  and_gate and_gate_h_u_cla32_and6579_y0(h_u_cla32_and6578_y0, h_u_cla32_and6577_y0, h_u_cla32_and6579_y0);
  and_gate and_gate_h_u_cla32_and6580_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6580_y0);
  and_gate and_gate_h_u_cla32_and6581_y0(h_u_cla32_and6580_y0, h_u_cla32_and6579_y0, h_u_cla32_and6581_y0);
  and_gate and_gate_h_u_cla32_and6582_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6582_y0);
  and_gate and_gate_h_u_cla32_and6583_y0(h_u_cla32_and6582_y0, h_u_cla32_and6581_y0, h_u_cla32_and6583_y0);
  and_gate and_gate_h_u_cla32_and6584_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6584_y0);
  and_gate and_gate_h_u_cla32_and6585_y0(h_u_cla32_and6584_y0, h_u_cla32_and6583_y0, h_u_cla32_and6585_y0);
  and_gate and_gate_h_u_cla32_and6586_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6586_y0);
  and_gate and_gate_h_u_cla32_and6587_y0(h_u_cla32_and6586_y0, h_u_cla32_and6585_y0, h_u_cla32_and6587_y0);
  and_gate and_gate_h_u_cla32_and6588_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6588_y0);
  and_gate and_gate_h_u_cla32_and6589_y0(h_u_cla32_and6588_y0, h_u_cla32_and6587_y0, h_u_cla32_and6589_y0);
  and_gate and_gate_h_u_cla32_and6590_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6590_y0);
  and_gate and_gate_h_u_cla32_and6591_y0(h_u_cla32_and6590_y0, h_u_cla32_and6589_y0, h_u_cla32_and6591_y0);
  and_gate and_gate_h_u_cla32_and6592_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6592_y0);
  and_gate and_gate_h_u_cla32_and6593_y0(h_u_cla32_and6592_y0, h_u_cla32_and6591_y0, h_u_cla32_and6593_y0);
  and_gate and_gate_h_u_cla32_and6594_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6594_y0);
  and_gate and_gate_h_u_cla32_and6595_y0(h_u_cla32_and6594_y0, h_u_cla32_and6593_y0, h_u_cla32_and6595_y0);
  and_gate and_gate_h_u_cla32_and6596_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6596_y0);
  and_gate and_gate_h_u_cla32_and6597_y0(h_u_cla32_and6596_y0, h_u_cla32_and6595_y0, h_u_cla32_and6597_y0);
  and_gate and_gate_h_u_cla32_and6598_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6598_y0);
  and_gate and_gate_h_u_cla32_and6599_y0(h_u_cla32_and6598_y0, h_u_cla32_and6597_y0, h_u_cla32_and6599_y0);
  and_gate and_gate_h_u_cla32_and6600_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6600_y0);
  and_gate and_gate_h_u_cla32_and6601_y0(h_u_cla32_and6600_y0, h_u_cla32_and6599_y0, h_u_cla32_and6601_y0);
  and_gate and_gate_h_u_cla32_and6602_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6602_y0);
  and_gate and_gate_h_u_cla32_and6603_y0(h_u_cla32_and6602_y0, h_u_cla32_and6601_y0, h_u_cla32_and6603_y0);
  and_gate and_gate_h_u_cla32_and6604_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and6604_y0);
  and_gate and_gate_h_u_cla32_and6605_y0(h_u_cla32_and6604_y0, h_u_cla32_and6603_y0, h_u_cla32_and6605_y0);
  and_gate and_gate_h_u_cla32_and6606_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6606_y0);
  and_gate and_gate_h_u_cla32_and6607_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6607_y0);
  and_gate and_gate_h_u_cla32_and6608_y0(h_u_cla32_and6607_y0, h_u_cla32_and6606_y0, h_u_cla32_and6608_y0);
  and_gate and_gate_h_u_cla32_and6609_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6609_y0);
  and_gate and_gate_h_u_cla32_and6610_y0(h_u_cla32_and6609_y0, h_u_cla32_and6608_y0, h_u_cla32_and6610_y0);
  and_gate and_gate_h_u_cla32_and6611_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6611_y0);
  and_gate and_gate_h_u_cla32_and6612_y0(h_u_cla32_and6611_y0, h_u_cla32_and6610_y0, h_u_cla32_and6612_y0);
  and_gate and_gate_h_u_cla32_and6613_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6613_y0);
  and_gate and_gate_h_u_cla32_and6614_y0(h_u_cla32_and6613_y0, h_u_cla32_and6612_y0, h_u_cla32_and6614_y0);
  and_gate and_gate_h_u_cla32_and6615_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6615_y0);
  and_gate and_gate_h_u_cla32_and6616_y0(h_u_cla32_and6615_y0, h_u_cla32_and6614_y0, h_u_cla32_and6616_y0);
  and_gate and_gate_h_u_cla32_and6617_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6617_y0);
  and_gate and_gate_h_u_cla32_and6618_y0(h_u_cla32_and6617_y0, h_u_cla32_and6616_y0, h_u_cla32_and6618_y0);
  and_gate and_gate_h_u_cla32_and6619_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6619_y0);
  and_gate and_gate_h_u_cla32_and6620_y0(h_u_cla32_and6619_y0, h_u_cla32_and6618_y0, h_u_cla32_and6620_y0);
  and_gate and_gate_h_u_cla32_and6621_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6621_y0);
  and_gate and_gate_h_u_cla32_and6622_y0(h_u_cla32_and6621_y0, h_u_cla32_and6620_y0, h_u_cla32_and6622_y0);
  and_gate and_gate_h_u_cla32_and6623_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6623_y0);
  and_gate and_gate_h_u_cla32_and6624_y0(h_u_cla32_and6623_y0, h_u_cla32_and6622_y0, h_u_cla32_and6624_y0);
  and_gate and_gate_h_u_cla32_and6625_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6625_y0);
  and_gate and_gate_h_u_cla32_and6626_y0(h_u_cla32_and6625_y0, h_u_cla32_and6624_y0, h_u_cla32_and6626_y0);
  and_gate and_gate_h_u_cla32_and6627_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6627_y0);
  and_gate and_gate_h_u_cla32_and6628_y0(h_u_cla32_and6627_y0, h_u_cla32_and6626_y0, h_u_cla32_and6628_y0);
  and_gate and_gate_h_u_cla32_and6629_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6629_y0);
  and_gate and_gate_h_u_cla32_and6630_y0(h_u_cla32_and6629_y0, h_u_cla32_and6628_y0, h_u_cla32_and6630_y0);
  and_gate and_gate_h_u_cla32_and6631_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6631_y0);
  and_gate and_gate_h_u_cla32_and6632_y0(h_u_cla32_and6631_y0, h_u_cla32_and6630_y0, h_u_cla32_and6632_y0);
  and_gate and_gate_h_u_cla32_and6633_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6633_y0);
  and_gate and_gate_h_u_cla32_and6634_y0(h_u_cla32_and6633_y0, h_u_cla32_and6632_y0, h_u_cla32_and6634_y0);
  and_gate and_gate_h_u_cla32_and6635_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6635_y0);
  and_gate and_gate_h_u_cla32_and6636_y0(h_u_cla32_and6635_y0, h_u_cla32_and6634_y0, h_u_cla32_and6636_y0);
  and_gate and_gate_h_u_cla32_and6637_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6637_y0);
  and_gate and_gate_h_u_cla32_and6638_y0(h_u_cla32_and6637_y0, h_u_cla32_and6636_y0, h_u_cla32_and6638_y0);
  and_gate and_gate_h_u_cla32_and6639_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and6639_y0);
  and_gate and_gate_h_u_cla32_and6640_y0(h_u_cla32_and6639_y0, h_u_cla32_and6638_y0, h_u_cla32_and6640_y0);
  and_gate and_gate_h_u_cla32_and6641_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6641_y0);
  and_gate and_gate_h_u_cla32_and6642_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6642_y0);
  and_gate and_gate_h_u_cla32_and6643_y0(h_u_cla32_and6642_y0, h_u_cla32_and6641_y0, h_u_cla32_and6643_y0);
  and_gate and_gate_h_u_cla32_and6644_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6644_y0);
  and_gate and_gate_h_u_cla32_and6645_y0(h_u_cla32_and6644_y0, h_u_cla32_and6643_y0, h_u_cla32_and6645_y0);
  and_gate and_gate_h_u_cla32_and6646_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6646_y0);
  and_gate and_gate_h_u_cla32_and6647_y0(h_u_cla32_and6646_y0, h_u_cla32_and6645_y0, h_u_cla32_and6647_y0);
  and_gate and_gate_h_u_cla32_and6648_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6648_y0);
  and_gate and_gate_h_u_cla32_and6649_y0(h_u_cla32_and6648_y0, h_u_cla32_and6647_y0, h_u_cla32_and6649_y0);
  and_gate and_gate_h_u_cla32_and6650_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6650_y0);
  and_gate and_gate_h_u_cla32_and6651_y0(h_u_cla32_and6650_y0, h_u_cla32_and6649_y0, h_u_cla32_and6651_y0);
  and_gate and_gate_h_u_cla32_and6652_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6652_y0);
  and_gate and_gate_h_u_cla32_and6653_y0(h_u_cla32_and6652_y0, h_u_cla32_and6651_y0, h_u_cla32_and6653_y0);
  and_gate and_gate_h_u_cla32_and6654_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6654_y0);
  and_gate and_gate_h_u_cla32_and6655_y0(h_u_cla32_and6654_y0, h_u_cla32_and6653_y0, h_u_cla32_and6655_y0);
  and_gate and_gate_h_u_cla32_and6656_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6656_y0);
  and_gate and_gate_h_u_cla32_and6657_y0(h_u_cla32_and6656_y0, h_u_cla32_and6655_y0, h_u_cla32_and6657_y0);
  and_gate and_gate_h_u_cla32_and6658_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6658_y0);
  and_gate and_gate_h_u_cla32_and6659_y0(h_u_cla32_and6658_y0, h_u_cla32_and6657_y0, h_u_cla32_and6659_y0);
  and_gate and_gate_h_u_cla32_and6660_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6660_y0);
  and_gate and_gate_h_u_cla32_and6661_y0(h_u_cla32_and6660_y0, h_u_cla32_and6659_y0, h_u_cla32_and6661_y0);
  and_gate and_gate_h_u_cla32_and6662_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6662_y0);
  and_gate and_gate_h_u_cla32_and6663_y0(h_u_cla32_and6662_y0, h_u_cla32_and6661_y0, h_u_cla32_and6663_y0);
  and_gate and_gate_h_u_cla32_and6664_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6664_y0);
  and_gate and_gate_h_u_cla32_and6665_y0(h_u_cla32_and6664_y0, h_u_cla32_and6663_y0, h_u_cla32_and6665_y0);
  and_gate and_gate_h_u_cla32_and6666_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6666_y0);
  and_gate and_gate_h_u_cla32_and6667_y0(h_u_cla32_and6666_y0, h_u_cla32_and6665_y0, h_u_cla32_and6667_y0);
  and_gate and_gate_h_u_cla32_and6668_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6668_y0);
  and_gate and_gate_h_u_cla32_and6669_y0(h_u_cla32_and6668_y0, h_u_cla32_and6667_y0, h_u_cla32_and6669_y0);
  and_gate and_gate_h_u_cla32_and6670_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6670_y0);
  and_gate and_gate_h_u_cla32_and6671_y0(h_u_cla32_and6670_y0, h_u_cla32_and6669_y0, h_u_cla32_and6671_y0);
  and_gate and_gate_h_u_cla32_and6672_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and6672_y0);
  and_gate and_gate_h_u_cla32_and6673_y0(h_u_cla32_and6672_y0, h_u_cla32_and6671_y0, h_u_cla32_and6673_y0);
  and_gate and_gate_h_u_cla32_and6674_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6674_y0);
  and_gate and_gate_h_u_cla32_and6675_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6675_y0);
  and_gate and_gate_h_u_cla32_and6676_y0(h_u_cla32_and6675_y0, h_u_cla32_and6674_y0, h_u_cla32_and6676_y0);
  and_gate and_gate_h_u_cla32_and6677_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6677_y0);
  and_gate and_gate_h_u_cla32_and6678_y0(h_u_cla32_and6677_y0, h_u_cla32_and6676_y0, h_u_cla32_and6678_y0);
  and_gate and_gate_h_u_cla32_and6679_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6679_y0);
  and_gate and_gate_h_u_cla32_and6680_y0(h_u_cla32_and6679_y0, h_u_cla32_and6678_y0, h_u_cla32_and6680_y0);
  and_gate and_gate_h_u_cla32_and6681_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6681_y0);
  and_gate and_gate_h_u_cla32_and6682_y0(h_u_cla32_and6681_y0, h_u_cla32_and6680_y0, h_u_cla32_and6682_y0);
  and_gate and_gate_h_u_cla32_and6683_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6683_y0);
  and_gate and_gate_h_u_cla32_and6684_y0(h_u_cla32_and6683_y0, h_u_cla32_and6682_y0, h_u_cla32_and6684_y0);
  and_gate and_gate_h_u_cla32_and6685_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6685_y0);
  and_gate and_gate_h_u_cla32_and6686_y0(h_u_cla32_and6685_y0, h_u_cla32_and6684_y0, h_u_cla32_and6686_y0);
  and_gate and_gate_h_u_cla32_and6687_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6687_y0);
  and_gate and_gate_h_u_cla32_and6688_y0(h_u_cla32_and6687_y0, h_u_cla32_and6686_y0, h_u_cla32_and6688_y0);
  and_gate and_gate_h_u_cla32_and6689_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6689_y0);
  and_gate and_gate_h_u_cla32_and6690_y0(h_u_cla32_and6689_y0, h_u_cla32_and6688_y0, h_u_cla32_and6690_y0);
  and_gate and_gate_h_u_cla32_and6691_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6691_y0);
  and_gate and_gate_h_u_cla32_and6692_y0(h_u_cla32_and6691_y0, h_u_cla32_and6690_y0, h_u_cla32_and6692_y0);
  and_gate and_gate_h_u_cla32_and6693_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6693_y0);
  and_gate and_gate_h_u_cla32_and6694_y0(h_u_cla32_and6693_y0, h_u_cla32_and6692_y0, h_u_cla32_and6694_y0);
  and_gate and_gate_h_u_cla32_and6695_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6695_y0);
  and_gate and_gate_h_u_cla32_and6696_y0(h_u_cla32_and6695_y0, h_u_cla32_and6694_y0, h_u_cla32_and6696_y0);
  and_gate and_gate_h_u_cla32_and6697_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6697_y0);
  and_gate and_gate_h_u_cla32_and6698_y0(h_u_cla32_and6697_y0, h_u_cla32_and6696_y0, h_u_cla32_and6698_y0);
  and_gate and_gate_h_u_cla32_and6699_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6699_y0);
  and_gate and_gate_h_u_cla32_and6700_y0(h_u_cla32_and6699_y0, h_u_cla32_and6698_y0, h_u_cla32_and6700_y0);
  and_gate and_gate_h_u_cla32_and6701_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6701_y0);
  and_gate and_gate_h_u_cla32_and6702_y0(h_u_cla32_and6701_y0, h_u_cla32_and6700_y0, h_u_cla32_and6702_y0);
  and_gate and_gate_h_u_cla32_and6703_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and6703_y0);
  and_gate and_gate_h_u_cla32_and6704_y0(h_u_cla32_and6703_y0, h_u_cla32_and6702_y0, h_u_cla32_and6704_y0);
  and_gate and_gate_h_u_cla32_and6705_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6705_y0);
  and_gate and_gate_h_u_cla32_and6706_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6706_y0);
  and_gate and_gate_h_u_cla32_and6707_y0(h_u_cla32_and6706_y0, h_u_cla32_and6705_y0, h_u_cla32_and6707_y0);
  and_gate and_gate_h_u_cla32_and6708_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6708_y0);
  and_gate and_gate_h_u_cla32_and6709_y0(h_u_cla32_and6708_y0, h_u_cla32_and6707_y0, h_u_cla32_and6709_y0);
  and_gate and_gate_h_u_cla32_and6710_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6710_y0);
  and_gate and_gate_h_u_cla32_and6711_y0(h_u_cla32_and6710_y0, h_u_cla32_and6709_y0, h_u_cla32_and6711_y0);
  and_gate and_gate_h_u_cla32_and6712_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6712_y0);
  and_gate and_gate_h_u_cla32_and6713_y0(h_u_cla32_and6712_y0, h_u_cla32_and6711_y0, h_u_cla32_and6713_y0);
  and_gate and_gate_h_u_cla32_and6714_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6714_y0);
  and_gate and_gate_h_u_cla32_and6715_y0(h_u_cla32_and6714_y0, h_u_cla32_and6713_y0, h_u_cla32_and6715_y0);
  and_gate and_gate_h_u_cla32_and6716_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6716_y0);
  and_gate and_gate_h_u_cla32_and6717_y0(h_u_cla32_and6716_y0, h_u_cla32_and6715_y0, h_u_cla32_and6717_y0);
  and_gate and_gate_h_u_cla32_and6718_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6718_y0);
  and_gate and_gate_h_u_cla32_and6719_y0(h_u_cla32_and6718_y0, h_u_cla32_and6717_y0, h_u_cla32_and6719_y0);
  and_gate and_gate_h_u_cla32_and6720_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6720_y0);
  and_gate and_gate_h_u_cla32_and6721_y0(h_u_cla32_and6720_y0, h_u_cla32_and6719_y0, h_u_cla32_and6721_y0);
  and_gate and_gate_h_u_cla32_and6722_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6722_y0);
  and_gate and_gate_h_u_cla32_and6723_y0(h_u_cla32_and6722_y0, h_u_cla32_and6721_y0, h_u_cla32_and6723_y0);
  and_gate and_gate_h_u_cla32_and6724_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6724_y0);
  and_gate and_gate_h_u_cla32_and6725_y0(h_u_cla32_and6724_y0, h_u_cla32_and6723_y0, h_u_cla32_and6725_y0);
  and_gate and_gate_h_u_cla32_and6726_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6726_y0);
  and_gate and_gate_h_u_cla32_and6727_y0(h_u_cla32_and6726_y0, h_u_cla32_and6725_y0, h_u_cla32_and6727_y0);
  and_gate and_gate_h_u_cla32_and6728_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6728_y0);
  and_gate and_gate_h_u_cla32_and6729_y0(h_u_cla32_and6728_y0, h_u_cla32_and6727_y0, h_u_cla32_and6729_y0);
  and_gate and_gate_h_u_cla32_and6730_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6730_y0);
  and_gate and_gate_h_u_cla32_and6731_y0(h_u_cla32_and6730_y0, h_u_cla32_and6729_y0, h_u_cla32_and6731_y0);
  and_gate and_gate_h_u_cla32_and6732_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and6732_y0);
  and_gate and_gate_h_u_cla32_and6733_y0(h_u_cla32_and6732_y0, h_u_cla32_and6731_y0, h_u_cla32_and6733_y0);
  and_gate and_gate_h_u_cla32_and6734_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6734_y0);
  and_gate and_gate_h_u_cla32_and6735_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6735_y0);
  and_gate and_gate_h_u_cla32_and6736_y0(h_u_cla32_and6735_y0, h_u_cla32_and6734_y0, h_u_cla32_and6736_y0);
  and_gate and_gate_h_u_cla32_and6737_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6737_y0);
  and_gate and_gate_h_u_cla32_and6738_y0(h_u_cla32_and6737_y0, h_u_cla32_and6736_y0, h_u_cla32_and6738_y0);
  and_gate and_gate_h_u_cla32_and6739_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6739_y0);
  and_gate and_gate_h_u_cla32_and6740_y0(h_u_cla32_and6739_y0, h_u_cla32_and6738_y0, h_u_cla32_and6740_y0);
  and_gate and_gate_h_u_cla32_and6741_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6741_y0);
  and_gate and_gate_h_u_cla32_and6742_y0(h_u_cla32_and6741_y0, h_u_cla32_and6740_y0, h_u_cla32_and6742_y0);
  and_gate and_gate_h_u_cla32_and6743_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6743_y0);
  and_gate and_gate_h_u_cla32_and6744_y0(h_u_cla32_and6743_y0, h_u_cla32_and6742_y0, h_u_cla32_and6744_y0);
  and_gate and_gate_h_u_cla32_and6745_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6745_y0);
  and_gate and_gate_h_u_cla32_and6746_y0(h_u_cla32_and6745_y0, h_u_cla32_and6744_y0, h_u_cla32_and6746_y0);
  and_gate and_gate_h_u_cla32_and6747_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6747_y0);
  and_gate and_gate_h_u_cla32_and6748_y0(h_u_cla32_and6747_y0, h_u_cla32_and6746_y0, h_u_cla32_and6748_y0);
  and_gate and_gate_h_u_cla32_and6749_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6749_y0);
  and_gate and_gate_h_u_cla32_and6750_y0(h_u_cla32_and6749_y0, h_u_cla32_and6748_y0, h_u_cla32_and6750_y0);
  and_gate and_gate_h_u_cla32_and6751_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6751_y0);
  and_gate and_gate_h_u_cla32_and6752_y0(h_u_cla32_and6751_y0, h_u_cla32_and6750_y0, h_u_cla32_and6752_y0);
  and_gate and_gate_h_u_cla32_and6753_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6753_y0);
  and_gate and_gate_h_u_cla32_and6754_y0(h_u_cla32_and6753_y0, h_u_cla32_and6752_y0, h_u_cla32_and6754_y0);
  and_gate and_gate_h_u_cla32_and6755_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6755_y0);
  and_gate and_gate_h_u_cla32_and6756_y0(h_u_cla32_and6755_y0, h_u_cla32_and6754_y0, h_u_cla32_and6756_y0);
  and_gate and_gate_h_u_cla32_and6757_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6757_y0);
  and_gate and_gate_h_u_cla32_and6758_y0(h_u_cla32_and6757_y0, h_u_cla32_and6756_y0, h_u_cla32_and6758_y0);
  and_gate and_gate_h_u_cla32_and6759_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and6759_y0);
  and_gate and_gate_h_u_cla32_and6760_y0(h_u_cla32_and6759_y0, h_u_cla32_and6758_y0, h_u_cla32_and6760_y0);
  and_gate and_gate_h_u_cla32_and6761_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6761_y0);
  and_gate and_gate_h_u_cla32_and6762_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6762_y0);
  and_gate and_gate_h_u_cla32_and6763_y0(h_u_cla32_and6762_y0, h_u_cla32_and6761_y0, h_u_cla32_and6763_y0);
  and_gate and_gate_h_u_cla32_and6764_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6764_y0);
  and_gate and_gate_h_u_cla32_and6765_y0(h_u_cla32_and6764_y0, h_u_cla32_and6763_y0, h_u_cla32_and6765_y0);
  and_gate and_gate_h_u_cla32_and6766_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6766_y0);
  and_gate and_gate_h_u_cla32_and6767_y0(h_u_cla32_and6766_y0, h_u_cla32_and6765_y0, h_u_cla32_and6767_y0);
  and_gate and_gate_h_u_cla32_and6768_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6768_y0);
  and_gate and_gate_h_u_cla32_and6769_y0(h_u_cla32_and6768_y0, h_u_cla32_and6767_y0, h_u_cla32_and6769_y0);
  and_gate and_gate_h_u_cla32_and6770_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6770_y0);
  and_gate and_gate_h_u_cla32_and6771_y0(h_u_cla32_and6770_y0, h_u_cla32_and6769_y0, h_u_cla32_and6771_y0);
  and_gate and_gate_h_u_cla32_and6772_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6772_y0);
  and_gate and_gate_h_u_cla32_and6773_y0(h_u_cla32_and6772_y0, h_u_cla32_and6771_y0, h_u_cla32_and6773_y0);
  and_gate and_gate_h_u_cla32_and6774_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6774_y0);
  and_gate and_gate_h_u_cla32_and6775_y0(h_u_cla32_and6774_y0, h_u_cla32_and6773_y0, h_u_cla32_and6775_y0);
  and_gate and_gate_h_u_cla32_and6776_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6776_y0);
  and_gate and_gate_h_u_cla32_and6777_y0(h_u_cla32_and6776_y0, h_u_cla32_and6775_y0, h_u_cla32_and6777_y0);
  and_gate and_gate_h_u_cla32_and6778_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6778_y0);
  and_gate and_gate_h_u_cla32_and6779_y0(h_u_cla32_and6778_y0, h_u_cla32_and6777_y0, h_u_cla32_and6779_y0);
  and_gate and_gate_h_u_cla32_and6780_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6780_y0);
  and_gate and_gate_h_u_cla32_and6781_y0(h_u_cla32_and6780_y0, h_u_cla32_and6779_y0, h_u_cla32_and6781_y0);
  and_gate and_gate_h_u_cla32_and6782_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6782_y0);
  and_gate and_gate_h_u_cla32_and6783_y0(h_u_cla32_and6782_y0, h_u_cla32_and6781_y0, h_u_cla32_and6783_y0);
  and_gate and_gate_h_u_cla32_and6784_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and6784_y0);
  and_gate and_gate_h_u_cla32_and6785_y0(h_u_cla32_and6784_y0, h_u_cla32_and6783_y0, h_u_cla32_and6785_y0);
  and_gate and_gate_h_u_cla32_and6786_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6786_y0);
  and_gate and_gate_h_u_cla32_and6787_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6787_y0);
  and_gate and_gate_h_u_cla32_and6788_y0(h_u_cla32_and6787_y0, h_u_cla32_and6786_y0, h_u_cla32_and6788_y0);
  and_gate and_gate_h_u_cla32_and6789_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6789_y0);
  and_gate and_gate_h_u_cla32_and6790_y0(h_u_cla32_and6789_y0, h_u_cla32_and6788_y0, h_u_cla32_and6790_y0);
  and_gate and_gate_h_u_cla32_and6791_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6791_y0);
  and_gate and_gate_h_u_cla32_and6792_y0(h_u_cla32_and6791_y0, h_u_cla32_and6790_y0, h_u_cla32_and6792_y0);
  and_gate and_gate_h_u_cla32_and6793_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6793_y0);
  and_gate and_gate_h_u_cla32_and6794_y0(h_u_cla32_and6793_y0, h_u_cla32_and6792_y0, h_u_cla32_and6794_y0);
  and_gate and_gate_h_u_cla32_and6795_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6795_y0);
  and_gate and_gate_h_u_cla32_and6796_y0(h_u_cla32_and6795_y0, h_u_cla32_and6794_y0, h_u_cla32_and6796_y0);
  and_gate and_gate_h_u_cla32_and6797_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6797_y0);
  and_gate and_gate_h_u_cla32_and6798_y0(h_u_cla32_and6797_y0, h_u_cla32_and6796_y0, h_u_cla32_and6798_y0);
  and_gate and_gate_h_u_cla32_and6799_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6799_y0);
  and_gate and_gate_h_u_cla32_and6800_y0(h_u_cla32_and6799_y0, h_u_cla32_and6798_y0, h_u_cla32_and6800_y0);
  and_gate and_gate_h_u_cla32_and6801_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6801_y0);
  and_gate and_gate_h_u_cla32_and6802_y0(h_u_cla32_and6801_y0, h_u_cla32_and6800_y0, h_u_cla32_and6802_y0);
  and_gate and_gate_h_u_cla32_and6803_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6803_y0);
  and_gate and_gate_h_u_cla32_and6804_y0(h_u_cla32_and6803_y0, h_u_cla32_and6802_y0, h_u_cla32_and6804_y0);
  and_gate and_gate_h_u_cla32_and6805_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6805_y0);
  and_gate and_gate_h_u_cla32_and6806_y0(h_u_cla32_and6805_y0, h_u_cla32_and6804_y0, h_u_cla32_and6806_y0);
  and_gate and_gate_h_u_cla32_and6807_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and6807_y0);
  and_gate and_gate_h_u_cla32_and6808_y0(h_u_cla32_and6807_y0, h_u_cla32_and6806_y0, h_u_cla32_and6808_y0);
  and_gate and_gate_h_u_cla32_and6809_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6809_y0);
  and_gate and_gate_h_u_cla32_and6810_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6810_y0);
  and_gate and_gate_h_u_cla32_and6811_y0(h_u_cla32_and6810_y0, h_u_cla32_and6809_y0, h_u_cla32_and6811_y0);
  and_gate and_gate_h_u_cla32_and6812_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6812_y0);
  and_gate and_gate_h_u_cla32_and6813_y0(h_u_cla32_and6812_y0, h_u_cla32_and6811_y0, h_u_cla32_and6813_y0);
  and_gate and_gate_h_u_cla32_and6814_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6814_y0);
  and_gate and_gate_h_u_cla32_and6815_y0(h_u_cla32_and6814_y0, h_u_cla32_and6813_y0, h_u_cla32_and6815_y0);
  and_gate and_gate_h_u_cla32_and6816_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6816_y0);
  and_gate and_gate_h_u_cla32_and6817_y0(h_u_cla32_and6816_y0, h_u_cla32_and6815_y0, h_u_cla32_and6817_y0);
  and_gate and_gate_h_u_cla32_and6818_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6818_y0);
  and_gate and_gate_h_u_cla32_and6819_y0(h_u_cla32_and6818_y0, h_u_cla32_and6817_y0, h_u_cla32_and6819_y0);
  and_gate and_gate_h_u_cla32_and6820_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6820_y0);
  and_gate and_gate_h_u_cla32_and6821_y0(h_u_cla32_and6820_y0, h_u_cla32_and6819_y0, h_u_cla32_and6821_y0);
  and_gate and_gate_h_u_cla32_and6822_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6822_y0);
  and_gate and_gate_h_u_cla32_and6823_y0(h_u_cla32_and6822_y0, h_u_cla32_and6821_y0, h_u_cla32_and6823_y0);
  and_gate and_gate_h_u_cla32_and6824_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6824_y0);
  and_gate and_gate_h_u_cla32_and6825_y0(h_u_cla32_and6824_y0, h_u_cla32_and6823_y0, h_u_cla32_and6825_y0);
  and_gate and_gate_h_u_cla32_and6826_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6826_y0);
  and_gate and_gate_h_u_cla32_and6827_y0(h_u_cla32_and6826_y0, h_u_cla32_and6825_y0, h_u_cla32_and6827_y0);
  and_gate and_gate_h_u_cla32_and6828_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and6828_y0);
  and_gate and_gate_h_u_cla32_and6829_y0(h_u_cla32_and6828_y0, h_u_cla32_and6827_y0, h_u_cla32_and6829_y0);
  and_gate and_gate_h_u_cla32_and6830_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6830_y0);
  and_gate and_gate_h_u_cla32_and6831_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6831_y0);
  and_gate and_gate_h_u_cla32_and6832_y0(h_u_cla32_and6831_y0, h_u_cla32_and6830_y0, h_u_cla32_and6832_y0);
  and_gate and_gate_h_u_cla32_and6833_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6833_y0);
  and_gate and_gate_h_u_cla32_and6834_y0(h_u_cla32_and6833_y0, h_u_cla32_and6832_y0, h_u_cla32_and6834_y0);
  and_gate and_gate_h_u_cla32_and6835_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6835_y0);
  and_gate and_gate_h_u_cla32_and6836_y0(h_u_cla32_and6835_y0, h_u_cla32_and6834_y0, h_u_cla32_and6836_y0);
  and_gate and_gate_h_u_cla32_and6837_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6837_y0);
  and_gate and_gate_h_u_cla32_and6838_y0(h_u_cla32_and6837_y0, h_u_cla32_and6836_y0, h_u_cla32_and6838_y0);
  and_gate and_gate_h_u_cla32_and6839_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6839_y0);
  and_gate and_gate_h_u_cla32_and6840_y0(h_u_cla32_and6839_y0, h_u_cla32_and6838_y0, h_u_cla32_and6840_y0);
  and_gate and_gate_h_u_cla32_and6841_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6841_y0);
  and_gate and_gate_h_u_cla32_and6842_y0(h_u_cla32_and6841_y0, h_u_cla32_and6840_y0, h_u_cla32_and6842_y0);
  and_gate and_gate_h_u_cla32_and6843_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6843_y0);
  and_gate and_gate_h_u_cla32_and6844_y0(h_u_cla32_and6843_y0, h_u_cla32_and6842_y0, h_u_cla32_and6844_y0);
  and_gate and_gate_h_u_cla32_and6845_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6845_y0);
  and_gate and_gate_h_u_cla32_and6846_y0(h_u_cla32_and6845_y0, h_u_cla32_and6844_y0, h_u_cla32_and6846_y0);
  and_gate and_gate_h_u_cla32_and6847_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and6847_y0);
  and_gate and_gate_h_u_cla32_and6848_y0(h_u_cla32_and6847_y0, h_u_cla32_and6846_y0, h_u_cla32_and6848_y0);
  and_gate and_gate_h_u_cla32_and6849_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6849_y0);
  and_gate and_gate_h_u_cla32_and6850_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6850_y0);
  and_gate and_gate_h_u_cla32_and6851_y0(h_u_cla32_and6850_y0, h_u_cla32_and6849_y0, h_u_cla32_and6851_y0);
  and_gate and_gate_h_u_cla32_and6852_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6852_y0);
  and_gate and_gate_h_u_cla32_and6853_y0(h_u_cla32_and6852_y0, h_u_cla32_and6851_y0, h_u_cla32_and6853_y0);
  and_gate and_gate_h_u_cla32_and6854_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6854_y0);
  and_gate and_gate_h_u_cla32_and6855_y0(h_u_cla32_and6854_y0, h_u_cla32_and6853_y0, h_u_cla32_and6855_y0);
  and_gate and_gate_h_u_cla32_and6856_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6856_y0);
  and_gate and_gate_h_u_cla32_and6857_y0(h_u_cla32_and6856_y0, h_u_cla32_and6855_y0, h_u_cla32_and6857_y0);
  and_gate and_gate_h_u_cla32_and6858_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6858_y0);
  and_gate and_gate_h_u_cla32_and6859_y0(h_u_cla32_and6858_y0, h_u_cla32_and6857_y0, h_u_cla32_and6859_y0);
  and_gate and_gate_h_u_cla32_and6860_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6860_y0);
  and_gate and_gate_h_u_cla32_and6861_y0(h_u_cla32_and6860_y0, h_u_cla32_and6859_y0, h_u_cla32_and6861_y0);
  and_gate and_gate_h_u_cla32_and6862_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6862_y0);
  and_gate and_gate_h_u_cla32_and6863_y0(h_u_cla32_and6862_y0, h_u_cla32_and6861_y0, h_u_cla32_and6863_y0);
  and_gate and_gate_h_u_cla32_and6864_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and6864_y0);
  and_gate and_gate_h_u_cla32_and6865_y0(h_u_cla32_and6864_y0, h_u_cla32_and6863_y0, h_u_cla32_and6865_y0);
  and_gate and_gate_h_u_cla32_and6866_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6866_y0);
  and_gate and_gate_h_u_cla32_and6867_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6867_y0);
  and_gate and_gate_h_u_cla32_and6868_y0(h_u_cla32_and6867_y0, h_u_cla32_and6866_y0, h_u_cla32_and6868_y0);
  and_gate and_gate_h_u_cla32_and6869_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6869_y0);
  and_gate and_gate_h_u_cla32_and6870_y0(h_u_cla32_and6869_y0, h_u_cla32_and6868_y0, h_u_cla32_and6870_y0);
  and_gate and_gate_h_u_cla32_and6871_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6871_y0);
  and_gate and_gate_h_u_cla32_and6872_y0(h_u_cla32_and6871_y0, h_u_cla32_and6870_y0, h_u_cla32_and6872_y0);
  and_gate and_gate_h_u_cla32_and6873_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6873_y0);
  and_gate and_gate_h_u_cla32_and6874_y0(h_u_cla32_and6873_y0, h_u_cla32_and6872_y0, h_u_cla32_and6874_y0);
  and_gate and_gate_h_u_cla32_and6875_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6875_y0);
  and_gate and_gate_h_u_cla32_and6876_y0(h_u_cla32_and6875_y0, h_u_cla32_and6874_y0, h_u_cla32_and6876_y0);
  and_gate and_gate_h_u_cla32_and6877_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6877_y0);
  and_gate and_gate_h_u_cla32_and6878_y0(h_u_cla32_and6877_y0, h_u_cla32_and6876_y0, h_u_cla32_and6878_y0);
  and_gate and_gate_h_u_cla32_and6879_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and6879_y0);
  and_gate and_gate_h_u_cla32_and6880_y0(h_u_cla32_and6879_y0, h_u_cla32_and6878_y0, h_u_cla32_and6880_y0);
  and_gate and_gate_h_u_cla32_and6881_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6881_y0);
  and_gate and_gate_h_u_cla32_and6882_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6882_y0);
  and_gate and_gate_h_u_cla32_and6883_y0(h_u_cla32_and6882_y0, h_u_cla32_and6881_y0, h_u_cla32_and6883_y0);
  and_gate and_gate_h_u_cla32_and6884_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6884_y0);
  and_gate and_gate_h_u_cla32_and6885_y0(h_u_cla32_and6884_y0, h_u_cla32_and6883_y0, h_u_cla32_and6885_y0);
  and_gate and_gate_h_u_cla32_and6886_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6886_y0);
  and_gate and_gate_h_u_cla32_and6887_y0(h_u_cla32_and6886_y0, h_u_cla32_and6885_y0, h_u_cla32_and6887_y0);
  and_gate and_gate_h_u_cla32_and6888_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6888_y0);
  and_gate and_gate_h_u_cla32_and6889_y0(h_u_cla32_and6888_y0, h_u_cla32_and6887_y0, h_u_cla32_and6889_y0);
  and_gate and_gate_h_u_cla32_and6890_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6890_y0);
  and_gate and_gate_h_u_cla32_and6891_y0(h_u_cla32_and6890_y0, h_u_cla32_and6889_y0, h_u_cla32_and6891_y0);
  and_gate and_gate_h_u_cla32_and6892_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and6892_y0);
  and_gate and_gate_h_u_cla32_and6893_y0(h_u_cla32_and6892_y0, h_u_cla32_and6891_y0, h_u_cla32_and6893_y0);
  and_gate and_gate_h_u_cla32_and6894_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6894_y0);
  and_gate and_gate_h_u_cla32_and6895_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6895_y0);
  and_gate and_gate_h_u_cla32_and6896_y0(h_u_cla32_and6895_y0, h_u_cla32_and6894_y0, h_u_cla32_and6896_y0);
  and_gate and_gate_h_u_cla32_and6897_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6897_y0);
  and_gate and_gate_h_u_cla32_and6898_y0(h_u_cla32_and6897_y0, h_u_cla32_and6896_y0, h_u_cla32_and6898_y0);
  and_gate and_gate_h_u_cla32_and6899_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6899_y0);
  and_gate and_gate_h_u_cla32_and6900_y0(h_u_cla32_and6899_y0, h_u_cla32_and6898_y0, h_u_cla32_and6900_y0);
  and_gate and_gate_h_u_cla32_and6901_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6901_y0);
  and_gate and_gate_h_u_cla32_and6902_y0(h_u_cla32_and6901_y0, h_u_cla32_and6900_y0, h_u_cla32_and6902_y0);
  and_gate and_gate_h_u_cla32_and6903_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and6903_y0);
  and_gate and_gate_h_u_cla32_and6904_y0(h_u_cla32_and6903_y0, h_u_cla32_and6902_y0, h_u_cla32_and6904_y0);
  and_gate and_gate_h_u_cla32_and6905_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6905_y0);
  and_gate and_gate_h_u_cla32_and6906_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6906_y0);
  and_gate and_gate_h_u_cla32_and6907_y0(h_u_cla32_and6906_y0, h_u_cla32_and6905_y0, h_u_cla32_and6907_y0);
  and_gate and_gate_h_u_cla32_and6908_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6908_y0);
  and_gate and_gate_h_u_cla32_and6909_y0(h_u_cla32_and6908_y0, h_u_cla32_and6907_y0, h_u_cla32_and6909_y0);
  and_gate and_gate_h_u_cla32_and6910_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6910_y0);
  and_gate and_gate_h_u_cla32_and6911_y0(h_u_cla32_and6910_y0, h_u_cla32_and6909_y0, h_u_cla32_and6911_y0);
  and_gate and_gate_h_u_cla32_and6912_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and6912_y0);
  and_gate and_gate_h_u_cla32_and6913_y0(h_u_cla32_and6912_y0, h_u_cla32_and6911_y0, h_u_cla32_and6913_y0);
  and_gate and_gate_h_u_cla32_and6914_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6914_y0);
  and_gate and_gate_h_u_cla32_and6915_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6915_y0);
  and_gate and_gate_h_u_cla32_and6916_y0(h_u_cla32_and6915_y0, h_u_cla32_and6914_y0, h_u_cla32_and6916_y0);
  and_gate and_gate_h_u_cla32_and6917_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6917_y0);
  and_gate and_gate_h_u_cla32_and6918_y0(h_u_cla32_and6917_y0, h_u_cla32_and6916_y0, h_u_cla32_and6918_y0);
  and_gate and_gate_h_u_cla32_and6919_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and6919_y0);
  and_gate and_gate_h_u_cla32_and6920_y0(h_u_cla32_and6919_y0, h_u_cla32_and6918_y0, h_u_cla32_and6920_y0);
  and_gate and_gate_h_u_cla32_and6921_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and6921_y0);
  and_gate and_gate_h_u_cla32_and6922_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and6922_y0);
  and_gate and_gate_h_u_cla32_and6923_y0(h_u_cla32_and6922_y0, h_u_cla32_and6921_y0, h_u_cla32_and6923_y0);
  and_gate and_gate_h_u_cla32_and6924_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and6924_y0);
  and_gate and_gate_h_u_cla32_and6925_y0(h_u_cla32_and6924_y0, h_u_cla32_and6923_y0, h_u_cla32_and6925_y0);
  and_gate and_gate_h_u_cla32_and6926_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and6926_y0);
  and_gate and_gate_h_u_cla32_and6927_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and6927_y0);
  and_gate and_gate_h_u_cla32_and6928_y0(h_u_cla32_and6927_y0, h_u_cla32_and6926_y0, h_u_cla32_and6928_y0);
  and_gate and_gate_h_u_cla32_and6929_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and6929_y0);
  or_gate or_gate_h_u_cla32_or351_y0(h_u_cla32_and6929_y0, h_u_cla32_and6253_y0, h_u_cla32_or351_y0);
  or_gate or_gate_h_u_cla32_or352_y0(h_u_cla32_or351_y0, h_u_cla32_and6304_y0, h_u_cla32_or352_y0);
  or_gate or_gate_h_u_cla32_or353_y0(h_u_cla32_or352_y0, h_u_cla32_and6353_y0, h_u_cla32_or353_y0);
  or_gate or_gate_h_u_cla32_or354_y0(h_u_cla32_or353_y0, h_u_cla32_and6400_y0, h_u_cla32_or354_y0);
  or_gate or_gate_h_u_cla32_or355_y0(h_u_cla32_or354_y0, h_u_cla32_and6445_y0, h_u_cla32_or355_y0);
  or_gate or_gate_h_u_cla32_or356_y0(h_u_cla32_or355_y0, h_u_cla32_and6488_y0, h_u_cla32_or356_y0);
  or_gate or_gate_h_u_cla32_or357_y0(h_u_cla32_or356_y0, h_u_cla32_and6529_y0, h_u_cla32_or357_y0);
  or_gate or_gate_h_u_cla32_or358_y0(h_u_cla32_or357_y0, h_u_cla32_and6568_y0, h_u_cla32_or358_y0);
  or_gate or_gate_h_u_cla32_or359_y0(h_u_cla32_or358_y0, h_u_cla32_and6605_y0, h_u_cla32_or359_y0);
  or_gate or_gate_h_u_cla32_or360_y0(h_u_cla32_or359_y0, h_u_cla32_and6640_y0, h_u_cla32_or360_y0);
  or_gate or_gate_h_u_cla32_or361_y0(h_u_cla32_or360_y0, h_u_cla32_and6673_y0, h_u_cla32_or361_y0);
  or_gate or_gate_h_u_cla32_or362_y0(h_u_cla32_or361_y0, h_u_cla32_and6704_y0, h_u_cla32_or362_y0);
  or_gate or_gate_h_u_cla32_or363_y0(h_u_cla32_or362_y0, h_u_cla32_and6733_y0, h_u_cla32_or363_y0);
  or_gate or_gate_h_u_cla32_or364_y0(h_u_cla32_or363_y0, h_u_cla32_and6760_y0, h_u_cla32_or364_y0);
  or_gate or_gate_h_u_cla32_or365_y0(h_u_cla32_or364_y0, h_u_cla32_and6785_y0, h_u_cla32_or365_y0);
  or_gate or_gate_h_u_cla32_or366_y0(h_u_cla32_or365_y0, h_u_cla32_and6808_y0, h_u_cla32_or366_y0);
  or_gate or_gate_h_u_cla32_or367_y0(h_u_cla32_or366_y0, h_u_cla32_and6829_y0, h_u_cla32_or367_y0);
  or_gate or_gate_h_u_cla32_or368_y0(h_u_cla32_or367_y0, h_u_cla32_and6848_y0, h_u_cla32_or368_y0);
  or_gate or_gate_h_u_cla32_or369_y0(h_u_cla32_or368_y0, h_u_cla32_and6865_y0, h_u_cla32_or369_y0);
  or_gate or_gate_h_u_cla32_or370_y0(h_u_cla32_or369_y0, h_u_cla32_and6880_y0, h_u_cla32_or370_y0);
  or_gate or_gate_h_u_cla32_or371_y0(h_u_cla32_or370_y0, h_u_cla32_and6893_y0, h_u_cla32_or371_y0);
  or_gate or_gate_h_u_cla32_or372_y0(h_u_cla32_or371_y0, h_u_cla32_and6904_y0, h_u_cla32_or372_y0);
  or_gate or_gate_h_u_cla32_or373_y0(h_u_cla32_or372_y0, h_u_cla32_and6913_y0, h_u_cla32_or373_y0);
  or_gate or_gate_h_u_cla32_or374_y0(h_u_cla32_or373_y0, h_u_cla32_and6920_y0, h_u_cla32_or374_y0);
  or_gate or_gate_h_u_cla32_or375_y0(h_u_cla32_or374_y0, h_u_cla32_and6925_y0, h_u_cla32_or375_y0);
  or_gate or_gate_h_u_cla32_or376_y0(h_u_cla32_or375_y0, h_u_cla32_and6928_y0, h_u_cla32_or376_y0);
  or_gate or_gate_h_u_cla32_or377_y0(h_u_cla32_pg_logic26_y1, h_u_cla32_or376_y0, h_u_cla32_or377_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic27_y0(a_27, b_27, h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_pg_logic27_y2);
  xor_gate xor_gate_h_u_cla32_xor27_y0(h_u_cla32_pg_logic27_y2, h_u_cla32_or377_y0, h_u_cla32_xor27_y0);
  and_gate and_gate_h_u_cla32_and6930_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and6930_y0);
  and_gate and_gate_h_u_cla32_and6931_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and6931_y0);
  and_gate and_gate_h_u_cla32_and6932_y0(h_u_cla32_and6931_y0, h_u_cla32_and6930_y0, h_u_cla32_and6932_y0);
  and_gate and_gate_h_u_cla32_and6933_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and6933_y0);
  and_gate and_gate_h_u_cla32_and6934_y0(h_u_cla32_and6933_y0, h_u_cla32_and6932_y0, h_u_cla32_and6934_y0);
  and_gate and_gate_h_u_cla32_and6935_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and6935_y0);
  and_gate and_gate_h_u_cla32_and6936_y0(h_u_cla32_and6935_y0, h_u_cla32_and6934_y0, h_u_cla32_and6936_y0);
  and_gate and_gate_h_u_cla32_and6937_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and6937_y0);
  and_gate and_gate_h_u_cla32_and6938_y0(h_u_cla32_and6937_y0, h_u_cla32_and6936_y0, h_u_cla32_and6938_y0);
  and_gate and_gate_h_u_cla32_and6939_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and6939_y0);
  and_gate and_gate_h_u_cla32_and6940_y0(h_u_cla32_and6939_y0, h_u_cla32_and6938_y0, h_u_cla32_and6940_y0);
  and_gate and_gate_h_u_cla32_and6941_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and6941_y0);
  and_gate and_gate_h_u_cla32_and6942_y0(h_u_cla32_and6941_y0, h_u_cla32_and6940_y0, h_u_cla32_and6942_y0);
  and_gate and_gate_h_u_cla32_and6943_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and6943_y0);
  and_gate and_gate_h_u_cla32_and6944_y0(h_u_cla32_and6943_y0, h_u_cla32_and6942_y0, h_u_cla32_and6944_y0);
  and_gate and_gate_h_u_cla32_and6945_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and6945_y0);
  and_gate and_gate_h_u_cla32_and6946_y0(h_u_cla32_and6945_y0, h_u_cla32_and6944_y0, h_u_cla32_and6946_y0);
  and_gate and_gate_h_u_cla32_and6947_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and6947_y0);
  and_gate and_gate_h_u_cla32_and6948_y0(h_u_cla32_and6947_y0, h_u_cla32_and6946_y0, h_u_cla32_and6948_y0);
  and_gate and_gate_h_u_cla32_and6949_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and6949_y0);
  and_gate and_gate_h_u_cla32_and6950_y0(h_u_cla32_and6949_y0, h_u_cla32_and6948_y0, h_u_cla32_and6950_y0);
  and_gate and_gate_h_u_cla32_and6951_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and6951_y0);
  and_gate and_gate_h_u_cla32_and6952_y0(h_u_cla32_and6951_y0, h_u_cla32_and6950_y0, h_u_cla32_and6952_y0);
  and_gate and_gate_h_u_cla32_and6953_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and6953_y0);
  and_gate and_gate_h_u_cla32_and6954_y0(h_u_cla32_and6953_y0, h_u_cla32_and6952_y0, h_u_cla32_and6954_y0);
  and_gate and_gate_h_u_cla32_and6955_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and6955_y0);
  and_gate and_gate_h_u_cla32_and6956_y0(h_u_cla32_and6955_y0, h_u_cla32_and6954_y0, h_u_cla32_and6956_y0);
  and_gate and_gate_h_u_cla32_and6957_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and6957_y0);
  and_gate and_gate_h_u_cla32_and6958_y0(h_u_cla32_and6957_y0, h_u_cla32_and6956_y0, h_u_cla32_and6958_y0);
  and_gate and_gate_h_u_cla32_and6959_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and6959_y0);
  and_gate and_gate_h_u_cla32_and6960_y0(h_u_cla32_and6959_y0, h_u_cla32_and6958_y0, h_u_cla32_and6960_y0);
  and_gate and_gate_h_u_cla32_and6961_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and6961_y0);
  and_gate and_gate_h_u_cla32_and6962_y0(h_u_cla32_and6961_y0, h_u_cla32_and6960_y0, h_u_cla32_and6962_y0);
  and_gate and_gate_h_u_cla32_and6963_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and6963_y0);
  and_gate and_gate_h_u_cla32_and6964_y0(h_u_cla32_and6963_y0, h_u_cla32_and6962_y0, h_u_cla32_and6964_y0);
  and_gate and_gate_h_u_cla32_and6965_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and6965_y0);
  and_gate and_gate_h_u_cla32_and6966_y0(h_u_cla32_and6965_y0, h_u_cla32_and6964_y0, h_u_cla32_and6966_y0);
  and_gate and_gate_h_u_cla32_and6967_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and6967_y0);
  and_gate and_gate_h_u_cla32_and6968_y0(h_u_cla32_and6967_y0, h_u_cla32_and6966_y0, h_u_cla32_and6968_y0);
  and_gate and_gate_h_u_cla32_and6969_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and6969_y0);
  and_gate and_gate_h_u_cla32_and6970_y0(h_u_cla32_and6969_y0, h_u_cla32_and6968_y0, h_u_cla32_and6970_y0);
  and_gate and_gate_h_u_cla32_and6971_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and6971_y0);
  and_gate and_gate_h_u_cla32_and6972_y0(h_u_cla32_and6971_y0, h_u_cla32_and6970_y0, h_u_cla32_and6972_y0);
  and_gate and_gate_h_u_cla32_and6973_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and6973_y0);
  and_gate and_gate_h_u_cla32_and6974_y0(h_u_cla32_and6973_y0, h_u_cla32_and6972_y0, h_u_cla32_and6974_y0);
  and_gate and_gate_h_u_cla32_and6975_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and6975_y0);
  and_gate and_gate_h_u_cla32_and6976_y0(h_u_cla32_and6975_y0, h_u_cla32_and6974_y0, h_u_cla32_and6976_y0);
  and_gate and_gate_h_u_cla32_and6977_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and6977_y0);
  and_gate and_gate_h_u_cla32_and6978_y0(h_u_cla32_and6977_y0, h_u_cla32_and6976_y0, h_u_cla32_and6978_y0);
  and_gate and_gate_h_u_cla32_and6979_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and6979_y0);
  and_gate and_gate_h_u_cla32_and6980_y0(h_u_cla32_and6979_y0, h_u_cla32_and6978_y0, h_u_cla32_and6980_y0);
  and_gate and_gate_h_u_cla32_and6981_y0(h_u_cla32_pg_logic26_y0, constant_wire_0, h_u_cla32_and6981_y0);
  and_gate and_gate_h_u_cla32_and6982_y0(h_u_cla32_and6981_y0, h_u_cla32_and6980_y0, h_u_cla32_and6982_y0);
  and_gate and_gate_h_u_cla32_and6983_y0(h_u_cla32_pg_logic27_y0, constant_wire_0, h_u_cla32_and6983_y0);
  and_gate and_gate_h_u_cla32_and6984_y0(h_u_cla32_and6983_y0, h_u_cla32_and6982_y0, h_u_cla32_and6984_y0);
  and_gate and_gate_h_u_cla32_and6985_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6985_y0);
  and_gate and_gate_h_u_cla32_and6986_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6986_y0);
  and_gate and_gate_h_u_cla32_and6987_y0(h_u_cla32_and6986_y0, h_u_cla32_and6985_y0, h_u_cla32_and6987_y0);
  and_gate and_gate_h_u_cla32_and6988_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6988_y0);
  and_gate and_gate_h_u_cla32_and6989_y0(h_u_cla32_and6988_y0, h_u_cla32_and6987_y0, h_u_cla32_and6989_y0);
  and_gate and_gate_h_u_cla32_and6990_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6990_y0);
  and_gate and_gate_h_u_cla32_and6991_y0(h_u_cla32_and6990_y0, h_u_cla32_and6989_y0, h_u_cla32_and6991_y0);
  and_gate and_gate_h_u_cla32_and6992_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6992_y0);
  and_gate and_gate_h_u_cla32_and6993_y0(h_u_cla32_and6992_y0, h_u_cla32_and6991_y0, h_u_cla32_and6993_y0);
  and_gate and_gate_h_u_cla32_and6994_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6994_y0);
  and_gate and_gate_h_u_cla32_and6995_y0(h_u_cla32_and6994_y0, h_u_cla32_and6993_y0, h_u_cla32_and6995_y0);
  and_gate and_gate_h_u_cla32_and6996_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6996_y0);
  and_gate and_gate_h_u_cla32_and6997_y0(h_u_cla32_and6996_y0, h_u_cla32_and6995_y0, h_u_cla32_and6997_y0);
  and_gate and_gate_h_u_cla32_and6998_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and6998_y0);
  and_gate and_gate_h_u_cla32_and6999_y0(h_u_cla32_and6998_y0, h_u_cla32_and6997_y0, h_u_cla32_and6999_y0);
  and_gate and_gate_h_u_cla32_and7000_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7000_y0);
  and_gate and_gate_h_u_cla32_and7001_y0(h_u_cla32_and7000_y0, h_u_cla32_and6999_y0, h_u_cla32_and7001_y0);
  and_gate and_gate_h_u_cla32_and7002_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7002_y0);
  and_gate and_gate_h_u_cla32_and7003_y0(h_u_cla32_and7002_y0, h_u_cla32_and7001_y0, h_u_cla32_and7003_y0);
  and_gate and_gate_h_u_cla32_and7004_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7004_y0);
  and_gate and_gate_h_u_cla32_and7005_y0(h_u_cla32_and7004_y0, h_u_cla32_and7003_y0, h_u_cla32_and7005_y0);
  and_gate and_gate_h_u_cla32_and7006_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7006_y0);
  and_gate and_gate_h_u_cla32_and7007_y0(h_u_cla32_and7006_y0, h_u_cla32_and7005_y0, h_u_cla32_and7007_y0);
  and_gate and_gate_h_u_cla32_and7008_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7008_y0);
  and_gate and_gate_h_u_cla32_and7009_y0(h_u_cla32_and7008_y0, h_u_cla32_and7007_y0, h_u_cla32_and7009_y0);
  and_gate and_gate_h_u_cla32_and7010_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7010_y0);
  and_gate and_gate_h_u_cla32_and7011_y0(h_u_cla32_and7010_y0, h_u_cla32_and7009_y0, h_u_cla32_and7011_y0);
  and_gate and_gate_h_u_cla32_and7012_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7012_y0);
  and_gate and_gate_h_u_cla32_and7013_y0(h_u_cla32_and7012_y0, h_u_cla32_and7011_y0, h_u_cla32_and7013_y0);
  and_gate and_gate_h_u_cla32_and7014_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7014_y0);
  and_gate and_gate_h_u_cla32_and7015_y0(h_u_cla32_and7014_y0, h_u_cla32_and7013_y0, h_u_cla32_and7015_y0);
  and_gate and_gate_h_u_cla32_and7016_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7016_y0);
  and_gate and_gate_h_u_cla32_and7017_y0(h_u_cla32_and7016_y0, h_u_cla32_and7015_y0, h_u_cla32_and7017_y0);
  and_gate and_gate_h_u_cla32_and7018_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7018_y0);
  and_gate and_gate_h_u_cla32_and7019_y0(h_u_cla32_and7018_y0, h_u_cla32_and7017_y0, h_u_cla32_and7019_y0);
  and_gate and_gate_h_u_cla32_and7020_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7020_y0);
  and_gate and_gate_h_u_cla32_and7021_y0(h_u_cla32_and7020_y0, h_u_cla32_and7019_y0, h_u_cla32_and7021_y0);
  and_gate and_gate_h_u_cla32_and7022_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7022_y0);
  and_gate and_gate_h_u_cla32_and7023_y0(h_u_cla32_and7022_y0, h_u_cla32_and7021_y0, h_u_cla32_and7023_y0);
  and_gate and_gate_h_u_cla32_and7024_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7024_y0);
  and_gate and_gate_h_u_cla32_and7025_y0(h_u_cla32_and7024_y0, h_u_cla32_and7023_y0, h_u_cla32_and7025_y0);
  and_gate and_gate_h_u_cla32_and7026_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7026_y0);
  and_gate and_gate_h_u_cla32_and7027_y0(h_u_cla32_and7026_y0, h_u_cla32_and7025_y0, h_u_cla32_and7027_y0);
  and_gate and_gate_h_u_cla32_and7028_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7028_y0);
  and_gate and_gate_h_u_cla32_and7029_y0(h_u_cla32_and7028_y0, h_u_cla32_and7027_y0, h_u_cla32_and7029_y0);
  and_gate and_gate_h_u_cla32_and7030_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7030_y0);
  and_gate and_gate_h_u_cla32_and7031_y0(h_u_cla32_and7030_y0, h_u_cla32_and7029_y0, h_u_cla32_and7031_y0);
  and_gate and_gate_h_u_cla32_and7032_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7032_y0);
  and_gate and_gate_h_u_cla32_and7033_y0(h_u_cla32_and7032_y0, h_u_cla32_and7031_y0, h_u_cla32_and7033_y0);
  and_gate and_gate_h_u_cla32_and7034_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7034_y0);
  and_gate and_gate_h_u_cla32_and7035_y0(h_u_cla32_and7034_y0, h_u_cla32_and7033_y0, h_u_cla32_and7035_y0);
  and_gate and_gate_h_u_cla32_and7036_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7036_y0);
  and_gate and_gate_h_u_cla32_and7037_y0(h_u_cla32_and7036_y0, h_u_cla32_and7035_y0, h_u_cla32_and7037_y0);
  and_gate and_gate_h_u_cla32_and7038_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7038_y0);
  and_gate and_gate_h_u_cla32_and7039_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7039_y0);
  and_gate and_gate_h_u_cla32_and7040_y0(h_u_cla32_and7039_y0, h_u_cla32_and7038_y0, h_u_cla32_and7040_y0);
  and_gate and_gate_h_u_cla32_and7041_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7041_y0);
  and_gate and_gate_h_u_cla32_and7042_y0(h_u_cla32_and7041_y0, h_u_cla32_and7040_y0, h_u_cla32_and7042_y0);
  and_gate and_gate_h_u_cla32_and7043_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7043_y0);
  and_gate and_gate_h_u_cla32_and7044_y0(h_u_cla32_and7043_y0, h_u_cla32_and7042_y0, h_u_cla32_and7044_y0);
  and_gate and_gate_h_u_cla32_and7045_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7045_y0);
  and_gate and_gate_h_u_cla32_and7046_y0(h_u_cla32_and7045_y0, h_u_cla32_and7044_y0, h_u_cla32_and7046_y0);
  and_gate and_gate_h_u_cla32_and7047_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7047_y0);
  and_gate and_gate_h_u_cla32_and7048_y0(h_u_cla32_and7047_y0, h_u_cla32_and7046_y0, h_u_cla32_and7048_y0);
  and_gate and_gate_h_u_cla32_and7049_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7049_y0);
  and_gate and_gate_h_u_cla32_and7050_y0(h_u_cla32_and7049_y0, h_u_cla32_and7048_y0, h_u_cla32_and7050_y0);
  and_gate and_gate_h_u_cla32_and7051_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7051_y0);
  and_gate and_gate_h_u_cla32_and7052_y0(h_u_cla32_and7051_y0, h_u_cla32_and7050_y0, h_u_cla32_and7052_y0);
  and_gate and_gate_h_u_cla32_and7053_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7053_y0);
  and_gate and_gate_h_u_cla32_and7054_y0(h_u_cla32_and7053_y0, h_u_cla32_and7052_y0, h_u_cla32_and7054_y0);
  and_gate and_gate_h_u_cla32_and7055_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7055_y0);
  and_gate and_gate_h_u_cla32_and7056_y0(h_u_cla32_and7055_y0, h_u_cla32_and7054_y0, h_u_cla32_and7056_y0);
  and_gate and_gate_h_u_cla32_and7057_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7057_y0);
  and_gate and_gate_h_u_cla32_and7058_y0(h_u_cla32_and7057_y0, h_u_cla32_and7056_y0, h_u_cla32_and7058_y0);
  and_gate and_gate_h_u_cla32_and7059_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7059_y0);
  and_gate and_gate_h_u_cla32_and7060_y0(h_u_cla32_and7059_y0, h_u_cla32_and7058_y0, h_u_cla32_and7060_y0);
  and_gate and_gate_h_u_cla32_and7061_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7061_y0);
  and_gate and_gate_h_u_cla32_and7062_y0(h_u_cla32_and7061_y0, h_u_cla32_and7060_y0, h_u_cla32_and7062_y0);
  and_gate and_gate_h_u_cla32_and7063_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7063_y0);
  and_gate and_gate_h_u_cla32_and7064_y0(h_u_cla32_and7063_y0, h_u_cla32_and7062_y0, h_u_cla32_and7064_y0);
  and_gate and_gate_h_u_cla32_and7065_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7065_y0);
  and_gate and_gate_h_u_cla32_and7066_y0(h_u_cla32_and7065_y0, h_u_cla32_and7064_y0, h_u_cla32_and7066_y0);
  and_gate and_gate_h_u_cla32_and7067_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7067_y0);
  and_gate and_gate_h_u_cla32_and7068_y0(h_u_cla32_and7067_y0, h_u_cla32_and7066_y0, h_u_cla32_and7068_y0);
  and_gate and_gate_h_u_cla32_and7069_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7069_y0);
  and_gate and_gate_h_u_cla32_and7070_y0(h_u_cla32_and7069_y0, h_u_cla32_and7068_y0, h_u_cla32_and7070_y0);
  and_gate and_gate_h_u_cla32_and7071_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7071_y0);
  and_gate and_gate_h_u_cla32_and7072_y0(h_u_cla32_and7071_y0, h_u_cla32_and7070_y0, h_u_cla32_and7072_y0);
  and_gate and_gate_h_u_cla32_and7073_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7073_y0);
  and_gate and_gate_h_u_cla32_and7074_y0(h_u_cla32_and7073_y0, h_u_cla32_and7072_y0, h_u_cla32_and7074_y0);
  and_gate and_gate_h_u_cla32_and7075_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7075_y0);
  and_gate and_gate_h_u_cla32_and7076_y0(h_u_cla32_and7075_y0, h_u_cla32_and7074_y0, h_u_cla32_and7076_y0);
  and_gate and_gate_h_u_cla32_and7077_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7077_y0);
  and_gate and_gate_h_u_cla32_and7078_y0(h_u_cla32_and7077_y0, h_u_cla32_and7076_y0, h_u_cla32_and7078_y0);
  and_gate and_gate_h_u_cla32_and7079_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7079_y0);
  and_gate and_gate_h_u_cla32_and7080_y0(h_u_cla32_and7079_y0, h_u_cla32_and7078_y0, h_u_cla32_and7080_y0);
  and_gate and_gate_h_u_cla32_and7081_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7081_y0);
  and_gate and_gate_h_u_cla32_and7082_y0(h_u_cla32_and7081_y0, h_u_cla32_and7080_y0, h_u_cla32_and7082_y0);
  and_gate and_gate_h_u_cla32_and7083_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7083_y0);
  and_gate and_gate_h_u_cla32_and7084_y0(h_u_cla32_and7083_y0, h_u_cla32_and7082_y0, h_u_cla32_and7084_y0);
  and_gate and_gate_h_u_cla32_and7085_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7085_y0);
  and_gate and_gate_h_u_cla32_and7086_y0(h_u_cla32_and7085_y0, h_u_cla32_and7084_y0, h_u_cla32_and7086_y0);
  and_gate and_gate_h_u_cla32_and7087_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7087_y0);
  and_gate and_gate_h_u_cla32_and7088_y0(h_u_cla32_and7087_y0, h_u_cla32_and7086_y0, h_u_cla32_and7088_y0);
  and_gate and_gate_h_u_cla32_and7089_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7089_y0);
  and_gate and_gate_h_u_cla32_and7090_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7090_y0);
  and_gate and_gate_h_u_cla32_and7091_y0(h_u_cla32_and7090_y0, h_u_cla32_and7089_y0, h_u_cla32_and7091_y0);
  and_gate and_gate_h_u_cla32_and7092_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7092_y0);
  and_gate and_gate_h_u_cla32_and7093_y0(h_u_cla32_and7092_y0, h_u_cla32_and7091_y0, h_u_cla32_and7093_y0);
  and_gate and_gate_h_u_cla32_and7094_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7094_y0);
  and_gate and_gate_h_u_cla32_and7095_y0(h_u_cla32_and7094_y0, h_u_cla32_and7093_y0, h_u_cla32_and7095_y0);
  and_gate and_gate_h_u_cla32_and7096_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7096_y0);
  and_gate and_gate_h_u_cla32_and7097_y0(h_u_cla32_and7096_y0, h_u_cla32_and7095_y0, h_u_cla32_and7097_y0);
  and_gate and_gate_h_u_cla32_and7098_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7098_y0);
  and_gate and_gate_h_u_cla32_and7099_y0(h_u_cla32_and7098_y0, h_u_cla32_and7097_y0, h_u_cla32_and7099_y0);
  and_gate and_gate_h_u_cla32_and7100_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7100_y0);
  and_gate and_gate_h_u_cla32_and7101_y0(h_u_cla32_and7100_y0, h_u_cla32_and7099_y0, h_u_cla32_and7101_y0);
  and_gate and_gate_h_u_cla32_and7102_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7102_y0);
  and_gate and_gate_h_u_cla32_and7103_y0(h_u_cla32_and7102_y0, h_u_cla32_and7101_y0, h_u_cla32_and7103_y0);
  and_gate and_gate_h_u_cla32_and7104_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7104_y0);
  and_gate and_gate_h_u_cla32_and7105_y0(h_u_cla32_and7104_y0, h_u_cla32_and7103_y0, h_u_cla32_and7105_y0);
  and_gate and_gate_h_u_cla32_and7106_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7106_y0);
  and_gate and_gate_h_u_cla32_and7107_y0(h_u_cla32_and7106_y0, h_u_cla32_and7105_y0, h_u_cla32_and7107_y0);
  and_gate and_gate_h_u_cla32_and7108_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7108_y0);
  and_gate and_gate_h_u_cla32_and7109_y0(h_u_cla32_and7108_y0, h_u_cla32_and7107_y0, h_u_cla32_and7109_y0);
  and_gate and_gate_h_u_cla32_and7110_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7110_y0);
  and_gate and_gate_h_u_cla32_and7111_y0(h_u_cla32_and7110_y0, h_u_cla32_and7109_y0, h_u_cla32_and7111_y0);
  and_gate and_gate_h_u_cla32_and7112_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7112_y0);
  and_gate and_gate_h_u_cla32_and7113_y0(h_u_cla32_and7112_y0, h_u_cla32_and7111_y0, h_u_cla32_and7113_y0);
  and_gate and_gate_h_u_cla32_and7114_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7114_y0);
  and_gate and_gate_h_u_cla32_and7115_y0(h_u_cla32_and7114_y0, h_u_cla32_and7113_y0, h_u_cla32_and7115_y0);
  and_gate and_gate_h_u_cla32_and7116_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7116_y0);
  and_gate and_gate_h_u_cla32_and7117_y0(h_u_cla32_and7116_y0, h_u_cla32_and7115_y0, h_u_cla32_and7117_y0);
  and_gate and_gate_h_u_cla32_and7118_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7118_y0);
  and_gate and_gate_h_u_cla32_and7119_y0(h_u_cla32_and7118_y0, h_u_cla32_and7117_y0, h_u_cla32_and7119_y0);
  and_gate and_gate_h_u_cla32_and7120_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7120_y0);
  and_gate and_gate_h_u_cla32_and7121_y0(h_u_cla32_and7120_y0, h_u_cla32_and7119_y0, h_u_cla32_and7121_y0);
  and_gate and_gate_h_u_cla32_and7122_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7122_y0);
  and_gate and_gate_h_u_cla32_and7123_y0(h_u_cla32_and7122_y0, h_u_cla32_and7121_y0, h_u_cla32_and7123_y0);
  and_gate and_gate_h_u_cla32_and7124_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7124_y0);
  and_gate and_gate_h_u_cla32_and7125_y0(h_u_cla32_and7124_y0, h_u_cla32_and7123_y0, h_u_cla32_and7125_y0);
  and_gate and_gate_h_u_cla32_and7126_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7126_y0);
  and_gate and_gate_h_u_cla32_and7127_y0(h_u_cla32_and7126_y0, h_u_cla32_and7125_y0, h_u_cla32_and7127_y0);
  and_gate and_gate_h_u_cla32_and7128_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7128_y0);
  and_gate and_gate_h_u_cla32_and7129_y0(h_u_cla32_and7128_y0, h_u_cla32_and7127_y0, h_u_cla32_and7129_y0);
  and_gate and_gate_h_u_cla32_and7130_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7130_y0);
  and_gate and_gate_h_u_cla32_and7131_y0(h_u_cla32_and7130_y0, h_u_cla32_and7129_y0, h_u_cla32_and7131_y0);
  and_gate and_gate_h_u_cla32_and7132_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7132_y0);
  and_gate and_gate_h_u_cla32_and7133_y0(h_u_cla32_and7132_y0, h_u_cla32_and7131_y0, h_u_cla32_and7133_y0);
  and_gate and_gate_h_u_cla32_and7134_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7134_y0);
  and_gate and_gate_h_u_cla32_and7135_y0(h_u_cla32_and7134_y0, h_u_cla32_and7133_y0, h_u_cla32_and7135_y0);
  and_gate and_gate_h_u_cla32_and7136_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7136_y0);
  and_gate and_gate_h_u_cla32_and7137_y0(h_u_cla32_and7136_y0, h_u_cla32_and7135_y0, h_u_cla32_and7137_y0);
  and_gate and_gate_h_u_cla32_and7138_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7138_y0);
  and_gate and_gate_h_u_cla32_and7139_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7139_y0);
  and_gate and_gate_h_u_cla32_and7140_y0(h_u_cla32_and7139_y0, h_u_cla32_and7138_y0, h_u_cla32_and7140_y0);
  and_gate and_gate_h_u_cla32_and7141_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7141_y0);
  and_gate and_gate_h_u_cla32_and7142_y0(h_u_cla32_and7141_y0, h_u_cla32_and7140_y0, h_u_cla32_and7142_y0);
  and_gate and_gate_h_u_cla32_and7143_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7143_y0);
  and_gate and_gate_h_u_cla32_and7144_y0(h_u_cla32_and7143_y0, h_u_cla32_and7142_y0, h_u_cla32_and7144_y0);
  and_gate and_gate_h_u_cla32_and7145_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7145_y0);
  and_gate and_gate_h_u_cla32_and7146_y0(h_u_cla32_and7145_y0, h_u_cla32_and7144_y0, h_u_cla32_and7146_y0);
  and_gate and_gate_h_u_cla32_and7147_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7147_y0);
  and_gate and_gate_h_u_cla32_and7148_y0(h_u_cla32_and7147_y0, h_u_cla32_and7146_y0, h_u_cla32_and7148_y0);
  and_gate and_gate_h_u_cla32_and7149_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7149_y0);
  and_gate and_gate_h_u_cla32_and7150_y0(h_u_cla32_and7149_y0, h_u_cla32_and7148_y0, h_u_cla32_and7150_y0);
  and_gate and_gate_h_u_cla32_and7151_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7151_y0);
  and_gate and_gate_h_u_cla32_and7152_y0(h_u_cla32_and7151_y0, h_u_cla32_and7150_y0, h_u_cla32_and7152_y0);
  and_gate and_gate_h_u_cla32_and7153_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7153_y0);
  and_gate and_gate_h_u_cla32_and7154_y0(h_u_cla32_and7153_y0, h_u_cla32_and7152_y0, h_u_cla32_and7154_y0);
  and_gate and_gate_h_u_cla32_and7155_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7155_y0);
  and_gate and_gate_h_u_cla32_and7156_y0(h_u_cla32_and7155_y0, h_u_cla32_and7154_y0, h_u_cla32_and7156_y0);
  and_gate and_gate_h_u_cla32_and7157_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7157_y0);
  and_gate and_gate_h_u_cla32_and7158_y0(h_u_cla32_and7157_y0, h_u_cla32_and7156_y0, h_u_cla32_and7158_y0);
  and_gate and_gate_h_u_cla32_and7159_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7159_y0);
  and_gate and_gate_h_u_cla32_and7160_y0(h_u_cla32_and7159_y0, h_u_cla32_and7158_y0, h_u_cla32_and7160_y0);
  and_gate and_gate_h_u_cla32_and7161_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7161_y0);
  and_gate and_gate_h_u_cla32_and7162_y0(h_u_cla32_and7161_y0, h_u_cla32_and7160_y0, h_u_cla32_and7162_y0);
  and_gate and_gate_h_u_cla32_and7163_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7163_y0);
  and_gate and_gate_h_u_cla32_and7164_y0(h_u_cla32_and7163_y0, h_u_cla32_and7162_y0, h_u_cla32_and7164_y0);
  and_gate and_gate_h_u_cla32_and7165_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7165_y0);
  and_gate and_gate_h_u_cla32_and7166_y0(h_u_cla32_and7165_y0, h_u_cla32_and7164_y0, h_u_cla32_and7166_y0);
  and_gate and_gate_h_u_cla32_and7167_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7167_y0);
  and_gate and_gate_h_u_cla32_and7168_y0(h_u_cla32_and7167_y0, h_u_cla32_and7166_y0, h_u_cla32_and7168_y0);
  and_gate and_gate_h_u_cla32_and7169_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7169_y0);
  and_gate and_gate_h_u_cla32_and7170_y0(h_u_cla32_and7169_y0, h_u_cla32_and7168_y0, h_u_cla32_and7170_y0);
  and_gate and_gate_h_u_cla32_and7171_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7171_y0);
  and_gate and_gate_h_u_cla32_and7172_y0(h_u_cla32_and7171_y0, h_u_cla32_and7170_y0, h_u_cla32_and7172_y0);
  and_gate and_gate_h_u_cla32_and7173_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7173_y0);
  and_gate and_gate_h_u_cla32_and7174_y0(h_u_cla32_and7173_y0, h_u_cla32_and7172_y0, h_u_cla32_and7174_y0);
  and_gate and_gate_h_u_cla32_and7175_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7175_y0);
  and_gate and_gate_h_u_cla32_and7176_y0(h_u_cla32_and7175_y0, h_u_cla32_and7174_y0, h_u_cla32_and7176_y0);
  and_gate and_gate_h_u_cla32_and7177_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7177_y0);
  and_gate and_gate_h_u_cla32_and7178_y0(h_u_cla32_and7177_y0, h_u_cla32_and7176_y0, h_u_cla32_and7178_y0);
  and_gate and_gate_h_u_cla32_and7179_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7179_y0);
  and_gate and_gate_h_u_cla32_and7180_y0(h_u_cla32_and7179_y0, h_u_cla32_and7178_y0, h_u_cla32_and7180_y0);
  and_gate and_gate_h_u_cla32_and7181_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7181_y0);
  and_gate and_gate_h_u_cla32_and7182_y0(h_u_cla32_and7181_y0, h_u_cla32_and7180_y0, h_u_cla32_and7182_y0);
  and_gate and_gate_h_u_cla32_and7183_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7183_y0);
  and_gate and_gate_h_u_cla32_and7184_y0(h_u_cla32_and7183_y0, h_u_cla32_and7182_y0, h_u_cla32_and7184_y0);
  and_gate and_gate_h_u_cla32_and7185_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7185_y0);
  and_gate and_gate_h_u_cla32_and7186_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7186_y0);
  and_gate and_gate_h_u_cla32_and7187_y0(h_u_cla32_and7186_y0, h_u_cla32_and7185_y0, h_u_cla32_and7187_y0);
  and_gate and_gate_h_u_cla32_and7188_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7188_y0);
  and_gate and_gate_h_u_cla32_and7189_y0(h_u_cla32_and7188_y0, h_u_cla32_and7187_y0, h_u_cla32_and7189_y0);
  and_gate and_gate_h_u_cla32_and7190_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7190_y0);
  and_gate and_gate_h_u_cla32_and7191_y0(h_u_cla32_and7190_y0, h_u_cla32_and7189_y0, h_u_cla32_and7191_y0);
  and_gate and_gate_h_u_cla32_and7192_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7192_y0);
  and_gate and_gate_h_u_cla32_and7193_y0(h_u_cla32_and7192_y0, h_u_cla32_and7191_y0, h_u_cla32_and7193_y0);
  and_gate and_gate_h_u_cla32_and7194_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7194_y0);
  and_gate and_gate_h_u_cla32_and7195_y0(h_u_cla32_and7194_y0, h_u_cla32_and7193_y0, h_u_cla32_and7195_y0);
  and_gate and_gate_h_u_cla32_and7196_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7196_y0);
  and_gate and_gate_h_u_cla32_and7197_y0(h_u_cla32_and7196_y0, h_u_cla32_and7195_y0, h_u_cla32_and7197_y0);
  and_gate and_gate_h_u_cla32_and7198_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7198_y0);
  and_gate and_gate_h_u_cla32_and7199_y0(h_u_cla32_and7198_y0, h_u_cla32_and7197_y0, h_u_cla32_and7199_y0);
  and_gate and_gate_h_u_cla32_and7200_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7200_y0);
  and_gate and_gate_h_u_cla32_and7201_y0(h_u_cla32_and7200_y0, h_u_cla32_and7199_y0, h_u_cla32_and7201_y0);
  and_gate and_gate_h_u_cla32_and7202_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7202_y0);
  and_gate and_gate_h_u_cla32_and7203_y0(h_u_cla32_and7202_y0, h_u_cla32_and7201_y0, h_u_cla32_and7203_y0);
  and_gate and_gate_h_u_cla32_and7204_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7204_y0);
  and_gate and_gate_h_u_cla32_and7205_y0(h_u_cla32_and7204_y0, h_u_cla32_and7203_y0, h_u_cla32_and7205_y0);
  and_gate and_gate_h_u_cla32_and7206_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7206_y0);
  and_gate and_gate_h_u_cla32_and7207_y0(h_u_cla32_and7206_y0, h_u_cla32_and7205_y0, h_u_cla32_and7207_y0);
  and_gate and_gate_h_u_cla32_and7208_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7208_y0);
  and_gate and_gate_h_u_cla32_and7209_y0(h_u_cla32_and7208_y0, h_u_cla32_and7207_y0, h_u_cla32_and7209_y0);
  and_gate and_gate_h_u_cla32_and7210_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7210_y0);
  and_gate and_gate_h_u_cla32_and7211_y0(h_u_cla32_and7210_y0, h_u_cla32_and7209_y0, h_u_cla32_and7211_y0);
  and_gate and_gate_h_u_cla32_and7212_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7212_y0);
  and_gate and_gate_h_u_cla32_and7213_y0(h_u_cla32_and7212_y0, h_u_cla32_and7211_y0, h_u_cla32_and7213_y0);
  and_gate and_gate_h_u_cla32_and7214_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7214_y0);
  and_gate and_gate_h_u_cla32_and7215_y0(h_u_cla32_and7214_y0, h_u_cla32_and7213_y0, h_u_cla32_and7215_y0);
  and_gate and_gate_h_u_cla32_and7216_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7216_y0);
  and_gate and_gate_h_u_cla32_and7217_y0(h_u_cla32_and7216_y0, h_u_cla32_and7215_y0, h_u_cla32_and7217_y0);
  and_gate and_gate_h_u_cla32_and7218_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7218_y0);
  and_gate and_gate_h_u_cla32_and7219_y0(h_u_cla32_and7218_y0, h_u_cla32_and7217_y0, h_u_cla32_and7219_y0);
  and_gate and_gate_h_u_cla32_and7220_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7220_y0);
  and_gate and_gate_h_u_cla32_and7221_y0(h_u_cla32_and7220_y0, h_u_cla32_and7219_y0, h_u_cla32_and7221_y0);
  and_gate and_gate_h_u_cla32_and7222_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7222_y0);
  and_gate and_gate_h_u_cla32_and7223_y0(h_u_cla32_and7222_y0, h_u_cla32_and7221_y0, h_u_cla32_and7223_y0);
  and_gate and_gate_h_u_cla32_and7224_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7224_y0);
  and_gate and_gate_h_u_cla32_and7225_y0(h_u_cla32_and7224_y0, h_u_cla32_and7223_y0, h_u_cla32_and7225_y0);
  and_gate and_gate_h_u_cla32_and7226_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7226_y0);
  and_gate and_gate_h_u_cla32_and7227_y0(h_u_cla32_and7226_y0, h_u_cla32_and7225_y0, h_u_cla32_and7227_y0);
  and_gate and_gate_h_u_cla32_and7228_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7228_y0);
  and_gate and_gate_h_u_cla32_and7229_y0(h_u_cla32_and7228_y0, h_u_cla32_and7227_y0, h_u_cla32_and7229_y0);
  and_gate and_gate_h_u_cla32_and7230_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7230_y0);
  and_gate and_gate_h_u_cla32_and7231_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7231_y0);
  and_gate and_gate_h_u_cla32_and7232_y0(h_u_cla32_and7231_y0, h_u_cla32_and7230_y0, h_u_cla32_and7232_y0);
  and_gate and_gate_h_u_cla32_and7233_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7233_y0);
  and_gate and_gate_h_u_cla32_and7234_y0(h_u_cla32_and7233_y0, h_u_cla32_and7232_y0, h_u_cla32_and7234_y0);
  and_gate and_gate_h_u_cla32_and7235_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7235_y0);
  and_gate and_gate_h_u_cla32_and7236_y0(h_u_cla32_and7235_y0, h_u_cla32_and7234_y0, h_u_cla32_and7236_y0);
  and_gate and_gate_h_u_cla32_and7237_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7237_y0);
  and_gate and_gate_h_u_cla32_and7238_y0(h_u_cla32_and7237_y0, h_u_cla32_and7236_y0, h_u_cla32_and7238_y0);
  and_gate and_gate_h_u_cla32_and7239_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7239_y0);
  and_gate and_gate_h_u_cla32_and7240_y0(h_u_cla32_and7239_y0, h_u_cla32_and7238_y0, h_u_cla32_and7240_y0);
  and_gate and_gate_h_u_cla32_and7241_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7241_y0);
  and_gate and_gate_h_u_cla32_and7242_y0(h_u_cla32_and7241_y0, h_u_cla32_and7240_y0, h_u_cla32_and7242_y0);
  and_gate and_gate_h_u_cla32_and7243_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7243_y0);
  and_gate and_gate_h_u_cla32_and7244_y0(h_u_cla32_and7243_y0, h_u_cla32_and7242_y0, h_u_cla32_and7244_y0);
  and_gate and_gate_h_u_cla32_and7245_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7245_y0);
  and_gate and_gate_h_u_cla32_and7246_y0(h_u_cla32_and7245_y0, h_u_cla32_and7244_y0, h_u_cla32_and7246_y0);
  and_gate and_gate_h_u_cla32_and7247_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7247_y0);
  and_gate and_gate_h_u_cla32_and7248_y0(h_u_cla32_and7247_y0, h_u_cla32_and7246_y0, h_u_cla32_and7248_y0);
  and_gate and_gate_h_u_cla32_and7249_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7249_y0);
  and_gate and_gate_h_u_cla32_and7250_y0(h_u_cla32_and7249_y0, h_u_cla32_and7248_y0, h_u_cla32_and7250_y0);
  and_gate and_gate_h_u_cla32_and7251_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7251_y0);
  and_gate and_gate_h_u_cla32_and7252_y0(h_u_cla32_and7251_y0, h_u_cla32_and7250_y0, h_u_cla32_and7252_y0);
  and_gate and_gate_h_u_cla32_and7253_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7253_y0);
  and_gate and_gate_h_u_cla32_and7254_y0(h_u_cla32_and7253_y0, h_u_cla32_and7252_y0, h_u_cla32_and7254_y0);
  and_gate and_gate_h_u_cla32_and7255_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7255_y0);
  and_gate and_gate_h_u_cla32_and7256_y0(h_u_cla32_and7255_y0, h_u_cla32_and7254_y0, h_u_cla32_and7256_y0);
  and_gate and_gate_h_u_cla32_and7257_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7257_y0);
  and_gate and_gate_h_u_cla32_and7258_y0(h_u_cla32_and7257_y0, h_u_cla32_and7256_y0, h_u_cla32_and7258_y0);
  and_gate and_gate_h_u_cla32_and7259_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7259_y0);
  and_gate and_gate_h_u_cla32_and7260_y0(h_u_cla32_and7259_y0, h_u_cla32_and7258_y0, h_u_cla32_and7260_y0);
  and_gate and_gate_h_u_cla32_and7261_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7261_y0);
  and_gate and_gate_h_u_cla32_and7262_y0(h_u_cla32_and7261_y0, h_u_cla32_and7260_y0, h_u_cla32_and7262_y0);
  and_gate and_gate_h_u_cla32_and7263_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7263_y0);
  and_gate and_gate_h_u_cla32_and7264_y0(h_u_cla32_and7263_y0, h_u_cla32_and7262_y0, h_u_cla32_and7264_y0);
  and_gate and_gate_h_u_cla32_and7265_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7265_y0);
  and_gate and_gate_h_u_cla32_and7266_y0(h_u_cla32_and7265_y0, h_u_cla32_and7264_y0, h_u_cla32_and7266_y0);
  and_gate and_gate_h_u_cla32_and7267_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7267_y0);
  and_gate and_gate_h_u_cla32_and7268_y0(h_u_cla32_and7267_y0, h_u_cla32_and7266_y0, h_u_cla32_and7268_y0);
  and_gate and_gate_h_u_cla32_and7269_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7269_y0);
  and_gate and_gate_h_u_cla32_and7270_y0(h_u_cla32_and7269_y0, h_u_cla32_and7268_y0, h_u_cla32_and7270_y0);
  and_gate and_gate_h_u_cla32_and7271_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and7271_y0);
  and_gate and_gate_h_u_cla32_and7272_y0(h_u_cla32_and7271_y0, h_u_cla32_and7270_y0, h_u_cla32_and7272_y0);
  and_gate and_gate_h_u_cla32_and7273_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7273_y0);
  and_gate and_gate_h_u_cla32_and7274_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7274_y0);
  and_gate and_gate_h_u_cla32_and7275_y0(h_u_cla32_and7274_y0, h_u_cla32_and7273_y0, h_u_cla32_and7275_y0);
  and_gate and_gate_h_u_cla32_and7276_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7276_y0);
  and_gate and_gate_h_u_cla32_and7277_y0(h_u_cla32_and7276_y0, h_u_cla32_and7275_y0, h_u_cla32_and7277_y0);
  and_gate and_gate_h_u_cla32_and7278_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7278_y0);
  and_gate and_gate_h_u_cla32_and7279_y0(h_u_cla32_and7278_y0, h_u_cla32_and7277_y0, h_u_cla32_and7279_y0);
  and_gate and_gate_h_u_cla32_and7280_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7280_y0);
  and_gate and_gate_h_u_cla32_and7281_y0(h_u_cla32_and7280_y0, h_u_cla32_and7279_y0, h_u_cla32_and7281_y0);
  and_gate and_gate_h_u_cla32_and7282_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7282_y0);
  and_gate and_gate_h_u_cla32_and7283_y0(h_u_cla32_and7282_y0, h_u_cla32_and7281_y0, h_u_cla32_and7283_y0);
  and_gate and_gate_h_u_cla32_and7284_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7284_y0);
  and_gate and_gate_h_u_cla32_and7285_y0(h_u_cla32_and7284_y0, h_u_cla32_and7283_y0, h_u_cla32_and7285_y0);
  and_gate and_gate_h_u_cla32_and7286_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7286_y0);
  and_gate and_gate_h_u_cla32_and7287_y0(h_u_cla32_and7286_y0, h_u_cla32_and7285_y0, h_u_cla32_and7287_y0);
  and_gate and_gate_h_u_cla32_and7288_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7288_y0);
  and_gate and_gate_h_u_cla32_and7289_y0(h_u_cla32_and7288_y0, h_u_cla32_and7287_y0, h_u_cla32_and7289_y0);
  and_gate and_gate_h_u_cla32_and7290_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7290_y0);
  and_gate and_gate_h_u_cla32_and7291_y0(h_u_cla32_and7290_y0, h_u_cla32_and7289_y0, h_u_cla32_and7291_y0);
  and_gate and_gate_h_u_cla32_and7292_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7292_y0);
  and_gate and_gate_h_u_cla32_and7293_y0(h_u_cla32_and7292_y0, h_u_cla32_and7291_y0, h_u_cla32_and7293_y0);
  and_gate and_gate_h_u_cla32_and7294_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7294_y0);
  and_gate and_gate_h_u_cla32_and7295_y0(h_u_cla32_and7294_y0, h_u_cla32_and7293_y0, h_u_cla32_and7295_y0);
  and_gate and_gate_h_u_cla32_and7296_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7296_y0);
  and_gate and_gate_h_u_cla32_and7297_y0(h_u_cla32_and7296_y0, h_u_cla32_and7295_y0, h_u_cla32_and7297_y0);
  and_gate and_gate_h_u_cla32_and7298_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7298_y0);
  and_gate and_gate_h_u_cla32_and7299_y0(h_u_cla32_and7298_y0, h_u_cla32_and7297_y0, h_u_cla32_and7299_y0);
  and_gate and_gate_h_u_cla32_and7300_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7300_y0);
  and_gate and_gate_h_u_cla32_and7301_y0(h_u_cla32_and7300_y0, h_u_cla32_and7299_y0, h_u_cla32_and7301_y0);
  and_gate and_gate_h_u_cla32_and7302_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7302_y0);
  and_gate and_gate_h_u_cla32_and7303_y0(h_u_cla32_and7302_y0, h_u_cla32_and7301_y0, h_u_cla32_and7303_y0);
  and_gate and_gate_h_u_cla32_and7304_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7304_y0);
  and_gate and_gate_h_u_cla32_and7305_y0(h_u_cla32_and7304_y0, h_u_cla32_and7303_y0, h_u_cla32_and7305_y0);
  and_gate and_gate_h_u_cla32_and7306_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7306_y0);
  and_gate and_gate_h_u_cla32_and7307_y0(h_u_cla32_and7306_y0, h_u_cla32_and7305_y0, h_u_cla32_and7307_y0);
  and_gate and_gate_h_u_cla32_and7308_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7308_y0);
  and_gate and_gate_h_u_cla32_and7309_y0(h_u_cla32_and7308_y0, h_u_cla32_and7307_y0, h_u_cla32_and7309_y0);
  and_gate and_gate_h_u_cla32_and7310_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7310_y0);
  and_gate and_gate_h_u_cla32_and7311_y0(h_u_cla32_and7310_y0, h_u_cla32_and7309_y0, h_u_cla32_and7311_y0);
  and_gate and_gate_h_u_cla32_and7312_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and7312_y0);
  and_gate and_gate_h_u_cla32_and7313_y0(h_u_cla32_and7312_y0, h_u_cla32_and7311_y0, h_u_cla32_and7313_y0);
  and_gate and_gate_h_u_cla32_and7314_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7314_y0);
  and_gate and_gate_h_u_cla32_and7315_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7315_y0);
  and_gate and_gate_h_u_cla32_and7316_y0(h_u_cla32_and7315_y0, h_u_cla32_and7314_y0, h_u_cla32_and7316_y0);
  and_gate and_gate_h_u_cla32_and7317_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7317_y0);
  and_gate and_gate_h_u_cla32_and7318_y0(h_u_cla32_and7317_y0, h_u_cla32_and7316_y0, h_u_cla32_and7318_y0);
  and_gate and_gate_h_u_cla32_and7319_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7319_y0);
  and_gate and_gate_h_u_cla32_and7320_y0(h_u_cla32_and7319_y0, h_u_cla32_and7318_y0, h_u_cla32_and7320_y0);
  and_gate and_gate_h_u_cla32_and7321_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7321_y0);
  and_gate and_gate_h_u_cla32_and7322_y0(h_u_cla32_and7321_y0, h_u_cla32_and7320_y0, h_u_cla32_and7322_y0);
  and_gate and_gate_h_u_cla32_and7323_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7323_y0);
  and_gate and_gate_h_u_cla32_and7324_y0(h_u_cla32_and7323_y0, h_u_cla32_and7322_y0, h_u_cla32_and7324_y0);
  and_gate and_gate_h_u_cla32_and7325_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7325_y0);
  and_gate and_gate_h_u_cla32_and7326_y0(h_u_cla32_and7325_y0, h_u_cla32_and7324_y0, h_u_cla32_and7326_y0);
  and_gate and_gate_h_u_cla32_and7327_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7327_y0);
  and_gate and_gate_h_u_cla32_and7328_y0(h_u_cla32_and7327_y0, h_u_cla32_and7326_y0, h_u_cla32_and7328_y0);
  and_gate and_gate_h_u_cla32_and7329_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7329_y0);
  and_gate and_gate_h_u_cla32_and7330_y0(h_u_cla32_and7329_y0, h_u_cla32_and7328_y0, h_u_cla32_and7330_y0);
  and_gate and_gate_h_u_cla32_and7331_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7331_y0);
  and_gate and_gate_h_u_cla32_and7332_y0(h_u_cla32_and7331_y0, h_u_cla32_and7330_y0, h_u_cla32_and7332_y0);
  and_gate and_gate_h_u_cla32_and7333_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7333_y0);
  and_gate and_gate_h_u_cla32_and7334_y0(h_u_cla32_and7333_y0, h_u_cla32_and7332_y0, h_u_cla32_and7334_y0);
  and_gate and_gate_h_u_cla32_and7335_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7335_y0);
  and_gate and_gate_h_u_cla32_and7336_y0(h_u_cla32_and7335_y0, h_u_cla32_and7334_y0, h_u_cla32_and7336_y0);
  and_gate and_gate_h_u_cla32_and7337_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7337_y0);
  and_gate and_gate_h_u_cla32_and7338_y0(h_u_cla32_and7337_y0, h_u_cla32_and7336_y0, h_u_cla32_and7338_y0);
  and_gate and_gate_h_u_cla32_and7339_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7339_y0);
  and_gate and_gate_h_u_cla32_and7340_y0(h_u_cla32_and7339_y0, h_u_cla32_and7338_y0, h_u_cla32_and7340_y0);
  and_gate and_gate_h_u_cla32_and7341_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7341_y0);
  and_gate and_gate_h_u_cla32_and7342_y0(h_u_cla32_and7341_y0, h_u_cla32_and7340_y0, h_u_cla32_and7342_y0);
  and_gate and_gate_h_u_cla32_and7343_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7343_y0);
  and_gate and_gate_h_u_cla32_and7344_y0(h_u_cla32_and7343_y0, h_u_cla32_and7342_y0, h_u_cla32_and7344_y0);
  and_gate and_gate_h_u_cla32_and7345_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7345_y0);
  and_gate and_gate_h_u_cla32_and7346_y0(h_u_cla32_and7345_y0, h_u_cla32_and7344_y0, h_u_cla32_and7346_y0);
  and_gate and_gate_h_u_cla32_and7347_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7347_y0);
  and_gate and_gate_h_u_cla32_and7348_y0(h_u_cla32_and7347_y0, h_u_cla32_and7346_y0, h_u_cla32_and7348_y0);
  and_gate and_gate_h_u_cla32_and7349_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7349_y0);
  and_gate and_gate_h_u_cla32_and7350_y0(h_u_cla32_and7349_y0, h_u_cla32_and7348_y0, h_u_cla32_and7350_y0);
  and_gate and_gate_h_u_cla32_and7351_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and7351_y0);
  and_gate and_gate_h_u_cla32_and7352_y0(h_u_cla32_and7351_y0, h_u_cla32_and7350_y0, h_u_cla32_and7352_y0);
  and_gate and_gate_h_u_cla32_and7353_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7353_y0);
  and_gate and_gate_h_u_cla32_and7354_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7354_y0);
  and_gate and_gate_h_u_cla32_and7355_y0(h_u_cla32_and7354_y0, h_u_cla32_and7353_y0, h_u_cla32_and7355_y0);
  and_gate and_gate_h_u_cla32_and7356_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7356_y0);
  and_gate and_gate_h_u_cla32_and7357_y0(h_u_cla32_and7356_y0, h_u_cla32_and7355_y0, h_u_cla32_and7357_y0);
  and_gate and_gate_h_u_cla32_and7358_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7358_y0);
  and_gate and_gate_h_u_cla32_and7359_y0(h_u_cla32_and7358_y0, h_u_cla32_and7357_y0, h_u_cla32_and7359_y0);
  and_gate and_gate_h_u_cla32_and7360_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7360_y0);
  and_gate and_gate_h_u_cla32_and7361_y0(h_u_cla32_and7360_y0, h_u_cla32_and7359_y0, h_u_cla32_and7361_y0);
  and_gate and_gate_h_u_cla32_and7362_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7362_y0);
  and_gate and_gate_h_u_cla32_and7363_y0(h_u_cla32_and7362_y0, h_u_cla32_and7361_y0, h_u_cla32_and7363_y0);
  and_gate and_gate_h_u_cla32_and7364_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7364_y0);
  and_gate and_gate_h_u_cla32_and7365_y0(h_u_cla32_and7364_y0, h_u_cla32_and7363_y0, h_u_cla32_and7365_y0);
  and_gate and_gate_h_u_cla32_and7366_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7366_y0);
  and_gate and_gate_h_u_cla32_and7367_y0(h_u_cla32_and7366_y0, h_u_cla32_and7365_y0, h_u_cla32_and7367_y0);
  and_gate and_gate_h_u_cla32_and7368_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7368_y0);
  and_gate and_gate_h_u_cla32_and7369_y0(h_u_cla32_and7368_y0, h_u_cla32_and7367_y0, h_u_cla32_and7369_y0);
  and_gate and_gate_h_u_cla32_and7370_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7370_y0);
  and_gate and_gate_h_u_cla32_and7371_y0(h_u_cla32_and7370_y0, h_u_cla32_and7369_y0, h_u_cla32_and7371_y0);
  and_gate and_gate_h_u_cla32_and7372_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7372_y0);
  and_gate and_gate_h_u_cla32_and7373_y0(h_u_cla32_and7372_y0, h_u_cla32_and7371_y0, h_u_cla32_and7373_y0);
  and_gate and_gate_h_u_cla32_and7374_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7374_y0);
  and_gate and_gate_h_u_cla32_and7375_y0(h_u_cla32_and7374_y0, h_u_cla32_and7373_y0, h_u_cla32_and7375_y0);
  and_gate and_gate_h_u_cla32_and7376_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7376_y0);
  and_gate and_gate_h_u_cla32_and7377_y0(h_u_cla32_and7376_y0, h_u_cla32_and7375_y0, h_u_cla32_and7377_y0);
  and_gate and_gate_h_u_cla32_and7378_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7378_y0);
  and_gate and_gate_h_u_cla32_and7379_y0(h_u_cla32_and7378_y0, h_u_cla32_and7377_y0, h_u_cla32_and7379_y0);
  and_gate and_gate_h_u_cla32_and7380_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7380_y0);
  and_gate and_gate_h_u_cla32_and7381_y0(h_u_cla32_and7380_y0, h_u_cla32_and7379_y0, h_u_cla32_and7381_y0);
  and_gate and_gate_h_u_cla32_and7382_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7382_y0);
  and_gate and_gate_h_u_cla32_and7383_y0(h_u_cla32_and7382_y0, h_u_cla32_and7381_y0, h_u_cla32_and7383_y0);
  and_gate and_gate_h_u_cla32_and7384_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7384_y0);
  and_gate and_gate_h_u_cla32_and7385_y0(h_u_cla32_and7384_y0, h_u_cla32_and7383_y0, h_u_cla32_and7385_y0);
  and_gate and_gate_h_u_cla32_and7386_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7386_y0);
  and_gate and_gate_h_u_cla32_and7387_y0(h_u_cla32_and7386_y0, h_u_cla32_and7385_y0, h_u_cla32_and7387_y0);
  and_gate and_gate_h_u_cla32_and7388_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and7388_y0);
  and_gate and_gate_h_u_cla32_and7389_y0(h_u_cla32_and7388_y0, h_u_cla32_and7387_y0, h_u_cla32_and7389_y0);
  and_gate and_gate_h_u_cla32_and7390_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7390_y0);
  and_gate and_gate_h_u_cla32_and7391_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7391_y0);
  and_gate and_gate_h_u_cla32_and7392_y0(h_u_cla32_and7391_y0, h_u_cla32_and7390_y0, h_u_cla32_and7392_y0);
  and_gate and_gate_h_u_cla32_and7393_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7393_y0);
  and_gate and_gate_h_u_cla32_and7394_y0(h_u_cla32_and7393_y0, h_u_cla32_and7392_y0, h_u_cla32_and7394_y0);
  and_gate and_gate_h_u_cla32_and7395_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7395_y0);
  and_gate and_gate_h_u_cla32_and7396_y0(h_u_cla32_and7395_y0, h_u_cla32_and7394_y0, h_u_cla32_and7396_y0);
  and_gate and_gate_h_u_cla32_and7397_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7397_y0);
  and_gate and_gate_h_u_cla32_and7398_y0(h_u_cla32_and7397_y0, h_u_cla32_and7396_y0, h_u_cla32_and7398_y0);
  and_gate and_gate_h_u_cla32_and7399_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7399_y0);
  and_gate and_gate_h_u_cla32_and7400_y0(h_u_cla32_and7399_y0, h_u_cla32_and7398_y0, h_u_cla32_and7400_y0);
  and_gate and_gate_h_u_cla32_and7401_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7401_y0);
  and_gate and_gate_h_u_cla32_and7402_y0(h_u_cla32_and7401_y0, h_u_cla32_and7400_y0, h_u_cla32_and7402_y0);
  and_gate and_gate_h_u_cla32_and7403_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7403_y0);
  and_gate and_gate_h_u_cla32_and7404_y0(h_u_cla32_and7403_y0, h_u_cla32_and7402_y0, h_u_cla32_and7404_y0);
  and_gate and_gate_h_u_cla32_and7405_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7405_y0);
  and_gate and_gate_h_u_cla32_and7406_y0(h_u_cla32_and7405_y0, h_u_cla32_and7404_y0, h_u_cla32_and7406_y0);
  and_gate and_gate_h_u_cla32_and7407_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7407_y0);
  and_gate and_gate_h_u_cla32_and7408_y0(h_u_cla32_and7407_y0, h_u_cla32_and7406_y0, h_u_cla32_and7408_y0);
  and_gate and_gate_h_u_cla32_and7409_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7409_y0);
  and_gate and_gate_h_u_cla32_and7410_y0(h_u_cla32_and7409_y0, h_u_cla32_and7408_y0, h_u_cla32_and7410_y0);
  and_gate and_gate_h_u_cla32_and7411_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7411_y0);
  and_gate and_gate_h_u_cla32_and7412_y0(h_u_cla32_and7411_y0, h_u_cla32_and7410_y0, h_u_cla32_and7412_y0);
  and_gate and_gate_h_u_cla32_and7413_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7413_y0);
  and_gate and_gate_h_u_cla32_and7414_y0(h_u_cla32_and7413_y0, h_u_cla32_and7412_y0, h_u_cla32_and7414_y0);
  and_gate and_gate_h_u_cla32_and7415_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7415_y0);
  and_gate and_gate_h_u_cla32_and7416_y0(h_u_cla32_and7415_y0, h_u_cla32_and7414_y0, h_u_cla32_and7416_y0);
  and_gate and_gate_h_u_cla32_and7417_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7417_y0);
  and_gate and_gate_h_u_cla32_and7418_y0(h_u_cla32_and7417_y0, h_u_cla32_and7416_y0, h_u_cla32_and7418_y0);
  and_gate and_gate_h_u_cla32_and7419_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7419_y0);
  and_gate and_gate_h_u_cla32_and7420_y0(h_u_cla32_and7419_y0, h_u_cla32_and7418_y0, h_u_cla32_and7420_y0);
  and_gate and_gate_h_u_cla32_and7421_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7421_y0);
  and_gate and_gate_h_u_cla32_and7422_y0(h_u_cla32_and7421_y0, h_u_cla32_and7420_y0, h_u_cla32_and7422_y0);
  and_gate and_gate_h_u_cla32_and7423_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and7423_y0);
  and_gate and_gate_h_u_cla32_and7424_y0(h_u_cla32_and7423_y0, h_u_cla32_and7422_y0, h_u_cla32_and7424_y0);
  and_gate and_gate_h_u_cla32_and7425_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7425_y0);
  and_gate and_gate_h_u_cla32_and7426_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7426_y0);
  and_gate and_gate_h_u_cla32_and7427_y0(h_u_cla32_and7426_y0, h_u_cla32_and7425_y0, h_u_cla32_and7427_y0);
  and_gate and_gate_h_u_cla32_and7428_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7428_y0);
  and_gate and_gate_h_u_cla32_and7429_y0(h_u_cla32_and7428_y0, h_u_cla32_and7427_y0, h_u_cla32_and7429_y0);
  and_gate and_gate_h_u_cla32_and7430_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7430_y0);
  and_gate and_gate_h_u_cla32_and7431_y0(h_u_cla32_and7430_y0, h_u_cla32_and7429_y0, h_u_cla32_and7431_y0);
  and_gate and_gate_h_u_cla32_and7432_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7432_y0);
  and_gate and_gate_h_u_cla32_and7433_y0(h_u_cla32_and7432_y0, h_u_cla32_and7431_y0, h_u_cla32_and7433_y0);
  and_gate and_gate_h_u_cla32_and7434_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7434_y0);
  and_gate and_gate_h_u_cla32_and7435_y0(h_u_cla32_and7434_y0, h_u_cla32_and7433_y0, h_u_cla32_and7435_y0);
  and_gate and_gate_h_u_cla32_and7436_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7436_y0);
  and_gate and_gate_h_u_cla32_and7437_y0(h_u_cla32_and7436_y0, h_u_cla32_and7435_y0, h_u_cla32_and7437_y0);
  and_gate and_gate_h_u_cla32_and7438_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7438_y0);
  and_gate and_gate_h_u_cla32_and7439_y0(h_u_cla32_and7438_y0, h_u_cla32_and7437_y0, h_u_cla32_and7439_y0);
  and_gate and_gate_h_u_cla32_and7440_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7440_y0);
  and_gate and_gate_h_u_cla32_and7441_y0(h_u_cla32_and7440_y0, h_u_cla32_and7439_y0, h_u_cla32_and7441_y0);
  and_gate and_gate_h_u_cla32_and7442_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7442_y0);
  and_gate and_gate_h_u_cla32_and7443_y0(h_u_cla32_and7442_y0, h_u_cla32_and7441_y0, h_u_cla32_and7443_y0);
  and_gate and_gate_h_u_cla32_and7444_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7444_y0);
  and_gate and_gate_h_u_cla32_and7445_y0(h_u_cla32_and7444_y0, h_u_cla32_and7443_y0, h_u_cla32_and7445_y0);
  and_gate and_gate_h_u_cla32_and7446_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7446_y0);
  and_gate and_gate_h_u_cla32_and7447_y0(h_u_cla32_and7446_y0, h_u_cla32_and7445_y0, h_u_cla32_and7447_y0);
  and_gate and_gate_h_u_cla32_and7448_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7448_y0);
  and_gate and_gate_h_u_cla32_and7449_y0(h_u_cla32_and7448_y0, h_u_cla32_and7447_y0, h_u_cla32_and7449_y0);
  and_gate and_gate_h_u_cla32_and7450_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7450_y0);
  and_gate and_gate_h_u_cla32_and7451_y0(h_u_cla32_and7450_y0, h_u_cla32_and7449_y0, h_u_cla32_and7451_y0);
  and_gate and_gate_h_u_cla32_and7452_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7452_y0);
  and_gate and_gate_h_u_cla32_and7453_y0(h_u_cla32_and7452_y0, h_u_cla32_and7451_y0, h_u_cla32_and7453_y0);
  and_gate and_gate_h_u_cla32_and7454_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7454_y0);
  and_gate and_gate_h_u_cla32_and7455_y0(h_u_cla32_and7454_y0, h_u_cla32_and7453_y0, h_u_cla32_and7455_y0);
  and_gate and_gate_h_u_cla32_and7456_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and7456_y0);
  and_gate and_gate_h_u_cla32_and7457_y0(h_u_cla32_and7456_y0, h_u_cla32_and7455_y0, h_u_cla32_and7457_y0);
  and_gate and_gate_h_u_cla32_and7458_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7458_y0);
  and_gate and_gate_h_u_cla32_and7459_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7459_y0);
  and_gate and_gate_h_u_cla32_and7460_y0(h_u_cla32_and7459_y0, h_u_cla32_and7458_y0, h_u_cla32_and7460_y0);
  and_gate and_gate_h_u_cla32_and7461_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7461_y0);
  and_gate and_gate_h_u_cla32_and7462_y0(h_u_cla32_and7461_y0, h_u_cla32_and7460_y0, h_u_cla32_and7462_y0);
  and_gate and_gate_h_u_cla32_and7463_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7463_y0);
  and_gate and_gate_h_u_cla32_and7464_y0(h_u_cla32_and7463_y0, h_u_cla32_and7462_y0, h_u_cla32_and7464_y0);
  and_gate and_gate_h_u_cla32_and7465_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7465_y0);
  and_gate and_gate_h_u_cla32_and7466_y0(h_u_cla32_and7465_y0, h_u_cla32_and7464_y0, h_u_cla32_and7466_y0);
  and_gate and_gate_h_u_cla32_and7467_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7467_y0);
  and_gate and_gate_h_u_cla32_and7468_y0(h_u_cla32_and7467_y0, h_u_cla32_and7466_y0, h_u_cla32_and7468_y0);
  and_gate and_gate_h_u_cla32_and7469_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7469_y0);
  and_gate and_gate_h_u_cla32_and7470_y0(h_u_cla32_and7469_y0, h_u_cla32_and7468_y0, h_u_cla32_and7470_y0);
  and_gate and_gate_h_u_cla32_and7471_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7471_y0);
  and_gate and_gate_h_u_cla32_and7472_y0(h_u_cla32_and7471_y0, h_u_cla32_and7470_y0, h_u_cla32_and7472_y0);
  and_gate and_gate_h_u_cla32_and7473_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7473_y0);
  and_gate and_gate_h_u_cla32_and7474_y0(h_u_cla32_and7473_y0, h_u_cla32_and7472_y0, h_u_cla32_and7474_y0);
  and_gate and_gate_h_u_cla32_and7475_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7475_y0);
  and_gate and_gate_h_u_cla32_and7476_y0(h_u_cla32_and7475_y0, h_u_cla32_and7474_y0, h_u_cla32_and7476_y0);
  and_gate and_gate_h_u_cla32_and7477_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7477_y0);
  and_gate and_gate_h_u_cla32_and7478_y0(h_u_cla32_and7477_y0, h_u_cla32_and7476_y0, h_u_cla32_and7478_y0);
  and_gate and_gate_h_u_cla32_and7479_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7479_y0);
  and_gate and_gate_h_u_cla32_and7480_y0(h_u_cla32_and7479_y0, h_u_cla32_and7478_y0, h_u_cla32_and7480_y0);
  and_gate and_gate_h_u_cla32_and7481_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7481_y0);
  and_gate and_gate_h_u_cla32_and7482_y0(h_u_cla32_and7481_y0, h_u_cla32_and7480_y0, h_u_cla32_and7482_y0);
  and_gate and_gate_h_u_cla32_and7483_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7483_y0);
  and_gate and_gate_h_u_cla32_and7484_y0(h_u_cla32_and7483_y0, h_u_cla32_and7482_y0, h_u_cla32_and7484_y0);
  and_gate and_gate_h_u_cla32_and7485_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7485_y0);
  and_gate and_gate_h_u_cla32_and7486_y0(h_u_cla32_and7485_y0, h_u_cla32_and7484_y0, h_u_cla32_and7486_y0);
  and_gate and_gate_h_u_cla32_and7487_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and7487_y0);
  and_gate and_gate_h_u_cla32_and7488_y0(h_u_cla32_and7487_y0, h_u_cla32_and7486_y0, h_u_cla32_and7488_y0);
  and_gate and_gate_h_u_cla32_and7489_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7489_y0);
  and_gate and_gate_h_u_cla32_and7490_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7490_y0);
  and_gate and_gate_h_u_cla32_and7491_y0(h_u_cla32_and7490_y0, h_u_cla32_and7489_y0, h_u_cla32_and7491_y0);
  and_gate and_gate_h_u_cla32_and7492_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7492_y0);
  and_gate and_gate_h_u_cla32_and7493_y0(h_u_cla32_and7492_y0, h_u_cla32_and7491_y0, h_u_cla32_and7493_y0);
  and_gate and_gate_h_u_cla32_and7494_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7494_y0);
  and_gate and_gate_h_u_cla32_and7495_y0(h_u_cla32_and7494_y0, h_u_cla32_and7493_y0, h_u_cla32_and7495_y0);
  and_gate and_gate_h_u_cla32_and7496_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7496_y0);
  and_gate and_gate_h_u_cla32_and7497_y0(h_u_cla32_and7496_y0, h_u_cla32_and7495_y0, h_u_cla32_and7497_y0);
  and_gate and_gate_h_u_cla32_and7498_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7498_y0);
  and_gate and_gate_h_u_cla32_and7499_y0(h_u_cla32_and7498_y0, h_u_cla32_and7497_y0, h_u_cla32_and7499_y0);
  and_gate and_gate_h_u_cla32_and7500_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7500_y0);
  and_gate and_gate_h_u_cla32_and7501_y0(h_u_cla32_and7500_y0, h_u_cla32_and7499_y0, h_u_cla32_and7501_y0);
  and_gate and_gate_h_u_cla32_and7502_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7502_y0);
  and_gate and_gate_h_u_cla32_and7503_y0(h_u_cla32_and7502_y0, h_u_cla32_and7501_y0, h_u_cla32_and7503_y0);
  and_gate and_gate_h_u_cla32_and7504_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7504_y0);
  and_gate and_gate_h_u_cla32_and7505_y0(h_u_cla32_and7504_y0, h_u_cla32_and7503_y0, h_u_cla32_and7505_y0);
  and_gate and_gate_h_u_cla32_and7506_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7506_y0);
  and_gate and_gate_h_u_cla32_and7507_y0(h_u_cla32_and7506_y0, h_u_cla32_and7505_y0, h_u_cla32_and7507_y0);
  and_gate and_gate_h_u_cla32_and7508_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7508_y0);
  and_gate and_gate_h_u_cla32_and7509_y0(h_u_cla32_and7508_y0, h_u_cla32_and7507_y0, h_u_cla32_and7509_y0);
  and_gate and_gate_h_u_cla32_and7510_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7510_y0);
  and_gate and_gate_h_u_cla32_and7511_y0(h_u_cla32_and7510_y0, h_u_cla32_and7509_y0, h_u_cla32_and7511_y0);
  and_gate and_gate_h_u_cla32_and7512_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7512_y0);
  and_gate and_gate_h_u_cla32_and7513_y0(h_u_cla32_and7512_y0, h_u_cla32_and7511_y0, h_u_cla32_and7513_y0);
  and_gate and_gate_h_u_cla32_and7514_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7514_y0);
  and_gate and_gate_h_u_cla32_and7515_y0(h_u_cla32_and7514_y0, h_u_cla32_and7513_y0, h_u_cla32_and7515_y0);
  and_gate and_gate_h_u_cla32_and7516_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and7516_y0);
  and_gate and_gate_h_u_cla32_and7517_y0(h_u_cla32_and7516_y0, h_u_cla32_and7515_y0, h_u_cla32_and7517_y0);
  and_gate and_gate_h_u_cla32_and7518_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7518_y0);
  and_gate and_gate_h_u_cla32_and7519_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7519_y0);
  and_gate and_gate_h_u_cla32_and7520_y0(h_u_cla32_and7519_y0, h_u_cla32_and7518_y0, h_u_cla32_and7520_y0);
  and_gate and_gate_h_u_cla32_and7521_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7521_y0);
  and_gate and_gate_h_u_cla32_and7522_y0(h_u_cla32_and7521_y0, h_u_cla32_and7520_y0, h_u_cla32_and7522_y0);
  and_gate and_gate_h_u_cla32_and7523_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7523_y0);
  and_gate and_gate_h_u_cla32_and7524_y0(h_u_cla32_and7523_y0, h_u_cla32_and7522_y0, h_u_cla32_and7524_y0);
  and_gate and_gate_h_u_cla32_and7525_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7525_y0);
  and_gate and_gate_h_u_cla32_and7526_y0(h_u_cla32_and7525_y0, h_u_cla32_and7524_y0, h_u_cla32_and7526_y0);
  and_gate and_gate_h_u_cla32_and7527_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7527_y0);
  and_gate and_gate_h_u_cla32_and7528_y0(h_u_cla32_and7527_y0, h_u_cla32_and7526_y0, h_u_cla32_and7528_y0);
  and_gate and_gate_h_u_cla32_and7529_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7529_y0);
  and_gate and_gate_h_u_cla32_and7530_y0(h_u_cla32_and7529_y0, h_u_cla32_and7528_y0, h_u_cla32_and7530_y0);
  and_gate and_gate_h_u_cla32_and7531_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7531_y0);
  and_gate and_gate_h_u_cla32_and7532_y0(h_u_cla32_and7531_y0, h_u_cla32_and7530_y0, h_u_cla32_and7532_y0);
  and_gate and_gate_h_u_cla32_and7533_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7533_y0);
  and_gate and_gate_h_u_cla32_and7534_y0(h_u_cla32_and7533_y0, h_u_cla32_and7532_y0, h_u_cla32_and7534_y0);
  and_gate and_gate_h_u_cla32_and7535_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7535_y0);
  and_gate and_gate_h_u_cla32_and7536_y0(h_u_cla32_and7535_y0, h_u_cla32_and7534_y0, h_u_cla32_and7536_y0);
  and_gate and_gate_h_u_cla32_and7537_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7537_y0);
  and_gate and_gate_h_u_cla32_and7538_y0(h_u_cla32_and7537_y0, h_u_cla32_and7536_y0, h_u_cla32_and7538_y0);
  and_gate and_gate_h_u_cla32_and7539_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7539_y0);
  and_gate and_gate_h_u_cla32_and7540_y0(h_u_cla32_and7539_y0, h_u_cla32_and7538_y0, h_u_cla32_and7540_y0);
  and_gate and_gate_h_u_cla32_and7541_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7541_y0);
  and_gate and_gate_h_u_cla32_and7542_y0(h_u_cla32_and7541_y0, h_u_cla32_and7540_y0, h_u_cla32_and7542_y0);
  and_gate and_gate_h_u_cla32_and7543_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and7543_y0);
  and_gate and_gate_h_u_cla32_and7544_y0(h_u_cla32_and7543_y0, h_u_cla32_and7542_y0, h_u_cla32_and7544_y0);
  and_gate and_gate_h_u_cla32_and7545_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7545_y0);
  and_gate and_gate_h_u_cla32_and7546_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7546_y0);
  and_gate and_gate_h_u_cla32_and7547_y0(h_u_cla32_and7546_y0, h_u_cla32_and7545_y0, h_u_cla32_and7547_y0);
  and_gate and_gate_h_u_cla32_and7548_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7548_y0);
  and_gate and_gate_h_u_cla32_and7549_y0(h_u_cla32_and7548_y0, h_u_cla32_and7547_y0, h_u_cla32_and7549_y0);
  and_gate and_gate_h_u_cla32_and7550_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7550_y0);
  and_gate and_gate_h_u_cla32_and7551_y0(h_u_cla32_and7550_y0, h_u_cla32_and7549_y0, h_u_cla32_and7551_y0);
  and_gate and_gate_h_u_cla32_and7552_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7552_y0);
  and_gate and_gate_h_u_cla32_and7553_y0(h_u_cla32_and7552_y0, h_u_cla32_and7551_y0, h_u_cla32_and7553_y0);
  and_gate and_gate_h_u_cla32_and7554_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7554_y0);
  and_gate and_gate_h_u_cla32_and7555_y0(h_u_cla32_and7554_y0, h_u_cla32_and7553_y0, h_u_cla32_and7555_y0);
  and_gate and_gate_h_u_cla32_and7556_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7556_y0);
  and_gate and_gate_h_u_cla32_and7557_y0(h_u_cla32_and7556_y0, h_u_cla32_and7555_y0, h_u_cla32_and7557_y0);
  and_gate and_gate_h_u_cla32_and7558_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7558_y0);
  and_gate and_gate_h_u_cla32_and7559_y0(h_u_cla32_and7558_y0, h_u_cla32_and7557_y0, h_u_cla32_and7559_y0);
  and_gate and_gate_h_u_cla32_and7560_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7560_y0);
  and_gate and_gate_h_u_cla32_and7561_y0(h_u_cla32_and7560_y0, h_u_cla32_and7559_y0, h_u_cla32_and7561_y0);
  and_gate and_gate_h_u_cla32_and7562_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7562_y0);
  and_gate and_gate_h_u_cla32_and7563_y0(h_u_cla32_and7562_y0, h_u_cla32_and7561_y0, h_u_cla32_and7563_y0);
  and_gate and_gate_h_u_cla32_and7564_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7564_y0);
  and_gate and_gate_h_u_cla32_and7565_y0(h_u_cla32_and7564_y0, h_u_cla32_and7563_y0, h_u_cla32_and7565_y0);
  and_gate and_gate_h_u_cla32_and7566_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7566_y0);
  and_gate and_gate_h_u_cla32_and7567_y0(h_u_cla32_and7566_y0, h_u_cla32_and7565_y0, h_u_cla32_and7567_y0);
  and_gate and_gate_h_u_cla32_and7568_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and7568_y0);
  and_gate and_gate_h_u_cla32_and7569_y0(h_u_cla32_and7568_y0, h_u_cla32_and7567_y0, h_u_cla32_and7569_y0);
  and_gate and_gate_h_u_cla32_and7570_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7570_y0);
  and_gate and_gate_h_u_cla32_and7571_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7571_y0);
  and_gate and_gate_h_u_cla32_and7572_y0(h_u_cla32_and7571_y0, h_u_cla32_and7570_y0, h_u_cla32_and7572_y0);
  and_gate and_gate_h_u_cla32_and7573_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7573_y0);
  and_gate and_gate_h_u_cla32_and7574_y0(h_u_cla32_and7573_y0, h_u_cla32_and7572_y0, h_u_cla32_and7574_y0);
  and_gate and_gate_h_u_cla32_and7575_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7575_y0);
  and_gate and_gate_h_u_cla32_and7576_y0(h_u_cla32_and7575_y0, h_u_cla32_and7574_y0, h_u_cla32_and7576_y0);
  and_gate and_gate_h_u_cla32_and7577_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7577_y0);
  and_gate and_gate_h_u_cla32_and7578_y0(h_u_cla32_and7577_y0, h_u_cla32_and7576_y0, h_u_cla32_and7578_y0);
  and_gate and_gate_h_u_cla32_and7579_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7579_y0);
  and_gate and_gate_h_u_cla32_and7580_y0(h_u_cla32_and7579_y0, h_u_cla32_and7578_y0, h_u_cla32_and7580_y0);
  and_gate and_gate_h_u_cla32_and7581_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7581_y0);
  and_gate and_gate_h_u_cla32_and7582_y0(h_u_cla32_and7581_y0, h_u_cla32_and7580_y0, h_u_cla32_and7582_y0);
  and_gate and_gate_h_u_cla32_and7583_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7583_y0);
  and_gate and_gate_h_u_cla32_and7584_y0(h_u_cla32_and7583_y0, h_u_cla32_and7582_y0, h_u_cla32_and7584_y0);
  and_gate and_gate_h_u_cla32_and7585_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7585_y0);
  and_gate and_gate_h_u_cla32_and7586_y0(h_u_cla32_and7585_y0, h_u_cla32_and7584_y0, h_u_cla32_and7586_y0);
  and_gate and_gate_h_u_cla32_and7587_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7587_y0);
  and_gate and_gate_h_u_cla32_and7588_y0(h_u_cla32_and7587_y0, h_u_cla32_and7586_y0, h_u_cla32_and7588_y0);
  and_gate and_gate_h_u_cla32_and7589_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7589_y0);
  and_gate and_gate_h_u_cla32_and7590_y0(h_u_cla32_and7589_y0, h_u_cla32_and7588_y0, h_u_cla32_and7590_y0);
  and_gate and_gate_h_u_cla32_and7591_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and7591_y0);
  and_gate and_gate_h_u_cla32_and7592_y0(h_u_cla32_and7591_y0, h_u_cla32_and7590_y0, h_u_cla32_and7592_y0);
  and_gate and_gate_h_u_cla32_and7593_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7593_y0);
  and_gate and_gate_h_u_cla32_and7594_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7594_y0);
  and_gate and_gate_h_u_cla32_and7595_y0(h_u_cla32_and7594_y0, h_u_cla32_and7593_y0, h_u_cla32_and7595_y0);
  and_gate and_gate_h_u_cla32_and7596_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7596_y0);
  and_gate and_gate_h_u_cla32_and7597_y0(h_u_cla32_and7596_y0, h_u_cla32_and7595_y0, h_u_cla32_and7597_y0);
  and_gate and_gate_h_u_cla32_and7598_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7598_y0);
  and_gate and_gate_h_u_cla32_and7599_y0(h_u_cla32_and7598_y0, h_u_cla32_and7597_y0, h_u_cla32_and7599_y0);
  and_gate and_gate_h_u_cla32_and7600_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7600_y0);
  and_gate and_gate_h_u_cla32_and7601_y0(h_u_cla32_and7600_y0, h_u_cla32_and7599_y0, h_u_cla32_and7601_y0);
  and_gate and_gate_h_u_cla32_and7602_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7602_y0);
  and_gate and_gate_h_u_cla32_and7603_y0(h_u_cla32_and7602_y0, h_u_cla32_and7601_y0, h_u_cla32_and7603_y0);
  and_gate and_gate_h_u_cla32_and7604_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7604_y0);
  and_gate and_gate_h_u_cla32_and7605_y0(h_u_cla32_and7604_y0, h_u_cla32_and7603_y0, h_u_cla32_and7605_y0);
  and_gate and_gate_h_u_cla32_and7606_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7606_y0);
  and_gate and_gate_h_u_cla32_and7607_y0(h_u_cla32_and7606_y0, h_u_cla32_and7605_y0, h_u_cla32_and7607_y0);
  and_gate and_gate_h_u_cla32_and7608_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7608_y0);
  and_gate and_gate_h_u_cla32_and7609_y0(h_u_cla32_and7608_y0, h_u_cla32_and7607_y0, h_u_cla32_and7609_y0);
  and_gate and_gate_h_u_cla32_and7610_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7610_y0);
  and_gate and_gate_h_u_cla32_and7611_y0(h_u_cla32_and7610_y0, h_u_cla32_and7609_y0, h_u_cla32_and7611_y0);
  and_gate and_gate_h_u_cla32_and7612_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and7612_y0);
  and_gate and_gate_h_u_cla32_and7613_y0(h_u_cla32_and7612_y0, h_u_cla32_and7611_y0, h_u_cla32_and7613_y0);
  and_gate and_gate_h_u_cla32_and7614_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7614_y0);
  and_gate and_gate_h_u_cla32_and7615_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7615_y0);
  and_gate and_gate_h_u_cla32_and7616_y0(h_u_cla32_and7615_y0, h_u_cla32_and7614_y0, h_u_cla32_and7616_y0);
  and_gate and_gate_h_u_cla32_and7617_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7617_y0);
  and_gate and_gate_h_u_cla32_and7618_y0(h_u_cla32_and7617_y0, h_u_cla32_and7616_y0, h_u_cla32_and7618_y0);
  and_gate and_gate_h_u_cla32_and7619_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7619_y0);
  and_gate and_gate_h_u_cla32_and7620_y0(h_u_cla32_and7619_y0, h_u_cla32_and7618_y0, h_u_cla32_and7620_y0);
  and_gate and_gate_h_u_cla32_and7621_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7621_y0);
  and_gate and_gate_h_u_cla32_and7622_y0(h_u_cla32_and7621_y0, h_u_cla32_and7620_y0, h_u_cla32_and7622_y0);
  and_gate and_gate_h_u_cla32_and7623_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7623_y0);
  and_gate and_gate_h_u_cla32_and7624_y0(h_u_cla32_and7623_y0, h_u_cla32_and7622_y0, h_u_cla32_and7624_y0);
  and_gate and_gate_h_u_cla32_and7625_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7625_y0);
  and_gate and_gate_h_u_cla32_and7626_y0(h_u_cla32_and7625_y0, h_u_cla32_and7624_y0, h_u_cla32_and7626_y0);
  and_gate and_gate_h_u_cla32_and7627_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7627_y0);
  and_gate and_gate_h_u_cla32_and7628_y0(h_u_cla32_and7627_y0, h_u_cla32_and7626_y0, h_u_cla32_and7628_y0);
  and_gate and_gate_h_u_cla32_and7629_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7629_y0);
  and_gate and_gate_h_u_cla32_and7630_y0(h_u_cla32_and7629_y0, h_u_cla32_and7628_y0, h_u_cla32_and7630_y0);
  and_gate and_gate_h_u_cla32_and7631_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and7631_y0);
  and_gate and_gate_h_u_cla32_and7632_y0(h_u_cla32_and7631_y0, h_u_cla32_and7630_y0, h_u_cla32_and7632_y0);
  and_gate and_gate_h_u_cla32_and7633_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7633_y0);
  and_gate and_gate_h_u_cla32_and7634_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7634_y0);
  and_gate and_gate_h_u_cla32_and7635_y0(h_u_cla32_and7634_y0, h_u_cla32_and7633_y0, h_u_cla32_and7635_y0);
  and_gate and_gate_h_u_cla32_and7636_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7636_y0);
  and_gate and_gate_h_u_cla32_and7637_y0(h_u_cla32_and7636_y0, h_u_cla32_and7635_y0, h_u_cla32_and7637_y0);
  and_gate and_gate_h_u_cla32_and7638_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7638_y0);
  and_gate and_gate_h_u_cla32_and7639_y0(h_u_cla32_and7638_y0, h_u_cla32_and7637_y0, h_u_cla32_and7639_y0);
  and_gate and_gate_h_u_cla32_and7640_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7640_y0);
  and_gate and_gate_h_u_cla32_and7641_y0(h_u_cla32_and7640_y0, h_u_cla32_and7639_y0, h_u_cla32_and7641_y0);
  and_gate and_gate_h_u_cla32_and7642_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7642_y0);
  and_gate and_gate_h_u_cla32_and7643_y0(h_u_cla32_and7642_y0, h_u_cla32_and7641_y0, h_u_cla32_and7643_y0);
  and_gate and_gate_h_u_cla32_and7644_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7644_y0);
  and_gate and_gate_h_u_cla32_and7645_y0(h_u_cla32_and7644_y0, h_u_cla32_and7643_y0, h_u_cla32_and7645_y0);
  and_gate and_gate_h_u_cla32_and7646_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7646_y0);
  and_gate and_gate_h_u_cla32_and7647_y0(h_u_cla32_and7646_y0, h_u_cla32_and7645_y0, h_u_cla32_and7647_y0);
  and_gate and_gate_h_u_cla32_and7648_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and7648_y0);
  and_gate and_gate_h_u_cla32_and7649_y0(h_u_cla32_and7648_y0, h_u_cla32_and7647_y0, h_u_cla32_and7649_y0);
  and_gate and_gate_h_u_cla32_and7650_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7650_y0);
  and_gate and_gate_h_u_cla32_and7651_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7651_y0);
  and_gate and_gate_h_u_cla32_and7652_y0(h_u_cla32_and7651_y0, h_u_cla32_and7650_y0, h_u_cla32_and7652_y0);
  and_gate and_gate_h_u_cla32_and7653_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7653_y0);
  and_gate and_gate_h_u_cla32_and7654_y0(h_u_cla32_and7653_y0, h_u_cla32_and7652_y0, h_u_cla32_and7654_y0);
  and_gate and_gate_h_u_cla32_and7655_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7655_y0);
  and_gate and_gate_h_u_cla32_and7656_y0(h_u_cla32_and7655_y0, h_u_cla32_and7654_y0, h_u_cla32_and7656_y0);
  and_gate and_gate_h_u_cla32_and7657_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7657_y0);
  and_gate and_gate_h_u_cla32_and7658_y0(h_u_cla32_and7657_y0, h_u_cla32_and7656_y0, h_u_cla32_and7658_y0);
  and_gate and_gate_h_u_cla32_and7659_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7659_y0);
  and_gate and_gate_h_u_cla32_and7660_y0(h_u_cla32_and7659_y0, h_u_cla32_and7658_y0, h_u_cla32_and7660_y0);
  and_gate and_gate_h_u_cla32_and7661_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7661_y0);
  and_gate and_gate_h_u_cla32_and7662_y0(h_u_cla32_and7661_y0, h_u_cla32_and7660_y0, h_u_cla32_and7662_y0);
  and_gate and_gate_h_u_cla32_and7663_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and7663_y0);
  and_gate and_gate_h_u_cla32_and7664_y0(h_u_cla32_and7663_y0, h_u_cla32_and7662_y0, h_u_cla32_and7664_y0);
  and_gate and_gate_h_u_cla32_and7665_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7665_y0);
  and_gate and_gate_h_u_cla32_and7666_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7666_y0);
  and_gate and_gate_h_u_cla32_and7667_y0(h_u_cla32_and7666_y0, h_u_cla32_and7665_y0, h_u_cla32_and7667_y0);
  and_gate and_gate_h_u_cla32_and7668_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7668_y0);
  and_gate and_gate_h_u_cla32_and7669_y0(h_u_cla32_and7668_y0, h_u_cla32_and7667_y0, h_u_cla32_and7669_y0);
  and_gate and_gate_h_u_cla32_and7670_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7670_y0);
  and_gate and_gate_h_u_cla32_and7671_y0(h_u_cla32_and7670_y0, h_u_cla32_and7669_y0, h_u_cla32_and7671_y0);
  and_gate and_gate_h_u_cla32_and7672_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7672_y0);
  and_gate and_gate_h_u_cla32_and7673_y0(h_u_cla32_and7672_y0, h_u_cla32_and7671_y0, h_u_cla32_and7673_y0);
  and_gate and_gate_h_u_cla32_and7674_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7674_y0);
  and_gate and_gate_h_u_cla32_and7675_y0(h_u_cla32_and7674_y0, h_u_cla32_and7673_y0, h_u_cla32_and7675_y0);
  and_gate and_gate_h_u_cla32_and7676_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and7676_y0);
  and_gate and_gate_h_u_cla32_and7677_y0(h_u_cla32_and7676_y0, h_u_cla32_and7675_y0, h_u_cla32_and7677_y0);
  and_gate and_gate_h_u_cla32_and7678_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and7678_y0);
  and_gate and_gate_h_u_cla32_and7679_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and7679_y0);
  and_gate and_gate_h_u_cla32_and7680_y0(h_u_cla32_and7679_y0, h_u_cla32_and7678_y0, h_u_cla32_and7680_y0);
  and_gate and_gate_h_u_cla32_and7681_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and7681_y0);
  and_gate and_gate_h_u_cla32_and7682_y0(h_u_cla32_and7681_y0, h_u_cla32_and7680_y0, h_u_cla32_and7682_y0);
  and_gate and_gate_h_u_cla32_and7683_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and7683_y0);
  and_gate and_gate_h_u_cla32_and7684_y0(h_u_cla32_and7683_y0, h_u_cla32_and7682_y0, h_u_cla32_and7684_y0);
  and_gate and_gate_h_u_cla32_and7685_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and7685_y0);
  and_gate and_gate_h_u_cla32_and7686_y0(h_u_cla32_and7685_y0, h_u_cla32_and7684_y0, h_u_cla32_and7686_y0);
  and_gate and_gate_h_u_cla32_and7687_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and7687_y0);
  and_gate and_gate_h_u_cla32_and7688_y0(h_u_cla32_and7687_y0, h_u_cla32_and7686_y0, h_u_cla32_and7688_y0);
  and_gate and_gate_h_u_cla32_and7689_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and7689_y0);
  and_gate and_gate_h_u_cla32_and7690_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and7690_y0);
  and_gate and_gate_h_u_cla32_and7691_y0(h_u_cla32_and7690_y0, h_u_cla32_and7689_y0, h_u_cla32_and7691_y0);
  and_gate and_gate_h_u_cla32_and7692_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and7692_y0);
  and_gate and_gate_h_u_cla32_and7693_y0(h_u_cla32_and7692_y0, h_u_cla32_and7691_y0, h_u_cla32_and7693_y0);
  and_gate and_gate_h_u_cla32_and7694_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and7694_y0);
  and_gate and_gate_h_u_cla32_and7695_y0(h_u_cla32_and7694_y0, h_u_cla32_and7693_y0, h_u_cla32_and7695_y0);
  and_gate and_gate_h_u_cla32_and7696_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and7696_y0);
  and_gate and_gate_h_u_cla32_and7697_y0(h_u_cla32_and7696_y0, h_u_cla32_and7695_y0, h_u_cla32_and7697_y0);
  and_gate and_gate_h_u_cla32_and7698_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and7698_y0);
  and_gate and_gate_h_u_cla32_and7699_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and7699_y0);
  and_gate and_gate_h_u_cla32_and7700_y0(h_u_cla32_and7699_y0, h_u_cla32_and7698_y0, h_u_cla32_and7700_y0);
  and_gate and_gate_h_u_cla32_and7701_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and7701_y0);
  and_gate and_gate_h_u_cla32_and7702_y0(h_u_cla32_and7701_y0, h_u_cla32_and7700_y0, h_u_cla32_and7702_y0);
  and_gate and_gate_h_u_cla32_and7703_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and7703_y0);
  and_gate and_gate_h_u_cla32_and7704_y0(h_u_cla32_and7703_y0, h_u_cla32_and7702_y0, h_u_cla32_and7704_y0);
  and_gate and_gate_h_u_cla32_and7705_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and7705_y0);
  and_gate and_gate_h_u_cla32_and7706_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and7706_y0);
  and_gate and_gate_h_u_cla32_and7707_y0(h_u_cla32_and7706_y0, h_u_cla32_and7705_y0, h_u_cla32_and7707_y0);
  and_gate and_gate_h_u_cla32_and7708_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and7708_y0);
  and_gate and_gate_h_u_cla32_and7709_y0(h_u_cla32_and7708_y0, h_u_cla32_and7707_y0, h_u_cla32_and7709_y0);
  and_gate and_gate_h_u_cla32_and7710_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and7710_y0);
  and_gate and_gate_h_u_cla32_and7711_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and7711_y0);
  and_gate and_gate_h_u_cla32_and7712_y0(h_u_cla32_and7711_y0, h_u_cla32_and7710_y0, h_u_cla32_and7712_y0);
  and_gate and_gate_h_u_cla32_and7713_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and7713_y0);
  or_gate or_gate_h_u_cla32_or378_y0(h_u_cla32_and7713_y0, h_u_cla32_and6984_y0, h_u_cla32_or378_y0);
  or_gate or_gate_h_u_cla32_or379_y0(h_u_cla32_or378_y0, h_u_cla32_and7037_y0, h_u_cla32_or379_y0);
  or_gate or_gate_h_u_cla32_or380_y0(h_u_cla32_or379_y0, h_u_cla32_and7088_y0, h_u_cla32_or380_y0);
  or_gate or_gate_h_u_cla32_or381_y0(h_u_cla32_or380_y0, h_u_cla32_and7137_y0, h_u_cla32_or381_y0);
  or_gate or_gate_h_u_cla32_or382_y0(h_u_cla32_or381_y0, h_u_cla32_and7184_y0, h_u_cla32_or382_y0);
  or_gate or_gate_h_u_cla32_or383_y0(h_u_cla32_or382_y0, h_u_cla32_and7229_y0, h_u_cla32_or383_y0);
  or_gate or_gate_h_u_cla32_or384_y0(h_u_cla32_or383_y0, h_u_cla32_and7272_y0, h_u_cla32_or384_y0);
  or_gate or_gate_h_u_cla32_or385_y0(h_u_cla32_or384_y0, h_u_cla32_and7313_y0, h_u_cla32_or385_y0);
  or_gate or_gate_h_u_cla32_or386_y0(h_u_cla32_or385_y0, h_u_cla32_and7352_y0, h_u_cla32_or386_y0);
  or_gate or_gate_h_u_cla32_or387_y0(h_u_cla32_or386_y0, h_u_cla32_and7389_y0, h_u_cla32_or387_y0);
  or_gate or_gate_h_u_cla32_or388_y0(h_u_cla32_or387_y0, h_u_cla32_and7424_y0, h_u_cla32_or388_y0);
  or_gate or_gate_h_u_cla32_or389_y0(h_u_cla32_or388_y0, h_u_cla32_and7457_y0, h_u_cla32_or389_y0);
  or_gate or_gate_h_u_cla32_or390_y0(h_u_cla32_or389_y0, h_u_cla32_and7488_y0, h_u_cla32_or390_y0);
  or_gate or_gate_h_u_cla32_or391_y0(h_u_cla32_or390_y0, h_u_cla32_and7517_y0, h_u_cla32_or391_y0);
  or_gate or_gate_h_u_cla32_or392_y0(h_u_cla32_or391_y0, h_u_cla32_and7544_y0, h_u_cla32_or392_y0);
  or_gate or_gate_h_u_cla32_or393_y0(h_u_cla32_or392_y0, h_u_cla32_and7569_y0, h_u_cla32_or393_y0);
  or_gate or_gate_h_u_cla32_or394_y0(h_u_cla32_or393_y0, h_u_cla32_and7592_y0, h_u_cla32_or394_y0);
  or_gate or_gate_h_u_cla32_or395_y0(h_u_cla32_or394_y0, h_u_cla32_and7613_y0, h_u_cla32_or395_y0);
  or_gate or_gate_h_u_cla32_or396_y0(h_u_cla32_or395_y0, h_u_cla32_and7632_y0, h_u_cla32_or396_y0);
  or_gate or_gate_h_u_cla32_or397_y0(h_u_cla32_or396_y0, h_u_cla32_and7649_y0, h_u_cla32_or397_y0);
  or_gate or_gate_h_u_cla32_or398_y0(h_u_cla32_or397_y0, h_u_cla32_and7664_y0, h_u_cla32_or398_y0);
  or_gate or_gate_h_u_cla32_or399_y0(h_u_cla32_or398_y0, h_u_cla32_and7677_y0, h_u_cla32_or399_y0);
  or_gate or_gate_h_u_cla32_or400_y0(h_u_cla32_or399_y0, h_u_cla32_and7688_y0, h_u_cla32_or400_y0);
  or_gate or_gate_h_u_cla32_or401_y0(h_u_cla32_or400_y0, h_u_cla32_and7697_y0, h_u_cla32_or401_y0);
  or_gate or_gate_h_u_cla32_or402_y0(h_u_cla32_or401_y0, h_u_cla32_and7704_y0, h_u_cla32_or402_y0);
  or_gate or_gate_h_u_cla32_or403_y0(h_u_cla32_or402_y0, h_u_cla32_and7709_y0, h_u_cla32_or403_y0);
  or_gate or_gate_h_u_cla32_or404_y0(h_u_cla32_or403_y0, h_u_cla32_and7712_y0, h_u_cla32_or404_y0);
  or_gate or_gate_h_u_cla32_or405_y0(h_u_cla32_pg_logic27_y1, h_u_cla32_or404_y0, h_u_cla32_or405_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic28_y0(a_28, b_28, h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_pg_logic28_y2);
  xor_gate xor_gate_h_u_cla32_xor28_y0(h_u_cla32_pg_logic28_y2, h_u_cla32_or405_y0, h_u_cla32_xor28_y0);
  and_gate and_gate_h_u_cla32_and7714_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and7714_y0);
  and_gate and_gate_h_u_cla32_and7715_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and7715_y0);
  and_gate and_gate_h_u_cla32_and7716_y0(h_u_cla32_and7715_y0, h_u_cla32_and7714_y0, h_u_cla32_and7716_y0);
  and_gate and_gate_h_u_cla32_and7717_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and7717_y0);
  and_gate and_gate_h_u_cla32_and7718_y0(h_u_cla32_and7717_y0, h_u_cla32_and7716_y0, h_u_cla32_and7718_y0);
  and_gate and_gate_h_u_cla32_and7719_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and7719_y0);
  and_gate and_gate_h_u_cla32_and7720_y0(h_u_cla32_and7719_y0, h_u_cla32_and7718_y0, h_u_cla32_and7720_y0);
  and_gate and_gate_h_u_cla32_and7721_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and7721_y0);
  and_gate and_gate_h_u_cla32_and7722_y0(h_u_cla32_and7721_y0, h_u_cla32_and7720_y0, h_u_cla32_and7722_y0);
  and_gate and_gate_h_u_cla32_and7723_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and7723_y0);
  and_gate and_gate_h_u_cla32_and7724_y0(h_u_cla32_and7723_y0, h_u_cla32_and7722_y0, h_u_cla32_and7724_y0);
  and_gate and_gate_h_u_cla32_and7725_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and7725_y0);
  and_gate and_gate_h_u_cla32_and7726_y0(h_u_cla32_and7725_y0, h_u_cla32_and7724_y0, h_u_cla32_and7726_y0);
  and_gate and_gate_h_u_cla32_and7727_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and7727_y0);
  and_gate and_gate_h_u_cla32_and7728_y0(h_u_cla32_and7727_y0, h_u_cla32_and7726_y0, h_u_cla32_and7728_y0);
  and_gate and_gate_h_u_cla32_and7729_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and7729_y0);
  and_gate and_gate_h_u_cla32_and7730_y0(h_u_cla32_and7729_y0, h_u_cla32_and7728_y0, h_u_cla32_and7730_y0);
  and_gate and_gate_h_u_cla32_and7731_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and7731_y0);
  and_gate and_gate_h_u_cla32_and7732_y0(h_u_cla32_and7731_y0, h_u_cla32_and7730_y0, h_u_cla32_and7732_y0);
  and_gate and_gate_h_u_cla32_and7733_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and7733_y0);
  and_gate and_gate_h_u_cla32_and7734_y0(h_u_cla32_and7733_y0, h_u_cla32_and7732_y0, h_u_cla32_and7734_y0);
  and_gate and_gate_h_u_cla32_and7735_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and7735_y0);
  and_gate and_gate_h_u_cla32_and7736_y0(h_u_cla32_and7735_y0, h_u_cla32_and7734_y0, h_u_cla32_and7736_y0);
  and_gate and_gate_h_u_cla32_and7737_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and7737_y0);
  and_gate and_gate_h_u_cla32_and7738_y0(h_u_cla32_and7737_y0, h_u_cla32_and7736_y0, h_u_cla32_and7738_y0);
  and_gate and_gate_h_u_cla32_and7739_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and7739_y0);
  and_gate and_gate_h_u_cla32_and7740_y0(h_u_cla32_and7739_y0, h_u_cla32_and7738_y0, h_u_cla32_and7740_y0);
  and_gate and_gate_h_u_cla32_and7741_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and7741_y0);
  and_gate and_gate_h_u_cla32_and7742_y0(h_u_cla32_and7741_y0, h_u_cla32_and7740_y0, h_u_cla32_and7742_y0);
  and_gate and_gate_h_u_cla32_and7743_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and7743_y0);
  and_gate and_gate_h_u_cla32_and7744_y0(h_u_cla32_and7743_y0, h_u_cla32_and7742_y0, h_u_cla32_and7744_y0);
  and_gate and_gate_h_u_cla32_and7745_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and7745_y0);
  and_gate and_gate_h_u_cla32_and7746_y0(h_u_cla32_and7745_y0, h_u_cla32_and7744_y0, h_u_cla32_and7746_y0);
  and_gate and_gate_h_u_cla32_and7747_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and7747_y0);
  and_gate and_gate_h_u_cla32_and7748_y0(h_u_cla32_and7747_y0, h_u_cla32_and7746_y0, h_u_cla32_and7748_y0);
  and_gate and_gate_h_u_cla32_and7749_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and7749_y0);
  and_gate and_gate_h_u_cla32_and7750_y0(h_u_cla32_and7749_y0, h_u_cla32_and7748_y0, h_u_cla32_and7750_y0);
  and_gate and_gate_h_u_cla32_and7751_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and7751_y0);
  and_gate and_gate_h_u_cla32_and7752_y0(h_u_cla32_and7751_y0, h_u_cla32_and7750_y0, h_u_cla32_and7752_y0);
  and_gate and_gate_h_u_cla32_and7753_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and7753_y0);
  and_gate and_gate_h_u_cla32_and7754_y0(h_u_cla32_and7753_y0, h_u_cla32_and7752_y0, h_u_cla32_and7754_y0);
  and_gate and_gate_h_u_cla32_and7755_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and7755_y0);
  and_gate and_gate_h_u_cla32_and7756_y0(h_u_cla32_and7755_y0, h_u_cla32_and7754_y0, h_u_cla32_and7756_y0);
  and_gate and_gate_h_u_cla32_and7757_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and7757_y0);
  and_gate and_gate_h_u_cla32_and7758_y0(h_u_cla32_and7757_y0, h_u_cla32_and7756_y0, h_u_cla32_and7758_y0);
  and_gate and_gate_h_u_cla32_and7759_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and7759_y0);
  and_gate and_gate_h_u_cla32_and7760_y0(h_u_cla32_and7759_y0, h_u_cla32_and7758_y0, h_u_cla32_and7760_y0);
  and_gate and_gate_h_u_cla32_and7761_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and7761_y0);
  and_gate and_gate_h_u_cla32_and7762_y0(h_u_cla32_and7761_y0, h_u_cla32_and7760_y0, h_u_cla32_and7762_y0);
  and_gate and_gate_h_u_cla32_and7763_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and7763_y0);
  and_gate and_gate_h_u_cla32_and7764_y0(h_u_cla32_and7763_y0, h_u_cla32_and7762_y0, h_u_cla32_and7764_y0);
  and_gate and_gate_h_u_cla32_and7765_y0(h_u_cla32_pg_logic26_y0, constant_wire_0, h_u_cla32_and7765_y0);
  and_gate and_gate_h_u_cla32_and7766_y0(h_u_cla32_and7765_y0, h_u_cla32_and7764_y0, h_u_cla32_and7766_y0);
  and_gate and_gate_h_u_cla32_and7767_y0(h_u_cla32_pg_logic27_y0, constant_wire_0, h_u_cla32_and7767_y0);
  and_gate and_gate_h_u_cla32_and7768_y0(h_u_cla32_and7767_y0, h_u_cla32_and7766_y0, h_u_cla32_and7768_y0);
  and_gate and_gate_h_u_cla32_and7769_y0(h_u_cla32_pg_logic28_y0, constant_wire_0, h_u_cla32_and7769_y0);
  and_gate and_gate_h_u_cla32_and7770_y0(h_u_cla32_and7769_y0, h_u_cla32_and7768_y0, h_u_cla32_and7770_y0);
  and_gate and_gate_h_u_cla32_and7771_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7771_y0);
  and_gate and_gate_h_u_cla32_and7772_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7772_y0);
  and_gate and_gate_h_u_cla32_and7773_y0(h_u_cla32_and7772_y0, h_u_cla32_and7771_y0, h_u_cla32_and7773_y0);
  and_gate and_gate_h_u_cla32_and7774_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7774_y0);
  and_gate and_gate_h_u_cla32_and7775_y0(h_u_cla32_and7774_y0, h_u_cla32_and7773_y0, h_u_cla32_and7775_y0);
  and_gate and_gate_h_u_cla32_and7776_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7776_y0);
  and_gate and_gate_h_u_cla32_and7777_y0(h_u_cla32_and7776_y0, h_u_cla32_and7775_y0, h_u_cla32_and7777_y0);
  and_gate and_gate_h_u_cla32_and7778_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7778_y0);
  and_gate and_gate_h_u_cla32_and7779_y0(h_u_cla32_and7778_y0, h_u_cla32_and7777_y0, h_u_cla32_and7779_y0);
  and_gate and_gate_h_u_cla32_and7780_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7780_y0);
  and_gate and_gate_h_u_cla32_and7781_y0(h_u_cla32_and7780_y0, h_u_cla32_and7779_y0, h_u_cla32_and7781_y0);
  and_gate and_gate_h_u_cla32_and7782_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7782_y0);
  and_gate and_gate_h_u_cla32_and7783_y0(h_u_cla32_and7782_y0, h_u_cla32_and7781_y0, h_u_cla32_and7783_y0);
  and_gate and_gate_h_u_cla32_and7784_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7784_y0);
  and_gate and_gate_h_u_cla32_and7785_y0(h_u_cla32_and7784_y0, h_u_cla32_and7783_y0, h_u_cla32_and7785_y0);
  and_gate and_gate_h_u_cla32_and7786_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7786_y0);
  and_gate and_gate_h_u_cla32_and7787_y0(h_u_cla32_and7786_y0, h_u_cla32_and7785_y0, h_u_cla32_and7787_y0);
  and_gate and_gate_h_u_cla32_and7788_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7788_y0);
  and_gate and_gate_h_u_cla32_and7789_y0(h_u_cla32_and7788_y0, h_u_cla32_and7787_y0, h_u_cla32_and7789_y0);
  and_gate and_gate_h_u_cla32_and7790_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7790_y0);
  and_gate and_gate_h_u_cla32_and7791_y0(h_u_cla32_and7790_y0, h_u_cla32_and7789_y0, h_u_cla32_and7791_y0);
  and_gate and_gate_h_u_cla32_and7792_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7792_y0);
  and_gate and_gate_h_u_cla32_and7793_y0(h_u_cla32_and7792_y0, h_u_cla32_and7791_y0, h_u_cla32_and7793_y0);
  and_gate and_gate_h_u_cla32_and7794_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7794_y0);
  and_gate and_gate_h_u_cla32_and7795_y0(h_u_cla32_and7794_y0, h_u_cla32_and7793_y0, h_u_cla32_and7795_y0);
  and_gate and_gate_h_u_cla32_and7796_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7796_y0);
  and_gate and_gate_h_u_cla32_and7797_y0(h_u_cla32_and7796_y0, h_u_cla32_and7795_y0, h_u_cla32_and7797_y0);
  and_gate and_gate_h_u_cla32_and7798_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7798_y0);
  and_gate and_gate_h_u_cla32_and7799_y0(h_u_cla32_and7798_y0, h_u_cla32_and7797_y0, h_u_cla32_and7799_y0);
  and_gate and_gate_h_u_cla32_and7800_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7800_y0);
  and_gate and_gate_h_u_cla32_and7801_y0(h_u_cla32_and7800_y0, h_u_cla32_and7799_y0, h_u_cla32_and7801_y0);
  and_gate and_gate_h_u_cla32_and7802_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7802_y0);
  and_gate and_gate_h_u_cla32_and7803_y0(h_u_cla32_and7802_y0, h_u_cla32_and7801_y0, h_u_cla32_and7803_y0);
  and_gate and_gate_h_u_cla32_and7804_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7804_y0);
  and_gate and_gate_h_u_cla32_and7805_y0(h_u_cla32_and7804_y0, h_u_cla32_and7803_y0, h_u_cla32_and7805_y0);
  and_gate and_gate_h_u_cla32_and7806_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7806_y0);
  and_gate and_gate_h_u_cla32_and7807_y0(h_u_cla32_and7806_y0, h_u_cla32_and7805_y0, h_u_cla32_and7807_y0);
  and_gate and_gate_h_u_cla32_and7808_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7808_y0);
  and_gate and_gate_h_u_cla32_and7809_y0(h_u_cla32_and7808_y0, h_u_cla32_and7807_y0, h_u_cla32_and7809_y0);
  and_gate and_gate_h_u_cla32_and7810_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7810_y0);
  and_gate and_gate_h_u_cla32_and7811_y0(h_u_cla32_and7810_y0, h_u_cla32_and7809_y0, h_u_cla32_and7811_y0);
  and_gate and_gate_h_u_cla32_and7812_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7812_y0);
  and_gate and_gate_h_u_cla32_and7813_y0(h_u_cla32_and7812_y0, h_u_cla32_and7811_y0, h_u_cla32_and7813_y0);
  and_gate and_gate_h_u_cla32_and7814_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7814_y0);
  and_gate and_gate_h_u_cla32_and7815_y0(h_u_cla32_and7814_y0, h_u_cla32_and7813_y0, h_u_cla32_and7815_y0);
  and_gate and_gate_h_u_cla32_and7816_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7816_y0);
  and_gate and_gate_h_u_cla32_and7817_y0(h_u_cla32_and7816_y0, h_u_cla32_and7815_y0, h_u_cla32_and7817_y0);
  and_gate and_gate_h_u_cla32_and7818_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7818_y0);
  and_gate and_gate_h_u_cla32_and7819_y0(h_u_cla32_and7818_y0, h_u_cla32_and7817_y0, h_u_cla32_and7819_y0);
  and_gate and_gate_h_u_cla32_and7820_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7820_y0);
  and_gate and_gate_h_u_cla32_and7821_y0(h_u_cla32_and7820_y0, h_u_cla32_and7819_y0, h_u_cla32_and7821_y0);
  and_gate and_gate_h_u_cla32_and7822_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7822_y0);
  and_gate and_gate_h_u_cla32_and7823_y0(h_u_cla32_and7822_y0, h_u_cla32_and7821_y0, h_u_cla32_and7823_y0);
  and_gate and_gate_h_u_cla32_and7824_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and7824_y0);
  and_gate and_gate_h_u_cla32_and7825_y0(h_u_cla32_and7824_y0, h_u_cla32_and7823_y0, h_u_cla32_and7825_y0);
  and_gate and_gate_h_u_cla32_and7826_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7826_y0);
  and_gate and_gate_h_u_cla32_and7827_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7827_y0);
  and_gate and_gate_h_u_cla32_and7828_y0(h_u_cla32_and7827_y0, h_u_cla32_and7826_y0, h_u_cla32_and7828_y0);
  and_gate and_gate_h_u_cla32_and7829_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7829_y0);
  and_gate and_gate_h_u_cla32_and7830_y0(h_u_cla32_and7829_y0, h_u_cla32_and7828_y0, h_u_cla32_and7830_y0);
  and_gate and_gate_h_u_cla32_and7831_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7831_y0);
  and_gate and_gate_h_u_cla32_and7832_y0(h_u_cla32_and7831_y0, h_u_cla32_and7830_y0, h_u_cla32_and7832_y0);
  and_gate and_gate_h_u_cla32_and7833_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7833_y0);
  and_gate and_gate_h_u_cla32_and7834_y0(h_u_cla32_and7833_y0, h_u_cla32_and7832_y0, h_u_cla32_and7834_y0);
  and_gate and_gate_h_u_cla32_and7835_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7835_y0);
  and_gate and_gate_h_u_cla32_and7836_y0(h_u_cla32_and7835_y0, h_u_cla32_and7834_y0, h_u_cla32_and7836_y0);
  and_gate and_gate_h_u_cla32_and7837_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7837_y0);
  and_gate and_gate_h_u_cla32_and7838_y0(h_u_cla32_and7837_y0, h_u_cla32_and7836_y0, h_u_cla32_and7838_y0);
  and_gate and_gate_h_u_cla32_and7839_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7839_y0);
  and_gate and_gate_h_u_cla32_and7840_y0(h_u_cla32_and7839_y0, h_u_cla32_and7838_y0, h_u_cla32_and7840_y0);
  and_gate and_gate_h_u_cla32_and7841_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7841_y0);
  and_gate and_gate_h_u_cla32_and7842_y0(h_u_cla32_and7841_y0, h_u_cla32_and7840_y0, h_u_cla32_and7842_y0);
  and_gate and_gate_h_u_cla32_and7843_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7843_y0);
  and_gate and_gate_h_u_cla32_and7844_y0(h_u_cla32_and7843_y0, h_u_cla32_and7842_y0, h_u_cla32_and7844_y0);
  and_gate and_gate_h_u_cla32_and7845_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7845_y0);
  and_gate and_gate_h_u_cla32_and7846_y0(h_u_cla32_and7845_y0, h_u_cla32_and7844_y0, h_u_cla32_and7846_y0);
  and_gate and_gate_h_u_cla32_and7847_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7847_y0);
  and_gate and_gate_h_u_cla32_and7848_y0(h_u_cla32_and7847_y0, h_u_cla32_and7846_y0, h_u_cla32_and7848_y0);
  and_gate and_gate_h_u_cla32_and7849_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7849_y0);
  and_gate and_gate_h_u_cla32_and7850_y0(h_u_cla32_and7849_y0, h_u_cla32_and7848_y0, h_u_cla32_and7850_y0);
  and_gate and_gate_h_u_cla32_and7851_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7851_y0);
  and_gate and_gate_h_u_cla32_and7852_y0(h_u_cla32_and7851_y0, h_u_cla32_and7850_y0, h_u_cla32_and7852_y0);
  and_gate and_gate_h_u_cla32_and7853_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7853_y0);
  and_gate and_gate_h_u_cla32_and7854_y0(h_u_cla32_and7853_y0, h_u_cla32_and7852_y0, h_u_cla32_and7854_y0);
  and_gate and_gate_h_u_cla32_and7855_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7855_y0);
  and_gate and_gate_h_u_cla32_and7856_y0(h_u_cla32_and7855_y0, h_u_cla32_and7854_y0, h_u_cla32_and7856_y0);
  and_gate and_gate_h_u_cla32_and7857_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7857_y0);
  and_gate and_gate_h_u_cla32_and7858_y0(h_u_cla32_and7857_y0, h_u_cla32_and7856_y0, h_u_cla32_and7858_y0);
  and_gate and_gate_h_u_cla32_and7859_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7859_y0);
  and_gate and_gate_h_u_cla32_and7860_y0(h_u_cla32_and7859_y0, h_u_cla32_and7858_y0, h_u_cla32_and7860_y0);
  and_gate and_gate_h_u_cla32_and7861_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7861_y0);
  and_gate and_gate_h_u_cla32_and7862_y0(h_u_cla32_and7861_y0, h_u_cla32_and7860_y0, h_u_cla32_and7862_y0);
  and_gate and_gate_h_u_cla32_and7863_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7863_y0);
  and_gate and_gate_h_u_cla32_and7864_y0(h_u_cla32_and7863_y0, h_u_cla32_and7862_y0, h_u_cla32_and7864_y0);
  and_gate and_gate_h_u_cla32_and7865_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7865_y0);
  and_gate and_gate_h_u_cla32_and7866_y0(h_u_cla32_and7865_y0, h_u_cla32_and7864_y0, h_u_cla32_and7866_y0);
  and_gate and_gate_h_u_cla32_and7867_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7867_y0);
  and_gate and_gate_h_u_cla32_and7868_y0(h_u_cla32_and7867_y0, h_u_cla32_and7866_y0, h_u_cla32_and7868_y0);
  and_gate and_gate_h_u_cla32_and7869_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7869_y0);
  and_gate and_gate_h_u_cla32_and7870_y0(h_u_cla32_and7869_y0, h_u_cla32_and7868_y0, h_u_cla32_and7870_y0);
  and_gate and_gate_h_u_cla32_and7871_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7871_y0);
  and_gate and_gate_h_u_cla32_and7872_y0(h_u_cla32_and7871_y0, h_u_cla32_and7870_y0, h_u_cla32_and7872_y0);
  and_gate and_gate_h_u_cla32_and7873_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7873_y0);
  and_gate and_gate_h_u_cla32_and7874_y0(h_u_cla32_and7873_y0, h_u_cla32_and7872_y0, h_u_cla32_and7874_y0);
  and_gate and_gate_h_u_cla32_and7875_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7875_y0);
  and_gate and_gate_h_u_cla32_and7876_y0(h_u_cla32_and7875_y0, h_u_cla32_and7874_y0, h_u_cla32_and7876_y0);
  and_gate and_gate_h_u_cla32_and7877_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and7877_y0);
  and_gate and_gate_h_u_cla32_and7878_y0(h_u_cla32_and7877_y0, h_u_cla32_and7876_y0, h_u_cla32_and7878_y0);
  and_gate and_gate_h_u_cla32_and7879_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7879_y0);
  and_gate and_gate_h_u_cla32_and7880_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7880_y0);
  and_gate and_gate_h_u_cla32_and7881_y0(h_u_cla32_and7880_y0, h_u_cla32_and7879_y0, h_u_cla32_and7881_y0);
  and_gate and_gate_h_u_cla32_and7882_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7882_y0);
  and_gate and_gate_h_u_cla32_and7883_y0(h_u_cla32_and7882_y0, h_u_cla32_and7881_y0, h_u_cla32_and7883_y0);
  and_gate and_gate_h_u_cla32_and7884_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7884_y0);
  and_gate and_gate_h_u_cla32_and7885_y0(h_u_cla32_and7884_y0, h_u_cla32_and7883_y0, h_u_cla32_and7885_y0);
  and_gate and_gate_h_u_cla32_and7886_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7886_y0);
  and_gate and_gate_h_u_cla32_and7887_y0(h_u_cla32_and7886_y0, h_u_cla32_and7885_y0, h_u_cla32_and7887_y0);
  and_gate and_gate_h_u_cla32_and7888_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7888_y0);
  and_gate and_gate_h_u_cla32_and7889_y0(h_u_cla32_and7888_y0, h_u_cla32_and7887_y0, h_u_cla32_and7889_y0);
  and_gate and_gate_h_u_cla32_and7890_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7890_y0);
  and_gate and_gate_h_u_cla32_and7891_y0(h_u_cla32_and7890_y0, h_u_cla32_and7889_y0, h_u_cla32_and7891_y0);
  and_gate and_gate_h_u_cla32_and7892_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7892_y0);
  and_gate and_gate_h_u_cla32_and7893_y0(h_u_cla32_and7892_y0, h_u_cla32_and7891_y0, h_u_cla32_and7893_y0);
  and_gate and_gate_h_u_cla32_and7894_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7894_y0);
  and_gate and_gate_h_u_cla32_and7895_y0(h_u_cla32_and7894_y0, h_u_cla32_and7893_y0, h_u_cla32_and7895_y0);
  and_gate and_gate_h_u_cla32_and7896_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7896_y0);
  and_gate and_gate_h_u_cla32_and7897_y0(h_u_cla32_and7896_y0, h_u_cla32_and7895_y0, h_u_cla32_and7897_y0);
  and_gate and_gate_h_u_cla32_and7898_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7898_y0);
  and_gate and_gate_h_u_cla32_and7899_y0(h_u_cla32_and7898_y0, h_u_cla32_and7897_y0, h_u_cla32_and7899_y0);
  and_gate and_gate_h_u_cla32_and7900_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7900_y0);
  and_gate and_gate_h_u_cla32_and7901_y0(h_u_cla32_and7900_y0, h_u_cla32_and7899_y0, h_u_cla32_and7901_y0);
  and_gate and_gate_h_u_cla32_and7902_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7902_y0);
  and_gate and_gate_h_u_cla32_and7903_y0(h_u_cla32_and7902_y0, h_u_cla32_and7901_y0, h_u_cla32_and7903_y0);
  and_gate and_gate_h_u_cla32_and7904_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7904_y0);
  and_gate and_gate_h_u_cla32_and7905_y0(h_u_cla32_and7904_y0, h_u_cla32_and7903_y0, h_u_cla32_and7905_y0);
  and_gate and_gate_h_u_cla32_and7906_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7906_y0);
  and_gate and_gate_h_u_cla32_and7907_y0(h_u_cla32_and7906_y0, h_u_cla32_and7905_y0, h_u_cla32_and7907_y0);
  and_gate and_gate_h_u_cla32_and7908_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7908_y0);
  and_gate and_gate_h_u_cla32_and7909_y0(h_u_cla32_and7908_y0, h_u_cla32_and7907_y0, h_u_cla32_and7909_y0);
  and_gate and_gate_h_u_cla32_and7910_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7910_y0);
  and_gate and_gate_h_u_cla32_and7911_y0(h_u_cla32_and7910_y0, h_u_cla32_and7909_y0, h_u_cla32_and7911_y0);
  and_gate and_gate_h_u_cla32_and7912_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7912_y0);
  and_gate and_gate_h_u_cla32_and7913_y0(h_u_cla32_and7912_y0, h_u_cla32_and7911_y0, h_u_cla32_and7913_y0);
  and_gate and_gate_h_u_cla32_and7914_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7914_y0);
  and_gate and_gate_h_u_cla32_and7915_y0(h_u_cla32_and7914_y0, h_u_cla32_and7913_y0, h_u_cla32_and7915_y0);
  and_gate and_gate_h_u_cla32_and7916_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7916_y0);
  and_gate and_gate_h_u_cla32_and7917_y0(h_u_cla32_and7916_y0, h_u_cla32_and7915_y0, h_u_cla32_and7917_y0);
  and_gate and_gate_h_u_cla32_and7918_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7918_y0);
  and_gate and_gate_h_u_cla32_and7919_y0(h_u_cla32_and7918_y0, h_u_cla32_and7917_y0, h_u_cla32_and7919_y0);
  and_gate and_gate_h_u_cla32_and7920_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7920_y0);
  and_gate and_gate_h_u_cla32_and7921_y0(h_u_cla32_and7920_y0, h_u_cla32_and7919_y0, h_u_cla32_and7921_y0);
  and_gate and_gate_h_u_cla32_and7922_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7922_y0);
  and_gate and_gate_h_u_cla32_and7923_y0(h_u_cla32_and7922_y0, h_u_cla32_and7921_y0, h_u_cla32_and7923_y0);
  and_gate and_gate_h_u_cla32_and7924_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7924_y0);
  and_gate and_gate_h_u_cla32_and7925_y0(h_u_cla32_and7924_y0, h_u_cla32_and7923_y0, h_u_cla32_and7925_y0);
  and_gate and_gate_h_u_cla32_and7926_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7926_y0);
  and_gate and_gate_h_u_cla32_and7927_y0(h_u_cla32_and7926_y0, h_u_cla32_and7925_y0, h_u_cla32_and7927_y0);
  and_gate and_gate_h_u_cla32_and7928_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and7928_y0);
  and_gate and_gate_h_u_cla32_and7929_y0(h_u_cla32_and7928_y0, h_u_cla32_and7927_y0, h_u_cla32_and7929_y0);
  and_gate and_gate_h_u_cla32_and7930_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7930_y0);
  and_gate and_gate_h_u_cla32_and7931_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7931_y0);
  and_gate and_gate_h_u_cla32_and7932_y0(h_u_cla32_and7931_y0, h_u_cla32_and7930_y0, h_u_cla32_and7932_y0);
  and_gate and_gate_h_u_cla32_and7933_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7933_y0);
  and_gate and_gate_h_u_cla32_and7934_y0(h_u_cla32_and7933_y0, h_u_cla32_and7932_y0, h_u_cla32_and7934_y0);
  and_gate and_gate_h_u_cla32_and7935_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7935_y0);
  and_gate and_gate_h_u_cla32_and7936_y0(h_u_cla32_and7935_y0, h_u_cla32_and7934_y0, h_u_cla32_and7936_y0);
  and_gate and_gate_h_u_cla32_and7937_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7937_y0);
  and_gate and_gate_h_u_cla32_and7938_y0(h_u_cla32_and7937_y0, h_u_cla32_and7936_y0, h_u_cla32_and7938_y0);
  and_gate and_gate_h_u_cla32_and7939_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7939_y0);
  and_gate and_gate_h_u_cla32_and7940_y0(h_u_cla32_and7939_y0, h_u_cla32_and7938_y0, h_u_cla32_and7940_y0);
  and_gate and_gate_h_u_cla32_and7941_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7941_y0);
  and_gate and_gate_h_u_cla32_and7942_y0(h_u_cla32_and7941_y0, h_u_cla32_and7940_y0, h_u_cla32_and7942_y0);
  and_gate and_gate_h_u_cla32_and7943_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7943_y0);
  and_gate and_gate_h_u_cla32_and7944_y0(h_u_cla32_and7943_y0, h_u_cla32_and7942_y0, h_u_cla32_and7944_y0);
  and_gate and_gate_h_u_cla32_and7945_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7945_y0);
  and_gate and_gate_h_u_cla32_and7946_y0(h_u_cla32_and7945_y0, h_u_cla32_and7944_y0, h_u_cla32_and7946_y0);
  and_gate and_gate_h_u_cla32_and7947_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7947_y0);
  and_gate and_gate_h_u_cla32_and7948_y0(h_u_cla32_and7947_y0, h_u_cla32_and7946_y0, h_u_cla32_and7948_y0);
  and_gate and_gate_h_u_cla32_and7949_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7949_y0);
  and_gate and_gate_h_u_cla32_and7950_y0(h_u_cla32_and7949_y0, h_u_cla32_and7948_y0, h_u_cla32_and7950_y0);
  and_gate and_gate_h_u_cla32_and7951_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7951_y0);
  and_gate and_gate_h_u_cla32_and7952_y0(h_u_cla32_and7951_y0, h_u_cla32_and7950_y0, h_u_cla32_and7952_y0);
  and_gate and_gate_h_u_cla32_and7953_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7953_y0);
  and_gate and_gate_h_u_cla32_and7954_y0(h_u_cla32_and7953_y0, h_u_cla32_and7952_y0, h_u_cla32_and7954_y0);
  and_gate and_gate_h_u_cla32_and7955_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7955_y0);
  and_gate and_gate_h_u_cla32_and7956_y0(h_u_cla32_and7955_y0, h_u_cla32_and7954_y0, h_u_cla32_and7956_y0);
  and_gate and_gate_h_u_cla32_and7957_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7957_y0);
  and_gate and_gate_h_u_cla32_and7958_y0(h_u_cla32_and7957_y0, h_u_cla32_and7956_y0, h_u_cla32_and7958_y0);
  and_gate and_gate_h_u_cla32_and7959_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7959_y0);
  and_gate and_gate_h_u_cla32_and7960_y0(h_u_cla32_and7959_y0, h_u_cla32_and7958_y0, h_u_cla32_and7960_y0);
  and_gate and_gate_h_u_cla32_and7961_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7961_y0);
  and_gate and_gate_h_u_cla32_and7962_y0(h_u_cla32_and7961_y0, h_u_cla32_and7960_y0, h_u_cla32_and7962_y0);
  and_gate and_gate_h_u_cla32_and7963_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7963_y0);
  and_gate and_gate_h_u_cla32_and7964_y0(h_u_cla32_and7963_y0, h_u_cla32_and7962_y0, h_u_cla32_and7964_y0);
  and_gate and_gate_h_u_cla32_and7965_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7965_y0);
  and_gate and_gate_h_u_cla32_and7966_y0(h_u_cla32_and7965_y0, h_u_cla32_and7964_y0, h_u_cla32_and7966_y0);
  and_gate and_gate_h_u_cla32_and7967_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7967_y0);
  and_gate and_gate_h_u_cla32_and7968_y0(h_u_cla32_and7967_y0, h_u_cla32_and7966_y0, h_u_cla32_and7968_y0);
  and_gate and_gate_h_u_cla32_and7969_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7969_y0);
  and_gate and_gate_h_u_cla32_and7970_y0(h_u_cla32_and7969_y0, h_u_cla32_and7968_y0, h_u_cla32_and7970_y0);
  and_gate and_gate_h_u_cla32_and7971_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7971_y0);
  and_gate and_gate_h_u_cla32_and7972_y0(h_u_cla32_and7971_y0, h_u_cla32_and7970_y0, h_u_cla32_and7972_y0);
  and_gate and_gate_h_u_cla32_and7973_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7973_y0);
  and_gate and_gate_h_u_cla32_and7974_y0(h_u_cla32_and7973_y0, h_u_cla32_and7972_y0, h_u_cla32_and7974_y0);
  and_gate and_gate_h_u_cla32_and7975_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7975_y0);
  and_gate and_gate_h_u_cla32_and7976_y0(h_u_cla32_and7975_y0, h_u_cla32_and7974_y0, h_u_cla32_and7976_y0);
  and_gate and_gate_h_u_cla32_and7977_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and7977_y0);
  and_gate and_gate_h_u_cla32_and7978_y0(h_u_cla32_and7977_y0, h_u_cla32_and7976_y0, h_u_cla32_and7978_y0);
  and_gate and_gate_h_u_cla32_and7979_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7979_y0);
  and_gate and_gate_h_u_cla32_and7980_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7980_y0);
  and_gate and_gate_h_u_cla32_and7981_y0(h_u_cla32_and7980_y0, h_u_cla32_and7979_y0, h_u_cla32_and7981_y0);
  and_gate and_gate_h_u_cla32_and7982_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7982_y0);
  and_gate and_gate_h_u_cla32_and7983_y0(h_u_cla32_and7982_y0, h_u_cla32_and7981_y0, h_u_cla32_and7983_y0);
  and_gate and_gate_h_u_cla32_and7984_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7984_y0);
  and_gate and_gate_h_u_cla32_and7985_y0(h_u_cla32_and7984_y0, h_u_cla32_and7983_y0, h_u_cla32_and7985_y0);
  and_gate and_gate_h_u_cla32_and7986_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7986_y0);
  and_gate and_gate_h_u_cla32_and7987_y0(h_u_cla32_and7986_y0, h_u_cla32_and7985_y0, h_u_cla32_and7987_y0);
  and_gate and_gate_h_u_cla32_and7988_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7988_y0);
  and_gate and_gate_h_u_cla32_and7989_y0(h_u_cla32_and7988_y0, h_u_cla32_and7987_y0, h_u_cla32_and7989_y0);
  and_gate and_gate_h_u_cla32_and7990_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7990_y0);
  and_gate and_gate_h_u_cla32_and7991_y0(h_u_cla32_and7990_y0, h_u_cla32_and7989_y0, h_u_cla32_and7991_y0);
  and_gate and_gate_h_u_cla32_and7992_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7992_y0);
  and_gate and_gate_h_u_cla32_and7993_y0(h_u_cla32_and7992_y0, h_u_cla32_and7991_y0, h_u_cla32_and7993_y0);
  and_gate and_gate_h_u_cla32_and7994_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7994_y0);
  and_gate and_gate_h_u_cla32_and7995_y0(h_u_cla32_and7994_y0, h_u_cla32_and7993_y0, h_u_cla32_and7995_y0);
  and_gate and_gate_h_u_cla32_and7996_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7996_y0);
  and_gate and_gate_h_u_cla32_and7997_y0(h_u_cla32_and7996_y0, h_u_cla32_and7995_y0, h_u_cla32_and7997_y0);
  and_gate and_gate_h_u_cla32_and7998_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and7998_y0);
  and_gate and_gate_h_u_cla32_and7999_y0(h_u_cla32_and7998_y0, h_u_cla32_and7997_y0, h_u_cla32_and7999_y0);
  and_gate and_gate_h_u_cla32_and8000_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8000_y0);
  and_gate and_gate_h_u_cla32_and8001_y0(h_u_cla32_and8000_y0, h_u_cla32_and7999_y0, h_u_cla32_and8001_y0);
  and_gate and_gate_h_u_cla32_and8002_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8002_y0);
  and_gate and_gate_h_u_cla32_and8003_y0(h_u_cla32_and8002_y0, h_u_cla32_and8001_y0, h_u_cla32_and8003_y0);
  and_gate and_gate_h_u_cla32_and8004_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8004_y0);
  and_gate and_gate_h_u_cla32_and8005_y0(h_u_cla32_and8004_y0, h_u_cla32_and8003_y0, h_u_cla32_and8005_y0);
  and_gate and_gate_h_u_cla32_and8006_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8006_y0);
  and_gate and_gate_h_u_cla32_and8007_y0(h_u_cla32_and8006_y0, h_u_cla32_and8005_y0, h_u_cla32_and8007_y0);
  and_gate and_gate_h_u_cla32_and8008_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8008_y0);
  and_gate and_gate_h_u_cla32_and8009_y0(h_u_cla32_and8008_y0, h_u_cla32_and8007_y0, h_u_cla32_and8009_y0);
  and_gate and_gate_h_u_cla32_and8010_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8010_y0);
  and_gate and_gate_h_u_cla32_and8011_y0(h_u_cla32_and8010_y0, h_u_cla32_and8009_y0, h_u_cla32_and8011_y0);
  and_gate and_gate_h_u_cla32_and8012_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8012_y0);
  and_gate and_gate_h_u_cla32_and8013_y0(h_u_cla32_and8012_y0, h_u_cla32_and8011_y0, h_u_cla32_and8013_y0);
  and_gate and_gate_h_u_cla32_and8014_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8014_y0);
  and_gate and_gate_h_u_cla32_and8015_y0(h_u_cla32_and8014_y0, h_u_cla32_and8013_y0, h_u_cla32_and8015_y0);
  and_gate and_gate_h_u_cla32_and8016_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8016_y0);
  and_gate and_gate_h_u_cla32_and8017_y0(h_u_cla32_and8016_y0, h_u_cla32_and8015_y0, h_u_cla32_and8017_y0);
  and_gate and_gate_h_u_cla32_and8018_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8018_y0);
  and_gate and_gate_h_u_cla32_and8019_y0(h_u_cla32_and8018_y0, h_u_cla32_and8017_y0, h_u_cla32_and8019_y0);
  and_gate and_gate_h_u_cla32_and8020_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8020_y0);
  and_gate and_gate_h_u_cla32_and8021_y0(h_u_cla32_and8020_y0, h_u_cla32_and8019_y0, h_u_cla32_and8021_y0);
  and_gate and_gate_h_u_cla32_and8022_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8022_y0);
  and_gate and_gate_h_u_cla32_and8023_y0(h_u_cla32_and8022_y0, h_u_cla32_and8021_y0, h_u_cla32_and8023_y0);
  and_gate and_gate_h_u_cla32_and8024_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8024_y0);
  and_gate and_gate_h_u_cla32_and8025_y0(h_u_cla32_and8024_y0, h_u_cla32_and8023_y0, h_u_cla32_and8025_y0);
  and_gate and_gate_h_u_cla32_and8026_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8026_y0);
  and_gate and_gate_h_u_cla32_and8027_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8027_y0);
  and_gate and_gate_h_u_cla32_and8028_y0(h_u_cla32_and8027_y0, h_u_cla32_and8026_y0, h_u_cla32_and8028_y0);
  and_gate and_gate_h_u_cla32_and8029_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8029_y0);
  and_gate and_gate_h_u_cla32_and8030_y0(h_u_cla32_and8029_y0, h_u_cla32_and8028_y0, h_u_cla32_and8030_y0);
  and_gate and_gate_h_u_cla32_and8031_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8031_y0);
  and_gate and_gate_h_u_cla32_and8032_y0(h_u_cla32_and8031_y0, h_u_cla32_and8030_y0, h_u_cla32_and8032_y0);
  and_gate and_gate_h_u_cla32_and8033_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8033_y0);
  and_gate and_gate_h_u_cla32_and8034_y0(h_u_cla32_and8033_y0, h_u_cla32_and8032_y0, h_u_cla32_and8034_y0);
  and_gate and_gate_h_u_cla32_and8035_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8035_y0);
  and_gate and_gate_h_u_cla32_and8036_y0(h_u_cla32_and8035_y0, h_u_cla32_and8034_y0, h_u_cla32_and8036_y0);
  and_gate and_gate_h_u_cla32_and8037_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8037_y0);
  and_gate and_gate_h_u_cla32_and8038_y0(h_u_cla32_and8037_y0, h_u_cla32_and8036_y0, h_u_cla32_and8038_y0);
  and_gate and_gate_h_u_cla32_and8039_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8039_y0);
  and_gate and_gate_h_u_cla32_and8040_y0(h_u_cla32_and8039_y0, h_u_cla32_and8038_y0, h_u_cla32_and8040_y0);
  and_gate and_gate_h_u_cla32_and8041_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8041_y0);
  and_gate and_gate_h_u_cla32_and8042_y0(h_u_cla32_and8041_y0, h_u_cla32_and8040_y0, h_u_cla32_and8042_y0);
  and_gate and_gate_h_u_cla32_and8043_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8043_y0);
  and_gate and_gate_h_u_cla32_and8044_y0(h_u_cla32_and8043_y0, h_u_cla32_and8042_y0, h_u_cla32_and8044_y0);
  and_gate and_gate_h_u_cla32_and8045_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8045_y0);
  and_gate and_gate_h_u_cla32_and8046_y0(h_u_cla32_and8045_y0, h_u_cla32_and8044_y0, h_u_cla32_and8046_y0);
  and_gate and_gate_h_u_cla32_and8047_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8047_y0);
  and_gate and_gate_h_u_cla32_and8048_y0(h_u_cla32_and8047_y0, h_u_cla32_and8046_y0, h_u_cla32_and8048_y0);
  and_gate and_gate_h_u_cla32_and8049_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8049_y0);
  and_gate and_gate_h_u_cla32_and8050_y0(h_u_cla32_and8049_y0, h_u_cla32_and8048_y0, h_u_cla32_and8050_y0);
  and_gate and_gate_h_u_cla32_and8051_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8051_y0);
  and_gate and_gate_h_u_cla32_and8052_y0(h_u_cla32_and8051_y0, h_u_cla32_and8050_y0, h_u_cla32_and8052_y0);
  and_gate and_gate_h_u_cla32_and8053_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8053_y0);
  and_gate and_gate_h_u_cla32_and8054_y0(h_u_cla32_and8053_y0, h_u_cla32_and8052_y0, h_u_cla32_and8054_y0);
  and_gate and_gate_h_u_cla32_and8055_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8055_y0);
  and_gate and_gate_h_u_cla32_and8056_y0(h_u_cla32_and8055_y0, h_u_cla32_and8054_y0, h_u_cla32_and8056_y0);
  and_gate and_gate_h_u_cla32_and8057_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8057_y0);
  and_gate and_gate_h_u_cla32_and8058_y0(h_u_cla32_and8057_y0, h_u_cla32_and8056_y0, h_u_cla32_and8058_y0);
  and_gate and_gate_h_u_cla32_and8059_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8059_y0);
  and_gate and_gate_h_u_cla32_and8060_y0(h_u_cla32_and8059_y0, h_u_cla32_and8058_y0, h_u_cla32_and8060_y0);
  and_gate and_gate_h_u_cla32_and8061_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8061_y0);
  and_gate and_gate_h_u_cla32_and8062_y0(h_u_cla32_and8061_y0, h_u_cla32_and8060_y0, h_u_cla32_and8062_y0);
  and_gate and_gate_h_u_cla32_and8063_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8063_y0);
  and_gate and_gate_h_u_cla32_and8064_y0(h_u_cla32_and8063_y0, h_u_cla32_and8062_y0, h_u_cla32_and8064_y0);
  and_gate and_gate_h_u_cla32_and8065_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8065_y0);
  and_gate and_gate_h_u_cla32_and8066_y0(h_u_cla32_and8065_y0, h_u_cla32_and8064_y0, h_u_cla32_and8066_y0);
  and_gate and_gate_h_u_cla32_and8067_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8067_y0);
  and_gate and_gate_h_u_cla32_and8068_y0(h_u_cla32_and8067_y0, h_u_cla32_and8066_y0, h_u_cla32_and8068_y0);
  and_gate and_gate_h_u_cla32_and8069_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8069_y0);
  and_gate and_gate_h_u_cla32_and8070_y0(h_u_cla32_and8069_y0, h_u_cla32_and8068_y0, h_u_cla32_and8070_y0);
  and_gate and_gate_h_u_cla32_and8071_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8071_y0);
  and_gate and_gate_h_u_cla32_and8072_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8072_y0);
  and_gate and_gate_h_u_cla32_and8073_y0(h_u_cla32_and8072_y0, h_u_cla32_and8071_y0, h_u_cla32_and8073_y0);
  and_gate and_gate_h_u_cla32_and8074_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8074_y0);
  and_gate and_gate_h_u_cla32_and8075_y0(h_u_cla32_and8074_y0, h_u_cla32_and8073_y0, h_u_cla32_and8075_y0);
  and_gate and_gate_h_u_cla32_and8076_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8076_y0);
  and_gate and_gate_h_u_cla32_and8077_y0(h_u_cla32_and8076_y0, h_u_cla32_and8075_y0, h_u_cla32_and8077_y0);
  and_gate and_gate_h_u_cla32_and8078_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8078_y0);
  and_gate and_gate_h_u_cla32_and8079_y0(h_u_cla32_and8078_y0, h_u_cla32_and8077_y0, h_u_cla32_and8079_y0);
  and_gate and_gate_h_u_cla32_and8080_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8080_y0);
  and_gate and_gate_h_u_cla32_and8081_y0(h_u_cla32_and8080_y0, h_u_cla32_and8079_y0, h_u_cla32_and8081_y0);
  and_gate and_gate_h_u_cla32_and8082_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8082_y0);
  and_gate and_gate_h_u_cla32_and8083_y0(h_u_cla32_and8082_y0, h_u_cla32_and8081_y0, h_u_cla32_and8083_y0);
  and_gate and_gate_h_u_cla32_and8084_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8084_y0);
  and_gate and_gate_h_u_cla32_and8085_y0(h_u_cla32_and8084_y0, h_u_cla32_and8083_y0, h_u_cla32_and8085_y0);
  and_gate and_gate_h_u_cla32_and8086_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8086_y0);
  and_gate and_gate_h_u_cla32_and8087_y0(h_u_cla32_and8086_y0, h_u_cla32_and8085_y0, h_u_cla32_and8087_y0);
  and_gate and_gate_h_u_cla32_and8088_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8088_y0);
  and_gate and_gate_h_u_cla32_and8089_y0(h_u_cla32_and8088_y0, h_u_cla32_and8087_y0, h_u_cla32_and8089_y0);
  and_gate and_gate_h_u_cla32_and8090_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8090_y0);
  and_gate and_gate_h_u_cla32_and8091_y0(h_u_cla32_and8090_y0, h_u_cla32_and8089_y0, h_u_cla32_and8091_y0);
  and_gate and_gate_h_u_cla32_and8092_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8092_y0);
  and_gate and_gate_h_u_cla32_and8093_y0(h_u_cla32_and8092_y0, h_u_cla32_and8091_y0, h_u_cla32_and8093_y0);
  and_gate and_gate_h_u_cla32_and8094_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8094_y0);
  and_gate and_gate_h_u_cla32_and8095_y0(h_u_cla32_and8094_y0, h_u_cla32_and8093_y0, h_u_cla32_and8095_y0);
  and_gate and_gate_h_u_cla32_and8096_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8096_y0);
  and_gate and_gate_h_u_cla32_and8097_y0(h_u_cla32_and8096_y0, h_u_cla32_and8095_y0, h_u_cla32_and8097_y0);
  and_gate and_gate_h_u_cla32_and8098_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8098_y0);
  and_gate and_gate_h_u_cla32_and8099_y0(h_u_cla32_and8098_y0, h_u_cla32_and8097_y0, h_u_cla32_and8099_y0);
  and_gate and_gate_h_u_cla32_and8100_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8100_y0);
  and_gate and_gate_h_u_cla32_and8101_y0(h_u_cla32_and8100_y0, h_u_cla32_and8099_y0, h_u_cla32_and8101_y0);
  and_gate and_gate_h_u_cla32_and8102_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8102_y0);
  and_gate and_gate_h_u_cla32_and8103_y0(h_u_cla32_and8102_y0, h_u_cla32_and8101_y0, h_u_cla32_and8103_y0);
  and_gate and_gate_h_u_cla32_and8104_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8104_y0);
  and_gate and_gate_h_u_cla32_and8105_y0(h_u_cla32_and8104_y0, h_u_cla32_and8103_y0, h_u_cla32_and8105_y0);
  and_gate and_gate_h_u_cla32_and8106_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8106_y0);
  and_gate and_gate_h_u_cla32_and8107_y0(h_u_cla32_and8106_y0, h_u_cla32_and8105_y0, h_u_cla32_and8107_y0);
  and_gate and_gate_h_u_cla32_and8108_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8108_y0);
  and_gate and_gate_h_u_cla32_and8109_y0(h_u_cla32_and8108_y0, h_u_cla32_and8107_y0, h_u_cla32_and8109_y0);
  and_gate and_gate_h_u_cla32_and8110_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8110_y0);
  and_gate and_gate_h_u_cla32_and8111_y0(h_u_cla32_and8110_y0, h_u_cla32_and8109_y0, h_u_cla32_and8111_y0);
  and_gate and_gate_h_u_cla32_and8112_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8112_y0);
  and_gate and_gate_h_u_cla32_and8113_y0(h_u_cla32_and8112_y0, h_u_cla32_and8111_y0, h_u_cla32_and8113_y0);
  and_gate and_gate_h_u_cla32_and8114_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8114_y0);
  and_gate and_gate_h_u_cla32_and8115_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8115_y0);
  and_gate and_gate_h_u_cla32_and8116_y0(h_u_cla32_and8115_y0, h_u_cla32_and8114_y0, h_u_cla32_and8116_y0);
  and_gate and_gate_h_u_cla32_and8117_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8117_y0);
  and_gate and_gate_h_u_cla32_and8118_y0(h_u_cla32_and8117_y0, h_u_cla32_and8116_y0, h_u_cla32_and8118_y0);
  and_gate and_gate_h_u_cla32_and8119_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8119_y0);
  and_gate and_gate_h_u_cla32_and8120_y0(h_u_cla32_and8119_y0, h_u_cla32_and8118_y0, h_u_cla32_and8120_y0);
  and_gate and_gate_h_u_cla32_and8121_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8121_y0);
  and_gate and_gate_h_u_cla32_and8122_y0(h_u_cla32_and8121_y0, h_u_cla32_and8120_y0, h_u_cla32_and8122_y0);
  and_gate and_gate_h_u_cla32_and8123_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8123_y0);
  and_gate and_gate_h_u_cla32_and8124_y0(h_u_cla32_and8123_y0, h_u_cla32_and8122_y0, h_u_cla32_and8124_y0);
  and_gate and_gate_h_u_cla32_and8125_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8125_y0);
  and_gate and_gate_h_u_cla32_and8126_y0(h_u_cla32_and8125_y0, h_u_cla32_and8124_y0, h_u_cla32_and8126_y0);
  and_gate and_gate_h_u_cla32_and8127_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8127_y0);
  and_gate and_gate_h_u_cla32_and8128_y0(h_u_cla32_and8127_y0, h_u_cla32_and8126_y0, h_u_cla32_and8128_y0);
  and_gate and_gate_h_u_cla32_and8129_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8129_y0);
  and_gate and_gate_h_u_cla32_and8130_y0(h_u_cla32_and8129_y0, h_u_cla32_and8128_y0, h_u_cla32_and8130_y0);
  and_gate and_gate_h_u_cla32_and8131_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8131_y0);
  and_gate and_gate_h_u_cla32_and8132_y0(h_u_cla32_and8131_y0, h_u_cla32_and8130_y0, h_u_cla32_and8132_y0);
  and_gate and_gate_h_u_cla32_and8133_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8133_y0);
  and_gate and_gate_h_u_cla32_and8134_y0(h_u_cla32_and8133_y0, h_u_cla32_and8132_y0, h_u_cla32_and8134_y0);
  and_gate and_gate_h_u_cla32_and8135_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8135_y0);
  and_gate and_gate_h_u_cla32_and8136_y0(h_u_cla32_and8135_y0, h_u_cla32_and8134_y0, h_u_cla32_and8136_y0);
  and_gate and_gate_h_u_cla32_and8137_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8137_y0);
  and_gate and_gate_h_u_cla32_and8138_y0(h_u_cla32_and8137_y0, h_u_cla32_and8136_y0, h_u_cla32_and8138_y0);
  and_gate and_gate_h_u_cla32_and8139_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8139_y0);
  and_gate and_gate_h_u_cla32_and8140_y0(h_u_cla32_and8139_y0, h_u_cla32_and8138_y0, h_u_cla32_and8140_y0);
  and_gate and_gate_h_u_cla32_and8141_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8141_y0);
  and_gate and_gate_h_u_cla32_and8142_y0(h_u_cla32_and8141_y0, h_u_cla32_and8140_y0, h_u_cla32_and8142_y0);
  and_gate and_gate_h_u_cla32_and8143_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8143_y0);
  and_gate and_gate_h_u_cla32_and8144_y0(h_u_cla32_and8143_y0, h_u_cla32_and8142_y0, h_u_cla32_and8144_y0);
  and_gate and_gate_h_u_cla32_and8145_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8145_y0);
  and_gate and_gate_h_u_cla32_and8146_y0(h_u_cla32_and8145_y0, h_u_cla32_and8144_y0, h_u_cla32_and8146_y0);
  and_gate and_gate_h_u_cla32_and8147_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8147_y0);
  and_gate and_gate_h_u_cla32_and8148_y0(h_u_cla32_and8147_y0, h_u_cla32_and8146_y0, h_u_cla32_and8148_y0);
  and_gate and_gate_h_u_cla32_and8149_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8149_y0);
  and_gate and_gate_h_u_cla32_and8150_y0(h_u_cla32_and8149_y0, h_u_cla32_and8148_y0, h_u_cla32_and8150_y0);
  and_gate and_gate_h_u_cla32_and8151_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8151_y0);
  and_gate and_gate_h_u_cla32_and8152_y0(h_u_cla32_and8151_y0, h_u_cla32_and8150_y0, h_u_cla32_and8152_y0);
  and_gate and_gate_h_u_cla32_and8153_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8153_y0);
  and_gate and_gate_h_u_cla32_and8154_y0(h_u_cla32_and8153_y0, h_u_cla32_and8152_y0, h_u_cla32_and8154_y0);
  and_gate and_gate_h_u_cla32_and8155_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8155_y0);
  and_gate and_gate_h_u_cla32_and8156_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8156_y0);
  and_gate and_gate_h_u_cla32_and8157_y0(h_u_cla32_and8156_y0, h_u_cla32_and8155_y0, h_u_cla32_and8157_y0);
  and_gate and_gate_h_u_cla32_and8158_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8158_y0);
  and_gate and_gate_h_u_cla32_and8159_y0(h_u_cla32_and8158_y0, h_u_cla32_and8157_y0, h_u_cla32_and8159_y0);
  and_gate and_gate_h_u_cla32_and8160_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8160_y0);
  and_gate and_gate_h_u_cla32_and8161_y0(h_u_cla32_and8160_y0, h_u_cla32_and8159_y0, h_u_cla32_and8161_y0);
  and_gate and_gate_h_u_cla32_and8162_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8162_y0);
  and_gate and_gate_h_u_cla32_and8163_y0(h_u_cla32_and8162_y0, h_u_cla32_and8161_y0, h_u_cla32_and8163_y0);
  and_gate and_gate_h_u_cla32_and8164_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8164_y0);
  and_gate and_gate_h_u_cla32_and8165_y0(h_u_cla32_and8164_y0, h_u_cla32_and8163_y0, h_u_cla32_and8165_y0);
  and_gate and_gate_h_u_cla32_and8166_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8166_y0);
  and_gate and_gate_h_u_cla32_and8167_y0(h_u_cla32_and8166_y0, h_u_cla32_and8165_y0, h_u_cla32_and8167_y0);
  and_gate and_gate_h_u_cla32_and8168_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8168_y0);
  and_gate and_gate_h_u_cla32_and8169_y0(h_u_cla32_and8168_y0, h_u_cla32_and8167_y0, h_u_cla32_and8169_y0);
  and_gate and_gate_h_u_cla32_and8170_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8170_y0);
  and_gate and_gate_h_u_cla32_and8171_y0(h_u_cla32_and8170_y0, h_u_cla32_and8169_y0, h_u_cla32_and8171_y0);
  and_gate and_gate_h_u_cla32_and8172_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8172_y0);
  and_gate and_gate_h_u_cla32_and8173_y0(h_u_cla32_and8172_y0, h_u_cla32_and8171_y0, h_u_cla32_and8173_y0);
  and_gate and_gate_h_u_cla32_and8174_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8174_y0);
  and_gate and_gate_h_u_cla32_and8175_y0(h_u_cla32_and8174_y0, h_u_cla32_and8173_y0, h_u_cla32_and8175_y0);
  and_gate and_gate_h_u_cla32_and8176_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8176_y0);
  and_gate and_gate_h_u_cla32_and8177_y0(h_u_cla32_and8176_y0, h_u_cla32_and8175_y0, h_u_cla32_and8177_y0);
  and_gate and_gate_h_u_cla32_and8178_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8178_y0);
  and_gate and_gate_h_u_cla32_and8179_y0(h_u_cla32_and8178_y0, h_u_cla32_and8177_y0, h_u_cla32_and8179_y0);
  and_gate and_gate_h_u_cla32_and8180_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8180_y0);
  and_gate and_gate_h_u_cla32_and8181_y0(h_u_cla32_and8180_y0, h_u_cla32_and8179_y0, h_u_cla32_and8181_y0);
  and_gate and_gate_h_u_cla32_and8182_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8182_y0);
  and_gate and_gate_h_u_cla32_and8183_y0(h_u_cla32_and8182_y0, h_u_cla32_and8181_y0, h_u_cla32_and8183_y0);
  and_gate and_gate_h_u_cla32_and8184_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8184_y0);
  and_gate and_gate_h_u_cla32_and8185_y0(h_u_cla32_and8184_y0, h_u_cla32_and8183_y0, h_u_cla32_and8185_y0);
  and_gate and_gate_h_u_cla32_and8186_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8186_y0);
  and_gate and_gate_h_u_cla32_and8187_y0(h_u_cla32_and8186_y0, h_u_cla32_and8185_y0, h_u_cla32_and8187_y0);
  and_gate and_gate_h_u_cla32_and8188_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8188_y0);
  and_gate and_gate_h_u_cla32_and8189_y0(h_u_cla32_and8188_y0, h_u_cla32_and8187_y0, h_u_cla32_and8189_y0);
  and_gate and_gate_h_u_cla32_and8190_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8190_y0);
  and_gate and_gate_h_u_cla32_and8191_y0(h_u_cla32_and8190_y0, h_u_cla32_and8189_y0, h_u_cla32_and8191_y0);
  and_gate and_gate_h_u_cla32_and8192_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and8192_y0);
  and_gate and_gate_h_u_cla32_and8193_y0(h_u_cla32_and8192_y0, h_u_cla32_and8191_y0, h_u_cla32_and8193_y0);
  and_gate and_gate_h_u_cla32_and8194_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8194_y0);
  and_gate and_gate_h_u_cla32_and8195_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8195_y0);
  and_gate and_gate_h_u_cla32_and8196_y0(h_u_cla32_and8195_y0, h_u_cla32_and8194_y0, h_u_cla32_and8196_y0);
  and_gate and_gate_h_u_cla32_and8197_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8197_y0);
  and_gate and_gate_h_u_cla32_and8198_y0(h_u_cla32_and8197_y0, h_u_cla32_and8196_y0, h_u_cla32_and8198_y0);
  and_gate and_gate_h_u_cla32_and8199_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8199_y0);
  and_gate and_gate_h_u_cla32_and8200_y0(h_u_cla32_and8199_y0, h_u_cla32_and8198_y0, h_u_cla32_and8200_y0);
  and_gate and_gate_h_u_cla32_and8201_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8201_y0);
  and_gate and_gate_h_u_cla32_and8202_y0(h_u_cla32_and8201_y0, h_u_cla32_and8200_y0, h_u_cla32_and8202_y0);
  and_gate and_gate_h_u_cla32_and8203_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8203_y0);
  and_gate and_gate_h_u_cla32_and8204_y0(h_u_cla32_and8203_y0, h_u_cla32_and8202_y0, h_u_cla32_and8204_y0);
  and_gate and_gate_h_u_cla32_and8205_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8205_y0);
  and_gate and_gate_h_u_cla32_and8206_y0(h_u_cla32_and8205_y0, h_u_cla32_and8204_y0, h_u_cla32_and8206_y0);
  and_gate and_gate_h_u_cla32_and8207_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8207_y0);
  and_gate and_gate_h_u_cla32_and8208_y0(h_u_cla32_and8207_y0, h_u_cla32_and8206_y0, h_u_cla32_and8208_y0);
  and_gate and_gate_h_u_cla32_and8209_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8209_y0);
  and_gate and_gate_h_u_cla32_and8210_y0(h_u_cla32_and8209_y0, h_u_cla32_and8208_y0, h_u_cla32_and8210_y0);
  and_gate and_gate_h_u_cla32_and8211_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8211_y0);
  and_gate and_gate_h_u_cla32_and8212_y0(h_u_cla32_and8211_y0, h_u_cla32_and8210_y0, h_u_cla32_and8212_y0);
  and_gate and_gate_h_u_cla32_and8213_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8213_y0);
  and_gate and_gate_h_u_cla32_and8214_y0(h_u_cla32_and8213_y0, h_u_cla32_and8212_y0, h_u_cla32_and8214_y0);
  and_gate and_gate_h_u_cla32_and8215_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8215_y0);
  and_gate and_gate_h_u_cla32_and8216_y0(h_u_cla32_and8215_y0, h_u_cla32_and8214_y0, h_u_cla32_and8216_y0);
  and_gate and_gate_h_u_cla32_and8217_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8217_y0);
  and_gate and_gate_h_u_cla32_and8218_y0(h_u_cla32_and8217_y0, h_u_cla32_and8216_y0, h_u_cla32_and8218_y0);
  and_gate and_gate_h_u_cla32_and8219_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8219_y0);
  and_gate and_gate_h_u_cla32_and8220_y0(h_u_cla32_and8219_y0, h_u_cla32_and8218_y0, h_u_cla32_and8220_y0);
  and_gate and_gate_h_u_cla32_and8221_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8221_y0);
  and_gate and_gate_h_u_cla32_and8222_y0(h_u_cla32_and8221_y0, h_u_cla32_and8220_y0, h_u_cla32_and8222_y0);
  and_gate and_gate_h_u_cla32_and8223_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8223_y0);
  and_gate and_gate_h_u_cla32_and8224_y0(h_u_cla32_and8223_y0, h_u_cla32_and8222_y0, h_u_cla32_and8224_y0);
  and_gate and_gate_h_u_cla32_and8225_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8225_y0);
  and_gate and_gate_h_u_cla32_and8226_y0(h_u_cla32_and8225_y0, h_u_cla32_and8224_y0, h_u_cla32_and8226_y0);
  and_gate and_gate_h_u_cla32_and8227_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8227_y0);
  and_gate and_gate_h_u_cla32_and8228_y0(h_u_cla32_and8227_y0, h_u_cla32_and8226_y0, h_u_cla32_and8228_y0);
  and_gate and_gate_h_u_cla32_and8229_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and8229_y0);
  and_gate and_gate_h_u_cla32_and8230_y0(h_u_cla32_and8229_y0, h_u_cla32_and8228_y0, h_u_cla32_and8230_y0);
  and_gate and_gate_h_u_cla32_and8231_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8231_y0);
  and_gate and_gate_h_u_cla32_and8232_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8232_y0);
  and_gate and_gate_h_u_cla32_and8233_y0(h_u_cla32_and8232_y0, h_u_cla32_and8231_y0, h_u_cla32_and8233_y0);
  and_gate and_gate_h_u_cla32_and8234_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8234_y0);
  and_gate and_gate_h_u_cla32_and8235_y0(h_u_cla32_and8234_y0, h_u_cla32_and8233_y0, h_u_cla32_and8235_y0);
  and_gate and_gate_h_u_cla32_and8236_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8236_y0);
  and_gate and_gate_h_u_cla32_and8237_y0(h_u_cla32_and8236_y0, h_u_cla32_and8235_y0, h_u_cla32_and8237_y0);
  and_gate and_gate_h_u_cla32_and8238_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8238_y0);
  and_gate and_gate_h_u_cla32_and8239_y0(h_u_cla32_and8238_y0, h_u_cla32_and8237_y0, h_u_cla32_and8239_y0);
  and_gate and_gate_h_u_cla32_and8240_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8240_y0);
  and_gate and_gate_h_u_cla32_and8241_y0(h_u_cla32_and8240_y0, h_u_cla32_and8239_y0, h_u_cla32_and8241_y0);
  and_gate and_gate_h_u_cla32_and8242_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8242_y0);
  and_gate and_gate_h_u_cla32_and8243_y0(h_u_cla32_and8242_y0, h_u_cla32_and8241_y0, h_u_cla32_and8243_y0);
  and_gate and_gate_h_u_cla32_and8244_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8244_y0);
  and_gate and_gate_h_u_cla32_and8245_y0(h_u_cla32_and8244_y0, h_u_cla32_and8243_y0, h_u_cla32_and8245_y0);
  and_gate and_gate_h_u_cla32_and8246_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8246_y0);
  and_gate and_gate_h_u_cla32_and8247_y0(h_u_cla32_and8246_y0, h_u_cla32_and8245_y0, h_u_cla32_and8247_y0);
  and_gate and_gate_h_u_cla32_and8248_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8248_y0);
  and_gate and_gate_h_u_cla32_and8249_y0(h_u_cla32_and8248_y0, h_u_cla32_and8247_y0, h_u_cla32_and8249_y0);
  and_gate and_gate_h_u_cla32_and8250_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8250_y0);
  and_gate and_gate_h_u_cla32_and8251_y0(h_u_cla32_and8250_y0, h_u_cla32_and8249_y0, h_u_cla32_and8251_y0);
  and_gate and_gate_h_u_cla32_and8252_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8252_y0);
  and_gate and_gate_h_u_cla32_and8253_y0(h_u_cla32_and8252_y0, h_u_cla32_and8251_y0, h_u_cla32_and8253_y0);
  and_gate and_gate_h_u_cla32_and8254_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8254_y0);
  and_gate and_gate_h_u_cla32_and8255_y0(h_u_cla32_and8254_y0, h_u_cla32_and8253_y0, h_u_cla32_and8255_y0);
  and_gate and_gate_h_u_cla32_and8256_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8256_y0);
  and_gate and_gate_h_u_cla32_and8257_y0(h_u_cla32_and8256_y0, h_u_cla32_and8255_y0, h_u_cla32_and8257_y0);
  and_gate and_gate_h_u_cla32_and8258_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8258_y0);
  and_gate and_gate_h_u_cla32_and8259_y0(h_u_cla32_and8258_y0, h_u_cla32_and8257_y0, h_u_cla32_and8259_y0);
  and_gate and_gate_h_u_cla32_and8260_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8260_y0);
  and_gate and_gate_h_u_cla32_and8261_y0(h_u_cla32_and8260_y0, h_u_cla32_and8259_y0, h_u_cla32_and8261_y0);
  and_gate and_gate_h_u_cla32_and8262_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8262_y0);
  and_gate and_gate_h_u_cla32_and8263_y0(h_u_cla32_and8262_y0, h_u_cla32_and8261_y0, h_u_cla32_and8263_y0);
  and_gate and_gate_h_u_cla32_and8264_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and8264_y0);
  and_gate and_gate_h_u_cla32_and8265_y0(h_u_cla32_and8264_y0, h_u_cla32_and8263_y0, h_u_cla32_and8265_y0);
  and_gate and_gate_h_u_cla32_and8266_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8266_y0);
  and_gate and_gate_h_u_cla32_and8267_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8267_y0);
  and_gate and_gate_h_u_cla32_and8268_y0(h_u_cla32_and8267_y0, h_u_cla32_and8266_y0, h_u_cla32_and8268_y0);
  and_gate and_gate_h_u_cla32_and8269_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8269_y0);
  and_gate and_gate_h_u_cla32_and8270_y0(h_u_cla32_and8269_y0, h_u_cla32_and8268_y0, h_u_cla32_and8270_y0);
  and_gate and_gate_h_u_cla32_and8271_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8271_y0);
  and_gate and_gate_h_u_cla32_and8272_y0(h_u_cla32_and8271_y0, h_u_cla32_and8270_y0, h_u_cla32_and8272_y0);
  and_gate and_gate_h_u_cla32_and8273_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8273_y0);
  and_gate and_gate_h_u_cla32_and8274_y0(h_u_cla32_and8273_y0, h_u_cla32_and8272_y0, h_u_cla32_and8274_y0);
  and_gate and_gate_h_u_cla32_and8275_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8275_y0);
  and_gate and_gate_h_u_cla32_and8276_y0(h_u_cla32_and8275_y0, h_u_cla32_and8274_y0, h_u_cla32_and8276_y0);
  and_gate and_gate_h_u_cla32_and8277_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8277_y0);
  and_gate and_gate_h_u_cla32_and8278_y0(h_u_cla32_and8277_y0, h_u_cla32_and8276_y0, h_u_cla32_and8278_y0);
  and_gate and_gate_h_u_cla32_and8279_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8279_y0);
  and_gate and_gate_h_u_cla32_and8280_y0(h_u_cla32_and8279_y0, h_u_cla32_and8278_y0, h_u_cla32_and8280_y0);
  and_gate and_gate_h_u_cla32_and8281_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8281_y0);
  and_gate and_gate_h_u_cla32_and8282_y0(h_u_cla32_and8281_y0, h_u_cla32_and8280_y0, h_u_cla32_and8282_y0);
  and_gate and_gate_h_u_cla32_and8283_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8283_y0);
  and_gate and_gate_h_u_cla32_and8284_y0(h_u_cla32_and8283_y0, h_u_cla32_and8282_y0, h_u_cla32_and8284_y0);
  and_gate and_gate_h_u_cla32_and8285_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8285_y0);
  and_gate and_gate_h_u_cla32_and8286_y0(h_u_cla32_and8285_y0, h_u_cla32_and8284_y0, h_u_cla32_and8286_y0);
  and_gate and_gate_h_u_cla32_and8287_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8287_y0);
  and_gate and_gate_h_u_cla32_and8288_y0(h_u_cla32_and8287_y0, h_u_cla32_and8286_y0, h_u_cla32_and8288_y0);
  and_gate and_gate_h_u_cla32_and8289_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8289_y0);
  and_gate and_gate_h_u_cla32_and8290_y0(h_u_cla32_and8289_y0, h_u_cla32_and8288_y0, h_u_cla32_and8290_y0);
  and_gate and_gate_h_u_cla32_and8291_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8291_y0);
  and_gate and_gate_h_u_cla32_and8292_y0(h_u_cla32_and8291_y0, h_u_cla32_and8290_y0, h_u_cla32_and8292_y0);
  and_gate and_gate_h_u_cla32_and8293_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8293_y0);
  and_gate and_gate_h_u_cla32_and8294_y0(h_u_cla32_and8293_y0, h_u_cla32_and8292_y0, h_u_cla32_and8294_y0);
  and_gate and_gate_h_u_cla32_and8295_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8295_y0);
  and_gate and_gate_h_u_cla32_and8296_y0(h_u_cla32_and8295_y0, h_u_cla32_and8294_y0, h_u_cla32_and8296_y0);
  and_gate and_gate_h_u_cla32_and8297_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and8297_y0);
  and_gate and_gate_h_u_cla32_and8298_y0(h_u_cla32_and8297_y0, h_u_cla32_and8296_y0, h_u_cla32_and8298_y0);
  and_gate and_gate_h_u_cla32_and8299_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8299_y0);
  and_gate and_gate_h_u_cla32_and8300_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8300_y0);
  and_gate and_gate_h_u_cla32_and8301_y0(h_u_cla32_and8300_y0, h_u_cla32_and8299_y0, h_u_cla32_and8301_y0);
  and_gate and_gate_h_u_cla32_and8302_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8302_y0);
  and_gate and_gate_h_u_cla32_and8303_y0(h_u_cla32_and8302_y0, h_u_cla32_and8301_y0, h_u_cla32_and8303_y0);
  and_gate and_gate_h_u_cla32_and8304_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8304_y0);
  and_gate and_gate_h_u_cla32_and8305_y0(h_u_cla32_and8304_y0, h_u_cla32_and8303_y0, h_u_cla32_and8305_y0);
  and_gate and_gate_h_u_cla32_and8306_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8306_y0);
  and_gate and_gate_h_u_cla32_and8307_y0(h_u_cla32_and8306_y0, h_u_cla32_and8305_y0, h_u_cla32_and8307_y0);
  and_gate and_gate_h_u_cla32_and8308_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8308_y0);
  and_gate and_gate_h_u_cla32_and8309_y0(h_u_cla32_and8308_y0, h_u_cla32_and8307_y0, h_u_cla32_and8309_y0);
  and_gate and_gate_h_u_cla32_and8310_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8310_y0);
  and_gate and_gate_h_u_cla32_and8311_y0(h_u_cla32_and8310_y0, h_u_cla32_and8309_y0, h_u_cla32_and8311_y0);
  and_gate and_gate_h_u_cla32_and8312_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8312_y0);
  and_gate and_gate_h_u_cla32_and8313_y0(h_u_cla32_and8312_y0, h_u_cla32_and8311_y0, h_u_cla32_and8313_y0);
  and_gate and_gate_h_u_cla32_and8314_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8314_y0);
  and_gate and_gate_h_u_cla32_and8315_y0(h_u_cla32_and8314_y0, h_u_cla32_and8313_y0, h_u_cla32_and8315_y0);
  and_gate and_gate_h_u_cla32_and8316_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8316_y0);
  and_gate and_gate_h_u_cla32_and8317_y0(h_u_cla32_and8316_y0, h_u_cla32_and8315_y0, h_u_cla32_and8317_y0);
  and_gate and_gate_h_u_cla32_and8318_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8318_y0);
  and_gate and_gate_h_u_cla32_and8319_y0(h_u_cla32_and8318_y0, h_u_cla32_and8317_y0, h_u_cla32_and8319_y0);
  and_gate and_gate_h_u_cla32_and8320_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8320_y0);
  and_gate and_gate_h_u_cla32_and8321_y0(h_u_cla32_and8320_y0, h_u_cla32_and8319_y0, h_u_cla32_and8321_y0);
  and_gate and_gate_h_u_cla32_and8322_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8322_y0);
  and_gate and_gate_h_u_cla32_and8323_y0(h_u_cla32_and8322_y0, h_u_cla32_and8321_y0, h_u_cla32_and8323_y0);
  and_gate and_gate_h_u_cla32_and8324_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8324_y0);
  and_gate and_gate_h_u_cla32_and8325_y0(h_u_cla32_and8324_y0, h_u_cla32_and8323_y0, h_u_cla32_and8325_y0);
  and_gate and_gate_h_u_cla32_and8326_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8326_y0);
  and_gate and_gate_h_u_cla32_and8327_y0(h_u_cla32_and8326_y0, h_u_cla32_and8325_y0, h_u_cla32_and8327_y0);
  and_gate and_gate_h_u_cla32_and8328_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and8328_y0);
  and_gate and_gate_h_u_cla32_and8329_y0(h_u_cla32_and8328_y0, h_u_cla32_and8327_y0, h_u_cla32_and8329_y0);
  and_gate and_gate_h_u_cla32_and8330_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8330_y0);
  and_gate and_gate_h_u_cla32_and8331_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8331_y0);
  and_gate and_gate_h_u_cla32_and8332_y0(h_u_cla32_and8331_y0, h_u_cla32_and8330_y0, h_u_cla32_and8332_y0);
  and_gate and_gate_h_u_cla32_and8333_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8333_y0);
  and_gate and_gate_h_u_cla32_and8334_y0(h_u_cla32_and8333_y0, h_u_cla32_and8332_y0, h_u_cla32_and8334_y0);
  and_gate and_gate_h_u_cla32_and8335_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8335_y0);
  and_gate and_gate_h_u_cla32_and8336_y0(h_u_cla32_and8335_y0, h_u_cla32_and8334_y0, h_u_cla32_and8336_y0);
  and_gate and_gate_h_u_cla32_and8337_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8337_y0);
  and_gate and_gate_h_u_cla32_and8338_y0(h_u_cla32_and8337_y0, h_u_cla32_and8336_y0, h_u_cla32_and8338_y0);
  and_gate and_gate_h_u_cla32_and8339_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8339_y0);
  and_gate and_gate_h_u_cla32_and8340_y0(h_u_cla32_and8339_y0, h_u_cla32_and8338_y0, h_u_cla32_and8340_y0);
  and_gate and_gate_h_u_cla32_and8341_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8341_y0);
  and_gate and_gate_h_u_cla32_and8342_y0(h_u_cla32_and8341_y0, h_u_cla32_and8340_y0, h_u_cla32_and8342_y0);
  and_gate and_gate_h_u_cla32_and8343_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8343_y0);
  and_gate and_gate_h_u_cla32_and8344_y0(h_u_cla32_and8343_y0, h_u_cla32_and8342_y0, h_u_cla32_and8344_y0);
  and_gate and_gate_h_u_cla32_and8345_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8345_y0);
  and_gate and_gate_h_u_cla32_and8346_y0(h_u_cla32_and8345_y0, h_u_cla32_and8344_y0, h_u_cla32_and8346_y0);
  and_gate and_gate_h_u_cla32_and8347_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8347_y0);
  and_gate and_gate_h_u_cla32_and8348_y0(h_u_cla32_and8347_y0, h_u_cla32_and8346_y0, h_u_cla32_and8348_y0);
  and_gate and_gate_h_u_cla32_and8349_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8349_y0);
  and_gate and_gate_h_u_cla32_and8350_y0(h_u_cla32_and8349_y0, h_u_cla32_and8348_y0, h_u_cla32_and8350_y0);
  and_gate and_gate_h_u_cla32_and8351_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8351_y0);
  and_gate and_gate_h_u_cla32_and8352_y0(h_u_cla32_and8351_y0, h_u_cla32_and8350_y0, h_u_cla32_and8352_y0);
  and_gate and_gate_h_u_cla32_and8353_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8353_y0);
  and_gate and_gate_h_u_cla32_and8354_y0(h_u_cla32_and8353_y0, h_u_cla32_and8352_y0, h_u_cla32_and8354_y0);
  and_gate and_gate_h_u_cla32_and8355_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8355_y0);
  and_gate and_gate_h_u_cla32_and8356_y0(h_u_cla32_and8355_y0, h_u_cla32_and8354_y0, h_u_cla32_and8356_y0);
  and_gate and_gate_h_u_cla32_and8357_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and8357_y0);
  and_gate and_gate_h_u_cla32_and8358_y0(h_u_cla32_and8357_y0, h_u_cla32_and8356_y0, h_u_cla32_and8358_y0);
  and_gate and_gate_h_u_cla32_and8359_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8359_y0);
  and_gate and_gate_h_u_cla32_and8360_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8360_y0);
  and_gate and_gate_h_u_cla32_and8361_y0(h_u_cla32_and8360_y0, h_u_cla32_and8359_y0, h_u_cla32_and8361_y0);
  and_gate and_gate_h_u_cla32_and8362_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8362_y0);
  and_gate and_gate_h_u_cla32_and8363_y0(h_u_cla32_and8362_y0, h_u_cla32_and8361_y0, h_u_cla32_and8363_y0);
  and_gate and_gate_h_u_cla32_and8364_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8364_y0);
  and_gate and_gate_h_u_cla32_and8365_y0(h_u_cla32_and8364_y0, h_u_cla32_and8363_y0, h_u_cla32_and8365_y0);
  and_gate and_gate_h_u_cla32_and8366_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8366_y0);
  and_gate and_gate_h_u_cla32_and8367_y0(h_u_cla32_and8366_y0, h_u_cla32_and8365_y0, h_u_cla32_and8367_y0);
  and_gate and_gate_h_u_cla32_and8368_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8368_y0);
  and_gate and_gate_h_u_cla32_and8369_y0(h_u_cla32_and8368_y0, h_u_cla32_and8367_y0, h_u_cla32_and8369_y0);
  and_gate and_gate_h_u_cla32_and8370_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8370_y0);
  and_gate and_gate_h_u_cla32_and8371_y0(h_u_cla32_and8370_y0, h_u_cla32_and8369_y0, h_u_cla32_and8371_y0);
  and_gate and_gate_h_u_cla32_and8372_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8372_y0);
  and_gate and_gate_h_u_cla32_and8373_y0(h_u_cla32_and8372_y0, h_u_cla32_and8371_y0, h_u_cla32_and8373_y0);
  and_gate and_gate_h_u_cla32_and8374_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8374_y0);
  and_gate and_gate_h_u_cla32_and8375_y0(h_u_cla32_and8374_y0, h_u_cla32_and8373_y0, h_u_cla32_and8375_y0);
  and_gate and_gate_h_u_cla32_and8376_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8376_y0);
  and_gate and_gate_h_u_cla32_and8377_y0(h_u_cla32_and8376_y0, h_u_cla32_and8375_y0, h_u_cla32_and8377_y0);
  and_gate and_gate_h_u_cla32_and8378_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8378_y0);
  and_gate and_gate_h_u_cla32_and8379_y0(h_u_cla32_and8378_y0, h_u_cla32_and8377_y0, h_u_cla32_and8379_y0);
  and_gate and_gate_h_u_cla32_and8380_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8380_y0);
  and_gate and_gate_h_u_cla32_and8381_y0(h_u_cla32_and8380_y0, h_u_cla32_and8379_y0, h_u_cla32_and8381_y0);
  and_gate and_gate_h_u_cla32_and8382_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8382_y0);
  and_gate and_gate_h_u_cla32_and8383_y0(h_u_cla32_and8382_y0, h_u_cla32_and8381_y0, h_u_cla32_and8383_y0);
  and_gate and_gate_h_u_cla32_and8384_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and8384_y0);
  and_gate and_gate_h_u_cla32_and8385_y0(h_u_cla32_and8384_y0, h_u_cla32_and8383_y0, h_u_cla32_and8385_y0);
  and_gate and_gate_h_u_cla32_and8386_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8386_y0);
  and_gate and_gate_h_u_cla32_and8387_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8387_y0);
  and_gate and_gate_h_u_cla32_and8388_y0(h_u_cla32_and8387_y0, h_u_cla32_and8386_y0, h_u_cla32_and8388_y0);
  and_gate and_gate_h_u_cla32_and8389_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8389_y0);
  and_gate and_gate_h_u_cla32_and8390_y0(h_u_cla32_and8389_y0, h_u_cla32_and8388_y0, h_u_cla32_and8390_y0);
  and_gate and_gate_h_u_cla32_and8391_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8391_y0);
  and_gate and_gate_h_u_cla32_and8392_y0(h_u_cla32_and8391_y0, h_u_cla32_and8390_y0, h_u_cla32_and8392_y0);
  and_gate and_gate_h_u_cla32_and8393_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8393_y0);
  and_gate and_gate_h_u_cla32_and8394_y0(h_u_cla32_and8393_y0, h_u_cla32_and8392_y0, h_u_cla32_and8394_y0);
  and_gate and_gate_h_u_cla32_and8395_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8395_y0);
  and_gate and_gate_h_u_cla32_and8396_y0(h_u_cla32_and8395_y0, h_u_cla32_and8394_y0, h_u_cla32_and8396_y0);
  and_gate and_gate_h_u_cla32_and8397_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8397_y0);
  and_gate and_gate_h_u_cla32_and8398_y0(h_u_cla32_and8397_y0, h_u_cla32_and8396_y0, h_u_cla32_and8398_y0);
  and_gate and_gate_h_u_cla32_and8399_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8399_y0);
  and_gate and_gate_h_u_cla32_and8400_y0(h_u_cla32_and8399_y0, h_u_cla32_and8398_y0, h_u_cla32_and8400_y0);
  and_gate and_gate_h_u_cla32_and8401_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8401_y0);
  and_gate and_gate_h_u_cla32_and8402_y0(h_u_cla32_and8401_y0, h_u_cla32_and8400_y0, h_u_cla32_and8402_y0);
  and_gate and_gate_h_u_cla32_and8403_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8403_y0);
  and_gate and_gate_h_u_cla32_and8404_y0(h_u_cla32_and8403_y0, h_u_cla32_and8402_y0, h_u_cla32_and8404_y0);
  and_gate and_gate_h_u_cla32_and8405_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8405_y0);
  and_gate and_gate_h_u_cla32_and8406_y0(h_u_cla32_and8405_y0, h_u_cla32_and8404_y0, h_u_cla32_and8406_y0);
  and_gate and_gate_h_u_cla32_and8407_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8407_y0);
  and_gate and_gate_h_u_cla32_and8408_y0(h_u_cla32_and8407_y0, h_u_cla32_and8406_y0, h_u_cla32_and8408_y0);
  and_gate and_gate_h_u_cla32_and8409_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and8409_y0);
  and_gate and_gate_h_u_cla32_and8410_y0(h_u_cla32_and8409_y0, h_u_cla32_and8408_y0, h_u_cla32_and8410_y0);
  and_gate and_gate_h_u_cla32_and8411_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8411_y0);
  and_gate and_gate_h_u_cla32_and8412_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8412_y0);
  and_gate and_gate_h_u_cla32_and8413_y0(h_u_cla32_and8412_y0, h_u_cla32_and8411_y0, h_u_cla32_and8413_y0);
  and_gate and_gate_h_u_cla32_and8414_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8414_y0);
  and_gate and_gate_h_u_cla32_and8415_y0(h_u_cla32_and8414_y0, h_u_cla32_and8413_y0, h_u_cla32_and8415_y0);
  and_gate and_gate_h_u_cla32_and8416_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8416_y0);
  and_gate and_gate_h_u_cla32_and8417_y0(h_u_cla32_and8416_y0, h_u_cla32_and8415_y0, h_u_cla32_and8417_y0);
  and_gate and_gate_h_u_cla32_and8418_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8418_y0);
  and_gate and_gate_h_u_cla32_and8419_y0(h_u_cla32_and8418_y0, h_u_cla32_and8417_y0, h_u_cla32_and8419_y0);
  and_gate and_gate_h_u_cla32_and8420_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8420_y0);
  and_gate and_gate_h_u_cla32_and8421_y0(h_u_cla32_and8420_y0, h_u_cla32_and8419_y0, h_u_cla32_and8421_y0);
  and_gate and_gate_h_u_cla32_and8422_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8422_y0);
  and_gate and_gate_h_u_cla32_and8423_y0(h_u_cla32_and8422_y0, h_u_cla32_and8421_y0, h_u_cla32_and8423_y0);
  and_gate and_gate_h_u_cla32_and8424_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8424_y0);
  and_gate and_gate_h_u_cla32_and8425_y0(h_u_cla32_and8424_y0, h_u_cla32_and8423_y0, h_u_cla32_and8425_y0);
  and_gate and_gate_h_u_cla32_and8426_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8426_y0);
  and_gate and_gate_h_u_cla32_and8427_y0(h_u_cla32_and8426_y0, h_u_cla32_and8425_y0, h_u_cla32_and8427_y0);
  and_gate and_gate_h_u_cla32_and8428_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8428_y0);
  and_gate and_gate_h_u_cla32_and8429_y0(h_u_cla32_and8428_y0, h_u_cla32_and8427_y0, h_u_cla32_and8429_y0);
  and_gate and_gate_h_u_cla32_and8430_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8430_y0);
  and_gate and_gate_h_u_cla32_and8431_y0(h_u_cla32_and8430_y0, h_u_cla32_and8429_y0, h_u_cla32_and8431_y0);
  and_gate and_gate_h_u_cla32_and8432_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and8432_y0);
  and_gate and_gate_h_u_cla32_and8433_y0(h_u_cla32_and8432_y0, h_u_cla32_and8431_y0, h_u_cla32_and8433_y0);
  and_gate and_gate_h_u_cla32_and8434_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8434_y0);
  and_gate and_gate_h_u_cla32_and8435_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8435_y0);
  and_gate and_gate_h_u_cla32_and8436_y0(h_u_cla32_and8435_y0, h_u_cla32_and8434_y0, h_u_cla32_and8436_y0);
  and_gate and_gate_h_u_cla32_and8437_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8437_y0);
  and_gate and_gate_h_u_cla32_and8438_y0(h_u_cla32_and8437_y0, h_u_cla32_and8436_y0, h_u_cla32_and8438_y0);
  and_gate and_gate_h_u_cla32_and8439_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8439_y0);
  and_gate and_gate_h_u_cla32_and8440_y0(h_u_cla32_and8439_y0, h_u_cla32_and8438_y0, h_u_cla32_and8440_y0);
  and_gate and_gate_h_u_cla32_and8441_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8441_y0);
  and_gate and_gate_h_u_cla32_and8442_y0(h_u_cla32_and8441_y0, h_u_cla32_and8440_y0, h_u_cla32_and8442_y0);
  and_gate and_gate_h_u_cla32_and8443_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8443_y0);
  and_gate and_gate_h_u_cla32_and8444_y0(h_u_cla32_and8443_y0, h_u_cla32_and8442_y0, h_u_cla32_and8444_y0);
  and_gate and_gate_h_u_cla32_and8445_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8445_y0);
  and_gate and_gate_h_u_cla32_and8446_y0(h_u_cla32_and8445_y0, h_u_cla32_and8444_y0, h_u_cla32_and8446_y0);
  and_gate and_gate_h_u_cla32_and8447_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8447_y0);
  and_gate and_gate_h_u_cla32_and8448_y0(h_u_cla32_and8447_y0, h_u_cla32_and8446_y0, h_u_cla32_and8448_y0);
  and_gate and_gate_h_u_cla32_and8449_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8449_y0);
  and_gate and_gate_h_u_cla32_and8450_y0(h_u_cla32_and8449_y0, h_u_cla32_and8448_y0, h_u_cla32_and8450_y0);
  and_gate and_gate_h_u_cla32_and8451_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8451_y0);
  and_gate and_gate_h_u_cla32_and8452_y0(h_u_cla32_and8451_y0, h_u_cla32_and8450_y0, h_u_cla32_and8452_y0);
  and_gate and_gate_h_u_cla32_and8453_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and8453_y0);
  and_gate and_gate_h_u_cla32_and8454_y0(h_u_cla32_and8453_y0, h_u_cla32_and8452_y0, h_u_cla32_and8454_y0);
  and_gate and_gate_h_u_cla32_and8455_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8455_y0);
  and_gate and_gate_h_u_cla32_and8456_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8456_y0);
  and_gate and_gate_h_u_cla32_and8457_y0(h_u_cla32_and8456_y0, h_u_cla32_and8455_y0, h_u_cla32_and8457_y0);
  and_gate and_gate_h_u_cla32_and8458_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8458_y0);
  and_gate and_gate_h_u_cla32_and8459_y0(h_u_cla32_and8458_y0, h_u_cla32_and8457_y0, h_u_cla32_and8459_y0);
  and_gate and_gate_h_u_cla32_and8460_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8460_y0);
  and_gate and_gate_h_u_cla32_and8461_y0(h_u_cla32_and8460_y0, h_u_cla32_and8459_y0, h_u_cla32_and8461_y0);
  and_gate and_gate_h_u_cla32_and8462_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8462_y0);
  and_gate and_gate_h_u_cla32_and8463_y0(h_u_cla32_and8462_y0, h_u_cla32_and8461_y0, h_u_cla32_and8463_y0);
  and_gate and_gate_h_u_cla32_and8464_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8464_y0);
  and_gate and_gate_h_u_cla32_and8465_y0(h_u_cla32_and8464_y0, h_u_cla32_and8463_y0, h_u_cla32_and8465_y0);
  and_gate and_gate_h_u_cla32_and8466_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8466_y0);
  and_gate and_gate_h_u_cla32_and8467_y0(h_u_cla32_and8466_y0, h_u_cla32_and8465_y0, h_u_cla32_and8467_y0);
  and_gate and_gate_h_u_cla32_and8468_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8468_y0);
  and_gate and_gate_h_u_cla32_and8469_y0(h_u_cla32_and8468_y0, h_u_cla32_and8467_y0, h_u_cla32_and8469_y0);
  and_gate and_gate_h_u_cla32_and8470_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8470_y0);
  and_gate and_gate_h_u_cla32_and8471_y0(h_u_cla32_and8470_y0, h_u_cla32_and8469_y0, h_u_cla32_and8471_y0);
  and_gate and_gate_h_u_cla32_and8472_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and8472_y0);
  and_gate and_gate_h_u_cla32_and8473_y0(h_u_cla32_and8472_y0, h_u_cla32_and8471_y0, h_u_cla32_and8473_y0);
  and_gate and_gate_h_u_cla32_and8474_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8474_y0);
  and_gate and_gate_h_u_cla32_and8475_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8475_y0);
  and_gate and_gate_h_u_cla32_and8476_y0(h_u_cla32_and8475_y0, h_u_cla32_and8474_y0, h_u_cla32_and8476_y0);
  and_gate and_gate_h_u_cla32_and8477_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8477_y0);
  and_gate and_gate_h_u_cla32_and8478_y0(h_u_cla32_and8477_y0, h_u_cla32_and8476_y0, h_u_cla32_and8478_y0);
  and_gate and_gate_h_u_cla32_and8479_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8479_y0);
  and_gate and_gate_h_u_cla32_and8480_y0(h_u_cla32_and8479_y0, h_u_cla32_and8478_y0, h_u_cla32_and8480_y0);
  and_gate and_gate_h_u_cla32_and8481_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8481_y0);
  and_gate and_gate_h_u_cla32_and8482_y0(h_u_cla32_and8481_y0, h_u_cla32_and8480_y0, h_u_cla32_and8482_y0);
  and_gate and_gate_h_u_cla32_and8483_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8483_y0);
  and_gate and_gate_h_u_cla32_and8484_y0(h_u_cla32_and8483_y0, h_u_cla32_and8482_y0, h_u_cla32_and8484_y0);
  and_gate and_gate_h_u_cla32_and8485_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8485_y0);
  and_gate and_gate_h_u_cla32_and8486_y0(h_u_cla32_and8485_y0, h_u_cla32_and8484_y0, h_u_cla32_and8486_y0);
  and_gate and_gate_h_u_cla32_and8487_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8487_y0);
  and_gate and_gate_h_u_cla32_and8488_y0(h_u_cla32_and8487_y0, h_u_cla32_and8486_y0, h_u_cla32_and8488_y0);
  and_gate and_gate_h_u_cla32_and8489_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and8489_y0);
  and_gate and_gate_h_u_cla32_and8490_y0(h_u_cla32_and8489_y0, h_u_cla32_and8488_y0, h_u_cla32_and8490_y0);
  and_gate and_gate_h_u_cla32_and8491_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8491_y0);
  and_gate and_gate_h_u_cla32_and8492_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8492_y0);
  and_gate and_gate_h_u_cla32_and8493_y0(h_u_cla32_and8492_y0, h_u_cla32_and8491_y0, h_u_cla32_and8493_y0);
  and_gate and_gate_h_u_cla32_and8494_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8494_y0);
  and_gate and_gate_h_u_cla32_and8495_y0(h_u_cla32_and8494_y0, h_u_cla32_and8493_y0, h_u_cla32_and8495_y0);
  and_gate and_gate_h_u_cla32_and8496_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8496_y0);
  and_gate and_gate_h_u_cla32_and8497_y0(h_u_cla32_and8496_y0, h_u_cla32_and8495_y0, h_u_cla32_and8497_y0);
  and_gate and_gate_h_u_cla32_and8498_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8498_y0);
  and_gate and_gate_h_u_cla32_and8499_y0(h_u_cla32_and8498_y0, h_u_cla32_and8497_y0, h_u_cla32_and8499_y0);
  and_gate and_gate_h_u_cla32_and8500_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8500_y0);
  and_gate and_gate_h_u_cla32_and8501_y0(h_u_cla32_and8500_y0, h_u_cla32_and8499_y0, h_u_cla32_and8501_y0);
  and_gate and_gate_h_u_cla32_and8502_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8502_y0);
  and_gate and_gate_h_u_cla32_and8503_y0(h_u_cla32_and8502_y0, h_u_cla32_and8501_y0, h_u_cla32_and8503_y0);
  and_gate and_gate_h_u_cla32_and8504_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and8504_y0);
  and_gate and_gate_h_u_cla32_and8505_y0(h_u_cla32_and8504_y0, h_u_cla32_and8503_y0, h_u_cla32_and8505_y0);
  and_gate and_gate_h_u_cla32_and8506_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8506_y0);
  and_gate and_gate_h_u_cla32_and8507_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8507_y0);
  and_gate and_gate_h_u_cla32_and8508_y0(h_u_cla32_and8507_y0, h_u_cla32_and8506_y0, h_u_cla32_and8508_y0);
  and_gate and_gate_h_u_cla32_and8509_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8509_y0);
  and_gate and_gate_h_u_cla32_and8510_y0(h_u_cla32_and8509_y0, h_u_cla32_and8508_y0, h_u_cla32_and8510_y0);
  and_gate and_gate_h_u_cla32_and8511_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8511_y0);
  and_gate and_gate_h_u_cla32_and8512_y0(h_u_cla32_and8511_y0, h_u_cla32_and8510_y0, h_u_cla32_and8512_y0);
  and_gate and_gate_h_u_cla32_and8513_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8513_y0);
  and_gate and_gate_h_u_cla32_and8514_y0(h_u_cla32_and8513_y0, h_u_cla32_and8512_y0, h_u_cla32_and8514_y0);
  and_gate and_gate_h_u_cla32_and8515_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8515_y0);
  and_gate and_gate_h_u_cla32_and8516_y0(h_u_cla32_and8515_y0, h_u_cla32_and8514_y0, h_u_cla32_and8516_y0);
  and_gate and_gate_h_u_cla32_and8517_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and8517_y0);
  and_gate and_gate_h_u_cla32_and8518_y0(h_u_cla32_and8517_y0, h_u_cla32_and8516_y0, h_u_cla32_and8518_y0);
  and_gate and_gate_h_u_cla32_and8519_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and8519_y0);
  and_gate and_gate_h_u_cla32_and8520_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and8520_y0);
  and_gate and_gate_h_u_cla32_and8521_y0(h_u_cla32_and8520_y0, h_u_cla32_and8519_y0, h_u_cla32_and8521_y0);
  and_gate and_gate_h_u_cla32_and8522_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and8522_y0);
  and_gate and_gate_h_u_cla32_and8523_y0(h_u_cla32_and8522_y0, h_u_cla32_and8521_y0, h_u_cla32_and8523_y0);
  and_gate and_gate_h_u_cla32_and8524_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and8524_y0);
  and_gate and_gate_h_u_cla32_and8525_y0(h_u_cla32_and8524_y0, h_u_cla32_and8523_y0, h_u_cla32_and8525_y0);
  and_gate and_gate_h_u_cla32_and8526_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and8526_y0);
  and_gate and_gate_h_u_cla32_and8527_y0(h_u_cla32_and8526_y0, h_u_cla32_and8525_y0, h_u_cla32_and8527_y0);
  and_gate and_gate_h_u_cla32_and8528_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and8528_y0);
  and_gate and_gate_h_u_cla32_and8529_y0(h_u_cla32_and8528_y0, h_u_cla32_and8527_y0, h_u_cla32_and8529_y0);
  and_gate and_gate_h_u_cla32_and8530_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and8530_y0);
  and_gate and_gate_h_u_cla32_and8531_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and8531_y0);
  and_gate and_gate_h_u_cla32_and8532_y0(h_u_cla32_and8531_y0, h_u_cla32_and8530_y0, h_u_cla32_and8532_y0);
  and_gate and_gate_h_u_cla32_and8533_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and8533_y0);
  and_gate and_gate_h_u_cla32_and8534_y0(h_u_cla32_and8533_y0, h_u_cla32_and8532_y0, h_u_cla32_and8534_y0);
  and_gate and_gate_h_u_cla32_and8535_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and8535_y0);
  and_gate and_gate_h_u_cla32_and8536_y0(h_u_cla32_and8535_y0, h_u_cla32_and8534_y0, h_u_cla32_and8536_y0);
  and_gate and_gate_h_u_cla32_and8537_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and8537_y0);
  and_gate and_gate_h_u_cla32_and8538_y0(h_u_cla32_and8537_y0, h_u_cla32_and8536_y0, h_u_cla32_and8538_y0);
  and_gate and_gate_h_u_cla32_and8539_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and8539_y0);
  and_gate and_gate_h_u_cla32_and8540_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and8540_y0);
  and_gate and_gate_h_u_cla32_and8541_y0(h_u_cla32_and8540_y0, h_u_cla32_and8539_y0, h_u_cla32_and8541_y0);
  and_gate and_gate_h_u_cla32_and8542_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and8542_y0);
  and_gate and_gate_h_u_cla32_and8543_y0(h_u_cla32_and8542_y0, h_u_cla32_and8541_y0, h_u_cla32_and8543_y0);
  and_gate and_gate_h_u_cla32_and8544_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and8544_y0);
  and_gate and_gate_h_u_cla32_and8545_y0(h_u_cla32_and8544_y0, h_u_cla32_and8543_y0, h_u_cla32_and8545_y0);
  and_gate and_gate_h_u_cla32_and8546_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and8546_y0);
  and_gate and_gate_h_u_cla32_and8547_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and8547_y0);
  and_gate and_gate_h_u_cla32_and8548_y0(h_u_cla32_and8547_y0, h_u_cla32_and8546_y0, h_u_cla32_and8548_y0);
  and_gate and_gate_h_u_cla32_and8549_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and8549_y0);
  and_gate and_gate_h_u_cla32_and8550_y0(h_u_cla32_and8549_y0, h_u_cla32_and8548_y0, h_u_cla32_and8550_y0);
  and_gate and_gate_h_u_cla32_and8551_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and8551_y0);
  and_gate and_gate_h_u_cla32_and8552_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and8552_y0);
  and_gate and_gate_h_u_cla32_and8553_y0(h_u_cla32_and8552_y0, h_u_cla32_and8551_y0, h_u_cla32_and8553_y0);
  and_gate and_gate_h_u_cla32_and8554_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and8554_y0);
  or_gate or_gate_h_u_cla32_or406_y0(h_u_cla32_and8554_y0, h_u_cla32_and7770_y0, h_u_cla32_or406_y0);
  or_gate or_gate_h_u_cla32_or407_y0(h_u_cla32_or406_y0, h_u_cla32_and7825_y0, h_u_cla32_or407_y0);
  or_gate or_gate_h_u_cla32_or408_y0(h_u_cla32_or407_y0, h_u_cla32_and7878_y0, h_u_cla32_or408_y0);
  or_gate or_gate_h_u_cla32_or409_y0(h_u_cla32_or408_y0, h_u_cla32_and7929_y0, h_u_cla32_or409_y0);
  or_gate or_gate_h_u_cla32_or410_y0(h_u_cla32_or409_y0, h_u_cla32_and7978_y0, h_u_cla32_or410_y0);
  or_gate or_gate_h_u_cla32_or411_y0(h_u_cla32_or410_y0, h_u_cla32_and8025_y0, h_u_cla32_or411_y0);
  or_gate or_gate_h_u_cla32_or412_y0(h_u_cla32_or411_y0, h_u_cla32_and8070_y0, h_u_cla32_or412_y0);
  or_gate or_gate_h_u_cla32_or413_y0(h_u_cla32_or412_y0, h_u_cla32_and8113_y0, h_u_cla32_or413_y0);
  or_gate or_gate_h_u_cla32_or414_y0(h_u_cla32_or413_y0, h_u_cla32_and8154_y0, h_u_cla32_or414_y0);
  or_gate or_gate_h_u_cla32_or415_y0(h_u_cla32_or414_y0, h_u_cla32_and8193_y0, h_u_cla32_or415_y0);
  or_gate or_gate_h_u_cla32_or416_y0(h_u_cla32_or415_y0, h_u_cla32_and8230_y0, h_u_cla32_or416_y0);
  or_gate or_gate_h_u_cla32_or417_y0(h_u_cla32_or416_y0, h_u_cla32_and8265_y0, h_u_cla32_or417_y0);
  or_gate or_gate_h_u_cla32_or418_y0(h_u_cla32_or417_y0, h_u_cla32_and8298_y0, h_u_cla32_or418_y0);
  or_gate or_gate_h_u_cla32_or419_y0(h_u_cla32_or418_y0, h_u_cla32_and8329_y0, h_u_cla32_or419_y0);
  or_gate or_gate_h_u_cla32_or420_y0(h_u_cla32_or419_y0, h_u_cla32_and8358_y0, h_u_cla32_or420_y0);
  or_gate or_gate_h_u_cla32_or421_y0(h_u_cla32_or420_y0, h_u_cla32_and8385_y0, h_u_cla32_or421_y0);
  or_gate or_gate_h_u_cla32_or422_y0(h_u_cla32_or421_y0, h_u_cla32_and8410_y0, h_u_cla32_or422_y0);
  or_gate or_gate_h_u_cla32_or423_y0(h_u_cla32_or422_y0, h_u_cla32_and8433_y0, h_u_cla32_or423_y0);
  or_gate or_gate_h_u_cla32_or424_y0(h_u_cla32_or423_y0, h_u_cla32_and8454_y0, h_u_cla32_or424_y0);
  or_gate or_gate_h_u_cla32_or425_y0(h_u_cla32_or424_y0, h_u_cla32_and8473_y0, h_u_cla32_or425_y0);
  or_gate or_gate_h_u_cla32_or426_y0(h_u_cla32_or425_y0, h_u_cla32_and8490_y0, h_u_cla32_or426_y0);
  or_gate or_gate_h_u_cla32_or427_y0(h_u_cla32_or426_y0, h_u_cla32_and8505_y0, h_u_cla32_or427_y0);
  or_gate or_gate_h_u_cla32_or428_y0(h_u_cla32_or427_y0, h_u_cla32_and8518_y0, h_u_cla32_or428_y0);
  or_gate or_gate_h_u_cla32_or429_y0(h_u_cla32_or428_y0, h_u_cla32_and8529_y0, h_u_cla32_or429_y0);
  or_gate or_gate_h_u_cla32_or430_y0(h_u_cla32_or429_y0, h_u_cla32_and8538_y0, h_u_cla32_or430_y0);
  or_gate or_gate_h_u_cla32_or431_y0(h_u_cla32_or430_y0, h_u_cla32_and8545_y0, h_u_cla32_or431_y0);
  or_gate or_gate_h_u_cla32_or432_y0(h_u_cla32_or431_y0, h_u_cla32_and8550_y0, h_u_cla32_or432_y0);
  or_gate or_gate_h_u_cla32_or433_y0(h_u_cla32_or432_y0, h_u_cla32_and8553_y0, h_u_cla32_or433_y0);
  or_gate or_gate_h_u_cla32_or434_y0(h_u_cla32_pg_logic28_y1, h_u_cla32_or433_y0, h_u_cla32_or434_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic29_y0(a_29, b_29, h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic29_y1, h_u_cla32_pg_logic29_y2);
  xor_gate xor_gate_h_u_cla32_xor29_y0(h_u_cla32_pg_logic29_y2, h_u_cla32_or434_y0, h_u_cla32_xor29_y0);
  and_gate and_gate_h_u_cla32_and8555_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and8555_y0);
  and_gate and_gate_h_u_cla32_and8556_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and8556_y0);
  and_gate and_gate_h_u_cla32_and8557_y0(h_u_cla32_and8556_y0, h_u_cla32_and8555_y0, h_u_cla32_and8557_y0);
  and_gate and_gate_h_u_cla32_and8558_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and8558_y0);
  and_gate and_gate_h_u_cla32_and8559_y0(h_u_cla32_and8558_y0, h_u_cla32_and8557_y0, h_u_cla32_and8559_y0);
  and_gate and_gate_h_u_cla32_and8560_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and8560_y0);
  and_gate and_gate_h_u_cla32_and8561_y0(h_u_cla32_and8560_y0, h_u_cla32_and8559_y0, h_u_cla32_and8561_y0);
  and_gate and_gate_h_u_cla32_and8562_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and8562_y0);
  and_gate and_gate_h_u_cla32_and8563_y0(h_u_cla32_and8562_y0, h_u_cla32_and8561_y0, h_u_cla32_and8563_y0);
  and_gate and_gate_h_u_cla32_and8564_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and8564_y0);
  and_gate and_gate_h_u_cla32_and8565_y0(h_u_cla32_and8564_y0, h_u_cla32_and8563_y0, h_u_cla32_and8565_y0);
  and_gate and_gate_h_u_cla32_and8566_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and8566_y0);
  and_gate and_gate_h_u_cla32_and8567_y0(h_u_cla32_and8566_y0, h_u_cla32_and8565_y0, h_u_cla32_and8567_y0);
  and_gate and_gate_h_u_cla32_and8568_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and8568_y0);
  and_gate and_gate_h_u_cla32_and8569_y0(h_u_cla32_and8568_y0, h_u_cla32_and8567_y0, h_u_cla32_and8569_y0);
  and_gate and_gate_h_u_cla32_and8570_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and8570_y0);
  and_gate and_gate_h_u_cla32_and8571_y0(h_u_cla32_and8570_y0, h_u_cla32_and8569_y0, h_u_cla32_and8571_y0);
  and_gate and_gate_h_u_cla32_and8572_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and8572_y0);
  and_gate and_gate_h_u_cla32_and8573_y0(h_u_cla32_and8572_y0, h_u_cla32_and8571_y0, h_u_cla32_and8573_y0);
  and_gate and_gate_h_u_cla32_and8574_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and8574_y0);
  and_gate and_gate_h_u_cla32_and8575_y0(h_u_cla32_and8574_y0, h_u_cla32_and8573_y0, h_u_cla32_and8575_y0);
  and_gate and_gate_h_u_cla32_and8576_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and8576_y0);
  and_gate and_gate_h_u_cla32_and8577_y0(h_u_cla32_and8576_y0, h_u_cla32_and8575_y0, h_u_cla32_and8577_y0);
  and_gate and_gate_h_u_cla32_and8578_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and8578_y0);
  and_gate and_gate_h_u_cla32_and8579_y0(h_u_cla32_and8578_y0, h_u_cla32_and8577_y0, h_u_cla32_and8579_y0);
  and_gate and_gate_h_u_cla32_and8580_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and8580_y0);
  and_gate and_gate_h_u_cla32_and8581_y0(h_u_cla32_and8580_y0, h_u_cla32_and8579_y0, h_u_cla32_and8581_y0);
  and_gate and_gate_h_u_cla32_and8582_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and8582_y0);
  and_gate and_gate_h_u_cla32_and8583_y0(h_u_cla32_and8582_y0, h_u_cla32_and8581_y0, h_u_cla32_and8583_y0);
  and_gate and_gate_h_u_cla32_and8584_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and8584_y0);
  and_gate and_gate_h_u_cla32_and8585_y0(h_u_cla32_and8584_y0, h_u_cla32_and8583_y0, h_u_cla32_and8585_y0);
  and_gate and_gate_h_u_cla32_and8586_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and8586_y0);
  and_gate and_gate_h_u_cla32_and8587_y0(h_u_cla32_and8586_y0, h_u_cla32_and8585_y0, h_u_cla32_and8587_y0);
  and_gate and_gate_h_u_cla32_and8588_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and8588_y0);
  and_gate and_gate_h_u_cla32_and8589_y0(h_u_cla32_and8588_y0, h_u_cla32_and8587_y0, h_u_cla32_and8589_y0);
  and_gate and_gate_h_u_cla32_and8590_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and8590_y0);
  and_gate and_gate_h_u_cla32_and8591_y0(h_u_cla32_and8590_y0, h_u_cla32_and8589_y0, h_u_cla32_and8591_y0);
  and_gate and_gate_h_u_cla32_and8592_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and8592_y0);
  and_gate and_gate_h_u_cla32_and8593_y0(h_u_cla32_and8592_y0, h_u_cla32_and8591_y0, h_u_cla32_and8593_y0);
  and_gate and_gate_h_u_cla32_and8594_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and8594_y0);
  and_gate and_gate_h_u_cla32_and8595_y0(h_u_cla32_and8594_y0, h_u_cla32_and8593_y0, h_u_cla32_and8595_y0);
  and_gate and_gate_h_u_cla32_and8596_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and8596_y0);
  and_gate and_gate_h_u_cla32_and8597_y0(h_u_cla32_and8596_y0, h_u_cla32_and8595_y0, h_u_cla32_and8597_y0);
  and_gate and_gate_h_u_cla32_and8598_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and8598_y0);
  and_gate and_gate_h_u_cla32_and8599_y0(h_u_cla32_and8598_y0, h_u_cla32_and8597_y0, h_u_cla32_and8599_y0);
  and_gate and_gate_h_u_cla32_and8600_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and8600_y0);
  and_gate and_gate_h_u_cla32_and8601_y0(h_u_cla32_and8600_y0, h_u_cla32_and8599_y0, h_u_cla32_and8601_y0);
  and_gate and_gate_h_u_cla32_and8602_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and8602_y0);
  and_gate and_gate_h_u_cla32_and8603_y0(h_u_cla32_and8602_y0, h_u_cla32_and8601_y0, h_u_cla32_and8603_y0);
  and_gate and_gate_h_u_cla32_and8604_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and8604_y0);
  and_gate and_gate_h_u_cla32_and8605_y0(h_u_cla32_and8604_y0, h_u_cla32_and8603_y0, h_u_cla32_and8605_y0);
  and_gate and_gate_h_u_cla32_and8606_y0(h_u_cla32_pg_logic26_y0, constant_wire_0, h_u_cla32_and8606_y0);
  and_gate and_gate_h_u_cla32_and8607_y0(h_u_cla32_and8606_y0, h_u_cla32_and8605_y0, h_u_cla32_and8607_y0);
  and_gate and_gate_h_u_cla32_and8608_y0(h_u_cla32_pg_logic27_y0, constant_wire_0, h_u_cla32_and8608_y0);
  and_gate and_gate_h_u_cla32_and8609_y0(h_u_cla32_and8608_y0, h_u_cla32_and8607_y0, h_u_cla32_and8609_y0);
  and_gate and_gate_h_u_cla32_and8610_y0(h_u_cla32_pg_logic28_y0, constant_wire_0, h_u_cla32_and8610_y0);
  and_gate and_gate_h_u_cla32_and8611_y0(h_u_cla32_and8610_y0, h_u_cla32_and8609_y0, h_u_cla32_and8611_y0);
  and_gate and_gate_h_u_cla32_and8612_y0(h_u_cla32_pg_logic29_y0, constant_wire_0, h_u_cla32_and8612_y0);
  and_gate and_gate_h_u_cla32_and8613_y0(h_u_cla32_and8612_y0, h_u_cla32_and8611_y0, h_u_cla32_and8613_y0);
  and_gate and_gate_h_u_cla32_and8614_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8614_y0);
  and_gate and_gate_h_u_cla32_and8615_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8615_y0);
  and_gate and_gate_h_u_cla32_and8616_y0(h_u_cla32_and8615_y0, h_u_cla32_and8614_y0, h_u_cla32_and8616_y0);
  and_gate and_gate_h_u_cla32_and8617_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8617_y0);
  and_gate and_gate_h_u_cla32_and8618_y0(h_u_cla32_and8617_y0, h_u_cla32_and8616_y0, h_u_cla32_and8618_y0);
  and_gate and_gate_h_u_cla32_and8619_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8619_y0);
  and_gate and_gate_h_u_cla32_and8620_y0(h_u_cla32_and8619_y0, h_u_cla32_and8618_y0, h_u_cla32_and8620_y0);
  and_gate and_gate_h_u_cla32_and8621_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8621_y0);
  and_gate and_gate_h_u_cla32_and8622_y0(h_u_cla32_and8621_y0, h_u_cla32_and8620_y0, h_u_cla32_and8622_y0);
  and_gate and_gate_h_u_cla32_and8623_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8623_y0);
  and_gate and_gate_h_u_cla32_and8624_y0(h_u_cla32_and8623_y0, h_u_cla32_and8622_y0, h_u_cla32_and8624_y0);
  and_gate and_gate_h_u_cla32_and8625_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8625_y0);
  and_gate and_gate_h_u_cla32_and8626_y0(h_u_cla32_and8625_y0, h_u_cla32_and8624_y0, h_u_cla32_and8626_y0);
  and_gate and_gate_h_u_cla32_and8627_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8627_y0);
  and_gate and_gate_h_u_cla32_and8628_y0(h_u_cla32_and8627_y0, h_u_cla32_and8626_y0, h_u_cla32_and8628_y0);
  and_gate and_gate_h_u_cla32_and8629_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8629_y0);
  and_gate and_gate_h_u_cla32_and8630_y0(h_u_cla32_and8629_y0, h_u_cla32_and8628_y0, h_u_cla32_and8630_y0);
  and_gate and_gate_h_u_cla32_and8631_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8631_y0);
  and_gate and_gate_h_u_cla32_and8632_y0(h_u_cla32_and8631_y0, h_u_cla32_and8630_y0, h_u_cla32_and8632_y0);
  and_gate and_gate_h_u_cla32_and8633_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8633_y0);
  and_gate and_gate_h_u_cla32_and8634_y0(h_u_cla32_and8633_y0, h_u_cla32_and8632_y0, h_u_cla32_and8634_y0);
  and_gate and_gate_h_u_cla32_and8635_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8635_y0);
  and_gate and_gate_h_u_cla32_and8636_y0(h_u_cla32_and8635_y0, h_u_cla32_and8634_y0, h_u_cla32_and8636_y0);
  and_gate and_gate_h_u_cla32_and8637_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8637_y0);
  and_gate and_gate_h_u_cla32_and8638_y0(h_u_cla32_and8637_y0, h_u_cla32_and8636_y0, h_u_cla32_and8638_y0);
  and_gate and_gate_h_u_cla32_and8639_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8639_y0);
  and_gate and_gate_h_u_cla32_and8640_y0(h_u_cla32_and8639_y0, h_u_cla32_and8638_y0, h_u_cla32_and8640_y0);
  and_gate and_gate_h_u_cla32_and8641_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8641_y0);
  and_gate and_gate_h_u_cla32_and8642_y0(h_u_cla32_and8641_y0, h_u_cla32_and8640_y0, h_u_cla32_and8642_y0);
  and_gate and_gate_h_u_cla32_and8643_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8643_y0);
  and_gate and_gate_h_u_cla32_and8644_y0(h_u_cla32_and8643_y0, h_u_cla32_and8642_y0, h_u_cla32_and8644_y0);
  and_gate and_gate_h_u_cla32_and8645_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8645_y0);
  and_gate and_gate_h_u_cla32_and8646_y0(h_u_cla32_and8645_y0, h_u_cla32_and8644_y0, h_u_cla32_and8646_y0);
  and_gate and_gate_h_u_cla32_and8647_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8647_y0);
  and_gate and_gate_h_u_cla32_and8648_y0(h_u_cla32_and8647_y0, h_u_cla32_and8646_y0, h_u_cla32_and8648_y0);
  and_gate and_gate_h_u_cla32_and8649_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8649_y0);
  and_gate and_gate_h_u_cla32_and8650_y0(h_u_cla32_and8649_y0, h_u_cla32_and8648_y0, h_u_cla32_and8650_y0);
  and_gate and_gate_h_u_cla32_and8651_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8651_y0);
  and_gate and_gate_h_u_cla32_and8652_y0(h_u_cla32_and8651_y0, h_u_cla32_and8650_y0, h_u_cla32_and8652_y0);
  and_gate and_gate_h_u_cla32_and8653_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8653_y0);
  and_gate and_gate_h_u_cla32_and8654_y0(h_u_cla32_and8653_y0, h_u_cla32_and8652_y0, h_u_cla32_and8654_y0);
  and_gate and_gate_h_u_cla32_and8655_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8655_y0);
  and_gate and_gate_h_u_cla32_and8656_y0(h_u_cla32_and8655_y0, h_u_cla32_and8654_y0, h_u_cla32_and8656_y0);
  and_gate and_gate_h_u_cla32_and8657_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8657_y0);
  and_gate and_gate_h_u_cla32_and8658_y0(h_u_cla32_and8657_y0, h_u_cla32_and8656_y0, h_u_cla32_and8658_y0);
  and_gate and_gate_h_u_cla32_and8659_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8659_y0);
  and_gate and_gate_h_u_cla32_and8660_y0(h_u_cla32_and8659_y0, h_u_cla32_and8658_y0, h_u_cla32_and8660_y0);
  and_gate and_gate_h_u_cla32_and8661_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8661_y0);
  and_gate and_gate_h_u_cla32_and8662_y0(h_u_cla32_and8661_y0, h_u_cla32_and8660_y0, h_u_cla32_and8662_y0);
  and_gate and_gate_h_u_cla32_and8663_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8663_y0);
  and_gate and_gate_h_u_cla32_and8664_y0(h_u_cla32_and8663_y0, h_u_cla32_and8662_y0, h_u_cla32_and8664_y0);
  and_gate and_gate_h_u_cla32_and8665_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8665_y0);
  and_gate and_gate_h_u_cla32_and8666_y0(h_u_cla32_and8665_y0, h_u_cla32_and8664_y0, h_u_cla32_and8666_y0);
  and_gate and_gate_h_u_cla32_and8667_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8667_y0);
  and_gate and_gate_h_u_cla32_and8668_y0(h_u_cla32_and8667_y0, h_u_cla32_and8666_y0, h_u_cla32_and8668_y0);
  and_gate and_gate_h_u_cla32_and8669_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and8669_y0);
  and_gate and_gate_h_u_cla32_and8670_y0(h_u_cla32_and8669_y0, h_u_cla32_and8668_y0, h_u_cla32_and8670_y0);
  and_gate and_gate_h_u_cla32_and8671_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8671_y0);
  and_gate and_gate_h_u_cla32_and8672_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8672_y0);
  and_gate and_gate_h_u_cla32_and8673_y0(h_u_cla32_and8672_y0, h_u_cla32_and8671_y0, h_u_cla32_and8673_y0);
  and_gate and_gate_h_u_cla32_and8674_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8674_y0);
  and_gate and_gate_h_u_cla32_and8675_y0(h_u_cla32_and8674_y0, h_u_cla32_and8673_y0, h_u_cla32_and8675_y0);
  and_gate and_gate_h_u_cla32_and8676_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8676_y0);
  and_gate and_gate_h_u_cla32_and8677_y0(h_u_cla32_and8676_y0, h_u_cla32_and8675_y0, h_u_cla32_and8677_y0);
  and_gate and_gate_h_u_cla32_and8678_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8678_y0);
  and_gate and_gate_h_u_cla32_and8679_y0(h_u_cla32_and8678_y0, h_u_cla32_and8677_y0, h_u_cla32_and8679_y0);
  and_gate and_gate_h_u_cla32_and8680_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8680_y0);
  and_gate and_gate_h_u_cla32_and8681_y0(h_u_cla32_and8680_y0, h_u_cla32_and8679_y0, h_u_cla32_and8681_y0);
  and_gate and_gate_h_u_cla32_and8682_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8682_y0);
  and_gate and_gate_h_u_cla32_and8683_y0(h_u_cla32_and8682_y0, h_u_cla32_and8681_y0, h_u_cla32_and8683_y0);
  and_gate and_gate_h_u_cla32_and8684_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8684_y0);
  and_gate and_gate_h_u_cla32_and8685_y0(h_u_cla32_and8684_y0, h_u_cla32_and8683_y0, h_u_cla32_and8685_y0);
  and_gate and_gate_h_u_cla32_and8686_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8686_y0);
  and_gate and_gate_h_u_cla32_and8687_y0(h_u_cla32_and8686_y0, h_u_cla32_and8685_y0, h_u_cla32_and8687_y0);
  and_gate and_gate_h_u_cla32_and8688_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8688_y0);
  and_gate and_gate_h_u_cla32_and8689_y0(h_u_cla32_and8688_y0, h_u_cla32_and8687_y0, h_u_cla32_and8689_y0);
  and_gate and_gate_h_u_cla32_and8690_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8690_y0);
  and_gate and_gate_h_u_cla32_and8691_y0(h_u_cla32_and8690_y0, h_u_cla32_and8689_y0, h_u_cla32_and8691_y0);
  and_gate and_gate_h_u_cla32_and8692_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8692_y0);
  and_gate and_gate_h_u_cla32_and8693_y0(h_u_cla32_and8692_y0, h_u_cla32_and8691_y0, h_u_cla32_and8693_y0);
  and_gate and_gate_h_u_cla32_and8694_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8694_y0);
  and_gate and_gate_h_u_cla32_and8695_y0(h_u_cla32_and8694_y0, h_u_cla32_and8693_y0, h_u_cla32_and8695_y0);
  and_gate and_gate_h_u_cla32_and8696_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8696_y0);
  and_gate and_gate_h_u_cla32_and8697_y0(h_u_cla32_and8696_y0, h_u_cla32_and8695_y0, h_u_cla32_and8697_y0);
  and_gate and_gate_h_u_cla32_and8698_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8698_y0);
  and_gate and_gate_h_u_cla32_and8699_y0(h_u_cla32_and8698_y0, h_u_cla32_and8697_y0, h_u_cla32_and8699_y0);
  and_gate and_gate_h_u_cla32_and8700_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8700_y0);
  and_gate and_gate_h_u_cla32_and8701_y0(h_u_cla32_and8700_y0, h_u_cla32_and8699_y0, h_u_cla32_and8701_y0);
  and_gate and_gate_h_u_cla32_and8702_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8702_y0);
  and_gate and_gate_h_u_cla32_and8703_y0(h_u_cla32_and8702_y0, h_u_cla32_and8701_y0, h_u_cla32_and8703_y0);
  and_gate and_gate_h_u_cla32_and8704_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8704_y0);
  and_gate and_gate_h_u_cla32_and8705_y0(h_u_cla32_and8704_y0, h_u_cla32_and8703_y0, h_u_cla32_and8705_y0);
  and_gate and_gate_h_u_cla32_and8706_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8706_y0);
  and_gate and_gate_h_u_cla32_and8707_y0(h_u_cla32_and8706_y0, h_u_cla32_and8705_y0, h_u_cla32_and8707_y0);
  and_gate and_gate_h_u_cla32_and8708_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8708_y0);
  and_gate and_gate_h_u_cla32_and8709_y0(h_u_cla32_and8708_y0, h_u_cla32_and8707_y0, h_u_cla32_and8709_y0);
  and_gate and_gate_h_u_cla32_and8710_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8710_y0);
  and_gate and_gate_h_u_cla32_and8711_y0(h_u_cla32_and8710_y0, h_u_cla32_and8709_y0, h_u_cla32_and8711_y0);
  and_gate and_gate_h_u_cla32_and8712_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8712_y0);
  and_gate and_gate_h_u_cla32_and8713_y0(h_u_cla32_and8712_y0, h_u_cla32_and8711_y0, h_u_cla32_and8713_y0);
  and_gate and_gate_h_u_cla32_and8714_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8714_y0);
  and_gate and_gate_h_u_cla32_and8715_y0(h_u_cla32_and8714_y0, h_u_cla32_and8713_y0, h_u_cla32_and8715_y0);
  and_gate and_gate_h_u_cla32_and8716_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8716_y0);
  and_gate and_gate_h_u_cla32_and8717_y0(h_u_cla32_and8716_y0, h_u_cla32_and8715_y0, h_u_cla32_and8717_y0);
  and_gate and_gate_h_u_cla32_and8718_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8718_y0);
  and_gate and_gate_h_u_cla32_and8719_y0(h_u_cla32_and8718_y0, h_u_cla32_and8717_y0, h_u_cla32_and8719_y0);
  and_gate and_gate_h_u_cla32_and8720_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8720_y0);
  and_gate and_gate_h_u_cla32_and8721_y0(h_u_cla32_and8720_y0, h_u_cla32_and8719_y0, h_u_cla32_and8721_y0);
  and_gate and_gate_h_u_cla32_and8722_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8722_y0);
  and_gate and_gate_h_u_cla32_and8723_y0(h_u_cla32_and8722_y0, h_u_cla32_and8721_y0, h_u_cla32_and8723_y0);
  and_gate and_gate_h_u_cla32_and8724_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and8724_y0);
  and_gate and_gate_h_u_cla32_and8725_y0(h_u_cla32_and8724_y0, h_u_cla32_and8723_y0, h_u_cla32_and8725_y0);
  and_gate and_gate_h_u_cla32_and8726_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8726_y0);
  and_gate and_gate_h_u_cla32_and8727_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8727_y0);
  and_gate and_gate_h_u_cla32_and8728_y0(h_u_cla32_and8727_y0, h_u_cla32_and8726_y0, h_u_cla32_and8728_y0);
  and_gate and_gate_h_u_cla32_and8729_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8729_y0);
  and_gate and_gate_h_u_cla32_and8730_y0(h_u_cla32_and8729_y0, h_u_cla32_and8728_y0, h_u_cla32_and8730_y0);
  and_gate and_gate_h_u_cla32_and8731_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8731_y0);
  and_gate and_gate_h_u_cla32_and8732_y0(h_u_cla32_and8731_y0, h_u_cla32_and8730_y0, h_u_cla32_and8732_y0);
  and_gate and_gate_h_u_cla32_and8733_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8733_y0);
  and_gate and_gate_h_u_cla32_and8734_y0(h_u_cla32_and8733_y0, h_u_cla32_and8732_y0, h_u_cla32_and8734_y0);
  and_gate and_gate_h_u_cla32_and8735_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8735_y0);
  and_gate and_gate_h_u_cla32_and8736_y0(h_u_cla32_and8735_y0, h_u_cla32_and8734_y0, h_u_cla32_and8736_y0);
  and_gate and_gate_h_u_cla32_and8737_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8737_y0);
  and_gate and_gate_h_u_cla32_and8738_y0(h_u_cla32_and8737_y0, h_u_cla32_and8736_y0, h_u_cla32_and8738_y0);
  and_gate and_gate_h_u_cla32_and8739_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8739_y0);
  and_gate and_gate_h_u_cla32_and8740_y0(h_u_cla32_and8739_y0, h_u_cla32_and8738_y0, h_u_cla32_and8740_y0);
  and_gate and_gate_h_u_cla32_and8741_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8741_y0);
  and_gate and_gate_h_u_cla32_and8742_y0(h_u_cla32_and8741_y0, h_u_cla32_and8740_y0, h_u_cla32_and8742_y0);
  and_gate and_gate_h_u_cla32_and8743_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8743_y0);
  and_gate and_gate_h_u_cla32_and8744_y0(h_u_cla32_and8743_y0, h_u_cla32_and8742_y0, h_u_cla32_and8744_y0);
  and_gate and_gate_h_u_cla32_and8745_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8745_y0);
  and_gate and_gate_h_u_cla32_and8746_y0(h_u_cla32_and8745_y0, h_u_cla32_and8744_y0, h_u_cla32_and8746_y0);
  and_gate and_gate_h_u_cla32_and8747_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8747_y0);
  and_gate and_gate_h_u_cla32_and8748_y0(h_u_cla32_and8747_y0, h_u_cla32_and8746_y0, h_u_cla32_and8748_y0);
  and_gate and_gate_h_u_cla32_and8749_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8749_y0);
  and_gate and_gate_h_u_cla32_and8750_y0(h_u_cla32_and8749_y0, h_u_cla32_and8748_y0, h_u_cla32_and8750_y0);
  and_gate and_gate_h_u_cla32_and8751_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8751_y0);
  and_gate and_gate_h_u_cla32_and8752_y0(h_u_cla32_and8751_y0, h_u_cla32_and8750_y0, h_u_cla32_and8752_y0);
  and_gate and_gate_h_u_cla32_and8753_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8753_y0);
  and_gate and_gate_h_u_cla32_and8754_y0(h_u_cla32_and8753_y0, h_u_cla32_and8752_y0, h_u_cla32_and8754_y0);
  and_gate and_gate_h_u_cla32_and8755_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8755_y0);
  and_gate and_gate_h_u_cla32_and8756_y0(h_u_cla32_and8755_y0, h_u_cla32_and8754_y0, h_u_cla32_and8756_y0);
  and_gate and_gate_h_u_cla32_and8757_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8757_y0);
  and_gate and_gate_h_u_cla32_and8758_y0(h_u_cla32_and8757_y0, h_u_cla32_and8756_y0, h_u_cla32_and8758_y0);
  and_gate and_gate_h_u_cla32_and8759_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8759_y0);
  and_gate and_gate_h_u_cla32_and8760_y0(h_u_cla32_and8759_y0, h_u_cla32_and8758_y0, h_u_cla32_and8760_y0);
  and_gate and_gate_h_u_cla32_and8761_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8761_y0);
  and_gate and_gate_h_u_cla32_and8762_y0(h_u_cla32_and8761_y0, h_u_cla32_and8760_y0, h_u_cla32_and8762_y0);
  and_gate and_gate_h_u_cla32_and8763_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8763_y0);
  and_gate and_gate_h_u_cla32_and8764_y0(h_u_cla32_and8763_y0, h_u_cla32_and8762_y0, h_u_cla32_and8764_y0);
  and_gate and_gate_h_u_cla32_and8765_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8765_y0);
  and_gate and_gate_h_u_cla32_and8766_y0(h_u_cla32_and8765_y0, h_u_cla32_and8764_y0, h_u_cla32_and8766_y0);
  and_gate and_gate_h_u_cla32_and8767_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8767_y0);
  and_gate and_gate_h_u_cla32_and8768_y0(h_u_cla32_and8767_y0, h_u_cla32_and8766_y0, h_u_cla32_and8768_y0);
  and_gate and_gate_h_u_cla32_and8769_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8769_y0);
  and_gate and_gate_h_u_cla32_and8770_y0(h_u_cla32_and8769_y0, h_u_cla32_and8768_y0, h_u_cla32_and8770_y0);
  and_gate and_gate_h_u_cla32_and8771_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8771_y0);
  and_gate and_gate_h_u_cla32_and8772_y0(h_u_cla32_and8771_y0, h_u_cla32_and8770_y0, h_u_cla32_and8772_y0);
  and_gate and_gate_h_u_cla32_and8773_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8773_y0);
  and_gate and_gate_h_u_cla32_and8774_y0(h_u_cla32_and8773_y0, h_u_cla32_and8772_y0, h_u_cla32_and8774_y0);
  and_gate and_gate_h_u_cla32_and8775_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8775_y0);
  and_gate and_gate_h_u_cla32_and8776_y0(h_u_cla32_and8775_y0, h_u_cla32_and8774_y0, h_u_cla32_and8776_y0);
  and_gate and_gate_h_u_cla32_and8777_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and8777_y0);
  and_gate and_gate_h_u_cla32_and8778_y0(h_u_cla32_and8777_y0, h_u_cla32_and8776_y0, h_u_cla32_and8778_y0);
  and_gate and_gate_h_u_cla32_and8779_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8779_y0);
  and_gate and_gate_h_u_cla32_and8780_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8780_y0);
  and_gate and_gate_h_u_cla32_and8781_y0(h_u_cla32_and8780_y0, h_u_cla32_and8779_y0, h_u_cla32_and8781_y0);
  and_gate and_gate_h_u_cla32_and8782_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8782_y0);
  and_gate and_gate_h_u_cla32_and8783_y0(h_u_cla32_and8782_y0, h_u_cla32_and8781_y0, h_u_cla32_and8783_y0);
  and_gate and_gate_h_u_cla32_and8784_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8784_y0);
  and_gate and_gate_h_u_cla32_and8785_y0(h_u_cla32_and8784_y0, h_u_cla32_and8783_y0, h_u_cla32_and8785_y0);
  and_gate and_gate_h_u_cla32_and8786_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8786_y0);
  and_gate and_gate_h_u_cla32_and8787_y0(h_u_cla32_and8786_y0, h_u_cla32_and8785_y0, h_u_cla32_and8787_y0);
  and_gate and_gate_h_u_cla32_and8788_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8788_y0);
  and_gate and_gate_h_u_cla32_and8789_y0(h_u_cla32_and8788_y0, h_u_cla32_and8787_y0, h_u_cla32_and8789_y0);
  and_gate and_gate_h_u_cla32_and8790_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8790_y0);
  and_gate and_gate_h_u_cla32_and8791_y0(h_u_cla32_and8790_y0, h_u_cla32_and8789_y0, h_u_cla32_and8791_y0);
  and_gate and_gate_h_u_cla32_and8792_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8792_y0);
  and_gate and_gate_h_u_cla32_and8793_y0(h_u_cla32_and8792_y0, h_u_cla32_and8791_y0, h_u_cla32_and8793_y0);
  and_gate and_gate_h_u_cla32_and8794_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8794_y0);
  and_gate and_gate_h_u_cla32_and8795_y0(h_u_cla32_and8794_y0, h_u_cla32_and8793_y0, h_u_cla32_and8795_y0);
  and_gate and_gate_h_u_cla32_and8796_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8796_y0);
  and_gate and_gate_h_u_cla32_and8797_y0(h_u_cla32_and8796_y0, h_u_cla32_and8795_y0, h_u_cla32_and8797_y0);
  and_gate and_gate_h_u_cla32_and8798_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8798_y0);
  and_gate and_gate_h_u_cla32_and8799_y0(h_u_cla32_and8798_y0, h_u_cla32_and8797_y0, h_u_cla32_and8799_y0);
  and_gate and_gate_h_u_cla32_and8800_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8800_y0);
  and_gate and_gate_h_u_cla32_and8801_y0(h_u_cla32_and8800_y0, h_u_cla32_and8799_y0, h_u_cla32_and8801_y0);
  and_gate and_gate_h_u_cla32_and8802_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8802_y0);
  and_gate and_gate_h_u_cla32_and8803_y0(h_u_cla32_and8802_y0, h_u_cla32_and8801_y0, h_u_cla32_and8803_y0);
  and_gate and_gate_h_u_cla32_and8804_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8804_y0);
  and_gate and_gate_h_u_cla32_and8805_y0(h_u_cla32_and8804_y0, h_u_cla32_and8803_y0, h_u_cla32_and8805_y0);
  and_gate and_gate_h_u_cla32_and8806_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8806_y0);
  and_gate and_gate_h_u_cla32_and8807_y0(h_u_cla32_and8806_y0, h_u_cla32_and8805_y0, h_u_cla32_and8807_y0);
  and_gate and_gate_h_u_cla32_and8808_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8808_y0);
  and_gate and_gate_h_u_cla32_and8809_y0(h_u_cla32_and8808_y0, h_u_cla32_and8807_y0, h_u_cla32_and8809_y0);
  and_gate and_gate_h_u_cla32_and8810_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8810_y0);
  and_gate and_gate_h_u_cla32_and8811_y0(h_u_cla32_and8810_y0, h_u_cla32_and8809_y0, h_u_cla32_and8811_y0);
  and_gate and_gate_h_u_cla32_and8812_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8812_y0);
  and_gate and_gate_h_u_cla32_and8813_y0(h_u_cla32_and8812_y0, h_u_cla32_and8811_y0, h_u_cla32_and8813_y0);
  and_gate and_gate_h_u_cla32_and8814_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8814_y0);
  and_gate and_gate_h_u_cla32_and8815_y0(h_u_cla32_and8814_y0, h_u_cla32_and8813_y0, h_u_cla32_and8815_y0);
  and_gate and_gate_h_u_cla32_and8816_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8816_y0);
  and_gate and_gate_h_u_cla32_and8817_y0(h_u_cla32_and8816_y0, h_u_cla32_and8815_y0, h_u_cla32_and8817_y0);
  and_gate and_gate_h_u_cla32_and8818_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8818_y0);
  and_gate and_gate_h_u_cla32_and8819_y0(h_u_cla32_and8818_y0, h_u_cla32_and8817_y0, h_u_cla32_and8819_y0);
  and_gate and_gate_h_u_cla32_and8820_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8820_y0);
  and_gate and_gate_h_u_cla32_and8821_y0(h_u_cla32_and8820_y0, h_u_cla32_and8819_y0, h_u_cla32_and8821_y0);
  and_gate and_gate_h_u_cla32_and8822_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8822_y0);
  and_gate and_gate_h_u_cla32_and8823_y0(h_u_cla32_and8822_y0, h_u_cla32_and8821_y0, h_u_cla32_and8823_y0);
  and_gate and_gate_h_u_cla32_and8824_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8824_y0);
  and_gate and_gate_h_u_cla32_and8825_y0(h_u_cla32_and8824_y0, h_u_cla32_and8823_y0, h_u_cla32_and8825_y0);
  and_gate and_gate_h_u_cla32_and8826_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8826_y0);
  and_gate and_gate_h_u_cla32_and8827_y0(h_u_cla32_and8826_y0, h_u_cla32_and8825_y0, h_u_cla32_and8827_y0);
  and_gate and_gate_h_u_cla32_and8828_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and8828_y0);
  and_gate and_gate_h_u_cla32_and8829_y0(h_u_cla32_and8828_y0, h_u_cla32_and8827_y0, h_u_cla32_and8829_y0);
  and_gate and_gate_h_u_cla32_and8830_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8830_y0);
  and_gate and_gate_h_u_cla32_and8831_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8831_y0);
  and_gate and_gate_h_u_cla32_and8832_y0(h_u_cla32_and8831_y0, h_u_cla32_and8830_y0, h_u_cla32_and8832_y0);
  and_gate and_gate_h_u_cla32_and8833_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8833_y0);
  and_gate and_gate_h_u_cla32_and8834_y0(h_u_cla32_and8833_y0, h_u_cla32_and8832_y0, h_u_cla32_and8834_y0);
  and_gate and_gate_h_u_cla32_and8835_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8835_y0);
  and_gate and_gate_h_u_cla32_and8836_y0(h_u_cla32_and8835_y0, h_u_cla32_and8834_y0, h_u_cla32_and8836_y0);
  and_gate and_gate_h_u_cla32_and8837_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8837_y0);
  and_gate and_gate_h_u_cla32_and8838_y0(h_u_cla32_and8837_y0, h_u_cla32_and8836_y0, h_u_cla32_and8838_y0);
  and_gate and_gate_h_u_cla32_and8839_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8839_y0);
  and_gate and_gate_h_u_cla32_and8840_y0(h_u_cla32_and8839_y0, h_u_cla32_and8838_y0, h_u_cla32_and8840_y0);
  and_gate and_gate_h_u_cla32_and8841_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8841_y0);
  and_gate and_gate_h_u_cla32_and8842_y0(h_u_cla32_and8841_y0, h_u_cla32_and8840_y0, h_u_cla32_and8842_y0);
  and_gate and_gate_h_u_cla32_and8843_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8843_y0);
  and_gate and_gate_h_u_cla32_and8844_y0(h_u_cla32_and8843_y0, h_u_cla32_and8842_y0, h_u_cla32_and8844_y0);
  and_gate and_gate_h_u_cla32_and8845_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8845_y0);
  and_gate and_gate_h_u_cla32_and8846_y0(h_u_cla32_and8845_y0, h_u_cla32_and8844_y0, h_u_cla32_and8846_y0);
  and_gate and_gate_h_u_cla32_and8847_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8847_y0);
  and_gate and_gate_h_u_cla32_and8848_y0(h_u_cla32_and8847_y0, h_u_cla32_and8846_y0, h_u_cla32_and8848_y0);
  and_gate and_gate_h_u_cla32_and8849_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8849_y0);
  and_gate and_gate_h_u_cla32_and8850_y0(h_u_cla32_and8849_y0, h_u_cla32_and8848_y0, h_u_cla32_and8850_y0);
  and_gate and_gate_h_u_cla32_and8851_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8851_y0);
  and_gate and_gate_h_u_cla32_and8852_y0(h_u_cla32_and8851_y0, h_u_cla32_and8850_y0, h_u_cla32_and8852_y0);
  and_gate and_gate_h_u_cla32_and8853_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8853_y0);
  and_gate and_gate_h_u_cla32_and8854_y0(h_u_cla32_and8853_y0, h_u_cla32_and8852_y0, h_u_cla32_and8854_y0);
  and_gate and_gate_h_u_cla32_and8855_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8855_y0);
  and_gate and_gate_h_u_cla32_and8856_y0(h_u_cla32_and8855_y0, h_u_cla32_and8854_y0, h_u_cla32_and8856_y0);
  and_gate and_gate_h_u_cla32_and8857_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8857_y0);
  and_gate and_gate_h_u_cla32_and8858_y0(h_u_cla32_and8857_y0, h_u_cla32_and8856_y0, h_u_cla32_and8858_y0);
  and_gate and_gate_h_u_cla32_and8859_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8859_y0);
  and_gate and_gate_h_u_cla32_and8860_y0(h_u_cla32_and8859_y0, h_u_cla32_and8858_y0, h_u_cla32_and8860_y0);
  and_gate and_gate_h_u_cla32_and8861_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8861_y0);
  and_gate and_gate_h_u_cla32_and8862_y0(h_u_cla32_and8861_y0, h_u_cla32_and8860_y0, h_u_cla32_and8862_y0);
  and_gate and_gate_h_u_cla32_and8863_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8863_y0);
  and_gate and_gate_h_u_cla32_and8864_y0(h_u_cla32_and8863_y0, h_u_cla32_and8862_y0, h_u_cla32_and8864_y0);
  and_gate and_gate_h_u_cla32_and8865_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8865_y0);
  and_gate and_gate_h_u_cla32_and8866_y0(h_u_cla32_and8865_y0, h_u_cla32_and8864_y0, h_u_cla32_and8866_y0);
  and_gate and_gate_h_u_cla32_and8867_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8867_y0);
  and_gate and_gate_h_u_cla32_and8868_y0(h_u_cla32_and8867_y0, h_u_cla32_and8866_y0, h_u_cla32_and8868_y0);
  and_gate and_gate_h_u_cla32_and8869_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8869_y0);
  and_gate and_gate_h_u_cla32_and8870_y0(h_u_cla32_and8869_y0, h_u_cla32_and8868_y0, h_u_cla32_and8870_y0);
  and_gate and_gate_h_u_cla32_and8871_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8871_y0);
  and_gate and_gate_h_u_cla32_and8872_y0(h_u_cla32_and8871_y0, h_u_cla32_and8870_y0, h_u_cla32_and8872_y0);
  and_gate and_gate_h_u_cla32_and8873_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8873_y0);
  and_gate and_gate_h_u_cla32_and8874_y0(h_u_cla32_and8873_y0, h_u_cla32_and8872_y0, h_u_cla32_and8874_y0);
  and_gate and_gate_h_u_cla32_and8875_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8875_y0);
  and_gate and_gate_h_u_cla32_and8876_y0(h_u_cla32_and8875_y0, h_u_cla32_and8874_y0, h_u_cla32_and8876_y0);
  and_gate and_gate_h_u_cla32_and8877_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and8877_y0);
  and_gate and_gate_h_u_cla32_and8878_y0(h_u_cla32_and8877_y0, h_u_cla32_and8876_y0, h_u_cla32_and8878_y0);
  and_gate and_gate_h_u_cla32_and8879_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8879_y0);
  and_gate and_gate_h_u_cla32_and8880_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8880_y0);
  and_gate and_gate_h_u_cla32_and8881_y0(h_u_cla32_and8880_y0, h_u_cla32_and8879_y0, h_u_cla32_and8881_y0);
  and_gate and_gate_h_u_cla32_and8882_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8882_y0);
  and_gate and_gate_h_u_cla32_and8883_y0(h_u_cla32_and8882_y0, h_u_cla32_and8881_y0, h_u_cla32_and8883_y0);
  and_gate and_gate_h_u_cla32_and8884_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8884_y0);
  and_gate and_gate_h_u_cla32_and8885_y0(h_u_cla32_and8884_y0, h_u_cla32_and8883_y0, h_u_cla32_and8885_y0);
  and_gate and_gate_h_u_cla32_and8886_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8886_y0);
  and_gate and_gate_h_u_cla32_and8887_y0(h_u_cla32_and8886_y0, h_u_cla32_and8885_y0, h_u_cla32_and8887_y0);
  and_gate and_gate_h_u_cla32_and8888_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8888_y0);
  and_gate and_gate_h_u_cla32_and8889_y0(h_u_cla32_and8888_y0, h_u_cla32_and8887_y0, h_u_cla32_and8889_y0);
  and_gate and_gate_h_u_cla32_and8890_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8890_y0);
  and_gate and_gate_h_u_cla32_and8891_y0(h_u_cla32_and8890_y0, h_u_cla32_and8889_y0, h_u_cla32_and8891_y0);
  and_gate and_gate_h_u_cla32_and8892_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8892_y0);
  and_gate and_gate_h_u_cla32_and8893_y0(h_u_cla32_and8892_y0, h_u_cla32_and8891_y0, h_u_cla32_and8893_y0);
  and_gate and_gate_h_u_cla32_and8894_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8894_y0);
  and_gate and_gate_h_u_cla32_and8895_y0(h_u_cla32_and8894_y0, h_u_cla32_and8893_y0, h_u_cla32_and8895_y0);
  and_gate and_gate_h_u_cla32_and8896_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8896_y0);
  and_gate and_gate_h_u_cla32_and8897_y0(h_u_cla32_and8896_y0, h_u_cla32_and8895_y0, h_u_cla32_and8897_y0);
  and_gate and_gate_h_u_cla32_and8898_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8898_y0);
  and_gate and_gate_h_u_cla32_and8899_y0(h_u_cla32_and8898_y0, h_u_cla32_and8897_y0, h_u_cla32_and8899_y0);
  and_gate and_gate_h_u_cla32_and8900_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8900_y0);
  and_gate and_gate_h_u_cla32_and8901_y0(h_u_cla32_and8900_y0, h_u_cla32_and8899_y0, h_u_cla32_and8901_y0);
  and_gate and_gate_h_u_cla32_and8902_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8902_y0);
  and_gate and_gate_h_u_cla32_and8903_y0(h_u_cla32_and8902_y0, h_u_cla32_and8901_y0, h_u_cla32_and8903_y0);
  and_gate and_gate_h_u_cla32_and8904_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8904_y0);
  and_gate and_gate_h_u_cla32_and8905_y0(h_u_cla32_and8904_y0, h_u_cla32_and8903_y0, h_u_cla32_and8905_y0);
  and_gate and_gate_h_u_cla32_and8906_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8906_y0);
  and_gate and_gate_h_u_cla32_and8907_y0(h_u_cla32_and8906_y0, h_u_cla32_and8905_y0, h_u_cla32_and8907_y0);
  and_gate and_gate_h_u_cla32_and8908_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8908_y0);
  and_gate and_gate_h_u_cla32_and8909_y0(h_u_cla32_and8908_y0, h_u_cla32_and8907_y0, h_u_cla32_and8909_y0);
  and_gate and_gate_h_u_cla32_and8910_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8910_y0);
  and_gate and_gate_h_u_cla32_and8911_y0(h_u_cla32_and8910_y0, h_u_cla32_and8909_y0, h_u_cla32_and8911_y0);
  and_gate and_gate_h_u_cla32_and8912_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8912_y0);
  and_gate and_gate_h_u_cla32_and8913_y0(h_u_cla32_and8912_y0, h_u_cla32_and8911_y0, h_u_cla32_and8913_y0);
  and_gate and_gate_h_u_cla32_and8914_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8914_y0);
  and_gate and_gate_h_u_cla32_and8915_y0(h_u_cla32_and8914_y0, h_u_cla32_and8913_y0, h_u_cla32_and8915_y0);
  and_gate and_gate_h_u_cla32_and8916_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8916_y0);
  and_gate and_gate_h_u_cla32_and8917_y0(h_u_cla32_and8916_y0, h_u_cla32_and8915_y0, h_u_cla32_and8917_y0);
  and_gate and_gate_h_u_cla32_and8918_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8918_y0);
  and_gate and_gate_h_u_cla32_and8919_y0(h_u_cla32_and8918_y0, h_u_cla32_and8917_y0, h_u_cla32_and8919_y0);
  and_gate and_gate_h_u_cla32_and8920_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8920_y0);
  and_gate and_gate_h_u_cla32_and8921_y0(h_u_cla32_and8920_y0, h_u_cla32_and8919_y0, h_u_cla32_and8921_y0);
  and_gate and_gate_h_u_cla32_and8922_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8922_y0);
  and_gate and_gate_h_u_cla32_and8923_y0(h_u_cla32_and8922_y0, h_u_cla32_and8921_y0, h_u_cla32_and8923_y0);
  and_gate and_gate_h_u_cla32_and8924_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and8924_y0);
  and_gate and_gate_h_u_cla32_and8925_y0(h_u_cla32_and8924_y0, h_u_cla32_and8923_y0, h_u_cla32_and8925_y0);
  and_gate and_gate_h_u_cla32_and8926_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8926_y0);
  and_gate and_gate_h_u_cla32_and8927_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8927_y0);
  and_gate and_gate_h_u_cla32_and8928_y0(h_u_cla32_and8927_y0, h_u_cla32_and8926_y0, h_u_cla32_and8928_y0);
  and_gate and_gate_h_u_cla32_and8929_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8929_y0);
  and_gate and_gate_h_u_cla32_and8930_y0(h_u_cla32_and8929_y0, h_u_cla32_and8928_y0, h_u_cla32_and8930_y0);
  and_gate and_gate_h_u_cla32_and8931_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8931_y0);
  and_gate and_gate_h_u_cla32_and8932_y0(h_u_cla32_and8931_y0, h_u_cla32_and8930_y0, h_u_cla32_and8932_y0);
  and_gate and_gate_h_u_cla32_and8933_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8933_y0);
  and_gate and_gate_h_u_cla32_and8934_y0(h_u_cla32_and8933_y0, h_u_cla32_and8932_y0, h_u_cla32_and8934_y0);
  and_gate and_gate_h_u_cla32_and8935_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8935_y0);
  and_gate and_gate_h_u_cla32_and8936_y0(h_u_cla32_and8935_y0, h_u_cla32_and8934_y0, h_u_cla32_and8936_y0);
  and_gate and_gate_h_u_cla32_and8937_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8937_y0);
  and_gate and_gate_h_u_cla32_and8938_y0(h_u_cla32_and8937_y0, h_u_cla32_and8936_y0, h_u_cla32_and8938_y0);
  and_gate and_gate_h_u_cla32_and8939_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8939_y0);
  and_gate and_gate_h_u_cla32_and8940_y0(h_u_cla32_and8939_y0, h_u_cla32_and8938_y0, h_u_cla32_and8940_y0);
  and_gate and_gate_h_u_cla32_and8941_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8941_y0);
  and_gate and_gate_h_u_cla32_and8942_y0(h_u_cla32_and8941_y0, h_u_cla32_and8940_y0, h_u_cla32_and8942_y0);
  and_gate and_gate_h_u_cla32_and8943_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8943_y0);
  and_gate and_gate_h_u_cla32_and8944_y0(h_u_cla32_and8943_y0, h_u_cla32_and8942_y0, h_u_cla32_and8944_y0);
  and_gate and_gate_h_u_cla32_and8945_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8945_y0);
  and_gate and_gate_h_u_cla32_and8946_y0(h_u_cla32_and8945_y0, h_u_cla32_and8944_y0, h_u_cla32_and8946_y0);
  and_gate and_gate_h_u_cla32_and8947_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8947_y0);
  and_gate and_gate_h_u_cla32_and8948_y0(h_u_cla32_and8947_y0, h_u_cla32_and8946_y0, h_u_cla32_and8948_y0);
  and_gate and_gate_h_u_cla32_and8949_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8949_y0);
  and_gate and_gate_h_u_cla32_and8950_y0(h_u_cla32_and8949_y0, h_u_cla32_and8948_y0, h_u_cla32_and8950_y0);
  and_gate and_gate_h_u_cla32_and8951_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8951_y0);
  and_gate and_gate_h_u_cla32_and8952_y0(h_u_cla32_and8951_y0, h_u_cla32_and8950_y0, h_u_cla32_and8952_y0);
  and_gate and_gate_h_u_cla32_and8953_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8953_y0);
  and_gate and_gate_h_u_cla32_and8954_y0(h_u_cla32_and8953_y0, h_u_cla32_and8952_y0, h_u_cla32_and8954_y0);
  and_gate and_gate_h_u_cla32_and8955_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8955_y0);
  and_gate and_gate_h_u_cla32_and8956_y0(h_u_cla32_and8955_y0, h_u_cla32_and8954_y0, h_u_cla32_and8956_y0);
  and_gate and_gate_h_u_cla32_and8957_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8957_y0);
  and_gate and_gate_h_u_cla32_and8958_y0(h_u_cla32_and8957_y0, h_u_cla32_and8956_y0, h_u_cla32_and8958_y0);
  and_gate and_gate_h_u_cla32_and8959_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8959_y0);
  and_gate and_gate_h_u_cla32_and8960_y0(h_u_cla32_and8959_y0, h_u_cla32_and8958_y0, h_u_cla32_and8960_y0);
  and_gate and_gate_h_u_cla32_and8961_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8961_y0);
  and_gate and_gate_h_u_cla32_and8962_y0(h_u_cla32_and8961_y0, h_u_cla32_and8960_y0, h_u_cla32_and8962_y0);
  and_gate and_gate_h_u_cla32_and8963_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8963_y0);
  and_gate and_gate_h_u_cla32_and8964_y0(h_u_cla32_and8963_y0, h_u_cla32_and8962_y0, h_u_cla32_and8964_y0);
  and_gate and_gate_h_u_cla32_and8965_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8965_y0);
  and_gate and_gate_h_u_cla32_and8966_y0(h_u_cla32_and8965_y0, h_u_cla32_and8964_y0, h_u_cla32_and8966_y0);
  and_gate and_gate_h_u_cla32_and8967_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8967_y0);
  and_gate and_gate_h_u_cla32_and8968_y0(h_u_cla32_and8967_y0, h_u_cla32_and8966_y0, h_u_cla32_and8968_y0);
  and_gate and_gate_h_u_cla32_and8969_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and8969_y0);
  and_gate and_gate_h_u_cla32_and8970_y0(h_u_cla32_and8969_y0, h_u_cla32_and8968_y0, h_u_cla32_and8970_y0);
  and_gate and_gate_h_u_cla32_and8971_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8971_y0);
  and_gate and_gate_h_u_cla32_and8972_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8972_y0);
  and_gate and_gate_h_u_cla32_and8973_y0(h_u_cla32_and8972_y0, h_u_cla32_and8971_y0, h_u_cla32_and8973_y0);
  and_gate and_gate_h_u_cla32_and8974_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8974_y0);
  and_gate and_gate_h_u_cla32_and8975_y0(h_u_cla32_and8974_y0, h_u_cla32_and8973_y0, h_u_cla32_and8975_y0);
  and_gate and_gate_h_u_cla32_and8976_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8976_y0);
  and_gate and_gate_h_u_cla32_and8977_y0(h_u_cla32_and8976_y0, h_u_cla32_and8975_y0, h_u_cla32_and8977_y0);
  and_gate and_gate_h_u_cla32_and8978_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8978_y0);
  and_gate and_gate_h_u_cla32_and8979_y0(h_u_cla32_and8978_y0, h_u_cla32_and8977_y0, h_u_cla32_and8979_y0);
  and_gate and_gate_h_u_cla32_and8980_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8980_y0);
  and_gate and_gate_h_u_cla32_and8981_y0(h_u_cla32_and8980_y0, h_u_cla32_and8979_y0, h_u_cla32_and8981_y0);
  and_gate and_gate_h_u_cla32_and8982_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8982_y0);
  and_gate and_gate_h_u_cla32_and8983_y0(h_u_cla32_and8982_y0, h_u_cla32_and8981_y0, h_u_cla32_and8983_y0);
  and_gate and_gate_h_u_cla32_and8984_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8984_y0);
  and_gate and_gate_h_u_cla32_and8985_y0(h_u_cla32_and8984_y0, h_u_cla32_and8983_y0, h_u_cla32_and8985_y0);
  and_gate and_gate_h_u_cla32_and8986_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8986_y0);
  and_gate and_gate_h_u_cla32_and8987_y0(h_u_cla32_and8986_y0, h_u_cla32_and8985_y0, h_u_cla32_and8987_y0);
  and_gate and_gate_h_u_cla32_and8988_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8988_y0);
  and_gate and_gate_h_u_cla32_and8989_y0(h_u_cla32_and8988_y0, h_u_cla32_and8987_y0, h_u_cla32_and8989_y0);
  and_gate and_gate_h_u_cla32_and8990_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8990_y0);
  and_gate and_gate_h_u_cla32_and8991_y0(h_u_cla32_and8990_y0, h_u_cla32_and8989_y0, h_u_cla32_and8991_y0);
  and_gate and_gate_h_u_cla32_and8992_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8992_y0);
  and_gate and_gate_h_u_cla32_and8993_y0(h_u_cla32_and8992_y0, h_u_cla32_and8991_y0, h_u_cla32_and8993_y0);
  and_gate and_gate_h_u_cla32_and8994_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8994_y0);
  and_gate and_gate_h_u_cla32_and8995_y0(h_u_cla32_and8994_y0, h_u_cla32_and8993_y0, h_u_cla32_and8995_y0);
  and_gate and_gate_h_u_cla32_and8996_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8996_y0);
  and_gate and_gate_h_u_cla32_and8997_y0(h_u_cla32_and8996_y0, h_u_cla32_and8995_y0, h_u_cla32_and8997_y0);
  and_gate and_gate_h_u_cla32_and8998_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and8998_y0);
  and_gate and_gate_h_u_cla32_and8999_y0(h_u_cla32_and8998_y0, h_u_cla32_and8997_y0, h_u_cla32_and8999_y0);
  and_gate and_gate_h_u_cla32_and9000_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9000_y0);
  and_gate and_gate_h_u_cla32_and9001_y0(h_u_cla32_and9000_y0, h_u_cla32_and8999_y0, h_u_cla32_and9001_y0);
  and_gate and_gate_h_u_cla32_and9002_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9002_y0);
  and_gate and_gate_h_u_cla32_and9003_y0(h_u_cla32_and9002_y0, h_u_cla32_and9001_y0, h_u_cla32_and9003_y0);
  and_gate and_gate_h_u_cla32_and9004_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9004_y0);
  and_gate and_gate_h_u_cla32_and9005_y0(h_u_cla32_and9004_y0, h_u_cla32_and9003_y0, h_u_cla32_and9005_y0);
  and_gate and_gate_h_u_cla32_and9006_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9006_y0);
  and_gate and_gate_h_u_cla32_and9007_y0(h_u_cla32_and9006_y0, h_u_cla32_and9005_y0, h_u_cla32_and9007_y0);
  and_gate and_gate_h_u_cla32_and9008_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9008_y0);
  and_gate and_gate_h_u_cla32_and9009_y0(h_u_cla32_and9008_y0, h_u_cla32_and9007_y0, h_u_cla32_and9009_y0);
  and_gate and_gate_h_u_cla32_and9010_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9010_y0);
  and_gate and_gate_h_u_cla32_and9011_y0(h_u_cla32_and9010_y0, h_u_cla32_and9009_y0, h_u_cla32_and9011_y0);
  and_gate and_gate_h_u_cla32_and9012_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9012_y0);
  and_gate and_gate_h_u_cla32_and9013_y0(h_u_cla32_and9012_y0, h_u_cla32_and9011_y0, h_u_cla32_and9013_y0);
  and_gate and_gate_h_u_cla32_and9014_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9014_y0);
  and_gate and_gate_h_u_cla32_and9015_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9015_y0);
  and_gate and_gate_h_u_cla32_and9016_y0(h_u_cla32_and9015_y0, h_u_cla32_and9014_y0, h_u_cla32_and9016_y0);
  and_gate and_gate_h_u_cla32_and9017_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9017_y0);
  and_gate and_gate_h_u_cla32_and9018_y0(h_u_cla32_and9017_y0, h_u_cla32_and9016_y0, h_u_cla32_and9018_y0);
  and_gate and_gate_h_u_cla32_and9019_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9019_y0);
  and_gate and_gate_h_u_cla32_and9020_y0(h_u_cla32_and9019_y0, h_u_cla32_and9018_y0, h_u_cla32_and9020_y0);
  and_gate and_gate_h_u_cla32_and9021_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9021_y0);
  and_gate and_gate_h_u_cla32_and9022_y0(h_u_cla32_and9021_y0, h_u_cla32_and9020_y0, h_u_cla32_and9022_y0);
  and_gate and_gate_h_u_cla32_and9023_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9023_y0);
  and_gate and_gate_h_u_cla32_and9024_y0(h_u_cla32_and9023_y0, h_u_cla32_and9022_y0, h_u_cla32_and9024_y0);
  and_gate and_gate_h_u_cla32_and9025_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9025_y0);
  and_gate and_gate_h_u_cla32_and9026_y0(h_u_cla32_and9025_y0, h_u_cla32_and9024_y0, h_u_cla32_and9026_y0);
  and_gate and_gate_h_u_cla32_and9027_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9027_y0);
  and_gate and_gate_h_u_cla32_and9028_y0(h_u_cla32_and9027_y0, h_u_cla32_and9026_y0, h_u_cla32_and9028_y0);
  and_gate and_gate_h_u_cla32_and9029_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9029_y0);
  and_gate and_gate_h_u_cla32_and9030_y0(h_u_cla32_and9029_y0, h_u_cla32_and9028_y0, h_u_cla32_and9030_y0);
  and_gate and_gate_h_u_cla32_and9031_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9031_y0);
  and_gate and_gate_h_u_cla32_and9032_y0(h_u_cla32_and9031_y0, h_u_cla32_and9030_y0, h_u_cla32_and9032_y0);
  and_gate and_gate_h_u_cla32_and9033_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9033_y0);
  and_gate and_gate_h_u_cla32_and9034_y0(h_u_cla32_and9033_y0, h_u_cla32_and9032_y0, h_u_cla32_and9034_y0);
  and_gate and_gate_h_u_cla32_and9035_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9035_y0);
  and_gate and_gate_h_u_cla32_and9036_y0(h_u_cla32_and9035_y0, h_u_cla32_and9034_y0, h_u_cla32_and9036_y0);
  and_gate and_gate_h_u_cla32_and9037_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9037_y0);
  and_gate and_gate_h_u_cla32_and9038_y0(h_u_cla32_and9037_y0, h_u_cla32_and9036_y0, h_u_cla32_and9038_y0);
  and_gate and_gate_h_u_cla32_and9039_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9039_y0);
  and_gate and_gate_h_u_cla32_and9040_y0(h_u_cla32_and9039_y0, h_u_cla32_and9038_y0, h_u_cla32_and9040_y0);
  and_gate and_gate_h_u_cla32_and9041_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9041_y0);
  and_gate and_gate_h_u_cla32_and9042_y0(h_u_cla32_and9041_y0, h_u_cla32_and9040_y0, h_u_cla32_and9042_y0);
  and_gate and_gate_h_u_cla32_and9043_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9043_y0);
  and_gate and_gate_h_u_cla32_and9044_y0(h_u_cla32_and9043_y0, h_u_cla32_and9042_y0, h_u_cla32_and9044_y0);
  and_gate and_gate_h_u_cla32_and9045_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9045_y0);
  and_gate and_gate_h_u_cla32_and9046_y0(h_u_cla32_and9045_y0, h_u_cla32_and9044_y0, h_u_cla32_and9046_y0);
  and_gate and_gate_h_u_cla32_and9047_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9047_y0);
  and_gate and_gate_h_u_cla32_and9048_y0(h_u_cla32_and9047_y0, h_u_cla32_and9046_y0, h_u_cla32_and9048_y0);
  and_gate and_gate_h_u_cla32_and9049_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9049_y0);
  and_gate and_gate_h_u_cla32_and9050_y0(h_u_cla32_and9049_y0, h_u_cla32_and9048_y0, h_u_cla32_and9050_y0);
  and_gate and_gate_h_u_cla32_and9051_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9051_y0);
  and_gate and_gate_h_u_cla32_and9052_y0(h_u_cla32_and9051_y0, h_u_cla32_and9050_y0, h_u_cla32_and9052_y0);
  and_gate and_gate_h_u_cla32_and9053_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9053_y0);
  and_gate and_gate_h_u_cla32_and9054_y0(h_u_cla32_and9053_y0, h_u_cla32_and9052_y0, h_u_cla32_and9054_y0);
  and_gate and_gate_h_u_cla32_and9055_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9055_y0);
  and_gate and_gate_h_u_cla32_and9056_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9056_y0);
  and_gate and_gate_h_u_cla32_and9057_y0(h_u_cla32_and9056_y0, h_u_cla32_and9055_y0, h_u_cla32_and9057_y0);
  and_gate and_gate_h_u_cla32_and9058_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9058_y0);
  and_gate and_gate_h_u_cla32_and9059_y0(h_u_cla32_and9058_y0, h_u_cla32_and9057_y0, h_u_cla32_and9059_y0);
  and_gate and_gate_h_u_cla32_and9060_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9060_y0);
  and_gate and_gate_h_u_cla32_and9061_y0(h_u_cla32_and9060_y0, h_u_cla32_and9059_y0, h_u_cla32_and9061_y0);
  and_gate and_gate_h_u_cla32_and9062_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9062_y0);
  and_gate and_gate_h_u_cla32_and9063_y0(h_u_cla32_and9062_y0, h_u_cla32_and9061_y0, h_u_cla32_and9063_y0);
  and_gate and_gate_h_u_cla32_and9064_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9064_y0);
  and_gate and_gate_h_u_cla32_and9065_y0(h_u_cla32_and9064_y0, h_u_cla32_and9063_y0, h_u_cla32_and9065_y0);
  and_gate and_gate_h_u_cla32_and9066_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9066_y0);
  and_gate and_gate_h_u_cla32_and9067_y0(h_u_cla32_and9066_y0, h_u_cla32_and9065_y0, h_u_cla32_and9067_y0);
  and_gate and_gate_h_u_cla32_and9068_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9068_y0);
  and_gate and_gate_h_u_cla32_and9069_y0(h_u_cla32_and9068_y0, h_u_cla32_and9067_y0, h_u_cla32_and9069_y0);
  and_gate and_gate_h_u_cla32_and9070_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9070_y0);
  and_gate and_gate_h_u_cla32_and9071_y0(h_u_cla32_and9070_y0, h_u_cla32_and9069_y0, h_u_cla32_and9071_y0);
  and_gate and_gate_h_u_cla32_and9072_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9072_y0);
  and_gate and_gate_h_u_cla32_and9073_y0(h_u_cla32_and9072_y0, h_u_cla32_and9071_y0, h_u_cla32_and9073_y0);
  and_gate and_gate_h_u_cla32_and9074_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9074_y0);
  and_gate and_gate_h_u_cla32_and9075_y0(h_u_cla32_and9074_y0, h_u_cla32_and9073_y0, h_u_cla32_and9075_y0);
  and_gate and_gate_h_u_cla32_and9076_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9076_y0);
  and_gate and_gate_h_u_cla32_and9077_y0(h_u_cla32_and9076_y0, h_u_cla32_and9075_y0, h_u_cla32_and9077_y0);
  and_gate and_gate_h_u_cla32_and9078_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9078_y0);
  and_gate and_gate_h_u_cla32_and9079_y0(h_u_cla32_and9078_y0, h_u_cla32_and9077_y0, h_u_cla32_and9079_y0);
  and_gate and_gate_h_u_cla32_and9080_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9080_y0);
  and_gate and_gate_h_u_cla32_and9081_y0(h_u_cla32_and9080_y0, h_u_cla32_and9079_y0, h_u_cla32_and9081_y0);
  and_gate and_gate_h_u_cla32_and9082_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9082_y0);
  and_gate and_gate_h_u_cla32_and9083_y0(h_u_cla32_and9082_y0, h_u_cla32_and9081_y0, h_u_cla32_and9083_y0);
  and_gate and_gate_h_u_cla32_and9084_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9084_y0);
  and_gate and_gate_h_u_cla32_and9085_y0(h_u_cla32_and9084_y0, h_u_cla32_and9083_y0, h_u_cla32_and9085_y0);
  and_gate and_gate_h_u_cla32_and9086_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9086_y0);
  and_gate and_gate_h_u_cla32_and9087_y0(h_u_cla32_and9086_y0, h_u_cla32_and9085_y0, h_u_cla32_and9087_y0);
  and_gate and_gate_h_u_cla32_and9088_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9088_y0);
  and_gate and_gate_h_u_cla32_and9089_y0(h_u_cla32_and9088_y0, h_u_cla32_and9087_y0, h_u_cla32_and9089_y0);
  and_gate and_gate_h_u_cla32_and9090_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9090_y0);
  and_gate and_gate_h_u_cla32_and9091_y0(h_u_cla32_and9090_y0, h_u_cla32_and9089_y0, h_u_cla32_and9091_y0);
  and_gate and_gate_h_u_cla32_and9092_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9092_y0);
  and_gate and_gate_h_u_cla32_and9093_y0(h_u_cla32_and9092_y0, h_u_cla32_and9091_y0, h_u_cla32_and9093_y0);
  and_gate and_gate_h_u_cla32_and9094_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9094_y0);
  and_gate and_gate_h_u_cla32_and9095_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9095_y0);
  and_gate and_gate_h_u_cla32_and9096_y0(h_u_cla32_and9095_y0, h_u_cla32_and9094_y0, h_u_cla32_and9096_y0);
  and_gate and_gate_h_u_cla32_and9097_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9097_y0);
  and_gate and_gate_h_u_cla32_and9098_y0(h_u_cla32_and9097_y0, h_u_cla32_and9096_y0, h_u_cla32_and9098_y0);
  and_gate and_gate_h_u_cla32_and9099_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9099_y0);
  and_gate and_gate_h_u_cla32_and9100_y0(h_u_cla32_and9099_y0, h_u_cla32_and9098_y0, h_u_cla32_and9100_y0);
  and_gate and_gate_h_u_cla32_and9101_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9101_y0);
  and_gate and_gate_h_u_cla32_and9102_y0(h_u_cla32_and9101_y0, h_u_cla32_and9100_y0, h_u_cla32_and9102_y0);
  and_gate and_gate_h_u_cla32_and9103_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9103_y0);
  and_gate and_gate_h_u_cla32_and9104_y0(h_u_cla32_and9103_y0, h_u_cla32_and9102_y0, h_u_cla32_and9104_y0);
  and_gate and_gate_h_u_cla32_and9105_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9105_y0);
  and_gate and_gate_h_u_cla32_and9106_y0(h_u_cla32_and9105_y0, h_u_cla32_and9104_y0, h_u_cla32_and9106_y0);
  and_gate and_gate_h_u_cla32_and9107_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9107_y0);
  and_gate and_gate_h_u_cla32_and9108_y0(h_u_cla32_and9107_y0, h_u_cla32_and9106_y0, h_u_cla32_and9108_y0);
  and_gate and_gate_h_u_cla32_and9109_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9109_y0);
  and_gate and_gate_h_u_cla32_and9110_y0(h_u_cla32_and9109_y0, h_u_cla32_and9108_y0, h_u_cla32_and9110_y0);
  and_gate and_gate_h_u_cla32_and9111_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9111_y0);
  and_gate and_gate_h_u_cla32_and9112_y0(h_u_cla32_and9111_y0, h_u_cla32_and9110_y0, h_u_cla32_and9112_y0);
  and_gate and_gate_h_u_cla32_and9113_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9113_y0);
  and_gate and_gate_h_u_cla32_and9114_y0(h_u_cla32_and9113_y0, h_u_cla32_and9112_y0, h_u_cla32_and9114_y0);
  and_gate and_gate_h_u_cla32_and9115_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9115_y0);
  and_gate and_gate_h_u_cla32_and9116_y0(h_u_cla32_and9115_y0, h_u_cla32_and9114_y0, h_u_cla32_and9116_y0);
  and_gate and_gate_h_u_cla32_and9117_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9117_y0);
  and_gate and_gate_h_u_cla32_and9118_y0(h_u_cla32_and9117_y0, h_u_cla32_and9116_y0, h_u_cla32_and9118_y0);
  and_gate and_gate_h_u_cla32_and9119_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9119_y0);
  and_gate and_gate_h_u_cla32_and9120_y0(h_u_cla32_and9119_y0, h_u_cla32_and9118_y0, h_u_cla32_and9120_y0);
  and_gate and_gate_h_u_cla32_and9121_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9121_y0);
  and_gate and_gate_h_u_cla32_and9122_y0(h_u_cla32_and9121_y0, h_u_cla32_and9120_y0, h_u_cla32_and9122_y0);
  and_gate and_gate_h_u_cla32_and9123_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9123_y0);
  and_gate and_gate_h_u_cla32_and9124_y0(h_u_cla32_and9123_y0, h_u_cla32_and9122_y0, h_u_cla32_and9124_y0);
  and_gate and_gate_h_u_cla32_and9125_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9125_y0);
  and_gate and_gate_h_u_cla32_and9126_y0(h_u_cla32_and9125_y0, h_u_cla32_and9124_y0, h_u_cla32_and9126_y0);
  and_gate and_gate_h_u_cla32_and9127_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9127_y0);
  and_gate and_gate_h_u_cla32_and9128_y0(h_u_cla32_and9127_y0, h_u_cla32_and9126_y0, h_u_cla32_and9128_y0);
  and_gate and_gate_h_u_cla32_and9129_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and9129_y0);
  and_gate and_gate_h_u_cla32_and9130_y0(h_u_cla32_and9129_y0, h_u_cla32_and9128_y0, h_u_cla32_and9130_y0);
  and_gate and_gate_h_u_cla32_and9131_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9131_y0);
  and_gate and_gate_h_u_cla32_and9132_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9132_y0);
  and_gate and_gate_h_u_cla32_and9133_y0(h_u_cla32_and9132_y0, h_u_cla32_and9131_y0, h_u_cla32_and9133_y0);
  and_gate and_gate_h_u_cla32_and9134_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9134_y0);
  and_gate and_gate_h_u_cla32_and9135_y0(h_u_cla32_and9134_y0, h_u_cla32_and9133_y0, h_u_cla32_and9135_y0);
  and_gate and_gate_h_u_cla32_and9136_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9136_y0);
  and_gate and_gate_h_u_cla32_and9137_y0(h_u_cla32_and9136_y0, h_u_cla32_and9135_y0, h_u_cla32_and9137_y0);
  and_gate and_gate_h_u_cla32_and9138_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9138_y0);
  and_gate and_gate_h_u_cla32_and9139_y0(h_u_cla32_and9138_y0, h_u_cla32_and9137_y0, h_u_cla32_and9139_y0);
  and_gate and_gate_h_u_cla32_and9140_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9140_y0);
  and_gate and_gate_h_u_cla32_and9141_y0(h_u_cla32_and9140_y0, h_u_cla32_and9139_y0, h_u_cla32_and9141_y0);
  and_gate and_gate_h_u_cla32_and9142_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9142_y0);
  and_gate and_gate_h_u_cla32_and9143_y0(h_u_cla32_and9142_y0, h_u_cla32_and9141_y0, h_u_cla32_and9143_y0);
  and_gate and_gate_h_u_cla32_and9144_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9144_y0);
  and_gate and_gate_h_u_cla32_and9145_y0(h_u_cla32_and9144_y0, h_u_cla32_and9143_y0, h_u_cla32_and9145_y0);
  and_gate and_gate_h_u_cla32_and9146_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9146_y0);
  and_gate and_gate_h_u_cla32_and9147_y0(h_u_cla32_and9146_y0, h_u_cla32_and9145_y0, h_u_cla32_and9147_y0);
  and_gate and_gate_h_u_cla32_and9148_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9148_y0);
  and_gate and_gate_h_u_cla32_and9149_y0(h_u_cla32_and9148_y0, h_u_cla32_and9147_y0, h_u_cla32_and9149_y0);
  and_gate and_gate_h_u_cla32_and9150_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9150_y0);
  and_gate and_gate_h_u_cla32_and9151_y0(h_u_cla32_and9150_y0, h_u_cla32_and9149_y0, h_u_cla32_and9151_y0);
  and_gate and_gate_h_u_cla32_and9152_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9152_y0);
  and_gate and_gate_h_u_cla32_and9153_y0(h_u_cla32_and9152_y0, h_u_cla32_and9151_y0, h_u_cla32_and9153_y0);
  and_gate and_gate_h_u_cla32_and9154_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9154_y0);
  and_gate and_gate_h_u_cla32_and9155_y0(h_u_cla32_and9154_y0, h_u_cla32_and9153_y0, h_u_cla32_and9155_y0);
  and_gate and_gate_h_u_cla32_and9156_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9156_y0);
  and_gate and_gate_h_u_cla32_and9157_y0(h_u_cla32_and9156_y0, h_u_cla32_and9155_y0, h_u_cla32_and9157_y0);
  and_gate and_gate_h_u_cla32_and9158_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9158_y0);
  and_gate and_gate_h_u_cla32_and9159_y0(h_u_cla32_and9158_y0, h_u_cla32_and9157_y0, h_u_cla32_and9159_y0);
  and_gate and_gate_h_u_cla32_and9160_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9160_y0);
  and_gate and_gate_h_u_cla32_and9161_y0(h_u_cla32_and9160_y0, h_u_cla32_and9159_y0, h_u_cla32_and9161_y0);
  and_gate and_gate_h_u_cla32_and9162_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9162_y0);
  and_gate and_gate_h_u_cla32_and9163_y0(h_u_cla32_and9162_y0, h_u_cla32_and9161_y0, h_u_cla32_and9163_y0);
  and_gate and_gate_h_u_cla32_and9164_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and9164_y0);
  and_gate and_gate_h_u_cla32_and9165_y0(h_u_cla32_and9164_y0, h_u_cla32_and9163_y0, h_u_cla32_and9165_y0);
  and_gate and_gate_h_u_cla32_and9166_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9166_y0);
  and_gate and_gate_h_u_cla32_and9167_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9167_y0);
  and_gate and_gate_h_u_cla32_and9168_y0(h_u_cla32_and9167_y0, h_u_cla32_and9166_y0, h_u_cla32_and9168_y0);
  and_gate and_gate_h_u_cla32_and9169_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9169_y0);
  and_gate and_gate_h_u_cla32_and9170_y0(h_u_cla32_and9169_y0, h_u_cla32_and9168_y0, h_u_cla32_and9170_y0);
  and_gate and_gate_h_u_cla32_and9171_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9171_y0);
  and_gate and_gate_h_u_cla32_and9172_y0(h_u_cla32_and9171_y0, h_u_cla32_and9170_y0, h_u_cla32_and9172_y0);
  and_gate and_gate_h_u_cla32_and9173_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9173_y0);
  and_gate and_gate_h_u_cla32_and9174_y0(h_u_cla32_and9173_y0, h_u_cla32_and9172_y0, h_u_cla32_and9174_y0);
  and_gate and_gate_h_u_cla32_and9175_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9175_y0);
  and_gate and_gate_h_u_cla32_and9176_y0(h_u_cla32_and9175_y0, h_u_cla32_and9174_y0, h_u_cla32_and9176_y0);
  and_gate and_gate_h_u_cla32_and9177_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9177_y0);
  and_gate and_gate_h_u_cla32_and9178_y0(h_u_cla32_and9177_y0, h_u_cla32_and9176_y0, h_u_cla32_and9178_y0);
  and_gate and_gate_h_u_cla32_and9179_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9179_y0);
  and_gate and_gate_h_u_cla32_and9180_y0(h_u_cla32_and9179_y0, h_u_cla32_and9178_y0, h_u_cla32_and9180_y0);
  and_gate and_gate_h_u_cla32_and9181_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9181_y0);
  and_gate and_gate_h_u_cla32_and9182_y0(h_u_cla32_and9181_y0, h_u_cla32_and9180_y0, h_u_cla32_and9182_y0);
  and_gate and_gate_h_u_cla32_and9183_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9183_y0);
  and_gate and_gate_h_u_cla32_and9184_y0(h_u_cla32_and9183_y0, h_u_cla32_and9182_y0, h_u_cla32_and9184_y0);
  and_gate and_gate_h_u_cla32_and9185_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9185_y0);
  and_gate and_gate_h_u_cla32_and9186_y0(h_u_cla32_and9185_y0, h_u_cla32_and9184_y0, h_u_cla32_and9186_y0);
  and_gate and_gate_h_u_cla32_and9187_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9187_y0);
  and_gate and_gate_h_u_cla32_and9188_y0(h_u_cla32_and9187_y0, h_u_cla32_and9186_y0, h_u_cla32_and9188_y0);
  and_gate and_gate_h_u_cla32_and9189_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9189_y0);
  and_gate and_gate_h_u_cla32_and9190_y0(h_u_cla32_and9189_y0, h_u_cla32_and9188_y0, h_u_cla32_and9190_y0);
  and_gate and_gate_h_u_cla32_and9191_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9191_y0);
  and_gate and_gate_h_u_cla32_and9192_y0(h_u_cla32_and9191_y0, h_u_cla32_and9190_y0, h_u_cla32_and9192_y0);
  and_gate and_gate_h_u_cla32_and9193_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9193_y0);
  and_gate and_gate_h_u_cla32_and9194_y0(h_u_cla32_and9193_y0, h_u_cla32_and9192_y0, h_u_cla32_and9194_y0);
  and_gate and_gate_h_u_cla32_and9195_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9195_y0);
  and_gate and_gate_h_u_cla32_and9196_y0(h_u_cla32_and9195_y0, h_u_cla32_and9194_y0, h_u_cla32_and9196_y0);
  and_gate and_gate_h_u_cla32_and9197_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and9197_y0);
  and_gate and_gate_h_u_cla32_and9198_y0(h_u_cla32_and9197_y0, h_u_cla32_and9196_y0, h_u_cla32_and9198_y0);
  and_gate and_gate_h_u_cla32_and9199_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9199_y0);
  and_gate and_gate_h_u_cla32_and9200_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9200_y0);
  and_gate and_gate_h_u_cla32_and9201_y0(h_u_cla32_and9200_y0, h_u_cla32_and9199_y0, h_u_cla32_and9201_y0);
  and_gate and_gate_h_u_cla32_and9202_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9202_y0);
  and_gate and_gate_h_u_cla32_and9203_y0(h_u_cla32_and9202_y0, h_u_cla32_and9201_y0, h_u_cla32_and9203_y0);
  and_gate and_gate_h_u_cla32_and9204_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9204_y0);
  and_gate and_gate_h_u_cla32_and9205_y0(h_u_cla32_and9204_y0, h_u_cla32_and9203_y0, h_u_cla32_and9205_y0);
  and_gate and_gate_h_u_cla32_and9206_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9206_y0);
  and_gate and_gate_h_u_cla32_and9207_y0(h_u_cla32_and9206_y0, h_u_cla32_and9205_y0, h_u_cla32_and9207_y0);
  and_gate and_gate_h_u_cla32_and9208_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9208_y0);
  and_gate and_gate_h_u_cla32_and9209_y0(h_u_cla32_and9208_y0, h_u_cla32_and9207_y0, h_u_cla32_and9209_y0);
  and_gate and_gate_h_u_cla32_and9210_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9210_y0);
  and_gate and_gate_h_u_cla32_and9211_y0(h_u_cla32_and9210_y0, h_u_cla32_and9209_y0, h_u_cla32_and9211_y0);
  and_gate and_gate_h_u_cla32_and9212_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9212_y0);
  and_gate and_gate_h_u_cla32_and9213_y0(h_u_cla32_and9212_y0, h_u_cla32_and9211_y0, h_u_cla32_and9213_y0);
  and_gate and_gate_h_u_cla32_and9214_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9214_y0);
  and_gate and_gate_h_u_cla32_and9215_y0(h_u_cla32_and9214_y0, h_u_cla32_and9213_y0, h_u_cla32_and9215_y0);
  and_gate and_gate_h_u_cla32_and9216_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9216_y0);
  and_gate and_gate_h_u_cla32_and9217_y0(h_u_cla32_and9216_y0, h_u_cla32_and9215_y0, h_u_cla32_and9217_y0);
  and_gate and_gate_h_u_cla32_and9218_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9218_y0);
  and_gate and_gate_h_u_cla32_and9219_y0(h_u_cla32_and9218_y0, h_u_cla32_and9217_y0, h_u_cla32_and9219_y0);
  and_gate and_gate_h_u_cla32_and9220_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9220_y0);
  and_gate and_gate_h_u_cla32_and9221_y0(h_u_cla32_and9220_y0, h_u_cla32_and9219_y0, h_u_cla32_and9221_y0);
  and_gate and_gate_h_u_cla32_and9222_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9222_y0);
  and_gate and_gate_h_u_cla32_and9223_y0(h_u_cla32_and9222_y0, h_u_cla32_and9221_y0, h_u_cla32_and9223_y0);
  and_gate and_gate_h_u_cla32_and9224_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9224_y0);
  and_gate and_gate_h_u_cla32_and9225_y0(h_u_cla32_and9224_y0, h_u_cla32_and9223_y0, h_u_cla32_and9225_y0);
  and_gate and_gate_h_u_cla32_and9226_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9226_y0);
  and_gate and_gate_h_u_cla32_and9227_y0(h_u_cla32_and9226_y0, h_u_cla32_and9225_y0, h_u_cla32_and9227_y0);
  and_gate and_gate_h_u_cla32_and9228_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and9228_y0);
  and_gate and_gate_h_u_cla32_and9229_y0(h_u_cla32_and9228_y0, h_u_cla32_and9227_y0, h_u_cla32_and9229_y0);
  and_gate and_gate_h_u_cla32_and9230_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9230_y0);
  and_gate and_gate_h_u_cla32_and9231_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9231_y0);
  and_gate and_gate_h_u_cla32_and9232_y0(h_u_cla32_and9231_y0, h_u_cla32_and9230_y0, h_u_cla32_and9232_y0);
  and_gate and_gate_h_u_cla32_and9233_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9233_y0);
  and_gate and_gate_h_u_cla32_and9234_y0(h_u_cla32_and9233_y0, h_u_cla32_and9232_y0, h_u_cla32_and9234_y0);
  and_gate and_gate_h_u_cla32_and9235_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9235_y0);
  and_gate and_gate_h_u_cla32_and9236_y0(h_u_cla32_and9235_y0, h_u_cla32_and9234_y0, h_u_cla32_and9236_y0);
  and_gate and_gate_h_u_cla32_and9237_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9237_y0);
  and_gate and_gate_h_u_cla32_and9238_y0(h_u_cla32_and9237_y0, h_u_cla32_and9236_y0, h_u_cla32_and9238_y0);
  and_gate and_gate_h_u_cla32_and9239_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9239_y0);
  and_gate and_gate_h_u_cla32_and9240_y0(h_u_cla32_and9239_y0, h_u_cla32_and9238_y0, h_u_cla32_and9240_y0);
  and_gate and_gate_h_u_cla32_and9241_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9241_y0);
  and_gate and_gate_h_u_cla32_and9242_y0(h_u_cla32_and9241_y0, h_u_cla32_and9240_y0, h_u_cla32_and9242_y0);
  and_gate and_gate_h_u_cla32_and9243_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9243_y0);
  and_gate and_gate_h_u_cla32_and9244_y0(h_u_cla32_and9243_y0, h_u_cla32_and9242_y0, h_u_cla32_and9244_y0);
  and_gate and_gate_h_u_cla32_and9245_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9245_y0);
  and_gate and_gate_h_u_cla32_and9246_y0(h_u_cla32_and9245_y0, h_u_cla32_and9244_y0, h_u_cla32_and9246_y0);
  and_gate and_gate_h_u_cla32_and9247_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9247_y0);
  and_gate and_gate_h_u_cla32_and9248_y0(h_u_cla32_and9247_y0, h_u_cla32_and9246_y0, h_u_cla32_and9248_y0);
  and_gate and_gate_h_u_cla32_and9249_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9249_y0);
  and_gate and_gate_h_u_cla32_and9250_y0(h_u_cla32_and9249_y0, h_u_cla32_and9248_y0, h_u_cla32_and9250_y0);
  and_gate and_gate_h_u_cla32_and9251_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9251_y0);
  and_gate and_gate_h_u_cla32_and9252_y0(h_u_cla32_and9251_y0, h_u_cla32_and9250_y0, h_u_cla32_and9252_y0);
  and_gate and_gate_h_u_cla32_and9253_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9253_y0);
  and_gate and_gate_h_u_cla32_and9254_y0(h_u_cla32_and9253_y0, h_u_cla32_and9252_y0, h_u_cla32_and9254_y0);
  and_gate and_gate_h_u_cla32_and9255_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9255_y0);
  and_gate and_gate_h_u_cla32_and9256_y0(h_u_cla32_and9255_y0, h_u_cla32_and9254_y0, h_u_cla32_and9256_y0);
  and_gate and_gate_h_u_cla32_and9257_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and9257_y0);
  and_gate and_gate_h_u_cla32_and9258_y0(h_u_cla32_and9257_y0, h_u_cla32_and9256_y0, h_u_cla32_and9258_y0);
  and_gate and_gate_h_u_cla32_and9259_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9259_y0);
  and_gate and_gate_h_u_cla32_and9260_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9260_y0);
  and_gate and_gate_h_u_cla32_and9261_y0(h_u_cla32_and9260_y0, h_u_cla32_and9259_y0, h_u_cla32_and9261_y0);
  and_gate and_gate_h_u_cla32_and9262_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9262_y0);
  and_gate and_gate_h_u_cla32_and9263_y0(h_u_cla32_and9262_y0, h_u_cla32_and9261_y0, h_u_cla32_and9263_y0);
  and_gate and_gate_h_u_cla32_and9264_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9264_y0);
  and_gate and_gate_h_u_cla32_and9265_y0(h_u_cla32_and9264_y0, h_u_cla32_and9263_y0, h_u_cla32_and9265_y0);
  and_gate and_gate_h_u_cla32_and9266_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9266_y0);
  and_gate and_gate_h_u_cla32_and9267_y0(h_u_cla32_and9266_y0, h_u_cla32_and9265_y0, h_u_cla32_and9267_y0);
  and_gate and_gate_h_u_cla32_and9268_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9268_y0);
  and_gate and_gate_h_u_cla32_and9269_y0(h_u_cla32_and9268_y0, h_u_cla32_and9267_y0, h_u_cla32_and9269_y0);
  and_gate and_gate_h_u_cla32_and9270_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9270_y0);
  and_gate and_gate_h_u_cla32_and9271_y0(h_u_cla32_and9270_y0, h_u_cla32_and9269_y0, h_u_cla32_and9271_y0);
  and_gate and_gate_h_u_cla32_and9272_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9272_y0);
  and_gate and_gate_h_u_cla32_and9273_y0(h_u_cla32_and9272_y0, h_u_cla32_and9271_y0, h_u_cla32_and9273_y0);
  and_gate and_gate_h_u_cla32_and9274_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9274_y0);
  and_gate and_gate_h_u_cla32_and9275_y0(h_u_cla32_and9274_y0, h_u_cla32_and9273_y0, h_u_cla32_and9275_y0);
  and_gate and_gate_h_u_cla32_and9276_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9276_y0);
  and_gate and_gate_h_u_cla32_and9277_y0(h_u_cla32_and9276_y0, h_u_cla32_and9275_y0, h_u_cla32_and9277_y0);
  and_gate and_gate_h_u_cla32_and9278_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9278_y0);
  and_gate and_gate_h_u_cla32_and9279_y0(h_u_cla32_and9278_y0, h_u_cla32_and9277_y0, h_u_cla32_and9279_y0);
  and_gate and_gate_h_u_cla32_and9280_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9280_y0);
  and_gate and_gate_h_u_cla32_and9281_y0(h_u_cla32_and9280_y0, h_u_cla32_and9279_y0, h_u_cla32_and9281_y0);
  and_gate and_gate_h_u_cla32_and9282_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9282_y0);
  and_gate and_gate_h_u_cla32_and9283_y0(h_u_cla32_and9282_y0, h_u_cla32_and9281_y0, h_u_cla32_and9283_y0);
  and_gate and_gate_h_u_cla32_and9284_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and9284_y0);
  and_gate and_gate_h_u_cla32_and9285_y0(h_u_cla32_and9284_y0, h_u_cla32_and9283_y0, h_u_cla32_and9285_y0);
  and_gate and_gate_h_u_cla32_and9286_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9286_y0);
  and_gate and_gate_h_u_cla32_and9287_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9287_y0);
  and_gate and_gate_h_u_cla32_and9288_y0(h_u_cla32_and9287_y0, h_u_cla32_and9286_y0, h_u_cla32_and9288_y0);
  and_gate and_gate_h_u_cla32_and9289_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9289_y0);
  and_gate and_gate_h_u_cla32_and9290_y0(h_u_cla32_and9289_y0, h_u_cla32_and9288_y0, h_u_cla32_and9290_y0);
  and_gate and_gate_h_u_cla32_and9291_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9291_y0);
  and_gate and_gate_h_u_cla32_and9292_y0(h_u_cla32_and9291_y0, h_u_cla32_and9290_y0, h_u_cla32_and9292_y0);
  and_gate and_gate_h_u_cla32_and9293_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9293_y0);
  and_gate and_gate_h_u_cla32_and9294_y0(h_u_cla32_and9293_y0, h_u_cla32_and9292_y0, h_u_cla32_and9294_y0);
  and_gate and_gate_h_u_cla32_and9295_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9295_y0);
  and_gate and_gate_h_u_cla32_and9296_y0(h_u_cla32_and9295_y0, h_u_cla32_and9294_y0, h_u_cla32_and9296_y0);
  and_gate and_gate_h_u_cla32_and9297_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9297_y0);
  and_gate and_gate_h_u_cla32_and9298_y0(h_u_cla32_and9297_y0, h_u_cla32_and9296_y0, h_u_cla32_and9298_y0);
  and_gate and_gate_h_u_cla32_and9299_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9299_y0);
  and_gate and_gate_h_u_cla32_and9300_y0(h_u_cla32_and9299_y0, h_u_cla32_and9298_y0, h_u_cla32_and9300_y0);
  and_gate and_gate_h_u_cla32_and9301_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9301_y0);
  and_gate and_gate_h_u_cla32_and9302_y0(h_u_cla32_and9301_y0, h_u_cla32_and9300_y0, h_u_cla32_and9302_y0);
  and_gate and_gate_h_u_cla32_and9303_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9303_y0);
  and_gate and_gate_h_u_cla32_and9304_y0(h_u_cla32_and9303_y0, h_u_cla32_and9302_y0, h_u_cla32_and9304_y0);
  and_gate and_gate_h_u_cla32_and9305_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9305_y0);
  and_gate and_gate_h_u_cla32_and9306_y0(h_u_cla32_and9305_y0, h_u_cla32_and9304_y0, h_u_cla32_and9306_y0);
  and_gate and_gate_h_u_cla32_and9307_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9307_y0);
  and_gate and_gate_h_u_cla32_and9308_y0(h_u_cla32_and9307_y0, h_u_cla32_and9306_y0, h_u_cla32_and9308_y0);
  and_gate and_gate_h_u_cla32_and9309_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and9309_y0);
  and_gate and_gate_h_u_cla32_and9310_y0(h_u_cla32_and9309_y0, h_u_cla32_and9308_y0, h_u_cla32_and9310_y0);
  and_gate and_gate_h_u_cla32_and9311_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9311_y0);
  and_gate and_gate_h_u_cla32_and9312_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9312_y0);
  and_gate and_gate_h_u_cla32_and9313_y0(h_u_cla32_and9312_y0, h_u_cla32_and9311_y0, h_u_cla32_and9313_y0);
  and_gate and_gate_h_u_cla32_and9314_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9314_y0);
  and_gate and_gate_h_u_cla32_and9315_y0(h_u_cla32_and9314_y0, h_u_cla32_and9313_y0, h_u_cla32_and9315_y0);
  and_gate and_gate_h_u_cla32_and9316_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9316_y0);
  and_gate and_gate_h_u_cla32_and9317_y0(h_u_cla32_and9316_y0, h_u_cla32_and9315_y0, h_u_cla32_and9317_y0);
  and_gate and_gate_h_u_cla32_and9318_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9318_y0);
  and_gate and_gate_h_u_cla32_and9319_y0(h_u_cla32_and9318_y0, h_u_cla32_and9317_y0, h_u_cla32_and9319_y0);
  and_gate and_gate_h_u_cla32_and9320_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9320_y0);
  and_gate and_gate_h_u_cla32_and9321_y0(h_u_cla32_and9320_y0, h_u_cla32_and9319_y0, h_u_cla32_and9321_y0);
  and_gate and_gate_h_u_cla32_and9322_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9322_y0);
  and_gate and_gate_h_u_cla32_and9323_y0(h_u_cla32_and9322_y0, h_u_cla32_and9321_y0, h_u_cla32_and9323_y0);
  and_gate and_gate_h_u_cla32_and9324_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9324_y0);
  and_gate and_gate_h_u_cla32_and9325_y0(h_u_cla32_and9324_y0, h_u_cla32_and9323_y0, h_u_cla32_and9325_y0);
  and_gate and_gate_h_u_cla32_and9326_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9326_y0);
  and_gate and_gate_h_u_cla32_and9327_y0(h_u_cla32_and9326_y0, h_u_cla32_and9325_y0, h_u_cla32_and9327_y0);
  and_gate and_gate_h_u_cla32_and9328_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9328_y0);
  and_gate and_gate_h_u_cla32_and9329_y0(h_u_cla32_and9328_y0, h_u_cla32_and9327_y0, h_u_cla32_and9329_y0);
  and_gate and_gate_h_u_cla32_and9330_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9330_y0);
  and_gate and_gate_h_u_cla32_and9331_y0(h_u_cla32_and9330_y0, h_u_cla32_and9329_y0, h_u_cla32_and9331_y0);
  and_gate and_gate_h_u_cla32_and9332_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and9332_y0);
  and_gate and_gate_h_u_cla32_and9333_y0(h_u_cla32_and9332_y0, h_u_cla32_and9331_y0, h_u_cla32_and9333_y0);
  and_gate and_gate_h_u_cla32_and9334_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9334_y0);
  and_gate and_gate_h_u_cla32_and9335_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9335_y0);
  and_gate and_gate_h_u_cla32_and9336_y0(h_u_cla32_and9335_y0, h_u_cla32_and9334_y0, h_u_cla32_and9336_y0);
  and_gate and_gate_h_u_cla32_and9337_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9337_y0);
  and_gate and_gate_h_u_cla32_and9338_y0(h_u_cla32_and9337_y0, h_u_cla32_and9336_y0, h_u_cla32_and9338_y0);
  and_gate and_gate_h_u_cla32_and9339_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9339_y0);
  and_gate and_gate_h_u_cla32_and9340_y0(h_u_cla32_and9339_y0, h_u_cla32_and9338_y0, h_u_cla32_and9340_y0);
  and_gate and_gate_h_u_cla32_and9341_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9341_y0);
  and_gate and_gate_h_u_cla32_and9342_y0(h_u_cla32_and9341_y0, h_u_cla32_and9340_y0, h_u_cla32_and9342_y0);
  and_gate and_gate_h_u_cla32_and9343_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9343_y0);
  and_gate and_gate_h_u_cla32_and9344_y0(h_u_cla32_and9343_y0, h_u_cla32_and9342_y0, h_u_cla32_and9344_y0);
  and_gate and_gate_h_u_cla32_and9345_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9345_y0);
  and_gate and_gate_h_u_cla32_and9346_y0(h_u_cla32_and9345_y0, h_u_cla32_and9344_y0, h_u_cla32_and9346_y0);
  and_gate and_gate_h_u_cla32_and9347_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9347_y0);
  and_gate and_gate_h_u_cla32_and9348_y0(h_u_cla32_and9347_y0, h_u_cla32_and9346_y0, h_u_cla32_and9348_y0);
  and_gate and_gate_h_u_cla32_and9349_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9349_y0);
  and_gate and_gate_h_u_cla32_and9350_y0(h_u_cla32_and9349_y0, h_u_cla32_and9348_y0, h_u_cla32_and9350_y0);
  and_gate and_gate_h_u_cla32_and9351_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9351_y0);
  and_gate and_gate_h_u_cla32_and9352_y0(h_u_cla32_and9351_y0, h_u_cla32_and9350_y0, h_u_cla32_and9352_y0);
  and_gate and_gate_h_u_cla32_and9353_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and9353_y0);
  and_gate and_gate_h_u_cla32_and9354_y0(h_u_cla32_and9353_y0, h_u_cla32_and9352_y0, h_u_cla32_and9354_y0);
  and_gate and_gate_h_u_cla32_and9355_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9355_y0);
  and_gate and_gate_h_u_cla32_and9356_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9356_y0);
  and_gate and_gate_h_u_cla32_and9357_y0(h_u_cla32_and9356_y0, h_u_cla32_and9355_y0, h_u_cla32_and9357_y0);
  and_gate and_gate_h_u_cla32_and9358_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9358_y0);
  and_gate and_gate_h_u_cla32_and9359_y0(h_u_cla32_and9358_y0, h_u_cla32_and9357_y0, h_u_cla32_and9359_y0);
  and_gate and_gate_h_u_cla32_and9360_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9360_y0);
  and_gate and_gate_h_u_cla32_and9361_y0(h_u_cla32_and9360_y0, h_u_cla32_and9359_y0, h_u_cla32_and9361_y0);
  and_gate and_gate_h_u_cla32_and9362_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9362_y0);
  and_gate and_gate_h_u_cla32_and9363_y0(h_u_cla32_and9362_y0, h_u_cla32_and9361_y0, h_u_cla32_and9363_y0);
  and_gate and_gate_h_u_cla32_and9364_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9364_y0);
  and_gate and_gate_h_u_cla32_and9365_y0(h_u_cla32_and9364_y0, h_u_cla32_and9363_y0, h_u_cla32_and9365_y0);
  and_gate and_gate_h_u_cla32_and9366_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9366_y0);
  and_gate and_gate_h_u_cla32_and9367_y0(h_u_cla32_and9366_y0, h_u_cla32_and9365_y0, h_u_cla32_and9367_y0);
  and_gate and_gate_h_u_cla32_and9368_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9368_y0);
  and_gate and_gate_h_u_cla32_and9369_y0(h_u_cla32_and9368_y0, h_u_cla32_and9367_y0, h_u_cla32_and9369_y0);
  and_gate and_gate_h_u_cla32_and9370_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9370_y0);
  and_gate and_gate_h_u_cla32_and9371_y0(h_u_cla32_and9370_y0, h_u_cla32_and9369_y0, h_u_cla32_and9371_y0);
  and_gate and_gate_h_u_cla32_and9372_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and9372_y0);
  and_gate and_gate_h_u_cla32_and9373_y0(h_u_cla32_and9372_y0, h_u_cla32_and9371_y0, h_u_cla32_and9373_y0);
  and_gate and_gate_h_u_cla32_and9374_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9374_y0);
  and_gate and_gate_h_u_cla32_and9375_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9375_y0);
  and_gate and_gate_h_u_cla32_and9376_y0(h_u_cla32_and9375_y0, h_u_cla32_and9374_y0, h_u_cla32_and9376_y0);
  and_gate and_gate_h_u_cla32_and9377_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9377_y0);
  and_gate and_gate_h_u_cla32_and9378_y0(h_u_cla32_and9377_y0, h_u_cla32_and9376_y0, h_u_cla32_and9378_y0);
  and_gate and_gate_h_u_cla32_and9379_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9379_y0);
  and_gate and_gate_h_u_cla32_and9380_y0(h_u_cla32_and9379_y0, h_u_cla32_and9378_y0, h_u_cla32_and9380_y0);
  and_gate and_gate_h_u_cla32_and9381_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9381_y0);
  and_gate and_gate_h_u_cla32_and9382_y0(h_u_cla32_and9381_y0, h_u_cla32_and9380_y0, h_u_cla32_and9382_y0);
  and_gate and_gate_h_u_cla32_and9383_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9383_y0);
  and_gate and_gate_h_u_cla32_and9384_y0(h_u_cla32_and9383_y0, h_u_cla32_and9382_y0, h_u_cla32_and9384_y0);
  and_gate and_gate_h_u_cla32_and9385_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9385_y0);
  and_gate and_gate_h_u_cla32_and9386_y0(h_u_cla32_and9385_y0, h_u_cla32_and9384_y0, h_u_cla32_and9386_y0);
  and_gate and_gate_h_u_cla32_and9387_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9387_y0);
  and_gate and_gate_h_u_cla32_and9388_y0(h_u_cla32_and9387_y0, h_u_cla32_and9386_y0, h_u_cla32_and9388_y0);
  and_gate and_gate_h_u_cla32_and9389_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and9389_y0);
  and_gate and_gate_h_u_cla32_and9390_y0(h_u_cla32_and9389_y0, h_u_cla32_and9388_y0, h_u_cla32_and9390_y0);
  and_gate and_gate_h_u_cla32_and9391_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9391_y0);
  and_gate and_gate_h_u_cla32_and9392_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9392_y0);
  and_gate and_gate_h_u_cla32_and9393_y0(h_u_cla32_and9392_y0, h_u_cla32_and9391_y0, h_u_cla32_and9393_y0);
  and_gate and_gate_h_u_cla32_and9394_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9394_y0);
  and_gate and_gate_h_u_cla32_and9395_y0(h_u_cla32_and9394_y0, h_u_cla32_and9393_y0, h_u_cla32_and9395_y0);
  and_gate and_gate_h_u_cla32_and9396_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9396_y0);
  and_gate and_gate_h_u_cla32_and9397_y0(h_u_cla32_and9396_y0, h_u_cla32_and9395_y0, h_u_cla32_and9397_y0);
  and_gate and_gate_h_u_cla32_and9398_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9398_y0);
  and_gate and_gate_h_u_cla32_and9399_y0(h_u_cla32_and9398_y0, h_u_cla32_and9397_y0, h_u_cla32_and9399_y0);
  and_gate and_gate_h_u_cla32_and9400_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9400_y0);
  and_gate and_gate_h_u_cla32_and9401_y0(h_u_cla32_and9400_y0, h_u_cla32_and9399_y0, h_u_cla32_and9401_y0);
  and_gate and_gate_h_u_cla32_and9402_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9402_y0);
  and_gate and_gate_h_u_cla32_and9403_y0(h_u_cla32_and9402_y0, h_u_cla32_and9401_y0, h_u_cla32_and9403_y0);
  and_gate and_gate_h_u_cla32_and9404_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and9404_y0);
  and_gate and_gate_h_u_cla32_and9405_y0(h_u_cla32_and9404_y0, h_u_cla32_and9403_y0, h_u_cla32_and9405_y0);
  and_gate and_gate_h_u_cla32_and9406_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9406_y0);
  and_gate and_gate_h_u_cla32_and9407_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9407_y0);
  and_gate and_gate_h_u_cla32_and9408_y0(h_u_cla32_and9407_y0, h_u_cla32_and9406_y0, h_u_cla32_and9408_y0);
  and_gate and_gate_h_u_cla32_and9409_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9409_y0);
  and_gate and_gate_h_u_cla32_and9410_y0(h_u_cla32_and9409_y0, h_u_cla32_and9408_y0, h_u_cla32_and9410_y0);
  and_gate and_gate_h_u_cla32_and9411_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9411_y0);
  and_gate and_gate_h_u_cla32_and9412_y0(h_u_cla32_and9411_y0, h_u_cla32_and9410_y0, h_u_cla32_and9412_y0);
  and_gate and_gate_h_u_cla32_and9413_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9413_y0);
  and_gate and_gate_h_u_cla32_and9414_y0(h_u_cla32_and9413_y0, h_u_cla32_and9412_y0, h_u_cla32_and9414_y0);
  and_gate and_gate_h_u_cla32_and9415_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9415_y0);
  and_gate and_gate_h_u_cla32_and9416_y0(h_u_cla32_and9415_y0, h_u_cla32_and9414_y0, h_u_cla32_and9416_y0);
  and_gate and_gate_h_u_cla32_and9417_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and9417_y0);
  and_gate and_gate_h_u_cla32_and9418_y0(h_u_cla32_and9417_y0, h_u_cla32_and9416_y0, h_u_cla32_and9418_y0);
  and_gate and_gate_h_u_cla32_and9419_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and9419_y0);
  and_gate and_gate_h_u_cla32_and9420_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and9420_y0);
  and_gate and_gate_h_u_cla32_and9421_y0(h_u_cla32_and9420_y0, h_u_cla32_and9419_y0, h_u_cla32_and9421_y0);
  and_gate and_gate_h_u_cla32_and9422_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and9422_y0);
  and_gate and_gate_h_u_cla32_and9423_y0(h_u_cla32_and9422_y0, h_u_cla32_and9421_y0, h_u_cla32_and9423_y0);
  and_gate and_gate_h_u_cla32_and9424_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and9424_y0);
  and_gate and_gate_h_u_cla32_and9425_y0(h_u_cla32_and9424_y0, h_u_cla32_and9423_y0, h_u_cla32_and9425_y0);
  and_gate and_gate_h_u_cla32_and9426_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and9426_y0);
  and_gate and_gate_h_u_cla32_and9427_y0(h_u_cla32_and9426_y0, h_u_cla32_and9425_y0, h_u_cla32_and9427_y0);
  and_gate and_gate_h_u_cla32_and9428_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and9428_y0);
  and_gate and_gate_h_u_cla32_and9429_y0(h_u_cla32_and9428_y0, h_u_cla32_and9427_y0, h_u_cla32_and9429_y0);
  and_gate and_gate_h_u_cla32_and9430_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and9430_y0);
  and_gate and_gate_h_u_cla32_and9431_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and9431_y0);
  and_gate and_gate_h_u_cla32_and9432_y0(h_u_cla32_and9431_y0, h_u_cla32_and9430_y0, h_u_cla32_and9432_y0);
  and_gate and_gate_h_u_cla32_and9433_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and9433_y0);
  and_gate and_gate_h_u_cla32_and9434_y0(h_u_cla32_and9433_y0, h_u_cla32_and9432_y0, h_u_cla32_and9434_y0);
  and_gate and_gate_h_u_cla32_and9435_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and9435_y0);
  and_gate and_gate_h_u_cla32_and9436_y0(h_u_cla32_and9435_y0, h_u_cla32_and9434_y0, h_u_cla32_and9436_y0);
  and_gate and_gate_h_u_cla32_and9437_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and9437_y0);
  and_gate and_gate_h_u_cla32_and9438_y0(h_u_cla32_and9437_y0, h_u_cla32_and9436_y0, h_u_cla32_and9438_y0);
  and_gate and_gate_h_u_cla32_and9439_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and9439_y0);
  and_gate and_gate_h_u_cla32_and9440_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and9440_y0);
  and_gate and_gate_h_u_cla32_and9441_y0(h_u_cla32_and9440_y0, h_u_cla32_and9439_y0, h_u_cla32_and9441_y0);
  and_gate and_gate_h_u_cla32_and9442_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and9442_y0);
  and_gate and_gate_h_u_cla32_and9443_y0(h_u_cla32_and9442_y0, h_u_cla32_and9441_y0, h_u_cla32_and9443_y0);
  and_gate and_gate_h_u_cla32_and9444_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and9444_y0);
  and_gate and_gate_h_u_cla32_and9445_y0(h_u_cla32_and9444_y0, h_u_cla32_and9443_y0, h_u_cla32_and9445_y0);
  and_gate and_gate_h_u_cla32_and9446_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and9446_y0);
  and_gate and_gate_h_u_cla32_and9447_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and9447_y0);
  and_gate and_gate_h_u_cla32_and9448_y0(h_u_cla32_and9447_y0, h_u_cla32_and9446_y0, h_u_cla32_and9448_y0);
  and_gate and_gate_h_u_cla32_and9449_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and9449_y0);
  and_gate and_gate_h_u_cla32_and9450_y0(h_u_cla32_and9449_y0, h_u_cla32_and9448_y0, h_u_cla32_and9450_y0);
  and_gate and_gate_h_u_cla32_and9451_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and9451_y0);
  and_gate and_gate_h_u_cla32_and9452_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and9452_y0);
  and_gate and_gate_h_u_cla32_and9453_y0(h_u_cla32_and9452_y0, h_u_cla32_and9451_y0, h_u_cla32_and9453_y0);
  and_gate and_gate_h_u_cla32_and9454_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_and9454_y0);
  or_gate or_gate_h_u_cla32_or435_y0(h_u_cla32_and9454_y0, h_u_cla32_and8613_y0, h_u_cla32_or435_y0);
  or_gate or_gate_h_u_cla32_or436_y0(h_u_cla32_or435_y0, h_u_cla32_and8670_y0, h_u_cla32_or436_y0);
  or_gate or_gate_h_u_cla32_or437_y0(h_u_cla32_or436_y0, h_u_cla32_and8725_y0, h_u_cla32_or437_y0);
  or_gate or_gate_h_u_cla32_or438_y0(h_u_cla32_or437_y0, h_u_cla32_and8778_y0, h_u_cla32_or438_y0);
  or_gate or_gate_h_u_cla32_or439_y0(h_u_cla32_or438_y0, h_u_cla32_and8829_y0, h_u_cla32_or439_y0);
  or_gate or_gate_h_u_cla32_or440_y0(h_u_cla32_or439_y0, h_u_cla32_and8878_y0, h_u_cla32_or440_y0);
  or_gate or_gate_h_u_cla32_or441_y0(h_u_cla32_or440_y0, h_u_cla32_and8925_y0, h_u_cla32_or441_y0);
  or_gate or_gate_h_u_cla32_or442_y0(h_u_cla32_or441_y0, h_u_cla32_and8970_y0, h_u_cla32_or442_y0);
  or_gate or_gate_h_u_cla32_or443_y0(h_u_cla32_or442_y0, h_u_cla32_and9013_y0, h_u_cla32_or443_y0);
  or_gate or_gate_h_u_cla32_or444_y0(h_u_cla32_or443_y0, h_u_cla32_and9054_y0, h_u_cla32_or444_y0);
  or_gate or_gate_h_u_cla32_or445_y0(h_u_cla32_or444_y0, h_u_cla32_and9093_y0, h_u_cla32_or445_y0);
  or_gate or_gate_h_u_cla32_or446_y0(h_u_cla32_or445_y0, h_u_cla32_and9130_y0, h_u_cla32_or446_y0);
  or_gate or_gate_h_u_cla32_or447_y0(h_u_cla32_or446_y0, h_u_cla32_and9165_y0, h_u_cla32_or447_y0);
  or_gate or_gate_h_u_cla32_or448_y0(h_u_cla32_or447_y0, h_u_cla32_and9198_y0, h_u_cla32_or448_y0);
  or_gate or_gate_h_u_cla32_or449_y0(h_u_cla32_or448_y0, h_u_cla32_and9229_y0, h_u_cla32_or449_y0);
  or_gate or_gate_h_u_cla32_or450_y0(h_u_cla32_or449_y0, h_u_cla32_and9258_y0, h_u_cla32_or450_y0);
  or_gate or_gate_h_u_cla32_or451_y0(h_u_cla32_or450_y0, h_u_cla32_and9285_y0, h_u_cla32_or451_y0);
  or_gate or_gate_h_u_cla32_or452_y0(h_u_cla32_or451_y0, h_u_cla32_and9310_y0, h_u_cla32_or452_y0);
  or_gate or_gate_h_u_cla32_or453_y0(h_u_cla32_or452_y0, h_u_cla32_and9333_y0, h_u_cla32_or453_y0);
  or_gate or_gate_h_u_cla32_or454_y0(h_u_cla32_or453_y0, h_u_cla32_and9354_y0, h_u_cla32_or454_y0);
  or_gate or_gate_h_u_cla32_or455_y0(h_u_cla32_or454_y0, h_u_cla32_and9373_y0, h_u_cla32_or455_y0);
  or_gate or_gate_h_u_cla32_or456_y0(h_u_cla32_or455_y0, h_u_cla32_and9390_y0, h_u_cla32_or456_y0);
  or_gate or_gate_h_u_cla32_or457_y0(h_u_cla32_or456_y0, h_u_cla32_and9405_y0, h_u_cla32_or457_y0);
  or_gate or_gate_h_u_cla32_or458_y0(h_u_cla32_or457_y0, h_u_cla32_and9418_y0, h_u_cla32_or458_y0);
  or_gate or_gate_h_u_cla32_or459_y0(h_u_cla32_or458_y0, h_u_cla32_and9429_y0, h_u_cla32_or459_y0);
  or_gate or_gate_h_u_cla32_or460_y0(h_u_cla32_or459_y0, h_u_cla32_and9438_y0, h_u_cla32_or460_y0);
  or_gate or_gate_h_u_cla32_or461_y0(h_u_cla32_or460_y0, h_u_cla32_and9445_y0, h_u_cla32_or461_y0);
  or_gate or_gate_h_u_cla32_or462_y0(h_u_cla32_or461_y0, h_u_cla32_and9450_y0, h_u_cla32_or462_y0);
  or_gate or_gate_h_u_cla32_or463_y0(h_u_cla32_or462_y0, h_u_cla32_and9453_y0, h_u_cla32_or463_y0);
  or_gate or_gate_h_u_cla32_or464_y0(h_u_cla32_pg_logic29_y1, h_u_cla32_or463_y0, h_u_cla32_or464_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic30_y0(a_30, b_30, h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic30_y1, h_u_cla32_pg_logic30_y2);
  xor_gate xor_gate_h_u_cla32_xor30_y0(h_u_cla32_pg_logic30_y2, h_u_cla32_or464_y0, h_u_cla32_xor30_y0);
  and_gate and_gate_h_u_cla32_and9455_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and9455_y0);
  and_gate and_gate_h_u_cla32_and9456_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and9456_y0);
  and_gate and_gate_h_u_cla32_and9457_y0(h_u_cla32_and9456_y0, h_u_cla32_and9455_y0, h_u_cla32_and9457_y0);
  and_gate and_gate_h_u_cla32_and9458_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and9458_y0);
  and_gate and_gate_h_u_cla32_and9459_y0(h_u_cla32_and9458_y0, h_u_cla32_and9457_y0, h_u_cla32_and9459_y0);
  and_gate and_gate_h_u_cla32_and9460_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and9460_y0);
  and_gate and_gate_h_u_cla32_and9461_y0(h_u_cla32_and9460_y0, h_u_cla32_and9459_y0, h_u_cla32_and9461_y0);
  and_gate and_gate_h_u_cla32_and9462_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and9462_y0);
  and_gate and_gate_h_u_cla32_and9463_y0(h_u_cla32_and9462_y0, h_u_cla32_and9461_y0, h_u_cla32_and9463_y0);
  and_gate and_gate_h_u_cla32_and9464_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and9464_y0);
  and_gate and_gate_h_u_cla32_and9465_y0(h_u_cla32_and9464_y0, h_u_cla32_and9463_y0, h_u_cla32_and9465_y0);
  and_gate and_gate_h_u_cla32_and9466_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and9466_y0);
  and_gate and_gate_h_u_cla32_and9467_y0(h_u_cla32_and9466_y0, h_u_cla32_and9465_y0, h_u_cla32_and9467_y0);
  and_gate and_gate_h_u_cla32_and9468_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and9468_y0);
  and_gate and_gate_h_u_cla32_and9469_y0(h_u_cla32_and9468_y0, h_u_cla32_and9467_y0, h_u_cla32_and9469_y0);
  and_gate and_gate_h_u_cla32_and9470_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and9470_y0);
  and_gate and_gate_h_u_cla32_and9471_y0(h_u_cla32_and9470_y0, h_u_cla32_and9469_y0, h_u_cla32_and9471_y0);
  and_gate and_gate_h_u_cla32_and9472_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and9472_y0);
  and_gate and_gate_h_u_cla32_and9473_y0(h_u_cla32_and9472_y0, h_u_cla32_and9471_y0, h_u_cla32_and9473_y0);
  and_gate and_gate_h_u_cla32_and9474_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and9474_y0);
  and_gate and_gate_h_u_cla32_and9475_y0(h_u_cla32_and9474_y0, h_u_cla32_and9473_y0, h_u_cla32_and9475_y0);
  and_gate and_gate_h_u_cla32_and9476_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and9476_y0);
  and_gate and_gate_h_u_cla32_and9477_y0(h_u_cla32_and9476_y0, h_u_cla32_and9475_y0, h_u_cla32_and9477_y0);
  and_gate and_gate_h_u_cla32_and9478_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and9478_y0);
  and_gate and_gate_h_u_cla32_and9479_y0(h_u_cla32_and9478_y0, h_u_cla32_and9477_y0, h_u_cla32_and9479_y0);
  and_gate and_gate_h_u_cla32_and9480_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and9480_y0);
  and_gate and_gate_h_u_cla32_and9481_y0(h_u_cla32_and9480_y0, h_u_cla32_and9479_y0, h_u_cla32_and9481_y0);
  and_gate and_gate_h_u_cla32_and9482_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and9482_y0);
  and_gate and_gate_h_u_cla32_and9483_y0(h_u_cla32_and9482_y0, h_u_cla32_and9481_y0, h_u_cla32_and9483_y0);
  and_gate and_gate_h_u_cla32_and9484_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and9484_y0);
  and_gate and_gate_h_u_cla32_and9485_y0(h_u_cla32_and9484_y0, h_u_cla32_and9483_y0, h_u_cla32_and9485_y0);
  and_gate and_gate_h_u_cla32_and9486_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and9486_y0);
  and_gate and_gate_h_u_cla32_and9487_y0(h_u_cla32_and9486_y0, h_u_cla32_and9485_y0, h_u_cla32_and9487_y0);
  and_gate and_gate_h_u_cla32_and9488_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and9488_y0);
  and_gate and_gate_h_u_cla32_and9489_y0(h_u_cla32_and9488_y0, h_u_cla32_and9487_y0, h_u_cla32_and9489_y0);
  and_gate and_gate_h_u_cla32_and9490_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and9490_y0);
  and_gate and_gate_h_u_cla32_and9491_y0(h_u_cla32_and9490_y0, h_u_cla32_and9489_y0, h_u_cla32_and9491_y0);
  and_gate and_gate_h_u_cla32_and9492_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and9492_y0);
  and_gate and_gate_h_u_cla32_and9493_y0(h_u_cla32_and9492_y0, h_u_cla32_and9491_y0, h_u_cla32_and9493_y0);
  and_gate and_gate_h_u_cla32_and9494_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and9494_y0);
  and_gate and_gate_h_u_cla32_and9495_y0(h_u_cla32_and9494_y0, h_u_cla32_and9493_y0, h_u_cla32_and9495_y0);
  and_gate and_gate_h_u_cla32_and9496_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and9496_y0);
  and_gate and_gate_h_u_cla32_and9497_y0(h_u_cla32_and9496_y0, h_u_cla32_and9495_y0, h_u_cla32_and9497_y0);
  and_gate and_gate_h_u_cla32_and9498_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and9498_y0);
  and_gate and_gate_h_u_cla32_and9499_y0(h_u_cla32_and9498_y0, h_u_cla32_and9497_y0, h_u_cla32_and9499_y0);
  and_gate and_gate_h_u_cla32_and9500_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and9500_y0);
  and_gate and_gate_h_u_cla32_and9501_y0(h_u_cla32_and9500_y0, h_u_cla32_and9499_y0, h_u_cla32_and9501_y0);
  and_gate and_gate_h_u_cla32_and9502_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and9502_y0);
  and_gate and_gate_h_u_cla32_and9503_y0(h_u_cla32_and9502_y0, h_u_cla32_and9501_y0, h_u_cla32_and9503_y0);
  and_gate and_gate_h_u_cla32_and9504_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and9504_y0);
  and_gate and_gate_h_u_cla32_and9505_y0(h_u_cla32_and9504_y0, h_u_cla32_and9503_y0, h_u_cla32_and9505_y0);
  and_gate and_gate_h_u_cla32_and9506_y0(h_u_cla32_pg_logic26_y0, constant_wire_0, h_u_cla32_and9506_y0);
  and_gate and_gate_h_u_cla32_and9507_y0(h_u_cla32_and9506_y0, h_u_cla32_and9505_y0, h_u_cla32_and9507_y0);
  and_gate and_gate_h_u_cla32_and9508_y0(h_u_cla32_pg_logic27_y0, constant_wire_0, h_u_cla32_and9508_y0);
  and_gate and_gate_h_u_cla32_and9509_y0(h_u_cla32_and9508_y0, h_u_cla32_and9507_y0, h_u_cla32_and9509_y0);
  and_gate and_gate_h_u_cla32_and9510_y0(h_u_cla32_pg_logic28_y0, constant_wire_0, h_u_cla32_and9510_y0);
  and_gate and_gate_h_u_cla32_and9511_y0(h_u_cla32_and9510_y0, h_u_cla32_and9509_y0, h_u_cla32_and9511_y0);
  and_gate and_gate_h_u_cla32_and9512_y0(h_u_cla32_pg_logic29_y0, constant_wire_0, h_u_cla32_and9512_y0);
  and_gate and_gate_h_u_cla32_and9513_y0(h_u_cla32_and9512_y0, h_u_cla32_and9511_y0, h_u_cla32_and9513_y0);
  and_gate and_gate_h_u_cla32_and9514_y0(h_u_cla32_pg_logic30_y0, constant_wire_0, h_u_cla32_and9514_y0);
  and_gate and_gate_h_u_cla32_and9515_y0(h_u_cla32_and9514_y0, h_u_cla32_and9513_y0, h_u_cla32_and9515_y0);
  and_gate and_gate_h_u_cla32_and9516_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9516_y0);
  and_gate and_gate_h_u_cla32_and9517_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9517_y0);
  and_gate and_gate_h_u_cla32_and9518_y0(h_u_cla32_and9517_y0, h_u_cla32_and9516_y0, h_u_cla32_and9518_y0);
  and_gate and_gate_h_u_cla32_and9519_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9519_y0);
  and_gate and_gate_h_u_cla32_and9520_y0(h_u_cla32_and9519_y0, h_u_cla32_and9518_y0, h_u_cla32_and9520_y0);
  and_gate and_gate_h_u_cla32_and9521_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9521_y0);
  and_gate and_gate_h_u_cla32_and9522_y0(h_u_cla32_and9521_y0, h_u_cla32_and9520_y0, h_u_cla32_and9522_y0);
  and_gate and_gate_h_u_cla32_and9523_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9523_y0);
  and_gate and_gate_h_u_cla32_and9524_y0(h_u_cla32_and9523_y0, h_u_cla32_and9522_y0, h_u_cla32_and9524_y0);
  and_gate and_gate_h_u_cla32_and9525_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9525_y0);
  and_gate and_gate_h_u_cla32_and9526_y0(h_u_cla32_and9525_y0, h_u_cla32_and9524_y0, h_u_cla32_and9526_y0);
  and_gate and_gate_h_u_cla32_and9527_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9527_y0);
  and_gate and_gate_h_u_cla32_and9528_y0(h_u_cla32_and9527_y0, h_u_cla32_and9526_y0, h_u_cla32_and9528_y0);
  and_gate and_gate_h_u_cla32_and9529_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9529_y0);
  and_gate and_gate_h_u_cla32_and9530_y0(h_u_cla32_and9529_y0, h_u_cla32_and9528_y0, h_u_cla32_and9530_y0);
  and_gate and_gate_h_u_cla32_and9531_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9531_y0);
  and_gate and_gate_h_u_cla32_and9532_y0(h_u_cla32_and9531_y0, h_u_cla32_and9530_y0, h_u_cla32_and9532_y0);
  and_gate and_gate_h_u_cla32_and9533_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9533_y0);
  and_gate and_gate_h_u_cla32_and9534_y0(h_u_cla32_and9533_y0, h_u_cla32_and9532_y0, h_u_cla32_and9534_y0);
  and_gate and_gate_h_u_cla32_and9535_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9535_y0);
  and_gate and_gate_h_u_cla32_and9536_y0(h_u_cla32_and9535_y0, h_u_cla32_and9534_y0, h_u_cla32_and9536_y0);
  and_gate and_gate_h_u_cla32_and9537_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9537_y0);
  and_gate and_gate_h_u_cla32_and9538_y0(h_u_cla32_and9537_y0, h_u_cla32_and9536_y0, h_u_cla32_and9538_y0);
  and_gate and_gate_h_u_cla32_and9539_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9539_y0);
  and_gate and_gate_h_u_cla32_and9540_y0(h_u_cla32_and9539_y0, h_u_cla32_and9538_y0, h_u_cla32_and9540_y0);
  and_gate and_gate_h_u_cla32_and9541_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9541_y0);
  and_gate and_gate_h_u_cla32_and9542_y0(h_u_cla32_and9541_y0, h_u_cla32_and9540_y0, h_u_cla32_and9542_y0);
  and_gate and_gate_h_u_cla32_and9543_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9543_y0);
  and_gate and_gate_h_u_cla32_and9544_y0(h_u_cla32_and9543_y0, h_u_cla32_and9542_y0, h_u_cla32_and9544_y0);
  and_gate and_gate_h_u_cla32_and9545_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9545_y0);
  and_gate and_gate_h_u_cla32_and9546_y0(h_u_cla32_and9545_y0, h_u_cla32_and9544_y0, h_u_cla32_and9546_y0);
  and_gate and_gate_h_u_cla32_and9547_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9547_y0);
  and_gate and_gate_h_u_cla32_and9548_y0(h_u_cla32_and9547_y0, h_u_cla32_and9546_y0, h_u_cla32_and9548_y0);
  and_gate and_gate_h_u_cla32_and9549_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9549_y0);
  and_gate and_gate_h_u_cla32_and9550_y0(h_u_cla32_and9549_y0, h_u_cla32_and9548_y0, h_u_cla32_and9550_y0);
  and_gate and_gate_h_u_cla32_and9551_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9551_y0);
  and_gate and_gate_h_u_cla32_and9552_y0(h_u_cla32_and9551_y0, h_u_cla32_and9550_y0, h_u_cla32_and9552_y0);
  and_gate and_gate_h_u_cla32_and9553_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9553_y0);
  and_gate and_gate_h_u_cla32_and9554_y0(h_u_cla32_and9553_y0, h_u_cla32_and9552_y0, h_u_cla32_and9554_y0);
  and_gate and_gate_h_u_cla32_and9555_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9555_y0);
  and_gate and_gate_h_u_cla32_and9556_y0(h_u_cla32_and9555_y0, h_u_cla32_and9554_y0, h_u_cla32_and9556_y0);
  and_gate and_gate_h_u_cla32_and9557_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9557_y0);
  and_gate and_gate_h_u_cla32_and9558_y0(h_u_cla32_and9557_y0, h_u_cla32_and9556_y0, h_u_cla32_and9558_y0);
  and_gate and_gate_h_u_cla32_and9559_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9559_y0);
  and_gate and_gate_h_u_cla32_and9560_y0(h_u_cla32_and9559_y0, h_u_cla32_and9558_y0, h_u_cla32_and9560_y0);
  and_gate and_gate_h_u_cla32_and9561_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9561_y0);
  and_gate and_gate_h_u_cla32_and9562_y0(h_u_cla32_and9561_y0, h_u_cla32_and9560_y0, h_u_cla32_and9562_y0);
  and_gate and_gate_h_u_cla32_and9563_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9563_y0);
  and_gate and_gate_h_u_cla32_and9564_y0(h_u_cla32_and9563_y0, h_u_cla32_and9562_y0, h_u_cla32_and9564_y0);
  and_gate and_gate_h_u_cla32_and9565_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9565_y0);
  and_gate and_gate_h_u_cla32_and9566_y0(h_u_cla32_and9565_y0, h_u_cla32_and9564_y0, h_u_cla32_and9566_y0);
  and_gate and_gate_h_u_cla32_and9567_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9567_y0);
  and_gate and_gate_h_u_cla32_and9568_y0(h_u_cla32_and9567_y0, h_u_cla32_and9566_y0, h_u_cla32_and9568_y0);
  and_gate and_gate_h_u_cla32_and9569_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9569_y0);
  and_gate and_gate_h_u_cla32_and9570_y0(h_u_cla32_and9569_y0, h_u_cla32_and9568_y0, h_u_cla32_and9570_y0);
  and_gate and_gate_h_u_cla32_and9571_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9571_y0);
  and_gate and_gate_h_u_cla32_and9572_y0(h_u_cla32_and9571_y0, h_u_cla32_and9570_y0, h_u_cla32_and9572_y0);
  and_gate and_gate_h_u_cla32_and9573_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and9573_y0);
  and_gate and_gate_h_u_cla32_and9574_y0(h_u_cla32_and9573_y0, h_u_cla32_and9572_y0, h_u_cla32_and9574_y0);
  and_gate and_gate_h_u_cla32_and9575_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9575_y0);
  and_gate and_gate_h_u_cla32_and9576_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9576_y0);
  and_gate and_gate_h_u_cla32_and9577_y0(h_u_cla32_and9576_y0, h_u_cla32_and9575_y0, h_u_cla32_and9577_y0);
  and_gate and_gate_h_u_cla32_and9578_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9578_y0);
  and_gate and_gate_h_u_cla32_and9579_y0(h_u_cla32_and9578_y0, h_u_cla32_and9577_y0, h_u_cla32_and9579_y0);
  and_gate and_gate_h_u_cla32_and9580_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9580_y0);
  and_gate and_gate_h_u_cla32_and9581_y0(h_u_cla32_and9580_y0, h_u_cla32_and9579_y0, h_u_cla32_and9581_y0);
  and_gate and_gate_h_u_cla32_and9582_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9582_y0);
  and_gate and_gate_h_u_cla32_and9583_y0(h_u_cla32_and9582_y0, h_u_cla32_and9581_y0, h_u_cla32_and9583_y0);
  and_gate and_gate_h_u_cla32_and9584_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9584_y0);
  and_gate and_gate_h_u_cla32_and9585_y0(h_u_cla32_and9584_y0, h_u_cla32_and9583_y0, h_u_cla32_and9585_y0);
  and_gate and_gate_h_u_cla32_and9586_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9586_y0);
  and_gate and_gate_h_u_cla32_and9587_y0(h_u_cla32_and9586_y0, h_u_cla32_and9585_y0, h_u_cla32_and9587_y0);
  and_gate and_gate_h_u_cla32_and9588_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9588_y0);
  and_gate and_gate_h_u_cla32_and9589_y0(h_u_cla32_and9588_y0, h_u_cla32_and9587_y0, h_u_cla32_and9589_y0);
  and_gate and_gate_h_u_cla32_and9590_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9590_y0);
  and_gate and_gate_h_u_cla32_and9591_y0(h_u_cla32_and9590_y0, h_u_cla32_and9589_y0, h_u_cla32_and9591_y0);
  and_gate and_gate_h_u_cla32_and9592_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9592_y0);
  and_gate and_gate_h_u_cla32_and9593_y0(h_u_cla32_and9592_y0, h_u_cla32_and9591_y0, h_u_cla32_and9593_y0);
  and_gate and_gate_h_u_cla32_and9594_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9594_y0);
  and_gate and_gate_h_u_cla32_and9595_y0(h_u_cla32_and9594_y0, h_u_cla32_and9593_y0, h_u_cla32_and9595_y0);
  and_gate and_gate_h_u_cla32_and9596_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9596_y0);
  and_gate and_gate_h_u_cla32_and9597_y0(h_u_cla32_and9596_y0, h_u_cla32_and9595_y0, h_u_cla32_and9597_y0);
  and_gate and_gate_h_u_cla32_and9598_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9598_y0);
  and_gate and_gate_h_u_cla32_and9599_y0(h_u_cla32_and9598_y0, h_u_cla32_and9597_y0, h_u_cla32_and9599_y0);
  and_gate and_gate_h_u_cla32_and9600_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9600_y0);
  and_gate and_gate_h_u_cla32_and9601_y0(h_u_cla32_and9600_y0, h_u_cla32_and9599_y0, h_u_cla32_and9601_y0);
  and_gate and_gate_h_u_cla32_and9602_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9602_y0);
  and_gate and_gate_h_u_cla32_and9603_y0(h_u_cla32_and9602_y0, h_u_cla32_and9601_y0, h_u_cla32_and9603_y0);
  and_gate and_gate_h_u_cla32_and9604_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9604_y0);
  and_gate and_gate_h_u_cla32_and9605_y0(h_u_cla32_and9604_y0, h_u_cla32_and9603_y0, h_u_cla32_and9605_y0);
  and_gate and_gate_h_u_cla32_and9606_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9606_y0);
  and_gate and_gate_h_u_cla32_and9607_y0(h_u_cla32_and9606_y0, h_u_cla32_and9605_y0, h_u_cla32_and9607_y0);
  and_gate and_gate_h_u_cla32_and9608_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9608_y0);
  and_gate and_gate_h_u_cla32_and9609_y0(h_u_cla32_and9608_y0, h_u_cla32_and9607_y0, h_u_cla32_and9609_y0);
  and_gate and_gate_h_u_cla32_and9610_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9610_y0);
  and_gate and_gate_h_u_cla32_and9611_y0(h_u_cla32_and9610_y0, h_u_cla32_and9609_y0, h_u_cla32_and9611_y0);
  and_gate and_gate_h_u_cla32_and9612_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9612_y0);
  and_gate and_gate_h_u_cla32_and9613_y0(h_u_cla32_and9612_y0, h_u_cla32_and9611_y0, h_u_cla32_and9613_y0);
  and_gate and_gate_h_u_cla32_and9614_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9614_y0);
  and_gate and_gate_h_u_cla32_and9615_y0(h_u_cla32_and9614_y0, h_u_cla32_and9613_y0, h_u_cla32_and9615_y0);
  and_gate and_gate_h_u_cla32_and9616_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9616_y0);
  and_gate and_gate_h_u_cla32_and9617_y0(h_u_cla32_and9616_y0, h_u_cla32_and9615_y0, h_u_cla32_and9617_y0);
  and_gate and_gate_h_u_cla32_and9618_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9618_y0);
  and_gate and_gate_h_u_cla32_and9619_y0(h_u_cla32_and9618_y0, h_u_cla32_and9617_y0, h_u_cla32_and9619_y0);
  and_gate and_gate_h_u_cla32_and9620_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9620_y0);
  and_gate and_gate_h_u_cla32_and9621_y0(h_u_cla32_and9620_y0, h_u_cla32_and9619_y0, h_u_cla32_and9621_y0);
  and_gate and_gate_h_u_cla32_and9622_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9622_y0);
  and_gate and_gate_h_u_cla32_and9623_y0(h_u_cla32_and9622_y0, h_u_cla32_and9621_y0, h_u_cla32_and9623_y0);
  and_gate and_gate_h_u_cla32_and9624_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9624_y0);
  and_gate and_gate_h_u_cla32_and9625_y0(h_u_cla32_and9624_y0, h_u_cla32_and9623_y0, h_u_cla32_and9625_y0);
  and_gate and_gate_h_u_cla32_and9626_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9626_y0);
  and_gate and_gate_h_u_cla32_and9627_y0(h_u_cla32_and9626_y0, h_u_cla32_and9625_y0, h_u_cla32_and9627_y0);
  and_gate and_gate_h_u_cla32_and9628_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9628_y0);
  and_gate and_gate_h_u_cla32_and9629_y0(h_u_cla32_and9628_y0, h_u_cla32_and9627_y0, h_u_cla32_and9629_y0);
  and_gate and_gate_h_u_cla32_and9630_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and9630_y0);
  and_gate and_gate_h_u_cla32_and9631_y0(h_u_cla32_and9630_y0, h_u_cla32_and9629_y0, h_u_cla32_and9631_y0);
  and_gate and_gate_h_u_cla32_and9632_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9632_y0);
  and_gate and_gate_h_u_cla32_and9633_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9633_y0);
  and_gate and_gate_h_u_cla32_and9634_y0(h_u_cla32_and9633_y0, h_u_cla32_and9632_y0, h_u_cla32_and9634_y0);
  and_gate and_gate_h_u_cla32_and9635_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9635_y0);
  and_gate and_gate_h_u_cla32_and9636_y0(h_u_cla32_and9635_y0, h_u_cla32_and9634_y0, h_u_cla32_and9636_y0);
  and_gate and_gate_h_u_cla32_and9637_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9637_y0);
  and_gate and_gate_h_u_cla32_and9638_y0(h_u_cla32_and9637_y0, h_u_cla32_and9636_y0, h_u_cla32_and9638_y0);
  and_gate and_gate_h_u_cla32_and9639_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9639_y0);
  and_gate and_gate_h_u_cla32_and9640_y0(h_u_cla32_and9639_y0, h_u_cla32_and9638_y0, h_u_cla32_and9640_y0);
  and_gate and_gate_h_u_cla32_and9641_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9641_y0);
  and_gate and_gate_h_u_cla32_and9642_y0(h_u_cla32_and9641_y0, h_u_cla32_and9640_y0, h_u_cla32_and9642_y0);
  and_gate and_gate_h_u_cla32_and9643_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9643_y0);
  and_gate and_gate_h_u_cla32_and9644_y0(h_u_cla32_and9643_y0, h_u_cla32_and9642_y0, h_u_cla32_and9644_y0);
  and_gate and_gate_h_u_cla32_and9645_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9645_y0);
  and_gate and_gate_h_u_cla32_and9646_y0(h_u_cla32_and9645_y0, h_u_cla32_and9644_y0, h_u_cla32_and9646_y0);
  and_gate and_gate_h_u_cla32_and9647_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9647_y0);
  and_gate and_gate_h_u_cla32_and9648_y0(h_u_cla32_and9647_y0, h_u_cla32_and9646_y0, h_u_cla32_and9648_y0);
  and_gate and_gate_h_u_cla32_and9649_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9649_y0);
  and_gate and_gate_h_u_cla32_and9650_y0(h_u_cla32_and9649_y0, h_u_cla32_and9648_y0, h_u_cla32_and9650_y0);
  and_gate and_gate_h_u_cla32_and9651_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9651_y0);
  and_gate and_gate_h_u_cla32_and9652_y0(h_u_cla32_and9651_y0, h_u_cla32_and9650_y0, h_u_cla32_and9652_y0);
  and_gate and_gate_h_u_cla32_and9653_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9653_y0);
  and_gate and_gate_h_u_cla32_and9654_y0(h_u_cla32_and9653_y0, h_u_cla32_and9652_y0, h_u_cla32_and9654_y0);
  and_gate and_gate_h_u_cla32_and9655_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9655_y0);
  and_gate and_gate_h_u_cla32_and9656_y0(h_u_cla32_and9655_y0, h_u_cla32_and9654_y0, h_u_cla32_and9656_y0);
  and_gate and_gate_h_u_cla32_and9657_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9657_y0);
  and_gate and_gate_h_u_cla32_and9658_y0(h_u_cla32_and9657_y0, h_u_cla32_and9656_y0, h_u_cla32_and9658_y0);
  and_gate and_gate_h_u_cla32_and9659_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9659_y0);
  and_gate and_gate_h_u_cla32_and9660_y0(h_u_cla32_and9659_y0, h_u_cla32_and9658_y0, h_u_cla32_and9660_y0);
  and_gate and_gate_h_u_cla32_and9661_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9661_y0);
  and_gate and_gate_h_u_cla32_and9662_y0(h_u_cla32_and9661_y0, h_u_cla32_and9660_y0, h_u_cla32_and9662_y0);
  and_gate and_gate_h_u_cla32_and9663_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9663_y0);
  and_gate and_gate_h_u_cla32_and9664_y0(h_u_cla32_and9663_y0, h_u_cla32_and9662_y0, h_u_cla32_and9664_y0);
  and_gate and_gate_h_u_cla32_and9665_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9665_y0);
  and_gate and_gate_h_u_cla32_and9666_y0(h_u_cla32_and9665_y0, h_u_cla32_and9664_y0, h_u_cla32_and9666_y0);
  and_gate and_gate_h_u_cla32_and9667_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9667_y0);
  and_gate and_gate_h_u_cla32_and9668_y0(h_u_cla32_and9667_y0, h_u_cla32_and9666_y0, h_u_cla32_and9668_y0);
  and_gate and_gate_h_u_cla32_and9669_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9669_y0);
  and_gate and_gate_h_u_cla32_and9670_y0(h_u_cla32_and9669_y0, h_u_cla32_and9668_y0, h_u_cla32_and9670_y0);
  and_gate and_gate_h_u_cla32_and9671_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9671_y0);
  and_gate and_gate_h_u_cla32_and9672_y0(h_u_cla32_and9671_y0, h_u_cla32_and9670_y0, h_u_cla32_and9672_y0);
  and_gate and_gate_h_u_cla32_and9673_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9673_y0);
  and_gate and_gate_h_u_cla32_and9674_y0(h_u_cla32_and9673_y0, h_u_cla32_and9672_y0, h_u_cla32_and9674_y0);
  and_gate and_gate_h_u_cla32_and9675_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9675_y0);
  and_gate and_gate_h_u_cla32_and9676_y0(h_u_cla32_and9675_y0, h_u_cla32_and9674_y0, h_u_cla32_and9676_y0);
  and_gate and_gate_h_u_cla32_and9677_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9677_y0);
  and_gate and_gate_h_u_cla32_and9678_y0(h_u_cla32_and9677_y0, h_u_cla32_and9676_y0, h_u_cla32_and9678_y0);
  and_gate and_gate_h_u_cla32_and9679_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9679_y0);
  and_gate and_gate_h_u_cla32_and9680_y0(h_u_cla32_and9679_y0, h_u_cla32_and9678_y0, h_u_cla32_and9680_y0);
  and_gate and_gate_h_u_cla32_and9681_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9681_y0);
  and_gate and_gate_h_u_cla32_and9682_y0(h_u_cla32_and9681_y0, h_u_cla32_and9680_y0, h_u_cla32_and9682_y0);
  and_gate and_gate_h_u_cla32_and9683_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9683_y0);
  and_gate and_gate_h_u_cla32_and9684_y0(h_u_cla32_and9683_y0, h_u_cla32_and9682_y0, h_u_cla32_and9684_y0);
  and_gate and_gate_h_u_cla32_and9685_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and9685_y0);
  and_gate and_gate_h_u_cla32_and9686_y0(h_u_cla32_and9685_y0, h_u_cla32_and9684_y0, h_u_cla32_and9686_y0);
  and_gate and_gate_h_u_cla32_and9687_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9687_y0);
  and_gate and_gate_h_u_cla32_and9688_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9688_y0);
  and_gate and_gate_h_u_cla32_and9689_y0(h_u_cla32_and9688_y0, h_u_cla32_and9687_y0, h_u_cla32_and9689_y0);
  and_gate and_gate_h_u_cla32_and9690_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9690_y0);
  and_gate and_gate_h_u_cla32_and9691_y0(h_u_cla32_and9690_y0, h_u_cla32_and9689_y0, h_u_cla32_and9691_y0);
  and_gate and_gate_h_u_cla32_and9692_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9692_y0);
  and_gate and_gate_h_u_cla32_and9693_y0(h_u_cla32_and9692_y0, h_u_cla32_and9691_y0, h_u_cla32_and9693_y0);
  and_gate and_gate_h_u_cla32_and9694_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9694_y0);
  and_gate and_gate_h_u_cla32_and9695_y0(h_u_cla32_and9694_y0, h_u_cla32_and9693_y0, h_u_cla32_and9695_y0);
  and_gate and_gate_h_u_cla32_and9696_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9696_y0);
  and_gate and_gate_h_u_cla32_and9697_y0(h_u_cla32_and9696_y0, h_u_cla32_and9695_y0, h_u_cla32_and9697_y0);
  and_gate and_gate_h_u_cla32_and9698_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9698_y0);
  and_gate and_gate_h_u_cla32_and9699_y0(h_u_cla32_and9698_y0, h_u_cla32_and9697_y0, h_u_cla32_and9699_y0);
  and_gate and_gate_h_u_cla32_and9700_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9700_y0);
  and_gate and_gate_h_u_cla32_and9701_y0(h_u_cla32_and9700_y0, h_u_cla32_and9699_y0, h_u_cla32_and9701_y0);
  and_gate and_gate_h_u_cla32_and9702_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9702_y0);
  and_gate and_gate_h_u_cla32_and9703_y0(h_u_cla32_and9702_y0, h_u_cla32_and9701_y0, h_u_cla32_and9703_y0);
  and_gate and_gate_h_u_cla32_and9704_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9704_y0);
  and_gate and_gate_h_u_cla32_and9705_y0(h_u_cla32_and9704_y0, h_u_cla32_and9703_y0, h_u_cla32_and9705_y0);
  and_gate and_gate_h_u_cla32_and9706_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9706_y0);
  and_gate and_gate_h_u_cla32_and9707_y0(h_u_cla32_and9706_y0, h_u_cla32_and9705_y0, h_u_cla32_and9707_y0);
  and_gate and_gate_h_u_cla32_and9708_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9708_y0);
  and_gate and_gate_h_u_cla32_and9709_y0(h_u_cla32_and9708_y0, h_u_cla32_and9707_y0, h_u_cla32_and9709_y0);
  and_gate and_gate_h_u_cla32_and9710_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9710_y0);
  and_gate and_gate_h_u_cla32_and9711_y0(h_u_cla32_and9710_y0, h_u_cla32_and9709_y0, h_u_cla32_and9711_y0);
  and_gate and_gate_h_u_cla32_and9712_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9712_y0);
  and_gate and_gate_h_u_cla32_and9713_y0(h_u_cla32_and9712_y0, h_u_cla32_and9711_y0, h_u_cla32_and9713_y0);
  and_gate and_gate_h_u_cla32_and9714_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9714_y0);
  and_gate and_gate_h_u_cla32_and9715_y0(h_u_cla32_and9714_y0, h_u_cla32_and9713_y0, h_u_cla32_and9715_y0);
  and_gate and_gate_h_u_cla32_and9716_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9716_y0);
  and_gate and_gate_h_u_cla32_and9717_y0(h_u_cla32_and9716_y0, h_u_cla32_and9715_y0, h_u_cla32_and9717_y0);
  and_gate and_gate_h_u_cla32_and9718_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9718_y0);
  and_gate and_gate_h_u_cla32_and9719_y0(h_u_cla32_and9718_y0, h_u_cla32_and9717_y0, h_u_cla32_and9719_y0);
  and_gate and_gate_h_u_cla32_and9720_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9720_y0);
  and_gate and_gate_h_u_cla32_and9721_y0(h_u_cla32_and9720_y0, h_u_cla32_and9719_y0, h_u_cla32_and9721_y0);
  and_gate and_gate_h_u_cla32_and9722_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9722_y0);
  and_gate and_gate_h_u_cla32_and9723_y0(h_u_cla32_and9722_y0, h_u_cla32_and9721_y0, h_u_cla32_and9723_y0);
  and_gate and_gate_h_u_cla32_and9724_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9724_y0);
  and_gate and_gate_h_u_cla32_and9725_y0(h_u_cla32_and9724_y0, h_u_cla32_and9723_y0, h_u_cla32_and9725_y0);
  and_gate and_gate_h_u_cla32_and9726_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9726_y0);
  and_gate and_gate_h_u_cla32_and9727_y0(h_u_cla32_and9726_y0, h_u_cla32_and9725_y0, h_u_cla32_and9727_y0);
  and_gate and_gate_h_u_cla32_and9728_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9728_y0);
  and_gate and_gate_h_u_cla32_and9729_y0(h_u_cla32_and9728_y0, h_u_cla32_and9727_y0, h_u_cla32_and9729_y0);
  and_gate and_gate_h_u_cla32_and9730_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9730_y0);
  and_gate and_gate_h_u_cla32_and9731_y0(h_u_cla32_and9730_y0, h_u_cla32_and9729_y0, h_u_cla32_and9731_y0);
  and_gate and_gate_h_u_cla32_and9732_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9732_y0);
  and_gate and_gate_h_u_cla32_and9733_y0(h_u_cla32_and9732_y0, h_u_cla32_and9731_y0, h_u_cla32_and9733_y0);
  and_gate and_gate_h_u_cla32_and9734_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9734_y0);
  and_gate and_gate_h_u_cla32_and9735_y0(h_u_cla32_and9734_y0, h_u_cla32_and9733_y0, h_u_cla32_and9735_y0);
  and_gate and_gate_h_u_cla32_and9736_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9736_y0);
  and_gate and_gate_h_u_cla32_and9737_y0(h_u_cla32_and9736_y0, h_u_cla32_and9735_y0, h_u_cla32_and9737_y0);
  and_gate and_gate_h_u_cla32_and9738_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and9738_y0);
  and_gate and_gate_h_u_cla32_and9739_y0(h_u_cla32_and9738_y0, h_u_cla32_and9737_y0, h_u_cla32_and9739_y0);
  and_gate and_gate_h_u_cla32_and9740_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9740_y0);
  and_gate and_gate_h_u_cla32_and9741_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9741_y0);
  and_gate and_gate_h_u_cla32_and9742_y0(h_u_cla32_and9741_y0, h_u_cla32_and9740_y0, h_u_cla32_and9742_y0);
  and_gate and_gate_h_u_cla32_and9743_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9743_y0);
  and_gate and_gate_h_u_cla32_and9744_y0(h_u_cla32_and9743_y0, h_u_cla32_and9742_y0, h_u_cla32_and9744_y0);
  and_gate and_gate_h_u_cla32_and9745_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9745_y0);
  and_gate and_gate_h_u_cla32_and9746_y0(h_u_cla32_and9745_y0, h_u_cla32_and9744_y0, h_u_cla32_and9746_y0);
  and_gate and_gate_h_u_cla32_and9747_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9747_y0);
  and_gate and_gate_h_u_cla32_and9748_y0(h_u_cla32_and9747_y0, h_u_cla32_and9746_y0, h_u_cla32_and9748_y0);
  and_gate and_gate_h_u_cla32_and9749_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9749_y0);
  and_gate and_gate_h_u_cla32_and9750_y0(h_u_cla32_and9749_y0, h_u_cla32_and9748_y0, h_u_cla32_and9750_y0);
  and_gate and_gate_h_u_cla32_and9751_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9751_y0);
  and_gate and_gate_h_u_cla32_and9752_y0(h_u_cla32_and9751_y0, h_u_cla32_and9750_y0, h_u_cla32_and9752_y0);
  and_gate and_gate_h_u_cla32_and9753_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9753_y0);
  and_gate and_gate_h_u_cla32_and9754_y0(h_u_cla32_and9753_y0, h_u_cla32_and9752_y0, h_u_cla32_and9754_y0);
  and_gate and_gate_h_u_cla32_and9755_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9755_y0);
  and_gate and_gate_h_u_cla32_and9756_y0(h_u_cla32_and9755_y0, h_u_cla32_and9754_y0, h_u_cla32_and9756_y0);
  and_gate and_gate_h_u_cla32_and9757_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9757_y0);
  and_gate and_gate_h_u_cla32_and9758_y0(h_u_cla32_and9757_y0, h_u_cla32_and9756_y0, h_u_cla32_and9758_y0);
  and_gate and_gate_h_u_cla32_and9759_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9759_y0);
  and_gate and_gate_h_u_cla32_and9760_y0(h_u_cla32_and9759_y0, h_u_cla32_and9758_y0, h_u_cla32_and9760_y0);
  and_gate and_gate_h_u_cla32_and9761_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9761_y0);
  and_gate and_gate_h_u_cla32_and9762_y0(h_u_cla32_and9761_y0, h_u_cla32_and9760_y0, h_u_cla32_and9762_y0);
  and_gate and_gate_h_u_cla32_and9763_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9763_y0);
  and_gate and_gate_h_u_cla32_and9764_y0(h_u_cla32_and9763_y0, h_u_cla32_and9762_y0, h_u_cla32_and9764_y0);
  and_gate and_gate_h_u_cla32_and9765_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9765_y0);
  and_gate and_gate_h_u_cla32_and9766_y0(h_u_cla32_and9765_y0, h_u_cla32_and9764_y0, h_u_cla32_and9766_y0);
  and_gate and_gate_h_u_cla32_and9767_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9767_y0);
  and_gate and_gate_h_u_cla32_and9768_y0(h_u_cla32_and9767_y0, h_u_cla32_and9766_y0, h_u_cla32_and9768_y0);
  and_gate and_gate_h_u_cla32_and9769_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9769_y0);
  and_gate and_gate_h_u_cla32_and9770_y0(h_u_cla32_and9769_y0, h_u_cla32_and9768_y0, h_u_cla32_and9770_y0);
  and_gate and_gate_h_u_cla32_and9771_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9771_y0);
  and_gate and_gate_h_u_cla32_and9772_y0(h_u_cla32_and9771_y0, h_u_cla32_and9770_y0, h_u_cla32_and9772_y0);
  and_gate and_gate_h_u_cla32_and9773_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9773_y0);
  and_gate and_gate_h_u_cla32_and9774_y0(h_u_cla32_and9773_y0, h_u_cla32_and9772_y0, h_u_cla32_and9774_y0);
  and_gate and_gate_h_u_cla32_and9775_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9775_y0);
  and_gate and_gate_h_u_cla32_and9776_y0(h_u_cla32_and9775_y0, h_u_cla32_and9774_y0, h_u_cla32_and9776_y0);
  and_gate and_gate_h_u_cla32_and9777_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9777_y0);
  and_gate and_gate_h_u_cla32_and9778_y0(h_u_cla32_and9777_y0, h_u_cla32_and9776_y0, h_u_cla32_and9778_y0);
  and_gate and_gate_h_u_cla32_and9779_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9779_y0);
  and_gate and_gate_h_u_cla32_and9780_y0(h_u_cla32_and9779_y0, h_u_cla32_and9778_y0, h_u_cla32_and9780_y0);
  and_gate and_gate_h_u_cla32_and9781_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9781_y0);
  and_gate and_gate_h_u_cla32_and9782_y0(h_u_cla32_and9781_y0, h_u_cla32_and9780_y0, h_u_cla32_and9782_y0);
  and_gate and_gate_h_u_cla32_and9783_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9783_y0);
  and_gate and_gate_h_u_cla32_and9784_y0(h_u_cla32_and9783_y0, h_u_cla32_and9782_y0, h_u_cla32_and9784_y0);
  and_gate and_gate_h_u_cla32_and9785_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9785_y0);
  and_gate and_gate_h_u_cla32_and9786_y0(h_u_cla32_and9785_y0, h_u_cla32_and9784_y0, h_u_cla32_and9786_y0);
  and_gate and_gate_h_u_cla32_and9787_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9787_y0);
  and_gate and_gate_h_u_cla32_and9788_y0(h_u_cla32_and9787_y0, h_u_cla32_and9786_y0, h_u_cla32_and9788_y0);
  and_gate and_gate_h_u_cla32_and9789_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and9789_y0);
  and_gate and_gate_h_u_cla32_and9790_y0(h_u_cla32_and9789_y0, h_u_cla32_and9788_y0, h_u_cla32_and9790_y0);
  and_gate and_gate_h_u_cla32_and9791_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9791_y0);
  and_gate and_gate_h_u_cla32_and9792_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9792_y0);
  and_gate and_gate_h_u_cla32_and9793_y0(h_u_cla32_and9792_y0, h_u_cla32_and9791_y0, h_u_cla32_and9793_y0);
  and_gate and_gate_h_u_cla32_and9794_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9794_y0);
  and_gate and_gate_h_u_cla32_and9795_y0(h_u_cla32_and9794_y0, h_u_cla32_and9793_y0, h_u_cla32_and9795_y0);
  and_gate and_gate_h_u_cla32_and9796_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9796_y0);
  and_gate and_gate_h_u_cla32_and9797_y0(h_u_cla32_and9796_y0, h_u_cla32_and9795_y0, h_u_cla32_and9797_y0);
  and_gate and_gate_h_u_cla32_and9798_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9798_y0);
  and_gate and_gate_h_u_cla32_and9799_y0(h_u_cla32_and9798_y0, h_u_cla32_and9797_y0, h_u_cla32_and9799_y0);
  and_gate and_gate_h_u_cla32_and9800_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9800_y0);
  and_gate and_gate_h_u_cla32_and9801_y0(h_u_cla32_and9800_y0, h_u_cla32_and9799_y0, h_u_cla32_and9801_y0);
  and_gate and_gate_h_u_cla32_and9802_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9802_y0);
  and_gate and_gate_h_u_cla32_and9803_y0(h_u_cla32_and9802_y0, h_u_cla32_and9801_y0, h_u_cla32_and9803_y0);
  and_gate and_gate_h_u_cla32_and9804_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9804_y0);
  and_gate and_gate_h_u_cla32_and9805_y0(h_u_cla32_and9804_y0, h_u_cla32_and9803_y0, h_u_cla32_and9805_y0);
  and_gate and_gate_h_u_cla32_and9806_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9806_y0);
  and_gate and_gate_h_u_cla32_and9807_y0(h_u_cla32_and9806_y0, h_u_cla32_and9805_y0, h_u_cla32_and9807_y0);
  and_gate and_gate_h_u_cla32_and9808_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9808_y0);
  and_gate and_gate_h_u_cla32_and9809_y0(h_u_cla32_and9808_y0, h_u_cla32_and9807_y0, h_u_cla32_and9809_y0);
  and_gate and_gate_h_u_cla32_and9810_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9810_y0);
  and_gate and_gate_h_u_cla32_and9811_y0(h_u_cla32_and9810_y0, h_u_cla32_and9809_y0, h_u_cla32_and9811_y0);
  and_gate and_gate_h_u_cla32_and9812_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9812_y0);
  and_gate and_gate_h_u_cla32_and9813_y0(h_u_cla32_and9812_y0, h_u_cla32_and9811_y0, h_u_cla32_and9813_y0);
  and_gate and_gate_h_u_cla32_and9814_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9814_y0);
  and_gate and_gate_h_u_cla32_and9815_y0(h_u_cla32_and9814_y0, h_u_cla32_and9813_y0, h_u_cla32_and9815_y0);
  and_gate and_gate_h_u_cla32_and9816_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9816_y0);
  and_gate and_gate_h_u_cla32_and9817_y0(h_u_cla32_and9816_y0, h_u_cla32_and9815_y0, h_u_cla32_and9817_y0);
  and_gate and_gate_h_u_cla32_and9818_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9818_y0);
  and_gate and_gate_h_u_cla32_and9819_y0(h_u_cla32_and9818_y0, h_u_cla32_and9817_y0, h_u_cla32_and9819_y0);
  and_gate and_gate_h_u_cla32_and9820_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9820_y0);
  and_gate and_gate_h_u_cla32_and9821_y0(h_u_cla32_and9820_y0, h_u_cla32_and9819_y0, h_u_cla32_and9821_y0);
  and_gate and_gate_h_u_cla32_and9822_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9822_y0);
  and_gate and_gate_h_u_cla32_and9823_y0(h_u_cla32_and9822_y0, h_u_cla32_and9821_y0, h_u_cla32_and9823_y0);
  and_gate and_gate_h_u_cla32_and9824_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9824_y0);
  and_gate and_gate_h_u_cla32_and9825_y0(h_u_cla32_and9824_y0, h_u_cla32_and9823_y0, h_u_cla32_and9825_y0);
  and_gate and_gate_h_u_cla32_and9826_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9826_y0);
  and_gate and_gate_h_u_cla32_and9827_y0(h_u_cla32_and9826_y0, h_u_cla32_and9825_y0, h_u_cla32_and9827_y0);
  and_gate and_gate_h_u_cla32_and9828_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9828_y0);
  and_gate and_gate_h_u_cla32_and9829_y0(h_u_cla32_and9828_y0, h_u_cla32_and9827_y0, h_u_cla32_and9829_y0);
  and_gate and_gate_h_u_cla32_and9830_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9830_y0);
  and_gate and_gate_h_u_cla32_and9831_y0(h_u_cla32_and9830_y0, h_u_cla32_and9829_y0, h_u_cla32_and9831_y0);
  and_gate and_gate_h_u_cla32_and9832_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9832_y0);
  and_gate and_gate_h_u_cla32_and9833_y0(h_u_cla32_and9832_y0, h_u_cla32_and9831_y0, h_u_cla32_and9833_y0);
  and_gate and_gate_h_u_cla32_and9834_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9834_y0);
  and_gate and_gate_h_u_cla32_and9835_y0(h_u_cla32_and9834_y0, h_u_cla32_and9833_y0, h_u_cla32_and9835_y0);
  and_gate and_gate_h_u_cla32_and9836_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9836_y0);
  and_gate and_gate_h_u_cla32_and9837_y0(h_u_cla32_and9836_y0, h_u_cla32_and9835_y0, h_u_cla32_and9837_y0);
  and_gate and_gate_h_u_cla32_and9838_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and9838_y0);
  and_gate and_gate_h_u_cla32_and9839_y0(h_u_cla32_and9838_y0, h_u_cla32_and9837_y0, h_u_cla32_and9839_y0);
  and_gate and_gate_h_u_cla32_and9840_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9840_y0);
  and_gate and_gate_h_u_cla32_and9841_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9841_y0);
  and_gate and_gate_h_u_cla32_and9842_y0(h_u_cla32_and9841_y0, h_u_cla32_and9840_y0, h_u_cla32_and9842_y0);
  and_gate and_gate_h_u_cla32_and9843_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9843_y0);
  and_gate and_gate_h_u_cla32_and9844_y0(h_u_cla32_and9843_y0, h_u_cla32_and9842_y0, h_u_cla32_and9844_y0);
  and_gate and_gate_h_u_cla32_and9845_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9845_y0);
  and_gate and_gate_h_u_cla32_and9846_y0(h_u_cla32_and9845_y0, h_u_cla32_and9844_y0, h_u_cla32_and9846_y0);
  and_gate and_gate_h_u_cla32_and9847_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9847_y0);
  and_gate and_gate_h_u_cla32_and9848_y0(h_u_cla32_and9847_y0, h_u_cla32_and9846_y0, h_u_cla32_and9848_y0);
  and_gate and_gate_h_u_cla32_and9849_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9849_y0);
  and_gate and_gate_h_u_cla32_and9850_y0(h_u_cla32_and9849_y0, h_u_cla32_and9848_y0, h_u_cla32_and9850_y0);
  and_gate and_gate_h_u_cla32_and9851_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9851_y0);
  and_gate and_gate_h_u_cla32_and9852_y0(h_u_cla32_and9851_y0, h_u_cla32_and9850_y0, h_u_cla32_and9852_y0);
  and_gate and_gate_h_u_cla32_and9853_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9853_y0);
  and_gate and_gate_h_u_cla32_and9854_y0(h_u_cla32_and9853_y0, h_u_cla32_and9852_y0, h_u_cla32_and9854_y0);
  and_gate and_gate_h_u_cla32_and9855_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9855_y0);
  and_gate and_gate_h_u_cla32_and9856_y0(h_u_cla32_and9855_y0, h_u_cla32_and9854_y0, h_u_cla32_and9856_y0);
  and_gate and_gate_h_u_cla32_and9857_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9857_y0);
  and_gate and_gate_h_u_cla32_and9858_y0(h_u_cla32_and9857_y0, h_u_cla32_and9856_y0, h_u_cla32_and9858_y0);
  and_gate and_gate_h_u_cla32_and9859_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9859_y0);
  and_gate and_gate_h_u_cla32_and9860_y0(h_u_cla32_and9859_y0, h_u_cla32_and9858_y0, h_u_cla32_and9860_y0);
  and_gate and_gate_h_u_cla32_and9861_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9861_y0);
  and_gate and_gate_h_u_cla32_and9862_y0(h_u_cla32_and9861_y0, h_u_cla32_and9860_y0, h_u_cla32_and9862_y0);
  and_gate and_gate_h_u_cla32_and9863_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9863_y0);
  and_gate and_gate_h_u_cla32_and9864_y0(h_u_cla32_and9863_y0, h_u_cla32_and9862_y0, h_u_cla32_and9864_y0);
  and_gate and_gate_h_u_cla32_and9865_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9865_y0);
  and_gate and_gate_h_u_cla32_and9866_y0(h_u_cla32_and9865_y0, h_u_cla32_and9864_y0, h_u_cla32_and9866_y0);
  and_gate and_gate_h_u_cla32_and9867_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9867_y0);
  and_gate and_gate_h_u_cla32_and9868_y0(h_u_cla32_and9867_y0, h_u_cla32_and9866_y0, h_u_cla32_and9868_y0);
  and_gate and_gate_h_u_cla32_and9869_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9869_y0);
  and_gate and_gate_h_u_cla32_and9870_y0(h_u_cla32_and9869_y0, h_u_cla32_and9868_y0, h_u_cla32_and9870_y0);
  and_gate and_gate_h_u_cla32_and9871_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9871_y0);
  and_gate and_gate_h_u_cla32_and9872_y0(h_u_cla32_and9871_y0, h_u_cla32_and9870_y0, h_u_cla32_and9872_y0);
  and_gate and_gate_h_u_cla32_and9873_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9873_y0);
  and_gate and_gate_h_u_cla32_and9874_y0(h_u_cla32_and9873_y0, h_u_cla32_and9872_y0, h_u_cla32_and9874_y0);
  and_gate and_gate_h_u_cla32_and9875_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9875_y0);
  and_gate and_gate_h_u_cla32_and9876_y0(h_u_cla32_and9875_y0, h_u_cla32_and9874_y0, h_u_cla32_and9876_y0);
  and_gate and_gate_h_u_cla32_and9877_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9877_y0);
  and_gate and_gate_h_u_cla32_and9878_y0(h_u_cla32_and9877_y0, h_u_cla32_and9876_y0, h_u_cla32_and9878_y0);
  and_gate and_gate_h_u_cla32_and9879_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9879_y0);
  and_gate and_gate_h_u_cla32_and9880_y0(h_u_cla32_and9879_y0, h_u_cla32_and9878_y0, h_u_cla32_and9880_y0);
  and_gate and_gate_h_u_cla32_and9881_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9881_y0);
  and_gate and_gate_h_u_cla32_and9882_y0(h_u_cla32_and9881_y0, h_u_cla32_and9880_y0, h_u_cla32_and9882_y0);
  and_gate and_gate_h_u_cla32_and9883_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9883_y0);
  and_gate and_gate_h_u_cla32_and9884_y0(h_u_cla32_and9883_y0, h_u_cla32_and9882_y0, h_u_cla32_and9884_y0);
  and_gate and_gate_h_u_cla32_and9885_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and9885_y0);
  and_gate and_gate_h_u_cla32_and9886_y0(h_u_cla32_and9885_y0, h_u_cla32_and9884_y0, h_u_cla32_and9886_y0);
  and_gate and_gate_h_u_cla32_and9887_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9887_y0);
  and_gate and_gate_h_u_cla32_and9888_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9888_y0);
  and_gate and_gate_h_u_cla32_and9889_y0(h_u_cla32_and9888_y0, h_u_cla32_and9887_y0, h_u_cla32_and9889_y0);
  and_gate and_gate_h_u_cla32_and9890_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9890_y0);
  and_gate and_gate_h_u_cla32_and9891_y0(h_u_cla32_and9890_y0, h_u_cla32_and9889_y0, h_u_cla32_and9891_y0);
  and_gate and_gate_h_u_cla32_and9892_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9892_y0);
  and_gate and_gate_h_u_cla32_and9893_y0(h_u_cla32_and9892_y0, h_u_cla32_and9891_y0, h_u_cla32_and9893_y0);
  and_gate and_gate_h_u_cla32_and9894_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9894_y0);
  and_gate and_gate_h_u_cla32_and9895_y0(h_u_cla32_and9894_y0, h_u_cla32_and9893_y0, h_u_cla32_and9895_y0);
  and_gate and_gate_h_u_cla32_and9896_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9896_y0);
  and_gate and_gate_h_u_cla32_and9897_y0(h_u_cla32_and9896_y0, h_u_cla32_and9895_y0, h_u_cla32_and9897_y0);
  and_gate and_gate_h_u_cla32_and9898_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9898_y0);
  and_gate and_gate_h_u_cla32_and9899_y0(h_u_cla32_and9898_y0, h_u_cla32_and9897_y0, h_u_cla32_and9899_y0);
  and_gate and_gate_h_u_cla32_and9900_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9900_y0);
  and_gate and_gate_h_u_cla32_and9901_y0(h_u_cla32_and9900_y0, h_u_cla32_and9899_y0, h_u_cla32_and9901_y0);
  and_gate and_gate_h_u_cla32_and9902_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9902_y0);
  and_gate and_gate_h_u_cla32_and9903_y0(h_u_cla32_and9902_y0, h_u_cla32_and9901_y0, h_u_cla32_and9903_y0);
  and_gate and_gate_h_u_cla32_and9904_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9904_y0);
  and_gate and_gate_h_u_cla32_and9905_y0(h_u_cla32_and9904_y0, h_u_cla32_and9903_y0, h_u_cla32_and9905_y0);
  and_gate and_gate_h_u_cla32_and9906_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9906_y0);
  and_gate and_gate_h_u_cla32_and9907_y0(h_u_cla32_and9906_y0, h_u_cla32_and9905_y0, h_u_cla32_and9907_y0);
  and_gate and_gate_h_u_cla32_and9908_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9908_y0);
  and_gate and_gate_h_u_cla32_and9909_y0(h_u_cla32_and9908_y0, h_u_cla32_and9907_y0, h_u_cla32_and9909_y0);
  and_gate and_gate_h_u_cla32_and9910_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9910_y0);
  and_gate and_gate_h_u_cla32_and9911_y0(h_u_cla32_and9910_y0, h_u_cla32_and9909_y0, h_u_cla32_and9911_y0);
  and_gate and_gate_h_u_cla32_and9912_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9912_y0);
  and_gate and_gate_h_u_cla32_and9913_y0(h_u_cla32_and9912_y0, h_u_cla32_and9911_y0, h_u_cla32_and9913_y0);
  and_gate and_gate_h_u_cla32_and9914_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9914_y0);
  and_gate and_gate_h_u_cla32_and9915_y0(h_u_cla32_and9914_y0, h_u_cla32_and9913_y0, h_u_cla32_and9915_y0);
  and_gate and_gate_h_u_cla32_and9916_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9916_y0);
  and_gate and_gate_h_u_cla32_and9917_y0(h_u_cla32_and9916_y0, h_u_cla32_and9915_y0, h_u_cla32_and9917_y0);
  and_gate and_gate_h_u_cla32_and9918_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9918_y0);
  and_gate and_gate_h_u_cla32_and9919_y0(h_u_cla32_and9918_y0, h_u_cla32_and9917_y0, h_u_cla32_and9919_y0);
  and_gate and_gate_h_u_cla32_and9920_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9920_y0);
  and_gate and_gate_h_u_cla32_and9921_y0(h_u_cla32_and9920_y0, h_u_cla32_and9919_y0, h_u_cla32_and9921_y0);
  and_gate and_gate_h_u_cla32_and9922_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9922_y0);
  and_gate and_gate_h_u_cla32_and9923_y0(h_u_cla32_and9922_y0, h_u_cla32_and9921_y0, h_u_cla32_and9923_y0);
  and_gate and_gate_h_u_cla32_and9924_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9924_y0);
  and_gate and_gate_h_u_cla32_and9925_y0(h_u_cla32_and9924_y0, h_u_cla32_and9923_y0, h_u_cla32_and9925_y0);
  and_gate and_gate_h_u_cla32_and9926_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9926_y0);
  and_gate and_gate_h_u_cla32_and9927_y0(h_u_cla32_and9926_y0, h_u_cla32_and9925_y0, h_u_cla32_and9927_y0);
  and_gate and_gate_h_u_cla32_and9928_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9928_y0);
  and_gate and_gate_h_u_cla32_and9929_y0(h_u_cla32_and9928_y0, h_u_cla32_and9927_y0, h_u_cla32_and9929_y0);
  and_gate and_gate_h_u_cla32_and9930_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and9930_y0);
  and_gate and_gate_h_u_cla32_and9931_y0(h_u_cla32_and9930_y0, h_u_cla32_and9929_y0, h_u_cla32_and9931_y0);
  and_gate and_gate_h_u_cla32_and9932_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9932_y0);
  and_gate and_gate_h_u_cla32_and9933_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9933_y0);
  and_gate and_gate_h_u_cla32_and9934_y0(h_u_cla32_and9933_y0, h_u_cla32_and9932_y0, h_u_cla32_and9934_y0);
  and_gate and_gate_h_u_cla32_and9935_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9935_y0);
  and_gate and_gate_h_u_cla32_and9936_y0(h_u_cla32_and9935_y0, h_u_cla32_and9934_y0, h_u_cla32_and9936_y0);
  and_gate and_gate_h_u_cla32_and9937_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9937_y0);
  and_gate and_gate_h_u_cla32_and9938_y0(h_u_cla32_and9937_y0, h_u_cla32_and9936_y0, h_u_cla32_and9938_y0);
  and_gate and_gate_h_u_cla32_and9939_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9939_y0);
  and_gate and_gate_h_u_cla32_and9940_y0(h_u_cla32_and9939_y0, h_u_cla32_and9938_y0, h_u_cla32_and9940_y0);
  and_gate and_gate_h_u_cla32_and9941_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9941_y0);
  and_gate and_gate_h_u_cla32_and9942_y0(h_u_cla32_and9941_y0, h_u_cla32_and9940_y0, h_u_cla32_and9942_y0);
  and_gate and_gate_h_u_cla32_and9943_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9943_y0);
  and_gate and_gate_h_u_cla32_and9944_y0(h_u_cla32_and9943_y0, h_u_cla32_and9942_y0, h_u_cla32_and9944_y0);
  and_gate and_gate_h_u_cla32_and9945_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9945_y0);
  and_gate and_gate_h_u_cla32_and9946_y0(h_u_cla32_and9945_y0, h_u_cla32_and9944_y0, h_u_cla32_and9946_y0);
  and_gate and_gate_h_u_cla32_and9947_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9947_y0);
  and_gate and_gate_h_u_cla32_and9948_y0(h_u_cla32_and9947_y0, h_u_cla32_and9946_y0, h_u_cla32_and9948_y0);
  and_gate and_gate_h_u_cla32_and9949_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9949_y0);
  and_gate and_gate_h_u_cla32_and9950_y0(h_u_cla32_and9949_y0, h_u_cla32_and9948_y0, h_u_cla32_and9950_y0);
  and_gate and_gate_h_u_cla32_and9951_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9951_y0);
  and_gate and_gate_h_u_cla32_and9952_y0(h_u_cla32_and9951_y0, h_u_cla32_and9950_y0, h_u_cla32_and9952_y0);
  and_gate and_gate_h_u_cla32_and9953_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9953_y0);
  and_gate and_gate_h_u_cla32_and9954_y0(h_u_cla32_and9953_y0, h_u_cla32_and9952_y0, h_u_cla32_and9954_y0);
  and_gate and_gate_h_u_cla32_and9955_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9955_y0);
  and_gate and_gate_h_u_cla32_and9956_y0(h_u_cla32_and9955_y0, h_u_cla32_and9954_y0, h_u_cla32_and9956_y0);
  and_gate and_gate_h_u_cla32_and9957_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9957_y0);
  and_gate and_gate_h_u_cla32_and9958_y0(h_u_cla32_and9957_y0, h_u_cla32_and9956_y0, h_u_cla32_and9958_y0);
  and_gate and_gate_h_u_cla32_and9959_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9959_y0);
  and_gate and_gate_h_u_cla32_and9960_y0(h_u_cla32_and9959_y0, h_u_cla32_and9958_y0, h_u_cla32_and9960_y0);
  and_gate and_gate_h_u_cla32_and9961_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9961_y0);
  and_gate and_gate_h_u_cla32_and9962_y0(h_u_cla32_and9961_y0, h_u_cla32_and9960_y0, h_u_cla32_and9962_y0);
  and_gate and_gate_h_u_cla32_and9963_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9963_y0);
  and_gate and_gate_h_u_cla32_and9964_y0(h_u_cla32_and9963_y0, h_u_cla32_and9962_y0, h_u_cla32_and9964_y0);
  and_gate and_gate_h_u_cla32_and9965_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9965_y0);
  and_gate and_gate_h_u_cla32_and9966_y0(h_u_cla32_and9965_y0, h_u_cla32_and9964_y0, h_u_cla32_and9966_y0);
  and_gate and_gate_h_u_cla32_and9967_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9967_y0);
  and_gate and_gate_h_u_cla32_and9968_y0(h_u_cla32_and9967_y0, h_u_cla32_and9966_y0, h_u_cla32_and9968_y0);
  and_gate and_gate_h_u_cla32_and9969_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9969_y0);
  and_gate and_gate_h_u_cla32_and9970_y0(h_u_cla32_and9969_y0, h_u_cla32_and9968_y0, h_u_cla32_and9970_y0);
  and_gate and_gate_h_u_cla32_and9971_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9971_y0);
  and_gate and_gate_h_u_cla32_and9972_y0(h_u_cla32_and9971_y0, h_u_cla32_and9970_y0, h_u_cla32_and9972_y0);
  and_gate and_gate_h_u_cla32_and9973_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and9973_y0);
  and_gate and_gate_h_u_cla32_and9974_y0(h_u_cla32_and9973_y0, h_u_cla32_and9972_y0, h_u_cla32_and9974_y0);
  and_gate and_gate_h_u_cla32_and9975_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9975_y0);
  and_gate and_gate_h_u_cla32_and9976_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9976_y0);
  and_gate and_gate_h_u_cla32_and9977_y0(h_u_cla32_and9976_y0, h_u_cla32_and9975_y0, h_u_cla32_and9977_y0);
  and_gate and_gate_h_u_cla32_and9978_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9978_y0);
  and_gate and_gate_h_u_cla32_and9979_y0(h_u_cla32_and9978_y0, h_u_cla32_and9977_y0, h_u_cla32_and9979_y0);
  and_gate and_gate_h_u_cla32_and9980_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9980_y0);
  and_gate and_gate_h_u_cla32_and9981_y0(h_u_cla32_and9980_y0, h_u_cla32_and9979_y0, h_u_cla32_and9981_y0);
  and_gate and_gate_h_u_cla32_and9982_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9982_y0);
  and_gate and_gate_h_u_cla32_and9983_y0(h_u_cla32_and9982_y0, h_u_cla32_and9981_y0, h_u_cla32_and9983_y0);
  and_gate and_gate_h_u_cla32_and9984_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9984_y0);
  and_gate and_gate_h_u_cla32_and9985_y0(h_u_cla32_and9984_y0, h_u_cla32_and9983_y0, h_u_cla32_and9985_y0);
  and_gate and_gate_h_u_cla32_and9986_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9986_y0);
  and_gate and_gate_h_u_cla32_and9987_y0(h_u_cla32_and9986_y0, h_u_cla32_and9985_y0, h_u_cla32_and9987_y0);
  and_gate and_gate_h_u_cla32_and9988_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9988_y0);
  and_gate and_gate_h_u_cla32_and9989_y0(h_u_cla32_and9988_y0, h_u_cla32_and9987_y0, h_u_cla32_and9989_y0);
  and_gate and_gate_h_u_cla32_and9990_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9990_y0);
  and_gate and_gate_h_u_cla32_and9991_y0(h_u_cla32_and9990_y0, h_u_cla32_and9989_y0, h_u_cla32_and9991_y0);
  and_gate and_gate_h_u_cla32_and9992_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9992_y0);
  and_gate and_gate_h_u_cla32_and9993_y0(h_u_cla32_and9992_y0, h_u_cla32_and9991_y0, h_u_cla32_and9993_y0);
  and_gate and_gate_h_u_cla32_and9994_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9994_y0);
  and_gate and_gate_h_u_cla32_and9995_y0(h_u_cla32_and9994_y0, h_u_cla32_and9993_y0, h_u_cla32_and9995_y0);
  and_gate and_gate_h_u_cla32_and9996_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9996_y0);
  and_gate and_gate_h_u_cla32_and9997_y0(h_u_cla32_and9996_y0, h_u_cla32_and9995_y0, h_u_cla32_and9997_y0);
  and_gate and_gate_h_u_cla32_and9998_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and9998_y0);
  and_gate and_gate_h_u_cla32_and9999_y0(h_u_cla32_and9998_y0, h_u_cla32_and9997_y0, h_u_cla32_and9999_y0);
  and_gate and_gate_h_u_cla32_and10000_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10000_y0);
  and_gate and_gate_h_u_cla32_and10001_y0(h_u_cla32_and10000_y0, h_u_cla32_and9999_y0, h_u_cla32_and10001_y0);
  and_gate and_gate_h_u_cla32_and10002_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10002_y0);
  and_gate and_gate_h_u_cla32_and10003_y0(h_u_cla32_and10002_y0, h_u_cla32_and10001_y0, h_u_cla32_and10003_y0);
  and_gate and_gate_h_u_cla32_and10004_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10004_y0);
  and_gate and_gate_h_u_cla32_and10005_y0(h_u_cla32_and10004_y0, h_u_cla32_and10003_y0, h_u_cla32_and10005_y0);
  and_gate and_gate_h_u_cla32_and10006_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10006_y0);
  and_gate and_gate_h_u_cla32_and10007_y0(h_u_cla32_and10006_y0, h_u_cla32_and10005_y0, h_u_cla32_and10007_y0);
  and_gate and_gate_h_u_cla32_and10008_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10008_y0);
  and_gate and_gate_h_u_cla32_and10009_y0(h_u_cla32_and10008_y0, h_u_cla32_and10007_y0, h_u_cla32_and10009_y0);
  and_gate and_gate_h_u_cla32_and10010_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10010_y0);
  and_gate and_gate_h_u_cla32_and10011_y0(h_u_cla32_and10010_y0, h_u_cla32_and10009_y0, h_u_cla32_and10011_y0);
  and_gate and_gate_h_u_cla32_and10012_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10012_y0);
  and_gate and_gate_h_u_cla32_and10013_y0(h_u_cla32_and10012_y0, h_u_cla32_and10011_y0, h_u_cla32_and10013_y0);
  and_gate and_gate_h_u_cla32_and10014_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10014_y0);
  and_gate and_gate_h_u_cla32_and10015_y0(h_u_cla32_and10014_y0, h_u_cla32_and10013_y0, h_u_cla32_and10015_y0);
  and_gate and_gate_h_u_cla32_and10016_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10016_y0);
  and_gate and_gate_h_u_cla32_and10017_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10017_y0);
  and_gate and_gate_h_u_cla32_and10018_y0(h_u_cla32_and10017_y0, h_u_cla32_and10016_y0, h_u_cla32_and10018_y0);
  and_gate and_gate_h_u_cla32_and10019_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10019_y0);
  and_gate and_gate_h_u_cla32_and10020_y0(h_u_cla32_and10019_y0, h_u_cla32_and10018_y0, h_u_cla32_and10020_y0);
  and_gate and_gate_h_u_cla32_and10021_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10021_y0);
  and_gate and_gate_h_u_cla32_and10022_y0(h_u_cla32_and10021_y0, h_u_cla32_and10020_y0, h_u_cla32_and10022_y0);
  and_gate and_gate_h_u_cla32_and10023_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10023_y0);
  and_gate and_gate_h_u_cla32_and10024_y0(h_u_cla32_and10023_y0, h_u_cla32_and10022_y0, h_u_cla32_and10024_y0);
  and_gate and_gate_h_u_cla32_and10025_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10025_y0);
  and_gate and_gate_h_u_cla32_and10026_y0(h_u_cla32_and10025_y0, h_u_cla32_and10024_y0, h_u_cla32_and10026_y0);
  and_gate and_gate_h_u_cla32_and10027_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10027_y0);
  and_gate and_gate_h_u_cla32_and10028_y0(h_u_cla32_and10027_y0, h_u_cla32_and10026_y0, h_u_cla32_and10028_y0);
  and_gate and_gate_h_u_cla32_and10029_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10029_y0);
  and_gate and_gate_h_u_cla32_and10030_y0(h_u_cla32_and10029_y0, h_u_cla32_and10028_y0, h_u_cla32_and10030_y0);
  and_gate and_gate_h_u_cla32_and10031_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10031_y0);
  and_gate and_gate_h_u_cla32_and10032_y0(h_u_cla32_and10031_y0, h_u_cla32_and10030_y0, h_u_cla32_and10032_y0);
  and_gate and_gate_h_u_cla32_and10033_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10033_y0);
  and_gate and_gate_h_u_cla32_and10034_y0(h_u_cla32_and10033_y0, h_u_cla32_and10032_y0, h_u_cla32_and10034_y0);
  and_gate and_gate_h_u_cla32_and10035_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10035_y0);
  and_gate and_gate_h_u_cla32_and10036_y0(h_u_cla32_and10035_y0, h_u_cla32_and10034_y0, h_u_cla32_and10036_y0);
  and_gate and_gate_h_u_cla32_and10037_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10037_y0);
  and_gate and_gate_h_u_cla32_and10038_y0(h_u_cla32_and10037_y0, h_u_cla32_and10036_y0, h_u_cla32_and10038_y0);
  and_gate and_gate_h_u_cla32_and10039_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10039_y0);
  and_gate and_gate_h_u_cla32_and10040_y0(h_u_cla32_and10039_y0, h_u_cla32_and10038_y0, h_u_cla32_and10040_y0);
  and_gate and_gate_h_u_cla32_and10041_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10041_y0);
  and_gate and_gate_h_u_cla32_and10042_y0(h_u_cla32_and10041_y0, h_u_cla32_and10040_y0, h_u_cla32_and10042_y0);
  and_gate and_gate_h_u_cla32_and10043_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10043_y0);
  and_gate and_gate_h_u_cla32_and10044_y0(h_u_cla32_and10043_y0, h_u_cla32_and10042_y0, h_u_cla32_and10044_y0);
  and_gate and_gate_h_u_cla32_and10045_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10045_y0);
  and_gate and_gate_h_u_cla32_and10046_y0(h_u_cla32_and10045_y0, h_u_cla32_and10044_y0, h_u_cla32_and10046_y0);
  and_gate and_gate_h_u_cla32_and10047_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10047_y0);
  and_gate and_gate_h_u_cla32_and10048_y0(h_u_cla32_and10047_y0, h_u_cla32_and10046_y0, h_u_cla32_and10048_y0);
  and_gate and_gate_h_u_cla32_and10049_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10049_y0);
  and_gate and_gate_h_u_cla32_and10050_y0(h_u_cla32_and10049_y0, h_u_cla32_and10048_y0, h_u_cla32_and10050_y0);
  and_gate and_gate_h_u_cla32_and10051_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10051_y0);
  and_gate and_gate_h_u_cla32_and10052_y0(h_u_cla32_and10051_y0, h_u_cla32_and10050_y0, h_u_cla32_and10052_y0);
  and_gate and_gate_h_u_cla32_and10053_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10053_y0);
  and_gate and_gate_h_u_cla32_and10054_y0(h_u_cla32_and10053_y0, h_u_cla32_and10052_y0, h_u_cla32_and10054_y0);
  and_gate and_gate_h_u_cla32_and10055_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10055_y0);
  and_gate and_gate_h_u_cla32_and10056_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10056_y0);
  and_gate and_gate_h_u_cla32_and10057_y0(h_u_cla32_and10056_y0, h_u_cla32_and10055_y0, h_u_cla32_and10057_y0);
  and_gate and_gate_h_u_cla32_and10058_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10058_y0);
  and_gate and_gate_h_u_cla32_and10059_y0(h_u_cla32_and10058_y0, h_u_cla32_and10057_y0, h_u_cla32_and10059_y0);
  and_gate and_gate_h_u_cla32_and10060_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10060_y0);
  and_gate and_gate_h_u_cla32_and10061_y0(h_u_cla32_and10060_y0, h_u_cla32_and10059_y0, h_u_cla32_and10061_y0);
  and_gate and_gate_h_u_cla32_and10062_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10062_y0);
  and_gate and_gate_h_u_cla32_and10063_y0(h_u_cla32_and10062_y0, h_u_cla32_and10061_y0, h_u_cla32_and10063_y0);
  and_gate and_gate_h_u_cla32_and10064_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10064_y0);
  and_gate and_gate_h_u_cla32_and10065_y0(h_u_cla32_and10064_y0, h_u_cla32_and10063_y0, h_u_cla32_and10065_y0);
  and_gate and_gate_h_u_cla32_and10066_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10066_y0);
  and_gate and_gate_h_u_cla32_and10067_y0(h_u_cla32_and10066_y0, h_u_cla32_and10065_y0, h_u_cla32_and10067_y0);
  and_gate and_gate_h_u_cla32_and10068_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10068_y0);
  and_gate and_gate_h_u_cla32_and10069_y0(h_u_cla32_and10068_y0, h_u_cla32_and10067_y0, h_u_cla32_and10069_y0);
  and_gate and_gate_h_u_cla32_and10070_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10070_y0);
  and_gate and_gate_h_u_cla32_and10071_y0(h_u_cla32_and10070_y0, h_u_cla32_and10069_y0, h_u_cla32_and10071_y0);
  and_gate and_gate_h_u_cla32_and10072_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10072_y0);
  and_gate and_gate_h_u_cla32_and10073_y0(h_u_cla32_and10072_y0, h_u_cla32_and10071_y0, h_u_cla32_and10073_y0);
  and_gate and_gate_h_u_cla32_and10074_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10074_y0);
  and_gate and_gate_h_u_cla32_and10075_y0(h_u_cla32_and10074_y0, h_u_cla32_and10073_y0, h_u_cla32_and10075_y0);
  and_gate and_gate_h_u_cla32_and10076_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10076_y0);
  and_gate and_gate_h_u_cla32_and10077_y0(h_u_cla32_and10076_y0, h_u_cla32_and10075_y0, h_u_cla32_and10077_y0);
  and_gate and_gate_h_u_cla32_and10078_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10078_y0);
  and_gate and_gate_h_u_cla32_and10079_y0(h_u_cla32_and10078_y0, h_u_cla32_and10077_y0, h_u_cla32_and10079_y0);
  and_gate and_gate_h_u_cla32_and10080_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10080_y0);
  and_gate and_gate_h_u_cla32_and10081_y0(h_u_cla32_and10080_y0, h_u_cla32_and10079_y0, h_u_cla32_and10081_y0);
  and_gate and_gate_h_u_cla32_and10082_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10082_y0);
  and_gate and_gate_h_u_cla32_and10083_y0(h_u_cla32_and10082_y0, h_u_cla32_and10081_y0, h_u_cla32_and10083_y0);
  and_gate and_gate_h_u_cla32_and10084_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10084_y0);
  and_gate and_gate_h_u_cla32_and10085_y0(h_u_cla32_and10084_y0, h_u_cla32_and10083_y0, h_u_cla32_and10085_y0);
  and_gate and_gate_h_u_cla32_and10086_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10086_y0);
  and_gate and_gate_h_u_cla32_and10087_y0(h_u_cla32_and10086_y0, h_u_cla32_and10085_y0, h_u_cla32_and10087_y0);
  and_gate and_gate_h_u_cla32_and10088_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10088_y0);
  and_gate and_gate_h_u_cla32_and10089_y0(h_u_cla32_and10088_y0, h_u_cla32_and10087_y0, h_u_cla32_and10089_y0);
  and_gate and_gate_h_u_cla32_and10090_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and10090_y0);
  and_gate and_gate_h_u_cla32_and10091_y0(h_u_cla32_and10090_y0, h_u_cla32_and10089_y0, h_u_cla32_and10091_y0);
  and_gate and_gate_h_u_cla32_and10092_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10092_y0);
  and_gate and_gate_h_u_cla32_and10093_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10093_y0);
  and_gate and_gate_h_u_cla32_and10094_y0(h_u_cla32_and10093_y0, h_u_cla32_and10092_y0, h_u_cla32_and10094_y0);
  and_gate and_gate_h_u_cla32_and10095_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10095_y0);
  and_gate and_gate_h_u_cla32_and10096_y0(h_u_cla32_and10095_y0, h_u_cla32_and10094_y0, h_u_cla32_and10096_y0);
  and_gate and_gate_h_u_cla32_and10097_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10097_y0);
  and_gate and_gate_h_u_cla32_and10098_y0(h_u_cla32_and10097_y0, h_u_cla32_and10096_y0, h_u_cla32_and10098_y0);
  and_gate and_gate_h_u_cla32_and10099_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10099_y0);
  and_gate and_gate_h_u_cla32_and10100_y0(h_u_cla32_and10099_y0, h_u_cla32_and10098_y0, h_u_cla32_and10100_y0);
  and_gate and_gate_h_u_cla32_and10101_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10101_y0);
  and_gate and_gate_h_u_cla32_and10102_y0(h_u_cla32_and10101_y0, h_u_cla32_and10100_y0, h_u_cla32_and10102_y0);
  and_gate and_gate_h_u_cla32_and10103_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10103_y0);
  and_gate and_gate_h_u_cla32_and10104_y0(h_u_cla32_and10103_y0, h_u_cla32_and10102_y0, h_u_cla32_and10104_y0);
  and_gate and_gate_h_u_cla32_and10105_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10105_y0);
  and_gate and_gate_h_u_cla32_and10106_y0(h_u_cla32_and10105_y0, h_u_cla32_and10104_y0, h_u_cla32_and10106_y0);
  and_gate and_gate_h_u_cla32_and10107_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10107_y0);
  and_gate and_gate_h_u_cla32_and10108_y0(h_u_cla32_and10107_y0, h_u_cla32_and10106_y0, h_u_cla32_and10108_y0);
  and_gate and_gate_h_u_cla32_and10109_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10109_y0);
  and_gate and_gate_h_u_cla32_and10110_y0(h_u_cla32_and10109_y0, h_u_cla32_and10108_y0, h_u_cla32_and10110_y0);
  and_gate and_gate_h_u_cla32_and10111_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10111_y0);
  and_gate and_gate_h_u_cla32_and10112_y0(h_u_cla32_and10111_y0, h_u_cla32_and10110_y0, h_u_cla32_and10112_y0);
  and_gate and_gate_h_u_cla32_and10113_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10113_y0);
  and_gate and_gate_h_u_cla32_and10114_y0(h_u_cla32_and10113_y0, h_u_cla32_and10112_y0, h_u_cla32_and10114_y0);
  and_gate and_gate_h_u_cla32_and10115_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10115_y0);
  and_gate and_gate_h_u_cla32_and10116_y0(h_u_cla32_and10115_y0, h_u_cla32_and10114_y0, h_u_cla32_and10116_y0);
  and_gate and_gate_h_u_cla32_and10117_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10117_y0);
  and_gate and_gate_h_u_cla32_and10118_y0(h_u_cla32_and10117_y0, h_u_cla32_and10116_y0, h_u_cla32_and10118_y0);
  and_gate and_gate_h_u_cla32_and10119_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10119_y0);
  and_gate and_gate_h_u_cla32_and10120_y0(h_u_cla32_and10119_y0, h_u_cla32_and10118_y0, h_u_cla32_and10120_y0);
  and_gate and_gate_h_u_cla32_and10121_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10121_y0);
  and_gate and_gate_h_u_cla32_and10122_y0(h_u_cla32_and10121_y0, h_u_cla32_and10120_y0, h_u_cla32_and10122_y0);
  and_gate and_gate_h_u_cla32_and10123_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10123_y0);
  and_gate and_gate_h_u_cla32_and10124_y0(h_u_cla32_and10123_y0, h_u_cla32_and10122_y0, h_u_cla32_and10124_y0);
  and_gate and_gate_h_u_cla32_and10125_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and10125_y0);
  and_gate and_gate_h_u_cla32_and10126_y0(h_u_cla32_and10125_y0, h_u_cla32_and10124_y0, h_u_cla32_and10126_y0);
  and_gate and_gate_h_u_cla32_and10127_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10127_y0);
  and_gate and_gate_h_u_cla32_and10128_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10128_y0);
  and_gate and_gate_h_u_cla32_and10129_y0(h_u_cla32_and10128_y0, h_u_cla32_and10127_y0, h_u_cla32_and10129_y0);
  and_gate and_gate_h_u_cla32_and10130_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10130_y0);
  and_gate and_gate_h_u_cla32_and10131_y0(h_u_cla32_and10130_y0, h_u_cla32_and10129_y0, h_u_cla32_and10131_y0);
  and_gate and_gate_h_u_cla32_and10132_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10132_y0);
  and_gate and_gate_h_u_cla32_and10133_y0(h_u_cla32_and10132_y0, h_u_cla32_and10131_y0, h_u_cla32_and10133_y0);
  and_gate and_gate_h_u_cla32_and10134_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10134_y0);
  and_gate and_gate_h_u_cla32_and10135_y0(h_u_cla32_and10134_y0, h_u_cla32_and10133_y0, h_u_cla32_and10135_y0);
  and_gate and_gate_h_u_cla32_and10136_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10136_y0);
  and_gate and_gate_h_u_cla32_and10137_y0(h_u_cla32_and10136_y0, h_u_cla32_and10135_y0, h_u_cla32_and10137_y0);
  and_gate and_gate_h_u_cla32_and10138_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10138_y0);
  and_gate and_gate_h_u_cla32_and10139_y0(h_u_cla32_and10138_y0, h_u_cla32_and10137_y0, h_u_cla32_and10139_y0);
  and_gate and_gate_h_u_cla32_and10140_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10140_y0);
  and_gate and_gate_h_u_cla32_and10141_y0(h_u_cla32_and10140_y0, h_u_cla32_and10139_y0, h_u_cla32_and10141_y0);
  and_gate and_gate_h_u_cla32_and10142_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10142_y0);
  and_gate and_gate_h_u_cla32_and10143_y0(h_u_cla32_and10142_y0, h_u_cla32_and10141_y0, h_u_cla32_and10143_y0);
  and_gate and_gate_h_u_cla32_and10144_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10144_y0);
  and_gate and_gate_h_u_cla32_and10145_y0(h_u_cla32_and10144_y0, h_u_cla32_and10143_y0, h_u_cla32_and10145_y0);
  and_gate and_gate_h_u_cla32_and10146_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10146_y0);
  and_gate and_gate_h_u_cla32_and10147_y0(h_u_cla32_and10146_y0, h_u_cla32_and10145_y0, h_u_cla32_and10147_y0);
  and_gate and_gate_h_u_cla32_and10148_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10148_y0);
  and_gate and_gate_h_u_cla32_and10149_y0(h_u_cla32_and10148_y0, h_u_cla32_and10147_y0, h_u_cla32_and10149_y0);
  and_gate and_gate_h_u_cla32_and10150_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10150_y0);
  and_gate and_gate_h_u_cla32_and10151_y0(h_u_cla32_and10150_y0, h_u_cla32_and10149_y0, h_u_cla32_and10151_y0);
  and_gate and_gate_h_u_cla32_and10152_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10152_y0);
  and_gate and_gate_h_u_cla32_and10153_y0(h_u_cla32_and10152_y0, h_u_cla32_and10151_y0, h_u_cla32_and10153_y0);
  and_gate and_gate_h_u_cla32_and10154_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10154_y0);
  and_gate and_gate_h_u_cla32_and10155_y0(h_u_cla32_and10154_y0, h_u_cla32_and10153_y0, h_u_cla32_and10155_y0);
  and_gate and_gate_h_u_cla32_and10156_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10156_y0);
  and_gate and_gate_h_u_cla32_and10157_y0(h_u_cla32_and10156_y0, h_u_cla32_and10155_y0, h_u_cla32_and10157_y0);
  and_gate and_gate_h_u_cla32_and10158_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and10158_y0);
  and_gate and_gate_h_u_cla32_and10159_y0(h_u_cla32_and10158_y0, h_u_cla32_and10157_y0, h_u_cla32_and10159_y0);
  and_gate and_gate_h_u_cla32_and10160_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10160_y0);
  and_gate and_gate_h_u_cla32_and10161_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10161_y0);
  and_gate and_gate_h_u_cla32_and10162_y0(h_u_cla32_and10161_y0, h_u_cla32_and10160_y0, h_u_cla32_and10162_y0);
  and_gate and_gate_h_u_cla32_and10163_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10163_y0);
  and_gate and_gate_h_u_cla32_and10164_y0(h_u_cla32_and10163_y0, h_u_cla32_and10162_y0, h_u_cla32_and10164_y0);
  and_gate and_gate_h_u_cla32_and10165_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10165_y0);
  and_gate and_gate_h_u_cla32_and10166_y0(h_u_cla32_and10165_y0, h_u_cla32_and10164_y0, h_u_cla32_and10166_y0);
  and_gate and_gate_h_u_cla32_and10167_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10167_y0);
  and_gate and_gate_h_u_cla32_and10168_y0(h_u_cla32_and10167_y0, h_u_cla32_and10166_y0, h_u_cla32_and10168_y0);
  and_gate and_gate_h_u_cla32_and10169_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10169_y0);
  and_gate and_gate_h_u_cla32_and10170_y0(h_u_cla32_and10169_y0, h_u_cla32_and10168_y0, h_u_cla32_and10170_y0);
  and_gate and_gate_h_u_cla32_and10171_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10171_y0);
  and_gate and_gate_h_u_cla32_and10172_y0(h_u_cla32_and10171_y0, h_u_cla32_and10170_y0, h_u_cla32_and10172_y0);
  and_gate and_gate_h_u_cla32_and10173_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10173_y0);
  and_gate and_gate_h_u_cla32_and10174_y0(h_u_cla32_and10173_y0, h_u_cla32_and10172_y0, h_u_cla32_and10174_y0);
  and_gate and_gate_h_u_cla32_and10175_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10175_y0);
  and_gate and_gate_h_u_cla32_and10176_y0(h_u_cla32_and10175_y0, h_u_cla32_and10174_y0, h_u_cla32_and10176_y0);
  and_gate and_gate_h_u_cla32_and10177_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10177_y0);
  and_gate and_gate_h_u_cla32_and10178_y0(h_u_cla32_and10177_y0, h_u_cla32_and10176_y0, h_u_cla32_and10178_y0);
  and_gate and_gate_h_u_cla32_and10179_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10179_y0);
  and_gate and_gate_h_u_cla32_and10180_y0(h_u_cla32_and10179_y0, h_u_cla32_and10178_y0, h_u_cla32_and10180_y0);
  and_gate and_gate_h_u_cla32_and10181_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10181_y0);
  and_gate and_gate_h_u_cla32_and10182_y0(h_u_cla32_and10181_y0, h_u_cla32_and10180_y0, h_u_cla32_and10182_y0);
  and_gate and_gate_h_u_cla32_and10183_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10183_y0);
  and_gate and_gate_h_u_cla32_and10184_y0(h_u_cla32_and10183_y0, h_u_cla32_and10182_y0, h_u_cla32_and10184_y0);
  and_gate and_gate_h_u_cla32_and10185_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10185_y0);
  and_gate and_gate_h_u_cla32_and10186_y0(h_u_cla32_and10185_y0, h_u_cla32_and10184_y0, h_u_cla32_and10186_y0);
  and_gate and_gate_h_u_cla32_and10187_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10187_y0);
  and_gate and_gate_h_u_cla32_and10188_y0(h_u_cla32_and10187_y0, h_u_cla32_and10186_y0, h_u_cla32_and10188_y0);
  and_gate and_gate_h_u_cla32_and10189_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and10189_y0);
  and_gate and_gate_h_u_cla32_and10190_y0(h_u_cla32_and10189_y0, h_u_cla32_and10188_y0, h_u_cla32_and10190_y0);
  and_gate and_gate_h_u_cla32_and10191_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10191_y0);
  and_gate and_gate_h_u_cla32_and10192_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10192_y0);
  and_gate and_gate_h_u_cla32_and10193_y0(h_u_cla32_and10192_y0, h_u_cla32_and10191_y0, h_u_cla32_and10193_y0);
  and_gate and_gate_h_u_cla32_and10194_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10194_y0);
  and_gate and_gate_h_u_cla32_and10195_y0(h_u_cla32_and10194_y0, h_u_cla32_and10193_y0, h_u_cla32_and10195_y0);
  and_gate and_gate_h_u_cla32_and10196_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10196_y0);
  and_gate and_gate_h_u_cla32_and10197_y0(h_u_cla32_and10196_y0, h_u_cla32_and10195_y0, h_u_cla32_and10197_y0);
  and_gate and_gate_h_u_cla32_and10198_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10198_y0);
  and_gate and_gate_h_u_cla32_and10199_y0(h_u_cla32_and10198_y0, h_u_cla32_and10197_y0, h_u_cla32_and10199_y0);
  and_gate and_gate_h_u_cla32_and10200_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10200_y0);
  and_gate and_gate_h_u_cla32_and10201_y0(h_u_cla32_and10200_y0, h_u_cla32_and10199_y0, h_u_cla32_and10201_y0);
  and_gate and_gate_h_u_cla32_and10202_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10202_y0);
  and_gate and_gate_h_u_cla32_and10203_y0(h_u_cla32_and10202_y0, h_u_cla32_and10201_y0, h_u_cla32_and10203_y0);
  and_gate and_gate_h_u_cla32_and10204_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10204_y0);
  and_gate and_gate_h_u_cla32_and10205_y0(h_u_cla32_and10204_y0, h_u_cla32_and10203_y0, h_u_cla32_and10205_y0);
  and_gate and_gate_h_u_cla32_and10206_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10206_y0);
  and_gate and_gate_h_u_cla32_and10207_y0(h_u_cla32_and10206_y0, h_u_cla32_and10205_y0, h_u_cla32_and10207_y0);
  and_gate and_gate_h_u_cla32_and10208_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10208_y0);
  and_gate and_gate_h_u_cla32_and10209_y0(h_u_cla32_and10208_y0, h_u_cla32_and10207_y0, h_u_cla32_and10209_y0);
  and_gate and_gate_h_u_cla32_and10210_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10210_y0);
  and_gate and_gate_h_u_cla32_and10211_y0(h_u_cla32_and10210_y0, h_u_cla32_and10209_y0, h_u_cla32_and10211_y0);
  and_gate and_gate_h_u_cla32_and10212_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10212_y0);
  and_gate and_gate_h_u_cla32_and10213_y0(h_u_cla32_and10212_y0, h_u_cla32_and10211_y0, h_u_cla32_and10213_y0);
  and_gate and_gate_h_u_cla32_and10214_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10214_y0);
  and_gate and_gate_h_u_cla32_and10215_y0(h_u_cla32_and10214_y0, h_u_cla32_and10213_y0, h_u_cla32_and10215_y0);
  and_gate and_gate_h_u_cla32_and10216_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10216_y0);
  and_gate and_gate_h_u_cla32_and10217_y0(h_u_cla32_and10216_y0, h_u_cla32_and10215_y0, h_u_cla32_and10217_y0);
  and_gate and_gate_h_u_cla32_and10218_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and10218_y0);
  and_gate and_gate_h_u_cla32_and10219_y0(h_u_cla32_and10218_y0, h_u_cla32_and10217_y0, h_u_cla32_and10219_y0);
  and_gate and_gate_h_u_cla32_and10220_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10220_y0);
  and_gate and_gate_h_u_cla32_and10221_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10221_y0);
  and_gate and_gate_h_u_cla32_and10222_y0(h_u_cla32_and10221_y0, h_u_cla32_and10220_y0, h_u_cla32_and10222_y0);
  and_gate and_gate_h_u_cla32_and10223_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10223_y0);
  and_gate and_gate_h_u_cla32_and10224_y0(h_u_cla32_and10223_y0, h_u_cla32_and10222_y0, h_u_cla32_and10224_y0);
  and_gate and_gate_h_u_cla32_and10225_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10225_y0);
  and_gate and_gate_h_u_cla32_and10226_y0(h_u_cla32_and10225_y0, h_u_cla32_and10224_y0, h_u_cla32_and10226_y0);
  and_gate and_gate_h_u_cla32_and10227_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10227_y0);
  and_gate and_gate_h_u_cla32_and10228_y0(h_u_cla32_and10227_y0, h_u_cla32_and10226_y0, h_u_cla32_and10228_y0);
  and_gate and_gate_h_u_cla32_and10229_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10229_y0);
  and_gate and_gate_h_u_cla32_and10230_y0(h_u_cla32_and10229_y0, h_u_cla32_and10228_y0, h_u_cla32_and10230_y0);
  and_gate and_gate_h_u_cla32_and10231_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10231_y0);
  and_gate and_gate_h_u_cla32_and10232_y0(h_u_cla32_and10231_y0, h_u_cla32_and10230_y0, h_u_cla32_and10232_y0);
  and_gate and_gate_h_u_cla32_and10233_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10233_y0);
  and_gate and_gate_h_u_cla32_and10234_y0(h_u_cla32_and10233_y0, h_u_cla32_and10232_y0, h_u_cla32_and10234_y0);
  and_gate and_gate_h_u_cla32_and10235_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10235_y0);
  and_gate and_gate_h_u_cla32_and10236_y0(h_u_cla32_and10235_y0, h_u_cla32_and10234_y0, h_u_cla32_and10236_y0);
  and_gate and_gate_h_u_cla32_and10237_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10237_y0);
  and_gate and_gate_h_u_cla32_and10238_y0(h_u_cla32_and10237_y0, h_u_cla32_and10236_y0, h_u_cla32_and10238_y0);
  and_gate and_gate_h_u_cla32_and10239_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10239_y0);
  and_gate and_gate_h_u_cla32_and10240_y0(h_u_cla32_and10239_y0, h_u_cla32_and10238_y0, h_u_cla32_and10240_y0);
  and_gate and_gate_h_u_cla32_and10241_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10241_y0);
  and_gate and_gate_h_u_cla32_and10242_y0(h_u_cla32_and10241_y0, h_u_cla32_and10240_y0, h_u_cla32_and10242_y0);
  and_gate and_gate_h_u_cla32_and10243_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10243_y0);
  and_gate and_gate_h_u_cla32_and10244_y0(h_u_cla32_and10243_y0, h_u_cla32_and10242_y0, h_u_cla32_and10244_y0);
  and_gate and_gate_h_u_cla32_and10245_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and10245_y0);
  and_gate and_gate_h_u_cla32_and10246_y0(h_u_cla32_and10245_y0, h_u_cla32_and10244_y0, h_u_cla32_and10246_y0);
  and_gate and_gate_h_u_cla32_and10247_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10247_y0);
  and_gate and_gate_h_u_cla32_and10248_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10248_y0);
  and_gate and_gate_h_u_cla32_and10249_y0(h_u_cla32_and10248_y0, h_u_cla32_and10247_y0, h_u_cla32_and10249_y0);
  and_gate and_gate_h_u_cla32_and10250_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10250_y0);
  and_gate and_gate_h_u_cla32_and10251_y0(h_u_cla32_and10250_y0, h_u_cla32_and10249_y0, h_u_cla32_and10251_y0);
  and_gate and_gate_h_u_cla32_and10252_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10252_y0);
  and_gate and_gate_h_u_cla32_and10253_y0(h_u_cla32_and10252_y0, h_u_cla32_and10251_y0, h_u_cla32_and10253_y0);
  and_gate and_gate_h_u_cla32_and10254_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10254_y0);
  and_gate and_gate_h_u_cla32_and10255_y0(h_u_cla32_and10254_y0, h_u_cla32_and10253_y0, h_u_cla32_and10255_y0);
  and_gate and_gate_h_u_cla32_and10256_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10256_y0);
  and_gate and_gate_h_u_cla32_and10257_y0(h_u_cla32_and10256_y0, h_u_cla32_and10255_y0, h_u_cla32_and10257_y0);
  and_gate and_gate_h_u_cla32_and10258_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10258_y0);
  and_gate and_gate_h_u_cla32_and10259_y0(h_u_cla32_and10258_y0, h_u_cla32_and10257_y0, h_u_cla32_and10259_y0);
  and_gate and_gate_h_u_cla32_and10260_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10260_y0);
  and_gate and_gate_h_u_cla32_and10261_y0(h_u_cla32_and10260_y0, h_u_cla32_and10259_y0, h_u_cla32_and10261_y0);
  and_gate and_gate_h_u_cla32_and10262_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10262_y0);
  and_gate and_gate_h_u_cla32_and10263_y0(h_u_cla32_and10262_y0, h_u_cla32_and10261_y0, h_u_cla32_and10263_y0);
  and_gate and_gate_h_u_cla32_and10264_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10264_y0);
  and_gate and_gate_h_u_cla32_and10265_y0(h_u_cla32_and10264_y0, h_u_cla32_and10263_y0, h_u_cla32_and10265_y0);
  and_gate and_gate_h_u_cla32_and10266_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10266_y0);
  and_gate and_gate_h_u_cla32_and10267_y0(h_u_cla32_and10266_y0, h_u_cla32_and10265_y0, h_u_cla32_and10267_y0);
  and_gate and_gate_h_u_cla32_and10268_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10268_y0);
  and_gate and_gate_h_u_cla32_and10269_y0(h_u_cla32_and10268_y0, h_u_cla32_and10267_y0, h_u_cla32_and10269_y0);
  and_gate and_gate_h_u_cla32_and10270_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and10270_y0);
  and_gate and_gate_h_u_cla32_and10271_y0(h_u_cla32_and10270_y0, h_u_cla32_and10269_y0, h_u_cla32_and10271_y0);
  and_gate and_gate_h_u_cla32_and10272_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10272_y0);
  and_gate and_gate_h_u_cla32_and10273_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10273_y0);
  and_gate and_gate_h_u_cla32_and10274_y0(h_u_cla32_and10273_y0, h_u_cla32_and10272_y0, h_u_cla32_and10274_y0);
  and_gate and_gate_h_u_cla32_and10275_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10275_y0);
  and_gate and_gate_h_u_cla32_and10276_y0(h_u_cla32_and10275_y0, h_u_cla32_and10274_y0, h_u_cla32_and10276_y0);
  and_gate and_gate_h_u_cla32_and10277_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10277_y0);
  and_gate and_gate_h_u_cla32_and10278_y0(h_u_cla32_and10277_y0, h_u_cla32_and10276_y0, h_u_cla32_and10278_y0);
  and_gate and_gate_h_u_cla32_and10279_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10279_y0);
  and_gate and_gate_h_u_cla32_and10280_y0(h_u_cla32_and10279_y0, h_u_cla32_and10278_y0, h_u_cla32_and10280_y0);
  and_gate and_gate_h_u_cla32_and10281_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10281_y0);
  and_gate and_gate_h_u_cla32_and10282_y0(h_u_cla32_and10281_y0, h_u_cla32_and10280_y0, h_u_cla32_and10282_y0);
  and_gate and_gate_h_u_cla32_and10283_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10283_y0);
  and_gate and_gate_h_u_cla32_and10284_y0(h_u_cla32_and10283_y0, h_u_cla32_and10282_y0, h_u_cla32_and10284_y0);
  and_gate and_gate_h_u_cla32_and10285_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10285_y0);
  and_gate and_gate_h_u_cla32_and10286_y0(h_u_cla32_and10285_y0, h_u_cla32_and10284_y0, h_u_cla32_and10286_y0);
  and_gate and_gate_h_u_cla32_and10287_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10287_y0);
  and_gate and_gate_h_u_cla32_and10288_y0(h_u_cla32_and10287_y0, h_u_cla32_and10286_y0, h_u_cla32_and10288_y0);
  and_gate and_gate_h_u_cla32_and10289_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10289_y0);
  and_gate and_gate_h_u_cla32_and10290_y0(h_u_cla32_and10289_y0, h_u_cla32_and10288_y0, h_u_cla32_and10290_y0);
  and_gate and_gate_h_u_cla32_and10291_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10291_y0);
  and_gate and_gate_h_u_cla32_and10292_y0(h_u_cla32_and10291_y0, h_u_cla32_and10290_y0, h_u_cla32_and10292_y0);
  and_gate and_gate_h_u_cla32_and10293_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and10293_y0);
  and_gate and_gate_h_u_cla32_and10294_y0(h_u_cla32_and10293_y0, h_u_cla32_and10292_y0, h_u_cla32_and10294_y0);
  and_gate and_gate_h_u_cla32_and10295_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10295_y0);
  and_gate and_gate_h_u_cla32_and10296_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10296_y0);
  and_gate and_gate_h_u_cla32_and10297_y0(h_u_cla32_and10296_y0, h_u_cla32_and10295_y0, h_u_cla32_and10297_y0);
  and_gate and_gate_h_u_cla32_and10298_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10298_y0);
  and_gate and_gate_h_u_cla32_and10299_y0(h_u_cla32_and10298_y0, h_u_cla32_and10297_y0, h_u_cla32_and10299_y0);
  and_gate and_gate_h_u_cla32_and10300_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10300_y0);
  and_gate and_gate_h_u_cla32_and10301_y0(h_u_cla32_and10300_y0, h_u_cla32_and10299_y0, h_u_cla32_and10301_y0);
  and_gate and_gate_h_u_cla32_and10302_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10302_y0);
  and_gate and_gate_h_u_cla32_and10303_y0(h_u_cla32_and10302_y0, h_u_cla32_and10301_y0, h_u_cla32_and10303_y0);
  and_gate and_gate_h_u_cla32_and10304_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10304_y0);
  and_gate and_gate_h_u_cla32_and10305_y0(h_u_cla32_and10304_y0, h_u_cla32_and10303_y0, h_u_cla32_and10305_y0);
  and_gate and_gate_h_u_cla32_and10306_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10306_y0);
  and_gate and_gate_h_u_cla32_and10307_y0(h_u_cla32_and10306_y0, h_u_cla32_and10305_y0, h_u_cla32_and10307_y0);
  and_gate and_gate_h_u_cla32_and10308_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10308_y0);
  and_gate and_gate_h_u_cla32_and10309_y0(h_u_cla32_and10308_y0, h_u_cla32_and10307_y0, h_u_cla32_and10309_y0);
  and_gate and_gate_h_u_cla32_and10310_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10310_y0);
  and_gate and_gate_h_u_cla32_and10311_y0(h_u_cla32_and10310_y0, h_u_cla32_and10309_y0, h_u_cla32_and10311_y0);
  and_gate and_gate_h_u_cla32_and10312_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10312_y0);
  and_gate and_gate_h_u_cla32_and10313_y0(h_u_cla32_and10312_y0, h_u_cla32_and10311_y0, h_u_cla32_and10313_y0);
  and_gate and_gate_h_u_cla32_and10314_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and10314_y0);
  and_gate and_gate_h_u_cla32_and10315_y0(h_u_cla32_and10314_y0, h_u_cla32_and10313_y0, h_u_cla32_and10315_y0);
  and_gate and_gate_h_u_cla32_and10316_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10316_y0);
  and_gate and_gate_h_u_cla32_and10317_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10317_y0);
  and_gate and_gate_h_u_cla32_and10318_y0(h_u_cla32_and10317_y0, h_u_cla32_and10316_y0, h_u_cla32_and10318_y0);
  and_gate and_gate_h_u_cla32_and10319_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10319_y0);
  and_gate and_gate_h_u_cla32_and10320_y0(h_u_cla32_and10319_y0, h_u_cla32_and10318_y0, h_u_cla32_and10320_y0);
  and_gate and_gate_h_u_cla32_and10321_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10321_y0);
  and_gate and_gate_h_u_cla32_and10322_y0(h_u_cla32_and10321_y0, h_u_cla32_and10320_y0, h_u_cla32_and10322_y0);
  and_gate and_gate_h_u_cla32_and10323_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10323_y0);
  and_gate and_gate_h_u_cla32_and10324_y0(h_u_cla32_and10323_y0, h_u_cla32_and10322_y0, h_u_cla32_and10324_y0);
  and_gate and_gate_h_u_cla32_and10325_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10325_y0);
  and_gate and_gate_h_u_cla32_and10326_y0(h_u_cla32_and10325_y0, h_u_cla32_and10324_y0, h_u_cla32_and10326_y0);
  and_gate and_gate_h_u_cla32_and10327_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10327_y0);
  and_gate and_gate_h_u_cla32_and10328_y0(h_u_cla32_and10327_y0, h_u_cla32_and10326_y0, h_u_cla32_and10328_y0);
  and_gate and_gate_h_u_cla32_and10329_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10329_y0);
  and_gate and_gate_h_u_cla32_and10330_y0(h_u_cla32_and10329_y0, h_u_cla32_and10328_y0, h_u_cla32_and10330_y0);
  and_gate and_gate_h_u_cla32_and10331_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10331_y0);
  and_gate and_gate_h_u_cla32_and10332_y0(h_u_cla32_and10331_y0, h_u_cla32_and10330_y0, h_u_cla32_and10332_y0);
  and_gate and_gate_h_u_cla32_and10333_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and10333_y0);
  and_gate and_gate_h_u_cla32_and10334_y0(h_u_cla32_and10333_y0, h_u_cla32_and10332_y0, h_u_cla32_and10334_y0);
  and_gate and_gate_h_u_cla32_and10335_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10335_y0);
  and_gate and_gate_h_u_cla32_and10336_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10336_y0);
  and_gate and_gate_h_u_cla32_and10337_y0(h_u_cla32_and10336_y0, h_u_cla32_and10335_y0, h_u_cla32_and10337_y0);
  and_gate and_gate_h_u_cla32_and10338_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10338_y0);
  and_gate and_gate_h_u_cla32_and10339_y0(h_u_cla32_and10338_y0, h_u_cla32_and10337_y0, h_u_cla32_and10339_y0);
  and_gate and_gate_h_u_cla32_and10340_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10340_y0);
  and_gate and_gate_h_u_cla32_and10341_y0(h_u_cla32_and10340_y0, h_u_cla32_and10339_y0, h_u_cla32_and10341_y0);
  and_gate and_gate_h_u_cla32_and10342_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10342_y0);
  and_gate and_gate_h_u_cla32_and10343_y0(h_u_cla32_and10342_y0, h_u_cla32_and10341_y0, h_u_cla32_and10343_y0);
  and_gate and_gate_h_u_cla32_and10344_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10344_y0);
  and_gate and_gate_h_u_cla32_and10345_y0(h_u_cla32_and10344_y0, h_u_cla32_and10343_y0, h_u_cla32_and10345_y0);
  and_gate and_gate_h_u_cla32_and10346_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10346_y0);
  and_gate and_gate_h_u_cla32_and10347_y0(h_u_cla32_and10346_y0, h_u_cla32_and10345_y0, h_u_cla32_and10347_y0);
  and_gate and_gate_h_u_cla32_and10348_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10348_y0);
  and_gate and_gate_h_u_cla32_and10349_y0(h_u_cla32_and10348_y0, h_u_cla32_and10347_y0, h_u_cla32_and10349_y0);
  and_gate and_gate_h_u_cla32_and10350_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and10350_y0);
  and_gate and_gate_h_u_cla32_and10351_y0(h_u_cla32_and10350_y0, h_u_cla32_and10349_y0, h_u_cla32_and10351_y0);
  and_gate and_gate_h_u_cla32_and10352_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10352_y0);
  and_gate and_gate_h_u_cla32_and10353_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10353_y0);
  and_gate and_gate_h_u_cla32_and10354_y0(h_u_cla32_and10353_y0, h_u_cla32_and10352_y0, h_u_cla32_and10354_y0);
  and_gate and_gate_h_u_cla32_and10355_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10355_y0);
  and_gate and_gate_h_u_cla32_and10356_y0(h_u_cla32_and10355_y0, h_u_cla32_and10354_y0, h_u_cla32_and10356_y0);
  and_gate and_gate_h_u_cla32_and10357_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10357_y0);
  and_gate and_gate_h_u_cla32_and10358_y0(h_u_cla32_and10357_y0, h_u_cla32_and10356_y0, h_u_cla32_and10358_y0);
  and_gate and_gate_h_u_cla32_and10359_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10359_y0);
  and_gate and_gate_h_u_cla32_and10360_y0(h_u_cla32_and10359_y0, h_u_cla32_and10358_y0, h_u_cla32_and10360_y0);
  and_gate and_gate_h_u_cla32_and10361_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10361_y0);
  and_gate and_gate_h_u_cla32_and10362_y0(h_u_cla32_and10361_y0, h_u_cla32_and10360_y0, h_u_cla32_and10362_y0);
  and_gate and_gate_h_u_cla32_and10363_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10363_y0);
  and_gate and_gate_h_u_cla32_and10364_y0(h_u_cla32_and10363_y0, h_u_cla32_and10362_y0, h_u_cla32_and10364_y0);
  and_gate and_gate_h_u_cla32_and10365_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and10365_y0);
  and_gate and_gate_h_u_cla32_and10366_y0(h_u_cla32_and10365_y0, h_u_cla32_and10364_y0, h_u_cla32_and10366_y0);
  and_gate and_gate_h_u_cla32_and10367_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10367_y0);
  and_gate and_gate_h_u_cla32_and10368_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10368_y0);
  and_gate and_gate_h_u_cla32_and10369_y0(h_u_cla32_and10368_y0, h_u_cla32_and10367_y0, h_u_cla32_and10369_y0);
  and_gate and_gate_h_u_cla32_and10370_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10370_y0);
  and_gate and_gate_h_u_cla32_and10371_y0(h_u_cla32_and10370_y0, h_u_cla32_and10369_y0, h_u_cla32_and10371_y0);
  and_gate and_gate_h_u_cla32_and10372_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10372_y0);
  and_gate and_gate_h_u_cla32_and10373_y0(h_u_cla32_and10372_y0, h_u_cla32_and10371_y0, h_u_cla32_and10373_y0);
  and_gate and_gate_h_u_cla32_and10374_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10374_y0);
  and_gate and_gate_h_u_cla32_and10375_y0(h_u_cla32_and10374_y0, h_u_cla32_and10373_y0, h_u_cla32_and10375_y0);
  and_gate and_gate_h_u_cla32_and10376_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10376_y0);
  and_gate and_gate_h_u_cla32_and10377_y0(h_u_cla32_and10376_y0, h_u_cla32_and10375_y0, h_u_cla32_and10377_y0);
  and_gate and_gate_h_u_cla32_and10378_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and10378_y0);
  and_gate and_gate_h_u_cla32_and10379_y0(h_u_cla32_and10378_y0, h_u_cla32_and10377_y0, h_u_cla32_and10379_y0);
  and_gate and_gate_h_u_cla32_and10380_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and10380_y0);
  and_gate and_gate_h_u_cla32_and10381_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and10381_y0);
  and_gate and_gate_h_u_cla32_and10382_y0(h_u_cla32_and10381_y0, h_u_cla32_and10380_y0, h_u_cla32_and10382_y0);
  and_gate and_gate_h_u_cla32_and10383_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and10383_y0);
  and_gate and_gate_h_u_cla32_and10384_y0(h_u_cla32_and10383_y0, h_u_cla32_and10382_y0, h_u_cla32_and10384_y0);
  and_gate and_gate_h_u_cla32_and10385_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and10385_y0);
  and_gate and_gate_h_u_cla32_and10386_y0(h_u_cla32_and10385_y0, h_u_cla32_and10384_y0, h_u_cla32_and10386_y0);
  and_gate and_gate_h_u_cla32_and10387_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and10387_y0);
  and_gate and_gate_h_u_cla32_and10388_y0(h_u_cla32_and10387_y0, h_u_cla32_and10386_y0, h_u_cla32_and10388_y0);
  and_gate and_gate_h_u_cla32_and10389_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and10389_y0);
  and_gate and_gate_h_u_cla32_and10390_y0(h_u_cla32_and10389_y0, h_u_cla32_and10388_y0, h_u_cla32_and10390_y0);
  and_gate and_gate_h_u_cla32_and10391_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and10391_y0);
  and_gate and_gate_h_u_cla32_and10392_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and10392_y0);
  and_gate and_gate_h_u_cla32_and10393_y0(h_u_cla32_and10392_y0, h_u_cla32_and10391_y0, h_u_cla32_and10393_y0);
  and_gate and_gate_h_u_cla32_and10394_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and10394_y0);
  and_gate and_gate_h_u_cla32_and10395_y0(h_u_cla32_and10394_y0, h_u_cla32_and10393_y0, h_u_cla32_and10395_y0);
  and_gate and_gate_h_u_cla32_and10396_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and10396_y0);
  and_gate and_gate_h_u_cla32_and10397_y0(h_u_cla32_and10396_y0, h_u_cla32_and10395_y0, h_u_cla32_and10397_y0);
  and_gate and_gate_h_u_cla32_and10398_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and10398_y0);
  and_gate and_gate_h_u_cla32_and10399_y0(h_u_cla32_and10398_y0, h_u_cla32_and10397_y0, h_u_cla32_and10399_y0);
  and_gate and_gate_h_u_cla32_and10400_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and10400_y0);
  and_gate and_gate_h_u_cla32_and10401_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and10401_y0);
  and_gate and_gate_h_u_cla32_and10402_y0(h_u_cla32_and10401_y0, h_u_cla32_and10400_y0, h_u_cla32_and10402_y0);
  and_gate and_gate_h_u_cla32_and10403_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and10403_y0);
  and_gate and_gate_h_u_cla32_and10404_y0(h_u_cla32_and10403_y0, h_u_cla32_and10402_y0, h_u_cla32_and10404_y0);
  and_gate and_gate_h_u_cla32_and10405_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and10405_y0);
  and_gate and_gate_h_u_cla32_and10406_y0(h_u_cla32_and10405_y0, h_u_cla32_and10404_y0, h_u_cla32_and10406_y0);
  and_gate and_gate_h_u_cla32_and10407_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and10407_y0);
  and_gate and_gate_h_u_cla32_and10408_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and10408_y0);
  and_gate and_gate_h_u_cla32_and10409_y0(h_u_cla32_and10408_y0, h_u_cla32_and10407_y0, h_u_cla32_and10409_y0);
  and_gate and_gate_h_u_cla32_and10410_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and10410_y0);
  and_gate and_gate_h_u_cla32_and10411_y0(h_u_cla32_and10410_y0, h_u_cla32_and10409_y0, h_u_cla32_and10411_y0);
  and_gate and_gate_h_u_cla32_and10412_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_and10412_y0);
  and_gate and_gate_h_u_cla32_and10413_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_and10413_y0);
  and_gate and_gate_h_u_cla32_and10414_y0(h_u_cla32_and10413_y0, h_u_cla32_and10412_y0, h_u_cla32_and10414_y0);
  and_gate and_gate_h_u_cla32_and10415_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic29_y1, h_u_cla32_and10415_y0);
  or_gate or_gate_h_u_cla32_or465_y0(h_u_cla32_and10415_y0, h_u_cla32_and9515_y0, h_u_cla32_or465_y0);
  or_gate or_gate_h_u_cla32_or466_y0(h_u_cla32_or465_y0, h_u_cla32_and9574_y0, h_u_cla32_or466_y0);
  or_gate or_gate_h_u_cla32_or467_y0(h_u_cla32_or466_y0, h_u_cla32_and9631_y0, h_u_cla32_or467_y0);
  or_gate or_gate_h_u_cla32_or468_y0(h_u_cla32_or467_y0, h_u_cla32_and9686_y0, h_u_cla32_or468_y0);
  or_gate or_gate_h_u_cla32_or469_y0(h_u_cla32_or468_y0, h_u_cla32_and9739_y0, h_u_cla32_or469_y0);
  or_gate or_gate_h_u_cla32_or470_y0(h_u_cla32_or469_y0, h_u_cla32_and9790_y0, h_u_cla32_or470_y0);
  or_gate or_gate_h_u_cla32_or471_y0(h_u_cla32_or470_y0, h_u_cla32_and9839_y0, h_u_cla32_or471_y0);
  or_gate or_gate_h_u_cla32_or472_y0(h_u_cla32_or471_y0, h_u_cla32_and9886_y0, h_u_cla32_or472_y0);
  or_gate or_gate_h_u_cla32_or473_y0(h_u_cla32_or472_y0, h_u_cla32_and9931_y0, h_u_cla32_or473_y0);
  or_gate or_gate_h_u_cla32_or474_y0(h_u_cla32_or473_y0, h_u_cla32_and9974_y0, h_u_cla32_or474_y0);
  or_gate or_gate_h_u_cla32_or475_y0(h_u_cla32_or474_y0, h_u_cla32_and10015_y0, h_u_cla32_or475_y0);
  or_gate or_gate_h_u_cla32_or476_y0(h_u_cla32_or475_y0, h_u_cla32_and10054_y0, h_u_cla32_or476_y0);
  or_gate or_gate_h_u_cla32_or477_y0(h_u_cla32_or476_y0, h_u_cla32_and10091_y0, h_u_cla32_or477_y0);
  or_gate or_gate_h_u_cla32_or478_y0(h_u_cla32_or477_y0, h_u_cla32_and10126_y0, h_u_cla32_or478_y0);
  or_gate or_gate_h_u_cla32_or479_y0(h_u_cla32_or478_y0, h_u_cla32_and10159_y0, h_u_cla32_or479_y0);
  or_gate or_gate_h_u_cla32_or480_y0(h_u_cla32_or479_y0, h_u_cla32_and10190_y0, h_u_cla32_or480_y0);
  or_gate or_gate_h_u_cla32_or481_y0(h_u_cla32_or480_y0, h_u_cla32_and10219_y0, h_u_cla32_or481_y0);
  or_gate or_gate_h_u_cla32_or482_y0(h_u_cla32_or481_y0, h_u_cla32_and10246_y0, h_u_cla32_or482_y0);
  or_gate or_gate_h_u_cla32_or483_y0(h_u_cla32_or482_y0, h_u_cla32_and10271_y0, h_u_cla32_or483_y0);
  or_gate or_gate_h_u_cla32_or484_y0(h_u_cla32_or483_y0, h_u_cla32_and10294_y0, h_u_cla32_or484_y0);
  or_gate or_gate_h_u_cla32_or485_y0(h_u_cla32_or484_y0, h_u_cla32_and10315_y0, h_u_cla32_or485_y0);
  or_gate or_gate_h_u_cla32_or486_y0(h_u_cla32_or485_y0, h_u_cla32_and10334_y0, h_u_cla32_or486_y0);
  or_gate or_gate_h_u_cla32_or487_y0(h_u_cla32_or486_y0, h_u_cla32_and10351_y0, h_u_cla32_or487_y0);
  or_gate or_gate_h_u_cla32_or488_y0(h_u_cla32_or487_y0, h_u_cla32_and10366_y0, h_u_cla32_or488_y0);
  or_gate or_gate_h_u_cla32_or489_y0(h_u_cla32_or488_y0, h_u_cla32_and10379_y0, h_u_cla32_or489_y0);
  or_gate or_gate_h_u_cla32_or490_y0(h_u_cla32_or489_y0, h_u_cla32_and10390_y0, h_u_cla32_or490_y0);
  or_gate or_gate_h_u_cla32_or491_y0(h_u_cla32_or490_y0, h_u_cla32_and10399_y0, h_u_cla32_or491_y0);
  or_gate or_gate_h_u_cla32_or492_y0(h_u_cla32_or491_y0, h_u_cla32_and10406_y0, h_u_cla32_or492_y0);
  or_gate or_gate_h_u_cla32_or493_y0(h_u_cla32_or492_y0, h_u_cla32_and10411_y0, h_u_cla32_or493_y0);
  or_gate or_gate_h_u_cla32_or494_y0(h_u_cla32_or493_y0, h_u_cla32_and10414_y0, h_u_cla32_or494_y0);
  or_gate or_gate_h_u_cla32_or495_y0(h_u_cla32_pg_logic30_y1, h_u_cla32_or494_y0, h_u_cla32_or495_y0);
  pg_logic pg_logic_h_u_cla32_pg_logic31_y0(a_31, b_31, h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic31_y1, h_u_cla32_pg_logic31_y2);
  xor_gate xor_gate_h_u_cla32_xor31_y0(h_u_cla32_pg_logic31_y2, h_u_cla32_or495_y0, h_u_cla32_xor31_y0);
  and_gate and_gate_h_u_cla32_and10416_y0(h_u_cla32_pg_logic0_y0, constant_wire_0, h_u_cla32_and10416_y0);
  and_gate and_gate_h_u_cla32_and10417_y0(h_u_cla32_pg_logic1_y0, constant_wire_0, h_u_cla32_and10417_y0);
  and_gate and_gate_h_u_cla32_and10418_y0(h_u_cla32_and10417_y0, h_u_cla32_and10416_y0, h_u_cla32_and10418_y0);
  and_gate and_gate_h_u_cla32_and10419_y0(h_u_cla32_pg_logic2_y0, constant_wire_0, h_u_cla32_and10419_y0);
  and_gate and_gate_h_u_cla32_and10420_y0(h_u_cla32_and10419_y0, h_u_cla32_and10418_y0, h_u_cla32_and10420_y0);
  and_gate and_gate_h_u_cla32_and10421_y0(h_u_cla32_pg_logic3_y0, constant_wire_0, h_u_cla32_and10421_y0);
  and_gate and_gate_h_u_cla32_and10422_y0(h_u_cla32_and10421_y0, h_u_cla32_and10420_y0, h_u_cla32_and10422_y0);
  and_gate and_gate_h_u_cla32_and10423_y0(h_u_cla32_pg_logic4_y0, constant_wire_0, h_u_cla32_and10423_y0);
  and_gate and_gate_h_u_cla32_and10424_y0(h_u_cla32_and10423_y0, h_u_cla32_and10422_y0, h_u_cla32_and10424_y0);
  and_gate and_gate_h_u_cla32_and10425_y0(h_u_cla32_pg_logic5_y0, constant_wire_0, h_u_cla32_and10425_y0);
  and_gate and_gate_h_u_cla32_and10426_y0(h_u_cla32_and10425_y0, h_u_cla32_and10424_y0, h_u_cla32_and10426_y0);
  and_gate and_gate_h_u_cla32_and10427_y0(h_u_cla32_pg_logic6_y0, constant_wire_0, h_u_cla32_and10427_y0);
  and_gate and_gate_h_u_cla32_and10428_y0(h_u_cla32_and10427_y0, h_u_cla32_and10426_y0, h_u_cla32_and10428_y0);
  and_gate and_gate_h_u_cla32_and10429_y0(h_u_cla32_pg_logic7_y0, constant_wire_0, h_u_cla32_and10429_y0);
  and_gate and_gate_h_u_cla32_and10430_y0(h_u_cla32_and10429_y0, h_u_cla32_and10428_y0, h_u_cla32_and10430_y0);
  and_gate and_gate_h_u_cla32_and10431_y0(h_u_cla32_pg_logic8_y0, constant_wire_0, h_u_cla32_and10431_y0);
  and_gate and_gate_h_u_cla32_and10432_y0(h_u_cla32_and10431_y0, h_u_cla32_and10430_y0, h_u_cla32_and10432_y0);
  and_gate and_gate_h_u_cla32_and10433_y0(h_u_cla32_pg_logic9_y0, constant_wire_0, h_u_cla32_and10433_y0);
  and_gate and_gate_h_u_cla32_and10434_y0(h_u_cla32_and10433_y0, h_u_cla32_and10432_y0, h_u_cla32_and10434_y0);
  and_gate and_gate_h_u_cla32_and10435_y0(h_u_cla32_pg_logic10_y0, constant_wire_0, h_u_cla32_and10435_y0);
  and_gate and_gate_h_u_cla32_and10436_y0(h_u_cla32_and10435_y0, h_u_cla32_and10434_y0, h_u_cla32_and10436_y0);
  and_gate and_gate_h_u_cla32_and10437_y0(h_u_cla32_pg_logic11_y0, constant_wire_0, h_u_cla32_and10437_y0);
  and_gate and_gate_h_u_cla32_and10438_y0(h_u_cla32_and10437_y0, h_u_cla32_and10436_y0, h_u_cla32_and10438_y0);
  and_gate and_gate_h_u_cla32_and10439_y0(h_u_cla32_pg_logic12_y0, constant_wire_0, h_u_cla32_and10439_y0);
  and_gate and_gate_h_u_cla32_and10440_y0(h_u_cla32_and10439_y0, h_u_cla32_and10438_y0, h_u_cla32_and10440_y0);
  and_gate and_gate_h_u_cla32_and10441_y0(h_u_cla32_pg_logic13_y0, constant_wire_0, h_u_cla32_and10441_y0);
  and_gate and_gate_h_u_cla32_and10442_y0(h_u_cla32_and10441_y0, h_u_cla32_and10440_y0, h_u_cla32_and10442_y0);
  and_gate and_gate_h_u_cla32_and10443_y0(h_u_cla32_pg_logic14_y0, constant_wire_0, h_u_cla32_and10443_y0);
  and_gate and_gate_h_u_cla32_and10444_y0(h_u_cla32_and10443_y0, h_u_cla32_and10442_y0, h_u_cla32_and10444_y0);
  and_gate and_gate_h_u_cla32_and10445_y0(h_u_cla32_pg_logic15_y0, constant_wire_0, h_u_cla32_and10445_y0);
  and_gate and_gate_h_u_cla32_and10446_y0(h_u_cla32_and10445_y0, h_u_cla32_and10444_y0, h_u_cla32_and10446_y0);
  and_gate and_gate_h_u_cla32_and10447_y0(h_u_cla32_pg_logic16_y0, constant_wire_0, h_u_cla32_and10447_y0);
  and_gate and_gate_h_u_cla32_and10448_y0(h_u_cla32_and10447_y0, h_u_cla32_and10446_y0, h_u_cla32_and10448_y0);
  and_gate and_gate_h_u_cla32_and10449_y0(h_u_cla32_pg_logic17_y0, constant_wire_0, h_u_cla32_and10449_y0);
  and_gate and_gate_h_u_cla32_and10450_y0(h_u_cla32_and10449_y0, h_u_cla32_and10448_y0, h_u_cla32_and10450_y0);
  and_gate and_gate_h_u_cla32_and10451_y0(h_u_cla32_pg_logic18_y0, constant_wire_0, h_u_cla32_and10451_y0);
  and_gate and_gate_h_u_cla32_and10452_y0(h_u_cla32_and10451_y0, h_u_cla32_and10450_y0, h_u_cla32_and10452_y0);
  and_gate and_gate_h_u_cla32_and10453_y0(h_u_cla32_pg_logic19_y0, constant_wire_0, h_u_cla32_and10453_y0);
  and_gate and_gate_h_u_cla32_and10454_y0(h_u_cla32_and10453_y0, h_u_cla32_and10452_y0, h_u_cla32_and10454_y0);
  and_gate and_gate_h_u_cla32_and10455_y0(h_u_cla32_pg_logic20_y0, constant_wire_0, h_u_cla32_and10455_y0);
  and_gate and_gate_h_u_cla32_and10456_y0(h_u_cla32_and10455_y0, h_u_cla32_and10454_y0, h_u_cla32_and10456_y0);
  and_gate and_gate_h_u_cla32_and10457_y0(h_u_cla32_pg_logic21_y0, constant_wire_0, h_u_cla32_and10457_y0);
  and_gate and_gate_h_u_cla32_and10458_y0(h_u_cla32_and10457_y0, h_u_cla32_and10456_y0, h_u_cla32_and10458_y0);
  and_gate and_gate_h_u_cla32_and10459_y0(h_u_cla32_pg_logic22_y0, constant_wire_0, h_u_cla32_and10459_y0);
  and_gate and_gate_h_u_cla32_and10460_y0(h_u_cla32_and10459_y0, h_u_cla32_and10458_y0, h_u_cla32_and10460_y0);
  and_gate and_gate_h_u_cla32_and10461_y0(h_u_cla32_pg_logic23_y0, constant_wire_0, h_u_cla32_and10461_y0);
  and_gate and_gate_h_u_cla32_and10462_y0(h_u_cla32_and10461_y0, h_u_cla32_and10460_y0, h_u_cla32_and10462_y0);
  and_gate and_gate_h_u_cla32_and10463_y0(h_u_cla32_pg_logic24_y0, constant_wire_0, h_u_cla32_and10463_y0);
  and_gate and_gate_h_u_cla32_and10464_y0(h_u_cla32_and10463_y0, h_u_cla32_and10462_y0, h_u_cla32_and10464_y0);
  and_gate and_gate_h_u_cla32_and10465_y0(h_u_cla32_pg_logic25_y0, constant_wire_0, h_u_cla32_and10465_y0);
  and_gate and_gate_h_u_cla32_and10466_y0(h_u_cla32_and10465_y0, h_u_cla32_and10464_y0, h_u_cla32_and10466_y0);
  and_gate and_gate_h_u_cla32_and10467_y0(h_u_cla32_pg_logic26_y0, constant_wire_0, h_u_cla32_and10467_y0);
  and_gate and_gate_h_u_cla32_and10468_y0(h_u_cla32_and10467_y0, h_u_cla32_and10466_y0, h_u_cla32_and10468_y0);
  and_gate and_gate_h_u_cla32_and10469_y0(h_u_cla32_pg_logic27_y0, constant_wire_0, h_u_cla32_and10469_y0);
  and_gate and_gate_h_u_cla32_and10470_y0(h_u_cla32_and10469_y0, h_u_cla32_and10468_y0, h_u_cla32_and10470_y0);
  and_gate and_gate_h_u_cla32_and10471_y0(h_u_cla32_pg_logic28_y0, constant_wire_0, h_u_cla32_and10471_y0);
  and_gate and_gate_h_u_cla32_and10472_y0(h_u_cla32_and10471_y0, h_u_cla32_and10470_y0, h_u_cla32_and10472_y0);
  and_gate and_gate_h_u_cla32_and10473_y0(h_u_cla32_pg_logic29_y0, constant_wire_0, h_u_cla32_and10473_y0);
  and_gate and_gate_h_u_cla32_and10474_y0(h_u_cla32_and10473_y0, h_u_cla32_and10472_y0, h_u_cla32_and10474_y0);
  and_gate and_gate_h_u_cla32_and10475_y0(h_u_cla32_pg_logic30_y0, constant_wire_0, h_u_cla32_and10475_y0);
  and_gate and_gate_h_u_cla32_and10476_y0(h_u_cla32_and10475_y0, h_u_cla32_and10474_y0, h_u_cla32_and10476_y0);
  and_gate and_gate_h_u_cla32_and10477_y0(h_u_cla32_pg_logic31_y0, constant_wire_0, h_u_cla32_and10477_y0);
  and_gate and_gate_h_u_cla32_and10478_y0(h_u_cla32_and10477_y0, h_u_cla32_and10476_y0, h_u_cla32_and10478_y0);
  and_gate and_gate_h_u_cla32_and10479_y0(h_u_cla32_pg_logic1_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10479_y0);
  and_gate and_gate_h_u_cla32_and10480_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10480_y0);
  and_gate and_gate_h_u_cla32_and10481_y0(h_u_cla32_and10480_y0, h_u_cla32_and10479_y0, h_u_cla32_and10481_y0);
  and_gate and_gate_h_u_cla32_and10482_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10482_y0);
  and_gate and_gate_h_u_cla32_and10483_y0(h_u_cla32_and10482_y0, h_u_cla32_and10481_y0, h_u_cla32_and10483_y0);
  and_gate and_gate_h_u_cla32_and10484_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10484_y0);
  and_gate and_gate_h_u_cla32_and10485_y0(h_u_cla32_and10484_y0, h_u_cla32_and10483_y0, h_u_cla32_and10485_y0);
  and_gate and_gate_h_u_cla32_and10486_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10486_y0);
  and_gate and_gate_h_u_cla32_and10487_y0(h_u_cla32_and10486_y0, h_u_cla32_and10485_y0, h_u_cla32_and10487_y0);
  and_gate and_gate_h_u_cla32_and10488_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10488_y0);
  and_gate and_gate_h_u_cla32_and10489_y0(h_u_cla32_and10488_y0, h_u_cla32_and10487_y0, h_u_cla32_and10489_y0);
  and_gate and_gate_h_u_cla32_and10490_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10490_y0);
  and_gate and_gate_h_u_cla32_and10491_y0(h_u_cla32_and10490_y0, h_u_cla32_and10489_y0, h_u_cla32_and10491_y0);
  and_gate and_gate_h_u_cla32_and10492_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10492_y0);
  and_gate and_gate_h_u_cla32_and10493_y0(h_u_cla32_and10492_y0, h_u_cla32_and10491_y0, h_u_cla32_and10493_y0);
  and_gate and_gate_h_u_cla32_and10494_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10494_y0);
  and_gate and_gate_h_u_cla32_and10495_y0(h_u_cla32_and10494_y0, h_u_cla32_and10493_y0, h_u_cla32_and10495_y0);
  and_gate and_gate_h_u_cla32_and10496_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10496_y0);
  and_gate and_gate_h_u_cla32_and10497_y0(h_u_cla32_and10496_y0, h_u_cla32_and10495_y0, h_u_cla32_and10497_y0);
  and_gate and_gate_h_u_cla32_and10498_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10498_y0);
  and_gate and_gate_h_u_cla32_and10499_y0(h_u_cla32_and10498_y0, h_u_cla32_and10497_y0, h_u_cla32_and10499_y0);
  and_gate and_gate_h_u_cla32_and10500_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10500_y0);
  and_gate and_gate_h_u_cla32_and10501_y0(h_u_cla32_and10500_y0, h_u_cla32_and10499_y0, h_u_cla32_and10501_y0);
  and_gate and_gate_h_u_cla32_and10502_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10502_y0);
  and_gate and_gate_h_u_cla32_and10503_y0(h_u_cla32_and10502_y0, h_u_cla32_and10501_y0, h_u_cla32_and10503_y0);
  and_gate and_gate_h_u_cla32_and10504_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10504_y0);
  and_gate and_gate_h_u_cla32_and10505_y0(h_u_cla32_and10504_y0, h_u_cla32_and10503_y0, h_u_cla32_and10505_y0);
  and_gate and_gate_h_u_cla32_and10506_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10506_y0);
  and_gate and_gate_h_u_cla32_and10507_y0(h_u_cla32_and10506_y0, h_u_cla32_and10505_y0, h_u_cla32_and10507_y0);
  and_gate and_gate_h_u_cla32_and10508_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10508_y0);
  and_gate and_gate_h_u_cla32_and10509_y0(h_u_cla32_and10508_y0, h_u_cla32_and10507_y0, h_u_cla32_and10509_y0);
  and_gate and_gate_h_u_cla32_and10510_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10510_y0);
  and_gate and_gate_h_u_cla32_and10511_y0(h_u_cla32_and10510_y0, h_u_cla32_and10509_y0, h_u_cla32_and10511_y0);
  and_gate and_gate_h_u_cla32_and10512_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10512_y0);
  and_gate and_gate_h_u_cla32_and10513_y0(h_u_cla32_and10512_y0, h_u_cla32_and10511_y0, h_u_cla32_and10513_y0);
  and_gate and_gate_h_u_cla32_and10514_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10514_y0);
  and_gate and_gate_h_u_cla32_and10515_y0(h_u_cla32_and10514_y0, h_u_cla32_and10513_y0, h_u_cla32_and10515_y0);
  and_gate and_gate_h_u_cla32_and10516_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10516_y0);
  and_gate and_gate_h_u_cla32_and10517_y0(h_u_cla32_and10516_y0, h_u_cla32_and10515_y0, h_u_cla32_and10517_y0);
  and_gate and_gate_h_u_cla32_and10518_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10518_y0);
  and_gate and_gate_h_u_cla32_and10519_y0(h_u_cla32_and10518_y0, h_u_cla32_and10517_y0, h_u_cla32_and10519_y0);
  and_gate and_gate_h_u_cla32_and10520_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10520_y0);
  and_gate and_gate_h_u_cla32_and10521_y0(h_u_cla32_and10520_y0, h_u_cla32_and10519_y0, h_u_cla32_and10521_y0);
  and_gate and_gate_h_u_cla32_and10522_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10522_y0);
  and_gate and_gate_h_u_cla32_and10523_y0(h_u_cla32_and10522_y0, h_u_cla32_and10521_y0, h_u_cla32_and10523_y0);
  and_gate and_gate_h_u_cla32_and10524_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10524_y0);
  and_gate and_gate_h_u_cla32_and10525_y0(h_u_cla32_and10524_y0, h_u_cla32_and10523_y0, h_u_cla32_and10525_y0);
  and_gate and_gate_h_u_cla32_and10526_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10526_y0);
  and_gate and_gate_h_u_cla32_and10527_y0(h_u_cla32_and10526_y0, h_u_cla32_and10525_y0, h_u_cla32_and10527_y0);
  and_gate and_gate_h_u_cla32_and10528_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10528_y0);
  and_gate and_gate_h_u_cla32_and10529_y0(h_u_cla32_and10528_y0, h_u_cla32_and10527_y0, h_u_cla32_and10529_y0);
  and_gate and_gate_h_u_cla32_and10530_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10530_y0);
  and_gate and_gate_h_u_cla32_and10531_y0(h_u_cla32_and10530_y0, h_u_cla32_and10529_y0, h_u_cla32_and10531_y0);
  and_gate and_gate_h_u_cla32_and10532_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10532_y0);
  and_gate and_gate_h_u_cla32_and10533_y0(h_u_cla32_and10532_y0, h_u_cla32_and10531_y0, h_u_cla32_and10533_y0);
  and_gate and_gate_h_u_cla32_and10534_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10534_y0);
  and_gate and_gate_h_u_cla32_and10535_y0(h_u_cla32_and10534_y0, h_u_cla32_and10533_y0, h_u_cla32_and10535_y0);
  and_gate and_gate_h_u_cla32_and10536_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10536_y0);
  and_gate and_gate_h_u_cla32_and10537_y0(h_u_cla32_and10536_y0, h_u_cla32_and10535_y0, h_u_cla32_and10537_y0);
  and_gate and_gate_h_u_cla32_and10538_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic0_y1, h_u_cla32_and10538_y0);
  and_gate and_gate_h_u_cla32_and10539_y0(h_u_cla32_and10538_y0, h_u_cla32_and10537_y0, h_u_cla32_and10539_y0);
  and_gate and_gate_h_u_cla32_and10540_y0(h_u_cla32_pg_logic2_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10540_y0);
  and_gate and_gate_h_u_cla32_and10541_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10541_y0);
  and_gate and_gate_h_u_cla32_and10542_y0(h_u_cla32_and10541_y0, h_u_cla32_and10540_y0, h_u_cla32_and10542_y0);
  and_gate and_gate_h_u_cla32_and10543_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10543_y0);
  and_gate and_gate_h_u_cla32_and10544_y0(h_u_cla32_and10543_y0, h_u_cla32_and10542_y0, h_u_cla32_and10544_y0);
  and_gate and_gate_h_u_cla32_and10545_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10545_y0);
  and_gate and_gate_h_u_cla32_and10546_y0(h_u_cla32_and10545_y0, h_u_cla32_and10544_y0, h_u_cla32_and10546_y0);
  and_gate and_gate_h_u_cla32_and10547_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10547_y0);
  and_gate and_gate_h_u_cla32_and10548_y0(h_u_cla32_and10547_y0, h_u_cla32_and10546_y0, h_u_cla32_and10548_y0);
  and_gate and_gate_h_u_cla32_and10549_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10549_y0);
  and_gate and_gate_h_u_cla32_and10550_y0(h_u_cla32_and10549_y0, h_u_cla32_and10548_y0, h_u_cla32_and10550_y0);
  and_gate and_gate_h_u_cla32_and10551_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10551_y0);
  and_gate and_gate_h_u_cla32_and10552_y0(h_u_cla32_and10551_y0, h_u_cla32_and10550_y0, h_u_cla32_and10552_y0);
  and_gate and_gate_h_u_cla32_and10553_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10553_y0);
  and_gate and_gate_h_u_cla32_and10554_y0(h_u_cla32_and10553_y0, h_u_cla32_and10552_y0, h_u_cla32_and10554_y0);
  and_gate and_gate_h_u_cla32_and10555_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10555_y0);
  and_gate and_gate_h_u_cla32_and10556_y0(h_u_cla32_and10555_y0, h_u_cla32_and10554_y0, h_u_cla32_and10556_y0);
  and_gate and_gate_h_u_cla32_and10557_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10557_y0);
  and_gate and_gate_h_u_cla32_and10558_y0(h_u_cla32_and10557_y0, h_u_cla32_and10556_y0, h_u_cla32_and10558_y0);
  and_gate and_gate_h_u_cla32_and10559_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10559_y0);
  and_gate and_gate_h_u_cla32_and10560_y0(h_u_cla32_and10559_y0, h_u_cla32_and10558_y0, h_u_cla32_and10560_y0);
  and_gate and_gate_h_u_cla32_and10561_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10561_y0);
  and_gate and_gate_h_u_cla32_and10562_y0(h_u_cla32_and10561_y0, h_u_cla32_and10560_y0, h_u_cla32_and10562_y0);
  and_gate and_gate_h_u_cla32_and10563_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10563_y0);
  and_gate and_gate_h_u_cla32_and10564_y0(h_u_cla32_and10563_y0, h_u_cla32_and10562_y0, h_u_cla32_and10564_y0);
  and_gate and_gate_h_u_cla32_and10565_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10565_y0);
  and_gate and_gate_h_u_cla32_and10566_y0(h_u_cla32_and10565_y0, h_u_cla32_and10564_y0, h_u_cla32_and10566_y0);
  and_gate and_gate_h_u_cla32_and10567_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10567_y0);
  and_gate and_gate_h_u_cla32_and10568_y0(h_u_cla32_and10567_y0, h_u_cla32_and10566_y0, h_u_cla32_and10568_y0);
  and_gate and_gate_h_u_cla32_and10569_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10569_y0);
  and_gate and_gate_h_u_cla32_and10570_y0(h_u_cla32_and10569_y0, h_u_cla32_and10568_y0, h_u_cla32_and10570_y0);
  and_gate and_gate_h_u_cla32_and10571_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10571_y0);
  and_gate and_gate_h_u_cla32_and10572_y0(h_u_cla32_and10571_y0, h_u_cla32_and10570_y0, h_u_cla32_and10572_y0);
  and_gate and_gate_h_u_cla32_and10573_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10573_y0);
  and_gate and_gate_h_u_cla32_and10574_y0(h_u_cla32_and10573_y0, h_u_cla32_and10572_y0, h_u_cla32_and10574_y0);
  and_gate and_gate_h_u_cla32_and10575_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10575_y0);
  and_gate and_gate_h_u_cla32_and10576_y0(h_u_cla32_and10575_y0, h_u_cla32_and10574_y0, h_u_cla32_and10576_y0);
  and_gate and_gate_h_u_cla32_and10577_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10577_y0);
  and_gate and_gate_h_u_cla32_and10578_y0(h_u_cla32_and10577_y0, h_u_cla32_and10576_y0, h_u_cla32_and10578_y0);
  and_gate and_gate_h_u_cla32_and10579_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10579_y0);
  and_gate and_gate_h_u_cla32_and10580_y0(h_u_cla32_and10579_y0, h_u_cla32_and10578_y0, h_u_cla32_and10580_y0);
  and_gate and_gate_h_u_cla32_and10581_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10581_y0);
  and_gate and_gate_h_u_cla32_and10582_y0(h_u_cla32_and10581_y0, h_u_cla32_and10580_y0, h_u_cla32_and10582_y0);
  and_gate and_gate_h_u_cla32_and10583_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10583_y0);
  and_gate and_gate_h_u_cla32_and10584_y0(h_u_cla32_and10583_y0, h_u_cla32_and10582_y0, h_u_cla32_and10584_y0);
  and_gate and_gate_h_u_cla32_and10585_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10585_y0);
  and_gate and_gate_h_u_cla32_and10586_y0(h_u_cla32_and10585_y0, h_u_cla32_and10584_y0, h_u_cla32_and10586_y0);
  and_gate and_gate_h_u_cla32_and10587_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10587_y0);
  and_gate and_gate_h_u_cla32_and10588_y0(h_u_cla32_and10587_y0, h_u_cla32_and10586_y0, h_u_cla32_and10588_y0);
  and_gate and_gate_h_u_cla32_and10589_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10589_y0);
  and_gate and_gate_h_u_cla32_and10590_y0(h_u_cla32_and10589_y0, h_u_cla32_and10588_y0, h_u_cla32_and10590_y0);
  and_gate and_gate_h_u_cla32_and10591_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10591_y0);
  and_gate and_gate_h_u_cla32_and10592_y0(h_u_cla32_and10591_y0, h_u_cla32_and10590_y0, h_u_cla32_and10592_y0);
  and_gate and_gate_h_u_cla32_and10593_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10593_y0);
  and_gate and_gate_h_u_cla32_and10594_y0(h_u_cla32_and10593_y0, h_u_cla32_and10592_y0, h_u_cla32_and10594_y0);
  and_gate and_gate_h_u_cla32_and10595_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10595_y0);
  and_gate and_gate_h_u_cla32_and10596_y0(h_u_cla32_and10595_y0, h_u_cla32_and10594_y0, h_u_cla32_and10596_y0);
  and_gate and_gate_h_u_cla32_and10597_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic1_y1, h_u_cla32_and10597_y0);
  and_gate and_gate_h_u_cla32_and10598_y0(h_u_cla32_and10597_y0, h_u_cla32_and10596_y0, h_u_cla32_and10598_y0);
  and_gate and_gate_h_u_cla32_and10599_y0(h_u_cla32_pg_logic3_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10599_y0);
  and_gate and_gate_h_u_cla32_and10600_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10600_y0);
  and_gate and_gate_h_u_cla32_and10601_y0(h_u_cla32_and10600_y0, h_u_cla32_and10599_y0, h_u_cla32_and10601_y0);
  and_gate and_gate_h_u_cla32_and10602_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10602_y0);
  and_gate and_gate_h_u_cla32_and10603_y0(h_u_cla32_and10602_y0, h_u_cla32_and10601_y0, h_u_cla32_and10603_y0);
  and_gate and_gate_h_u_cla32_and10604_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10604_y0);
  and_gate and_gate_h_u_cla32_and10605_y0(h_u_cla32_and10604_y0, h_u_cla32_and10603_y0, h_u_cla32_and10605_y0);
  and_gate and_gate_h_u_cla32_and10606_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10606_y0);
  and_gate and_gate_h_u_cla32_and10607_y0(h_u_cla32_and10606_y0, h_u_cla32_and10605_y0, h_u_cla32_and10607_y0);
  and_gate and_gate_h_u_cla32_and10608_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10608_y0);
  and_gate and_gate_h_u_cla32_and10609_y0(h_u_cla32_and10608_y0, h_u_cla32_and10607_y0, h_u_cla32_and10609_y0);
  and_gate and_gate_h_u_cla32_and10610_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10610_y0);
  and_gate and_gate_h_u_cla32_and10611_y0(h_u_cla32_and10610_y0, h_u_cla32_and10609_y0, h_u_cla32_and10611_y0);
  and_gate and_gate_h_u_cla32_and10612_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10612_y0);
  and_gate and_gate_h_u_cla32_and10613_y0(h_u_cla32_and10612_y0, h_u_cla32_and10611_y0, h_u_cla32_and10613_y0);
  and_gate and_gate_h_u_cla32_and10614_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10614_y0);
  and_gate and_gate_h_u_cla32_and10615_y0(h_u_cla32_and10614_y0, h_u_cla32_and10613_y0, h_u_cla32_and10615_y0);
  and_gate and_gate_h_u_cla32_and10616_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10616_y0);
  and_gate and_gate_h_u_cla32_and10617_y0(h_u_cla32_and10616_y0, h_u_cla32_and10615_y0, h_u_cla32_and10617_y0);
  and_gate and_gate_h_u_cla32_and10618_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10618_y0);
  and_gate and_gate_h_u_cla32_and10619_y0(h_u_cla32_and10618_y0, h_u_cla32_and10617_y0, h_u_cla32_and10619_y0);
  and_gate and_gate_h_u_cla32_and10620_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10620_y0);
  and_gate and_gate_h_u_cla32_and10621_y0(h_u_cla32_and10620_y0, h_u_cla32_and10619_y0, h_u_cla32_and10621_y0);
  and_gate and_gate_h_u_cla32_and10622_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10622_y0);
  and_gate and_gate_h_u_cla32_and10623_y0(h_u_cla32_and10622_y0, h_u_cla32_and10621_y0, h_u_cla32_and10623_y0);
  and_gate and_gate_h_u_cla32_and10624_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10624_y0);
  and_gate and_gate_h_u_cla32_and10625_y0(h_u_cla32_and10624_y0, h_u_cla32_and10623_y0, h_u_cla32_and10625_y0);
  and_gate and_gate_h_u_cla32_and10626_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10626_y0);
  and_gate and_gate_h_u_cla32_and10627_y0(h_u_cla32_and10626_y0, h_u_cla32_and10625_y0, h_u_cla32_and10627_y0);
  and_gate and_gate_h_u_cla32_and10628_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10628_y0);
  and_gate and_gate_h_u_cla32_and10629_y0(h_u_cla32_and10628_y0, h_u_cla32_and10627_y0, h_u_cla32_and10629_y0);
  and_gate and_gate_h_u_cla32_and10630_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10630_y0);
  and_gate and_gate_h_u_cla32_and10631_y0(h_u_cla32_and10630_y0, h_u_cla32_and10629_y0, h_u_cla32_and10631_y0);
  and_gate and_gate_h_u_cla32_and10632_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10632_y0);
  and_gate and_gate_h_u_cla32_and10633_y0(h_u_cla32_and10632_y0, h_u_cla32_and10631_y0, h_u_cla32_and10633_y0);
  and_gate and_gate_h_u_cla32_and10634_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10634_y0);
  and_gate and_gate_h_u_cla32_and10635_y0(h_u_cla32_and10634_y0, h_u_cla32_and10633_y0, h_u_cla32_and10635_y0);
  and_gate and_gate_h_u_cla32_and10636_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10636_y0);
  and_gate and_gate_h_u_cla32_and10637_y0(h_u_cla32_and10636_y0, h_u_cla32_and10635_y0, h_u_cla32_and10637_y0);
  and_gate and_gate_h_u_cla32_and10638_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10638_y0);
  and_gate and_gate_h_u_cla32_and10639_y0(h_u_cla32_and10638_y0, h_u_cla32_and10637_y0, h_u_cla32_and10639_y0);
  and_gate and_gate_h_u_cla32_and10640_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10640_y0);
  and_gate and_gate_h_u_cla32_and10641_y0(h_u_cla32_and10640_y0, h_u_cla32_and10639_y0, h_u_cla32_and10641_y0);
  and_gate and_gate_h_u_cla32_and10642_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10642_y0);
  and_gate and_gate_h_u_cla32_and10643_y0(h_u_cla32_and10642_y0, h_u_cla32_and10641_y0, h_u_cla32_and10643_y0);
  and_gate and_gate_h_u_cla32_and10644_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10644_y0);
  and_gate and_gate_h_u_cla32_and10645_y0(h_u_cla32_and10644_y0, h_u_cla32_and10643_y0, h_u_cla32_and10645_y0);
  and_gate and_gate_h_u_cla32_and10646_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10646_y0);
  and_gate and_gate_h_u_cla32_and10647_y0(h_u_cla32_and10646_y0, h_u_cla32_and10645_y0, h_u_cla32_and10647_y0);
  and_gate and_gate_h_u_cla32_and10648_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10648_y0);
  and_gate and_gate_h_u_cla32_and10649_y0(h_u_cla32_and10648_y0, h_u_cla32_and10647_y0, h_u_cla32_and10649_y0);
  and_gate and_gate_h_u_cla32_and10650_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10650_y0);
  and_gate and_gate_h_u_cla32_and10651_y0(h_u_cla32_and10650_y0, h_u_cla32_and10649_y0, h_u_cla32_and10651_y0);
  and_gate and_gate_h_u_cla32_and10652_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10652_y0);
  and_gate and_gate_h_u_cla32_and10653_y0(h_u_cla32_and10652_y0, h_u_cla32_and10651_y0, h_u_cla32_and10653_y0);
  and_gate and_gate_h_u_cla32_and10654_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic2_y1, h_u_cla32_and10654_y0);
  and_gate and_gate_h_u_cla32_and10655_y0(h_u_cla32_and10654_y0, h_u_cla32_and10653_y0, h_u_cla32_and10655_y0);
  and_gate and_gate_h_u_cla32_and10656_y0(h_u_cla32_pg_logic4_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10656_y0);
  and_gate and_gate_h_u_cla32_and10657_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10657_y0);
  and_gate and_gate_h_u_cla32_and10658_y0(h_u_cla32_and10657_y0, h_u_cla32_and10656_y0, h_u_cla32_and10658_y0);
  and_gate and_gate_h_u_cla32_and10659_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10659_y0);
  and_gate and_gate_h_u_cla32_and10660_y0(h_u_cla32_and10659_y0, h_u_cla32_and10658_y0, h_u_cla32_and10660_y0);
  and_gate and_gate_h_u_cla32_and10661_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10661_y0);
  and_gate and_gate_h_u_cla32_and10662_y0(h_u_cla32_and10661_y0, h_u_cla32_and10660_y0, h_u_cla32_and10662_y0);
  and_gate and_gate_h_u_cla32_and10663_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10663_y0);
  and_gate and_gate_h_u_cla32_and10664_y0(h_u_cla32_and10663_y0, h_u_cla32_and10662_y0, h_u_cla32_and10664_y0);
  and_gate and_gate_h_u_cla32_and10665_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10665_y0);
  and_gate and_gate_h_u_cla32_and10666_y0(h_u_cla32_and10665_y0, h_u_cla32_and10664_y0, h_u_cla32_and10666_y0);
  and_gate and_gate_h_u_cla32_and10667_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10667_y0);
  and_gate and_gate_h_u_cla32_and10668_y0(h_u_cla32_and10667_y0, h_u_cla32_and10666_y0, h_u_cla32_and10668_y0);
  and_gate and_gate_h_u_cla32_and10669_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10669_y0);
  and_gate and_gate_h_u_cla32_and10670_y0(h_u_cla32_and10669_y0, h_u_cla32_and10668_y0, h_u_cla32_and10670_y0);
  and_gate and_gate_h_u_cla32_and10671_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10671_y0);
  and_gate and_gate_h_u_cla32_and10672_y0(h_u_cla32_and10671_y0, h_u_cla32_and10670_y0, h_u_cla32_and10672_y0);
  and_gate and_gate_h_u_cla32_and10673_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10673_y0);
  and_gate and_gate_h_u_cla32_and10674_y0(h_u_cla32_and10673_y0, h_u_cla32_and10672_y0, h_u_cla32_and10674_y0);
  and_gate and_gate_h_u_cla32_and10675_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10675_y0);
  and_gate and_gate_h_u_cla32_and10676_y0(h_u_cla32_and10675_y0, h_u_cla32_and10674_y0, h_u_cla32_and10676_y0);
  and_gate and_gate_h_u_cla32_and10677_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10677_y0);
  and_gate and_gate_h_u_cla32_and10678_y0(h_u_cla32_and10677_y0, h_u_cla32_and10676_y0, h_u_cla32_and10678_y0);
  and_gate and_gate_h_u_cla32_and10679_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10679_y0);
  and_gate and_gate_h_u_cla32_and10680_y0(h_u_cla32_and10679_y0, h_u_cla32_and10678_y0, h_u_cla32_and10680_y0);
  and_gate and_gate_h_u_cla32_and10681_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10681_y0);
  and_gate and_gate_h_u_cla32_and10682_y0(h_u_cla32_and10681_y0, h_u_cla32_and10680_y0, h_u_cla32_and10682_y0);
  and_gate and_gate_h_u_cla32_and10683_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10683_y0);
  and_gate and_gate_h_u_cla32_and10684_y0(h_u_cla32_and10683_y0, h_u_cla32_and10682_y0, h_u_cla32_and10684_y0);
  and_gate and_gate_h_u_cla32_and10685_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10685_y0);
  and_gate and_gate_h_u_cla32_and10686_y0(h_u_cla32_and10685_y0, h_u_cla32_and10684_y0, h_u_cla32_and10686_y0);
  and_gate and_gate_h_u_cla32_and10687_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10687_y0);
  and_gate and_gate_h_u_cla32_and10688_y0(h_u_cla32_and10687_y0, h_u_cla32_and10686_y0, h_u_cla32_and10688_y0);
  and_gate and_gate_h_u_cla32_and10689_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10689_y0);
  and_gate and_gate_h_u_cla32_and10690_y0(h_u_cla32_and10689_y0, h_u_cla32_and10688_y0, h_u_cla32_and10690_y0);
  and_gate and_gate_h_u_cla32_and10691_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10691_y0);
  and_gate and_gate_h_u_cla32_and10692_y0(h_u_cla32_and10691_y0, h_u_cla32_and10690_y0, h_u_cla32_and10692_y0);
  and_gate and_gate_h_u_cla32_and10693_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10693_y0);
  and_gate and_gate_h_u_cla32_and10694_y0(h_u_cla32_and10693_y0, h_u_cla32_and10692_y0, h_u_cla32_and10694_y0);
  and_gate and_gate_h_u_cla32_and10695_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10695_y0);
  and_gate and_gate_h_u_cla32_and10696_y0(h_u_cla32_and10695_y0, h_u_cla32_and10694_y0, h_u_cla32_and10696_y0);
  and_gate and_gate_h_u_cla32_and10697_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10697_y0);
  and_gate and_gate_h_u_cla32_and10698_y0(h_u_cla32_and10697_y0, h_u_cla32_and10696_y0, h_u_cla32_and10698_y0);
  and_gate and_gate_h_u_cla32_and10699_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10699_y0);
  and_gate and_gate_h_u_cla32_and10700_y0(h_u_cla32_and10699_y0, h_u_cla32_and10698_y0, h_u_cla32_and10700_y0);
  and_gate and_gate_h_u_cla32_and10701_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10701_y0);
  and_gate and_gate_h_u_cla32_and10702_y0(h_u_cla32_and10701_y0, h_u_cla32_and10700_y0, h_u_cla32_and10702_y0);
  and_gate and_gate_h_u_cla32_and10703_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10703_y0);
  and_gate and_gate_h_u_cla32_and10704_y0(h_u_cla32_and10703_y0, h_u_cla32_and10702_y0, h_u_cla32_and10704_y0);
  and_gate and_gate_h_u_cla32_and10705_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10705_y0);
  and_gate and_gate_h_u_cla32_and10706_y0(h_u_cla32_and10705_y0, h_u_cla32_and10704_y0, h_u_cla32_and10706_y0);
  and_gate and_gate_h_u_cla32_and10707_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10707_y0);
  and_gate and_gate_h_u_cla32_and10708_y0(h_u_cla32_and10707_y0, h_u_cla32_and10706_y0, h_u_cla32_and10708_y0);
  and_gate and_gate_h_u_cla32_and10709_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic3_y1, h_u_cla32_and10709_y0);
  and_gate and_gate_h_u_cla32_and10710_y0(h_u_cla32_and10709_y0, h_u_cla32_and10708_y0, h_u_cla32_and10710_y0);
  and_gate and_gate_h_u_cla32_and10711_y0(h_u_cla32_pg_logic5_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10711_y0);
  and_gate and_gate_h_u_cla32_and10712_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10712_y0);
  and_gate and_gate_h_u_cla32_and10713_y0(h_u_cla32_and10712_y0, h_u_cla32_and10711_y0, h_u_cla32_and10713_y0);
  and_gate and_gate_h_u_cla32_and10714_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10714_y0);
  and_gate and_gate_h_u_cla32_and10715_y0(h_u_cla32_and10714_y0, h_u_cla32_and10713_y0, h_u_cla32_and10715_y0);
  and_gate and_gate_h_u_cla32_and10716_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10716_y0);
  and_gate and_gate_h_u_cla32_and10717_y0(h_u_cla32_and10716_y0, h_u_cla32_and10715_y0, h_u_cla32_and10717_y0);
  and_gate and_gate_h_u_cla32_and10718_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10718_y0);
  and_gate and_gate_h_u_cla32_and10719_y0(h_u_cla32_and10718_y0, h_u_cla32_and10717_y0, h_u_cla32_and10719_y0);
  and_gate and_gate_h_u_cla32_and10720_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10720_y0);
  and_gate and_gate_h_u_cla32_and10721_y0(h_u_cla32_and10720_y0, h_u_cla32_and10719_y0, h_u_cla32_and10721_y0);
  and_gate and_gate_h_u_cla32_and10722_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10722_y0);
  and_gate and_gate_h_u_cla32_and10723_y0(h_u_cla32_and10722_y0, h_u_cla32_and10721_y0, h_u_cla32_and10723_y0);
  and_gate and_gate_h_u_cla32_and10724_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10724_y0);
  and_gate and_gate_h_u_cla32_and10725_y0(h_u_cla32_and10724_y0, h_u_cla32_and10723_y0, h_u_cla32_and10725_y0);
  and_gate and_gate_h_u_cla32_and10726_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10726_y0);
  and_gate and_gate_h_u_cla32_and10727_y0(h_u_cla32_and10726_y0, h_u_cla32_and10725_y0, h_u_cla32_and10727_y0);
  and_gate and_gate_h_u_cla32_and10728_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10728_y0);
  and_gate and_gate_h_u_cla32_and10729_y0(h_u_cla32_and10728_y0, h_u_cla32_and10727_y0, h_u_cla32_and10729_y0);
  and_gate and_gate_h_u_cla32_and10730_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10730_y0);
  and_gate and_gate_h_u_cla32_and10731_y0(h_u_cla32_and10730_y0, h_u_cla32_and10729_y0, h_u_cla32_and10731_y0);
  and_gate and_gate_h_u_cla32_and10732_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10732_y0);
  and_gate and_gate_h_u_cla32_and10733_y0(h_u_cla32_and10732_y0, h_u_cla32_and10731_y0, h_u_cla32_and10733_y0);
  and_gate and_gate_h_u_cla32_and10734_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10734_y0);
  and_gate and_gate_h_u_cla32_and10735_y0(h_u_cla32_and10734_y0, h_u_cla32_and10733_y0, h_u_cla32_and10735_y0);
  and_gate and_gate_h_u_cla32_and10736_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10736_y0);
  and_gate and_gate_h_u_cla32_and10737_y0(h_u_cla32_and10736_y0, h_u_cla32_and10735_y0, h_u_cla32_and10737_y0);
  and_gate and_gate_h_u_cla32_and10738_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10738_y0);
  and_gate and_gate_h_u_cla32_and10739_y0(h_u_cla32_and10738_y0, h_u_cla32_and10737_y0, h_u_cla32_and10739_y0);
  and_gate and_gate_h_u_cla32_and10740_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10740_y0);
  and_gate and_gate_h_u_cla32_and10741_y0(h_u_cla32_and10740_y0, h_u_cla32_and10739_y0, h_u_cla32_and10741_y0);
  and_gate and_gate_h_u_cla32_and10742_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10742_y0);
  and_gate and_gate_h_u_cla32_and10743_y0(h_u_cla32_and10742_y0, h_u_cla32_and10741_y0, h_u_cla32_and10743_y0);
  and_gate and_gate_h_u_cla32_and10744_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10744_y0);
  and_gate and_gate_h_u_cla32_and10745_y0(h_u_cla32_and10744_y0, h_u_cla32_and10743_y0, h_u_cla32_and10745_y0);
  and_gate and_gate_h_u_cla32_and10746_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10746_y0);
  and_gate and_gate_h_u_cla32_and10747_y0(h_u_cla32_and10746_y0, h_u_cla32_and10745_y0, h_u_cla32_and10747_y0);
  and_gate and_gate_h_u_cla32_and10748_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10748_y0);
  and_gate and_gate_h_u_cla32_and10749_y0(h_u_cla32_and10748_y0, h_u_cla32_and10747_y0, h_u_cla32_and10749_y0);
  and_gate and_gate_h_u_cla32_and10750_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10750_y0);
  and_gate and_gate_h_u_cla32_and10751_y0(h_u_cla32_and10750_y0, h_u_cla32_and10749_y0, h_u_cla32_and10751_y0);
  and_gate and_gate_h_u_cla32_and10752_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10752_y0);
  and_gate and_gate_h_u_cla32_and10753_y0(h_u_cla32_and10752_y0, h_u_cla32_and10751_y0, h_u_cla32_and10753_y0);
  and_gate and_gate_h_u_cla32_and10754_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10754_y0);
  and_gate and_gate_h_u_cla32_and10755_y0(h_u_cla32_and10754_y0, h_u_cla32_and10753_y0, h_u_cla32_and10755_y0);
  and_gate and_gate_h_u_cla32_and10756_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10756_y0);
  and_gate and_gate_h_u_cla32_and10757_y0(h_u_cla32_and10756_y0, h_u_cla32_and10755_y0, h_u_cla32_and10757_y0);
  and_gate and_gate_h_u_cla32_and10758_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10758_y0);
  and_gate and_gate_h_u_cla32_and10759_y0(h_u_cla32_and10758_y0, h_u_cla32_and10757_y0, h_u_cla32_and10759_y0);
  and_gate and_gate_h_u_cla32_and10760_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10760_y0);
  and_gate and_gate_h_u_cla32_and10761_y0(h_u_cla32_and10760_y0, h_u_cla32_and10759_y0, h_u_cla32_and10761_y0);
  and_gate and_gate_h_u_cla32_and10762_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic4_y1, h_u_cla32_and10762_y0);
  and_gate and_gate_h_u_cla32_and10763_y0(h_u_cla32_and10762_y0, h_u_cla32_and10761_y0, h_u_cla32_and10763_y0);
  and_gate and_gate_h_u_cla32_and10764_y0(h_u_cla32_pg_logic6_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10764_y0);
  and_gate and_gate_h_u_cla32_and10765_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10765_y0);
  and_gate and_gate_h_u_cla32_and10766_y0(h_u_cla32_and10765_y0, h_u_cla32_and10764_y0, h_u_cla32_and10766_y0);
  and_gate and_gate_h_u_cla32_and10767_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10767_y0);
  and_gate and_gate_h_u_cla32_and10768_y0(h_u_cla32_and10767_y0, h_u_cla32_and10766_y0, h_u_cla32_and10768_y0);
  and_gate and_gate_h_u_cla32_and10769_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10769_y0);
  and_gate and_gate_h_u_cla32_and10770_y0(h_u_cla32_and10769_y0, h_u_cla32_and10768_y0, h_u_cla32_and10770_y0);
  and_gate and_gate_h_u_cla32_and10771_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10771_y0);
  and_gate and_gate_h_u_cla32_and10772_y0(h_u_cla32_and10771_y0, h_u_cla32_and10770_y0, h_u_cla32_and10772_y0);
  and_gate and_gate_h_u_cla32_and10773_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10773_y0);
  and_gate and_gate_h_u_cla32_and10774_y0(h_u_cla32_and10773_y0, h_u_cla32_and10772_y0, h_u_cla32_and10774_y0);
  and_gate and_gate_h_u_cla32_and10775_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10775_y0);
  and_gate and_gate_h_u_cla32_and10776_y0(h_u_cla32_and10775_y0, h_u_cla32_and10774_y0, h_u_cla32_and10776_y0);
  and_gate and_gate_h_u_cla32_and10777_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10777_y0);
  and_gate and_gate_h_u_cla32_and10778_y0(h_u_cla32_and10777_y0, h_u_cla32_and10776_y0, h_u_cla32_and10778_y0);
  and_gate and_gate_h_u_cla32_and10779_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10779_y0);
  and_gate and_gate_h_u_cla32_and10780_y0(h_u_cla32_and10779_y0, h_u_cla32_and10778_y0, h_u_cla32_and10780_y0);
  and_gate and_gate_h_u_cla32_and10781_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10781_y0);
  and_gate and_gate_h_u_cla32_and10782_y0(h_u_cla32_and10781_y0, h_u_cla32_and10780_y0, h_u_cla32_and10782_y0);
  and_gate and_gate_h_u_cla32_and10783_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10783_y0);
  and_gate and_gate_h_u_cla32_and10784_y0(h_u_cla32_and10783_y0, h_u_cla32_and10782_y0, h_u_cla32_and10784_y0);
  and_gate and_gate_h_u_cla32_and10785_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10785_y0);
  and_gate and_gate_h_u_cla32_and10786_y0(h_u_cla32_and10785_y0, h_u_cla32_and10784_y0, h_u_cla32_and10786_y0);
  and_gate and_gate_h_u_cla32_and10787_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10787_y0);
  and_gate and_gate_h_u_cla32_and10788_y0(h_u_cla32_and10787_y0, h_u_cla32_and10786_y0, h_u_cla32_and10788_y0);
  and_gate and_gate_h_u_cla32_and10789_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10789_y0);
  and_gate and_gate_h_u_cla32_and10790_y0(h_u_cla32_and10789_y0, h_u_cla32_and10788_y0, h_u_cla32_and10790_y0);
  and_gate and_gate_h_u_cla32_and10791_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10791_y0);
  and_gate and_gate_h_u_cla32_and10792_y0(h_u_cla32_and10791_y0, h_u_cla32_and10790_y0, h_u_cla32_and10792_y0);
  and_gate and_gate_h_u_cla32_and10793_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10793_y0);
  and_gate and_gate_h_u_cla32_and10794_y0(h_u_cla32_and10793_y0, h_u_cla32_and10792_y0, h_u_cla32_and10794_y0);
  and_gate and_gate_h_u_cla32_and10795_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10795_y0);
  and_gate and_gate_h_u_cla32_and10796_y0(h_u_cla32_and10795_y0, h_u_cla32_and10794_y0, h_u_cla32_and10796_y0);
  and_gate and_gate_h_u_cla32_and10797_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10797_y0);
  and_gate and_gate_h_u_cla32_and10798_y0(h_u_cla32_and10797_y0, h_u_cla32_and10796_y0, h_u_cla32_and10798_y0);
  and_gate and_gate_h_u_cla32_and10799_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10799_y0);
  and_gate and_gate_h_u_cla32_and10800_y0(h_u_cla32_and10799_y0, h_u_cla32_and10798_y0, h_u_cla32_and10800_y0);
  and_gate and_gate_h_u_cla32_and10801_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10801_y0);
  and_gate and_gate_h_u_cla32_and10802_y0(h_u_cla32_and10801_y0, h_u_cla32_and10800_y0, h_u_cla32_and10802_y0);
  and_gate and_gate_h_u_cla32_and10803_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10803_y0);
  and_gate and_gate_h_u_cla32_and10804_y0(h_u_cla32_and10803_y0, h_u_cla32_and10802_y0, h_u_cla32_and10804_y0);
  and_gate and_gate_h_u_cla32_and10805_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10805_y0);
  and_gate and_gate_h_u_cla32_and10806_y0(h_u_cla32_and10805_y0, h_u_cla32_and10804_y0, h_u_cla32_and10806_y0);
  and_gate and_gate_h_u_cla32_and10807_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10807_y0);
  and_gate and_gate_h_u_cla32_and10808_y0(h_u_cla32_and10807_y0, h_u_cla32_and10806_y0, h_u_cla32_and10808_y0);
  and_gate and_gate_h_u_cla32_and10809_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10809_y0);
  and_gate and_gate_h_u_cla32_and10810_y0(h_u_cla32_and10809_y0, h_u_cla32_and10808_y0, h_u_cla32_and10810_y0);
  and_gate and_gate_h_u_cla32_and10811_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10811_y0);
  and_gate and_gate_h_u_cla32_and10812_y0(h_u_cla32_and10811_y0, h_u_cla32_and10810_y0, h_u_cla32_and10812_y0);
  and_gate and_gate_h_u_cla32_and10813_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic5_y1, h_u_cla32_and10813_y0);
  and_gate and_gate_h_u_cla32_and10814_y0(h_u_cla32_and10813_y0, h_u_cla32_and10812_y0, h_u_cla32_and10814_y0);
  and_gate and_gate_h_u_cla32_and10815_y0(h_u_cla32_pg_logic7_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10815_y0);
  and_gate and_gate_h_u_cla32_and10816_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10816_y0);
  and_gate and_gate_h_u_cla32_and10817_y0(h_u_cla32_and10816_y0, h_u_cla32_and10815_y0, h_u_cla32_and10817_y0);
  and_gate and_gate_h_u_cla32_and10818_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10818_y0);
  and_gate and_gate_h_u_cla32_and10819_y0(h_u_cla32_and10818_y0, h_u_cla32_and10817_y0, h_u_cla32_and10819_y0);
  and_gate and_gate_h_u_cla32_and10820_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10820_y0);
  and_gate and_gate_h_u_cla32_and10821_y0(h_u_cla32_and10820_y0, h_u_cla32_and10819_y0, h_u_cla32_and10821_y0);
  and_gate and_gate_h_u_cla32_and10822_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10822_y0);
  and_gate and_gate_h_u_cla32_and10823_y0(h_u_cla32_and10822_y0, h_u_cla32_and10821_y0, h_u_cla32_and10823_y0);
  and_gate and_gate_h_u_cla32_and10824_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10824_y0);
  and_gate and_gate_h_u_cla32_and10825_y0(h_u_cla32_and10824_y0, h_u_cla32_and10823_y0, h_u_cla32_and10825_y0);
  and_gate and_gate_h_u_cla32_and10826_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10826_y0);
  and_gate and_gate_h_u_cla32_and10827_y0(h_u_cla32_and10826_y0, h_u_cla32_and10825_y0, h_u_cla32_and10827_y0);
  and_gate and_gate_h_u_cla32_and10828_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10828_y0);
  and_gate and_gate_h_u_cla32_and10829_y0(h_u_cla32_and10828_y0, h_u_cla32_and10827_y0, h_u_cla32_and10829_y0);
  and_gate and_gate_h_u_cla32_and10830_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10830_y0);
  and_gate and_gate_h_u_cla32_and10831_y0(h_u_cla32_and10830_y0, h_u_cla32_and10829_y0, h_u_cla32_and10831_y0);
  and_gate and_gate_h_u_cla32_and10832_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10832_y0);
  and_gate and_gate_h_u_cla32_and10833_y0(h_u_cla32_and10832_y0, h_u_cla32_and10831_y0, h_u_cla32_and10833_y0);
  and_gate and_gate_h_u_cla32_and10834_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10834_y0);
  and_gate and_gate_h_u_cla32_and10835_y0(h_u_cla32_and10834_y0, h_u_cla32_and10833_y0, h_u_cla32_and10835_y0);
  and_gate and_gate_h_u_cla32_and10836_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10836_y0);
  and_gate and_gate_h_u_cla32_and10837_y0(h_u_cla32_and10836_y0, h_u_cla32_and10835_y0, h_u_cla32_and10837_y0);
  and_gate and_gate_h_u_cla32_and10838_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10838_y0);
  and_gate and_gate_h_u_cla32_and10839_y0(h_u_cla32_and10838_y0, h_u_cla32_and10837_y0, h_u_cla32_and10839_y0);
  and_gate and_gate_h_u_cla32_and10840_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10840_y0);
  and_gate and_gate_h_u_cla32_and10841_y0(h_u_cla32_and10840_y0, h_u_cla32_and10839_y0, h_u_cla32_and10841_y0);
  and_gate and_gate_h_u_cla32_and10842_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10842_y0);
  and_gate and_gate_h_u_cla32_and10843_y0(h_u_cla32_and10842_y0, h_u_cla32_and10841_y0, h_u_cla32_and10843_y0);
  and_gate and_gate_h_u_cla32_and10844_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10844_y0);
  and_gate and_gate_h_u_cla32_and10845_y0(h_u_cla32_and10844_y0, h_u_cla32_and10843_y0, h_u_cla32_and10845_y0);
  and_gate and_gate_h_u_cla32_and10846_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10846_y0);
  and_gate and_gate_h_u_cla32_and10847_y0(h_u_cla32_and10846_y0, h_u_cla32_and10845_y0, h_u_cla32_and10847_y0);
  and_gate and_gate_h_u_cla32_and10848_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10848_y0);
  and_gate and_gate_h_u_cla32_and10849_y0(h_u_cla32_and10848_y0, h_u_cla32_and10847_y0, h_u_cla32_and10849_y0);
  and_gate and_gate_h_u_cla32_and10850_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10850_y0);
  and_gate and_gate_h_u_cla32_and10851_y0(h_u_cla32_and10850_y0, h_u_cla32_and10849_y0, h_u_cla32_and10851_y0);
  and_gate and_gate_h_u_cla32_and10852_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10852_y0);
  and_gate and_gate_h_u_cla32_and10853_y0(h_u_cla32_and10852_y0, h_u_cla32_and10851_y0, h_u_cla32_and10853_y0);
  and_gate and_gate_h_u_cla32_and10854_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10854_y0);
  and_gate and_gate_h_u_cla32_and10855_y0(h_u_cla32_and10854_y0, h_u_cla32_and10853_y0, h_u_cla32_and10855_y0);
  and_gate and_gate_h_u_cla32_and10856_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10856_y0);
  and_gate and_gate_h_u_cla32_and10857_y0(h_u_cla32_and10856_y0, h_u_cla32_and10855_y0, h_u_cla32_and10857_y0);
  and_gate and_gate_h_u_cla32_and10858_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10858_y0);
  and_gate and_gate_h_u_cla32_and10859_y0(h_u_cla32_and10858_y0, h_u_cla32_and10857_y0, h_u_cla32_and10859_y0);
  and_gate and_gate_h_u_cla32_and10860_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10860_y0);
  and_gate and_gate_h_u_cla32_and10861_y0(h_u_cla32_and10860_y0, h_u_cla32_and10859_y0, h_u_cla32_and10861_y0);
  and_gate and_gate_h_u_cla32_and10862_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic6_y1, h_u_cla32_and10862_y0);
  and_gate and_gate_h_u_cla32_and10863_y0(h_u_cla32_and10862_y0, h_u_cla32_and10861_y0, h_u_cla32_and10863_y0);
  and_gate and_gate_h_u_cla32_and10864_y0(h_u_cla32_pg_logic8_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10864_y0);
  and_gate and_gate_h_u_cla32_and10865_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10865_y0);
  and_gate and_gate_h_u_cla32_and10866_y0(h_u_cla32_and10865_y0, h_u_cla32_and10864_y0, h_u_cla32_and10866_y0);
  and_gate and_gate_h_u_cla32_and10867_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10867_y0);
  and_gate and_gate_h_u_cla32_and10868_y0(h_u_cla32_and10867_y0, h_u_cla32_and10866_y0, h_u_cla32_and10868_y0);
  and_gate and_gate_h_u_cla32_and10869_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10869_y0);
  and_gate and_gate_h_u_cla32_and10870_y0(h_u_cla32_and10869_y0, h_u_cla32_and10868_y0, h_u_cla32_and10870_y0);
  and_gate and_gate_h_u_cla32_and10871_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10871_y0);
  and_gate and_gate_h_u_cla32_and10872_y0(h_u_cla32_and10871_y0, h_u_cla32_and10870_y0, h_u_cla32_and10872_y0);
  and_gate and_gate_h_u_cla32_and10873_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10873_y0);
  and_gate and_gate_h_u_cla32_and10874_y0(h_u_cla32_and10873_y0, h_u_cla32_and10872_y0, h_u_cla32_and10874_y0);
  and_gate and_gate_h_u_cla32_and10875_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10875_y0);
  and_gate and_gate_h_u_cla32_and10876_y0(h_u_cla32_and10875_y0, h_u_cla32_and10874_y0, h_u_cla32_and10876_y0);
  and_gate and_gate_h_u_cla32_and10877_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10877_y0);
  and_gate and_gate_h_u_cla32_and10878_y0(h_u_cla32_and10877_y0, h_u_cla32_and10876_y0, h_u_cla32_and10878_y0);
  and_gate and_gate_h_u_cla32_and10879_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10879_y0);
  and_gate and_gate_h_u_cla32_and10880_y0(h_u_cla32_and10879_y0, h_u_cla32_and10878_y0, h_u_cla32_and10880_y0);
  and_gate and_gate_h_u_cla32_and10881_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10881_y0);
  and_gate and_gate_h_u_cla32_and10882_y0(h_u_cla32_and10881_y0, h_u_cla32_and10880_y0, h_u_cla32_and10882_y0);
  and_gate and_gate_h_u_cla32_and10883_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10883_y0);
  and_gate and_gate_h_u_cla32_and10884_y0(h_u_cla32_and10883_y0, h_u_cla32_and10882_y0, h_u_cla32_and10884_y0);
  and_gate and_gate_h_u_cla32_and10885_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10885_y0);
  and_gate and_gate_h_u_cla32_and10886_y0(h_u_cla32_and10885_y0, h_u_cla32_and10884_y0, h_u_cla32_and10886_y0);
  and_gate and_gate_h_u_cla32_and10887_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10887_y0);
  and_gate and_gate_h_u_cla32_and10888_y0(h_u_cla32_and10887_y0, h_u_cla32_and10886_y0, h_u_cla32_and10888_y0);
  and_gate and_gate_h_u_cla32_and10889_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10889_y0);
  and_gate and_gate_h_u_cla32_and10890_y0(h_u_cla32_and10889_y0, h_u_cla32_and10888_y0, h_u_cla32_and10890_y0);
  and_gate and_gate_h_u_cla32_and10891_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10891_y0);
  and_gate and_gate_h_u_cla32_and10892_y0(h_u_cla32_and10891_y0, h_u_cla32_and10890_y0, h_u_cla32_and10892_y0);
  and_gate and_gate_h_u_cla32_and10893_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10893_y0);
  and_gate and_gate_h_u_cla32_and10894_y0(h_u_cla32_and10893_y0, h_u_cla32_and10892_y0, h_u_cla32_and10894_y0);
  and_gate and_gate_h_u_cla32_and10895_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10895_y0);
  and_gate and_gate_h_u_cla32_and10896_y0(h_u_cla32_and10895_y0, h_u_cla32_and10894_y0, h_u_cla32_and10896_y0);
  and_gate and_gate_h_u_cla32_and10897_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10897_y0);
  and_gate and_gate_h_u_cla32_and10898_y0(h_u_cla32_and10897_y0, h_u_cla32_and10896_y0, h_u_cla32_and10898_y0);
  and_gate and_gate_h_u_cla32_and10899_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10899_y0);
  and_gate and_gate_h_u_cla32_and10900_y0(h_u_cla32_and10899_y0, h_u_cla32_and10898_y0, h_u_cla32_and10900_y0);
  and_gate and_gate_h_u_cla32_and10901_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10901_y0);
  and_gate and_gate_h_u_cla32_and10902_y0(h_u_cla32_and10901_y0, h_u_cla32_and10900_y0, h_u_cla32_and10902_y0);
  and_gate and_gate_h_u_cla32_and10903_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10903_y0);
  and_gate and_gate_h_u_cla32_and10904_y0(h_u_cla32_and10903_y0, h_u_cla32_and10902_y0, h_u_cla32_and10904_y0);
  and_gate and_gate_h_u_cla32_and10905_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10905_y0);
  and_gate and_gate_h_u_cla32_and10906_y0(h_u_cla32_and10905_y0, h_u_cla32_and10904_y0, h_u_cla32_and10906_y0);
  and_gate and_gate_h_u_cla32_and10907_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10907_y0);
  and_gate and_gate_h_u_cla32_and10908_y0(h_u_cla32_and10907_y0, h_u_cla32_and10906_y0, h_u_cla32_and10908_y0);
  and_gate and_gate_h_u_cla32_and10909_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic7_y1, h_u_cla32_and10909_y0);
  and_gate and_gate_h_u_cla32_and10910_y0(h_u_cla32_and10909_y0, h_u_cla32_and10908_y0, h_u_cla32_and10910_y0);
  and_gate and_gate_h_u_cla32_and10911_y0(h_u_cla32_pg_logic9_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10911_y0);
  and_gate and_gate_h_u_cla32_and10912_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10912_y0);
  and_gate and_gate_h_u_cla32_and10913_y0(h_u_cla32_and10912_y0, h_u_cla32_and10911_y0, h_u_cla32_and10913_y0);
  and_gate and_gate_h_u_cla32_and10914_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10914_y0);
  and_gate and_gate_h_u_cla32_and10915_y0(h_u_cla32_and10914_y0, h_u_cla32_and10913_y0, h_u_cla32_and10915_y0);
  and_gate and_gate_h_u_cla32_and10916_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10916_y0);
  and_gate and_gate_h_u_cla32_and10917_y0(h_u_cla32_and10916_y0, h_u_cla32_and10915_y0, h_u_cla32_and10917_y0);
  and_gate and_gate_h_u_cla32_and10918_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10918_y0);
  and_gate and_gate_h_u_cla32_and10919_y0(h_u_cla32_and10918_y0, h_u_cla32_and10917_y0, h_u_cla32_and10919_y0);
  and_gate and_gate_h_u_cla32_and10920_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10920_y0);
  and_gate and_gate_h_u_cla32_and10921_y0(h_u_cla32_and10920_y0, h_u_cla32_and10919_y0, h_u_cla32_and10921_y0);
  and_gate and_gate_h_u_cla32_and10922_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10922_y0);
  and_gate and_gate_h_u_cla32_and10923_y0(h_u_cla32_and10922_y0, h_u_cla32_and10921_y0, h_u_cla32_and10923_y0);
  and_gate and_gate_h_u_cla32_and10924_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10924_y0);
  and_gate and_gate_h_u_cla32_and10925_y0(h_u_cla32_and10924_y0, h_u_cla32_and10923_y0, h_u_cla32_and10925_y0);
  and_gate and_gate_h_u_cla32_and10926_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10926_y0);
  and_gate and_gate_h_u_cla32_and10927_y0(h_u_cla32_and10926_y0, h_u_cla32_and10925_y0, h_u_cla32_and10927_y0);
  and_gate and_gate_h_u_cla32_and10928_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10928_y0);
  and_gate and_gate_h_u_cla32_and10929_y0(h_u_cla32_and10928_y0, h_u_cla32_and10927_y0, h_u_cla32_and10929_y0);
  and_gate and_gate_h_u_cla32_and10930_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10930_y0);
  and_gate and_gate_h_u_cla32_and10931_y0(h_u_cla32_and10930_y0, h_u_cla32_and10929_y0, h_u_cla32_and10931_y0);
  and_gate and_gate_h_u_cla32_and10932_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10932_y0);
  and_gate and_gate_h_u_cla32_and10933_y0(h_u_cla32_and10932_y0, h_u_cla32_and10931_y0, h_u_cla32_and10933_y0);
  and_gate and_gate_h_u_cla32_and10934_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10934_y0);
  and_gate and_gate_h_u_cla32_and10935_y0(h_u_cla32_and10934_y0, h_u_cla32_and10933_y0, h_u_cla32_and10935_y0);
  and_gate and_gate_h_u_cla32_and10936_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10936_y0);
  and_gate and_gate_h_u_cla32_and10937_y0(h_u_cla32_and10936_y0, h_u_cla32_and10935_y0, h_u_cla32_and10937_y0);
  and_gate and_gate_h_u_cla32_and10938_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10938_y0);
  and_gate and_gate_h_u_cla32_and10939_y0(h_u_cla32_and10938_y0, h_u_cla32_and10937_y0, h_u_cla32_and10939_y0);
  and_gate and_gate_h_u_cla32_and10940_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10940_y0);
  and_gate and_gate_h_u_cla32_and10941_y0(h_u_cla32_and10940_y0, h_u_cla32_and10939_y0, h_u_cla32_and10941_y0);
  and_gate and_gate_h_u_cla32_and10942_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10942_y0);
  and_gate and_gate_h_u_cla32_and10943_y0(h_u_cla32_and10942_y0, h_u_cla32_and10941_y0, h_u_cla32_and10943_y0);
  and_gate and_gate_h_u_cla32_and10944_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10944_y0);
  and_gate and_gate_h_u_cla32_and10945_y0(h_u_cla32_and10944_y0, h_u_cla32_and10943_y0, h_u_cla32_and10945_y0);
  and_gate and_gate_h_u_cla32_and10946_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10946_y0);
  and_gate and_gate_h_u_cla32_and10947_y0(h_u_cla32_and10946_y0, h_u_cla32_and10945_y0, h_u_cla32_and10947_y0);
  and_gate and_gate_h_u_cla32_and10948_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10948_y0);
  and_gate and_gate_h_u_cla32_and10949_y0(h_u_cla32_and10948_y0, h_u_cla32_and10947_y0, h_u_cla32_and10949_y0);
  and_gate and_gate_h_u_cla32_and10950_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10950_y0);
  and_gate and_gate_h_u_cla32_and10951_y0(h_u_cla32_and10950_y0, h_u_cla32_and10949_y0, h_u_cla32_and10951_y0);
  and_gate and_gate_h_u_cla32_and10952_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10952_y0);
  and_gate and_gate_h_u_cla32_and10953_y0(h_u_cla32_and10952_y0, h_u_cla32_and10951_y0, h_u_cla32_and10953_y0);
  and_gate and_gate_h_u_cla32_and10954_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic8_y1, h_u_cla32_and10954_y0);
  and_gate and_gate_h_u_cla32_and10955_y0(h_u_cla32_and10954_y0, h_u_cla32_and10953_y0, h_u_cla32_and10955_y0);
  and_gate and_gate_h_u_cla32_and10956_y0(h_u_cla32_pg_logic10_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10956_y0);
  and_gate and_gate_h_u_cla32_and10957_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10957_y0);
  and_gate and_gate_h_u_cla32_and10958_y0(h_u_cla32_and10957_y0, h_u_cla32_and10956_y0, h_u_cla32_and10958_y0);
  and_gate and_gate_h_u_cla32_and10959_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10959_y0);
  and_gate and_gate_h_u_cla32_and10960_y0(h_u_cla32_and10959_y0, h_u_cla32_and10958_y0, h_u_cla32_and10960_y0);
  and_gate and_gate_h_u_cla32_and10961_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10961_y0);
  and_gate and_gate_h_u_cla32_and10962_y0(h_u_cla32_and10961_y0, h_u_cla32_and10960_y0, h_u_cla32_and10962_y0);
  and_gate and_gate_h_u_cla32_and10963_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10963_y0);
  and_gate and_gate_h_u_cla32_and10964_y0(h_u_cla32_and10963_y0, h_u_cla32_and10962_y0, h_u_cla32_and10964_y0);
  and_gate and_gate_h_u_cla32_and10965_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10965_y0);
  and_gate and_gate_h_u_cla32_and10966_y0(h_u_cla32_and10965_y0, h_u_cla32_and10964_y0, h_u_cla32_and10966_y0);
  and_gate and_gate_h_u_cla32_and10967_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10967_y0);
  and_gate and_gate_h_u_cla32_and10968_y0(h_u_cla32_and10967_y0, h_u_cla32_and10966_y0, h_u_cla32_and10968_y0);
  and_gate and_gate_h_u_cla32_and10969_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10969_y0);
  and_gate and_gate_h_u_cla32_and10970_y0(h_u_cla32_and10969_y0, h_u_cla32_and10968_y0, h_u_cla32_and10970_y0);
  and_gate and_gate_h_u_cla32_and10971_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10971_y0);
  and_gate and_gate_h_u_cla32_and10972_y0(h_u_cla32_and10971_y0, h_u_cla32_and10970_y0, h_u_cla32_and10972_y0);
  and_gate and_gate_h_u_cla32_and10973_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10973_y0);
  and_gate and_gate_h_u_cla32_and10974_y0(h_u_cla32_and10973_y0, h_u_cla32_and10972_y0, h_u_cla32_and10974_y0);
  and_gate and_gate_h_u_cla32_and10975_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10975_y0);
  and_gate and_gate_h_u_cla32_and10976_y0(h_u_cla32_and10975_y0, h_u_cla32_and10974_y0, h_u_cla32_and10976_y0);
  and_gate and_gate_h_u_cla32_and10977_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10977_y0);
  and_gate and_gate_h_u_cla32_and10978_y0(h_u_cla32_and10977_y0, h_u_cla32_and10976_y0, h_u_cla32_and10978_y0);
  and_gate and_gate_h_u_cla32_and10979_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10979_y0);
  and_gate and_gate_h_u_cla32_and10980_y0(h_u_cla32_and10979_y0, h_u_cla32_and10978_y0, h_u_cla32_and10980_y0);
  and_gate and_gate_h_u_cla32_and10981_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10981_y0);
  and_gate and_gate_h_u_cla32_and10982_y0(h_u_cla32_and10981_y0, h_u_cla32_and10980_y0, h_u_cla32_and10982_y0);
  and_gate and_gate_h_u_cla32_and10983_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10983_y0);
  and_gate and_gate_h_u_cla32_and10984_y0(h_u_cla32_and10983_y0, h_u_cla32_and10982_y0, h_u_cla32_and10984_y0);
  and_gate and_gate_h_u_cla32_and10985_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10985_y0);
  and_gate and_gate_h_u_cla32_and10986_y0(h_u_cla32_and10985_y0, h_u_cla32_and10984_y0, h_u_cla32_and10986_y0);
  and_gate and_gate_h_u_cla32_and10987_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10987_y0);
  and_gate and_gate_h_u_cla32_and10988_y0(h_u_cla32_and10987_y0, h_u_cla32_and10986_y0, h_u_cla32_and10988_y0);
  and_gate and_gate_h_u_cla32_and10989_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10989_y0);
  and_gate and_gate_h_u_cla32_and10990_y0(h_u_cla32_and10989_y0, h_u_cla32_and10988_y0, h_u_cla32_and10990_y0);
  and_gate and_gate_h_u_cla32_and10991_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10991_y0);
  and_gate and_gate_h_u_cla32_and10992_y0(h_u_cla32_and10991_y0, h_u_cla32_and10990_y0, h_u_cla32_and10992_y0);
  and_gate and_gate_h_u_cla32_and10993_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10993_y0);
  and_gate and_gate_h_u_cla32_and10994_y0(h_u_cla32_and10993_y0, h_u_cla32_and10992_y0, h_u_cla32_and10994_y0);
  and_gate and_gate_h_u_cla32_and10995_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10995_y0);
  and_gate and_gate_h_u_cla32_and10996_y0(h_u_cla32_and10995_y0, h_u_cla32_and10994_y0, h_u_cla32_and10996_y0);
  and_gate and_gate_h_u_cla32_and10997_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic9_y1, h_u_cla32_and10997_y0);
  and_gate and_gate_h_u_cla32_and10998_y0(h_u_cla32_and10997_y0, h_u_cla32_and10996_y0, h_u_cla32_and10998_y0);
  and_gate and_gate_h_u_cla32_and10999_y0(h_u_cla32_pg_logic11_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and10999_y0);
  and_gate and_gate_h_u_cla32_and11000_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11000_y0);
  and_gate and_gate_h_u_cla32_and11001_y0(h_u_cla32_and11000_y0, h_u_cla32_and10999_y0, h_u_cla32_and11001_y0);
  and_gate and_gate_h_u_cla32_and11002_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11002_y0);
  and_gate and_gate_h_u_cla32_and11003_y0(h_u_cla32_and11002_y0, h_u_cla32_and11001_y0, h_u_cla32_and11003_y0);
  and_gate and_gate_h_u_cla32_and11004_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11004_y0);
  and_gate and_gate_h_u_cla32_and11005_y0(h_u_cla32_and11004_y0, h_u_cla32_and11003_y0, h_u_cla32_and11005_y0);
  and_gate and_gate_h_u_cla32_and11006_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11006_y0);
  and_gate and_gate_h_u_cla32_and11007_y0(h_u_cla32_and11006_y0, h_u_cla32_and11005_y0, h_u_cla32_and11007_y0);
  and_gate and_gate_h_u_cla32_and11008_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11008_y0);
  and_gate and_gate_h_u_cla32_and11009_y0(h_u_cla32_and11008_y0, h_u_cla32_and11007_y0, h_u_cla32_and11009_y0);
  and_gate and_gate_h_u_cla32_and11010_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11010_y0);
  and_gate and_gate_h_u_cla32_and11011_y0(h_u_cla32_and11010_y0, h_u_cla32_and11009_y0, h_u_cla32_and11011_y0);
  and_gate and_gate_h_u_cla32_and11012_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11012_y0);
  and_gate and_gate_h_u_cla32_and11013_y0(h_u_cla32_and11012_y0, h_u_cla32_and11011_y0, h_u_cla32_and11013_y0);
  and_gate and_gate_h_u_cla32_and11014_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11014_y0);
  and_gate and_gate_h_u_cla32_and11015_y0(h_u_cla32_and11014_y0, h_u_cla32_and11013_y0, h_u_cla32_and11015_y0);
  and_gate and_gate_h_u_cla32_and11016_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11016_y0);
  and_gate and_gate_h_u_cla32_and11017_y0(h_u_cla32_and11016_y0, h_u_cla32_and11015_y0, h_u_cla32_and11017_y0);
  and_gate and_gate_h_u_cla32_and11018_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11018_y0);
  and_gate and_gate_h_u_cla32_and11019_y0(h_u_cla32_and11018_y0, h_u_cla32_and11017_y0, h_u_cla32_and11019_y0);
  and_gate and_gate_h_u_cla32_and11020_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11020_y0);
  and_gate and_gate_h_u_cla32_and11021_y0(h_u_cla32_and11020_y0, h_u_cla32_and11019_y0, h_u_cla32_and11021_y0);
  and_gate and_gate_h_u_cla32_and11022_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11022_y0);
  and_gate and_gate_h_u_cla32_and11023_y0(h_u_cla32_and11022_y0, h_u_cla32_and11021_y0, h_u_cla32_and11023_y0);
  and_gate and_gate_h_u_cla32_and11024_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11024_y0);
  and_gate and_gate_h_u_cla32_and11025_y0(h_u_cla32_and11024_y0, h_u_cla32_and11023_y0, h_u_cla32_and11025_y0);
  and_gate and_gate_h_u_cla32_and11026_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11026_y0);
  and_gate and_gate_h_u_cla32_and11027_y0(h_u_cla32_and11026_y0, h_u_cla32_and11025_y0, h_u_cla32_and11027_y0);
  and_gate and_gate_h_u_cla32_and11028_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11028_y0);
  and_gate and_gate_h_u_cla32_and11029_y0(h_u_cla32_and11028_y0, h_u_cla32_and11027_y0, h_u_cla32_and11029_y0);
  and_gate and_gate_h_u_cla32_and11030_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11030_y0);
  and_gate and_gate_h_u_cla32_and11031_y0(h_u_cla32_and11030_y0, h_u_cla32_and11029_y0, h_u_cla32_and11031_y0);
  and_gate and_gate_h_u_cla32_and11032_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11032_y0);
  and_gate and_gate_h_u_cla32_and11033_y0(h_u_cla32_and11032_y0, h_u_cla32_and11031_y0, h_u_cla32_and11033_y0);
  and_gate and_gate_h_u_cla32_and11034_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11034_y0);
  and_gate and_gate_h_u_cla32_and11035_y0(h_u_cla32_and11034_y0, h_u_cla32_and11033_y0, h_u_cla32_and11035_y0);
  and_gate and_gate_h_u_cla32_and11036_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11036_y0);
  and_gate and_gate_h_u_cla32_and11037_y0(h_u_cla32_and11036_y0, h_u_cla32_and11035_y0, h_u_cla32_and11037_y0);
  and_gate and_gate_h_u_cla32_and11038_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic10_y1, h_u_cla32_and11038_y0);
  and_gate and_gate_h_u_cla32_and11039_y0(h_u_cla32_and11038_y0, h_u_cla32_and11037_y0, h_u_cla32_and11039_y0);
  and_gate and_gate_h_u_cla32_and11040_y0(h_u_cla32_pg_logic12_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11040_y0);
  and_gate and_gate_h_u_cla32_and11041_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11041_y0);
  and_gate and_gate_h_u_cla32_and11042_y0(h_u_cla32_and11041_y0, h_u_cla32_and11040_y0, h_u_cla32_and11042_y0);
  and_gate and_gate_h_u_cla32_and11043_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11043_y0);
  and_gate and_gate_h_u_cla32_and11044_y0(h_u_cla32_and11043_y0, h_u_cla32_and11042_y0, h_u_cla32_and11044_y0);
  and_gate and_gate_h_u_cla32_and11045_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11045_y0);
  and_gate and_gate_h_u_cla32_and11046_y0(h_u_cla32_and11045_y0, h_u_cla32_and11044_y0, h_u_cla32_and11046_y0);
  and_gate and_gate_h_u_cla32_and11047_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11047_y0);
  and_gate and_gate_h_u_cla32_and11048_y0(h_u_cla32_and11047_y0, h_u_cla32_and11046_y0, h_u_cla32_and11048_y0);
  and_gate and_gate_h_u_cla32_and11049_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11049_y0);
  and_gate and_gate_h_u_cla32_and11050_y0(h_u_cla32_and11049_y0, h_u_cla32_and11048_y0, h_u_cla32_and11050_y0);
  and_gate and_gate_h_u_cla32_and11051_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11051_y0);
  and_gate and_gate_h_u_cla32_and11052_y0(h_u_cla32_and11051_y0, h_u_cla32_and11050_y0, h_u_cla32_and11052_y0);
  and_gate and_gate_h_u_cla32_and11053_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11053_y0);
  and_gate and_gate_h_u_cla32_and11054_y0(h_u_cla32_and11053_y0, h_u_cla32_and11052_y0, h_u_cla32_and11054_y0);
  and_gate and_gate_h_u_cla32_and11055_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11055_y0);
  and_gate and_gate_h_u_cla32_and11056_y0(h_u_cla32_and11055_y0, h_u_cla32_and11054_y0, h_u_cla32_and11056_y0);
  and_gate and_gate_h_u_cla32_and11057_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11057_y0);
  and_gate and_gate_h_u_cla32_and11058_y0(h_u_cla32_and11057_y0, h_u_cla32_and11056_y0, h_u_cla32_and11058_y0);
  and_gate and_gate_h_u_cla32_and11059_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11059_y0);
  and_gate and_gate_h_u_cla32_and11060_y0(h_u_cla32_and11059_y0, h_u_cla32_and11058_y0, h_u_cla32_and11060_y0);
  and_gate and_gate_h_u_cla32_and11061_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11061_y0);
  and_gate and_gate_h_u_cla32_and11062_y0(h_u_cla32_and11061_y0, h_u_cla32_and11060_y0, h_u_cla32_and11062_y0);
  and_gate and_gate_h_u_cla32_and11063_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11063_y0);
  and_gate and_gate_h_u_cla32_and11064_y0(h_u_cla32_and11063_y0, h_u_cla32_and11062_y0, h_u_cla32_and11064_y0);
  and_gate and_gate_h_u_cla32_and11065_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11065_y0);
  and_gate and_gate_h_u_cla32_and11066_y0(h_u_cla32_and11065_y0, h_u_cla32_and11064_y0, h_u_cla32_and11066_y0);
  and_gate and_gate_h_u_cla32_and11067_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11067_y0);
  and_gate and_gate_h_u_cla32_and11068_y0(h_u_cla32_and11067_y0, h_u_cla32_and11066_y0, h_u_cla32_and11068_y0);
  and_gate and_gate_h_u_cla32_and11069_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11069_y0);
  and_gate and_gate_h_u_cla32_and11070_y0(h_u_cla32_and11069_y0, h_u_cla32_and11068_y0, h_u_cla32_and11070_y0);
  and_gate and_gate_h_u_cla32_and11071_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11071_y0);
  and_gate and_gate_h_u_cla32_and11072_y0(h_u_cla32_and11071_y0, h_u_cla32_and11070_y0, h_u_cla32_and11072_y0);
  and_gate and_gate_h_u_cla32_and11073_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11073_y0);
  and_gate and_gate_h_u_cla32_and11074_y0(h_u_cla32_and11073_y0, h_u_cla32_and11072_y0, h_u_cla32_and11074_y0);
  and_gate and_gate_h_u_cla32_and11075_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11075_y0);
  and_gate and_gate_h_u_cla32_and11076_y0(h_u_cla32_and11075_y0, h_u_cla32_and11074_y0, h_u_cla32_and11076_y0);
  and_gate and_gate_h_u_cla32_and11077_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic11_y1, h_u_cla32_and11077_y0);
  and_gate and_gate_h_u_cla32_and11078_y0(h_u_cla32_and11077_y0, h_u_cla32_and11076_y0, h_u_cla32_and11078_y0);
  and_gate and_gate_h_u_cla32_and11079_y0(h_u_cla32_pg_logic13_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11079_y0);
  and_gate and_gate_h_u_cla32_and11080_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11080_y0);
  and_gate and_gate_h_u_cla32_and11081_y0(h_u_cla32_and11080_y0, h_u_cla32_and11079_y0, h_u_cla32_and11081_y0);
  and_gate and_gate_h_u_cla32_and11082_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11082_y0);
  and_gate and_gate_h_u_cla32_and11083_y0(h_u_cla32_and11082_y0, h_u_cla32_and11081_y0, h_u_cla32_and11083_y0);
  and_gate and_gate_h_u_cla32_and11084_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11084_y0);
  and_gate and_gate_h_u_cla32_and11085_y0(h_u_cla32_and11084_y0, h_u_cla32_and11083_y0, h_u_cla32_and11085_y0);
  and_gate and_gate_h_u_cla32_and11086_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11086_y0);
  and_gate and_gate_h_u_cla32_and11087_y0(h_u_cla32_and11086_y0, h_u_cla32_and11085_y0, h_u_cla32_and11087_y0);
  and_gate and_gate_h_u_cla32_and11088_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11088_y0);
  and_gate and_gate_h_u_cla32_and11089_y0(h_u_cla32_and11088_y0, h_u_cla32_and11087_y0, h_u_cla32_and11089_y0);
  and_gate and_gate_h_u_cla32_and11090_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11090_y0);
  and_gate and_gate_h_u_cla32_and11091_y0(h_u_cla32_and11090_y0, h_u_cla32_and11089_y0, h_u_cla32_and11091_y0);
  and_gate and_gate_h_u_cla32_and11092_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11092_y0);
  and_gate and_gate_h_u_cla32_and11093_y0(h_u_cla32_and11092_y0, h_u_cla32_and11091_y0, h_u_cla32_and11093_y0);
  and_gate and_gate_h_u_cla32_and11094_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11094_y0);
  and_gate and_gate_h_u_cla32_and11095_y0(h_u_cla32_and11094_y0, h_u_cla32_and11093_y0, h_u_cla32_and11095_y0);
  and_gate and_gate_h_u_cla32_and11096_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11096_y0);
  and_gate and_gate_h_u_cla32_and11097_y0(h_u_cla32_and11096_y0, h_u_cla32_and11095_y0, h_u_cla32_and11097_y0);
  and_gate and_gate_h_u_cla32_and11098_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11098_y0);
  and_gate and_gate_h_u_cla32_and11099_y0(h_u_cla32_and11098_y0, h_u_cla32_and11097_y0, h_u_cla32_and11099_y0);
  and_gate and_gate_h_u_cla32_and11100_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11100_y0);
  and_gate and_gate_h_u_cla32_and11101_y0(h_u_cla32_and11100_y0, h_u_cla32_and11099_y0, h_u_cla32_and11101_y0);
  and_gate and_gate_h_u_cla32_and11102_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11102_y0);
  and_gate and_gate_h_u_cla32_and11103_y0(h_u_cla32_and11102_y0, h_u_cla32_and11101_y0, h_u_cla32_and11103_y0);
  and_gate and_gate_h_u_cla32_and11104_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11104_y0);
  and_gate and_gate_h_u_cla32_and11105_y0(h_u_cla32_and11104_y0, h_u_cla32_and11103_y0, h_u_cla32_and11105_y0);
  and_gate and_gate_h_u_cla32_and11106_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11106_y0);
  and_gate and_gate_h_u_cla32_and11107_y0(h_u_cla32_and11106_y0, h_u_cla32_and11105_y0, h_u_cla32_and11107_y0);
  and_gate and_gate_h_u_cla32_and11108_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11108_y0);
  and_gate and_gate_h_u_cla32_and11109_y0(h_u_cla32_and11108_y0, h_u_cla32_and11107_y0, h_u_cla32_and11109_y0);
  and_gate and_gate_h_u_cla32_and11110_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11110_y0);
  and_gate and_gate_h_u_cla32_and11111_y0(h_u_cla32_and11110_y0, h_u_cla32_and11109_y0, h_u_cla32_and11111_y0);
  and_gate and_gate_h_u_cla32_and11112_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11112_y0);
  and_gate and_gate_h_u_cla32_and11113_y0(h_u_cla32_and11112_y0, h_u_cla32_and11111_y0, h_u_cla32_and11113_y0);
  and_gate and_gate_h_u_cla32_and11114_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic12_y1, h_u_cla32_and11114_y0);
  and_gate and_gate_h_u_cla32_and11115_y0(h_u_cla32_and11114_y0, h_u_cla32_and11113_y0, h_u_cla32_and11115_y0);
  and_gate and_gate_h_u_cla32_and11116_y0(h_u_cla32_pg_logic14_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11116_y0);
  and_gate and_gate_h_u_cla32_and11117_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11117_y0);
  and_gate and_gate_h_u_cla32_and11118_y0(h_u_cla32_and11117_y0, h_u_cla32_and11116_y0, h_u_cla32_and11118_y0);
  and_gate and_gate_h_u_cla32_and11119_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11119_y0);
  and_gate and_gate_h_u_cla32_and11120_y0(h_u_cla32_and11119_y0, h_u_cla32_and11118_y0, h_u_cla32_and11120_y0);
  and_gate and_gate_h_u_cla32_and11121_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11121_y0);
  and_gate and_gate_h_u_cla32_and11122_y0(h_u_cla32_and11121_y0, h_u_cla32_and11120_y0, h_u_cla32_and11122_y0);
  and_gate and_gate_h_u_cla32_and11123_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11123_y0);
  and_gate and_gate_h_u_cla32_and11124_y0(h_u_cla32_and11123_y0, h_u_cla32_and11122_y0, h_u_cla32_and11124_y0);
  and_gate and_gate_h_u_cla32_and11125_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11125_y0);
  and_gate and_gate_h_u_cla32_and11126_y0(h_u_cla32_and11125_y0, h_u_cla32_and11124_y0, h_u_cla32_and11126_y0);
  and_gate and_gate_h_u_cla32_and11127_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11127_y0);
  and_gate and_gate_h_u_cla32_and11128_y0(h_u_cla32_and11127_y0, h_u_cla32_and11126_y0, h_u_cla32_and11128_y0);
  and_gate and_gate_h_u_cla32_and11129_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11129_y0);
  and_gate and_gate_h_u_cla32_and11130_y0(h_u_cla32_and11129_y0, h_u_cla32_and11128_y0, h_u_cla32_and11130_y0);
  and_gate and_gate_h_u_cla32_and11131_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11131_y0);
  and_gate and_gate_h_u_cla32_and11132_y0(h_u_cla32_and11131_y0, h_u_cla32_and11130_y0, h_u_cla32_and11132_y0);
  and_gate and_gate_h_u_cla32_and11133_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11133_y0);
  and_gate and_gate_h_u_cla32_and11134_y0(h_u_cla32_and11133_y0, h_u_cla32_and11132_y0, h_u_cla32_and11134_y0);
  and_gate and_gate_h_u_cla32_and11135_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11135_y0);
  and_gate and_gate_h_u_cla32_and11136_y0(h_u_cla32_and11135_y0, h_u_cla32_and11134_y0, h_u_cla32_and11136_y0);
  and_gate and_gate_h_u_cla32_and11137_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11137_y0);
  and_gate and_gate_h_u_cla32_and11138_y0(h_u_cla32_and11137_y0, h_u_cla32_and11136_y0, h_u_cla32_and11138_y0);
  and_gate and_gate_h_u_cla32_and11139_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11139_y0);
  and_gate and_gate_h_u_cla32_and11140_y0(h_u_cla32_and11139_y0, h_u_cla32_and11138_y0, h_u_cla32_and11140_y0);
  and_gate and_gate_h_u_cla32_and11141_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11141_y0);
  and_gate and_gate_h_u_cla32_and11142_y0(h_u_cla32_and11141_y0, h_u_cla32_and11140_y0, h_u_cla32_and11142_y0);
  and_gate and_gate_h_u_cla32_and11143_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11143_y0);
  and_gate and_gate_h_u_cla32_and11144_y0(h_u_cla32_and11143_y0, h_u_cla32_and11142_y0, h_u_cla32_and11144_y0);
  and_gate and_gate_h_u_cla32_and11145_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11145_y0);
  and_gate and_gate_h_u_cla32_and11146_y0(h_u_cla32_and11145_y0, h_u_cla32_and11144_y0, h_u_cla32_and11146_y0);
  and_gate and_gate_h_u_cla32_and11147_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11147_y0);
  and_gate and_gate_h_u_cla32_and11148_y0(h_u_cla32_and11147_y0, h_u_cla32_and11146_y0, h_u_cla32_and11148_y0);
  and_gate and_gate_h_u_cla32_and11149_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic13_y1, h_u_cla32_and11149_y0);
  and_gate and_gate_h_u_cla32_and11150_y0(h_u_cla32_and11149_y0, h_u_cla32_and11148_y0, h_u_cla32_and11150_y0);
  and_gate and_gate_h_u_cla32_and11151_y0(h_u_cla32_pg_logic15_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11151_y0);
  and_gate and_gate_h_u_cla32_and11152_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11152_y0);
  and_gate and_gate_h_u_cla32_and11153_y0(h_u_cla32_and11152_y0, h_u_cla32_and11151_y0, h_u_cla32_and11153_y0);
  and_gate and_gate_h_u_cla32_and11154_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11154_y0);
  and_gate and_gate_h_u_cla32_and11155_y0(h_u_cla32_and11154_y0, h_u_cla32_and11153_y0, h_u_cla32_and11155_y0);
  and_gate and_gate_h_u_cla32_and11156_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11156_y0);
  and_gate and_gate_h_u_cla32_and11157_y0(h_u_cla32_and11156_y0, h_u_cla32_and11155_y0, h_u_cla32_and11157_y0);
  and_gate and_gate_h_u_cla32_and11158_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11158_y0);
  and_gate and_gate_h_u_cla32_and11159_y0(h_u_cla32_and11158_y0, h_u_cla32_and11157_y0, h_u_cla32_and11159_y0);
  and_gate and_gate_h_u_cla32_and11160_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11160_y0);
  and_gate and_gate_h_u_cla32_and11161_y0(h_u_cla32_and11160_y0, h_u_cla32_and11159_y0, h_u_cla32_and11161_y0);
  and_gate and_gate_h_u_cla32_and11162_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11162_y0);
  and_gate and_gate_h_u_cla32_and11163_y0(h_u_cla32_and11162_y0, h_u_cla32_and11161_y0, h_u_cla32_and11163_y0);
  and_gate and_gate_h_u_cla32_and11164_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11164_y0);
  and_gate and_gate_h_u_cla32_and11165_y0(h_u_cla32_and11164_y0, h_u_cla32_and11163_y0, h_u_cla32_and11165_y0);
  and_gate and_gate_h_u_cla32_and11166_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11166_y0);
  and_gate and_gate_h_u_cla32_and11167_y0(h_u_cla32_and11166_y0, h_u_cla32_and11165_y0, h_u_cla32_and11167_y0);
  and_gate and_gate_h_u_cla32_and11168_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11168_y0);
  and_gate and_gate_h_u_cla32_and11169_y0(h_u_cla32_and11168_y0, h_u_cla32_and11167_y0, h_u_cla32_and11169_y0);
  and_gate and_gate_h_u_cla32_and11170_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11170_y0);
  and_gate and_gate_h_u_cla32_and11171_y0(h_u_cla32_and11170_y0, h_u_cla32_and11169_y0, h_u_cla32_and11171_y0);
  and_gate and_gate_h_u_cla32_and11172_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11172_y0);
  and_gate and_gate_h_u_cla32_and11173_y0(h_u_cla32_and11172_y0, h_u_cla32_and11171_y0, h_u_cla32_and11173_y0);
  and_gate and_gate_h_u_cla32_and11174_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11174_y0);
  and_gate and_gate_h_u_cla32_and11175_y0(h_u_cla32_and11174_y0, h_u_cla32_and11173_y0, h_u_cla32_and11175_y0);
  and_gate and_gate_h_u_cla32_and11176_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11176_y0);
  and_gate and_gate_h_u_cla32_and11177_y0(h_u_cla32_and11176_y0, h_u_cla32_and11175_y0, h_u_cla32_and11177_y0);
  and_gate and_gate_h_u_cla32_and11178_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11178_y0);
  and_gate and_gate_h_u_cla32_and11179_y0(h_u_cla32_and11178_y0, h_u_cla32_and11177_y0, h_u_cla32_and11179_y0);
  and_gate and_gate_h_u_cla32_and11180_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11180_y0);
  and_gate and_gate_h_u_cla32_and11181_y0(h_u_cla32_and11180_y0, h_u_cla32_and11179_y0, h_u_cla32_and11181_y0);
  and_gate and_gate_h_u_cla32_and11182_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic14_y1, h_u_cla32_and11182_y0);
  and_gate and_gate_h_u_cla32_and11183_y0(h_u_cla32_and11182_y0, h_u_cla32_and11181_y0, h_u_cla32_and11183_y0);
  and_gate and_gate_h_u_cla32_and11184_y0(h_u_cla32_pg_logic16_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11184_y0);
  and_gate and_gate_h_u_cla32_and11185_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11185_y0);
  and_gate and_gate_h_u_cla32_and11186_y0(h_u_cla32_and11185_y0, h_u_cla32_and11184_y0, h_u_cla32_and11186_y0);
  and_gate and_gate_h_u_cla32_and11187_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11187_y0);
  and_gate and_gate_h_u_cla32_and11188_y0(h_u_cla32_and11187_y0, h_u_cla32_and11186_y0, h_u_cla32_and11188_y0);
  and_gate and_gate_h_u_cla32_and11189_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11189_y0);
  and_gate and_gate_h_u_cla32_and11190_y0(h_u_cla32_and11189_y0, h_u_cla32_and11188_y0, h_u_cla32_and11190_y0);
  and_gate and_gate_h_u_cla32_and11191_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11191_y0);
  and_gate and_gate_h_u_cla32_and11192_y0(h_u_cla32_and11191_y0, h_u_cla32_and11190_y0, h_u_cla32_and11192_y0);
  and_gate and_gate_h_u_cla32_and11193_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11193_y0);
  and_gate and_gate_h_u_cla32_and11194_y0(h_u_cla32_and11193_y0, h_u_cla32_and11192_y0, h_u_cla32_and11194_y0);
  and_gate and_gate_h_u_cla32_and11195_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11195_y0);
  and_gate and_gate_h_u_cla32_and11196_y0(h_u_cla32_and11195_y0, h_u_cla32_and11194_y0, h_u_cla32_and11196_y0);
  and_gate and_gate_h_u_cla32_and11197_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11197_y0);
  and_gate and_gate_h_u_cla32_and11198_y0(h_u_cla32_and11197_y0, h_u_cla32_and11196_y0, h_u_cla32_and11198_y0);
  and_gate and_gate_h_u_cla32_and11199_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11199_y0);
  and_gate and_gate_h_u_cla32_and11200_y0(h_u_cla32_and11199_y0, h_u_cla32_and11198_y0, h_u_cla32_and11200_y0);
  and_gate and_gate_h_u_cla32_and11201_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11201_y0);
  and_gate and_gate_h_u_cla32_and11202_y0(h_u_cla32_and11201_y0, h_u_cla32_and11200_y0, h_u_cla32_and11202_y0);
  and_gate and_gate_h_u_cla32_and11203_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11203_y0);
  and_gate and_gate_h_u_cla32_and11204_y0(h_u_cla32_and11203_y0, h_u_cla32_and11202_y0, h_u_cla32_and11204_y0);
  and_gate and_gate_h_u_cla32_and11205_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11205_y0);
  and_gate and_gate_h_u_cla32_and11206_y0(h_u_cla32_and11205_y0, h_u_cla32_and11204_y0, h_u_cla32_and11206_y0);
  and_gate and_gate_h_u_cla32_and11207_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11207_y0);
  and_gate and_gate_h_u_cla32_and11208_y0(h_u_cla32_and11207_y0, h_u_cla32_and11206_y0, h_u_cla32_and11208_y0);
  and_gate and_gate_h_u_cla32_and11209_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11209_y0);
  and_gate and_gate_h_u_cla32_and11210_y0(h_u_cla32_and11209_y0, h_u_cla32_and11208_y0, h_u_cla32_and11210_y0);
  and_gate and_gate_h_u_cla32_and11211_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11211_y0);
  and_gate and_gate_h_u_cla32_and11212_y0(h_u_cla32_and11211_y0, h_u_cla32_and11210_y0, h_u_cla32_and11212_y0);
  and_gate and_gate_h_u_cla32_and11213_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic15_y1, h_u_cla32_and11213_y0);
  and_gate and_gate_h_u_cla32_and11214_y0(h_u_cla32_and11213_y0, h_u_cla32_and11212_y0, h_u_cla32_and11214_y0);
  and_gate and_gate_h_u_cla32_and11215_y0(h_u_cla32_pg_logic17_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11215_y0);
  and_gate and_gate_h_u_cla32_and11216_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11216_y0);
  and_gate and_gate_h_u_cla32_and11217_y0(h_u_cla32_and11216_y0, h_u_cla32_and11215_y0, h_u_cla32_and11217_y0);
  and_gate and_gate_h_u_cla32_and11218_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11218_y0);
  and_gate and_gate_h_u_cla32_and11219_y0(h_u_cla32_and11218_y0, h_u_cla32_and11217_y0, h_u_cla32_and11219_y0);
  and_gate and_gate_h_u_cla32_and11220_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11220_y0);
  and_gate and_gate_h_u_cla32_and11221_y0(h_u_cla32_and11220_y0, h_u_cla32_and11219_y0, h_u_cla32_and11221_y0);
  and_gate and_gate_h_u_cla32_and11222_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11222_y0);
  and_gate and_gate_h_u_cla32_and11223_y0(h_u_cla32_and11222_y0, h_u_cla32_and11221_y0, h_u_cla32_and11223_y0);
  and_gate and_gate_h_u_cla32_and11224_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11224_y0);
  and_gate and_gate_h_u_cla32_and11225_y0(h_u_cla32_and11224_y0, h_u_cla32_and11223_y0, h_u_cla32_and11225_y0);
  and_gate and_gate_h_u_cla32_and11226_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11226_y0);
  and_gate and_gate_h_u_cla32_and11227_y0(h_u_cla32_and11226_y0, h_u_cla32_and11225_y0, h_u_cla32_and11227_y0);
  and_gate and_gate_h_u_cla32_and11228_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11228_y0);
  and_gate and_gate_h_u_cla32_and11229_y0(h_u_cla32_and11228_y0, h_u_cla32_and11227_y0, h_u_cla32_and11229_y0);
  and_gate and_gate_h_u_cla32_and11230_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11230_y0);
  and_gate and_gate_h_u_cla32_and11231_y0(h_u_cla32_and11230_y0, h_u_cla32_and11229_y0, h_u_cla32_and11231_y0);
  and_gate and_gate_h_u_cla32_and11232_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11232_y0);
  and_gate and_gate_h_u_cla32_and11233_y0(h_u_cla32_and11232_y0, h_u_cla32_and11231_y0, h_u_cla32_and11233_y0);
  and_gate and_gate_h_u_cla32_and11234_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11234_y0);
  and_gate and_gate_h_u_cla32_and11235_y0(h_u_cla32_and11234_y0, h_u_cla32_and11233_y0, h_u_cla32_and11235_y0);
  and_gate and_gate_h_u_cla32_and11236_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11236_y0);
  and_gate and_gate_h_u_cla32_and11237_y0(h_u_cla32_and11236_y0, h_u_cla32_and11235_y0, h_u_cla32_and11237_y0);
  and_gate and_gate_h_u_cla32_and11238_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11238_y0);
  and_gate and_gate_h_u_cla32_and11239_y0(h_u_cla32_and11238_y0, h_u_cla32_and11237_y0, h_u_cla32_and11239_y0);
  and_gate and_gate_h_u_cla32_and11240_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11240_y0);
  and_gate and_gate_h_u_cla32_and11241_y0(h_u_cla32_and11240_y0, h_u_cla32_and11239_y0, h_u_cla32_and11241_y0);
  and_gate and_gate_h_u_cla32_and11242_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic16_y1, h_u_cla32_and11242_y0);
  and_gate and_gate_h_u_cla32_and11243_y0(h_u_cla32_and11242_y0, h_u_cla32_and11241_y0, h_u_cla32_and11243_y0);
  and_gate and_gate_h_u_cla32_and11244_y0(h_u_cla32_pg_logic18_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11244_y0);
  and_gate and_gate_h_u_cla32_and11245_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11245_y0);
  and_gate and_gate_h_u_cla32_and11246_y0(h_u_cla32_and11245_y0, h_u_cla32_and11244_y0, h_u_cla32_and11246_y0);
  and_gate and_gate_h_u_cla32_and11247_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11247_y0);
  and_gate and_gate_h_u_cla32_and11248_y0(h_u_cla32_and11247_y0, h_u_cla32_and11246_y0, h_u_cla32_and11248_y0);
  and_gate and_gate_h_u_cla32_and11249_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11249_y0);
  and_gate and_gate_h_u_cla32_and11250_y0(h_u_cla32_and11249_y0, h_u_cla32_and11248_y0, h_u_cla32_and11250_y0);
  and_gate and_gate_h_u_cla32_and11251_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11251_y0);
  and_gate and_gate_h_u_cla32_and11252_y0(h_u_cla32_and11251_y0, h_u_cla32_and11250_y0, h_u_cla32_and11252_y0);
  and_gate and_gate_h_u_cla32_and11253_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11253_y0);
  and_gate and_gate_h_u_cla32_and11254_y0(h_u_cla32_and11253_y0, h_u_cla32_and11252_y0, h_u_cla32_and11254_y0);
  and_gate and_gate_h_u_cla32_and11255_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11255_y0);
  and_gate and_gate_h_u_cla32_and11256_y0(h_u_cla32_and11255_y0, h_u_cla32_and11254_y0, h_u_cla32_and11256_y0);
  and_gate and_gate_h_u_cla32_and11257_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11257_y0);
  and_gate and_gate_h_u_cla32_and11258_y0(h_u_cla32_and11257_y0, h_u_cla32_and11256_y0, h_u_cla32_and11258_y0);
  and_gate and_gate_h_u_cla32_and11259_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11259_y0);
  and_gate and_gate_h_u_cla32_and11260_y0(h_u_cla32_and11259_y0, h_u_cla32_and11258_y0, h_u_cla32_and11260_y0);
  and_gate and_gate_h_u_cla32_and11261_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11261_y0);
  and_gate and_gate_h_u_cla32_and11262_y0(h_u_cla32_and11261_y0, h_u_cla32_and11260_y0, h_u_cla32_and11262_y0);
  and_gate and_gate_h_u_cla32_and11263_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11263_y0);
  and_gate and_gate_h_u_cla32_and11264_y0(h_u_cla32_and11263_y0, h_u_cla32_and11262_y0, h_u_cla32_and11264_y0);
  and_gate and_gate_h_u_cla32_and11265_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11265_y0);
  and_gate and_gate_h_u_cla32_and11266_y0(h_u_cla32_and11265_y0, h_u_cla32_and11264_y0, h_u_cla32_and11266_y0);
  and_gate and_gate_h_u_cla32_and11267_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11267_y0);
  and_gate and_gate_h_u_cla32_and11268_y0(h_u_cla32_and11267_y0, h_u_cla32_and11266_y0, h_u_cla32_and11268_y0);
  and_gate and_gate_h_u_cla32_and11269_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic17_y1, h_u_cla32_and11269_y0);
  and_gate and_gate_h_u_cla32_and11270_y0(h_u_cla32_and11269_y0, h_u_cla32_and11268_y0, h_u_cla32_and11270_y0);
  and_gate and_gate_h_u_cla32_and11271_y0(h_u_cla32_pg_logic19_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11271_y0);
  and_gate and_gate_h_u_cla32_and11272_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11272_y0);
  and_gate and_gate_h_u_cla32_and11273_y0(h_u_cla32_and11272_y0, h_u_cla32_and11271_y0, h_u_cla32_and11273_y0);
  and_gate and_gate_h_u_cla32_and11274_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11274_y0);
  and_gate and_gate_h_u_cla32_and11275_y0(h_u_cla32_and11274_y0, h_u_cla32_and11273_y0, h_u_cla32_and11275_y0);
  and_gate and_gate_h_u_cla32_and11276_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11276_y0);
  and_gate and_gate_h_u_cla32_and11277_y0(h_u_cla32_and11276_y0, h_u_cla32_and11275_y0, h_u_cla32_and11277_y0);
  and_gate and_gate_h_u_cla32_and11278_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11278_y0);
  and_gate and_gate_h_u_cla32_and11279_y0(h_u_cla32_and11278_y0, h_u_cla32_and11277_y0, h_u_cla32_and11279_y0);
  and_gate and_gate_h_u_cla32_and11280_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11280_y0);
  and_gate and_gate_h_u_cla32_and11281_y0(h_u_cla32_and11280_y0, h_u_cla32_and11279_y0, h_u_cla32_and11281_y0);
  and_gate and_gate_h_u_cla32_and11282_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11282_y0);
  and_gate and_gate_h_u_cla32_and11283_y0(h_u_cla32_and11282_y0, h_u_cla32_and11281_y0, h_u_cla32_and11283_y0);
  and_gate and_gate_h_u_cla32_and11284_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11284_y0);
  and_gate and_gate_h_u_cla32_and11285_y0(h_u_cla32_and11284_y0, h_u_cla32_and11283_y0, h_u_cla32_and11285_y0);
  and_gate and_gate_h_u_cla32_and11286_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11286_y0);
  and_gate and_gate_h_u_cla32_and11287_y0(h_u_cla32_and11286_y0, h_u_cla32_and11285_y0, h_u_cla32_and11287_y0);
  and_gate and_gate_h_u_cla32_and11288_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11288_y0);
  and_gate and_gate_h_u_cla32_and11289_y0(h_u_cla32_and11288_y0, h_u_cla32_and11287_y0, h_u_cla32_and11289_y0);
  and_gate and_gate_h_u_cla32_and11290_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11290_y0);
  and_gate and_gate_h_u_cla32_and11291_y0(h_u_cla32_and11290_y0, h_u_cla32_and11289_y0, h_u_cla32_and11291_y0);
  and_gate and_gate_h_u_cla32_and11292_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11292_y0);
  and_gate and_gate_h_u_cla32_and11293_y0(h_u_cla32_and11292_y0, h_u_cla32_and11291_y0, h_u_cla32_and11293_y0);
  and_gate and_gate_h_u_cla32_and11294_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic18_y1, h_u_cla32_and11294_y0);
  and_gate and_gate_h_u_cla32_and11295_y0(h_u_cla32_and11294_y0, h_u_cla32_and11293_y0, h_u_cla32_and11295_y0);
  and_gate and_gate_h_u_cla32_and11296_y0(h_u_cla32_pg_logic20_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11296_y0);
  and_gate and_gate_h_u_cla32_and11297_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11297_y0);
  and_gate and_gate_h_u_cla32_and11298_y0(h_u_cla32_and11297_y0, h_u_cla32_and11296_y0, h_u_cla32_and11298_y0);
  and_gate and_gate_h_u_cla32_and11299_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11299_y0);
  and_gate and_gate_h_u_cla32_and11300_y0(h_u_cla32_and11299_y0, h_u_cla32_and11298_y0, h_u_cla32_and11300_y0);
  and_gate and_gate_h_u_cla32_and11301_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11301_y0);
  and_gate and_gate_h_u_cla32_and11302_y0(h_u_cla32_and11301_y0, h_u_cla32_and11300_y0, h_u_cla32_and11302_y0);
  and_gate and_gate_h_u_cla32_and11303_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11303_y0);
  and_gate and_gate_h_u_cla32_and11304_y0(h_u_cla32_and11303_y0, h_u_cla32_and11302_y0, h_u_cla32_and11304_y0);
  and_gate and_gate_h_u_cla32_and11305_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11305_y0);
  and_gate and_gate_h_u_cla32_and11306_y0(h_u_cla32_and11305_y0, h_u_cla32_and11304_y0, h_u_cla32_and11306_y0);
  and_gate and_gate_h_u_cla32_and11307_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11307_y0);
  and_gate and_gate_h_u_cla32_and11308_y0(h_u_cla32_and11307_y0, h_u_cla32_and11306_y0, h_u_cla32_and11308_y0);
  and_gate and_gate_h_u_cla32_and11309_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11309_y0);
  and_gate and_gate_h_u_cla32_and11310_y0(h_u_cla32_and11309_y0, h_u_cla32_and11308_y0, h_u_cla32_and11310_y0);
  and_gate and_gate_h_u_cla32_and11311_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11311_y0);
  and_gate and_gate_h_u_cla32_and11312_y0(h_u_cla32_and11311_y0, h_u_cla32_and11310_y0, h_u_cla32_and11312_y0);
  and_gate and_gate_h_u_cla32_and11313_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11313_y0);
  and_gate and_gate_h_u_cla32_and11314_y0(h_u_cla32_and11313_y0, h_u_cla32_and11312_y0, h_u_cla32_and11314_y0);
  and_gate and_gate_h_u_cla32_and11315_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11315_y0);
  and_gate and_gate_h_u_cla32_and11316_y0(h_u_cla32_and11315_y0, h_u_cla32_and11314_y0, h_u_cla32_and11316_y0);
  and_gate and_gate_h_u_cla32_and11317_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic19_y1, h_u_cla32_and11317_y0);
  and_gate and_gate_h_u_cla32_and11318_y0(h_u_cla32_and11317_y0, h_u_cla32_and11316_y0, h_u_cla32_and11318_y0);
  and_gate and_gate_h_u_cla32_and11319_y0(h_u_cla32_pg_logic21_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11319_y0);
  and_gate and_gate_h_u_cla32_and11320_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11320_y0);
  and_gate and_gate_h_u_cla32_and11321_y0(h_u_cla32_and11320_y0, h_u_cla32_and11319_y0, h_u_cla32_and11321_y0);
  and_gate and_gate_h_u_cla32_and11322_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11322_y0);
  and_gate and_gate_h_u_cla32_and11323_y0(h_u_cla32_and11322_y0, h_u_cla32_and11321_y0, h_u_cla32_and11323_y0);
  and_gate and_gate_h_u_cla32_and11324_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11324_y0);
  and_gate and_gate_h_u_cla32_and11325_y0(h_u_cla32_and11324_y0, h_u_cla32_and11323_y0, h_u_cla32_and11325_y0);
  and_gate and_gate_h_u_cla32_and11326_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11326_y0);
  and_gate and_gate_h_u_cla32_and11327_y0(h_u_cla32_and11326_y0, h_u_cla32_and11325_y0, h_u_cla32_and11327_y0);
  and_gate and_gate_h_u_cla32_and11328_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11328_y0);
  and_gate and_gate_h_u_cla32_and11329_y0(h_u_cla32_and11328_y0, h_u_cla32_and11327_y0, h_u_cla32_and11329_y0);
  and_gate and_gate_h_u_cla32_and11330_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11330_y0);
  and_gate and_gate_h_u_cla32_and11331_y0(h_u_cla32_and11330_y0, h_u_cla32_and11329_y0, h_u_cla32_and11331_y0);
  and_gate and_gate_h_u_cla32_and11332_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11332_y0);
  and_gate and_gate_h_u_cla32_and11333_y0(h_u_cla32_and11332_y0, h_u_cla32_and11331_y0, h_u_cla32_and11333_y0);
  and_gate and_gate_h_u_cla32_and11334_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11334_y0);
  and_gate and_gate_h_u_cla32_and11335_y0(h_u_cla32_and11334_y0, h_u_cla32_and11333_y0, h_u_cla32_and11335_y0);
  and_gate and_gate_h_u_cla32_and11336_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11336_y0);
  and_gate and_gate_h_u_cla32_and11337_y0(h_u_cla32_and11336_y0, h_u_cla32_and11335_y0, h_u_cla32_and11337_y0);
  and_gate and_gate_h_u_cla32_and11338_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic20_y1, h_u_cla32_and11338_y0);
  and_gate and_gate_h_u_cla32_and11339_y0(h_u_cla32_and11338_y0, h_u_cla32_and11337_y0, h_u_cla32_and11339_y0);
  and_gate and_gate_h_u_cla32_and11340_y0(h_u_cla32_pg_logic22_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11340_y0);
  and_gate and_gate_h_u_cla32_and11341_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11341_y0);
  and_gate and_gate_h_u_cla32_and11342_y0(h_u_cla32_and11341_y0, h_u_cla32_and11340_y0, h_u_cla32_and11342_y0);
  and_gate and_gate_h_u_cla32_and11343_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11343_y0);
  and_gate and_gate_h_u_cla32_and11344_y0(h_u_cla32_and11343_y0, h_u_cla32_and11342_y0, h_u_cla32_and11344_y0);
  and_gate and_gate_h_u_cla32_and11345_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11345_y0);
  and_gate and_gate_h_u_cla32_and11346_y0(h_u_cla32_and11345_y0, h_u_cla32_and11344_y0, h_u_cla32_and11346_y0);
  and_gate and_gate_h_u_cla32_and11347_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11347_y0);
  and_gate and_gate_h_u_cla32_and11348_y0(h_u_cla32_and11347_y0, h_u_cla32_and11346_y0, h_u_cla32_and11348_y0);
  and_gate and_gate_h_u_cla32_and11349_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11349_y0);
  and_gate and_gate_h_u_cla32_and11350_y0(h_u_cla32_and11349_y0, h_u_cla32_and11348_y0, h_u_cla32_and11350_y0);
  and_gate and_gate_h_u_cla32_and11351_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11351_y0);
  and_gate and_gate_h_u_cla32_and11352_y0(h_u_cla32_and11351_y0, h_u_cla32_and11350_y0, h_u_cla32_and11352_y0);
  and_gate and_gate_h_u_cla32_and11353_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11353_y0);
  and_gate and_gate_h_u_cla32_and11354_y0(h_u_cla32_and11353_y0, h_u_cla32_and11352_y0, h_u_cla32_and11354_y0);
  and_gate and_gate_h_u_cla32_and11355_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11355_y0);
  and_gate and_gate_h_u_cla32_and11356_y0(h_u_cla32_and11355_y0, h_u_cla32_and11354_y0, h_u_cla32_and11356_y0);
  and_gate and_gate_h_u_cla32_and11357_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic21_y1, h_u_cla32_and11357_y0);
  and_gate and_gate_h_u_cla32_and11358_y0(h_u_cla32_and11357_y0, h_u_cla32_and11356_y0, h_u_cla32_and11358_y0);
  and_gate and_gate_h_u_cla32_and11359_y0(h_u_cla32_pg_logic23_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11359_y0);
  and_gate and_gate_h_u_cla32_and11360_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11360_y0);
  and_gate and_gate_h_u_cla32_and11361_y0(h_u_cla32_and11360_y0, h_u_cla32_and11359_y0, h_u_cla32_and11361_y0);
  and_gate and_gate_h_u_cla32_and11362_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11362_y0);
  and_gate and_gate_h_u_cla32_and11363_y0(h_u_cla32_and11362_y0, h_u_cla32_and11361_y0, h_u_cla32_and11363_y0);
  and_gate and_gate_h_u_cla32_and11364_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11364_y0);
  and_gate and_gate_h_u_cla32_and11365_y0(h_u_cla32_and11364_y0, h_u_cla32_and11363_y0, h_u_cla32_and11365_y0);
  and_gate and_gate_h_u_cla32_and11366_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11366_y0);
  and_gate and_gate_h_u_cla32_and11367_y0(h_u_cla32_and11366_y0, h_u_cla32_and11365_y0, h_u_cla32_and11367_y0);
  and_gate and_gate_h_u_cla32_and11368_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11368_y0);
  and_gate and_gate_h_u_cla32_and11369_y0(h_u_cla32_and11368_y0, h_u_cla32_and11367_y0, h_u_cla32_and11369_y0);
  and_gate and_gate_h_u_cla32_and11370_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11370_y0);
  and_gate and_gate_h_u_cla32_and11371_y0(h_u_cla32_and11370_y0, h_u_cla32_and11369_y0, h_u_cla32_and11371_y0);
  and_gate and_gate_h_u_cla32_and11372_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11372_y0);
  and_gate and_gate_h_u_cla32_and11373_y0(h_u_cla32_and11372_y0, h_u_cla32_and11371_y0, h_u_cla32_and11373_y0);
  and_gate and_gate_h_u_cla32_and11374_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic22_y1, h_u_cla32_and11374_y0);
  and_gate and_gate_h_u_cla32_and11375_y0(h_u_cla32_and11374_y0, h_u_cla32_and11373_y0, h_u_cla32_and11375_y0);
  and_gate and_gate_h_u_cla32_and11376_y0(h_u_cla32_pg_logic24_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11376_y0);
  and_gate and_gate_h_u_cla32_and11377_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11377_y0);
  and_gate and_gate_h_u_cla32_and11378_y0(h_u_cla32_and11377_y0, h_u_cla32_and11376_y0, h_u_cla32_and11378_y0);
  and_gate and_gate_h_u_cla32_and11379_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11379_y0);
  and_gate and_gate_h_u_cla32_and11380_y0(h_u_cla32_and11379_y0, h_u_cla32_and11378_y0, h_u_cla32_and11380_y0);
  and_gate and_gate_h_u_cla32_and11381_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11381_y0);
  and_gate and_gate_h_u_cla32_and11382_y0(h_u_cla32_and11381_y0, h_u_cla32_and11380_y0, h_u_cla32_and11382_y0);
  and_gate and_gate_h_u_cla32_and11383_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11383_y0);
  and_gate and_gate_h_u_cla32_and11384_y0(h_u_cla32_and11383_y0, h_u_cla32_and11382_y0, h_u_cla32_and11384_y0);
  and_gate and_gate_h_u_cla32_and11385_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11385_y0);
  and_gate and_gate_h_u_cla32_and11386_y0(h_u_cla32_and11385_y0, h_u_cla32_and11384_y0, h_u_cla32_and11386_y0);
  and_gate and_gate_h_u_cla32_and11387_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11387_y0);
  and_gate and_gate_h_u_cla32_and11388_y0(h_u_cla32_and11387_y0, h_u_cla32_and11386_y0, h_u_cla32_and11388_y0);
  and_gate and_gate_h_u_cla32_and11389_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic23_y1, h_u_cla32_and11389_y0);
  and_gate and_gate_h_u_cla32_and11390_y0(h_u_cla32_and11389_y0, h_u_cla32_and11388_y0, h_u_cla32_and11390_y0);
  and_gate and_gate_h_u_cla32_and11391_y0(h_u_cla32_pg_logic25_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11391_y0);
  and_gate and_gate_h_u_cla32_and11392_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11392_y0);
  and_gate and_gate_h_u_cla32_and11393_y0(h_u_cla32_and11392_y0, h_u_cla32_and11391_y0, h_u_cla32_and11393_y0);
  and_gate and_gate_h_u_cla32_and11394_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11394_y0);
  and_gate and_gate_h_u_cla32_and11395_y0(h_u_cla32_and11394_y0, h_u_cla32_and11393_y0, h_u_cla32_and11395_y0);
  and_gate and_gate_h_u_cla32_and11396_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11396_y0);
  and_gate and_gate_h_u_cla32_and11397_y0(h_u_cla32_and11396_y0, h_u_cla32_and11395_y0, h_u_cla32_and11397_y0);
  and_gate and_gate_h_u_cla32_and11398_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11398_y0);
  and_gate and_gate_h_u_cla32_and11399_y0(h_u_cla32_and11398_y0, h_u_cla32_and11397_y0, h_u_cla32_and11399_y0);
  and_gate and_gate_h_u_cla32_and11400_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11400_y0);
  and_gate and_gate_h_u_cla32_and11401_y0(h_u_cla32_and11400_y0, h_u_cla32_and11399_y0, h_u_cla32_and11401_y0);
  and_gate and_gate_h_u_cla32_and11402_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic24_y1, h_u_cla32_and11402_y0);
  and_gate and_gate_h_u_cla32_and11403_y0(h_u_cla32_and11402_y0, h_u_cla32_and11401_y0, h_u_cla32_and11403_y0);
  and_gate and_gate_h_u_cla32_and11404_y0(h_u_cla32_pg_logic26_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and11404_y0);
  and_gate and_gate_h_u_cla32_and11405_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and11405_y0);
  and_gate and_gate_h_u_cla32_and11406_y0(h_u_cla32_and11405_y0, h_u_cla32_and11404_y0, h_u_cla32_and11406_y0);
  and_gate and_gate_h_u_cla32_and11407_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and11407_y0);
  and_gate and_gate_h_u_cla32_and11408_y0(h_u_cla32_and11407_y0, h_u_cla32_and11406_y0, h_u_cla32_and11408_y0);
  and_gate and_gate_h_u_cla32_and11409_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and11409_y0);
  and_gate and_gate_h_u_cla32_and11410_y0(h_u_cla32_and11409_y0, h_u_cla32_and11408_y0, h_u_cla32_and11410_y0);
  and_gate and_gate_h_u_cla32_and11411_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and11411_y0);
  and_gate and_gate_h_u_cla32_and11412_y0(h_u_cla32_and11411_y0, h_u_cla32_and11410_y0, h_u_cla32_and11412_y0);
  and_gate and_gate_h_u_cla32_and11413_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic25_y1, h_u_cla32_and11413_y0);
  and_gate and_gate_h_u_cla32_and11414_y0(h_u_cla32_and11413_y0, h_u_cla32_and11412_y0, h_u_cla32_and11414_y0);
  and_gate and_gate_h_u_cla32_and11415_y0(h_u_cla32_pg_logic27_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and11415_y0);
  and_gate and_gate_h_u_cla32_and11416_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and11416_y0);
  and_gate and_gate_h_u_cla32_and11417_y0(h_u_cla32_and11416_y0, h_u_cla32_and11415_y0, h_u_cla32_and11417_y0);
  and_gate and_gate_h_u_cla32_and11418_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and11418_y0);
  and_gate and_gate_h_u_cla32_and11419_y0(h_u_cla32_and11418_y0, h_u_cla32_and11417_y0, h_u_cla32_and11419_y0);
  and_gate and_gate_h_u_cla32_and11420_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and11420_y0);
  and_gate and_gate_h_u_cla32_and11421_y0(h_u_cla32_and11420_y0, h_u_cla32_and11419_y0, h_u_cla32_and11421_y0);
  and_gate and_gate_h_u_cla32_and11422_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic26_y1, h_u_cla32_and11422_y0);
  and_gate and_gate_h_u_cla32_and11423_y0(h_u_cla32_and11422_y0, h_u_cla32_and11421_y0, h_u_cla32_and11423_y0);
  and_gate and_gate_h_u_cla32_and11424_y0(h_u_cla32_pg_logic28_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and11424_y0);
  and_gate and_gate_h_u_cla32_and11425_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and11425_y0);
  and_gate and_gate_h_u_cla32_and11426_y0(h_u_cla32_and11425_y0, h_u_cla32_and11424_y0, h_u_cla32_and11426_y0);
  and_gate and_gate_h_u_cla32_and11427_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and11427_y0);
  and_gate and_gate_h_u_cla32_and11428_y0(h_u_cla32_and11427_y0, h_u_cla32_and11426_y0, h_u_cla32_and11428_y0);
  and_gate and_gate_h_u_cla32_and11429_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic27_y1, h_u_cla32_and11429_y0);
  and_gate and_gate_h_u_cla32_and11430_y0(h_u_cla32_and11429_y0, h_u_cla32_and11428_y0, h_u_cla32_and11430_y0);
  and_gate and_gate_h_u_cla32_and11431_y0(h_u_cla32_pg_logic29_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_and11431_y0);
  and_gate and_gate_h_u_cla32_and11432_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_and11432_y0);
  and_gate and_gate_h_u_cla32_and11433_y0(h_u_cla32_and11432_y0, h_u_cla32_and11431_y0, h_u_cla32_and11433_y0);
  and_gate and_gate_h_u_cla32_and11434_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic28_y1, h_u_cla32_and11434_y0);
  and_gate and_gate_h_u_cla32_and11435_y0(h_u_cla32_and11434_y0, h_u_cla32_and11433_y0, h_u_cla32_and11435_y0);
  and_gate and_gate_h_u_cla32_and11436_y0(h_u_cla32_pg_logic30_y0, h_u_cla32_pg_logic29_y1, h_u_cla32_and11436_y0);
  and_gate and_gate_h_u_cla32_and11437_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic29_y1, h_u_cla32_and11437_y0);
  and_gate and_gate_h_u_cla32_and11438_y0(h_u_cla32_and11437_y0, h_u_cla32_and11436_y0, h_u_cla32_and11438_y0);
  and_gate and_gate_h_u_cla32_and11439_y0(h_u_cla32_pg_logic31_y0, h_u_cla32_pg_logic30_y1, h_u_cla32_and11439_y0);
  or_gate or_gate_h_u_cla32_or496_y0(h_u_cla32_and11439_y0, h_u_cla32_and10478_y0, h_u_cla32_or496_y0);
  or_gate or_gate_h_u_cla32_or497_y0(h_u_cla32_or496_y0, h_u_cla32_and10539_y0, h_u_cla32_or497_y0);
  or_gate or_gate_h_u_cla32_or498_y0(h_u_cla32_or497_y0, h_u_cla32_and10598_y0, h_u_cla32_or498_y0);
  or_gate or_gate_h_u_cla32_or499_y0(h_u_cla32_or498_y0, h_u_cla32_and10655_y0, h_u_cla32_or499_y0);
  or_gate or_gate_h_u_cla32_or500_y0(h_u_cla32_or499_y0, h_u_cla32_and10710_y0, h_u_cla32_or500_y0);
  or_gate or_gate_h_u_cla32_or501_y0(h_u_cla32_or500_y0, h_u_cla32_and10763_y0, h_u_cla32_or501_y0);
  or_gate or_gate_h_u_cla32_or502_y0(h_u_cla32_or501_y0, h_u_cla32_and10814_y0, h_u_cla32_or502_y0);
  or_gate or_gate_h_u_cla32_or503_y0(h_u_cla32_or502_y0, h_u_cla32_and10863_y0, h_u_cla32_or503_y0);
  or_gate or_gate_h_u_cla32_or504_y0(h_u_cla32_or503_y0, h_u_cla32_and10910_y0, h_u_cla32_or504_y0);
  or_gate or_gate_h_u_cla32_or505_y0(h_u_cla32_or504_y0, h_u_cla32_and10955_y0, h_u_cla32_or505_y0);
  or_gate or_gate_h_u_cla32_or506_y0(h_u_cla32_or505_y0, h_u_cla32_and10998_y0, h_u_cla32_or506_y0);
  or_gate or_gate_h_u_cla32_or507_y0(h_u_cla32_or506_y0, h_u_cla32_and11039_y0, h_u_cla32_or507_y0);
  or_gate or_gate_h_u_cla32_or508_y0(h_u_cla32_or507_y0, h_u_cla32_and11078_y0, h_u_cla32_or508_y0);
  or_gate or_gate_h_u_cla32_or509_y0(h_u_cla32_or508_y0, h_u_cla32_and11115_y0, h_u_cla32_or509_y0);
  or_gate or_gate_h_u_cla32_or510_y0(h_u_cla32_or509_y0, h_u_cla32_and11150_y0, h_u_cla32_or510_y0);
  or_gate or_gate_h_u_cla32_or511_y0(h_u_cla32_or510_y0, h_u_cla32_and11183_y0, h_u_cla32_or511_y0);
  or_gate or_gate_h_u_cla32_or512_y0(h_u_cla32_or511_y0, h_u_cla32_and11214_y0, h_u_cla32_or512_y0);
  or_gate or_gate_h_u_cla32_or513_y0(h_u_cla32_or512_y0, h_u_cla32_and11243_y0, h_u_cla32_or513_y0);
  or_gate or_gate_h_u_cla32_or514_y0(h_u_cla32_or513_y0, h_u_cla32_and11270_y0, h_u_cla32_or514_y0);
  or_gate or_gate_h_u_cla32_or515_y0(h_u_cla32_or514_y0, h_u_cla32_and11295_y0, h_u_cla32_or515_y0);
  or_gate or_gate_h_u_cla32_or516_y0(h_u_cla32_or515_y0, h_u_cla32_and11318_y0, h_u_cla32_or516_y0);
  or_gate or_gate_h_u_cla32_or517_y0(h_u_cla32_or516_y0, h_u_cla32_and11339_y0, h_u_cla32_or517_y0);
  or_gate or_gate_h_u_cla32_or518_y0(h_u_cla32_or517_y0, h_u_cla32_and11358_y0, h_u_cla32_or518_y0);
  or_gate or_gate_h_u_cla32_or519_y0(h_u_cla32_or518_y0, h_u_cla32_and11375_y0, h_u_cla32_or519_y0);
  or_gate or_gate_h_u_cla32_or520_y0(h_u_cla32_or519_y0, h_u_cla32_and11390_y0, h_u_cla32_or520_y0);
  or_gate or_gate_h_u_cla32_or521_y0(h_u_cla32_or520_y0, h_u_cla32_and11403_y0, h_u_cla32_or521_y0);
  or_gate or_gate_h_u_cla32_or522_y0(h_u_cla32_or521_y0, h_u_cla32_and11414_y0, h_u_cla32_or522_y0);
  or_gate or_gate_h_u_cla32_or523_y0(h_u_cla32_or522_y0, h_u_cla32_and11423_y0, h_u_cla32_or523_y0);
  or_gate or_gate_h_u_cla32_or524_y0(h_u_cla32_or523_y0, h_u_cla32_and11430_y0, h_u_cla32_or524_y0);
  or_gate or_gate_h_u_cla32_or525_y0(h_u_cla32_or524_y0, h_u_cla32_and11435_y0, h_u_cla32_or525_y0);
  or_gate or_gate_h_u_cla32_or526_y0(h_u_cla32_or525_y0, h_u_cla32_and11438_y0, h_u_cla32_or526_y0);
  or_gate or_gate_h_u_cla32_or527_y0(h_u_cla32_pg_logic31_y1, h_u_cla32_or526_y0, h_u_cla32_or527_y0);

  assign out[0] = h_u_cla32_xor0_y0;
  assign out[1] = h_u_cla32_xor1_y0;
  assign out[2] = h_u_cla32_xor2_y0;
  assign out[3] = h_u_cla32_xor3_y0;
  assign out[4] = h_u_cla32_xor4_y0;
  assign out[5] = h_u_cla32_xor5_y0;
  assign out[6] = h_u_cla32_xor6_y0;
  assign out[7] = h_u_cla32_xor7_y0;
  assign out[8] = h_u_cla32_xor8_y0;
  assign out[9] = h_u_cla32_xor9_y0;
  assign out[10] = h_u_cla32_xor10_y0;
  assign out[11] = h_u_cla32_xor11_y0;
  assign out[12] = h_u_cla32_xor12_y0;
  assign out[13] = h_u_cla32_xor13_y0;
  assign out[14] = h_u_cla32_xor14_y0;
  assign out[15] = h_u_cla32_xor15_y0;
  assign out[16] = h_u_cla32_xor16_y0;
  assign out[17] = h_u_cla32_xor17_y0;
  assign out[18] = h_u_cla32_xor18_y0;
  assign out[19] = h_u_cla32_xor19_y0;
  assign out[20] = h_u_cla32_xor20_y0;
  assign out[21] = h_u_cla32_xor21_y0;
  assign out[22] = h_u_cla32_xor22_y0;
  assign out[23] = h_u_cla32_xor23_y0;
  assign out[24] = h_u_cla32_xor24_y0;
  assign out[25] = h_u_cla32_xor25_y0;
  assign out[26] = h_u_cla32_xor26_y0;
  assign out[27] = h_u_cla32_xor27_y0;
  assign out[28] = h_u_cla32_xor28_y0;
  assign out[29] = h_u_cla32_xor29_y0;
  assign out[30] = h_u_cla32_xor30_y0;
  assign out[31] = h_u_cla32_xor31_y0;
  assign out[32] = h_u_cla32_or527_y0;
endmodule