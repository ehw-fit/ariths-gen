module s_cla24(input [23:0] a, input [23:0] b, output [24:0] s_cla24_out);
  wire s_cla24_pg_logic0_or0;
  wire s_cla24_pg_logic0_and0;
  wire s_cla24_pg_logic0_xor0;
  wire s_cla24_pg_logic1_or0;
  wire s_cla24_pg_logic1_and0;
  wire s_cla24_pg_logic1_xor0;
  wire s_cla24_xor1;
  wire s_cla24_and0;
  wire s_cla24_or0;
  wire s_cla24_pg_logic2_or0;
  wire s_cla24_pg_logic2_and0;
  wire s_cla24_pg_logic2_xor0;
  wire s_cla24_xor2;
  wire s_cla24_and1;
  wire s_cla24_and2;
  wire s_cla24_and3;
  wire s_cla24_and4;
  wire s_cla24_or1;
  wire s_cla24_or2;
  wire s_cla24_pg_logic3_or0;
  wire s_cla24_pg_logic3_and0;
  wire s_cla24_pg_logic3_xor0;
  wire s_cla24_xor3;
  wire s_cla24_and5;
  wire s_cla24_and6;
  wire s_cla24_and7;
  wire s_cla24_and8;
  wire s_cla24_and9;
  wire s_cla24_and10;
  wire s_cla24_and11;
  wire s_cla24_or3;
  wire s_cla24_or4;
  wire s_cla24_or5;
  wire s_cla24_pg_logic4_or0;
  wire s_cla24_pg_logic4_and0;
  wire s_cla24_pg_logic4_xor0;
  wire s_cla24_xor4;
  wire s_cla24_and12;
  wire s_cla24_or6;
  wire s_cla24_pg_logic5_or0;
  wire s_cla24_pg_logic5_and0;
  wire s_cla24_pg_logic5_xor0;
  wire s_cla24_xor5;
  wire s_cla24_and13;
  wire s_cla24_and14;
  wire s_cla24_and15;
  wire s_cla24_or7;
  wire s_cla24_or8;
  wire s_cla24_pg_logic6_or0;
  wire s_cla24_pg_logic6_and0;
  wire s_cla24_pg_logic6_xor0;
  wire s_cla24_xor6;
  wire s_cla24_and16;
  wire s_cla24_and17;
  wire s_cla24_and18;
  wire s_cla24_and19;
  wire s_cla24_and20;
  wire s_cla24_and21;
  wire s_cla24_or9;
  wire s_cla24_or10;
  wire s_cla24_or11;
  wire s_cla24_pg_logic7_or0;
  wire s_cla24_pg_logic7_and0;
  wire s_cla24_pg_logic7_xor0;
  wire s_cla24_xor7;
  wire s_cla24_and22;
  wire s_cla24_and23;
  wire s_cla24_and24;
  wire s_cla24_and25;
  wire s_cla24_and26;
  wire s_cla24_and27;
  wire s_cla24_and28;
  wire s_cla24_and29;
  wire s_cla24_and30;
  wire s_cla24_and31;
  wire s_cla24_or12;
  wire s_cla24_or13;
  wire s_cla24_or14;
  wire s_cla24_or15;
  wire s_cla24_pg_logic8_or0;
  wire s_cla24_pg_logic8_and0;
  wire s_cla24_pg_logic8_xor0;
  wire s_cla24_xor8;
  wire s_cla24_and32;
  wire s_cla24_or16;
  wire s_cla24_pg_logic9_or0;
  wire s_cla24_pg_logic9_and0;
  wire s_cla24_pg_logic9_xor0;
  wire s_cla24_xor9;
  wire s_cla24_and33;
  wire s_cla24_and34;
  wire s_cla24_and35;
  wire s_cla24_or17;
  wire s_cla24_or18;
  wire s_cla24_pg_logic10_or0;
  wire s_cla24_pg_logic10_and0;
  wire s_cla24_pg_logic10_xor0;
  wire s_cla24_xor10;
  wire s_cla24_and36;
  wire s_cla24_and37;
  wire s_cla24_and38;
  wire s_cla24_and39;
  wire s_cla24_and40;
  wire s_cla24_and41;
  wire s_cla24_or19;
  wire s_cla24_or20;
  wire s_cla24_or21;
  wire s_cla24_pg_logic11_or0;
  wire s_cla24_pg_logic11_and0;
  wire s_cla24_pg_logic11_xor0;
  wire s_cla24_xor11;
  wire s_cla24_and42;
  wire s_cla24_and43;
  wire s_cla24_and44;
  wire s_cla24_and45;
  wire s_cla24_and46;
  wire s_cla24_and47;
  wire s_cla24_and48;
  wire s_cla24_and49;
  wire s_cla24_and50;
  wire s_cla24_and51;
  wire s_cla24_or22;
  wire s_cla24_or23;
  wire s_cla24_or24;
  wire s_cla24_or25;
  wire s_cla24_pg_logic12_or0;
  wire s_cla24_pg_logic12_and0;
  wire s_cla24_pg_logic12_xor0;
  wire s_cla24_xor12;
  wire s_cla24_and52;
  wire s_cla24_or26;
  wire s_cla24_pg_logic13_or0;
  wire s_cla24_pg_logic13_and0;
  wire s_cla24_pg_logic13_xor0;
  wire s_cla24_xor13;
  wire s_cla24_and53;
  wire s_cla24_and54;
  wire s_cla24_and55;
  wire s_cla24_or27;
  wire s_cla24_or28;
  wire s_cla24_pg_logic14_or0;
  wire s_cla24_pg_logic14_and0;
  wire s_cla24_pg_logic14_xor0;
  wire s_cla24_xor14;
  wire s_cla24_and56;
  wire s_cla24_and57;
  wire s_cla24_and58;
  wire s_cla24_and59;
  wire s_cla24_and60;
  wire s_cla24_and61;
  wire s_cla24_or29;
  wire s_cla24_or30;
  wire s_cla24_or31;
  wire s_cla24_pg_logic15_or0;
  wire s_cla24_pg_logic15_and0;
  wire s_cla24_pg_logic15_xor0;
  wire s_cla24_xor15;
  wire s_cla24_and62;
  wire s_cla24_and63;
  wire s_cla24_and64;
  wire s_cla24_and65;
  wire s_cla24_and66;
  wire s_cla24_and67;
  wire s_cla24_and68;
  wire s_cla24_and69;
  wire s_cla24_and70;
  wire s_cla24_and71;
  wire s_cla24_or32;
  wire s_cla24_or33;
  wire s_cla24_or34;
  wire s_cla24_or35;
  wire s_cla24_pg_logic16_or0;
  wire s_cla24_pg_logic16_and0;
  wire s_cla24_pg_logic16_xor0;
  wire s_cla24_xor16;
  wire s_cla24_and72;
  wire s_cla24_or36;
  wire s_cla24_pg_logic17_or0;
  wire s_cla24_pg_logic17_and0;
  wire s_cla24_pg_logic17_xor0;
  wire s_cla24_xor17;
  wire s_cla24_and73;
  wire s_cla24_and74;
  wire s_cla24_and75;
  wire s_cla24_or37;
  wire s_cla24_or38;
  wire s_cla24_pg_logic18_or0;
  wire s_cla24_pg_logic18_and0;
  wire s_cla24_pg_logic18_xor0;
  wire s_cla24_xor18;
  wire s_cla24_and76;
  wire s_cla24_and77;
  wire s_cla24_and78;
  wire s_cla24_and79;
  wire s_cla24_and80;
  wire s_cla24_and81;
  wire s_cla24_or39;
  wire s_cla24_or40;
  wire s_cla24_or41;
  wire s_cla24_pg_logic19_or0;
  wire s_cla24_pg_logic19_and0;
  wire s_cla24_pg_logic19_xor0;
  wire s_cla24_xor19;
  wire s_cla24_and82;
  wire s_cla24_and83;
  wire s_cla24_and84;
  wire s_cla24_and85;
  wire s_cla24_and86;
  wire s_cla24_and87;
  wire s_cla24_and88;
  wire s_cla24_and89;
  wire s_cla24_and90;
  wire s_cla24_and91;
  wire s_cla24_or42;
  wire s_cla24_or43;
  wire s_cla24_or44;
  wire s_cla24_or45;
  wire s_cla24_pg_logic20_or0;
  wire s_cla24_pg_logic20_and0;
  wire s_cla24_pg_logic20_xor0;
  wire s_cla24_xor20;
  wire s_cla24_and92;
  wire s_cla24_or46;
  wire s_cla24_pg_logic21_or0;
  wire s_cla24_pg_logic21_and0;
  wire s_cla24_pg_logic21_xor0;
  wire s_cla24_xor21;
  wire s_cla24_and93;
  wire s_cla24_and94;
  wire s_cla24_and95;
  wire s_cla24_or47;
  wire s_cla24_or48;
  wire s_cla24_pg_logic22_or0;
  wire s_cla24_pg_logic22_and0;
  wire s_cla24_pg_logic22_xor0;
  wire s_cla24_xor22;
  wire s_cla24_and96;
  wire s_cla24_and97;
  wire s_cla24_and98;
  wire s_cla24_and99;
  wire s_cla24_and100;
  wire s_cla24_and101;
  wire s_cla24_or49;
  wire s_cla24_or50;
  wire s_cla24_or51;
  wire s_cla24_pg_logic23_or0;
  wire s_cla24_pg_logic23_and0;
  wire s_cla24_pg_logic23_xor0;
  wire s_cla24_xor23;
  wire s_cla24_and102;
  wire s_cla24_and103;
  wire s_cla24_and104;
  wire s_cla24_and105;
  wire s_cla24_and106;
  wire s_cla24_and107;
  wire s_cla24_and108;
  wire s_cla24_and109;
  wire s_cla24_and110;
  wire s_cla24_and111;
  wire s_cla24_or52;
  wire s_cla24_or53;
  wire s_cla24_or54;
  wire s_cla24_or55;
  wire s_cla24_xor24;
  wire s_cla24_xor25;

  assign s_cla24_pg_logic0_or0 = a[0] | b[0];
  assign s_cla24_pg_logic0_and0 = a[0] & b[0];
  assign s_cla24_pg_logic0_xor0 = a[0] ^ b[0];
  assign s_cla24_pg_logic1_or0 = a[1] | b[1];
  assign s_cla24_pg_logic1_and0 = a[1] & b[1];
  assign s_cla24_pg_logic1_xor0 = a[1] ^ b[1];
  assign s_cla24_xor1 = s_cla24_pg_logic1_xor0 ^ s_cla24_pg_logic0_and0;
  assign s_cla24_and0 = s_cla24_pg_logic0_and0 & s_cla24_pg_logic1_or0;
  assign s_cla24_or0 = s_cla24_pg_logic1_and0 | s_cla24_and0;
  assign s_cla24_pg_logic2_or0 = a[2] | b[2];
  assign s_cla24_pg_logic2_and0 = a[2] & b[2];
  assign s_cla24_pg_logic2_xor0 = a[2] ^ b[2];
  assign s_cla24_xor2 = s_cla24_pg_logic2_xor0 ^ s_cla24_or0;
  assign s_cla24_and1 = s_cla24_pg_logic2_or0 & s_cla24_pg_logic0_or0;
  assign s_cla24_and2 = s_cla24_pg_logic0_and0 & s_cla24_pg_logic2_or0;
  assign s_cla24_and3 = s_cla24_and2 & s_cla24_pg_logic1_or0;
  assign s_cla24_and4 = s_cla24_pg_logic1_and0 & s_cla24_pg_logic2_or0;
  assign s_cla24_or1 = s_cla24_and3 | s_cla24_and4;
  assign s_cla24_or2 = s_cla24_pg_logic2_and0 | s_cla24_or1;
  assign s_cla24_pg_logic3_or0 = a[3] | b[3];
  assign s_cla24_pg_logic3_and0 = a[3] & b[3];
  assign s_cla24_pg_logic3_xor0 = a[3] ^ b[3];
  assign s_cla24_xor3 = s_cla24_pg_logic3_xor0 ^ s_cla24_or2;
  assign s_cla24_and5 = s_cla24_pg_logic3_or0 & s_cla24_pg_logic1_or0;
  assign s_cla24_and6 = s_cla24_pg_logic0_and0 & s_cla24_pg_logic2_or0;
  assign s_cla24_and7 = s_cla24_pg_logic3_or0 & s_cla24_pg_logic1_or0;
  assign s_cla24_and8 = s_cla24_and6 & s_cla24_and7;
  assign s_cla24_and9 = s_cla24_pg_logic1_and0 & s_cla24_pg_logic3_or0;
  assign s_cla24_and10 = s_cla24_and9 & s_cla24_pg_logic2_or0;
  assign s_cla24_and11 = s_cla24_pg_logic2_and0 & s_cla24_pg_logic3_or0;
  assign s_cla24_or3 = s_cla24_and8 | s_cla24_and11;
  assign s_cla24_or4 = s_cla24_and10 | s_cla24_or3;
  assign s_cla24_or5 = s_cla24_pg_logic3_and0 | s_cla24_or4;
  assign s_cla24_pg_logic4_or0 = a[4] | b[4];
  assign s_cla24_pg_logic4_and0 = a[4] & b[4];
  assign s_cla24_pg_logic4_xor0 = a[4] ^ b[4];
  assign s_cla24_xor4 = s_cla24_pg_logic4_xor0 ^ s_cla24_or5;
  assign s_cla24_and12 = s_cla24_or5 & s_cla24_pg_logic4_or0;
  assign s_cla24_or6 = s_cla24_pg_logic4_and0 | s_cla24_and12;
  assign s_cla24_pg_logic5_or0 = a[5] | b[5];
  assign s_cla24_pg_logic5_and0 = a[5] & b[5];
  assign s_cla24_pg_logic5_xor0 = a[5] ^ b[5];
  assign s_cla24_xor5 = s_cla24_pg_logic5_xor0 ^ s_cla24_or6;
  assign s_cla24_and13 = s_cla24_or5 & s_cla24_pg_logic5_or0;
  assign s_cla24_and14 = s_cla24_and13 & s_cla24_pg_logic4_or0;
  assign s_cla24_and15 = s_cla24_pg_logic4_and0 & s_cla24_pg_logic5_or0;
  assign s_cla24_or7 = s_cla24_and14 | s_cla24_and15;
  assign s_cla24_or8 = s_cla24_pg_logic5_and0 | s_cla24_or7;
  assign s_cla24_pg_logic6_or0 = a[6] | b[6];
  assign s_cla24_pg_logic6_and0 = a[6] & b[6];
  assign s_cla24_pg_logic6_xor0 = a[6] ^ b[6];
  assign s_cla24_xor6 = s_cla24_pg_logic6_xor0 ^ s_cla24_or8;
  assign s_cla24_and16 = s_cla24_or5 & s_cla24_pg_logic5_or0;
  assign s_cla24_and17 = s_cla24_pg_logic6_or0 & s_cla24_pg_logic4_or0;
  assign s_cla24_and18 = s_cla24_and16 & s_cla24_and17;
  assign s_cla24_and19 = s_cla24_pg_logic4_and0 & s_cla24_pg_logic6_or0;
  assign s_cla24_and20 = s_cla24_and19 & s_cla24_pg_logic5_or0;
  assign s_cla24_and21 = s_cla24_pg_logic5_and0 & s_cla24_pg_logic6_or0;
  assign s_cla24_or9 = s_cla24_and18 | s_cla24_and20;
  assign s_cla24_or10 = s_cla24_or9 | s_cla24_and21;
  assign s_cla24_or11 = s_cla24_pg_logic6_and0 | s_cla24_or10;
  assign s_cla24_pg_logic7_or0 = a[7] | b[7];
  assign s_cla24_pg_logic7_and0 = a[7] & b[7];
  assign s_cla24_pg_logic7_xor0 = a[7] ^ b[7];
  assign s_cla24_xor7 = s_cla24_pg_logic7_xor0 ^ s_cla24_or11;
  assign s_cla24_and22 = s_cla24_or5 & s_cla24_pg_logic6_or0;
  assign s_cla24_and23 = s_cla24_pg_logic7_or0 & s_cla24_pg_logic5_or0;
  assign s_cla24_and24 = s_cla24_and22 & s_cla24_and23;
  assign s_cla24_and25 = s_cla24_and24 & s_cla24_pg_logic4_or0;
  assign s_cla24_and26 = s_cla24_pg_logic4_and0 & s_cla24_pg_logic6_or0;
  assign s_cla24_and27 = s_cla24_pg_logic7_or0 & s_cla24_pg_logic5_or0;
  assign s_cla24_and28 = s_cla24_and26 & s_cla24_and27;
  assign s_cla24_and29 = s_cla24_pg_logic5_and0 & s_cla24_pg_logic7_or0;
  assign s_cla24_and30 = s_cla24_and29 & s_cla24_pg_logic6_or0;
  assign s_cla24_and31 = s_cla24_pg_logic6_and0 & s_cla24_pg_logic7_or0;
  assign s_cla24_or12 = s_cla24_and25 | s_cla24_and30;
  assign s_cla24_or13 = s_cla24_and28 | s_cla24_and31;
  assign s_cla24_or14 = s_cla24_or12 | s_cla24_or13;
  assign s_cla24_or15 = s_cla24_pg_logic7_and0 | s_cla24_or14;
  assign s_cla24_pg_logic8_or0 = a[8] | b[8];
  assign s_cla24_pg_logic8_and0 = a[8] & b[8];
  assign s_cla24_pg_logic8_xor0 = a[8] ^ b[8];
  assign s_cla24_xor8 = s_cla24_pg_logic8_xor0 ^ s_cla24_or15;
  assign s_cla24_and32 = s_cla24_or15 & s_cla24_pg_logic8_or0;
  assign s_cla24_or16 = s_cla24_pg_logic8_and0 | s_cla24_and32;
  assign s_cla24_pg_logic9_or0 = a[9] | b[9];
  assign s_cla24_pg_logic9_and0 = a[9] & b[9];
  assign s_cla24_pg_logic9_xor0 = a[9] ^ b[9];
  assign s_cla24_xor9 = s_cla24_pg_logic9_xor0 ^ s_cla24_or16;
  assign s_cla24_and33 = s_cla24_or15 & s_cla24_pg_logic9_or0;
  assign s_cla24_and34 = s_cla24_and33 & s_cla24_pg_logic8_or0;
  assign s_cla24_and35 = s_cla24_pg_logic8_and0 & s_cla24_pg_logic9_or0;
  assign s_cla24_or17 = s_cla24_and34 | s_cla24_and35;
  assign s_cla24_or18 = s_cla24_pg_logic9_and0 | s_cla24_or17;
  assign s_cla24_pg_logic10_or0 = a[10] | b[10];
  assign s_cla24_pg_logic10_and0 = a[10] & b[10];
  assign s_cla24_pg_logic10_xor0 = a[10] ^ b[10];
  assign s_cla24_xor10 = s_cla24_pg_logic10_xor0 ^ s_cla24_or18;
  assign s_cla24_and36 = s_cla24_or15 & s_cla24_pg_logic9_or0;
  assign s_cla24_and37 = s_cla24_pg_logic10_or0 & s_cla24_pg_logic8_or0;
  assign s_cla24_and38 = s_cla24_and36 & s_cla24_and37;
  assign s_cla24_and39 = s_cla24_pg_logic8_and0 & s_cla24_pg_logic10_or0;
  assign s_cla24_and40 = s_cla24_and39 & s_cla24_pg_logic9_or0;
  assign s_cla24_and41 = s_cla24_pg_logic9_and0 & s_cla24_pg_logic10_or0;
  assign s_cla24_or19 = s_cla24_and38 | s_cla24_and40;
  assign s_cla24_or20 = s_cla24_or19 | s_cla24_and41;
  assign s_cla24_or21 = s_cla24_pg_logic10_and0 | s_cla24_or20;
  assign s_cla24_pg_logic11_or0 = a[11] | b[11];
  assign s_cla24_pg_logic11_and0 = a[11] & b[11];
  assign s_cla24_pg_logic11_xor0 = a[11] ^ b[11];
  assign s_cla24_xor11 = s_cla24_pg_logic11_xor0 ^ s_cla24_or21;
  assign s_cla24_and42 = s_cla24_or15 & s_cla24_pg_logic10_or0;
  assign s_cla24_and43 = s_cla24_pg_logic11_or0 & s_cla24_pg_logic9_or0;
  assign s_cla24_and44 = s_cla24_and42 & s_cla24_and43;
  assign s_cla24_and45 = s_cla24_and44 & s_cla24_pg_logic8_or0;
  assign s_cla24_and46 = s_cla24_pg_logic8_and0 & s_cla24_pg_logic10_or0;
  assign s_cla24_and47 = s_cla24_pg_logic11_or0 & s_cla24_pg_logic9_or0;
  assign s_cla24_and48 = s_cla24_and46 & s_cla24_and47;
  assign s_cla24_and49 = s_cla24_pg_logic9_and0 & s_cla24_pg_logic11_or0;
  assign s_cla24_and50 = s_cla24_and49 & s_cla24_pg_logic10_or0;
  assign s_cla24_and51 = s_cla24_pg_logic10_and0 & s_cla24_pg_logic11_or0;
  assign s_cla24_or22 = s_cla24_and45 | s_cla24_and50;
  assign s_cla24_or23 = s_cla24_and48 | s_cla24_and51;
  assign s_cla24_or24 = s_cla24_or22 | s_cla24_or23;
  assign s_cla24_or25 = s_cla24_pg_logic11_and0 | s_cla24_or24;
  assign s_cla24_pg_logic12_or0 = a[12] | b[12];
  assign s_cla24_pg_logic12_and0 = a[12] & b[12];
  assign s_cla24_pg_logic12_xor0 = a[12] ^ b[12];
  assign s_cla24_xor12 = s_cla24_pg_logic12_xor0 ^ s_cla24_or25;
  assign s_cla24_and52 = s_cla24_or25 & s_cla24_pg_logic12_or0;
  assign s_cla24_or26 = s_cla24_pg_logic12_and0 | s_cla24_and52;
  assign s_cla24_pg_logic13_or0 = a[13] | b[13];
  assign s_cla24_pg_logic13_and0 = a[13] & b[13];
  assign s_cla24_pg_logic13_xor0 = a[13] ^ b[13];
  assign s_cla24_xor13 = s_cla24_pg_logic13_xor0 ^ s_cla24_or26;
  assign s_cla24_and53 = s_cla24_or25 & s_cla24_pg_logic13_or0;
  assign s_cla24_and54 = s_cla24_and53 & s_cla24_pg_logic12_or0;
  assign s_cla24_and55 = s_cla24_pg_logic12_and0 & s_cla24_pg_logic13_or0;
  assign s_cla24_or27 = s_cla24_and54 | s_cla24_and55;
  assign s_cla24_or28 = s_cla24_pg_logic13_and0 | s_cla24_or27;
  assign s_cla24_pg_logic14_or0 = a[14] | b[14];
  assign s_cla24_pg_logic14_and0 = a[14] & b[14];
  assign s_cla24_pg_logic14_xor0 = a[14] ^ b[14];
  assign s_cla24_xor14 = s_cla24_pg_logic14_xor0 ^ s_cla24_or28;
  assign s_cla24_and56 = s_cla24_or25 & s_cla24_pg_logic13_or0;
  assign s_cla24_and57 = s_cla24_pg_logic14_or0 & s_cla24_pg_logic12_or0;
  assign s_cla24_and58 = s_cla24_and56 & s_cla24_and57;
  assign s_cla24_and59 = s_cla24_pg_logic12_and0 & s_cla24_pg_logic14_or0;
  assign s_cla24_and60 = s_cla24_and59 & s_cla24_pg_logic13_or0;
  assign s_cla24_and61 = s_cla24_pg_logic13_and0 & s_cla24_pg_logic14_or0;
  assign s_cla24_or29 = s_cla24_and58 | s_cla24_and60;
  assign s_cla24_or30 = s_cla24_or29 | s_cla24_and61;
  assign s_cla24_or31 = s_cla24_pg_logic14_and0 | s_cla24_or30;
  assign s_cla24_pg_logic15_or0 = a[15] | b[15];
  assign s_cla24_pg_logic15_and0 = a[15] & b[15];
  assign s_cla24_pg_logic15_xor0 = a[15] ^ b[15];
  assign s_cla24_xor15 = s_cla24_pg_logic15_xor0 ^ s_cla24_or31;
  assign s_cla24_and62 = s_cla24_or25 & s_cla24_pg_logic14_or0;
  assign s_cla24_and63 = s_cla24_pg_logic15_or0 & s_cla24_pg_logic13_or0;
  assign s_cla24_and64 = s_cla24_and62 & s_cla24_and63;
  assign s_cla24_and65 = s_cla24_and64 & s_cla24_pg_logic12_or0;
  assign s_cla24_and66 = s_cla24_pg_logic12_and0 & s_cla24_pg_logic14_or0;
  assign s_cla24_and67 = s_cla24_pg_logic15_or0 & s_cla24_pg_logic13_or0;
  assign s_cla24_and68 = s_cla24_and66 & s_cla24_and67;
  assign s_cla24_and69 = s_cla24_pg_logic13_and0 & s_cla24_pg_logic15_or0;
  assign s_cla24_and70 = s_cla24_and69 & s_cla24_pg_logic14_or0;
  assign s_cla24_and71 = s_cla24_pg_logic14_and0 & s_cla24_pg_logic15_or0;
  assign s_cla24_or32 = s_cla24_and65 | s_cla24_and70;
  assign s_cla24_or33 = s_cla24_and68 | s_cla24_and71;
  assign s_cla24_or34 = s_cla24_or32 | s_cla24_or33;
  assign s_cla24_or35 = s_cla24_pg_logic15_and0 | s_cla24_or34;
  assign s_cla24_pg_logic16_or0 = a[16] | b[16];
  assign s_cla24_pg_logic16_and0 = a[16] & b[16];
  assign s_cla24_pg_logic16_xor0 = a[16] ^ b[16];
  assign s_cla24_xor16 = s_cla24_pg_logic16_xor0 ^ s_cla24_or35;
  assign s_cla24_and72 = s_cla24_or35 & s_cla24_pg_logic16_or0;
  assign s_cla24_or36 = s_cla24_pg_logic16_and0 | s_cla24_and72;
  assign s_cla24_pg_logic17_or0 = a[17] | b[17];
  assign s_cla24_pg_logic17_and0 = a[17] & b[17];
  assign s_cla24_pg_logic17_xor0 = a[17] ^ b[17];
  assign s_cla24_xor17 = s_cla24_pg_logic17_xor0 ^ s_cla24_or36;
  assign s_cla24_and73 = s_cla24_or35 & s_cla24_pg_logic17_or0;
  assign s_cla24_and74 = s_cla24_and73 & s_cla24_pg_logic16_or0;
  assign s_cla24_and75 = s_cla24_pg_logic16_and0 & s_cla24_pg_logic17_or0;
  assign s_cla24_or37 = s_cla24_and74 | s_cla24_and75;
  assign s_cla24_or38 = s_cla24_pg_logic17_and0 | s_cla24_or37;
  assign s_cla24_pg_logic18_or0 = a[18] | b[18];
  assign s_cla24_pg_logic18_and0 = a[18] & b[18];
  assign s_cla24_pg_logic18_xor0 = a[18] ^ b[18];
  assign s_cla24_xor18 = s_cla24_pg_logic18_xor0 ^ s_cla24_or38;
  assign s_cla24_and76 = s_cla24_or35 & s_cla24_pg_logic17_or0;
  assign s_cla24_and77 = s_cla24_pg_logic18_or0 & s_cla24_pg_logic16_or0;
  assign s_cla24_and78 = s_cla24_and76 & s_cla24_and77;
  assign s_cla24_and79 = s_cla24_pg_logic16_and0 & s_cla24_pg_logic18_or0;
  assign s_cla24_and80 = s_cla24_and79 & s_cla24_pg_logic17_or0;
  assign s_cla24_and81 = s_cla24_pg_logic17_and0 & s_cla24_pg_logic18_or0;
  assign s_cla24_or39 = s_cla24_and78 | s_cla24_and80;
  assign s_cla24_or40 = s_cla24_or39 | s_cla24_and81;
  assign s_cla24_or41 = s_cla24_pg_logic18_and0 | s_cla24_or40;
  assign s_cla24_pg_logic19_or0 = a[19] | b[19];
  assign s_cla24_pg_logic19_and0 = a[19] & b[19];
  assign s_cla24_pg_logic19_xor0 = a[19] ^ b[19];
  assign s_cla24_xor19 = s_cla24_pg_logic19_xor0 ^ s_cla24_or41;
  assign s_cla24_and82 = s_cla24_or35 & s_cla24_pg_logic18_or0;
  assign s_cla24_and83 = s_cla24_pg_logic19_or0 & s_cla24_pg_logic17_or0;
  assign s_cla24_and84 = s_cla24_and82 & s_cla24_and83;
  assign s_cla24_and85 = s_cla24_and84 & s_cla24_pg_logic16_or0;
  assign s_cla24_and86 = s_cla24_pg_logic16_and0 & s_cla24_pg_logic18_or0;
  assign s_cla24_and87 = s_cla24_pg_logic19_or0 & s_cla24_pg_logic17_or0;
  assign s_cla24_and88 = s_cla24_and86 & s_cla24_and87;
  assign s_cla24_and89 = s_cla24_pg_logic17_and0 & s_cla24_pg_logic19_or0;
  assign s_cla24_and90 = s_cla24_and89 & s_cla24_pg_logic18_or0;
  assign s_cla24_and91 = s_cla24_pg_logic18_and0 & s_cla24_pg_logic19_or0;
  assign s_cla24_or42 = s_cla24_and85 | s_cla24_and90;
  assign s_cla24_or43 = s_cla24_and88 | s_cla24_and91;
  assign s_cla24_or44 = s_cla24_or42 | s_cla24_or43;
  assign s_cla24_or45 = s_cla24_pg_logic19_and0 | s_cla24_or44;
  assign s_cla24_pg_logic20_or0 = a[20] | b[20];
  assign s_cla24_pg_logic20_and0 = a[20] & b[20];
  assign s_cla24_pg_logic20_xor0 = a[20] ^ b[20];
  assign s_cla24_xor20 = s_cla24_pg_logic20_xor0 ^ s_cla24_or45;
  assign s_cla24_and92 = s_cla24_or45 & s_cla24_pg_logic20_or0;
  assign s_cla24_or46 = s_cla24_pg_logic20_and0 | s_cla24_and92;
  assign s_cla24_pg_logic21_or0 = a[21] | b[21];
  assign s_cla24_pg_logic21_and0 = a[21] & b[21];
  assign s_cla24_pg_logic21_xor0 = a[21] ^ b[21];
  assign s_cla24_xor21 = s_cla24_pg_logic21_xor0 ^ s_cla24_or46;
  assign s_cla24_and93 = s_cla24_or45 & s_cla24_pg_logic21_or0;
  assign s_cla24_and94 = s_cla24_and93 & s_cla24_pg_logic20_or0;
  assign s_cla24_and95 = s_cla24_pg_logic20_and0 & s_cla24_pg_logic21_or0;
  assign s_cla24_or47 = s_cla24_and94 | s_cla24_and95;
  assign s_cla24_or48 = s_cla24_pg_logic21_and0 | s_cla24_or47;
  assign s_cla24_pg_logic22_or0 = a[22] | b[22];
  assign s_cla24_pg_logic22_and0 = a[22] & b[22];
  assign s_cla24_pg_logic22_xor0 = a[22] ^ b[22];
  assign s_cla24_xor22 = s_cla24_pg_logic22_xor0 ^ s_cla24_or48;
  assign s_cla24_and96 = s_cla24_or45 & s_cla24_pg_logic21_or0;
  assign s_cla24_and97 = s_cla24_pg_logic22_or0 & s_cla24_pg_logic20_or0;
  assign s_cla24_and98 = s_cla24_and96 & s_cla24_and97;
  assign s_cla24_and99 = s_cla24_pg_logic20_and0 & s_cla24_pg_logic22_or0;
  assign s_cla24_and100 = s_cla24_and99 & s_cla24_pg_logic21_or0;
  assign s_cla24_and101 = s_cla24_pg_logic21_and0 & s_cla24_pg_logic22_or0;
  assign s_cla24_or49 = s_cla24_and98 | s_cla24_and100;
  assign s_cla24_or50 = s_cla24_or49 | s_cla24_and101;
  assign s_cla24_or51 = s_cla24_pg_logic22_and0 | s_cla24_or50;
  assign s_cla24_pg_logic23_or0 = a[23] | b[23];
  assign s_cla24_pg_logic23_and0 = a[23] & b[23];
  assign s_cla24_pg_logic23_xor0 = a[23] ^ b[23];
  assign s_cla24_xor23 = s_cla24_pg_logic23_xor0 ^ s_cla24_or51;
  assign s_cla24_and102 = s_cla24_or45 & s_cla24_pg_logic22_or0;
  assign s_cla24_and103 = s_cla24_pg_logic23_or0 & s_cla24_pg_logic21_or0;
  assign s_cla24_and104 = s_cla24_and102 & s_cla24_and103;
  assign s_cla24_and105 = s_cla24_and104 & s_cla24_pg_logic20_or0;
  assign s_cla24_and106 = s_cla24_pg_logic20_and0 & s_cla24_pg_logic22_or0;
  assign s_cla24_and107 = s_cla24_pg_logic23_or0 & s_cla24_pg_logic21_or0;
  assign s_cla24_and108 = s_cla24_and106 & s_cla24_and107;
  assign s_cla24_and109 = s_cla24_pg_logic21_and0 & s_cla24_pg_logic23_or0;
  assign s_cla24_and110 = s_cla24_and109 & s_cla24_pg_logic22_or0;
  assign s_cla24_and111 = s_cla24_pg_logic22_and0 & s_cla24_pg_logic23_or0;
  assign s_cla24_or52 = s_cla24_and105 | s_cla24_and110;
  assign s_cla24_or53 = s_cla24_and108 | s_cla24_and111;
  assign s_cla24_or54 = s_cla24_or52 | s_cla24_or53;
  assign s_cla24_or55 = s_cla24_pg_logic23_and0 | s_cla24_or54;
  assign s_cla24_xor24 = a[23] ^ b[23];
  assign s_cla24_xor25 = s_cla24_xor24 ^ s_cla24_or55;

  assign s_cla24_out[0] = s_cla24_pg_logic0_xor0;
  assign s_cla24_out[1] = s_cla24_xor1;
  assign s_cla24_out[2] = s_cla24_xor2;
  assign s_cla24_out[3] = s_cla24_xor3;
  assign s_cla24_out[4] = s_cla24_xor4;
  assign s_cla24_out[5] = s_cla24_xor5;
  assign s_cla24_out[6] = s_cla24_xor6;
  assign s_cla24_out[7] = s_cla24_xor7;
  assign s_cla24_out[8] = s_cla24_xor8;
  assign s_cla24_out[9] = s_cla24_xor9;
  assign s_cla24_out[10] = s_cla24_xor10;
  assign s_cla24_out[11] = s_cla24_xor11;
  assign s_cla24_out[12] = s_cla24_xor12;
  assign s_cla24_out[13] = s_cla24_xor13;
  assign s_cla24_out[14] = s_cla24_xor14;
  assign s_cla24_out[15] = s_cla24_xor15;
  assign s_cla24_out[16] = s_cla24_xor16;
  assign s_cla24_out[17] = s_cla24_xor17;
  assign s_cla24_out[18] = s_cla24_xor18;
  assign s_cla24_out[19] = s_cla24_xor19;
  assign s_cla24_out[20] = s_cla24_xor20;
  assign s_cla24_out[21] = s_cla24_xor21;
  assign s_cla24_out[22] = s_cla24_xor22;
  assign s_cla24_out[23] = s_cla24_xor23;
  assign s_cla24_out[24] = s_cla24_xor25;
endmodule