module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module nor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a | _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module constant_wire_value_0(input a, input b, output constant_wire_0);
  wire constant_wire_value_0_a;
  wire constant_wire_value_0_b;

  assign constant_wire_value_0_a = a;
  assign constant_wire_value_0_b = b;

  xor_gate xor_gate_constant_wire_value_0_y0(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y0);
  xnor_gate xnor_gate_constant_wire_value_0_y1(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y1);
  nor_gate nor_gate_constant_wire_0(constant_wire_value_0_y0, constant_wire_value_0_y1, constant_wire_0);
endmodule

module pg_logic(input a, input b, output pg_logic_y0, output pg_logic_y1, output pg_logic_y2);
  wire pg_logic_a;
  wire pg_logic_b;

  assign pg_logic_a = a;
  assign pg_logic_b = b;

  or_gate or_gate_pg_logic_y0(pg_logic_a, pg_logic_b, pg_logic_y0);
  and_gate and_gate_pg_logic_y1(pg_logic_a, pg_logic_b, pg_logic_y1);
  xor_gate xor_gate_pg_logic_y2(pg_logic_a, pg_logic_b, pg_logic_y2);
endmodule

module h_u_cla12(input [11:0] a, input [11:0] b, output [12:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire constant_wire_0;
  wire h_u_cla12_pg_logic0_y0;
  wire h_u_cla12_pg_logic0_y1;
  wire h_u_cla12_pg_logic0_y2;
  wire h_u_cla12_xor0_y0;
  wire h_u_cla12_and0_y0;
  wire h_u_cla12_or0_y0;
  wire h_u_cla12_pg_logic1_y0;
  wire h_u_cla12_pg_logic1_y1;
  wire h_u_cla12_pg_logic1_y2;
  wire h_u_cla12_xor1_y0;
  wire h_u_cla12_and1_y0;
  wire h_u_cla12_and2_y0;
  wire h_u_cla12_and3_y0;
  wire h_u_cla12_and4_y0;
  wire h_u_cla12_or1_y0;
  wire h_u_cla12_or2_y0;
  wire h_u_cla12_pg_logic2_y0;
  wire h_u_cla12_pg_logic2_y1;
  wire h_u_cla12_pg_logic2_y2;
  wire h_u_cla12_xor2_y0;
  wire h_u_cla12_and5_y0;
  wire h_u_cla12_and6_y0;
  wire h_u_cla12_and7_y0;
  wire h_u_cla12_and8_y0;
  wire h_u_cla12_and9_y0;
  wire h_u_cla12_and10_y0;
  wire h_u_cla12_and11_y0;
  wire h_u_cla12_and12_y0;
  wire h_u_cla12_and13_y0;
  wire h_u_cla12_or3_y0;
  wire h_u_cla12_or4_y0;
  wire h_u_cla12_or5_y0;
  wire h_u_cla12_pg_logic3_y0;
  wire h_u_cla12_pg_logic3_y1;
  wire h_u_cla12_pg_logic3_y2;
  wire h_u_cla12_xor3_y0;
  wire h_u_cla12_and14_y0;
  wire h_u_cla12_and15_y0;
  wire h_u_cla12_and16_y0;
  wire h_u_cla12_and17_y0;
  wire h_u_cla12_and18_y0;
  wire h_u_cla12_and19_y0;
  wire h_u_cla12_and20_y0;
  wire h_u_cla12_and21_y0;
  wire h_u_cla12_and22_y0;
  wire h_u_cla12_and23_y0;
  wire h_u_cla12_and24_y0;
  wire h_u_cla12_and25_y0;
  wire h_u_cla12_and26_y0;
  wire h_u_cla12_and27_y0;
  wire h_u_cla12_and28_y0;
  wire h_u_cla12_and29_y0;
  wire h_u_cla12_or6_y0;
  wire h_u_cla12_or7_y0;
  wire h_u_cla12_or8_y0;
  wire h_u_cla12_or9_y0;
  wire h_u_cla12_pg_logic4_y0;
  wire h_u_cla12_pg_logic4_y1;
  wire h_u_cla12_pg_logic4_y2;
  wire h_u_cla12_xor4_y0;
  wire h_u_cla12_and30_y0;
  wire h_u_cla12_and31_y0;
  wire h_u_cla12_and32_y0;
  wire h_u_cla12_and33_y0;
  wire h_u_cla12_and34_y0;
  wire h_u_cla12_and35_y0;
  wire h_u_cla12_and36_y0;
  wire h_u_cla12_and37_y0;
  wire h_u_cla12_and38_y0;
  wire h_u_cla12_and39_y0;
  wire h_u_cla12_and40_y0;
  wire h_u_cla12_and41_y0;
  wire h_u_cla12_and42_y0;
  wire h_u_cla12_and43_y0;
  wire h_u_cla12_and44_y0;
  wire h_u_cla12_and45_y0;
  wire h_u_cla12_and46_y0;
  wire h_u_cla12_and47_y0;
  wire h_u_cla12_and48_y0;
  wire h_u_cla12_and49_y0;
  wire h_u_cla12_and50_y0;
  wire h_u_cla12_and51_y0;
  wire h_u_cla12_and52_y0;
  wire h_u_cla12_and53_y0;
  wire h_u_cla12_and54_y0;
  wire h_u_cla12_or10_y0;
  wire h_u_cla12_or11_y0;
  wire h_u_cla12_or12_y0;
  wire h_u_cla12_or13_y0;
  wire h_u_cla12_or14_y0;
  wire h_u_cla12_pg_logic5_y0;
  wire h_u_cla12_pg_logic5_y1;
  wire h_u_cla12_pg_logic5_y2;
  wire h_u_cla12_xor5_y0;
  wire h_u_cla12_and55_y0;
  wire h_u_cla12_and56_y0;
  wire h_u_cla12_and57_y0;
  wire h_u_cla12_and58_y0;
  wire h_u_cla12_and59_y0;
  wire h_u_cla12_and60_y0;
  wire h_u_cla12_and61_y0;
  wire h_u_cla12_and62_y0;
  wire h_u_cla12_and63_y0;
  wire h_u_cla12_and64_y0;
  wire h_u_cla12_and65_y0;
  wire h_u_cla12_and66_y0;
  wire h_u_cla12_and67_y0;
  wire h_u_cla12_and68_y0;
  wire h_u_cla12_and69_y0;
  wire h_u_cla12_and70_y0;
  wire h_u_cla12_and71_y0;
  wire h_u_cla12_and72_y0;
  wire h_u_cla12_and73_y0;
  wire h_u_cla12_and74_y0;
  wire h_u_cla12_and75_y0;
  wire h_u_cla12_and76_y0;
  wire h_u_cla12_and77_y0;
  wire h_u_cla12_and78_y0;
  wire h_u_cla12_and79_y0;
  wire h_u_cla12_and80_y0;
  wire h_u_cla12_and81_y0;
  wire h_u_cla12_and82_y0;
  wire h_u_cla12_and83_y0;
  wire h_u_cla12_and84_y0;
  wire h_u_cla12_and85_y0;
  wire h_u_cla12_and86_y0;
  wire h_u_cla12_and87_y0;
  wire h_u_cla12_and88_y0;
  wire h_u_cla12_and89_y0;
  wire h_u_cla12_and90_y0;
  wire h_u_cla12_or15_y0;
  wire h_u_cla12_or16_y0;
  wire h_u_cla12_or17_y0;
  wire h_u_cla12_or18_y0;
  wire h_u_cla12_or19_y0;
  wire h_u_cla12_or20_y0;
  wire h_u_cla12_pg_logic6_y0;
  wire h_u_cla12_pg_logic6_y1;
  wire h_u_cla12_pg_logic6_y2;
  wire h_u_cla12_xor6_y0;
  wire h_u_cla12_and91_y0;
  wire h_u_cla12_and92_y0;
  wire h_u_cla12_and93_y0;
  wire h_u_cla12_and94_y0;
  wire h_u_cla12_and95_y0;
  wire h_u_cla12_and96_y0;
  wire h_u_cla12_and97_y0;
  wire h_u_cla12_and98_y0;
  wire h_u_cla12_and99_y0;
  wire h_u_cla12_and100_y0;
  wire h_u_cla12_and101_y0;
  wire h_u_cla12_and102_y0;
  wire h_u_cla12_and103_y0;
  wire h_u_cla12_and104_y0;
  wire h_u_cla12_and105_y0;
  wire h_u_cla12_and106_y0;
  wire h_u_cla12_and107_y0;
  wire h_u_cla12_and108_y0;
  wire h_u_cla12_and109_y0;
  wire h_u_cla12_and110_y0;
  wire h_u_cla12_and111_y0;
  wire h_u_cla12_and112_y0;
  wire h_u_cla12_and113_y0;
  wire h_u_cla12_and114_y0;
  wire h_u_cla12_and115_y0;
  wire h_u_cla12_and116_y0;
  wire h_u_cla12_and117_y0;
  wire h_u_cla12_and118_y0;
  wire h_u_cla12_and119_y0;
  wire h_u_cla12_and120_y0;
  wire h_u_cla12_and121_y0;
  wire h_u_cla12_and122_y0;
  wire h_u_cla12_and123_y0;
  wire h_u_cla12_and124_y0;
  wire h_u_cla12_and125_y0;
  wire h_u_cla12_and126_y0;
  wire h_u_cla12_and127_y0;
  wire h_u_cla12_and128_y0;
  wire h_u_cla12_and129_y0;
  wire h_u_cla12_and130_y0;
  wire h_u_cla12_and131_y0;
  wire h_u_cla12_and132_y0;
  wire h_u_cla12_and133_y0;
  wire h_u_cla12_and134_y0;
  wire h_u_cla12_and135_y0;
  wire h_u_cla12_and136_y0;
  wire h_u_cla12_and137_y0;
  wire h_u_cla12_and138_y0;
  wire h_u_cla12_and139_y0;
  wire h_u_cla12_or21_y0;
  wire h_u_cla12_or22_y0;
  wire h_u_cla12_or23_y0;
  wire h_u_cla12_or24_y0;
  wire h_u_cla12_or25_y0;
  wire h_u_cla12_or26_y0;
  wire h_u_cla12_or27_y0;
  wire h_u_cla12_pg_logic7_y0;
  wire h_u_cla12_pg_logic7_y1;
  wire h_u_cla12_pg_logic7_y2;
  wire h_u_cla12_xor7_y0;
  wire h_u_cla12_and140_y0;
  wire h_u_cla12_and141_y0;
  wire h_u_cla12_and142_y0;
  wire h_u_cla12_and143_y0;
  wire h_u_cla12_and144_y0;
  wire h_u_cla12_and145_y0;
  wire h_u_cla12_and146_y0;
  wire h_u_cla12_and147_y0;
  wire h_u_cla12_and148_y0;
  wire h_u_cla12_and149_y0;
  wire h_u_cla12_and150_y0;
  wire h_u_cla12_and151_y0;
  wire h_u_cla12_and152_y0;
  wire h_u_cla12_and153_y0;
  wire h_u_cla12_and154_y0;
  wire h_u_cla12_and155_y0;
  wire h_u_cla12_and156_y0;
  wire h_u_cla12_and157_y0;
  wire h_u_cla12_and158_y0;
  wire h_u_cla12_and159_y0;
  wire h_u_cla12_and160_y0;
  wire h_u_cla12_and161_y0;
  wire h_u_cla12_and162_y0;
  wire h_u_cla12_and163_y0;
  wire h_u_cla12_and164_y0;
  wire h_u_cla12_and165_y0;
  wire h_u_cla12_and166_y0;
  wire h_u_cla12_and167_y0;
  wire h_u_cla12_and168_y0;
  wire h_u_cla12_and169_y0;
  wire h_u_cla12_and170_y0;
  wire h_u_cla12_and171_y0;
  wire h_u_cla12_and172_y0;
  wire h_u_cla12_and173_y0;
  wire h_u_cla12_and174_y0;
  wire h_u_cla12_and175_y0;
  wire h_u_cla12_and176_y0;
  wire h_u_cla12_and177_y0;
  wire h_u_cla12_and178_y0;
  wire h_u_cla12_and179_y0;
  wire h_u_cla12_and180_y0;
  wire h_u_cla12_and181_y0;
  wire h_u_cla12_and182_y0;
  wire h_u_cla12_and183_y0;
  wire h_u_cla12_and184_y0;
  wire h_u_cla12_and185_y0;
  wire h_u_cla12_and186_y0;
  wire h_u_cla12_and187_y0;
  wire h_u_cla12_and188_y0;
  wire h_u_cla12_and189_y0;
  wire h_u_cla12_and190_y0;
  wire h_u_cla12_and191_y0;
  wire h_u_cla12_and192_y0;
  wire h_u_cla12_and193_y0;
  wire h_u_cla12_and194_y0;
  wire h_u_cla12_and195_y0;
  wire h_u_cla12_and196_y0;
  wire h_u_cla12_and197_y0;
  wire h_u_cla12_and198_y0;
  wire h_u_cla12_and199_y0;
  wire h_u_cla12_and200_y0;
  wire h_u_cla12_and201_y0;
  wire h_u_cla12_and202_y0;
  wire h_u_cla12_and203_y0;
  wire h_u_cla12_or28_y0;
  wire h_u_cla12_or29_y0;
  wire h_u_cla12_or30_y0;
  wire h_u_cla12_or31_y0;
  wire h_u_cla12_or32_y0;
  wire h_u_cla12_or33_y0;
  wire h_u_cla12_or34_y0;
  wire h_u_cla12_or35_y0;
  wire h_u_cla12_pg_logic8_y0;
  wire h_u_cla12_pg_logic8_y1;
  wire h_u_cla12_pg_logic8_y2;
  wire h_u_cla12_xor8_y0;
  wire h_u_cla12_and204_y0;
  wire h_u_cla12_and205_y0;
  wire h_u_cla12_and206_y0;
  wire h_u_cla12_and207_y0;
  wire h_u_cla12_and208_y0;
  wire h_u_cla12_and209_y0;
  wire h_u_cla12_and210_y0;
  wire h_u_cla12_and211_y0;
  wire h_u_cla12_and212_y0;
  wire h_u_cla12_and213_y0;
  wire h_u_cla12_and214_y0;
  wire h_u_cla12_and215_y0;
  wire h_u_cla12_and216_y0;
  wire h_u_cla12_and217_y0;
  wire h_u_cla12_and218_y0;
  wire h_u_cla12_and219_y0;
  wire h_u_cla12_and220_y0;
  wire h_u_cla12_and221_y0;
  wire h_u_cla12_and222_y0;
  wire h_u_cla12_and223_y0;
  wire h_u_cla12_and224_y0;
  wire h_u_cla12_and225_y0;
  wire h_u_cla12_and226_y0;
  wire h_u_cla12_and227_y0;
  wire h_u_cla12_and228_y0;
  wire h_u_cla12_and229_y0;
  wire h_u_cla12_and230_y0;
  wire h_u_cla12_and231_y0;
  wire h_u_cla12_and232_y0;
  wire h_u_cla12_and233_y0;
  wire h_u_cla12_and234_y0;
  wire h_u_cla12_and235_y0;
  wire h_u_cla12_and236_y0;
  wire h_u_cla12_and237_y0;
  wire h_u_cla12_and238_y0;
  wire h_u_cla12_and239_y0;
  wire h_u_cla12_and240_y0;
  wire h_u_cla12_and241_y0;
  wire h_u_cla12_and242_y0;
  wire h_u_cla12_and243_y0;
  wire h_u_cla12_and244_y0;
  wire h_u_cla12_and245_y0;
  wire h_u_cla12_and246_y0;
  wire h_u_cla12_and247_y0;
  wire h_u_cla12_and248_y0;
  wire h_u_cla12_and249_y0;
  wire h_u_cla12_and250_y0;
  wire h_u_cla12_and251_y0;
  wire h_u_cla12_and252_y0;
  wire h_u_cla12_and253_y0;
  wire h_u_cla12_and254_y0;
  wire h_u_cla12_and255_y0;
  wire h_u_cla12_and256_y0;
  wire h_u_cla12_and257_y0;
  wire h_u_cla12_and258_y0;
  wire h_u_cla12_and259_y0;
  wire h_u_cla12_and260_y0;
  wire h_u_cla12_and261_y0;
  wire h_u_cla12_and262_y0;
  wire h_u_cla12_and263_y0;
  wire h_u_cla12_and264_y0;
  wire h_u_cla12_and265_y0;
  wire h_u_cla12_and266_y0;
  wire h_u_cla12_and267_y0;
  wire h_u_cla12_and268_y0;
  wire h_u_cla12_and269_y0;
  wire h_u_cla12_and270_y0;
  wire h_u_cla12_and271_y0;
  wire h_u_cla12_and272_y0;
  wire h_u_cla12_and273_y0;
  wire h_u_cla12_and274_y0;
  wire h_u_cla12_and275_y0;
  wire h_u_cla12_and276_y0;
  wire h_u_cla12_and277_y0;
  wire h_u_cla12_and278_y0;
  wire h_u_cla12_and279_y0;
  wire h_u_cla12_and280_y0;
  wire h_u_cla12_and281_y0;
  wire h_u_cla12_and282_y0;
  wire h_u_cla12_and283_y0;
  wire h_u_cla12_and284_y0;
  wire h_u_cla12_or36_y0;
  wire h_u_cla12_or37_y0;
  wire h_u_cla12_or38_y0;
  wire h_u_cla12_or39_y0;
  wire h_u_cla12_or40_y0;
  wire h_u_cla12_or41_y0;
  wire h_u_cla12_or42_y0;
  wire h_u_cla12_or43_y0;
  wire h_u_cla12_or44_y0;
  wire h_u_cla12_pg_logic9_y0;
  wire h_u_cla12_pg_logic9_y1;
  wire h_u_cla12_pg_logic9_y2;
  wire h_u_cla12_xor9_y0;
  wire h_u_cla12_and285_y0;
  wire h_u_cla12_and286_y0;
  wire h_u_cla12_and287_y0;
  wire h_u_cla12_and288_y0;
  wire h_u_cla12_and289_y0;
  wire h_u_cla12_and290_y0;
  wire h_u_cla12_and291_y0;
  wire h_u_cla12_and292_y0;
  wire h_u_cla12_and293_y0;
  wire h_u_cla12_and294_y0;
  wire h_u_cla12_and295_y0;
  wire h_u_cla12_and296_y0;
  wire h_u_cla12_and297_y0;
  wire h_u_cla12_and298_y0;
  wire h_u_cla12_and299_y0;
  wire h_u_cla12_and300_y0;
  wire h_u_cla12_and301_y0;
  wire h_u_cla12_and302_y0;
  wire h_u_cla12_and303_y0;
  wire h_u_cla12_and304_y0;
  wire h_u_cla12_and305_y0;
  wire h_u_cla12_and306_y0;
  wire h_u_cla12_and307_y0;
  wire h_u_cla12_and308_y0;
  wire h_u_cla12_and309_y0;
  wire h_u_cla12_and310_y0;
  wire h_u_cla12_and311_y0;
  wire h_u_cla12_and312_y0;
  wire h_u_cla12_and313_y0;
  wire h_u_cla12_and314_y0;
  wire h_u_cla12_and315_y0;
  wire h_u_cla12_and316_y0;
  wire h_u_cla12_and317_y0;
  wire h_u_cla12_and318_y0;
  wire h_u_cla12_and319_y0;
  wire h_u_cla12_and320_y0;
  wire h_u_cla12_and321_y0;
  wire h_u_cla12_and322_y0;
  wire h_u_cla12_and323_y0;
  wire h_u_cla12_and324_y0;
  wire h_u_cla12_and325_y0;
  wire h_u_cla12_and326_y0;
  wire h_u_cla12_and327_y0;
  wire h_u_cla12_and328_y0;
  wire h_u_cla12_and329_y0;
  wire h_u_cla12_and330_y0;
  wire h_u_cla12_and331_y0;
  wire h_u_cla12_and332_y0;
  wire h_u_cla12_and333_y0;
  wire h_u_cla12_and334_y0;
  wire h_u_cla12_and335_y0;
  wire h_u_cla12_and336_y0;
  wire h_u_cla12_and337_y0;
  wire h_u_cla12_and338_y0;
  wire h_u_cla12_and339_y0;
  wire h_u_cla12_and340_y0;
  wire h_u_cla12_and341_y0;
  wire h_u_cla12_and342_y0;
  wire h_u_cla12_and343_y0;
  wire h_u_cla12_and344_y0;
  wire h_u_cla12_and345_y0;
  wire h_u_cla12_and346_y0;
  wire h_u_cla12_and347_y0;
  wire h_u_cla12_and348_y0;
  wire h_u_cla12_and349_y0;
  wire h_u_cla12_and350_y0;
  wire h_u_cla12_and351_y0;
  wire h_u_cla12_and352_y0;
  wire h_u_cla12_and353_y0;
  wire h_u_cla12_and354_y0;
  wire h_u_cla12_and355_y0;
  wire h_u_cla12_and356_y0;
  wire h_u_cla12_and357_y0;
  wire h_u_cla12_and358_y0;
  wire h_u_cla12_and359_y0;
  wire h_u_cla12_and360_y0;
  wire h_u_cla12_and361_y0;
  wire h_u_cla12_and362_y0;
  wire h_u_cla12_and363_y0;
  wire h_u_cla12_and364_y0;
  wire h_u_cla12_and365_y0;
  wire h_u_cla12_and366_y0;
  wire h_u_cla12_and367_y0;
  wire h_u_cla12_and368_y0;
  wire h_u_cla12_and369_y0;
  wire h_u_cla12_and370_y0;
  wire h_u_cla12_and371_y0;
  wire h_u_cla12_and372_y0;
  wire h_u_cla12_and373_y0;
  wire h_u_cla12_and374_y0;
  wire h_u_cla12_and375_y0;
  wire h_u_cla12_and376_y0;
  wire h_u_cla12_and377_y0;
  wire h_u_cla12_and378_y0;
  wire h_u_cla12_and379_y0;
  wire h_u_cla12_and380_y0;
  wire h_u_cla12_and381_y0;
  wire h_u_cla12_and382_y0;
  wire h_u_cla12_and383_y0;
  wire h_u_cla12_and384_y0;
  wire h_u_cla12_or45_y0;
  wire h_u_cla12_or46_y0;
  wire h_u_cla12_or47_y0;
  wire h_u_cla12_or48_y0;
  wire h_u_cla12_or49_y0;
  wire h_u_cla12_or50_y0;
  wire h_u_cla12_or51_y0;
  wire h_u_cla12_or52_y0;
  wire h_u_cla12_or53_y0;
  wire h_u_cla12_or54_y0;
  wire h_u_cla12_pg_logic10_y0;
  wire h_u_cla12_pg_logic10_y1;
  wire h_u_cla12_pg_logic10_y2;
  wire h_u_cla12_xor10_y0;
  wire h_u_cla12_and385_y0;
  wire h_u_cla12_and386_y0;
  wire h_u_cla12_and387_y0;
  wire h_u_cla12_and388_y0;
  wire h_u_cla12_and389_y0;
  wire h_u_cla12_and390_y0;
  wire h_u_cla12_and391_y0;
  wire h_u_cla12_and392_y0;
  wire h_u_cla12_and393_y0;
  wire h_u_cla12_and394_y0;
  wire h_u_cla12_and395_y0;
  wire h_u_cla12_and396_y0;
  wire h_u_cla12_and397_y0;
  wire h_u_cla12_and398_y0;
  wire h_u_cla12_and399_y0;
  wire h_u_cla12_and400_y0;
  wire h_u_cla12_and401_y0;
  wire h_u_cla12_and402_y0;
  wire h_u_cla12_and403_y0;
  wire h_u_cla12_and404_y0;
  wire h_u_cla12_and405_y0;
  wire h_u_cla12_and406_y0;
  wire h_u_cla12_and407_y0;
  wire h_u_cla12_and408_y0;
  wire h_u_cla12_and409_y0;
  wire h_u_cla12_and410_y0;
  wire h_u_cla12_and411_y0;
  wire h_u_cla12_and412_y0;
  wire h_u_cla12_and413_y0;
  wire h_u_cla12_and414_y0;
  wire h_u_cla12_and415_y0;
  wire h_u_cla12_and416_y0;
  wire h_u_cla12_and417_y0;
  wire h_u_cla12_and418_y0;
  wire h_u_cla12_and419_y0;
  wire h_u_cla12_and420_y0;
  wire h_u_cla12_and421_y0;
  wire h_u_cla12_and422_y0;
  wire h_u_cla12_and423_y0;
  wire h_u_cla12_and424_y0;
  wire h_u_cla12_and425_y0;
  wire h_u_cla12_and426_y0;
  wire h_u_cla12_and427_y0;
  wire h_u_cla12_and428_y0;
  wire h_u_cla12_and429_y0;
  wire h_u_cla12_and430_y0;
  wire h_u_cla12_and431_y0;
  wire h_u_cla12_and432_y0;
  wire h_u_cla12_and433_y0;
  wire h_u_cla12_and434_y0;
  wire h_u_cla12_and435_y0;
  wire h_u_cla12_and436_y0;
  wire h_u_cla12_and437_y0;
  wire h_u_cla12_and438_y0;
  wire h_u_cla12_and439_y0;
  wire h_u_cla12_and440_y0;
  wire h_u_cla12_and441_y0;
  wire h_u_cla12_and442_y0;
  wire h_u_cla12_and443_y0;
  wire h_u_cla12_and444_y0;
  wire h_u_cla12_and445_y0;
  wire h_u_cla12_and446_y0;
  wire h_u_cla12_and447_y0;
  wire h_u_cla12_and448_y0;
  wire h_u_cla12_and449_y0;
  wire h_u_cla12_and450_y0;
  wire h_u_cla12_and451_y0;
  wire h_u_cla12_and452_y0;
  wire h_u_cla12_and453_y0;
  wire h_u_cla12_and454_y0;
  wire h_u_cla12_and455_y0;
  wire h_u_cla12_and456_y0;
  wire h_u_cla12_and457_y0;
  wire h_u_cla12_and458_y0;
  wire h_u_cla12_and459_y0;
  wire h_u_cla12_and460_y0;
  wire h_u_cla12_and461_y0;
  wire h_u_cla12_and462_y0;
  wire h_u_cla12_and463_y0;
  wire h_u_cla12_and464_y0;
  wire h_u_cla12_and465_y0;
  wire h_u_cla12_and466_y0;
  wire h_u_cla12_and467_y0;
  wire h_u_cla12_and468_y0;
  wire h_u_cla12_and469_y0;
  wire h_u_cla12_and470_y0;
  wire h_u_cla12_and471_y0;
  wire h_u_cla12_and472_y0;
  wire h_u_cla12_and473_y0;
  wire h_u_cla12_and474_y0;
  wire h_u_cla12_and475_y0;
  wire h_u_cla12_and476_y0;
  wire h_u_cla12_and477_y0;
  wire h_u_cla12_and478_y0;
  wire h_u_cla12_and479_y0;
  wire h_u_cla12_and480_y0;
  wire h_u_cla12_and481_y0;
  wire h_u_cla12_and482_y0;
  wire h_u_cla12_and483_y0;
  wire h_u_cla12_and484_y0;
  wire h_u_cla12_and485_y0;
  wire h_u_cla12_and486_y0;
  wire h_u_cla12_and487_y0;
  wire h_u_cla12_and488_y0;
  wire h_u_cla12_and489_y0;
  wire h_u_cla12_and490_y0;
  wire h_u_cla12_and491_y0;
  wire h_u_cla12_and492_y0;
  wire h_u_cla12_and493_y0;
  wire h_u_cla12_and494_y0;
  wire h_u_cla12_and495_y0;
  wire h_u_cla12_and496_y0;
  wire h_u_cla12_and497_y0;
  wire h_u_cla12_and498_y0;
  wire h_u_cla12_and499_y0;
  wire h_u_cla12_and500_y0;
  wire h_u_cla12_and501_y0;
  wire h_u_cla12_and502_y0;
  wire h_u_cla12_and503_y0;
  wire h_u_cla12_and504_y0;
  wire h_u_cla12_and505_y0;
  wire h_u_cla12_or55_y0;
  wire h_u_cla12_or56_y0;
  wire h_u_cla12_or57_y0;
  wire h_u_cla12_or58_y0;
  wire h_u_cla12_or59_y0;
  wire h_u_cla12_or60_y0;
  wire h_u_cla12_or61_y0;
  wire h_u_cla12_or62_y0;
  wire h_u_cla12_or63_y0;
  wire h_u_cla12_or64_y0;
  wire h_u_cla12_or65_y0;
  wire h_u_cla12_pg_logic11_y0;
  wire h_u_cla12_pg_logic11_y1;
  wire h_u_cla12_pg_logic11_y2;
  wire h_u_cla12_xor11_y0;
  wire h_u_cla12_and506_y0;
  wire h_u_cla12_and507_y0;
  wire h_u_cla12_and508_y0;
  wire h_u_cla12_and509_y0;
  wire h_u_cla12_and510_y0;
  wire h_u_cla12_and511_y0;
  wire h_u_cla12_and512_y0;
  wire h_u_cla12_and513_y0;
  wire h_u_cla12_and514_y0;
  wire h_u_cla12_and515_y0;
  wire h_u_cla12_and516_y0;
  wire h_u_cla12_and517_y0;
  wire h_u_cla12_and518_y0;
  wire h_u_cla12_and519_y0;
  wire h_u_cla12_and520_y0;
  wire h_u_cla12_and521_y0;
  wire h_u_cla12_and522_y0;
  wire h_u_cla12_and523_y0;
  wire h_u_cla12_and524_y0;
  wire h_u_cla12_and525_y0;
  wire h_u_cla12_and526_y0;
  wire h_u_cla12_and527_y0;
  wire h_u_cla12_and528_y0;
  wire h_u_cla12_and529_y0;
  wire h_u_cla12_and530_y0;
  wire h_u_cla12_and531_y0;
  wire h_u_cla12_and532_y0;
  wire h_u_cla12_and533_y0;
  wire h_u_cla12_and534_y0;
  wire h_u_cla12_and535_y0;
  wire h_u_cla12_and536_y0;
  wire h_u_cla12_and537_y0;
  wire h_u_cla12_and538_y0;
  wire h_u_cla12_and539_y0;
  wire h_u_cla12_and540_y0;
  wire h_u_cla12_and541_y0;
  wire h_u_cla12_and542_y0;
  wire h_u_cla12_and543_y0;
  wire h_u_cla12_and544_y0;
  wire h_u_cla12_and545_y0;
  wire h_u_cla12_and546_y0;
  wire h_u_cla12_and547_y0;
  wire h_u_cla12_and548_y0;
  wire h_u_cla12_and549_y0;
  wire h_u_cla12_and550_y0;
  wire h_u_cla12_and551_y0;
  wire h_u_cla12_and552_y0;
  wire h_u_cla12_and553_y0;
  wire h_u_cla12_and554_y0;
  wire h_u_cla12_and555_y0;
  wire h_u_cla12_and556_y0;
  wire h_u_cla12_and557_y0;
  wire h_u_cla12_and558_y0;
  wire h_u_cla12_and559_y0;
  wire h_u_cla12_and560_y0;
  wire h_u_cla12_and561_y0;
  wire h_u_cla12_and562_y0;
  wire h_u_cla12_and563_y0;
  wire h_u_cla12_and564_y0;
  wire h_u_cla12_and565_y0;
  wire h_u_cla12_and566_y0;
  wire h_u_cla12_and567_y0;
  wire h_u_cla12_and568_y0;
  wire h_u_cla12_and569_y0;
  wire h_u_cla12_and570_y0;
  wire h_u_cla12_and571_y0;
  wire h_u_cla12_and572_y0;
  wire h_u_cla12_and573_y0;
  wire h_u_cla12_and574_y0;
  wire h_u_cla12_and575_y0;
  wire h_u_cla12_and576_y0;
  wire h_u_cla12_and577_y0;
  wire h_u_cla12_and578_y0;
  wire h_u_cla12_and579_y0;
  wire h_u_cla12_and580_y0;
  wire h_u_cla12_and581_y0;
  wire h_u_cla12_and582_y0;
  wire h_u_cla12_and583_y0;
  wire h_u_cla12_and584_y0;
  wire h_u_cla12_and585_y0;
  wire h_u_cla12_and586_y0;
  wire h_u_cla12_and587_y0;
  wire h_u_cla12_and588_y0;
  wire h_u_cla12_and589_y0;
  wire h_u_cla12_and590_y0;
  wire h_u_cla12_and591_y0;
  wire h_u_cla12_and592_y0;
  wire h_u_cla12_and593_y0;
  wire h_u_cla12_and594_y0;
  wire h_u_cla12_and595_y0;
  wire h_u_cla12_and596_y0;
  wire h_u_cla12_and597_y0;
  wire h_u_cla12_and598_y0;
  wire h_u_cla12_and599_y0;
  wire h_u_cla12_and600_y0;
  wire h_u_cla12_and601_y0;
  wire h_u_cla12_and602_y0;
  wire h_u_cla12_and603_y0;
  wire h_u_cla12_and604_y0;
  wire h_u_cla12_and605_y0;
  wire h_u_cla12_and606_y0;
  wire h_u_cla12_and607_y0;
  wire h_u_cla12_and608_y0;
  wire h_u_cla12_and609_y0;
  wire h_u_cla12_and610_y0;
  wire h_u_cla12_and611_y0;
  wire h_u_cla12_and612_y0;
  wire h_u_cla12_and613_y0;
  wire h_u_cla12_and614_y0;
  wire h_u_cla12_and615_y0;
  wire h_u_cla12_and616_y0;
  wire h_u_cla12_and617_y0;
  wire h_u_cla12_and618_y0;
  wire h_u_cla12_and619_y0;
  wire h_u_cla12_and620_y0;
  wire h_u_cla12_and621_y0;
  wire h_u_cla12_and622_y0;
  wire h_u_cla12_and623_y0;
  wire h_u_cla12_and624_y0;
  wire h_u_cla12_and625_y0;
  wire h_u_cla12_and626_y0;
  wire h_u_cla12_and627_y0;
  wire h_u_cla12_and628_y0;
  wire h_u_cla12_and629_y0;
  wire h_u_cla12_and630_y0;
  wire h_u_cla12_and631_y0;
  wire h_u_cla12_and632_y0;
  wire h_u_cla12_and633_y0;
  wire h_u_cla12_and634_y0;
  wire h_u_cla12_and635_y0;
  wire h_u_cla12_and636_y0;
  wire h_u_cla12_and637_y0;
  wire h_u_cla12_and638_y0;
  wire h_u_cla12_and639_y0;
  wire h_u_cla12_and640_y0;
  wire h_u_cla12_and641_y0;
  wire h_u_cla12_and642_y0;
  wire h_u_cla12_and643_y0;
  wire h_u_cla12_and644_y0;
  wire h_u_cla12_and645_y0;
  wire h_u_cla12_and646_y0;
  wire h_u_cla12_and647_y0;
  wire h_u_cla12_and648_y0;
  wire h_u_cla12_and649_y0;
  wire h_u_cla12_or66_y0;
  wire h_u_cla12_or67_y0;
  wire h_u_cla12_or68_y0;
  wire h_u_cla12_or69_y0;
  wire h_u_cla12_or70_y0;
  wire h_u_cla12_or71_y0;
  wire h_u_cla12_or72_y0;
  wire h_u_cla12_or73_y0;
  wire h_u_cla12_or74_y0;
  wire h_u_cla12_or75_y0;
  wire h_u_cla12_or76_y0;
  wire h_u_cla12_or77_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  constant_wire_value_0 constant_wire_value_0_constant_wire_0(a_0, b_0, constant_wire_0);
  pg_logic pg_logic_h_u_cla12_pg_logic0_y0(a_0, b_0, h_u_cla12_pg_logic0_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_pg_logic0_y2);
  xor_gate xor_gate_h_u_cla12_xor0_y0(h_u_cla12_pg_logic0_y2, constant_wire_0, h_u_cla12_xor0_y0);
  and_gate and_gate_h_u_cla12_and0_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and0_y0);
  or_gate or_gate_h_u_cla12_or0_y0(h_u_cla12_pg_logic0_y1, h_u_cla12_and0_y0, h_u_cla12_or0_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic1_y0(a_1, b_1, h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_pg_logic1_y2);
  xor_gate xor_gate_h_u_cla12_xor1_y0(h_u_cla12_pg_logic1_y2, h_u_cla12_or0_y0, h_u_cla12_xor1_y0);
  and_gate and_gate_h_u_cla12_and1_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and1_y0);
  and_gate and_gate_h_u_cla12_and2_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and2_y0);
  and_gate and_gate_h_u_cla12_and3_y0(h_u_cla12_and2_y0, h_u_cla12_and1_y0, h_u_cla12_and3_y0);
  and_gate and_gate_h_u_cla12_and4_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and4_y0);
  or_gate or_gate_h_u_cla12_or1_y0(h_u_cla12_and4_y0, h_u_cla12_and3_y0, h_u_cla12_or1_y0);
  or_gate or_gate_h_u_cla12_or2_y0(h_u_cla12_pg_logic1_y1, h_u_cla12_or1_y0, h_u_cla12_or2_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic2_y0(a_2, b_2, h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_pg_logic2_y2);
  xor_gate xor_gate_h_u_cla12_xor2_y0(h_u_cla12_pg_logic2_y2, h_u_cla12_or2_y0, h_u_cla12_xor2_y0);
  and_gate and_gate_h_u_cla12_and5_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and5_y0);
  and_gate and_gate_h_u_cla12_and6_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and6_y0);
  and_gate and_gate_h_u_cla12_and7_y0(h_u_cla12_and6_y0, h_u_cla12_and5_y0, h_u_cla12_and7_y0);
  and_gate and_gate_h_u_cla12_and8_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and8_y0);
  and_gate and_gate_h_u_cla12_and9_y0(h_u_cla12_and8_y0, h_u_cla12_and7_y0, h_u_cla12_and9_y0);
  and_gate and_gate_h_u_cla12_and10_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and10_y0);
  and_gate and_gate_h_u_cla12_and11_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and11_y0);
  and_gate and_gate_h_u_cla12_and12_y0(h_u_cla12_and11_y0, h_u_cla12_and10_y0, h_u_cla12_and12_y0);
  and_gate and_gate_h_u_cla12_and13_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and13_y0);
  or_gate or_gate_h_u_cla12_or3_y0(h_u_cla12_and13_y0, h_u_cla12_and9_y0, h_u_cla12_or3_y0);
  or_gate or_gate_h_u_cla12_or4_y0(h_u_cla12_or3_y0, h_u_cla12_and12_y0, h_u_cla12_or4_y0);
  or_gate or_gate_h_u_cla12_or5_y0(h_u_cla12_pg_logic2_y1, h_u_cla12_or4_y0, h_u_cla12_or5_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic3_y0(a_3, b_3, h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_pg_logic3_y2);
  xor_gate xor_gate_h_u_cla12_xor3_y0(h_u_cla12_pg_logic3_y2, h_u_cla12_or5_y0, h_u_cla12_xor3_y0);
  and_gate and_gate_h_u_cla12_and14_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and14_y0);
  and_gate and_gate_h_u_cla12_and15_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and15_y0);
  and_gate and_gate_h_u_cla12_and16_y0(h_u_cla12_and15_y0, h_u_cla12_and14_y0, h_u_cla12_and16_y0);
  and_gate and_gate_h_u_cla12_and17_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and17_y0);
  and_gate and_gate_h_u_cla12_and18_y0(h_u_cla12_and17_y0, h_u_cla12_and16_y0, h_u_cla12_and18_y0);
  and_gate and_gate_h_u_cla12_and19_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and19_y0);
  and_gate and_gate_h_u_cla12_and20_y0(h_u_cla12_and19_y0, h_u_cla12_and18_y0, h_u_cla12_and20_y0);
  and_gate and_gate_h_u_cla12_and21_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and21_y0);
  and_gate and_gate_h_u_cla12_and22_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and22_y0);
  and_gate and_gate_h_u_cla12_and23_y0(h_u_cla12_and22_y0, h_u_cla12_and21_y0, h_u_cla12_and23_y0);
  and_gate and_gate_h_u_cla12_and24_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and24_y0);
  and_gate and_gate_h_u_cla12_and25_y0(h_u_cla12_and24_y0, h_u_cla12_and23_y0, h_u_cla12_and25_y0);
  and_gate and_gate_h_u_cla12_and26_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and26_y0);
  and_gate and_gate_h_u_cla12_and27_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and27_y0);
  and_gate and_gate_h_u_cla12_and28_y0(h_u_cla12_and27_y0, h_u_cla12_and26_y0, h_u_cla12_and28_y0);
  and_gate and_gate_h_u_cla12_and29_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and29_y0);
  or_gate or_gate_h_u_cla12_or6_y0(h_u_cla12_and29_y0, h_u_cla12_and20_y0, h_u_cla12_or6_y0);
  or_gate or_gate_h_u_cla12_or7_y0(h_u_cla12_or6_y0, h_u_cla12_and25_y0, h_u_cla12_or7_y0);
  or_gate or_gate_h_u_cla12_or8_y0(h_u_cla12_or7_y0, h_u_cla12_and28_y0, h_u_cla12_or8_y0);
  or_gate or_gate_h_u_cla12_or9_y0(h_u_cla12_pg_logic3_y1, h_u_cla12_or8_y0, h_u_cla12_or9_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic4_y0(a_4, b_4, h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_pg_logic4_y2);
  xor_gate xor_gate_h_u_cla12_xor4_y0(h_u_cla12_pg_logic4_y2, h_u_cla12_or9_y0, h_u_cla12_xor4_y0);
  and_gate and_gate_h_u_cla12_and30_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and30_y0);
  and_gate and_gate_h_u_cla12_and31_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and31_y0);
  and_gate and_gate_h_u_cla12_and32_y0(h_u_cla12_and31_y0, h_u_cla12_and30_y0, h_u_cla12_and32_y0);
  and_gate and_gate_h_u_cla12_and33_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and33_y0);
  and_gate and_gate_h_u_cla12_and34_y0(h_u_cla12_and33_y0, h_u_cla12_and32_y0, h_u_cla12_and34_y0);
  and_gate and_gate_h_u_cla12_and35_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and35_y0);
  and_gate and_gate_h_u_cla12_and36_y0(h_u_cla12_and35_y0, h_u_cla12_and34_y0, h_u_cla12_and36_y0);
  and_gate and_gate_h_u_cla12_and37_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and37_y0);
  and_gate and_gate_h_u_cla12_and38_y0(h_u_cla12_and37_y0, h_u_cla12_and36_y0, h_u_cla12_and38_y0);
  and_gate and_gate_h_u_cla12_and39_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and39_y0);
  and_gate and_gate_h_u_cla12_and40_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and40_y0);
  and_gate and_gate_h_u_cla12_and41_y0(h_u_cla12_and40_y0, h_u_cla12_and39_y0, h_u_cla12_and41_y0);
  and_gate and_gate_h_u_cla12_and42_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and42_y0);
  and_gate and_gate_h_u_cla12_and43_y0(h_u_cla12_and42_y0, h_u_cla12_and41_y0, h_u_cla12_and43_y0);
  and_gate and_gate_h_u_cla12_and44_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and44_y0);
  and_gate and_gate_h_u_cla12_and45_y0(h_u_cla12_and44_y0, h_u_cla12_and43_y0, h_u_cla12_and45_y0);
  and_gate and_gate_h_u_cla12_and46_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and46_y0);
  and_gate and_gate_h_u_cla12_and47_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and47_y0);
  and_gate and_gate_h_u_cla12_and48_y0(h_u_cla12_and47_y0, h_u_cla12_and46_y0, h_u_cla12_and48_y0);
  and_gate and_gate_h_u_cla12_and49_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and49_y0);
  and_gate and_gate_h_u_cla12_and50_y0(h_u_cla12_and49_y0, h_u_cla12_and48_y0, h_u_cla12_and50_y0);
  and_gate and_gate_h_u_cla12_and51_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and51_y0);
  and_gate and_gate_h_u_cla12_and52_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and52_y0);
  and_gate and_gate_h_u_cla12_and53_y0(h_u_cla12_and52_y0, h_u_cla12_and51_y0, h_u_cla12_and53_y0);
  and_gate and_gate_h_u_cla12_and54_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and54_y0);
  or_gate or_gate_h_u_cla12_or10_y0(h_u_cla12_and54_y0, h_u_cla12_and38_y0, h_u_cla12_or10_y0);
  or_gate or_gate_h_u_cla12_or11_y0(h_u_cla12_or10_y0, h_u_cla12_and45_y0, h_u_cla12_or11_y0);
  or_gate or_gate_h_u_cla12_or12_y0(h_u_cla12_or11_y0, h_u_cla12_and50_y0, h_u_cla12_or12_y0);
  or_gate or_gate_h_u_cla12_or13_y0(h_u_cla12_or12_y0, h_u_cla12_and53_y0, h_u_cla12_or13_y0);
  or_gate or_gate_h_u_cla12_or14_y0(h_u_cla12_pg_logic4_y1, h_u_cla12_or13_y0, h_u_cla12_or14_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic5_y0(a_5, b_5, h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_pg_logic5_y2);
  xor_gate xor_gate_h_u_cla12_xor5_y0(h_u_cla12_pg_logic5_y2, h_u_cla12_or14_y0, h_u_cla12_xor5_y0);
  and_gate and_gate_h_u_cla12_and55_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and55_y0);
  and_gate and_gate_h_u_cla12_and56_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and56_y0);
  and_gate and_gate_h_u_cla12_and57_y0(h_u_cla12_and56_y0, h_u_cla12_and55_y0, h_u_cla12_and57_y0);
  and_gate and_gate_h_u_cla12_and58_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and58_y0);
  and_gate and_gate_h_u_cla12_and59_y0(h_u_cla12_and58_y0, h_u_cla12_and57_y0, h_u_cla12_and59_y0);
  and_gate and_gate_h_u_cla12_and60_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and60_y0);
  and_gate and_gate_h_u_cla12_and61_y0(h_u_cla12_and60_y0, h_u_cla12_and59_y0, h_u_cla12_and61_y0);
  and_gate and_gate_h_u_cla12_and62_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and62_y0);
  and_gate and_gate_h_u_cla12_and63_y0(h_u_cla12_and62_y0, h_u_cla12_and61_y0, h_u_cla12_and63_y0);
  and_gate and_gate_h_u_cla12_and64_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and64_y0);
  and_gate and_gate_h_u_cla12_and65_y0(h_u_cla12_and64_y0, h_u_cla12_and63_y0, h_u_cla12_and65_y0);
  and_gate and_gate_h_u_cla12_and66_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and66_y0);
  and_gate and_gate_h_u_cla12_and67_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and67_y0);
  and_gate and_gate_h_u_cla12_and68_y0(h_u_cla12_and67_y0, h_u_cla12_and66_y0, h_u_cla12_and68_y0);
  and_gate and_gate_h_u_cla12_and69_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and69_y0);
  and_gate and_gate_h_u_cla12_and70_y0(h_u_cla12_and69_y0, h_u_cla12_and68_y0, h_u_cla12_and70_y0);
  and_gate and_gate_h_u_cla12_and71_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and71_y0);
  and_gate and_gate_h_u_cla12_and72_y0(h_u_cla12_and71_y0, h_u_cla12_and70_y0, h_u_cla12_and72_y0);
  and_gate and_gate_h_u_cla12_and73_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and73_y0);
  and_gate and_gate_h_u_cla12_and74_y0(h_u_cla12_and73_y0, h_u_cla12_and72_y0, h_u_cla12_and74_y0);
  and_gate and_gate_h_u_cla12_and75_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and75_y0);
  and_gate and_gate_h_u_cla12_and76_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and76_y0);
  and_gate and_gate_h_u_cla12_and77_y0(h_u_cla12_and76_y0, h_u_cla12_and75_y0, h_u_cla12_and77_y0);
  and_gate and_gate_h_u_cla12_and78_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and78_y0);
  and_gate and_gate_h_u_cla12_and79_y0(h_u_cla12_and78_y0, h_u_cla12_and77_y0, h_u_cla12_and79_y0);
  and_gate and_gate_h_u_cla12_and80_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and80_y0);
  and_gate and_gate_h_u_cla12_and81_y0(h_u_cla12_and80_y0, h_u_cla12_and79_y0, h_u_cla12_and81_y0);
  and_gate and_gate_h_u_cla12_and82_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and82_y0);
  and_gate and_gate_h_u_cla12_and83_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and83_y0);
  and_gate and_gate_h_u_cla12_and84_y0(h_u_cla12_and83_y0, h_u_cla12_and82_y0, h_u_cla12_and84_y0);
  and_gate and_gate_h_u_cla12_and85_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and85_y0);
  and_gate and_gate_h_u_cla12_and86_y0(h_u_cla12_and85_y0, h_u_cla12_and84_y0, h_u_cla12_and86_y0);
  and_gate and_gate_h_u_cla12_and87_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and87_y0);
  and_gate and_gate_h_u_cla12_and88_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and88_y0);
  and_gate and_gate_h_u_cla12_and89_y0(h_u_cla12_and88_y0, h_u_cla12_and87_y0, h_u_cla12_and89_y0);
  and_gate and_gate_h_u_cla12_and90_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and90_y0);
  or_gate or_gate_h_u_cla12_or15_y0(h_u_cla12_and90_y0, h_u_cla12_and65_y0, h_u_cla12_or15_y0);
  or_gate or_gate_h_u_cla12_or16_y0(h_u_cla12_or15_y0, h_u_cla12_and74_y0, h_u_cla12_or16_y0);
  or_gate or_gate_h_u_cla12_or17_y0(h_u_cla12_or16_y0, h_u_cla12_and81_y0, h_u_cla12_or17_y0);
  or_gate or_gate_h_u_cla12_or18_y0(h_u_cla12_or17_y0, h_u_cla12_and86_y0, h_u_cla12_or18_y0);
  or_gate or_gate_h_u_cla12_or19_y0(h_u_cla12_or18_y0, h_u_cla12_and89_y0, h_u_cla12_or19_y0);
  or_gate or_gate_h_u_cla12_or20_y0(h_u_cla12_pg_logic5_y1, h_u_cla12_or19_y0, h_u_cla12_or20_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic6_y0(a_6, b_6, h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_pg_logic6_y2);
  xor_gate xor_gate_h_u_cla12_xor6_y0(h_u_cla12_pg_logic6_y2, h_u_cla12_or20_y0, h_u_cla12_xor6_y0);
  and_gate and_gate_h_u_cla12_and91_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and91_y0);
  and_gate and_gate_h_u_cla12_and92_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and92_y0);
  and_gate and_gate_h_u_cla12_and93_y0(h_u_cla12_and92_y0, h_u_cla12_and91_y0, h_u_cla12_and93_y0);
  and_gate and_gate_h_u_cla12_and94_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and94_y0);
  and_gate and_gate_h_u_cla12_and95_y0(h_u_cla12_and94_y0, h_u_cla12_and93_y0, h_u_cla12_and95_y0);
  and_gate and_gate_h_u_cla12_and96_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and96_y0);
  and_gate and_gate_h_u_cla12_and97_y0(h_u_cla12_and96_y0, h_u_cla12_and95_y0, h_u_cla12_and97_y0);
  and_gate and_gate_h_u_cla12_and98_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and98_y0);
  and_gate and_gate_h_u_cla12_and99_y0(h_u_cla12_and98_y0, h_u_cla12_and97_y0, h_u_cla12_and99_y0);
  and_gate and_gate_h_u_cla12_and100_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and100_y0);
  and_gate and_gate_h_u_cla12_and101_y0(h_u_cla12_and100_y0, h_u_cla12_and99_y0, h_u_cla12_and101_y0);
  and_gate and_gate_h_u_cla12_and102_y0(h_u_cla12_pg_logic6_y0, constant_wire_0, h_u_cla12_and102_y0);
  and_gate and_gate_h_u_cla12_and103_y0(h_u_cla12_and102_y0, h_u_cla12_and101_y0, h_u_cla12_and103_y0);
  and_gate and_gate_h_u_cla12_and104_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and104_y0);
  and_gate and_gate_h_u_cla12_and105_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and105_y0);
  and_gate and_gate_h_u_cla12_and106_y0(h_u_cla12_and105_y0, h_u_cla12_and104_y0, h_u_cla12_and106_y0);
  and_gate and_gate_h_u_cla12_and107_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and107_y0);
  and_gate and_gate_h_u_cla12_and108_y0(h_u_cla12_and107_y0, h_u_cla12_and106_y0, h_u_cla12_and108_y0);
  and_gate and_gate_h_u_cla12_and109_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and109_y0);
  and_gate and_gate_h_u_cla12_and110_y0(h_u_cla12_and109_y0, h_u_cla12_and108_y0, h_u_cla12_and110_y0);
  and_gate and_gate_h_u_cla12_and111_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and111_y0);
  and_gate and_gate_h_u_cla12_and112_y0(h_u_cla12_and111_y0, h_u_cla12_and110_y0, h_u_cla12_and112_y0);
  and_gate and_gate_h_u_cla12_and113_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and113_y0);
  and_gate and_gate_h_u_cla12_and114_y0(h_u_cla12_and113_y0, h_u_cla12_and112_y0, h_u_cla12_and114_y0);
  and_gate and_gate_h_u_cla12_and115_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and115_y0);
  and_gate and_gate_h_u_cla12_and116_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and116_y0);
  and_gate and_gate_h_u_cla12_and117_y0(h_u_cla12_and116_y0, h_u_cla12_and115_y0, h_u_cla12_and117_y0);
  and_gate and_gate_h_u_cla12_and118_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and118_y0);
  and_gate and_gate_h_u_cla12_and119_y0(h_u_cla12_and118_y0, h_u_cla12_and117_y0, h_u_cla12_and119_y0);
  and_gate and_gate_h_u_cla12_and120_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and120_y0);
  and_gate and_gate_h_u_cla12_and121_y0(h_u_cla12_and120_y0, h_u_cla12_and119_y0, h_u_cla12_and121_y0);
  and_gate and_gate_h_u_cla12_and122_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and122_y0);
  and_gate and_gate_h_u_cla12_and123_y0(h_u_cla12_and122_y0, h_u_cla12_and121_y0, h_u_cla12_and123_y0);
  and_gate and_gate_h_u_cla12_and124_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and124_y0);
  and_gate and_gate_h_u_cla12_and125_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and125_y0);
  and_gate and_gate_h_u_cla12_and126_y0(h_u_cla12_and125_y0, h_u_cla12_and124_y0, h_u_cla12_and126_y0);
  and_gate and_gate_h_u_cla12_and127_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and127_y0);
  and_gate and_gate_h_u_cla12_and128_y0(h_u_cla12_and127_y0, h_u_cla12_and126_y0, h_u_cla12_and128_y0);
  and_gate and_gate_h_u_cla12_and129_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and129_y0);
  and_gate and_gate_h_u_cla12_and130_y0(h_u_cla12_and129_y0, h_u_cla12_and128_y0, h_u_cla12_and130_y0);
  and_gate and_gate_h_u_cla12_and131_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and131_y0);
  and_gate and_gate_h_u_cla12_and132_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and132_y0);
  and_gate and_gate_h_u_cla12_and133_y0(h_u_cla12_and132_y0, h_u_cla12_and131_y0, h_u_cla12_and133_y0);
  and_gate and_gate_h_u_cla12_and134_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and134_y0);
  and_gate and_gate_h_u_cla12_and135_y0(h_u_cla12_and134_y0, h_u_cla12_and133_y0, h_u_cla12_and135_y0);
  and_gate and_gate_h_u_cla12_and136_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and136_y0);
  and_gate and_gate_h_u_cla12_and137_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and137_y0);
  and_gate and_gate_h_u_cla12_and138_y0(h_u_cla12_and137_y0, h_u_cla12_and136_y0, h_u_cla12_and138_y0);
  and_gate and_gate_h_u_cla12_and139_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and139_y0);
  or_gate or_gate_h_u_cla12_or21_y0(h_u_cla12_and139_y0, h_u_cla12_and103_y0, h_u_cla12_or21_y0);
  or_gate or_gate_h_u_cla12_or22_y0(h_u_cla12_or21_y0, h_u_cla12_and114_y0, h_u_cla12_or22_y0);
  or_gate or_gate_h_u_cla12_or23_y0(h_u_cla12_or22_y0, h_u_cla12_and123_y0, h_u_cla12_or23_y0);
  or_gate or_gate_h_u_cla12_or24_y0(h_u_cla12_or23_y0, h_u_cla12_and130_y0, h_u_cla12_or24_y0);
  or_gate or_gate_h_u_cla12_or25_y0(h_u_cla12_or24_y0, h_u_cla12_and135_y0, h_u_cla12_or25_y0);
  or_gate or_gate_h_u_cla12_or26_y0(h_u_cla12_or25_y0, h_u_cla12_and138_y0, h_u_cla12_or26_y0);
  or_gate or_gate_h_u_cla12_or27_y0(h_u_cla12_pg_logic6_y1, h_u_cla12_or26_y0, h_u_cla12_or27_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic7_y0(a_7, b_7, h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_pg_logic7_y2);
  xor_gate xor_gate_h_u_cla12_xor7_y0(h_u_cla12_pg_logic7_y2, h_u_cla12_or27_y0, h_u_cla12_xor7_y0);
  and_gate and_gate_h_u_cla12_and140_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and140_y0);
  and_gate and_gate_h_u_cla12_and141_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and141_y0);
  and_gate and_gate_h_u_cla12_and142_y0(h_u_cla12_and141_y0, h_u_cla12_and140_y0, h_u_cla12_and142_y0);
  and_gate and_gate_h_u_cla12_and143_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and143_y0);
  and_gate and_gate_h_u_cla12_and144_y0(h_u_cla12_and143_y0, h_u_cla12_and142_y0, h_u_cla12_and144_y0);
  and_gate and_gate_h_u_cla12_and145_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and145_y0);
  and_gate and_gate_h_u_cla12_and146_y0(h_u_cla12_and145_y0, h_u_cla12_and144_y0, h_u_cla12_and146_y0);
  and_gate and_gate_h_u_cla12_and147_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and147_y0);
  and_gate and_gate_h_u_cla12_and148_y0(h_u_cla12_and147_y0, h_u_cla12_and146_y0, h_u_cla12_and148_y0);
  and_gate and_gate_h_u_cla12_and149_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and149_y0);
  and_gate and_gate_h_u_cla12_and150_y0(h_u_cla12_and149_y0, h_u_cla12_and148_y0, h_u_cla12_and150_y0);
  and_gate and_gate_h_u_cla12_and151_y0(h_u_cla12_pg_logic6_y0, constant_wire_0, h_u_cla12_and151_y0);
  and_gate and_gate_h_u_cla12_and152_y0(h_u_cla12_and151_y0, h_u_cla12_and150_y0, h_u_cla12_and152_y0);
  and_gate and_gate_h_u_cla12_and153_y0(h_u_cla12_pg_logic7_y0, constant_wire_0, h_u_cla12_and153_y0);
  and_gate and_gate_h_u_cla12_and154_y0(h_u_cla12_and153_y0, h_u_cla12_and152_y0, h_u_cla12_and154_y0);
  and_gate and_gate_h_u_cla12_and155_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and155_y0);
  and_gate and_gate_h_u_cla12_and156_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and156_y0);
  and_gate and_gate_h_u_cla12_and157_y0(h_u_cla12_and156_y0, h_u_cla12_and155_y0, h_u_cla12_and157_y0);
  and_gate and_gate_h_u_cla12_and158_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and158_y0);
  and_gate and_gate_h_u_cla12_and159_y0(h_u_cla12_and158_y0, h_u_cla12_and157_y0, h_u_cla12_and159_y0);
  and_gate and_gate_h_u_cla12_and160_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and160_y0);
  and_gate and_gate_h_u_cla12_and161_y0(h_u_cla12_and160_y0, h_u_cla12_and159_y0, h_u_cla12_and161_y0);
  and_gate and_gate_h_u_cla12_and162_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and162_y0);
  and_gate and_gate_h_u_cla12_and163_y0(h_u_cla12_and162_y0, h_u_cla12_and161_y0, h_u_cla12_and163_y0);
  and_gate and_gate_h_u_cla12_and164_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and164_y0);
  and_gate and_gate_h_u_cla12_and165_y0(h_u_cla12_and164_y0, h_u_cla12_and163_y0, h_u_cla12_and165_y0);
  and_gate and_gate_h_u_cla12_and166_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and166_y0);
  and_gate and_gate_h_u_cla12_and167_y0(h_u_cla12_and166_y0, h_u_cla12_and165_y0, h_u_cla12_and167_y0);
  and_gate and_gate_h_u_cla12_and168_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and168_y0);
  and_gate and_gate_h_u_cla12_and169_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and169_y0);
  and_gate and_gate_h_u_cla12_and170_y0(h_u_cla12_and169_y0, h_u_cla12_and168_y0, h_u_cla12_and170_y0);
  and_gate and_gate_h_u_cla12_and171_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and171_y0);
  and_gate and_gate_h_u_cla12_and172_y0(h_u_cla12_and171_y0, h_u_cla12_and170_y0, h_u_cla12_and172_y0);
  and_gate and_gate_h_u_cla12_and173_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and173_y0);
  and_gate and_gate_h_u_cla12_and174_y0(h_u_cla12_and173_y0, h_u_cla12_and172_y0, h_u_cla12_and174_y0);
  and_gate and_gate_h_u_cla12_and175_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and175_y0);
  and_gate and_gate_h_u_cla12_and176_y0(h_u_cla12_and175_y0, h_u_cla12_and174_y0, h_u_cla12_and176_y0);
  and_gate and_gate_h_u_cla12_and177_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and177_y0);
  and_gate and_gate_h_u_cla12_and178_y0(h_u_cla12_and177_y0, h_u_cla12_and176_y0, h_u_cla12_and178_y0);
  and_gate and_gate_h_u_cla12_and179_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and179_y0);
  and_gate and_gate_h_u_cla12_and180_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and180_y0);
  and_gate and_gate_h_u_cla12_and181_y0(h_u_cla12_and180_y0, h_u_cla12_and179_y0, h_u_cla12_and181_y0);
  and_gate and_gate_h_u_cla12_and182_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and182_y0);
  and_gate and_gate_h_u_cla12_and183_y0(h_u_cla12_and182_y0, h_u_cla12_and181_y0, h_u_cla12_and183_y0);
  and_gate and_gate_h_u_cla12_and184_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and184_y0);
  and_gate and_gate_h_u_cla12_and185_y0(h_u_cla12_and184_y0, h_u_cla12_and183_y0, h_u_cla12_and185_y0);
  and_gate and_gate_h_u_cla12_and186_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and186_y0);
  and_gate and_gate_h_u_cla12_and187_y0(h_u_cla12_and186_y0, h_u_cla12_and185_y0, h_u_cla12_and187_y0);
  and_gate and_gate_h_u_cla12_and188_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and188_y0);
  and_gate and_gate_h_u_cla12_and189_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and189_y0);
  and_gate and_gate_h_u_cla12_and190_y0(h_u_cla12_and189_y0, h_u_cla12_and188_y0, h_u_cla12_and190_y0);
  and_gate and_gate_h_u_cla12_and191_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and191_y0);
  and_gate and_gate_h_u_cla12_and192_y0(h_u_cla12_and191_y0, h_u_cla12_and190_y0, h_u_cla12_and192_y0);
  and_gate and_gate_h_u_cla12_and193_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and193_y0);
  and_gate and_gate_h_u_cla12_and194_y0(h_u_cla12_and193_y0, h_u_cla12_and192_y0, h_u_cla12_and194_y0);
  and_gate and_gate_h_u_cla12_and195_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and195_y0);
  and_gate and_gate_h_u_cla12_and196_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and196_y0);
  and_gate and_gate_h_u_cla12_and197_y0(h_u_cla12_and196_y0, h_u_cla12_and195_y0, h_u_cla12_and197_y0);
  and_gate and_gate_h_u_cla12_and198_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and198_y0);
  and_gate and_gate_h_u_cla12_and199_y0(h_u_cla12_and198_y0, h_u_cla12_and197_y0, h_u_cla12_and199_y0);
  and_gate and_gate_h_u_cla12_and200_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and200_y0);
  and_gate and_gate_h_u_cla12_and201_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and201_y0);
  and_gate and_gate_h_u_cla12_and202_y0(h_u_cla12_and201_y0, h_u_cla12_and200_y0, h_u_cla12_and202_y0);
  and_gate and_gate_h_u_cla12_and203_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and203_y0);
  or_gate or_gate_h_u_cla12_or28_y0(h_u_cla12_and203_y0, h_u_cla12_and154_y0, h_u_cla12_or28_y0);
  or_gate or_gate_h_u_cla12_or29_y0(h_u_cla12_or28_y0, h_u_cla12_and167_y0, h_u_cla12_or29_y0);
  or_gate or_gate_h_u_cla12_or30_y0(h_u_cla12_or29_y0, h_u_cla12_and178_y0, h_u_cla12_or30_y0);
  or_gate or_gate_h_u_cla12_or31_y0(h_u_cla12_or30_y0, h_u_cla12_and187_y0, h_u_cla12_or31_y0);
  or_gate or_gate_h_u_cla12_or32_y0(h_u_cla12_or31_y0, h_u_cla12_and194_y0, h_u_cla12_or32_y0);
  or_gate or_gate_h_u_cla12_or33_y0(h_u_cla12_or32_y0, h_u_cla12_and199_y0, h_u_cla12_or33_y0);
  or_gate or_gate_h_u_cla12_or34_y0(h_u_cla12_or33_y0, h_u_cla12_and202_y0, h_u_cla12_or34_y0);
  or_gate or_gate_h_u_cla12_or35_y0(h_u_cla12_pg_logic7_y1, h_u_cla12_or34_y0, h_u_cla12_or35_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic8_y0(a_8, b_8, h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_pg_logic8_y2);
  xor_gate xor_gate_h_u_cla12_xor8_y0(h_u_cla12_pg_logic8_y2, h_u_cla12_or35_y0, h_u_cla12_xor8_y0);
  and_gate and_gate_h_u_cla12_and204_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and204_y0);
  and_gate and_gate_h_u_cla12_and205_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and205_y0);
  and_gate and_gate_h_u_cla12_and206_y0(h_u_cla12_and205_y0, h_u_cla12_and204_y0, h_u_cla12_and206_y0);
  and_gate and_gate_h_u_cla12_and207_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and207_y0);
  and_gate and_gate_h_u_cla12_and208_y0(h_u_cla12_and207_y0, h_u_cla12_and206_y0, h_u_cla12_and208_y0);
  and_gate and_gate_h_u_cla12_and209_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and209_y0);
  and_gate and_gate_h_u_cla12_and210_y0(h_u_cla12_and209_y0, h_u_cla12_and208_y0, h_u_cla12_and210_y0);
  and_gate and_gate_h_u_cla12_and211_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and211_y0);
  and_gate and_gate_h_u_cla12_and212_y0(h_u_cla12_and211_y0, h_u_cla12_and210_y0, h_u_cla12_and212_y0);
  and_gate and_gate_h_u_cla12_and213_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and213_y0);
  and_gate and_gate_h_u_cla12_and214_y0(h_u_cla12_and213_y0, h_u_cla12_and212_y0, h_u_cla12_and214_y0);
  and_gate and_gate_h_u_cla12_and215_y0(h_u_cla12_pg_logic6_y0, constant_wire_0, h_u_cla12_and215_y0);
  and_gate and_gate_h_u_cla12_and216_y0(h_u_cla12_and215_y0, h_u_cla12_and214_y0, h_u_cla12_and216_y0);
  and_gate and_gate_h_u_cla12_and217_y0(h_u_cla12_pg_logic7_y0, constant_wire_0, h_u_cla12_and217_y0);
  and_gate and_gate_h_u_cla12_and218_y0(h_u_cla12_and217_y0, h_u_cla12_and216_y0, h_u_cla12_and218_y0);
  and_gate and_gate_h_u_cla12_and219_y0(h_u_cla12_pg_logic8_y0, constant_wire_0, h_u_cla12_and219_y0);
  and_gate and_gate_h_u_cla12_and220_y0(h_u_cla12_and219_y0, h_u_cla12_and218_y0, h_u_cla12_and220_y0);
  and_gate and_gate_h_u_cla12_and221_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and221_y0);
  and_gate and_gate_h_u_cla12_and222_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and222_y0);
  and_gate and_gate_h_u_cla12_and223_y0(h_u_cla12_and222_y0, h_u_cla12_and221_y0, h_u_cla12_and223_y0);
  and_gate and_gate_h_u_cla12_and224_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and224_y0);
  and_gate and_gate_h_u_cla12_and225_y0(h_u_cla12_and224_y0, h_u_cla12_and223_y0, h_u_cla12_and225_y0);
  and_gate and_gate_h_u_cla12_and226_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and226_y0);
  and_gate and_gate_h_u_cla12_and227_y0(h_u_cla12_and226_y0, h_u_cla12_and225_y0, h_u_cla12_and227_y0);
  and_gate and_gate_h_u_cla12_and228_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and228_y0);
  and_gate and_gate_h_u_cla12_and229_y0(h_u_cla12_and228_y0, h_u_cla12_and227_y0, h_u_cla12_and229_y0);
  and_gate and_gate_h_u_cla12_and230_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and230_y0);
  and_gate and_gate_h_u_cla12_and231_y0(h_u_cla12_and230_y0, h_u_cla12_and229_y0, h_u_cla12_and231_y0);
  and_gate and_gate_h_u_cla12_and232_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and232_y0);
  and_gate and_gate_h_u_cla12_and233_y0(h_u_cla12_and232_y0, h_u_cla12_and231_y0, h_u_cla12_and233_y0);
  and_gate and_gate_h_u_cla12_and234_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and234_y0);
  and_gate and_gate_h_u_cla12_and235_y0(h_u_cla12_and234_y0, h_u_cla12_and233_y0, h_u_cla12_and235_y0);
  and_gate and_gate_h_u_cla12_and236_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and236_y0);
  and_gate and_gate_h_u_cla12_and237_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and237_y0);
  and_gate and_gate_h_u_cla12_and238_y0(h_u_cla12_and237_y0, h_u_cla12_and236_y0, h_u_cla12_and238_y0);
  and_gate and_gate_h_u_cla12_and239_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and239_y0);
  and_gate and_gate_h_u_cla12_and240_y0(h_u_cla12_and239_y0, h_u_cla12_and238_y0, h_u_cla12_and240_y0);
  and_gate and_gate_h_u_cla12_and241_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and241_y0);
  and_gate and_gate_h_u_cla12_and242_y0(h_u_cla12_and241_y0, h_u_cla12_and240_y0, h_u_cla12_and242_y0);
  and_gate and_gate_h_u_cla12_and243_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and243_y0);
  and_gate and_gate_h_u_cla12_and244_y0(h_u_cla12_and243_y0, h_u_cla12_and242_y0, h_u_cla12_and244_y0);
  and_gate and_gate_h_u_cla12_and245_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and245_y0);
  and_gate and_gate_h_u_cla12_and246_y0(h_u_cla12_and245_y0, h_u_cla12_and244_y0, h_u_cla12_and246_y0);
  and_gate and_gate_h_u_cla12_and247_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and247_y0);
  and_gate and_gate_h_u_cla12_and248_y0(h_u_cla12_and247_y0, h_u_cla12_and246_y0, h_u_cla12_and248_y0);
  and_gate and_gate_h_u_cla12_and249_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and249_y0);
  and_gate and_gate_h_u_cla12_and250_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and250_y0);
  and_gate and_gate_h_u_cla12_and251_y0(h_u_cla12_and250_y0, h_u_cla12_and249_y0, h_u_cla12_and251_y0);
  and_gate and_gate_h_u_cla12_and252_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and252_y0);
  and_gate and_gate_h_u_cla12_and253_y0(h_u_cla12_and252_y0, h_u_cla12_and251_y0, h_u_cla12_and253_y0);
  and_gate and_gate_h_u_cla12_and254_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and254_y0);
  and_gate and_gate_h_u_cla12_and255_y0(h_u_cla12_and254_y0, h_u_cla12_and253_y0, h_u_cla12_and255_y0);
  and_gate and_gate_h_u_cla12_and256_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and256_y0);
  and_gate and_gate_h_u_cla12_and257_y0(h_u_cla12_and256_y0, h_u_cla12_and255_y0, h_u_cla12_and257_y0);
  and_gate and_gate_h_u_cla12_and258_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and258_y0);
  and_gate and_gate_h_u_cla12_and259_y0(h_u_cla12_and258_y0, h_u_cla12_and257_y0, h_u_cla12_and259_y0);
  and_gate and_gate_h_u_cla12_and260_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and260_y0);
  and_gate and_gate_h_u_cla12_and261_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and261_y0);
  and_gate and_gate_h_u_cla12_and262_y0(h_u_cla12_and261_y0, h_u_cla12_and260_y0, h_u_cla12_and262_y0);
  and_gate and_gate_h_u_cla12_and263_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and263_y0);
  and_gate and_gate_h_u_cla12_and264_y0(h_u_cla12_and263_y0, h_u_cla12_and262_y0, h_u_cla12_and264_y0);
  and_gate and_gate_h_u_cla12_and265_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and265_y0);
  and_gate and_gate_h_u_cla12_and266_y0(h_u_cla12_and265_y0, h_u_cla12_and264_y0, h_u_cla12_and266_y0);
  and_gate and_gate_h_u_cla12_and267_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and267_y0);
  and_gate and_gate_h_u_cla12_and268_y0(h_u_cla12_and267_y0, h_u_cla12_and266_y0, h_u_cla12_and268_y0);
  and_gate and_gate_h_u_cla12_and269_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and269_y0);
  and_gate and_gate_h_u_cla12_and270_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and270_y0);
  and_gate and_gate_h_u_cla12_and271_y0(h_u_cla12_and270_y0, h_u_cla12_and269_y0, h_u_cla12_and271_y0);
  and_gate and_gate_h_u_cla12_and272_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and272_y0);
  and_gate and_gate_h_u_cla12_and273_y0(h_u_cla12_and272_y0, h_u_cla12_and271_y0, h_u_cla12_and273_y0);
  and_gate and_gate_h_u_cla12_and274_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and274_y0);
  and_gate and_gate_h_u_cla12_and275_y0(h_u_cla12_and274_y0, h_u_cla12_and273_y0, h_u_cla12_and275_y0);
  and_gate and_gate_h_u_cla12_and276_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and276_y0);
  and_gate and_gate_h_u_cla12_and277_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and277_y0);
  and_gate and_gate_h_u_cla12_and278_y0(h_u_cla12_and277_y0, h_u_cla12_and276_y0, h_u_cla12_and278_y0);
  and_gate and_gate_h_u_cla12_and279_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and279_y0);
  and_gate and_gate_h_u_cla12_and280_y0(h_u_cla12_and279_y0, h_u_cla12_and278_y0, h_u_cla12_and280_y0);
  and_gate and_gate_h_u_cla12_and281_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and281_y0);
  and_gate and_gate_h_u_cla12_and282_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and282_y0);
  and_gate and_gate_h_u_cla12_and283_y0(h_u_cla12_and282_y0, h_u_cla12_and281_y0, h_u_cla12_and283_y0);
  and_gate and_gate_h_u_cla12_and284_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and284_y0);
  or_gate or_gate_h_u_cla12_or36_y0(h_u_cla12_and284_y0, h_u_cla12_and220_y0, h_u_cla12_or36_y0);
  or_gate or_gate_h_u_cla12_or37_y0(h_u_cla12_or36_y0, h_u_cla12_and235_y0, h_u_cla12_or37_y0);
  or_gate or_gate_h_u_cla12_or38_y0(h_u_cla12_or37_y0, h_u_cla12_and248_y0, h_u_cla12_or38_y0);
  or_gate or_gate_h_u_cla12_or39_y0(h_u_cla12_or38_y0, h_u_cla12_and259_y0, h_u_cla12_or39_y0);
  or_gate or_gate_h_u_cla12_or40_y0(h_u_cla12_or39_y0, h_u_cla12_and268_y0, h_u_cla12_or40_y0);
  or_gate or_gate_h_u_cla12_or41_y0(h_u_cla12_or40_y0, h_u_cla12_and275_y0, h_u_cla12_or41_y0);
  or_gate or_gate_h_u_cla12_or42_y0(h_u_cla12_or41_y0, h_u_cla12_and280_y0, h_u_cla12_or42_y0);
  or_gate or_gate_h_u_cla12_or43_y0(h_u_cla12_or42_y0, h_u_cla12_and283_y0, h_u_cla12_or43_y0);
  or_gate or_gate_h_u_cla12_or44_y0(h_u_cla12_pg_logic8_y1, h_u_cla12_or43_y0, h_u_cla12_or44_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic9_y0(a_9, b_9, h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic9_y1, h_u_cla12_pg_logic9_y2);
  xor_gate xor_gate_h_u_cla12_xor9_y0(h_u_cla12_pg_logic9_y2, h_u_cla12_or44_y0, h_u_cla12_xor9_y0);
  and_gate and_gate_h_u_cla12_and285_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and285_y0);
  and_gate and_gate_h_u_cla12_and286_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and286_y0);
  and_gate and_gate_h_u_cla12_and287_y0(h_u_cla12_and286_y0, h_u_cla12_and285_y0, h_u_cla12_and287_y0);
  and_gate and_gate_h_u_cla12_and288_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and288_y0);
  and_gate and_gate_h_u_cla12_and289_y0(h_u_cla12_and288_y0, h_u_cla12_and287_y0, h_u_cla12_and289_y0);
  and_gate and_gate_h_u_cla12_and290_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and290_y0);
  and_gate and_gate_h_u_cla12_and291_y0(h_u_cla12_and290_y0, h_u_cla12_and289_y0, h_u_cla12_and291_y0);
  and_gate and_gate_h_u_cla12_and292_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and292_y0);
  and_gate and_gate_h_u_cla12_and293_y0(h_u_cla12_and292_y0, h_u_cla12_and291_y0, h_u_cla12_and293_y0);
  and_gate and_gate_h_u_cla12_and294_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and294_y0);
  and_gate and_gate_h_u_cla12_and295_y0(h_u_cla12_and294_y0, h_u_cla12_and293_y0, h_u_cla12_and295_y0);
  and_gate and_gate_h_u_cla12_and296_y0(h_u_cla12_pg_logic6_y0, constant_wire_0, h_u_cla12_and296_y0);
  and_gate and_gate_h_u_cla12_and297_y0(h_u_cla12_and296_y0, h_u_cla12_and295_y0, h_u_cla12_and297_y0);
  and_gate and_gate_h_u_cla12_and298_y0(h_u_cla12_pg_logic7_y0, constant_wire_0, h_u_cla12_and298_y0);
  and_gate and_gate_h_u_cla12_and299_y0(h_u_cla12_and298_y0, h_u_cla12_and297_y0, h_u_cla12_and299_y0);
  and_gate and_gate_h_u_cla12_and300_y0(h_u_cla12_pg_logic8_y0, constant_wire_0, h_u_cla12_and300_y0);
  and_gate and_gate_h_u_cla12_and301_y0(h_u_cla12_and300_y0, h_u_cla12_and299_y0, h_u_cla12_and301_y0);
  and_gate and_gate_h_u_cla12_and302_y0(h_u_cla12_pg_logic9_y0, constant_wire_0, h_u_cla12_and302_y0);
  and_gate and_gate_h_u_cla12_and303_y0(h_u_cla12_and302_y0, h_u_cla12_and301_y0, h_u_cla12_and303_y0);
  and_gate and_gate_h_u_cla12_and304_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and304_y0);
  and_gate and_gate_h_u_cla12_and305_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and305_y0);
  and_gate and_gate_h_u_cla12_and306_y0(h_u_cla12_and305_y0, h_u_cla12_and304_y0, h_u_cla12_and306_y0);
  and_gate and_gate_h_u_cla12_and307_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and307_y0);
  and_gate and_gate_h_u_cla12_and308_y0(h_u_cla12_and307_y0, h_u_cla12_and306_y0, h_u_cla12_and308_y0);
  and_gate and_gate_h_u_cla12_and309_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and309_y0);
  and_gate and_gate_h_u_cla12_and310_y0(h_u_cla12_and309_y0, h_u_cla12_and308_y0, h_u_cla12_and310_y0);
  and_gate and_gate_h_u_cla12_and311_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and311_y0);
  and_gate and_gate_h_u_cla12_and312_y0(h_u_cla12_and311_y0, h_u_cla12_and310_y0, h_u_cla12_and312_y0);
  and_gate and_gate_h_u_cla12_and313_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and313_y0);
  and_gate and_gate_h_u_cla12_and314_y0(h_u_cla12_and313_y0, h_u_cla12_and312_y0, h_u_cla12_and314_y0);
  and_gate and_gate_h_u_cla12_and315_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and315_y0);
  and_gate and_gate_h_u_cla12_and316_y0(h_u_cla12_and315_y0, h_u_cla12_and314_y0, h_u_cla12_and316_y0);
  and_gate and_gate_h_u_cla12_and317_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and317_y0);
  and_gate and_gate_h_u_cla12_and318_y0(h_u_cla12_and317_y0, h_u_cla12_and316_y0, h_u_cla12_and318_y0);
  and_gate and_gate_h_u_cla12_and319_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and319_y0);
  and_gate and_gate_h_u_cla12_and320_y0(h_u_cla12_and319_y0, h_u_cla12_and318_y0, h_u_cla12_and320_y0);
  and_gate and_gate_h_u_cla12_and321_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and321_y0);
  and_gate and_gate_h_u_cla12_and322_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and322_y0);
  and_gate and_gate_h_u_cla12_and323_y0(h_u_cla12_and322_y0, h_u_cla12_and321_y0, h_u_cla12_and323_y0);
  and_gate and_gate_h_u_cla12_and324_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and324_y0);
  and_gate and_gate_h_u_cla12_and325_y0(h_u_cla12_and324_y0, h_u_cla12_and323_y0, h_u_cla12_and325_y0);
  and_gate and_gate_h_u_cla12_and326_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and326_y0);
  and_gate and_gate_h_u_cla12_and327_y0(h_u_cla12_and326_y0, h_u_cla12_and325_y0, h_u_cla12_and327_y0);
  and_gate and_gate_h_u_cla12_and328_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and328_y0);
  and_gate and_gate_h_u_cla12_and329_y0(h_u_cla12_and328_y0, h_u_cla12_and327_y0, h_u_cla12_and329_y0);
  and_gate and_gate_h_u_cla12_and330_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and330_y0);
  and_gate and_gate_h_u_cla12_and331_y0(h_u_cla12_and330_y0, h_u_cla12_and329_y0, h_u_cla12_and331_y0);
  and_gate and_gate_h_u_cla12_and332_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and332_y0);
  and_gate and_gate_h_u_cla12_and333_y0(h_u_cla12_and332_y0, h_u_cla12_and331_y0, h_u_cla12_and333_y0);
  and_gate and_gate_h_u_cla12_and334_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and334_y0);
  and_gate and_gate_h_u_cla12_and335_y0(h_u_cla12_and334_y0, h_u_cla12_and333_y0, h_u_cla12_and335_y0);
  and_gate and_gate_h_u_cla12_and336_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and336_y0);
  and_gate and_gate_h_u_cla12_and337_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and337_y0);
  and_gate and_gate_h_u_cla12_and338_y0(h_u_cla12_and337_y0, h_u_cla12_and336_y0, h_u_cla12_and338_y0);
  and_gate and_gate_h_u_cla12_and339_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and339_y0);
  and_gate and_gate_h_u_cla12_and340_y0(h_u_cla12_and339_y0, h_u_cla12_and338_y0, h_u_cla12_and340_y0);
  and_gate and_gate_h_u_cla12_and341_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and341_y0);
  and_gate and_gate_h_u_cla12_and342_y0(h_u_cla12_and341_y0, h_u_cla12_and340_y0, h_u_cla12_and342_y0);
  and_gate and_gate_h_u_cla12_and343_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and343_y0);
  and_gate and_gate_h_u_cla12_and344_y0(h_u_cla12_and343_y0, h_u_cla12_and342_y0, h_u_cla12_and344_y0);
  and_gate and_gate_h_u_cla12_and345_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and345_y0);
  and_gate and_gate_h_u_cla12_and346_y0(h_u_cla12_and345_y0, h_u_cla12_and344_y0, h_u_cla12_and346_y0);
  and_gate and_gate_h_u_cla12_and347_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and347_y0);
  and_gate and_gate_h_u_cla12_and348_y0(h_u_cla12_and347_y0, h_u_cla12_and346_y0, h_u_cla12_and348_y0);
  and_gate and_gate_h_u_cla12_and349_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and349_y0);
  and_gate and_gate_h_u_cla12_and350_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and350_y0);
  and_gate and_gate_h_u_cla12_and351_y0(h_u_cla12_and350_y0, h_u_cla12_and349_y0, h_u_cla12_and351_y0);
  and_gate and_gate_h_u_cla12_and352_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and352_y0);
  and_gate and_gate_h_u_cla12_and353_y0(h_u_cla12_and352_y0, h_u_cla12_and351_y0, h_u_cla12_and353_y0);
  and_gate and_gate_h_u_cla12_and354_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and354_y0);
  and_gate and_gate_h_u_cla12_and355_y0(h_u_cla12_and354_y0, h_u_cla12_and353_y0, h_u_cla12_and355_y0);
  and_gate and_gate_h_u_cla12_and356_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and356_y0);
  and_gate and_gate_h_u_cla12_and357_y0(h_u_cla12_and356_y0, h_u_cla12_and355_y0, h_u_cla12_and357_y0);
  and_gate and_gate_h_u_cla12_and358_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and358_y0);
  and_gate and_gate_h_u_cla12_and359_y0(h_u_cla12_and358_y0, h_u_cla12_and357_y0, h_u_cla12_and359_y0);
  and_gate and_gate_h_u_cla12_and360_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and360_y0);
  and_gate and_gate_h_u_cla12_and361_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and361_y0);
  and_gate and_gate_h_u_cla12_and362_y0(h_u_cla12_and361_y0, h_u_cla12_and360_y0, h_u_cla12_and362_y0);
  and_gate and_gate_h_u_cla12_and363_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and363_y0);
  and_gate and_gate_h_u_cla12_and364_y0(h_u_cla12_and363_y0, h_u_cla12_and362_y0, h_u_cla12_and364_y0);
  and_gate and_gate_h_u_cla12_and365_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and365_y0);
  and_gate and_gate_h_u_cla12_and366_y0(h_u_cla12_and365_y0, h_u_cla12_and364_y0, h_u_cla12_and366_y0);
  and_gate and_gate_h_u_cla12_and367_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and367_y0);
  and_gate and_gate_h_u_cla12_and368_y0(h_u_cla12_and367_y0, h_u_cla12_and366_y0, h_u_cla12_and368_y0);
  and_gate and_gate_h_u_cla12_and369_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and369_y0);
  and_gate and_gate_h_u_cla12_and370_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and370_y0);
  and_gate and_gate_h_u_cla12_and371_y0(h_u_cla12_and370_y0, h_u_cla12_and369_y0, h_u_cla12_and371_y0);
  and_gate and_gate_h_u_cla12_and372_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and372_y0);
  and_gate and_gate_h_u_cla12_and373_y0(h_u_cla12_and372_y0, h_u_cla12_and371_y0, h_u_cla12_and373_y0);
  and_gate and_gate_h_u_cla12_and374_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and374_y0);
  and_gate and_gate_h_u_cla12_and375_y0(h_u_cla12_and374_y0, h_u_cla12_and373_y0, h_u_cla12_and375_y0);
  and_gate and_gate_h_u_cla12_and376_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and376_y0);
  and_gate and_gate_h_u_cla12_and377_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and377_y0);
  and_gate and_gate_h_u_cla12_and378_y0(h_u_cla12_and377_y0, h_u_cla12_and376_y0, h_u_cla12_and378_y0);
  and_gate and_gate_h_u_cla12_and379_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and379_y0);
  and_gate and_gate_h_u_cla12_and380_y0(h_u_cla12_and379_y0, h_u_cla12_and378_y0, h_u_cla12_and380_y0);
  and_gate and_gate_h_u_cla12_and381_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and381_y0);
  and_gate and_gate_h_u_cla12_and382_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and382_y0);
  and_gate and_gate_h_u_cla12_and383_y0(h_u_cla12_and382_y0, h_u_cla12_and381_y0, h_u_cla12_and383_y0);
  and_gate and_gate_h_u_cla12_and384_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_and384_y0);
  or_gate or_gate_h_u_cla12_or45_y0(h_u_cla12_and384_y0, h_u_cla12_and303_y0, h_u_cla12_or45_y0);
  or_gate or_gate_h_u_cla12_or46_y0(h_u_cla12_or45_y0, h_u_cla12_and320_y0, h_u_cla12_or46_y0);
  or_gate or_gate_h_u_cla12_or47_y0(h_u_cla12_or46_y0, h_u_cla12_and335_y0, h_u_cla12_or47_y0);
  or_gate or_gate_h_u_cla12_or48_y0(h_u_cla12_or47_y0, h_u_cla12_and348_y0, h_u_cla12_or48_y0);
  or_gate or_gate_h_u_cla12_or49_y0(h_u_cla12_or48_y0, h_u_cla12_and359_y0, h_u_cla12_or49_y0);
  or_gate or_gate_h_u_cla12_or50_y0(h_u_cla12_or49_y0, h_u_cla12_and368_y0, h_u_cla12_or50_y0);
  or_gate or_gate_h_u_cla12_or51_y0(h_u_cla12_or50_y0, h_u_cla12_and375_y0, h_u_cla12_or51_y0);
  or_gate or_gate_h_u_cla12_or52_y0(h_u_cla12_or51_y0, h_u_cla12_and380_y0, h_u_cla12_or52_y0);
  or_gate or_gate_h_u_cla12_or53_y0(h_u_cla12_or52_y0, h_u_cla12_and383_y0, h_u_cla12_or53_y0);
  or_gate or_gate_h_u_cla12_or54_y0(h_u_cla12_pg_logic9_y1, h_u_cla12_or53_y0, h_u_cla12_or54_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic10_y0(a_10, b_10, h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic10_y1, h_u_cla12_pg_logic10_y2);
  xor_gate xor_gate_h_u_cla12_xor10_y0(h_u_cla12_pg_logic10_y2, h_u_cla12_or54_y0, h_u_cla12_xor10_y0);
  and_gate and_gate_h_u_cla12_and385_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and385_y0);
  and_gate and_gate_h_u_cla12_and386_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and386_y0);
  and_gate and_gate_h_u_cla12_and387_y0(h_u_cla12_and386_y0, h_u_cla12_and385_y0, h_u_cla12_and387_y0);
  and_gate and_gate_h_u_cla12_and388_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and388_y0);
  and_gate and_gate_h_u_cla12_and389_y0(h_u_cla12_and388_y0, h_u_cla12_and387_y0, h_u_cla12_and389_y0);
  and_gate and_gate_h_u_cla12_and390_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and390_y0);
  and_gate and_gate_h_u_cla12_and391_y0(h_u_cla12_and390_y0, h_u_cla12_and389_y0, h_u_cla12_and391_y0);
  and_gate and_gate_h_u_cla12_and392_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and392_y0);
  and_gate and_gate_h_u_cla12_and393_y0(h_u_cla12_and392_y0, h_u_cla12_and391_y0, h_u_cla12_and393_y0);
  and_gate and_gate_h_u_cla12_and394_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and394_y0);
  and_gate and_gate_h_u_cla12_and395_y0(h_u_cla12_and394_y0, h_u_cla12_and393_y0, h_u_cla12_and395_y0);
  and_gate and_gate_h_u_cla12_and396_y0(h_u_cla12_pg_logic6_y0, constant_wire_0, h_u_cla12_and396_y0);
  and_gate and_gate_h_u_cla12_and397_y0(h_u_cla12_and396_y0, h_u_cla12_and395_y0, h_u_cla12_and397_y0);
  and_gate and_gate_h_u_cla12_and398_y0(h_u_cla12_pg_logic7_y0, constant_wire_0, h_u_cla12_and398_y0);
  and_gate and_gate_h_u_cla12_and399_y0(h_u_cla12_and398_y0, h_u_cla12_and397_y0, h_u_cla12_and399_y0);
  and_gate and_gate_h_u_cla12_and400_y0(h_u_cla12_pg_logic8_y0, constant_wire_0, h_u_cla12_and400_y0);
  and_gate and_gate_h_u_cla12_and401_y0(h_u_cla12_and400_y0, h_u_cla12_and399_y0, h_u_cla12_and401_y0);
  and_gate and_gate_h_u_cla12_and402_y0(h_u_cla12_pg_logic9_y0, constant_wire_0, h_u_cla12_and402_y0);
  and_gate and_gate_h_u_cla12_and403_y0(h_u_cla12_and402_y0, h_u_cla12_and401_y0, h_u_cla12_and403_y0);
  and_gate and_gate_h_u_cla12_and404_y0(h_u_cla12_pg_logic10_y0, constant_wire_0, h_u_cla12_and404_y0);
  and_gate and_gate_h_u_cla12_and405_y0(h_u_cla12_and404_y0, h_u_cla12_and403_y0, h_u_cla12_and405_y0);
  and_gate and_gate_h_u_cla12_and406_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and406_y0);
  and_gate and_gate_h_u_cla12_and407_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and407_y0);
  and_gate and_gate_h_u_cla12_and408_y0(h_u_cla12_and407_y0, h_u_cla12_and406_y0, h_u_cla12_and408_y0);
  and_gate and_gate_h_u_cla12_and409_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and409_y0);
  and_gate and_gate_h_u_cla12_and410_y0(h_u_cla12_and409_y0, h_u_cla12_and408_y0, h_u_cla12_and410_y0);
  and_gate and_gate_h_u_cla12_and411_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and411_y0);
  and_gate and_gate_h_u_cla12_and412_y0(h_u_cla12_and411_y0, h_u_cla12_and410_y0, h_u_cla12_and412_y0);
  and_gate and_gate_h_u_cla12_and413_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and413_y0);
  and_gate and_gate_h_u_cla12_and414_y0(h_u_cla12_and413_y0, h_u_cla12_and412_y0, h_u_cla12_and414_y0);
  and_gate and_gate_h_u_cla12_and415_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and415_y0);
  and_gate and_gate_h_u_cla12_and416_y0(h_u_cla12_and415_y0, h_u_cla12_and414_y0, h_u_cla12_and416_y0);
  and_gate and_gate_h_u_cla12_and417_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and417_y0);
  and_gate and_gate_h_u_cla12_and418_y0(h_u_cla12_and417_y0, h_u_cla12_and416_y0, h_u_cla12_and418_y0);
  and_gate and_gate_h_u_cla12_and419_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and419_y0);
  and_gate and_gate_h_u_cla12_and420_y0(h_u_cla12_and419_y0, h_u_cla12_and418_y0, h_u_cla12_and420_y0);
  and_gate and_gate_h_u_cla12_and421_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and421_y0);
  and_gate and_gate_h_u_cla12_and422_y0(h_u_cla12_and421_y0, h_u_cla12_and420_y0, h_u_cla12_and422_y0);
  and_gate and_gate_h_u_cla12_and423_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and423_y0);
  and_gate and_gate_h_u_cla12_and424_y0(h_u_cla12_and423_y0, h_u_cla12_and422_y0, h_u_cla12_and424_y0);
  and_gate and_gate_h_u_cla12_and425_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and425_y0);
  and_gate and_gate_h_u_cla12_and426_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and426_y0);
  and_gate and_gate_h_u_cla12_and427_y0(h_u_cla12_and426_y0, h_u_cla12_and425_y0, h_u_cla12_and427_y0);
  and_gate and_gate_h_u_cla12_and428_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and428_y0);
  and_gate and_gate_h_u_cla12_and429_y0(h_u_cla12_and428_y0, h_u_cla12_and427_y0, h_u_cla12_and429_y0);
  and_gate and_gate_h_u_cla12_and430_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and430_y0);
  and_gate and_gate_h_u_cla12_and431_y0(h_u_cla12_and430_y0, h_u_cla12_and429_y0, h_u_cla12_and431_y0);
  and_gate and_gate_h_u_cla12_and432_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and432_y0);
  and_gate and_gate_h_u_cla12_and433_y0(h_u_cla12_and432_y0, h_u_cla12_and431_y0, h_u_cla12_and433_y0);
  and_gate and_gate_h_u_cla12_and434_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and434_y0);
  and_gate and_gate_h_u_cla12_and435_y0(h_u_cla12_and434_y0, h_u_cla12_and433_y0, h_u_cla12_and435_y0);
  and_gate and_gate_h_u_cla12_and436_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and436_y0);
  and_gate and_gate_h_u_cla12_and437_y0(h_u_cla12_and436_y0, h_u_cla12_and435_y0, h_u_cla12_and437_y0);
  and_gate and_gate_h_u_cla12_and438_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and438_y0);
  and_gate and_gate_h_u_cla12_and439_y0(h_u_cla12_and438_y0, h_u_cla12_and437_y0, h_u_cla12_and439_y0);
  and_gate and_gate_h_u_cla12_and440_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and440_y0);
  and_gate and_gate_h_u_cla12_and441_y0(h_u_cla12_and440_y0, h_u_cla12_and439_y0, h_u_cla12_and441_y0);
  and_gate and_gate_h_u_cla12_and442_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and442_y0);
  and_gate and_gate_h_u_cla12_and443_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and443_y0);
  and_gate and_gate_h_u_cla12_and444_y0(h_u_cla12_and443_y0, h_u_cla12_and442_y0, h_u_cla12_and444_y0);
  and_gate and_gate_h_u_cla12_and445_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and445_y0);
  and_gate and_gate_h_u_cla12_and446_y0(h_u_cla12_and445_y0, h_u_cla12_and444_y0, h_u_cla12_and446_y0);
  and_gate and_gate_h_u_cla12_and447_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and447_y0);
  and_gate and_gate_h_u_cla12_and448_y0(h_u_cla12_and447_y0, h_u_cla12_and446_y0, h_u_cla12_and448_y0);
  and_gate and_gate_h_u_cla12_and449_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and449_y0);
  and_gate and_gate_h_u_cla12_and450_y0(h_u_cla12_and449_y0, h_u_cla12_and448_y0, h_u_cla12_and450_y0);
  and_gate and_gate_h_u_cla12_and451_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and451_y0);
  and_gate and_gate_h_u_cla12_and452_y0(h_u_cla12_and451_y0, h_u_cla12_and450_y0, h_u_cla12_and452_y0);
  and_gate and_gate_h_u_cla12_and453_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and453_y0);
  and_gate and_gate_h_u_cla12_and454_y0(h_u_cla12_and453_y0, h_u_cla12_and452_y0, h_u_cla12_and454_y0);
  and_gate and_gate_h_u_cla12_and455_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and455_y0);
  and_gate and_gate_h_u_cla12_and456_y0(h_u_cla12_and455_y0, h_u_cla12_and454_y0, h_u_cla12_and456_y0);
  and_gate and_gate_h_u_cla12_and457_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and457_y0);
  and_gate and_gate_h_u_cla12_and458_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and458_y0);
  and_gate and_gate_h_u_cla12_and459_y0(h_u_cla12_and458_y0, h_u_cla12_and457_y0, h_u_cla12_and459_y0);
  and_gate and_gate_h_u_cla12_and460_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and460_y0);
  and_gate and_gate_h_u_cla12_and461_y0(h_u_cla12_and460_y0, h_u_cla12_and459_y0, h_u_cla12_and461_y0);
  and_gate and_gate_h_u_cla12_and462_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and462_y0);
  and_gate and_gate_h_u_cla12_and463_y0(h_u_cla12_and462_y0, h_u_cla12_and461_y0, h_u_cla12_and463_y0);
  and_gate and_gate_h_u_cla12_and464_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and464_y0);
  and_gate and_gate_h_u_cla12_and465_y0(h_u_cla12_and464_y0, h_u_cla12_and463_y0, h_u_cla12_and465_y0);
  and_gate and_gate_h_u_cla12_and466_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and466_y0);
  and_gate and_gate_h_u_cla12_and467_y0(h_u_cla12_and466_y0, h_u_cla12_and465_y0, h_u_cla12_and467_y0);
  and_gate and_gate_h_u_cla12_and468_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and468_y0);
  and_gate and_gate_h_u_cla12_and469_y0(h_u_cla12_and468_y0, h_u_cla12_and467_y0, h_u_cla12_and469_y0);
  and_gate and_gate_h_u_cla12_and470_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and470_y0);
  and_gate and_gate_h_u_cla12_and471_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and471_y0);
  and_gate and_gate_h_u_cla12_and472_y0(h_u_cla12_and471_y0, h_u_cla12_and470_y0, h_u_cla12_and472_y0);
  and_gate and_gate_h_u_cla12_and473_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and473_y0);
  and_gate and_gate_h_u_cla12_and474_y0(h_u_cla12_and473_y0, h_u_cla12_and472_y0, h_u_cla12_and474_y0);
  and_gate and_gate_h_u_cla12_and475_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and475_y0);
  and_gate and_gate_h_u_cla12_and476_y0(h_u_cla12_and475_y0, h_u_cla12_and474_y0, h_u_cla12_and476_y0);
  and_gate and_gate_h_u_cla12_and477_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and477_y0);
  and_gate and_gate_h_u_cla12_and478_y0(h_u_cla12_and477_y0, h_u_cla12_and476_y0, h_u_cla12_and478_y0);
  and_gate and_gate_h_u_cla12_and479_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and479_y0);
  and_gate and_gate_h_u_cla12_and480_y0(h_u_cla12_and479_y0, h_u_cla12_and478_y0, h_u_cla12_and480_y0);
  and_gate and_gate_h_u_cla12_and481_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and481_y0);
  and_gate and_gate_h_u_cla12_and482_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and482_y0);
  and_gate and_gate_h_u_cla12_and483_y0(h_u_cla12_and482_y0, h_u_cla12_and481_y0, h_u_cla12_and483_y0);
  and_gate and_gate_h_u_cla12_and484_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and484_y0);
  and_gate and_gate_h_u_cla12_and485_y0(h_u_cla12_and484_y0, h_u_cla12_and483_y0, h_u_cla12_and485_y0);
  and_gate and_gate_h_u_cla12_and486_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and486_y0);
  and_gate and_gate_h_u_cla12_and487_y0(h_u_cla12_and486_y0, h_u_cla12_and485_y0, h_u_cla12_and487_y0);
  and_gate and_gate_h_u_cla12_and488_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and488_y0);
  and_gate and_gate_h_u_cla12_and489_y0(h_u_cla12_and488_y0, h_u_cla12_and487_y0, h_u_cla12_and489_y0);
  and_gate and_gate_h_u_cla12_and490_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and490_y0);
  and_gate and_gate_h_u_cla12_and491_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and491_y0);
  and_gate and_gate_h_u_cla12_and492_y0(h_u_cla12_and491_y0, h_u_cla12_and490_y0, h_u_cla12_and492_y0);
  and_gate and_gate_h_u_cla12_and493_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and493_y0);
  and_gate and_gate_h_u_cla12_and494_y0(h_u_cla12_and493_y0, h_u_cla12_and492_y0, h_u_cla12_and494_y0);
  and_gate and_gate_h_u_cla12_and495_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and495_y0);
  and_gate and_gate_h_u_cla12_and496_y0(h_u_cla12_and495_y0, h_u_cla12_and494_y0, h_u_cla12_and496_y0);
  and_gate and_gate_h_u_cla12_and497_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and497_y0);
  and_gate and_gate_h_u_cla12_and498_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and498_y0);
  and_gate and_gate_h_u_cla12_and499_y0(h_u_cla12_and498_y0, h_u_cla12_and497_y0, h_u_cla12_and499_y0);
  and_gate and_gate_h_u_cla12_and500_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and500_y0);
  and_gate and_gate_h_u_cla12_and501_y0(h_u_cla12_and500_y0, h_u_cla12_and499_y0, h_u_cla12_and501_y0);
  and_gate and_gate_h_u_cla12_and502_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_and502_y0);
  and_gate and_gate_h_u_cla12_and503_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_and503_y0);
  and_gate and_gate_h_u_cla12_and504_y0(h_u_cla12_and503_y0, h_u_cla12_and502_y0, h_u_cla12_and504_y0);
  and_gate and_gate_h_u_cla12_and505_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic9_y1, h_u_cla12_and505_y0);
  or_gate or_gate_h_u_cla12_or55_y0(h_u_cla12_and505_y0, h_u_cla12_and405_y0, h_u_cla12_or55_y0);
  or_gate or_gate_h_u_cla12_or56_y0(h_u_cla12_or55_y0, h_u_cla12_and424_y0, h_u_cla12_or56_y0);
  or_gate or_gate_h_u_cla12_or57_y0(h_u_cla12_or56_y0, h_u_cla12_and441_y0, h_u_cla12_or57_y0);
  or_gate or_gate_h_u_cla12_or58_y0(h_u_cla12_or57_y0, h_u_cla12_and456_y0, h_u_cla12_or58_y0);
  or_gate or_gate_h_u_cla12_or59_y0(h_u_cla12_or58_y0, h_u_cla12_and469_y0, h_u_cla12_or59_y0);
  or_gate or_gate_h_u_cla12_or60_y0(h_u_cla12_or59_y0, h_u_cla12_and480_y0, h_u_cla12_or60_y0);
  or_gate or_gate_h_u_cla12_or61_y0(h_u_cla12_or60_y0, h_u_cla12_and489_y0, h_u_cla12_or61_y0);
  or_gate or_gate_h_u_cla12_or62_y0(h_u_cla12_or61_y0, h_u_cla12_and496_y0, h_u_cla12_or62_y0);
  or_gate or_gate_h_u_cla12_or63_y0(h_u_cla12_or62_y0, h_u_cla12_and501_y0, h_u_cla12_or63_y0);
  or_gate or_gate_h_u_cla12_or64_y0(h_u_cla12_or63_y0, h_u_cla12_and504_y0, h_u_cla12_or64_y0);
  or_gate or_gate_h_u_cla12_or65_y0(h_u_cla12_pg_logic10_y1, h_u_cla12_or64_y0, h_u_cla12_or65_y0);
  pg_logic pg_logic_h_u_cla12_pg_logic11_y0(a_11, b_11, h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic11_y1, h_u_cla12_pg_logic11_y2);
  xor_gate xor_gate_h_u_cla12_xor11_y0(h_u_cla12_pg_logic11_y2, h_u_cla12_or65_y0, h_u_cla12_xor11_y0);
  and_gate and_gate_h_u_cla12_and506_y0(h_u_cla12_pg_logic0_y0, constant_wire_0, h_u_cla12_and506_y0);
  and_gate and_gate_h_u_cla12_and507_y0(h_u_cla12_pg_logic1_y0, constant_wire_0, h_u_cla12_and507_y0);
  and_gate and_gate_h_u_cla12_and508_y0(h_u_cla12_and507_y0, h_u_cla12_and506_y0, h_u_cla12_and508_y0);
  and_gate and_gate_h_u_cla12_and509_y0(h_u_cla12_pg_logic2_y0, constant_wire_0, h_u_cla12_and509_y0);
  and_gate and_gate_h_u_cla12_and510_y0(h_u_cla12_and509_y0, h_u_cla12_and508_y0, h_u_cla12_and510_y0);
  and_gate and_gate_h_u_cla12_and511_y0(h_u_cla12_pg_logic3_y0, constant_wire_0, h_u_cla12_and511_y0);
  and_gate and_gate_h_u_cla12_and512_y0(h_u_cla12_and511_y0, h_u_cla12_and510_y0, h_u_cla12_and512_y0);
  and_gate and_gate_h_u_cla12_and513_y0(h_u_cla12_pg_logic4_y0, constant_wire_0, h_u_cla12_and513_y0);
  and_gate and_gate_h_u_cla12_and514_y0(h_u_cla12_and513_y0, h_u_cla12_and512_y0, h_u_cla12_and514_y0);
  and_gate and_gate_h_u_cla12_and515_y0(h_u_cla12_pg_logic5_y0, constant_wire_0, h_u_cla12_and515_y0);
  and_gate and_gate_h_u_cla12_and516_y0(h_u_cla12_and515_y0, h_u_cla12_and514_y0, h_u_cla12_and516_y0);
  and_gate and_gate_h_u_cla12_and517_y0(h_u_cla12_pg_logic6_y0, constant_wire_0, h_u_cla12_and517_y0);
  and_gate and_gate_h_u_cla12_and518_y0(h_u_cla12_and517_y0, h_u_cla12_and516_y0, h_u_cla12_and518_y0);
  and_gate and_gate_h_u_cla12_and519_y0(h_u_cla12_pg_logic7_y0, constant_wire_0, h_u_cla12_and519_y0);
  and_gate and_gate_h_u_cla12_and520_y0(h_u_cla12_and519_y0, h_u_cla12_and518_y0, h_u_cla12_and520_y0);
  and_gate and_gate_h_u_cla12_and521_y0(h_u_cla12_pg_logic8_y0, constant_wire_0, h_u_cla12_and521_y0);
  and_gate and_gate_h_u_cla12_and522_y0(h_u_cla12_and521_y0, h_u_cla12_and520_y0, h_u_cla12_and522_y0);
  and_gate and_gate_h_u_cla12_and523_y0(h_u_cla12_pg_logic9_y0, constant_wire_0, h_u_cla12_and523_y0);
  and_gate and_gate_h_u_cla12_and524_y0(h_u_cla12_and523_y0, h_u_cla12_and522_y0, h_u_cla12_and524_y0);
  and_gate and_gate_h_u_cla12_and525_y0(h_u_cla12_pg_logic10_y0, constant_wire_0, h_u_cla12_and525_y0);
  and_gate and_gate_h_u_cla12_and526_y0(h_u_cla12_and525_y0, h_u_cla12_and524_y0, h_u_cla12_and526_y0);
  and_gate and_gate_h_u_cla12_and527_y0(h_u_cla12_pg_logic11_y0, constant_wire_0, h_u_cla12_and527_y0);
  and_gate and_gate_h_u_cla12_and528_y0(h_u_cla12_and527_y0, h_u_cla12_and526_y0, h_u_cla12_and528_y0);
  and_gate and_gate_h_u_cla12_and529_y0(h_u_cla12_pg_logic1_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and529_y0);
  and_gate and_gate_h_u_cla12_and530_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and530_y0);
  and_gate and_gate_h_u_cla12_and531_y0(h_u_cla12_and530_y0, h_u_cla12_and529_y0, h_u_cla12_and531_y0);
  and_gate and_gate_h_u_cla12_and532_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and532_y0);
  and_gate and_gate_h_u_cla12_and533_y0(h_u_cla12_and532_y0, h_u_cla12_and531_y0, h_u_cla12_and533_y0);
  and_gate and_gate_h_u_cla12_and534_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and534_y0);
  and_gate and_gate_h_u_cla12_and535_y0(h_u_cla12_and534_y0, h_u_cla12_and533_y0, h_u_cla12_and535_y0);
  and_gate and_gate_h_u_cla12_and536_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and536_y0);
  and_gate and_gate_h_u_cla12_and537_y0(h_u_cla12_and536_y0, h_u_cla12_and535_y0, h_u_cla12_and537_y0);
  and_gate and_gate_h_u_cla12_and538_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and538_y0);
  and_gate and_gate_h_u_cla12_and539_y0(h_u_cla12_and538_y0, h_u_cla12_and537_y0, h_u_cla12_and539_y0);
  and_gate and_gate_h_u_cla12_and540_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and540_y0);
  and_gate and_gate_h_u_cla12_and541_y0(h_u_cla12_and540_y0, h_u_cla12_and539_y0, h_u_cla12_and541_y0);
  and_gate and_gate_h_u_cla12_and542_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and542_y0);
  and_gate and_gate_h_u_cla12_and543_y0(h_u_cla12_and542_y0, h_u_cla12_and541_y0, h_u_cla12_and543_y0);
  and_gate and_gate_h_u_cla12_and544_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and544_y0);
  and_gate and_gate_h_u_cla12_and545_y0(h_u_cla12_and544_y0, h_u_cla12_and543_y0, h_u_cla12_and545_y0);
  and_gate and_gate_h_u_cla12_and546_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and546_y0);
  and_gate and_gate_h_u_cla12_and547_y0(h_u_cla12_and546_y0, h_u_cla12_and545_y0, h_u_cla12_and547_y0);
  and_gate and_gate_h_u_cla12_and548_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic0_y1, h_u_cla12_and548_y0);
  and_gate and_gate_h_u_cla12_and549_y0(h_u_cla12_and548_y0, h_u_cla12_and547_y0, h_u_cla12_and549_y0);
  and_gate and_gate_h_u_cla12_and550_y0(h_u_cla12_pg_logic2_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and550_y0);
  and_gate and_gate_h_u_cla12_and551_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and551_y0);
  and_gate and_gate_h_u_cla12_and552_y0(h_u_cla12_and551_y0, h_u_cla12_and550_y0, h_u_cla12_and552_y0);
  and_gate and_gate_h_u_cla12_and553_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and553_y0);
  and_gate and_gate_h_u_cla12_and554_y0(h_u_cla12_and553_y0, h_u_cla12_and552_y0, h_u_cla12_and554_y0);
  and_gate and_gate_h_u_cla12_and555_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and555_y0);
  and_gate and_gate_h_u_cla12_and556_y0(h_u_cla12_and555_y0, h_u_cla12_and554_y0, h_u_cla12_and556_y0);
  and_gate and_gate_h_u_cla12_and557_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and557_y0);
  and_gate and_gate_h_u_cla12_and558_y0(h_u_cla12_and557_y0, h_u_cla12_and556_y0, h_u_cla12_and558_y0);
  and_gate and_gate_h_u_cla12_and559_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and559_y0);
  and_gate and_gate_h_u_cla12_and560_y0(h_u_cla12_and559_y0, h_u_cla12_and558_y0, h_u_cla12_and560_y0);
  and_gate and_gate_h_u_cla12_and561_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and561_y0);
  and_gate and_gate_h_u_cla12_and562_y0(h_u_cla12_and561_y0, h_u_cla12_and560_y0, h_u_cla12_and562_y0);
  and_gate and_gate_h_u_cla12_and563_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and563_y0);
  and_gate and_gate_h_u_cla12_and564_y0(h_u_cla12_and563_y0, h_u_cla12_and562_y0, h_u_cla12_and564_y0);
  and_gate and_gate_h_u_cla12_and565_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and565_y0);
  and_gate and_gate_h_u_cla12_and566_y0(h_u_cla12_and565_y0, h_u_cla12_and564_y0, h_u_cla12_and566_y0);
  and_gate and_gate_h_u_cla12_and567_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic1_y1, h_u_cla12_and567_y0);
  and_gate and_gate_h_u_cla12_and568_y0(h_u_cla12_and567_y0, h_u_cla12_and566_y0, h_u_cla12_and568_y0);
  and_gate and_gate_h_u_cla12_and569_y0(h_u_cla12_pg_logic3_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and569_y0);
  and_gate and_gate_h_u_cla12_and570_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and570_y0);
  and_gate and_gate_h_u_cla12_and571_y0(h_u_cla12_and570_y0, h_u_cla12_and569_y0, h_u_cla12_and571_y0);
  and_gate and_gate_h_u_cla12_and572_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and572_y0);
  and_gate and_gate_h_u_cla12_and573_y0(h_u_cla12_and572_y0, h_u_cla12_and571_y0, h_u_cla12_and573_y0);
  and_gate and_gate_h_u_cla12_and574_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and574_y0);
  and_gate and_gate_h_u_cla12_and575_y0(h_u_cla12_and574_y0, h_u_cla12_and573_y0, h_u_cla12_and575_y0);
  and_gate and_gate_h_u_cla12_and576_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and576_y0);
  and_gate and_gate_h_u_cla12_and577_y0(h_u_cla12_and576_y0, h_u_cla12_and575_y0, h_u_cla12_and577_y0);
  and_gate and_gate_h_u_cla12_and578_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and578_y0);
  and_gate and_gate_h_u_cla12_and579_y0(h_u_cla12_and578_y0, h_u_cla12_and577_y0, h_u_cla12_and579_y0);
  and_gate and_gate_h_u_cla12_and580_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and580_y0);
  and_gate and_gate_h_u_cla12_and581_y0(h_u_cla12_and580_y0, h_u_cla12_and579_y0, h_u_cla12_and581_y0);
  and_gate and_gate_h_u_cla12_and582_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and582_y0);
  and_gate and_gate_h_u_cla12_and583_y0(h_u_cla12_and582_y0, h_u_cla12_and581_y0, h_u_cla12_and583_y0);
  and_gate and_gate_h_u_cla12_and584_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic2_y1, h_u_cla12_and584_y0);
  and_gate and_gate_h_u_cla12_and585_y0(h_u_cla12_and584_y0, h_u_cla12_and583_y0, h_u_cla12_and585_y0);
  and_gate and_gate_h_u_cla12_and586_y0(h_u_cla12_pg_logic4_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and586_y0);
  and_gate and_gate_h_u_cla12_and587_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and587_y0);
  and_gate and_gate_h_u_cla12_and588_y0(h_u_cla12_and587_y0, h_u_cla12_and586_y0, h_u_cla12_and588_y0);
  and_gate and_gate_h_u_cla12_and589_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and589_y0);
  and_gate and_gate_h_u_cla12_and590_y0(h_u_cla12_and589_y0, h_u_cla12_and588_y0, h_u_cla12_and590_y0);
  and_gate and_gate_h_u_cla12_and591_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and591_y0);
  and_gate and_gate_h_u_cla12_and592_y0(h_u_cla12_and591_y0, h_u_cla12_and590_y0, h_u_cla12_and592_y0);
  and_gate and_gate_h_u_cla12_and593_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and593_y0);
  and_gate and_gate_h_u_cla12_and594_y0(h_u_cla12_and593_y0, h_u_cla12_and592_y0, h_u_cla12_and594_y0);
  and_gate and_gate_h_u_cla12_and595_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and595_y0);
  and_gate and_gate_h_u_cla12_and596_y0(h_u_cla12_and595_y0, h_u_cla12_and594_y0, h_u_cla12_and596_y0);
  and_gate and_gate_h_u_cla12_and597_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and597_y0);
  and_gate and_gate_h_u_cla12_and598_y0(h_u_cla12_and597_y0, h_u_cla12_and596_y0, h_u_cla12_and598_y0);
  and_gate and_gate_h_u_cla12_and599_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic3_y1, h_u_cla12_and599_y0);
  and_gate and_gate_h_u_cla12_and600_y0(h_u_cla12_and599_y0, h_u_cla12_and598_y0, h_u_cla12_and600_y0);
  and_gate and_gate_h_u_cla12_and601_y0(h_u_cla12_pg_logic5_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and601_y0);
  and_gate and_gate_h_u_cla12_and602_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and602_y0);
  and_gate and_gate_h_u_cla12_and603_y0(h_u_cla12_and602_y0, h_u_cla12_and601_y0, h_u_cla12_and603_y0);
  and_gate and_gate_h_u_cla12_and604_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and604_y0);
  and_gate and_gate_h_u_cla12_and605_y0(h_u_cla12_and604_y0, h_u_cla12_and603_y0, h_u_cla12_and605_y0);
  and_gate and_gate_h_u_cla12_and606_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and606_y0);
  and_gate and_gate_h_u_cla12_and607_y0(h_u_cla12_and606_y0, h_u_cla12_and605_y0, h_u_cla12_and607_y0);
  and_gate and_gate_h_u_cla12_and608_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and608_y0);
  and_gate and_gate_h_u_cla12_and609_y0(h_u_cla12_and608_y0, h_u_cla12_and607_y0, h_u_cla12_and609_y0);
  and_gate and_gate_h_u_cla12_and610_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and610_y0);
  and_gate and_gate_h_u_cla12_and611_y0(h_u_cla12_and610_y0, h_u_cla12_and609_y0, h_u_cla12_and611_y0);
  and_gate and_gate_h_u_cla12_and612_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic4_y1, h_u_cla12_and612_y0);
  and_gate and_gate_h_u_cla12_and613_y0(h_u_cla12_and612_y0, h_u_cla12_and611_y0, h_u_cla12_and613_y0);
  and_gate and_gate_h_u_cla12_and614_y0(h_u_cla12_pg_logic6_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and614_y0);
  and_gate and_gate_h_u_cla12_and615_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and615_y0);
  and_gate and_gate_h_u_cla12_and616_y0(h_u_cla12_and615_y0, h_u_cla12_and614_y0, h_u_cla12_and616_y0);
  and_gate and_gate_h_u_cla12_and617_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and617_y0);
  and_gate and_gate_h_u_cla12_and618_y0(h_u_cla12_and617_y0, h_u_cla12_and616_y0, h_u_cla12_and618_y0);
  and_gate and_gate_h_u_cla12_and619_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and619_y0);
  and_gate and_gate_h_u_cla12_and620_y0(h_u_cla12_and619_y0, h_u_cla12_and618_y0, h_u_cla12_and620_y0);
  and_gate and_gate_h_u_cla12_and621_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and621_y0);
  and_gate and_gate_h_u_cla12_and622_y0(h_u_cla12_and621_y0, h_u_cla12_and620_y0, h_u_cla12_and622_y0);
  and_gate and_gate_h_u_cla12_and623_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic5_y1, h_u_cla12_and623_y0);
  and_gate and_gate_h_u_cla12_and624_y0(h_u_cla12_and623_y0, h_u_cla12_and622_y0, h_u_cla12_and624_y0);
  and_gate and_gate_h_u_cla12_and625_y0(h_u_cla12_pg_logic7_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and625_y0);
  and_gate and_gate_h_u_cla12_and626_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and626_y0);
  and_gate and_gate_h_u_cla12_and627_y0(h_u_cla12_and626_y0, h_u_cla12_and625_y0, h_u_cla12_and627_y0);
  and_gate and_gate_h_u_cla12_and628_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and628_y0);
  and_gate and_gate_h_u_cla12_and629_y0(h_u_cla12_and628_y0, h_u_cla12_and627_y0, h_u_cla12_and629_y0);
  and_gate and_gate_h_u_cla12_and630_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and630_y0);
  and_gate and_gate_h_u_cla12_and631_y0(h_u_cla12_and630_y0, h_u_cla12_and629_y0, h_u_cla12_and631_y0);
  and_gate and_gate_h_u_cla12_and632_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic6_y1, h_u_cla12_and632_y0);
  and_gate and_gate_h_u_cla12_and633_y0(h_u_cla12_and632_y0, h_u_cla12_and631_y0, h_u_cla12_and633_y0);
  and_gate and_gate_h_u_cla12_and634_y0(h_u_cla12_pg_logic8_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and634_y0);
  and_gate and_gate_h_u_cla12_and635_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and635_y0);
  and_gate and_gate_h_u_cla12_and636_y0(h_u_cla12_and635_y0, h_u_cla12_and634_y0, h_u_cla12_and636_y0);
  and_gate and_gate_h_u_cla12_and637_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and637_y0);
  and_gate and_gate_h_u_cla12_and638_y0(h_u_cla12_and637_y0, h_u_cla12_and636_y0, h_u_cla12_and638_y0);
  and_gate and_gate_h_u_cla12_and639_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic7_y1, h_u_cla12_and639_y0);
  and_gate and_gate_h_u_cla12_and640_y0(h_u_cla12_and639_y0, h_u_cla12_and638_y0, h_u_cla12_and640_y0);
  and_gate and_gate_h_u_cla12_and641_y0(h_u_cla12_pg_logic9_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_and641_y0);
  and_gate and_gate_h_u_cla12_and642_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_and642_y0);
  and_gate and_gate_h_u_cla12_and643_y0(h_u_cla12_and642_y0, h_u_cla12_and641_y0, h_u_cla12_and643_y0);
  and_gate and_gate_h_u_cla12_and644_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic8_y1, h_u_cla12_and644_y0);
  and_gate and_gate_h_u_cla12_and645_y0(h_u_cla12_and644_y0, h_u_cla12_and643_y0, h_u_cla12_and645_y0);
  and_gate and_gate_h_u_cla12_and646_y0(h_u_cla12_pg_logic10_y0, h_u_cla12_pg_logic9_y1, h_u_cla12_and646_y0);
  and_gate and_gate_h_u_cla12_and647_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic9_y1, h_u_cla12_and647_y0);
  and_gate and_gate_h_u_cla12_and648_y0(h_u_cla12_and647_y0, h_u_cla12_and646_y0, h_u_cla12_and648_y0);
  and_gate and_gate_h_u_cla12_and649_y0(h_u_cla12_pg_logic11_y0, h_u_cla12_pg_logic10_y1, h_u_cla12_and649_y0);
  or_gate or_gate_h_u_cla12_or66_y0(h_u_cla12_and649_y0, h_u_cla12_and528_y0, h_u_cla12_or66_y0);
  or_gate or_gate_h_u_cla12_or67_y0(h_u_cla12_or66_y0, h_u_cla12_and549_y0, h_u_cla12_or67_y0);
  or_gate or_gate_h_u_cla12_or68_y0(h_u_cla12_or67_y0, h_u_cla12_and568_y0, h_u_cla12_or68_y0);
  or_gate or_gate_h_u_cla12_or69_y0(h_u_cla12_or68_y0, h_u_cla12_and585_y0, h_u_cla12_or69_y0);
  or_gate or_gate_h_u_cla12_or70_y0(h_u_cla12_or69_y0, h_u_cla12_and600_y0, h_u_cla12_or70_y0);
  or_gate or_gate_h_u_cla12_or71_y0(h_u_cla12_or70_y0, h_u_cla12_and613_y0, h_u_cla12_or71_y0);
  or_gate or_gate_h_u_cla12_or72_y0(h_u_cla12_or71_y0, h_u_cla12_and624_y0, h_u_cla12_or72_y0);
  or_gate or_gate_h_u_cla12_or73_y0(h_u_cla12_or72_y0, h_u_cla12_and633_y0, h_u_cla12_or73_y0);
  or_gate or_gate_h_u_cla12_or74_y0(h_u_cla12_or73_y0, h_u_cla12_and640_y0, h_u_cla12_or74_y0);
  or_gate or_gate_h_u_cla12_or75_y0(h_u_cla12_or74_y0, h_u_cla12_and645_y0, h_u_cla12_or75_y0);
  or_gate or_gate_h_u_cla12_or76_y0(h_u_cla12_or75_y0, h_u_cla12_and648_y0, h_u_cla12_or76_y0);
  or_gate or_gate_h_u_cla12_or77_y0(h_u_cla12_pg_logic11_y1, h_u_cla12_or76_y0, h_u_cla12_or77_y0);

  assign out[0] = h_u_cla12_xor0_y0;
  assign out[1] = h_u_cla12_xor1_y0;
  assign out[2] = h_u_cla12_xor2_y0;
  assign out[3] = h_u_cla12_xor3_y0;
  assign out[4] = h_u_cla12_xor4_y0;
  assign out[5] = h_u_cla12_xor5_y0;
  assign out[6] = h_u_cla12_xor6_y0;
  assign out[7] = h_u_cla12_xor7_y0;
  assign out[8] = h_u_cla12_xor8_y0;
  assign out[9] = h_u_cla12_xor9_y0;
  assign out[10] = h_u_cla12_xor10_y0;
  assign out[11] = h_u_cla12_xor11_y0;
  assign out[12] = h_u_cla12_or77_y0;
endmodule