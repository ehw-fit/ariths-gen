module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module h_u_rca32(input [31:0] a, input [31:0] b, output [32:0] h_u_rca32_out);
  wire [0:0] h_u_rca32_ha_xor0;
  wire [0:0] h_u_rca32_ha_and0;
  wire [0:0] h_u_rca32_fa1_xor1;
  wire [0:0] h_u_rca32_fa1_or0;
  wire [0:0] h_u_rca32_fa2_xor1;
  wire [0:0] h_u_rca32_fa2_or0;
  wire [0:0] h_u_rca32_fa3_xor1;
  wire [0:0] h_u_rca32_fa3_or0;
  wire [0:0] h_u_rca32_fa4_xor1;
  wire [0:0] h_u_rca32_fa4_or0;
  wire [0:0] h_u_rca32_fa5_xor1;
  wire [0:0] h_u_rca32_fa5_or0;
  wire [0:0] h_u_rca32_fa6_xor1;
  wire [0:0] h_u_rca32_fa6_or0;
  wire [0:0] h_u_rca32_fa7_xor1;
  wire [0:0] h_u_rca32_fa7_or0;
  wire [0:0] h_u_rca32_fa8_xor1;
  wire [0:0] h_u_rca32_fa8_or0;
  wire [0:0] h_u_rca32_fa9_xor1;
  wire [0:0] h_u_rca32_fa9_or0;
  wire [0:0] h_u_rca32_fa10_xor1;
  wire [0:0] h_u_rca32_fa10_or0;
  wire [0:0] h_u_rca32_fa11_xor1;
  wire [0:0] h_u_rca32_fa11_or0;
  wire [0:0] h_u_rca32_fa12_xor1;
  wire [0:0] h_u_rca32_fa12_or0;
  wire [0:0] h_u_rca32_fa13_xor1;
  wire [0:0] h_u_rca32_fa13_or0;
  wire [0:0] h_u_rca32_fa14_xor1;
  wire [0:0] h_u_rca32_fa14_or0;
  wire [0:0] h_u_rca32_fa15_xor1;
  wire [0:0] h_u_rca32_fa15_or0;
  wire [0:0] h_u_rca32_fa16_xor1;
  wire [0:0] h_u_rca32_fa16_or0;
  wire [0:0] h_u_rca32_fa17_xor1;
  wire [0:0] h_u_rca32_fa17_or0;
  wire [0:0] h_u_rca32_fa18_xor1;
  wire [0:0] h_u_rca32_fa18_or0;
  wire [0:0] h_u_rca32_fa19_xor1;
  wire [0:0] h_u_rca32_fa19_or0;
  wire [0:0] h_u_rca32_fa20_xor1;
  wire [0:0] h_u_rca32_fa20_or0;
  wire [0:0] h_u_rca32_fa21_xor1;
  wire [0:0] h_u_rca32_fa21_or0;
  wire [0:0] h_u_rca32_fa22_xor1;
  wire [0:0] h_u_rca32_fa22_or0;
  wire [0:0] h_u_rca32_fa23_xor1;
  wire [0:0] h_u_rca32_fa23_or0;
  wire [0:0] h_u_rca32_fa24_xor1;
  wire [0:0] h_u_rca32_fa24_or0;
  wire [0:0] h_u_rca32_fa25_xor1;
  wire [0:0] h_u_rca32_fa25_or0;
  wire [0:0] h_u_rca32_fa26_xor1;
  wire [0:0] h_u_rca32_fa26_or0;
  wire [0:0] h_u_rca32_fa27_xor1;
  wire [0:0] h_u_rca32_fa27_or0;
  wire [0:0] h_u_rca32_fa28_xor1;
  wire [0:0] h_u_rca32_fa28_or0;
  wire [0:0] h_u_rca32_fa29_xor1;
  wire [0:0] h_u_rca32_fa29_or0;
  wire [0:0] h_u_rca32_fa30_xor1;
  wire [0:0] h_u_rca32_fa30_or0;
  wire [0:0] h_u_rca32_fa31_xor1;
  wire [0:0] h_u_rca32_fa31_or0;

  ha ha_h_u_rca32_ha_out(.a(a[0]), .b(b[0]), .ha_xor0(h_u_rca32_ha_xor0), .ha_and0(h_u_rca32_ha_and0));
  fa fa_h_u_rca32_fa1_out(.a(a[1]), .b(b[1]), .cin(h_u_rca32_ha_and0[0]), .fa_xor1(h_u_rca32_fa1_xor1), .fa_or0(h_u_rca32_fa1_or0));
  fa fa_h_u_rca32_fa2_out(.a(a[2]), .b(b[2]), .cin(h_u_rca32_fa1_or0[0]), .fa_xor1(h_u_rca32_fa2_xor1), .fa_or0(h_u_rca32_fa2_or0));
  fa fa_h_u_rca32_fa3_out(.a(a[3]), .b(b[3]), .cin(h_u_rca32_fa2_or0[0]), .fa_xor1(h_u_rca32_fa3_xor1), .fa_or0(h_u_rca32_fa3_or0));
  fa fa_h_u_rca32_fa4_out(.a(a[4]), .b(b[4]), .cin(h_u_rca32_fa3_or0[0]), .fa_xor1(h_u_rca32_fa4_xor1), .fa_or0(h_u_rca32_fa4_or0));
  fa fa_h_u_rca32_fa5_out(.a(a[5]), .b(b[5]), .cin(h_u_rca32_fa4_or0[0]), .fa_xor1(h_u_rca32_fa5_xor1), .fa_or0(h_u_rca32_fa5_or0));
  fa fa_h_u_rca32_fa6_out(.a(a[6]), .b(b[6]), .cin(h_u_rca32_fa5_or0[0]), .fa_xor1(h_u_rca32_fa6_xor1), .fa_or0(h_u_rca32_fa6_or0));
  fa fa_h_u_rca32_fa7_out(.a(a[7]), .b(b[7]), .cin(h_u_rca32_fa6_or0[0]), .fa_xor1(h_u_rca32_fa7_xor1), .fa_or0(h_u_rca32_fa7_or0));
  fa fa_h_u_rca32_fa8_out(.a(a[8]), .b(b[8]), .cin(h_u_rca32_fa7_or0[0]), .fa_xor1(h_u_rca32_fa8_xor1), .fa_or0(h_u_rca32_fa8_or0));
  fa fa_h_u_rca32_fa9_out(.a(a[9]), .b(b[9]), .cin(h_u_rca32_fa8_or0[0]), .fa_xor1(h_u_rca32_fa9_xor1), .fa_or0(h_u_rca32_fa9_or0));
  fa fa_h_u_rca32_fa10_out(.a(a[10]), .b(b[10]), .cin(h_u_rca32_fa9_or0[0]), .fa_xor1(h_u_rca32_fa10_xor1), .fa_or0(h_u_rca32_fa10_or0));
  fa fa_h_u_rca32_fa11_out(.a(a[11]), .b(b[11]), .cin(h_u_rca32_fa10_or0[0]), .fa_xor1(h_u_rca32_fa11_xor1), .fa_or0(h_u_rca32_fa11_or0));
  fa fa_h_u_rca32_fa12_out(.a(a[12]), .b(b[12]), .cin(h_u_rca32_fa11_or0[0]), .fa_xor1(h_u_rca32_fa12_xor1), .fa_or0(h_u_rca32_fa12_or0));
  fa fa_h_u_rca32_fa13_out(.a(a[13]), .b(b[13]), .cin(h_u_rca32_fa12_or0[0]), .fa_xor1(h_u_rca32_fa13_xor1), .fa_or0(h_u_rca32_fa13_or0));
  fa fa_h_u_rca32_fa14_out(.a(a[14]), .b(b[14]), .cin(h_u_rca32_fa13_or0[0]), .fa_xor1(h_u_rca32_fa14_xor1), .fa_or0(h_u_rca32_fa14_or0));
  fa fa_h_u_rca32_fa15_out(.a(a[15]), .b(b[15]), .cin(h_u_rca32_fa14_or0[0]), .fa_xor1(h_u_rca32_fa15_xor1), .fa_or0(h_u_rca32_fa15_or0));
  fa fa_h_u_rca32_fa16_out(.a(a[16]), .b(b[16]), .cin(h_u_rca32_fa15_or0[0]), .fa_xor1(h_u_rca32_fa16_xor1), .fa_or0(h_u_rca32_fa16_or0));
  fa fa_h_u_rca32_fa17_out(.a(a[17]), .b(b[17]), .cin(h_u_rca32_fa16_or0[0]), .fa_xor1(h_u_rca32_fa17_xor1), .fa_or0(h_u_rca32_fa17_or0));
  fa fa_h_u_rca32_fa18_out(.a(a[18]), .b(b[18]), .cin(h_u_rca32_fa17_or0[0]), .fa_xor1(h_u_rca32_fa18_xor1), .fa_or0(h_u_rca32_fa18_or0));
  fa fa_h_u_rca32_fa19_out(.a(a[19]), .b(b[19]), .cin(h_u_rca32_fa18_or0[0]), .fa_xor1(h_u_rca32_fa19_xor1), .fa_or0(h_u_rca32_fa19_or0));
  fa fa_h_u_rca32_fa20_out(.a(a[20]), .b(b[20]), .cin(h_u_rca32_fa19_or0[0]), .fa_xor1(h_u_rca32_fa20_xor1), .fa_or0(h_u_rca32_fa20_or0));
  fa fa_h_u_rca32_fa21_out(.a(a[21]), .b(b[21]), .cin(h_u_rca32_fa20_or0[0]), .fa_xor1(h_u_rca32_fa21_xor1), .fa_or0(h_u_rca32_fa21_or0));
  fa fa_h_u_rca32_fa22_out(.a(a[22]), .b(b[22]), .cin(h_u_rca32_fa21_or0[0]), .fa_xor1(h_u_rca32_fa22_xor1), .fa_or0(h_u_rca32_fa22_or0));
  fa fa_h_u_rca32_fa23_out(.a(a[23]), .b(b[23]), .cin(h_u_rca32_fa22_or0[0]), .fa_xor1(h_u_rca32_fa23_xor1), .fa_or0(h_u_rca32_fa23_or0));
  fa fa_h_u_rca32_fa24_out(.a(a[24]), .b(b[24]), .cin(h_u_rca32_fa23_or0[0]), .fa_xor1(h_u_rca32_fa24_xor1), .fa_or0(h_u_rca32_fa24_or0));
  fa fa_h_u_rca32_fa25_out(.a(a[25]), .b(b[25]), .cin(h_u_rca32_fa24_or0[0]), .fa_xor1(h_u_rca32_fa25_xor1), .fa_or0(h_u_rca32_fa25_or0));
  fa fa_h_u_rca32_fa26_out(.a(a[26]), .b(b[26]), .cin(h_u_rca32_fa25_or0[0]), .fa_xor1(h_u_rca32_fa26_xor1), .fa_or0(h_u_rca32_fa26_or0));
  fa fa_h_u_rca32_fa27_out(.a(a[27]), .b(b[27]), .cin(h_u_rca32_fa26_or0[0]), .fa_xor1(h_u_rca32_fa27_xor1), .fa_or0(h_u_rca32_fa27_or0));
  fa fa_h_u_rca32_fa28_out(.a(a[28]), .b(b[28]), .cin(h_u_rca32_fa27_or0[0]), .fa_xor1(h_u_rca32_fa28_xor1), .fa_or0(h_u_rca32_fa28_or0));
  fa fa_h_u_rca32_fa29_out(.a(a[29]), .b(b[29]), .cin(h_u_rca32_fa28_or0[0]), .fa_xor1(h_u_rca32_fa29_xor1), .fa_or0(h_u_rca32_fa29_or0));
  fa fa_h_u_rca32_fa30_out(.a(a[30]), .b(b[30]), .cin(h_u_rca32_fa29_or0[0]), .fa_xor1(h_u_rca32_fa30_xor1), .fa_or0(h_u_rca32_fa30_or0));
  fa fa_h_u_rca32_fa31_out(.a(a[31]), .b(b[31]), .cin(h_u_rca32_fa30_or0[0]), .fa_xor1(h_u_rca32_fa31_xor1), .fa_or0(h_u_rca32_fa31_or0));

  assign h_u_rca32_out[0] = h_u_rca32_ha_xor0[0];
  assign h_u_rca32_out[1] = h_u_rca32_fa1_xor1[0];
  assign h_u_rca32_out[2] = h_u_rca32_fa2_xor1[0];
  assign h_u_rca32_out[3] = h_u_rca32_fa3_xor1[0];
  assign h_u_rca32_out[4] = h_u_rca32_fa4_xor1[0];
  assign h_u_rca32_out[5] = h_u_rca32_fa5_xor1[0];
  assign h_u_rca32_out[6] = h_u_rca32_fa6_xor1[0];
  assign h_u_rca32_out[7] = h_u_rca32_fa7_xor1[0];
  assign h_u_rca32_out[8] = h_u_rca32_fa8_xor1[0];
  assign h_u_rca32_out[9] = h_u_rca32_fa9_xor1[0];
  assign h_u_rca32_out[10] = h_u_rca32_fa10_xor1[0];
  assign h_u_rca32_out[11] = h_u_rca32_fa11_xor1[0];
  assign h_u_rca32_out[12] = h_u_rca32_fa12_xor1[0];
  assign h_u_rca32_out[13] = h_u_rca32_fa13_xor1[0];
  assign h_u_rca32_out[14] = h_u_rca32_fa14_xor1[0];
  assign h_u_rca32_out[15] = h_u_rca32_fa15_xor1[0];
  assign h_u_rca32_out[16] = h_u_rca32_fa16_xor1[0];
  assign h_u_rca32_out[17] = h_u_rca32_fa17_xor1[0];
  assign h_u_rca32_out[18] = h_u_rca32_fa18_xor1[0];
  assign h_u_rca32_out[19] = h_u_rca32_fa19_xor1[0];
  assign h_u_rca32_out[20] = h_u_rca32_fa20_xor1[0];
  assign h_u_rca32_out[21] = h_u_rca32_fa21_xor1[0];
  assign h_u_rca32_out[22] = h_u_rca32_fa22_xor1[0];
  assign h_u_rca32_out[23] = h_u_rca32_fa23_xor1[0];
  assign h_u_rca32_out[24] = h_u_rca32_fa24_xor1[0];
  assign h_u_rca32_out[25] = h_u_rca32_fa25_xor1[0];
  assign h_u_rca32_out[26] = h_u_rca32_fa26_xor1[0];
  assign h_u_rca32_out[27] = h_u_rca32_fa27_xor1[0];
  assign h_u_rca32_out[28] = h_u_rca32_fa28_xor1[0];
  assign h_u_rca32_out[29] = h_u_rca32_fa29_xor1[0];
  assign h_u_rca32_out[30] = h_u_rca32_fa30_xor1[0];
  assign h_u_rca32_out[31] = h_u_rca32_fa31_xor1[0];
  assign h_u_rca32_out[32] = h_u_rca32_fa31_or0[0];
endmodule