module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_cin;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module h_s_arrmul16(input [15:0] a, input [15:0] b, output [31:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire constant_wire_1;
  wire h_s_arrmul16_and0_0_y0;
  wire h_s_arrmul16_and1_0_y0;
  wire h_s_arrmul16_and2_0_y0;
  wire h_s_arrmul16_and3_0_y0;
  wire h_s_arrmul16_and4_0_y0;
  wire h_s_arrmul16_and5_0_y0;
  wire h_s_arrmul16_and6_0_y0;
  wire h_s_arrmul16_and7_0_y0;
  wire h_s_arrmul16_and8_0_y0;
  wire h_s_arrmul16_and9_0_y0;
  wire h_s_arrmul16_and10_0_y0;
  wire h_s_arrmul16_and11_0_y0;
  wire h_s_arrmul16_and12_0_y0;
  wire h_s_arrmul16_and13_0_y0;
  wire h_s_arrmul16_and14_0_y0;
  wire h_s_arrmul16_nand15_0_y0;
  wire h_s_arrmul16_and0_1_y0;
  wire h_s_arrmul16_ha0_1_y0;
  wire h_s_arrmul16_ha0_1_y1;
  wire h_s_arrmul16_and1_1_y0;
  wire h_s_arrmul16_fa1_1_y2;
  wire h_s_arrmul16_fa1_1_y4;
  wire h_s_arrmul16_and2_1_y0;
  wire h_s_arrmul16_fa2_1_y2;
  wire h_s_arrmul16_fa2_1_y4;
  wire h_s_arrmul16_and3_1_y0;
  wire h_s_arrmul16_fa3_1_y2;
  wire h_s_arrmul16_fa3_1_y4;
  wire h_s_arrmul16_and4_1_y0;
  wire h_s_arrmul16_fa4_1_y2;
  wire h_s_arrmul16_fa4_1_y4;
  wire h_s_arrmul16_and5_1_y0;
  wire h_s_arrmul16_fa5_1_y2;
  wire h_s_arrmul16_fa5_1_y4;
  wire h_s_arrmul16_and6_1_y0;
  wire h_s_arrmul16_fa6_1_y2;
  wire h_s_arrmul16_fa6_1_y4;
  wire h_s_arrmul16_and7_1_y0;
  wire h_s_arrmul16_fa7_1_y2;
  wire h_s_arrmul16_fa7_1_y4;
  wire h_s_arrmul16_and8_1_y0;
  wire h_s_arrmul16_fa8_1_y2;
  wire h_s_arrmul16_fa8_1_y4;
  wire h_s_arrmul16_and9_1_y0;
  wire h_s_arrmul16_fa9_1_y2;
  wire h_s_arrmul16_fa9_1_y4;
  wire h_s_arrmul16_and10_1_y0;
  wire h_s_arrmul16_fa10_1_y2;
  wire h_s_arrmul16_fa10_1_y4;
  wire h_s_arrmul16_and11_1_y0;
  wire h_s_arrmul16_fa11_1_y2;
  wire h_s_arrmul16_fa11_1_y4;
  wire h_s_arrmul16_and12_1_y0;
  wire h_s_arrmul16_fa12_1_y2;
  wire h_s_arrmul16_fa12_1_y4;
  wire h_s_arrmul16_and13_1_y0;
  wire h_s_arrmul16_fa13_1_y2;
  wire h_s_arrmul16_fa13_1_y4;
  wire h_s_arrmul16_and14_1_y0;
  wire h_s_arrmul16_fa14_1_y2;
  wire h_s_arrmul16_fa14_1_y4;
  wire h_s_arrmul16_nand15_1_y0;
  wire h_s_arrmul16_fa15_1_y2;
  wire h_s_arrmul16_fa15_1_y4;
  wire h_s_arrmul16_and0_2_y0;
  wire h_s_arrmul16_ha0_2_y0;
  wire h_s_arrmul16_ha0_2_y1;
  wire h_s_arrmul16_and1_2_y0;
  wire h_s_arrmul16_fa1_2_y2;
  wire h_s_arrmul16_fa1_2_y4;
  wire h_s_arrmul16_and2_2_y0;
  wire h_s_arrmul16_fa2_2_y2;
  wire h_s_arrmul16_fa2_2_y4;
  wire h_s_arrmul16_and3_2_y0;
  wire h_s_arrmul16_fa3_2_y2;
  wire h_s_arrmul16_fa3_2_y4;
  wire h_s_arrmul16_and4_2_y0;
  wire h_s_arrmul16_fa4_2_y2;
  wire h_s_arrmul16_fa4_2_y4;
  wire h_s_arrmul16_and5_2_y0;
  wire h_s_arrmul16_fa5_2_y2;
  wire h_s_arrmul16_fa5_2_y4;
  wire h_s_arrmul16_and6_2_y0;
  wire h_s_arrmul16_fa6_2_y2;
  wire h_s_arrmul16_fa6_2_y4;
  wire h_s_arrmul16_and7_2_y0;
  wire h_s_arrmul16_fa7_2_y2;
  wire h_s_arrmul16_fa7_2_y4;
  wire h_s_arrmul16_and8_2_y0;
  wire h_s_arrmul16_fa8_2_y2;
  wire h_s_arrmul16_fa8_2_y4;
  wire h_s_arrmul16_and9_2_y0;
  wire h_s_arrmul16_fa9_2_y2;
  wire h_s_arrmul16_fa9_2_y4;
  wire h_s_arrmul16_and10_2_y0;
  wire h_s_arrmul16_fa10_2_y2;
  wire h_s_arrmul16_fa10_2_y4;
  wire h_s_arrmul16_and11_2_y0;
  wire h_s_arrmul16_fa11_2_y2;
  wire h_s_arrmul16_fa11_2_y4;
  wire h_s_arrmul16_and12_2_y0;
  wire h_s_arrmul16_fa12_2_y2;
  wire h_s_arrmul16_fa12_2_y4;
  wire h_s_arrmul16_and13_2_y0;
  wire h_s_arrmul16_fa13_2_y2;
  wire h_s_arrmul16_fa13_2_y4;
  wire h_s_arrmul16_and14_2_y0;
  wire h_s_arrmul16_fa14_2_y2;
  wire h_s_arrmul16_fa14_2_y4;
  wire h_s_arrmul16_nand15_2_y0;
  wire h_s_arrmul16_fa15_2_y2;
  wire h_s_arrmul16_fa15_2_y4;
  wire h_s_arrmul16_and0_3_y0;
  wire h_s_arrmul16_ha0_3_y0;
  wire h_s_arrmul16_ha0_3_y1;
  wire h_s_arrmul16_and1_3_y0;
  wire h_s_arrmul16_fa1_3_y2;
  wire h_s_arrmul16_fa1_3_y4;
  wire h_s_arrmul16_and2_3_y0;
  wire h_s_arrmul16_fa2_3_y2;
  wire h_s_arrmul16_fa2_3_y4;
  wire h_s_arrmul16_and3_3_y0;
  wire h_s_arrmul16_fa3_3_y2;
  wire h_s_arrmul16_fa3_3_y4;
  wire h_s_arrmul16_and4_3_y0;
  wire h_s_arrmul16_fa4_3_y2;
  wire h_s_arrmul16_fa4_3_y4;
  wire h_s_arrmul16_and5_3_y0;
  wire h_s_arrmul16_fa5_3_y2;
  wire h_s_arrmul16_fa5_3_y4;
  wire h_s_arrmul16_and6_3_y0;
  wire h_s_arrmul16_fa6_3_y2;
  wire h_s_arrmul16_fa6_3_y4;
  wire h_s_arrmul16_and7_3_y0;
  wire h_s_arrmul16_fa7_3_y2;
  wire h_s_arrmul16_fa7_3_y4;
  wire h_s_arrmul16_and8_3_y0;
  wire h_s_arrmul16_fa8_3_y2;
  wire h_s_arrmul16_fa8_3_y4;
  wire h_s_arrmul16_and9_3_y0;
  wire h_s_arrmul16_fa9_3_y2;
  wire h_s_arrmul16_fa9_3_y4;
  wire h_s_arrmul16_and10_3_y0;
  wire h_s_arrmul16_fa10_3_y2;
  wire h_s_arrmul16_fa10_3_y4;
  wire h_s_arrmul16_and11_3_y0;
  wire h_s_arrmul16_fa11_3_y2;
  wire h_s_arrmul16_fa11_3_y4;
  wire h_s_arrmul16_and12_3_y0;
  wire h_s_arrmul16_fa12_3_y2;
  wire h_s_arrmul16_fa12_3_y4;
  wire h_s_arrmul16_and13_3_y0;
  wire h_s_arrmul16_fa13_3_y2;
  wire h_s_arrmul16_fa13_3_y4;
  wire h_s_arrmul16_and14_3_y0;
  wire h_s_arrmul16_fa14_3_y2;
  wire h_s_arrmul16_fa14_3_y4;
  wire h_s_arrmul16_nand15_3_y0;
  wire h_s_arrmul16_fa15_3_y2;
  wire h_s_arrmul16_fa15_3_y4;
  wire h_s_arrmul16_and0_4_y0;
  wire h_s_arrmul16_ha0_4_y0;
  wire h_s_arrmul16_ha0_4_y1;
  wire h_s_arrmul16_and1_4_y0;
  wire h_s_arrmul16_fa1_4_y2;
  wire h_s_arrmul16_fa1_4_y4;
  wire h_s_arrmul16_and2_4_y0;
  wire h_s_arrmul16_fa2_4_y2;
  wire h_s_arrmul16_fa2_4_y4;
  wire h_s_arrmul16_and3_4_y0;
  wire h_s_arrmul16_fa3_4_y2;
  wire h_s_arrmul16_fa3_4_y4;
  wire h_s_arrmul16_and4_4_y0;
  wire h_s_arrmul16_fa4_4_y2;
  wire h_s_arrmul16_fa4_4_y4;
  wire h_s_arrmul16_and5_4_y0;
  wire h_s_arrmul16_fa5_4_y2;
  wire h_s_arrmul16_fa5_4_y4;
  wire h_s_arrmul16_and6_4_y0;
  wire h_s_arrmul16_fa6_4_y2;
  wire h_s_arrmul16_fa6_4_y4;
  wire h_s_arrmul16_and7_4_y0;
  wire h_s_arrmul16_fa7_4_y2;
  wire h_s_arrmul16_fa7_4_y4;
  wire h_s_arrmul16_and8_4_y0;
  wire h_s_arrmul16_fa8_4_y2;
  wire h_s_arrmul16_fa8_4_y4;
  wire h_s_arrmul16_and9_4_y0;
  wire h_s_arrmul16_fa9_4_y2;
  wire h_s_arrmul16_fa9_4_y4;
  wire h_s_arrmul16_and10_4_y0;
  wire h_s_arrmul16_fa10_4_y2;
  wire h_s_arrmul16_fa10_4_y4;
  wire h_s_arrmul16_and11_4_y0;
  wire h_s_arrmul16_fa11_4_y2;
  wire h_s_arrmul16_fa11_4_y4;
  wire h_s_arrmul16_and12_4_y0;
  wire h_s_arrmul16_fa12_4_y2;
  wire h_s_arrmul16_fa12_4_y4;
  wire h_s_arrmul16_and13_4_y0;
  wire h_s_arrmul16_fa13_4_y2;
  wire h_s_arrmul16_fa13_4_y4;
  wire h_s_arrmul16_and14_4_y0;
  wire h_s_arrmul16_fa14_4_y2;
  wire h_s_arrmul16_fa14_4_y4;
  wire h_s_arrmul16_nand15_4_y0;
  wire h_s_arrmul16_fa15_4_y2;
  wire h_s_arrmul16_fa15_4_y4;
  wire h_s_arrmul16_and0_5_y0;
  wire h_s_arrmul16_ha0_5_y0;
  wire h_s_arrmul16_ha0_5_y1;
  wire h_s_arrmul16_and1_5_y0;
  wire h_s_arrmul16_fa1_5_y2;
  wire h_s_arrmul16_fa1_5_y4;
  wire h_s_arrmul16_and2_5_y0;
  wire h_s_arrmul16_fa2_5_y2;
  wire h_s_arrmul16_fa2_5_y4;
  wire h_s_arrmul16_and3_5_y0;
  wire h_s_arrmul16_fa3_5_y2;
  wire h_s_arrmul16_fa3_5_y4;
  wire h_s_arrmul16_and4_5_y0;
  wire h_s_arrmul16_fa4_5_y2;
  wire h_s_arrmul16_fa4_5_y4;
  wire h_s_arrmul16_and5_5_y0;
  wire h_s_arrmul16_fa5_5_y2;
  wire h_s_arrmul16_fa5_5_y4;
  wire h_s_arrmul16_and6_5_y0;
  wire h_s_arrmul16_fa6_5_y2;
  wire h_s_arrmul16_fa6_5_y4;
  wire h_s_arrmul16_and7_5_y0;
  wire h_s_arrmul16_fa7_5_y2;
  wire h_s_arrmul16_fa7_5_y4;
  wire h_s_arrmul16_and8_5_y0;
  wire h_s_arrmul16_fa8_5_y2;
  wire h_s_arrmul16_fa8_5_y4;
  wire h_s_arrmul16_and9_5_y0;
  wire h_s_arrmul16_fa9_5_y2;
  wire h_s_arrmul16_fa9_5_y4;
  wire h_s_arrmul16_and10_5_y0;
  wire h_s_arrmul16_fa10_5_y2;
  wire h_s_arrmul16_fa10_5_y4;
  wire h_s_arrmul16_and11_5_y0;
  wire h_s_arrmul16_fa11_5_y2;
  wire h_s_arrmul16_fa11_5_y4;
  wire h_s_arrmul16_and12_5_y0;
  wire h_s_arrmul16_fa12_5_y2;
  wire h_s_arrmul16_fa12_5_y4;
  wire h_s_arrmul16_and13_5_y0;
  wire h_s_arrmul16_fa13_5_y2;
  wire h_s_arrmul16_fa13_5_y4;
  wire h_s_arrmul16_and14_5_y0;
  wire h_s_arrmul16_fa14_5_y2;
  wire h_s_arrmul16_fa14_5_y4;
  wire h_s_arrmul16_nand15_5_y0;
  wire h_s_arrmul16_fa15_5_y2;
  wire h_s_arrmul16_fa15_5_y4;
  wire h_s_arrmul16_and0_6_y0;
  wire h_s_arrmul16_ha0_6_y0;
  wire h_s_arrmul16_ha0_6_y1;
  wire h_s_arrmul16_and1_6_y0;
  wire h_s_arrmul16_fa1_6_y2;
  wire h_s_arrmul16_fa1_6_y4;
  wire h_s_arrmul16_and2_6_y0;
  wire h_s_arrmul16_fa2_6_y2;
  wire h_s_arrmul16_fa2_6_y4;
  wire h_s_arrmul16_and3_6_y0;
  wire h_s_arrmul16_fa3_6_y2;
  wire h_s_arrmul16_fa3_6_y4;
  wire h_s_arrmul16_and4_6_y0;
  wire h_s_arrmul16_fa4_6_y2;
  wire h_s_arrmul16_fa4_6_y4;
  wire h_s_arrmul16_and5_6_y0;
  wire h_s_arrmul16_fa5_6_y2;
  wire h_s_arrmul16_fa5_6_y4;
  wire h_s_arrmul16_and6_6_y0;
  wire h_s_arrmul16_fa6_6_y2;
  wire h_s_arrmul16_fa6_6_y4;
  wire h_s_arrmul16_and7_6_y0;
  wire h_s_arrmul16_fa7_6_y2;
  wire h_s_arrmul16_fa7_6_y4;
  wire h_s_arrmul16_and8_6_y0;
  wire h_s_arrmul16_fa8_6_y2;
  wire h_s_arrmul16_fa8_6_y4;
  wire h_s_arrmul16_and9_6_y0;
  wire h_s_arrmul16_fa9_6_y2;
  wire h_s_arrmul16_fa9_6_y4;
  wire h_s_arrmul16_and10_6_y0;
  wire h_s_arrmul16_fa10_6_y2;
  wire h_s_arrmul16_fa10_6_y4;
  wire h_s_arrmul16_and11_6_y0;
  wire h_s_arrmul16_fa11_6_y2;
  wire h_s_arrmul16_fa11_6_y4;
  wire h_s_arrmul16_and12_6_y0;
  wire h_s_arrmul16_fa12_6_y2;
  wire h_s_arrmul16_fa12_6_y4;
  wire h_s_arrmul16_and13_6_y0;
  wire h_s_arrmul16_fa13_6_y2;
  wire h_s_arrmul16_fa13_6_y4;
  wire h_s_arrmul16_and14_6_y0;
  wire h_s_arrmul16_fa14_6_y2;
  wire h_s_arrmul16_fa14_6_y4;
  wire h_s_arrmul16_nand15_6_y0;
  wire h_s_arrmul16_fa15_6_y2;
  wire h_s_arrmul16_fa15_6_y4;
  wire h_s_arrmul16_and0_7_y0;
  wire h_s_arrmul16_ha0_7_y0;
  wire h_s_arrmul16_ha0_7_y1;
  wire h_s_arrmul16_and1_7_y0;
  wire h_s_arrmul16_fa1_7_y2;
  wire h_s_arrmul16_fa1_7_y4;
  wire h_s_arrmul16_and2_7_y0;
  wire h_s_arrmul16_fa2_7_y2;
  wire h_s_arrmul16_fa2_7_y4;
  wire h_s_arrmul16_and3_7_y0;
  wire h_s_arrmul16_fa3_7_y2;
  wire h_s_arrmul16_fa3_7_y4;
  wire h_s_arrmul16_and4_7_y0;
  wire h_s_arrmul16_fa4_7_y2;
  wire h_s_arrmul16_fa4_7_y4;
  wire h_s_arrmul16_and5_7_y0;
  wire h_s_arrmul16_fa5_7_y2;
  wire h_s_arrmul16_fa5_7_y4;
  wire h_s_arrmul16_and6_7_y0;
  wire h_s_arrmul16_fa6_7_y2;
  wire h_s_arrmul16_fa6_7_y4;
  wire h_s_arrmul16_and7_7_y0;
  wire h_s_arrmul16_fa7_7_y2;
  wire h_s_arrmul16_fa7_7_y4;
  wire h_s_arrmul16_and8_7_y0;
  wire h_s_arrmul16_fa8_7_y2;
  wire h_s_arrmul16_fa8_7_y4;
  wire h_s_arrmul16_and9_7_y0;
  wire h_s_arrmul16_fa9_7_y2;
  wire h_s_arrmul16_fa9_7_y4;
  wire h_s_arrmul16_and10_7_y0;
  wire h_s_arrmul16_fa10_7_y2;
  wire h_s_arrmul16_fa10_7_y4;
  wire h_s_arrmul16_and11_7_y0;
  wire h_s_arrmul16_fa11_7_y2;
  wire h_s_arrmul16_fa11_7_y4;
  wire h_s_arrmul16_and12_7_y0;
  wire h_s_arrmul16_fa12_7_y2;
  wire h_s_arrmul16_fa12_7_y4;
  wire h_s_arrmul16_and13_7_y0;
  wire h_s_arrmul16_fa13_7_y2;
  wire h_s_arrmul16_fa13_7_y4;
  wire h_s_arrmul16_and14_7_y0;
  wire h_s_arrmul16_fa14_7_y2;
  wire h_s_arrmul16_fa14_7_y4;
  wire h_s_arrmul16_nand15_7_y0;
  wire h_s_arrmul16_fa15_7_y2;
  wire h_s_arrmul16_fa15_7_y4;
  wire h_s_arrmul16_and0_8_y0;
  wire h_s_arrmul16_ha0_8_y0;
  wire h_s_arrmul16_ha0_8_y1;
  wire h_s_arrmul16_and1_8_y0;
  wire h_s_arrmul16_fa1_8_y2;
  wire h_s_arrmul16_fa1_8_y4;
  wire h_s_arrmul16_and2_8_y0;
  wire h_s_arrmul16_fa2_8_y2;
  wire h_s_arrmul16_fa2_8_y4;
  wire h_s_arrmul16_and3_8_y0;
  wire h_s_arrmul16_fa3_8_y2;
  wire h_s_arrmul16_fa3_8_y4;
  wire h_s_arrmul16_and4_8_y0;
  wire h_s_arrmul16_fa4_8_y2;
  wire h_s_arrmul16_fa4_8_y4;
  wire h_s_arrmul16_and5_8_y0;
  wire h_s_arrmul16_fa5_8_y2;
  wire h_s_arrmul16_fa5_8_y4;
  wire h_s_arrmul16_and6_8_y0;
  wire h_s_arrmul16_fa6_8_y2;
  wire h_s_arrmul16_fa6_8_y4;
  wire h_s_arrmul16_and7_8_y0;
  wire h_s_arrmul16_fa7_8_y2;
  wire h_s_arrmul16_fa7_8_y4;
  wire h_s_arrmul16_and8_8_y0;
  wire h_s_arrmul16_fa8_8_y2;
  wire h_s_arrmul16_fa8_8_y4;
  wire h_s_arrmul16_and9_8_y0;
  wire h_s_arrmul16_fa9_8_y2;
  wire h_s_arrmul16_fa9_8_y4;
  wire h_s_arrmul16_and10_8_y0;
  wire h_s_arrmul16_fa10_8_y2;
  wire h_s_arrmul16_fa10_8_y4;
  wire h_s_arrmul16_and11_8_y0;
  wire h_s_arrmul16_fa11_8_y2;
  wire h_s_arrmul16_fa11_8_y4;
  wire h_s_arrmul16_and12_8_y0;
  wire h_s_arrmul16_fa12_8_y2;
  wire h_s_arrmul16_fa12_8_y4;
  wire h_s_arrmul16_and13_8_y0;
  wire h_s_arrmul16_fa13_8_y2;
  wire h_s_arrmul16_fa13_8_y4;
  wire h_s_arrmul16_and14_8_y0;
  wire h_s_arrmul16_fa14_8_y2;
  wire h_s_arrmul16_fa14_8_y4;
  wire h_s_arrmul16_nand15_8_y0;
  wire h_s_arrmul16_fa15_8_y2;
  wire h_s_arrmul16_fa15_8_y4;
  wire h_s_arrmul16_and0_9_y0;
  wire h_s_arrmul16_ha0_9_y0;
  wire h_s_arrmul16_ha0_9_y1;
  wire h_s_arrmul16_and1_9_y0;
  wire h_s_arrmul16_fa1_9_y2;
  wire h_s_arrmul16_fa1_9_y4;
  wire h_s_arrmul16_and2_9_y0;
  wire h_s_arrmul16_fa2_9_y2;
  wire h_s_arrmul16_fa2_9_y4;
  wire h_s_arrmul16_and3_9_y0;
  wire h_s_arrmul16_fa3_9_y2;
  wire h_s_arrmul16_fa3_9_y4;
  wire h_s_arrmul16_and4_9_y0;
  wire h_s_arrmul16_fa4_9_y2;
  wire h_s_arrmul16_fa4_9_y4;
  wire h_s_arrmul16_and5_9_y0;
  wire h_s_arrmul16_fa5_9_y2;
  wire h_s_arrmul16_fa5_9_y4;
  wire h_s_arrmul16_and6_9_y0;
  wire h_s_arrmul16_fa6_9_y2;
  wire h_s_arrmul16_fa6_9_y4;
  wire h_s_arrmul16_and7_9_y0;
  wire h_s_arrmul16_fa7_9_y2;
  wire h_s_arrmul16_fa7_9_y4;
  wire h_s_arrmul16_and8_9_y0;
  wire h_s_arrmul16_fa8_9_y2;
  wire h_s_arrmul16_fa8_9_y4;
  wire h_s_arrmul16_and9_9_y0;
  wire h_s_arrmul16_fa9_9_y2;
  wire h_s_arrmul16_fa9_9_y4;
  wire h_s_arrmul16_and10_9_y0;
  wire h_s_arrmul16_fa10_9_y2;
  wire h_s_arrmul16_fa10_9_y4;
  wire h_s_arrmul16_and11_9_y0;
  wire h_s_arrmul16_fa11_9_y2;
  wire h_s_arrmul16_fa11_9_y4;
  wire h_s_arrmul16_and12_9_y0;
  wire h_s_arrmul16_fa12_9_y2;
  wire h_s_arrmul16_fa12_9_y4;
  wire h_s_arrmul16_and13_9_y0;
  wire h_s_arrmul16_fa13_9_y2;
  wire h_s_arrmul16_fa13_9_y4;
  wire h_s_arrmul16_and14_9_y0;
  wire h_s_arrmul16_fa14_9_y2;
  wire h_s_arrmul16_fa14_9_y4;
  wire h_s_arrmul16_nand15_9_y0;
  wire h_s_arrmul16_fa15_9_y2;
  wire h_s_arrmul16_fa15_9_y4;
  wire h_s_arrmul16_and0_10_y0;
  wire h_s_arrmul16_ha0_10_y0;
  wire h_s_arrmul16_ha0_10_y1;
  wire h_s_arrmul16_and1_10_y0;
  wire h_s_arrmul16_fa1_10_y2;
  wire h_s_arrmul16_fa1_10_y4;
  wire h_s_arrmul16_and2_10_y0;
  wire h_s_arrmul16_fa2_10_y2;
  wire h_s_arrmul16_fa2_10_y4;
  wire h_s_arrmul16_and3_10_y0;
  wire h_s_arrmul16_fa3_10_y2;
  wire h_s_arrmul16_fa3_10_y4;
  wire h_s_arrmul16_and4_10_y0;
  wire h_s_arrmul16_fa4_10_y2;
  wire h_s_arrmul16_fa4_10_y4;
  wire h_s_arrmul16_and5_10_y0;
  wire h_s_arrmul16_fa5_10_y2;
  wire h_s_arrmul16_fa5_10_y4;
  wire h_s_arrmul16_and6_10_y0;
  wire h_s_arrmul16_fa6_10_y2;
  wire h_s_arrmul16_fa6_10_y4;
  wire h_s_arrmul16_and7_10_y0;
  wire h_s_arrmul16_fa7_10_y2;
  wire h_s_arrmul16_fa7_10_y4;
  wire h_s_arrmul16_and8_10_y0;
  wire h_s_arrmul16_fa8_10_y2;
  wire h_s_arrmul16_fa8_10_y4;
  wire h_s_arrmul16_and9_10_y0;
  wire h_s_arrmul16_fa9_10_y2;
  wire h_s_arrmul16_fa9_10_y4;
  wire h_s_arrmul16_and10_10_y0;
  wire h_s_arrmul16_fa10_10_y2;
  wire h_s_arrmul16_fa10_10_y4;
  wire h_s_arrmul16_and11_10_y0;
  wire h_s_arrmul16_fa11_10_y2;
  wire h_s_arrmul16_fa11_10_y4;
  wire h_s_arrmul16_and12_10_y0;
  wire h_s_arrmul16_fa12_10_y2;
  wire h_s_arrmul16_fa12_10_y4;
  wire h_s_arrmul16_and13_10_y0;
  wire h_s_arrmul16_fa13_10_y2;
  wire h_s_arrmul16_fa13_10_y4;
  wire h_s_arrmul16_and14_10_y0;
  wire h_s_arrmul16_fa14_10_y2;
  wire h_s_arrmul16_fa14_10_y4;
  wire h_s_arrmul16_nand15_10_y0;
  wire h_s_arrmul16_fa15_10_y2;
  wire h_s_arrmul16_fa15_10_y4;
  wire h_s_arrmul16_and0_11_y0;
  wire h_s_arrmul16_ha0_11_y0;
  wire h_s_arrmul16_ha0_11_y1;
  wire h_s_arrmul16_and1_11_y0;
  wire h_s_arrmul16_fa1_11_y2;
  wire h_s_arrmul16_fa1_11_y4;
  wire h_s_arrmul16_and2_11_y0;
  wire h_s_arrmul16_fa2_11_y2;
  wire h_s_arrmul16_fa2_11_y4;
  wire h_s_arrmul16_and3_11_y0;
  wire h_s_arrmul16_fa3_11_y2;
  wire h_s_arrmul16_fa3_11_y4;
  wire h_s_arrmul16_and4_11_y0;
  wire h_s_arrmul16_fa4_11_y2;
  wire h_s_arrmul16_fa4_11_y4;
  wire h_s_arrmul16_and5_11_y0;
  wire h_s_arrmul16_fa5_11_y2;
  wire h_s_arrmul16_fa5_11_y4;
  wire h_s_arrmul16_and6_11_y0;
  wire h_s_arrmul16_fa6_11_y2;
  wire h_s_arrmul16_fa6_11_y4;
  wire h_s_arrmul16_and7_11_y0;
  wire h_s_arrmul16_fa7_11_y2;
  wire h_s_arrmul16_fa7_11_y4;
  wire h_s_arrmul16_and8_11_y0;
  wire h_s_arrmul16_fa8_11_y2;
  wire h_s_arrmul16_fa8_11_y4;
  wire h_s_arrmul16_and9_11_y0;
  wire h_s_arrmul16_fa9_11_y2;
  wire h_s_arrmul16_fa9_11_y4;
  wire h_s_arrmul16_and10_11_y0;
  wire h_s_arrmul16_fa10_11_y2;
  wire h_s_arrmul16_fa10_11_y4;
  wire h_s_arrmul16_and11_11_y0;
  wire h_s_arrmul16_fa11_11_y2;
  wire h_s_arrmul16_fa11_11_y4;
  wire h_s_arrmul16_and12_11_y0;
  wire h_s_arrmul16_fa12_11_y2;
  wire h_s_arrmul16_fa12_11_y4;
  wire h_s_arrmul16_and13_11_y0;
  wire h_s_arrmul16_fa13_11_y2;
  wire h_s_arrmul16_fa13_11_y4;
  wire h_s_arrmul16_and14_11_y0;
  wire h_s_arrmul16_fa14_11_y2;
  wire h_s_arrmul16_fa14_11_y4;
  wire h_s_arrmul16_nand15_11_y0;
  wire h_s_arrmul16_fa15_11_y2;
  wire h_s_arrmul16_fa15_11_y4;
  wire h_s_arrmul16_and0_12_y0;
  wire h_s_arrmul16_ha0_12_y0;
  wire h_s_arrmul16_ha0_12_y1;
  wire h_s_arrmul16_and1_12_y0;
  wire h_s_arrmul16_fa1_12_y2;
  wire h_s_arrmul16_fa1_12_y4;
  wire h_s_arrmul16_and2_12_y0;
  wire h_s_arrmul16_fa2_12_y2;
  wire h_s_arrmul16_fa2_12_y4;
  wire h_s_arrmul16_and3_12_y0;
  wire h_s_arrmul16_fa3_12_y2;
  wire h_s_arrmul16_fa3_12_y4;
  wire h_s_arrmul16_and4_12_y0;
  wire h_s_arrmul16_fa4_12_y2;
  wire h_s_arrmul16_fa4_12_y4;
  wire h_s_arrmul16_and5_12_y0;
  wire h_s_arrmul16_fa5_12_y2;
  wire h_s_arrmul16_fa5_12_y4;
  wire h_s_arrmul16_and6_12_y0;
  wire h_s_arrmul16_fa6_12_y2;
  wire h_s_arrmul16_fa6_12_y4;
  wire h_s_arrmul16_and7_12_y0;
  wire h_s_arrmul16_fa7_12_y2;
  wire h_s_arrmul16_fa7_12_y4;
  wire h_s_arrmul16_and8_12_y0;
  wire h_s_arrmul16_fa8_12_y2;
  wire h_s_arrmul16_fa8_12_y4;
  wire h_s_arrmul16_and9_12_y0;
  wire h_s_arrmul16_fa9_12_y2;
  wire h_s_arrmul16_fa9_12_y4;
  wire h_s_arrmul16_and10_12_y0;
  wire h_s_arrmul16_fa10_12_y2;
  wire h_s_arrmul16_fa10_12_y4;
  wire h_s_arrmul16_and11_12_y0;
  wire h_s_arrmul16_fa11_12_y2;
  wire h_s_arrmul16_fa11_12_y4;
  wire h_s_arrmul16_and12_12_y0;
  wire h_s_arrmul16_fa12_12_y2;
  wire h_s_arrmul16_fa12_12_y4;
  wire h_s_arrmul16_and13_12_y0;
  wire h_s_arrmul16_fa13_12_y2;
  wire h_s_arrmul16_fa13_12_y4;
  wire h_s_arrmul16_and14_12_y0;
  wire h_s_arrmul16_fa14_12_y2;
  wire h_s_arrmul16_fa14_12_y4;
  wire h_s_arrmul16_nand15_12_y0;
  wire h_s_arrmul16_fa15_12_y2;
  wire h_s_arrmul16_fa15_12_y4;
  wire h_s_arrmul16_and0_13_y0;
  wire h_s_arrmul16_ha0_13_y0;
  wire h_s_arrmul16_ha0_13_y1;
  wire h_s_arrmul16_and1_13_y0;
  wire h_s_arrmul16_fa1_13_y2;
  wire h_s_arrmul16_fa1_13_y4;
  wire h_s_arrmul16_and2_13_y0;
  wire h_s_arrmul16_fa2_13_y2;
  wire h_s_arrmul16_fa2_13_y4;
  wire h_s_arrmul16_and3_13_y0;
  wire h_s_arrmul16_fa3_13_y2;
  wire h_s_arrmul16_fa3_13_y4;
  wire h_s_arrmul16_and4_13_y0;
  wire h_s_arrmul16_fa4_13_y2;
  wire h_s_arrmul16_fa4_13_y4;
  wire h_s_arrmul16_and5_13_y0;
  wire h_s_arrmul16_fa5_13_y2;
  wire h_s_arrmul16_fa5_13_y4;
  wire h_s_arrmul16_and6_13_y0;
  wire h_s_arrmul16_fa6_13_y2;
  wire h_s_arrmul16_fa6_13_y4;
  wire h_s_arrmul16_and7_13_y0;
  wire h_s_arrmul16_fa7_13_y2;
  wire h_s_arrmul16_fa7_13_y4;
  wire h_s_arrmul16_and8_13_y0;
  wire h_s_arrmul16_fa8_13_y2;
  wire h_s_arrmul16_fa8_13_y4;
  wire h_s_arrmul16_and9_13_y0;
  wire h_s_arrmul16_fa9_13_y2;
  wire h_s_arrmul16_fa9_13_y4;
  wire h_s_arrmul16_and10_13_y0;
  wire h_s_arrmul16_fa10_13_y2;
  wire h_s_arrmul16_fa10_13_y4;
  wire h_s_arrmul16_and11_13_y0;
  wire h_s_arrmul16_fa11_13_y2;
  wire h_s_arrmul16_fa11_13_y4;
  wire h_s_arrmul16_and12_13_y0;
  wire h_s_arrmul16_fa12_13_y2;
  wire h_s_arrmul16_fa12_13_y4;
  wire h_s_arrmul16_and13_13_y0;
  wire h_s_arrmul16_fa13_13_y2;
  wire h_s_arrmul16_fa13_13_y4;
  wire h_s_arrmul16_and14_13_y0;
  wire h_s_arrmul16_fa14_13_y2;
  wire h_s_arrmul16_fa14_13_y4;
  wire h_s_arrmul16_nand15_13_y0;
  wire h_s_arrmul16_fa15_13_y2;
  wire h_s_arrmul16_fa15_13_y4;
  wire h_s_arrmul16_and0_14_y0;
  wire h_s_arrmul16_ha0_14_y0;
  wire h_s_arrmul16_ha0_14_y1;
  wire h_s_arrmul16_and1_14_y0;
  wire h_s_arrmul16_fa1_14_y2;
  wire h_s_arrmul16_fa1_14_y4;
  wire h_s_arrmul16_and2_14_y0;
  wire h_s_arrmul16_fa2_14_y2;
  wire h_s_arrmul16_fa2_14_y4;
  wire h_s_arrmul16_and3_14_y0;
  wire h_s_arrmul16_fa3_14_y2;
  wire h_s_arrmul16_fa3_14_y4;
  wire h_s_arrmul16_and4_14_y0;
  wire h_s_arrmul16_fa4_14_y2;
  wire h_s_arrmul16_fa4_14_y4;
  wire h_s_arrmul16_and5_14_y0;
  wire h_s_arrmul16_fa5_14_y2;
  wire h_s_arrmul16_fa5_14_y4;
  wire h_s_arrmul16_and6_14_y0;
  wire h_s_arrmul16_fa6_14_y2;
  wire h_s_arrmul16_fa6_14_y4;
  wire h_s_arrmul16_and7_14_y0;
  wire h_s_arrmul16_fa7_14_y2;
  wire h_s_arrmul16_fa7_14_y4;
  wire h_s_arrmul16_and8_14_y0;
  wire h_s_arrmul16_fa8_14_y2;
  wire h_s_arrmul16_fa8_14_y4;
  wire h_s_arrmul16_and9_14_y0;
  wire h_s_arrmul16_fa9_14_y2;
  wire h_s_arrmul16_fa9_14_y4;
  wire h_s_arrmul16_and10_14_y0;
  wire h_s_arrmul16_fa10_14_y2;
  wire h_s_arrmul16_fa10_14_y4;
  wire h_s_arrmul16_and11_14_y0;
  wire h_s_arrmul16_fa11_14_y2;
  wire h_s_arrmul16_fa11_14_y4;
  wire h_s_arrmul16_and12_14_y0;
  wire h_s_arrmul16_fa12_14_y2;
  wire h_s_arrmul16_fa12_14_y4;
  wire h_s_arrmul16_and13_14_y0;
  wire h_s_arrmul16_fa13_14_y2;
  wire h_s_arrmul16_fa13_14_y4;
  wire h_s_arrmul16_and14_14_y0;
  wire h_s_arrmul16_fa14_14_y2;
  wire h_s_arrmul16_fa14_14_y4;
  wire h_s_arrmul16_nand15_14_y0;
  wire h_s_arrmul16_fa15_14_y2;
  wire h_s_arrmul16_fa15_14_y4;
  wire h_s_arrmul16_nand0_15_y0;
  wire h_s_arrmul16_ha0_15_y0;
  wire h_s_arrmul16_ha0_15_y1;
  wire h_s_arrmul16_nand1_15_y0;
  wire h_s_arrmul16_fa1_15_y2;
  wire h_s_arrmul16_fa1_15_y4;
  wire h_s_arrmul16_nand2_15_y0;
  wire h_s_arrmul16_fa2_15_y2;
  wire h_s_arrmul16_fa2_15_y4;
  wire h_s_arrmul16_nand3_15_y0;
  wire h_s_arrmul16_fa3_15_y2;
  wire h_s_arrmul16_fa3_15_y4;
  wire h_s_arrmul16_nand4_15_y0;
  wire h_s_arrmul16_fa4_15_y2;
  wire h_s_arrmul16_fa4_15_y4;
  wire h_s_arrmul16_nand5_15_y0;
  wire h_s_arrmul16_fa5_15_y2;
  wire h_s_arrmul16_fa5_15_y4;
  wire h_s_arrmul16_nand6_15_y0;
  wire h_s_arrmul16_fa6_15_y2;
  wire h_s_arrmul16_fa6_15_y4;
  wire h_s_arrmul16_nand7_15_y0;
  wire h_s_arrmul16_fa7_15_y2;
  wire h_s_arrmul16_fa7_15_y4;
  wire h_s_arrmul16_nand8_15_y0;
  wire h_s_arrmul16_fa8_15_y2;
  wire h_s_arrmul16_fa8_15_y4;
  wire h_s_arrmul16_nand9_15_y0;
  wire h_s_arrmul16_fa9_15_y2;
  wire h_s_arrmul16_fa9_15_y4;
  wire h_s_arrmul16_nand10_15_y0;
  wire h_s_arrmul16_fa10_15_y2;
  wire h_s_arrmul16_fa10_15_y4;
  wire h_s_arrmul16_nand11_15_y0;
  wire h_s_arrmul16_fa11_15_y2;
  wire h_s_arrmul16_fa11_15_y4;
  wire h_s_arrmul16_nand12_15_y0;
  wire h_s_arrmul16_fa12_15_y2;
  wire h_s_arrmul16_fa12_15_y4;
  wire h_s_arrmul16_nand13_15_y0;
  wire h_s_arrmul16_fa13_15_y2;
  wire h_s_arrmul16_fa13_15_y4;
  wire h_s_arrmul16_nand14_15_y0;
  wire h_s_arrmul16_fa14_15_y2;
  wire h_s_arrmul16_fa14_15_y4;
  wire h_s_arrmul16_and15_15_y0;
  wire h_s_arrmul16_fa15_15_y2;
  wire h_s_arrmul16_fa15_15_y4;
  wire h_s_arrmul16_xor16_15_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_arrmul16_and0_0_y0(a_0, b_0, h_s_arrmul16_and0_0_y0);
  and_gate and_gate_h_s_arrmul16_and1_0_y0(a_1, b_0, h_s_arrmul16_and1_0_y0);
  and_gate and_gate_h_s_arrmul16_and2_0_y0(a_2, b_0, h_s_arrmul16_and2_0_y0);
  and_gate and_gate_h_s_arrmul16_and3_0_y0(a_3, b_0, h_s_arrmul16_and3_0_y0);
  and_gate and_gate_h_s_arrmul16_and4_0_y0(a_4, b_0, h_s_arrmul16_and4_0_y0);
  and_gate and_gate_h_s_arrmul16_and5_0_y0(a_5, b_0, h_s_arrmul16_and5_0_y0);
  and_gate and_gate_h_s_arrmul16_and6_0_y0(a_6, b_0, h_s_arrmul16_and6_0_y0);
  and_gate and_gate_h_s_arrmul16_and7_0_y0(a_7, b_0, h_s_arrmul16_and7_0_y0);
  and_gate and_gate_h_s_arrmul16_and8_0_y0(a_8, b_0, h_s_arrmul16_and8_0_y0);
  and_gate and_gate_h_s_arrmul16_and9_0_y0(a_9, b_0, h_s_arrmul16_and9_0_y0);
  and_gate and_gate_h_s_arrmul16_and10_0_y0(a_10, b_0, h_s_arrmul16_and10_0_y0);
  and_gate and_gate_h_s_arrmul16_and11_0_y0(a_11, b_0, h_s_arrmul16_and11_0_y0);
  and_gate and_gate_h_s_arrmul16_and12_0_y0(a_12, b_0, h_s_arrmul16_and12_0_y0);
  and_gate and_gate_h_s_arrmul16_and13_0_y0(a_13, b_0, h_s_arrmul16_and13_0_y0);
  and_gate and_gate_h_s_arrmul16_and14_0_y0(a_14, b_0, h_s_arrmul16_and14_0_y0);
  nand_gate nand_gate_h_s_arrmul16_nand15_0_y0(a_15, b_0, h_s_arrmul16_nand15_0_y0);
  and_gate and_gate_h_s_arrmul16_and0_1_y0(a_0, b_1, h_s_arrmul16_and0_1_y0);
  ha ha_h_s_arrmul16_ha0_1_y0(h_s_arrmul16_and0_1_y0, h_s_arrmul16_and1_0_y0, h_s_arrmul16_ha0_1_y0, h_s_arrmul16_ha0_1_y1);
  and_gate and_gate_h_s_arrmul16_and1_1_y0(a_1, b_1, h_s_arrmul16_and1_1_y0);
  fa fa_h_s_arrmul16_fa1_1_y2(h_s_arrmul16_and1_1_y0, h_s_arrmul16_and2_0_y0, h_s_arrmul16_ha0_1_y1, h_s_arrmul16_fa1_1_y2, h_s_arrmul16_fa1_1_y4);
  and_gate and_gate_h_s_arrmul16_and2_1_y0(a_2, b_1, h_s_arrmul16_and2_1_y0);
  fa fa_h_s_arrmul16_fa2_1_y2(h_s_arrmul16_and2_1_y0, h_s_arrmul16_and3_0_y0, h_s_arrmul16_fa1_1_y4, h_s_arrmul16_fa2_1_y2, h_s_arrmul16_fa2_1_y4);
  and_gate and_gate_h_s_arrmul16_and3_1_y0(a_3, b_1, h_s_arrmul16_and3_1_y0);
  fa fa_h_s_arrmul16_fa3_1_y2(h_s_arrmul16_and3_1_y0, h_s_arrmul16_and4_0_y0, h_s_arrmul16_fa2_1_y4, h_s_arrmul16_fa3_1_y2, h_s_arrmul16_fa3_1_y4);
  and_gate and_gate_h_s_arrmul16_and4_1_y0(a_4, b_1, h_s_arrmul16_and4_1_y0);
  fa fa_h_s_arrmul16_fa4_1_y2(h_s_arrmul16_and4_1_y0, h_s_arrmul16_and5_0_y0, h_s_arrmul16_fa3_1_y4, h_s_arrmul16_fa4_1_y2, h_s_arrmul16_fa4_1_y4);
  and_gate and_gate_h_s_arrmul16_and5_1_y0(a_5, b_1, h_s_arrmul16_and5_1_y0);
  fa fa_h_s_arrmul16_fa5_1_y2(h_s_arrmul16_and5_1_y0, h_s_arrmul16_and6_0_y0, h_s_arrmul16_fa4_1_y4, h_s_arrmul16_fa5_1_y2, h_s_arrmul16_fa5_1_y4);
  and_gate and_gate_h_s_arrmul16_and6_1_y0(a_6, b_1, h_s_arrmul16_and6_1_y0);
  fa fa_h_s_arrmul16_fa6_1_y2(h_s_arrmul16_and6_1_y0, h_s_arrmul16_and7_0_y0, h_s_arrmul16_fa5_1_y4, h_s_arrmul16_fa6_1_y2, h_s_arrmul16_fa6_1_y4);
  and_gate and_gate_h_s_arrmul16_and7_1_y0(a_7, b_1, h_s_arrmul16_and7_1_y0);
  fa fa_h_s_arrmul16_fa7_1_y2(h_s_arrmul16_and7_1_y0, h_s_arrmul16_and8_0_y0, h_s_arrmul16_fa6_1_y4, h_s_arrmul16_fa7_1_y2, h_s_arrmul16_fa7_1_y4);
  and_gate and_gate_h_s_arrmul16_and8_1_y0(a_8, b_1, h_s_arrmul16_and8_1_y0);
  fa fa_h_s_arrmul16_fa8_1_y2(h_s_arrmul16_and8_1_y0, h_s_arrmul16_and9_0_y0, h_s_arrmul16_fa7_1_y4, h_s_arrmul16_fa8_1_y2, h_s_arrmul16_fa8_1_y4);
  and_gate and_gate_h_s_arrmul16_and9_1_y0(a_9, b_1, h_s_arrmul16_and9_1_y0);
  fa fa_h_s_arrmul16_fa9_1_y2(h_s_arrmul16_and9_1_y0, h_s_arrmul16_and10_0_y0, h_s_arrmul16_fa8_1_y4, h_s_arrmul16_fa9_1_y2, h_s_arrmul16_fa9_1_y4);
  and_gate and_gate_h_s_arrmul16_and10_1_y0(a_10, b_1, h_s_arrmul16_and10_1_y0);
  fa fa_h_s_arrmul16_fa10_1_y2(h_s_arrmul16_and10_1_y0, h_s_arrmul16_and11_0_y0, h_s_arrmul16_fa9_1_y4, h_s_arrmul16_fa10_1_y2, h_s_arrmul16_fa10_1_y4);
  and_gate and_gate_h_s_arrmul16_and11_1_y0(a_11, b_1, h_s_arrmul16_and11_1_y0);
  fa fa_h_s_arrmul16_fa11_1_y2(h_s_arrmul16_and11_1_y0, h_s_arrmul16_and12_0_y0, h_s_arrmul16_fa10_1_y4, h_s_arrmul16_fa11_1_y2, h_s_arrmul16_fa11_1_y4);
  and_gate and_gate_h_s_arrmul16_and12_1_y0(a_12, b_1, h_s_arrmul16_and12_1_y0);
  fa fa_h_s_arrmul16_fa12_1_y2(h_s_arrmul16_and12_1_y0, h_s_arrmul16_and13_0_y0, h_s_arrmul16_fa11_1_y4, h_s_arrmul16_fa12_1_y2, h_s_arrmul16_fa12_1_y4);
  and_gate and_gate_h_s_arrmul16_and13_1_y0(a_13, b_1, h_s_arrmul16_and13_1_y0);
  fa fa_h_s_arrmul16_fa13_1_y2(h_s_arrmul16_and13_1_y0, h_s_arrmul16_and14_0_y0, h_s_arrmul16_fa12_1_y4, h_s_arrmul16_fa13_1_y2, h_s_arrmul16_fa13_1_y4);
  and_gate and_gate_h_s_arrmul16_and14_1_y0(a_14, b_1, h_s_arrmul16_and14_1_y0);
  fa fa_h_s_arrmul16_fa14_1_y2(h_s_arrmul16_and14_1_y0, h_s_arrmul16_nand15_0_y0, h_s_arrmul16_fa13_1_y4, h_s_arrmul16_fa14_1_y2, h_s_arrmul16_fa14_1_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_1_y0(a_15, b_1, h_s_arrmul16_nand15_1_y0);
  fa fa_h_s_arrmul16_fa15_1_y2(h_s_arrmul16_nand15_1_y0, constant_wire_1, h_s_arrmul16_fa14_1_y4, h_s_arrmul16_fa15_1_y2, h_s_arrmul16_fa15_1_y4);
  and_gate and_gate_h_s_arrmul16_and0_2_y0(a_0, b_2, h_s_arrmul16_and0_2_y0);
  ha ha_h_s_arrmul16_ha0_2_y0(h_s_arrmul16_and0_2_y0, h_s_arrmul16_fa1_1_y2, h_s_arrmul16_ha0_2_y0, h_s_arrmul16_ha0_2_y1);
  and_gate and_gate_h_s_arrmul16_and1_2_y0(a_1, b_2, h_s_arrmul16_and1_2_y0);
  fa fa_h_s_arrmul16_fa1_2_y2(h_s_arrmul16_and1_2_y0, h_s_arrmul16_fa2_1_y2, h_s_arrmul16_ha0_2_y1, h_s_arrmul16_fa1_2_y2, h_s_arrmul16_fa1_2_y4);
  and_gate and_gate_h_s_arrmul16_and2_2_y0(a_2, b_2, h_s_arrmul16_and2_2_y0);
  fa fa_h_s_arrmul16_fa2_2_y2(h_s_arrmul16_and2_2_y0, h_s_arrmul16_fa3_1_y2, h_s_arrmul16_fa1_2_y4, h_s_arrmul16_fa2_2_y2, h_s_arrmul16_fa2_2_y4);
  and_gate and_gate_h_s_arrmul16_and3_2_y0(a_3, b_2, h_s_arrmul16_and3_2_y0);
  fa fa_h_s_arrmul16_fa3_2_y2(h_s_arrmul16_and3_2_y0, h_s_arrmul16_fa4_1_y2, h_s_arrmul16_fa2_2_y4, h_s_arrmul16_fa3_2_y2, h_s_arrmul16_fa3_2_y4);
  and_gate and_gate_h_s_arrmul16_and4_2_y0(a_4, b_2, h_s_arrmul16_and4_2_y0);
  fa fa_h_s_arrmul16_fa4_2_y2(h_s_arrmul16_and4_2_y0, h_s_arrmul16_fa5_1_y2, h_s_arrmul16_fa3_2_y4, h_s_arrmul16_fa4_2_y2, h_s_arrmul16_fa4_2_y4);
  and_gate and_gate_h_s_arrmul16_and5_2_y0(a_5, b_2, h_s_arrmul16_and5_2_y0);
  fa fa_h_s_arrmul16_fa5_2_y2(h_s_arrmul16_and5_2_y0, h_s_arrmul16_fa6_1_y2, h_s_arrmul16_fa4_2_y4, h_s_arrmul16_fa5_2_y2, h_s_arrmul16_fa5_2_y4);
  and_gate and_gate_h_s_arrmul16_and6_2_y0(a_6, b_2, h_s_arrmul16_and6_2_y0);
  fa fa_h_s_arrmul16_fa6_2_y2(h_s_arrmul16_and6_2_y0, h_s_arrmul16_fa7_1_y2, h_s_arrmul16_fa5_2_y4, h_s_arrmul16_fa6_2_y2, h_s_arrmul16_fa6_2_y4);
  and_gate and_gate_h_s_arrmul16_and7_2_y0(a_7, b_2, h_s_arrmul16_and7_2_y0);
  fa fa_h_s_arrmul16_fa7_2_y2(h_s_arrmul16_and7_2_y0, h_s_arrmul16_fa8_1_y2, h_s_arrmul16_fa6_2_y4, h_s_arrmul16_fa7_2_y2, h_s_arrmul16_fa7_2_y4);
  and_gate and_gate_h_s_arrmul16_and8_2_y0(a_8, b_2, h_s_arrmul16_and8_2_y0);
  fa fa_h_s_arrmul16_fa8_2_y2(h_s_arrmul16_and8_2_y0, h_s_arrmul16_fa9_1_y2, h_s_arrmul16_fa7_2_y4, h_s_arrmul16_fa8_2_y2, h_s_arrmul16_fa8_2_y4);
  and_gate and_gate_h_s_arrmul16_and9_2_y0(a_9, b_2, h_s_arrmul16_and9_2_y0);
  fa fa_h_s_arrmul16_fa9_2_y2(h_s_arrmul16_and9_2_y0, h_s_arrmul16_fa10_1_y2, h_s_arrmul16_fa8_2_y4, h_s_arrmul16_fa9_2_y2, h_s_arrmul16_fa9_2_y4);
  and_gate and_gate_h_s_arrmul16_and10_2_y0(a_10, b_2, h_s_arrmul16_and10_2_y0);
  fa fa_h_s_arrmul16_fa10_2_y2(h_s_arrmul16_and10_2_y0, h_s_arrmul16_fa11_1_y2, h_s_arrmul16_fa9_2_y4, h_s_arrmul16_fa10_2_y2, h_s_arrmul16_fa10_2_y4);
  and_gate and_gate_h_s_arrmul16_and11_2_y0(a_11, b_2, h_s_arrmul16_and11_2_y0);
  fa fa_h_s_arrmul16_fa11_2_y2(h_s_arrmul16_and11_2_y0, h_s_arrmul16_fa12_1_y2, h_s_arrmul16_fa10_2_y4, h_s_arrmul16_fa11_2_y2, h_s_arrmul16_fa11_2_y4);
  and_gate and_gate_h_s_arrmul16_and12_2_y0(a_12, b_2, h_s_arrmul16_and12_2_y0);
  fa fa_h_s_arrmul16_fa12_2_y2(h_s_arrmul16_and12_2_y0, h_s_arrmul16_fa13_1_y2, h_s_arrmul16_fa11_2_y4, h_s_arrmul16_fa12_2_y2, h_s_arrmul16_fa12_2_y4);
  and_gate and_gate_h_s_arrmul16_and13_2_y0(a_13, b_2, h_s_arrmul16_and13_2_y0);
  fa fa_h_s_arrmul16_fa13_2_y2(h_s_arrmul16_and13_2_y0, h_s_arrmul16_fa14_1_y2, h_s_arrmul16_fa12_2_y4, h_s_arrmul16_fa13_2_y2, h_s_arrmul16_fa13_2_y4);
  and_gate and_gate_h_s_arrmul16_and14_2_y0(a_14, b_2, h_s_arrmul16_and14_2_y0);
  fa fa_h_s_arrmul16_fa14_2_y2(h_s_arrmul16_and14_2_y0, h_s_arrmul16_fa15_1_y2, h_s_arrmul16_fa13_2_y4, h_s_arrmul16_fa14_2_y2, h_s_arrmul16_fa14_2_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_2_y0(a_15, b_2, h_s_arrmul16_nand15_2_y0);
  fa fa_h_s_arrmul16_fa15_2_y2(h_s_arrmul16_nand15_2_y0, h_s_arrmul16_fa15_1_y4, h_s_arrmul16_fa14_2_y4, h_s_arrmul16_fa15_2_y2, h_s_arrmul16_fa15_2_y4);
  and_gate and_gate_h_s_arrmul16_and0_3_y0(a_0, b_3, h_s_arrmul16_and0_3_y0);
  ha ha_h_s_arrmul16_ha0_3_y0(h_s_arrmul16_and0_3_y0, h_s_arrmul16_fa1_2_y2, h_s_arrmul16_ha0_3_y0, h_s_arrmul16_ha0_3_y1);
  and_gate and_gate_h_s_arrmul16_and1_3_y0(a_1, b_3, h_s_arrmul16_and1_3_y0);
  fa fa_h_s_arrmul16_fa1_3_y2(h_s_arrmul16_and1_3_y0, h_s_arrmul16_fa2_2_y2, h_s_arrmul16_ha0_3_y1, h_s_arrmul16_fa1_3_y2, h_s_arrmul16_fa1_3_y4);
  and_gate and_gate_h_s_arrmul16_and2_3_y0(a_2, b_3, h_s_arrmul16_and2_3_y0);
  fa fa_h_s_arrmul16_fa2_3_y2(h_s_arrmul16_and2_3_y0, h_s_arrmul16_fa3_2_y2, h_s_arrmul16_fa1_3_y4, h_s_arrmul16_fa2_3_y2, h_s_arrmul16_fa2_3_y4);
  and_gate and_gate_h_s_arrmul16_and3_3_y0(a_3, b_3, h_s_arrmul16_and3_3_y0);
  fa fa_h_s_arrmul16_fa3_3_y2(h_s_arrmul16_and3_3_y0, h_s_arrmul16_fa4_2_y2, h_s_arrmul16_fa2_3_y4, h_s_arrmul16_fa3_3_y2, h_s_arrmul16_fa3_3_y4);
  and_gate and_gate_h_s_arrmul16_and4_3_y0(a_4, b_3, h_s_arrmul16_and4_3_y0);
  fa fa_h_s_arrmul16_fa4_3_y2(h_s_arrmul16_and4_3_y0, h_s_arrmul16_fa5_2_y2, h_s_arrmul16_fa3_3_y4, h_s_arrmul16_fa4_3_y2, h_s_arrmul16_fa4_3_y4);
  and_gate and_gate_h_s_arrmul16_and5_3_y0(a_5, b_3, h_s_arrmul16_and5_3_y0);
  fa fa_h_s_arrmul16_fa5_3_y2(h_s_arrmul16_and5_3_y0, h_s_arrmul16_fa6_2_y2, h_s_arrmul16_fa4_3_y4, h_s_arrmul16_fa5_3_y2, h_s_arrmul16_fa5_3_y4);
  and_gate and_gate_h_s_arrmul16_and6_3_y0(a_6, b_3, h_s_arrmul16_and6_3_y0);
  fa fa_h_s_arrmul16_fa6_3_y2(h_s_arrmul16_and6_3_y0, h_s_arrmul16_fa7_2_y2, h_s_arrmul16_fa5_3_y4, h_s_arrmul16_fa6_3_y2, h_s_arrmul16_fa6_3_y4);
  and_gate and_gate_h_s_arrmul16_and7_3_y0(a_7, b_3, h_s_arrmul16_and7_3_y0);
  fa fa_h_s_arrmul16_fa7_3_y2(h_s_arrmul16_and7_3_y0, h_s_arrmul16_fa8_2_y2, h_s_arrmul16_fa6_3_y4, h_s_arrmul16_fa7_3_y2, h_s_arrmul16_fa7_3_y4);
  and_gate and_gate_h_s_arrmul16_and8_3_y0(a_8, b_3, h_s_arrmul16_and8_3_y0);
  fa fa_h_s_arrmul16_fa8_3_y2(h_s_arrmul16_and8_3_y0, h_s_arrmul16_fa9_2_y2, h_s_arrmul16_fa7_3_y4, h_s_arrmul16_fa8_3_y2, h_s_arrmul16_fa8_3_y4);
  and_gate and_gate_h_s_arrmul16_and9_3_y0(a_9, b_3, h_s_arrmul16_and9_3_y0);
  fa fa_h_s_arrmul16_fa9_3_y2(h_s_arrmul16_and9_3_y0, h_s_arrmul16_fa10_2_y2, h_s_arrmul16_fa8_3_y4, h_s_arrmul16_fa9_3_y2, h_s_arrmul16_fa9_3_y4);
  and_gate and_gate_h_s_arrmul16_and10_3_y0(a_10, b_3, h_s_arrmul16_and10_3_y0);
  fa fa_h_s_arrmul16_fa10_3_y2(h_s_arrmul16_and10_3_y0, h_s_arrmul16_fa11_2_y2, h_s_arrmul16_fa9_3_y4, h_s_arrmul16_fa10_3_y2, h_s_arrmul16_fa10_3_y4);
  and_gate and_gate_h_s_arrmul16_and11_3_y0(a_11, b_3, h_s_arrmul16_and11_3_y0);
  fa fa_h_s_arrmul16_fa11_3_y2(h_s_arrmul16_and11_3_y0, h_s_arrmul16_fa12_2_y2, h_s_arrmul16_fa10_3_y4, h_s_arrmul16_fa11_3_y2, h_s_arrmul16_fa11_3_y4);
  and_gate and_gate_h_s_arrmul16_and12_3_y0(a_12, b_3, h_s_arrmul16_and12_3_y0);
  fa fa_h_s_arrmul16_fa12_3_y2(h_s_arrmul16_and12_3_y0, h_s_arrmul16_fa13_2_y2, h_s_arrmul16_fa11_3_y4, h_s_arrmul16_fa12_3_y2, h_s_arrmul16_fa12_3_y4);
  and_gate and_gate_h_s_arrmul16_and13_3_y0(a_13, b_3, h_s_arrmul16_and13_3_y0);
  fa fa_h_s_arrmul16_fa13_3_y2(h_s_arrmul16_and13_3_y0, h_s_arrmul16_fa14_2_y2, h_s_arrmul16_fa12_3_y4, h_s_arrmul16_fa13_3_y2, h_s_arrmul16_fa13_3_y4);
  and_gate and_gate_h_s_arrmul16_and14_3_y0(a_14, b_3, h_s_arrmul16_and14_3_y0);
  fa fa_h_s_arrmul16_fa14_3_y2(h_s_arrmul16_and14_3_y0, h_s_arrmul16_fa15_2_y2, h_s_arrmul16_fa13_3_y4, h_s_arrmul16_fa14_3_y2, h_s_arrmul16_fa14_3_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_3_y0(a_15, b_3, h_s_arrmul16_nand15_3_y0);
  fa fa_h_s_arrmul16_fa15_3_y2(h_s_arrmul16_nand15_3_y0, h_s_arrmul16_fa15_2_y4, h_s_arrmul16_fa14_3_y4, h_s_arrmul16_fa15_3_y2, h_s_arrmul16_fa15_3_y4);
  and_gate and_gate_h_s_arrmul16_and0_4_y0(a_0, b_4, h_s_arrmul16_and0_4_y0);
  ha ha_h_s_arrmul16_ha0_4_y0(h_s_arrmul16_and0_4_y0, h_s_arrmul16_fa1_3_y2, h_s_arrmul16_ha0_4_y0, h_s_arrmul16_ha0_4_y1);
  and_gate and_gate_h_s_arrmul16_and1_4_y0(a_1, b_4, h_s_arrmul16_and1_4_y0);
  fa fa_h_s_arrmul16_fa1_4_y2(h_s_arrmul16_and1_4_y0, h_s_arrmul16_fa2_3_y2, h_s_arrmul16_ha0_4_y1, h_s_arrmul16_fa1_4_y2, h_s_arrmul16_fa1_4_y4);
  and_gate and_gate_h_s_arrmul16_and2_4_y0(a_2, b_4, h_s_arrmul16_and2_4_y0);
  fa fa_h_s_arrmul16_fa2_4_y2(h_s_arrmul16_and2_4_y0, h_s_arrmul16_fa3_3_y2, h_s_arrmul16_fa1_4_y4, h_s_arrmul16_fa2_4_y2, h_s_arrmul16_fa2_4_y4);
  and_gate and_gate_h_s_arrmul16_and3_4_y0(a_3, b_4, h_s_arrmul16_and3_4_y0);
  fa fa_h_s_arrmul16_fa3_4_y2(h_s_arrmul16_and3_4_y0, h_s_arrmul16_fa4_3_y2, h_s_arrmul16_fa2_4_y4, h_s_arrmul16_fa3_4_y2, h_s_arrmul16_fa3_4_y4);
  and_gate and_gate_h_s_arrmul16_and4_4_y0(a_4, b_4, h_s_arrmul16_and4_4_y0);
  fa fa_h_s_arrmul16_fa4_4_y2(h_s_arrmul16_and4_4_y0, h_s_arrmul16_fa5_3_y2, h_s_arrmul16_fa3_4_y4, h_s_arrmul16_fa4_4_y2, h_s_arrmul16_fa4_4_y4);
  and_gate and_gate_h_s_arrmul16_and5_4_y0(a_5, b_4, h_s_arrmul16_and5_4_y0);
  fa fa_h_s_arrmul16_fa5_4_y2(h_s_arrmul16_and5_4_y0, h_s_arrmul16_fa6_3_y2, h_s_arrmul16_fa4_4_y4, h_s_arrmul16_fa5_4_y2, h_s_arrmul16_fa5_4_y4);
  and_gate and_gate_h_s_arrmul16_and6_4_y0(a_6, b_4, h_s_arrmul16_and6_4_y0);
  fa fa_h_s_arrmul16_fa6_4_y2(h_s_arrmul16_and6_4_y0, h_s_arrmul16_fa7_3_y2, h_s_arrmul16_fa5_4_y4, h_s_arrmul16_fa6_4_y2, h_s_arrmul16_fa6_4_y4);
  and_gate and_gate_h_s_arrmul16_and7_4_y0(a_7, b_4, h_s_arrmul16_and7_4_y0);
  fa fa_h_s_arrmul16_fa7_4_y2(h_s_arrmul16_and7_4_y0, h_s_arrmul16_fa8_3_y2, h_s_arrmul16_fa6_4_y4, h_s_arrmul16_fa7_4_y2, h_s_arrmul16_fa7_4_y4);
  and_gate and_gate_h_s_arrmul16_and8_4_y0(a_8, b_4, h_s_arrmul16_and8_4_y0);
  fa fa_h_s_arrmul16_fa8_4_y2(h_s_arrmul16_and8_4_y0, h_s_arrmul16_fa9_3_y2, h_s_arrmul16_fa7_4_y4, h_s_arrmul16_fa8_4_y2, h_s_arrmul16_fa8_4_y4);
  and_gate and_gate_h_s_arrmul16_and9_4_y0(a_9, b_4, h_s_arrmul16_and9_4_y0);
  fa fa_h_s_arrmul16_fa9_4_y2(h_s_arrmul16_and9_4_y0, h_s_arrmul16_fa10_3_y2, h_s_arrmul16_fa8_4_y4, h_s_arrmul16_fa9_4_y2, h_s_arrmul16_fa9_4_y4);
  and_gate and_gate_h_s_arrmul16_and10_4_y0(a_10, b_4, h_s_arrmul16_and10_4_y0);
  fa fa_h_s_arrmul16_fa10_4_y2(h_s_arrmul16_and10_4_y0, h_s_arrmul16_fa11_3_y2, h_s_arrmul16_fa9_4_y4, h_s_arrmul16_fa10_4_y2, h_s_arrmul16_fa10_4_y4);
  and_gate and_gate_h_s_arrmul16_and11_4_y0(a_11, b_4, h_s_arrmul16_and11_4_y0);
  fa fa_h_s_arrmul16_fa11_4_y2(h_s_arrmul16_and11_4_y0, h_s_arrmul16_fa12_3_y2, h_s_arrmul16_fa10_4_y4, h_s_arrmul16_fa11_4_y2, h_s_arrmul16_fa11_4_y4);
  and_gate and_gate_h_s_arrmul16_and12_4_y0(a_12, b_4, h_s_arrmul16_and12_4_y0);
  fa fa_h_s_arrmul16_fa12_4_y2(h_s_arrmul16_and12_4_y0, h_s_arrmul16_fa13_3_y2, h_s_arrmul16_fa11_4_y4, h_s_arrmul16_fa12_4_y2, h_s_arrmul16_fa12_4_y4);
  and_gate and_gate_h_s_arrmul16_and13_4_y0(a_13, b_4, h_s_arrmul16_and13_4_y0);
  fa fa_h_s_arrmul16_fa13_4_y2(h_s_arrmul16_and13_4_y0, h_s_arrmul16_fa14_3_y2, h_s_arrmul16_fa12_4_y4, h_s_arrmul16_fa13_4_y2, h_s_arrmul16_fa13_4_y4);
  and_gate and_gate_h_s_arrmul16_and14_4_y0(a_14, b_4, h_s_arrmul16_and14_4_y0);
  fa fa_h_s_arrmul16_fa14_4_y2(h_s_arrmul16_and14_4_y0, h_s_arrmul16_fa15_3_y2, h_s_arrmul16_fa13_4_y4, h_s_arrmul16_fa14_4_y2, h_s_arrmul16_fa14_4_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_4_y0(a_15, b_4, h_s_arrmul16_nand15_4_y0);
  fa fa_h_s_arrmul16_fa15_4_y2(h_s_arrmul16_nand15_4_y0, h_s_arrmul16_fa15_3_y4, h_s_arrmul16_fa14_4_y4, h_s_arrmul16_fa15_4_y2, h_s_arrmul16_fa15_4_y4);
  and_gate and_gate_h_s_arrmul16_and0_5_y0(a_0, b_5, h_s_arrmul16_and0_5_y0);
  ha ha_h_s_arrmul16_ha0_5_y0(h_s_arrmul16_and0_5_y0, h_s_arrmul16_fa1_4_y2, h_s_arrmul16_ha0_5_y0, h_s_arrmul16_ha0_5_y1);
  and_gate and_gate_h_s_arrmul16_and1_5_y0(a_1, b_5, h_s_arrmul16_and1_5_y0);
  fa fa_h_s_arrmul16_fa1_5_y2(h_s_arrmul16_and1_5_y0, h_s_arrmul16_fa2_4_y2, h_s_arrmul16_ha0_5_y1, h_s_arrmul16_fa1_5_y2, h_s_arrmul16_fa1_5_y4);
  and_gate and_gate_h_s_arrmul16_and2_5_y0(a_2, b_5, h_s_arrmul16_and2_5_y0);
  fa fa_h_s_arrmul16_fa2_5_y2(h_s_arrmul16_and2_5_y0, h_s_arrmul16_fa3_4_y2, h_s_arrmul16_fa1_5_y4, h_s_arrmul16_fa2_5_y2, h_s_arrmul16_fa2_5_y4);
  and_gate and_gate_h_s_arrmul16_and3_5_y0(a_3, b_5, h_s_arrmul16_and3_5_y0);
  fa fa_h_s_arrmul16_fa3_5_y2(h_s_arrmul16_and3_5_y0, h_s_arrmul16_fa4_4_y2, h_s_arrmul16_fa2_5_y4, h_s_arrmul16_fa3_5_y2, h_s_arrmul16_fa3_5_y4);
  and_gate and_gate_h_s_arrmul16_and4_5_y0(a_4, b_5, h_s_arrmul16_and4_5_y0);
  fa fa_h_s_arrmul16_fa4_5_y2(h_s_arrmul16_and4_5_y0, h_s_arrmul16_fa5_4_y2, h_s_arrmul16_fa3_5_y4, h_s_arrmul16_fa4_5_y2, h_s_arrmul16_fa4_5_y4);
  and_gate and_gate_h_s_arrmul16_and5_5_y0(a_5, b_5, h_s_arrmul16_and5_5_y0);
  fa fa_h_s_arrmul16_fa5_5_y2(h_s_arrmul16_and5_5_y0, h_s_arrmul16_fa6_4_y2, h_s_arrmul16_fa4_5_y4, h_s_arrmul16_fa5_5_y2, h_s_arrmul16_fa5_5_y4);
  and_gate and_gate_h_s_arrmul16_and6_5_y0(a_6, b_5, h_s_arrmul16_and6_5_y0);
  fa fa_h_s_arrmul16_fa6_5_y2(h_s_arrmul16_and6_5_y0, h_s_arrmul16_fa7_4_y2, h_s_arrmul16_fa5_5_y4, h_s_arrmul16_fa6_5_y2, h_s_arrmul16_fa6_5_y4);
  and_gate and_gate_h_s_arrmul16_and7_5_y0(a_7, b_5, h_s_arrmul16_and7_5_y0);
  fa fa_h_s_arrmul16_fa7_5_y2(h_s_arrmul16_and7_5_y0, h_s_arrmul16_fa8_4_y2, h_s_arrmul16_fa6_5_y4, h_s_arrmul16_fa7_5_y2, h_s_arrmul16_fa7_5_y4);
  and_gate and_gate_h_s_arrmul16_and8_5_y0(a_8, b_5, h_s_arrmul16_and8_5_y0);
  fa fa_h_s_arrmul16_fa8_5_y2(h_s_arrmul16_and8_5_y0, h_s_arrmul16_fa9_4_y2, h_s_arrmul16_fa7_5_y4, h_s_arrmul16_fa8_5_y2, h_s_arrmul16_fa8_5_y4);
  and_gate and_gate_h_s_arrmul16_and9_5_y0(a_9, b_5, h_s_arrmul16_and9_5_y0);
  fa fa_h_s_arrmul16_fa9_5_y2(h_s_arrmul16_and9_5_y0, h_s_arrmul16_fa10_4_y2, h_s_arrmul16_fa8_5_y4, h_s_arrmul16_fa9_5_y2, h_s_arrmul16_fa9_5_y4);
  and_gate and_gate_h_s_arrmul16_and10_5_y0(a_10, b_5, h_s_arrmul16_and10_5_y0);
  fa fa_h_s_arrmul16_fa10_5_y2(h_s_arrmul16_and10_5_y0, h_s_arrmul16_fa11_4_y2, h_s_arrmul16_fa9_5_y4, h_s_arrmul16_fa10_5_y2, h_s_arrmul16_fa10_5_y4);
  and_gate and_gate_h_s_arrmul16_and11_5_y0(a_11, b_5, h_s_arrmul16_and11_5_y0);
  fa fa_h_s_arrmul16_fa11_5_y2(h_s_arrmul16_and11_5_y0, h_s_arrmul16_fa12_4_y2, h_s_arrmul16_fa10_5_y4, h_s_arrmul16_fa11_5_y2, h_s_arrmul16_fa11_5_y4);
  and_gate and_gate_h_s_arrmul16_and12_5_y0(a_12, b_5, h_s_arrmul16_and12_5_y0);
  fa fa_h_s_arrmul16_fa12_5_y2(h_s_arrmul16_and12_5_y0, h_s_arrmul16_fa13_4_y2, h_s_arrmul16_fa11_5_y4, h_s_arrmul16_fa12_5_y2, h_s_arrmul16_fa12_5_y4);
  and_gate and_gate_h_s_arrmul16_and13_5_y0(a_13, b_5, h_s_arrmul16_and13_5_y0);
  fa fa_h_s_arrmul16_fa13_5_y2(h_s_arrmul16_and13_5_y0, h_s_arrmul16_fa14_4_y2, h_s_arrmul16_fa12_5_y4, h_s_arrmul16_fa13_5_y2, h_s_arrmul16_fa13_5_y4);
  and_gate and_gate_h_s_arrmul16_and14_5_y0(a_14, b_5, h_s_arrmul16_and14_5_y0);
  fa fa_h_s_arrmul16_fa14_5_y2(h_s_arrmul16_and14_5_y0, h_s_arrmul16_fa15_4_y2, h_s_arrmul16_fa13_5_y4, h_s_arrmul16_fa14_5_y2, h_s_arrmul16_fa14_5_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_5_y0(a_15, b_5, h_s_arrmul16_nand15_5_y0);
  fa fa_h_s_arrmul16_fa15_5_y2(h_s_arrmul16_nand15_5_y0, h_s_arrmul16_fa15_4_y4, h_s_arrmul16_fa14_5_y4, h_s_arrmul16_fa15_5_y2, h_s_arrmul16_fa15_5_y4);
  and_gate and_gate_h_s_arrmul16_and0_6_y0(a_0, b_6, h_s_arrmul16_and0_6_y0);
  ha ha_h_s_arrmul16_ha0_6_y0(h_s_arrmul16_and0_6_y0, h_s_arrmul16_fa1_5_y2, h_s_arrmul16_ha0_6_y0, h_s_arrmul16_ha0_6_y1);
  and_gate and_gate_h_s_arrmul16_and1_6_y0(a_1, b_6, h_s_arrmul16_and1_6_y0);
  fa fa_h_s_arrmul16_fa1_6_y2(h_s_arrmul16_and1_6_y0, h_s_arrmul16_fa2_5_y2, h_s_arrmul16_ha0_6_y1, h_s_arrmul16_fa1_6_y2, h_s_arrmul16_fa1_6_y4);
  and_gate and_gate_h_s_arrmul16_and2_6_y0(a_2, b_6, h_s_arrmul16_and2_6_y0);
  fa fa_h_s_arrmul16_fa2_6_y2(h_s_arrmul16_and2_6_y0, h_s_arrmul16_fa3_5_y2, h_s_arrmul16_fa1_6_y4, h_s_arrmul16_fa2_6_y2, h_s_arrmul16_fa2_6_y4);
  and_gate and_gate_h_s_arrmul16_and3_6_y0(a_3, b_6, h_s_arrmul16_and3_6_y0);
  fa fa_h_s_arrmul16_fa3_6_y2(h_s_arrmul16_and3_6_y0, h_s_arrmul16_fa4_5_y2, h_s_arrmul16_fa2_6_y4, h_s_arrmul16_fa3_6_y2, h_s_arrmul16_fa3_6_y4);
  and_gate and_gate_h_s_arrmul16_and4_6_y0(a_4, b_6, h_s_arrmul16_and4_6_y0);
  fa fa_h_s_arrmul16_fa4_6_y2(h_s_arrmul16_and4_6_y0, h_s_arrmul16_fa5_5_y2, h_s_arrmul16_fa3_6_y4, h_s_arrmul16_fa4_6_y2, h_s_arrmul16_fa4_6_y4);
  and_gate and_gate_h_s_arrmul16_and5_6_y0(a_5, b_6, h_s_arrmul16_and5_6_y0);
  fa fa_h_s_arrmul16_fa5_6_y2(h_s_arrmul16_and5_6_y0, h_s_arrmul16_fa6_5_y2, h_s_arrmul16_fa4_6_y4, h_s_arrmul16_fa5_6_y2, h_s_arrmul16_fa5_6_y4);
  and_gate and_gate_h_s_arrmul16_and6_6_y0(a_6, b_6, h_s_arrmul16_and6_6_y0);
  fa fa_h_s_arrmul16_fa6_6_y2(h_s_arrmul16_and6_6_y0, h_s_arrmul16_fa7_5_y2, h_s_arrmul16_fa5_6_y4, h_s_arrmul16_fa6_6_y2, h_s_arrmul16_fa6_6_y4);
  and_gate and_gate_h_s_arrmul16_and7_6_y0(a_7, b_6, h_s_arrmul16_and7_6_y0);
  fa fa_h_s_arrmul16_fa7_6_y2(h_s_arrmul16_and7_6_y0, h_s_arrmul16_fa8_5_y2, h_s_arrmul16_fa6_6_y4, h_s_arrmul16_fa7_6_y2, h_s_arrmul16_fa7_6_y4);
  and_gate and_gate_h_s_arrmul16_and8_6_y0(a_8, b_6, h_s_arrmul16_and8_6_y0);
  fa fa_h_s_arrmul16_fa8_6_y2(h_s_arrmul16_and8_6_y0, h_s_arrmul16_fa9_5_y2, h_s_arrmul16_fa7_6_y4, h_s_arrmul16_fa8_6_y2, h_s_arrmul16_fa8_6_y4);
  and_gate and_gate_h_s_arrmul16_and9_6_y0(a_9, b_6, h_s_arrmul16_and9_6_y0);
  fa fa_h_s_arrmul16_fa9_6_y2(h_s_arrmul16_and9_6_y0, h_s_arrmul16_fa10_5_y2, h_s_arrmul16_fa8_6_y4, h_s_arrmul16_fa9_6_y2, h_s_arrmul16_fa9_6_y4);
  and_gate and_gate_h_s_arrmul16_and10_6_y0(a_10, b_6, h_s_arrmul16_and10_6_y0);
  fa fa_h_s_arrmul16_fa10_6_y2(h_s_arrmul16_and10_6_y0, h_s_arrmul16_fa11_5_y2, h_s_arrmul16_fa9_6_y4, h_s_arrmul16_fa10_6_y2, h_s_arrmul16_fa10_6_y4);
  and_gate and_gate_h_s_arrmul16_and11_6_y0(a_11, b_6, h_s_arrmul16_and11_6_y0);
  fa fa_h_s_arrmul16_fa11_6_y2(h_s_arrmul16_and11_6_y0, h_s_arrmul16_fa12_5_y2, h_s_arrmul16_fa10_6_y4, h_s_arrmul16_fa11_6_y2, h_s_arrmul16_fa11_6_y4);
  and_gate and_gate_h_s_arrmul16_and12_6_y0(a_12, b_6, h_s_arrmul16_and12_6_y0);
  fa fa_h_s_arrmul16_fa12_6_y2(h_s_arrmul16_and12_6_y0, h_s_arrmul16_fa13_5_y2, h_s_arrmul16_fa11_6_y4, h_s_arrmul16_fa12_6_y2, h_s_arrmul16_fa12_6_y4);
  and_gate and_gate_h_s_arrmul16_and13_6_y0(a_13, b_6, h_s_arrmul16_and13_6_y0);
  fa fa_h_s_arrmul16_fa13_6_y2(h_s_arrmul16_and13_6_y0, h_s_arrmul16_fa14_5_y2, h_s_arrmul16_fa12_6_y4, h_s_arrmul16_fa13_6_y2, h_s_arrmul16_fa13_6_y4);
  and_gate and_gate_h_s_arrmul16_and14_6_y0(a_14, b_6, h_s_arrmul16_and14_6_y0);
  fa fa_h_s_arrmul16_fa14_6_y2(h_s_arrmul16_and14_6_y0, h_s_arrmul16_fa15_5_y2, h_s_arrmul16_fa13_6_y4, h_s_arrmul16_fa14_6_y2, h_s_arrmul16_fa14_6_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_6_y0(a_15, b_6, h_s_arrmul16_nand15_6_y0);
  fa fa_h_s_arrmul16_fa15_6_y2(h_s_arrmul16_nand15_6_y0, h_s_arrmul16_fa15_5_y4, h_s_arrmul16_fa14_6_y4, h_s_arrmul16_fa15_6_y2, h_s_arrmul16_fa15_6_y4);
  and_gate and_gate_h_s_arrmul16_and0_7_y0(a_0, b_7, h_s_arrmul16_and0_7_y0);
  ha ha_h_s_arrmul16_ha0_7_y0(h_s_arrmul16_and0_7_y0, h_s_arrmul16_fa1_6_y2, h_s_arrmul16_ha0_7_y0, h_s_arrmul16_ha0_7_y1);
  and_gate and_gate_h_s_arrmul16_and1_7_y0(a_1, b_7, h_s_arrmul16_and1_7_y0);
  fa fa_h_s_arrmul16_fa1_7_y2(h_s_arrmul16_and1_7_y0, h_s_arrmul16_fa2_6_y2, h_s_arrmul16_ha0_7_y1, h_s_arrmul16_fa1_7_y2, h_s_arrmul16_fa1_7_y4);
  and_gate and_gate_h_s_arrmul16_and2_7_y0(a_2, b_7, h_s_arrmul16_and2_7_y0);
  fa fa_h_s_arrmul16_fa2_7_y2(h_s_arrmul16_and2_7_y0, h_s_arrmul16_fa3_6_y2, h_s_arrmul16_fa1_7_y4, h_s_arrmul16_fa2_7_y2, h_s_arrmul16_fa2_7_y4);
  and_gate and_gate_h_s_arrmul16_and3_7_y0(a_3, b_7, h_s_arrmul16_and3_7_y0);
  fa fa_h_s_arrmul16_fa3_7_y2(h_s_arrmul16_and3_7_y0, h_s_arrmul16_fa4_6_y2, h_s_arrmul16_fa2_7_y4, h_s_arrmul16_fa3_7_y2, h_s_arrmul16_fa3_7_y4);
  and_gate and_gate_h_s_arrmul16_and4_7_y0(a_4, b_7, h_s_arrmul16_and4_7_y0);
  fa fa_h_s_arrmul16_fa4_7_y2(h_s_arrmul16_and4_7_y0, h_s_arrmul16_fa5_6_y2, h_s_arrmul16_fa3_7_y4, h_s_arrmul16_fa4_7_y2, h_s_arrmul16_fa4_7_y4);
  and_gate and_gate_h_s_arrmul16_and5_7_y0(a_5, b_7, h_s_arrmul16_and5_7_y0);
  fa fa_h_s_arrmul16_fa5_7_y2(h_s_arrmul16_and5_7_y0, h_s_arrmul16_fa6_6_y2, h_s_arrmul16_fa4_7_y4, h_s_arrmul16_fa5_7_y2, h_s_arrmul16_fa5_7_y4);
  and_gate and_gate_h_s_arrmul16_and6_7_y0(a_6, b_7, h_s_arrmul16_and6_7_y0);
  fa fa_h_s_arrmul16_fa6_7_y2(h_s_arrmul16_and6_7_y0, h_s_arrmul16_fa7_6_y2, h_s_arrmul16_fa5_7_y4, h_s_arrmul16_fa6_7_y2, h_s_arrmul16_fa6_7_y4);
  and_gate and_gate_h_s_arrmul16_and7_7_y0(a_7, b_7, h_s_arrmul16_and7_7_y0);
  fa fa_h_s_arrmul16_fa7_7_y2(h_s_arrmul16_and7_7_y0, h_s_arrmul16_fa8_6_y2, h_s_arrmul16_fa6_7_y4, h_s_arrmul16_fa7_7_y2, h_s_arrmul16_fa7_7_y4);
  and_gate and_gate_h_s_arrmul16_and8_7_y0(a_8, b_7, h_s_arrmul16_and8_7_y0);
  fa fa_h_s_arrmul16_fa8_7_y2(h_s_arrmul16_and8_7_y0, h_s_arrmul16_fa9_6_y2, h_s_arrmul16_fa7_7_y4, h_s_arrmul16_fa8_7_y2, h_s_arrmul16_fa8_7_y4);
  and_gate and_gate_h_s_arrmul16_and9_7_y0(a_9, b_7, h_s_arrmul16_and9_7_y0);
  fa fa_h_s_arrmul16_fa9_7_y2(h_s_arrmul16_and9_7_y0, h_s_arrmul16_fa10_6_y2, h_s_arrmul16_fa8_7_y4, h_s_arrmul16_fa9_7_y2, h_s_arrmul16_fa9_7_y4);
  and_gate and_gate_h_s_arrmul16_and10_7_y0(a_10, b_7, h_s_arrmul16_and10_7_y0);
  fa fa_h_s_arrmul16_fa10_7_y2(h_s_arrmul16_and10_7_y0, h_s_arrmul16_fa11_6_y2, h_s_arrmul16_fa9_7_y4, h_s_arrmul16_fa10_7_y2, h_s_arrmul16_fa10_7_y4);
  and_gate and_gate_h_s_arrmul16_and11_7_y0(a_11, b_7, h_s_arrmul16_and11_7_y0);
  fa fa_h_s_arrmul16_fa11_7_y2(h_s_arrmul16_and11_7_y0, h_s_arrmul16_fa12_6_y2, h_s_arrmul16_fa10_7_y4, h_s_arrmul16_fa11_7_y2, h_s_arrmul16_fa11_7_y4);
  and_gate and_gate_h_s_arrmul16_and12_7_y0(a_12, b_7, h_s_arrmul16_and12_7_y0);
  fa fa_h_s_arrmul16_fa12_7_y2(h_s_arrmul16_and12_7_y0, h_s_arrmul16_fa13_6_y2, h_s_arrmul16_fa11_7_y4, h_s_arrmul16_fa12_7_y2, h_s_arrmul16_fa12_7_y4);
  and_gate and_gate_h_s_arrmul16_and13_7_y0(a_13, b_7, h_s_arrmul16_and13_7_y0);
  fa fa_h_s_arrmul16_fa13_7_y2(h_s_arrmul16_and13_7_y0, h_s_arrmul16_fa14_6_y2, h_s_arrmul16_fa12_7_y4, h_s_arrmul16_fa13_7_y2, h_s_arrmul16_fa13_7_y4);
  and_gate and_gate_h_s_arrmul16_and14_7_y0(a_14, b_7, h_s_arrmul16_and14_7_y0);
  fa fa_h_s_arrmul16_fa14_7_y2(h_s_arrmul16_and14_7_y0, h_s_arrmul16_fa15_6_y2, h_s_arrmul16_fa13_7_y4, h_s_arrmul16_fa14_7_y2, h_s_arrmul16_fa14_7_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_7_y0(a_15, b_7, h_s_arrmul16_nand15_7_y0);
  fa fa_h_s_arrmul16_fa15_7_y2(h_s_arrmul16_nand15_7_y0, h_s_arrmul16_fa15_6_y4, h_s_arrmul16_fa14_7_y4, h_s_arrmul16_fa15_7_y2, h_s_arrmul16_fa15_7_y4);
  and_gate and_gate_h_s_arrmul16_and0_8_y0(a_0, b_8, h_s_arrmul16_and0_8_y0);
  ha ha_h_s_arrmul16_ha0_8_y0(h_s_arrmul16_and0_8_y0, h_s_arrmul16_fa1_7_y2, h_s_arrmul16_ha0_8_y0, h_s_arrmul16_ha0_8_y1);
  and_gate and_gate_h_s_arrmul16_and1_8_y0(a_1, b_8, h_s_arrmul16_and1_8_y0);
  fa fa_h_s_arrmul16_fa1_8_y2(h_s_arrmul16_and1_8_y0, h_s_arrmul16_fa2_7_y2, h_s_arrmul16_ha0_8_y1, h_s_arrmul16_fa1_8_y2, h_s_arrmul16_fa1_8_y4);
  and_gate and_gate_h_s_arrmul16_and2_8_y0(a_2, b_8, h_s_arrmul16_and2_8_y0);
  fa fa_h_s_arrmul16_fa2_8_y2(h_s_arrmul16_and2_8_y0, h_s_arrmul16_fa3_7_y2, h_s_arrmul16_fa1_8_y4, h_s_arrmul16_fa2_8_y2, h_s_arrmul16_fa2_8_y4);
  and_gate and_gate_h_s_arrmul16_and3_8_y0(a_3, b_8, h_s_arrmul16_and3_8_y0);
  fa fa_h_s_arrmul16_fa3_8_y2(h_s_arrmul16_and3_8_y0, h_s_arrmul16_fa4_7_y2, h_s_arrmul16_fa2_8_y4, h_s_arrmul16_fa3_8_y2, h_s_arrmul16_fa3_8_y4);
  and_gate and_gate_h_s_arrmul16_and4_8_y0(a_4, b_8, h_s_arrmul16_and4_8_y0);
  fa fa_h_s_arrmul16_fa4_8_y2(h_s_arrmul16_and4_8_y0, h_s_arrmul16_fa5_7_y2, h_s_arrmul16_fa3_8_y4, h_s_arrmul16_fa4_8_y2, h_s_arrmul16_fa4_8_y4);
  and_gate and_gate_h_s_arrmul16_and5_8_y0(a_5, b_8, h_s_arrmul16_and5_8_y0);
  fa fa_h_s_arrmul16_fa5_8_y2(h_s_arrmul16_and5_8_y0, h_s_arrmul16_fa6_7_y2, h_s_arrmul16_fa4_8_y4, h_s_arrmul16_fa5_8_y2, h_s_arrmul16_fa5_8_y4);
  and_gate and_gate_h_s_arrmul16_and6_8_y0(a_6, b_8, h_s_arrmul16_and6_8_y0);
  fa fa_h_s_arrmul16_fa6_8_y2(h_s_arrmul16_and6_8_y0, h_s_arrmul16_fa7_7_y2, h_s_arrmul16_fa5_8_y4, h_s_arrmul16_fa6_8_y2, h_s_arrmul16_fa6_8_y4);
  and_gate and_gate_h_s_arrmul16_and7_8_y0(a_7, b_8, h_s_arrmul16_and7_8_y0);
  fa fa_h_s_arrmul16_fa7_8_y2(h_s_arrmul16_and7_8_y0, h_s_arrmul16_fa8_7_y2, h_s_arrmul16_fa6_8_y4, h_s_arrmul16_fa7_8_y2, h_s_arrmul16_fa7_8_y4);
  and_gate and_gate_h_s_arrmul16_and8_8_y0(a_8, b_8, h_s_arrmul16_and8_8_y0);
  fa fa_h_s_arrmul16_fa8_8_y2(h_s_arrmul16_and8_8_y0, h_s_arrmul16_fa9_7_y2, h_s_arrmul16_fa7_8_y4, h_s_arrmul16_fa8_8_y2, h_s_arrmul16_fa8_8_y4);
  and_gate and_gate_h_s_arrmul16_and9_8_y0(a_9, b_8, h_s_arrmul16_and9_8_y0);
  fa fa_h_s_arrmul16_fa9_8_y2(h_s_arrmul16_and9_8_y0, h_s_arrmul16_fa10_7_y2, h_s_arrmul16_fa8_8_y4, h_s_arrmul16_fa9_8_y2, h_s_arrmul16_fa9_8_y4);
  and_gate and_gate_h_s_arrmul16_and10_8_y0(a_10, b_8, h_s_arrmul16_and10_8_y0);
  fa fa_h_s_arrmul16_fa10_8_y2(h_s_arrmul16_and10_8_y0, h_s_arrmul16_fa11_7_y2, h_s_arrmul16_fa9_8_y4, h_s_arrmul16_fa10_8_y2, h_s_arrmul16_fa10_8_y4);
  and_gate and_gate_h_s_arrmul16_and11_8_y0(a_11, b_8, h_s_arrmul16_and11_8_y0);
  fa fa_h_s_arrmul16_fa11_8_y2(h_s_arrmul16_and11_8_y0, h_s_arrmul16_fa12_7_y2, h_s_arrmul16_fa10_8_y4, h_s_arrmul16_fa11_8_y2, h_s_arrmul16_fa11_8_y4);
  and_gate and_gate_h_s_arrmul16_and12_8_y0(a_12, b_8, h_s_arrmul16_and12_8_y0);
  fa fa_h_s_arrmul16_fa12_8_y2(h_s_arrmul16_and12_8_y0, h_s_arrmul16_fa13_7_y2, h_s_arrmul16_fa11_8_y4, h_s_arrmul16_fa12_8_y2, h_s_arrmul16_fa12_8_y4);
  and_gate and_gate_h_s_arrmul16_and13_8_y0(a_13, b_8, h_s_arrmul16_and13_8_y0);
  fa fa_h_s_arrmul16_fa13_8_y2(h_s_arrmul16_and13_8_y0, h_s_arrmul16_fa14_7_y2, h_s_arrmul16_fa12_8_y4, h_s_arrmul16_fa13_8_y2, h_s_arrmul16_fa13_8_y4);
  and_gate and_gate_h_s_arrmul16_and14_8_y0(a_14, b_8, h_s_arrmul16_and14_8_y0);
  fa fa_h_s_arrmul16_fa14_8_y2(h_s_arrmul16_and14_8_y0, h_s_arrmul16_fa15_7_y2, h_s_arrmul16_fa13_8_y4, h_s_arrmul16_fa14_8_y2, h_s_arrmul16_fa14_8_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_8_y0(a_15, b_8, h_s_arrmul16_nand15_8_y0);
  fa fa_h_s_arrmul16_fa15_8_y2(h_s_arrmul16_nand15_8_y0, h_s_arrmul16_fa15_7_y4, h_s_arrmul16_fa14_8_y4, h_s_arrmul16_fa15_8_y2, h_s_arrmul16_fa15_8_y4);
  and_gate and_gate_h_s_arrmul16_and0_9_y0(a_0, b_9, h_s_arrmul16_and0_9_y0);
  ha ha_h_s_arrmul16_ha0_9_y0(h_s_arrmul16_and0_9_y0, h_s_arrmul16_fa1_8_y2, h_s_arrmul16_ha0_9_y0, h_s_arrmul16_ha0_9_y1);
  and_gate and_gate_h_s_arrmul16_and1_9_y0(a_1, b_9, h_s_arrmul16_and1_9_y0);
  fa fa_h_s_arrmul16_fa1_9_y2(h_s_arrmul16_and1_9_y0, h_s_arrmul16_fa2_8_y2, h_s_arrmul16_ha0_9_y1, h_s_arrmul16_fa1_9_y2, h_s_arrmul16_fa1_9_y4);
  and_gate and_gate_h_s_arrmul16_and2_9_y0(a_2, b_9, h_s_arrmul16_and2_9_y0);
  fa fa_h_s_arrmul16_fa2_9_y2(h_s_arrmul16_and2_9_y0, h_s_arrmul16_fa3_8_y2, h_s_arrmul16_fa1_9_y4, h_s_arrmul16_fa2_9_y2, h_s_arrmul16_fa2_9_y4);
  and_gate and_gate_h_s_arrmul16_and3_9_y0(a_3, b_9, h_s_arrmul16_and3_9_y0);
  fa fa_h_s_arrmul16_fa3_9_y2(h_s_arrmul16_and3_9_y0, h_s_arrmul16_fa4_8_y2, h_s_arrmul16_fa2_9_y4, h_s_arrmul16_fa3_9_y2, h_s_arrmul16_fa3_9_y4);
  and_gate and_gate_h_s_arrmul16_and4_9_y0(a_4, b_9, h_s_arrmul16_and4_9_y0);
  fa fa_h_s_arrmul16_fa4_9_y2(h_s_arrmul16_and4_9_y0, h_s_arrmul16_fa5_8_y2, h_s_arrmul16_fa3_9_y4, h_s_arrmul16_fa4_9_y2, h_s_arrmul16_fa4_9_y4);
  and_gate and_gate_h_s_arrmul16_and5_9_y0(a_5, b_9, h_s_arrmul16_and5_9_y0);
  fa fa_h_s_arrmul16_fa5_9_y2(h_s_arrmul16_and5_9_y0, h_s_arrmul16_fa6_8_y2, h_s_arrmul16_fa4_9_y4, h_s_arrmul16_fa5_9_y2, h_s_arrmul16_fa5_9_y4);
  and_gate and_gate_h_s_arrmul16_and6_9_y0(a_6, b_9, h_s_arrmul16_and6_9_y0);
  fa fa_h_s_arrmul16_fa6_9_y2(h_s_arrmul16_and6_9_y0, h_s_arrmul16_fa7_8_y2, h_s_arrmul16_fa5_9_y4, h_s_arrmul16_fa6_9_y2, h_s_arrmul16_fa6_9_y4);
  and_gate and_gate_h_s_arrmul16_and7_9_y0(a_7, b_9, h_s_arrmul16_and7_9_y0);
  fa fa_h_s_arrmul16_fa7_9_y2(h_s_arrmul16_and7_9_y0, h_s_arrmul16_fa8_8_y2, h_s_arrmul16_fa6_9_y4, h_s_arrmul16_fa7_9_y2, h_s_arrmul16_fa7_9_y4);
  and_gate and_gate_h_s_arrmul16_and8_9_y0(a_8, b_9, h_s_arrmul16_and8_9_y0);
  fa fa_h_s_arrmul16_fa8_9_y2(h_s_arrmul16_and8_9_y0, h_s_arrmul16_fa9_8_y2, h_s_arrmul16_fa7_9_y4, h_s_arrmul16_fa8_9_y2, h_s_arrmul16_fa8_9_y4);
  and_gate and_gate_h_s_arrmul16_and9_9_y0(a_9, b_9, h_s_arrmul16_and9_9_y0);
  fa fa_h_s_arrmul16_fa9_9_y2(h_s_arrmul16_and9_9_y0, h_s_arrmul16_fa10_8_y2, h_s_arrmul16_fa8_9_y4, h_s_arrmul16_fa9_9_y2, h_s_arrmul16_fa9_9_y4);
  and_gate and_gate_h_s_arrmul16_and10_9_y0(a_10, b_9, h_s_arrmul16_and10_9_y0);
  fa fa_h_s_arrmul16_fa10_9_y2(h_s_arrmul16_and10_9_y0, h_s_arrmul16_fa11_8_y2, h_s_arrmul16_fa9_9_y4, h_s_arrmul16_fa10_9_y2, h_s_arrmul16_fa10_9_y4);
  and_gate and_gate_h_s_arrmul16_and11_9_y0(a_11, b_9, h_s_arrmul16_and11_9_y0);
  fa fa_h_s_arrmul16_fa11_9_y2(h_s_arrmul16_and11_9_y0, h_s_arrmul16_fa12_8_y2, h_s_arrmul16_fa10_9_y4, h_s_arrmul16_fa11_9_y2, h_s_arrmul16_fa11_9_y4);
  and_gate and_gate_h_s_arrmul16_and12_9_y0(a_12, b_9, h_s_arrmul16_and12_9_y0);
  fa fa_h_s_arrmul16_fa12_9_y2(h_s_arrmul16_and12_9_y0, h_s_arrmul16_fa13_8_y2, h_s_arrmul16_fa11_9_y4, h_s_arrmul16_fa12_9_y2, h_s_arrmul16_fa12_9_y4);
  and_gate and_gate_h_s_arrmul16_and13_9_y0(a_13, b_9, h_s_arrmul16_and13_9_y0);
  fa fa_h_s_arrmul16_fa13_9_y2(h_s_arrmul16_and13_9_y0, h_s_arrmul16_fa14_8_y2, h_s_arrmul16_fa12_9_y4, h_s_arrmul16_fa13_9_y2, h_s_arrmul16_fa13_9_y4);
  and_gate and_gate_h_s_arrmul16_and14_9_y0(a_14, b_9, h_s_arrmul16_and14_9_y0);
  fa fa_h_s_arrmul16_fa14_9_y2(h_s_arrmul16_and14_9_y0, h_s_arrmul16_fa15_8_y2, h_s_arrmul16_fa13_9_y4, h_s_arrmul16_fa14_9_y2, h_s_arrmul16_fa14_9_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_9_y0(a_15, b_9, h_s_arrmul16_nand15_9_y0);
  fa fa_h_s_arrmul16_fa15_9_y2(h_s_arrmul16_nand15_9_y0, h_s_arrmul16_fa15_8_y4, h_s_arrmul16_fa14_9_y4, h_s_arrmul16_fa15_9_y2, h_s_arrmul16_fa15_9_y4);
  and_gate and_gate_h_s_arrmul16_and0_10_y0(a_0, b_10, h_s_arrmul16_and0_10_y0);
  ha ha_h_s_arrmul16_ha0_10_y0(h_s_arrmul16_and0_10_y0, h_s_arrmul16_fa1_9_y2, h_s_arrmul16_ha0_10_y0, h_s_arrmul16_ha0_10_y1);
  and_gate and_gate_h_s_arrmul16_and1_10_y0(a_1, b_10, h_s_arrmul16_and1_10_y0);
  fa fa_h_s_arrmul16_fa1_10_y2(h_s_arrmul16_and1_10_y0, h_s_arrmul16_fa2_9_y2, h_s_arrmul16_ha0_10_y1, h_s_arrmul16_fa1_10_y2, h_s_arrmul16_fa1_10_y4);
  and_gate and_gate_h_s_arrmul16_and2_10_y0(a_2, b_10, h_s_arrmul16_and2_10_y0);
  fa fa_h_s_arrmul16_fa2_10_y2(h_s_arrmul16_and2_10_y0, h_s_arrmul16_fa3_9_y2, h_s_arrmul16_fa1_10_y4, h_s_arrmul16_fa2_10_y2, h_s_arrmul16_fa2_10_y4);
  and_gate and_gate_h_s_arrmul16_and3_10_y0(a_3, b_10, h_s_arrmul16_and3_10_y0);
  fa fa_h_s_arrmul16_fa3_10_y2(h_s_arrmul16_and3_10_y0, h_s_arrmul16_fa4_9_y2, h_s_arrmul16_fa2_10_y4, h_s_arrmul16_fa3_10_y2, h_s_arrmul16_fa3_10_y4);
  and_gate and_gate_h_s_arrmul16_and4_10_y0(a_4, b_10, h_s_arrmul16_and4_10_y0);
  fa fa_h_s_arrmul16_fa4_10_y2(h_s_arrmul16_and4_10_y0, h_s_arrmul16_fa5_9_y2, h_s_arrmul16_fa3_10_y4, h_s_arrmul16_fa4_10_y2, h_s_arrmul16_fa4_10_y4);
  and_gate and_gate_h_s_arrmul16_and5_10_y0(a_5, b_10, h_s_arrmul16_and5_10_y0);
  fa fa_h_s_arrmul16_fa5_10_y2(h_s_arrmul16_and5_10_y0, h_s_arrmul16_fa6_9_y2, h_s_arrmul16_fa4_10_y4, h_s_arrmul16_fa5_10_y2, h_s_arrmul16_fa5_10_y4);
  and_gate and_gate_h_s_arrmul16_and6_10_y0(a_6, b_10, h_s_arrmul16_and6_10_y0);
  fa fa_h_s_arrmul16_fa6_10_y2(h_s_arrmul16_and6_10_y0, h_s_arrmul16_fa7_9_y2, h_s_arrmul16_fa5_10_y4, h_s_arrmul16_fa6_10_y2, h_s_arrmul16_fa6_10_y4);
  and_gate and_gate_h_s_arrmul16_and7_10_y0(a_7, b_10, h_s_arrmul16_and7_10_y0);
  fa fa_h_s_arrmul16_fa7_10_y2(h_s_arrmul16_and7_10_y0, h_s_arrmul16_fa8_9_y2, h_s_arrmul16_fa6_10_y4, h_s_arrmul16_fa7_10_y2, h_s_arrmul16_fa7_10_y4);
  and_gate and_gate_h_s_arrmul16_and8_10_y0(a_8, b_10, h_s_arrmul16_and8_10_y0);
  fa fa_h_s_arrmul16_fa8_10_y2(h_s_arrmul16_and8_10_y0, h_s_arrmul16_fa9_9_y2, h_s_arrmul16_fa7_10_y4, h_s_arrmul16_fa8_10_y2, h_s_arrmul16_fa8_10_y4);
  and_gate and_gate_h_s_arrmul16_and9_10_y0(a_9, b_10, h_s_arrmul16_and9_10_y0);
  fa fa_h_s_arrmul16_fa9_10_y2(h_s_arrmul16_and9_10_y0, h_s_arrmul16_fa10_9_y2, h_s_arrmul16_fa8_10_y4, h_s_arrmul16_fa9_10_y2, h_s_arrmul16_fa9_10_y4);
  and_gate and_gate_h_s_arrmul16_and10_10_y0(a_10, b_10, h_s_arrmul16_and10_10_y0);
  fa fa_h_s_arrmul16_fa10_10_y2(h_s_arrmul16_and10_10_y0, h_s_arrmul16_fa11_9_y2, h_s_arrmul16_fa9_10_y4, h_s_arrmul16_fa10_10_y2, h_s_arrmul16_fa10_10_y4);
  and_gate and_gate_h_s_arrmul16_and11_10_y0(a_11, b_10, h_s_arrmul16_and11_10_y0);
  fa fa_h_s_arrmul16_fa11_10_y2(h_s_arrmul16_and11_10_y0, h_s_arrmul16_fa12_9_y2, h_s_arrmul16_fa10_10_y4, h_s_arrmul16_fa11_10_y2, h_s_arrmul16_fa11_10_y4);
  and_gate and_gate_h_s_arrmul16_and12_10_y0(a_12, b_10, h_s_arrmul16_and12_10_y0);
  fa fa_h_s_arrmul16_fa12_10_y2(h_s_arrmul16_and12_10_y0, h_s_arrmul16_fa13_9_y2, h_s_arrmul16_fa11_10_y4, h_s_arrmul16_fa12_10_y2, h_s_arrmul16_fa12_10_y4);
  and_gate and_gate_h_s_arrmul16_and13_10_y0(a_13, b_10, h_s_arrmul16_and13_10_y0);
  fa fa_h_s_arrmul16_fa13_10_y2(h_s_arrmul16_and13_10_y0, h_s_arrmul16_fa14_9_y2, h_s_arrmul16_fa12_10_y4, h_s_arrmul16_fa13_10_y2, h_s_arrmul16_fa13_10_y4);
  and_gate and_gate_h_s_arrmul16_and14_10_y0(a_14, b_10, h_s_arrmul16_and14_10_y0);
  fa fa_h_s_arrmul16_fa14_10_y2(h_s_arrmul16_and14_10_y0, h_s_arrmul16_fa15_9_y2, h_s_arrmul16_fa13_10_y4, h_s_arrmul16_fa14_10_y2, h_s_arrmul16_fa14_10_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_10_y0(a_15, b_10, h_s_arrmul16_nand15_10_y0);
  fa fa_h_s_arrmul16_fa15_10_y2(h_s_arrmul16_nand15_10_y0, h_s_arrmul16_fa15_9_y4, h_s_arrmul16_fa14_10_y4, h_s_arrmul16_fa15_10_y2, h_s_arrmul16_fa15_10_y4);
  and_gate and_gate_h_s_arrmul16_and0_11_y0(a_0, b_11, h_s_arrmul16_and0_11_y0);
  ha ha_h_s_arrmul16_ha0_11_y0(h_s_arrmul16_and0_11_y0, h_s_arrmul16_fa1_10_y2, h_s_arrmul16_ha0_11_y0, h_s_arrmul16_ha0_11_y1);
  and_gate and_gate_h_s_arrmul16_and1_11_y0(a_1, b_11, h_s_arrmul16_and1_11_y0);
  fa fa_h_s_arrmul16_fa1_11_y2(h_s_arrmul16_and1_11_y0, h_s_arrmul16_fa2_10_y2, h_s_arrmul16_ha0_11_y1, h_s_arrmul16_fa1_11_y2, h_s_arrmul16_fa1_11_y4);
  and_gate and_gate_h_s_arrmul16_and2_11_y0(a_2, b_11, h_s_arrmul16_and2_11_y0);
  fa fa_h_s_arrmul16_fa2_11_y2(h_s_arrmul16_and2_11_y0, h_s_arrmul16_fa3_10_y2, h_s_arrmul16_fa1_11_y4, h_s_arrmul16_fa2_11_y2, h_s_arrmul16_fa2_11_y4);
  and_gate and_gate_h_s_arrmul16_and3_11_y0(a_3, b_11, h_s_arrmul16_and3_11_y0);
  fa fa_h_s_arrmul16_fa3_11_y2(h_s_arrmul16_and3_11_y0, h_s_arrmul16_fa4_10_y2, h_s_arrmul16_fa2_11_y4, h_s_arrmul16_fa3_11_y2, h_s_arrmul16_fa3_11_y4);
  and_gate and_gate_h_s_arrmul16_and4_11_y0(a_4, b_11, h_s_arrmul16_and4_11_y0);
  fa fa_h_s_arrmul16_fa4_11_y2(h_s_arrmul16_and4_11_y0, h_s_arrmul16_fa5_10_y2, h_s_arrmul16_fa3_11_y4, h_s_arrmul16_fa4_11_y2, h_s_arrmul16_fa4_11_y4);
  and_gate and_gate_h_s_arrmul16_and5_11_y0(a_5, b_11, h_s_arrmul16_and5_11_y0);
  fa fa_h_s_arrmul16_fa5_11_y2(h_s_arrmul16_and5_11_y0, h_s_arrmul16_fa6_10_y2, h_s_arrmul16_fa4_11_y4, h_s_arrmul16_fa5_11_y2, h_s_arrmul16_fa5_11_y4);
  and_gate and_gate_h_s_arrmul16_and6_11_y0(a_6, b_11, h_s_arrmul16_and6_11_y0);
  fa fa_h_s_arrmul16_fa6_11_y2(h_s_arrmul16_and6_11_y0, h_s_arrmul16_fa7_10_y2, h_s_arrmul16_fa5_11_y4, h_s_arrmul16_fa6_11_y2, h_s_arrmul16_fa6_11_y4);
  and_gate and_gate_h_s_arrmul16_and7_11_y0(a_7, b_11, h_s_arrmul16_and7_11_y0);
  fa fa_h_s_arrmul16_fa7_11_y2(h_s_arrmul16_and7_11_y0, h_s_arrmul16_fa8_10_y2, h_s_arrmul16_fa6_11_y4, h_s_arrmul16_fa7_11_y2, h_s_arrmul16_fa7_11_y4);
  and_gate and_gate_h_s_arrmul16_and8_11_y0(a_8, b_11, h_s_arrmul16_and8_11_y0);
  fa fa_h_s_arrmul16_fa8_11_y2(h_s_arrmul16_and8_11_y0, h_s_arrmul16_fa9_10_y2, h_s_arrmul16_fa7_11_y4, h_s_arrmul16_fa8_11_y2, h_s_arrmul16_fa8_11_y4);
  and_gate and_gate_h_s_arrmul16_and9_11_y0(a_9, b_11, h_s_arrmul16_and9_11_y0);
  fa fa_h_s_arrmul16_fa9_11_y2(h_s_arrmul16_and9_11_y0, h_s_arrmul16_fa10_10_y2, h_s_arrmul16_fa8_11_y4, h_s_arrmul16_fa9_11_y2, h_s_arrmul16_fa9_11_y4);
  and_gate and_gate_h_s_arrmul16_and10_11_y0(a_10, b_11, h_s_arrmul16_and10_11_y0);
  fa fa_h_s_arrmul16_fa10_11_y2(h_s_arrmul16_and10_11_y0, h_s_arrmul16_fa11_10_y2, h_s_arrmul16_fa9_11_y4, h_s_arrmul16_fa10_11_y2, h_s_arrmul16_fa10_11_y4);
  and_gate and_gate_h_s_arrmul16_and11_11_y0(a_11, b_11, h_s_arrmul16_and11_11_y0);
  fa fa_h_s_arrmul16_fa11_11_y2(h_s_arrmul16_and11_11_y0, h_s_arrmul16_fa12_10_y2, h_s_arrmul16_fa10_11_y4, h_s_arrmul16_fa11_11_y2, h_s_arrmul16_fa11_11_y4);
  and_gate and_gate_h_s_arrmul16_and12_11_y0(a_12, b_11, h_s_arrmul16_and12_11_y0);
  fa fa_h_s_arrmul16_fa12_11_y2(h_s_arrmul16_and12_11_y0, h_s_arrmul16_fa13_10_y2, h_s_arrmul16_fa11_11_y4, h_s_arrmul16_fa12_11_y2, h_s_arrmul16_fa12_11_y4);
  and_gate and_gate_h_s_arrmul16_and13_11_y0(a_13, b_11, h_s_arrmul16_and13_11_y0);
  fa fa_h_s_arrmul16_fa13_11_y2(h_s_arrmul16_and13_11_y0, h_s_arrmul16_fa14_10_y2, h_s_arrmul16_fa12_11_y4, h_s_arrmul16_fa13_11_y2, h_s_arrmul16_fa13_11_y4);
  and_gate and_gate_h_s_arrmul16_and14_11_y0(a_14, b_11, h_s_arrmul16_and14_11_y0);
  fa fa_h_s_arrmul16_fa14_11_y2(h_s_arrmul16_and14_11_y0, h_s_arrmul16_fa15_10_y2, h_s_arrmul16_fa13_11_y4, h_s_arrmul16_fa14_11_y2, h_s_arrmul16_fa14_11_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_11_y0(a_15, b_11, h_s_arrmul16_nand15_11_y0);
  fa fa_h_s_arrmul16_fa15_11_y2(h_s_arrmul16_nand15_11_y0, h_s_arrmul16_fa15_10_y4, h_s_arrmul16_fa14_11_y4, h_s_arrmul16_fa15_11_y2, h_s_arrmul16_fa15_11_y4);
  and_gate and_gate_h_s_arrmul16_and0_12_y0(a_0, b_12, h_s_arrmul16_and0_12_y0);
  ha ha_h_s_arrmul16_ha0_12_y0(h_s_arrmul16_and0_12_y0, h_s_arrmul16_fa1_11_y2, h_s_arrmul16_ha0_12_y0, h_s_arrmul16_ha0_12_y1);
  and_gate and_gate_h_s_arrmul16_and1_12_y0(a_1, b_12, h_s_arrmul16_and1_12_y0);
  fa fa_h_s_arrmul16_fa1_12_y2(h_s_arrmul16_and1_12_y0, h_s_arrmul16_fa2_11_y2, h_s_arrmul16_ha0_12_y1, h_s_arrmul16_fa1_12_y2, h_s_arrmul16_fa1_12_y4);
  and_gate and_gate_h_s_arrmul16_and2_12_y0(a_2, b_12, h_s_arrmul16_and2_12_y0);
  fa fa_h_s_arrmul16_fa2_12_y2(h_s_arrmul16_and2_12_y0, h_s_arrmul16_fa3_11_y2, h_s_arrmul16_fa1_12_y4, h_s_arrmul16_fa2_12_y2, h_s_arrmul16_fa2_12_y4);
  and_gate and_gate_h_s_arrmul16_and3_12_y0(a_3, b_12, h_s_arrmul16_and3_12_y0);
  fa fa_h_s_arrmul16_fa3_12_y2(h_s_arrmul16_and3_12_y0, h_s_arrmul16_fa4_11_y2, h_s_arrmul16_fa2_12_y4, h_s_arrmul16_fa3_12_y2, h_s_arrmul16_fa3_12_y4);
  and_gate and_gate_h_s_arrmul16_and4_12_y0(a_4, b_12, h_s_arrmul16_and4_12_y0);
  fa fa_h_s_arrmul16_fa4_12_y2(h_s_arrmul16_and4_12_y0, h_s_arrmul16_fa5_11_y2, h_s_arrmul16_fa3_12_y4, h_s_arrmul16_fa4_12_y2, h_s_arrmul16_fa4_12_y4);
  and_gate and_gate_h_s_arrmul16_and5_12_y0(a_5, b_12, h_s_arrmul16_and5_12_y0);
  fa fa_h_s_arrmul16_fa5_12_y2(h_s_arrmul16_and5_12_y0, h_s_arrmul16_fa6_11_y2, h_s_arrmul16_fa4_12_y4, h_s_arrmul16_fa5_12_y2, h_s_arrmul16_fa5_12_y4);
  and_gate and_gate_h_s_arrmul16_and6_12_y0(a_6, b_12, h_s_arrmul16_and6_12_y0);
  fa fa_h_s_arrmul16_fa6_12_y2(h_s_arrmul16_and6_12_y0, h_s_arrmul16_fa7_11_y2, h_s_arrmul16_fa5_12_y4, h_s_arrmul16_fa6_12_y2, h_s_arrmul16_fa6_12_y4);
  and_gate and_gate_h_s_arrmul16_and7_12_y0(a_7, b_12, h_s_arrmul16_and7_12_y0);
  fa fa_h_s_arrmul16_fa7_12_y2(h_s_arrmul16_and7_12_y0, h_s_arrmul16_fa8_11_y2, h_s_arrmul16_fa6_12_y4, h_s_arrmul16_fa7_12_y2, h_s_arrmul16_fa7_12_y4);
  and_gate and_gate_h_s_arrmul16_and8_12_y0(a_8, b_12, h_s_arrmul16_and8_12_y0);
  fa fa_h_s_arrmul16_fa8_12_y2(h_s_arrmul16_and8_12_y0, h_s_arrmul16_fa9_11_y2, h_s_arrmul16_fa7_12_y4, h_s_arrmul16_fa8_12_y2, h_s_arrmul16_fa8_12_y4);
  and_gate and_gate_h_s_arrmul16_and9_12_y0(a_9, b_12, h_s_arrmul16_and9_12_y0);
  fa fa_h_s_arrmul16_fa9_12_y2(h_s_arrmul16_and9_12_y0, h_s_arrmul16_fa10_11_y2, h_s_arrmul16_fa8_12_y4, h_s_arrmul16_fa9_12_y2, h_s_arrmul16_fa9_12_y4);
  and_gate and_gate_h_s_arrmul16_and10_12_y0(a_10, b_12, h_s_arrmul16_and10_12_y0);
  fa fa_h_s_arrmul16_fa10_12_y2(h_s_arrmul16_and10_12_y0, h_s_arrmul16_fa11_11_y2, h_s_arrmul16_fa9_12_y4, h_s_arrmul16_fa10_12_y2, h_s_arrmul16_fa10_12_y4);
  and_gate and_gate_h_s_arrmul16_and11_12_y0(a_11, b_12, h_s_arrmul16_and11_12_y0);
  fa fa_h_s_arrmul16_fa11_12_y2(h_s_arrmul16_and11_12_y0, h_s_arrmul16_fa12_11_y2, h_s_arrmul16_fa10_12_y4, h_s_arrmul16_fa11_12_y2, h_s_arrmul16_fa11_12_y4);
  and_gate and_gate_h_s_arrmul16_and12_12_y0(a_12, b_12, h_s_arrmul16_and12_12_y0);
  fa fa_h_s_arrmul16_fa12_12_y2(h_s_arrmul16_and12_12_y0, h_s_arrmul16_fa13_11_y2, h_s_arrmul16_fa11_12_y4, h_s_arrmul16_fa12_12_y2, h_s_arrmul16_fa12_12_y4);
  and_gate and_gate_h_s_arrmul16_and13_12_y0(a_13, b_12, h_s_arrmul16_and13_12_y0);
  fa fa_h_s_arrmul16_fa13_12_y2(h_s_arrmul16_and13_12_y0, h_s_arrmul16_fa14_11_y2, h_s_arrmul16_fa12_12_y4, h_s_arrmul16_fa13_12_y2, h_s_arrmul16_fa13_12_y4);
  and_gate and_gate_h_s_arrmul16_and14_12_y0(a_14, b_12, h_s_arrmul16_and14_12_y0);
  fa fa_h_s_arrmul16_fa14_12_y2(h_s_arrmul16_and14_12_y0, h_s_arrmul16_fa15_11_y2, h_s_arrmul16_fa13_12_y4, h_s_arrmul16_fa14_12_y2, h_s_arrmul16_fa14_12_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_12_y0(a_15, b_12, h_s_arrmul16_nand15_12_y0);
  fa fa_h_s_arrmul16_fa15_12_y2(h_s_arrmul16_nand15_12_y0, h_s_arrmul16_fa15_11_y4, h_s_arrmul16_fa14_12_y4, h_s_arrmul16_fa15_12_y2, h_s_arrmul16_fa15_12_y4);
  and_gate and_gate_h_s_arrmul16_and0_13_y0(a_0, b_13, h_s_arrmul16_and0_13_y0);
  ha ha_h_s_arrmul16_ha0_13_y0(h_s_arrmul16_and0_13_y0, h_s_arrmul16_fa1_12_y2, h_s_arrmul16_ha0_13_y0, h_s_arrmul16_ha0_13_y1);
  and_gate and_gate_h_s_arrmul16_and1_13_y0(a_1, b_13, h_s_arrmul16_and1_13_y0);
  fa fa_h_s_arrmul16_fa1_13_y2(h_s_arrmul16_and1_13_y0, h_s_arrmul16_fa2_12_y2, h_s_arrmul16_ha0_13_y1, h_s_arrmul16_fa1_13_y2, h_s_arrmul16_fa1_13_y4);
  and_gate and_gate_h_s_arrmul16_and2_13_y0(a_2, b_13, h_s_arrmul16_and2_13_y0);
  fa fa_h_s_arrmul16_fa2_13_y2(h_s_arrmul16_and2_13_y0, h_s_arrmul16_fa3_12_y2, h_s_arrmul16_fa1_13_y4, h_s_arrmul16_fa2_13_y2, h_s_arrmul16_fa2_13_y4);
  and_gate and_gate_h_s_arrmul16_and3_13_y0(a_3, b_13, h_s_arrmul16_and3_13_y0);
  fa fa_h_s_arrmul16_fa3_13_y2(h_s_arrmul16_and3_13_y0, h_s_arrmul16_fa4_12_y2, h_s_arrmul16_fa2_13_y4, h_s_arrmul16_fa3_13_y2, h_s_arrmul16_fa3_13_y4);
  and_gate and_gate_h_s_arrmul16_and4_13_y0(a_4, b_13, h_s_arrmul16_and4_13_y0);
  fa fa_h_s_arrmul16_fa4_13_y2(h_s_arrmul16_and4_13_y0, h_s_arrmul16_fa5_12_y2, h_s_arrmul16_fa3_13_y4, h_s_arrmul16_fa4_13_y2, h_s_arrmul16_fa4_13_y4);
  and_gate and_gate_h_s_arrmul16_and5_13_y0(a_5, b_13, h_s_arrmul16_and5_13_y0);
  fa fa_h_s_arrmul16_fa5_13_y2(h_s_arrmul16_and5_13_y0, h_s_arrmul16_fa6_12_y2, h_s_arrmul16_fa4_13_y4, h_s_arrmul16_fa5_13_y2, h_s_arrmul16_fa5_13_y4);
  and_gate and_gate_h_s_arrmul16_and6_13_y0(a_6, b_13, h_s_arrmul16_and6_13_y0);
  fa fa_h_s_arrmul16_fa6_13_y2(h_s_arrmul16_and6_13_y0, h_s_arrmul16_fa7_12_y2, h_s_arrmul16_fa5_13_y4, h_s_arrmul16_fa6_13_y2, h_s_arrmul16_fa6_13_y4);
  and_gate and_gate_h_s_arrmul16_and7_13_y0(a_7, b_13, h_s_arrmul16_and7_13_y0);
  fa fa_h_s_arrmul16_fa7_13_y2(h_s_arrmul16_and7_13_y0, h_s_arrmul16_fa8_12_y2, h_s_arrmul16_fa6_13_y4, h_s_arrmul16_fa7_13_y2, h_s_arrmul16_fa7_13_y4);
  and_gate and_gate_h_s_arrmul16_and8_13_y0(a_8, b_13, h_s_arrmul16_and8_13_y0);
  fa fa_h_s_arrmul16_fa8_13_y2(h_s_arrmul16_and8_13_y0, h_s_arrmul16_fa9_12_y2, h_s_arrmul16_fa7_13_y4, h_s_arrmul16_fa8_13_y2, h_s_arrmul16_fa8_13_y4);
  and_gate and_gate_h_s_arrmul16_and9_13_y0(a_9, b_13, h_s_arrmul16_and9_13_y0);
  fa fa_h_s_arrmul16_fa9_13_y2(h_s_arrmul16_and9_13_y0, h_s_arrmul16_fa10_12_y2, h_s_arrmul16_fa8_13_y4, h_s_arrmul16_fa9_13_y2, h_s_arrmul16_fa9_13_y4);
  and_gate and_gate_h_s_arrmul16_and10_13_y0(a_10, b_13, h_s_arrmul16_and10_13_y0);
  fa fa_h_s_arrmul16_fa10_13_y2(h_s_arrmul16_and10_13_y0, h_s_arrmul16_fa11_12_y2, h_s_arrmul16_fa9_13_y4, h_s_arrmul16_fa10_13_y2, h_s_arrmul16_fa10_13_y4);
  and_gate and_gate_h_s_arrmul16_and11_13_y0(a_11, b_13, h_s_arrmul16_and11_13_y0);
  fa fa_h_s_arrmul16_fa11_13_y2(h_s_arrmul16_and11_13_y0, h_s_arrmul16_fa12_12_y2, h_s_arrmul16_fa10_13_y4, h_s_arrmul16_fa11_13_y2, h_s_arrmul16_fa11_13_y4);
  and_gate and_gate_h_s_arrmul16_and12_13_y0(a_12, b_13, h_s_arrmul16_and12_13_y0);
  fa fa_h_s_arrmul16_fa12_13_y2(h_s_arrmul16_and12_13_y0, h_s_arrmul16_fa13_12_y2, h_s_arrmul16_fa11_13_y4, h_s_arrmul16_fa12_13_y2, h_s_arrmul16_fa12_13_y4);
  and_gate and_gate_h_s_arrmul16_and13_13_y0(a_13, b_13, h_s_arrmul16_and13_13_y0);
  fa fa_h_s_arrmul16_fa13_13_y2(h_s_arrmul16_and13_13_y0, h_s_arrmul16_fa14_12_y2, h_s_arrmul16_fa12_13_y4, h_s_arrmul16_fa13_13_y2, h_s_arrmul16_fa13_13_y4);
  and_gate and_gate_h_s_arrmul16_and14_13_y0(a_14, b_13, h_s_arrmul16_and14_13_y0);
  fa fa_h_s_arrmul16_fa14_13_y2(h_s_arrmul16_and14_13_y0, h_s_arrmul16_fa15_12_y2, h_s_arrmul16_fa13_13_y4, h_s_arrmul16_fa14_13_y2, h_s_arrmul16_fa14_13_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_13_y0(a_15, b_13, h_s_arrmul16_nand15_13_y0);
  fa fa_h_s_arrmul16_fa15_13_y2(h_s_arrmul16_nand15_13_y0, h_s_arrmul16_fa15_12_y4, h_s_arrmul16_fa14_13_y4, h_s_arrmul16_fa15_13_y2, h_s_arrmul16_fa15_13_y4);
  and_gate and_gate_h_s_arrmul16_and0_14_y0(a_0, b_14, h_s_arrmul16_and0_14_y0);
  ha ha_h_s_arrmul16_ha0_14_y0(h_s_arrmul16_and0_14_y0, h_s_arrmul16_fa1_13_y2, h_s_arrmul16_ha0_14_y0, h_s_arrmul16_ha0_14_y1);
  and_gate and_gate_h_s_arrmul16_and1_14_y0(a_1, b_14, h_s_arrmul16_and1_14_y0);
  fa fa_h_s_arrmul16_fa1_14_y2(h_s_arrmul16_and1_14_y0, h_s_arrmul16_fa2_13_y2, h_s_arrmul16_ha0_14_y1, h_s_arrmul16_fa1_14_y2, h_s_arrmul16_fa1_14_y4);
  and_gate and_gate_h_s_arrmul16_and2_14_y0(a_2, b_14, h_s_arrmul16_and2_14_y0);
  fa fa_h_s_arrmul16_fa2_14_y2(h_s_arrmul16_and2_14_y0, h_s_arrmul16_fa3_13_y2, h_s_arrmul16_fa1_14_y4, h_s_arrmul16_fa2_14_y2, h_s_arrmul16_fa2_14_y4);
  and_gate and_gate_h_s_arrmul16_and3_14_y0(a_3, b_14, h_s_arrmul16_and3_14_y0);
  fa fa_h_s_arrmul16_fa3_14_y2(h_s_arrmul16_and3_14_y0, h_s_arrmul16_fa4_13_y2, h_s_arrmul16_fa2_14_y4, h_s_arrmul16_fa3_14_y2, h_s_arrmul16_fa3_14_y4);
  and_gate and_gate_h_s_arrmul16_and4_14_y0(a_4, b_14, h_s_arrmul16_and4_14_y0);
  fa fa_h_s_arrmul16_fa4_14_y2(h_s_arrmul16_and4_14_y0, h_s_arrmul16_fa5_13_y2, h_s_arrmul16_fa3_14_y4, h_s_arrmul16_fa4_14_y2, h_s_arrmul16_fa4_14_y4);
  and_gate and_gate_h_s_arrmul16_and5_14_y0(a_5, b_14, h_s_arrmul16_and5_14_y0);
  fa fa_h_s_arrmul16_fa5_14_y2(h_s_arrmul16_and5_14_y0, h_s_arrmul16_fa6_13_y2, h_s_arrmul16_fa4_14_y4, h_s_arrmul16_fa5_14_y2, h_s_arrmul16_fa5_14_y4);
  and_gate and_gate_h_s_arrmul16_and6_14_y0(a_6, b_14, h_s_arrmul16_and6_14_y0);
  fa fa_h_s_arrmul16_fa6_14_y2(h_s_arrmul16_and6_14_y0, h_s_arrmul16_fa7_13_y2, h_s_arrmul16_fa5_14_y4, h_s_arrmul16_fa6_14_y2, h_s_arrmul16_fa6_14_y4);
  and_gate and_gate_h_s_arrmul16_and7_14_y0(a_7, b_14, h_s_arrmul16_and7_14_y0);
  fa fa_h_s_arrmul16_fa7_14_y2(h_s_arrmul16_and7_14_y0, h_s_arrmul16_fa8_13_y2, h_s_arrmul16_fa6_14_y4, h_s_arrmul16_fa7_14_y2, h_s_arrmul16_fa7_14_y4);
  and_gate and_gate_h_s_arrmul16_and8_14_y0(a_8, b_14, h_s_arrmul16_and8_14_y0);
  fa fa_h_s_arrmul16_fa8_14_y2(h_s_arrmul16_and8_14_y0, h_s_arrmul16_fa9_13_y2, h_s_arrmul16_fa7_14_y4, h_s_arrmul16_fa8_14_y2, h_s_arrmul16_fa8_14_y4);
  and_gate and_gate_h_s_arrmul16_and9_14_y0(a_9, b_14, h_s_arrmul16_and9_14_y0);
  fa fa_h_s_arrmul16_fa9_14_y2(h_s_arrmul16_and9_14_y0, h_s_arrmul16_fa10_13_y2, h_s_arrmul16_fa8_14_y4, h_s_arrmul16_fa9_14_y2, h_s_arrmul16_fa9_14_y4);
  and_gate and_gate_h_s_arrmul16_and10_14_y0(a_10, b_14, h_s_arrmul16_and10_14_y0);
  fa fa_h_s_arrmul16_fa10_14_y2(h_s_arrmul16_and10_14_y0, h_s_arrmul16_fa11_13_y2, h_s_arrmul16_fa9_14_y4, h_s_arrmul16_fa10_14_y2, h_s_arrmul16_fa10_14_y4);
  and_gate and_gate_h_s_arrmul16_and11_14_y0(a_11, b_14, h_s_arrmul16_and11_14_y0);
  fa fa_h_s_arrmul16_fa11_14_y2(h_s_arrmul16_and11_14_y0, h_s_arrmul16_fa12_13_y2, h_s_arrmul16_fa10_14_y4, h_s_arrmul16_fa11_14_y2, h_s_arrmul16_fa11_14_y4);
  and_gate and_gate_h_s_arrmul16_and12_14_y0(a_12, b_14, h_s_arrmul16_and12_14_y0);
  fa fa_h_s_arrmul16_fa12_14_y2(h_s_arrmul16_and12_14_y0, h_s_arrmul16_fa13_13_y2, h_s_arrmul16_fa11_14_y4, h_s_arrmul16_fa12_14_y2, h_s_arrmul16_fa12_14_y4);
  and_gate and_gate_h_s_arrmul16_and13_14_y0(a_13, b_14, h_s_arrmul16_and13_14_y0);
  fa fa_h_s_arrmul16_fa13_14_y2(h_s_arrmul16_and13_14_y0, h_s_arrmul16_fa14_13_y2, h_s_arrmul16_fa12_14_y4, h_s_arrmul16_fa13_14_y2, h_s_arrmul16_fa13_14_y4);
  and_gate and_gate_h_s_arrmul16_and14_14_y0(a_14, b_14, h_s_arrmul16_and14_14_y0);
  fa fa_h_s_arrmul16_fa14_14_y2(h_s_arrmul16_and14_14_y0, h_s_arrmul16_fa15_13_y2, h_s_arrmul16_fa13_14_y4, h_s_arrmul16_fa14_14_y2, h_s_arrmul16_fa14_14_y4);
  nand_gate nand_gate_h_s_arrmul16_nand15_14_y0(a_15, b_14, h_s_arrmul16_nand15_14_y0);
  fa fa_h_s_arrmul16_fa15_14_y2(h_s_arrmul16_nand15_14_y0, h_s_arrmul16_fa15_13_y4, h_s_arrmul16_fa14_14_y4, h_s_arrmul16_fa15_14_y2, h_s_arrmul16_fa15_14_y4);
  nand_gate nand_gate_h_s_arrmul16_nand0_15_y0(a_0, b_15, h_s_arrmul16_nand0_15_y0);
  ha ha_h_s_arrmul16_ha0_15_y0(h_s_arrmul16_nand0_15_y0, h_s_arrmul16_fa1_14_y2, h_s_arrmul16_ha0_15_y0, h_s_arrmul16_ha0_15_y1);
  nand_gate nand_gate_h_s_arrmul16_nand1_15_y0(a_1, b_15, h_s_arrmul16_nand1_15_y0);
  fa fa_h_s_arrmul16_fa1_15_y2(h_s_arrmul16_nand1_15_y0, h_s_arrmul16_fa2_14_y2, h_s_arrmul16_ha0_15_y1, h_s_arrmul16_fa1_15_y2, h_s_arrmul16_fa1_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand2_15_y0(a_2, b_15, h_s_arrmul16_nand2_15_y0);
  fa fa_h_s_arrmul16_fa2_15_y2(h_s_arrmul16_nand2_15_y0, h_s_arrmul16_fa3_14_y2, h_s_arrmul16_fa1_15_y4, h_s_arrmul16_fa2_15_y2, h_s_arrmul16_fa2_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand3_15_y0(a_3, b_15, h_s_arrmul16_nand3_15_y0);
  fa fa_h_s_arrmul16_fa3_15_y2(h_s_arrmul16_nand3_15_y0, h_s_arrmul16_fa4_14_y2, h_s_arrmul16_fa2_15_y4, h_s_arrmul16_fa3_15_y2, h_s_arrmul16_fa3_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand4_15_y0(a_4, b_15, h_s_arrmul16_nand4_15_y0);
  fa fa_h_s_arrmul16_fa4_15_y2(h_s_arrmul16_nand4_15_y0, h_s_arrmul16_fa5_14_y2, h_s_arrmul16_fa3_15_y4, h_s_arrmul16_fa4_15_y2, h_s_arrmul16_fa4_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand5_15_y0(a_5, b_15, h_s_arrmul16_nand5_15_y0);
  fa fa_h_s_arrmul16_fa5_15_y2(h_s_arrmul16_nand5_15_y0, h_s_arrmul16_fa6_14_y2, h_s_arrmul16_fa4_15_y4, h_s_arrmul16_fa5_15_y2, h_s_arrmul16_fa5_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand6_15_y0(a_6, b_15, h_s_arrmul16_nand6_15_y0);
  fa fa_h_s_arrmul16_fa6_15_y2(h_s_arrmul16_nand6_15_y0, h_s_arrmul16_fa7_14_y2, h_s_arrmul16_fa5_15_y4, h_s_arrmul16_fa6_15_y2, h_s_arrmul16_fa6_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand7_15_y0(a_7, b_15, h_s_arrmul16_nand7_15_y0);
  fa fa_h_s_arrmul16_fa7_15_y2(h_s_arrmul16_nand7_15_y0, h_s_arrmul16_fa8_14_y2, h_s_arrmul16_fa6_15_y4, h_s_arrmul16_fa7_15_y2, h_s_arrmul16_fa7_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand8_15_y0(a_8, b_15, h_s_arrmul16_nand8_15_y0);
  fa fa_h_s_arrmul16_fa8_15_y2(h_s_arrmul16_nand8_15_y0, h_s_arrmul16_fa9_14_y2, h_s_arrmul16_fa7_15_y4, h_s_arrmul16_fa8_15_y2, h_s_arrmul16_fa8_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand9_15_y0(a_9, b_15, h_s_arrmul16_nand9_15_y0);
  fa fa_h_s_arrmul16_fa9_15_y2(h_s_arrmul16_nand9_15_y0, h_s_arrmul16_fa10_14_y2, h_s_arrmul16_fa8_15_y4, h_s_arrmul16_fa9_15_y2, h_s_arrmul16_fa9_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand10_15_y0(a_10, b_15, h_s_arrmul16_nand10_15_y0);
  fa fa_h_s_arrmul16_fa10_15_y2(h_s_arrmul16_nand10_15_y0, h_s_arrmul16_fa11_14_y2, h_s_arrmul16_fa9_15_y4, h_s_arrmul16_fa10_15_y2, h_s_arrmul16_fa10_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand11_15_y0(a_11, b_15, h_s_arrmul16_nand11_15_y0);
  fa fa_h_s_arrmul16_fa11_15_y2(h_s_arrmul16_nand11_15_y0, h_s_arrmul16_fa12_14_y2, h_s_arrmul16_fa10_15_y4, h_s_arrmul16_fa11_15_y2, h_s_arrmul16_fa11_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand12_15_y0(a_12, b_15, h_s_arrmul16_nand12_15_y0);
  fa fa_h_s_arrmul16_fa12_15_y2(h_s_arrmul16_nand12_15_y0, h_s_arrmul16_fa13_14_y2, h_s_arrmul16_fa11_15_y4, h_s_arrmul16_fa12_15_y2, h_s_arrmul16_fa12_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand13_15_y0(a_13, b_15, h_s_arrmul16_nand13_15_y0);
  fa fa_h_s_arrmul16_fa13_15_y2(h_s_arrmul16_nand13_15_y0, h_s_arrmul16_fa14_14_y2, h_s_arrmul16_fa12_15_y4, h_s_arrmul16_fa13_15_y2, h_s_arrmul16_fa13_15_y4);
  nand_gate nand_gate_h_s_arrmul16_nand14_15_y0(a_14, b_15, h_s_arrmul16_nand14_15_y0);
  fa fa_h_s_arrmul16_fa14_15_y2(h_s_arrmul16_nand14_15_y0, h_s_arrmul16_fa15_14_y2, h_s_arrmul16_fa13_15_y4, h_s_arrmul16_fa14_15_y2, h_s_arrmul16_fa14_15_y4);
  and_gate and_gate_h_s_arrmul16_and15_15_y0(a_15, b_15, h_s_arrmul16_and15_15_y0);
  fa fa_h_s_arrmul16_fa15_15_y2(h_s_arrmul16_and15_15_y0, h_s_arrmul16_fa15_14_y4, h_s_arrmul16_fa14_15_y4, h_s_arrmul16_fa15_15_y2, h_s_arrmul16_fa15_15_y4);
  xor_gate xor_gate_h_s_arrmul16_xor16_15_y0(h_s_arrmul16_fa15_15_y4, constant_wire_1, h_s_arrmul16_xor16_15_y0);

  assign out[0] = h_s_arrmul16_and0_0_y0;
  assign out[1] = h_s_arrmul16_ha0_1_y0;
  assign out[2] = h_s_arrmul16_ha0_2_y0;
  assign out[3] = h_s_arrmul16_ha0_3_y0;
  assign out[4] = h_s_arrmul16_ha0_4_y0;
  assign out[5] = h_s_arrmul16_ha0_5_y0;
  assign out[6] = h_s_arrmul16_ha0_6_y0;
  assign out[7] = h_s_arrmul16_ha0_7_y0;
  assign out[8] = h_s_arrmul16_ha0_8_y0;
  assign out[9] = h_s_arrmul16_ha0_9_y0;
  assign out[10] = h_s_arrmul16_ha0_10_y0;
  assign out[11] = h_s_arrmul16_ha0_11_y0;
  assign out[12] = h_s_arrmul16_ha0_12_y0;
  assign out[13] = h_s_arrmul16_ha0_13_y0;
  assign out[14] = h_s_arrmul16_ha0_14_y0;
  assign out[15] = h_s_arrmul16_ha0_15_y0;
  assign out[16] = h_s_arrmul16_fa1_15_y2;
  assign out[17] = h_s_arrmul16_fa2_15_y2;
  assign out[18] = h_s_arrmul16_fa3_15_y2;
  assign out[19] = h_s_arrmul16_fa4_15_y2;
  assign out[20] = h_s_arrmul16_fa5_15_y2;
  assign out[21] = h_s_arrmul16_fa6_15_y2;
  assign out[22] = h_s_arrmul16_fa7_15_y2;
  assign out[23] = h_s_arrmul16_fa8_15_y2;
  assign out[24] = h_s_arrmul16_fa9_15_y2;
  assign out[25] = h_s_arrmul16_fa10_15_y2;
  assign out[26] = h_s_arrmul16_fa11_15_y2;
  assign out[27] = h_s_arrmul16_fa12_15_y2;
  assign out[28] = h_s_arrmul16_fa13_15_y2;
  assign out[29] = h_s_arrmul16_fa14_15_y2;
  assign out[30] = h_s_arrmul16_fa15_15_y2;
  assign out[31] = h_s_arrmul16_xor16_15_y0;
endmodule