module f_u_dadda_cla32(input [31:0] a, input [31:0] b, output [63:0] f_u_dadda_cla32_out);
  wire f_u_dadda_cla32_and_28_0;
  wire f_u_dadda_cla32_and_27_1;
  wire f_u_dadda_cla32_ha0_xor0;
  wire f_u_dadda_cla32_ha0_and0;
  wire f_u_dadda_cla32_and_29_0;
  wire f_u_dadda_cla32_and_28_1;
  wire f_u_dadda_cla32_fa0_xor0;
  wire f_u_dadda_cla32_fa0_and0;
  wire f_u_dadda_cla32_fa0_xor1;
  wire f_u_dadda_cla32_fa0_and1;
  wire f_u_dadda_cla32_fa0_or0;
  wire f_u_dadda_cla32_and_27_2;
  wire f_u_dadda_cla32_and_26_3;
  wire f_u_dadda_cla32_ha1_xor0;
  wire f_u_dadda_cla32_ha1_and0;
  wire f_u_dadda_cla32_and_30_0;
  wire f_u_dadda_cla32_fa1_xor0;
  wire f_u_dadda_cla32_fa1_and0;
  wire f_u_dadda_cla32_fa1_xor1;
  wire f_u_dadda_cla32_fa1_and1;
  wire f_u_dadda_cla32_fa1_or0;
  wire f_u_dadda_cla32_and_29_1;
  wire f_u_dadda_cla32_and_28_2;
  wire f_u_dadda_cla32_and_27_3;
  wire f_u_dadda_cla32_fa2_xor0;
  wire f_u_dadda_cla32_fa2_and0;
  wire f_u_dadda_cla32_fa2_xor1;
  wire f_u_dadda_cla32_fa2_and1;
  wire f_u_dadda_cla32_fa2_or0;
  wire f_u_dadda_cla32_and_26_4;
  wire f_u_dadda_cla32_and_25_5;
  wire f_u_dadda_cla32_ha2_xor0;
  wire f_u_dadda_cla32_ha2_and0;
  wire f_u_dadda_cla32_fa3_xor0;
  wire f_u_dadda_cla32_fa3_and0;
  wire f_u_dadda_cla32_fa3_xor1;
  wire f_u_dadda_cla32_fa3_and1;
  wire f_u_dadda_cla32_fa3_or0;
  wire f_u_dadda_cla32_and_31_0;
  wire f_u_dadda_cla32_and_30_1;
  wire f_u_dadda_cla32_and_29_2;
  wire f_u_dadda_cla32_fa4_xor0;
  wire f_u_dadda_cla32_fa4_and0;
  wire f_u_dadda_cla32_fa4_xor1;
  wire f_u_dadda_cla32_fa4_and1;
  wire f_u_dadda_cla32_fa4_or0;
  wire f_u_dadda_cla32_and_28_3;
  wire f_u_dadda_cla32_and_27_4;
  wire f_u_dadda_cla32_and_26_5;
  wire f_u_dadda_cla32_fa5_xor0;
  wire f_u_dadda_cla32_fa5_and0;
  wire f_u_dadda_cla32_fa5_xor1;
  wire f_u_dadda_cla32_fa5_and1;
  wire f_u_dadda_cla32_fa5_or0;
  wire f_u_dadda_cla32_and_25_6;
  wire f_u_dadda_cla32_and_24_7;
  wire f_u_dadda_cla32_ha3_xor0;
  wire f_u_dadda_cla32_ha3_and0;
  wire f_u_dadda_cla32_fa6_xor0;
  wire f_u_dadda_cla32_fa6_and0;
  wire f_u_dadda_cla32_fa6_xor1;
  wire f_u_dadda_cla32_fa6_and1;
  wire f_u_dadda_cla32_fa6_or0;
  wire f_u_dadda_cla32_and_31_1;
  wire f_u_dadda_cla32_and_30_2;
  wire f_u_dadda_cla32_fa7_xor0;
  wire f_u_dadda_cla32_fa7_and0;
  wire f_u_dadda_cla32_fa7_xor1;
  wire f_u_dadda_cla32_fa7_and1;
  wire f_u_dadda_cla32_fa7_or0;
  wire f_u_dadda_cla32_and_29_3;
  wire f_u_dadda_cla32_and_28_4;
  wire f_u_dadda_cla32_and_27_5;
  wire f_u_dadda_cla32_fa8_xor0;
  wire f_u_dadda_cla32_fa8_and0;
  wire f_u_dadda_cla32_fa8_xor1;
  wire f_u_dadda_cla32_fa8_and1;
  wire f_u_dadda_cla32_fa8_or0;
  wire f_u_dadda_cla32_and_26_6;
  wire f_u_dadda_cla32_and_25_7;
  wire f_u_dadda_cla32_ha4_xor0;
  wire f_u_dadda_cla32_ha4_and0;
  wire f_u_dadda_cla32_fa9_xor0;
  wire f_u_dadda_cla32_fa9_and0;
  wire f_u_dadda_cla32_fa9_xor1;
  wire f_u_dadda_cla32_fa9_and1;
  wire f_u_dadda_cla32_fa9_or0;
  wire f_u_dadda_cla32_and_31_2;
  wire f_u_dadda_cla32_and_30_3;
  wire f_u_dadda_cla32_fa10_xor0;
  wire f_u_dadda_cla32_fa10_and0;
  wire f_u_dadda_cla32_fa10_xor1;
  wire f_u_dadda_cla32_fa10_and1;
  wire f_u_dadda_cla32_fa10_or0;
  wire f_u_dadda_cla32_and_29_4;
  wire f_u_dadda_cla32_and_28_5;
  wire f_u_dadda_cla32_and_27_6;
  wire f_u_dadda_cla32_fa11_xor0;
  wire f_u_dadda_cla32_fa11_and0;
  wire f_u_dadda_cla32_fa11_xor1;
  wire f_u_dadda_cla32_fa11_and1;
  wire f_u_dadda_cla32_fa11_or0;
  wire f_u_dadda_cla32_fa12_xor0;
  wire f_u_dadda_cla32_fa12_and0;
  wire f_u_dadda_cla32_fa12_xor1;
  wire f_u_dadda_cla32_fa12_and1;
  wire f_u_dadda_cla32_fa12_or0;
  wire f_u_dadda_cla32_and_31_3;
  wire f_u_dadda_cla32_and_30_4;
  wire f_u_dadda_cla32_and_29_5;
  wire f_u_dadda_cla32_fa13_xor0;
  wire f_u_dadda_cla32_fa13_and0;
  wire f_u_dadda_cla32_fa13_xor1;
  wire f_u_dadda_cla32_fa13_and1;
  wire f_u_dadda_cla32_fa13_or0;
  wire f_u_dadda_cla32_and_31_4;
  wire f_u_dadda_cla32_fa14_xor0;
  wire f_u_dadda_cla32_fa14_and0;
  wire f_u_dadda_cla32_fa14_xor1;
  wire f_u_dadda_cla32_fa14_and1;
  wire f_u_dadda_cla32_fa14_or0;
  wire f_u_dadda_cla32_and_6_0;
  wire f_u_dadda_cla32_and_5_1;
  wire f_u_dadda_cla32_ha5_xor0;
  wire f_u_dadda_cla32_ha5_and0;
  wire f_u_dadda_cla32_and_7_0;
  wire f_u_dadda_cla32_and_6_1;
  wire f_u_dadda_cla32_fa15_xor0;
  wire f_u_dadda_cla32_fa15_and0;
  wire f_u_dadda_cla32_fa15_xor1;
  wire f_u_dadda_cla32_fa15_and1;
  wire f_u_dadda_cla32_fa15_or0;
  wire f_u_dadda_cla32_and_5_2;
  wire f_u_dadda_cla32_and_4_3;
  wire f_u_dadda_cla32_ha6_xor0;
  wire f_u_dadda_cla32_ha6_and0;
  wire f_u_dadda_cla32_and_8_0;
  wire f_u_dadda_cla32_fa16_xor0;
  wire f_u_dadda_cla32_fa16_and0;
  wire f_u_dadda_cla32_fa16_xor1;
  wire f_u_dadda_cla32_fa16_and1;
  wire f_u_dadda_cla32_fa16_or0;
  wire f_u_dadda_cla32_and_7_1;
  wire f_u_dadda_cla32_and_6_2;
  wire f_u_dadda_cla32_and_5_3;
  wire f_u_dadda_cla32_fa17_xor0;
  wire f_u_dadda_cla32_fa17_and0;
  wire f_u_dadda_cla32_fa17_xor1;
  wire f_u_dadda_cla32_fa17_and1;
  wire f_u_dadda_cla32_fa17_or0;
  wire f_u_dadda_cla32_and_4_4;
  wire f_u_dadda_cla32_and_3_5;
  wire f_u_dadda_cla32_ha7_xor0;
  wire f_u_dadda_cla32_ha7_and0;
  wire f_u_dadda_cla32_fa18_xor0;
  wire f_u_dadda_cla32_fa18_and0;
  wire f_u_dadda_cla32_fa18_xor1;
  wire f_u_dadda_cla32_fa18_and1;
  wire f_u_dadda_cla32_fa18_or0;
  wire f_u_dadda_cla32_and_9_0;
  wire f_u_dadda_cla32_and_8_1;
  wire f_u_dadda_cla32_and_7_2;
  wire f_u_dadda_cla32_fa19_xor0;
  wire f_u_dadda_cla32_fa19_and0;
  wire f_u_dadda_cla32_fa19_xor1;
  wire f_u_dadda_cla32_fa19_and1;
  wire f_u_dadda_cla32_fa19_or0;
  wire f_u_dadda_cla32_and_6_3;
  wire f_u_dadda_cla32_and_5_4;
  wire f_u_dadda_cla32_and_4_5;
  wire f_u_dadda_cla32_fa20_xor0;
  wire f_u_dadda_cla32_fa20_and0;
  wire f_u_dadda_cla32_fa20_xor1;
  wire f_u_dadda_cla32_fa20_and1;
  wire f_u_dadda_cla32_fa20_or0;
  wire f_u_dadda_cla32_and_3_6;
  wire f_u_dadda_cla32_and_2_7;
  wire f_u_dadda_cla32_ha8_xor0;
  wire f_u_dadda_cla32_ha8_and0;
  wire f_u_dadda_cla32_fa21_xor0;
  wire f_u_dadda_cla32_fa21_and0;
  wire f_u_dadda_cla32_fa21_xor1;
  wire f_u_dadda_cla32_fa21_and1;
  wire f_u_dadda_cla32_fa21_or0;
  wire f_u_dadda_cla32_and_10_0;
  wire f_u_dadda_cla32_and_9_1;
  wire f_u_dadda_cla32_fa22_xor0;
  wire f_u_dadda_cla32_fa22_and0;
  wire f_u_dadda_cla32_fa22_xor1;
  wire f_u_dadda_cla32_fa22_and1;
  wire f_u_dadda_cla32_fa22_or0;
  wire f_u_dadda_cla32_and_8_2;
  wire f_u_dadda_cla32_and_7_3;
  wire f_u_dadda_cla32_and_6_4;
  wire f_u_dadda_cla32_fa23_xor0;
  wire f_u_dadda_cla32_fa23_and0;
  wire f_u_dadda_cla32_fa23_xor1;
  wire f_u_dadda_cla32_fa23_and1;
  wire f_u_dadda_cla32_fa23_or0;
  wire f_u_dadda_cla32_and_5_5;
  wire f_u_dadda_cla32_and_4_6;
  wire f_u_dadda_cla32_and_3_7;
  wire f_u_dadda_cla32_fa24_xor0;
  wire f_u_dadda_cla32_fa24_and0;
  wire f_u_dadda_cla32_fa24_xor1;
  wire f_u_dadda_cla32_fa24_and1;
  wire f_u_dadda_cla32_fa24_or0;
  wire f_u_dadda_cla32_and_2_8;
  wire f_u_dadda_cla32_and_1_9;
  wire f_u_dadda_cla32_ha9_xor0;
  wire f_u_dadda_cla32_ha9_and0;
  wire f_u_dadda_cla32_fa25_xor0;
  wire f_u_dadda_cla32_fa25_and0;
  wire f_u_dadda_cla32_fa25_xor1;
  wire f_u_dadda_cla32_fa25_and1;
  wire f_u_dadda_cla32_fa25_or0;
  wire f_u_dadda_cla32_and_11_0;
  wire f_u_dadda_cla32_fa26_xor0;
  wire f_u_dadda_cla32_fa26_and0;
  wire f_u_dadda_cla32_fa26_xor1;
  wire f_u_dadda_cla32_fa26_and1;
  wire f_u_dadda_cla32_fa26_or0;
  wire f_u_dadda_cla32_and_10_1;
  wire f_u_dadda_cla32_and_9_2;
  wire f_u_dadda_cla32_and_8_3;
  wire f_u_dadda_cla32_fa27_xor0;
  wire f_u_dadda_cla32_fa27_and0;
  wire f_u_dadda_cla32_fa27_xor1;
  wire f_u_dadda_cla32_fa27_and1;
  wire f_u_dadda_cla32_fa27_or0;
  wire f_u_dadda_cla32_and_7_4;
  wire f_u_dadda_cla32_and_6_5;
  wire f_u_dadda_cla32_and_5_6;
  wire f_u_dadda_cla32_fa28_xor0;
  wire f_u_dadda_cla32_fa28_and0;
  wire f_u_dadda_cla32_fa28_xor1;
  wire f_u_dadda_cla32_fa28_and1;
  wire f_u_dadda_cla32_fa28_or0;
  wire f_u_dadda_cla32_and_4_7;
  wire f_u_dadda_cla32_and_3_8;
  wire f_u_dadda_cla32_and_2_9;
  wire f_u_dadda_cla32_fa29_xor0;
  wire f_u_dadda_cla32_fa29_and0;
  wire f_u_dadda_cla32_fa29_xor1;
  wire f_u_dadda_cla32_fa29_and1;
  wire f_u_dadda_cla32_fa29_or0;
  wire f_u_dadda_cla32_and_1_10;
  wire f_u_dadda_cla32_and_0_11;
  wire f_u_dadda_cla32_ha10_xor0;
  wire f_u_dadda_cla32_ha10_and0;
  wire f_u_dadda_cla32_fa30_xor0;
  wire f_u_dadda_cla32_fa30_and0;
  wire f_u_dadda_cla32_fa30_xor1;
  wire f_u_dadda_cla32_fa30_and1;
  wire f_u_dadda_cla32_fa30_or0;
  wire f_u_dadda_cla32_fa31_xor0;
  wire f_u_dadda_cla32_fa31_and0;
  wire f_u_dadda_cla32_fa31_xor1;
  wire f_u_dadda_cla32_fa31_and1;
  wire f_u_dadda_cla32_fa31_or0;
  wire f_u_dadda_cla32_and_12_0;
  wire f_u_dadda_cla32_and_11_1;
  wire f_u_dadda_cla32_and_10_2;
  wire f_u_dadda_cla32_fa32_xor0;
  wire f_u_dadda_cla32_fa32_and0;
  wire f_u_dadda_cla32_fa32_xor1;
  wire f_u_dadda_cla32_fa32_and1;
  wire f_u_dadda_cla32_fa32_or0;
  wire f_u_dadda_cla32_and_9_3;
  wire f_u_dadda_cla32_and_8_4;
  wire f_u_dadda_cla32_and_7_5;
  wire f_u_dadda_cla32_fa33_xor0;
  wire f_u_dadda_cla32_fa33_and0;
  wire f_u_dadda_cla32_fa33_xor1;
  wire f_u_dadda_cla32_fa33_and1;
  wire f_u_dadda_cla32_fa33_or0;
  wire f_u_dadda_cla32_and_6_6;
  wire f_u_dadda_cla32_and_5_7;
  wire f_u_dadda_cla32_and_4_8;
  wire f_u_dadda_cla32_fa34_xor0;
  wire f_u_dadda_cla32_fa34_and0;
  wire f_u_dadda_cla32_fa34_xor1;
  wire f_u_dadda_cla32_fa34_and1;
  wire f_u_dadda_cla32_fa34_or0;
  wire f_u_dadda_cla32_and_3_9;
  wire f_u_dadda_cla32_and_2_10;
  wire f_u_dadda_cla32_and_1_11;
  wire f_u_dadda_cla32_fa35_xor0;
  wire f_u_dadda_cla32_fa35_and0;
  wire f_u_dadda_cla32_fa35_xor1;
  wire f_u_dadda_cla32_fa35_and1;
  wire f_u_dadda_cla32_fa35_or0;
  wire f_u_dadda_cla32_and_0_12;
  wire f_u_dadda_cla32_ha11_xor0;
  wire f_u_dadda_cla32_ha11_and0;
  wire f_u_dadda_cla32_fa36_xor0;
  wire f_u_dadda_cla32_fa36_and0;
  wire f_u_dadda_cla32_fa36_xor1;
  wire f_u_dadda_cla32_fa36_and1;
  wire f_u_dadda_cla32_fa36_or0;
  wire f_u_dadda_cla32_fa37_xor0;
  wire f_u_dadda_cla32_fa37_and0;
  wire f_u_dadda_cla32_fa37_xor1;
  wire f_u_dadda_cla32_fa37_and1;
  wire f_u_dadda_cla32_fa37_or0;
  wire f_u_dadda_cla32_and_13_0;
  wire f_u_dadda_cla32_and_12_1;
  wire f_u_dadda_cla32_fa38_xor0;
  wire f_u_dadda_cla32_fa38_and0;
  wire f_u_dadda_cla32_fa38_xor1;
  wire f_u_dadda_cla32_fa38_and1;
  wire f_u_dadda_cla32_fa38_or0;
  wire f_u_dadda_cla32_and_11_2;
  wire f_u_dadda_cla32_and_10_3;
  wire f_u_dadda_cla32_and_9_4;
  wire f_u_dadda_cla32_fa39_xor0;
  wire f_u_dadda_cla32_fa39_and0;
  wire f_u_dadda_cla32_fa39_xor1;
  wire f_u_dadda_cla32_fa39_and1;
  wire f_u_dadda_cla32_fa39_or0;
  wire f_u_dadda_cla32_and_8_5;
  wire f_u_dadda_cla32_and_7_6;
  wire f_u_dadda_cla32_and_6_7;
  wire f_u_dadda_cla32_fa40_xor0;
  wire f_u_dadda_cla32_fa40_and0;
  wire f_u_dadda_cla32_fa40_xor1;
  wire f_u_dadda_cla32_fa40_and1;
  wire f_u_dadda_cla32_fa40_or0;
  wire f_u_dadda_cla32_and_5_8;
  wire f_u_dadda_cla32_and_4_9;
  wire f_u_dadda_cla32_and_3_10;
  wire f_u_dadda_cla32_fa41_xor0;
  wire f_u_dadda_cla32_fa41_and0;
  wire f_u_dadda_cla32_fa41_xor1;
  wire f_u_dadda_cla32_fa41_and1;
  wire f_u_dadda_cla32_fa41_or0;
  wire f_u_dadda_cla32_and_2_11;
  wire f_u_dadda_cla32_and_1_12;
  wire f_u_dadda_cla32_and_0_13;
  wire f_u_dadda_cla32_fa42_xor0;
  wire f_u_dadda_cla32_fa42_and0;
  wire f_u_dadda_cla32_fa42_xor1;
  wire f_u_dadda_cla32_fa42_and1;
  wire f_u_dadda_cla32_fa42_or0;
  wire f_u_dadda_cla32_ha12_xor0;
  wire f_u_dadda_cla32_ha12_and0;
  wire f_u_dadda_cla32_fa43_xor0;
  wire f_u_dadda_cla32_fa43_and0;
  wire f_u_dadda_cla32_fa43_xor1;
  wire f_u_dadda_cla32_fa43_and1;
  wire f_u_dadda_cla32_fa43_or0;
  wire f_u_dadda_cla32_fa44_xor0;
  wire f_u_dadda_cla32_fa44_and0;
  wire f_u_dadda_cla32_fa44_xor1;
  wire f_u_dadda_cla32_fa44_and1;
  wire f_u_dadda_cla32_fa44_or0;
  wire f_u_dadda_cla32_and_14_0;
  wire f_u_dadda_cla32_fa45_xor0;
  wire f_u_dadda_cla32_fa45_and0;
  wire f_u_dadda_cla32_fa45_xor1;
  wire f_u_dadda_cla32_fa45_and1;
  wire f_u_dadda_cla32_fa45_or0;
  wire f_u_dadda_cla32_and_13_1;
  wire f_u_dadda_cla32_and_12_2;
  wire f_u_dadda_cla32_and_11_3;
  wire f_u_dadda_cla32_fa46_xor0;
  wire f_u_dadda_cla32_fa46_and0;
  wire f_u_dadda_cla32_fa46_xor1;
  wire f_u_dadda_cla32_fa46_and1;
  wire f_u_dadda_cla32_fa46_or0;
  wire f_u_dadda_cla32_and_10_4;
  wire f_u_dadda_cla32_and_9_5;
  wire f_u_dadda_cla32_and_8_6;
  wire f_u_dadda_cla32_fa47_xor0;
  wire f_u_dadda_cla32_fa47_and0;
  wire f_u_dadda_cla32_fa47_xor1;
  wire f_u_dadda_cla32_fa47_and1;
  wire f_u_dadda_cla32_fa47_or0;
  wire f_u_dadda_cla32_and_7_7;
  wire f_u_dadda_cla32_and_6_8;
  wire f_u_dadda_cla32_and_5_9;
  wire f_u_dadda_cla32_fa48_xor0;
  wire f_u_dadda_cla32_fa48_and0;
  wire f_u_dadda_cla32_fa48_xor1;
  wire f_u_dadda_cla32_fa48_and1;
  wire f_u_dadda_cla32_fa48_or0;
  wire f_u_dadda_cla32_and_4_10;
  wire f_u_dadda_cla32_and_3_11;
  wire f_u_dadda_cla32_and_2_12;
  wire f_u_dadda_cla32_fa49_xor0;
  wire f_u_dadda_cla32_fa49_and0;
  wire f_u_dadda_cla32_fa49_xor1;
  wire f_u_dadda_cla32_fa49_and1;
  wire f_u_dadda_cla32_fa49_or0;
  wire f_u_dadda_cla32_and_1_13;
  wire f_u_dadda_cla32_and_0_14;
  wire f_u_dadda_cla32_fa50_xor0;
  wire f_u_dadda_cla32_fa50_and0;
  wire f_u_dadda_cla32_fa50_xor1;
  wire f_u_dadda_cla32_fa50_and1;
  wire f_u_dadda_cla32_fa50_or0;
  wire f_u_dadda_cla32_ha13_xor0;
  wire f_u_dadda_cla32_ha13_and0;
  wire f_u_dadda_cla32_fa51_xor0;
  wire f_u_dadda_cla32_fa51_and0;
  wire f_u_dadda_cla32_fa51_xor1;
  wire f_u_dadda_cla32_fa51_and1;
  wire f_u_dadda_cla32_fa51_or0;
  wire f_u_dadda_cla32_fa52_xor0;
  wire f_u_dadda_cla32_fa52_and0;
  wire f_u_dadda_cla32_fa52_xor1;
  wire f_u_dadda_cla32_fa52_and1;
  wire f_u_dadda_cla32_fa52_or0;
  wire f_u_dadda_cla32_fa53_xor0;
  wire f_u_dadda_cla32_fa53_and0;
  wire f_u_dadda_cla32_fa53_xor1;
  wire f_u_dadda_cla32_fa53_and1;
  wire f_u_dadda_cla32_fa53_or0;
  wire f_u_dadda_cla32_and_15_0;
  wire f_u_dadda_cla32_and_14_1;
  wire f_u_dadda_cla32_and_13_2;
  wire f_u_dadda_cla32_fa54_xor0;
  wire f_u_dadda_cla32_fa54_and0;
  wire f_u_dadda_cla32_fa54_xor1;
  wire f_u_dadda_cla32_fa54_and1;
  wire f_u_dadda_cla32_fa54_or0;
  wire f_u_dadda_cla32_and_12_3;
  wire f_u_dadda_cla32_and_11_4;
  wire f_u_dadda_cla32_and_10_5;
  wire f_u_dadda_cla32_fa55_xor0;
  wire f_u_dadda_cla32_fa55_and0;
  wire f_u_dadda_cla32_fa55_xor1;
  wire f_u_dadda_cla32_fa55_and1;
  wire f_u_dadda_cla32_fa55_or0;
  wire f_u_dadda_cla32_and_9_6;
  wire f_u_dadda_cla32_and_8_7;
  wire f_u_dadda_cla32_and_7_8;
  wire f_u_dadda_cla32_fa56_xor0;
  wire f_u_dadda_cla32_fa56_and0;
  wire f_u_dadda_cla32_fa56_xor1;
  wire f_u_dadda_cla32_fa56_and1;
  wire f_u_dadda_cla32_fa56_or0;
  wire f_u_dadda_cla32_and_6_9;
  wire f_u_dadda_cla32_and_5_10;
  wire f_u_dadda_cla32_and_4_11;
  wire f_u_dadda_cla32_fa57_xor0;
  wire f_u_dadda_cla32_fa57_and0;
  wire f_u_dadda_cla32_fa57_xor1;
  wire f_u_dadda_cla32_fa57_and1;
  wire f_u_dadda_cla32_fa57_or0;
  wire f_u_dadda_cla32_and_3_12;
  wire f_u_dadda_cla32_and_2_13;
  wire f_u_dadda_cla32_and_1_14;
  wire f_u_dadda_cla32_fa58_xor0;
  wire f_u_dadda_cla32_fa58_and0;
  wire f_u_dadda_cla32_fa58_xor1;
  wire f_u_dadda_cla32_fa58_and1;
  wire f_u_dadda_cla32_fa58_or0;
  wire f_u_dadda_cla32_and_0_15;
  wire f_u_dadda_cla32_fa59_xor0;
  wire f_u_dadda_cla32_fa59_and0;
  wire f_u_dadda_cla32_fa59_xor1;
  wire f_u_dadda_cla32_fa59_and1;
  wire f_u_dadda_cla32_fa59_or0;
  wire f_u_dadda_cla32_ha14_xor0;
  wire f_u_dadda_cla32_ha14_and0;
  wire f_u_dadda_cla32_fa60_xor0;
  wire f_u_dadda_cla32_fa60_and0;
  wire f_u_dadda_cla32_fa60_xor1;
  wire f_u_dadda_cla32_fa60_and1;
  wire f_u_dadda_cla32_fa60_or0;
  wire f_u_dadda_cla32_fa61_xor0;
  wire f_u_dadda_cla32_fa61_and0;
  wire f_u_dadda_cla32_fa61_xor1;
  wire f_u_dadda_cla32_fa61_and1;
  wire f_u_dadda_cla32_fa61_or0;
  wire f_u_dadda_cla32_fa62_xor0;
  wire f_u_dadda_cla32_fa62_and0;
  wire f_u_dadda_cla32_fa62_xor1;
  wire f_u_dadda_cla32_fa62_and1;
  wire f_u_dadda_cla32_fa62_or0;
  wire f_u_dadda_cla32_and_16_0;
  wire f_u_dadda_cla32_and_15_1;
  wire f_u_dadda_cla32_fa63_xor0;
  wire f_u_dadda_cla32_fa63_and0;
  wire f_u_dadda_cla32_fa63_xor1;
  wire f_u_dadda_cla32_fa63_and1;
  wire f_u_dadda_cla32_fa63_or0;
  wire f_u_dadda_cla32_and_14_2;
  wire f_u_dadda_cla32_and_13_3;
  wire f_u_dadda_cla32_and_12_4;
  wire f_u_dadda_cla32_fa64_xor0;
  wire f_u_dadda_cla32_fa64_and0;
  wire f_u_dadda_cla32_fa64_xor1;
  wire f_u_dadda_cla32_fa64_and1;
  wire f_u_dadda_cla32_fa64_or0;
  wire f_u_dadda_cla32_and_11_5;
  wire f_u_dadda_cla32_and_10_6;
  wire f_u_dadda_cla32_and_9_7;
  wire f_u_dadda_cla32_fa65_xor0;
  wire f_u_dadda_cla32_fa65_and0;
  wire f_u_dadda_cla32_fa65_xor1;
  wire f_u_dadda_cla32_fa65_and1;
  wire f_u_dadda_cla32_fa65_or0;
  wire f_u_dadda_cla32_and_8_8;
  wire f_u_dadda_cla32_and_7_9;
  wire f_u_dadda_cla32_and_6_10;
  wire f_u_dadda_cla32_fa66_xor0;
  wire f_u_dadda_cla32_fa66_and0;
  wire f_u_dadda_cla32_fa66_xor1;
  wire f_u_dadda_cla32_fa66_and1;
  wire f_u_dadda_cla32_fa66_or0;
  wire f_u_dadda_cla32_and_5_11;
  wire f_u_dadda_cla32_and_4_12;
  wire f_u_dadda_cla32_and_3_13;
  wire f_u_dadda_cla32_fa67_xor0;
  wire f_u_dadda_cla32_fa67_and0;
  wire f_u_dadda_cla32_fa67_xor1;
  wire f_u_dadda_cla32_fa67_and1;
  wire f_u_dadda_cla32_fa67_or0;
  wire f_u_dadda_cla32_and_2_14;
  wire f_u_dadda_cla32_and_1_15;
  wire f_u_dadda_cla32_and_0_16;
  wire f_u_dadda_cla32_fa68_xor0;
  wire f_u_dadda_cla32_fa68_and0;
  wire f_u_dadda_cla32_fa68_xor1;
  wire f_u_dadda_cla32_fa68_and1;
  wire f_u_dadda_cla32_fa68_or0;
  wire f_u_dadda_cla32_fa69_xor0;
  wire f_u_dadda_cla32_fa69_and0;
  wire f_u_dadda_cla32_fa69_xor1;
  wire f_u_dadda_cla32_fa69_and1;
  wire f_u_dadda_cla32_fa69_or0;
  wire f_u_dadda_cla32_ha15_xor0;
  wire f_u_dadda_cla32_ha15_and0;
  wire f_u_dadda_cla32_fa70_xor0;
  wire f_u_dadda_cla32_fa70_and0;
  wire f_u_dadda_cla32_fa70_xor1;
  wire f_u_dadda_cla32_fa70_and1;
  wire f_u_dadda_cla32_fa70_or0;
  wire f_u_dadda_cla32_fa71_xor0;
  wire f_u_dadda_cla32_fa71_and0;
  wire f_u_dadda_cla32_fa71_xor1;
  wire f_u_dadda_cla32_fa71_and1;
  wire f_u_dadda_cla32_fa71_or0;
  wire f_u_dadda_cla32_fa72_xor0;
  wire f_u_dadda_cla32_fa72_and0;
  wire f_u_dadda_cla32_fa72_xor1;
  wire f_u_dadda_cla32_fa72_and1;
  wire f_u_dadda_cla32_fa72_or0;
  wire f_u_dadda_cla32_and_17_0;
  wire f_u_dadda_cla32_fa73_xor0;
  wire f_u_dadda_cla32_fa73_and0;
  wire f_u_dadda_cla32_fa73_xor1;
  wire f_u_dadda_cla32_fa73_and1;
  wire f_u_dadda_cla32_fa73_or0;
  wire f_u_dadda_cla32_and_16_1;
  wire f_u_dadda_cla32_and_15_2;
  wire f_u_dadda_cla32_and_14_3;
  wire f_u_dadda_cla32_fa74_xor0;
  wire f_u_dadda_cla32_fa74_and0;
  wire f_u_dadda_cla32_fa74_xor1;
  wire f_u_dadda_cla32_fa74_and1;
  wire f_u_dadda_cla32_fa74_or0;
  wire f_u_dadda_cla32_and_13_4;
  wire f_u_dadda_cla32_and_12_5;
  wire f_u_dadda_cla32_and_11_6;
  wire f_u_dadda_cla32_fa75_xor0;
  wire f_u_dadda_cla32_fa75_and0;
  wire f_u_dadda_cla32_fa75_xor1;
  wire f_u_dadda_cla32_fa75_and1;
  wire f_u_dadda_cla32_fa75_or0;
  wire f_u_dadda_cla32_and_10_7;
  wire f_u_dadda_cla32_and_9_8;
  wire f_u_dadda_cla32_and_8_9;
  wire f_u_dadda_cla32_fa76_xor0;
  wire f_u_dadda_cla32_fa76_and0;
  wire f_u_dadda_cla32_fa76_xor1;
  wire f_u_dadda_cla32_fa76_and1;
  wire f_u_dadda_cla32_fa76_or0;
  wire f_u_dadda_cla32_and_7_10;
  wire f_u_dadda_cla32_and_6_11;
  wire f_u_dadda_cla32_and_5_12;
  wire f_u_dadda_cla32_fa77_xor0;
  wire f_u_dadda_cla32_fa77_and0;
  wire f_u_dadda_cla32_fa77_xor1;
  wire f_u_dadda_cla32_fa77_and1;
  wire f_u_dadda_cla32_fa77_or0;
  wire f_u_dadda_cla32_and_4_13;
  wire f_u_dadda_cla32_and_3_14;
  wire f_u_dadda_cla32_and_2_15;
  wire f_u_dadda_cla32_fa78_xor0;
  wire f_u_dadda_cla32_fa78_and0;
  wire f_u_dadda_cla32_fa78_xor1;
  wire f_u_dadda_cla32_fa78_and1;
  wire f_u_dadda_cla32_fa78_or0;
  wire f_u_dadda_cla32_and_1_16;
  wire f_u_dadda_cla32_and_0_17;
  wire f_u_dadda_cla32_fa79_xor0;
  wire f_u_dadda_cla32_fa79_and0;
  wire f_u_dadda_cla32_fa79_xor1;
  wire f_u_dadda_cla32_fa79_and1;
  wire f_u_dadda_cla32_fa79_or0;
  wire f_u_dadda_cla32_fa80_xor0;
  wire f_u_dadda_cla32_fa80_and0;
  wire f_u_dadda_cla32_fa80_xor1;
  wire f_u_dadda_cla32_fa80_and1;
  wire f_u_dadda_cla32_fa80_or0;
  wire f_u_dadda_cla32_ha16_xor0;
  wire f_u_dadda_cla32_ha16_and0;
  wire f_u_dadda_cla32_fa81_xor0;
  wire f_u_dadda_cla32_fa81_and0;
  wire f_u_dadda_cla32_fa81_xor1;
  wire f_u_dadda_cla32_fa81_and1;
  wire f_u_dadda_cla32_fa81_or0;
  wire f_u_dadda_cla32_fa82_xor0;
  wire f_u_dadda_cla32_fa82_and0;
  wire f_u_dadda_cla32_fa82_xor1;
  wire f_u_dadda_cla32_fa82_and1;
  wire f_u_dadda_cla32_fa82_or0;
  wire f_u_dadda_cla32_fa83_xor0;
  wire f_u_dadda_cla32_fa83_and0;
  wire f_u_dadda_cla32_fa83_xor1;
  wire f_u_dadda_cla32_fa83_and1;
  wire f_u_dadda_cla32_fa83_or0;
  wire f_u_dadda_cla32_fa84_xor0;
  wire f_u_dadda_cla32_fa84_and0;
  wire f_u_dadda_cla32_fa84_xor1;
  wire f_u_dadda_cla32_fa84_and1;
  wire f_u_dadda_cla32_fa84_or0;
  wire f_u_dadda_cla32_and_18_0;
  wire f_u_dadda_cla32_and_17_1;
  wire f_u_dadda_cla32_and_16_2;
  wire f_u_dadda_cla32_fa85_xor0;
  wire f_u_dadda_cla32_fa85_and0;
  wire f_u_dadda_cla32_fa85_xor1;
  wire f_u_dadda_cla32_fa85_and1;
  wire f_u_dadda_cla32_fa85_or0;
  wire f_u_dadda_cla32_and_15_3;
  wire f_u_dadda_cla32_and_14_4;
  wire f_u_dadda_cla32_and_13_5;
  wire f_u_dadda_cla32_fa86_xor0;
  wire f_u_dadda_cla32_fa86_and0;
  wire f_u_dadda_cla32_fa86_xor1;
  wire f_u_dadda_cla32_fa86_and1;
  wire f_u_dadda_cla32_fa86_or0;
  wire f_u_dadda_cla32_and_12_6;
  wire f_u_dadda_cla32_and_11_7;
  wire f_u_dadda_cla32_and_10_8;
  wire f_u_dadda_cla32_fa87_xor0;
  wire f_u_dadda_cla32_fa87_and0;
  wire f_u_dadda_cla32_fa87_xor1;
  wire f_u_dadda_cla32_fa87_and1;
  wire f_u_dadda_cla32_fa87_or0;
  wire f_u_dadda_cla32_and_9_9;
  wire f_u_dadda_cla32_and_8_10;
  wire f_u_dadda_cla32_and_7_11;
  wire f_u_dadda_cla32_fa88_xor0;
  wire f_u_dadda_cla32_fa88_and0;
  wire f_u_dadda_cla32_fa88_xor1;
  wire f_u_dadda_cla32_fa88_and1;
  wire f_u_dadda_cla32_fa88_or0;
  wire f_u_dadda_cla32_and_6_12;
  wire f_u_dadda_cla32_and_5_13;
  wire f_u_dadda_cla32_and_4_14;
  wire f_u_dadda_cla32_fa89_xor0;
  wire f_u_dadda_cla32_fa89_and0;
  wire f_u_dadda_cla32_fa89_xor1;
  wire f_u_dadda_cla32_fa89_and1;
  wire f_u_dadda_cla32_fa89_or0;
  wire f_u_dadda_cla32_and_3_15;
  wire f_u_dadda_cla32_and_2_16;
  wire f_u_dadda_cla32_and_1_17;
  wire f_u_dadda_cla32_fa90_xor0;
  wire f_u_dadda_cla32_fa90_and0;
  wire f_u_dadda_cla32_fa90_xor1;
  wire f_u_dadda_cla32_fa90_and1;
  wire f_u_dadda_cla32_fa90_or0;
  wire f_u_dadda_cla32_and_0_18;
  wire f_u_dadda_cla32_fa91_xor0;
  wire f_u_dadda_cla32_fa91_and0;
  wire f_u_dadda_cla32_fa91_xor1;
  wire f_u_dadda_cla32_fa91_and1;
  wire f_u_dadda_cla32_fa91_or0;
  wire f_u_dadda_cla32_fa92_xor0;
  wire f_u_dadda_cla32_fa92_and0;
  wire f_u_dadda_cla32_fa92_xor1;
  wire f_u_dadda_cla32_fa92_and1;
  wire f_u_dadda_cla32_fa92_or0;
  wire f_u_dadda_cla32_ha17_xor0;
  wire f_u_dadda_cla32_ha17_and0;
  wire f_u_dadda_cla32_fa93_xor0;
  wire f_u_dadda_cla32_fa93_and0;
  wire f_u_dadda_cla32_fa93_xor1;
  wire f_u_dadda_cla32_fa93_and1;
  wire f_u_dadda_cla32_fa93_or0;
  wire f_u_dadda_cla32_fa94_xor0;
  wire f_u_dadda_cla32_fa94_and0;
  wire f_u_dadda_cla32_fa94_xor1;
  wire f_u_dadda_cla32_fa94_and1;
  wire f_u_dadda_cla32_fa94_or0;
  wire f_u_dadda_cla32_fa95_xor0;
  wire f_u_dadda_cla32_fa95_and0;
  wire f_u_dadda_cla32_fa95_xor1;
  wire f_u_dadda_cla32_fa95_and1;
  wire f_u_dadda_cla32_fa95_or0;
  wire f_u_dadda_cla32_fa96_xor0;
  wire f_u_dadda_cla32_fa96_and0;
  wire f_u_dadda_cla32_fa96_xor1;
  wire f_u_dadda_cla32_fa96_and1;
  wire f_u_dadda_cla32_fa96_or0;
  wire f_u_dadda_cla32_and_19_0;
  wire f_u_dadda_cla32_and_18_1;
  wire f_u_dadda_cla32_fa97_xor0;
  wire f_u_dadda_cla32_fa97_and0;
  wire f_u_dadda_cla32_fa97_xor1;
  wire f_u_dadda_cla32_fa97_and1;
  wire f_u_dadda_cla32_fa97_or0;
  wire f_u_dadda_cla32_and_17_2;
  wire f_u_dadda_cla32_and_16_3;
  wire f_u_dadda_cla32_and_15_4;
  wire f_u_dadda_cla32_fa98_xor0;
  wire f_u_dadda_cla32_fa98_and0;
  wire f_u_dadda_cla32_fa98_xor1;
  wire f_u_dadda_cla32_fa98_and1;
  wire f_u_dadda_cla32_fa98_or0;
  wire f_u_dadda_cla32_and_14_5;
  wire f_u_dadda_cla32_and_13_6;
  wire f_u_dadda_cla32_and_12_7;
  wire f_u_dadda_cla32_fa99_xor0;
  wire f_u_dadda_cla32_fa99_and0;
  wire f_u_dadda_cla32_fa99_xor1;
  wire f_u_dadda_cla32_fa99_and1;
  wire f_u_dadda_cla32_fa99_or0;
  wire f_u_dadda_cla32_and_11_8;
  wire f_u_dadda_cla32_and_10_9;
  wire f_u_dadda_cla32_and_9_10;
  wire f_u_dadda_cla32_fa100_xor0;
  wire f_u_dadda_cla32_fa100_and0;
  wire f_u_dadda_cla32_fa100_xor1;
  wire f_u_dadda_cla32_fa100_and1;
  wire f_u_dadda_cla32_fa100_or0;
  wire f_u_dadda_cla32_and_8_11;
  wire f_u_dadda_cla32_and_7_12;
  wire f_u_dadda_cla32_and_6_13;
  wire f_u_dadda_cla32_fa101_xor0;
  wire f_u_dadda_cla32_fa101_and0;
  wire f_u_dadda_cla32_fa101_xor1;
  wire f_u_dadda_cla32_fa101_and1;
  wire f_u_dadda_cla32_fa101_or0;
  wire f_u_dadda_cla32_and_5_14;
  wire f_u_dadda_cla32_and_4_15;
  wire f_u_dadda_cla32_and_3_16;
  wire f_u_dadda_cla32_fa102_xor0;
  wire f_u_dadda_cla32_fa102_and0;
  wire f_u_dadda_cla32_fa102_xor1;
  wire f_u_dadda_cla32_fa102_and1;
  wire f_u_dadda_cla32_fa102_or0;
  wire f_u_dadda_cla32_and_2_17;
  wire f_u_dadda_cla32_and_1_18;
  wire f_u_dadda_cla32_and_0_19;
  wire f_u_dadda_cla32_fa103_xor0;
  wire f_u_dadda_cla32_fa103_and0;
  wire f_u_dadda_cla32_fa103_xor1;
  wire f_u_dadda_cla32_fa103_and1;
  wire f_u_dadda_cla32_fa103_or0;
  wire f_u_dadda_cla32_fa104_xor0;
  wire f_u_dadda_cla32_fa104_and0;
  wire f_u_dadda_cla32_fa104_xor1;
  wire f_u_dadda_cla32_fa104_and1;
  wire f_u_dadda_cla32_fa104_or0;
  wire f_u_dadda_cla32_fa105_xor0;
  wire f_u_dadda_cla32_fa105_and0;
  wire f_u_dadda_cla32_fa105_xor1;
  wire f_u_dadda_cla32_fa105_and1;
  wire f_u_dadda_cla32_fa105_or0;
  wire f_u_dadda_cla32_ha18_xor0;
  wire f_u_dadda_cla32_ha18_and0;
  wire f_u_dadda_cla32_fa106_xor0;
  wire f_u_dadda_cla32_fa106_and0;
  wire f_u_dadda_cla32_fa106_xor1;
  wire f_u_dadda_cla32_fa106_and1;
  wire f_u_dadda_cla32_fa106_or0;
  wire f_u_dadda_cla32_fa107_xor0;
  wire f_u_dadda_cla32_fa107_and0;
  wire f_u_dadda_cla32_fa107_xor1;
  wire f_u_dadda_cla32_fa107_and1;
  wire f_u_dadda_cla32_fa107_or0;
  wire f_u_dadda_cla32_fa108_xor0;
  wire f_u_dadda_cla32_fa108_and0;
  wire f_u_dadda_cla32_fa108_xor1;
  wire f_u_dadda_cla32_fa108_and1;
  wire f_u_dadda_cla32_fa108_or0;
  wire f_u_dadda_cla32_fa109_xor0;
  wire f_u_dadda_cla32_fa109_and0;
  wire f_u_dadda_cla32_fa109_xor1;
  wire f_u_dadda_cla32_fa109_and1;
  wire f_u_dadda_cla32_fa109_or0;
  wire f_u_dadda_cla32_and_20_0;
  wire f_u_dadda_cla32_fa110_xor0;
  wire f_u_dadda_cla32_fa110_and0;
  wire f_u_dadda_cla32_fa110_xor1;
  wire f_u_dadda_cla32_fa110_and1;
  wire f_u_dadda_cla32_fa110_or0;
  wire f_u_dadda_cla32_and_19_1;
  wire f_u_dadda_cla32_and_18_2;
  wire f_u_dadda_cla32_and_17_3;
  wire f_u_dadda_cla32_fa111_xor0;
  wire f_u_dadda_cla32_fa111_and0;
  wire f_u_dadda_cla32_fa111_xor1;
  wire f_u_dadda_cla32_fa111_and1;
  wire f_u_dadda_cla32_fa111_or0;
  wire f_u_dadda_cla32_and_16_4;
  wire f_u_dadda_cla32_and_15_5;
  wire f_u_dadda_cla32_and_14_6;
  wire f_u_dadda_cla32_fa112_xor0;
  wire f_u_dadda_cla32_fa112_and0;
  wire f_u_dadda_cla32_fa112_xor1;
  wire f_u_dadda_cla32_fa112_and1;
  wire f_u_dadda_cla32_fa112_or0;
  wire f_u_dadda_cla32_and_13_7;
  wire f_u_dadda_cla32_and_12_8;
  wire f_u_dadda_cla32_and_11_9;
  wire f_u_dadda_cla32_fa113_xor0;
  wire f_u_dadda_cla32_fa113_and0;
  wire f_u_dadda_cla32_fa113_xor1;
  wire f_u_dadda_cla32_fa113_and1;
  wire f_u_dadda_cla32_fa113_or0;
  wire f_u_dadda_cla32_and_10_10;
  wire f_u_dadda_cla32_and_9_11;
  wire f_u_dadda_cla32_and_8_12;
  wire f_u_dadda_cla32_fa114_xor0;
  wire f_u_dadda_cla32_fa114_and0;
  wire f_u_dadda_cla32_fa114_xor1;
  wire f_u_dadda_cla32_fa114_and1;
  wire f_u_dadda_cla32_fa114_or0;
  wire f_u_dadda_cla32_and_7_13;
  wire f_u_dadda_cla32_and_6_14;
  wire f_u_dadda_cla32_and_5_15;
  wire f_u_dadda_cla32_fa115_xor0;
  wire f_u_dadda_cla32_fa115_and0;
  wire f_u_dadda_cla32_fa115_xor1;
  wire f_u_dadda_cla32_fa115_and1;
  wire f_u_dadda_cla32_fa115_or0;
  wire f_u_dadda_cla32_and_4_16;
  wire f_u_dadda_cla32_and_3_17;
  wire f_u_dadda_cla32_and_2_18;
  wire f_u_dadda_cla32_fa116_xor0;
  wire f_u_dadda_cla32_fa116_and0;
  wire f_u_dadda_cla32_fa116_xor1;
  wire f_u_dadda_cla32_fa116_and1;
  wire f_u_dadda_cla32_fa116_or0;
  wire f_u_dadda_cla32_and_1_19;
  wire f_u_dadda_cla32_and_0_20;
  wire f_u_dadda_cla32_fa117_xor0;
  wire f_u_dadda_cla32_fa117_and0;
  wire f_u_dadda_cla32_fa117_xor1;
  wire f_u_dadda_cla32_fa117_and1;
  wire f_u_dadda_cla32_fa117_or0;
  wire f_u_dadda_cla32_fa118_xor0;
  wire f_u_dadda_cla32_fa118_and0;
  wire f_u_dadda_cla32_fa118_xor1;
  wire f_u_dadda_cla32_fa118_and1;
  wire f_u_dadda_cla32_fa118_or0;
  wire f_u_dadda_cla32_fa119_xor0;
  wire f_u_dadda_cla32_fa119_and0;
  wire f_u_dadda_cla32_fa119_xor1;
  wire f_u_dadda_cla32_fa119_and1;
  wire f_u_dadda_cla32_fa119_or0;
  wire f_u_dadda_cla32_ha19_xor0;
  wire f_u_dadda_cla32_ha19_and0;
  wire f_u_dadda_cla32_fa120_xor0;
  wire f_u_dadda_cla32_fa120_and0;
  wire f_u_dadda_cla32_fa120_xor1;
  wire f_u_dadda_cla32_fa120_and1;
  wire f_u_dadda_cla32_fa120_or0;
  wire f_u_dadda_cla32_fa121_xor0;
  wire f_u_dadda_cla32_fa121_and0;
  wire f_u_dadda_cla32_fa121_xor1;
  wire f_u_dadda_cla32_fa121_and1;
  wire f_u_dadda_cla32_fa121_or0;
  wire f_u_dadda_cla32_fa122_xor0;
  wire f_u_dadda_cla32_fa122_and0;
  wire f_u_dadda_cla32_fa122_xor1;
  wire f_u_dadda_cla32_fa122_and1;
  wire f_u_dadda_cla32_fa122_or0;
  wire f_u_dadda_cla32_fa123_xor0;
  wire f_u_dadda_cla32_fa123_and0;
  wire f_u_dadda_cla32_fa123_xor1;
  wire f_u_dadda_cla32_fa123_and1;
  wire f_u_dadda_cla32_fa123_or0;
  wire f_u_dadda_cla32_fa124_xor0;
  wire f_u_dadda_cla32_fa124_and0;
  wire f_u_dadda_cla32_fa124_xor1;
  wire f_u_dadda_cla32_fa124_and1;
  wire f_u_dadda_cla32_fa124_or0;
  wire f_u_dadda_cla32_and_21_0;
  wire f_u_dadda_cla32_and_20_1;
  wire f_u_dadda_cla32_and_19_2;
  wire f_u_dadda_cla32_fa125_xor0;
  wire f_u_dadda_cla32_fa125_and0;
  wire f_u_dadda_cla32_fa125_xor1;
  wire f_u_dadda_cla32_fa125_and1;
  wire f_u_dadda_cla32_fa125_or0;
  wire f_u_dadda_cla32_and_18_3;
  wire f_u_dadda_cla32_and_17_4;
  wire f_u_dadda_cla32_and_16_5;
  wire f_u_dadda_cla32_fa126_xor0;
  wire f_u_dadda_cla32_fa126_and0;
  wire f_u_dadda_cla32_fa126_xor1;
  wire f_u_dadda_cla32_fa126_and1;
  wire f_u_dadda_cla32_fa126_or0;
  wire f_u_dadda_cla32_and_15_6;
  wire f_u_dadda_cla32_and_14_7;
  wire f_u_dadda_cla32_and_13_8;
  wire f_u_dadda_cla32_fa127_xor0;
  wire f_u_dadda_cla32_fa127_and0;
  wire f_u_dadda_cla32_fa127_xor1;
  wire f_u_dadda_cla32_fa127_and1;
  wire f_u_dadda_cla32_fa127_or0;
  wire f_u_dadda_cla32_and_12_9;
  wire f_u_dadda_cla32_and_11_10;
  wire f_u_dadda_cla32_and_10_11;
  wire f_u_dadda_cla32_fa128_xor0;
  wire f_u_dadda_cla32_fa128_and0;
  wire f_u_dadda_cla32_fa128_xor1;
  wire f_u_dadda_cla32_fa128_and1;
  wire f_u_dadda_cla32_fa128_or0;
  wire f_u_dadda_cla32_and_9_12;
  wire f_u_dadda_cla32_and_8_13;
  wire f_u_dadda_cla32_and_7_14;
  wire f_u_dadda_cla32_fa129_xor0;
  wire f_u_dadda_cla32_fa129_and0;
  wire f_u_dadda_cla32_fa129_xor1;
  wire f_u_dadda_cla32_fa129_and1;
  wire f_u_dadda_cla32_fa129_or0;
  wire f_u_dadda_cla32_and_6_15;
  wire f_u_dadda_cla32_and_5_16;
  wire f_u_dadda_cla32_and_4_17;
  wire f_u_dadda_cla32_fa130_xor0;
  wire f_u_dadda_cla32_fa130_and0;
  wire f_u_dadda_cla32_fa130_xor1;
  wire f_u_dadda_cla32_fa130_and1;
  wire f_u_dadda_cla32_fa130_or0;
  wire f_u_dadda_cla32_and_3_18;
  wire f_u_dadda_cla32_and_2_19;
  wire f_u_dadda_cla32_and_1_20;
  wire f_u_dadda_cla32_fa131_xor0;
  wire f_u_dadda_cla32_fa131_and0;
  wire f_u_dadda_cla32_fa131_xor1;
  wire f_u_dadda_cla32_fa131_and1;
  wire f_u_dadda_cla32_fa131_or0;
  wire f_u_dadda_cla32_and_0_21;
  wire f_u_dadda_cla32_fa132_xor0;
  wire f_u_dadda_cla32_fa132_and0;
  wire f_u_dadda_cla32_fa132_xor1;
  wire f_u_dadda_cla32_fa132_and1;
  wire f_u_dadda_cla32_fa132_or0;
  wire f_u_dadda_cla32_fa133_xor0;
  wire f_u_dadda_cla32_fa133_and0;
  wire f_u_dadda_cla32_fa133_xor1;
  wire f_u_dadda_cla32_fa133_and1;
  wire f_u_dadda_cla32_fa133_or0;
  wire f_u_dadda_cla32_fa134_xor0;
  wire f_u_dadda_cla32_fa134_and0;
  wire f_u_dadda_cla32_fa134_xor1;
  wire f_u_dadda_cla32_fa134_and1;
  wire f_u_dadda_cla32_fa134_or0;
  wire f_u_dadda_cla32_ha20_xor0;
  wire f_u_dadda_cla32_ha20_and0;
  wire f_u_dadda_cla32_fa135_xor0;
  wire f_u_dadda_cla32_fa135_and0;
  wire f_u_dadda_cla32_fa135_xor1;
  wire f_u_dadda_cla32_fa135_and1;
  wire f_u_dadda_cla32_fa135_or0;
  wire f_u_dadda_cla32_fa136_xor0;
  wire f_u_dadda_cla32_fa136_and0;
  wire f_u_dadda_cla32_fa136_xor1;
  wire f_u_dadda_cla32_fa136_and1;
  wire f_u_dadda_cla32_fa136_or0;
  wire f_u_dadda_cla32_fa137_xor0;
  wire f_u_dadda_cla32_fa137_and0;
  wire f_u_dadda_cla32_fa137_xor1;
  wire f_u_dadda_cla32_fa137_and1;
  wire f_u_dadda_cla32_fa137_or0;
  wire f_u_dadda_cla32_fa138_xor0;
  wire f_u_dadda_cla32_fa138_and0;
  wire f_u_dadda_cla32_fa138_xor1;
  wire f_u_dadda_cla32_fa138_and1;
  wire f_u_dadda_cla32_fa138_or0;
  wire f_u_dadda_cla32_fa139_xor0;
  wire f_u_dadda_cla32_fa139_and0;
  wire f_u_dadda_cla32_fa139_xor1;
  wire f_u_dadda_cla32_fa139_and1;
  wire f_u_dadda_cla32_fa139_or0;
  wire f_u_dadda_cla32_and_22_0;
  wire f_u_dadda_cla32_and_21_1;
  wire f_u_dadda_cla32_fa140_xor0;
  wire f_u_dadda_cla32_fa140_and0;
  wire f_u_dadda_cla32_fa140_xor1;
  wire f_u_dadda_cla32_fa140_and1;
  wire f_u_dadda_cla32_fa140_or0;
  wire f_u_dadda_cla32_and_20_2;
  wire f_u_dadda_cla32_and_19_3;
  wire f_u_dadda_cla32_and_18_4;
  wire f_u_dadda_cla32_fa141_xor0;
  wire f_u_dadda_cla32_fa141_and0;
  wire f_u_dadda_cla32_fa141_xor1;
  wire f_u_dadda_cla32_fa141_and1;
  wire f_u_dadda_cla32_fa141_or0;
  wire f_u_dadda_cla32_and_17_5;
  wire f_u_dadda_cla32_and_16_6;
  wire f_u_dadda_cla32_and_15_7;
  wire f_u_dadda_cla32_fa142_xor0;
  wire f_u_dadda_cla32_fa142_and0;
  wire f_u_dadda_cla32_fa142_xor1;
  wire f_u_dadda_cla32_fa142_and1;
  wire f_u_dadda_cla32_fa142_or0;
  wire f_u_dadda_cla32_and_14_8;
  wire f_u_dadda_cla32_and_13_9;
  wire f_u_dadda_cla32_and_12_10;
  wire f_u_dadda_cla32_fa143_xor0;
  wire f_u_dadda_cla32_fa143_and0;
  wire f_u_dadda_cla32_fa143_xor1;
  wire f_u_dadda_cla32_fa143_and1;
  wire f_u_dadda_cla32_fa143_or0;
  wire f_u_dadda_cla32_and_11_11;
  wire f_u_dadda_cla32_and_10_12;
  wire f_u_dadda_cla32_and_9_13;
  wire f_u_dadda_cla32_fa144_xor0;
  wire f_u_dadda_cla32_fa144_and0;
  wire f_u_dadda_cla32_fa144_xor1;
  wire f_u_dadda_cla32_fa144_and1;
  wire f_u_dadda_cla32_fa144_or0;
  wire f_u_dadda_cla32_and_8_14;
  wire f_u_dadda_cla32_and_7_15;
  wire f_u_dadda_cla32_and_6_16;
  wire f_u_dadda_cla32_fa145_xor0;
  wire f_u_dadda_cla32_fa145_and0;
  wire f_u_dadda_cla32_fa145_xor1;
  wire f_u_dadda_cla32_fa145_and1;
  wire f_u_dadda_cla32_fa145_or0;
  wire f_u_dadda_cla32_and_5_17;
  wire f_u_dadda_cla32_and_4_18;
  wire f_u_dadda_cla32_and_3_19;
  wire f_u_dadda_cla32_fa146_xor0;
  wire f_u_dadda_cla32_fa146_and0;
  wire f_u_dadda_cla32_fa146_xor1;
  wire f_u_dadda_cla32_fa146_and1;
  wire f_u_dadda_cla32_fa146_or0;
  wire f_u_dadda_cla32_and_2_20;
  wire f_u_dadda_cla32_and_1_21;
  wire f_u_dadda_cla32_and_0_22;
  wire f_u_dadda_cla32_fa147_xor0;
  wire f_u_dadda_cla32_fa147_and0;
  wire f_u_dadda_cla32_fa147_xor1;
  wire f_u_dadda_cla32_fa147_and1;
  wire f_u_dadda_cla32_fa147_or0;
  wire f_u_dadda_cla32_fa148_xor0;
  wire f_u_dadda_cla32_fa148_and0;
  wire f_u_dadda_cla32_fa148_xor1;
  wire f_u_dadda_cla32_fa148_and1;
  wire f_u_dadda_cla32_fa148_or0;
  wire f_u_dadda_cla32_fa149_xor0;
  wire f_u_dadda_cla32_fa149_and0;
  wire f_u_dadda_cla32_fa149_xor1;
  wire f_u_dadda_cla32_fa149_and1;
  wire f_u_dadda_cla32_fa149_or0;
  wire f_u_dadda_cla32_fa150_xor0;
  wire f_u_dadda_cla32_fa150_and0;
  wire f_u_dadda_cla32_fa150_xor1;
  wire f_u_dadda_cla32_fa150_and1;
  wire f_u_dadda_cla32_fa150_or0;
  wire f_u_dadda_cla32_ha21_xor0;
  wire f_u_dadda_cla32_ha21_and0;
  wire f_u_dadda_cla32_fa151_xor0;
  wire f_u_dadda_cla32_fa151_and0;
  wire f_u_dadda_cla32_fa151_xor1;
  wire f_u_dadda_cla32_fa151_and1;
  wire f_u_dadda_cla32_fa151_or0;
  wire f_u_dadda_cla32_fa152_xor0;
  wire f_u_dadda_cla32_fa152_and0;
  wire f_u_dadda_cla32_fa152_xor1;
  wire f_u_dadda_cla32_fa152_and1;
  wire f_u_dadda_cla32_fa152_or0;
  wire f_u_dadda_cla32_fa153_xor0;
  wire f_u_dadda_cla32_fa153_and0;
  wire f_u_dadda_cla32_fa153_xor1;
  wire f_u_dadda_cla32_fa153_and1;
  wire f_u_dadda_cla32_fa153_or0;
  wire f_u_dadda_cla32_fa154_xor0;
  wire f_u_dadda_cla32_fa154_and0;
  wire f_u_dadda_cla32_fa154_xor1;
  wire f_u_dadda_cla32_fa154_and1;
  wire f_u_dadda_cla32_fa154_or0;
  wire f_u_dadda_cla32_fa155_xor0;
  wire f_u_dadda_cla32_fa155_and0;
  wire f_u_dadda_cla32_fa155_xor1;
  wire f_u_dadda_cla32_fa155_and1;
  wire f_u_dadda_cla32_fa155_or0;
  wire f_u_dadda_cla32_and_23_0;
  wire f_u_dadda_cla32_fa156_xor0;
  wire f_u_dadda_cla32_fa156_and0;
  wire f_u_dadda_cla32_fa156_xor1;
  wire f_u_dadda_cla32_fa156_and1;
  wire f_u_dadda_cla32_fa156_or0;
  wire f_u_dadda_cla32_and_22_1;
  wire f_u_dadda_cla32_and_21_2;
  wire f_u_dadda_cla32_and_20_3;
  wire f_u_dadda_cla32_fa157_xor0;
  wire f_u_dadda_cla32_fa157_and0;
  wire f_u_dadda_cla32_fa157_xor1;
  wire f_u_dadda_cla32_fa157_and1;
  wire f_u_dadda_cla32_fa157_or0;
  wire f_u_dadda_cla32_and_19_4;
  wire f_u_dadda_cla32_and_18_5;
  wire f_u_dadda_cla32_and_17_6;
  wire f_u_dadda_cla32_fa158_xor0;
  wire f_u_dadda_cla32_fa158_and0;
  wire f_u_dadda_cla32_fa158_xor1;
  wire f_u_dadda_cla32_fa158_and1;
  wire f_u_dadda_cla32_fa158_or0;
  wire f_u_dadda_cla32_and_16_7;
  wire f_u_dadda_cla32_and_15_8;
  wire f_u_dadda_cla32_and_14_9;
  wire f_u_dadda_cla32_fa159_xor0;
  wire f_u_dadda_cla32_fa159_and0;
  wire f_u_dadda_cla32_fa159_xor1;
  wire f_u_dadda_cla32_fa159_and1;
  wire f_u_dadda_cla32_fa159_or0;
  wire f_u_dadda_cla32_and_13_10;
  wire f_u_dadda_cla32_and_12_11;
  wire f_u_dadda_cla32_and_11_12;
  wire f_u_dadda_cla32_fa160_xor0;
  wire f_u_dadda_cla32_fa160_and0;
  wire f_u_dadda_cla32_fa160_xor1;
  wire f_u_dadda_cla32_fa160_and1;
  wire f_u_dadda_cla32_fa160_or0;
  wire f_u_dadda_cla32_and_10_13;
  wire f_u_dadda_cla32_and_9_14;
  wire f_u_dadda_cla32_and_8_15;
  wire f_u_dadda_cla32_fa161_xor0;
  wire f_u_dadda_cla32_fa161_and0;
  wire f_u_dadda_cla32_fa161_xor1;
  wire f_u_dadda_cla32_fa161_and1;
  wire f_u_dadda_cla32_fa161_or0;
  wire f_u_dadda_cla32_and_7_16;
  wire f_u_dadda_cla32_and_6_17;
  wire f_u_dadda_cla32_and_5_18;
  wire f_u_dadda_cla32_fa162_xor0;
  wire f_u_dadda_cla32_fa162_and0;
  wire f_u_dadda_cla32_fa162_xor1;
  wire f_u_dadda_cla32_fa162_and1;
  wire f_u_dadda_cla32_fa162_or0;
  wire f_u_dadda_cla32_and_4_19;
  wire f_u_dadda_cla32_and_3_20;
  wire f_u_dadda_cla32_and_2_21;
  wire f_u_dadda_cla32_fa163_xor0;
  wire f_u_dadda_cla32_fa163_and0;
  wire f_u_dadda_cla32_fa163_xor1;
  wire f_u_dadda_cla32_fa163_and1;
  wire f_u_dadda_cla32_fa163_or0;
  wire f_u_dadda_cla32_and_1_22;
  wire f_u_dadda_cla32_and_0_23;
  wire f_u_dadda_cla32_fa164_xor0;
  wire f_u_dadda_cla32_fa164_and0;
  wire f_u_dadda_cla32_fa164_xor1;
  wire f_u_dadda_cla32_fa164_and1;
  wire f_u_dadda_cla32_fa164_or0;
  wire f_u_dadda_cla32_fa165_xor0;
  wire f_u_dadda_cla32_fa165_and0;
  wire f_u_dadda_cla32_fa165_xor1;
  wire f_u_dadda_cla32_fa165_and1;
  wire f_u_dadda_cla32_fa165_or0;
  wire f_u_dadda_cla32_fa166_xor0;
  wire f_u_dadda_cla32_fa166_and0;
  wire f_u_dadda_cla32_fa166_xor1;
  wire f_u_dadda_cla32_fa166_and1;
  wire f_u_dadda_cla32_fa166_or0;
  wire f_u_dadda_cla32_fa167_xor0;
  wire f_u_dadda_cla32_fa167_and0;
  wire f_u_dadda_cla32_fa167_xor1;
  wire f_u_dadda_cla32_fa167_and1;
  wire f_u_dadda_cla32_fa167_or0;
  wire f_u_dadda_cla32_ha22_xor0;
  wire f_u_dadda_cla32_ha22_and0;
  wire f_u_dadda_cla32_fa168_xor0;
  wire f_u_dadda_cla32_fa168_and0;
  wire f_u_dadda_cla32_fa168_xor1;
  wire f_u_dadda_cla32_fa168_and1;
  wire f_u_dadda_cla32_fa168_or0;
  wire f_u_dadda_cla32_fa169_xor0;
  wire f_u_dadda_cla32_fa169_and0;
  wire f_u_dadda_cla32_fa169_xor1;
  wire f_u_dadda_cla32_fa169_and1;
  wire f_u_dadda_cla32_fa169_or0;
  wire f_u_dadda_cla32_fa170_xor0;
  wire f_u_dadda_cla32_fa170_and0;
  wire f_u_dadda_cla32_fa170_xor1;
  wire f_u_dadda_cla32_fa170_and1;
  wire f_u_dadda_cla32_fa170_or0;
  wire f_u_dadda_cla32_fa171_xor0;
  wire f_u_dadda_cla32_fa171_and0;
  wire f_u_dadda_cla32_fa171_xor1;
  wire f_u_dadda_cla32_fa171_and1;
  wire f_u_dadda_cla32_fa171_or0;
  wire f_u_dadda_cla32_fa172_xor0;
  wire f_u_dadda_cla32_fa172_and0;
  wire f_u_dadda_cla32_fa172_xor1;
  wire f_u_dadda_cla32_fa172_and1;
  wire f_u_dadda_cla32_fa172_or0;
  wire f_u_dadda_cla32_fa173_xor0;
  wire f_u_dadda_cla32_fa173_and0;
  wire f_u_dadda_cla32_fa173_xor1;
  wire f_u_dadda_cla32_fa173_and1;
  wire f_u_dadda_cla32_fa173_or0;
  wire f_u_dadda_cla32_and_24_0;
  wire f_u_dadda_cla32_and_23_1;
  wire f_u_dadda_cla32_and_22_2;
  wire f_u_dadda_cla32_fa174_xor0;
  wire f_u_dadda_cla32_fa174_and0;
  wire f_u_dadda_cla32_fa174_xor1;
  wire f_u_dadda_cla32_fa174_and1;
  wire f_u_dadda_cla32_fa174_or0;
  wire f_u_dadda_cla32_and_21_3;
  wire f_u_dadda_cla32_and_20_4;
  wire f_u_dadda_cla32_and_19_5;
  wire f_u_dadda_cla32_fa175_xor0;
  wire f_u_dadda_cla32_fa175_and0;
  wire f_u_dadda_cla32_fa175_xor1;
  wire f_u_dadda_cla32_fa175_and1;
  wire f_u_dadda_cla32_fa175_or0;
  wire f_u_dadda_cla32_and_18_6;
  wire f_u_dadda_cla32_and_17_7;
  wire f_u_dadda_cla32_and_16_8;
  wire f_u_dadda_cla32_fa176_xor0;
  wire f_u_dadda_cla32_fa176_and0;
  wire f_u_dadda_cla32_fa176_xor1;
  wire f_u_dadda_cla32_fa176_and1;
  wire f_u_dadda_cla32_fa176_or0;
  wire f_u_dadda_cla32_and_15_9;
  wire f_u_dadda_cla32_and_14_10;
  wire f_u_dadda_cla32_and_13_11;
  wire f_u_dadda_cla32_fa177_xor0;
  wire f_u_dadda_cla32_fa177_and0;
  wire f_u_dadda_cla32_fa177_xor1;
  wire f_u_dadda_cla32_fa177_and1;
  wire f_u_dadda_cla32_fa177_or0;
  wire f_u_dadda_cla32_and_12_12;
  wire f_u_dadda_cla32_and_11_13;
  wire f_u_dadda_cla32_and_10_14;
  wire f_u_dadda_cla32_fa178_xor0;
  wire f_u_dadda_cla32_fa178_and0;
  wire f_u_dadda_cla32_fa178_xor1;
  wire f_u_dadda_cla32_fa178_and1;
  wire f_u_dadda_cla32_fa178_or0;
  wire f_u_dadda_cla32_and_9_15;
  wire f_u_dadda_cla32_and_8_16;
  wire f_u_dadda_cla32_and_7_17;
  wire f_u_dadda_cla32_fa179_xor0;
  wire f_u_dadda_cla32_fa179_and0;
  wire f_u_dadda_cla32_fa179_xor1;
  wire f_u_dadda_cla32_fa179_and1;
  wire f_u_dadda_cla32_fa179_or0;
  wire f_u_dadda_cla32_and_6_18;
  wire f_u_dadda_cla32_and_5_19;
  wire f_u_dadda_cla32_and_4_20;
  wire f_u_dadda_cla32_fa180_xor0;
  wire f_u_dadda_cla32_fa180_and0;
  wire f_u_dadda_cla32_fa180_xor1;
  wire f_u_dadda_cla32_fa180_and1;
  wire f_u_dadda_cla32_fa180_or0;
  wire f_u_dadda_cla32_and_3_21;
  wire f_u_dadda_cla32_and_2_22;
  wire f_u_dadda_cla32_and_1_23;
  wire f_u_dadda_cla32_fa181_xor0;
  wire f_u_dadda_cla32_fa181_and0;
  wire f_u_dadda_cla32_fa181_xor1;
  wire f_u_dadda_cla32_fa181_and1;
  wire f_u_dadda_cla32_fa181_or0;
  wire f_u_dadda_cla32_and_0_24;
  wire f_u_dadda_cla32_fa182_xor0;
  wire f_u_dadda_cla32_fa182_and0;
  wire f_u_dadda_cla32_fa182_xor1;
  wire f_u_dadda_cla32_fa182_and1;
  wire f_u_dadda_cla32_fa182_or0;
  wire f_u_dadda_cla32_fa183_xor0;
  wire f_u_dadda_cla32_fa183_and0;
  wire f_u_dadda_cla32_fa183_xor1;
  wire f_u_dadda_cla32_fa183_and1;
  wire f_u_dadda_cla32_fa183_or0;
  wire f_u_dadda_cla32_fa184_xor0;
  wire f_u_dadda_cla32_fa184_and0;
  wire f_u_dadda_cla32_fa184_xor1;
  wire f_u_dadda_cla32_fa184_and1;
  wire f_u_dadda_cla32_fa184_or0;
  wire f_u_dadda_cla32_fa185_xor0;
  wire f_u_dadda_cla32_fa185_and0;
  wire f_u_dadda_cla32_fa185_xor1;
  wire f_u_dadda_cla32_fa185_and1;
  wire f_u_dadda_cla32_fa185_or0;
  wire f_u_dadda_cla32_ha23_xor0;
  wire f_u_dadda_cla32_ha23_and0;
  wire f_u_dadda_cla32_fa186_xor0;
  wire f_u_dadda_cla32_fa186_and0;
  wire f_u_dadda_cla32_fa186_xor1;
  wire f_u_dadda_cla32_fa186_and1;
  wire f_u_dadda_cla32_fa186_or0;
  wire f_u_dadda_cla32_fa187_xor0;
  wire f_u_dadda_cla32_fa187_and0;
  wire f_u_dadda_cla32_fa187_xor1;
  wire f_u_dadda_cla32_fa187_and1;
  wire f_u_dadda_cla32_fa187_or0;
  wire f_u_dadda_cla32_fa188_xor0;
  wire f_u_dadda_cla32_fa188_and0;
  wire f_u_dadda_cla32_fa188_xor1;
  wire f_u_dadda_cla32_fa188_and1;
  wire f_u_dadda_cla32_fa188_or0;
  wire f_u_dadda_cla32_fa189_xor0;
  wire f_u_dadda_cla32_fa189_and0;
  wire f_u_dadda_cla32_fa189_xor1;
  wire f_u_dadda_cla32_fa189_and1;
  wire f_u_dadda_cla32_fa189_or0;
  wire f_u_dadda_cla32_fa190_xor0;
  wire f_u_dadda_cla32_fa190_and0;
  wire f_u_dadda_cla32_fa190_xor1;
  wire f_u_dadda_cla32_fa190_and1;
  wire f_u_dadda_cla32_fa190_or0;
  wire f_u_dadda_cla32_fa191_xor0;
  wire f_u_dadda_cla32_fa191_and0;
  wire f_u_dadda_cla32_fa191_xor1;
  wire f_u_dadda_cla32_fa191_and1;
  wire f_u_dadda_cla32_fa191_or0;
  wire f_u_dadda_cla32_and_25_0;
  wire f_u_dadda_cla32_and_24_1;
  wire f_u_dadda_cla32_fa192_xor0;
  wire f_u_dadda_cla32_fa192_and0;
  wire f_u_dadda_cla32_fa192_xor1;
  wire f_u_dadda_cla32_fa192_and1;
  wire f_u_dadda_cla32_fa192_or0;
  wire f_u_dadda_cla32_and_23_2;
  wire f_u_dadda_cla32_and_22_3;
  wire f_u_dadda_cla32_and_21_4;
  wire f_u_dadda_cla32_fa193_xor0;
  wire f_u_dadda_cla32_fa193_and0;
  wire f_u_dadda_cla32_fa193_xor1;
  wire f_u_dadda_cla32_fa193_and1;
  wire f_u_dadda_cla32_fa193_or0;
  wire f_u_dadda_cla32_and_20_5;
  wire f_u_dadda_cla32_and_19_6;
  wire f_u_dadda_cla32_and_18_7;
  wire f_u_dadda_cla32_fa194_xor0;
  wire f_u_dadda_cla32_fa194_and0;
  wire f_u_dadda_cla32_fa194_xor1;
  wire f_u_dadda_cla32_fa194_and1;
  wire f_u_dadda_cla32_fa194_or0;
  wire f_u_dadda_cla32_and_17_8;
  wire f_u_dadda_cla32_and_16_9;
  wire f_u_dadda_cla32_and_15_10;
  wire f_u_dadda_cla32_fa195_xor0;
  wire f_u_dadda_cla32_fa195_and0;
  wire f_u_dadda_cla32_fa195_xor1;
  wire f_u_dadda_cla32_fa195_and1;
  wire f_u_dadda_cla32_fa195_or0;
  wire f_u_dadda_cla32_and_14_11;
  wire f_u_dadda_cla32_and_13_12;
  wire f_u_dadda_cla32_and_12_13;
  wire f_u_dadda_cla32_fa196_xor0;
  wire f_u_dadda_cla32_fa196_and0;
  wire f_u_dadda_cla32_fa196_xor1;
  wire f_u_dadda_cla32_fa196_and1;
  wire f_u_dadda_cla32_fa196_or0;
  wire f_u_dadda_cla32_and_11_14;
  wire f_u_dadda_cla32_and_10_15;
  wire f_u_dadda_cla32_and_9_16;
  wire f_u_dadda_cla32_fa197_xor0;
  wire f_u_dadda_cla32_fa197_and0;
  wire f_u_dadda_cla32_fa197_xor1;
  wire f_u_dadda_cla32_fa197_and1;
  wire f_u_dadda_cla32_fa197_or0;
  wire f_u_dadda_cla32_and_8_17;
  wire f_u_dadda_cla32_and_7_18;
  wire f_u_dadda_cla32_and_6_19;
  wire f_u_dadda_cla32_fa198_xor0;
  wire f_u_dadda_cla32_fa198_and0;
  wire f_u_dadda_cla32_fa198_xor1;
  wire f_u_dadda_cla32_fa198_and1;
  wire f_u_dadda_cla32_fa198_or0;
  wire f_u_dadda_cla32_and_5_20;
  wire f_u_dadda_cla32_and_4_21;
  wire f_u_dadda_cla32_and_3_22;
  wire f_u_dadda_cla32_fa199_xor0;
  wire f_u_dadda_cla32_fa199_and0;
  wire f_u_dadda_cla32_fa199_xor1;
  wire f_u_dadda_cla32_fa199_and1;
  wire f_u_dadda_cla32_fa199_or0;
  wire f_u_dadda_cla32_and_2_23;
  wire f_u_dadda_cla32_and_1_24;
  wire f_u_dadda_cla32_and_0_25;
  wire f_u_dadda_cla32_fa200_xor0;
  wire f_u_dadda_cla32_fa200_and0;
  wire f_u_dadda_cla32_fa200_xor1;
  wire f_u_dadda_cla32_fa200_and1;
  wire f_u_dadda_cla32_fa200_or0;
  wire f_u_dadda_cla32_fa201_xor0;
  wire f_u_dadda_cla32_fa201_and0;
  wire f_u_dadda_cla32_fa201_xor1;
  wire f_u_dadda_cla32_fa201_and1;
  wire f_u_dadda_cla32_fa201_or0;
  wire f_u_dadda_cla32_fa202_xor0;
  wire f_u_dadda_cla32_fa202_and0;
  wire f_u_dadda_cla32_fa202_xor1;
  wire f_u_dadda_cla32_fa202_and1;
  wire f_u_dadda_cla32_fa202_or0;
  wire f_u_dadda_cla32_fa203_xor0;
  wire f_u_dadda_cla32_fa203_and0;
  wire f_u_dadda_cla32_fa203_xor1;
  wire f_u_dadda_cla32_fa203_and1;
  wire f_u_dadda_cla32_fa203_or0;
  wire f_u_dadda_cla32_fa204_xor0;
  wire f_u_dadda_cla32_fa204_and0;
  wire f_u_dadda_cla32_fa204_xor1;
  wire f_u_dadda_cla32_fa204_and1;
  wire f_u_dadda_cla32_fa204_or0;
  wire f_u_dadda_cla32_ha24_xor0;
  wire f_u_dadda_cla32_ha24_and0;
  wire f_u_dadda_cla32_fa205_xor0;
  wire f_u_dadda_cla32_fa205_and0;
  wire f_u_dadda_cla32_fa205_xor1;
  wire f_u_dadda_cla32_fa205_and1;
  wire f_u_dadda_cla32_fa205_or0;
  wire f_u_dadda_cla32_fa206_xor0;
  wire f_u_dadda_cla32_fa206_and0;
  wire f_u_dadda_cla32_fa206_xor1;
  wire f_u_dadda_cla32_fa206_and1;
  wire f_u_dadda_cla32_fa206_or0;
  wire f_u_dadda_cla32_fa207_xor0;
  wire f_u_dadda_cla32_fa207_and0;
  wire f_u_dadda_cla32_fa207_xor1;
  wire f_u_dadda_cla32_fa207_and1;
  wire f_u_dadda_cla32_fa207_or0;
  wire f_u_dadda_cla32_fa208_xor0;
  wire f_u_dadda_cla32_fa208_and0;
  wire f_u_dadda_cla32_fa208_xor1;
  wire f_u_dadda_cla32_fa208_and1;
  wire f_u_dadda_cla32_fa208_or0;
  wire f_u_dadda_cla32_fa209_xor0;
  wire f_u_dadda_cla32_fa209_and0;
  wire f_u_dadda_cla32_fa209_xor1;
  wire f_u_dadda_cla32_fa209_and1;
  wire f_u_dadda_cla32_fa209_or0;
  wire f_u_dadda_cla32_fa210_xor0;
  wire f_u_dadda_cla32_fa210_and0;
  wire f_u_dadda_cla32_fa210_xor1;
  wire f_u_dadda_cla32_fa210_and1;
  wire f_u_dadda_cla32_fa210_or0;
  wire f_u_dadda_cla32_and_26_0;
  wire f_u_dadda_cla32_fa211_xor0;
  wire f_u_dadda_cla32_fa211_and0;
  wire f_u_dadda_cla32_fa211_xor1;
  wire f_u_dadda_cla32_fa211_and1;
  wire f_u_dadda_cla32_fa211_or0;
  wire f_u_dadda_cla32_and_25_1;
  wire f_u_dadda_cla32_and_24_2;
  wire f_u_dadda_cla32_and_23_3;
  wire f_u_dadda_cla32_fa212_xor0;
  wire f_u_dadda_cla32_fa212_and0;
  wire f_u_dadda_cla32_fa212_xor1;
  wire f_u_dadda_cla32_fa212_and1;
  wire f_u_dadda_cla32_fa212_or0;
  wire f_u_dadda_cla32_and_22_4;
  wire f_u_dadda_cla32_and_21_5;
  wire f_u_dadda_cla32_and_20_6;
  wire f_u_dadda_cla32_fa213_xor0;
  wire f_u_dadda_cla32_fa213_and0;
  wire f_u_dadda_cla32_fa213_xor1;
  wire f_u_dadda_cla32_fa213_and1;
  wire f_u_dadda_cla32_fa213_or0;
  wire f_u_dadda_cla32_and_19_7;
  wire f_u_dadda_cla32_and_18_8;
  wire f_u_dadda_cla32_and_17_9;
  wire f_u_dadda_cla32_fa214_xor0;
  wire f_u_dadda_cla32_fa214_and0;
  wire f_u_dadda_cla32_fa214_xor1;
  wire f_u_dadda_cla32_fa214_and1;
  wire f_u_dadda_cla32_fa214_or0;
  wire f_u_dadda_cla32_and_16_10;
  wire f_u_dadda_cla32_and_15_11;
  wire f_u_dadda_cla32_and_14_12;
  wire f_u_dadda_cla32_fa215_xor0;
  wire f_u_dadda_cla32_fa215_and0;
  wire f_u_dadda_cla32_fa215_xor1;
  wire f_u_dadda_cla32_fa215_and1;
  wire f_u_dadda_cla32_fa215_or0;
  wire f_u_dadda_cla32_and_13_13;
  wire f_u_dadda_cla32_and_12_14;
  wire f_u_dadda_cla32_and_11_15;
  wire f_u_dadda_cla32_fa216_xor0;
  wire f_u_dadda_cla32_fa216_and0;
  wire f_u_dadda_cla32_fa216_xor1;
  wire f_u_dadda_cla32_fa216_and1;
  wire f_u_dadda_cla32_fa216_or0;
  wire f_u_dadda_cla32_and_10_16;
  wire f_u_dadda_cla32_and_9_17;
  wire f_u_dadda_cla32_and_8_18;
  wire f_u_dadda_cla32_fa217_xor0;
  wire f_u_dadda_cla32_fa217_and0;
  wire f_u_dadda_cla32_fa217_xor1;
  wire f_u_dadda_cla32_fa217_and1;
  wire f_u_dadda_cla32_fa217_or0;
  wire f_u_dadda_cla32_and_7_19;
  wire f_u_dadda_cla32_and_6_20;
  wire f_u_dadda_cla32_and_5_21;
  wire f_u_dadda_cla32_fa218_xor0;
  wire f_u_dadda_cla32_fa218_and0;
  wire f_u_dadda_cla32_fa218_xor1;
  wire f_u_dadda_cla32_fa218_and1;
  wire f_u_dadda_cla32_fa218_or0;
  wire f_u_dadda_cla32_and_4_22;
  wire f_u_dadda_cla32_and_3_23;
  wire f_u_dadda_cla32_and_2_24;
  wire f_u_dadda_cla32_fa219_xor0;
  wire f_u_dadda_cla32_fa219_and0;
  wire f_u_dadda_cla32_fa219_xor1;
  wire f_u_dadda_cla32_fa219_and1;
  wire f_u_dadda_cla32_fa219_or0;
  wire f_u_dadda_cla32_and_1_25;
  wire f_u_dadda_cla32_and_0_26;
  wire f_u_dadda_cla32_fa220_xor0;
  wire f_u_dadda_cla32_fa220_and0;
  wire f_u_dadda_cla32_fa220_xor1;
  wire f_u_dadda_cla32_fa220_and1;
  wire f_u_dadda_cla32_fa220_or0;
  wire f_u_dadda_cla32_fa221_xor0;
  wire f_u_dadda_cla32_fa221_and0;
  wire f_u_dadda_cla32_fa221_xor1;
  wire f_u_dadda_cla32_fa221_and1;
  wire f_u_dadda_cla32_fa221_or0;
  wire f_u_dadda_cla32_fa222_xor0;
  wire f_u_dadda_cla32_fa222_and0;
  wire f_u_dadda_cla32_fa222_xor1;
  wire f_u_dadda_cla32_fa222_and1;
  wire f_u_dadda_cla32_fa222_or0;
  wire f_u_dadda_cla32_fa223_xor0;
  wire f_u_dadda_cla32_fa223_and0;
  wire f_u_dadda_cla32_fa223_xor1;
  wire f_u_dadda_cla32_fa223_and1;
  wire f_u_dadda_cla32_fa223_or0;
  wire f_u_dadda_cla32_fa224_xor0;
  wire f_u_dadda_cla32_fa224_and0;
  wire f_u_dadda_cla32_fa224_xor1;
  wire f_u_dadda_cla32_fa224_and1;
  wire f_u_dadda_cla32_fa224_or0;
  wire f_u_dadda_cla32_ha25_xor0;
  wire f_u_dadda_cla32_ha25_and0;
  wire f_u_dadda_cla32_fa225_xor0;
  wire f_u_dadda_cla32_fa225_and0;
  wire f_u_dadda_cla32_fa225_xor1;
  wire f_u_dadda_cla32_fa225_and1;
  wire f_u_dadda_cla32_fa225_or0;
  wire f_u_dadda_cla32_fa226_xor0;
  wire f_u_dadda_cla32_fa226_and0;
  wire f_u_dadda_cla32_fa226_xor1;
  wire f_u_dadda_cla32_fa226_and1;
  wire f_u_dadda_cla32_fa226_or0;
  wire f_u_dadda_cla32_fa227_xor0;
  wire f_u_dadda_cla32_fa227_and0;
  wire f_u_dadda_cla32_fa227_xor1;
  wire f_u_dadda_cla32_fa227_and1;
  wire f_u_dadda_cla32_fa227_or0;
  wire f_u_dadda_cla32_fa228_xor0;
  wire f_u_dadda_cla32_fa228_and0;
  wire f_u_dadda_cla32_fa228_xor1;
  wire f_u_dadda_cla32_fa228_and1;
  wire f_u_dadda_cla32_fa228_or0;
  wire f_u_dadda_cla32_fa229_xor0;
  wire f_u_dadda_cla32_fa229_and0;
  wire f_u_dadda_cla32_fa229_xor1;
  wire f_u_dadda_cla32_fa229_and1;
  wire f_u_dadda_cla32_fa229_or0;
  wire f_u_dadda_cla32_fa230_xor0;
  wire f_u_dadda_cla32_fa230_and0;
  wire f_u_dadda_cla32_fa230_xor1;
  wire f_u_dadda_cla32_fa230_and1;
  wire f_u_dadda_cla32_fa230_or0;
  wire f_u_dadda_cla32_fa231_xor0;
  wire f_u_dadda_cla32_fa231_and0;
  wire f_u_dadda_cla32_fa231_xor1;
  wire f_u_dadda_cla32_fa231_and1;
  wire f_u_dadda_cla32_fa231_or0;
  wire f_u_dadda_cla32_and_27_0;
  wire f_u_dadda_cla32_and_26_1;
  wire f_u_dadda_cla32_and_25_2;
  wire f_u_dadda_cla32_fa232_xor0;
  wire f_u_dadda_cla32_fa232_and0;
  wire f_u_dadda_cla32_fa232_xor1;
  wire f_u_dadda_cla32_fa232_and1;
  wire f_u_dadda_cla32_fa232_or0;
  wire f_u_dadda_cla32_and_24_3;
  wire f_u_dadda_cla32_and_23_4;
  wire f_u_dadda_cla32_and_22_5;
  wire f_u_dadda_cla32_fa233_xor0;
  wire f_u_dadda_cla32_fa233_and0;
  wire f_u_dadda_cla32_fa233_xor1;
  wire f_u_dadda_cla32_fa233_and1;
  wire f_u_dadda_cla32_fa233_or0;
  wire f_u_dadda_cla32_and_21_6;
  wire f_u_dadda_cla32_and_20_7;
  wire f_u_dadda_cla32_and_19_8;
  wire f_u_dadda_cla32_fa234_xor0;
  wire f_u_dadda_cla32_fa234_and0;
  wire f_u_dadda_cla32_fa234_xor1;
  wire f_u_dadda_cla32_fa234_and1;
  wire f_u_dadda_cla32_fa234_or0;
  wire f_u_dadda_cla32_and_18_9;
  wire f_u_dadda_cla32_and_17_10;
  wire f_u_dadda_cla32_and_16_11;
  wire f_u_dadda_cla32_fa235_xor0;
  wire f_u_dadda_cla32_fa235_and0;
  wire f_u_dadda_cla32_fa235_xor1;
  wire f_u_dadda_cla32_fa235_and1;
  wire f_u_dadda_cla32_fa235_or0;
  wire f_u_dadda_cla32_and_15_12;
  wire f_u_dadda_cla32_and_14_13;
  wire f_u_dadda_cla32_and_13_14;
  wire f_u_dadda_cla32_fa236_xor0;
  wire f_u_dadda_cla32_fa236_and0;
  wire f_u_dadda_cla32_fa236_xor1;
  wire f_u_dadda_cla32_fa236_and1;
  wire f_u_dadda_cla32_fa236_or0;
  wire f_u_dadda_cla32_and_12_15;
  wire f_u_dadda_cla32_and_11_16;
  wire f_u_dadda_cla32_and_10_17;
  wire f_u_dadda_cla32_fa237_xor0;
  wire f_u_dadda_cla32_fa237_and0;
  wire f_u_dadda_cla32_fa237_xor1;
  wire f_u_dadda_cla32_fa237_and1;
  wire f_u_dadda_cla32_fa237_or0;
  wire f_u_dadda_cla32_and_9_18;
  wire f_u_dadda_cla32_and_8_19;
  wire f_u_dadda_cla32_and_7_20;
  wire f_u_dadda_cla32_fa238_xor0;
  wire f_u_dadda_cla32_fa238_and0;
  wire f_u_dadda_cla32_fa238_xor1;
  wire f_u_dadda_cla32_fa238_and1;
  wire f_u_dadda_cla32_fa238_or0;
  wire f_u_dadda_cla32_and_6_21;
  wire f_u_dadda_cla32_and_5_22;
  wire f_u_dadda_cla32_and_4_23;
  wire f_u_dadda_cla32_fa239_xor0;
  wire f_u_dadda_cla32_fa239_and0;
  wire f_u_dadda_cla32_fa239_xor1;
  wire f_u_dadda_cla32_fa239_and1;
  wire f_u_dadda_cla32_fa239_or0;
  wire f_u_dadda_cla32_and_3_24;
  wire f_u_dadda_cla32_and_2_25;
  wire f_u_dadda_cla32_and_1_26;
  wire f_u_dadda_cla32_fa240_xor0;
  wire f_u_dadda_cla32_fa240_and0;
  wire f_u_dadda_cla32_fa240_xor1;
  wire f_u_dadda_cla32_fa240_and1;
  wire f_u_dadda_cla32_fa240_or0;
  wire f_u_dadda_cla32_and_0_27;
  wire f_u_dadda_cla32_fa241_xor0;
  wire f_u_dadda_cla32_fa241_and0;
  wire f_u_dadda_cla32_fa241_xor1;
  wire f_u_dadda_cla32_fa241_and1;
  wire f_u_dadda_cla32_fa241_or0;
  wire f_u_dadda_cla32_fa242_xor0;
  wire f_u_dadda_cla32_fa242_and0;
  wire f_u_dadda_cla32_fa242_xor1;
  wire f_u_dadda_cla32_fa242_and1;
  wire f_u_dadda_cla32_fa242_or0;
  wire f_u_dadda_cla32_fa243_xor0;
  wire f_u_dadda_cla32_fa243_and0;
  wire f_u_dadda_cla32_fa243_xor1;
  wire f_u_dadda_cla32_fa243_and1;
  wire f_u_dadda_cla32_fa243_or0;
  wire f_u_dadda_cla32_fa244_xor0;
  wire f_u_dadda_cla32_fa244_and0;
  wire f_u_dadda_cla32_fa244_xor1;
  wire f_u_dadda_cla32_fa244_and1;
  wire f_u_dadda_cla32_fa244_or0;
  wire f_u_dadda_cla32_fa245_xor0;
  wire f_u_dadda_cla32_fa245_and0;
  wire f_u_dadda_cla32_fa245_xor1;
  wire f_u_dadda_cla32_fa245_and1;
  wire f_u_dadda_cla32_fa245_or0;
  wire f_u_dadda_cla32_ha26_xor0;
  wire f_u_dadda_cla32_ha26_and0;
  wire f_u_dadda_cla32_fa246_xor0;
  wire f_u_dadda_cla32_fa246_and0;
  wire f_u_dadda_cla32_fa246_xor1;
  wire f_u_dadda_cla32_fa246_and1;
  wire f_u_dadda_cla32_fa246_or0;
  wire f_u_dadda_cla32_fa247_xor0;
  wire f_u_dadda_cla32_fa247_and0;
  wire f_u_dadda_cla32_fa247_xor1;
  wire f_u_dadda_cla32_fa247_and1;
  wire f_u_dadda_cla32_fa247_or0;
  wire f_u_dadda_cla32_fa248_xor0;
  wire f_u_dadda_cla32_fa248_and0;
  wire f_u_dadda_cla32_fa248_xor1;
  wire f_u_dadda_cla32_fa248_and1;
  wire f_u_dadda_cla32_fa248_or0;
  wire f_u_dadda_cla32_fa249_xor0;
  wire f_u_dadda_cla32_fa249_and0;
  wire f_u_dadda_cla32_fa249_xor1;
  wire f_u_dadda_cla32_fa249_and1;
  wire f_u_dadda_cla32_fa249_or0;
  wire f_u_dadda_cla32_fa250_xor0;
  wire f_u_dadda_cla32_fa250_and0;
  wire f_u_dadda_cla32_fa250_xor1;
  wire f_u_dadda_cla32_fa250_and1;
  wire f_u_dadda_cla32_fa250_or0;
  wire f_u_dadda_cla32_fa251_xor0;
  wire f_u_dadda_cla32_fa251_and0;
  wire f_u_dadda_cla32_fa251_xor1;
  wire f_u_dadda_cla32_fa251_and1;
  wire f_u_dadda_cla32_fa251_or0;
  wire f_u_dadda_cla32_fa252_xor0;
  wire f_u_dadda_cla32_fa252_and0;
  wire f_u_dadda_cla32_fa252_xor1;
  wire f_u_dadda_cla32_fa252_and1;
  wire f_u_dadda_cla32_fa252_or0;
  wire f_u_dadda_cla32_and_26_2;
  wire f_u_dadda_cla32_and_25_3;
  wire f_u_dadda_cla32_fa253_xor0;
  wire f_u_dadda_cla32_fa253_and0;
  wire f_u_dadda_cla32_fa253_xor1;
  wire f_u_dadda_cla32_fa253_and1;
  wire f_u_dadda_cla32_fa253_or0;
  wire f_u_dadda_cla32_and_24_4;
  wire f_u_dadda_cla32_and_23_5;
  wire f_u_dadda_cla32_and_22_6;
  wire f_u_dadda_cla32_fa254_xor0;
  wire f_u_dadda_cla32_fa254_and0;
  wire f_u_dadda_cla32_fa254_xor1;
  wire f_u_dadda_cla32_fa254_and1;
  wire f_u_dadda_cla32_fa254_or0;
  wire f_u_dadda_cla32_and_21_7;
  wire f_u_dadda_cla32_and_20_8;
  wire f_u_dadda_cla32_and_19_9;
  wire f_u_dadda_cla32_fa255_xor0;
  wire f_u_dadda_cla32_fa255_and0;
  wire f_u_dadda_cla32_fa255_xor1;
  wire f_u_dadda_cla32_fa255_and1;
  wire f_u_dadda_cla32_fa255_or0;
  wire f_u_dadda_cla32_and_18_10;
  wire f_u_dadda_cla32_and_17_11;
  wire f_u_dadda_cla32_and_16_12;
  wire f_u_dadda_cla32_fa256_xor0;
  wire f_u_dadda_cla32_fa256_and0;
  wire f_u_dadda_cla32_fa256_xor1;
  wire f_u_dadda_cla32_fa256_and1;
  wire f_u_dadda_cla32_fa256_or0;
  wire f_u_dadda_cla32_and_15_13;
  wire f_u_dadda_cla32_and_14_14;
  wire f_u_dadda_cla32_and_13_15;
  wire f_u_dadda_cla32_fa257_xor0;
  wire f_u_dadda_cla32_fa257_and0;
  wire f_u_dadda_cla32_fa257_xor1;
  wire f_u_dadda_cla32_fa257_and1;
  wire f_u_dadda_cla32_fa257_or0;
  wire f_u_dadda_cla32_and_12_16;
  wire f_u_dadda_cla32_and_11_17;
  wire f_u_dadda_cla32_and_10_18;
  wire f_u_dadda_cla32_fa258_xor0;
  wire f_u_dadda_cla32_fa258_and0;
  wire f_u_dadda_cla32_fa258_xor1;
  wire f_u_dadda_cla32_fa258_and1;
  wire f_u_dadda_cla32_fa258_or0;
  wire f_u_dadda_cla32_and_9_19;
  wire f_u_dadda_cla32_and_8_20;
  wire f_u_dadda_cla32_and_7_21;
  wire f_u_dadda_cla32_fa259_xor0;
  wire f_u_dadda_cla32_fa259_and0;
  wire f_u_dadda_cla32_fa259_xor1;
  wire f_u_dadda_cla32_fa259_and1;
  wire f_u_dadda_cla32_fa259_or0;
  wire f_u_dadda_cla32_and_6_22;
  wire f_u_dadda_cla32_and_5_23;
  wire f_u_dadda_cla32_and_4_24;
  wire f_u_dadda_cla32_fa260_xor0;
  wire f_u_dadda_cla32_fa260_and0;
  wire f_u_dadda_cla32_fa260_xor1;
  wire f_u_dadda_cla32_fa260_and1;
  wire f_u_dadda_cla32_fa260_or0;
  wire f_u_dadda_cla32_and_3_25;
  wire f_u_dadda_cla32_and_2_26;
  wire f_u_dadda_cla32_and_1_27;
  wire f_u_dadda_cla32_fa261_xor0;
  wire f_u_dadda_cla32_fa261_and0;
  wire f_u_dadda_cla32_fa261_xor1;
  wire f_u_dadda_cla32_fa261_and1;
  wire f_u_dadda_cla32_fa261_or0;
  wire f_u_dadda_cla32_and_0_28;
  wire f_u_dadda_cla32_fa262_xor0;
  wire f_u_dadda_cla32_fa262_and0;
  wire f_u_dadda_cla32_fa262_xor1;
  wire f_u_dadda_cla32_fa262_and1;
  wire f_u_dadda_cla32_fa262_or0;
  wire f_u_dadda_cla32_fa263_xor0;
  wire f_u_dadda_cla32_fa263_and0;
  wire f_u_dadda_cla32_fa263_xor1;
  wire f_u_dadda_cla32_fa263_and1;
  wire f_u_dadda_cla32_fa263_or0;
  wire f_u_dadda_cla32_fa264_xor0;
  wire f_u_dadda_cla32_fa264_and0;
  wire f_u_dadda_cla32_fa264_xor1;
  wire f_u_dadda_cla32_fa264_and1;
  wire f_u_dadda_cla32_fa264_or0;
  wire f_u_dadda_cla32_fa265_xor0;
  wire f_u_dadda_cla32_fa265_and0;
  wire f_u_dadda_cla32_fa265_xor1;
  wire f_u_dadda_cla32_fa265_and1;
  wire f_u_dadda_cla32_fa265_or0;
  wire f_u_dadda_cla32_fa266_xor0;
  wire f_u_dadda_cla32_fa266_and0;
  wire f_u_dadda_cla32_fa266_xor1;
  wire f_u_dadda_cla32_fa266_and1;
  wire f_u_dadda_cla32_fa266_or0;
  wire f_u_dadda_cla32_fa267_xor0;
  wire f_u_dadda_cla32_fa267_and0;
  wire f_u_dadda_cla32_fa267_xor1;
  wire f_u_dadda_cla32_fa267_and1;
  wire f_u_dadda_cla32_fa267_or0;
  wire f_u_dadda_cla32_fa268_xor0;
  wire f_u_dadda_cla32_fa268_and0;
  wire f_u_dadda_cla32_fa268_xor1;
  wire f_u_dadda_cla32_fa268_and1;
  wire f_u_dadda_cla32_fa268_or0;
  wire f_u_dadda_cla32_fa269_xor0;
  wire f_u_dadda_cla32_fa269_and0;
  wire f_u_dadda_cla32_fa269_xor1;
  wire f_u_dadda_cla32_fa269_and1;
  wire f_u_dadda_cla32_fa269_or0;
  wire f_u_dadda_cla32_fa270_xor0;
  wire f_u_dadda_cla32_fa270_and0;
  wire f_u_dadda_cla32_fa270_xor1;
  wire f_u_dadda_cla32_fa270_and1;
  wire f_u_dadda_cla32_fa270_or0;
  wire f_u_dadda_cla32_fa271_xor0;
  wire f_u_dadda_cla32_fa271_and0;
  wire f_u_dadda_cla32_fa271_xor1;
  wire f_u_dadda_cla32_fa271_and1;
  wire f_u_dadda_cla32_fa271_or0;
  wire f_u_dadda_cla32_fa272_xor0;
  wire f_u_dadda_cla32_fa272_and0;
  wire f_u_dadda_cla32_fa272_xor1;
  wire f_u_dadda_cla32_fa272_and1;
  wire f_u_dadda_cla32_fa272_or0;
  wire f_u_dadda_cla32_fa273_xor0;
  wire f_u_dadda_cla32_fa273_and0;
  wire f_u_dadda_cla32_fa273_xor1;
  wire f_u_dadda_cla32_fa273_and1;
  wire f_u_dadda_cla32_fa273_or0;
  wire f_u_dadda_cla32_fa274_xor0;
  wire f_u_dadda_cla32_fa274_and0;
  wire f_u_dadda_cla32_fa274_xor1;
  wire f_u_dadda_cla32_fa274_and1;
  wire f_u_dadda_cla32_fa274_or0;
  wire f_u_dadda_cla32_and_25_4;
  wire f_u_dadda_cla32_and_24_5;
  wire f_u_dadda_cla32_fa275_xor0;
  wire f_u_dadda_cla32_fa275_and0;
  wire f_u_dadda_cla32_fa275_xor1;
  wire f_u_dadda_cla32_fa275_and1;
  wire f_u_dadda_cla32_fa275_or0;
  wire f_u_dadda_cla32_and_23_6;
  wire f_u_dadda_cla32_and_22_7;
  wire f_u_dadda_cla32_and_21_8;
  wire f_u_dadda_cla32_fa276_xor0;
  wire f_u_dadda_cla32_fa276_and0;
  wire f_u_dadda_cla32_fa276_xor1;
  wire f_u_dadda_cla32_fa276_and1;
  wire f_u_dadda_cla32_fa276_or0;
  wire f_u_dadda_cla32_and_20_9;
  wire f_u_dadda_cla32_and_19_10;
  wire f_u_dadda_cla32_and_18_11;
  wire f_u_dadda_cla32_fa277_xor0;
  wire f_u_dadda_cla32_fa277_and0;
  wire f_u_dadda_cla32_fa277_xor1;
  wire f_u_dadda_cla32_fa277_and1;
  wire f_u_dadda_cla32_fa277_or0;
  wire f_u_dadda_cla32_and_17_12;
  wire f_u_dadda_cla32_and_16_13;
  wire f_u_dadda_cla32_and_15_14;
  wire f_u_dadda_cla32_fa278_xor0;
  wire f_u_dadda_cla32_fa278_and0;
  wire f_u_dadda_cla32_fa278_xor1;
  wire f_u_dadda_cla32_fa278_and1;
  wire f_u_dadda_cla32_fa278_or0;
  wire f_u_dadda_cla32_and_14_15;
  wire f_u_dadda_cla32_and_13_16;
  wire f_u_dadda_cla32_and_12_17;
  wire f_u_dadda_cla32_fa279_xor0;
  wire f_u_dadda_cla32_fa279_and0;
  wire f_u_dadda_cla32_fa279_xor1;
  wire f_u_dadda_cla32_fa279_and1;
  wire f_u_dadda_cla32_fa279_or0;
  wire f_u_dadda_cla32_and_11_18;
  wire f_u_dadda_cla32_and_10_19;
  wire f_u_dadda_cla32_and_9_20;
  wire f_u_dadda_cla32_fa280_xor0;
  wire f_u_dadda_cla32_fa280_and0;
  wire f_u_dadda_cla32_fa280_xor1;
  wire f_u_dadda_cla32_fa280_and1;
  wire f_u_dadda_cla32_fa280_or0;
  wire f_u_dadda_cla32_and_8_21;
  wire f_u_dadda_cla32_and_7_22;
  wire f_u_dadda_cla32_and_6_23;
  wire f_u_dadda_cla32_fa281_xor0;
  wire f_u_dadda_cla32_fa281_and0;
  wire f_u_dadda_cla32_fa281_xor1;
  wire f_u_dadda_cla32_fa281_and1;
  wire f_u_dadda_cla32_fa281_or0;
  wire f_u_dadda_cla32_and_5_24;
  wire f_u_dadda_cla32_and_4_25;
  wire f_u_dadda_cla32_and_3_26;
  wire f_u_dadda_cla32_fa282_xor0;
  wire f_u_dadda_cla32_fa282_and0;
  wire f_u_dadda_cla32_fa282_xor1;
  wire f_u_dadda_cla32_fa282_and1;
  wire f_u_dadda_cla32_fa282_or0;
  wire f_u_dadda_cla32_and_2_27;
  wire f_u_dadda_cla32_and_1_28;
  wire f_u_dadda_cla32_and_0_29;
  wire f_u_dadda_cla32_fa283_xor0;
  wire f_u_dadda_cla32_fa283_and0;
  wire f_u_dadda_cla32_fa283_xor1;
  wire f_u_dadda_cla32_fa283_and1;
  wire f_u_dadda_cla32_fa283_or0;
  wire f_u_dadda_cla32_fa284_xor0;
  wire f_u_dadda_cla32_fa284_and0;
  wire f_u_dadda_cla32_fa284_xor1;
  wire f_u_dadda_cla32_fa284_and1;
  wire f_u_dadda_cla32_fa284_or0;
  wire f_u_dadda_cla32_fa285_xor0;
  wire f_u_dadda_cla32_fa285_and0;
  wire f_u_dadda_cla32_fa285_xor1;
  wire f_u_dadda_cla32_fa285_and1;
  wire f_u_dadda_cla32_fa285_or0;
  wire f_u_dadda_cla32_fa286_xor0;
  wire f_u_dadda_cla32_fa286_and0;
  wire f_u_dadda_cla32_fa286_xor1;
  wire f_u_dadda_cla32_fa286_and1;
  wire f_u_dadda_cla32_fa286_or0;
  wire f_u_dadda_cla32_fa287_xor0;
  wire f_u_dadda_cla32_fa287_and0;
  wire f_u_dadda_cla32_fa287_xor1;
  wire f_u_dadda_cla32_fa287_and1;
  wire f_u_dadda_cla32_fa287_or0;
  wire f_u_dadda_cla32_fa288_xor0;
  wire f_u_dadda_cla32_fa288_and0;
  wire f_u_dadda_cla32_fa288_xor1;
  wire f_u_dadda_cla32_fa288_and1;
  wire f_u_dadda_cla32_fa288_or0;
  wire f_u_dadda_cla32_fa289_xor0;
  wire f_u_dadda_cla32_fa289_and0;
  wire f_u_dadda_cla32_fa289_xor1;
  wire f_u_dadda_cla32_fa289_and1;
  wire f_u_dadda_cla32_fa289_or0;
  wire f_u_dadda_cla32_fa290_xor0;
  wire f_u_dadda_cla32_fa290_and0;
  wire f_u_dadda_cla32_fa290_xor1;
  wire f_u_dadda_cla32_fa290_and1;
  wire f_u_dadda_cla32_fa290_or0;
  wire f_u_dadda_cla32_fa291_xor0;
  wire f_u_dadda_cla32_fa291_and0;
  wire f_u_dadda_cla32_fa291_xor1;
  wire f_u_dadda_cla32_fa291_and1;
  wire f_u_dadda_cla32_fa291_or0;
  wire f_u_dadda_cla32_fa292_xor0;
  wire f_u_dadda_cla32_fa292_and0;
  wire f_u_dadda_cla32_fa292_xor1;
  wire f_u_dadda_cla32_fa292_and1;
  wire f_u_dadda_cla32_fa292_or0;
  wire f_u_dadda_cla32_fa293_xor0;
  wire f_u_dadda_cla32_fa293_and0;
  wire f_u_dadda_cla32_fa293_xor1;
  wire f_u_dadda_cla32_fa293_and1;
  wire f_u_dadda_cla32_fa293_or0;
  wire f_u_dadda_cla32_fa294_xor0;
  wire f_u_dadda_cla32_fa294_and0;
  wire f_u_dadda_cla32_fa294_xor1;
  wire f_u_dadda_cla32_fa294_and1;
  wire f_u_dadda_cla32_fa294_or0;
  wire f_u_dadda_cla32_fa295_xor0;
  wire f_u_dadda_cla32_fa295_and0;
  wire f_u_dadda_cla32_fa295_xor1;
  wire f_u_dadda_cla32_fa295_and1;
  wire f_u_dadda_cla32_fa295_or0;
  wire f_u_dadda_cla32_fa296_xor0;
  wire f_u_dadda_cla32_fa296_and0;
  wire f_u_dadda_cla32_fa296_xor1;
  wire f_u_dadda_cla32_fa296_and1;
  wire f_u_dadda_cla32_fa296_or0;
  wire f_u_dadda_cla32_and_24_6;
  wire f_u_dadda_cla32_and_23_7;
  wire f_u_dadda_cla32_fa297_xor0;
  wire f_u_dadda_cla32_fa297_and0;
  wire f_u_dadda_cla32_fa297_xor1;
  wire f_u_dadda_cla32_fa297_and1;
  wire f_u_dadda_cla32_fa297_or0;
  wire f_u_dadda_cla32_and_22_8;
  wire f_u_dadda_cla32_and_21_9;
  wire f_u_dadda_cla32_and_20_10;
  wire f_u_dadda_cla32_fa298_xor0;
  wire f_u_dadda_cla32_fa298_and0;
  wire f_u_dadda_cla32_fa298_xor1;
  wire f_u_dadda_cla32_fa298_and1;
  wire f_u_dadda_cla32_fa298_or0;
  wire f_u_dadda_cla32_and_19_11;
  wire f_u_dadda_cla32_and_18_12;
  wire f_u_dadda_cla32_and_17_13;
  wire f_u_dadda_cla32_fa299_xor0;
  wire f_u_dadda_cla32_fa299_and0;
  wire f_u_dadda_cla32_fa299_xor1;
  wire f_u_dadda_cla32_fa299_and1;
  wire f_u_dadda_cla32_fa299_or0;
  wire f_u_dadda_cla32_and_16_14;
  wire f_u_dadda_cla32_and_15_15;
  wire f_u_dadda_cla32_and_14_16;
  wire f_u_dadda_cla32_fa300_xor0;
  wire f_u_dadda_cla32_fa300_and0;
  wire f_u_dadda_cla32_fa300_xor1;
  wire f_u_dadda_cla32_fa300_and1;
  wire f_u_dadda_cla32_fa300_or0;
  wire f_u_dadda_cla32_and_13_17;
  wire f_u_dadda_cla32_and_12_18;
  wire f_u_dadda_cla32_and_11_19;
  wire f_u_dadda_cla32_fa301_xor0;
  wire f_u_dadda_cla32_fa301_and0;
  wire f_u_dadda_cla32_fa301_xor1;
  wire f_u_dadda_cla32_fa301_and1;
  wire f_u_dadda_cla32_fa301_or0;
  wire f_u_dadda_cla32_and_10_20;
  wire f_u_dadda_cla32_and_9_21;
  wire f_u_dadda_cla32_and_8_22;
  wire f_u_dadda_cla32_fa302_xor0;
  wire f_u_dadda_cla32_fa302_and0;
  wire f_u_dadda_cla32_fa302_xor1;
  wire f_u_dadda_cla32_fa302_and1;
  wire f_u_dadda_cla32_fa302_or0;
  wire f_u_dadda_cla32_and_7_23;
  wire f_u_dadda_cla32_and_6_24;
  wire f_u_dadda_cla32_and_5_25;
  wire f_u_dadda_cla32_fa303_xor0;
  wire f_u_dadda_cla32_fa303_and0;
  wire f_u_dadda_cla32_fa303_xor1;
  wire f_u_dadda_cla32_fa303_and1;
  wire f_u_dadda_cla32_fa303_or0;
  wire f_u_dadda_cla32_and_4_26;
  wire f_u_dadda_cla32_and_3_27;
  wire f_u_dadda_cla32_and_2_28;
  wire f_u_dadda_cla32_fa304_xor0;
  wire f_u_dadda_cla32_fa304_and0;
  wire f_u_dadda_cla32_fa304_xor1;
  wire f_u_dadda_cla32_fa304_and1;
  wire f_u_dadda_cla32_fa304_or0;
  wire f_u_dadda_cla32_and_1_29;
  wire f_u_dadda_cla32_and_0_30;
  wire f_u_dadda_cla32_fa305_xor0;
  wire f_u_dadda_cla32_fa305_and0;
  wire f_u_dadda_cla32_fa305_xor1;
  wire f_u_dadda_cla32_fa305_and1;
  wire f_u_dadda_cla32_fa305_or0;
  wire f_u_dadda_cla32_fa306_xor0;
  wire f_u_dadda_cla32_fa306_and0;
  wire f_u_dadda_cla32_fa306_xor1;
  wire f_u_dadda_cla32_fa306_and1;
  wire f_u_dadda_cla32_fa306_or0;
  wire f_u_dadda_cla32_fa307_xor0;
  wire f_u_dadda_cla32_fa307_and0;
  wire f_u_dadda_cla32_fa307_xor1;
  wire f_u_dadda_cla32_fa307_and1;
  wire f_u_dadda_cla32_fa307_or0;
  wire f_u_dadda_cla32_fa308_xor0;
  wire f_u_dadda_cla32_fa308_and0;
  wire f_u_dadda_cla32_fa308_xor1;
  wire f_u_dadda_cla32_fa308_and1;
  wire f_u_dadda_cla32_fa308_or0;
  wire f_u_dadda_cla32_fa309_xor0;
  wire f_u_dadda_cla32_fa309_and0;
  wire f_u_dadda_cla32_fa309_xor1;
  wire f_u_dadda_cla32_fa309_and1;
  wire f_u_dadda_cla32_fa309_or0;
  wire f_u_dadda_cla32_fa310_xor0;
  wire f_u_dadda_cla32_fa310_and0;
  wire f_u_dadda_cla32_fa310_xor1;
  wire f_u_dadda_cla32_fa310_and1;
  wire f_u_dadda_cla32_fa310_or0;
  wire f_u_dadda_cla32_fa311_xor0;
  wire f_u_dadda_cla32_fa311_and0;
  wire f_u_dadda_cla32_fa311_xor1;
  wire f_u_dadda_cla32_fa311_and1;
  wire f_u_dadda_cla32_fa311_or0;
  wire f_u_dadda_cla32_fa312_xor0;
  wire f_u_dadda_cla32_fa312_and0;
  wire f_u_dadda_cla32_fa312_xor1;
  wire f_u_dadda_cla32_fa312_and1;
  wire f_u_dadda_cla32_fa312_or0;
  wire f_u_dadda_cla32_fa313_xor0;
  wire f_u_dadda_cla32_fa313_and0;
  wire f_u_dadda_cla32_fa313_xor1;
  wire f_u_dadda_cla32_fa313_and1;
  wire f_u_dadda_cla32_fa313_or0;
  wire f_u_dadda_cla32_fa314_xor0;
  wire f_u_dadda_cla32_fa314_and0;
  wire f_u_dadda_cla32_fa314_xor1;
  wire f_u_dadda_cla32_fa314_and1;
  wire f_u_dadda_cla32_fa314_or0;
  wire f_u_dadda_cla32_fa315_xor0;
  wire f_u_dadda_cla32_fa315_and0;
  wire f_u_dadda_cla32_fa315_xor1;
  wire f_u_dadda_cla32_fa315_and1;
  wire f_u_dadda_cla32_fa315_or0;
  wire f_u_dadda_cla32_fa316_xor0;
  wire f_u_dadda_cla32_fa316_and0;
  wire f_u_dadda_cla32_fa316_xor1;
  wire f_u_dadda_cla32_fa316_and1;
  wire f_u_dadda_cla32_fa316_or0;
  wire f_u_dadda_cla32_fa317_xor0;
  wire f_u_dadda_cla32_fa317_and0;
  wire f_u_dadda_cla32_fa317_xor1;
  wire f_u_dadda_cla32_fa317_and1;
  wire f_u_dadda_cla32_fa317_or0;
  wire f_u_dadda_cla32_fa318_xor0;
  wire f_u_dadda_cla32_fa318_and0;
  wire f_u_dadda_cla32_fa318_xor1;
  wire f_u_dadda_cla32_fa318_and1;
  wire f_u_dadda_cla32_fa318_or0;
  wire f_u_dadda_cla32_and_23_8;
  wire f_u_dadda_cla32_and_22_9;
  wire f_u_dadda_cla32_fa319_xor0;
  wire f_u_dadda_cla32_fa319_and0;
  wire f_u_dadda_cla32_fa319_xor1;
  wire f_u_dadda_cla32_fa319_and1;
  wire f_u_dadda_cla32_fa319_or0;
  wire f_u_dadda_cla32_and_21_10;
  wire f_u_dadda_cla32_and_20_11;
  wire f_u_dadda_cla32_and_19_12;
  wire f_u_dadda_cla32_fa320_xor0;
  wire f_u_dadda_cla32_fa320_and0;
  wire f_u_dadda_cla32_fa320_xor1;
  wire f_u_dadda_cla32_fa320_and1;
  wire f_u_dadda_cla32_fa320_or0;
  wire f_u_dadda_cla32_and_18_13;
  wire f_u_dadda_cla32_and_17_14;
  wire f_u_dadda_cla32_and_16_15;
  wire f_u_dadda_cla32_fa321_xor0;
  wire f_u_dadda_cla32_fa321_and0;
  wire f_u_dadda_cla32_fa321_xor1;
  wire f_u_dadda_cla32_fa321_and1;
  wire f_u_dadda_cla32_fa321_or0;
  wire f_u_dadda_cla32_and_15_16;
  wire f_u_dadda_cla32_and_14_17;
  wire f_u_dadda_cla32_and_13_18;
  wire f_u_dadda_cla32_fa322_xor0;
  wire f_u_dadda_cla32_fa322_and0;
  wire f_u_dadda_cla32_fa322_xor1;
  wire f_u_dadda_cla32_fa322_and1;
  wire f_u_dadda_cla32_fa322_or0;
  wire f_u_dadda_cla32_and_12_19;
  wire f_u_dadda_cla32_and_11_20;
  wire f_u_dadda_cla32_and_10_21;
  wire f_u_dadda_cla32_fa323_xor0;
  wire f_u_dadda_cla32_fa323_and0;
  wire f_u_dadda_cla32_fa323_xor1;
  wire f_u_dadda_cla32_fa323_and1;
  wire f_u_dadda_cla32_fa323_or0;
  wire f_u_dadda_cla32_and_9_22;
  wire f_u_dadda_cla32_and_8_23;
  wire f_u_dadda_cla32_and_7_24;
  wire f_u_dadda_cla32_fa324_xor0;
  wire f_u_dadda_cla32_fa324_and0;
  wire f_u_dadda_cla32_fa324_xor1;
  wire f_u_dadda_cla32_fa324_and1;
  wire f_u_dadda_cla32_fa324_or0;
  wire f_u_dadda_cla32_and_6_25;
  wire f_u_dadda_cla32_and_5_26;
  wire f_u_dadda_cla32_and_4_27;
  wire f_u_dadda_cla32_fa325_xor0;
  wire f_u_dadda_cla32_fa325_and0;
  wire f_u_dadda_cla32_fa325_xor1;
  wire f_u_dadda_cla32_fa325_and1;
  wire f_u_dadda_cla32_fa325_or0;
  wire f_u_dadda_cla32_and_3_28;
  wire f_u_dadda_cla32_and_2_29;
  wire f_u_dadda_cla32_and_1_30;
  wire f_u_dadda_cla32_fa326_xor0;
  wire f_u_dadda_cla32_fa326_and0;
  wire f_u_dadda_cla32_fa326_xor1;
  wire f_u_dadda_cla32_fa326_and1;
  wire f_u_dadda_cla32_fa326_or0;
  wire f_u_dadda_cla32_and_0_31;
  wire f_u_dadda_cla32_fa327_xor0;
  wire f_u_dadda_cla32_fa327_and0;
  wire f_u_dadda_cla32_fa327_xor1;
  wire f_u_dadda_cla32_fa327_and1;
  wire f_u_dadda_cla32_fa327_or0;
  wire f_u_dadda_cla32_fa328_xor0;
  wire f_u_dadda_cla32_fa328_and0;
  wire f_u_dadda_cla32_fa328_xor1;
  wire f_u_dadda_cla32_fa328_and1;
  wire f_u_dadda_cla32_fa328_or0;
  wire f_u_dadda_cla32_fa329_xor0;
  wire f_u_dadda_cla32_fa329_and0;
  wire f_u_dadda_cla32_fa329_xor1;
  wire f_u_dadda_cla32_fa329_and1;
  wire f_u_dadda_cla32_fa329_or0;
  wire f_u_dadda_cla32_fa330_xor0;
  wire f_u_dadda_cla32_fa330_and0;
  wire f_u_dadda_cla32_fa330_xor1;
  wire f_u_dadda_cla32_fa330_and1;
  wire f_u_dadda_cla32_fa330_or0;
  wire f_u_dadda_cla32_fa331_xor0;
  wire f_u_dadda_cla32_fa331_and0;
  wire f_u_dadda_cla32_fa331_xor1;
  wire f_u_dadda_cla32_fa331_and1;
  wire f_u_dadda_cla32_fa331_or0;
  wire f_u_dadda_cla32_fa332_xor0;
  wire f_u_dadda_cla32_fa332_and0;
  wire f_u_dadda_cla32_fa332_xor1;
  wire f_u_dadda_cla32_fa332_and1;
  wire f_u_dadda_cla32_fa332_or0;
  wire f_u_dadda_cla32_fa333_xor0;
  wire f_u_dadda_cla32_fa333_and0;
  wire f_u_dadda_cla32_fa333_xor1;
  wire f_u_dadda_cla32_fa333_and1;
  wire f_u_dadda_cla32_fa333_or0;
  wire f_u_dadda_cla32_fa334_xor0;
  wire f_u_dadda_cla32_fa334_and0;
  wire f_u_dadda_cla32_fa334_xor1;
  wire f_u_dadda_cla32_fa334_and1;
  wire f_u_dadda_cla32_fa334_or0;
  wire f_u_dadda_cla32_fa335_xor0;
  wire f_u_dadda_cla32_fa335_and0;
  wire f_u_dadda_cla32_fa335_xor1;
  wire f_u_dadda_cla32_fa335_and1;
  wire f_u_dadda_cla32_fa335_or0;
  wire f_u_dadda_cla32_fa336_xor0;
  wire f_u_dadda_cla32_fa336_and0;
  wire f_u_dadda_cla32_fa336_xor1;
  wire f_u_dadda_cla32_fa336_and1;
  wire f_u_dadda_cla32_fa336_or0;
  wire f_u_dadda_cla32_fa337_xor0;
  wire f_u_dadda_cla32_fa337_and0;
  wire f_u_dadda_cla32_fa337_xor1;
  wire f_u_dadda_cla32_fa337_and1;
  wire f_u_dadda_cla32_fa337_or0;
  wire f_u_dadda_cla32_fa338_xor0;
  wire f_u_dadda_cla32_fa338_and0;
  wire f_u_dadda_cla32_fa338_xor1;
  wire f_u_dadda_cla32_fa338_and1;
  wire f_u_dadda_cla32_fa338_or0;
  wire f_u_dadda_cla32_fa339_xor0;
  wire f_u_dadda_cla32_fa339_and0;
  wire f_u_dadda_cla32_fa339_xor1;
  wire f_u_dadda_cla32_fa339_and1;
  wire f_u_dadda_cla32_fa339_or0;
  wire f_u_dadda_cla32_fa340_xor0;
  wire f_u_dadda_cla32_fa340_and0;
  wire f_u_dadda_cla32_fa340_xor1;
  wire f_u_dadda_cla32_fa340_and1;
  wire f_u_dadda_cla32_fa340_or0;
  wire f_u_dadda_cla32_and_24_8;
  wire f_u_dadda_cla32_and_23_9;
  wire f_u_dadda_cla32_fa341_xor0;
  wire f_u_dadda_cla32_fa341_and0;
  wire f_u_dadda_cla32_fa341_xor1;
  wire f_u_dadda_cla32_fa341_and1;
  wire f_u_dadda_cla32_fa341_or0;
  wire f_u_dadda_cla32_and_22_10;
  wire f_u_dadda_cla32_and_21_11;
  wire f_u_dadda_cla32_and_20_12;
  wire f_u_dadda_cla32_fa342_xor0;
  wire f_u_dadda_cla32_fa342_and0;
  wire f_u_dadda_cla32_fa342_xor1;
  wire f_u_dadda_cla32_fa342_and1;
  wire f_u_dadda_cla32_fa342_or0;
  wire f_u_dadda_cla32_and_19_13;
  wire f_u_dadda_cla32_and_18_14;
  wire f_u_dadda_cla32_and_17_15;
  wire f_u_dadda_cla32_fa343_xor0;
  wire f_u_dadda_cla32_fa343_and0;
  wire f_u_dadda_cla32_fa343_xor1;
  wire f_u_dadda_cla32_fa343_and1;
  wire f_u_dadda_cla32_fa343_or0;
  wire f_u_dadda_cla32_and_16_16;
  wire f_u_dadda_cla32_and_15_17;
  wire f_u_dadda_cla32_and_14_18;
  wire f_u_dadda_cla32_fa344_xor0;
  wire f_u_dadda_cla32_fa344_and0;
  wire f_u_dadda_cla32_fa344_xor1;
  wire f_u_dadda_cla32_fa344_and1;
  wire f_u_dadda_cla32_fa344_or0;
  wire f_u_dadda_cla32_and_13_19;
  wire f_u_dadda_cla32_and_12_20;
  wire f_u_dadda_cla32_and_11_21;
  wire f_u_dadda_cla32_fa345_xor0;
  wire f_u_dadda_cla32_fa345_and0;
  wire f_u_dadda_cla32_fa345_xor1;
  wire f_u_dadda_cla32_fa345_and1;
  wire f_u_dadda_cla32_fa345_or0;
  wire f_u_dadda_cla32_and_10_22;
  wire f_u_dadda_cla32_and_9_23;
  wire f_u_dadda_cla32_and_8_24;
  wire f_u_dadda_cla32_fa346_xor0;
  wire f_u_dadda_cla32_fa346_and0;
  wire f_u_dadda_cla32_fa346_xor1;
  wire f_u_dadda_cla32_fa346_and1;
  wire f_u_dadda_cla32_fa346_or0;
  wire f_u_dadda_cla32_and_7_25;
  wire f_u_dadda_cla32_and_6_26;
  wire f_u_dadda_cla32_and_5_27;
  wire f_u_dadda_cla32_fa347_xor0;
  wire f_u_dadda_cla32_fa347_and0;
  wire f_u_dadda_cla32_fa347_xor1;
  wire f_u_dadda_cla32_fa347_and1;
  wire f_u_dadda_cla32_fa347_or0;
  wire f_u_dadda_cla32_and_4_28;
  wire f_u_dadda_cla32_and_3_29;
  wire f_u_dadda_cla32_and_2_30;
  wire f_u_dadda_cla32_fa348_xor0;
  wire f_u_dadda_cla32_fa348_and0;
  wire f_u_dadda_cla32_fa348_xor1;
  wire f_u_dadda_cla32_fa348_and1;
  wire f_u_dadda_cla32_fa348_or0;
  wire f_u_dadda_cla32_and_1_31;
  wire f_u_dadda_cla32_fa349_xor0;
  wire f_u_dadda_cla32_fa349_and0;
  wire f_u_dadda_cla32_fa349_xor1;
  wire f_u_dadda_cla32_fa349_and1;
  wire f_u_dadda_cla32_fa349_or0;
  wire f_u_dadda_cla32_fa350_xor0;
  wire f_u_dadda_cla32_fa350_and0;
  wire f_u_dadda_cla32_fa350_xor1;
  wire f_u_dadda_cla32_fa350_and1;
  wire f_u_dadda_cla32_fa350_or0;
  wire f_u_dadda_cla32_fa351_xor0;
  wire f_u_dadda_cla32_fa351_and0;
  wire f_u_dadda_cla32_fa351_xor1;
  wire f_u_dadda_cla32_fa351_and1;
  wire f_u_dadda_cla32_fa351_or0;
  wire f_u_dadda_cla32_fa352_xor0;
  wire f_u_dadda_cla32_fa352_and0;
  wire f_u_dadda_cla32_fa352_xor1;
  wire f_u_dadda_cla32_fa352_and1;
  wire f_u_dadda_cla32_fa352_or0;
  wire f_u_dadda_cla32_fa353_xor0;
  wire f_u_dadda_cla32_fa353_and0;
  wire f_u_dadda_cla32_fa353_xor1;
  wire f_u_dadda_cla32_fa353_and1;
  wire f_u_dadda_cla32_fa353_or0;
  wire f_u_dadda_cla32_fa354_xor0;
  wire f_u_dadda_cla32_fa354_and0;
  wire f_u_dadda_cla32_fa354_xor1;
  wire f_u_dadda_cla32_fa354_and1;
  wire f_u_dadda_cla32_fa354_or0;
  wire f_u_dadda_cla32_fa355_xor0;
  wire f_u_dadda_cla32_fa355_and0;
  wire f_u_dadda_cla32_fa355_xor1;
  wire f_u_dadda_cla32_fa355_and1;
  wire f_u_dadda_cla32_fa355_or0;
  wire f_u_dadda_cla32_fa356_xor0;
  wire f_u_dadda_cla32_fa356_and0;
  wire f_u_dadda_cla32_fa356_xor1;
  wire f_u_dadda_cla32_fa356_and1;
  wire f_u_dadda_cla32_fa356_or0;
  wire f_u_dadda_cla32_fa357_xor0;
  wire f_u_dadda_cla32_fa357_and0;
  wire f_u_dadda_cla32_fa357_xor1;
  wire f_u_dadda_cla32_fa357_and1;
  wire f_u_dadda_cla32_fa357_or0;
  wire f_u_dadda_cla32_fa358_xor0;
  wire f_u_dadda_cla32_fa358_and0;
  wire f_u_dadda_cla32_fa358_xor1;
  wire f_u_dadda_cla32_fa358_and1;
  wire f_u_dadda_cla32_fa358_or0;
  wire f_u_dadda_cla32_fa359_xor0;
  wire f_u_dadda_cla32_fa359_and0;
  wire f_u_dadda_cla32_fa359_xor1;
  wire f_u_dadda_cla32_fa359_and1;
  wire f_u_dadda_cla32_fa359_or0;
  wire f_u_dadda_cla32_fa360_xor0;
  wire f_u_dadda_cla32_fa360_and0;
  wire f_u_dadda_cla32_fa360_xor1;
  wire f_u_dadda_cla32_fa360_and1;
  wire f_u_dadda_cla32_fa360_or0;
  wire f_u_dadda_cla32_fa361_xor0;
  wire f_u_dadda_cla32_fa361_and0;
  wire f_u_dadda_cla32_fa361_xor1;
  wire f_u_dadda_cla32_fa361_and1;
  wire f_u_dadda_cla32_fa361_or0;
  wire f_u_dadda_cla32_fa362_xor0;
  wire f_u_dadda_cla32_fa362_and0;
  wire f_u_dadda_cla32_fa362_xor1;
  wire f_u_dadda_cla32_fa362_and1;
  wire f_u_dadda_cla32_fa362_or0;
  wire f_u_dadda_cla32_and_26_7;
  wire f_u_dadda_cla32_and_25_8;
  wire f_u_dadda_cla32_fa363_xor0;
  wire f_u_dadda_cla32_fa363_and0;
  wire f_u_dadda_cla32_fa363_xor1;
  wire f_u_dadda_cla32_fa363_and1;
  wire f_u_dadda_cla32_fa363_or0;
  wire f_u_dadda_cla32_and_24_9;
  wire f_u_dadda_cla32_and_23_10;
  wire f_u_dadda_cla32_and_22_11;
  wire f_u_dadda_cla32_fa364_xor0;
  wire f_u_dadda_cla32_fa364_and0;
  wire f_u_dadda_cla32_fa364_xor1;
  wire f_u_dadda_cla32_fa364_and1;
  wire f_u_dadda_cla32_fa364_or0;
  wire f_u_dadda_cla32_and_21_12;
  wire f_u_dadda_cla32_and_20_13;
  wire f_u_dadda_cla32_and_19_14;
  wire f_u_dadda_cla32_fa365_xor0;
  wire f_u_dadda_cla32_fa365_and0;
  wire f_u_dadda_cla32_fa365_xor1;
  wire f_u_dadda_cla32_fa365_and1;
  wire f_u_dadda_cla32_fa365_or0;
  wire f_u_dadda_cla32_and_18_15;
  wire f_u_dadda_cla32_and_17_16;
  wire f_u_dadda_cla32_and_16_17;
  wire f_u_dadda_cla32_fa366_xor0;
  wire f_u_dadda_cla32_fa366_and0;
  wire f_u_dadda_cla32_fa366_xor1;
  wire f_u_dadda_cla32_fa366_and1;
  wire f_u_dadda_cla32_fa366_or0;
  wire f_u_dadda_cla32_and_15_18;
  wire f_u_dadda_cla32_and_14_19;
  wire f_u_dadda_cla32_and_13_20;
  wire f_u_dadda_cla32_fa367_xor0;
  wire f_u_dadda_cla32_fa367_and0;
  wire f_u_dadda_cla32_fa367_xor1;
  wire f_u_dadda_cla32_fa367_and1;
  wire f_u_dadda_cla32_fa367_or0;
  wire f_u_dadda_cla32_and_12_21;
  wire f_u_dadda_cla32_and_11_22;
  wire f_u_dadda_cla32_and_10_23;
  wire f_u_dadda_cla32_fa368_xor0;
  wire f_u_dadda_cla32_fa368_and0;
  wire f_u_dadda_cla32_fa368_xor1;
  wire f_u_dadda_cla32_fa368_and1;
  wire f_u_dadda_cla32_fa368_or0;
  wire f_u_dadda_cla32_and_9_24;
  wire f_u_dadda_cla32_and_8_25;
  wire f_u_dadda_cla32_and_7_26;
  wire f_u_dadda_cla32_fa369_xor0;
  wire f_u_dadda_cla32_fa369_and0;
  wire f_u_dadda_cla32_fa369_xor1;
  wire f_u_dadda_cla32_fa369_and1;
  wire f_u_dadda_cla32_fa369_or0;
  wire f_u_dadda_cla32_and_6_27;
  wire f_u_dadda_cla32_and_5_28;
  wire f_u_dadda_cla32_and_4_29;
  wire f_u_dadda_cla32_fa370_xor0;
  wire f_u_dadda_cla32_fa370_and0;
  wire f_u_dadda_cla32_fa370_xor1;
  wire f_u_dadda_cla32_fa370_and1;
  wire f_u_dadda_cla32_fa370_or0;
  wire f_u_dadda_cla32_and_3_30;
  wire f_u_dadda_cla32_and_2_31;
  wire f_u_dadda_cla32_fa371_xor0;
  wire f_u_dadda_cla32_fa371_and0;
  wire f_u_dadda_cla32_fa371_xor1;
  wire f_u_dadda_cla32_fa371_and1;
  wire f_u_dadda_cla32_fa371_or0;
  wire f_u_dadda_cla32_fa372_xor0;
  wire f_u_dadda_cla32_fa372_and0;
  wire f_u_dadda_cla32_fa372_xor1;
  wire f_u_dadda_cla32_fa372_and1;
  wire f_u_dadda_cla32_fa372_or0;
  wire f_u_dadda_cla32_fa373_xor0;
  wire f_u_dadda_cla32_fa373_and0;
  wire f_u_dadda_cla32_fa373_xor1;
  wire f_u_dadda_cla32_fa373_and1;
  wire f_u_dadda_cla32_fa373_or0;
  wire f_u_dadda_cla32_fa374_xor0;
  wire f_u_dadda_cla32_fa374_and0;
  wire f_u_dadda_cla32_fa374_xor1;
  wire f_u_dadda_cla32_fa374_and1;
  wire f_u_dadda_cla32_fa374_or0;
  wire f_u_dadda_cla32_fa375_xor0;
  wire f_u_dadda_cla32_fa375_and0;
  wire f_u_dadda_cla32_fa375_xor1;
  wire f_u_dadda_cla32_fa375_and1;
  wire f_u_dadda_cla32_fa375_or0;
  wire f_u_dadda_cla32_fa376_xor0;
  wire f_u_dadda_cla32_fa376_and0;
  wire f_u_dadda_cla32_fa376_xor1;
  wire f_u_dadda_cla32_fa376_and1;
  wire f_u_dadda_cla32_fa376_or0;
  wire f_u_dadda_cla32_fa377_xor0;
  wire f_u_dadda_cla32_fa377_and0;
  wire f_u_dadda_cla32_fa377_xor1;
  wire f_u_dadda_cla32_fa377_and1;
  wire f_u_dadda_cla32_fa377_or0;
  wire f_u_dadda_cla32_fa378_xor0;
  wire f_u_dadda_cla32_fa378_and0;
  wire f_u_dadda_cla32_fa378_xor1;
  wire f_u_dadda_cla32_fa378_and1;
  wire f_u_dadda_cla32_fa378_or0;
  wire f_u_dadda_cla32_fa379_xor0;
  wire f_u_dadda_cla32_fa379_and0;
  wire f_u_dadda_cla32_fa379_xor1;
  wire f_u_dadda_cla32_fa379_and1;
  wire f_u_dadda_cla32_fa379_or0;
  wire f_u_dadda_cla32_fa380_xor0;
  wire f_u_dadda_cla32_fa380_and0;
  wire f_u_dadda_cla32_fa380_xor1;
  wire f_u_dadda_cla32_fa380_and1;
  wire f_u_dadda_cla32_fa380_or0;
  wire f_u_dadda_cla32_fa381_xor0;
  wire f_u_dadda_cla32_fa381_and0;
  wire f_u_dadda_cla32_fa381_xor1;
  wire f_u_dadda_cla32_fa381_and1;
  wire f_u_dadda_cla32_fa381_or0;
  wire f_u_dadda_cla32_fa382_xor0;
  wire f_u_dadda_cla32_fa382_and0;
  wire f_u_dadda_cla32_fa382_xor1;
  wire f_u_dadda_cla32_fa382_and1;
  wire f_u_dadda_cla32_fa382_or0;
  wire f_u_dadda_cla32_fa383_xor0;
  wire f_u_dadda_cla32_fa383_and0;
  wire f_u_dadda_cla32_fa383_xor1;
  wire f_u_dadda_cla32_fa383_and1;
  wire f_u_dadda_cla32_fa383_or0;
  wire f_u_dadda_cla32_fa384_xor0;
  wire f_u_dadda_cla32_fa384_and0;
  wire f_u_dadda_cla32_fa384_xor1;
  wire f_u_dadda_cla32_fa384_and1;
  wire f_u_dadda_cla32_fa384_or0;
  wire f_u_dadda_cla32_and_28_6;
  wire f_u_dadda_cla32_and_27_7;
  wire f_u_dadda_cla32_fa385_xor0;
  wire f_u_dadda_cla32_fa385_and0;
  wire f_u_dadda_cla32_fa385_xor1;
  wire f_u_dadda_cla32_fa385_and1;
  wire f_u_dadda_cla32_fa385_or0;
  wire f_u_dadda_cla32_and_26_8;
  wire f_u_dadda_cla32_and_25_9;
  wire f_u_dadda_cla32_and_24_10;
  wire f_u_dadda_cla32_fa386_xor0;
  wire f_u_dadda_cla32_fa386_and0;
  wire f_u_dadda_cla32_fa386_xor1;
  wire f_u_dadda_cla32_fa386_and1;
  wire f_u_dadda_cla32_fa386_or0;
  wire f_u_dadda_cla32_and_23_11;
  wire f_u_dadda_cla32_and_22_12;
  wire f_u_dadda_cla32_and_21_13;
  wire f_u_dadda_cla32_fa387_xor0;
  wire f_u_dadda_cla32_fa387_and0;
  wire f_u_dadda_cla32_fa387_xor1;
  wire f_u_dadda_cla32_fa387_and1;
  wire f_u_dadda_cla32_fa387_or0;
  wire f_u_dadda_cla32_and_20_14;
  wire f_u_dadda_cla32_and_19_15;
  wire f_u_dadda_cla32_and_18_16;
  wire f_u_dadda_cla32_fa388_xor0;
  wire f_u_dadda_cla32_fa388_and0;
  wire f_u_dadda_cla32_fa388_xor1;
  wire f_u_dadda_cla32_fa388_and1;
  wire f_u_dadda_cla32_fa388_or0;
  wire f_u_dadda_cla32_and_17_17;
  wire f_u_dadda_cla32_and_16_18;
  wire f_u_dadda_cla32_and_15_19;
  wire f_u_dadda_cla32_fa389_xor0;
  wire f_u_dadda_cla32_fa389_and0;
  wire f_u_dadda_cla32_fa389_xor1;
  wire f_u_dadda_cla32_fa389_and1;
  wire f_u_dadda_cla32_fa389_or0;
  wire f_u_dadda_cla32_and_14_20;
  wire f_u_dadda_cla32_and_13_21;
  wire f_u_dadda_cla32_and_12_22;
  wire f_u_dadda_cla32_fa390_xor0;
  wire f_u_dadda_cla32_fa390_and0;
  wire f_u_dadda_cla32_fa390_xor1;
  wire f_u_dadda_cla32_fa390_and1;
  wire f_u_dadda_cla32_fa390_or0;
  wire f_u_dadda_cla32_and_11_23;
  wire f_u_dadda_cla32_and_10_24;
  wire f_u_dadda_cla32_and_9_25;
  wire f_u_dadda_cla32_fa391_xor0;
  wire f_u_dadda_cla32_fa391_and0;
  wire f_u_dadda_cla32_fa391_xor1;
  wire f_u_dadda_cla32_fa391_and1;
  wire f_u_dadda_cla32_fa391_or0;
  wire f_u_dadda_cla32_and_8_26;
  wire f_u_dadda_cla32_and_7_27;
  wire f_u_dadda_cla32_and_6_28;
  wire f_u_dadda_cla32_fa392_xor0;
  wire f_u_dadda_cla32_fa392_and0;
  wire f_u_dadda_cla32_fa392_xor1;
  wire f_u_dadda_cla32_fa392_and1;
  wire f_u_dadda_cla32_fa392_or0;
  wire f_u_dadda_cla32_and_5_29;
  wire f_u_dadda_cla32_and_4_30;
  wire f_u_dadda_cla32_and_3_31;
  wire f_u_dadda_cla32_fa393_xor0;
  wire f_u_dadda_cla32_fa393_and0;
  wire f_u_dadda_cla32_fa393_xor1;
  wire f_u_dadda_cla32_fa393_and1;
  wire f_u_dadda_cla32_fa393_or0;
  wire f_u_dadda_cla32_fa394_xor0;
  wire f_u_dadda_cla32_fa394_and0;
  wire f_u_dadda_cla32_fa394_xor1;
  wire f_u_dadda_cla32_fa394_and1;
  wire f_u_dadda_cla32_fa394_or0;
  wire f_u_dadda_cla32_fa395_xor0;
  wire f_u_dadda_cla32_fa395_and0;
  wire f_u_dadda_cla32_fa395_xor1;
  wire f_u_dadda_cla32_fa395_and1;
  wire f_u_dadda_cla32_fa395_or0;
  wire f_u_dadda_cla32_fa396_xor0;
  wire f_u_dadda_cla32_fa396_and0;
  wire f_u_dadda_cla32_fa396_xor1;
  wire f_u_dadda_cla32_fa396_and1;
  wire f_u_dadda_cla32_fa396_or0;
  wire f_u_dadda_cla32_fa397_xor0;
  wire f_u_dadda_cla32_fa397_and0;
  wire f_u_dadda_cla32_fa397_xor1;
  wire f_u_dadda_cla32_fa397_and1;
  wire f_u_dadda_cla32_fa397_or0;
  wire f_u_dadda_cla32_fa398_xor0;
  wire f_u_dadda_cla32_fa398_and0;
  wire f_u_dadda_cla32_fa398_xor1;
  wire f_u_dadda_cla32_fa398_and1;
  wire f_u_dadda_cla32_fa398_or0;
  wire f_u_dadda_cla32_fa399_xor0;
  wire f_u_dadda_cla32_fa399_and0;
  wire f_u_dadda_cla32_fa399_xor1;
  wire f_u_dadda_cla32_fa399_and1;
  wire f_u_dadda_cla32_fa399_or0;
  wire f_u_dadda_cla32_fa400_xor0;
  wire f_u_dadda_cla32_fa400_and0;
  wire f_u_dadda_cla32_fa400_xor1;
  wire f_u_dadda_cla32_fa400_and1;
  wire f_u_dadda_cla32_fa400_or0;
  wire f_u_dadda_cla32_fa401_xor0;
  wire f_u_dadda_cla32_fa401_and0;
  wire f_u_dadda_cla32_fa401_xor1;
  wire f_u_dadda_cla32_fa401_and1;
  wire f_u_dadda_cla32_fa401_or0;
  wire f_u_dadda_cla32_fa402_xor0;
  wire f_u_dadda_cla32_fa402_and0;
  wire f_u_dadda_cla32_fa402_xor1;
  wire f_u_dadda_cla32_fa402_and1;
  wire f_u_dadda_cla32_fa402_or0;
  wire f_u_dadda_cla32_fa403_xor0;
  wire f_u_dadda_cla32_fa403_and0;
  wire f_u_dadda_cla32_fa403_xor1;
  wire f_u_dadda_cla32_fa403_and1;
  wire f_u_dadda_cla32_fa403_or0;
  wire f_u_dadda_cla32_fa404_xor0;
  wire f_u_dadda_cla32_fa404_and0;
  wire f_u_dadda_cla32_fa404_xor1;
  wire f_u_dadda_cla32_fa404_and1;
  wire f_u_dadda_cla32_fa404_or0;
  wire f_u_dadda_cla32_fa405_xor0;
  wire f_u_dadda_cla32_fa405_and0;
  wire f_u_dadda_cla32_fa405_xor1;
  wire f_u_dadda_cla32_fa405_and1;
  wire f_u_dadda_cla32_fa405_or0;
  wire f_u_dadda_cla32_fa406_xor0;
  wire f_u_dadda_cla32_fa406_and0;
  wire f_u_dadda_cla32_fa406_xor1;
  wire f_u_dadda_cla32_fa406_and1;
  wire f_u_dadda_cla32_fa406_or0;
  wire f_u_dadda_cla32_and_30_5;
  wire f_u_dadda_cla32_and_29_6;
  wire f_u_dadda_cla32_fa407_xor0;
  wire f_u_dadda_cla32_fa407_and0;
  wire f_u_dadda_cla32_fa407_xor1;
  wire f_u_dadda_cla32_fa407_and1;
  wire f_u_dadda_cla32_fa407_or0;
  wire f_u_dadda_cla32_and_28_7;
  wire f_u_dadda_cla32_and_27_8;
  wire f_u_dadda_cla32_and_26_9;
  wire f_u_dadda_cla32_fa408_xor0;
  wire f_u_dadda_cla32_fa408_and0;
  wire f_u_dadda_cla32_fa408_xor1;
  wire f_u_dadda_cla32_fa408_and1;
  wire f_u_dadda_cla32_fa408_or0;
  wire f_u_dadda_cla32_and_25_10;
  wire f_u_dadda_cla32_and_24_11;
  wire f_u_dadda_cla32_and_23_12;
  wire f_u_dadda_cla32_fa409_xor0;
  wire f_u_dadda_cla32_fa409_and0;
  wire f_u_dadda_cla32_fa409_xor1;
  wire f_u_dadda_cla32_fa409_and1;
  wire f_u_dadda_cla32_fa409_or0;
  wire f_u_dadda_cla32_and_22_13;
  wire f_u_dadda_cla32_and_21_14;
  wire f_u_dadda_cla32_and_20_15;
  wire f_u_dadda_cla32_fa410_xor0;
  wire f_u_dadda_cla32_fa410_and0;
  wire f_u_dadda_cla32_fa410_xor1;
  wire f_u_dadda_cla32_fa410_and1;
  wire f_u_dadda_cla32_fa410_or0;
  wire f_u_dadda_cla32_and_19_16;
  wire f_u_dadda_cla32_and_18_17;
  wire f_u_dadda_cla32_and_17_18;
  wire f_u_dadda_cla32_fa411_xor0;
  wire f_u_dadda_cla32_fa411_and0;
  wire f_u_dadda_cla32_fa411_xor1;
  wire f_u_dadda_cla32_fa411_and1;
  wire f_u_dadda_cla32_fa411_or0;
  wire f_u_dadda_cla32_and_16_19;
  wire f_u_dadda_cla32_and_15_20;
  wire f_u_dadda_cla32_and_14_21;
  wire f_u_dadda_cla32_fa412_xor0;
  wire f_u_dadda_cla32_fa412_and0;
  wire f_u_dadda_cla32_fa412_xor1;
  wire f_u_dadda_cla32_fa412_and1;
  wire f_u_dadda_cla32_fa412_or0;
  wire f_u_dadda_cla32_and_13_22;
  wire f_u_dadda_cla32_and_12_23;
  wire f_u_dadda_cla32_and_11_24;
  wire f_u_dadda_cla32_fa413_xor0;
  wire f_u_dadda_cla32_fa413_and0;
  wire f_u_dadda_cla32_fa413_xor1;
  wire f_u_dadda_cla32_fa413_and1;
  wire f_u_dadda_cla32_fa413_or0;
  wire f_u_dadda_cla32_and_10_25;
  wire f_u_dadda_cla32_and_9_26;
  wire f_u_dadda_cla32_and_8_27;
  wire f_u_dadda_cla32_fa414_xor0;
  wire f_u_dadda_cla32_fa414_and0;
  wire f_u_dadda_cla32_fa414_xor1;
  wire f_u_dadda_cla32_fa414_and1;
  wire f_u_dadda_cla32_fa414_or0;
  wire f_u_dadda_cla32_and_7_28;
  wire f_u_dadda_cla32_and_6_29;
  wire f_u_dadda_cla32_and_5_30;
  wire f_u_dadda_cla32_fa415_xor0;
  wire f_u_dadda_cla32_fa415_and0;
  wire f_u_dadda_cla32_fa415_xor1;
  wire f_u_dadda_cla32_fa415_and1;
  wire f_u_dadda_cla32_fa415_or0;
  wire f_u_dadda_cla32_and_4_31;
  wire f_u_dadda_cla32_fa416_xor0;
  wire f_u_dadda_cla32_fa416_and0;
  wire f_u_dadda_cla32_fa416_xor1;
  wire f_u_dadda_cla32_fa416_and1;
  wire f_u_dadda_cla32_fa416_or0;
  wire f_u_dadda_cla32_fa417_xor0;
  wire f_u_dadda_cla32_fa417_and0;
  wire f_u_dadda_cla32_fa417_xor1;
  wire f_u_dadda_cla32_fa417_and1;
  wire f_u_dadda_cla32_fa417_or0;
  wire f_u_dadda_cla32_fa418_xor0;
  wire f_u_dadda_cla32_fa418_and0;
  wire f_u_dadda_cla32_fa418_xor1;
  wire f_u_dadda_cla32_fa418_and1;
  wire f_u_dadda_cla32_fa418_or0;
  wire f_u_dadda_cla32_fa419_xor0;
  wire f_u_dadda_cla32_fa419_and0;
  wire f_u_dadda_cla32_fa419_xor1;
  wire f_u_dadda_cla32_fa419_and1;
  wire f_u_dadda_cla32_fa419_or0;
  wire f_u_dadda_cla32_fa420_xor0;
  wire f_u_dadda_cla32_fa420_and0;
  wire f_u_dadda_cla32_fa420_xor1;
  wire f_u_dadda_cla32_fa420_and1;
  wire f_u_dadda_cla32_fa420_or0;
  wire f_u_dadda_cla32_fa421_xor0;
  wire f_u_dadda_cla32_fa421_and0;
  wire f_u_dadda_cla32_fa421_xor1;
  wire f_u_dadda_cla32_fa421_and1;
  wire f_u_dadda_cla32_fa421_or0;
  wire f_u_dadda_cla32_fa422_xor0;
  wire f_u_dadda_cla32_fa422_and0;
  wire f_u_dadda_cla32_fa422_xor1;
  wire f_u_dadda_cla32_fa422_and1;
  wire f_u_dadda_cla32_fa422_or0;
  wire f_u_dadda_cla32_fa423_xor0;
  wire f_u_dadda_cla32_fa423_and0;
  wire f_u_dadda_cla32_fa423_xor1;
  wire f_u_dadda_cla32_fa423_and1;
  wire f_u_dadda_cla32_fa423_or0;
  wire f_u_dadda_cla32_fa424_xor0;
  wire f_u_dadda_cla32_fa424_and0;
  wire f_u_dadda_cla32_fa424_xor1;
  wire f_u_dadda_cla32_fa424_and1;
  wire f_u_dadda_cla32_fa424_or0;
  wire f_u_dadda_cla32_fa425_xor0;
  wire f_u_dadda_cla32_fa425_and0;
  wire f_u_dadda_cla32_fa425_xor1;
  wire f_u_dadda_cla32_fa425_and1;
  wire f_u_dadda_cla32_fa425_or0;
  wire f_u_dadda_cla32_fa426_xor0;
  wire f_u_dadda_cla32_fa426_and0;
  wire f_u_dadda_cla32_fa426_xor1;
  wire f_u_dadda_cla32_fa426_and1;
  wire f_u_dadda_cla32_fa426_or0;
  wire f_u_dadda_cla32_fa427_xor0;
  wire f_u_dadda_cla32_fa427_and0;
  wire f_u_dadda_cla32_fa427_xor1;
  wire f_u_dadda_cla32_fa427_and1;
  wire f_u_dadda_cla32_fa427_or0;
  wire f_u_dadda_cla32_fa428_xor0;
  wire f_u_dadda_cla32_fa428_and0;
  wire f_u_dadda_cla32_fa428_xor1;
  wire f_u_dadda_cla32_fa428_and1;
  wire f_u_dadda_cla32_fa428_or0;
  wire f_u_dadda_cla32_and_31_5;
  wire f_u_dadda_cla32_fa429_xor0;
  wire f_u_dadda_cla32_fa429_and0;
  wire f_u_dadda_cla32_fa429_xor1;
  wire f_u_dadda_cla32_fa429_and1;
  wire f_u_dadda_cla32_fa429_or0;
  wire f_u_dadda_cla32_and_30_6;
  wire f_u_dadda_cla32_and_29_7;
  wire f_u_dadda_cla32_and_28_8;
  wire f_u_dadda_cla32_fa430_xor0;
  wire f_u_dadda_cla32_fa430_and0;
  wire f_u_dadda_cla32_fa430_xor1;
  wire f_u_dadda_cla32_fa430_and1;
  wire f_u_dadda_cla32_fa430_or0;
  wire f_u_dadda_cla32_and_27_9;
  wire f_u_dadda_cla32_and_26_10;
  wire f_u_dadda_cla32_and_25_11;
  wire f_u_dadda_cla32_fa431_xor0;
  wire f_u_dadda_cla32_fa431_and0;
  wire f_u_dadda_cla32_fa431_xor1;
  wire f_u_dadda_cla32_fa431_and1;
  wire f_u_dadda_cla32_fa431_or0;
  wire f_u_dadda_cla32_and_24_12;
  wire f_u_dadda_cla32_and_23_13;
  wire f_u_dadda_cla32_and_22_14;
  wire f_u_dadda_cla32_fa432_xor0;
  wire f_u_dadda_cla32_fa432_and0;
  wire f_u_dadda_cla32_fa432_xor1;
  wire f_u_dadda_cla32_fa432_and1;
  wire f_u_dadda_cla32_fa432_or0;
  wire f_u_dadda_cla32_and_21_15;
  wire f_u_dadda_cla32_and_20_16;
  wire f_u_dadda_cla32_and_19_17;
  wire f_u_dadda_cla32_fa433_xor0;
  wire f_u_dadda_cla32_fa433_and0;
  wire f_u_dadda_cla32_fa433_xor1;
  wire f_u_dadda_cla32_fa433_and1;
  wire f_u_dadda_cla32_fa433_or0;
  wire f_u_dadda_cla32_and_18_18;
  wire f_u_dadda_cla32_and_17_19;
  wire f_u_dadda_cla32_and_16_20;
  wire f_u_dadda_cla32_fa434_xor0;
  wire f_u_dadda_cla32_fa434_and0;
  wire f_u_dadda_cla32_fa434_xor1;
  wire f_u_dadda_cla32_fa434_and1;
  wire f_u_dadda_cla32_fa434_or0;
  wire f_u_dadda_cla32_and_15_21;
  wire f_u_dadda_cla32_and_14_22;
  wire f_u_dadda_cla32_and_13_23;
  wire f_u_dadda_cla32_fa435_xor0;
  wire f_u_dadda_cla32_fa435_and0;
  wire f_u_dadda_cla32_fa435_xor1;
  wire f_u_dadda_cla32_fa435_and1;
  wire f_u_dadda_cla32_fa435_or0;
  wire f_u_dadda_cla32_and_12_24;
  wire f_u_dadda_cla32_and_11_25;
  wire f_u_dadda_cla32_and_10_26;
  wire f_u_dadda_cla32_fa436_xor0;
  wire f_u_dadda_cla32_fa436_and0;
  wire f_u_dadda_cla32_fa436_xor1;
  wire f_u_dadda_cla32_fa436_and1;
  wire f_u_dadda_cla32_fa436_or0;
  wire f_u_dadda_cla32_and_9_27;
  wire f_u_dadda_cla32_and_8_28;
  wire f_u_dadda_cla32_and_7_29;
  wire f_u_dadda_cla32_fa437_xor0;
  wire f_u_dadda_cla32_fa437_and0;
  wire f_u_dadda_cla32_fa437_xor1;
  wire f_u_dadda_cla32_fa437_and1;
  wire f_u_dadda_cla32_fa437_or0;
  wire f_u_dadda_cla32_and_6_30;
  wire f_u_dadda_cla32_and_5_31;
  wire f_u_dadda_cla32_fa438_xor0;
  wire f_u_dadda_cla32_fa438_and0;
  wire f_u_dadda_cla32_fa438_xor1;
  wire f_u_dadda_cla32_fa438_and1;
  wire f_u_dadda_cla32_fa438_or0;
  wire f_u_dadda_cla32_fa439_xor0;
  wire f_u_dadda_cla32_fa439_and0;
  wire f_u_dadda_cla32_fa439_xor1;
  wire f_u_dadda_cla32_fa439_and1;
  wire f_u_dadda_cla32_fa439_or0;
  wire f_u_dadda_cla32_fa440_xor0;
  wire f_u_dadda_cla32_fa440_and0;
  wire f_u_dadda_cla32_fa440_xor1;
  wire f_u_dadda_cla32_fa440_and1;
  wire f_u_dadda_cla32_fa440_or0;
  wire f_u_dadda_cla32_fa441_xor0;
  wire f_u_dadda_cla32_fa441_and0;
  wire f_u_dadda_cla32_fa441_xor1;
  wire f_u_dadda_cla32_fa441_and1;
  wire f_u_dadda_cla32_fa441_or0;
  wire f_u_dadda_cla32_fa442_xor0;
  wire f_u_dadda_cla32_fa442_and0;
  wire f_u_dadda_cla32_fa442_xor1;
  wire f_u_dadda_cla32_fa442_and1;
  wire f_u_dadda_cla32_fa442_or0;
  wire f_u_dadda_cla32_fa443_xor0;
  wire f_u_dadda_cla32_fa443_and0;
  wire f_u_dadda_cla32_fa443_xor1;
  wire f_u_dadda_cla32_fa443_and1;
  wire f_u_dadda_cla32_fa443_or0;
  wire f_u_dadda_cla32_fa444_xor0;
  wire f_u_dadda_cla32_fa444_and0;
  wire f_u_dadda_cla32_fa444_xor1;
  wire f_u_dadda_cla32_fa444_and1;
  wire f_u_dadda_cla32_fa444_or0;
  wire f_u_dadda_cla32_fa445_xor0;
  wire f_u_dadda_cla32_fa445_and0;
  wire f_u_dadda_cla32_fa445_xor1;
  wire f_u_dadda_cla32_fa445_and1;
  wire f_u_dadda_cla32_fa445_or0;
  wire f_u_dadda_cla32_fa446_xor0;
  wire f_u_dadda_cla32_fa446_and0;
  wire f_u_dadda_cla32_fa446_xor1;
  wire f_u_dadda_cla32_fa446_and1;
  wire f_u_dadda_cla32_fa446_or0;
  wire f_u_dadda_cla32_fa447_xor0;
  wire f_u_dadda_cla32_fa447_and0;
  wire f_u_dadda_cla32_fa447_xor1;
  wire f_u_dadda_cla32_fa447_and1;
  wire f_u_dadda_cla32_fa447_or0;
  wire f_u_dadda_cla32_fa448_xor0;
  wire f_u_dadda_cla32_fa448_and0;
  wire f_u_dadda_cla32_fa448_xor1;
  wire f_u_dadda_cla32_fa448_and1;
  wire f_u_dadda_cla32_fa448_or0;
  wire f_u_dadda_cla32_fa449_xor0;
  wire f_u_dadda_cla32_fa449_and0;
  wire f_u_dadda_cla32_fa449_xor1;
  wire f_u_dadda_cla32_fa449_and1;
  wire f_u_dadda_cla32_fa449_or0;
  wire f_u_dadda_cla32_fa450_xor0;
  wire f_u_dadda_cla32_fa450_and0;
  wire f_u_dadda_cla32_fa450_xor1;
  wire f_u_dadda_cla32_fa450_and1;
  wire f_u_dadda_cla32_fa450_or0;
  wire f_u_dadda_cla32_and_31_6;
  wire f_u_dadda_cla32_and_30_7;
  wire f_u_dadda_cla32_fa451_xor0;
  wire f_u_dadda_cla32_fa451_and0;
  wire f_u_dadda_cla32_fa451_xor1;
  wire f_u_dadda_cla32_fa451_and1;
  wire f_u_dadda_cla32_fa451_or0;
  wire f_u_dadda_cla32_and_29_8;
  wire f_u_dadda_cla32_and_28_9;
  wire f_u_dadda_cla32_and_27_10;
  wire f_u_dadda_cla32_fa452_xor0;
  wire f_u_dadda_cla32_fa452_and0;
  wire f_u_dadda_cla32_fa452_xor1;
  wire f_u_dadda_cla32_fa452_and1;
  wire f_u_dadda_cla32_fa452_or0;
  wire f_u_dadda_cla32_and_26_11;
  wire f_u_dadda_cla32_and_25_12;
  wire f_u_dadda_cla32_and_24_13;
  wire f_u_dadda_cla32_fa453_xor0;
  wire f_u_dadda_cla32_fa453_and0;
  wire f_u_dadda_cla32_fa453_xor1;
  wire f_u_dadda_cla32_fa453_and1;
  wire f_u_dadda_cla32_fa453_or0;
  wire f_u_dadda_cla32_and_23_14;
  wire f_u_dadda_cla32_and_22_15;
  wire f_u_dadda_cla32_and_21_16;
  wire f_u_dadda_cla32_fa454_xor0;
  wire f_u_dadda_cla32_fa454_and0;
  wire f_u_dadda_cla32_fa454_xor1;
  wire f_u_dadda_cla32_fa454_and1;
  wire f_u_dadda_cla32_fa454_or0;
  wire f_u_dadda_cla32_and_20_17;
  wire f_u_dadda_cla32_and_19_18;
  wire f_u_dadda_cla32_and_18_19;
  wire f_u_dadda_cla32_fa455_xor0;
  wire f_u_dadda_cla32_fa455_and0;
  wire f_u_dadda_cla32_fa455_xor1;
  wire f_u_dadda_cla32_fa455_and1;
  wire f_u_dadda_cla32_fa455_or0;
  wire f_u_dadda_cla32_and_17_20;
  wire f_u_dadda_cla32_and_16_21;
  wire f_u_dadda_cla32_and_15_22;
  wire f_u_dadda_cla32_fa456_xor0;
  wire f_u_dadda_cla32_fa456_and0;
  wire f_u_dadda_cla32_fa456_xor1;
  wire f_u_dadda_cla32_fa456_and1;
  wire f_u_dadda_cla32_fa456_or0;
  wire f_u_dadda_cla32_and_14_23;
  wire f_u_dadda_cla32_and_13_24;
  wire f_u_dadda_cla32_and_12_25;
  wire f_u_dadda_cla32_fa457_xor0;
  wire f_u_dadda_cla32_fa457_and0;
  wire f_u_dadda_cla32_fa457_xor1;
  wire f_u_dadda_cla32_fa457_and1;
  wire f_u_dadda_cla32_fa457_or0;
  wire f_u_dadda_cla32_and_11_26;
  wire f_u_dadda_cla32_and_10_27;
  wire f_u_dadda_cla32_and_9_28;
  wire f_u_dadda_cla32_fa458_xor0;
  wire f_u_dadda_cla32_fa458_and0;
  wire f_u_dadda_cla32_fa458_xor1;
  wire f_u_dadda_cla32_fa458_and1;
  wire f_u_dadda_cla32_fa458_or0;
  wire f_u_dadda_cla32_and_8_29;
  wire f_u_dadda_cla32_and_7_30;
  wire f_u_dadda_cla32_and_6_31;
  wire f_u_dadda_cla32_fa459_xor0;
  wire f_u_dadda_cla32_fa459_and0;
  wire f_u_dadda_cla32_fa459_xor1;
  wire f_u_dadda_cla32_fa459_and1;
  wire f_u_dadda_cla32_fa459_or0;
  wire f_u_dadda_cla32_fa460_xor0;
  wire f_u_dadda_cla32_fa460_and0;
  wire f_u_dadda_cla32_fa460_xor1;
  wire f_u_dadda_cla32_fa460_and1;
  wire f_u_dadda_cla32_fa460_or0;
  wire f_u_dadda_cla32_fa461_xor0;
  wire f_u_dadda_cla32_fa461_and0;
  wire f_u_dadda_cla32_fa461_xor1;
  wire f_u_dadda_cla32_fa461_and1;
  wire f_u_dadda_cla32_fa461_or0;
  wire f_u_dadda_cla32_fa462_xor0;
  wire f_u_dadda_cla32_fa462_and0;
  wire f_u_dadda_cla32_fa462_xor1;
  wire f_u_dadda_cla32_fa462_and1;
  wire f_u_dadda_cla32_fa462_or0;
  wire f_u_dadda_cla32_fa463_xor0;
  wire f_u_dadda_cla32_fa463_and0;
  wire f_u_dadda_cla32_fa463_xor1;
  wire f_u_dadda_cla32_fa463_and1;
  wire f_u_dadda_cla32_fa463_or0;
  wire f_u_dadda_cla32_fa464_xor0;
  wire f_u_dadda_cla32_fa464_and0;
  wire f_u_dadda_cla32_fa464_xor1;
  wire f_u_dadda_cla32_fa464_and1;
  wire f_u_dadda_cla32_fa464_or0;
  wire f_u_dadda_cla32_fa465_xor0;
  wire f_u_dadda_cla32_fa465_and0;
  wire f_u_dadda_cla32_fa465_xor1;
  wire f_u_dadda_cla32_fa465_and1;
  wire f_u_dadda_cla32_fa465_or0;
  wire f_u_dadda_cla32_fa466_xor0;
  wire f_u_dadda_cla32_fa466_and0;
  wire f_u_dadda_cla32_fa466_xor1;
  wire f_u_dadda_cla32_fa466_and1;
  wire f_u_dadda_cla32_fa466_or0;
  wire f_u_dadda_cla32_fa467_xor0;
  wire f_u_dadda_cla32_fa467_and0;
  wire f_u_dadda_cla32_fa467_xor1;
  wire f_u_dadda_cla32_fa467_and1;
  wire f_u_dadda_cla32_fa467_or0;
  wire f_u_dadda_cla32_fa468_xor0;
  wire f_u_dadda_cla32_fa468_and0;
  wire f_u_dadda_cla32_fa468_xor1;
  wire f_u_dadda_cla32_fa468_and1;
  wire f_u_dadda_cla32_fa468_or0;
  wire f_u_dadda_cla32_fa469_xor0;
  wire f_u_dadda_cla32_fa469_and0;
  wire f_u_dadda_cla32_fa469_xor1;
  wire f_u_dadda_cla32_fa469_and1;
  wire f_u_dadda_cla32_fa469_or0;
  wire f_u_dadda_cla32_fa470_xor0;
  wire f_u_dadda_cla32_fa470_and0;
  wire f_u_dadda_cla32_fa470_xor1;
  wire f_u_dadda_cla32_fa470_and1;
  wire f_u_dadda_cla32_fa470_or0;
  wire f_u_dadda_cla32_fa471_xor0;
  wire f_u_dadda_cla32_fa471_and0;
  wire f_u_dadda_cla32_fa471_xor1;
  wire f_u_dadda_cla32_fa471_and1;
  wire f_u_dadda_cla32_fa471_or0;
  wire f_u_dadda_cla32_and_31_7;
  wire f_u_dadda_cla32_and_30_8;
  wire f_u_dadda_cla32_and_29_9;
  wire f_u_dadda_cla32_fa472_xor0;
  wire f_u_dadda_cla32_fa472_and0;
  wire f_u_dadda_cla32_fa472_xor1;
  wire f_u_dadda_cla32_fa472_and1;
  wire f_u_dadda_cla32_fa472_or0;
  wire f_u_dadda_cla32_and_28_10;
  wire f_u_dadda_cla32_and_27_11;
  wire f_u_dadda_cla32_and_26_12;
  wire f_u_dadda_cla32_fa473_xor0;
  wire f_u_dadda_cla32_fa473_and0;
  wire f_u_dadda_cla32_fa473_xor1;
  wire f_u_dadda_cla32_fa473_and1;
  wire f_u_dadda_cla32_fa473_or0;
  wire f_u_dadda_cla32_and_25_13;
  wire f_u_dadda_cla32_and_24_14;
  wire f_u_dadda_cla32_and_23_15;
  wire f_u_dadda_cla32_fa474_xor0;
  wire f_u_dadda_cla32_fa474_and0;
  wire f_u_dadda_cla32_fa474_xor1;
  wire f_u_dadda_cla32_fa474_and1;
  wire f_u_dadda_cla32_fa474_or0;
  wire f_u_dadda_cla32_and_22_16;
  wire f_u_dadda_cla32_and_21_17;
  wire f_u_dadda_cla32_and_20_18;
  wire f_u_dadda_cla32_fa475_xor0;
  wire f_u_dadda_cla32_fa475_and0;
  wire f_u_dadda_cla32_fa475_xor1;
  wire f_u_dadda_cla32_fa475_and1;
  wire f_u_dadda_cla32_fa475_or0;
  wire f_u_dadda_cla32_and_19_19;
  wire f_u_dadda_cla32_and_18_20;
  wire f_u_dadda_cla32_and_17_21;
  wire f_u_dadda_cla32_fa476_xor0;
  wire f_u_dadda_cla32_fa476_and0;
  wire f_u_dadda_cla32_fa476_xor1;
  wire f_u_dadda_cla32_fa476_and1;
  wire f_u_dadda_cla32_fa476_or0;
  wire f_u_dadda_cla32_and_16_22;
  wire f_u_dadda_cla32_and_15_23;
  wire f_u_dadda_cla32_and_14_24;
  wire f_u_dadda_cla32_fa477_xor0;
  wire f_u_dadda_cla32_fa477_and0;
  wire f_u_dadda_cla32_fa477_xor1;
  wire f_u_dadda_cla32_fa477_and1;
  wire f_u_dadda_cla32_fa477_or0;
  wire f_u_dadda_cla32_and_13_25;
  wire f_u_dadda_cla32_and_12_26;
  wire f_u_dadda_cla32_and_11_27;
  wire f_u_dadda_cla32_fa478_xor0;
  wire f_u_dadda_cla32_fa478_and0;
  wire f_u_dadda_cla32_fa478_xor1;
  wire f_u_dadda_cla32_fa478_and1;
  wire f_u_dadda_cla32_fa478_or0;
  wire f_u_dadda_cla32_and_10_28;
  wire f_u_dadda_cla32_and_9_29;
  wire f_u_dadda_cla32_and_8_30;
  wire f_u_dadda_cla32_fa479_xor0;
  wire f_u_dadda_cla32_fa479_and0;
  wire f_u_dadda_cla32_fa479_xor1;
  wire f_u_dadda_cla32_fa479_and1;
  wire f_u_dadda_cla32_fa479_or0;
  wire f_u_dadda_cla32_and_7_31;
  wire f_u_dadda_cla32_fa480_xor0;
  wire f_u_dadda_cla32_fa480_and0;
  wire f_u_dadda_cla32_fa480_xor1;
  wire f_u_dadda_cla32_fa480_and1;
  wire f_u_dadda_cla32_fa480_or0;
  wire f_u_dadda_cla32_fa481_xor0;
  wire f_u_dadda_cla32_fa481_and0;
  wire f_u_dadda_cla32_fa481_xor1;
  wire f_u_dadda_cla32_fa481_and1;
  wire f_u_dadda_cla32_fa481_or0;
  wire f_u_dadda_cla32_fa482_xor0;
  wire f_u_dadda_cla32_fa482_and0;
  wire f_u_dadda_cla32_fa482_xor1;
  wire f_u_dadda_cla32_fa482_and1;
  wire f_u_dadda_cla32_fa482_or0;
  wire f_u_dadda_cla32_fa483_xor0;
  wire f_u_dadda_cla32_fa483_and0;
  wire f_u_dadda_cla32_fa483_xor1;
  wire f_u_dadda_cla32_fa483_and1;
  wire f_u_dadda_cla32_fa483_or0;
  wire f_u_dadda_cla32_fa484_xor0;
  wire f_u_dadda_cla32_fa484_and0;
  wire f_u_dadda_cla32_fa484_xor1;
  wire f_u_dadda_cla32_fa484_and1;
  wire f_u_dadda_cla32_fa484_or0;
  wire f_u_dadda_cla32_fa485_xor0;
  wire f_u_dadda_cla32_fa485_and0;
  wire f_u_dadda_cla32_fa485_xor1;
  wire f_u_dadda_cla32_fa485_and1;
  wire f_u_dadda_cla32_fa485_or0;
  wire f_u_dadda_cla32_fa486_xor0;
  wire f_u_dadda_cla32_fa486_and0;
  wire f_u_dadda_cla32_fa486_xor1;
  wire f_u_dadda_cla32_fa486_and1;
  wire f_u_dadda_cla32_fa486_or0;
  wire f_u_dadda_cla32_fa487_xor0;
  wire f_u_dadda_cla32_fa487_and0;
  wire f_u_dadda_cla32_fa487_xor1;
  wire f_u_dadda_cla32_fa487_and1;
  wire f_u_dadda_cla32_fa487_or0;
  wire f_u_dadda_cla32_fa488_xor0;
  wire f_u_dadda_cla32_fa488_and0;
  wire f_u_dadda_cla32_fa488_xor1;
  wire f_u_dadda_cla32_fa488_and1;
  wire f_u_dadda_cla32_fa488_or0;
  wire f_u_dadda_cla32_fa489_xor0;
  wire f_u_dadda_cla32_fa489_and0;
  wire f_u_dadda_cla32_fa489_xor1;
  wire f_u_dadda_cla32_fa489_and1;
  wire f_u_dadda_cla32_fa489_or0;
  wire f_u_dadda_cla32_fa490_xor0;
  wire f_u_dadda_cla32_fa490_and0;
  wire f_u_dadda_cla32_fa490_xor1;
  wire f_u_dadda_cla32_fa490_and1;
  wire f_u_dadda_cla32_fa490_or0;
  wire f_u_dadda_cla32_and_31_8;
  wire f_u_dadda_cla32_fa491_xor0;
  wire f_u_dadda_cla32_fa491_and0;
  wire f_u_dadda_cla32_fa491_xor1;
  wire f_u_dadda_cla32_fa491_and1;
  wire f_u_dadda_cla32_fa491_or0;
  wire f_u_dadda_cla32_and_30_9;
  wire f_u_dadda_cla32_and_29_10;
  wire f_u_dadda_cla32_and_28_11;
  wire f_u_dadda_cla32_fa492_xor0;
  wire f_u_dadda_cla32_fa492_and0;
  wire f_u_dadda_cla32_fa492_xor1;
  wire f_u_dadda_cla32_fa492_and1;
  wire f_u_dadda_cla32_fa492_or0;
  wire f_u_dadda_cla32_and_27_12;
  wire f_u_dadda_cla32_and_26_13;
  wire f_u_dadda_cla32_and_25_14;
  wire f_u_dadda_cla32_fa493_xor0;
  wire f_u_dadda_cla32_fa493_and0;
  wire f_u_dadda_cla32_fa493_xor1;
  wire f_u_dadda_cla32_fa493_and1;
  wire f_u_dadda_cla32_fa493_or0;
  wire f_u_dadda_cla32_and_24_15;
  wire f_u_dadda_cla32_and_23_16;
  wire f_u_dadda_cla32_and_22_17;
  wire f_u_dadda_cla32_fa494_xor0;
  wire f_u_dadda_cla32_fa494_and0;
  wire f_u_dadda_cla32_fa494_xor1;
  wire f_u_dadda_cla32_fa494_and1;
  wire f_u_dadda_cla32_fa494_or0;
  wire f_u_dadda_cla32_and_21_18;
  wire f_u_dadda_cla32_and_20_19;
  wire f_u_dadda_cla32_and_19_20;
  wire f_u_dadda_cla32_fa495_xor0;
  wire f_u_dadda_cla32_fa495_and0;
  wire f_u_dadda_cla32_fa495_xor1;
  wire f_u_dadda_cla32_fa495_and1;
  wire f_u_dadda_cla32_fa495_or0;
  wire f_u_dadda_cla32_and_18_21;
  wire f_u_dadda_cla32_and_17_22;
  wire f_u_dadda_cla32_and_16_23;
  wire f_u_dadda_cla32_fa496_xor0;
  wire f_u_dadda_cla32_fa496_and0;
  wire f_u_dadda_cla32_fa496_xor1;
  wire f_u_dadda_cla32_fa496_and1;
  wire f_u_dadda_cla32_fa496_or0;
  wire f_u_dadda_cla32_and_15_24;
  wire f_u_dadda_cla32_and_14_25;
  wire f_u_dadda_cla32_and_13_26;
  wire f_u_dadda_cla32_fa497_xor0;
  wire f_u_dadda_cla32_fa497_and0;
  wire f_u_dadda_cla32_fa497_xor1;
  wire f_u_dadda_cla32_fa497_and1;
  wire f_u_dadda_cla32_fa497_or0;
  wire f_u_dadda_cla32_and_12_27;
  wire f_u_dadda_cla32_and_11_28;
  wire f_u_dadda_cla32_and_10_29;
  wire f_u_dadda_cla32_fa498_xor0;
  wire f_u_dadda_cla32_fa498_and0;
  wire f_u_dadda_cla32_fa498_xor1;
  wire f_u_dadda_cla32_fa498_and1;
  wire f_u_dadda_cla32_fa498_or0;
  wire f_u_dadda_cla32_and_9_30;
  wire f_u_dadda_cla32_and_8_31;
  wire f_u_dadda_cla32_fa499_xor0;
  wire f_u_dadda_cla32_fa499_and0;
  wire f_u_dadda_cla32_fa499_xor1;
  wire f_u_dadda_cla32_fa499_and1;
  wire f_u_dadda_cla32_fa499_or0;
  wire f_u_dadda_cla32_fa500_xor0;
  wire f_u_dadda_cla32_fa500_and0;
  wire f_u_dadda_cla32_fa500_xor1;
  wire f_u_dadda_cla32_fa500_and1;
  wire f_u_dadda_cla32_fa500_or0;
  wire f_u_dadda_cla32_fa501_xor0;
  wire f_u_dadda_cla32_fa501_and0;
  wire f_u_dadda_cla32_fa501_xor1;
  wire f_u_dadda_cla32_fa501_and1;
  wire f_u_dadda_cla32_fa501_or0;
  wire f_u_dadda_cla32_fa502_xor0;
  wire f_u_dadda_cla32_fa502_and0;
  wire f_u_dadda_cla32_fa502_xor1;
  wire f_u_dadda_cla32_fa502_and1;
  wire f_u_dadda_cla32_fa502_or0;
  wire f_u_dadda_cla32_fa503_xor0;
  wire f_u_dadda_cla32_fa503_and0;
  wire f_u_dadda_cla32_fa503_xor1;
  wire f_u_dadda_cla32_fa503_and1;
  wire f_u_dadda_cla32_fa503_or0;
  wire f_u_dadda_cla32_fa504_xor0;
  wire f_u_dadda_cla32_fa504_and0;
  wire f_u_dadda_cla32_fa504_xor1;
  wire f_u_dadda_cla32_fa504_and1;
  wire f_u_dadda_cla32_fa504_or0;
  wire f_u_dadda_cla32_fa505_xor0;
  wire f_u_dadda_cla32_fa505_and0;
  wire f_u_dadda_cla32_fa505_xor1;
  wire f_u_dadda_cla32_fa505_and1;
  wire f_u_dadda_cla32_fa505_or0;
  wire f_u_dadda_cla32_fa506_xor0;
  wire f_u_dadda_cla32_fa506_and0;
  wire f_u_dadda_cla32_fa506_xor1;
  wire f_u_dadda_cla32_fa506_and1;
  wire f_u_dadda_cla32_fa506_or0;
  wire f_u_dadda_cla32_fa507_xor0;
  wire f_u_dadda_cla32_fa507_and0;
  wire f_u_dadda_cla32_fa507_xor1;
  wire f_u_dadda_cla32_fa507_and1;
  wire f_u_dadda_cla32_fa507_or0;
  wire f_u_dadda_cla32_fa508_xor0;
  wire f_u_dadda_cla32_fa508_and0;
  wire f_u_dadda_cla32_fa508_xor1;
  wire f_u_dadda_cla32_fa508_and1;
  wire f_u_dadda_cla32_fa508_or0;
  wire f_u_dadda_cla32_fa509_xor0;
  wire f_u_dadda_cla32_fa509_and0;
  wire f_u_dadda_cla32_fa509_xor1;
  wire f_u_dadda_cla32_fa509_and1;
  wire f_u_dadda_cla32_fa509_or0;
  wire f_u_dadda_cla32_and_31_9;
  wire f_u_dadda_cla32_and_30_10;
  wire f_u_dadda_cla32_fa510_xor0;
  wire f_u_dadda_cla32_fa510_and0;
  wire f_u_dadda_cla32_fa510_xor1;
  wire f_u_dadda_cla32_fa510_and1;
  wire f_u_dadda_cla32_fa510_or0;
  wire f_u_dadda_cla32_and_29_11;
  wire f_u_dadda_cla32_and_28_12;
  wire f_u_dadda_cla32_and_27_13;
  wire f_u_dadda_cla32_fa511_xor0;
  wire f_u_dadda_cla32_fa511_and0;
  wire f_u_dadda_cla32_fa511_xor1;
  wire f_u_dadda_cla32_fa511_and1;
  wire f_u_dadda_cla32_fa511_or0;
  wire f_u_dadda_cla32_and_26_14;
  wire f_u_dadda_cla32_and_25_15;
  wire f_u_dadda_cla32_and_24_16;
  wire f_u_dadda_cla32_fa512_xor0;
  wire f_u_dadda_cla32_fa512_and0;
  wire f_u_dadda_cla32_fa512_xor1;
  wire f_u_dadda_cla32_fa512_and1;
  wire f_u_dadda_cla32_fa512_or0;
  wire f_u_dadda_cla32_and_23_17;
  wire f_u_dadda_cla32_and_22_18;
  wire f_u_dadda_cla32_and_21_19;
  wire f_u_dadda_cla32_fa513_xor0;
  wire f_u_dadda_cla32_fa513_and0;
  wire f_u_dadda_cla32_fa513_xor1;
  wire f_u_dadda_cla32_fa513_and1;
  wire f_u_dadda_cla32_fa513_or0;
  wire f_u_dadda_cla32_and_20_20;
  wire f_u_dadda_cla32_and_19_21;
  wire f_u_dadda_cla32_and_18_22;
  wire f_u_dadda_cla32_fa514_xor0;
  wire f_u_dadda_cla32_fa514_and0;
  wire f_u_dadda_cla32_fa514_xor1;
  wire f_u_dadda_cla32_fa514_and1;
  wire f_u_dadda_cla32_fa514_or0;
  wire f_u_dadda_cla32_and_17_23;
  wire f_u_dadda_cla32_and_16_24;
  wire f_u_dadda_cla32_and_15_25;
  wire f_u_dadda_cla32_fa515_xor0;
  wire f_u_dadda_cla32_fa515_and0;
  wire f_u_dadda_cla32_fa515_xor1;
  wire f_u_dadda_cla32_fa515_and1;
  wire f_u_dadda_cla32_fa515_or0;
  wire f_u_dadda_cla32_and_14_26;
  wire f_u_dadda_cla32_and_13_27;
  wire f_u_dadda_cla32_and_12_28;
  wire f_u_dadda_cla32_fa516_xor0;
  wire f_u_dadda_cla32_fa516_and0;
  wire f_u_dadda_cla32_fa516_xor1;
  wire f_u_dadda_cla32_fa516_and1;
  wire f_u_dadda_cla32_fa516_or0;
  wire f_u_dadda_cla32_and_11_29;
  wire f_u_dadda_cla32_and_10_30;
  wire f_u_dadda_cla32_and_9_31;
  wire f_u_dadda_cla32_fa517_xor0;
  wire f_u_dadda_cla32_fa517_and0;
  wire f_u_dadda_cla32_fa517_xor1;
  wire f_u_dadda_cla32_fa517_and1;
  wire f_u_dadda_cla32_fa517_or0;
  wire f_u_dadda_cla32_fa518_xor0;
  wire f_u_dadda_cla32_fa518_and0;
  wire f_u_dadda_cla32_fa518_xor1;
  wire f_u_dadda_cla32_fa518_and1;
  wire f_u_dadda_cla32_fa518_or0;
  wire f_u_dadda_cla32_fa519_xor0;
  wire f_u_dadda_cla32_fa519_and0;
  wire f_u_dadda_cla32_fa519_xor1;
  wire f_u_dadda_cla32_fa519_and1;
  wire f_u_dadda_cla32_fa519_or0;
  wire f_u_dadda_cla32_fa520_xor0;
  wire f_u_dadda_cla32_fa520_and0;
  wire f_u_dadda_cla32_fa520_xor1;
  wire f_u_dadda_cla32_fa520_and1;
  wire f_u_dadda_cla32_fa520_or0;
  wire f_u_dadda_cla32_fa521_xor0;
  wire f_u_dadda_cla32_fa521_and0;
  wire f_u_dadda_cla32_fa521_xor1;
  wire f_u_dadda_cla32_fa521_and1;
  wire f_u_dadda_cla32_fa521_or0;
  wire f_u_dadda_cla32_fa522_xor0;
  wire f_u_dadda_cla32_fa522_and0;
  wire f_u_dadda_cla32_fa522_xor1;
  wire f_u_dadda_cla32_fa522_and1;
  wire f_u_dadda_cla32_fa522_or0;
  wire f_u_dadda_cla32_fa523_xor0;
  wire f_u_dadda_cla32_fa523_and0;
  wire f_u_dadda_cla32_fa523_xor1;
  wire f_u_dadda_cla32_fa523_and1;
  wire f_u_dadda_cla32_fa523_or0;
  wire f_u_dadda_cla32_fa524_xor0;
  wire f_u_dadda_cla32_fa524_and0;
  wire f_u_dadda_cla32_fa524_xor1;
  wire f_u_dadda_cla32_fa524_and1;
  wire f_u_dadda_cla32_fa524_or0;
  wire f_u_dadda_cla32_fa525_xor0;
  wire f_u_dadda_cla32_fa525_and0;
  wire f_u_dadda_cla32_fa525_xor1;
  wire f_u_dadda_cla32_fa525_and1;
  wire f_u_dadda_cla32_fa525_or0;
  wire f_u_dadda_cla32_fa526_xor0;
  wire f_u_dadda_cla32_fa526_and0;
  wire f_u_dadda_cla32_fa526_xor1;
  wire f_u_dadda_cla32_fa526_and1;
  wire f_u_dadda_cla32_fa526_or0;
  wire f_u_dadda_cla32_fa527_xor0;
  wire f_u_dadda_cla32_fa527_and0;
  wire f_u_dadda_cla32_fa527_xor1;
  wire f_u_dadda_cla32_fa527_and1;
  wire f_u_dadda_cla32_fa527_or0;
  wire f_u_dadda_cla32_and_31_10;
  wire f_u_dadda_cla32_and_30_11;
  wire f_u_dadda_cla32_and_29_12;
  wire f_u_dadda_cla32_fa528_xor0;
  wire f_u_dadda_cla32_fa528_and0;
  wire f_u_dadda_cla32_fa528_xor1;
  wire f_u_dadda_cla32_fa528_and1;
  wire f_u_dadda_cla32_fa528_or0;
  wire f_u_dadda_cla32_and_28_13;
  wire f_u_dadda_cla32_and_27_14;
  wire f_u_dadda_cla32_and_26_15;
  wire f_u_dadda_cla32_fa529_xor0;
  wire f_u_dadda_cla32_fa529_and0;
  wire f_u_dadda_cla32_fa529_xor1;
  wire f_u_dadda_cla32_fa529_and1;
  wire f_u_dadda_cla32_fa529_or0;
  wire f_u_dadda_cla32_and_25_16;
  wire f_u_dadda_cla32_and_24_17;
  wire f_u_dadda_cla32_and_23_18;
  wire f_u_dadda_cla32_fa530_xor0;
  wire f_u_dadda_cla32_fa530_and0;
  wire f_u_dadda_cla32_fa530_xor1;
  wire f_u_dadda_cla32_fa530_and1;
  wire f_u_dadda_cla32_fa530_or0;
  wire f_u_dadda_cla32_and_22_19;
  wire f_u_dadda_cla32_and_21_20;
  wire f_u_dadda_cla32_and_20_21;
  wire f_u_dadda_cla32_fa531_xor0;
  wire f_u_dadda_cla32_fa531_and0;
  wire f_u_dadda_cla32_fa531_xor1;
  wire f_u_dadda_cla32_fa531_and1;
  wire f_u_dadda_cla32_fa531_or0;
  wire f_u_dadda_cla32_and_19_22;
  wire f_u_dadda_cla32_and_18_23;
  wire f_u_dadda_cla32_and_17_24;
  wire f_u_dadda_cla32_fa532_xor0;
  wire f_u_dadda_cla32_fa532_and0;
  wire f_u_dadda_cla32_fa532_xor1;
  wire f_u_dadda_cla32_fa532_and1;
  wire f_u_dadda_cla32_fa532_or0;
  wire f_u_dadda_cla32_and_16_25;
  wire f_u_dadda_cla32_and_15_26;
  wire f_u_dadda_cla32_and_14_27;
  wire f_u_dadda_cla32_fa533_xor0;
  wire f_u_dadda_cla32_fa533_and0;
  wire f_u_dadda_cla32_fa533_xor1;
  wire f_u_dadda_cla32_fa533_and1;
  wire f_u_dadda_cla32_fa533_or0;
  wire f_u_dadda_cla32_and_13_28;
  wire f_u_dadda_cla32_and_12_29;
  wire f_u_dadda_cla32_and_11_30;
  wire f_u_dadda_cla32_fa534_xor0;
  wire f_u_dadda_cla32_fa534_and0;
  wire f_u_dadda_cla32_fa534_xor1;
  wire f_u_dadda_cla32_fa534_and1;
  wire f_u_dadda_cla32_fa534_or0;
  wire f_u_dadda_cla32_and_10_31;
  wire f_u_dadda_cla32_fa535_xor0;
  wire f_u_dadda_cla32_fa535_and0;
  wire f_u_dadda_cla32_fa535_xor1;
  wire f_u_dadda_cla32_fa535_and1;
  wire f_u_dadda_cla32_fa535_or0;
  wire f_u_dadda_cla32_fa536_xor0;
  wire f_u_dadda_cla32_fa536_and0;
  wire f_u_dadda_cla32_fa536_xor1;
  wire f_u_dadda_cla32_fa536_and1;
  wire f_u_dadda_cla32_fa536_or0;
  wire f_u_dadda_cla32_fa537_xor0;
  wire f_u_dadda_cla32_fa537_and0;
  wire f_u_dadda_cla32_fa537_xor1;
  wire f_u_dadda_cla32_fa537_and1;
  wire f_u_dadda_cla32_fa537_or0;
  wire f_u_dadda_cla32_fa538_xor0;
  wire f_u_dadda_cla32_fa538_and0;
  wire f_u_dadda_cla32_fa538_xor1;
  wire f_u_dadda_cla32_fa538_and1;
  wire f_u_dadda_cla32_fa538_or0;
  wire f_u_dadda_cla32_fa539_xor0;
  wire f_u_dadda_cla32_fa539_and0;
  wire f_u_dadda_cla32_fa539_xor1;
  wire f_u_dadda_cla32_fa539_and1;
  wire f_u_dadda_cla32_fa539_or0;
  wire f_u_dadda_cla32_fa540_xor0;
  wire f_u_dadda_cla32_fa540_and0;
  wire f_u_dadda_cla32_fa540_xor1;
  wire f_u_dadda_cla32_fa540_and1;
  wire f_u_dadda_cla32_fa540_or0;
  wire f_u_dadda_cla32_fa541_xor0;
  wire f_u_dadda_cla32_fa541_and0;
  wire f_u_dadda_cla32_fa541_xor1;
  wire f_u_dadda_cla32_fa541_and1;
  wire f_u_dadda_cla32_fa541_or0;
  wire f_u_dadda_cla32_fa542_xor0;
  wire f_u_dadda_cla32_fa542_and0;
  wire f_u_dadda_cla32_fa542_xor1;
  wire f_u_dadda_cla32_fa542_and1;
  wire f_u_dadda_cla32_fa542_or0;
  wire f_u_dadda_cla32_fa543_xor0;
  wire f_u_dadda_cla32_fa543_and0;
  wire f_u_dadda_cla32_fa543_xor1;
  wire f_u_dadda_cla32_fa543_and1;
  wire f_u_dadda_cla32_fa543_or0;
  wire f_u_dadda_cla32_and_31_11;
  wire f_u_dadda_cla32_fa544_xor0;
  wire f_u_dadda_cla32_fa544_and0;
  wire f_u_dadda_cla32_fa544_xor1;
  wire f_u_dadda_cla32_fa544_and1;
  wire f_u_dadda_cla32_fa544_or0;
  wire f_u_dadda_cla32_and_30_12;
  wire f_u_dadda_cla32_and_29_13;
  wire f_u_dadda_cla32_and_28_14;
  wire f_u_dadda_cla32_fa545_xor0;
  wire f_u_dadda_cla32_fa545_and0;
  wire f_u_dadda_cla32_fa545_xor1;
  wire f_u_dadda_cla32_fa545_and1;
  wire f_u_dadda_cla32_fa545_or0;
  wire f_u_dadda_cla32_and_27_15;
  wire f_u_dadda_cla32_and_26_16;
  wire f_u_dadda_cla32_and_25_17;
  wire f_u_dadda_cla32_fa546_xor0;
  wire f_u_dadda_cla32_fa546_and0;
  wire f_u_dadda_cla32_fa546_xor1;
  wire f_u_dadda_cla32_fa546_and1;
  wire f_u_dadda_cla32_fa546_or0;
  wire f_u_dadda_cla32_and_24_18;
  wire f_u_dadda_cla32_and_23_19;
  wire f_u_dadda_cla32_and_22_20;
  wire f_u_dadda_cla32_fa547_xor0;
  wire f_u_dadda_cla32_fa547_and0;
  wire f_u_dadda_cla32_fa547_xor1;
  wire f_u_dadda_cla32_fa547_and1;
  wire f_u_dadda_cla32_fa547_or0;
  wire f_u_dadda_cla32_and_21_21;
  wire f_u_dadda_cla32_and_20_22;
  wire f_u_dadda_cla32_and_19_23;
  wire f_u_dadda_cla32_fa548_xor0;
  wire f_u_dadda_cla32_fa548_and0;
  wire f_u_dadda_cla32_fa548_xor1;
  wire f_u_dadda_cla32_fa548_and1;
  wire f_u_dadda_cla32_fa548_or0;
  wire f_u_dadda_cla32_and_18_24;
  wire f_u_dadda_cla32_and_17_25;
  wire f_u_dadda_cla32_and_16_26;
  wire f_u_dadda_cla32_fa549_xor0;
  wire f_u_dadda_cla32_fa549_and0;
  wire f_u_dadda_cla32_fa549_xor1;
  wire f_u_dadda_cla32_fa549_and1;
  wire f_u_dadda_cla32_fa549_or0;
  wire f_u_dadda_cla32_and_15_27;
  wire f_u_dadda_cla32_and_14_28;
  wire f_u_dadda_cla32_and_13_29;
  wire f_u_dadda_cla32_fa550_xor0;
  wire f_u_dadda_cla32_fa550_and0;
  wire f_u_dadda_cla32_fa550_xor1;
  wire f_u_dadda_cla32_fa550_and1;
  wire f_u_dadda_cla32_fa550_or0;
  wire f_u_dadda_cla32_and_12_30;
  wire f_u_dadda_cla32_and_11_31;
  wire f_u_dadda_cla32_fa551_xor0;
  wire f_u_dadda_cla32_fa551_and0;
  wire f_u_dadda_cla32_fa551_xor1;
  wire f_u_dadda_cla32_fa551_and1;
  wire f_u_dadda_cla32_fa551_or0;
  wire f_u_dadda_cla32_fa552_xor0;
  wire f_u_dadda_cla32_fa552_and0;
  wire f_u_dadda_cla32_fa552_xor1;
  wire f_u_dadda_cla32_fa552_and1;
  wire f_u_dadda_cla32_fa552_or0;
  wire f_u_dadda_cla32_fa553_xor0;
  wire f_u_dadda_cla32_fa553_and0;
  wire f_u_dadda_cla32_fa553_xor1;
  wire f_u_dadda_cla32_fa553_and1;
  wire f_u_dadda_cla32_fa553_or0;
  wire f_u_dadda_cla32_fa554_xor0;
  wire f_u_dadda_cla32_fa554_and0;
  wire f_u_dadda_cla32_fa554_xor1;
  wire f_u_dadda_cla32_fa554_and1;
  wire f_u_dadda_cla32_fa554_or0;
  wire f_u_dadda_cla32_fa555_xor0;
  wire f_u_dadda_cla32_fa555_and0;
  wire f_u_dadda_cla32_fa555_xor1;
  wire f_u_dadda_cla32_fa555_and1;
  wire f_u_dadda_cla32_fa555_or0;
  wire f_u_dadda_cla32_fa556_xor0;
  wire f_u_dadda_cla32_fa556_and0;
  wire f_u_dadda_cla32_fa556_xor1;
  wire f_u_dadda_cla32_fa556_and1;
  wire f_u_dadda_cla32_fa556_or0;
  wire f_u_dadda_cla32_fa557_xor0;
  wire f_u_dadda_cla32_fa557_and0;
  wire f_u_dadda_cla32_fa557_xor1;
  wire f_u_dadda_cla32_fa557_and1;
  wire f_u_dadda_cla32_fa557_or0;
  wire f_u_dadda_cla32_fa558_xor0;
  wire f_u_dadda_cla32_fa558_and0;
  wire f_u_dadda_cla32_fa558_xor1;
  wire f_u_dadda_cla32_fa558_and1;
  wire f_u_dadda_cla32_fa558_or0;
  wire f_u_dadda_cla32_fa559_xor0;
  wire f_u_dadda_cla32_fa559_and0;
  wire f_u_dadda_cla32_fa559_xor1;
  wire f_u_dadda_cla32_fa559_and1;
  wire f_u_dadda_cla32_fa559_or0;
  wire f_u_dadda_cla32_and_31_12;
  wire f_u_dadda_cla32_and_30_13;
  wire f_u_dadda_cla32_fa560_xor0;
  wire f_u_dadda_cla32_fa560_and0;
  wire f_u_dadda_cla32_fa560_xor1;
  wire f_u_dadda_cla32_fa560_and1;
  wire f_u_dadda_cla32_fa560_or0;
  wire f_u_dadda_cla32_and_29_14;
  wire f_u_dadda_cla32_and_28_15;
  wire f_u_dadda_cla32_and_27_16;
  wire f_u_dadda_cla32_fa561_xor0;
  wire f_u_dadda_cla32_fa561_and0;
  wire f_u_dadda_cla32_fa561_xor1;
  wire f_u_dadda_cla32_fa561_and1;
  wire f_u_dadda_cla32_fa561_or0;
  wire f_u_dadda_cla32_and_26_17;
  wire f_u_dadda_cla32_and_25_18;
  wire f_u_dadda_cla32_and_24_19;
  wire f_u_dadda_cla32_fa562_xor0;
  wire f_u_dadda_cla32_fa562_and0;
  wire f_u_dadda_cla32_fa562_xor1;
  wire f_u_dadda_cla32_fa562_and1;
  wire f_u_dadda_cla32_fa562_or0;
  wire f_u_dadda_cla32_and_23_20;
  wire f_u_dadda_cla32_and_22_21;
  wire f_u_dadda_cla32_and_21_22;
  wire f_u_dadda_cla32_fa563_xor0;
  wire f_u_dadda_cla32_fa563_and0;
  wire f_u_dadda_cla32_fa563_xor1;
  wire f_u_dadda_cla32_fa563_and1;
  wire f_u_dadda_cla32_fa563_or0;
  wire f_u_dadda_cla32_and_20_23;
  wire f_u_dadda_cla32_and_19_24;
  wire f_u_dadda_cla32_and_18_25;
  wire f_u_dadda_cla32_fa564_xor0;
  wire f_u_dadda_cla32_fa564_and0;
  wire f_u_dadda_cla32_fa564_xor1;
  wire f_u_dadda_cla32_fa564_and1;
  wire f_u_dadda_cla32_fa564_or0;
  wire f_u_dadda_cla32_and_17_26;
  wire f_u_dadda_cla32_and_16_27;
  wire f_u_dadda_cla32_and_15_28;
  wire f_u_dadda_cla32_fa565_xor0;
  wire f_u_dadda_cla32_fa565_and0;
  wire f_u_dadda_cla32_fa565_xor1;
  wire f_u_dadda_cla32_fa565_and1;
  wire f_u_dadda_cla32_fa565_or0;
  wire f_u_dadda_cla32_and_14_29;
  wire f_u_dadda_cla32_and_13_30;
  wire f_u_dadda_cla32_and_12_31;
  wire f_u_dadda_cla32_fa566_xor0;
  wire f_u_dadda_cla32_fa566_and0;
  wire f_u_dadda_cla32_fa566_xor1;
  wire f_u_dadda_cla32_fa566_and1;
  wire f_u_dadda_cla32_fa566_or0;
  wire f_u_dadda_cla32_fa567_xor0;
  wire f_u_dadda_cla32_fa567_and0;
  wire f_u_dadda_cla32_fa567_xor1;
  wire f_u_dadda_cla32_fa567_and1;
  wire f_u_dadda_cla32_fa567_or0;
  wire f_u_dadda_cla32_fa568_xor0;
  wire f_u_dadda_cla32_fa568_and0;
  wire f_u_dadda_cla32_fa568_xor1;
  wire f_u_dadda_cla32_fa568_and1;
  wire f_u_dadda_cla32_fa568_or0;
  wire f_u_dadda_cla32_fa569_xor0;
  wire f_u_dadda_cla32_fa569_and0;
  wire f_u_dadda_cla32_fa569_xor1;
  wire f_u_dadda_cla32_fa569_and1;
  wire f_u_dadda_cla32_fa569_or0;
  wire f_u_dadda_cla32_fa570_xor0;
  wire f_u_dadda_cla32_fa570_and0;
  wire f_u_dadda_cla32_fa570_xor1;
  wire f_u_dadda_cla32_fa570_and1;
  wire f_u_dadda_cla32_fa570_or0;
  wire f_u_dadda_cla32_fa571_xor0;
  wire f_u_dadda_cla32_fa571_and0;
  wire f_u_dadda_cla32_fa571_xor1;
  wire f_u_dadda_cla32_fa571_and1;
  wire f_u_dadda_cla32_fa571_or0;
  wire f_u_dadda_cla32_fa572_xor0;
  wire f_u_dadda_cla32_fa572_and0;
  wire f_u_dadda_cla32_fa572_xor1;
  wire f_u_dadda_cla32_fa572_and1;
  wire f_u_dadda_cla32_fa572_or0;
  wire f_u_dadda_cla32_fa573_xor0;
  wire f_u_dadda_cla32_fa573_and0;
  wire f_u_dadda_cla32_fa573_xor1;
  wire f_u_dadda_cla32_fa573_and1;
  wire f_u_dadda_cla32_fa573_or0;
  wire f_u_dadda_cla32_fa574_xor0;
  wire f_u_dadda_cla32_fa574_and0;
  wire f_u_dadda_cla32_fa574_xor1;
  wire f_u_dadda_cla32_fa574_and1;
  wire f_u_dadda_cla32_fa574_or0;
  wire f_u_dadda_cla32_and_31_13;
  wire f_u_dadda_cla32_and_30_14;
  wire f_u_dadda_cla32_and_29_15;
  wire f_u_dadda_cla32_fa575_xor0;
  wire f_u_dadda_cla32_fa575_and0;
  wire f_u_dadda_cla32_fa575_xor1;
  wire f_u_dadda_cla32_fa575_and1;
  wire f_u_dadda_cla32_fa575_or0;
  wire f_u_dadda_cla32_and_28_16;
  wire f_u_dadda_cla32_and_27_17;
  wire f_u_dadda_cla32_and_26_18;
  wire f_u_dadda_cla32_fa576_xor0;
  wire f_u_dadda_cla32_fa576_and0;
  wire f_u_dadda_cla32_fa576_xor1;
  wire f_u_dadda_cla32_fa576_and1;
  wire f_u_dadda_cla32_fa576_or0;
  wire f_u_dadda_cla32_and_25_19;
  wire f_u_dadda_cla32_and_24_20;
  wire f_u_dadda_cla32_and_23_21;
  wire f_u_dadda_cla32_fa577_xor0;
  wire f_u_dadda_cla32_fa577_and0;
  wire f_u_dadda_cla32_fa577_xor1;
  wire f_u_dadda_cla32_fa577_and1;
  wire f_u_dadda_cla32_fa577_or0;
  wire f_u_dadda_cla32_and_22_22;
  wire f_u_dadda_cla32_and_21_23;
  wire f_u_dadda_cla32_and_20_24;
  wire f_u_dadda_cla32_fa578_xor0;
  wire f_u_dadda_cla32_fa578_and0;
  wire f_u_dadda_cla32_fa578_xor1;
  wire f_u_dadda_cla32_fa578_and1;
  wire f_u_dadda_cla32_fa578_or0;
  wire f_u_dadda_cla32_and_19_25;
  wire f_u_dadda_cla32_and_18_26;
  wire f_u_dadda_cla32_and_17_27;
  wire f_u_dadda_cla32_fa579_xor0;
  wire f_u_dadda_cla32_fa579_and0;
  wire f_u_dadda_cla32_fa579_xor1;
  wire f_u_dadda_cla32_fa579_and1;
  wire f_u_dadda_cla32_fa579_or0;
  wire f_u_dadda_cla32_and_16_28;
  wire f_u_dadda_cla32_and_15_29;
  wire f_u_dadda_cla32_and_14_30;
  wire f_u_dadda_cla32_fa580_xor0;
  wire f_u_dadda_cla32_fa580_and0;
  wire f_u_dadda_cla32_fa580_xor1;
  wire f_u_dadda_cla32_fa580_and1;
  wire f_u_dadda_cla32_fa580_or0;
  wire f_u_dadda_cla32_and_13_31;
  wire f_u_dadda_cla32_fa581_xor0;
  wire f_u_dadda_cla32_fa581_and0;
  wire f_u_dadda_cla32_fa581_xor1;
  wire f_u_dadda_cla32_fa581_and1;
  wire f_u_dadda_cla32_fa581_or0;
  wire f_u_dadda_cla32_fa582_xor0;
  wire f_u_dadda_cla32_fa582_and0;
  wire f_u_dadda_cla32_fa582_xor1;
  wire f_u_dadda_cla32_fa582_and1;
  wire f_u_dadda_cla32_fa582_or0;
  wire f_u_dadda_cla32_fa583_xor0;
  wire f_u_dadda_cla32_fa583_and0;
  wire f_u_dadda_cla32_fa583_xor1;
  wire f_u_dadda_cla32_fa583_and1;
  wire f_u_dadda_cla32_fa583_or0;
  wire f_u_dadda_cla32_fa584_xor0;
  wire f_u_dadda_cla32_fa584_and0;
  wire f_u_dadda_cla32_fa584_xor1;
  wire f_u_dadda_cla32_fa584_and1;
  wire f_u_dadda_cla32_fa584_or0;
  wire f_u_dadda_cla32_fa585_xor0;
  wire f_u_dadda_cla32_fa585_and0;
  wire f_u_dadda_cla32_fa585_xor1;
  wire f_u_dadda_cla32_fa585_and1;
  wire f_u_dadda_cla32_fa585_or0;
  wire f_u_dadda_cla32_fa586_xor0;
  wire f_u_dadda_cla32_fa586_and0;
  wire f_u_dadda_cla32_fa586_xor1;
  wire f_u_dadda_cla32_fa586_and1;
  wire f_u_dadda_cla32_fa586_or0;
  wire f_u_dadda_cla32_fa587_xor0;
  wire f_u_dadda_cla32_fa587_and0;
  wire f_u_dadda_cla32_fa587_xor1;
  wire f_u_dadda_cla32_fa587_and1;
  wire f_u_dadda_cla32_fa587_or0;
  wire f_u_dadda_cla32_and_31_14;
  wire f_u_dadda_cla32_fa588_xor0;
  wire f_u_dadda_cla32_fa588_and0;
  wire f_u_dadda_cla32_fa588_xor1;
  wire f_u_dadda_cla32_fa588_and1;
  wire f_u_dadda_cla32_fa588_or0;
  wire f_u_dadda_cla32_and_30_15;
  wire f_u_dadda_cla32_and_29_16;
  wire f_u_dadda_cla32_and_28_17;
  wire f_u_dadda_cla32_fa589_xor0;
  wire f_u_dadda_cla32_fa589_and0;
  wire f_u_dadda_cla32_fa589_xor1;
  wire f_u_dadda_cla32_fa589_and1;
  wire f_u_dadda_cla32_fa589_or0;
  wire f_u_dadda_cla32_and_27_18;
  wire f_u_dadda_cla32_and_26_19;
  wire f_u_dadda_cla32_and_25_20;
  wire f_u_dadda_cla32_fa590_xor0;
  wire f_u_dadda_cla32_fa590_and0;
  wire f_u_dadda_cla32_fa590_xor1;
  wire f_u_dadda_cla32_fa590_and1;
  wire f_u_dadda_cla32_fa590_or0;
  wire f_u_dadda_cla32_and_24_21;
  wire f_u_dadda_cla32_and_23_22;
  wire f_u_dadda_cla32_and_22_23;
  wire f_u_dadda_cla32_fa591_xor0;
  wire f_u_dadda_cla32_fa591_and0;
  wire f_u_dadda_cla32_fa591_xor1;
  wire f_u_dadda_cla32_fa591_and1;
  wire f_u_dadda_cla32_fa591_or0;
  wire f_u_dadda_cla32_and_21_24;
  wire f_u_dadda_cla32_and_20_25;
  wire f_u_dadda_cla32_and_19_26;
  wire f_u_dadda_cla32_fa592_xor0;
  wire f_u_dadda_cla32_fa592_and0;
  wire f_u_dadda_cla32_fa592_xor1;
  wire f_u_dadda_cla32_fa592_and1;
  wire f_u_dadda_cla32_fa592_or0;
  wire f_u_dadda_cla32_and_18_27;
  wire f_u_dadda_cla32_and_17_28;
  wire f_u_dadda_cla32_and_16_29;
  wire f_u_dadda_cla32_fa593_xor0;
  wire f_u_dadda_cla32_fa593_and0;
  wire f_u_dadda_cla32_fa593_xor1;
  wire f_u_dadda_cla32_fa593_and1;
  wire f_u_dadda_cla32_fa593_or0;
  wire f_u_dadda_cla32_and_15_30;
  wire f_u_dadda_cla32_and_14_31;
  wire f_u_dadda_cla32_fa594_xor0;
  wire f_u_dadda_cla32_fa594_and0;
  wire f_u_dadda_cla32_fa594_xor1;
  wire f_u_dadda_cla32_fa594_and1;
  wire f_u_dadda_cla32_fa594_or0;
  wire f_u_dadda_cla32_fa595_xor0;
  wire f_u_dadda_cla32_fa595_and0;
  wire f_u_dadda_cla32_fa595_xor1;
  wire f_u_dadda_cla32_fa595_and1;
  wire f_u_dadda_cla32_fa595_or0;
  wire f_u_dadda_cla32_fa596_xor0;
  wire f_u_dadda_cla32_fa596_and0;
  wire f_u_dadda_cla32_fa596_xor1;
  wire f_u_dadda_cla32_fa596_and1;
  wire f_u_dadda_cla32_fa596_or0;
  wire f_u_dadda_cla32_fa597_xor0;
  wire f_u_dadda_cla32_fa597_and0;
  wire f_u_dadda_cla32_fa597_xor1;
  wire f_u_dadda_cla32_fa597_and1;
  wire f_u_dadda_cla32_fa597_or0;
  wire f_u_dadda_cla32_fa598_xor0;
  wire f_u_dadda_cla32_fa598_and0;
  wire f_u_dadda_cla32_fa598_xor1;
  wire f_u_dadda_cla32_fa598_and1;
  wire f_u_dadda_cla32_fa598_or0;
  wire f_u_dadda_cla32_fa599_xor0;
  wire f_u_dadda_cla32_fa599_and0;
  wire f_u_dadda_cla32_fa599_xor1;
  wire f_u_dadda_cla32_fa599_and1;
  wire f_u_dadda_cla32_fa599_or0;
  wire f_u_dadda_cla32_fa600_xor0;
  wire f_u_dadda_cla32_fa600_and0;
  wire f_u_dadda_cla32_fa600_xor1;
  wire f_u_dadda_cla32_fa600_and1;
  wire f_u_dadda_cla32_fa600_or0;
  wire f_u_dadda_cla32_and_31_15;
  wire f_u_dadda_cla32_and_30_16;
  wire f_u_dadda_cla32_fa601_xor0;
  wire f_u_dadda_cla32_fa601_and0;
  wire f_u_dadda_cla32_fa601_xor1;
  wire f_u_dadda_cla32_fa601_and1;
  wire f_u_dadda_cla32_fa601_or0;
  wire f_u_dadda_cla32_and_29_17;
  wire f_u_dadda_cla32_and_28_18;
  wire f_u_dadda_cla32_and_27_19;
  wire f_u_dadda_cla32_fa602_xor0;
  wire f_u_dadda_cla32_fa602_and0;
  wire f_u_dadda_cla32_fa602_xor1;
  wire f_u_dadda_cla32_fa602_and1;
  wire f_u_dadda_cla32_fa602_or0;
  wire f_u_dadda_cla32_and_26_20;
  wire f_u_dadda_cla32_and_25_21;
  wire f_u_dadda_cla32_and_24_22;
  wire f_u_dadda_cla32_fa603_xor0;
  wire f_u_dadda_cla32_fa603_and0;
  wire f_u_dadda_cla32_fa603_xor1;
  wire f_u_dadda_cla32_fa603_and1;
  wire f_u_dadda_cla32_fa603_or0;
  wire f_u_dadda_cla32_and_23_23;
  wire f_u_dadda_cla32_and_22_24;
  wire f_u_dadda_cla32_and_21_25;
  wire f_u_dadda_cla32_fa604_xor0;
  wire f_u_dadda_cla32_fa604_and0;
  wire f_u_dadda_cla32_fa604_xor1;
  wire f_u_dadda_cla32_fa604_and1;
  wire f_u_dadda_cla32_fa604_or0;
  wire f_u_dadda_cla32_and_20_26;
  wire f_u_dadda_cla32_and_19_27;
  wire f_u_dadda_cla32_and_18_28;
  wire f_u_dadda_cla32_fa605_xor0;
  wire f_u_dadda_cla32_fa605_and0;
  wire f_u_dadda_cla32_fa605_xor1;
  wire f_u_dadda_cla32_fa605_and1;
  wire f_u_dadda_cla32_fa605_or0;
  wire f_u_dadda_cla32_and_17_29;
  wire f_u_dadda_cla32_and_16_30;
  wire f_u_dadda_cla32_and_15_31;
  wire f_u_dadda_cla32_fa606_xor0;
  wire f_u_dadda_cla32_fa606_and0;
  wire f_u_dadda_cla32_fa606_xor1;
  wire f_u_dadda_cla32_fa606_and1;
  wire f_u_dadda_cla32_fa606_or0;
  wire f_u_dadda_cla32_fa607_xor0;
  wire f_u_dadda_cla32_fa607_and0;
  wire f_u_dadda_cla32_fa607_xor1;
  wire f_u_dadda_cla32_fa607_and1;
  wire f_u_dadda_cla32_fa607_or0;
  wire f_u_dadda_cla32_fa608_xor0;
  wire f_u_dadda_cla32_fa608_and0;
  wire f_u_dadda_cla32_fa608_xor1;
  wire f_u_dadda_cla32_fa608_and1;
  wire f_u_dadda_cla32_fa608_or0;
  wire f_u_dadda_cla32_fa609_xor0;
  wire f_u_dadda_cla32_fa609_and0;
  wire f_u_dadda_cla32_fa609_xor1;
  wire f_u_dadda_cla32_fa609_and1;
  wire f_u_dadda_cla32_fa609_or0;
  wire f_u_dadda_cla32_fa610_xor0;
  wire f_u_dadda_cla32_fa610_and0;
  wire f_u_dadda_cla32_fa610_xor1;
  wire f_u_dadda_cla32_fa610_and1;
  wire f_u_dadda_cla32_fa610_or0;
  wire f_u_dadda_cla32_fa611_xor0;
  wire f_u_dadda_cla32_fa611_and0;
  wire f_u_dadda_cla32_fa611_xor1;
  wire f_u_dadda_cla32_fa611_and1;
  wire f_u_dadda_cla32_fa611_or0;
  wire f_u_dadda_cla32_fa612_xor0;
  wire f_u_dadda_cla32_fa612_and0;
  wire f_u_dadda_cla32_fa612_xor1;
  wire f_u_dadda_cla32_fa612_and1;
  wire f_u_dadda_cla32_fa612_or0;
  wire f_u_dadda_cla32_and_31_16;
  wire f_u_dadda_cla32_and_30_17;
  wire f_u_dadda_cla32_and_29_18;
  wire f_u_dadda_cla32_fa613_xor0;
  wire f_u_dadda_cla32_fa613_and0;
  wire f_u_dadda_cla32_fa613_xor1;
  wire f_u_dadda_cla32_fa613_and1;
  wire f_u_dadda_cla32_fa613_or0;
  wire f_u_dadda_cla32_and_28_19;
  wire f_u_dadda_cla32_and_27_20;
  wire f_u_dadda_cla32_and_26_21;
  wire f_u_dadda_cla32_fa614_xor0;
  wire f_u_dadda_cla32_fa614_and0;
  wire f_u_dadda_cla32_fa614_xor1;
  wire f_u_dadda_cla32_fa614_and1;
  wire f_u_dadda_cla32_fa614_or0;
  wire f_u_dadda_cla32_and_25_22;
  wire f_u_dadda_cla32_and_24_23;
  wire f_u_dadda_cla32_and_23_24;
  wire f_u_dadda_cla32_fa615_xor0;
  wire f_u_dadda_cla32_fa615_and0;
  wire f_u_dadda_cla32_fa615_xor1;
  wire f_u_dadda_cla32_fa615_and1;
  wire f_u_dadda_cla32_fa615_or0;
  wire f_u_dadda_cla32_and_22_25;
  wire f_u_dadda_cla32_and_21_26;
  wire f_u_dadda_cla32_and_20_27;
  wire f_u_dadda_cla32_fa616_xor0;
  wire f_u_dadda_cla32_fa616_and0;
  wire f_u_dadda_cla32_fa616_xor1;
  wire f_u_dadda_cla32_fa616_and1;
  wire f_u_dadda_cla32_fa616_or0;
  wire f_u_dadda_cla32_and_19_28;
  wire f_u_dadda_cla32_and_18_29;
  wire f_u_dadda_cla32_and_17_30;
  wire f_u_dadda_cla32_fa617_xor0;
  wire f_u_dadda_cla32_fa617_and0;
  wire f_u_dadda_cla32_fa617_xor1;
  wire f_u_dadda_cla32_fa617_and1;
  wire f_u_dadda_cla32_fa617_or0;
  wire f_u_dadda_cla32_and_16_31;
  wire f_u_dadda_cla32_fa618_xor0;
  wire f_u_dadda_cla32_fa618_and0;
  wire f_u_dadda_cla32_fa618_xor1;
  wire f_u_dadda_cla32_fa618_and1;
  wire f_u_dadda_cla32_fa618_or0;
  wire f_u_dadda_cla32_fa619_xor0;
  wire f_u_dadda_cla32_fa619_and0;
  wire f_u_dadda_cla32_fa619_xor1;
  wire f_u_dadda_cla32_fa619_and1;
  wire f_u_dadda_cla32_fa619_or0;
  wire f_u_dadda_cla32_fa620_xor0;
  wire f_u_dadda_cla32_fa620_and0;
  wire f_u_dadda_cla32_fa620_xor1;
  wire f_u_dadda_cla32_fa620_and1;
  wire f_u_dadda_cla32_fa620_or0;
  wire f_u_dadda_cla32_fa621_xor0;
  wire f_u_dadda_cla32_fa621_and0;
  wire f_u_dadda_cla32_fa621_xor1;
  wire f_u_dadda_cla32_fa621_and1;
  wire f_u_dadda_cla32_fa621_or0;
  wire f_u_dadda_cla32_fa622_xor0;
  wire f_u_dadda_cla32_fa622_and0;
  wire f_u_dadda_cla32_fa622_xor1;
  wire f_u_dadda_cla32_fa622_and1;
  wire f_u_dadda_cla32_fa622_or0;
  wire f_u_dadda_cla32_and_31_17;
  wire f_u_dadda_cla32_fa623_xor0;
  wire f_u_dadda_cla32_fa623_and0;
  wire f_u_dadda_cla32_fa623_xor1;
  wire f_u_dadda_cla32_fa623_and1;
  wire f_u_dadda_cla32_fa623_or0;
  wire f_u_dadda_cla32_and_30_18;
  wire f_u_dadda_cla32_and_29_19;
  wire f_u_dadda_cla32_and_28_20;
  wire f_u_dadda_cla32_fa624_xor0;
  wire f_u_dadda_cla32_fa624_and0;
  wire f_u_dadda_cla32_fa624_xor1;
  wire f_u_dadda_cla32_fa624_and1;
  wire f_u_dadda_cla32_fa624_or0;
  wire f_u_dadda_cla32_and_27_21;
  wire f_u_dadda_cla32_and_26_22;
  wire f_u_dadda_cla32_and_25_23;
  wire f_u_dadda_cla32_fa625_xor0;
  wire f_u_dadda_cla32_fa625_and0;
  wire f_u_dadda_cla32_fa625_xor1;
  wire f_u_dadda_cla32_fa625_and1;
  wire f_u_dadda_cla32_fa625_or0;
  wire f_u_dadda_cla32_and_24_24;
  wire f_u_dadda_cla32_and_23_25;
  wire f_u_dadda_cla32_and_22_26;
  wire f_u_dadda_cla32_fa626_xor0;
  wire f_u_dadda_cla32_fa626_and0;
  wire f_u_dadda_cla32_fa626_xor1;
  wire f_u_dadda_cla32_fa626_and1;
  wire f_u_dadda_cla32_fa626_or0;
  wire f_u_dadda_cla32_and_21_27;
  wire f_u_dadda_cla32_and_20_28;
  wire f_u_dadda_cla32_and_19_29;
  wire f_u_dadda_cla32_fa627_xor0;
  wire f_u_dadda_cla32_fa627_and0;
  wire f_u_dadda_cla32_fa627_xor1;
  wire f_u_dadda_cla32_fa627_and1;
  wire f_u_dadda_cla32_fa627_or0;
  wire f_u_dadda_cla32_and_18_30;
  wire f_u_dadda_cla32_and_17_31;
  wire f_u_dadda_cla32_fa628_xor0;
  wire f_u_dadda_cla32_fa628_and0;
  wire f_u_dadda_cla32_fa628_xor1;
  wire f_u_dadda_cla32_fa628_and1;
  wire f_u_dadda_cla32_fa628_or0;
  wire f_u_dadda_cla32_fa629_xor0;
  wire f_u_dadda_cla32_fa629_and0;
  wire f_u_dadda_cla32_fa629_xor1;
  wire f_u_dadda_cla32_fa629_and1;
  wire f_u_dadda_cla32_fa629_or0;
  wire f_u_dadda_cla32_fa630_xor0;
  wire f_u_dadda_cla32_fa630_and0;
  wire f_u_dadda_cla32_fa630_xor1;
  wire f_u_dadda_cla32_fa630_and1;
  wire f_u_dadda_cla32_fa630_or0;
  wire f_u_dadda_cla32_fa631_xor0;
  wire f_u_dadda_cla32_fa631_and0;
  wire f_u_dadda_cla32_fa631_xor1;
  wire f_u_dadda_cla32_fa631_and1;
  wire f_u_dadda_cla32_fa631_or0;
  wire f_u_dadda_cla32_fa632_xor0;
  wire f_u_dadda_cla32_fa632_and0;
  wire f_u_dadda_cla32_fa632_xor1;
  wire f_u_dadda_cla32_fa632_and1;
  wire f_u_dadda_cla32_fa632_or0;
  wire f_u_dadda_cla32_and_31_18;
  wire f_u_dadda_cla32_and_30_19;
  wire f_u_dadda_cla32_fa633_xor0;
  wire f_u_dadda_cla32_fa633_and0;
  wire f_u_dadda_cla32_fa633_xor1;
  wire f_u_dadda_cla32_fa633_and1;
  wire f_u_dadda_cla32_fa633_or0;
  wire f_u_dadda_cla32_and_29_20;
  wire f_u_dadda_cla32_and_28_21;
  wire f_u_dadda_cla32_and_27_22;
  wire f_u_dadda_cla32_fa634_xor0;
  wire f_u_dadda_cla32_fa634_and0;
  wire f_u_dadda_cla32_fa634_xor1;
  wire f_u_dadda_cla32_fa634_and1;
  wire f_u_dadda_cla32_fa634_or0;
  wire f_u_dadda_cla32_and_26_23;
  wire f_u_dadda_cla32_and_25_24;
  wire f_u_dadda_cla32_and_24_25;
  wire f_u_dadda_cla32_fa635_xor0;
  wire f_u_dadda_cla32_fa635_and0;
  wire f_u_dadda_cla32_fa635_xor1;
  wire f_u_dadda_cla32_fa635_and1;
  wire f_u_dadda_cla32_fa635_or0;
  wire f_u_dadda_cla32_and_23_26;
  wire f_u_dadda_cla32_and_22_27;
  wire f_u_dadda_cla32_and_21_28;
  wire f_u_dadda_cla32_fa636_xor0;
  wire f_u_dadda_cla32_fa636_and0;
  wire f_u_dadda_cla32_fa636_xor1;
  wire f_u_dadda_cla32_fa636_and1;
  wire f_u_dadda_cla32_fa636_or0;
  wire f_u_dadda_cla32_and_20_29;
  wire f_u_dadda_cla32_and_19_30;
  wire f_u_dadda_cla32_and_18_31;
  wire f_u_dadda_cla32_fa637_xor0;
  wire f_u_dadda_cla32_fa637_and0;
  wire f_u_dadda_cla32_fa637_xor1;
  wire f_u_dadda_cla32_fa637_and1;
  wire f_u_dadda_cla32_fa637_or0;
  wire f_u_dadda_cla32_fa638_xor0;
  wire f_u_dadda_cla32_fa638_and0;
  wire f_u_dadda_cla32_fa638_xor1;
  wire f_u_dadda_cla32_fa638_and1;
  wire f_u_dadda_cla32_fa638_or0;
  wire f_u_dadda_cla32_fa639_xor0;
  wire f_u_dadda_cla32_fa639_and0;
  wire f_u_dadda_cla32_fa639_xor1;
  wire f_u_dadda_cla32_fa639_and1;
  wire f_u_dadda_cla32_fa639_or0;
  wire f_u_dadda_cla32_fa640_xor0;
  wire f_u_dadda_cla32_fa640_and0;
  wire f_u_dadda_cla32_fa640_xor1;
  wire f_u_dadda_cla32_fa640_and1;
  wire f_u_dadda_cla32_fa640_or0;
  wire f_u_dadda_cla32_fa641_xor0;
  wire f_u_dadda_cla32_fa641_and0;
  wire f_u_dadda_cla32_fa641_xor1;
  wire f_u_dadda_cla32_fa641_and1;
  wire f_u_dadda_cla32_fa641_or0;
  wire f_u_dadda_cla32_and_31_19;
  wire f_u_dadda_cla32_and_30_20;
  wire f_u_dadda_cla32_and_29_21;
  wire f_u_dadda_cla32_fa642_xor0;
  wire f_u_dadda_cla32_fa642_and0;
  wire f_u_dadda_cla32_fa642_xor1;
  wire f_u_dadda_cla32_fa642_and1;
  wire f_u_dadda_cla32_fa642_or0;
  wire f_u_dadda_cla32_and_28_22;
  wire f_u_dadda_cla32_and_27_23;
  wire f_u_dadda_cla32_and_26_24;
  wire f_u_dadda_cla32_fa643_xor0;
  wire f_u_dadda_cla32_fa643_and0;
  wire f_u_dadda_cla32_fa643_xor1;
  wire f_u_dadda_cla32_fa643_and1;
  wire f_u_dadda_cla32_fa643_or0;
  wire f_u_dadda_cla32_and_25_25;
  wire f_u_dadda_cla32_and_24_26;
  wire f_u_dadda_cla32_and_23_27;
  wire f_u_dadda_cla32_fa644_xor0;
  wire f_u_dadda_cla32_fa644_and0;
  wire f_u_dadda_cla32_fa644_xor1;
  wire f_u_dadda_cla32_fa644_and1;
  wire f_u_dadda_cla32_fa644_or0;
  wire f_u_dadda_cla32_and_22_28;
  wire f_u_dadda_cla32_and_21_29;
  wire f_u_dadda_cla32_and_20_30;
  wire f_u_dadda_cla32_fa645_xor0;
  wire f_u_dadda_cla32_fa645_and0;
  wire f_u_dadda_cla32_fa645_xor1;
  wire f_u_dadda_cla32_fa645_and1;
  wire f_u_dadda_cla32_fa645_or0;
  wire f_u_dadda_cla32_and_19_31;
  wire f_u_dadda_cla32_fa646_xor0;
  wire f_u_dadda_cla32_fa646_and0;
  wire f_u_dadda_cla32_fa646_xor1;
  wire f_u_dadda_cla32_fa646_and1;
  wire f_u_dadda_cla32_fa646_or0;
  wire f_u_dadda_cla32_fa647_xor0;
  wire f_u_dadda_cla32_fa647_and0;
  wire f_u_dadda_cla32_fa647_xor1;
  wire f_u_dadda_cla32_fa647_and1;
  wire f_u_dadda_cla32_fa647_or0;
  wire f_u_dadda_cla32_fa648_xor0;
  wire f_u_dadda_cla32_fa648_and0;
  wire f_u_dadda_cla32_fa648_xor1;
  wire f_u_dadda_cla32_fa648_and1;
  wire f_u_dadda_cla32_fa648_or0;
  wire f_u_dadda_cla32_and_31_20;
  wire f_u_dadda_cla32_fa649_xor0;
  wire f_u_dadda_cla32_fa649_and0;
  wire f_u_dadda_cla32_fa649_xor1;
  wire f_u_dadda_cla32_fa649_and1;
  wire f_u_dadda_cla32_fa649_or0;
  wire f_u_dadda_cla32_and_30_21;
  wire f_u_dadda_cla32_and_29_22;
  wire f_u_dadda_cla32_and_28_23;
  wire f_u_dadda_cla32_fa650_xor0;
  wire f_u_dadda_cla32_fa650_and0;
  wire f_u_dadda_cla32_fa650_xor1;
  wire f_u_dadda_cla32_fa650_and1;
  wire f_u_dadda_cla32_fa650_or0;
  wire f_u_dadda_cla32_and_27_24;
  wire f_u_dadda_cla32_and_26_25;
  wire f_u_dadda_cla32_and_25_26;
  wire f_u_dadda_cla32_fa651_xor0;
  wire f_u_dadda_cla32_fa651_and0;
  wire f_u_dadda_cla32_fa651_xor1;
  wire f_u_dadda_cla32_fa651_and1;
  wire f_u_dadda_cla32_fa651_or0;
  wire f_u_dadda_cla32_and_24_27;
  wire f_u_dadda_cla32_and_23_28;
  wire f_u_dadda_cla32_and_22_29;
  wire f_u_dadda_cla32_fa652_xor0;
  wire f_u_dadda_cla32_fa652_and0;
  wire f_u_dadda_cla32_fa652_xor1;
  wire f_u_dadda_cla32_fa652_and1;
  wire f_u_dadda_cla32_fa652_or0;
  wire f_u_dadda_cla32_and_21_30;
  wire f_u_dadda_cla32_and_20_31;
  wire f_u_dadda_cla32_fa653_xor0;
  wire f_u_dadda_cla32_fa653_and0;
  wire f_u_dadda_cla32_fa653_xor1;
  wire f_u_dadda_cla32_fa653_and1;
  wire f_u_dadda_cla32_fa653_or0;
  wire f_u_dadda_cla32_fa654_xor0;
  wire f_u_dadda_cla32_fa654_and0;
  wire f_u_dadda_cla32_fa654_xor1;
  wire f_u_dadda_cla32_fa654_and1;
  wire f_u_dadda_cla32_fa654_or0;
  wire f_u_dadda_cla32_fa655_xor0;
  wire f_u_dadda_cla32_fa655_and0;
  wire f_u_dadda_cla32_fa655_xor1;
  wire f_u_dadda_cla32_fa655_and1;
  wire f_u_dadda_cla32_fa655_or0;
  wire f_u_dadda_cla32_and_31_21;
  wire f_u_dadda_cla32_and_30_22;
  wire f_u_dadda_cla32_fa656_xor0;
  wire f_u_dadda_cla32_fa656_and0;
  wire f_u_dadda_cla32_fa656_xor1;
  wire f_u_dadda_cla32_fa656_and1;
  wire f_u_dadda_cla32_fa656_or0;
  wire f_u_dadda_cla32_and_29_23;
  wire f_u_dadda_cla32_and_28_24;
  wire f_u_dadda_cla32_and_27_25;
  wire f_u_dadda_cla32_fa657_xor0;
  wire f_u_dadda_cla32_fa657_and0;
  wire f_u_dadda_cla32_fa657_xor1;
  wire f_u_dadda_cla32_fa657_and1;
  wire f_u_dadda_cla32_fa657_or0;
  wire f_u_dadda_cla32_and_26_26;
  wire f_u_dadda_cla32_and_25_27;
  wire f_u_dadda_cla32_and_24_28;
  wire f_u_dadda_cla32_fa658_xor0;
  wire f_u_dadda_cla32_fa658_and0;
  wire f_u_dadda_cla32_fa658_xor1;
  wire f_u_dadda_cla32_fa658_and1;
  wire f_u_dadda_cla32_fa658_or0;
  wire f_u_dadda_cla32_and_23_29;
  wire f_u_dadda_cla32_and_22_30;
  wire f_u_dadda_cla32_and_21_31;
  wire f_u_dadda_cla32_fa659_xor0;
  wire f_u_dadda_cla32_fa659_and0;
  wire f_u_dadda_cla32_fa659_xor1;
  wire f_u_dadda_cla32_fa659_and1;
  wire f_u_dadda_cla32_fa659_or0;
  wire f_u_dadda_cla32_fa660_xor0;
  wire f_u_dadda_cla32_fa660_and0;
  wire f_u_dadda_cla32_fa660_xor1;
  wire f_u_dadda_cla32_fa660_and1;
  wire f_u_dadda_cla32_fa660_or0;
  wire f_u_dadda_cla32_fa661_xor0;
  wire f_u_dadda_cla32_fa661_and0;
  wire f_u_dadda_cla32_fa661_xor1;
  wire f_u_dadda_cla32_fa661_and1;
  wire f_u_dadda_cla32_fa661_or0;
  wire f_u_dadda_cla32_and_31_22;
  wire f_u_dadda_cla32_and_30_23;
  wire f_u_dadda_cla32_and_29_24;
  wire f_u_dadda_cla32_fa662_xor0;
  wire f_u_dadda_cla32_fa662_and0;
  wire f_u_dadda_cla32_fa662_xor1;
  wire f_u_dadda_cla32_fa662_and1;
  wire f_u_dadda_cla32_fa662_or0;
  wire f_u_dadda_cla32_and_28_25;
  wire f_u_dadda_cla32_and_27_26;
  wire f_u_dadda_cla32_and_26_27;
  wire f_u_dadda_cla32_fa663_xor0;
  wire f_u_dadda_cla32_fa663_and0;
  wire f_u_dadda_cla32_fa663_xor1;
  wire f_u_dadda_cla32_fa663_and1;
  wire f_u_dadda_cla32_fa663_or0;
  wire f_u_dadda_cla32_and_25_28;
  wire f_u_dadda_cla32_and_24_29;
  wire f_u_dadda_cla32_and_23_30;
  wire f_u_dadda_cla32_fa664_xor0;
  wire f_u_dadda_cla32_fa664_and0;
  wire f_u_dadda_cla32_fa664_xor1;
  wire f_u_dadda_cla32_fa664_and1;
  wire f_u_dadda_cla32_fa664_or0;
  wire f_u_dadda_cla32_fa665_xor0;
  wire f_u_dadda_cla32_fa665_and0;
  wire f_u_dadda_cla32_fa665_xor1;
  wire f_u_dadda_cla32_fa665_and1;
  wire f_u_dadda_cla32_fa665_or0;
  wire f_u_dadda_cla32_and_31_23;
  wire f_u_dadda_cla32_fa666_xor0;
  wire f_u_dadda_cla32_fa666_and0;
  wire f_u_dadda_cla32_fa666_xor1;
  wire f_u_dadda_cla32_fa666_and1;
  wire f_u_dadda_cla32_fa666_or0;
  wire f_u_dadda_cla32_and_30_24;
  wire f_u_dadda_cla32_and_29_25;
  wire f_u_dadda_cla32_and_28_26;
  wire f_u_dadda_cla32_fa667_xor0;
  wire f_u_dadda_cla32_fa667_and0;
  wire f_u_dadda_cla32_fa667_xor1;
  wire f_u_dadda_cla32_fa667_and1;
  wire f_u_dadda_cla32_fa667_or0;
  wire f_u_dadda_cla32_and_27_27;
  wire f_u_dadda_cla32_and_26_28;
  wire f_u_dadda_cla32_and_25_29;
  wire f_u_dadda_cla32_fa668_xor0;
  wire f_u_dadda_cla32_fa668_and0;
  wire f_u_dadda_cla32_fa668_xor1;
  wire f_u_dadda_cla32_fa668_and1;
  wire f_u_dadda_cla32_fa668_or0;
  wire f_u_dadda_cla32_fa669_xor0;
  wire f_u_dadda_cla32_fa669_and0;
  wire f_u_dadda_cla32_fa669_xor1;
  wire f_u_dadda_cla32_fa669_and1;
  wire f_u_dadda_cla32_fa669_or0;
  wire f_u_dadda_cla32_and_31_24;
  wire f_u_dadda_cla32_and_30_25;
  wire f_u_dadda_cla32_fa670_xor0;
  wire f_u_dadda_cla32_fa670_and0;
  wire f_u_dadda_cla32_fa670_xor1;
  wire f_u_dadda_cla32_fa670_and1;
  wire f_u_dadda_cla32_fa670_or0;
  wire f_u_dadda_cla32_and_29_26;
  wire f_u_dadda_cla32_and_28_27;
  wire f_u_dadda_cla32_and_27_28;
  wire f_u_dadda_cla32_fa671_xor0;
  wire f_u_dadda_cla32_fa671_and0;
  wire f_u_dadda_cla32_fa671_xor1;
  wire f_u_dadda_cla32_fa671_and1;
  wire f_u_dadda_cla32_fa671_or0;
  wire f_u_dadda_cla32_fa672_xor0;
  wire f_u_dadda_cla32_fa672_and0;
  wire f_u_dadda_cla32_fa672_xor1;
  wire f_u_dadda_cla32_fa672_and1;
  wire f_u_dadda_cla32_fa672_or0;
  wire f_u_dadda_cla32_and_31_25;
  wire f_u_dadda_cla32_and_30_26;
  wire f_u_dadda_cla32_and_29_27;
  wire f_u_dadda_cla32_fa673_xor0;
  wire f_u_dadda_cla32_fa673_and0;
  wire f_u_dadda_cla32_fa673_xor1;
  wire f_u_dadda_cla32_fa673_and1;
  wire f_u_dadda_cla32_fa673_or0;
  wire f_u_dadda_cla32_and_31_26;
  wire f_u_dadda_cla32_fa674_xor0;
  wire f_u_dadda_cla32_fa674_and0;
  wire f_u_dadda_cla32_fa674_xor1;
  wire f_u_dadda_cla32_fa674_and1;
  wire f_u_dadda_cla32_fa674_or0;
  wire f_u_dadda_cla32_and_4_0;
  wire f_u_dadda_cla32_and_3_1;
  wire f_u_dadda_cla32_ha27_xor0;
  wire f_u_dadda_cla32_ha27_and0;
  wire f_u_dadda_cla32_and_5_0;
  wire f_u_dadda_cla32_and_4_1;
  wire f_u_dadda_cla32_fa675_xor0;
  wire f_u_dadda_cla32_fa675_and0;
  wire f_u_dadda_cla32_fa675_xor1;
  wire f_u_dadda_cla32_fa675_and1;
  wire f_u_dadda_cla32_fa675_or0;
  wire f_u_dadda_cla32_and_3_2;
  wire f_u_dadda_cla32_and_2_3;
  wire f_u_dadda_cla32_ha28_xor0;
  wire f_u_dadda_cla32_ha28_and0;
  wire f_u_dadda_cla32_and_4_2;
  wire f_u_dadda_cla32_fa676_xor0;
  wire f_u_dadda_cla32_fa676_and0;
  wire f_u_dadda_cla32_fa676_xor1;
  wire f_u_dadda_cla32_fa676_and1;
  wire f_u_dadda_cla32_fa676_or0;
  wire f_u_dadda_cla32_and_3_3;
  wire f_u_dadda_cla32_and_2_4;
  wire f_u_dadda_cla32_and_1_5;
  wire f_u_dadda_cla32_fa677_xor0;
  wire f_u_dadda_cla32_fa677_and0;
  wire f_u_dadda_cla32_fa677_xor1;
  wire f_u_dadda_cla32_fa677_and1;
  wire f_u_dadda_cla32_fa677_or0;
  wire f_u_dadda_cla32_and_3_4;
  wire f_u_dadda_cla32_fa678_xor0;
  wire f_u_dadda_cla32_fa678_and0;
  wire f_u_dadda_cla32_fa678_xor1;
  wire f_u_dadda_cla32_fa678_and1;
  wire f_u_dadda_cla32_fa678_or0;
  wire f_u_dadda_cla32_and_2_5;
  wire f_u_dadda_cla32_and_1_6;
  wire f_u_dadda_cla32_and_0_7;
  wire f_u_dadda_cla32_fa679_xor0;
  wire f_u_dadda_cla32_fa679_and0;
  wire f_u_dadda_cla32_fa679_xor1;
  wire f_u_dadda_cla32_fa679_and1;
  wire f_u_dadda_cla32_fa679_or0;
  wire f_u_dadda_cla32_and_2_6;
  wire f_u_dadda_cla32_fa680_xor0;
  wire f_u_dadda_cla32_fa680_and0;
  wire f_u_dadda_cla32_fa680_xor1;
  wire f_u_dadda_cla32_fa680_and1;
  wire f_u_dadda_cla32_fa680_or0;
  wire f_u_dadda_cla32_and_1_7;
  wire f_u_dadda_cla32_and_0_8;
  wire f_u_dadda_cla32_fa681_xor0;
  wire f_u_dadda_cla32_fa681_and0;
  wire f_u_dadda_cla32_fa681_xor1;
  wire f_u_dadda_cla32_fa681_and1;
  wire f_u_dadda_cla32_fa681_or0;
  wire f_u_dadda_cla32_and_1_8;
  wire f_u_dadda_cla32_fa682_xor0;
  wire f_u_dadda_cla32_fa682_and0;
  wire f_u_dadda_cla32_fa682_xor1;
  wire f_u_dadda_cla32_fa682_and1;
  wire f_u_dadda_cla32_fa682_or0;
  wire f_u_dadda_cla32_and_0_9;
  wire f_u_dadda_cla32_fa683_xor0;
  wire f_u_dadda_cla32_fa683_and0;
  wire f_u_dadda_cla32_fa683_xor1;
  wire f_u_dadda_cla32_fa683_and1;
  wire f_u_dadda_cla32_fa683_or0;
  wire f_u_dadda_cla32_and_0_10;
  wire f_u_dadda_cla32_fa684_xor0;
  wire f_u_dadda_cla32_fa684_and0;
  wire f_u_dadda_cla32_fa684_xor1;
  wire f_u_dadda_cla32_fa684_and1;
  wire f_u_dadda_cla32_fa684_or0;
  wire f_u_dadda_cla32_fa685_xor0;
  wire f_u_dadda_cla32_fa685_and0;
  wire f_u_dadda_cla32_fa685_xor1;
  wire f_u_dadda_cla32_fa685_and1;
  wire f_u_dadda_cla32_fa685_or0;
  wire f_u_dadda_cla32_fa686_xor0;
  wire f_u_dadda_cla32_fa686_and0;
  wire f_u_dadda_cla32_fa686_xor1;
  wire f_u_dadda_cla32_fa686_and1;
  wire f_u_dadda_cla32_fa686_or0;
  wire f_u_dadda_cla32_fa687_xor0;
  wire f_u_dadda_cla32_fa687_and0;
  wire f_u_dadda_cla32_fa687_xor1;
  wire f_u_dadda_cla32_fa687_and1;
  wire f_u_dadda_cla32_fa687_or0;
  wire f_u_dadda_cla32_fa688_xor0;
  wire f_u_dadda_cla32_fa688_and0;
  wire f_u_dadda_cla32_fa688_xor1;
  wire f_u_dadda_cla32_fa688_and1;
  wire f_u_dadda_cla32_fa688_or0;
  wire f_u_dadda_cla32_fa689_xor0;
  wire f_u_dadda_cla32_fa689_and0;
  wire f_u_dadda_cla32_fa689_xor1;
  wire f_u_dadda_cla32_fa689_and1;
  wire f_u_dadda_cla32_fa689_or0;
  wire f_u_dadda_cla32_fa690_xor0;
  wire f_u_dadda_cla32_fa690_and0;
  wire f_u_dadda_cla32_fa690_xor1;
  wire f_u_dadda_cla32_fa690_and1;
  wire f_u_dadda_cla32_fa690_or0;
  wire f_u_dadda_cla32_fa691_xor0;
  wire f_u_dadda_cla32_fa691_and0;
  wire f_u_dadda_cla32_fa691_xor1;
  wire f_u_dadda_cla32_fa691_and1;
  wire f_u_dadda_cla32_fa691_or0;
  wire f_u_dadda_cla32_fa692_xor0;
  wire f_u_dadda_cla32_fa692_and0;
  wire f_u_dadda_cla32_fa692_xor1;
  wire f_u_dadda_cla32_fa692_and1;
  wire f_u_dadda_cla32_fa692_or0;
  wire f_u_dadda_cla32_fa693_xor0;
  wire f_u_dadda_cla32_fa693_and0;
  wire f_u_dadda_cla32_fa693_xor1;
  wire f_u_dadda_cla32_fa693_and1;
  wire f_u_dadda_cla32_fa693_or0;
  wire f_u_dadda_cla32_fa694_xor0;
  wire f_u_dadda_cla32_fa694_and0;
  wire f_u_dadda_cla32_fa694_xor1;
  wire f_u_dadda_cla32_fa694_and1;
  wire f_u_dadda_cla32_fa694_or0;
  wire f_u_dadda_cla32_fa695_xor0;
  wire f_u_dadda_cla32_fa695_and0;
  wire f_u_dadda_cla32_fa695_xor1;
  wire f_u_dadda_cla32_fa695_and1;
  wire f_u_dadda_cla32_fa695_or0;
  wire f_u_dadda_cla32_fa696_xor0;
  wire f_u_dadda_cla32_fa696_and0;
  wire f_u_dadda_cla32_fa696_xor1;
  wire f_u_dadda_cla32_fa696_and1;
  wire f_u_dadda_cla32_fa696_or0;
  wire f_u_dadda_cla32_fa697_xor0;
  wire f_u_dadda_cla32_fa697_and0;
  wire f_u_dadda_cla32_fa697_xor1;
  wire f_u_dadda_cla32_fa697_and1;
  wire f_u_dadda_cla32_fa697_or0;
  wire f_u_dadda_cla32_fa698_xor0;
  wire f_u_dadda_cla32_fa698_and0;
  wire f_u_dadda_cla32_fa698_xor1;
  wire f_u_dadda_cla32_fa698_and1;
  wire f_u_dadda_cla32_fa698_or0;
  wire f_u_dadda_cla32_fa699_xor0;
  wire f_u_dadda_cla32_fa699_and0;
  wire f_u_dadda_cla32_fa699_xor1;
  wire f_u_dadda_cla32_fa699_and1;
  wire f_u_dadda_cla32_fa699_or0;
  wire f_u_dadda_cla32_fa700_xor0;
  wire f_u_dadda_cla32_fa700_and0;
  wire f_u_dadda_cla32_fa700_xor1;
  wire f_u_dadda_cla32_fa700_and1;
  wire f_u_dadda_cla32_fa700_or0;
  wire f_u_dadda_cla32_fa701_xor0;
  wire f_u_dadda_cla32_fa701_and0;
  wire f_u_dadda_cla32_fa701_xor1;
  wire f_u_dadda_cla32_fa701_and1;
  wire f_u_dadda_cla32_fa701_or0;
  wire f_u_dadda_cla32_fa702_xor0;
  wire f_u_dadda_cla32_fa702_and0;
  wire f_u_dadda_cla32_fa702_xor1;
  wire f_u_dadda_cla32_fa702_and1;
  wire f_u_dadda_cla32_fa702_or0;
  wire f_u_dadda_cla32_fa703_xor0;
  wire f_u_dadda_cla32_fa703_and0;
  wire f_u_dadda_cla32_fa703_xor1;
  wire f_u_dadda_cla32_fa703_and1;
  wire f_u_dadda_cla32_fa703_or0;
  wire f_u_dadda_cla32_fa704_xor0;
  wire f_u_dadda_cla32_fa704_and0;
  wire f_u_dadda_cla32_fa704_xor1;
  wire f_u_dadda_cla32_fa704_and1;
  wire f_u_dadda_cla32_fa704_or0;
  wire f_u_dadda_cla32_fa705_xor0;
  wire f_u_dadda_cla32_fa705_and0;
  wire f_u_dadda_cla32_fa705_xor1;
  wire f_u_dadda_cla32_fa705_and1;
  wire f_u_dadda_cla32_fa705_or0;
  wire f_u_dadda_cla32_fa706_xor0;
  wire f_u_dadda_cla32_fa706_and0;
  wire f_u_dadda_cla32_fa706_xor1;
  wire f_u_dadda_cla32_fa706_and1;
  wire f_u_dadda_cla32_fa706_or0;
  wire f_u_dadda_cla32_fa707_xor0;
  wire f_u_dadda_cla32_fa707_and0;
  wire f_u_dadda_cla32_fa707_xor1;
  wire f_u_dadda_cla32_fa707_and1;
  wire f_u_dadda_cla32_fa707_or0;
  wire f_u_dadda_cla32_fa708_xor0;
  wire f_u_dadda_cla32_fa708_and0;
  wire f_u_dadda_cla32_fa708_xor1;
  wire f_u_dadda_cla32_fa708_and1;
  wire f_u_dadda_cla32_fa708_or0;
  wire f_u_dadda_cla32_fa709_xor0;
  wire f_u_dadda_cla32_fa709_and0;
  wire f_u_dadda_cla32_fa709_xor1;
  wire f_u_dadda_cla32_fa709_and1;
  wire f_u_dadda_cla32_fa709_or0;
  wire f_u_dadda_cla32_fa710_xor0;
  wire f_u_dadda_cla32_fa710_and0;
  wire f_u_dadda_cla32_fa710_xor1;
  wire f_u_dadda_cla32_fa710_and1;
  wire f_u_dadda_cla32_fa710_or0;
  wire f_u_dadda_cla32_fa711_xor0;
  wire f_u_dadda_cla32_fa711_and0;
  wire f_u_dadda_cla32_fa711_xor1;
  wire f_u_dadda_cla32_fa711_and1;
  wire f_u_dadda_cla32_fa711_or0;
  wire f_u_dadda_cla32_fa712_xor0;
  wire f_u_dadda_cla32_fa712_and0;
  wire f_u_dadda_cla32_fa712_xor1;
  wire f_u_dadda_cla32_fa712_and1;
  wire f_u_dadda_cla32_fa712_or0;
  wire f_u_dadda_cla32_fa713_xor0;
  wire f_u_dadda_cla32_fa713_and0;
  wire f_u_dadda_cla32_fa713_xor1;
  wire f_u_dadda_cla32_fa713_and1;
  wire f_u_dadda_cla32_fa713_or0;
  wire f_u_dadda_cla32_fa714_xor0;
  wire f_u_dadda_cla32_fa714_and0;
  wire f_u_dadda_cla32_fa714_xor1;
  wire f_u_dadda_cla32_fa714_and1;
  wire f_u_dadda_cla32_fa714_or0;
  wire f_u_dadda_cla32_fa715_xor0;
  wire f_u_dadda_cla32_fa715_and0;
  wire f_u_dadda_cla32_fa715_xor1;
  wire f_u_dadda_cla32_fa715_and1;
  wire f_u_dadda_cla32_fa715_or0;
  wire f_u_dadda_cla32_fa716_xor0;
  wire f_u_dadda_cla32_fa716_and0;
  wire f_u_dadda_cla32_fa716_xor1;
  wire f_u_dadda_cla32_fa716_and1;
  wire f_u_dadda_cla32_fa716_or0;
  wire f_u_dadda_cla32_fa717_xor0;
  wire f_u_dadda_cla32_fa717_and0;
  wire f_u_dadda_cla32_fa717_xor1;
  wire f_u_dadda_cla32_fa717_and1;
  wire f_u_dadda_cla32_fa717_or0;
  wire f_u_dadda_cla32_fa718_xor0;
  wire f_u_dadda_cla32_fa718_and0;
  wire f_u_dadda_cla32_fa718_xor1;
  wire f_u_dadda_cla32_fa718_and1;
  wire f_u_dadda_cla32_fa718_or0;
  wire f_u_dadda_cla32_fa719_xor0;
  wire f_u_dadda_cla32_fa719_and0;
  wire f_u_dadda_cla32_fa719_xor1;
  wire f_u_dadda_cla32_fa719_and1;
  wire f_u_dadda_cla32_fa719_or0;
  wire f_u_dadda_cla32_fa720_xor0;
  wire f_u_dadda_cla32_fa720_and0;
  wire f_u_dadda_cla32_fa720_xor1;
  wire f_u_dadda_cla32_fa720_and1;
  wire f_u_dadda_cla32_fa720_or0;
  wire f_u_dadda_cla32_fa721_xor0;
  wire f_u_dadda_cla32_fa721_and0;
  wire f_u_dadda_cla32_fa721_xor1;
  wire f_u_dadda_cla32_fa721_and1;
  wire f_u_dadda_cla32_fa721_or0;
  wire f_u_dadda_cla32_fa722_xor0;
  wire f_u_dadda_cla32_fa722_and0;
  wire f_u_dadda_cla32_fa722_xor1;
  wire f_u_dadda_cla32_fa722_and1;
  wire f_u_dadda_cla32_fa722_or0;
  wire f_u_dadda_cla32_fa723_xor0;
  wire f_u_dadda_cla32_fa723_and0;
  wire f_u_dadda_cla32_fa723_xor1;
  wire f_u_dadda_cla32_fa723_and1;
  wire f_u_dadda_cla32_fa723_or0;
  wire f_u_dadda_cla32_fa724_xor0;
  wire f_u_dadda_cla32_fa724_and0;
  wire f_u_dadda_cla32_fa724_xor1;
  wire f_u_dadda_cla32_fa724_and1;
  wire f_u_dadda_cla32_fa724_or0;
  wire f_u_dadda_cla32_fa725_xor0;
  wire f_u_dadda_cla32_fa725_and0;
  wire f_u_dadda_cla32_fa725_xor1;
  wire f_u_dadda_cla32_fa725_and1;
  wire f_u_dadda_cla32_fa725_or0;
  wire f_u_dadda_cla32_fa726_xor0;
  wire f_u_dadda_cla32_fa726_and0;
  wire f_u_dadda_cla32_fa726_xor1;
  wire f_u_dadda_cla32_fa726_and1;
  wire f_u_dadda_cla32_fa726_or0;
  wire f_u_dadda_cla32_fa727_xor0;
  wire f_u_dadda_cla32_fa727_and0;
  wire f_u_dadda_cla32_fa727_xor1;
  wire f_u_dadda_cla32_fa727_and1;
  wire f_u_dadda_cla32_fa727_or0;
  wire f_u_dadda_cla32_fa728_xor0;
  wire f_u_dadda_cla32_fa728_and0;
  wire f_u_dadda_cla32_fa728_xor1;
  wire f_u_dadda_cla32_fa728_and1;
  wire f_u_dadda_cla32_fa728_or0;
  wire f_u_dadda_cla32_fa729_xor0;
  wire f_u_dadda_cla32_fa729_and0;
  wire f_u_dadda_cla32_fa729_xor1;
  wire f_u_dadda_cla32_fa729_and1;
  wire f_u_dadda_cla32_fa729_or0;
  wire f_u_dadda_cla32_fa730_xor0;
  wire f_u_dadda_cla32_fa730_and0;
  wire f_u_dadda_cla32_fa730_xor1;
  wire f_u_dadda_cla32_fa730_and1;
  wire f_u_dadda_cla32_fa730_or0;
  wire f_u_dadda_cla32_fa731_xor0;
  wire f_u_dadda_cla32_fa731_and0;
  wire f_u_dadda_cla32_fa731_xor1;
  wire f_u_dadda_cla32_fa731_and1;
  wire f_u_dadda_cla32_fa731_or0;
  wire f_u_dadda_cla32_fa732_xor0;
  wire f_u_dadda_cla32_fa732_and0;
  wire f_u_dadda_cla32_fa732_xor1;
  wire f_u_dadda_cla32_fa732_and1;
  wire f_u_dadda_cla32_fa732_or0;
  wire f_u_dadda_cla32_fa733_xor0;
  wire f_u_dadda_cla32_fa733_and0;
  wire f_u_dadda_cla32_fa733_xor1;
  wire f_u_dadda_cla32_fa733_and1;
  wire f_u_dadda_cla32_fa733_or0;
  wire f_u_dadda_cla32_fa734_xor0;
  wire f_u_dadda_cla32_fa734_and0;
  wire f_u_dadda_cla32_fa734_xor1;
  wire f_u_dadda_cla32_fa734_and1;
  wire f_u_dadda_cla32_fa734_or0;
  wire f_u_dadda_cla32_fa735_xor0;
  wire f_u_dadda_cla32_fa735_and0;
  wire f_u_dadda_cla32_fa735_xor1;
  wire f_u_dadda_cla32_fa735_and1;
  wire f_u_dadda_cla32_fa735_or0;
  wire f_u_dadda_cla32_fa736_xor0;
  wire f_u_dadda_cla32_fa736_and0;
  wire f_u_dadda_cla32_fa736_xor1;
  wire f_u_dadda_cla32_fa736_and1;
  wire f_u_dadda_cla32_fa736_or0;
  wire f_u_dadda_cla32_fa737_xor0;
  wire f_u_dadda_cla32_fa737_and0;
  wire f_u_dadda_cla32_fa737_xor1;
  wire f_u_dadda_cla32_fa737_and1;
  wire f_u_dadda_cla32_fa737_or0;
  wire f_u_dadda_cla32_fa738_xor0;
  wire f_u_dadda_cla32_fa738_and0;
  wire f_u_dadda_cla32_fa738_xor1;
  wire f_u_dadda_cla32_fa738_and1;
  wire f_u_dadda_cla32_fa738_or0;
  wire f_u_dadda_cla32_fa739_xor0;
  wire f_u_dadda_cla32_fa739_and0;
  wire f_u_dadda_cla32_fa739_xor1;
  wire f_u_dadda_cla32_fa739_and1;
  wire f_u_dadda_cla32_fa739_or0;
  wire f_u_dadda_cla32_fa740_xor0;
  wire f_u_dadda_cla32_fa740_and0;
  wire f_u_dadda_cla32_fa740_xor1;
  wire f_u_dadda_cla32_fa740_and1;
  wire f_u_dadda_cla32_fa740_or0;
  wire f_u_dadda_cla32_fa741_xor0;
  wire f_u_dadda_cla32_fa741_and0;
  wire f_u_dadda_cla32_fa741_xor1;
  wire f_u_dadda_cla32_fa741_and1;
  wire f_u_dadda_cla32_fa741_or0;
  wire f_u_dadda_cla32_fa742_xor0;
  wire f_u_dadda_cla32_fa742_and0;
  wire f_u_dadda_cla32_fa742_xor1;
  wire f_u_dadda_cla32_fa742_and1;
  wire f_u_dadda_cla32_fa742_or0;
  wire f_u_dadda_cla32_fa743_xor0;
  wire f_u_dadda_cla32_fa743_and0;
  wire f_u_dadda_cla32_fa743_xor1;
  wire f_u_dadda_cla32_fa743_and1;
  wire f_u_dadda_cla32_fa743_or0;
  wire f_u_dadda_cla32_fa744_xor0;
  wire f_u_dadda_cla32_fa744_and0;
  wire f_u_dadda_cla32_fa744_xor1;
  wire f_u_dadda_cla32_fa744_and1;
  wire f_u_dadda_cla32_fa744_or0;
  wire f_u_dadda_cla32_fa745_xor0;
  wire f_u_dadda_cla32_fa745_and0;
  wire f_u_dadda_cla32_fa745_xor1;
  wire f_u_dadda_cla32_fa745_and1;
  wire f_u_dadda_cla32_fa745_or0;
  wire f_u_dadda_cla32_fa746_xor0;
  wire f_u_dadda_cla32_fa746_and0;
  wire f_u_dadda_cla32_fa746_xor1;
  wire f_u_dadda_cla32_fa746_and1;
  wire f_u_dadda_cla32_fa746_or0;
  wire f_u_dadda_cla32_fa747_xor0;
  wire f_u_dadda_cla32_fa747_and0;
  wire f_u_dadda_cla32_fa747_xor1;
  wire f_u_dadda_cla32_fa747_and1;
  wire f_u_dadda_cla32_fa747_or0;
  wire f_u_dadda_cla32_fa748_xor0;
  wire f_u_dadda_cla32_fa748_and0;
  wire f_u_dadda_cla32_fa748_xor1;
  wire f_u_dadda_cla32_fa748_and1;
  wire f_u_dadda_cla32_fa748_or0;
  wire f_u_dadda_cla32_fa749_xor0;
  wire f_u_dadda_cla32_fa749_and0;
  wire f_u_dadda_cla32_fa749_xor1;
  wire f_u_dadda_cla32_fa749_and1;
  wire f_u_dadda_cla32_fa749_or0;
  wire f_u_dadda_cla32_fa750_xor0;
  wire f_u_dadda_cla32_fa750_and0;
  wire f_u_dadda_cla32_fa750_xor1;
  wire f_u_dadda_cla32_fa750_and1;
  wire f_u_dadda_cla32_fa750_or0;
  wire f_u_dadda_cla32_fa751_xor0;
  wire f_u_dadda_cla32_fa751_and0;
  wire f_u_dadda_cla32_fa751_xor1;
  wire f_u_dadda_cla32_fa751_and1;
  wire f_u_dadda_cla32_fa751_or0;
  wire f_u_dadda_cla32_fa752_xor0;
  wire f_u_dadda_cla32_fa752_and0;
  wire f_u_dadda_cla32_fa752_xor1;
  wire f_u_dadda_cla32_fa752_and1;
  wire f_u_dadda_cla32_fa752_or0;
  wire f_u_dadda_cla32_fa753_xor0;
  wire f_u_dadda_cla32_fa753_and0;
  wire f_u_dadda_cla32_fa753_xor1;
  wire f_u_dadda_cla32_fa753_and1;
  wire f_u_dadda_cla32_fa753_or0;
  wire f_u_dadda_cla32_fa754_xor0;
  wire f_u_dadda_cla32_fa754_and0;
  wire f_u_dadda_cla32_fa754_xor1;
  wire f_u_dadda_cla32_fa754_and1;
  wire f_u_dadda_cla32_fa754_or0;
  wire f_u_dadda_cla32_fa755_xor0;
  wire f_u_dadda_cla32_fa755_and0;
  wire f_u_dadda_cla32_fa755_xor1;
  wire f_u_dadda_cla32_fa755_and1;
  wire f_u_dadda_cla32_fa755_or0;
  wire f_u_dadda_cla32_fa756_xor0;
  wire f_u_dadda_cla32_fa756_and0;
  wire f_u_dadda_cla32_fa756_xor1;
  wire f_u_dadda_cla32_fa756_and1;
  wire f_u_dadda_cla32_fa756_or0;
  wire f_u_dadda_cla32_fa757_xor0;
  wire f_u_dadda_cla32_fa757_and0;
  wire f_u_dadda_cla32_fa757_xor1;
  wire f_u_dadda_cla32_fa757_and1;
  wire f_u_dadda_cla32_fa757_or0;
  wire f_u_dadda_cla32_fa758_xor0;
  wire f_u_dadda_cla32_fa758_and0;
  wire f_u_dadda_cla32_fa758_xor1;
  wire f_u_dadda_cla32_fa758_and1;
  wire f_u_dadda_cla32_fa758_or0;
  wire f_u_dadda_cla32_fa759_xor0;
  wire f_u_dadda_cla32_fa759_and0;
  wire f_u_dadda_cla32_fa759_xor1;
  wire f_u_dadda_cla32_fa759_and1;
  wire f_u_dadda_cla32_fa759_or0;
  wire f_u_dadda_cla32_fa760_xor0;
  wire f_u_dadda_cla32_fa760_and0;
  wire f_u_dadda_cla32_fa760_xor1;
  wire f_u_dadda_cla32_fa760_and1;
  wire f_u_dadda_cla32_fa760_or0;
  wire f_u_dadda_cla32_fa761_xor0;
  wire f_u_dadda_cla32_fa761_and0;
  wire f_u_dadda_cla32_fa761_xor1;
  wire f_u_dadda_cla32_fa761_and1;
  wire f_u_dadda_cla32_fa761_or0;
  wire f_u_dadda_cla32_fa762_xor0;
  wire f_u_dadda_cla32_fa762_and0;
  wire f_u_dadda_cla32_fa762_xor1;
  wire f_u_dadda_cla32_fa762_and1;
  wire f_u_dadda_cla32_fa762_or0;
  wire f_u_dadda_cla32_fa763_xor0;
  wire f_u_dadda_cla32_fa763_and0;
  wire f_u_dadda_cla32_fa763_xor1;
  wire f_u_dadda_cla32_fa763_and1;
  wire f_u_dadda_cla32_fa763_or0;
  wire f_u_dadda_cla32_fa764_xor0;
  wire f_u_dadda_cla32_fa764_and0;
  wire f_u_dadda_cla32_fa764_xor1;
  wire f_u_dadda_cla32_fa764_and1;
  wire f_u_dadda_cla32_fa764_or0;
  wire f_u_dadda_cla32_fa765_xor0;
  wire f_u_dadda_cla32_fa765_and0;
  wire f_u_dadda_cla32_fa765_xor1;
  wire f_u_dadda_cla32_fa765_and1;
  wire f_u_dadda_cla32_fa765_or0;
  wire f_u_dadda_cla32_fa766_xor0;
  wire f_u_dadda_cla32_fa766_and0;
  wire f_u_dadda_cla32_fa766_xor1;
  wire f_u_dadda_cla32_fa766_and1;
  wire f_u_dadda_cla32_fa766_or0;
  wire f_u_dadda_cla32_fa767_xor0;
  wire f_u_dadda_cla32_fa767_and0;
  wire f_u_dadda_cla32_fa767_xor1;
  wire f_u_dadda_cla32_fa767_and1;
  wire f_u_dadda_cla32_fa767_or0;
  wire f_u_dadda_cla32_fa768_xor0;
  wire f_u_dadda_cla32_fa768_and0;
  wire f_u_dadda_cla32_fa768_xor1;
  wire f_u_dadda_cla32_fa768_and1;
  wire f_u_dadda_cla32_fa768_or0;
  wire f_u_dadda_cla32_fa769_xor0;
  wire f_u_dadda_cla32_fa769_and0;
  wire f_u_dadda_cla32_fa769_xor1;
  wire f_u_dadda_cla32_fa769_and1;
  wire f_u_dadda_cla32_fa769_or0;
  wire f_u_dadda_cla32_and_22_31;
  wire f_u_dadda_cla32_fa770_xor0;
  wire f_u_dadda_cla32_fa770_and0;
  wire f_u_dadda_cla32_fa770_xor1;
  wire f_u_dadda_cla32_fa770_and1;
  wire f_u_dadda_cla32_fa770_or0;
  wire f_u_dadda_cla32_fa771_xor0;
  wire f_u_dadda_cla32_fa771_and0;
  wire f_u_dadda_cla32_fa771_xor1;
  wire f_u_dadda_cla32_fa771_and1;
  wire f_u_dadda_cla32_fa771_or0;
  wire f_u_dadda_cla32_and_24_30;
  wire f_u_dadda_cla32_fa772_xor0;
  wire f_u_dadda_cla32_fa772_and0;
  wire f_u_dadda_cla32_fa772_xor1;
  wire f_u_dadda_cla32_fa772_and1;
  wire f_u_dadda_cla32_fa772_or0;
  wire f_u_dadda_cla32_and_23_31;
  wire f_u_dadda_cla32_fa773_xor0;
  wire f_u_dadda_cla32_fa773_and0;
  wire f_u_dadda_cla32_fa773_xor1;
  wire f_u_dadda_cla32_fa773_and1;
  wire f_u_dadda_cla32_fa773_or0;
  wire f_u_dadda_cla32_and_26_29;
  wire f_u_dadda_cla32_fa774_xor0;
  wire f_u_dadda_cla32_fa774_and0;
  wire f_u_dadda_cla32_fa774_xor1;
  wire f_u_dadda_cla32_fa774_and1;
  wire f_u_dadda_cla32_fa774_or0;
  wire f_u_dadda_cla32_and_25_30;
  wire f_u_dadda_cla32_and_24_31;
  wire f_u_dadda_cla32_fa775_xor0;
  wire f_u_dadda_cla32_fa775_and0;
  wire f_u_dadda_cla32_fa775_xor1;
  wire f_u_dadda_cla32_fa775_and1;
  wire f_u_dadda_cla32_fa775_or0;
  wire f_u_dadda_cla32_and_28_28;
  wire f_u_dadda_cla32_fa776_xor0;
  wire f_u_dadda_cla32_fa776_and0;
  wire f_u_dadda_cla32_fa776_xor1;
  wire f_u_dadda_cla32_fa776_and1;
  wire f_u_dadda_cla32_fa776_or0;
  wire f_u_dadda_cla32_and_27_29;
  wire f_u_dadda_cla32_and_26_30;
  wire f_u_dadda_cla32_and_25_31;
  wire f_u_dadda_cla32_fa777_xor0;
  wire f_u_dadda_cla32_fa777_and0;
  wire f_u_dadda_cla32_fa777_xor1;
  wire f_u_dadda_cla32_fa777_and1;
  wire f_u_dadda_cla32_fa777_or0;
  wire f_u_dadda_cla32_and_30_27;
  wire f_u_dadda_cla32_fa778_xor0;
  wire f_u_dadda_cla32_fa778_and0;
  wire f_u_dadda_cla32_fa778_xor1;
  wire f_u_dadda_cla32_fa778_and1;
  wire f_u_dadda_cla32_fa778_or0;
  wire f_u_dadda_cla32_and_29_28;
  wire f_u_dadda_cla32_and_28_29;
  wire f_u_dadda_cla32_and_27_30;
  wire f_u_dadda_cla32_fa779_xor0;
  wire f_u_dadda_cla32_fa779_and0;
  wire f_u_dadda_cla32_fa779_xor1;
  wire f_u_dadda_cla32_fa779_and1;
  wire f_u_dadda_cla32_fa779_or0;
  wire f_u_dadda_cla32_fa780_xor0;
  wire f_u_dadda_cla32_fa780_and0;
  wire f_u_dadda_cla32_fa780_xor1;
  wire f_u_dadda_cla32_fa780_and1;
  wire f_u_dadda_cla32_fa780_or0;
  wire f_u_dadda_cla32_and_31_27;
  wire f_u_dadda_cla32_and_30_28;
  wire f_u_dadda_cla32_and_29_29;
  wire f_u_dadda_cla32_fa781_xor0;
  wire f_u_dadda_cla32_fa781_and0;
  wire f_u_dadda_cla32_fa781_xor1;
  wire f_u_dadda_cla32_fa781_and1;
  wire f_u_dadda_cla32_fa781_or0;
  wire f_u_dadda_cla32_and_31_28;
  wire f_u_dadda_cla32_fa782_xor0;
  wire f_u_dadda_cla32_fa782_and0;
  wire f_u_dadda_cla32_fa782_xor1;
  wire f_u_dadda_cla32_fa782_and1;
  wire f_u_dadda_cla32_fa782_or0;
  wire f_u_dadda_cla32_and_3_0;
  wire f_u_dadda_cla32_and_2_1;
  wire f_u_dadda_cla32_ha29_xor0;
  wire f_u_dadda_cla32_ha29_and0;
  wire f_u_dadda_cla32_and_2_2;
  wire f_u_dadda_cla32_and_1_3;
  wire f_u_dadda_cla32_fa783_xor0;
  wire f_u_dadda_cla32_fa783_and0;
  wire f_u_dadda_cla32_fa783_xor1;
  wire f_u_dadda_cla32_fa783_and1;
  wire f_u_dadda_cla32_fa783_or0;
  wire f_u_dadda_cla32_and_1_4;
  wire f_u_dadda_cla32_and_0_5;
  wire f_u_dadda_cla32_fa784_xor0;
  wire f_u_dadda_cla32_fa784_and0;
  wire f_u_dadda_cla32_fa784_xor1;
  wire f_u_dadda_cla32_fa784_and1;
  wire f_u_dadda_cla32_fa784_or0;
  wire f_u_dadda_cla32_and_0_6;
  wire f_u_dadda_cla32_fa785_xor0;
  wire f_u_dadda_cla32_fa785_and0;
  wire f_u_dadda_cla32_fa785_xor1;
  wire f_u_dadda_cla32_fa785_and1;
  wire f_u_dadda_cla32_fa785_or0;
  wire f_u_dadda_cla32_fa786_xor0;
  wire f_u_dadda_cla32_fa786_and0;
  wire f_u_dadda_cla32_fa786_xor1;
  wire f_u_dadda_cla32_fa786_and1;
  wire f_u_dadda_cla32_fa786_or0;
  wire f_u_dadda_cla32_fa787_xor0;
  wire f_u_dadda_cla32_fa787_and0;
  wire f_u_dadda_cla32_fa787_xor1;
  wire f_u_dadda_cla32_fa787_and1;
  wire f_u_dadda_cla32_fa787_or0;
  wire f_u_dadda_cla32_fa788_xor0;
  wire f_u_dadda_cla32_fa788_and0;
  wire f_u_dadda_cla32_fa788_xor1;
  wire f_u_dadda_cla32_fa788_and1;
  wire f_u_dadda_cla32_fa788_or0;
  wire f_u_dadda_cla32_fa789_xor0;
  wire f_u_dadda_cla32_fa789_and0;
  wire f_u_dadda_cla32_fa789_xor1;
  wire f_u_dadda_cla32_fa789_and1;
  wire f_u_dadda_cla32_fa789_or0;
  wire f_u_dadda_cla32_fa790_xor0;
  wire f_u_dadda_cla32_fa790_and0;
  wire f_u_dadda_cla32_fa790_xor1;
  wire f_u_dadda_cla32_fa790_and1;
  wire f_u_dadda_cla32_fa790_or0;
  wire f_u_dadda_cla32_fa791_xor0;
  wire f_u_dadda_cla32_fa791_and0;
  wire f_u_dadda_cla32_fa791_xor1;
  wire f_u_dadda_cla32_fa791_and1;
  wire f_u_dadda_cla32_fa791_or0;
  wire f_u_dadda_cla32_fa792_xor0;
  wire f_u_dadda_cla32_fa792_and0;
  wire f_u_dadda_cla32_fa792_xor1;
  wire f_u_dadda_cla32_fa792_and1;
  wire f_u_dadda_cla32_fa792_or0;
  wire f_u_dadda_cla32_fa793_xor0;
  wire f_u_dadda_cla32_fa793_and0;
  wire f_u_dadda_cla32_fa793_xor1;
  wire f_u_dadda_cla32_fa793_and1;
  wire f_u_dadda_cla32_fa793_or0;
  wire f_u_dadda_cla32_fa794_xor0;
  wire f_u_dadda_cla32_fa794_and0;
  wire f_u_dadda_cla32_fa794_xor1;
  wire f_u_dadda_cla32_fa794_and1;
  wire f_u_dadda_cla32_fa794_or0;
  wire f_u_dadda_cla32_fa795_xor0;
  wire f_u_dadda_cla32_fa795_and0;
  wire f_u_dadda_cla32_fa795_xor1;
  wire f_u_dadda_cla32_fa795_and1;
  wire f_u_dadda_cla32_fa795_or0;
  wire f_u_dadda_cla32_fa796_xor0;
  wire f_u_dadda_cla32_fa796_and0;
  wire f_u_dadda_cla32_fa796_xor1;
  wire f_u_dadda_cla32_fa796_and1;
  wire f_u_dadda_cla32_fa796_or0;
  wire f_u_dadda_cla32_fa797_xor0;
  wire f_u_dadda_cla32_fa797_and0;
  wire f_u_dadda_cla32_fa797_xor1;
  wire f_u_dadda_cla32_fa797_and1;
  wire f_u_dadda_cla32_fa797_or0;
  wire f_u_dadda_cla32_fa798_xor0;
  wire f_u_dadda_cla32_fa798_and0;
  wire f_u_dadda_cla32_fa798_xor1;
  wire f_u_dadda_cla32_fa798_and1;
  wire f_u_dadda_cla32_fa798_or0;
  wire f_u_dadda_cla32_fa799_xor0;
  wire f_u_dadda_cla32_fa799_and0;
  wire f_u_dadda_cla32_fa799_xor1;
  wire f_u_dadda_cla32_fa799_and1;
  wire f_u_dadda_cla32_fa799_or0;
  wire f_u_dadda_cla32_fa800_xor0;
  wire f_u_dadda_cla32_fa800_and0;
  wire f_u_dadda_cla32_fa800_xor1;
  wire f_u_dadda_cla32_fa800_and1;
  wire f_u_dadda_cla32_fa800_or0;
  wire f_u_dadda_cla32_fa801_xor0;
  wire f_u_dadda_cla32_fa801_and0;
  wire f_u_dadda_cla32_fa801_xor1;
  wire f_u_dadda_cla32_fa801_and1;
  wire f_u_dadda_cla32_fa801_or0;
  wire f_u_dadda_cla32_fa802_xor0;
  wire f_u_dadda_cla32_fa802_and0;
  wire f_u_dadda_cla32_fa802_xor1;
  wire f_u_dadda_cla32_fa802_and1;
  wire f_u_dadda_cla32_fa802_or0;
  wire f_u_dadda_cla32_fa803_xor0;
  wire f_u_dadda_cla32_fa803_and0;
  wire f_u_dadda_cla32_fa803_xor1;
  wire f_u_dadda_cla32_fa803_and1;
  wire f_u_dadda_cla32_fa803_or0;
  wire f_u_dadda_cla32_fa804_xor0;
  wire f_u_dadda_cla32_fa804_and0;
  wire f_u_dadda_cla32_fa804_xor1;
  wire f_u_dadda_cla32_fa804_and1;
  wire f_u_dadda_cla32_fa804_or0;
  wire f_u_dadda_cla32_fa805_xor0;
  wire f_u_dadda_cla32_fa805_and0;
  wire f_u_dadda_cla32_fa805_xor1;
  wire f_u_dadda_cla32_fa805_and1;
  wire f_u_dadda_cla32_fa805_or0;
  wire f_u_dadda_cla32_fa806_xor0;
  wire f_u_dadda_cla32_fa806_and0;
  wire f_u_dadda_cla32_fa806_xor1;
  wire f_u_dadda_cla32_fa806_and1;
  wire f_u_dadda_cla32_fa806_or0;
  wire f_u_dadda_cla32_fa807_xor0;
  wire f_u_dadda_cla32_fa807_and0;
  wire f_u_dadda_cla32_fa807_xor1;
  wire f_u_dadda_cla32_fa807_and1;
  wire f_u_dadda_cla32_fa807_or0;
  wire f_u_dadda_cla32_fa808_xor0;
  wire f_u_dadda_cla32_fa808_and0;
  wire f_u_dadda_cla32_fa808_xor1;
  wire f_u_dadda_cla32_fa808_and1;
  wire f_u_dadda_cla32_fa808_or0;
  wire f_u_dadda_cla32_fa809_xor0;
  wire f_u_dadda_cla32_fa809_and0;
  wire f_u_dadda_cla32_fa809_xor1;
  wire f_u_dadda_cla32_fa809_and1;
  wire f_u_dadda_cla32_fa809_or0;
  wire f_u_dadda_cla32_fa810_xor0;
  wire f_u_dadda_cla32_fa810_and0;
  wire f_u_dadda_cla32_fa810_xor1;
  wire f_u_dadda_cla32_fa810_and1;
  wire f_u_dadda_cla32_fa810_or0;
  wire f_u_dadda_cla32_fa811_xor0;
  wire f_u_dadda_cla32_fa811_and0;
  wire f_u_dadda_cla32_fa811_xor1;
  wire f_u_dadda_cla32_fa811_and1;
  wire f_u_dadda_cla32_fa811_or0;
  wire f_u_dadda_cla32_fa812_xor0;
  wire f_u_dadda_cla32_fa812_and0;
  wire f_u_dadda_cla32_fa812_xor1;
  wire f_u_dadda_cla32_fa812_and1;
  wire f_u_dadda_cla32_fa812_or0;
  wire f_u_dadda_cla32_fa813_xor0;
  wire f_u_dadda_cla32_fa813_and0;
  wire f_u_dadda_cla32_fa813_xor1;
  wire f_u_dadda_cla32_fa813_and1;
  wire f_u_dadda_cla32_fa813_or0;
  wire f_u_dadda_cla32_fa814_xor0;
  wire f_u_dadda_cla32_fa814_and0;
  wire f_u_dadda_cla32_fa814_xor1;
  wire f_u_dadda_cla32_fa814_and1;
  wire f_u_dadda_cla32_fa814_or0;
  wire f_u_dadda_cla32_fa815_xor0;
  wire f_u_dadda_cla32_fa815_and0;
  wire f_u_dadda_cla32_fa815_xor1;
  wire f_u_dadda_cla32_fa815_and1;
  wire f_u_dadda_cla32_fa815_or0;
  wire f_u_dadda_cla32_fa816_xor0;
  wire f_u_dadda_cla32_fa816_and0;
  wire f_u_dadda_cla32_fa816_xor1;
  wire f_u_dadda_cla32_fa816_and1;
  wire f_u_dadda_cla32_fa816_or0;
  wire f_u_dadda_cla32_fa817_xor0;
  wire f_u_dadda_cla32_fa817_and0;
  wire f_u_dadda_cla32_fa817_xor1;
  wire f_u_dadda_cla32_fa817_and1;
  wire f_u_dadda_cla32_fa817_or0;
  wire f_u_dadda_cla32_fa818_xor0;
  wire f_u_dadda_cla32_fa818_and0;
  wire f_u_dadda_cla32_fa818_xor1;
  wire f_u_dadda_cla32_fa818_and1;
  wire f_u_dadda_cla32_fa818_or0;
  wire f_u_dadda_cla32_fa819_xor0;
  wire f_u_dadda_cla32_fa819_and0;
  wire f_u_dadda_cla32_fa819_xor1;
  wire f_u_dadda_cla32_fa819_and1;
  wire f_u_dadda_cla32_fa819_or0;
  wire f_u_dadda_cla32_fa820_xor0;
  wire f_u_dadda_cla32_fa820_and0;
  wire f_u_dadda_cla32_fa820_xor1;
  wire f_u_dadda_cla32_fa820_and1;
  wire f_u_dadda_cla32_fa820_or0;
  wire f_u_dadda_cla32_fa821_xor0;
  wire f_u_dadda_cla32_fa821_and0;
  wire f_u_dadda_cla32_fa821_xor1;
  wire f_u_dadda_cla32_fa821_and1;
  wire f_u_dadda_cla32_fa821_or0;
  wire f_u_dadda_cla32_fa822_xor0;
  wire f_u_dadda_cla32_fa822_and0;
  wire f_u_dadda_cla32_fa822_xor1;
  wire f_u_dadda_cla32_fa822_and1;
  wire f_u_dadda_cla32_fa822_or0;
  wire f_u_dadda_cla32_fa823_xor0;
  wire f_u_dadda_cla32_fa823_and0;
  wire f_u_dadda_cla32_fa823_xor1;
  wire f_u_dadda_cla32_fa823_and1;
  wire f_u_dadda_cla32_fa823_or0;
  wire f_u_dadda_cla32_fa824_xor0;
  wire f_u_dadda_cla32_fa824_and0;
  wire f_u_dadda_cla32_fa824_xor1;
  wire f_u_dadda_cla32_fa824_and1;
  wire f_u_dadda_cla32_fa824_or0;
  wire f_u_dadda_cla32_fa825_xor0;
  wire f_u_dadda_cla32_fa825_and0;
  wire f_u_dadda_cla32_fa825_xor1;
  wire f_u_dadda_cla32_fa825_and1;
  wire f_u_dadda_cla32_fa825_or0;
  wire f_u_dadda_cla32_fa826_xor0;
  wire f_u_dadda_cla32_fa826_and0;
  wire f_u_dadda_cla32_fa826_xor1;
  wire f_u_dadda_cla32_fa826_and1;
  wire f_u_dadda_cla32_fa826_or0;
  wire f_u_dadda_cla32_fa827_xor0;
  wire f_u_dadda_cla32_fa827_and0;
  wire f_u_dadda_cla32_fa827_xor1;
  wire f_u_dadda_cla32_fa827_and1;
  wire f_u_dadda_cla32_fa827_or0;
  wire f_u_dadda_cla32_fa828_xor0;
  wire f_u_dadda_cla32_fa828_and0;
  wire f_u_dadda_cla32_fa828_xor1;
  wire f_u_dadda_cla32_fa828_and1;
  wire f_u_dadda_cla32_fa828_or0;
  wire f_u_dadda_cla32_fa829_xor0;
  wire f_u_dadda_cla32_fa829_and0;
  wire f_u_dadda_cla32_fa829_xor1;
  wire f_u_dadda_cla32_fa829_and1;
  wire f_u_dadda_cla32_fa829_or0;
  wire f_u_dadda_cla32_fa830_xor0;
  wire f_u_dadda_cla32_fa830_and0;
  wire f_u_dadda_cla32_fa830_xor1;
  wire f_u_dadda_cla32_fa830_and1;
  wire f_u_dadda_cla32_fa830_or0;
  wire f_u_dadda_cla32_fa831_xor0;
  wire f_u_dadda_cla32_fa831_and0;
  wire f_u_dadda_cla32_fa831_xor1;
  wire f_u_dadda_cla32_fa831_and1;
  wire f_u_dadda_cla32_fa831_or0;
  wire f_u_dadda_cla32_fa832_xor0;
  wire f_u_dadda_cla32_fa832_and0;
  wire f_u_dadda_cla32_fa832_xor1;
  wire f_u_dadda_cla32_fa832_and1;
  wire f_u_dadda_cla32_fa832_or0;
  wire f_u_dadda_cla32_fa833_xor0;
  wire f_u_dadda_cla32_fa833_and0;
  wire f_u_dadda_cla32_fa833_xor1;
  wire f_u_dadda_cla32_fa833_and1;
  wire f_u_dadda_cla32_fa833_or0;
  wire f_u_dadda_cla32_fa834_xor0;
  wire f_u_dadda_cla32_fa834_and0;
  wire f_u_dadda_cla32_fa834_xor1;
  wire f_u_dadda_cla32_fa834_and1;
  wire f_u_dadda_cla32_fa834_or0;
  wire f_u_dadda_cla32_fa835_xor0;
  wire f_u_dadda_cla32_fa835_and0;
  wire f_u_dadda_cla32_fa835_xor1;
  wire f_u_dadda_cla32_fa835_and1;
  wire f_u_dadda_cla32_fa835_or0;
  wire f_u_dadda_cla32_and_26_31;
  wire f_u_dadda_cla32_fa836_xor0;
  wire f_u_dadda_cla32_fa836_and0;
  wire f_u_dadda_cla32_fa836_xor1;
  wire f_u_dadda_cla32_fa836_and1;
  wire f_u_dadda_cla32_fa836_or0;
  wire f_u_dadda_cla32_and_28_30;
  wire f_u_dadda_cla32_and_27_31;
  wire f_u_dadda_cla32_fa837_xor0;
  wire f_u_dadda_cla32_fa837_and0;
  wire f_u_dadda_cla32_fa837_xor1;
  wire f_u_dadda_cla32_fa837_and1;
  wire f_u_dadda_cla32_fa837_or0;
  wire f_u_dadda_cla32_and_30_29;
  wire f_u_dadda_cla32_and_29_30;
  wire f_u_dadda_cla32_fa838_xor0;
  wire f_u_dadda_cla32_fa838_and0;
  wire f_u_dadda_cla32_fa838_xor1;
  wire f_u_dadda_cla32_fa838_and1;
  wire f_u_dadda_cla32_fa838_or0;
  wire f_u_dadda_cla32_and_31_29;
  wire f_u_dadda_cla32_fa839_xor0;
  wire f_u_dadda_cla32_fa839_and0;
  wire f_u_dadda_cla32_fa839_xor1;
  wire f_u_dadda_cla32_fa839_and1;
  wire f_u_dadda_cla32_fa839_or0;
  wire f_u_dadda_cla32_and_2_0;
  wire f_u_dadda_cla32_and_1_1;
  wire f_u_dadda_cla32_ha30_xor0;
  wire f_u_dadda_cla32_ha30_and0;
  wire f_u_dadda_cla32_and_1_2;
  wire f_u_dadda_cla32_and_0_3;
  wire f_u_dadda_cla32_fa840_xor0;
  wire f_u_dadda_cla32_fa840_and0;
  wire f_u_dadda_cla32_fa840_xor1;
  wire f_u_dadda_cla32_fa840_and1;
  wire f_u_dadda_cla32_fa840_or0;
  wire f_u_dadda_cla32_and_0_4;
  wire f_u_dadda_cla32_fa841_xor0;
  wire f_u_dadda_cla32_fa841_and0;
  wire f_u_dadda_cla32_fa841_xor1;
  wire f_u_dadda_cla32_fa841_and1;
  wire f_u_dadda_cla32_fa841_or0;
  wire f_u_dadda_cla32_fa842_xor0;
  wire f_u_dadda_cla32_fa842_and0;
  wire f_u_dadda_cla32_fa842_xor1;
  wire f_u_dadda_cla32_fa842_and1;
  wire f_u_dadda_cla32_fa842_or0;
  wire f_u_dadda_cla32_fa843_xor0;
  wire f_u_dadda_cla32_fa843_and0;
  wire f_u_dadda_cla32_fa843_xor1;
  wire f_u_dadda_cla32_fa843_and1;
  wire f_u_dadda_cla32_fa843_or0;
  wire f_u_dadda_cla32_fa844_xor0;
  wire f_u_dadda_cla32_fa844_and0;
  wire f_u_dadda_cla32_fa844_xor1;
  wire f_u_dadda_cla32_fa844_and1;
  wire f_u_dadda_cla32_fa844_or0;
  wire f_u_dadda_cla32_fa845_xor0;
  wire f_u_dadda_cla32_fa845_and0;
  wire f_u_dadda_cla32_fa845_xor1;
  wire f_u_dadda_cla32_fa845_and1;
  wire f_u_dadda_cla32_fa845_or0;
  wire f_u_dadda_cla32_fa846_xor0;
  wire f_u_dadda_cla32_fa846_and0;
  wire f_u_dadda_cla32_fa846_xor1;
  wire f_u_dadda_cla32_fa846_and1;
  wire f_u_dadda_cla32_fa846_or0;
  wire f_u_dadda_cla32_fa847_xor0;
  wire f_u_dadda_cla32_fa847_and0;
  wire f_u_dadda_cla32_fa847_xor1;
  wire f_u_dadda_cla32_fa847_and1;
  wire f_u_dadda_cla32_fa847_or0;
  wire f_u_dadda_cla32_fa848_xor0;
  wire f_u_dadda_cla32_fa848_and0;
  wire f_u_dadda_cla32_fa848_xor1;
  wire f_u_dadda_cla32_fa848_and1;
  wire f_u_dadda_cla32_fa848_or0;
  wire f_u_dadda_cla32_fa849_xor0;
  wire f_u_dadda_cla32_fa849_and0;
  wire f_u_dadda_cla32_fa849_xor1;
  wire f_u_dadda_cla32_fa849_and1;
  wire f_u_dadda_cla32_fa849_or0;
  wire f_u_dadda_cla32_fa850_xor0;
  wire f_u_dadda_cla32_fa850_and0;
  wire f_u_dadda_cla32_fa850_xor1;
  wire f_u_dadda_cla32_fa850_and1;
  wire f_u_dadda_cla32_fa850_or0;
  wire f_u_dadda_cla32_fa851_xor0;
  wire f_u_dadda_cla32_fa851_and0;
  wire f_u_dadda_cla32_fa851_xor1;
  wire f_u_dadda_cla32_fa851_and1;
  wire f_u_dadda_cla32_fa851_or0;
  wire f_u_dadda_cla32_fa852_xor0;
  wire f_u_dadda_cla32_fa852_and0;
  wire f_u_dadda_cla32_fa852_xor1;
  wire f_u_dadda_cla32_fa852_and1;
  wire f_u_dadda_cla32_fa852_or0;
  wire f_u_dadda_cla32_fa853_xor0;
  wire f_u_dadda_cla32_fa853_and0;
  wire f_u_dadda_cla32_fa853_xor1;
  wire f_u_dadda_cla32_fa853_and1;
  wire f_u_dadda_cla32_fa853_or0;
  wire f_u_dadda_cla32_fa854_xor0;
  wire f_u_dadda_cla32_fa854_and0;
  wire f_u_dadda_cla32_fa854_xor1;
  wire f_u_dadda_cla32_fa854_and1;
  wire f_u_dadda_cla32_fa854_or0;
  wire f_u_dadda_cla32_fa855_xor0;
  wire f_u_dadda_cla32_fa855_and0;
  wire f_u_dadda_cla32_fa855_xor1;
  wire f_u_dadda_cla32_fa855_and1;
  wire f_u_dadda_cla32_fa855_or0;
  wire f_u_dadda_cla32_fa856_xor0;
  wire f_u_dadda_cla32_fa856_and0;
  wire f_u_dadda_cla32_fa856_xor1;
  wire f_u_dadda_cla32_fa856_and1;
  wire f_u_dadda_cla32_fa856_or0;
  wire f_u_dadda_cla32_fa857_xor0;
  wire f_u_dadda_cla32_fa857_and0;
  wire f_u_dadda_cla32_fa857_xor1;
  wire f_u_dadda_cla32_fa857_and1;
  wire f_u_dadda_cla32_fa857_or0;
  wire f_u_dadda_cla32_fa858_xor0;
  wire f_u_dadda_cla32_fa858_and0;
  wire f_u_dadda_cla32_fa858_xor1;
  wire f_u_dadda_cla32_fa858_and1;
  wire f_u_dadda_cla32_fa858_or0;
  wire f_u_dadda_cla32_fa859_xor0;
  wire f_u_dadda_cla32_fa859_and0;
  wire f_u_dadda_cla32_fa859_xor1;
  wire f_u_dadda_cla32_fa859_and1;
  wire f_u_dadda_cla32_fa859_or0;
  wire f_u_dadda_cla32_fa860_xor0;
  wire f_u_dadda_cla32_fa860_and0;
  wire f_u_dadda_cla32_fa860_xor1;
  wire f_u_dadda_cla32_fa860_and1;
  wire f_u_dadda_cla32_fa860_or0;
  wire f_u_dadda_cla32_fa861_xor0;
  wire f_u_dadda_cla32_fa861_and0;
  wire f_u_dadda_cla32_fa861_xor1;
  wire f_u_dadda_cla32_fa861_and1;
  wire f_u_dadda_cla32_fa861_or0;
  wire f_u_dadda_cla32_fa862_xor0;
  wire f_u_dadda_cla32_fa862_and0;
  wire f_u_dadda_cla32_fa862_xor1;
  wire f_u_dadda_cla32_fa862_and1;
  wire f_u_dadda_cla32_fa862_or0;
  wire f_u_dadda_cla32_fa863_xor0;
  wire f_u_dadda_cla32_fa863_and0;
  wire f_u_dadda_cla32_fa863_xor1;
  wire f_u_dadda_cla32_fa863_and1;
  wire f_u_dadda_cla32_fa863_or0;
  wire f_u_dadda_cla32_fa864_xor0;
  wire f_u_dadda_cla32_fa864_and0;
  wire f_u_dadda_cla32_fa864_xor1;
  wire f_u_dadda_cla32_fa864_and1;
  wire f_u_dadda_cla32_fa864_or0;
  wire f_u_dadda_cla32_fa865_xor0;
  wire f_u_dadda_cla32_fa865_and0;
  wire f_u_dadda_cla32_fa865_xor1;
  wire f_u_dadda_cla32_fa865_and1;
  wire f_u_dadda_cla32_fa865_or0;
  wire f_u_dadda_cla32_fa866_xor0;
  wire f_u_dadda_cla32_fa866_and0;
  wire f_u_dadda_cla32_fa866_xor1;
  wire f_u_dadda_cla32_fa866_and1;
  wire f_u_dadda_cla32_fa866_or0;
  wire f_u_dadda_cla32_fa867_xor0;
  wire f_u_dadda_cla32_fa867_and0;
  wire f_u_dadda_cla32_fa867_xor1;
  wire f_u_dadda_cla32_fa867_and1;
  wire f_u_dadda_cla32_fa867_or0;
  wire f_u_dadda_cla32_fa868_xor0;
  wire f_u_dadda_cla32_fa868_and0;
  wire f_u_dadda_cla32_fa868_xor1;
  wire f_u_dadda_cla32_fa868_and1;
  wire f_u_dadda_cla32_fa868_or0;
  wire f_u_dadda_cla32_fa869_xor0;
  wire f_u_dadda_cla32_fa869_and0;
  wire f_u_dadda_cla32_fa869_xor1;
  wire f_u_dadda_cla32_fa869_and1;
  wire f_u_dadda_cla32_fa869_or0;
  wire f_u_dadda_cla32_fa870_xor0;
  wire f_u_dadda_cla32_fa870_and0;
  wire f_u_dadda_cla32_fa870_xor1;
  wire f_u_dadda_cla32_fa870_and1;
  wire f_u_dadda_cla32_fa870_or0;
  wire f_u_dadda_cla32_fa871_xor0;
  wire f_u_dadda_cla32_fa871_and0;
  wire f_u_dadda_cla32_fa871_xor1;
  wire f_u_dadda_cla32_fa871_and1;
  wire f_u_dadda_cla32_fa871_or0;
  wire f_u_dadda_cla32_fa872_xor0;
  wire f_u_dadda_cla32_fa872_and0;
  wire f_u_dadda_cla32_fa872_xor1;
  wire f_u_dadda_cla32_fa872_and1;
  wire f_u_dadda_cla32_fa872_or0;
  wire f_u_dadda_cla32_fa873_xor0;
  wire f_u_dadda_cla32_fa873_and0;
  wire f_u_dadda_cla32_fa873_xor1;
  wire f_u_dadda_cla32_fa873_and1;
  wire f_u_dadda_cla32_fa873_or0;
  wire f_u_dadda_cla32_fa874_xor0;
  wire f_u_dadda_cla32_fa874_and0;
  wire f_u_dadda_cla32_fa874_xor1;
  wire f_u_dadda_cla32_fa874_and1;
  wire f_u_dadda_cla32_fa874_or0;
  wire f_u_dadda_cla32_fa875_xor0;
  wire f_u_dadda_cla32_fa875_and0;
  wire f_u_dadda_cla32_fa875_xor1;
  wire f_u_dadda_cla32_fa875_and1;
  wire f_u_dadda_cla32_fa875_or0;
  wire f_u_dadda_cla32_fa876_xor0;
  wire f_u_dadda_cla32_fa876_and0;
  wire f_u_dadda_cla32_fa876_xor1;
  wire f_u_dadda_cla32_fa876_and1;
  wire f_u_dadda_cla32_fa876_or0;
  wire f_u_dadda_cla32_fa877_xor0;
  wire f_u_dadda_cla32_fa877_and0;
  wire f_u_dadda_cla32_fa877_xor1;
  wire f_u_dadda_cla32_fa877_and1;
  wire f_u_dadda_cla32_fa877_or0;
  wire f_u_dadda_cla32_fa878_xor0;
  wire f_u_dadda_cla32_fa878_and0;
  wire f_u_dadda_cla32_fa878_xor1;
  wire f_u_dadda_cla32_fa878_and1;
  wire f_u_dadda_cla32_fa878_or0;
  wire f_u_dadda_cla32_fa879_xor0;
  wire f_u_dadda_cla32_fa879_and0;
  wire f_u_dadda_cla32_fa879_xor1;
  wire f_u_dadda_cla32_fa879_and1;
  wire f_u_dadda_cla32_fa879_or0;
  wire f_u_dadda_cla32_fa880_xor0;
  wire f_u_dadda_cla32_fa880_and0;
  wire f_u_dadda_cla32_fa880_xor1;
  wire f_u_dadda_cla32_fa880_and1;
  wire f_u_dadda_cla32_fa880_or0;
  wire f_u_dadda_cla32_fa881_xor0;
  wire f_u_dadda_cla32_fa881_and0;
  wire f_u_dadda_cla32_fa881_xor1;
  wire f_u_dadda_cla32_fa881_and1;
  wire f_u_dadda_cla32_fa881_or0;
  wire f_u_dadda_cla32_fa882_xor0;
  wire f_u_dadda_cla32_fa882_and0;
  wire f_u_dadda_cla32_fa882_xor1;
  wire f_u_dadda_cla32_fa882_and1;
  wire f_u_dadda_cla32_fa882_or0;
  wire f_u_dadda_cla32_fa883_xor0;
  wire f_u_dadda_cla32_fa883_and0;
  wire f_u_dadda_cla32_fa883_xor1;
  wire f_u_dadda_cla32_fa883_and1;
  wire f_u_dadda_cla32_fa883_or0;
  wire f_u_dadda_cla32_fa884_xor0;
  wire f_u_dadda_cla32_fa884_and0;
  wire f_u_dadda_cla32_fa884_xor1;
  wire f_u_dadda_cla32_fa884_and1;
  wire f_u_dadda_cla32_fa884_or0;
  wire f_u_dadda_cla32_fa885_xor0;
  wire f_u_dadda_cla32_fa885_and0;
  wire f_u_dadda_cla32_fa885_xor1;
  wire f_u_dadda_cla32_fa885_and1;
  wire f_u_dadda_cla32_fa885_or0;
  wire f_u_dadda_cla32_fa886_xor0;
  wire f_u_dadda_cla32_fa886_and0;
  wire f_u_dadda_cla32_fa886_xor1;
  wire f_u_dadda_cla32_fa886_and1;
  wire f_u_dadda_cla32_fa886_or0;
  wire f_u_dadda_cla32_fa887_xor0;
  wire f_u_dadda_cla32_fa887_and0;
  wire f_u_dadda_cla32_fa887_xor1;
  wire f_u_dadda_cla32_fa887_and1;
  wire f_u_dadda_cla32_fa887_or0;
  wire f_u_dadda_cla32_fa888_xor0;
  wire f_u_dadda_cla32_fa888_and0;
  wire f_u_dadda_cla32_fa888_xor1;
  wire f_u_dadda_cla32_fa888_and1;
  wire f_u_dadda_cla32_fa888_or0;
  wire f_u_dadda_cla32_fa889_xor0;
  wire f_u_dadda_cla32_fa889_and0;
  wire f_u_dadda_cla32_fa889_xor1;
  wire f_u_dadda_cla32_fa889_and1;
  wire f_u_dadda_cla32_fa889_or0;
  wire f_u_dadda_cla32_fa890_xor0;
  wire f_u_dadda_cla32_fa890_and0;
  wire f_u_dadda_cla32_fa890_xor1;
  wire f_u_dadda_cla32_fa890_and1;
  wire f_u_dadda_cla32_fa890_or0;
  wire f_u_dadda_cla32_fa891_xor0;
  wire f_u_dadda_cla32_fa891_and0;
  wire f_u_dadda_cla32_fa891_xor1;
  wire f_u_dadda_cla32_fa891_and1;
  wire f_u_dadda_cla32_fa891_or0;
  wire f_u_dadda_cla32_fa892_xor0;
  wire f_u_dadda_cla32_fa892_and0;
  wire f_u_dadda_cla32_fa892_xor1;
  wire f_u_dadda_cla32_fa892_and1;
  wire f_u_dadda_cla32_fa892_or0;
  wire f_u_dadda_cla32_fa893_xor0;
  wire f_u_dadda_cla32_fa893_and0;
  wire f_u_dadda_cla32_fa893_xor1;
  wire f_u_dadda_cla32_fa893_and1;
  wire f_u_dadda_cla32_fa893_or0;
  wire f_u_dadda_cla32_fa894_xor0;
  wire f_u_dadda_cla32_fa894_and0;
  wire f_u_dadda_cla32_fa894_xor1;
  wire f_u_dadda_cla32_fa894_and1;
  wire f_u_dadda_cla32_fa894_or0;
  wire f_u_dadda_cla32_fa895_xor0;
  wire f_u_dadda_cla32_fa895_and0;
  wire f_u_dadda_cla32_fa895_xor1;
  wire f_u_dadda_cla32_fa895_and1;
  wire f_u_dadda_cla32_fa895_or0;
  wire f_u_dadda_cla32_and_28_31;
  wire f_u_dadda_cla32_fa896_xor0;
  wire f_u_dadda_cla32_fa896_and0;
  wire f_u_dadda_cla32_fa896_xor1;
  wire f_u_dadda_cla32_fa896_and1;
  wire f_u_dadda_cla32_fa896_or0;
  wire f_u_dadda_cla32_and_30_30;
  wire f_u_dadda_cla32_and_29_31;
  wire f_u_dadda_cla32_fa897_xor0;
  wire f_u_dadda_cla32_fa897_and0;
  wire f_u_dadda_cla32_fa897_xor1;
  wire f_u_dadda_cla32_fa897_and1;
  wire f_u_dadda_cla32_fa897_or0;
  wire f_u_dadda_cla32_and_31_30;
  wire f_u_dadda_cla32_fa898_xor0;
  wire f_u_dadda_cla32_fa898_and0;
  wire f_u_dadda_cla32_fa898_xor1;
  wire f_u_dadda_cla32_fa898_and1;
  wire f_u_dadda_cla32_fa898_or0;
  wire f_u_dadda_cla32_and_0_0;
  wire f_u_dadda_cla32_and_1_0;
  wire f_u_dadda_cla32_and_0_2;
  wire f_u_dadda_cla32_and_30_31;
  wire f_u_dadda_cla32_and_0_1;
  wire f_u_dadda_cla32_and_31_31;
  wire f_u_dadda_cla32_u_cla62_pg_logic0_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic0_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic0_xor0;
  wire f_u_dadda_cla32_u_cla62_pg_logic1_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic1_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic1_xor0;
  wire f_u_dadda_cla32_u_cla62_xor1;
  wire f_u_dadda_cla32_u_cla62_and0;
  wire f_u_dadda_cla32_u_cla62_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic2_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic2_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic2_xor0;
  wire f_u_dadda_cla32_u_cla62_xor2;
  wire f_u_dadda_cla32_u_cla62_and1;
  wire f_u_dadda_cla32_u_cla62_and2;
  wire f_u_dadda_cla32_u_cla62_and3;
  wire f_u_dadda_cla32_u_cla62_and4;
  wire f_u_dadda_cla32_u_cla62_or1;
  wire f_u_dadda_cla32_u_cla62_or2;
  wire f_u_dadda_cla32_u_cla62_pg_logic3_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic3_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic3_xor0;
  wire f_u_dadda_cla32_u_cla62_xor3;
  wire f_u_dadda_cla32_u_cla62_and5;
  wire f_u_dadda_cla32_u_cla62_and6;
  wire f_u_dadda_cla32_u_cla62_and7;
  wire f_u_dadda_cla32_u_cla62_and8;
  wire f_u_dadda_cla32_u_cla62_and9;
  wire f_u_dadda_cla32_u_cla62_and10;
  wire f_u_dadda_cla32_u_cla62_and11;
  wire f_u_dadda_cla32_u_cla62_or3;
  wire f_u_dadda_cla32_u_cla62_or4;
  wire f_u_dadda_cla32_u_cla62_or5;
  wire f_u_dadda_cla32_u_cla62_pg_logic4_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic4_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic4_xor0;
  wire f_u_dadda_cla32_u_cla62_xor4;
  wire f_u_dadda_cla32_u_cla62_and12;
  wire f_u_dadda_cla32_u_cla62_or6;
  wire f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic5_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic5_xor0;
  wire f_u_dadda_cla32_u_cla62_xor5;
  wire f_u_dadda_cla32_u_cla62_and13;
  wire f_u_dadda_cla32_u_cla62_and14;
  wire f_u_dadda_cla32_u_cla62_and15;
  wire f_u_dadda_cla32_u_cla62_or7;
  wire f_u_dadda_cla32_u_cla62_or8;
  wire f_u_dadda_cla32_u_cla62_pg_logic6_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic6_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic6_xor0;
  wire f_u_dadda_cla32_u_cla62_xor6;
  wire f_u_dadda_cla32_u_cla62_and16;
  wire f_u_dadda_cla32_u_cla62_and17;
  wire f_u_dadda_cla32_u_cla62_and18;
  wire f_u_dadda_cla32_u_cla62_and19;
  wire f_u_dadda_cla32_u_cla62_and20;
  wire f_u_dadda_cla32_u_cla62_and21;
  wire f_u_dadda_cla32_u_cla62_or9;
  wire f_u_dadda_cla32_u_cla62_or10;
  wire f_u_dadda_cla32_u_cla62_or11;
  wire f_u_dadda_cla32_u_cla62_pg_logic7_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic7_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic7_xor0;
  wire f_u_dadda_cla32_u_cla62_xor7;
  wire f_u_dadda_cla32_u_cla62_and22;
  wire f_u_dadda_cla32_u_cla62_and23;
  wire f_u_dadda_cla32_u_cla62_and24;
  wire f_u_dadda_cla32_u_cla62_and25;
  wire f_u_dadda_cla32_u_cla62_and26;
  wire f_u_dadda_cla32_u_cla62_and27;
  wire f_u_dadda_cla32_u_cla62_and28;
  wire f_u_dadda_cla32_u_cla62_and29;
  wire f_u_dadda_cla32_u_cla62_and30;
  wire f_u_dadda_cla32_u_cla62_and31;
  wire f_u_dadda_cla32_u_cla62_or12;
  wire f_u_dadda_cla32_u_cla62_or13;
  wire f_u_dadda_cla32_u_cla62_or14;
  wire f_u_dadda_cla32_u_cla62_or15;
  wire f_u_dadda_cla32_u_cla62_pg_logic8_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic8_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic8_xor0;
  wire f_u_dadda_cla32_u_cla62_xor8;
  wire f_u_dadda_cla32_u_cla62_and32;
  wire f_u_dadda_cla32_u_cla62_or16;
  wire f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic9_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic9_xor0;
  wire f_u_dadda_cla32_u_cla62_xor9;
  wire f_u_dadda_cla32_u_cla62_and33;
  wire f_u_dadda_cla32_u_cla62_and34;
  wire f_u_dadda_cla32_u_cla62_and35;
  wire f_u_dadda_cla32_u_cla62_or17;
  wire f_u_dadda_cla32_u_cla62_or18;
  wire f_u_dadda_cla32_u_cla62_pg_logic10_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic10_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic10_xor0;
  wire f_u_dadda_cla32_u_cla62_xor10;
  wire f_u_dadda_cla32_u_cla62_and36;
  wire f_u_dadda_cla32_u_cla62_and37;
  wire f_u_dadda_cla32_u_cla62_and38;
  wire f_u_dadda_cla32_u_cla62_and39;
  wire f_u_dadda_cla32_u_cla62_and40;
  wire f_u_dadda_cla32_u_cla62_and41;
  wire f_u_dadda_cla32_u_cla62_or19;
  wire f_u_dadda_cla32_u_cla62_or20;
  wire f_u_dadda_cla32_u_cla62_or21;
  wire f_u_dadda_cla32_u_cla62_pg_logic11_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic11_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic11_xor0;
  wire f_u_dadda_cla32_u_cla62_xor11;
  wire f_u_dadda_cla32_u_cla62_and42;
  wire f_u_dadda_cla32_u_cla62_and43;
  wire f_u_dadda_cla32_u_cla62_and44;
  wire f_u_dadda_cla32_u_cla62_and45;
  wire f_u_dadda_cla32_u_cla62_and46;
  wire f_u_dadda_cla32_u_cla62_and47;
  wire f_u_dadda_cla32_u_cla62_and48;
  wire f_u_dadda_cla32_u_cla62_and49;
  wire f_u_dadda_cla32_u_cla62_and50;
  wire f_u_dadda_cla32_u_cla62_and51;
  wire f_u_dadda_cla32_u_cla62_or22;
  wire f_u_dadda_cla32_u_cla62_or23;
  wire f_u_dadda_cla32_u_cla62_or24;
  wire f_u_dadda_cla32_u_cla62_or25;
  wire f_u_dadda_cla32_u_cla62_pg_logic12_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic12_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic12_xor0;
  wire f_u_dadda_cla32_u_cla62_xor12;
  wire f_u_dadda_cla32_u_cla62_and52;
  wire f_u_dadda_cla32_u_cla62_or26;
  wire f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic13_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic13_xor0;
  wire f_u_dadda_cla32_u_cla62_xor13;
  wire f_u_dadda_cla32_u_cla62_and53;
  wire f_u_dadda_cla32_u_cla62_and54;
  wire f_u_dadda_cla32_u_cla62_and55;
  wire f_u_dadda_cla32_u_cla62_or27;
  wire f_u_dadda_cla32_u_cla62_or28;
  wire f_u_dadda_cla32_u_cla62_pg_logic14_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic14_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic14_xor0;
  wire f_u_dadda_cla32_u_cla62_xor14;
  wire f_u_dadda_cla32_u_cla62_and56;
  wire f_u_dadda_cla32_u_cla62_and57;
  wire f_u_dadda_cla32_u_cla62_and58;
  wire f_u_dadda_cla32_u_cla62_and59;
  wire f_u_dadda_cla32_u_cla62_and60;
  wire f_u_dadda_cla32_u_cla62_and61;
  wire f_u_dadda_cla32_u_cla62_or29;
  wire f_u_dadda_cla32_u_cla62_or30;
  wire f_u_dadda_cla32_u_cla62_or31;
  wire f_u_dadda_cla32_u_cla62_pg_logic15_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic15_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic15_xor0;
  wire f_u_dadda_cla32_u_cla62_xor15;
  wire f_u_dadda_cla32_u_cla62_and62;
  wire f_u_dadda_cla32_u_cla62_and63;
  wire f_u_dadda_cla32_u_cla62_and64;
  wire f_u_dadda_cla32_u_cla62_and65;
  wire f_u_dadda_cla32_u_cla62_and66;
  wire f_u_dadda_cla32_u_cla62_and67;
  wire f_u_dadda_cla32_u_cla62_and68;
  wire f_u_dadda_cla32_u_cla62_and69;
  wire f_u_dadda_cla32_u_cla62_and70;
  wire f_u_dadda_cla32_u_cla62_and71;
  wire f_u_dadda_cla32_u_cla62_or32;
  wire f_u_dadda_cla32_u_cla62_or33;
  wire f_u_dadda_cla32_u_cla62_or34;
  wire f_u_dadda_cla32_u_cla62_or35;
  wire f_u_dadda_cla32_u_cla62_pg_logic16_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic16_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic16_xor0;
  wire f_u_dadda_cla32_u_cla62_xor16;
  wire f_u_dadda_cla32_u_cla62_and72;
  wire f_u_dadda_cla32_u_cla62_or36;
  wire f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic17_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic17_xor0;
  wire f_u_dadda_cla32_u_cla62_xor17;
  wire f_u_dadda_cla32_u_cla62_and73;
  wire f_u_dadda_cla32_u_cla62_and74;
  wire f_u_dadda_cla32_u_cla62_and75;
  wire f_u_dadda_cla32_u_cla62_or37;
  wire f_u_dadda_cla32_u_cla62_or38;
  wire f_u_dadda_cla32_u_cla62_pg_logic18_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic18_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic18_xor0;
  wire f_u_dadda_cla32_u_cla62_xor18;
  wire f_u_dadda_cla32_u_cla62_and76;
  wire f_u_dadda_cla32_u_cla62_and77;
  wire f_u_dadda_cla32_u_cla62_and78;
  wire f_u_dadda_cla32_u_cla62_and79;
  wire f_u_dadda_cla32_u_cla62_and80;
  wire f_u_dadda_cla32_u_cla62_and81;
  wire f_u_dadda_cla32_u_cla62_or39;
  wire f_u_dadda_cla32_u_cla62_or40;
  wire f_u_dadda_cla32_u_cla62_or41;
  wire f_u_dadda_cla32_u_cla62_pg_logic19_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic19_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic19_xor0;
  wire f_u_dadda_cla32_u_cla62_xor19;
  wire f_u_dadda_cla32_u_cla62_and82;
  wire f_u_dadda_cla32_u_cla62_and83;
  wire f_u_dadda_cla32_u_cla62_and84;
  wire f_u_dadda_cla32_u_cla62_and85;
  wire f_u_dadda_cla32_u_cla62_and86;
  wire f_u_dadda_cla32_u_cla62_and87;
  wire f_u_dadda_cla32_u_cla62_and88;
  wire f_u_dadda_cla32_u_cla62_and89;
  wire f_u_dadda_cla32_u_cla62_and90;
  wire f_u_dadda_cla32_u_cla62_and91;
  wire f_u_dadda_cla32_u_cla62_or42;
  wire f_u_dadda_cla32_u_cla62_or43;
  wire f_u_dadda_cla32_u_cla62_or44;
  wire f_u_dadda_cla32_u_cla62_or45;
  wire f_u_dadda_cla32_u_cla62_pg_logic20_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic20_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic20_xor0;
  wire f_u_dadda_cla32_u_cla62_xor20;
  wire f_u_dadda_cla32_u_cla62_and92;
  wire f_u_dadda_cla32_u_cla62_or46;
  wire f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic21_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic21_xor0;
  wire f_u_dadda_cla32_u_cla62_xor21;
  wire f_u_dadda_cla32_u_cla62_and93;
  wire f_u_dadda_cla32_u_cla62_and94;
  wire f_u_dadda_cla32_u_cla62_and95;
  wire f_u_dadda_cla32_u_cla62_or47;
  wire f_u_dadda_cla32_u_cla62_or48;
  wire f_u_dadda_cla32_u_cla62_pg_logic22_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic22_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic22_xor0;
  wire f_u_dadda_cla32_u_cla62_xor22;
  wire f_u_dadda_cla32_u_cla62_and96;
  wire f_u_dadda_cla32_u_cla62_and97;
  wire f_u_dadda_cla32_u_cla62_and98;
  wire f_u_dadda_cla32_u_cla62_and99;
  wire f_u_dadda_cla32_u_cla62_and100;
  wire f_u_dadda_cla32_u_cla62_and101;
  wire f_u_dadda_cla32_u_cla62_or49;
  wire f_u_dadda_cla32_u_cla62_or50;
  wire f_u_dadda_cla32_u_cla62_or51;
  wire f_u_dadda_cla32_u_cla62_pg_logic23_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic23_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic23_xor0;
  wire f_u_dadda_cla32_u_cla62_xor23;
  wire f_u_dadda_cla32_u_cla62_and102;
  wire f_u_dadda_cla32_u_cla62_and103;
  wire f_u_dadda_cla32_u_cla62_and104;
  wire f_u_dadda_cla32_u_cla62_and105;
  wire f_u_dadda_cla32_u_cla62_and106;
  wire f_u_dadda_cla32_u_cla62_and107;
  wire f_u_dadda_cla32_u_cla62_and108;
  wire f_u_dadda_cla32_u_cla62_and109;
  wire f_u_dadda_cla32_u_cla62_and110;
  wire f_u_dadda_cla32_u_cla62_and111;
  wire f_u_dadda_cla32_u_cla62_or52;
  wire f_u_dadda_cla32_u_cla62_or53;
  wire f_u_dadda_cla32_u_cla62_or54;
  wire f_u_dadda_cla32_u_cla62_or55;
  wire f_u_dadda_cla32_u_cla62_pg_logic24_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic24_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic24_xor0;
  wire f_u_dadda_cla32_u_cla62_xor24;
  wire f_u_dadda_cla32_u_cla62_and112;
  wire f_u_dadda_cla32_u_cla62_or56;
  wire f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic25_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic25_xor0;
  wire f_u_dadda_cla32_u_cla62_xor25;
  wire f_u_dadda_cla32_u_cla62_and113;
  wire f_u_dadda_cla32_u_cla62_and114;
  wire f_u_dadda_cla32_u_cla62_and115;
  wire f_u_dadda_cla32_u_cla62_or57;
  wire f_u_dadda_cla32_u_cla62_or58;
  wire f_u_dadda_cla32_u_cla62_pg_logic26_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic26_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic26_xor0;
  wire f_u_dadda_cla32_u_cla62_xor26;
  wire f_u_dadda_cla32_u_cla62_and116;
  wire f_u_dadda_cla32_u_cla62_and117;
  wire f_u_dadda_cla32_u_cla62_and118;
  wire f_u_dadda_cla32_u_cla62_and119;
  wire f_u_dadda_cla32_u_cla62_and120;
  wire f_u_dadda_cla32_u_cla62_and121;
  wire f_u_dadda_cla32_u_cla62_or59;
  wire f_u_dadda_cla32_u_cla62_or60;
  wire f_u_dadda_cla32_u_cla62_or61;
  wire f_u_dadda_cla32_u_cla62_pg_logic27_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic27_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic27_xor0;
  wire f_u_dadda_cla32_u_cla62_xor27;
  wire f_u_dadda_cla32_u_cla62_and122;
  wire f_u_dadda_cla32_u_cla62_and123;
  wire f_u_dadda_cla32_u_cla62_and124;
  wire f_u_dadda_cla32_u_cla62_and125;
  wire f_u_dadda_cla32_u_cla62_and126;
  wire f_u_dadda_cla32_u_cla62_and127;
  wire f_u_dadda_cla32_u_cla62_and128;
  wire f_u_dadda_cla32_u_cla62_and129;
  wire f_u_dadda_cla32_u_cla62_and130;
  wire f_u_dadda_cla32_u_cla62_and131;
  wire f_u_dadda_cla32_u_cla62_or62;
  wire f_u_dadda_cla32_u_cla62_or63;
  wire f_u_dadda_cla32_u_cla62_or64;
  wire f_u_dadda_cla32_u_cla62_or65;
  wire f_u_dadda_cla32_u_cla62_pg_logic28_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic28_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic28_xor0;
  wire f_u_dadda_cla32_u_cla62_xor28;
  wire f_u_dadda_cla32_u_cla62_and132;
  wire f_u_dadda_cla32_u_cla62_or66;
  wire f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic29_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic29_xor0;
  wire f_u_dadda_cla32_u_cla62_xor29;
  wire f_u_dadda_cla32_u_cla62_and133;
  wire f_u_dadda_cla32_u_cla62_and134;
  wire f_u_dadda_cla32_u_cla62_and135;
  wire f_u_dadda_cla32_u_cla62_or67;
  wire f_u_dadda_cla32_u_cla62_or68;
  wire f_u_dadda_cla32_u_cla62_pg_logic30_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic30_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic30_xor0;
  wire f_u_dadda_cla32_u_cla62_xor30;
  wire f_u_dadda_cla32_u_cla62_and136;
  wire f_u_dadda_cla32_u_cla62_and137;
  wire f_u_dadda_cla32_u_cla62_and138;
  wire f_u_dadda_cla32_u_cla62_and139;
  wire f_u_dadda_cla32_u_cla62_and140;
  wire f_u_dadda_cla32_u_cla62_and141;
  wire f_u_dadda_cla32_u_cla62_or69;
  wire f_u_dadda_cla32_u_cla62_or70;
  wire f_u_dadda_cla32_u_cla62_or71;
  wire f_u_dadda_cla32_u_cla62_pg_logic31_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic31_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic31_xor0;
  wire f_u_dadda_cla32_u_cla62_xor31;
  wire f_u_dadda_cla32_u_cla62_and142;
  wire f_u_dadda_cla32_u_cla62_and143;
  wire f_u_dadda_cla32_u_cla62_and144;
  wire f_u_dadda_cla32_u_cla62_and145;
  wire f_u_dadda_cla32_u_cla62_and146;
  wire f_u_dadda_cla32_u_cla62_and147;
  wire f_u_dadda_cla32_u_cla62_and148;
  wire f_u_dadda_cla32_u_cla62_and149;
  wire f_u_dadda_cla32_u_cla62_and150;
  wire f_u_dadda_cla32_u_cla62_and151;
  wire f_u_dadda_cla32_u_cla62_or72;
  wire f_u_dadda_cla32_u_cla62_or73;
  wire f_u_dadda_cla32_u_cla62_or74;
  wire f_u_dadda_cla32_u_cla62_or75;
  wire f_u_dadda_cla32_u_cla62_pg_logic32_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic32_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic32_xor0;
  wire f_u_dadda_cla32_u_cla62_xor32;
  wire f_u_dadda_cla32_u_cla62_and152;
  wire f_u_dadda_cla32_u_cla62_or76;
  wire f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic33_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic33_xor0;
  wire f_u_dadda_cla32_u_cla62_xor33;
  wire f_u_dadda_cla32_u_cla62_and153;
  wire f_u_dadda_cla32_u_cla62_and154;
  wire f_u_dadda_cla32_u_cla62_and155;
  wire f_u_dadda_cla32_u_cla62_or77;
  wire f_u_dadda_cla32_u_cla62_or78;
  wire f_u_dadda_cla32_u_cla62_pg_logic34_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic34_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic34_xor0;
  wire f_u_dadda_cla32_u_cla62_xor34;
  wire f_u_dadda_cla32_u_cla62_and156;
  wire f_u_dadda_cla32_u_cla62_and157;
  wire f_u_dadda_cla32_u_cla62_and158;
  wire f_u_dadda_cla32_u_cla62_and159;
  wire f_u_dadda_cla32_u_cla62_and160;
  wire f_u_dadda_cla32_u_cla62_and161;
  wire f_u_dadda_cla32_u_cla62_or79;
  wire f_u_dadda_cla32_u_cla62_or80;
  wire f_u_dadda_cla32_u_cla62_or81;
  wire f_u_dadda_cla32_u_cla62_pg_logic35_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic35_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic35_xor0;
  wire f_u_dadda_cla32_u_cla62_xor35;
  wire f_u_dadda_cla32_u_cla62_and162;
  wire f_u_dadda_cla32_u_cla62_and163;
  wire f_u_dadda_cla32_u_cla62_and164;
  wire f_u_dadda_cla32_u_cla62_and165;
  wire f_u_dadda_cla32_u_cla62_and166;
  wire f_u_dadda_cla32_u_cla62_and167;
  wire f_u_dadda_cla32_u_cla62_and168;
  wire f_u_dadda_cla32_u_cla62_and169;
  wire f_u_dadda_cla32_u_cla62_and170;
  wire f_u_dadda_cla32_u_cla62_and171;
  wire f_u_dadda_cla32_u_cla62_or82;
  wire f_u_dadda_cla32_u_cla62_or83;
  wire f_u_dadda_cla32_u_cla62_or84;
  wire f_u_dadda_cla32_u_cla62_or85;
  wire f_u_dadda_cla32_u_cla62_pg_logic36_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic36_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic36_xor0;
  wire f_u_dadda_cla32_u_cla62_xor36;
  wire f_u_dadda_cla32_u_cla62_and172;
  wire f_u_dadda_cla32_u_cla62_or86;
  wire f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic37_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic37_xor0;
  wire f_u_dadda_cla32_u_cla62_xor37;
  wire f_u_dadda_cla32_u_cla62_and173;
  wire f_u_dadda_cla32_u_cla62_and174;
  wire f_u_dadda_cla32_u_cla62_and175;
  wire f_u_dadda_cla32_u_cla62_or87;
  wire f_u_dadda_cla32_u_cla62_or88;
  wire f_u_dadda_cla32_u_cla62_pg_logic38_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic38_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic38_xor0;
  wire f_u_dadda_cla32_u_cla62_xor38;
  wire f_u_dadda_cla32_u_cla62_and176;
  wire f_u_dadda_cla32_u_cla62_and177;
  wire f_u_dadda_cla32_u_cla62_and178;
  wire f_u_dadda_cla32_u_cla62_and179;
  wire f_u_dadda_cla32_u_cla62_and180;
  wire f_u_dadda_cla32_u_cla62_and181;
  wire f_u_dadda_cla32_u_cla62_or89;
  wire f_u_dadda_cla32_u_cla62_or90;
  wire f_u_dadda_cla32_u_cla62_or91;
  wire f_u_dadda_cla32_u_cla62_pg_logic39_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic39_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic39_xor0;
  wire f_u_dadda_cla32_u_cla62_xor39;
  wire f_u_dadda_cla32_u_cla62_and182;
  wire f_u_dadda_cla32_u_cla62_and183;
  wire f_u_dadda_cla32_u_cla62_and184;
  wire f_u_dadda_cla32_u_cla62_and185;
  wire f_u_dadda_cla32_u_cla62_and186;
  wire f_u_dadda_cla32_u_cla62_and187;
  wire f_u_dadda_cla32_u_cla62_and188;
  wire f_u_dadda_cla32_u_cla62_and189;
  wire f_u_dadda_cla32_u_cla62_and190;
  wire f_u_dadda_cla32_u_cla62_and191;
  wire f_u_dadda_cla32_u_cla62_or92;
  wire f_u_dadda_cla32_u_cla62_or93;
  wire f_u_dadda_cla32_u_cla62_or94;
  wire f_u_dadda_cla32_u_cla62_or95;
  wire f_u_dadda_cla32_u_cla62_pg_logic40_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic40_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic40_xor0;
  wire f_u_dadda_cla32_u_cla62_xor40;
  wire f_u_dadda_cla32_u_cla62_and192;
  wire f_u_dadda_cla32_u_cla62_or96;
  wire f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic41_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic41_xor0;
  wire f_u_dadda_cla32_u_cla62_xor41;
  wire f_u_dadda_cla32_u_cla62_and193;
  wire f_u_dadda_cla32_u_cla62_and194;
  wire f_u_dadda_cla32_u_cla62_and195;
  wire f_u_dadda_cla32_u_cla62_or97;
  wire f_u_dadda_cla32_u_cla62_or98;
  wire f_u_dadda_cla32_u_cla62_pg_logic42_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic42_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic42_xor0;
  wire f_u_dadda_cla32_u_cla62_xor42;
  wire f_u_dadda_cla32_u_cla62_and196;
  wire f_u_dadda_cla32_u_cla62_and197;
  wire f_u_dadda_cla32_u_cla62_and198;
  wire f_u_dadda_cla32_u_cla62_and199;
  wire f_u_dadda_cla32_u_cla62_and200;
  wire f_u_dadda_cla32_u_cla62_and201;
  wire f_u_dadda_cla32_u_cla62_or99;
  wire f_u_dadda_cla32_u_cla62_or100;
  wire f_u_dadda_cla32_u_cla62_or101;
  wire f_u_dadda_cla32_u_cla62_pg_logic43_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic43_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic43_xor0;
  wire f_u_dadda_cla32_u_cla62_xor43;
  wire f_u_dadda_cla32_u_cla62_and202;
  wire f_u_dadda_cla32_u_cla62_and203;
  wire f_u_dadda_cla32_u_cla62_and204;
  wire f_u_dadda_cla32_u_cla62_and205;
  wire f_u_dadda_cla32_u_cla62_and206;
  wire f_u_dadda_cla32_u_cla62_and207;
  wire f_u_dadda_cla32_u_cla62_and208;
  wire f_u_dadda_cla32_u_cla62_and209;
  wire f_u_dadda_cla32_u_cla62_and210;
  wire f_u_dadda_cla32_u_cla62_and211;
  wire f_u_dadda_cla32_u_cla62_or102;
  wire f_u_dadda_cla32_u_cla62_or103;
  wire f_u_dadda_cla32_u_cla62_or104;
  wire f_u_dadda_cla32_u_cla62_or105;
  wire f_u_dadda_cla32_u_cla62_pg_logic44_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic44_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic44_xor0;
  wire f_u_dadda_cla32_u_cla62_xor44;
  wire f_u_dadda_cla32_u_cla62_and212;
  wire f_u_dadda_cla32_u_cla62_or106;
  wire f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic45_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic45_xor0;
  wire f_u_dadda_cla32_u_cla62_xor45;
  wire f_u_dadda_cla32_u_cla62_and213;
  wire f_u_dadda_cla32_u_cla62_and214;
  wire f_u_dadda_cla32_u_cla62_and215;
  wire f_u_dadda_cla32_u_cla62_or107;
  wire f_u_dadda_cla32_u_cla62_or108;
  wire f_u_dadda_cla32_u_cla62_pg_logic46_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic46_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic46_xor0;
  wire f_u_dadda_cla32_u_cla62_xor46;
  wire f_u_dadda_cla32_u_cla62_and216;
  wire f_u_dadda_cla32_u_cla62_and217;
  wire f_u_dadda_cla32_u_cla62_and218;
  wire f_u_dadda_cla32_u_cla62_and219;
  wire f_u_dadda_cla32_u_cla62_and220;
  wire f_u_dadda_cla32_u_cla62_and221;
  wire f_u_dadda_cla32_u_cla62_or109;
  wire f_u_dadda_cla32_u_cla62_or110;
  wire f_u_dadda_cla32_u_cla62_or111;
  wire f_u_dadda_cla32_u_cla62_pg_logic47_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic47_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic47_xor0;
  wire f_u_dadda_cla32_u_cla62_xor47;
  wire f_u_dadda_cla32_u_cla62_and222;
  wire f_u_dadda_cla32_u_cla62_and223;
  wire f_u_dadda_cla32_u_cla62_and224;
  wire f_u_dadda_cla32_u_cla62_and225;
  wire f_u_dadda_cla32_u_cla62_and226;
  wire f_u_dadda_cla32_u_cla62_and227;
  wire f_u_dadda_cla32_u_cla62_and228;
  wire f_u_dadda_cla32_u_cla62_and229;
  wire f_u_dadda_cla32_u_cla62_and230;
  wire f_u_dadda_cla32_u_cla62_and231;
  wire f_u_dadda_cla32_u_cla62_or112;
  wire f_u_dadda_cla32_u_cla62_or113;
  wire f_u_dadda_cla32_u_cla62_or114;
  wire f_u_dadda_cla32_u_cla62_or115;
  wire f_u_dadda_cla32_u_cla62_pg_logic48_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic48_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic48_xor0;
  wire f_u_dadda_cla32_u_cla62_xor48;
  wire f_u_dadda_cla32_u_cla62_and232;
  wire f_u_dadda_cla32_u_cla62_or116;
  wire f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic49_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic49_xor0;
  wire f_u_dadda_cla32_u_cla62_xor49;
  wire f_u_dadda_cla32_u_cla62_and233;
  wire f_u_dadda_cla32_u_cla62_and234;
  wire f_u_dadda_cla32_u_cla62_and235;
  wire f_u_dadda_cla32_u_cla62_or117;
  wire f_u_dadda_cla32_u_cla62_or118;
  wire f_u_dadda_cla32_u_cla62_pg_logic50_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic50_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic50_xor0;
  wire f_u_dadda_cla32_u_cla62_xor50;
  wire f_u_dadda_cla32_u_cla62_and236;
  wire f_u_dadda_cla32_u_cla62_and237;
  wire f_u_dadda_cla32_u_cla62_and238;
  wire f_u_dadda_cla32_u_cla62_and239;
  wire f_u_dadda_cla32_u_cla62_and240;
  wire f_u_dadda_cla32_u_cla62_and241;
  wire f_u_dadda_cla32_u_cla62_or119;
  wire f_u_dadda_cla32_u_cla62_or120;
  wire f_u_dadda_cla32_u_cla62_or121;
  wire f_u_dadda_cla32_u_cla62_pg_logic51_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic51_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic51_xor0;
  wire f_u_dadda_cla32_u_cla62_xor51;
  wire f_u_dadda_cla32_u_cla62_and242;
  wire f_u_dadda_cla32_u_cla62_and243;
  wire f_u_dadda_cla32_u_cla62_and244;
  wire f_u_dadda_cla32_u_cla62_and245;
  wire f_u_dadda_cla32_u_cla62_and246;
  wire f_u_dadda_cla32_u_cla62_and247;
  wire f_u_dadda_cla32_u_cla62_and248;
  wire f_u_dadda_cla32_u_cla62_and249;
  wire f_u_dadda_cla32_u_cla62_and250;
  wire f_u_dadda_cla32_u_cla62_and251;
  wire f_u_dadda_cla32_u_cla62_or122;
  wire f_u_dadda_cla32_u_cla62_or123;
  wire f_u_dadda_cla32_u_cla62_or124;
  wire f_u_dadda_cla32_u_cla62_or125;
  wire f_u_dadda_cla32_u_cla62_pg_logic52_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic52_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic52_xor0;
  wire f_u_dadda_cla32_u_cla62_xor52;
  wire f_u_dadda_cla32_u_cla62_and252;
  wire f_u_dadda_cla32_u_cla62_or126;
  wire f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic53_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic53_xor0;
  wire f_u_dadda_cla32_u_cla62_xor53;
  wire f_u_dadda_cla32_u_cla62_and253;
  wire f_u_dadda_cla32_u_cla62_and254;
  wire f_u_dadda_cla32_u_cla62_and255;
  wire f_u_dadda_cla32_u_cla62_or127;
  wire f_u_dadda_cla32_u_cla62_or128;
  wire f_u_dadda_cla32_u_cla62_pg_logic54_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic54_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic54_xor0;
  wire f_u_dadda_cla32_u_cla62_xor54;
  wire f_u_dadda_cla32_u_cla62_and256;
  wire f_u_dadda_cla32_u_cla62_and257;
  wire f_u_dadda_cla32_u_cla62_and258;
  wire f_u_dadda_cla32_u_cla62_and259;
  wire f_u_dadda_cla32_u_cla62_and260;
  wire f_u_dadda_cla32_u_cla62_and261;
  wire f_u_dadda_cla32_u_cla62_or129;
  wire f_u_dadda_cla32_u_cla62_or130;
  wire f_u_dadda_cla32_u_cla62_or131;
  wire f_u_dadda_cla32_u_cla62_pg_logic55_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic55_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic55_xor0;
  wire f_u_dadda_cla32_u_cla62_xor55;
  wire f_u_dadda_cla32_u_cla62_and262;
  wire f_u_dadda_cla32_u_cla62_and263;
  wire f_u_dadda_cla32_u_cla62_and264;
  wire f_u_dadda_cla32_u_cla62_and265;
  wire f_u_dadda_cla32_u_cla62_and266;
  wire f_u_dadda_cla32_u_cla62_and267;
  wire f_u_dadda_cla32_u_cla62_and268;
  wire f_u_dadda_cla32_u_cla62_and269;
  wire f_u_dadda_cla32_u_cla62_and270;
  wire f_u_dadda_cla32_u_cla62_and271;
  wire f_u_dadda_cla32_u_cla62_or132;
  wire f_u_dadda_cla32_u_cla62_or133;
  wire f_u_dadda_cla32_u_cla62_or134;
  wire f_u_dadda_cla32_u_cla62_or135;
  wire f_u_dadda_cla32_u_cla62_pg_logic56_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic56_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic56_xor0;
  wire f_u_dadda_cla32_u_cla62_xor56;
  wire f_u_dadda_cla32_u_cla62_and272;
  wire f_u_dadda_cla32_u_cla62_or136;
  wire f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic57_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic57_xor0;
  wire f_u_dadda_cla32_u_cla62_xor57;
  wire f_u_dadda_cla32_u_cla62_and273;
  wire f_u_dadda_cla32_u_cla62_and274;
  wire f_u_dadda_cla32_u_cla62_and275;
  wire f_u_dadda_cla32_u_cla62_or137;
  wire f_u_dadda_cla32_u_cla62_or138;
  wire f_u_dadda_cla32_u_cla62_pg_logic58_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic58_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic58_xor0;
  wire f_u_dadda_cla32_u_cla62_xor58;
  wire f_u_dadda_cla32_u_cla62_and276;
  wire f_u_dadda_cla32_u_cla62_and277;
  wire f_u_dadda_cla32_u_cla62_and278;
  wire f_u_dadda_cla32_u_cla62_and279;
  wire f_u_dadda_cla32_u_cla62_and280;
  wire f_u_dadda_cla32_u_cla62_and281;
  wire f_u_dadda_cla32_u_cla62_or139;
  wire f_u_dadda_cla32_u_cla62_or140;
  wire f_u_dadda_cla32_u_cla62_or141;
  wire f_u_dadda_cla32_u_cla62_pg_logic59_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic59_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic59_xor0;
  wire f_u_dadda_cla32_u_cla62_xor59;
  wire f_u_dadda_cla32_u_cla62_and282;
  wire f_u_dadda_cla32_u_cla62_and283;
  wire f_u_dadda_cla32_u_cla62_and284;
  wire f_u_dadda_cla32_u_cla62_and285;
  wire f_u_dadda_cla32_u_cla62_and286;
  wire f_u_dadda_cla32_u_cla62_and287;
  wire f_u_dadda_cla32_u_cla62_and288;
  wire f_u_dadda_cla32_u_cla62_and289;
  wire f_u_dadda_cla32_u_cla62_and290;
  wire f_u_dadda_cla32_u_cla62_and291;
  wire f_u_dadda_cla32_u_cla62_or142;
  wire f_u_dadda_cla32_u_cla62_or143;
  wire f_u_dadda_cla32_u_cla62_or144;
  wire f_u_dadda_cla32_u_cla62_or145;
  wire f_u_dadda_cla32_u_cla62_pg_logic60_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic60_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic60_xor0;
  wire f_u_dadda_cla32_u_cla62_xor60;
  wire f_u_dadda_cla32_u_cla62_and292;
  wire f_u_dadda_cla32_u_cla62_or146;
  wire f_u_dadda_cla32_u_cla62_pg_logic61_or0;
  wire f_u_dadda_cla32_u_cla62_pg_logic61_and0;
  wire f_u_dadda_cla32_u_cla62_pg_logic61_xor0;
  wire f_u_dadda_cla32_u_cla62_xor61;
  wire f_u_dadda_cla32_u_cla62_and293;
  wire f_u_dadda_cla32_u_cla62_and294;
  wire f_u_dadda_cla32_u_cla62_and295;
  wire f_u_dadda_cla32_u_cla62_or147;
  wire f_u_dadda_cla32_u_cla62_or148;

  assign f_u_dadda_cla32_and_28_0 = a[28] & b[0];
  assign f_u_dadda_cla32_and_27_1 = a[27] & b[1];
  assign f_u_dadda_cla32_ha0_xor0 = f_u_dadda_cla32_and_28_0 ^ f_u_dadda_cla32_and_27_1;
  assign f_u_dadda_cla32_ha0_and0 = f_u_dadda_cla32_and_28_0 & f_u_dadda_cla32_and_27_1;
  assign f_u_dadda_cla32_and_29_0 = a[29] & b[0];
  assign f_u_dadda_cla32_and_28_1 = a[28] & b[1];
  assign f_u_dadda_cla32_fa0_xor0 = f_u_dadda_cla32_ha0_and0 ^ f_u_dadda_cla32_and_29_0;
  assign f_u_dadda_cla32_fa0_and0 = f_u_dadda_cla32_ha0_and0 & f_u_dadda_cla32_and_29_0;
  assign f_u_dadda_cla32_fa0_xor1 = f_u_dadda_cla32_fa0_xor0 ^ f_u_dadda_cla32_and_28_1;
  assign f_u_dadda_cla32_fa0_and1 = f_u_dadda_cla32_fa0_xor0 & f_u_dadda_cla32_and_28_1;
  assign f_u_dadda_cla32_fa0_or0 = f_u_dadda_cla32_fa0_and0 | f_u_dadda_cla32_fa0_and1;
  assign f_u_dadda_cla32_and_27_2 = a[27] & b[2];
  assign f_u_dadda_cla32_and_26_3 = a[26] & b[3];
  assign f_u_dadda_cla32_ha1_xor0 = f_u_dadda_cla32_and_27_2 ^ f_u_dadda_cla32_and_26_3;
  assign f_u_dadda_cla32_ha1_and0 = f_u_dadda_cla32_and_27_2 & f_u_dadda_cla32_and_26_3;
  assign f_u_dadda_cla32_and_30_0 = a[30] & b[0];
  assign f_u_dadda_cla32_fa1_xor0 = f_u_dadda_cla32_ha1_and0 ^ f_u_dadda_cla32_fa0_or0;
  assign f_u_dadda_cla32_fa1_and0 = f_u_dadda_cla32_ha1_and0 & f_u_dadda_cla32_fa0_or0;
  assign f_u_dadda_cla32_fa1_xor1 = f_u_dadda_cla32_fa1_xor0 ^ f_u_dadda_cla32_and_30_0;
  assign f_u_dadda_cla32_fa1_and1 = f_u_dadda_cla32_fa1_xor0 & f_u_dadda_cla32_and_30_0;
  assign f_u_dadda_cla32_fa1_or0 = f_u_dadda_cla32_fa1_and0 | f_u_dadda_cla32_fa1_and1;
  assign f_u_dadda_cla32_and_29_1 = a[29] & b[1];
  assign f_u_dadda_cla32_and_28_2 = a[28] & b[2];
  assign f_u_dadda_cla32_and_27_3 = a[27] & b[3];
  assign f_u_dadda_cla32_fa2_xor0 = f_u_dadda_cla32_and_29_1 ^ f_u_dadda_cla32_and_28_2;
  assign f_u_dadda_cla32_fa2_and0 = f_u_dadda_cla32_and_29_1 & f_u_dadda_cla32_and_28_2;
  assign f_u_dadda_cla32_fa2_xor1 = f_u_dadda_cla32_fa2_xor0 ^ f_u_dadda_cla32_and_27_3;
  assign f_u_dadda_cla32_fa2_and1 = f_u_dadda_cla32_fa2_xor0 & f_u_dadda_cla32_and_27_3;
  assign f_u_dadda_cla32_fa2_or0 = f_u_dadda_cla32_fa2_and0 | f_u_dadda_cla32_fa2_and1;
  assign f_u_dadda_cla32_and_26_4 = a[26] & b[4];
  assign f_u_dadda_cla32_and_25_5 = a[25] & b[5];
  assign f_u_dadda_cla32_ha2_xor0 = f_u_dadda_cla32_and_26_4 ^ f_u_dadda_cla32_and_25_5;
  assign f_u_dadda_cla32_ha2_and0 = f_u_dadda_cla32_and_26_4 & f_u_dadda_cla32_and_25_5;
  assign f_u_dadda_cla32_fa3_xor0 = f_u_dadda_cla32_ha2_and0 ^ f_u_dadda_cla32_fa2_or0;
  assign f_u_dadda_cla32_fa3_and0 = f_u_dadda_cla32_ha2_and0 & f_u_dadda_cla32_fa2_or0;
  assign f_u_dadda_cla32_fa3_xor1 = f_u_dadda_cla32_fa3_xor0 ^ f_u_dadda_cla32_fa1_or0;
  assign f_u_dadda_cla32_fa3_and1 = f_u_dadda_cla32_fa3_xor0 & f_u_dadda_cla32_fa1_or0;
  assign f_u_dadda_cla32_fa3_or0 = f_u_dadda_cla32_fa3_and0 | f_u_dadda_cla32_fa3_and1;
  assign f_u_dadda_cla32_and_31_0 = a[31] & b[0];
  assign f_u_dadda_cla32_and_30_1 = a[30] & b[1];
  assign f_u_dadda_cla32_and_29_2 = a[29] & b[2];
  assign f_u_dadda_cla32_fa4_xor0 = f_u_dadda_cla32_and_31_0 ^ f_u_dadda_cla32_and_30_1;
  assign f_u_dadda_cla32_fa4_and0 = f_u_dadda_cla32_and_31_0 & f_u_dadda_cla32_and_30_1;
  assign f_u_dadda_cla32_fa4_xor1 = f_u_dadda_cla32_fa4_xor0 ^ f_u_dadda_cla32_and_29_2;
  assign f_u_dadda_cla32_fa4_and1 = f_u_dadda_cla32_fa4_xor0 & f_u_dadda_cla32_and_29_2;
  assign f_u_dadda_cla32_fa4_or0 = f_u_dadda_cla32_fa4_and0 | f_u_dadda_cla32_fa4_and1;
  assign f_u_dadda_cla32_and_28_3 = a[28] & b[3];
  assign f_u_dadda_cla32_and_27_4 = a[27] & b[4];
  assign f_u_dadda_cla32_and_26_5 = a[26] & b[5];
  assign f_u_dadda_cla32_fa5_xor0 = f_u_dadda_cla32_and_28_3 ^ f_u_dadda_cla32_and_27_4;
  assign f_u_dadda_cla32_fa5_and0 = f_u_dadda_cla32_and_28_3 & f_u_dadda_cla32_and_27_4;
  assign f_u_dadda_cla32_fa5_xor1 = f_u_dadda_cla32_fa5_xor0 ^ f_u_dadda_cla32_and_26_5;
  assign f_u_dadda_cla32_fa5_and1 = f_u_dadda_cla32_fa5_xor0 & f_u_dadda_cla32_and_26_5;
  assign f_u_dadda_cla32_fa5_or0 = f_u_dadda_cla32_fa5_and0 | f_u_dadda_cla32_fa5_and1;
  assign f_u_dadda_cla32_and_25_6 = a[25] & b[6];
  assign f_u_dadda_cla32_and_24_7 = a[24] & b[7];
  assign f_u_dadda_cla32_ha3_xor0 = f_u_dadda_cla32_and_25_6 ^ f_u_dadda_cla32_and_24_7;
  assign f_u_dadda_cla32_ha3_and0 = f_u_dadda_cla32_and_25_6 & f_u_dadda_cla32_and_24_7;
  assign f_u_dadda_cla32_fa6_xor0 = f_u_dadda_cla32_ha3_and0 ^ f_u_dadda_cla32_fa5_or0;
  assign f_u_dadda_cla32_fa6_and0 = f_u_dadda_cla32_ha3_and0 & f_u_dadda_cla32_fa5_or0;
  assign f_u_dadda_cla32_fa6_xor1 = f_u_dadda_cla32_fa6_xor0 ^ f_u_dadda_cla32_fa4_or0;
  assign f_u_dadda_cla32_fa6_and1 = f_u_dadda_cla32_fa6_xor0 & f_u_dadda_cla32_fa4_or0;
  assign f_u_dadda_cla32_fa6_or0 = f_u_dadda_cla32_fa6_and0 | f_u_dadda_cla32_fa6_and1;
  assign f_u_dadda_cla32_and_31_1 = a[31] & b[1];
  assign f_u_dadda_cla32_and_30_2 = a[30] & b[2];
  assign f_u_dadda_cla32_fa7_xor0 = f_u_dadda_cla32_fa3_or0 ^ f_u_dadda_cla32_and_31_1;
  assign f_u_dadda_cla32_fa7_and0 = f_u_dadda_cla32_fa3_or0 & f_u_dadda_cla32_and_31_1;
  assign f_u_dadda_cla32_fa7_xor1 = f_u_dadda_cla32_fa7_xor0 ^ f_u_dadda_cla32_and_30_2;
  assign f_u_dadda_cla32_fa7_and1 = f_u_dadda_cla32_fa7_xor0 & f_u_dadda_cla32_and_30_2;
  assign f_u_dadda_cla32_fa7_or0 = f_u_dadda_cla32_fa7_and0 | f_u_dadda_cla32_fa7_and1;
  assign f_u_dadda_cla32_and_29_3 = a[29] & b[3];
  assign f_u_dadda_cla32_and_28_4 = a[28] & b[4];
  assign f_u_dadda_cla32_and_27_5 = a[27] & b[5];
  assign f_u_dadda_cla32_fa8_xor0 = f_u_dadda_cla32_and_29_3 ^ f_u_dadda_cla32_and_28_4;
  assign f_u_dadda_cla32_fa8_and0 = f_u_dadda_cla32_and_29_3 & f_u_dadda_cla32_and_28_4;
  assign f_u_dadda_cla32_fa8_xor1 = f_u_dadda_cla32_fa8_xor0 ^ f_u_dadda_cla32_and_27_5;
  assign f_u_dadda_cla32_fa8_and1 = f_u_dadda_cla32_fa8_xor0 & f_u_dadda_cla32_and_27_5;
  assign f_u_dadda_cla32_fa8_or0 = f_u_dadda_cla32_fa8_and0 | f_u_dadda_cla32_fa8_and1;
  assign f_u_dadda_cla32_and_26_6 = a[26] & b[6];
  assign f_u_dadda_cla32_and_25_7 = a[25] & b[7];
  assign f_u_dadda_cla32_ha4_xor0 = f_u_dadda_cla32_and_26_6 ^ f_u_dadda_cla32_and_25_7;
  assign f_u_dadda_cla32_ha4_and0 = f_u_dadda_cla32_and_26_6 & f_u_dadda_cla32_and_25_7;
  assign f_u_dadda_cla32_fa9_xor0 = f_u_dadda_cla32_ha4_and0 ^ f_u_dadda_cla32_fa8_or0;
  assign f_u_dadda_cla32_fa9_and0 = f_u_dadda_cla32_ha4_and0 & f_u_dadda_cla32_fa8_or0;
  assign f_u_dadda_cla32_fa9_xor1 = f_u_dadda_cla32_fa9_xor0 ^ f_u_dadda_cla32_fa7_or0;
  assign f_u_dadda_cla32_fa9_and1 = f_u_dadda_cla32_fa9_xor0 & f_u_dadda_cla32_fa7_or0;
  assign f_u_dadda_cla32_fa9_or0 = f_u_dadda_cla32_fa9_and0 | f_u_dadda_cla32_fa9_and1;
  assign f_u_dadda_cla32_and_31_2 = a[31] & b[2];
  assign f_u_dadda_cla32_and_30_3 = a[30] & b[3];
  assign f_u_dadda_cla32_fa10_xor0 = f_u_dadda_cla32_fa6_or0 ^ f_u_dadda_cla32_and_31_2;
  assign f_u_dadda_cla32_fa10_and0 = f_u_dadda_cla32_fa6_or0 & f_u_dadda_cla32_and_31_2;
  assign f_u_dadda_cla32_fa10_xor1 = f_u_dadda_cla32_fa10_xor0 ^ f_u_dadda_cla32_and_30_3;
  assign f_u_dadda_cla32_fa10_and1 = f_u_dadda_cla32_fa10_xor0 & f_u_dadda_cla32_and_30_3;
  assign f_u_dadda_cla32_fa10_or0 = f_u_dadda_cla32_fa10_and0 | f_u_dadda_cla32_fa10_and1;
  assign f_u_dadda_cla32_and_29_4 = a[29] & b[4];
  assign f_u_dadda_cla32_and_28_5 = a[28] & b[5];
  assign f_u_dadda_cla32_and_27_6 = a[27] & b[6];
  assign f_u_dadda_cla32_fa11_xor0 = f_u_dadda_cla32_and_29_4 ^ f_u_dadda_cla32_and_28_5;
  assign f_u_dadda_cla32_fa11_and0 = f_u_dadda_cla32_and_29_4 & f_u_dadda_cla32_and_28_5;
  assign f_u_dadda_cla32_fa11_xor1 = f_u_dadda_cla32_fa11_xor0 ^ f_u_dadda_cla32_and_27_6;
  assign f_u_dadda_cla32_fa11_and1 = f_u_dadda_cla32_fa11_xor0 & f_u_dadda_cla32_and_27_6;
  assign f_u_dadda_cla32_fa11_or0 = f_u_dadda_cla32_fa11_and0 | f_u_dadda_cla32_fa11_and1;
  assign f_u_dadda_cla32_fa12_xor0 = f_u_dadda_cla32_fa11_or0 ^ f_u_dadda_cla32_fa10_or0;
  assign f_u_dadda_cla32_fa12_and0 = f_u_dadda_cla32_fa11_or0 & f_u_dadda_cla32_fa10_or0;
  assign f_u_dadda_cla32_fa12_xor1 = f_u_dadda_cla32_fa12_xor0 ^ f_u_dadda_cla32_fa9_or0;
  assign f_u_dadda_cla32_fa12_and1 = f_u_dadda_cla32_fa12_xor0 & f_u_dadda_cla32_fa9_or0;
  assign f_u_dadda_cla32_fa12_or0 = f_u_dadda_cla32_fa12_and0 | f_u_dadda_cla32_fa12_and1;
  assign f_u_dadda_cla32_and_31_3 = a[31] & b[3];
  assign f_u_dadda_cla32_and_30_4 = a[30] & b[4];
  assign f_u_dadda_cla32_and_29_5 = a[29] & b[5];
  assign f_u_dadda_cla32_fa13_xor0 = f_u_dadda_cla32_and_31_3 ^ f_u_dadda_cla32_and_30_4;
  assign f_u_dadda_cla32_fa13_and0 = f_u_dadda_cla32_and_31_3 & f_u_dadda_cla32_and_30_4;
  assign f_u_dadda_cla32_fa13_xor1 = f_u_dadda_cla32_fa13_xor0 ^ f_u_dadda_cla32_and_29_5;
  assign f_u_dadda_cla32_fa13_and1 = f_u_dadda_cla32_fa13_xor0 & f_u_dadda_cla32_and_29_5;
  assign f_u_dadda_cla32_fa13_or0 = f_u_dadda_cla32_fa13_and0 | f_u_dadda_cla32_fa13_and1;
  assign f_u_dadda_cla32_and_31_4 = a[31] & b[4];
  assign f_u_dadda_cla32_fa14_xor0 = f_u_dadda_cla32_fa13_or0 ^ f_u_dadda_cla32_fa12_or0;
  assign f_u_dadda_cla32_fa14_and0 = f_u_dadda_cla32_fa13_or0 & f_u_dadda_cla32_fa12_or0;
  assign f_u_dadda_cla32_fa14_xor1 = f_u_dadda_cla32_fa14_xor0 ^ f_u_dadda_cla32_and_31_4;
  assign f_u_dadda_cla32_fa14_and1 = f_u_dadda_cla32_fa14_xor0 & f_u_dadda_cla32_and_31_4;
  assign f_u_dadda_cla32_fa14_or0 = f_u_dadda_cla32_fa14_and0 | f_u_dadda_cla32_fa14_and1;
  assign f_u_dadda_cla32_and_6_0 = a[6] & b[0];
  assign f_u_dadda_cla32_and_5_1 = a[5] & b[1];
  assign f_u_dadda_cla32_ha5_xor0 = f_u_dadda_cla32_and_6_0 ^ f_u_dadda_cla32_and_5_1;
  assign f_u_dadda_cla32_ha5_and0 = f_u_dadda_cla32_and_6_0 & f_u_dadda_cla32_and_5_1;
  assign f_u_dadda_cla32_and_7_0 = a[7] & b[0];
  assign f_u_dadda_cla32_and_6_1 = a[6] & b[1];
  assign f_u_dadda_cla32_fa15_xor0 = f_u_dadda_cla32_ha5_and0 ^ f_u_dadda_cla32_and_7_0;
  assign f_u_dadda_cla32_fa15_and0 = f_u_dadda_cla32_ha5_and0 & f_u_dadda_cla32_and_7_0;
  assign f_u_dadda_cla32_fa15_xor1 = f_u_dadda_cla32_fa15_xor0 ^ f_u_dadda_cla32_and_6_1;
  assign f_u_dadda_cla32_fa15_and1 = f_u_dadda_cla32_fa15_xor0 & f_u_dadda_cla32_and_6_1;
  assign f_u_dadda_cla32_fa15_or0 = f_u_dadda_cla32_fa15_and0 | f_u_dadda_cla32_fa15_and1;
  assign f_u_dadda_cla32_and_5_2 = a[5] & b[2];
  assign f_u_dadda_cla32_and_4_3 = a[4] & b[3];
  assign f_u_dadda_cla32_ha6_xor0 = f_u_dadda_cla32_and_5_2 ^ f_u_dadda_cla32_and_4_3;
  assign f_u_dadda_cla32_ha6_and0 = f_u_dadda_cla32_and_5_2 & f_u_dadda_cla32_and_4_3;
  assign f_u_dadda_cla32_and_8_0 = a[8] & b[0];
  assign f_u_dadda_cla32_fa16_xor0 = f_u_dadda_cla32_ha6_and0 ^ f_u_dadda_cla32_fa15_or0;
  assign f_u_dadda_cla32_fa16_and0 = f_u_dadda_cla32_ha6_and0 & f_u_dadda_cla32_fa15_or0;
  assign f_u_dadda_cla32_fa16_xor1 = f_u_dadda_cla32_fa16_xor0 ^ f_u_dadda_cla32_and_8_0;
  assign f_u_dadda_cla32_fa16_and1 = f_u_dadda_cla32_fa16_xor0 & f_u_dadda_cla32_and_8_0;
  assign f_u_dadda_cla32_fa16_or0 = f_u_dadda_cla32_fa16_and0 | f_u_dadda_cla32_fa16_and1;
  assign f_u_dadda_cla32_and_7_1 = a[7] & b[1];
  assign f_u_dadda_cla32_and_6_2 = a[6] & b[2];
  assign f_u_dadda_cla32_and_5_3 = a[5] & b[3];
  assign f_u_dadda_cla32_fa17_xor0 = f_u_dadda_cla32_and_7_1 ^ f_u_dadda_cla32_and_6_2;
  assign f_u_dadda_cla32_fa17_and0 = f_u_dadda_cla32_and_7_1 & f_u_dadda_cla32_and_6_2;
  assign f_u_dadda_cla32_fa17_xor1 = f_u_dadda_cla32_fa17_xor0 ^ f_u_dadda_cla32_and_5_3;
  assign f_u_dadda_cla32_fa17_and1 = f_u_dadda_cla32_fa17_xor0 & f_u_dadda_cla32_and_5_3;
  assign f_u_dadda_cla32_fa17_or0 = f_u_dadda_cla32_fa17_and0 | f_u_dadda_cla32_fa17_and1;
  assign f_u_dadda_cla32_and_4_4 = a[4] & b[4];
  assign f_u_dadda_cla32_and_3_5 = a[3] & b[5];
  assign f_u_dadda_cla32_ha7_xor0 = f_u_dadda_cla32_and_4_4 ^ f_u_dadda_cla32_and_3_5;
  assign f_u_dadda_cla32_ha7_and0 = f_u_dadda_cla32_and_4_4 & f_u_dadda_cla32_and_3_5;
  assign f_u_dadda_cla32_fa18_xor0 = f_u_dadda_cla32_ha7_and0 ^ f_u_dadda_cla32_fa17_or0;
  assign f_u_dadda_cla32_fa18_and0 = f_u_dadda_cla32_ha7_and0 & f_u_dadda_cla32_fa17_or0;
  assign f_u_dadda_cla32_fa18_xor1 = f_u_dadda_cla32_fa18_xor0 ^ f_u_dadda_cla32_fa16_or0;
  assign f_u_dadda_cla32_fa18_and1 = f_u_dadda_cla32_fa18_xor0 & f_u_dadda_cla32_fa16_or0;
  assign f_u_dadda_cla32_fa18_or0 = f_u_dadda_cla32_fa18_and0 | f_u_dadda_cla32_fa18_and1;
  assign f_u_dadda_cla32_and_9_0 = a[9] & b[0];
  assign f_u_dadda_cla32_and_8_1 = a[8] & b[1];
  assign f_u_dadda_cla32_and_7_2 = a[7] & b[2];
  assign f_u_dadda_cla32_fa19_xor0 = f_u_dadda_cla32_and_9_0 ^ f_u_dadda_cla32_and_8_1;
  assign f_u_dadda_cla32_fa19_and0 = f_u_dadda_cla32_and_9_0 & f_u_dadda_cla32_and_8_1;
  assign f_u_dadda_cla32_fa19_xor1 = f_u_dadda_cla32_fa19_xor0 ^ f_u_dadda_cla32_and_7_2;
  assign f_u_dadda_cla32_fa19_and1 = f_u_dadda_cla32_fa19_xor0 & f_u_dadda_cla32_and_7_2;
  assign f_u_dadda_cla32_fa19_or0 = f_u_dadda_cla32_fa19_and0 | f_u_dadda_cla32_fa19_and1;
  assign f_u_dadda_cla32_and_6_3 = a[6] & b[3];
  assign f_u_dadda_cla32_and_5_4 = a[5] & b[4];
  assign f_u_dadda_cla32_and_4_5 = a[4] & b[5];
  assign f_u_dadda_cla32_fa20_xor0 = f_u_dadda_cla32_and_6_3 ^ f_u_dadda_cla32_and_5_4;
  assign f_u_dadda_cla32_fa20_and0 = f_u_dadda_cla32_and_6_3 & f_u_dadda_cla32_and_5_4;
  assign f_u_dadda_cla32_fa20_xor1 = f_u_dadda_cla32_fa20_xor0 ^ f_u_dadda_cla32_and_4_5;
  assign f_u_dadda_cla32_fa20_and1 = f_u_dadda_cla32_fa20_xor0 & f_u_dadda_cla32_and_4_5;
  assign f_u_dadda_cla32_fa20_or0 = f_u_dadda_cla32_fa20_and0 | f_u_dadda_cla32_fa20_and1;
  assign f_u_dadda_cla32_and_3_6 = a[3] & b[6];
  assign f_u_dadda_cla32_and_2_7 = a[2] & b[7];
  assign f_u_dadda_cla32_ha8_xor0 = f_u_dadda_cla32_and_3_6 ^ f_u_dadda_cla32_and_2_7;
  assign f_u_dadda_cla32_ha8_and0 = f_u_dadda_cla32_and_3_6 & f_u_dadda_cla32_and_2_7;
  assign f_u_dadda_cla32_fa21_xor0 = f_u_dadda_cla32_ha8_and0 ^ f_u_dadda_cla32_fa20_or0;
  assign f_u_dadda_cla32_fa21_and0 = f_u_dadda_cla32_ha8_and0 & f_u_dadda_cla32_fa20_or0;
  assign f_u_dadda_cla32_fa21_xor1 = f_u_dadda_cla32_fa21_xor0 ^ f_u_dadda_cla32_fa19_or0;
  assign f_u_dadda_cla32_fa21_and1 = f_u_dadda_cla32_fa21_xor0 & f_u_dadda_cla32_fa19_or0;
  assign f_u_dadda_cla32_fa21_or0 = f_u_dadda_cla32_fa21_and0 | f_u_dadda_cla32_fa21_and1;
  assign f_u_dadda_cla32_and_10_0 = a[10] & b[0];
  assign f_u_dadda_cla32_and_9_1 = a[9] & b[1];
  assign f_u_dadda_cla32_fa22_xor0 = f_u_dadda_cla32_fa18_or0 ^ f_u_dadda_cla32_and_10_0;
  assign f_u_dadda_cla32_fa22_and0 = f_u_dadda_cla32_fa18_or0 & f_u_dadda_cla32_and_10_0;
  assign f_u_dadda_cla32_fa22_xor1 = f_u_dadda_cla32_fa22_xor0 ^ f_u_dadda_cla32_and_9_1;
  assign f_u_dadda_cla32_fa22_and1 = f_u_dadda_cla32_fa22_xor0 & f_u_dadda_cla32_and_9_1;
  assign f_u_dadda_cla32_fa22_or0 = f_u_dadda_cla32_fa22_and0 | f_u_dadda_cla32_fa22_and1;
  assign f_u_dadda_cla32_and_8_2 = a[8] & b[2];
  assign f_u_dadda_cla32_and_7_3 = a[7] & b[3];
  assign f_u_dadda_cla32_and_6_4 = a[6] & b[4];
  assign f_u_dadda_cla32_fa23_xor0 = f_u_dadda_cla32_and_8_2 ^ f_u_dadda_cla32_and_7_3;
  assign f_u_dadda_cla32_fa23_and0 = f_u_dadda_cla32_and_8_2 & f_u_dadda_cla32_and_7_3;
  assign f_u_dadda_cla32_fa23_xor1 = f_u_dadda_cla32_fa23_xor0 ^ f_u_dadda_cla32_and_6_4;
  assign f_u_dadda_cla32_fa23_and1 = f_u_dadda_cla32_fa23_xor0 & f_u_dadda_cla32_and_6_4;
  assign f_u_dadda_cla32_fa23_or0 = f_u_dadda_cla32_fa23_and0 | f_u_dadda_cla32_fa23_and1;
  assign f_u_dadda_cla32_and_5_5 = a[5] & b[5];
  assign f_u_dadda_cla32_and_4_6 = a[4] & b[6];
  assign f_u_dadda_cla32_and_3_7 = a[3] & b[7];
  assign f_u_dadda_cla32_fa24_xor0 = f_u_dadda_cla32_and_5_5 ^ f_u_dadda_cla32_and_4_6;
  assign f_u_dadda_cla32_fa24_and0 = f_u_dadda_cla32_and_5_5 & f_u_dadda_cla32_and_4_6;
  assign f_u_dadda_cla32_fa24_xor1 = f_u_dadda_cla32_fa24_xor0 ^ f_u_dadda_cla32_and_3_7;
  assign f_u_dadda_cla32_fa24_and1 = f_u_dadda_cla32_fa24_xor0 & f_u_dadda_cla32_and_3_7;
  assign f_u_dadda_cla32_fa24_or0 = f_u_dadda_cla32_fa24_and0 | f_u_dadda_cla32_fa24_and1;
  assign f_u_dadda_cla32_and_2_8 = a[2] & b[8];
  assign f_u_dadda_cla32_and_1_9 = a[1] & b[9];
  assign f_u_dadda_cla32_ha9_xor0 = f_u_dadda_cla32_and_2_8 ^ f_u_dadda_cla32_and_1_9;
  assign f_u_dadda_cla32_ha9_and0 = f_u_dadda_cla32_and_2_8 & f_u_dadda_cla32_and_1_9;
  assign f_u_dadda_cla32_fa25_xor0 = f_u_dadda_cla32_ha9_and0 ^ f_u_dadda_cla32_fa24_or0;
  assign f_u_dadda_cla32_fa25_and0 = f_u_dadda_cla32_ha9_and0 & f_u_dadda_cla32_fa24_or0;
  assign f_u_dadda_cla32_fa25_xor1 = f_u_dadda_cla32_fa25_xor0 ^ f_u_dadda_cla32_fa23_or0;
  assign f_u_dadda_cla32_fa25_and1 = f_u_dadda_cla32_fa25_xor0 & f_u_dadda_cla32_fa23_or0;
  assign f_u_dadda_cla32_fa25_or0 = f_u_dadda_cla32_fa25_and0 | f_u_dadda_cla32_fa25_and1;
  assign f_u_dadda_cla32_and_11_0 = a[11] & b[0];
  assign f_u_dadda_cla32_fa26_xor0 = f_u_dadda_cla32_fa22_or0 ^ f_u_dadda_cla32_fa21_or0;
  assign f_u_dadda_cla32_fa26_and0 = f_u_dadda_cla32_fa22_or0 & f_u_dadda_cla32_fa21_or0;
  assign f_u_dadda_cla32_fa26_xor1 = f_u_dadda_cla32_fa26_xor0 ^ f_u_dadda_cla32_and_11_0;
  assign f_u_dadda_cla32_fa26_and1 = f_u_dadda_cla32_fa26_xor0 & f_u_dadda_cla32_and_11_0;
  assign f_u_dadda_cla32_fa26_or0 = f_u_dadda_cla32_fa26_and0 | f_u_dadda_cla32_fa26_and1;
  assign f_u_dadda_cla32_and_10_1 = a[10] & b[1];
  assign f_u_dadda_cla32_and_9_2 = a[9] & b[2];
  assign f_u_dadda_cla32_and_8_3 = a[8] & b[3];
  assign f_u_dadda_cla32_fa27_xor0 = f_u_dadda_cla32_and_10_1 ^ f_u_dadda_cla32_and_9_2;
  assign f_u_dadda_cla32_fa27_and0 = f_u_dadda_cla32_and_10_1 & f_u_dadda_cla32_and_9_2;
  assign f_u_dadda_cla32_fa27_xor1 = f_u_dadda_cla32_fa27_xor0 ^ f_u_dadda_cla32_and_8_3;
  assign f_u_dadda_cla32_fa27_and1 = f_u_dadda_cla32_fa27_xor0 & f_u_dadda_cla32_and_8_3;
  assign f_u_dadda_cla32_fa27_or0 = f_u_dadda_cla32_fa27_and0 | f_u_dadda_cla32_fa27_and1;
  assign f_u_dadda_cla32_and_7_4 = a[7] & b[4];
  assign f_u_dadda_cla32_and_6_5 = a[6] & b[5];
  assign f_u_dadda_cla32_and_5_6 = a[5] & b[6];
  assign f_u_dadda_cla32_fa28_xor0 = f_u_dadda_cla32_and_7_4 ^ f_u_dadda_cla32_and_6_5;
  assign f_u_dadda_cla32_fa28_and0 = f_u_dadda_cla32_and_7_4 & f_u_dadda_cla32_and_6_5;
  assign f_u_dadda_cla32_fa28_xor1 = f_u_dadda_cla32_fa28_xor0 ^ f_u_dadda_cla32_and_5_6;
  assign f_u_dadda_cla32_fa28_and1 = f_u_dadda_cla32_fa28_xor0 & f_u_dadda_cla32_and_5_6;
  assign f_u_dadda_cla32_fa28_or0 = f_u_dadda_cla32_fa28_and0 | f_u_dadda_cla32_fa28_and1;
  assign f_u_dadda_cla32_and_4_7 = a[4] & b[7];
  assign f_u_dadda_cla32_and_3_8 = a[3] & b[8];
  assign f_u_dadda_cla32_and_2_9 = a[2] & b[9];
  assign f_u_dadda_cla32_fa29_xor0 = f_u_dadda_cla32_and_4_7 ^ f_u_dadda_cla32_and_3_8;
  assign f_u_dadda_cla32_fa29_and0 = f_u_dadda_cla32_and_4_7 & f_u_dadda_cla32_and_3_8;
  assign f_u_dadda_cla32_fa29_xor1 = f_u_dadda_cla32_fa29_xor0 ^ f_u_dadda_cla32_and_2_9;
  assign f_u_dadda_cla32_fa29_and1 = f_u_dadda_cla32_fa29_xor0 & f_u_dadda_cla32_and_2_9;
  assign f_u_dadda_cla32_fa29_or0 = f_u_dadda_cla32_fa29_and0 | f_u_dadda_cla32_fa29_and1;
  assign f_u_dadda_cla32_and_1_10 = a[1] & b[10];
  assign f_u_dadda_cla32_and_0_11 = a[0] & b[11];
  assign f_u_dadda_cla32_ha10_xor0 = f_u_dadda_cla32_and_1_10 ^ f_u_dadda_cla32_and_0_11;
  assign f_u_dadda_cla32_ha10_and0 = f_u_dadda_cla32_and_1_10 & f_u_dadda_cla32_and_0_11;
  assign f_u_dadda_cla32_fa30_xor0 = f_u_dadda_cla32_ha10_and0 ^ f_u_dadda_cla32_fa29_or0;
  assign f_u_dadda_cla32_fa30_and0 = f_u_dadda_cla32_ha10_and0 & f_u_dadda_cla32_fa29_or0;
  assign f_u_dadda_cla32_fa30_xor1 = f_u_dadda_cla32_fa30_xor0 ^ f_u_dadda_cla32_fa28_or0;
  assign f_u_dadda_cla32_fa30_and1 = f_u_dadda_cla32_fa30_xor0 & f_u_dadda_cla32_fa28_or0;
  assign f_u_dadda_cla32_fa30_or0 = f_u_dadda_cla32_fa30_and0 | f_u_dadda_cla32_fa30_and1;
  assign f_u_dadda_cla32_fa31_xor0 = f_u_dadda_cla32_fa27_or0 ^ f_u_dadda_cla32_fa26_or0;
  assign f_u_dadda_cla32_fa31_and0 = f_u_dadda_cla32_fa27_or0 & f_u_dadda_cla32_fa26_or0;
  assign f_u_dadda_cla32_fa31_xor1 = f_u_dadda_cla32_fa31_xor0 ^ f_u_dadda_cla32_fa25_or0;
  assign f_u_dadda_cla32_fa31_and1 = f_u_dadda_cla32_fa31_xor0 & f_u_dadda_cla32_fa25_or0;
  assign f_u_dadda_cla32_fa31_or0 = f_u_dadda_cla32_fa31_and0 | f_u_dadda_cla32_fa31_and1;
  assign f_u_dadda_cla32_and_12_0 = a[12] & b[0];
  assign f_u_dadda_cla32_and_11_1 = a[11] & b[1];
  assign f_u_dadda_cla32_and_10_2 = a[10] & b[2];
  assign f_u_dadda_cla32_fa32_xor0 = f_u_dadda_cla32_and_12_0 ^ f_u_dadda_cla32_and_11_1;
  assign f_u_dadda_cla32_fa32_and0 = f_u_dadda_cla32_and_12_0 & f_u_dadda_cla32_and_11_1;
  assign f_u_dadda_cla32_fa32_xor1 = f_u_dadda_cla32_fa32_xor0 ^ f_u_dadda_cla32_and_10_2;
  assign f_u_dadda_cla32_fa32_and1 = f_u_dadda_cla32_fa32_xor0 & f_u_dadda_cla32_and_10_2;
  assign f_u_dadda_cla32_fa32_or0 = f_u_dadda_cla32_fa32_and0 | f_u_dadda_cla32_fa32_and1;
  assign f_u_dadda_cla32_and_9_3 = a[9] & b[3];
  assign f_u_dadda_cla32_and_8_4 = a[8] & b[4];
  assign f_u_dadda_cla32_and_7_5 = a[7] & b[5];
  assign f_u_dadda_cla32_fa33_xor0 = f_u_dadda_cla32_and_9_3 ^ f_u_dadda_cla32_and_8_4;
  assign f_u_dadda_cla32_fa33_and0 = f_u_dadda_cla32_and_9_3 & f_u_dadda_cla32_and_8_4;
  assign f_u_dadda_cla32_fa33_xor1 = f_u_dadda_cla32_fa33_xor0 ^ f_u_dadda_cla32_and_7_5;
  assign f_u_dadda_cla32_fa33_and1 = f_u_dadda_cla32_fa33_xor0 & f_u_dadda_cla32_and_7_5;
  assign f_u_dadda_cla32_fa33_or0 = f_u_dadda_cla32_fa33_and0 | f_u_dadda_cla32_fa33_and1;
  assign f_u_dadda_cla32_and_6_6 = a[6] & b[6];
  assign f_u_dadda_cla32_and_5_7 = a[5] & b[7];
  assign f_u_dadda_cla32_and_4_8 = a[4] & b[8];
  assign f_u_dadda_cla32_fa34_xor0 = f_u_dadda_cla32_and_6_6 ^ f_u_dadda_cla32_and_5_7;
  assign f_u_dadda_cla32_fa34_and0 = f_u_dadda_cla32_and_6_6 & f_u_dadda_cla32_and_5_7;
  assign f_u_dadda_cla32_fa34_xor1 = f_u_dadda_cla32_fa34_xor0 ^ f_u_dadda_cla32_and_4_8;
  assign f_u_dadda_cla32_fa34_and1 = f_u_dadda_cla32_fa34_xor0 & f_u_dadda_cla32_and_4_8;
  assign f_u_dadda_cla32_fa34_or0 = f_u_dadda_cla32_fa34_and0 | f_u_dadda_cla32_fa34_and1;
  assign f_u_dadda_cla32_and_3_9 = a[3] & b[9];
  assign f_u_dadda_cla32_and_2_10 = a[2] & b[10];
  assign f_u_dadda_cla32_and_1_11 = a[1] & b[11];
  assign f_u_dadda_cla32_fa35_xor0 = f_u_dadda_cla32_and_3_9 ^ f_u_dadda_cla32_and_2_10;
  assign f_u_dadda_cla32_fa35_and0 = f_u_dadda_cla32_and_3_9 & f_u_dadda_cla32_and_2_10;
  assign f_u_dadda_cla32_fa35_xor1 = f_u_dadda_cla32_fa35_xor0 ^ f_u_dadda_cla32_and_1_11;
  assign f_u_dadda_cla32_fa35_and1 = f_u_dadda_cla32_fa35_xor0 & f_u_dadda_cla32_and_1_11;
  assign f_u_dadda_cla32_fa35_or0 = f_u_dadda_cla32_fa35_and0 | f_u_dadda_cla32_fa35_and1;
  assign f_u_dadda_cla32_and_0_12 = a[0] & b[12];
  assign f_u_dadda_cla32_ha11_xor0 = f_u_dadda_cla32_and_0_12 ^ f_u_dadda_cla32_fa30_xor1;
  assign f_u_dadda_cla32_ha11_and0 = f_u_dadda_cla32_and_0_12 & f_u_dadda_cla32_fa30_xor1;
  assign f_u_dadda_cla32_fa36_xor0 = f_u_dadda_cla32_ha11_and0 ^ f_u_dadda_cla32_fa35_or0;
  assign f_u_dadda_cla32_fa36_and0 = f_u_dadda_cla32_ha11_and0 & f_u_dadda_cla32_fa35_or0;
  assign f_u_dadda_cla32_fa36_xor1 = f_u_dadda_cla32_fa36_xor0 ^ f_u_dadda_cla32_fa34_or0;
  assign f_u_dadda_cla32_fa36_and1 = f_u_dadda_cla32_fa36_xor0 & f_u_dadda_cla32_fa34_or0;
  assign f_u_dadda_cla32_fa36_or0 = f_u_dadda_cla32_fa36_and0 | f_u_dadda_cla32_fa36_and1;
  assign f_u_dadda_cla32_fa37_xor0 = f_u_dadda_cla32_fa33_or0 ^ f_u_dadda_cla32_fa32_or0;
  assign f_u_dadda_cla32_fa37_and0 = f_u_dadda_cla32_fa33_or0 & f_u_dadda_cla32_fa32_or0;
  assign f_u_dadda_cla32_fa37_xor1 = f_u_dadda_cla32_fa37_xor0 ^ f_u_dadda_cla32_fa31_or0;
  assign f_u_dadda_cla32_fa37_and1 = f_u_dadda_cla32_fa37_xor0 & f_u_dadda_cla32_fa31_or0;
  assign f_u_dadda_cla32_fa37_or0 = f_u_dadda_cla32_fa37_and0 | f_u_dadda_cla32_fa37_and1;
  assign f_u_dadda_cla32_and_13_0 = a[13] & b[0];
  assign f_u_dadda_cla32_and_12_1 = a[12] & b[1];
  assign f_u_dadda_cla32_fa38_xor0 = f_u_dadda_cla32_fa30_or0 ^ f_u_dadda_cla32_and_13_0;
  assign f_u_dadda_cla32_fa38_and0 = f_u_dadda_cla32_fa30_or0 & f_u_dadda_cla32_and_13_0;
  assign f_u_dadda_cla32_fa38_xor1 = f_u_dadda_cla32_fa38_xor0 ^ f_u_dadda_cla32_and_12_1;
  assign f_u_dadda_cla32_fa38_and1 = f_u_dadda_cla32_fa38_xor0 & f_u_dadda_cla32_and_12_1;
  assign f_u_dadda_cla32_fa38_or0 = f_u_dadda_cla32_fa38_and0 | f_u_dadda_cla32_fa38_and1;
  assign f_u_dadda_cla32_and_11_2 = a[11] & b[2];
  assign f_u_dadda_cla32_and_10_3 = a[10] & b[3];
  assign f_u_dadda_cla32_and_9_4 = a[9] & b[4];
  assign f_u_dadda_cla32_fa39_xor0 = f_u_dadda_cla32_and_11_2 ^ f_u_dadda_cla32_and_10_3;
  assign f_u_dadda_cla32_fa39_and0 = f_u_dadda_cla32_and_11_2 & f_u_dadda_cla32_and_10_3;
  assign f_u_dadda_cla32_fa39_xor1 = f_u_dadda_cla32_fa39_xor0 ^ f_u_dadda_cla32_and_9_4;
  assign f_u_dadda_cla32_fa39_and1 = f_u_dadda_cla32_fa39_xor0 & f_u_dadda_cla32_and_9_4;
  assign f_u_dadda_cla32_fa39_or0 = f_u_dadda_cla32_fa39_and0 | f_u_dadda_cla32_fa39_and1;
  assign f_u_dadda_cla32_and_8_5 = a[8] & b[5];
  assign f_u_dadda_cla32_and_7_6 = a[7] & b[6];
  assign f_u_dadda_cla32_and_6_7 = a[6] & b[7];
  assign f_u_dadda_cla32_fa40_xor0 = f_u_dadda_cla32_and_8_5 ^ f_u_dadda_cla32_and_7_6;
  assign f_u_dadda_cla32_fa40_and0 = f_u_dadda_cla32_and_8_5 & f_u_dadda_cla32_and_7_6;
  assign f_u_dadda_cla32_fa40_xor1 = f_u_dadda_cla32_fa40_xor0 ^ f_u_dadda_cla32_and_6_7;
  assign f_u_dadda_cla32_fa40_and1 = f_u_dadda_cla32_fa40_xor0 & f_u_dadda_cla32_and_6_7;
  assign f_u_dadda_cla32_fa40_or0 = f_u_dadda_cla32_fa40_and0 | f_u_dadda_cla32_fa40_and1;
  assign f_u_dadda_cla32_and_5_8 = a[5] & b[8];
  assign f_u_dadda_cla32_and_4_9 = a[4] & b[9];
  assign f_u_dadda_cla32_and_3_10 = a[3] & b[10];
  assign f_u_dadda_cla32_fa41_xor0 = f_u_dadda_cla32_and_5_8 ^ f_u_dadda_cla32_and_4_9;
  assign f_u_dadda_cla32_fa41_and0 = f_u_dadda_cla32_and_5_8 & f_u_dadda_cla32_and_4_9;
  assign f_u_dadda_cla32_fa41_xor1 = f_u_dadda_cla32_fa41_xor0 ^ f_u_dadda_cla32_and_3_10;
  assign f_u_dadda_cla32_fa41_and1 = f_u_dadda_cla32_fa41_xor0 & f_u_dadda_cla32_and_3_10;
  assign f_u_dadda_cla32_fa41_or0 = f_u_dadda_cla32_fa41_and0 | f_u_dadda_cla32_fa41_and1;
  assign f_u_dadda_cla32_and_2_11 = a[2] & b[11];
  assign f_u_dadda_cla32_and_1_12 = a[1] & b[12];
  assign f_u_dadda_cla32_and_0_13 = a[0] & b[13];
  assign f_u_dadda_cla32_fa42_xor0 = f_u_dadda_cla32_and_2_11 ^ f_u_dadda_cla32_and_1_12;
  assign f_u_dadda_cla32_fa42_and0 = f_u_dadda_cla32_and_2_11 & f_u_dadda_cla32_and_1_12;
  assign f_u_dadda_cla32_fa42_xor1 = f_u_dadda_cla32_fa42_xor0 ^ f_u_dadda_cla32_and_0_13;
  assign f_u_dadda_cla32_fa42_and1 = f_u_dadda_cla32_fa42_xor0 & f_u_dadda_cla32_and_0_13;
  assign f_u_dadda_cla32_fa42_or0 = f_u_dadda_cla32_fa42_and0 | f_u_dadda_cla32_fa42_and1;
  assign f_u_dadda_cla32_ha12_xor0 = f_u_dadda_cla32_fa36_xor1 ^ f_u_dadda_cla32_fa37_xor1;
  assign f_u_dadda_cla32_ha12_and0 = f_u_dadda_cla32_fa36_xor1 & f_u_dadda_cla32_fa37_xor1;
  assign f_u_dadda_cla32_fa43_xor0 = f_u_dadda_cla32_ha12_and0 ^ f_u_dadda_cla32_fa42_or0;
  assign f_u_dadda_cla32_fa43_and0 = f_u_dadda_cla32_ha12_and0 & f_u_dadda_cla32_fa42_or0;
  assign f_u_dadda_cla32_fa43_xor1 = f_u_dadda_cla32_fa43_xor0 ^ f_u_dadda_cla32_fa41_or0;
  assign f_u_dadda_cla32_fa43_and1 = f_u_dadda_cla32_fa43_xor0 & f_u_dadda_cla32_fa41_or0;
  assign f_u_dadda_cla32_fa43_or0 = f_u_dadda_cla32_fa43_and0 | f_u_dadda_cla32_fa43_and1;
  assign f_u_dadda_cla32_fa44_xor0 = f_u_dadda_cla32_fa40_or0 ^ f_u_dadda_cla32_fa39_or0;
  assign f_u_dadda_cla32_fa44_and0 = f_u_dadda_cla32_fa40_or0 & f_u_dadda_cla32_fa39_or0;
  assign f_u_dadda_cla32_fa44_xor1 = f_u_dadda_cla32_fa44_xor0 ^ f_u_dadda_cla32_fa38_or0;
  assign f_u_dadda_cla32_fa44_and1 = f_u_dadda_cla32_fa44_xor0 & f_u_dadda_cla32_fa38_or0;
  assign f_u_dadda_cla32_fa44_or0 = f_u_dadda_cla32_fa44_and0 | f_u_dadda_cla32_fa44_and1;
  assign f_u_dadda_cla32_and_14_0 = a[14] & b[0];
  assign f_u_dadda_cla32_fa45_xor0 = f_u_dadda_cla32_fa37_or0 ^ f_u_dadda_cla32_fa36_or0;
  assign f_u_dadda_cla32_fa45_and0 = f_u_dadda_cla32_fa37_or0 & f_u_dadda_cla32_fa36_or0;
  assign f_u_dadda_cla32_fa45_xor1 = f_u_dadda_cla32_fa45_xor0 ^ f_u_dadda_cla32_and_14_0;
  assign f_u_dadda_cla32_fa45_and1 = f_u_dadda_cla32_fa45_xor0 & f_u_dadda_cla32_and_14_0;
  assign f_u_dadda_cla32_fa45_or0 = f_u_dadda_cla32_fa45_and0 | f_u_dadda_cla32_fa45_and1;
  assign f_u_dadda_cla32_and_13_1 = a[13] & b[1];
  assign f_u_dadda_cla32_and_12_2 = a[12] & b[2];
  assign f_u_dadda_cla32_and_11_3 = a[11] & b[3];
  assign f_u_dadda_cla32_fa46_xor0 = f_u_dadda_cla32_and_13_1 ^ f_u_dadda_cla32_and_12_2;
  assign f_u_dadda_cla32_fa46_and0 = f_u_dadda_cla32_and_13_1 & f_u_dadda_cla32_and_12_2;
  assign f_u_dadda_cla32_fa46_xor1 = f_u_dadda_cla32_fa46_xor0 ^ f_u_dadda_cla32_and_11_3;
  assign f_u_dadda_cla32_fa46_and1 = f_u_dadda_cla32_fa46_xor0 & f_u_dadda_cla32_and_11_3;
  assign f_u_dadda_cla32_fa46_or0 = f_u_dadda_cla32_fa46_and0 | f_u_dadda_cla32_fa46_and1;
  assign f_u_dadda_cla32_and_10_4 = a[10] & b[4];
  assign f_u_dadda_cla32_and_9_5 = a[9] & b[5];
  assign f_u_dadda_cla32_and_8_6 = a[8] & b[6];
  assign f_u_dadda_cla32_fa47_xor0 = f_u_dadda_cla32_and_10_4 ^ f_u_dadda_cla32_and_9_5;
  assign f_u_dadda_cla32_fa47_and0 = f_u_dadda_cla32_and_10_4 & f_u_dadda_cla32_and_9_5;
  assign f_u_dadda_cla32_fa47_xor1 = f_u_dadda_cla32_fa47_xor0 ^ f_u_dadda_cla32_and_8_6;
  assign f_u_dadda_cla32_fa47_and1 = f_u_dadda_cla32_fa47_xor0 & f_u_dadda_cla32_and_8_6;
  assign f_u_dadda_cla32_fa47_or0 = f_u_dadda_cla32_fa47_and0 | f_u_dadda_cla32_fa47_and1;
  assign f_u_dadda_cla32_and_7_7 = a[7] & b[7];
  assign f_u_dadda_cla32_and_6_8 = a[6] & b[8];
  assign f_u_dadda_cla32_and_5_9 = a[5] & b[9];
  assign f_u_dadda_cla32_fa48_xor0 = f_u_dadda_cla32_and_7_7 ^ f_u_dadda_cla32_and_6_8;
  assign f_u_dadda_cla32_fa48_and0 = f_u_dadda_cla32_and_7_7 & f_u_dadda_cla32_and_6_8;
  assign f_u_dadda_cla32_fa48_xor1 = f_u_dadda_cla32_fa48_xor0 ^ f_u_dadda_cla32_and_5_9;
  assign f_u_dadda_cla32_fa48_and1 = f_u_dadda_cla32_fa48_xor0 & f_u_dadda_cla32_and_5_9;
  assign f_u_dadda_cla32_fa48_or0 = f_u_dadda_cla32_fa48_and0 | f_u_dadda_cla32_fa48_and1;
  assign f_u_dadda_cla32_and_4_10 = a[4] & b[10];
  assign f_u_dadda_cla32_and_3_11 = a[3] & b[11];
  assign f_u_dadda_cla32_and_2_12 = a[2] & b[12];
  assign f_u_dadda_cla32_fa49_xor0 = f_u_dadda_cla32_and_4_10 ^ f_u_dadda_cla32_and_3_11;
  assign f_u_dadda_cla32_fa49_and0 = f_u_dadda_cla32_and_4_10 & f_u_dadda_cla32_and_3_11;
  assign f_u_dadda_cla32_fa49_xor1 = f_u_dadda_cla32_fa49_xor0 ^ f_u_dadda_cla32_and_2_12;
  assign f_u_dadda_cla32_fa49_and1 = f_u_dadda_cla32_fa49_xor0 & f_u_dadda_cla32_and_2_12;
  assign f_u_dadda_cla32_fa49_or0 = f_u_dadda_cla32_fa49_and0 | f_u_dadda_cla32_fa49_and1;
  assign f_u_dadda_cla32_and_1_13 = a[1] & b[13];
  assign f_u_dadda_cla32_and_0_14 = a[0] & b[14];
  assign f_u_dadda_cla32_fa50_xor0 = f_u_dadda_cla32_and_1_13 ^ f_u_dadda_cla32_and_0_14;
  assign f_u_dadda_cla32_fa50_and0 = f_u_dadda_cla32_and_1_13 & f_u_dadda_cla32_and_0_14;
  assign f_u_dadda_cla32_fa50_xor1 = f_u_dadda_cla32_fa50_xor0 ^ f_u_dadda_cla32_fa43_xor1;
  assign f_u_dadda_cla32_fa50_and1 = f_u_dadda_cla32_fa50_xor0 & f_u_dadda_cla32_fa43_xor1;
  assign f_u_dadda_cla32_fa50_or0 = f_u_dadda_cla32_fa50_and0 | f_u_dadda_cla32_fa50_and1;
  assign f_u_dadda_cla32_ha13_xor0 = f_u_dadda_cla32_fa44_xor1 ^ f_u_dadda_cla32_fa45_xor1;
  assign f_u_dadda_cla32_ha13_and0 = f_u_dadda_cla32_fa44_xor1 & f_u_dadda_cla32_fa45_xor1;
  assign f_u_dadda_cla32_fa51_xor0 = f_u_dadda_cla32_ha13_and0 ^ f_u_dadda_cla32_fa50_or0;
  assign f_u_dadda_cla32_fa51_and0 = f_u_dadda_cla32_ha13_and0 & f_u_dadda_cla32_fa50_or0;
  assign f_u_dadda_cla32_fa51_xor1 = f_u_dadda_cla32_fa51_xor0 ^ f_u_dadda_cla32_fa49_or0;
  assign f_u_dadda_cla32_fa51_and1 = f_u_dadda_cla32_fa51_xor0 & f_u_dadda_cla32_fa49_or0;
  assign f_u_dadda_cla32_fa51_or0 = f_u_dadda_cla32_fa51_and0 | f_u_dadda_cla32_fa51_and1;
  assign f_u_dadda_cla32_fa52_xor0 = f_u_dadda_cla32_fa48_or0 ^ f_u_dadda_cla32_fa47_or0;
  assign f_u_dadda_cla32_fa52_and0 = f_u_dadda_cla32_fa48_or0 & f_u_dadda_cla32_fa47_or0;
  assign f_u_dadda_cla32_fa52_xor1 = f_u_dadda_cla32_fa52_xor0 ^ f_u_dadda_cla32_fa46_or0;
  assign f_u_dadda_cla32_fa52_and1 = f_u_dadda_cla32_fa52_xor0 & f_u_dadda_cla32_fa46_or0;
  assign f_u_dadda_cla32_fa52_or0 = f_u_dadda_cla32_fa52_and0 | f_u_dadda_cla32_fa52_and1;
  assign f_u_dadda_cla32_fa53_xor0 = f_u_dadda_cla32_fa45_or0 ^ f_u_dadda_cla32_fa44_or0;
  assign f_u_dadda_cla32_fa53_and0 = f_u_dadda_cla32_fa45_or0 & f_u_dadda_cla32_fa44_or0;
  assign f_u_dadda_cla32_fa53_xor1 = f_u_dadda_cla32_fa53_xor0 ^ f_u_dadda_cla32_fa43_or0;
  assign f_u_dadda_cla32_fa53_and1 = f_u_dadda_cla32_fa53_xor0 & f_u_dadda_cla32_fa43_or0;
  assign f_u_dadda_cla32_fa53_or0 = f_u_dadda_cla32_fa53_and0 | f_u_dadda_cla32_fa53_and1;
  assign f_u_dadda_cla32_and_15_0 = a[15] & b[0];
  assign f_u_dadda_cla32_and_14_1 = a[14] & b[1];
  assign f_u_dadda_cla32_and_13_2 = a[13] & b[2];
  assign f_u_dadda_cla32_fa54_xor0 = f_u_dadda_cla32_and_15_0 ^ f_u_dadda_cla32_and_14_1;
  assign f_u_dadda_cla32_fa54_and0 = f_u_dadda_cla32_and_15_0 & f_u_dadda_cla32_and_14_1;
  assign f_u_dadda_cla32_fa54_xor1 = f_u_dadda_cla32_fa54_xor0 ^ f_u_dadda_cla32_and_13_2;
  assign f_u_dadda_cla32_fa54_and1 = f_u_dadda_cla32_fa54_xor0 & f_u_dadda_cla32_and_13_2;
  assign f_u_dadda_cla32_fa54_or0 = f_u_dadda_cla32_fa54_and0 | f_u_dadda_cla32_fa54_and1;
  assign f_u_dadda_cla32_and_12_3 = a[12] & b[3];
  assign f_u_dadda_cla32_and_11_4 = a[11] & b[4];
  assign f_u_dadda_cla32_and_10_5 = a[10] & b[5];
  assign f_u_dadda_cla32_fa55_xor0 = f_u_dadda_cla32_and_12_3 ^ f_u_dadda_cla32_and_11_4;
  assign f_u_dadda_cla32_fa55_and0 = f_u_dadda_cla32_and_12_3 & f_u_dadda_cla32_and_11_4;
  assign f_u_dadda_cla32_fa55_xor1 = f_u_dadda_cla32_fa55_xor0 ^ f_u_dadda_cla32_and_10_5;
  assign f_u_dadda_cla32_fa55_and1 = f_u_dadda_cla32_fa55_xor0 & f_u_dadda_cla32_and_10_5;
  assign f_u_dadda_cla32_fa55_or0 = f_u_dadda_cla32_fa55_and0 | f_u_dadda_cla32_fa55_and1;
  assign f_u_dadda_cla32_and_9_6 = a[9] & b[6];
  assign f_u_dadda_cla32_and_8_7 = a[8] & b[7];
  assign f_u_dadda_cla32_and_7_8 = a[7] & b[8];
  assign f_u_dadda_cla32_fa56_xor0 = f_u_dadda_cla32_and_9_6 ^ f_u_dadda_cla32_and_8_7;
  assign f_u_dadda_cla32_fa56_and0 = f_u_dadda_cla32_and_9_6 & f_u_dadda_cla32_and_8_7;
  assign f_u_dadda_cla32_fa56_xor1 = f_u_dadda_cla32_fa56_xor0 ^ f_u_dadda_cla32_and_7_8;
  assign f_u_dadda_cla32_fa56_and1 = f_u_dadda_cla32_fa56_xor0 & f_u_dadda_cla32_and_7_8;
  assign f_u_dadda_cla32_fa56_or0 = f_u_dadda_cla32_fa56_and0 | f_u_dadda_cla32_fa56_and1;
  assign f_u_dadda_cla32_and_6_9 = a[6] & b[9];
  assign f_u_dadda_cla32_and_5_10 = a[5] & b[10];
  assign f_u_dadda_cla32_and_4_11 = a[4] & b[11];
  assign f_u_dadda_cla32_fa57_xor0 = f_u_dadda_cla32_and_6_9 ^ f_u_dadda_cla32_and_5_10;
  assign f_u_dadda_cla32_fa57_and0 = f_u_dadda_cla32_and_6_9 & f_u_dadda_cla32_and_5_10;
  assign f_u_dadda_cla32_fa57_xor1 = f_u_dadda_cla32_fa57_xor0 ^ f_u_dadda_cla32_and_4_11;
  assign f_u_dadda_cla32_fa57_and1 = f_u_dadda_cla32_fa57_xor0 & f_u_dadda_cla32_and_4_11;
  assign f_u_dadda_cla32_fa57_or0 = f_u_dadda_cla32_fa57_and0 | f_u_dadda_cla32_fa57_and1;
  assign f_u_dadda_cla32_and_3_12 = a[3] & b[12];
  assign f_u_dadda_cla32_and_2_13 = a[2] & b[13];
  assign f_u_dadda_cla32_and_1_14 = a[1] & b[14];
  assign f_u_dadda_cla32_fa58_xor0 = f_u_dadda_cla32_and_3_12 ^ f_u_dadda_cla32_and_2_13;
  assign f_u_dadda_cla32_fa58_and0 = f_u_dadda_cla32_and_3_12 & f_u_dadda_cla32_and_2_13;
  assign f_u_dadda_cla32_fa58_xor1 = f_u_dadda_cla32_fa58_xor0 ^ f_u_dadda_cla32_and_1_14;
  assign f_u_dadda_cla32_fa58_and1 = f_u_dadda_cla32_fa58_xor0 & f_u_dadda_cla32_and_1_14;
  assign f_u_dadda_cla32_fa58_or0 = f_u_dadda_cla32_fa58_and0 | f_u_dadda_cla32_fa58_and1;
  assign f_u_dadda_cla32_and_0_15 = a[0] & b[15];
  assign f_u_dadda_cla32_fa59_xor0 = f_u_dadda_cla32_and_0_15 ^ f_u_dadda_cla32_fa51_xor1;
  assign f_u_dadda_cla32_fa59_and0 = f_u_dadda_cla32_and_0_15 & f_u_dadda_cla32_fa51_xor1;
  assign f_u_dadda_cla32_fa59_xor1 = f_u_dadda_cla32_fa59_xor0 ^ f_u_dadda_cla32_fa52_xor1;
  assign f_u_dadda_cla32_fa59_and1 = f_u_dadda_cla32_fa59_xor0 & f_u_dadda_cla32_fa52_xor1;
  assign f_u_dadda_cla32_fa59_or0 = f_u_dadda_cla32_fa59_and0 | f_u_dadda_cla32_fa59_and1;
  assign f_u_dadda_cla32_ha14_xor0 = f_u_dadda_cla32_fa53_xor1 ^ f_u_dadda_cla32_fa54_xor1;
  assign f_u_dadda_cla32_ha14_and0 = f_u_dadda_cla32_fa53_xor1 & f_u_dadda_cla32_fa54_xor1;
  assign f_u_dadda_cla32_fa60_xor0 = f_u_dadda_cla32_ha14_and0 ^ f_u_dadda_cla32_fa59_or0;
  assign f_u_dadda_cla32_fa60_and0 = f_u_dadda_cla32_ha14_and0 & f_u_dadda_cla32_fa59_or0;
  assign f_u_dadda_cla32_fa60_xor1 = f_u_dadda_cla32_fa60_xor0 ^ f_u_dadda_cla32_fa58_or0;
  assign f_u_dadda_cla32_fa60_and1 = f_u_dadda_cla32_fa60_xor0 & f_u_dadda_cla32_fa58_or0;
  assign f_u_dadda_cla32_fa60_or0 = f_u_dadda_cla32_fa60_and0 | f_u_dadda_cla32_fa60_and1;
  assign f_u_dadda_cla32_fa61_xor0 = f_u_dadda_cla32_fa57_or0 ^ f_u_dadda_cla32_fa56_or0;
  assign f_u_dadda_cla32_fa61_and0 = f_u_dadda_cla32_fa57_or0 & f_u_dadda_cla32_fa56_or0;
  assign f_u_dadda_cla32_fa61_xor1 = f_u_dadda_cla32_fa61_xor0 ^ f_u_dadda_cla32_fa55_or0;
  assign f_u_dadda_cla32_fa61_and1 = f_u_dadda_cla32_fa61_xor0 & f_u_dadda_cla32_fa55_or0;
  assign f_u_dadda_cla32_fa61_or0 = f_u_dadda_cla32_fa61_and0 | f_u_dadda_cla32_fa61_and1;
  assign f_u_dadda_cla32_fa62_xor0 = f_u_dadda_cla32_fa54_or0 ^ f_u_dadda_cla32_fa53_or0;
  assign f_u_dadda_cla32_fa62_and0 = f_u_dadda_cla32_fa54_or0 & f_u_dadda_cla32_fa53_or0;
  assign f_u_dadda_cla32_fa62_xor1 = f_u_dadda_cla32_fa62_xor0 ^ f_u_dadda_cla32_fa52_or0;
  assign f_u_dadda_cla32_fa62_and1 = f_u_dadda_cla32_fa62_xor0 & f_u_dadda_cla32_fa52_or0;
  assign f_u_dadda_cla32_fa62_or0 = f_u_dadda_cla32_fa62_and0 | f_u_dadda_cla32_fa62_and1;
  assign f_u_dadda_cla32_and_16_0 = a[16] & b[0];
  assign f_u_dadda_cla32_and_15_1 = a[15] & b[1];
  assign f_u_dadda_cla32_fa63_xor0 = f_u_dadda_cla32_fa51_or0 ^ f_u_dadda_cla32_and_16_0;
  assign f_u_dadda_cla32_fa63_and0 = f_u_dadda_cla32_fa51_or0 & f_u_dadda_cla32_and_16_0;
  assign f_u_dadda_cla32_fa63_xor1 = f_u_dadda_cla32_fa63_xor0 ^ f_u_dadda_cla32_and_15_1;
  assign f_u_dadda_cla32_fa63_and1 = f_u_dadda_cla32_fa63_xor0 & f_u_dadda_cla32_and_15_1;
  assign f_u_dadda_cla32_fa63_or0 = f_u_dadda_cla32_fa63_and0 | f_u_dadda_cla32_fa63_and1;
  assign f_u_dadda_cla32_and_14_2 = a[14] & b[2];
  assign f_u_dadda_cla32_and_13_3 = a[13] & b[3];
  assign f_u_dadda_cla32_and_12_4 = a[12] & b[4];
  assign f_u_dadda_cla32_fa64_xor0 = f_u_dadda_cla32_and_14_2 ^ f_u_dadda_cla32_and_13_3;
  assign f_u_dadda_cla32_fa64_and0 = f_u_dadda_cla32_and_14_2 & f_u_dadda_cla32_and_13_3;
  assign f_u_dadda_cla32_fa64_xor1 = f_u_dadda_cla32_fa64_xor0 ^ f_u_dadda_cla32_and_12_4;
  assign f_u_dadda_cla32_fa64_and1 = f_u_dadda_cla32_fa64_xor0 & f_u_dadda_cla32_and_12_4;
  assign f_u_dadda_cla32_fa64_or0 = f_u_dadda_cla32_fa64_and0 | f_u_dadda_cla32_fa64_and1;
  assign f_u_dadda_cla32_and_11_5 = a[11] & b[5];
  assign f_u_dadda_cla32_and_10_6 = a[10] & b[6];
  assign f_u_dadda_cla32_and_9_7 = a[9] & b[7];
  assign f_u_dadda_cla32_fa65_xor0 = f_u_dadda_cla32_and_11_5 ^ f_u_dadda_cla32_and_10_6;
  assign f_u_dadda_cla32_fa65_and0 = f_u_dadda_cla32_and_11_5 & f_u_dadda_cla32_and_10_6;
  assign f_u_dadda_cla32_fa65_xor1 = f_u_dadda_cla32_fa65_xor0 ^ f_u_dadda_cla32_and_9_7;
  assign f_u_dadda_cla32_fa65_and1 = f_u_dadda_cla32_fa65_xor0 & f_u_dadda_cla32_and_9_7;
  assign f_u_dadda_cla32_fa65_or0 = f_u_dadda_cla32_fa65_and0 | f_u_dadda_cla32_fa65_and1;
  assign f_u_dadda_cla32_and_8_8 = a[8] & b[8];
  assign f_u_dadda_cla32_and_7_9 = a[7] & b[9];
  assign f_u_dadda_cla32_and_6_10 = a[6] & b[10];
  assign f_u_dadda_cla32_fa66_xor0 = f_u_dadda_cla32_and_8_8 ^ f_u_dadda_cla32_and_7_9;
  assign f_u_dadda_cla32_fa66_and0 = f_u_dadda_cla32_and_8_8 & f_u_dadda_cla32_and_7_9;
  assign f_u_dadda_cla32_fa66_xor1 = f_u_dadda_cla32_fa66_xor0 ^ f_u_dadda_cla32_and_6_10;
  assign f_u_dadda_cla32_fa66_and1 = f_u_dadda_cla32_fa66_xor0 & f_u_dadda_cla32_and_6_10;
  assign f_u_dadda_cla32_fa66_or0 = f_u_dadda_cla32_fa66_and0 | f_u_dadda_cla32_fa66_and1;
  assign f_u_dadda_cla32_and_5_11 = a[5] & b[11];
  assign f_u_dadda_cla32_and_4_12 = a[4] & b[12];
  assign f_u_dadda_cla32_and_3_13 = a[3] & b[13];
  assign f_u_dadda_cla32_fa67_xor0 = f_u_dadda_cla32_and_5_11 ^ f_u_dadda_cla32_and_4_12;
  assign f_u_dadda_cla32_fa67_and0 = f_u_dadda_cla32_and_5_11 & f_u_dadda_cla32_and_4_12;
  assign f_u_dadda_cla32_fa67_xor1 = f_u_dadda_cla32_fa67_xor0 ^ f_u_dadda_cla32_and_3_13;
  assign f_u_dadda_cla32_fa67_and1 = f_u_dadda_cla32_fa67_xor0 & f_u_dadda_cla32_and_3_13;
  assign f_u_dadda_cla32_fa67_or0 = f_u_dadda_cla32_fa67_and0 | f_u_dadda_cla32_fa67_and1;
  assign f_u_dadda_cla32_and_2_14 = a[2] & b[14];
  assign f_u_dadda_cla32_and_1_15 = a[1] & b[15];
  assign f_u_dadda_cla32_and_0_16 = a[0] & b[16];
  assign f_u_dadda_cla32_fa68_xor0 = f_u_dadda_cla32_and_2_14 ^ f_u_dadda_cla32_and_1_15;
  assign f_u_dadda_cla32_fa68_and0 = f_u_dadda_cla32_and_2_14 & f_u_dadda_cla32_and_1_15;
  assign f_u_dadda_cla32_fa68_xor1 = f_u_dadda_cla32_fa68_xor0 ^ f_u_dadda_cla32_and_0_16;
  assign f_u_dadda_cla32_fa68_and1 = f_u_dadda_cla32_fa68_xor0 & f_u_dadda_cla32_and_0_16;
  assign f_u_dadda_cla32_fa68_or0 = f_u_dadda_cla32_fa68_and0 | f_u_dadda_cla32_fa68_and1;
  assign f_u_dadda_cla32_fa69_xor0 = f_u_dadda_cla32_fa60_xor1 ^ f_u_dadda_cla32_fa61_xor1;
  assign f_u_dadda_cla32_fa69_and0 = f_u_dadda_cla32_fa60_xor1 & f_u_dadda_cla32_fa61_xor1;
  assign f_u_dadda_cla32_fa69_xor1 = f_u_dadda_cla32_fa69_xor0 ^ f_u_dadda_cla32_fa62_xor1;
  assign f_u_dadda_cla32_fa69_and1 = f_u_dadda_cla32_fa69_xor0 & f_u_dadda_cla32_fa62_xor1;
  assign f_u_dadda_cla32_fa69_or0 = f_u_dadda_cla32_fa69_and0 | f_u_dadda_cla32_fa69_and1;
  assign f_u_dadda_cla32_ha15_xor0 = f_u_dadda_cla32_fa63_xor1 ^ f_u_dadda_cla32_fa64_xor1;
  assign f_u_dadda_cla32_ha15_and0 = f_u_dadda_cla32_fa63_xor1 & f_u_dadda_cla32_fa64_xor1;
  assign f_u_dadda_cla32_fa70_xor0 = f_u_dadda_cla32_ha15_and0 ^ f_u_dadda_cla32_fa69_or0;
  assign f_u_dadda_cla32_fa70_and0 = f_u_dadda_cla32_ha15_and0 & f_u_dadda_cla32_fa69_or0;
  assign f_u_dadda_cla32_fa70_xor1 = f_u_dadda_cla32_fa70_xor0 ^ f_u_dadda_cla32_fa68_or0;
  assign f_u_dadda_cla32_fa70_and1 = f_u_dadda_cla32_fa70_xor0 & f_u_dadda_cla32_fa68_or0;
  assign f_u_dadda_cla32_fa70_or0 = f_u_dadda_cla32_fa70_and0 | f_u_dadda_cla32_fa70_and1;
  assign f_u_dadda_cla32_fa71_xor0 = f_u_dadda_cla32_fa67_or0 ^ f_u_dadda_cla32_fa66_or0;
  assign f_u_dadda_cla32_fa71_and0 = f_u_dadda_cla32_fa67_or0 & f_u_dadda_cla32_fa66_or0;
  assign f_u_dadda_cla32_fa71_xor1 = f_u_dadda_cla32_fa71_xor0 ^ f_u_dadda_cla32_fa65_or0;
  assign f_u_dadda_cla32_fa71_and1 = f_u_dadda_cla32_fa71_xor0 & f_u_dadda_cla32_fa65_or0;
  assign f_u_dadda_cla32_fa71_or0 = f_u_dadda_cla32_fa71_and0 | f_u_dadda_cla32_fa71_and1;
  assign f_u_dadda_cla32_fa72_xor0 = f_u_dadda_cla32_fa64_or0 ^ f_u_dadda_cla32_fa63_or0;
  assign f_u_dadda_cla32_fa72_and0 = f_u_dadda_cla32_fa64_or0 & f_u_dadda_cla32_fa63_or0;
  assign f_u_dadda_cla32_fa72_xor1 = f_u_dadda_cla32_fa72_xor0 ^ f_u_dadda_cla32_fa62_or0;
  assign f_u_dadda_cla32_fa72_and1 = f_u_dadda_cla32_fa72_xor0 & f_u_dadda_cla32_fa62_or0;
  assign f_u_dadda_cla32_fa72_or0 = f_u_dadda_cla32_fa72_and0 | f_u_dadda_cla32_fa72_and1;
  assign f_u_dadda_cla32_and_17_0 = a[17] & b[0];
  assign f_u_dadda_cla32_fa73_xor0 = f_u_dadda_cla32_fa61_or0 ^ f_u_dadda_cla32_fa60_or0;
  assign f_u_dadda_cla32_fa73_and0 = f_u_dadda_cla32_fa61_or0 & f_u_dadda_cla32_fa60_or0;
  assign f_u_dadda_cla32_fa73_xor1 = f_u_dadda_cla32_fa73_xor0 ^ f_u_dadda_cla32_and_17_0;
  assign f_u_dadda_cla32_fa73_and1 = f_u_dadda_cla32_fa73_xor0 & f_u_dadda_cla32_and_17_0;
  assign f_u_dadda_cla32_fa73_or0 = f_u_dadda_cla32_fa73_and0 | f_u_dadda_cla32_fa73_and1;
  assign f_u_dadda_cla32_and_16_1 = a[16] & b[1];
  assign f_u_dadda_cla32_and_15_2 = a[15] & b[2];
  assign f_u_dadda_cla32_and_14_3 = a[14] & b[3];
  assign f_u_dadda_cla32_fa74_xor0 = f_u_dadda_cla32_and_16_1 ^ f_u_dadda_cla32_and_15_2;
  assign f_u_dadda_cla32_fa74_and0 = f_u_dadda_cla32_and_16_1 & f_u_dadda_cla32_and_15_2;
  assign f_u_dadda_cla32_fa74_xor1 = f_u_dadda_cla32_fa74_xor0 ^ f_u_dadda_cla32_and_14_3;
  assign f_u_dadda_cla32_fa74_and1 = f_u_dadda_cla32_fa74_xor0 & f_u_dadda_cla32_and_14_3;
  assign f_u_dadda_cla32_fa74_or0 = f_u_dadda_cla32_fa74_and0 | f_u_dadda_cla32_fa74_and1;
  assign f_u_dadda_cla32_and_13_4 = a[13] & b[4];
  assign f_u_dadda_cla32_and_12_5 = a[12] & b[5];
  assign f_u_dadda_cla32_and_11_6 = a[11] & b[6];
  assign f_u_dadda_cla32_fa75_xor0 = f_u_dadda_cla32_and_13_4 ^ f_u_dadda_cla32_and_12_5;
  assign f_u_dadda_cla32_fa75_and0 = f_u_dadda_cla32_and_13_4 & f_u_dadda_cla32_and_12_5;
  assign f_u_dadda_cla32_fa75_xor1 = f_u_dadda_cla32_fa75_xor0 ^ f_u_dadda_cla32_and_11_6;
  assign f_u_dadda_cla32_fa75_and1 = f_u_dadda_cla32_fa75_xor0 & f_u_dadda_cla32_and_11_6;
  assign f_u_dadda_cla32_fa75_or0 = f_u_dadda_cla32_fa75_and0 | f_u_dadda_cla32_fa75_and1;
  assign f_u_dadda_cla32_and_10_7 = a[10] & b[7];
  assign f_u_dadda_cla32_and_9_8 = a[9] & b[8];
  assign f_u_dadda_cla32_and_8_9 = a[8] & b[9];
  assign f_u_dadda_cla32_fa76_xor0 = f_u_dadda_cla32_and_10_7 ^ f_u_dadda_cla32_and_9_8;
  assign f_u_dadda_cla32_fa76_and0 = f_u_dadda_cla32_and_10_7 & f_u_dadda_cla32_and_9_8;
  assign f_u_dadda_cla32_fa76_xor1 = f_u_dadda_cla32_fa76_xor0 ^ f_u_dadda_cla32_and_8_9;
  assign f_u_dadda_cla32_fa76_and1 = f_u_dadda_cla32_fa76_xor0 & f_u_dadda_cla32_and_8_9;
  assign f_u_dadda_cla32_fa76_or0 = f_u_dadda_cla32_fa76_and0 | f_u_dadda_cla32_fa76_and1;
  assign f_u_dadda_cla32_and_7_10 = a[7] & b[10];
  assign f_u_dadda_cla32_and_6_11 = a[6] & b[11];
  assign f_u_dadda_cla32_and_5_12 = a[5] & b[12];
  assign f_u_dadda_cla32_fa77_xor0 = f_u_dadda_cla32_and_7_10 ^ f_u_dadda_cla32_and_6_11;
  assign f_u_dadda_cla32_fa77_and0 = f_u_dadda_cla32_and_7_10 & f_u_dadda_cla32_and_6_11;
  assign f_u_dadda_cla32_fa77_xor1 = f_u_dadda_cla32_fa77_xor0 ^ f_u_dadda_cla32_and_5_12;
  assign f_u_dadda_cla32_fa77_and1 = f_u_dadda_cla32_fa77_xor0 & f_u_dadda_cla32_and_5_12;
  assign f_u_dadda_cla32_fa77_or0 = f_u_dadda_cla32_fa77_and0 | f_u_dadda_cla32_fa77_and1;
  assign f_u_dadda_cla32_and_4_13 = a[4] & b[13];
  assign f_u_dadda_cla32_and_3_14 = a[3] & b[14];
  assign f_u_dadda_cla32_and_2_15 = a[2] & b[15];
  assign f_u_dadda_cla32_fa78_xor0 = f_u_dadda_cla32_and_4_13 ^ f_u_dadda_cla32_and_3_14;
  assign f_u_dadda_cla32_fa78_and0 = f_u_dadda_cla32_and_4_13 & f_u_dadda_cla32_and_3_14;
  assign f_u_dadda_cla32_fa78_xor1 = f_u_dadda_cla32_fa78_xor0 ^ f_u_dadda_cla32_and_2_15;
  assign f_u_dadda_cla32_fa78_and1 = f_u_dadda_cla32_fa78_xor0 & f_u_dadda_cla32_and_2_15;
  assign f_u_dadda_cla32_fa78_or0 = f_u_dadda_cla32_fa78_and0 | f_u_dadda_cla32_fa78_and1;
  assign f_u_dadda_cla32_and_1_16 = a[1] & b[16];
  assign f_u_dadda_cla32_and_0_17 = a[0] & b[17];
  assign f_u_dadda_cla32_fa79_xor0 = f_u_dadda_cla32_and_1_16 ^ f_u_dadda_cla32_and_0_17;
  assign f_u_dadda_cla32_fa79_and0 = f_u_dadda_cla32_and_1_16 & f_u_dadda_cla32_and_0_17;
  assign f_u_dadda_cla32_fa79_xor1 = f_u_dadda_cla32_fa79_xor0 ^ f_u_dadda_cla32_fa70_xor1;
  assign f_u_dadda_cla32_fa79_and1 = f_u_dadda_cla32_fa79_xor0 & f_u_dadda_cla32_fa70_xor1;
  assign f_u_dadda_cla32_fa79_or0 = f_u_dadda_cla32_fa79_and0 | f_u_dadda_cla32_fa79_and1;
  assign f_u_dadda_cla32_fa80_xor0 = f_u_dadda_cla32_fa71_xor1 ^ f_u_dadda_cla32_fa72_xor1;
  assign f_u_dadda_cla32_fa80_and0 = f_u_dadda_cla32_fa71_xor1 & f_u_dadda_cla32_fa72_xor1;
  assign f_u_dadda_cla32_fa80_xor1 = f_u_dadda_cla32_fa80_xor0 ^ f_u_dadda_cla32_fa73_xor1;
  assign f_u_dadda_cla32_fa80_and1 = f_u_dadda_cla32_fa80_xor0 & f_u_dadda_cla32_fa73_xor1;
  assign f_u_dadda_cla32_fa80_or0 = f_u_dadda_cla32_fa80_and0 | f_u_dadda_cla32_fa80_and1;
  assign f_u_dadda_cla32_ha16_xor0 = f_u_dadda_cla32_fa74_xor1 ^ f_u_dadda_cla32_fa75_xor1;
  assign f_u_dadda_cla32_ha16_and0 = f_u_dadda_cla32_fa74_xor1 & f_u_dadda_cla32_fa75_xor1;
  assign f_u_dadda_cla32_fa81_xor0 = f_u_dadda_cla32_ha16_and0 ^ f_u_dadda_cla32_fa80_or0;
  assign f_u_dadda_cla32_fa81_and0 = f_u_dadda_cla32_ha16_and0 & f_u_dadda_cla32_fa80_or0;
  assign f_u_dadda_cla32_fa81_xor1 = f_u_dadda_cla32_fa81_xor0 ^ f_u_dadda_cla32_fa79_or0;
  assign f_u_dadda_cla32_fa81_and1 = f_u_dadda_cla32_fa81_xor0 & f_u_dadda_cla32_fa79_or0;
  assign f_u_dadda_cla32_fa81_or0 = f_u_dadda_cla32_fa81_and0 | f_u_dadda_cla32_fa81_and1;
  assign f_u_dadda_cla32_fa82_xor0 = f_u_dadda_cla32_fa78_or0 ^ f_u_dadda_cla32_fa77_or0;
  assign f_u_dadda_cla32_fa82_and0 = f_u_dadda_cla32_fa78_or0 & f_u_dadda_cla32_fa77_or0;
  assign f_u_dadda_cla32_fa82_xor1 = f_u_dadda_cla32_fa82_xor0 ^ f_u_dadda_cla32_fa76_or0;
  assign f_u_dadda_cla32_fa82_and1 = f_u_dadda_cla32_fa82_xor0 & f_u_dadda_cla32_fa76_or0;
  assign f_u_dadda_cla32_fa82_or0 = f_u_dadda_cla32_fa82_and0 | f_u_dadda_cla32_fa82_and1;
  assign f_u_dadda_cla32_fa83_xor0 = f_u_dadda_cla32_fa75_or0 ^ f_u_dadda_cla32_fa74_or0;
  assign f_u_dadda_cla32_fa83_and0 = f_u_dadda_cla32_fa75_or0 & f_u_dadda_cla32_fa74_or0;
  assign f_u_dadda_cla32_fa83_xor1 = f_u_dadda_cla32_fa83_xor0 ^ f_u_dadda_cla32_fa73_or0;
  assign f_u_dadda_cla32_fa83_and1 = f_u_dadda_cla32_fa83_xor0 & f_u_dadda_cla32_fa73_or0;
  assign f_u_dadda_cla32_fa83_or0 = f_u_dadda_cla32_fa83_and0 | f_u_dadda_cla32_fa83_and1;
  assign f_u_dadda_cla32_fa84_xor0 = f_u_dadda_cla32_fa72_or0 ^ f_u_dadda_cla32_fa71_or0;
  assign f_u_dadda_cla32_fa84_and0 = f_u_dadda_cla32_fa72_or0 & f_u_dadda_cla32_fa71_or0;
  assign f_u_dadda_cla32_fa84_xor1 = f_u_dadda_cla32_fa84_xor0 ^ f_u_dadda_cla32_fa70_or0;
  assign f_u_dadda_cla32_fa84_and1 = f_u_dadda_cla32_fa84_xor0 & f_u_dadda_cla32_fa70_or0;
  assign f_u_dadda_cla32_fa84_or0 = f_u_dadda_cla32_fa84_and0 | f_u_dadda_cla32_fa84_and1;
  assign f_u_dadda_cla32_and_18_0 = a[18] & b[0];
  assign f_u_dadda_cla32_and_17_1 = a[17] & b[1];
  assign f_u_dadda_cla32_and_16_2 = a[16] & b[2];
  assign f_u_dadda_cla32_fa85_xor0 = f_u_dadda_cla32_and_18_0 ^ f_u_dadda_cla32_and_17_1;
  assign f_u_dadda_cla32_fa85_and0 = f_u_dadda_cla32_and_18_0 & f_u_dadda_cla32_and_17_1;
  assign f_u_dadda_cla32_fa85_xor1 = f_u_dadda_cla32_fa85_xor0 ^ f_u_dadda_cla32_and_16_2;
  assign f_u_dadda_cla32_fa85_and1 = f_u_dadda_cla32_fa85_xor0 & f_u_dadda_cla32_and_16_2;
  assign f_u_dadda_cla32_fa85_or0 = f_u_dadda_cla32_fa85_and0 | f_u_dadda_cla32_fa85_and1;
  assign f_u_dadda_cla32_and_15_3 = a[15] & b[3];
  assign f_u_dadda_cla32_and_14_4 = a[14] & b[4];
  assign f_u_dadda_cla32_and_13_5 = a[13] & b[5];
  assign f_u_dadda_cla32_fa86_xor0 = f_u_dadda_cla32_and_15_3 ^ f_u_dadda_cla32_and_14_4;
  assign f_u_dadda_cla32_fa86_and0 = f_u_dadda_cla32_and_15_3 & f_u_dadda_cla32_and_14_4;
  assign f_u_dadda_cla32_fa86_xor1 = f_u_dadda_cla32_fa86_xor0 ^ f_u_dadda_cla32_and_13_5;
  assign f_u_dadda_cla32_fa86_and1 = f_u_dadda_cla32_fa86_xor0 & f_u_dadda_cla32_and_13_5;
  assign f_u_dadda_cla32_fa86_or0 = f_u_dadda_cla32_fa86_and0 | f_u_dadda_cla32_fa86_and1;
  assign f_u_dadda_cla32_and_12_6 = a[12] & b[6];
  assign f_u_dadda_cla32_and_11_7 = a[11] & b[7];
  assign f_u_dadda_cla32_and_10_8 = a[10] & b[8];
  assign f_u_dadda_cla32_fa87_xor0 = f_u_dadda_cla32_and_12_6 ^ f_u_dadda_cla32_and_11_7;
  assign f_u_dadda_cla32_fa87_and0 = f_u_dadda_cla32_and_12_6 & f_u_dadda_cla32_and_11_7;
  assign f_u_dadda_cla32_fa87_xor1 = f_u_dadda_cla32_fa87_xor0 ^ f_u_dadda_cla32_and_10_8;
  assign f_u_dadda_cla32_fa87_and1 = f_u_dadda_cla32_fa87_xor0 & f_u_dadda_cla32_and_10_8;
  assign f_u_dadda_cla32_fa87_or0 = f_u_dadda_cla32_fa87_and0 | f_u_dadda_cla32_fa87_and1;
  assign f_u_dadda_cla32_and_9_9 = a[9] & b[9];
  assign f_u_dadda_cla32_and_8_10 = a[8] & b[10];
  assign f_u_dadda_cla32_and_7_11 = a[7] & b[11];
  assign f_u_dadda_cla32_fa88_xor0 = f_u_dadda_cla32_and_9_9 ^ f_u_dadda_cla32_and_8_10;
  assign f_u_dadda_cla32_fa88_and0 = f_u_dadda_cla32_and_9_9 & f_u_dadda_cla32_and_8_10;
  assign f_u_dadda_cla32_fa88_xor1 = f_u_dadda_cla32_fa88_xor0 ^ f_u_dadda_cla32_and_7_11;
  assign f_u_dadda_cla32_fa88_and1 = f_u_dadda_cla32_fa88_xor0 & f_u_dadda_cla32_and_7_11;
  assign f_u_dadda_cla32_fa88_or0 = f_u_dadda_cla32_fa88_and0 | f_u_dadda_cla32_fa88_and1;
  assign f_u_dadda_cla32_and_6_12 = a[6] & b[12];
  assign f_u_dadda_cla32_and_5_13 = a[5] & b[13];
  assign f_u_dadda_cla32_and_4_14 = a[4] & b[14];
  assign f_u_dadda_cla32_fa89_xor0 = f_u_dadda_cla32_and_6_12 ^ f_u_dadda_cla32_and_5_13;
  assign f_u_dadda_cla32_fa89_and0 = f_u_dadda_cla32_and_6_12 & f_u_dadda_cla32_and_5_13;
  assign f_u_dadda_cla32_fa89_xor1 = f_u_dadda_cla32_fa89_xor0 ^ f_u_dadda_cla32_and_4_14;
  assign f_u_dadda_cla32_fa89_and1 = f_u_dadda_cla32_fa89_xor0 & f_u_dadda_cla32_and_4_14;
  assign f_u_dadda_cla32_fa89_or0 = f_u_dadda_cla32_fa89_and0 | f_u_dadda_cla32_fa89_and1;
  assign f_u_dadda_cla32_and_3_15 = a[3] & b[15];
  assign f_u_dadda_cla32_and_2_16 = a[2] & b[16];
  assign f_u_dadda_cla32_and_1_17 = a[1] & b[17];
  assign f_u_dadda_cla32_fa90_xor0 = f_u_dadda_cla32_and_3_15 ^ f_u_dadda_cla32_and_2_16;
  assign f_u_dadda_cla32_fa90_and0 = f_u_dadda_cla32_and_3_15 & f_u_dadda_cla32_and_2_16;
  assign f_u_dadda_cla32_fa90_xor1 = f_u_dadda_cla32_fa90_xor0 ^ f_u_dadda_cla32_and_1_17;
  assign f_u_dadda_cla32_fa90_and1 = f_u_dadda_cla32_fa90_xor0 & f_u_dadda_cla32_and_1_17;
  assign f_u_dadda_cla32_fa90_or0 = f_u_dadda_cla32_fa90_and0 | f_u_dadda_cla32_fa90_and1;
  assign f_u_dadda_cla32_and_0_18 = a[0] & b[18];
  assign f_u_dadda_cla32_fa91_xor0 = f_u_dadda_cla32_and_0_18 ^ f_u_dadda_cla32_fa81_xor1;
  assign f_u_dadda_cla32_fa91_and0 = f_u_dadda_cla32_and_0_18 & f_u_dadda_cla32_fa81_xor1;
  assign f_u_dadda_cla32_fa91_xor1 = f_u_dadda_cla32_fa91_xor0 ^ f_u_dadda_cla32_fa82_xor1;
  assign f_u_dadda_cla32_fa91_and1 = f_u_dadda_cla32_fa91_xor0 & f_u_dadda_cla32_fa82_xor1;
  assign f_u_dadda_cla32_fa91_or0 = f_u_dadda_cla32_fa91_and0 | f_u_dadda_cla32_fa91_and1;
  assign f_u_dadda_cla32_fa92_xor0 = f_u_dadda_cla32_fa83_xor1 ^ f_u_dadda_cla32_fa84_xor1;
  assign f_u_dadda_cla32_fa92_and0 = f_u_dadda_cla32_fa83_xor1 & f_u_dadda_cla32_fa84_xor1;
  assign f_u_dadda_cla32_fa92_xor1 = f_u_dadda_cla32_fa92_xor0 ^ f_u_dadda_cla32_fa85_xor1;
  assign f_u_dadda_cla32_fa92_and1 = f_u_dadda_cla32_fa92_xor0 & f_u_dadda_cla32_fa85_xor1;
  assign f_u_dadda_cla32_fa92_or0 = f_u_dadda_cla32_fa92_and0 | f_u_dadda_cla32_fa92_and1;
  assign f_u_dadda_cla32_ha17_xor0 = f_u_dadda_cla32_fa86_xor1 ^ f_u_dadda_cla32_fa87_xor1;
  assign f_u_dadda_cla32_ha17_and0 = f_u_dadda_cla32_fa86_xor1 & f_u_dadda_cla32_fa87_xor1;
  assign f_u_dadda_cla32_fa93_xor0 = f_u_dadda_cla32_ha17_and0 ^ f_u_dadda_cla32_fa92_or0;
  assign f_u_dadda_cla32_fa93_and0 = f_u_dadda_cla32_ha17_and0 & f_u_dadda_cla32_fa92_or0;
  assign f_u_dadda_cla32_fa93_xor1 = f_u_dadda_cla32_fa93_xor0 ^ f_u_dadda_cla32_fa91_or0;
  assign f_u_dadda_cla32_fa93_and1 = f_u_dadda_cla32_fa93_xor0 & f_u_dadda_cla32_fa91_or0;
  assign f_u_dadda_cla32_fa93_or0 = f_u_dadda_cla32_fa93_and0 | f_u_dadda_cla32_fa93_and1;
  assign f_u_dadda_cla32_fa94_xor0 = f_u_dadda_cla32_fa90_or0 ^ f_u_dadda_cla32_fa89_or0;
  assign f_u_dadda_cla32_fa94_and0 = f_u_dadda_cla32_fa90_or0 & f_u_dadda_cla32_fa89_or0;
  assign f_u_dadda_cla32_fa94_xor1 = f_u_dadda_cla32_fa94_xor0 ^ f_u_dadda_cla32_fa88_or0;
  assign f_u_dadda_cla32_fa94_and1 = f_u_dadda_cla32_fa94_xor0 & f_u_dadda_cla32_fa88_or0;
  assign f_u_dadda_cla32_fa94_or0 = f_u_dadda_cla32_fa94_and0 | f_u_dadda_cla32_fa94_and1;
  assign f_u_dadda_cla32_fa95_xor0 = f_u_dadda_cla32_fa87_or0 ^ f_u_dadda_cla32_fa86_or0;
  assign f_u_dadda_cla32_fa95_and0 = f_u_dadda_cla32_fa87_or0 & f_u_dadda_cla32_fa86_or0;
  assign f_u_dadda_cla32_fa95_xor1 = f_u_dadda_cla32_fa95_xor0 ^ f_u_dadda_cla32_fa85_or0;
  assign f_u_dadda_cla32_fa95_and1 = f_u_dadda_cla32_fa95_xor0 & f_u_dadda_cla32_fa85_or0;
  assign f_u_dadda_cla32_fa95_or0 = f_u_dadda_cla32_fa95_and0 | f_u_dadda_cla32_fa95_and1;
  assign f_u_dadda_cla32_fa96_xor0 = f_u_dadda_cla32_fa84_or0 ^ f_u_dadda_cla32_fa83_or0;
  assign f_u_dadda_cla32_fa96_and0 = f_u_dadda_cla32_fa84_or0 & f_u_dadda_cla32_fa83_or0;
  assign f_u_dadda_cla32_fa96_xor1 = f_u_dadda_cla32_fa96_xor0 ^ f_u_dadda_cla32_fa82_or0;
  assign f_u_dadda_cla32_fa96_and1 = f_u_dadda_cla32_fa96_xor0 & f_u_dadda_cla32_fa82_or0;
  assign f_u_dadda_cla32_fa96_or0 = f_u_dadda_cla32_fa96_and0 | f_u_dadda_cla32_fa96_and1;
  assign f_u_dadda_cla32_and_19_0 = a[19] & b[0];
  assign f_u_dadda_cla32_and_18_1 = a[18] & b[1];
  assign f_u_dadda_cla32_fa97_xor0 = f_u_dadda_cla32_fa81_or0 ^ f_u_dadda_cla32_and_19_0;
  assign f_u_dadda_cla32_fa97_and0 = f_u_dadda_cla32_fa81_or0 & f_u_dadda_cla32_and_19_0;
  assign f_u_dadda_cla32_fa97_xor1 = f_u_dadda_cla32_fa97_xor0 ^ f_u_dadda_cla32_and_18_1;
  assign f_u_dadda_cla32_fa97_and1 = f_u_dadda_cla32_fa97_xor0 & f_u_dadda_cla32_and_18_1;
  assign f_u_dadda_cla32_fa97_or0 = f_u_dadda_cla32_fa97_and0 | f_u_dadda_cla32_fa97_and1;
  assign f_u_dadda_cla32_and_17_2 = a[17] & b[2];
  assign f_u_dadda_cla32_and_16_3 = a[16] & b[3];
  assign f_u_dadda_cla32_and_15_4 = a[15] & b[4];
  assign f_u_dadda_cla32_fa98_xor0 = f_u_dadda_cla32_and_17_2 ^ f_u_dadda_cla32_and_16_3;
  assign f_u_dadda_cla32_fa98_and0 = f_u_dadda_cla32_and_17_2 & f_u_dadda_cla32_and_16_3;
  assign f_u_dadda_cla32_fa98_xor1 = f_u_dadda_cla32_fa98_xor0 ^ f_u_dadda_cla32_and_15_4;
  assign f_u_dadda_cla32_fa98_and1 = f_u_dadda_cla32_fa98_xor0 & f_u_dadda_cla32_and_15_4;
  assign f_u_dadda_cla32_fa98_or0 = f_u_dadda_cla32_fa98_and0 | f_u_dadda_cla32_fa98_and1;
  assign f_u_dadda_cla32_and_14_5 = a[14] & b[5];
  assign f_u_dadda_cla32_and_13_6 = a[13] & b[6];
  assign f_u_dadda_cla32_and_12_7 = a[12] & b[7];
  assign f_u_dadda_cla32_fa99_xor0 = f_u_dadda_cla32_and_14_5 ^ f_u_dadda_cla32_and_13_6;
  assign f_u_dadda_cla32_fa99_and0 = f_u_dadda_cla32_and_14_5 & f_u_dadda_cla32_and_13_6;
  assign f_u_dadda_cla32_fa99_xor1 = f_u_dadda_cla32_fa99_xor0 ^ f_u_dadda_cla32_and_12_7;
  assign f_u_dadda_cla32_fa99_and1 = f_u_dadda_cla32_fa99_xor0 & f_u_dadda_cla32_and_12_7;
  assign f_u_dadda_cla32_fa99_or0 = f_u_dadda_cla32_fa99_and0 | f_u_dadda_cla32_fa99_and1;
  assign f_u_dadda_cla32_and_11_8 = a[11] & b[8];
  assign f_u_dadda_cla32_and_10_9 = a[10] & b[9];
  assign f_u_dadda_cla32_and_9_10 = a[9] & b[10];
  assign f_u_dadda_cla32_fa100_xor0 = f_u_dadda_cla32_and_11_8 ^ f_u_dadda_cla32_and_10_9;
  assign f_u_dadda_cla32_fa100_and0 = f_u_dadda_cla32_and_11_8 & f_u_dadda_cla32_and_10_9;
  assign f_u_dadda_cla32_fa100_xor1 = f_u_dadda_cla32_fa100_xor0 ^ f_u_dadda_cla32_and_9_10;
  assign f_u_dadda_cla32_fa100_and1 = f_u_dadda_cla32_fa100_xor0 & f_u_dadda_cla32_and_9_10;
  assign f_u_dadda_cla32_fa100_or0 = f_u_dadda_cla32_fa100_and0 | f_u_dadda_cla32_fa100_and1;
  assign f_u_dadda_cla32_and_8_11 = a[8] & b[11];
  assign f_u_dadda_cla32_and_7_12 = a[7] & b[12];
  assign f_u_dadda_cla32_and_6_13 = a[6] & b[13];
  assign f_u_dadda_cla32_fa101_xor0 = f_u_dadda_cla32_and_8_11 ^ f_u_dadda_cla32_and_7_12;
  assign f_u_dadda_cla32_fa101_and0 = f_u_dadda_cla32_and_8_11 & f_u_dadda_cla32_and_7_12;
  assign f_u_dadda_cla32_fa101_xor1 = f_u_dadda_cla32_fa101_xor0 ^ f_u_dadda_cla32_and_6_13;
  assign f_u_dadda_cla32_fa101_and1 = f_u_dadda_cla32_fa101_xor0 & f_u_dadda_cla32_and_6_13;
  assign f_u_dadda_cla32_fa101_or0 = f_u_dadda_cla32_fa101_and0 | f_u_dadda_cla32_fa101_and1;
  assign f_u_dadda_cla32_and_5_14 = a[5] & b[14];
  assign f_u_dadda_cla32_and_4_15 = a[4] & b[15];
  assign f_u_dadda_cla32_and_3_16 = a[3] & b[16];
  assign f_u_dadda_cla32_fa102_xor0 = f_u_dadda_cla32_and_5_14 ^ f_u_dadda_cla32_and_4_15;
  assign f_u_dadda_cla32_fa102_and0 = f_u_dadda_cla32_and_5_14 & f_u_dadda_cla32_and_4_15;
  assign f_u_dadda_cla32_fa102_xor1 = f_u_dadda_cla32_fa102_xor0 ^ f_u_dadda_cla32_and_3_16;
  assign f_u_dadda_cla32_fa102_and1 = f_u_dadda_cla32_fa102_xor0 & f_u_dadda_cla32_and_3_16;
  assign f_u_dadda_cla32_fa102_or0 = f_u_dadda_cla32_fa102_and0 | f_u_dadda_cla32_fa102_and1;
  assign f_u_dadda_cla32_and_2_17 = a[2] & b[17];
  assign f_u_dadda_cla32_and_1_18 = a[1] & b[18];
  assign f_u_dadda_cla32_and_0_19 = a[0] & b[19];
  assign f_u_dadda_cla32_fa103_xor0 = f_u_dadda_cla32_and_2_17 ^ f_u_dadda_cla32_and_1_18;
  assign f_u_dadda_cla32_fa103_and0 = f_u_dadda_cla32_and_2_17 & f_u_dadda_cla32_and_1_18;
  assign f_u_dadda_cla32_fa103_xor1 = f_u_dadda_cla32_fa103_xor0 ^ f_u_dadda_cla32_and_0_19;
  assign f_u_dadda_cla32_fa103_and1 = f_u_dadda_cla32_fa103_xor0 & f_u_dadda_cla32_and_0_19;
  assign f_u_dadda_cla32_fa103_or0 = f_u_dadda_cla32_fa103_and0 | f_u_dadda_cla32_fa103_and1;
  assign f_u_dadda_cla32_fa104_xor0 = f_u_dadda_cla32_fa93_xor1 ^ f_u_dadda_cla32_fa94_xor1;
  assign f_u_dadda_cla32_fa104_and0 = f_u_dadda_cla32_fa93_xor1 & f_u_dadda_cla32_fa94_xor1;
  assign f_u_dadda_cla32_fa104_xor1 = f_u_dadda_cla32_fa104_xor0 ^ f_u_dadda_cla32_fa95_xor1;
  assign f_u_dadda_cla32_fa104_and1 = f_u_dadda_cla32_fa104_xor0 & f_u_dadda_cla32_fa95_xor1;
  assign f_u_dadda_cla32_fa104_or0 = f_u_dadda_cla32_fa104_and0 | f_u_dadda_cla32_fa104_and1;
  assign f_u_dadda_cla32_fa105_xor0 = f_u_dadda_cla32_fa96_xor1 ^ f_u_dadda_cla32_fa97_xor1;
  assign f_u_dadda_cla32_fa105_and0 = f_u_dadda_cla32_fa96_xor1 & f_u_dadda_cla32_fa97_xor1;
  assign f_u_dadda_cla32_fa105_xor1 = f_u_dadda_cla32_fa105_xor0 ^ f_u_dadda_cla32_fa98_xor1;
  assign f_u_dadda_cla32_fa105_and1 = f_u_dadda_cla32_fa105_xor0 & f_u_dadda_cla32_fa98_xor1;
  assign f_u_dadda_cla32_fa105_or0 = f_u_dadda_cla32_fa105_and0 | f_u_dadda_cla32_fa105_and1;
  assign f_u_dadda_cla32_ha18_xor0 = f_u_dadda_cla32_fa99_xor1 ^ f_u_dadda_cla32_fa100_xor1;
  assign f_u_dadda_cla32_ha18_and0 = f_u_dadda_cla32_fa99_xor1 & f_u_dadda_cla32_fa100_xor1;
  assign f_u_dadda_cla32_fa106_xor0 = f_u_dadda_cla32_ha18_and0 ^ f_u_dadda_cla32_fa105_or0;
  assign f_u_dadda_cla32_fa106_and0 = f_u_dadda_cla32_ha18_and0 & f_u_dadda_cla32_fa105_or0;
  assign f_u_dadda_cla32_fa106_xor1 = f_u_dadda_cla32_fa106_xor0 ^ f_u_dadda_cla32_fa104_or0;
  assign f_u_dadda_cla32_fa106_and1 = f_u_dadda_cla32_fa106_xor0 & f_u_dadda_cla32_fa104_or0;
  assign f_u_dadda_cla32_fa106_or0 = f_u_dadda_cla32_fa106_and0 | f_u_dadda_cla32_fa106_and1;
  assign f_u_dadda_cla32_fa107_xor0 = f_u_dadda_cla32_fa103_or0 ^ f_u_dadda_cla32_fa102_or0;
  assign f_u_dadda_cla32_fa107_and0 = f_u_dadda_cla32_fa103_or0 & f_u_dadda_cla32_fa102_or0;
  assign f_u_dadda_cla32_fa107_xor1 = f_u_dadda_cla32_fa107_xor0 ^ f_u_dadda_cla32_fa101_or0;
  assign f_u_dadda_cla32_fa107_and1 = f_u_dadda_cla32_fa107_xor0 & f_u_dadda_cla32_fa101_or0;
  assign f_u_dadda_cla32_fa107_or0 = f_u_dadda_cla32_fa107_and0 | f_u_dadda_cla32_fa107_and1;
  assign f_u_dadda_cla32_fa108_xor0 = f_u_dadda_cla32_fa100_or0 ^ f_u_dadda_cla32_fa99_or0;
  assign f_u_dadda_cla32_fa108_and0 = f_u_dadda_cla32_fa100_or0 & f_u_dadda_cla32_fa99_or0;
  assign f_u_dadda_cla32_fa108_xor1 = f_u_dadda_cla32_fa108_xor0 ^ f_u_dadda_cla32_fa98_or0;
  assign f_u_dadda_cla32_fa108_and1 = f_u_dadda_cla32_fa108_xor0 & f_u_dadda_cla32_fa98_or0;
  assign f_u_dadda_cla32_fa108_or0 = f_u_dadda_cla32_fa108_and0 | f_u_dadda_cla32_fa108_and1;
  assign f_u_dadda_cla32_fa109_xor0 = f_u_dadda_cla32_fa97_or0 ^ f_u_dadda_cla32_fa96_or0;
  assign f_u_dadda_cla32_fa109_and0 = f_u_dadda_cla32_fa97_or0 & f_u_dadda_cla32_fa96_or0;
  assign f_u_dadda_cla32_fa109_xor1 = f_u_dadda_cla32_fa109_xor0 ^ f_u_dadda_cla32_fa95_or0;
  assign f_u_dadda_cla32_fa109_and1 = f_u_dadda_cla32_fa109_xor0 & f_u_dadda_cla32_fa95_or0;
  assign f_u_dadda_cla32_fa109_or0 = f_u_dadda_cla32_fa109_and0 | f_u_dadda_cla32_fa109_and1;
  assign f_u_dadda_cla32_and_20_0 = a[20] & b[0];
  assign f_u_dadda_cla32_fa110_xor0 = f_u_dadda_cla32_fa94_or0 ^ f_u_dadda_cla32_fa93_or0;
  assign f_u_dadda_cla32_fa110_and0 = f_u_dadda_cla32_fa94_or0 & f_u_dadda_cla32_fa93_or0;
  assign f_u_dadda_cla32_fa110_xor1 = f_u_dadda_cla32_fa110_xor0 ^ f_u_dadda_cla32_and_20_0;
  assign f_u_dadda_cla32_fa110_and1 = f_u_dadda_cla32_fa110_xor0 & f_u_dadda_cla32_and_20_0;
  assign f_u_dadda_cla32_fa110_or0 = f_u_dadda_cla32_fa110_and0 | f_u_dadda_cla32_fa110_and1;
  assign f_u_dadda_cla32_and_19_1 = a[19] & b[1];
  assign f_u_dadda_cla32_and_18_2 = a[18] & b[2];
  assign f_u_dadda_cla32_and_17_3 = a[17] & b[3];
  assign f_u_dadda_cla32_fa111_xor0 = f_u_dadda_cla32_and_19_1 ^ f_u_dadda_cla32_and_18_2;
  assign f_u_dadda_cla32_fa111_and0 = f_u_dadda_cla32_and_19_1 & f_u_dadda_cla32_and_18_2;
  assign f_u_dadda_cla32_fa111_xor1 = f_u_dadda_cla32_fa111_xor0 ^ f_u_dadda_cla32_and_17_3;
  assign f_u_dadda_cla32_fa111_and1 = f_u_dadda_cla32_fa111_xor0 & f_u_dadda_cla32_and_17_3;
  assign f_u_dadda_cla32_fa111_or0 = f_u_dadda_cla32_fa111_and0 | f_u_dadda_cla32_fa111_and1;
  assign f_u_dadda_cla32_and_16_4 = a[16] & b[4];
  assign f_u_dadda_cla32_and_15_5 = a[15] & b[5];
  assign f_u_dadda_cla32_and_14_6 = a[14] & b[6];
  assign f_u_dadda_cla32_fa112_xor0 = f_u_dadda_cla32_and_16_4 ^ f_u_dadda_cla32_and_15_5;
  assign f_u_dadda_cla32_fa112_and0 = f_u_dadda_cla32_and_16_4 & f_u_dadda_cla32_and_15_5;
  assign f_u_dadda_cla32_fa112_xor1 = f_u_dadda_cla32_fa112_xor0 ^ f_u_dadda_cla32_and_14_6;
  assign f_u_dadda_cla32_fa112_and1 = f_u_dadda_cla32_fa112_xor0 & f_u_dadda_cla32_and_14_6;
  assign f_u_dadda_cla32_fa112_or0 = f_u_dadda_cla32_fa112_and0 | f_u_dadda_cla32_fa112_and1;
  assign f_u_dadda_cla32_and_13_7 = a[13] & b[7];
  assign f_u_dadda_cla32_and_12_8 = a[12] & b[8];
  assign f_u_dadda_cla32_and_11_9 = a[11] & b[9];
  assign f_u_dadda_cla32_fa113_xor0 = f_u_dadda_cla32_and_13_7 ^ f_u_dadda_cla32_and_12_8;
  assign f_u_dadda_cla32_fa113_and0 = f_u_dadda_cla32_and_13_7 & f_u_dadda_cla32_and_12_8;
  assign f_u_dadda_cla32_fa113_xor1 = f_u_dadda_cla32_fa113_xor0 ^ f_u_dadda_cla32_and_11_9;
  assign f_u_dadda_cla32_fa113_and1 = f_u_dadda_cla32_fa113_xor0 & f_u_dadda_cla32_and_11_9;
  assign f_u_dadda_cla32_fa113_or0 = f_u_dadda_cla32_fa113_and0 | f_u_dadda_cla32_fa113_and1;
  assign f_u_dadda_cla32_and_10_10 = a[10] & b[10];
  assign f_u_dadda_cla32_and_9_11 = a[9] & b[11];
  assign f_u_dadda_cla32_and_8_12 = a[8] & b[12];
  assign f_u_dadda_cla32_fa114_xor0 = f_u_dadda_cla32_and_10_10 ^ f_u_dadda_cla32_and_9_11;
  assign f_u_dadda_cla32_fa114_and0 = f_u_dadda_cla32_and_10_10 & f_u_dadda_cla32_and_9_11;
  assign f_u_dadda_cla32_fa114_xor1 = f_u_dadda_cla32_fa114_xor0 ^ f_u_dadda_cla32_and_8_12;
  assign f_u_dadda_cla32_fa114_and1 = f_u_dadda_cla32_fa114_xor0 & f_u_dadda_cla32_and_8_12;
  assign f_u_dadda_cla32_fa114_or0 = f_u_dadda_cla32_fa114_and0 | f_u_dadda_cla32_fa114_and1;
  assign f_u_dadda_cla32_and_7_13 = a[7] & b[13];
  assign f_u_dadda_cla32_and_6_14 = a[6] & b[14];
  assign f_u_dadda_cla32_and_5_15 = a[5] & b[15];
  assign f_u_dadda_cla32_fa115_xor0 = f_u_dadda_cla32_and_7_13 ^ f_u_dadda_cla32_and_6_14;
  assign f_u_dadda_cla32_fa115_and0 = f_u_dadda_cla32_and_7_13 & f_u_dadda_cla32_and_6_14;
  assign f_u_dadda_cla32_fa115_xor1 = f_u_dadda_cla32_fa115_xor0 ^ f_u_dadda_cla32_and_5_15;
  assign f_u_dadda_cla32_fa115_and1 = f_u_dadda_cla32_fa115_xor0 & f_u_dadda_cla32_and_5_15;
  assign f_u_dadda_cla32_fa115_or0 = f_u_dadda_cla32_fa115_and0 | f_u_dadda_cla32_fa115_and1;
  assign f_u_dadda_cla32_and_4_16 = a[4] & b[16];
  assign f_u_dadda_cla32_and_3_17 = a[3] & b[17];
  assign f_u_dadda_cla32_and_2_18 = a[2] & b[18];
  assign f_u_dadda_cla32_fa116_xor0 = f_u_dadda_cla32_and_4_16 ^ f_u_dadda_cla32_and_3_17;
  assign f_u_dadda_cla32_fa116_and0 = f_u_dadda_cla32_and_4_16 & f_u_dadda_cla32_and_3_17;
  assign f_u_dadda_cla32_fa116_xor1 = f_u_dadda_cla32_fa116_xor0 ^ f_u_dadda_cla32_and_2_18;
  assign f_u_dadda_cla32_fa116_and1 = f_u_dadda_cla32_fa116_xor0 & f_u_dadda_cla32_and_2_18;
  assign f_u_dadda_cla32_fa116_or0 = f_u_dadda_cla32_fa116_and0 | f_u_dadda_cla32_fa116_and1;
  assign f_u_dadda_cla32_and_1_19 = a[1] & b[19];
  assign f_u_dadda_cla32_and_0_20 = a[0] & b[20];
  assign f_u_dadda_cla32_fa117_xor0 = f_u_dadda_cla32_and_1_19 ^ f_u_dadda_cla32_and_0_20;
  assign f_u_dadda_cla32_fa117_and0 = f_u_dadda_cla32_and_1_19 & f_u_dadda_cla32_and_0_20;
  assign f_u_dadda_cla32_fa117_xor1 = f_u_dadda_cla32_fa117_xor0 ^ f_u_dadda_cla32_fa106_xor1;
  assign f_u_dadda_cla32_fa117_and1 = f_u_dadda_cla32_fa117_xor0 & f_u_dadda_cla32_fa106_xor1;
  assign f_u_dadda_cla32_fa117_or0 = f_u_dadda_cla32_fa117_and0 | f_u_dadda_cla32_fa117_and1;
  assign f_u_dadda_cla32_fa118_xor0 = f_u_dadda_cla32_fa107_xor1 ^ f_u_dadda_cla32_fa108_xor1;
  assign f_u_dadda_cla32_fa118_and0 = f_u_dadda_cla32_fa107_xor1 & f_u_dadda_cla32_fa108_xor1;
  assign f_u_dadda_cla32_fa118_xor1 = f_u_dadda_cla32_fa118_xor0 ^ f_u_dadda_cla32_fa109_xor1;
  assign f_u_dadda_cla32_fa118_and1 = f_u_dadda_cla32_fa118_xor0 & f_u_dadda_cla32_fa109_xor1;
  assign f_u_dadda_cla32_fa118_or0 = f_u_dadda_cla32_fa118_and0 | f_u_dadda_cla32_fa118_and1;
  assign f_u_dadda_cla32_fa119_xor0 = f_u_dadda_cla32_fa110_xor1 ^ f_u_dadda_cla32_fa111_xor1;
  assign f_u_dadda_cla32_fa119_and0 = f_u_dadda_cla32_fa110_xor1 & f_u_dadda_cla32_fa111_xor1;
  assign f_u_dadda_cla32_fa119_xor1 = f_u_dadda_cla32_fa119_xor0 ^ f_u_dadda_cla32_fa112_xor1;
  assign f_u_dadda_cla32_fa119_and1 = f_u_dadda_cla32_fa119_xor0 & f_u_dadda_cla32_fa112_xor1;
  assign f_u_dadda_cla32_fa119_or0 = f_u_dadda_cla32_fa119_and0 | f_u_dadda_cla32_fa119_and1;
  assign f_u_dadda_cla32_ha19_xor0 = f_u_dadda_cla32_fa113_xor1 ^ f_u_dadda_cla32_fa114_xor1;
  assign f_u_dadda_cla32_ha19_and0 = f_u_dadda_cla32_fa113_xor1 & f_u_dadda_cla32_fa114_xor1;
  assign f_u_dadda_cla32_fa120_xor0 = f_u_dadda_cla32_ha19_and0 ^ f_u_dadda_cla32_fa119_or0;
  assign f_u_dadda_cla32_fa120_and0 = f_u_dadda_cla32_ha19_and0 & f_u_dadda_cla32_fa119_or0;
  assign f_u_dadda_cla32_fa120_xor1 = f_u_dadda_cla32_fa120_xor0 ^ f_u_dadda_cla32_fa118_or0;
  assign f_u_dadda_cla32_fa120_and1 = f_u_dadda_cla32_fa120_xor0 & f_u_dadda_cla32_fa118_or0;
  assign f_u_dadda_cla32_fa120_or0 = f_u_dadda_cla32_fa120_and0 | f_u_dadda_cla32_fa120_and1;
  assign f_u_dadda_cla32_fa121_xor0 = f_u_dadda_cla32_fa117_or0 ^ f_u_dadda_cla32_fa116_or0;
  assign f_u_dadda_cla32_fa121_and0 = f_u_dadda_cla32_fa117_or0 & f_u_dadda_cla32_fa116_or0;
  assign f_u_dadda_cla32_fa121_xor1 = f_u_dadda_cla32_fa121_xor0 ^ f_u_dadda_cla32_fa115_or0;
  assign f_u_dadda_cla32_fa121_and1 = f_u_dadda_cla32_fa121_xor0 & f_u_dadda_cla32_fa115_or0;
  assign f_u_dadda_cla32_fa121_or0 = f_u_dadda_cla32_fa121_and0 | f_u_dadda_cla32_fa121_and1;
  assign f_u_dadda_cla32_fa122_xor0 = f_u_dadda_cla32_fa114_or0 ^ f_u_dadda_cla32_fa113_or0;
  assign f_u_dadda_cla32_fa122_and0 = f_u_dadda_cla32_fa114_or0 & f_u_dadda_cla32_fa113_or0;
  assign f_u_dadda_cla32_fa122_xor1 = f_u_dadda_cla32_fa122_xor0 ^ f_u_dadda_cla32_fa112_or0;
  assign f_u_dadda_cla32_fa122_and1 = f_u_dadda_cla32_fa122_xor0 & f_u_dadda_cla32_fa112_or0;
  assign f_u_dadda_cla32_fa122_or0 = f_u_dadda_cla32_fa122_and0 | f_u_dadda_cla32_fa122_and1;
  assign f_u_dadda_cla32_fa123_xor0 = f_u_dadda_cla32_fa111_or0 ^ f_u_dadda_cla32_fa110_or0;
  assign f_u_dadda_cla32_fa123_and0 = f_u_dadda_cla32_fa111_or0 & f_u_dadda_cla32_fa110_or0;
  assign f_u_dadda_cla32_fa123_xor1 = f_u_dadda_cla32_fa123_xor0 ^ f_u_dadda_cla32_fa109_or0;
  assign f_u_dadda_cla32_fa123_and1 = f_u_dadda_cla32_fa123_xor0 & f_u_dadda_cla32_fa109_or0;
  assign f_u_dadda_cla32_fa123_or0 = f_u_dadda_cla32_fa123_and0 | f_u_dadda_cla32_fa123_and1;
  assign f_u_dadda_cla32_fa124_xor0 = f_u_dadda_cla32_fa108_or0 ^ f_u_dadda_cla32_fa107_or0;
  assign f_u_dadda_cla32_fa124_and0 = f_u_dadda_cla32_fa108_or0 & f_u_dadda_cla32_fa107_or0;
  assign f_u_dadda_cla32_fa124_xor1 = f_u_dadda_cla32_fa124_xor0 ^ f_u_dadda_cla32_fa106_or0;
  assign f_u_dadda_cla32_fa124_and1 = f_u_dadda_cla32_fa124_xor0 & f_u_dadda_cla32_fa106_or0;
  assign f_u_dadda_cla32_fa124_or0 = f_u_dadda_cla32_fa124_and0 | f_u_dadda_cla32_fa124_and1;
  assign f_u_dadda_cla32_and_21_0 = a[21] & b[0];
  assign f_u_dadda_cla32_and_20_1 = a[20] & b[1];
  assign f_u_dadda_cla32_and_19_2 = a[19] & b[2];
  assign f_u_dadda_cla32_fa125_xor0 = f_u_dadda_cla32_and_21_0 ^ f_u_dadda_cla32_and_20_1;
  assign f_u_dadda_cla32_fa125_and0 = f_u_dadda_cla32_and_21_0 & f_u_dadda_cla32_and_20_1;
  assign f_u_dadda_cla32_fa125_xor1 = f_u_dadda_cla32_fa125_xor0 ^ f_u_dadda_cla32_and_19_2;
  assign f_u_dadda_cla32_fa125_and1 = f_u_dadda_cla32_fa125_xor0 & f_u_dadda_cla32_and_19_2;
  assign f_u_dadda_cla32_fa125_or0 = f_u_dadda_cla32_fa125_and0 | f_u_dadda_cla32_fa125_and1;
  assign f_u_dadda_cla32_and_18_3 = a[18] & b[3];
  assign f_u_dadda_cla32_and_17_4 = a[17] & b[4];
  assign f_u_dadda_cla32_and_16_5 = a[16] & b[5];
  assign f_u_dadda_cla32_fa126_xor0 = f_u_dadda_cla32_and_18_3 ^ f_u_dadda_cla32_and_17_4;
  assign f_u_dadda_cla32_fa126_and0 = f_u_dadda_cla32_and_18_3 & f_u_dadda_cla32_and_17_4;
  assign f_u_dadda_cla32_fa126_xor1 = f_u_dadda_cla32_fa126_xor0 ^ f_u_dadda_cla32_and_16_5;
  assign f_u_dadda_cla32_fa126_and1 = f_u_dadda_cla32_fa126_xor0 & f_u_dadda_cla32_and_16_5;
  assign f_u_dadda_cla32_fa126_or0 = f_u_dadda_cla32_fa126_and0 | f_u_dadda_cla32_fa126_and1;
  assign f_u_dadda_cla32_and_15_6 = a[15] & b[6];
  assign f_u_dadda_cla32_and_14_7 = a[14] & b[7];
  assign f_u_dadda_cla32_and_13_8 = a[13] & b[8];
  assign f_u_dadda_cla32_fa127_xor0 = f_u_dadda_cla32_and_15_6 ^ f_u_dadda_cla32_and_14_7;
  assign f_u_dadda_cla32_fa127_and0 = f_u_dadda_cla32_and_15_6 & f_u_dadda_cla32_and_14_7;
  assign f_u_dadda_cla32_fa127_xor1 = f_u_dadda_cla32_fa127_xor0 ^ f_u_dadda_cla32_and_13_8;
  assign f_u_dadda_cla32_fa127_and1 = f_u_dadda_cla32_fa127_xor0 & f_u_dadda_cla32_and_13_8;
  assign f_u_dadda_cla32_fa127_or0 = f_u_dadda_cla32_fa127_and0 | f_u_dadda_cla32_fa127_and1;
  assign f_u_dadda_cla32_and_12_9 = a[12] & b[9];
  assign f_u_dadda_cla32_and_11_10 = a[11] & b[10];
  assign f_u_dadda_cla32_and_10_11 = a[10] & b[11];
  assign f_u_dadda_cla32_fa128_xor0 = f_u_dadda_cla32_and_12_9 ^ f_u_dadda_cla32_and_11_10;
  assign f_u_dadda_cla32_fa128_and0 = f_u_dadda_cla32_and_12_9 & f_u_dadda_cla32_and_11_10;
  assign f_u_dadda_cla32_fa128_xor1 = f_u_dadda_cla32_fa128_xor0 ^ f_u_dadda_cla32_and_10_11;
  assign f_u_dadda_cla32_fa128_and1 = f_u_dadda_cla32_fa128_xor0 & f_u_dadda_cla32_and_10_11;
  assign f_u_dadda_cla32_fa128_or0 = f_u_dadda_cla32_fa128_and0 | f_u_dadda_cla32_fa128_and1;
  assign f_u_dadda_cla32_and_9_12 = a[9] & b[12];
  assign f_u_dadda_cla32_and_8_13 = a[8] & b[13];
  assign f_u_dadda_cla32_and_7_14 = a[7] & b[14];
  assign f_u_dadda_cla32_fa129_xor0 = f_u_dadda_cla32_and_9_12 ^ f_u_dadda_cla32_and_8_13;
  assign f_u_dadda_cla32_fa129_and0 = f_u_dadda_cla32_and_9_12 & f_u_dadda_cla32_and_8_13;
  assign f_u_dadda_cla32_fa129_xor1 = f_u_dadda_cla32_fa129_xor0 ^ f_u_dadda_cla32_and_7_14;
  assign f_u_dadda_cla32_fa129_and1 = f_u_dadda_cla32_fa129_xor0 & f_u_dadda_cla32_and_7_14;
  assign f_u_dadda_cla32_fa129_or0 = f_u_dadda_cla32_fa129_and0 | f_u_dadda_cla32_fa129_and1;
  assign f_u_dadda_cla32_and_6_15 = a[6] & b[15];
  assign f_u_dadda_cla32_and_5_16 = a[5] & b[16];
  assign f_u_dadda_cla32_and_4_17 = a[4] & b[17];
  assign f_u_dadda_cla32_fa130_xor0 = f_u_dadda_cla32_and_6_15 ^ f_u_dadda_cla32_and_5_16;
  assign f_u_dadda_cla32_fa130_and0 = f_u_dadda_cla32_and_6_15 & f_u_dadda_cla32_and_5_16;
  assign f_u_dadda_cla32_fa130_xor1 = f_u_dadda_cla32_fa130_xor0 ^ f_u_dadda_cla32_and_4_17;
  assign f_u_dadda_cla32_fa130_and1 = f_u_dadda_cla32_fa130_xor0 & f_u_dadda_cla32_and_4_17;
  assign f_u_dadda_cla32_fa130_or0 = f_u_dadda_cla32_fa130_and0 | f_u_dadda_cla32_fa130_and1;
  assign f_u_dadda_cla32_and_3_18 = a[3] & b[18];
  assign f_u_dadda_cla32_and_2_19 = a[2] & b[19];
  assign f_u_dadda_cla32_and_1_20 = a[1] & b[20];
  assign f_u_dadda_cla32_fa131_xor0 = f_u_dadda_cla32_and_3_18 ^ f_u_dadda_cla32_and_2_19;
  assign f_u_dadda_cla32_fa131_and0 = f_u_dadda_cla32_and_3_18 & f_u_dadda_cla32_and_2_19;
  assign f_u_dadda_cla32_fa131_xor1 = f_u_dadda_cla32_fa131_xor0 ^ f_u_dadda_cla32_and_1_20;
  assign f_u_dadda_cla32_fa131_and1 = f_u_dadda_cla32_fa131_xor0 & f_u_dadda_cla32_and_1_20;
  assign f_u_dadda_cla32_fa131_or0 = f_u_dadda_cla32_fa131_and0 | f_u_dadda_cla32_fa131_and1;
  assign f_u_dadda_cla32_and_0_21 = a[0] & b[21];
  assign f_u_dadda_cla32_fa132_xor0 = f_u_dadda_cla32_and_0_21 ^ f_u_dadda_cla32_fa120_xor1;
  assign f_u_dadda_cla32_fa132_and0 = f_u_dadda_cla32_and_0_21 & f_u_dadda_cla32_fa120_xor1;
  assign f_u_dadda_cla32_fa132_xor1 = f_u_dadda_cla32_fa132_xor0 ^ f_u_dadda_cla32_fa121_xor1;
  assign f_u_dadda_cla32_fa132_and1 = f_u_dadda_cla32_fa132_xor0 & f_u_dadda_cla32_fa121_xor1;
  assign f_u_dadda_cla32_fa132_or0 = f_u_dadda_cla32_fa132_and0 | f_u_dadda_cla32_fa132_and1;
  assign f_u_dadda_cla32_fa133_xor0 = f_u_dadda_cla32_fa122_xor1 ^ f_u_dadda_cla32_fa123_xor1;
  assign f_u_dadda_cla32_fa133_and0 = f_u_dadda_cla32_fa122_xor1 & f_u_dadda_cla32_fa123_xor1;
  assign f_u_dadda_cla32_fa133_xor1 = f_u_dadda_cla32_fa133_xor0 ^ f_u_dadda_cla32_fa124_xor1;
  assign f_u_dadda_cla32_fa133_and1 = f_u_dadda_cla32_fa133_xor0 & f_u_dadda_cla32_fa124_xor1;
  assign f_u_dadda_cla32_fa133_or0 = f_u_dadda_cla32_fa133_and0 | f_u_dadda_cla32_fa133_and1;
  assign f_u_dadda_cla32_fa134_xor0 = f_u_dadda_cla32_fa125_xor1 ^ f_u_dadda_cla32_fa126_xor1;
  assign f_u_dadda_cla32_fa134_and0 = f_u_dadda_cla32_fa125_xor1 & f_u_dadda_cla32_fa126_xor1;
  assign f_u_dadda_cla32_fa134_xor1 = f_u_dadda_cla32_fa134_xor0 ^ f_u_dadda_cla32_fa127_xor1;
  assign f_u_dadda_cla32_fa134_and1 = f_u_dadda_cla32_fa134_xor0 & f_u_dadda_cla32_fa127_xor1;
  assign f_u_dadda_cla32_fa134_or0 = f_u_dadda_cla32_fa134_and0 | f_u_dadda_cla32_fa134_and1;
  assign f_u_dadda_cla32_ha20_xor0 = f_u_dadda_cla32_fa128_xor1 ^ f_u_dadda_cla32_fa129_xor1;
  assign f_u_dadda_cla32_ha20_and0 = f_u_dadda_cla32_fa128_xor1 & f_u_dadda_cla32_fa129_xor1;
  assign f_u_dadda_cla32_fa135_xor0 = f_u_dadda_cla32_ha20_and0 ^ f_u_dadda_cla32_fa134_or0;
  assign f_u_dadda_cla32_fa135_and0 = f_u_dadda_cla32_ha20_and0 & f_u_dadda_cla32_fa134_or0;
  assign f_u_dadda_cla32_fa135_xor1 = f_u_dadda_cla32_fa135_xor0 ^ f_u_dadda_cla32_fa133_or0;
  assign f_u_dadda_cla32_fa135_and1 = f_u_dadda_cla32_fa135_xor0 & f_u_dadda_cla32_fa133_or0;
  assign f_u_dadda_cla32_fa135_or0 = f_u_dadda_cla32_fa135_and0 | f_u_dadda_cla32_fa135_and1;
  assign f_u_dadda_cla32_fa136_xor0 = f_u_dadda_cla32_fa132_or0 ^ f_u_dadda_cla32_fa131_or0;
  assign f_u_dadda_cla32_fa136_and0 = f_u_dadda_cla32_fa132_or0 & f_u_dadda_cla32_fa131_or0;
  assign f_u_dadda_cla32_fa136_xor1 = f_u_dadda_cla32_fa136_xor0 ^ f_u_dadda_cla32_fa130_or0;
  assign f_u_dadda_cla32_fa136_and1 = f_u_dadda_cla32_fa136_xor0 & f_u_dadda_cla32_fa130_or0;
  assign f_u_dadda_cla32_fa136_or0 = f_u_dadda_cla32_fa136_and0 | f_u_dadda_cla32_fa136_and1;
  assign f_u_dadda_cla32_fa137_xor0 = f_u_dadda_cla32_fa129_or0 ^ f_u_dadda_cla32_fa128_or0;
  assign f_u_dadda_cla32_fa137_and0 = f_u_dadda_cla32_fa129_or0 & f_u_dadda_cla32_fa128_or0;
  assign f_u_dadda_cla32_fa137_xor1 = f_u_dadda_cla32_fa137_xor0 ^ f_u_dadda_cla32_fa127_or0;
  assign f_u_dadda_cla32_fa137_and1 = f_u_dadda_cla32_fa137_xor0 & f_u_dadda_cla32_fa127_or0;
  assign f_u_dadda_cla32_fa137_or0 = f_u_dadda_cla32_fa137_and0 | f_u_dadda_cla32_fa137_and1;
  assign f_u_dadda_cla32_fa138_xor0 = f_u_dadda_cla32_fa126_or0 ^ f_u_dadda_cla32_fa125_or0;
  assign f_u_dadda_cla32_fa138_and0 = f_u_dadda_cla32_fa126_or0 & f_u_dadda_cla32_fa125_or0;
  assign f_u_dadda_cla32_fa138_xor1 = f_u_dadda_cla32_fa138_xor0 ^ f_u_dadda_cla32_fa124_or0;
  assign f_u_dadda_cla32_fa138_and1 = f_u_dadda_cla32_fa138_xor0 & f_u_dadda_cla32_fa124_or0;
  assign f_u_dadda_cla32_fa138_or0 = f_u_dadda_cla32_fa138_and0 | f_u_dadda_cla32_fa138_and1;
  assign f_u_dadda_cla32_fa139_xor0 = f_u_dadda_cla32_fa123_or0 ^ f_u_dadda_cla32_fa122_or0;
  assign f_u_dadda_cla32_fa139_and0 = f_u_dadda_cla32_fa123_or0 & f_u_dadda_cla32_fa122_or0;
  assign f_u_dadda_cla32_fa139_xor1 = f_u_dadda_cla32_fa139_xor0 ^ f_u_dadda_cla32_fa121_or0;
  assign f_u_dadda_cla32_fa139_and1 = f_u_dadda_cla32_fa139_xor0 & f_u_dadda_cla32_fa121_or0;
  assign f_u_dadda_cla32_fa139_or0 = f_u_dadda_cla32_fa139_and0 | f_u_dadda_cla32_fa139_and1;
  assign f_u_dadda_cla32_and_22_0 = a[22] & b[0];
  assign f_u_dadda_cla32_and_21_1 = a[21] & b[1];
  assign f_u_dadda_cla32_fa140_xor0 = f_u_dadda_cla32_fa120_or0 ^ f_u_dadda_cla32_and_22_0;
  assign f_u_dadda_cla32_fa140_and0 = f_u_dadda_cla32_fa120_or0 & f_u_dadda_cla32_and_22_0;
  assign f_u_dadda_cla32_fa140_xor1 = f_u_dadda_cla32_fa140_xor0 ^ f_u_dadda_cla32_and_21_1;
  assign f_u_dadda_cla32_fa140_and1 = f_u_dadda_cla32_fa140_xor0 & f_u_dadda_cla32_and_21_1;
  assign f_u_dadda_cla32_fa140_or0 = f_u_dadda_cla32_fa140_and0 | f_u_dadda_cla32_fa140_and1;
  assign f_u_dadda_cla32_and_20_2 = a[20] & b[2];
  assign f_u_dadda_cla32_and_19_3 = a[19] & b[3];
  assign f_u_dadda_cla32_and_18_4 = a[18] & b[4];
  assign f_u_dadda_cla32_fa141_xor0 = f_u_dadda_cla32_and_20_2 ^ f_u_dadda_cla32_and_19_3;
  assign f_u_dadda_cla32_fa141_and0 = f_u_dadda_cla32_and_20_2 & f_u_dadda_cla32_and_19_3;
  assign f_u_dadda_cla32_fa141_xor1 = f_u_dadda_cla32_fa141_xor0 ^ f_u_dadda_cla32_and_18_4;
  assign f_u_dadda_cla32_fa141_and1 = f_u_dadda_cla32_fa141_xor0 & f_u_dadda_cla32_and_18_4;
  assign f_u_dadda_cla32_fa141_or0 = f_u_dadda_cla32_fa141_and0 | f_u_dadda_cla32_fa141_and1;
  assign f_u_dadda_cla32_and_17_5 = a[17] & b[5];
  assign f_u_dadda_cla32_and_16_6 = a[16] & b[6];
  assign f_u_dadda_cla32_and_15_7 = a[15] & b[7];
  assign f_u_dadda_cla32_fa142_xor0 = f_u_dadda_cla32_and_17_5 ^ f_u_dadda_cla32_and_16_6;
  assign f_u_dadda_cla32_fa142_and0 = f_u_dadda_cla32_and_17_5 & f_u_dadda_cla32_and_16_6;
  assign f_u_dadda_cla32_fa142_xor1 = f_u_dadda_cla32_fa142_xor0 ^ f_u_dadda_cla32_and_15_7;
  assign f_u_dadda_cla32_fa142_and1 = f_u_dadda_cla32_fa142_xor0 & f_u_dadda_cla32_and_15_7;
  assign f_u_dadda_cla32_fa142_or0 = f_u_dadda_cla32_fa142_and0 | f_u_dadda_cla32_fa142_and1;
  assign f_u_dadda_cla32_and_14_8 = a[14] & b[8];
  assign f_u_dadda_cla32_and_13_9 = a[13] & b[9];
  assign f_u_dadda_cla32_and_12_10 = a[12] & b[10];
  assign f_u_dadda_cla32_fa143_xor0 = f_u_dadda_cla32_and_14_8 ^ f_u_dadda_cla32_and_13_9;
  assign f_u_dadda_cla32_fa143_and0 = f_u_dadda_cla32_and_14_8 & f_u_dadda_cla32_and_13_9;
  assign f_u_dadda_cla32_fa143_xor1 = f_u_dadda_cla32_fa143_xor0 ^ f_u_dadda_cla32_and_12_10;
  assign f_u_dadda_cla32_fa143_and1 = f_u_dadda_cla32_fa143_xor0 & f_u_dadda_cla32_and_12_10;
  assign f_u_dadda_cla32_fa143_or0 = f_u_dadda_cla32_fa143_and0 | f_u_dadda_cla32_fa143_and1;
  assign f_u_dadda_cla32_and_11_11 = a[11] & b[11];
  assign f_u_dadda_cla32_and_10_12 = a[10] & b[12];
  assign f_u_dadda_cla32_and_9_13 = a[9] & b[13];
  assign f_u_dadda_cla32_fa144_xor0 = f_u_dadda_cla32_and_11_11 ^ f_u_dadda_cla32_and_10_12;
  assign f_u_dadda_cla32_fa144_and0 = f_u_dadda_cla32_and_11_11 & f_u_dadda_cla32_and_10_12;
  assign f_u_dadda_cla32_fa144_xor1 = f_u_dadda_cla32_fa144_xor0 ^ f_u_dadda_cla32_and_9_13;
  assign f_u_dadda_cla32_fa144_and1 = f_u_dadda_cla32_fa144_xor0 & f_u_dadda_cla32_and_9_13;
  assign f_u_dadda_cla32_fa144_or0 = f_u_dadda_cla32_fa144_and0 | f_u_dadda_cla32_fa144_and1;
  assign f_u_dadda_cla32_and_8_14 = a[8] & b[14];
  assign f_u_dadda_cla32_and_7_15 = a[7] & b[15];
  assign f_u_dadda_cla32_and_6_16 = a[6] & b[16];
  assign f_u_dadda_cla32_fa145_xor0 = f_u_dadda_cla32_and_8_14 ^ f_u_dadda_cla32_and_7_15;
  assign f_u_dadda_cla32_fa145_and0 = f_u_dadda_cla32_and_8_14 & f_u_dadda_cla32_and_7_15;
  assign f_u_dadda_cla32_fa145_xor1 = f_u_dadda_cla32_fa145_xor0 ^ f_u_dadda_cla32_and_6_16;
  assign f_u_dadda_cla32_fa145_and1 = f_u_dadda_cla32_fa145_xor0 & f_u_dadda_cla32_and_6_16;
  assign f_u_dadda_cla32_fa145_or0 = f_u_dadda_cla32_fa145_and0 | f_u_dadda_cla32_fa145_and1;
  assign f_u_dadda_cla32_and_5_17 = a[5] & b[17];
  assign f_u_dadda_cla32_and_4_18 = a[4] & b[18];
  assign f_u_dadda_cla32_and_3_19 = a[3] & b[19];
  assign f_u_dadda_cla32_fa146_xor0 = f_u_dadda_cla32_and_5_17 ^ f_u_dadda_cla32_and_4_18;
  assign f_u_dadda_cla32_fa146_and0 = f_u_dadda_cla32_and_5_17 & f_u_dadda_cla32_and_4_18;
  assign f_u_dadda_cla32_fa146_xor1 = f_u_dadda_cla32_fa146_xor0 ^ f_u_dadda_cla32_and_3_19;
  assign f_u_dadda_cla32_fa146_and1 = f_u_dadda_cla32_fa146_xor0 & f_u_dadda_cla32_and_3_19;
  assign f_u_dadda_cla32_fa146_or0 = f_u_dadda_cla32_fa146_and0 | f_u_dadda_cla32_fa146_and1;
  assign f_u_dadda_cla32_and_2_20 = a[2] & b[20];
  assign f_u_dadda_cla32_and_1_21 = a[1] & b[21];
  assign f_u_dadda_cla32_and_0_22 = a[0] & b[22];
  assign f_u_dadda_cla32_fa147_xor0 = f_u_dadda_cla32_and_2_20 ^ f_u_dadda_cla32_and_1_21;
  assign f_u_dadda_cla32_fa147_and0 = f_u_dadda_cla32_and_2_20 & f_u_dadda_cla32_and_1_21;
  assign f_u_dadda_cla32_fa147_xor1 = f_u_dadda_cla32_fa147_xor0 ^ f_u_dadda_cla32_and_0_22;
  assign f_u_dadda_cla32_fa147_and1 = f_u_dadda_cla32_fa147_xor0 & f_u_dadda_cla32_and_0_22;
  assign f_u_dadda_cla32_fa147_or0 = f_u_dadda_cla32_fa147_and0 | f_u_dadda_cla32_fa147_and1;
  assign f_u_dadda_cla32_fa148_xor0 = f_u_dadda_cla32_fa135_xor1 ^ f_u_dadda_cla32_fa136_xor1;
  assign f_u_dadda_cla32_fa148_and0 = f_u_dadda_cla32_fa135_xor1 & f_u_dadda_cla32_fa136_xor1;
  assign f_u_dadda_cla32_fa148_xor1 = f_u_dadda_cla32_fa148_xor0 ^ f_u_dadda_cla32_fa137_xor1;
  assign f_u_dadda_cla32_fa148_and1 = f_u_dadda_cla32_fa148_xor0 & f_u_dadda_cla32_fa137_xor1;
  assign f_u_dadda_cla32_fa148_or0 = f_u_dadda_cla32_fa148_and0 | f_u_dadda_cla32_fa148_and1;
  assign f_u_dadda_cla32_fa149_xor0 = f_u_dadda_cla32_fa138_xor1 ^ f_u_dadda_cla32_fa139_xor1;
  assign f_u_dadda_cla32_fa149_and0 = f_u_dadda_cla32_fa138_xor1 & f_u_dadda_cla32_fa139_xor1;
  assign f_u_dadda_cla32_fa149_xor1 = f_u_dadda_cla32_fa149_xor0 ^ f_u_dadda_cla32_fa140_xor1;
  assign f_u_dadda_cla32_fa149_and1 = f_u_dadda_cla32_fa149_xor0 & f_u_dadda_cla32_fa140_xor1;
  assign f_u_dadda_cla32_fa149_or0 = f_u_dadda_cla32_fa149_and0 | f_u_dadda_cla32_fa149_and1;
  assign f_u_dadda_cla32_fa150_xor0 = f_u_dadda_cla32_fa141_xor1 ^ f_u_dadda_cla32_fa142_xor1;
  assign f_u_dadda_cla32_fa150_and0 = f_u_dadda_cla32_fa141_xor1 & f_u_dadda_cla32_fa142_xor1;
  assign f_u_dadda_cla32_fa150_xor1 = f_u_dadda_cla32_fa150_xor0 ^ f_u_dadda_cla32_fa143_xor1;
  assign f_u_dadda_cla32_fa150_and1 = f_u_dadda_cla32_fa150_xor0 & f_u_dadda_cla32_fa143_xor1;
  assign f_u_dadda_cla32_fa150_or0 = f_u_dadda_cla32_fa150_and0 | f_u_dadda_cla32_fa150_and1;
  assign f_u_dadda_cla32_ha21_xor0 = f_u_dadda_cla32_fa144_xor1 ^ f_u_dadda_cla32_fa145_xor1;
  assign f_u_dadda_cla32_ha21_and0 = f_u_dadda_cla32_fa144_xor1 & f_u_dadda_cla32_fa145_xor1;
  assign f_u_dadda_cla32_fa151_xor0 = f_u_dadda_cla32_ha21_and0 ^ f_u_dadda_cla32_fa150_or0;
  assign f_u_dadda_cla32_fa151_and0 = f_u_dadda_cla32_ha21_and0 & f_u_dadda_cla32_fa150_or0;
  assign f_u_dadda_cla32_fa151_xor1 = f_u_dadda_cla32_fa151_xor0 ^ f_u_dadda_cla32_fa149_or0;
  assign f_u_dadda_cla32_fa151_and1 = f_u_dadda_cla32_fa151_xor0 & f_u_dadda_cla32_fa149_or0;
  assign f_u_dadda_cla32_fa151_or0 = f_u_dadda_cla32_fa151_and0 | f_u_dadda_cla32_fa151_and1;
  assign f_u_dadda_cla32_fa152_xor0 = f_u_dadda_cla32_fa148_or0 ^ f_u_dadda_cla32_fa147_or0;
  assign f_u_dadda_cla32_fa152_and0 = f_u_dadda_cla32_fa148_or0 & f_u_dadda_cla32_fa147_or0;
  assign f_u_dadda_cla32_fa152_xor1 = f_u_dadda_cla32_fa152_xor0 ^ f_u_dadda_cla32_fa146_or0;
  assign f_u_dadda_cla32_fa152_and1 = f_u_dadda_cla32_fa152_xor0 & f_u_dadda_cla32_fa146_or0;
  assign f_u_dadda_cla32_fa152_or0 = f_u_dadda_cla32_fa152_and0 | f_u_dadda_cla32_fa152_and1;
  assign f_u_dadda_cla32_fa153_xor0 = f_u_dadda_cla32_fa145_or0 ^ f_u_dadda_cla32_fa144_or0;
  assign f_u_dadda_cla32_fa153_and0 = f_u_dadda_cla32_fa145_or0 & f_u_dadda_cla32_fa144_or0;
  assign f_u_dadda_cla32_fa153_xor1 = f_u_dadda_cla32_fa153_xor0 ^ f_u_dadda_cla32_fa143_or0;
  assign f_u_dadda_cla32_fa153_and1 = f_u_dadda_cla32_fa153_xor0 & f_u_dadda_cla32_fa143_or0;
  assign f_u_dadda_cla32_fa153_or0 = f_u_dadda_cla32_fa153_and0 | f_u_dadda_cla32_fa153_and1;
  assign f_u_dadda_cla32_fa154_xor0 = f_u_dadda_cla32_fa142_or0 ^ f_u_dadda_cla32_fa141_or0;
  assign f_u_dadda_cla32_fa154_and0 = f_u_dadda_cla32_fa142_or0 & f_u_dadda_cla32_fa141_or0;
  assign f_u_dadda_cla32_fa154_xor1 = f_u_dadda_cla32_fa154_xor0 ^ f_u_dadda_cla32_fa140_or0;
  assign f_u_dadda_cla32_fa154_and1 = f_u_dadda_cla32_fa154_xor0 & f_u_dadda_cla32_fa140_or0;
  assign f_u_dadda_cla32_fa154_or0 = f_u_dadda_cla32_fa154_and0 | f_u_dadda_cla32_fa154_and1;
  assign f_u_dadda_cla32_fa155_xor0 = f_u_dadda_cla32_fa139_or0 ^ f_u_dadda_cla32_fa138_or0;
  assign f_u_dadda_cla32_fa155_and0 = f_u_dadda_cla32_fa139_or0 & f_u_dadda_cla32_fa138_or0;
  assign f_u_dadda_cla32_fa155_xor1 = f_u_dadda_cla32_fa155_xor0 ^ f_u_dadda_cla32_fa137_or0;
  assign f_u_dadda_cla32_fa155_and1 = f_u_dadda_cla32_fa155_xor0 & f_u_dadda_cla32_fa137_or0;
  assign f_u_dadda_cla32_fa155_or0 = f_u_dadda_cla32_fa155_and0 | f_u_dadda_cla32_fa155_and1;
  assign f_u_dadda_cla32_and_23_0 = a[23] & b[0];
  assign f_u_dadda_cla32_fa156_xor0 = f_u_dadda_cla32_fa136_or0 ^ f_u_dadda_cla32_fa135_or0;
  assign f_u_dadda_cla32_fa156_and0 = f_u_dadda_cla32_fa136_or0 & f_u_dadda_cla32_fa135_or0;
  assign f_u_dadda_cla32_fa156_xor1 = f_u_dadda_cla32_fa156_xor0 ^ f_u_dadda_cla32_and_23_0;
  assign f_u_dadda_cla32_fa156_and1 = f_u_dadda_cla32_fa156_xor0 & f_u_dadda_cla32_and_23_0;
  assign f_u_dadda_cla32_fa156_or0 = f_u_dadda_cla32_fa156_and0 | f_u_dadda_cla32_fa156_and1;
  assign f_u_dadda_cla32_and_22_1 = a[22] & b[1];
  assign f_u_dadda_cla32_and_21_2 = a[21] & b[2];
  assign f_u_dadda_cla32_and_20_3 = a[20] & b[3];
  assign f_u_dadda_cla32_fa157_xor0 = f_u_dadda_cla32_and_22_1 ^ f_u_dadda_cla32_and_21_2;
  assign f_u_dadda_cla32_fa157_and0 = f_u_dadda_cla32_and_22_1 & f_u_dadda_cla32_and_21_2;
  assign f_u_dadda_cla32_fa157_xor1 = f_u_dadda_cla32_fa157_xor0 ^ f_u_dadda_cla32_and_20_3;
  assign f_u_dadda_cla32_fa157_and1 = f_u_dadda_cla32_fa157_xor0 & f_u_dadda_cla32_and_20_3;
  assign f_u_dadda_cla32_fa157_or0 = f_u_dadda_cla32_fa157_and0 | f_u_dadda_cla32_fa157_and1;
  assign f_u_dadda_cla32_and_19_4 = a[19] & b[4];
  assign f_u_dadda_cla32_and_18_5 = a[18] & b[5];
  assign f_u_dadda_cla32_and_17_6 = a[17] & b[6];
  assign f_u_dadda_cla32_fa158_xor0 = f_u_dadda_cla32_and_19_4 ^ f_u_dadda_cla32_and_18_5;
  assign f_u_dadda_cla32_fa158_and0 = f_u_dadda_cla32_and_19_4 & f_u_dadda_cla32_and_18_5;
  assign f_u_dadda_cla32_fa158_xor1 = f_u_dadda_cla32_fa158_xor0 ^ f_u_dadda_cla32_and_17_6;
  assign f_u_dadda_cla32_fa158_and1 = f_u_dadda_cla32_fa158_xor0 & f_u_dadda_cla32_and_17_6;
  assign f_u_dadda_cla32_fa158_or0 = f_u_dadda_cla32_fa158_and0 | f_u_dadda_cla32_fa158_and1;
  assign f_u_dadda_cla32_and_16_7 = a[16] & b[7];
  assign f_u_dadda_cla32_and_15_8 = a[15] & b[8];
  assign f_u_dadda_cla32_and_14_9 = a[14] & b[9];
  assign f_u_dadda_cla32_fa159_xor0 = f_u_dadda_cla32_and_16_7 ^ f_u_dadda_cla32_and_15_8;
  assign f_u_dadda_cla32_fa159_and0 = f_u_dadda_cla32_and_16_7 & f_u_dadda_cla32_and_15_8;
  assign f_u_dadda_cla32_fa159_xor1 = f_u_dadda_cla32_fa159_xor0 ^ f_u_dadda_cla32_and_14_9;
  assign f_u_dadda_cla32_fa159_and1 = f_u_dadda_cla32_fa159_xor0 & f_u_dadda_cla32_and_14_9;
  assign f_u_dadda_cla32_fa159_or0 = f_u_dadda_cla32_fa159_and0 | f_u_dadda_cla32_fa159_and1;
  assign f_u_dadda_cla32_and_13_10 = a[13] & b[10];
  assign f_u_dadda_cla32_and_12_11 = a[12] & b[11];
  assign f_u_dadda_cla32_and_11_12 = a[11] & b[12];
  assign f_u_dadda_cla32_fa160_xor0 = f_u_dadda_cla32_and_13_10 ^ f_u_dadda_cla32_and_12_11;
  assign f_u_dadda_cla32_fa160_and0 = f_u_dadda_cla32_and_13_10 & f_u_dadda_cla32_and_12_11;
  assign f_u_dadda_cla32_fa160_xor1 = f_u_dadda_cla32_fa160_xor0 ^ f_u_dadda_cla32_and_11_12;
  assign f_u_dadda_cla32_fa160_and1 = f_u_dadda_cla32_fa160_xor0 & f_u_dadda_cla32_and_11_12;
  assign f_u_dadda_cla32_fa160_or0 = f_u_dadda_cla32_fa160_and0 | f_u_dadda_cla32_fa160_and1;
  assign f_u_dadda_cla32_and_10_13 = a[10] & b[13];
  assign f_u_dadda_cla32_and_9_14 = a[9] & b[14];
  assign f_u_dadda_cla32_and_8_15 = a[8] & b[15];
  assign f_u_dadda_cla32_fa161_xor0 = f_u_dadda_cla32_and_10_13 ^ f_u_dadda_cla32_and_9_14;
  assign f_u_dadda_cla32_fa161_and0 = f_u_dadda_cla32_and_10_13 & f_u_dadda_cla32_and_9_14;
  assign f_u_dadda_cla32_fa161_xor1 = f_u_dadda_cla32_fa161_xor0 ^ f_u_dadda_cla32_and_8_15;
  assign f_u_dadda_cla32_fa161_and1 = f_u_dadda_cla32_fa161_xor0 & f_u_dadda_cla32_and_8_15;
  assign f_u_dadda_cla32_fa161_or0 = f_u_dadda_cla32_fa161_and0 | f_u_dadda_cla32_fa161_and1;
  assign f_u_dadda_cla32_and_7_16 = a[7] & b[16];
  assign f_u_dadda_cla32_and_6_17 = a[6] & b[17];
  assign f_u_dadda_cla32_and_5_18 = a[5] & b[18];
  assign f_u_dadda_cla32_fa162_xor0 = f_u_dadda_cla32_and_7_16 ^ f_u_dadda_cla32_and_6_17;
  assign f_u_dadda_cla32_fa162_and0 = f_u_dadda_cla32_and_7_16 & f_u_dadda_cla32_and_6_17;
  assign f_u_dadda_cla32_fa162_xor1 = f_u_dadda_cla32_fa162_xor0 ^ f_u_dadda_cla32_and_5_18;
  assign f_u_dadda_cla32_fa162_and1 = f_u_dadda_cla32_fa162_xor0 & f_u_dadda_cla32_and_5_18;
  assign f_u_dadda_cla32_fa162_or0 = f_u_dadda_cla32_fa162_and0 | f_u_dadda_cla32_fa162_and1;
  assign f_u_dadda_cla32_and_4_19 = a[4] & b[19];
  assign f_u_dadda_cla32_and_3_20 = a[3] & b[20];
  assign f_u_dadda_cla32_and_2_21 = a[2] & b[21];
  assign f_u_dadda_cla32_fa163_xor0 = f_u_dadda_cla32_and_4_19 ^ f_u_dadda_cla32_and_3_20;
  assign f_u_dadda_cla32_fa163_and0 = f_u_dadda_cla32_and_4_19 & f_u_dadda_cla32_and_3_20;
  assign f_u_dadda_cla32_fa163_xor1 = f_u_dadda_cla32_fa163_xor0 ^ f_u_dadda_cla32_and_2_21;
  assign f_u_dadda_cla32_fa163_and1 = f_u_dadda_cla32_fa163_xor0 & f_u_dadda_cla32_and_2_21;
  assign f_u_dadda_cla32_fa163_or0 = f_u_dadda_cla32_fa163_and0 | f_u_dadda_cla32_fa163_and1;
  assign f_u_dadda_cla32_and_1_22 = a[1] & b[22];
  assign f_u_dadda_cla32_and_0_23 = a[0] & b[23];
  assign f_u_dadda_cla32_fa164_xor0 = f_u_dadda_cla32_and_1_22 ^ f_u_dadda_cla32_and_0_23;
  assign f_u_dadda_cla32_fa164_and0 = f_u_dadda_cla32_and_1_22 & f_u_dadda_cla32_and_0_23;
  assign f_u_dadda_cla32_fa164_xor1 = f_u_dadda_cla32_fa164_xor0 ^ f_u_dadda_cla32_fa151_xor1;
  assign f_u_dadda_cla32_fa164_and1 = f_u_dadda_cla32_fa164_xor0 & f_u_dadda_cla32_fa151_xor1;
  assign f_u_dadda_cla32_fa164_or0 = f_u_dadda_cla32_fa164_and0 | f_u_dadda_cla32_fa164_and1;
  assign f_u_dadda_cla32_fa165_xor0 = f_u_dadda_cla32_fa152_xor1 ^ f_u_dadda_cla32_fa153_xor1;
  assign f_u_dadda_cla32_fa165_and0 = f_u_dadda_cla32_fa152_xor1 & f_u_dadda_cla32_fa153_xor1;
  assign f_u_dadda_cla32_fa165_xor1 = f_u_dadda_cla32_fa165_xor0 ^ f_u_dadda_cla32_fa154_xor1;
  assign f_u_dadda_cla32_fa165_and1 = f_u_dadda_cla32_fa165_xor0 & f_u_dadda_cla32_fa154_xor1;
  assign f_u_dadda_cla32_fa165_or0 = f_u_dadda_cla32_fa165_and0 | f_u_dadda_cla32_fa165_and1;
  assign f_u_dadda_cla32_fa166_xor0 = f_u_dadda_cla32_fa155_xor1 ^ f_u_dadda_cla32_fa156_xor1;
  assign f_u_dadda_cla32_fa166_and0 = f_u_dadda_cla32_fa155_xor1 & f_u_dadda_cla32_fa156_xor1;
  assign f_u_dadda_cla32_fa166_xor1 = f_u_dadda_cla32_fa166_xor0 ^ f_u_dadda_cla32_fa157_xor1;
  assign f_u_dadda_cla32_fa166_and1 = f_u_dadda_cla32_fa166_xor0 & f_u_dadda_cla32_fa157_xor1;
  assign f_u_dadda_cla32_fa166_or0 = f_u_dadda_cla32_fa166_and0 | f_u_dadda_cla32_fa166_and1;
  assign f_u_dadda_cla32_fa167_xor0 = f_u_dadda_cla32_fa158_xor1 ^ f_u_dadda_cla32_fa159_xor1;
  assign f_u_dadda_cla32_fa167_and0 = f_u_dadda_cla32_fa158_xor1 & f_u_dadda_cla32_fa159_xor1;
  assign f_u_dadda_cla32_fa167_xor1 = f_u_dadda_cla32_fa167_xor0 ^ f_u_dadda_cla32_fa160_xor1;
  assign f_u_dadda_cla32_fa167_and1 = f_u_dadda_cla32_fa167_xor0 & f_u_dadda_cla32_fa160_xor1;
  assign f_u_dadda_cla32_fa167_or0 = f_u_dadda_cla32_fa167_and0 | f_u_dadda_cla32_fa167_and1;
  assign f_u_dadda_cla32_ha22_xor0 = f_u_dadda_cla32_fa161_xor1 ^ f_u_dadda_cla32_fa162_xor1;
  assign f_u_dadda_cla32_ha22_and0 = f_u_dadda_cla32_fa161_xor1 & f_u_dadda_cla32_fa162_xor1;
  assign f_u_dadda_cla32_fa168_xor0 = f_u_dadda_cla32_ha22_and0 ^ f_u_dadda_cla32_fa167_or0;
  assign f_u_dadda_cla32_fa168_and0 = f_u_dadda_cla32_ha22_and0 & f_u_dadda_cla32_fa167_or0;
  assign f_u_dadda_cla32_fa168_xor1 = f_u_dadda_cla32_fa168_xor0 ^ f_u_dadda_cla32_fa166_or0;
  assign f_u_dadda_cla32_fa168_and1 = f_u_dadda_cla32_fa168_xor0 & f_u_dadda_cla32_fa166_or0;
  assign f_u_dadda_cla32_fa168_or0 = f_u_dadda_cla32_fa168_and0 | f_u_dadda_cla32_fa168_and1;
  assign f_u_dadda_cla32_fa169_xor0 = f_u_dadda_cla32_fa165_or0 ^ f_u_dadda_cla32_fa164_or0;
  assign f_u_dadda_cla32_fa169_and0 = f_u_dadda_cla32_fa165_or0 & f_u_dadda_cla32_fa164_or0;
  assign f_u_dadda_cla32_fa169_xor1 = f_u_dadda_cla32_fa169_xor0 ^ f_u_dadda_cla32_fa163_or0;
  assign f_u_dadda_cla32_fa169_and1 = f_u_dadda_cla32_fa169_xor0 & f_u_dadda_cla32_fa163_or0;
  assign f_u_dadda_cla32_fa169_or0 = f_u_dadda_cla32_fa169_and0 | f_u_dadda_cla32_fa169_and1;
  assign f_u_dadda_cla32_fa170_xor0 = f_u_dadda_cla32_fa162_or0 ^ f_u_dadda_cla32_fa161_or0;
  assign f_u_dadda_cla32_fa170_and0 = f_u_dadda_cla32_fa162_or0 & f_u_dadda_cla32_fa161_or0;
  assign f_u_dadda_cla32_fa170_xor1 = f_u_dadda_cla32_fa170_xor0 ^ f_u_dadda_cla32_fa160_or0;
  assign f_u_dadda_cla32_fa170_and1 = f_u_dadda_cla32_fa170_xor0 & f_u_dadda_cla32_fa160_or0;
  assign f_u_dadda_cla32_fa170_or0 = f_u_dadda_cla32_fa170_and0 | f_u_dadda_cla32_fa170_and1;
  assign f_u_dadda_cla32_fa171_xor0 = f_u_dadda_cla32_fa159_or0 ^ f_u_dadda_cla32_fa158_or0;
  assign f_u_dadda_cla32_fa171_and0 = f_u_dadda_cla32_fa159_or0 & f_u_dadda_cla32_fa158_or0;
  assign f_u_dadda_cla32_fa171_xor1 = f_u_dadda_cla32_fa171_xor0 ^ f_u_dadda_cla32_fa157_or0;
  assign f_u_dadda_cla32_fa171_and1 = f_u_dadda_cla32_fa171_xor0 & f_u_dadda_cla32_fa157_or0;
  assign f_u_dadda_cla32_fa171_or0 = f_u_dadda_cla32_fa171_and0 | f_u_dadda_cla32_fa171_and1;
  assign f_u_dadda_cla32_fa172_xor0 = f_u_dadda_cla32_fa156_or0 ^ f_u_dadda_cla32_fa155_or0;
  assign f_u_dadda_cla32_fa172_and0 = f_u_dadda_cla32_fa156_or0 & f_u_dadda_cla32_fa155_or0;
  assign f_u_dadda_cla32_fa172_xor1 = f_u_dadda_cla32_fa172_xor0 ^ f_u_dadda_cla32_fa154_or0;
  assign f_u_dadda_cla32_fa172_and1 = f_u_dadda_cla32_fa172_xor0 & f_u_dadda_cla32_fa154_or0;
  assign f_u_dadda_cla32_fa172_or0 = f_u_dadda_cla32_fa172_and0 | f_u_dadda_cla32_fa172_and1;
  assign f_u_dadda_cla32_fa173_xor0 = f_u_dadda_cla32_fa153_or0 ^ f_u_dadda_cla32_fa152_or0;
  assign f_u_dadda_cla32_fa173_and0 = f_u_dadda_cla32_fa153_or0 & f_u_dadda_cla32_fa152_or0;
  assign f_u_dadda_cla32_fa173_xor1 = f_u_dadda_cla32_fa173_xor0 ^ f_u_dadda_cla32_fa151_or0;
  assign f_u_dadda_cla32_fa173_and1 = f_u_dadda_cla32_fa173_xor0 & f_u_dadda_cla32_fa151_or0;
  assign f_u_dadda_cla32_fa173_or0 = f_u_dadda_cla32_fa173_and0 | f_u_dadda_cla32_fa173_and1;
  assign f_u_dadda_cla32_and_24_0 = a[24] & b[0];
  assign f_u_dadda_cla32_and_23_1 = a[23] & b[1];
  assign f_u_dadda_cla32_and_22_2 = a[22] & b[2];
  assign f_u_dadda_cla32_fa174_xor0 = f_u_dadda_cla32_and_24_0 ^ f_u_dadda_cla32_and_23_1;
  assign f_u_dadda_cla32_fa174_and0 = f_u_dadda_cla32_and_24_0 & f_u_dadda_cla32_and_23_1;
  assign f_u_dadda_cla32_fa174_xor1 = f_u_dadda_cla32_fa174_xor0 ^ f_u_dadda_cla32_and_22_2;
  assign f_u_dadda_cla32_fa174_and1 = f_u_dadda_cla32_fa174_xor0 & f_u_dadda_cla32_and_22_2;
  assign f_u_dadda_cla32_fa174_or0 = f_u_dadda_cla32_fa174_and0 | f_u_dadda_cla32_fa174_and1;
  assign f_u_dadda_cla32_and_21_3 = a[21] & b[3];
  assign f_u_dadda_cla32_and_20_4 = a[20] & b[4];
  assign f_u_dadda_cla32_and_19_5 = a[19] & b[5];
  assign f_u_dadda_cla32_fa175_xor0 = f_u_dadda_cla32_and_21_3 ^ f_u_dadda_cla32_and_20_4;
  assign f_u_dadda_cla32_fa175_and0 = f_u_dadda_cla32_and_21_3 & f_u_dadda_cla32_and_20_4;
  assign f_u_dadda_cla32_fa175_xor1 = f_u_dadda_cla32_fa175_xor0 ^ f_u_dadda_cla32_and_19_5;
  assign f_u_dadda_cla32_fa175_and1 = f_u_dadda_cla32_fa175_xor0 & f_u_dadda_cla32_and_19_5;
  assign f_u_dadda_cla32_fa175_or0 = f_u_dadda_cla32_fa175_and0 | f_u_dadda_cla32_fa175_and1;
  assign f_u_dadda_cla32_and_18_6 = a[18] & b[6];
  assign f_u_dadda_cla32_and_17_7 = a[17] & b[7];
  assign f_u_dadda_cla32_and_16_8 = a[16] & b[8];
  assign f_u_dadda_cla32_fa176_xor0 = f_u_dadda_cla32_and_18_6 ^ f_u_dadda_cla32_and_17_7;
  assign f_u_dadda_cla32_fa176_and0 = f_u_dadda_cla32_and_18_6 & f_u_dadda_cla32_and_17_7;
  assign f_u_dadda_cla32_fa176_xor1 = f_u_dadda_cla32_fa176_xor0 ^ f_u_dadda_cla32_and_16_8;
  assign f_u_dadda_cla32_fa176_and1 = f_u_dadda_cla32_fa176_xor0 & f_u_dadda_cla32_and_16_8;
  assign f_u_dadda_cla32_fa176_or0 = f_u_dadda_cla32_fa176_and0 | f_u_dadda_cla32_fa176_and1;
  assign f_u_dadda_cla32_and_15_9 = a[15] & b[9];
  assign f_u_dadda_cla32_and_14_10 = a[14] & b[10];
  assign f_u_dadda_cla32_and_13_11 = a[13] & b[11];
  assign f_u_dadda_cla32_fa177_xor0 = f_u_dadda_cla32_and_15_9 ^ f_u_dadda_cla32_and_14_10;
  assign f_u_dadda_cla32_fa177_and0 = f_u_dadda_cla32_and_15_9 & f_u_dadda_cla32_and_14_10;
  assign f_u_dadda_cla32_fa177_xor1 = f_u_dadda_cla32_fa177_xor0 ^ f_u_dadda_cla32_and_13_11;
  assign f_u_dadda_cla32_fa177_and1 = f_u_dadda_cla32_fa177_xor0 & f_u_dadda_cla32_and_13_11;
  assign f_u_dadda_cla32_fa177_or0 = f_u_dadda_cla32_fa177_and0 | f_u_dadda_cla32_fa177_and1;
  assign f_u_dadda_cla32_and_12_12 = a[12] & b[12];
  assign f_u_dadda_cla32_and_11_13 = a[11] & b[13];
  assign f_u_dadda_cla32_and_10_14 = a[10] & b[14];
  assign f_u_dadda_cla32_fa178_xor0 = f_u_dadda_cla32_and_12_12 ^ f_u_dadda_cla32_and_11_13;
  assign f_u_dadda_cla32_fa178_and0 = f_u_dadda_cla32_and_12_12 & f_u_dadda_cla32_and_11_13;
  assign f_u_dadda_cla32_fa178_xor1 = f_u_dadda_cla32_fa178_xor0 ^ f_u_dadda_cla32_and_10_14;
  assign f_u_dadda_cla32_fa178_and1 = f_u_dadda_cla32_fa178_xor0 & f_u_dadda_cla32_and_10_14;
  assign f_u_dadda_cla32_fa178_or0 = f_u_dadda_cla32_fa178_and0 | f_u_dadda_cla32_fa178_and1;
  assign f_u_dadda_cla32_and_9_15 = a[9] & b[15];
  assign f_u_dadda_cla32_and_8_16 = a[8] & b[16];
  assign f_u_dadda_cla32_and_7_17 = a[7] & b[17];
  assign f_u_dadda_cla32_fa179_xor0 = f_u_dadda_cla32_and_9_15 ^ f_u_dadda_cla32_and_8_16;
  assign f_u_dadda_cla32_fa179_and0 = f_u_dadda_cla32_and_9_15 & f_u_dadda_cla32_and_8_16;
  assign f_u_dadda_cla32_fa179_xor1 = f_u_dadda_cla32_fa179_xor0 ^ f_u_dadda_cla32_and_7_17;
  assign f_u_dadda_cla32_fa179_and1 = f_u_dadda_cla32_fa179_xor0 & f_u_dadda_cla32_and_7_17;
  assign f_u_dadda_cla32_fa179_or0 = f_u_dadda_cla32_fa179_and0 | f_u_dadda_cla32_fa179_and1;
  assign f_u_dadda_cla32_and_6_18 = a[6] & b[18];
  assign f_u_dadda_cla32_and_5_19 = a[5] & b[19];
  assign f_u_dadda_cla32_and_4_20 = a[4] & b[20];
  assign f_u_dadda_cla32_fa180_xor0 = f_u_dadda_cla32_and_6_18 ^ f_u_dadda_cla32_and_5_19;
  assign f_u_dadda_cla32_fa180_and0 = f_u_dadda_cla32_and_6_18 & f_u_dadda_cla32_and_5_19;
  assign f_u_dadda_cla32_fa180_xor1 = f_u_dadda_cla32_fa180_xor0 ^ f_u_dadda_cla32_and_4_20;
  assign f_u_dadda_cla32_fa180_and1 = f_u_dadda_cla32_fa180_xor0 & f_u_dadda_cla32_and_4_20;
  assign f_u_dadda_cla32_fa180_or0 = f_u_dadda_cla32_fa180_and0 | f_u_dadda_cla32_fa180_and1;
  assign f_u_dadda_cla32_and_3_21 = a[3] & b[21];
  assign f_u_dadda_cla32_and_2_22 = a[2] & b[22];
  assign f_u_dadda_cla32_and_1_23 = a[1] & b[23];
  assign f_u_dadda_cla32_fa181_xor0 = f_u_dadda_cla32_and_3_21 ^ f_u_dadda_cla32_and_2_22;
  assign f_u_dadda_cla32_fa181_and0 = f_u_dadda_cla32_and_3_21 & f_u_dadda_cla32_and_2_22;
  assign f_u_dadda_cla32_fa181_xor1 = f_u_dadda_cla32_fa181_xor0 ^ f_u_dadda_cla32_and_1_23;
  assign f_u_dadda_cla32_fa181_and1 = f_u_dadda_cla32_fa181_xor0 & f_u_dadda_cla32_and_1_23;
  assign f_u_dadda_cla32_fa181_or0 = f_u_dadda_cla32_fa181_and0 | f_u_dadda_cla32_fa181_and1;
  assign f_u_dadda_cla32_and_0_24 = a[0] & b[24];
  assign f_u_dadda_cla32_fa182_xor0 = f_u_dadda_cla32_and_0_24 ^ f_u_dadda_cla32_fa168_xor1;
  assign f_u_dadda_cla32_fa182_and0 = f_u_dadda_cla32_and_0_24 & f_u_dadda_cla32_fa168_xor1;
  assign f_u_dadda_cla32_fa182_xor1 = f_u_dadda_cla32_fa182_xor0 ^ f_u_dadda_cla32_fa169_xor1;
  assign f_u_dadda_cla32_fa182_and1 = f_u_dadda_cla32_fa182_xor0 & f_u_dadda_cla32_fa169_xor1;
  assign f_u_dadda_cla32_fa182_or0 = f_u_dadda_cla32_fa182_and0 | f_u_dadda_cla32_fa182_and1;
  assign f_u_dadda_cla32_fa183_xor0 = f_u_dadda_cla32_fa170_xor1 ^ f_u_dadda_cla32_fa171_xor1;
  assign f_u_dadda_cla32_fa183_and0 = f_u_dadda_cla32_fa170_xor1 & f_u_dadda_cla32_fa171_xor1;
  assign f_u_dadda_cla32_fa183_xor1 = f_u_dadda_cla32_fa183_xor0 ^ f_u_dadda_cla32_fa172_xor1;
  assign f_u_dadda_cla32_fa183_and1 = f_u_dadda_cla32_fa183_xor0 & f_u_dadda_cla32_fa172_xor1;
  assign f_u_dadda_cla32_fa183_or0 = f_u_dadda_cla32_fa183_and0 | f_u_dadda_cla32_fa183_and1;
  assign f_u_dadda_cla32_fa184_xor0 = f_u_dadda_cla32_fa173_xor1 ^ f_u_dadda_cla32_fa174_xor1;
  assign f_u_dadda_cla32_fa184_and0 = f_u_dadda_cla32_fa173_xor1 & f_u_dadda_cla32_fa174_xor1;
  assign f_u_dadda_cla32_fa184_xor1 = f_u_dadda_cla32_fa184_xor0 ^ f_u_dadda_cla32_fa175_xor1;
  assign f_u_dadda_cla32_fa184_and1 = f_u_dadda_cla32_fa184_xor0 & f_u_dadda_cla32_fa175_xor1;
  assign f_u_dadda_cla32_fa184_or0 = f_u_dadda_cla32_fa184_and0 | f_u_dadda_cla32_fa184_and1;
  assign f_u_dadda_cla32_fa185_xor0 = f_u_dadda_cla32_fa176_xor1 ^ f_u_dadda_cla32_fa177_xor1;
  assign f_u_dadda_cla32_fa185_and0 = f_u_dadda_cla32_fa176_xor1 & f_u_dadda_cla32_fa177_xor1;
  assign f_u_dadda_cla32_fa185_xor1 = f_u_dadda_cla32_fa185_xor0 ^ f_u_dadda_cla32_fa178_xor1;
  assign f_u_dadda_cla32_fa185_and1 = f_u_dadda_cla32_fa185_xor0 & f_u_dadda_cla32_fa178_xor1;
  assign f_u_dadda_cla32_fa185_or0 = f_u_dadda_cla32_fa185_and0 | f_u_dadda_cla32_fa185_and1;
  assign f_u_dadda_cla32_ha23_xor0 = f_u_dadda_cla32_fa179_xor1 ^ f_u_dadda_cla32_fa180_xor1;
  assign f_u_dadda_cla32_ha23_and0 = f_u_dadda_cla32_fa179_xor1 & f_u_dadda_cla32_fa180_xor1;
  assign f_u_dadda_cla32_fa186_xor0 = f_u_dadda_cla32_ha23_and0 ^ f_u_dadda_cla32_fa185_or0;
  assign f_u_dadda_cla32_fa186_and0 = f_u_dadda_cla32_ha23_and0 & f_u_dadda_cla32_fa185_or0;
  assign f_u_dadda_cla32_fa186_xor1 = f_u_dadda_cla32_fa186_xor0 ^ f_u_dadda_cla32_fa184_or0;
  assign f_u_dadda_cla32_fa186_and1 = f_u_dadda_cla32_fa186_xor0 & f_u_dadda_cla32_fa184_or0;
  assign f_u_dadda_cla32_fa186_or0 = f_u_dadda_cla32_fa186_and0 | f_u_dadda_cla32_fa186_and1;
  assign f_u_dadda_cla32_fa187_xor0 = f_u_dadda_cla32_fa183_or0 ^ f_u_dadda_cla32_fa182_or0;
  assign f_u_dadda_cla32_fa187_and0 = f_u_dadda_cla32_fa183_or0 & f_u_dadda_cla32_fa182_or0;
  assign f_u_dadda_cla32_fa187_xor1 = f_u_dadda_cla32_fa187_xor0 ^ f_u_dadda_cla32_fa181_or0;
  assign f_u_dadda_cla32_fa187_and1 = f_u_dadda_cla32_fa187_xor0 & f_u_dadda_cla32_fa181_or0;
  assign f_u_dadda_cla32_fa187_or0 = f_u_dadda_cla32_fa187_and0 | f_u_dadda_cla32_fa187_and1;
  assign f_u_dadda_cla32_fa188_xor0 = f_u_dadda_cla32_fa180_or0 ^ f_u_dadda_cla32_fa179_or0;
  assign f_u_dadda_cla32_fa188_and0 = f_u_dadda_cla32_fa180_or0 & f_u_dadda_cla32_fa179_or0;
  assign f_u_dadda_cla32_fa188_xor1 = f_u_dadda_cla32_fa188_xor0 ^ f_u_dadda_cla32_fa178_or0;
  assign f_u_dadda_cla32_fa188_and1 = f_u_dadda_cla32_fa188_xor0 & f_u_dadda_cla32_fa178_or0;
  assign f_u_dadda_cla32_fa188_or0 = f_u_dadda_cla32_fa188_and0 | f_u_dadda_cla32_fa188_and1;
  assign f_u_dadda_cla32_fa189_xor0 = f_u_dadda_cla32_fa177_or0 ^ f_u_dadda_cla32_fa176_or0;
  assign f_u_dadda_cla32_fa189_and0 = f_u_dadda_cla32_fa177_or0 & f_u_dadda_cla32_fa176_or0;
  assign f_u_dadda_cla32_fa189_xor1 = f_u_dadda_cla32_fa189_xor0 ^ f_u_dadda_cla32_fa175_or0;
  assign f_u_dadda_cla32_fa189_and1 = f_u_dadda_cla32_fa189_xor0 & f_u_dadda_cla32_fa175_or0;
  assign f_u_dadda_cla32_fa189_or0 = f_u_dadda_cla32_fa189_and0 | f_u_dadda_cla32_fa189_and1;
  assign f_u_dadda_cla32_fa190_xor0 = f_u_dadda_cla32_fa174_or0 ^ f_u_dadda_cla32_fa173_or0;
  assign f_u_dadda_cla32_fa190_and0 = f_u_dadda_cla32_fa174_or0 & f_u_dadda_cla32_fa173_or0;
  assign f_u_dadda_cla32_fa190_xor1 = f_u_dadda_cla32_fa190_xor0 ^ f_u_dadda_cla32_fa172_or0;
  assign f_u_dadda_cla32_fa190_and1 = f_u_dadda_cla32_fa190_xor0 & f_u_dadda_cla32_fa172_or0;
  assign f_u_dadda_cla32_fa190_or0 = f_u_dadda_cla32_fa190_and0 | f_u_dadda_cla32_fa190_and1;
  assign f_u_dadda_cla32_fa191_xor0 = f_u_dadda_cla32_fa171_or0 ^ f_u_dadda_cla32_fa170_or0;
  assign f_u_dadda_cla32_fa191_and0 = f_u_dadda_cla32_fa171_or0 & f_u_dadda_cla32_fa170_or0;
  assign f_u_dadda_cla32_fa191_xor1 = f_u_dadda_cla32_fa191_xor0 ^ f_u_dadda_cla32_fa169_or0;
  assign f_u_dadda_cla32_fa191_and1 = f_u_dadda_cla32_fa191_xor0 & f_u_dadda_cla32_fa169_or0;
  assign f_u_dadda_cla32_fa191_or0 = f_u_dadda_cla32_fa191_and0 | f_u_dadda_cla32_fa191_and1;
  assign f_u_dadda_cla32_and_25_0 = a[25] & b[0];
  assign f_u_dadda_cla32_and_24_1 = a[24] & b[1];
  assign f_u_dadda_cla32_fa192_xor0 = f_u_dadda_cla32_fa168_or0 ^ f_u_dadda_cla32_and_25_0;
  assign f_u_dadda_cla32_fa192_and0 = f_u_dadda_cla32_fa168_or0 & f_u_dadda_cla32_and_25_0;
  assign f_u_dadda_cla32_fa192_xor1 = f_u_dadda_cla32_fa192_xor0 ^ f_u_dadda_cla32_and_24_1;
  assign f_u_dadda_cla32_fa192_and1 = f_u_dadda_cla32_fa192_xor0 & f_u_dadda_cla32_and_24_1;
  assign f_u_dadda_cla32_fa192_or0 = f_u_dadda_cla32_fa192_and0 | f_u_dadda_cla32_fa192_and1;
  assign f_u_dadda_cla32_and_23_2 = a[23] & b[2];
  assign f_u_dadda_cla32_and_22_3 = a[22] & b[3];
  assign f_u_dadda_cla32_and_21_4 = a[21] & b[4];
  assign f_u_dadda_cla32_fa193_xor0 = f_u_dadda_cla32_and_23_2 ^ f_u_dadda_cla32_and_22_3;
  assign f_u_dadda_cla32_fa193_and0 = f_u_dadda_cla32_and_23_2 & f_u_dadda_cla32_and_22_3;
  assign f_u_dadda_cla32_fa193_xor1 = f_u_dadda_cla32_fa193_xor0 ^ f_u_dadda_cla32_and_21_4;
  assign f_u_dadda_cla32_fa193_and1 = f_u_dadda_cla32_fa193_xor0 & f_u_dadda_cla32_and_21_4;
  assign f_u_dadda_cla32_fa193_or0 = f_u_dadda_cla32_fa193_and0 | f_u_dadda_cla32_fa193_and1;
  assign f_u_dadda_cla32_and_20_5 = a[20] & b[5];
  assign f_u_dadda_cla32_and_19_6 = a[19] & b[6];
  assign f_u_dadda_cla32_and_18_7 = a[18] & b[7];
  assign f_u_dadda_cla32_fa194_xor0 = f_u_dadda_cla32_and_20_5 ^ f_u_dadda_cla32_and_19_6;
  assign f_u_dadda_cla32_fa194_and0 = f_u_dadda_cla32_and_20_5 & f_u_dadda_cla32_and_19_6;
  assign f_u_dadda_cla32_fa194_xor1 = f_u_dadda_cla32_fa194_xor0 ^ f_u_dadda_cla32_and_18_7;
  assign f_u_dadda_cla32_fa194_and1 = f_u_dadda_cla32_fa194_xor0 & f_u_dadda_cla32_and_18_7;
  assign f_u_dadda_cla32_fa194_or0 = f_u_dadda_cla32_fa194_and0 | f_u_dadda_cla32_fa194_and1;
  assign f_u_dadda_cla32_and_17_8 = a[17] & b[8];
  assign f_u_dadda_cla32_and_16_9 = a[16] & b[9];
  assign f_u_dadda_cla32_and_15_10 = a[15] & b[10];
  assign f_u_dadda_cla32_fa195_xor0 = f_u_dadda_cla32_and_17_8 ^ f_u_dadda_cla32_and_16_9;
  assign f_u_dadda_cla32_fa195_and0 = f_u_dadda_cla32_and_17_8 & f_u_dadda_cla32_and_16_9;
  assign f_u_dadda_cla32_fa195_xor1 = f_u_dadda_cla32_fa195_xor0 ^ f_u_dadda_cla32_and_15_10;
  assign f_u_dadda_cla32_fa195_and1 = f_u_dadda_cla32_fa195_xor0 & f_u_dadda_cla32_and_15_10;
  assign f_u_dadda_cla32_fa195_or0 = f_u_dadda_cla32_fa195_and0 | f_u_dadda_cla32_fa195_and1;
  assign f_u_dadda_cla32_and_14_11 = a[14] & b[11];
  assign f_u_dadda_cla32_and_13_12 = a[13] & b[12];
  assign f_u_dadda_cla32_and_12_13 = a[12] & b[13];
  assign f_u_dadda_cla32_fa196_xor0 = f_u_dadda_cla32_and_14_11 ^ f_u_dadda_cla32_and_13_12;
  assign f_u_dadda_cla32_fa196_and0 = f_u_dadda_cla32_and_14_11 & f_u_dadda_cla32_and_13_12;
  assign f_u_dadda_cla32_fa196_xor1 = f_u_dadda_cla32_fa196_xor0 ^ f_u_dadda_cla32_and_12_13;
  assign f_u_dadda_cla32_fa196_and1 = f_u_dadda_cla32_fa196_xor0 & f_u_dadda_cla32_and_12_13;
  assign f_u_dadda_cla32_fa196_or0 = f_u_dadda_cla32_fa196_and0 | f_u_dadda_cla32_fa196_and1;
  assign f_u_dadda_cla32_and_11_14 = a[11] & b[14];
  assign f_u_dadda_cla32_and_10_15 = a[10] & b[15];
  assign f_u_dadda_cla32_and_9_16 = a[9] & b[16];
  assign f_u_dadda_cla32_fa197_xor0 = f_u_dadda_cla32_and_11_14 ^ f_u_dadda_cla32_and_10_15;
  assign f_u_dadda_cla32_fa197_and0 = f_u_dadda_cla32_and_11_14 & f_u_dadda_cla32_and_10_15;
  assign f_u_dadda_cla32_fa197_xor1 = f_u_dadda_cla32_fa197_xor0 ^ f_u_dadda_cla32_and_9_16;
  assign f_u_dadda_cla32_fa197_and1 = f_u_dadda_cla32_fa197_xor0 & f_u_dadda_cla32_and_9_16;
  assign f_u_dadda_cla32_fa197_or0 = f_u_dadda_cla32_fa197_and0 | f_u_dadda_cla32_fa197_and1;
  assign f_u_dadda_cla32_and_8_17 = a[8] & b[17];
  assign f_u_dadda_cla32_and_7_18 = a[7] & b[18];
  assign f_u_dadda_cla32_and_6_19 = a[6] & b[19];
  assign f_u_dadda_cla32_fa198_xor0 = f_u_dadda_cla32_and_8_17 ^ f_u_dadda_cla32_and_7_18;
  assign f_u_dadda_cla32_fa198_and0 = f_u_dadda_cla32_and_8_17 & f_u_dadda_cla32_and_7_18;
  assign f_u_dadda_cla32_fa198_xor1 = f_u_dadda_cla32_fa198_xor0 ^ f_u_dadda_cla32_and_6_19;
  assign f_u_dadda_cla32_fa198_and1 = f_u_dadda_cla32_fa198_xor0 & f_u_dadda_cla32_and_6_19;
  assign f_u_dadda_cla32_fa198_or0 = f_u_dadda_cla32_fa198_and0 | f_u_dadda_cla32_fa198_and1;
  assign f_u_dadda_cla32_and_5_20 = a[5] & b[20];
  assign f_u_dadda_cla32_and_4_21 = a[4] & b[21];
  assign f_u_dadda_cla32_and_3_22 = a[3] & b[22];
  assign f_u_dadda_cla32_fa199_xor0 = f_u_dadda_cla32_and_5_20 ^ f_u_dadda_cla32_and_4_21;
  assign f_u_dadda_cla32_fa199_and0 = f_u_dadda_cla32_and_5_20 & f_u_dadda_cla32_and_4_21;
  assign f_u_dadda_cla32_fa199_xor1 = f_u_dadda_cla32_fa199_xor0 ^ f_u_dadda_cla32_and_3_22;
  assign f_u_dadda_cla32_fa199_and1 = f_u_dadda_cla32_fa199_xor0 & f_u_dadda_cla32_and_3_22;
  assign f_u_dadda_cla32_fa199_or0 = f_u_dadda_cla32_fa199_and0 | f_u_dadda_cla32_fa199_and1;
  assign f_u_dadda_cla32_and_2_23 = a[2] & b[23];
  assign f_u_dadda_cla32_and_1_24 = a[1] & b[24];
  assign f_u_dadda_cla32_and_0_25 = a[0] & b[25];
  assign f_u_dadda_cla32_fa200_xor0 = f_u_dadda_cla32_and_2_23 ^ f_u_dadda_cla32_and_1_24;
  assign f_u_dadda_cla32_fa200_and0 = f_u_dadda_cla32_and_2_23 & f_u_dadda_cla32_and_1_24;
  assign f_u_dadda_cla32_fa200_xor1 = f_u_dadda_cla32_fa200_xor0 ^ f_u_dadda_cla32_and_0_25;
  assign f_u_dadda_cla32_fa200_and1 = f_u_dadda_cla32_fa200_xor0 & f_u_dadda_cla32_and_0_25;
  assign f_u_dadda_cla32_fa200_or0 = f_u_dadda_cla32_fa200_and0 | f_u_dadda_cla32_fa200_and1;
  assign f_u_dadda_cla32_fa201_xor0 = f_u_dadda_cla32_fa186_xor1 ^ f_u_dadda_cla32_fa187_xor1;
  assign f_u_dadda_cla32_fa201_and0 = f_u_dadda_cla32_fa186_xor1 & f_u_dadda_cla32_fa187_xor1;
  assign f_u_dadda_cla32_fa201_xor1 = f_u_dadda_cla32_fa201_xor0 ^ f_u_dadda_cla32_fa188_xor1;
  assign f_u_dadda_cla32_fa201_and1 = f_u_dadda_cla32_fa201_xor0 & f_u_dadda_cla32_fa188_xor1;
  assign f_u_dadda_cla32_fa201_or0 = f_u_dadda_cla32_fa201_and0 | f_u_dadda_cla32_fa201_and1;
  assign f_u_dadda_cla32_fa202_xor0 = f_u_dadda_cla32_fa189_xor1 ^ f_u_dadda_cla32_fa190_xor1;
  assign f_u_dadda_cla32_fa202_and0 = f_u_dadda_cla32_fa189_xor1 & f_u_dadda_cla32_fa190_xor1;
  assign f_u_dadda_cla32_fa202_xor1 = f_u_dadda_cla32_fa202_xor0 ^ f_u_dadda_cla32_fa191_xor1;
  assign f_u_dadda_cla32_fa202_and1 = f_u_dadda_cla32_fa202_xor0 & f_u_dadda_cla32_fa191_xor1;
  assign f_u_dadda_cla32_fa202_or0 = f_u_dadda_cla32_fa202_and0 | f_u_dadda_cla32_fa202_and1;
  assign f_u_dadda_cla32_fa203_xor0 = f_u_dadda_cla32_fa192_xor1 ^ f_u_dadda_cla32_fa193_xor1;
  assign f_u_dadda_cla32_fa203_and0 = f_u_dadda_cla32_fa192_xor1 & f_u_dadda_cla32_fa193_xor1;
  assign f_u_dadda_cla32_fa203_xor1 = f_u_dadda_cla32_fa203_xor0 ^ f_u_dadda_cla32_fa194_xor1;
  assign f_u_dadda_cla32_fa203_and1 = f_u_dadda_cla32_fa203_xor0 & f_u_dadda_cla32_fa194_xor1;
  assign f_u_dadda_cla32_fa203_or0 = f_u_dadda_cla32_fa203_and0 | f_u_dadda_cla32_fa203_and1;
  assign f_u_dadda_cla32_fa204_xor0 = f_u_dadda_cla32_fa195_xor1 ^ f_u_dadda_cla32_fa196_xor1;
  assign f_u_dadda_cla32_fa204_and0 = f_u_dadda_cla32_fa195_xor1 & f_u_dadda_cla32_fa196_xor1;
  assign f_u_dadda_cla32_fa204_xor1 = f_u_dadda_cla32_fa204_xor0 ^ f_u_dadda_cla32_fa197_xor1;
  assign f_u_dadda_cla32_fa204_and1 = f_u_dadda_cla32_fa204_xor0 & f_u_dadda_cla32_fa197_xor1;
  assign f_u_dadda_cla32_fa204_or0 = f_u_dadda_cla32_fa204_and0 | f_u_dadda_cla32_fa204_and1;
  assign f_u_dadda_cla32_ha24_xor0 = f_u_dadda_cla32_fa198_xor1 ^ f_u_dadda_cla32_fa199_xor1;
  assign f_u_dadda_cla32_ha24_and0 = f_u_dadda_cla32_fa198_xor1 & f_u_dadda_cla32_fa199_xor1;
  assign f_u_dadda_cla32_fa205_xor0 = f_u_dadda_cla32_ha24_and0 ^ f_u_dadda_cla32_fa204_or0;
  assign f_u_dadda_cla32_fa205_and0 = f_u_dadda_cla32_ha24_and0 & f_u_dadda_cla32_fa204_or0;
  assign f_u_dadda_cla32_fa205_xor1 = f_u_dadda_cla32_fa205_xor0 ^ f_u_dadda_cla32_fa203_or0;
  assign f_u_dadda_cla32_fa205_and1 = f_u_dadda_cla32_fa205_xor0 & f_u_dadda_cla32_fa203_or0;
  assign f_u_dadda_cla32_fa205_or0 = f_u_dadda_cla32_fa205_and0 | f_u_dadda_cla32_fa205_and1;
  assign f_u_dadda_cla32_fa206_xor0 = f_u_dadda_cla32_fa202_or0 ^ f_u_dadda_cla32_fa201_or0;
  assign f_u_dadda_cla32_fa206_and0 = f_u_dadda_cla32_fa202_or0 & f_u_dadda_cla32_fa201_or0;
  assign f_u_dadda_cla32_fa206_xor1 = f_u_dadda_cla32_fa206_xor0 ^ f_u_dadda_cla32_fa200_or0;
  assign f_u_dadda_cla32_fa206_and1 = f_u_dadda_cla32_fa206_xor0 & f_u_dadda_cla32_fa200_or0;
  assign f_u_dadda_cla32_fa206_or0 = f_u_dadda_cla32_fa206_and0 | f_u_dadda_cla32_fa206_and1;
  assign f_u_dadda_cla32_fa207_xor0 = f_u_dadda_cla32_fa199_or0 ^ f_u_dadda_cla32_fa198_or0;
  assign f_u_dadda_cla32_fa207_and0 = f_u_dadda_cla32_fa199_or0 & f_u_dadda_cla32_fa198_or0;
  assign f_u_dadda_cla32_fa207_xor1 = f_u_dadda_cla32_fa207_xor0 ^ f_u_dadda_cla32_fa197_or0;
  assign f_u_dadda_cla32_fa207_and1 = f_u_dadda_cla32_fa207_xor0 & f_u_dadda_cla32_fa197_or0;
  assign f_u_dadda_cla32_fa207_or0 = f_u_dadda_cla32_fa207_and0 | f_u_dadda_cla32_fa207_and1;
  assign f_u_dadda_cla32_fa208_xor0 = f_u_dadda_cla32_fa196_or0 ^ f_u_dadda_cla32_fa195_or0;
  assign f_u_dadda_cla32_fa208_and0 = f_u_dadda_cla32_fa196_or0 & f_u_dadda_cla32_fa195_or0;
  assign f_u_dadda_cla32_fa208_xor1 = f_u_dadda_cla32_fa208_xor0 ^ f_u_dadda_cla32_fa194_or0;
  assign f_u_dadda_cla32_fa208_and1 = f_u_dadda_cla32_fa208_xor0 & f_u_dadda_cla32_fa194_or0;
  assign f_u_dadda_cla32_fa208_or0 = f_u_dadda_cla32_fa208_and0 | f_u_dadda_cla32_fa208_and1;
  assign f_u_dadda_cla32_fa209_xor0 = f_u_dadda_cla32_fa193_or0 ^ f_u_dadda_cla32_fa192_or0;
  assign f_u_dadda_cla32_fa209_and0 = f_u_dadda_cla32_fa193_or0 & f_u_dadda_cla32_fa192_or0;
  assign f_u_dadda_cla32_fa209_xor1 = f_u_dadda_cla32_fa209_xor0 ^ f_u_dadda_cla32_fa191_or0;
  assign f_u_dadda_cla32_fa209_and1 = f_u_dadda_cla32_fa209_xor0 & f_u_dadda_cla32_fa191_or0;
  assign f_u_dadda_cla32_fa209_or0 = f_u_dadda_cla32_fa209_and0 | f_u_dadda_cla32_fa209_and1;
  assign f_u_dadda_cla32_fa210_xor0 = f_u_dadda_cla32_fa190_or0 ^ f_u_dadda_cla32_fa189_or0;
  assign f_u_dadda_cla32_fa210_and0 = f_u_dadda_cla32_fa190_or0 & f_u_dadda_cla32_fa189_or0;
  assign f_u_dadda_cla32_fa210_xor1 = f_u_dadda_cla32_fa210_xor0 ^ f_u_dadda_cla32_fa188_or0;
  assign f_u_dadda_cla32_fa210_and1 = f_u_dadda_cla32_fa210_xor0 & f_u_dadda_cla32_fa188_or0;
  assign f_u_dadda_cla32_fa210_or0 = f_u_dadda_cla32_fa210_and0 | f_u_dadda_cla32_fa210_and1;
  assign f_u_dadda_cla32_and_26_0 = a[26] & b[0];
  assign f_u_dadda_cla32_fa211_xor0 = f_u_dadda_cla32_fa187_or0 ^ f_u_dadda_cla32_fa186_or0;
  assign f_u_dadda_cla32_fa211_and0 = f_u_dadda_cla32_fa187_or0 & f_u_dadda_cla32_fa186_or0;
  assign f_u_dadda_cla32_fa211_xor1 = f_u_dadda_cla32_fa211_xor0 ^ f_u_dadda_cla32_and_26_0;
  assign f_u_dadda_cla32_fa211_and1 = f_u_dadda_cla32_fa211_xor0 & f_u_dadda_cla32_and_26_0;
  assign f_u_dadda_cla32_fa211_or0 = f_u_dadda_cla32_fa211_and0 | f_u_dadda_cla32_fa211_and1;
  assign f_u_dadda_cla32_and_25_1 = a[25] & b[1];
  assign f_u_dadda_cla32_and_24_2 = a[24] & b[2];
  assign f_u_dadda_cla32_and_23_3 = a[23] & b[3];
  assign f_u_dadda_cla32_fa212_xor0 = f_u_dadda_cla32_and_25_1 ^ f_u_dadda_cla32_and_24_2;
  assign f_u_dadda_cla32_fa212_and0 = f_u_dadda_cla32_and_25_1 & f_u_dadda_cla32_and_24_2;
  assign f_u_dadda_cla32_fa212_xor1 = f_u_dadda_cla32_fa212_xor0 ^ f_u_dadda_cla32_and_23_3;
  assign f_u_dadda_cla32_fa212_and1 = f_u_dadda_cla32_fa212_xor0 & f_u_dadda_cla32_and_23_3;
  assign f_u_dadda_cla32_fa212_or0 = f_u_dadda_cla32_fa212_and0 | f_u_dadda_cla32_fa212_and1;
  assign f_u_dadda_cla32_and_22_4 = a[22] & b[4];
  assign f_u_dadda_cla32_and_21_5 = a[21] & b[5];
  assign f_u_dadda_cla32_and_20_6 = a[20] & b[6];
  assign f_u_dadda_cla32_fa213_xor0 = f_u_dadda_cla32_and_22_4 ^ f_u_dadda_cla32_and_21_5;
  assign f_u_dadda_cla32_fa213_and0 = f_u_dadda_cla32_and_22_4 & f_u_dadda_cla32_and_21_5;
  assign f_u_dadda_cla32_fa213_xor1 = f_u_dadda_cla32_fa213_xor0 ^ f_u_dadda_cla32_and_20_6;
  assign f_u_dadda_cla32_fa213_and1 = f_u_dadda_cla32_fa213_xor0 & f_u_dadda_cla32_and_20_6;
  assign f_u_dadda_cla32_fa213_or0 = f_u_dadda_cla32_fa213_and0 | f_u_dadda_cla32_fa213_and1;
  assign f_u_dadda_cla32_and_19_7 = a[19] & b[7];
  assign f_u_dadda_cla32_and_18_8 = a[18] & b[8];
  assign f_u_dadda_cla32_and_17_9 = a[17] & b[9];
  assign f_u_dadda_cla32_fa214_xor0 = f_u_dadda_cla32_and_19_7 ^ f_u_dadda_cla32_and_18_8;
  assign f_u_dadda_cla32_fa214_and0 = f_u_dadda_cla32_and_19_7 & f_u_dadda_cla32_and_18_8;
  assign f_u_dadda_cla32_fa214_xor1 = f_u_dadda_cla32_fa214_xor0 ^ f_u_dadda_cla32_and_17_9;
  assign f_u_dadda_cla32_fa214_and1 = f_u_dadda_cla32_fa214_xor0 & f_u_dadda_cla32_and_17_9;
  assign f_u_dadda_cla32_fa214_or0 = f_u_dadda_cla32_fa214_and0 | f_u_dadda_cla32_fa214_and1;
  assign f_u_dadda_cla32_and_16_10 = a[16] & b[10];
  assign f_u_dadda_cla32_and_15_11 = a[15] & b[11];
  assign f_u_dadda_cla32_and_14_12 = a[14] & b[12];
  assign f_u_dadda_cla32_fa215_xor0 = f_u_dadda_cla32_and_16_10 ^ f_u_dadda_cla32_and_15_11;
  assign f_u_dadda_cla32_fa215_and0 = f_u_dadda_cla32_and_16_10 & f_u_dadda_cla32_and_15_11;
  assign f_u_dadda_cla32_fa215_xor1 = f_u_dadda_cla32_fa215_xor0 ^ f_u_dadda_cla32_and_14_12;
  assign f_u_dadda_cla32_fa215_and1 = f_u_dadda_cla32_fa215_xor0 & f_u_dadda_cla32_and_14_12;
  assign f_u_dadda_cla32_fa215_or0 = f_u_dadda_cla32_fa215_and0 | f_u_dadda_cla32_fa215_and1;
  assign f_u_dadda_cla32_and_13_13 = a[13] & b[13];
  assign f_u_dadda_cla32_and_12_14 = a[12] & b[14];
  assign f_u_dadda_cla32_and_11_15 = a[11] & b[15];
  assign f_u_dadda_cla32_fa216_xor0 = f_u_dadda_cla32_and_13_13 ^ f_u_dadda_cla32_and_12_14;
  assign f_u_dadda_cla32_fa216_and0 = f_u_dadda_cla32_and_13_13 & f_u_dadda_cla32_and_12_14;
  assign f_u_dadda_cla32_fa216_xor1 = f_u_dadda_cla32_fa216_xor0 ^ f_u_dadda_cla32_and_11_15;
  assign f_u_dadda_cla32_fa216_and1 = f_u_dadda_cla32_fa216_xor0 & f_u_dadda_cla32_and_11_15;
  assign f_u_dadda_cla32_fa216_or0 = f_u_dadda_cla32_fa216_and0 | f_u_dadda_cla32_fa216_and1;
  assign f_u_dadda_cla32_and_10_16 = a[10] & b[16];
  assign f_u_dadda_cla32_and_9_17 = a[9] & b[17];
  assign f_u_dadda_cla32_and_8_18 = a[8] & b[18];
  assign f_u_dadda_cla32_fa217_xor0 = f_u_dadda_cla32_and_10_16 ^ f_u_dadda_cla32_and_9_17;
  assign f_u_dadda_cla32_fa217_and0 = f_u_dadda_cla32_and_10_16 & f_u_dadda_cla32_and_9_17;
  assign f_u_dadda_cla32_fa217_xor1 = f_u_dadda_cla32_fa217_xor0 ^ f_u_dadda_cla32_and_8_18;
  assign f_u_dadda_cla32_fa217_and1 = f_u_dadda_cla32_fa217_xor0 & f_u_dadda_cla32_and_8_18;
  assign f_u_dadda_cla32_fa217_or0 = f_u_dadda_cla32_fa217_and0 | f_u_dadda_cla32_fa217_and1;
  assign f_u_dadda_cla32_and_7_19 = a[7] & b[19];
  assign f_u_dadda_cla32_and_6_20 = a[6] & b[20];
  assign f_u_dadda_cla32_and_5_21 = a[5] & b[21];
  assign f_u_dadda_cla32_fa218_xor0 = f_u_dadda_cla32_and_7_19 ^ f_u_dadda_cla32_and_6_20;
  assign f_u_dadda_cla32_fa218_and0 = f_u_dadda_cla32_and_7_19 & f_u_dadda_cla32_and_6_20;
  assign f_u_dadda_cla32_fa218_xor1 = f_u_dadda_cla32_fa218_xor0 ^ f_u_dadda_cla32_and_5_21;
  assign f_u_dadda_cla32_fa218_and1 = f_u_dadda_cla32_fa218_xor0 & f_u_dadda_cla32_and_5_21;
  assign f_u_dadda_cla32_fa218_or0 = f_u_dadda_cla32_fa218_and0 | f_u_dadda_cla32_fa218_and1;
  assign f_u_dadda_cla32_and_4_22 = a[4] & b[22];
  assign f_u_dadda_cla32_and_3_23 = a[3] & b[23];
  assign f_u_dadda_cla32_and_2_24 = a[2] & b[24];
  assign f_u_dadda_cla32_fa219_xor0 = f_u_dadda_cla32_and_4_22 ^ f_u_dadda_cla32_and_3_23;
  assign f_u_dadda_cla32_fa219_and0 = f_u_dadda_cla32_and_4_22 & f_u_dadda_cla32_and_3_23;
  assign f_u_dadda_cla32_fa219_xor1 = f_u_dadda_cla32_fa219_xor0 ^ f_u_dadda_cla32_and_2_24;
  assign f_u_dadda_cla32_fa219_and1 = f_u_dadda_cla32_fa219_xor0 & f_u_dadda_cla32_and_2_24;
  assign f_u_dadda_cla32_fa219_or0 = f_u_dadda_cla32_fa219_and0 | f_u_dadda_cla32_fa219_and1;
  assign f_u_dadda_cla32_and_1_25 = a[1] & b[25];
  assign f_u_dadda_cla32_and_0_26 = a[0] & b[26];
  assign f_u_dadda_cla32_fa220_xor0 = f_u_dadda_cla32_and_1_25 ^ f_u_dadda_cla32_and_0_26;
  assign f_u_dadda_cla32_fa220_and0 = f_u_dadda_cla32_and_1_25 & f_u_dadda_cla32_and_0_26;
  assign f_u_dadda_cla32_fa220_xor1 = f_u_dadda_cla32_fa220_xor0 ^ f_u_dadda_cla32_fa205_xor1;
  assign f_u_dadda_cla32_fa220_and1 = f_u_dadda_cla32_fa220_xor0 & f_u_dadda_cla32_fa205_xor1;
  assign f_u_dadda_cla32_fa220_or0 = f_u_dadda_cla32_fa220_and0 | f_u_dadda_cla32_fa220_and1;
  assign f_u_dadda_cla32_fa221_xor0 = f_u_dadda_cla32_fa206_xor1 ^ f_u_dadda_cla32_fa207_xor1;
  assign f_u_dadda_cla32_fa221_and0 = f_u_dadda_cla32_fa206_xor1 & f_u_dadda_cla32_fa207_xor1;
  assign f_u_dadda_cla32_fa221_xor1 = f_u_dadda_cla32_fa221_xor0 ^ f_u_dadda_cla32_fa208_xor1;
  assign f_u_dadda_cla32_fa221_and1 = f_u_dadda_cla32_fa221_xor0 & f_u_dadda_cla32_fa208_xor1;
  assign f_u_dadda_cla32_fa221_or0 = f_u_dadda_cla32_fa221_and0 | f_u_dadda_cla32_fa221_and1;
  assign f_u_dadda_cla32_fa222_xor0 = f_u_dadda_cla32_fa209_xor1 ^ f_u_dadda_cla32_fa210_xor1;
  assign f_u_dadda_cla32_fa222_and0 = f_u_dadda_cla32_fa209_xor1 & f_u_dadda_cla32_fa210_xor1;
  assign f_u_dadda_cla32_fa222_xor1 = f_u_dadda_cla32_fa222_xor0 ^ f_u_dadda_cla32_fa211_xor1;
  assign f_u_dadda_cla32_fa222_and1 = f_u_dadda_cla32_fa222_xor0 & f_u_dadda_cla32_fa211_xor1;
  assign f_u_dadda_cla32_fa222_or0 = f_u_dadda_cla32_fa222_and0 | f_u_dadda_cla32_fa222_and1;
  assign f_u_dadda_cla32_fa223_xor0 = f_u_dadda_cla32_fa212_xor1 ^ f_u_dadda_cla32_fa213_xor1;
  assign f_u_dadda_cla32_fa223_and0 = f_u_dadda_cla32_fa212_xor1 & f_u_dadda_cla32_fa213_xor1;
  assign f_u_dadda_cla32_fa223_xor1 = f_u_dadda_cla32_fa223_xor0 ^ f_u_dadda_cla32_fa214_xor1;
  assign f_u_dadda_cla32_fa223_and1 = f_u_dadda_cla32_fa223_xor0 & f_u_dadda_cla32_fa214_xor1;
  assign f_u_dadda_cla32_fa223_or0 = f_u_dadda_cla32_fa223_and0 | f_u_dadda_cla32_fa223_and1;
  assign f_u_dadda_cla32_fa224_xor0 = f_u_dadda_cla32_fa215_xor1 ^ f_u_dadda_cla32_fa216_xor1;
  assign f_u_dadda_cla32_fa224_and0 = f_u_dadda_cla32_fa215_xor1 & f_u_dadda_cla32_fa216_xor1;
  assign f_u_dadda_cla32_fa224_xor1 = f_u_dadda_cla32_fa224_xor0 ^ f_u_dadda_cla32_fa217_xor1;
  assign f_u_dadda_cla32_fa224_and1 = f_u_dadda_cla32_fa224_xor0 & f_u_dadda_cla32_fa217_xor1;
  assign f_u_dadda_cla32_fa224_or0 = f_u_dadda_cla32_fa224_and0 | f_u_dadda_cla32_fa224_and1;
  assign f_u_dadda_cla32_ha25_xor0 = f_u_dadda_cla32_fa218_xor1 ^ f_u_dadda_cla32_fa219_xor1;
  assign f_u_dadda_cla32_ha25_and0 = f_u_dadda_cla32_fa218_xor1 & f_u_dadda_cla32_fa219_xor1;
  assign f_u_dadda_cla32_fa225_xor0 = f_u_dadda_cla32_ha25_and0 ^ f_u_dadda_cla32_fa224_or0;
  assign f_u_dadda_cla32_fa225_and0 = f_u_dadda_cla32_ha25_and0 & f_u_dadda_cla32_fa224_or0;
  assign f_u_dadda_cla32_fa225_xor1 = f_u_dadda_cla32_fa225_xor0 ^ f_u_dadda_cla32_fa223_or0;
  assign f_u_dadda_cla32_fa225_and1 = f_u_dadda_cla32_fa225_xor0 & f_u_dadda_cla32_fa223_or0;
  assign f_u_dadda_cla32_fa225_or0 = f_u_dadda_cla32_fa225_and0 | f_u_dadda_cla32_fa225_and1;
  assign f_u_dadda_cla32_fa226_xor0 = f_u_dadda_cla32_fa222_or0 ^ f_u_dadda_cla32_fa221_or0;
  assign f_u_dadda_cla32_fa226_and0 = f_u_dadda_cla32_fa222_or0 & f_u_dadda_cla32_fa221_or0;
  assign f_u_dadda_cla32_fa226_xor1 = f_u_dadda_cla32_fa226_xor0 ^ f_u_dadda_cla32_fa220_or0;
  assign f_u_dadda_cla32_fa226_and1 = f_u_dadda_cla32_fa226_xor0 & f_u_dadda_cla32_fa220_or0;
  assign f_u_dadda_cla32_fa226_or0 = f_u_dadda_cla32_fa226_and0 | f_u_dadda_cla32_fa226_and1;
  assign f_u_dadda_cla32_fa227_xor0 = f_u_dadda_cla32_fa219_or0 ^ f_u_dadda_cla32_fa218_or0;
  assign f_u_dadda_cla32_fa227_and0 = f_u_dadda_cla32_fa219_or0 & f_u_dadda_cla32_fa218_or0;
  assign f_u_dadda_cla32_fa227_xor1 = f_u_dadda_cla32_fa227_xor0 ^ f_u_dadda_cla32_fa217_or0;
  assign f_u_dadda_cla32_fa227_and1 = f_u_dadda_cla32_fa227_xor0 & f_u_dadda_cla32_fa217_or0;
  assign f_u_dadda_cla32_fa227_or0 = f_u_dadda_cla32_fa227_and0 | f_u_dadda_cla32_fa227_and1;
  assign f_u_dadda_cla32_fa228_xor0 = f_u_dadda_cla32_fa216_or0 ^ f_u_dadda_cla32_fa215_or0;
  assign f_u_dadda_cla32_fa228_and0 = f_u_dadda_cla32_fa216_or0 & f_u_dadda_cla32_fa215_or0;
  assign f_u_dadda_cla32_fa228_xor1 = f_u_dadda_cla32_fa228_xor0 ^ f_u_dadda_cla32_fa214_or0;
  assign f_u_dadda_cla32_fa228_and1 = f_u_dadda_cla32_fa228_xor0 & f_u_dadda_cla32_fa214_or0;
  assign f_u_dadda_cla32_fa228_or0 = f_u_dadda_cla32_fa228_and0 | f_u_dadda_cla32_fa228_and1;
  assign f_u_dadda_cla32_fa229_xor0 = f_u_dadda_cla32_fa213_or0 ^ f_u_dadda_cla32_fa212_or0;
  assign f_u_dadda_cla32_fa229_and0 = f_u_dadda_cla32_fa213_or0 & f_u_dadda_cla32_fa212_or0;
  assign f_u_dadda_cla32_fa229_xor1 = f_u_dadda_cla32_fa229_xor0 ^ f_u_dadda_cla32_fa211_or0;
  assign f_u_dadda_cla32_fa229_and1 = f_u_dadda_cla32_fa229_xor0 & f_u_dadda_cla32_fa211_or0;
  assign f_u_dadda_cla32_fa229_or0 = f_u_dadda_cla32_fa229_and0 | f_u_dadda_cla32_fa229_and1;
  assign f_u_dadda_cla32_fa230_xor0 = f_u_dadda_cla32_fa210_or0 ^ f_u_dadda_cla32_fa209_or0;
  assign f_u_dadda_cla32_fa230_and0 = f_u_dadda_cla32_fa210_or0 & f_u_dadda_cla32_fa209_or0;
  assign f_u_dadda_cla32_fa230_xor1 = f_u_dadda_cla32_fa230_xor0 ^ f_u_dadda_cla32_fa208_or0;
  assign f_u_dadda_cla32_fa230_and1 = f_u_dadda_cla32_fa230_xor0 & f_u_dadda_cla32_fa208_or0;
  assign f_u_dadda_cla32_fa230_or0 = f_u_dadda_cla32_fa230_and0 | f_u_dadda_cla32_fa230_and1;
  assign f_u_dadda_cla32_fa231_xor0 = f_u_dadda_cla32_fa207_or0 ^ f_u_dadda_cla32_fa206_or0;
  assign f_u_dadda_cla32_fa231_and0 = f_u_dadda_cla32_fa207_or0 & f_u_dadda_cla32_fa206_or0;
  assign f_u_dadda_cla32_fa231_xor1 = f_u_dadda_cla32_fa231_xor0 ^ f_u_dadda_cla32_fa205_or0;
  assign f_u_dadda_cla32_fa231_and1 = f_u_dadda_cla32_fa231_xor0 & f_u_dadda_cla32_fa205_or0;
  assign f_u_dadda_cla32_fa231_or0 = f_u_dadda_cla32_fa231_and0 | f_u_dadda_cla32_fa231_and1;
  assign f_u_dadda_cla32_and_27_0 = a[27] & b[0];
  assign f_u_dadda_cla32_and_26_1 = a[26] & b[1];
  assign f_u_dadda_cla32_and_25_2 = a[25] & b[2];
  assign f_u_dadda_cla32_fa232_xor0 = f_u_dadda_cla32_and_27_0 ^ f_u_dadda_cla32_and_26_1;
  assign f_u_dadda_cla32_fa232_and0 = f_u_dadda_cla32_and_27_0 & f_u_dadda_cla32_and_26_1;
  assign f_u_dadda_cla32_fa232_xor1 = f_u_dadda_cla32_fa232_xor0 ^ f_u_dadda_cla32_and_25_2;
  assign f_u_dadda_cla32_fa232_and1 = f_u_dadda_cla32_fa232_xor0 & f_u_dadda_cla32_and_25_2;
  assign f_u_dadda_cla32_fa232_or0 = f_u_dadda_cla32_fa232_and0 | f_u_dadda_cla32_fa232_and1;
  assign f_u_dadda_cla32_and_24_3 = a[24] & b[3];
  assign f_u_dadda_cla32_and_23_4 = a[23] & b[4];
  assign f_u_dadda_cla32_and_22_5 = a[22] & b[5];
  assign f_u_dadda_cla32_fa233_xor0 = f_u_dadda_cla32_and_24_3 ^ f_u_dadda_cla32_and_23_4;
  assign f_u_dadda_cla32_fa233_and0 = f_u_dadda_cla32_and_24_3 & f_u_dadda_cla32_and_23_4;
  assign f_u_dadda_cla32_fa233_xor1 = f_u_dadda_cla32_fa233_xor0 ^ f_u_dadda_cla32_and_22_5;
  assign f_u_dadda_cla32_fa233_and1 = f_u_dadda_cla32_fa233_xor0 & f_u_dadda_cla32_and_22_5;
  assign f_u_dadda_cla32_fa233_or0 = f_u_dadda_cla32_fa233_and0 | f_u_dadda_cla32_fa233_and1;
  assign f_u_dadda_cla32_and_21_6 = a[21] & b[6];
  assign f_u_dadda_cla32_and_20_7 = a[20] & b[7];
  assign f_u_dadda_cla32_and_19_8 = a[19] & b[8];
  assign f_u_dadda_cla32_fa234_xor0 = f_u_dadda_cla32_and_21_6 ^ f_u_dadda_cla32_and_20_7;
  assign f_u_dadda_cla32_fa234_and0 = f_u_dadda_cla32_and_21_6 & f_u_dadda_cla32_and_20_7;
  assign f_u_dadda_cla32_fa234_xor1 = f_u_dadda_cla32_fa234_xor0 ^ f_u_dadda_cla32_and_19_8;
  assign f_u_dadda_cla32_fa234_and1 = f_u_dadda_cla32_fa234_xor0 & f_u_dadda_cla32_and_19_8;
  assign f_u_dadda_cla32_fa234_or0 = f_u_dadda_cla32_fa234_and0 | f_u_dadda_cla32_fa234_and1;
  assign f_u_dadda_cla32_and_18_9 = a[18] & b[9];
  assign f_u_dadda_cla32_and_17_10 = a[17] & b[10];
  assign f_u_dadda_cla32_and_16_11 = a[16] & b[11];
  assign f_u_dadda_cla32_fa235_xor0 = f_u_dadda_cla32_and_18_9 ^ f_u_dadda_cla32_and_17_10;
  assign f_u_dadda_cla32_fa235_and0 = f_u_dadda_cla32_and_18_9 & f_u_dadda_cla32_and_17_10;
  assign f_u_dadda_cla32_fa235_xor1 = f_u_dadda_cla32_fa235_xor0 ^ f_u_dadda_cla32_and_16_11;
  assign f_u_dadda_cla32_fa235_and1 = f_u_dadda_cla32_fa235_xor0 & f_u_dadda_cla32_and_16_11;
  assign f_u_dadda_cla32_fa235_or0 = f_u_dadda_cla32_fa235_and0 | f_u_dadda_cla32_fa235_and1;
  assign f_u_dadda_cla32_and_15_12 = a[15] & b[12];
  assign f_u_dadda_cla32_and_14_13 = a[14] & b[13];
  assign f_u_dadda_cla32_and_13_14 = a[13] & b[14];
  assign f_u_dadda_cla32_fa236_xor0 = f_u_dadda_cla32_and_15_12 ^ f_u_dadda_cla32_and_14_13;
  assign f_u_dadda_cla32_fa236_and0 = f_u_dadda_cla32_and_15_12 & f_u_dadda_cla32_and_14_13;
  assign f_u_dadda_cla32_fa236_xor1 = f_u_dadda_cla32_fa236_xor0 ^ f_u_dadda_cla32_and_13_14;
  assign f_u_dadda_cla32_fa236_and1 = f_u_dadda_cla32_fa236_xor0 & f_u_dadda_cla32_and_13_14;
  assign f_u_dadda_cla32_fa236_or0 = f_u_dadda_cla32_fa236_and0 | f_u_dadda_cla32_fa236_and1;
  assign f_u_dadda_cla32_and_12_15 = a[12] & b[15];
  assign f_u_dadda_cla32_and_11_16 = a[11] & b[16];
  assign f_u_dadda_cla32_and_10_17 = a[10] & b[17];
  assign f_u_dadda_cla32_fa237_xor0 = f_u_dadda_cla32_and_12_15 ^ f_u_dadda_cla32_and_11_16;
  assign f_u_dadda_cla32_fa237_and0 = f_u_dadda_cla32_and_12_15 & f_u_dadda_cla32_and_11_16;
  assign f_u_dadda_cla32_fa237_xor1 = f_u_dadda_cla32_fa237_xor0 ^ f_u_dadda_cla32_and_10_17;
  assign f_u_dadda_cla32_fa237_and1 = f_u_dadda_cla32_fa237_xor0 & f_u_dadda_cla32_and_10_17;
  assign f_u_dadda_cla32_fa237_or0 = f_u_dadda_cla32_fa237_and0 | f_u_dadda_cla32_fa237_and1;
  assign f_u_dadda_cla32_and_9_18 = a[9] & b[18];
  assign f_u_dadda_cla32_and_8_19 = a[8] & b[19];
  assign f_u_dadda_cla32_and_7_20 = a[7] & b[20];
  assign f_u_dadda_cla32_fa238_xor0 = f_u_dadda_cla32_and_9_18 ^ f_u_dadda_cla32_and_8_19;
  assign f_u_dadda_cla32_fa238_and0 = f_u_dadda_cla32_and_9_18 & f_u_dadda_cla32_and_8_19;
  assign f_u_dadda_cla32_fa238_xor1 = f_u_dadda_cla32_fa238_xor0 ^ f_u_dadda_cla32_and_7_20;
  assign f_u_dadda_cla32_fa238_and1 = f_u_dadda_cla32_fa238_xor0 & f_u_dadda_cla32_and_7_20;
  assign f_u_dadda_cla32_fa238_or0 = f_u_dadda_cla32_fa238_and0 | f_u_dadda_cla32_fa238_and1;
  assign f_u_dadda_cla32_and_6_21 = a[6] & b[21];
  assign f_u_dadda_cla32_and_5_22 = a[5] & b[22];
  assign f_u_dadda_cla32_and_4_23 = a[4] & b[23];
  assign f_u_dadda_cla32_fa239_xor0 = f_u_dadda_cla32_and_6_21 ^ f_u_dadda_cla32_and_5_22;
  assign f_u_dadda_cla32_fa239_and0 = f_u_dadda_cla32_and_6_21 & f_u_dadda_cla32_and_5_22;
  assign f_u_dadda_cla32_fa239_xor1 = f_u_dadda_cla32_fa239_xor0 ^ f_u_dadda_cla32_and_4_23;
  assign f_u_dadda_cla32_fa239_and1 = f_u_dadda_cla32_fa239_xor0 & f_u_dadda_cla32_and_4_23;
  assign f_u_dadda_cla32_fa239_or0 = f_u_dadda_cla32_fa239_and0 | f_u_dadda_cla32_fa239_and1;
  assign f_u_dadda_cla32_and_3_24 = a[3] & b[24];
  assign f_u_dadda_cla32_and_2_25 = a[2] & b[25];
  assign f_u_dadda_cla32_and_1_26 = a[1] & b[26];
  assign f_u_dadda_cla32_fa240_xor0 = f_u_dadda_cla32_and_3_24 ^ f_u_dadda_cla32_and_2_25;
  assign f_u_dadda_cla32_fa240_and0 = f_u_dadda_cla32_and_3_24 & f_u_dadda_cla32_and_2_25;
  assign f_u_dadda_cla32_fa240_xor1 = f_u_dadda_cla32_fa240_xor0 ^ f_u_dadda_cla32_and_1_26;
  assign f_u_dadda_cla32_fa240_and1 = f_u_dadda_cla32_fa240_xor0 & f_u_dadda_cla32_and_1_26;
  assign f_u_dadda_cla32_fa240_or0 = f_u_dadda_cla32_fa240_and0 | f_u_dadda_cla32_fa240_and1;
  assign f_u_dadda_cla32_and_0_27 = a[0] & b[27];
  assign f_u_dadda_cla32_fa241_xor0 = f_u_dadda_cla32_and_0_27 ^ f_u_dadda_cla32_fa225_xor1;
  assign f_u_dadda_cla32_fa241_and0 = f_u_dadda_cla32_and_0_27 & f_u_dadda_cla32_fa225_xor1;
  assign f_u_dadda_cla32_fa241_xor1 = f_u_dadda_cla32_fa241_xor0 ^ f_u_dadda_cla32_fa226_xor1;
  assign f_u_dadda_cla32_fa241_and1 = f_u_dadda_cla32_fa241_xor0 & f_u_dadda_cla32_fa226_xor1;
  assign f_u_dadda_cla32_fa241_or0 = f_u_dadda_cla32_fa241_and0 | f_u_dadda_cla32_fa241_and1;
  assign f_u_dadda_cla32_fa242_xor0 = f_u_dadda_cla32_fa227_xor1 ^ f_u_dadda_cla32_fa228_xor1;
  assign f_u_dadda_cla32_fa242_and0 = f_u_dadda_cla32_fa227_xor1 & f_u_dadda_cla32_fa228_xor1;
  assign f_u_dadda_cla32_fa242_xor1 = f_u_dadda_cla32_fa242_xor0 ^ f_u_dadda_cla32_fa229_xor1;
  assign f_u_dadda_cla32_fa242_and1 = f_u_dadda_cla32_fa242_xor0 & f_u_dadda_cla32_fa229_xor1;
  assign f_u_dadda_cla32_fa242_or0 = f_u_dadda_cla32_fa242_and0 | f_u_dadda_cla32_fa242_and1;
  assign f_u_dadda_cla32_fa243_xor0 = f_u_dadda_cla32_fa230_xor1 ^ f_u_dadda_cla32_fa231_xor1;
  assign f_u_dadda_cla32_fa243_and0 = f_u_dadda_cla32_fa230_xor1 & f_u_dadda_cla32_fa231_xor1;
  assign f_u_dadda_cla32_fa243_xor1 = f_u_dadda_cla32_fa243_xor0 ^ f_u_dadda_cla32_fa232_xor1;
  assign f_u_dadda_cla32_fa243_and1 = f_u_dadda_cla32_fa243_xor0 & f_u_dadda_cla32_fa232_xor1;
  assign f_u_dadda_cla32_fa243_or0 = f_u_dadda_cla32_fa243_and0 | f_u_dadda_cla32_fa243_and1;
  assign f_u_dadda_cla32_fa244_xor0 = f_u_dadda_cla32_fa233_xor1 ^ f_u_dadda_cla32_fa234_xor1;
  assign f_u_dadda_cla32_fa244_and0 = f_u_dadda_cla32_fa233_xor1 & f_u_dadda_cla32_fa234_xor1;
  assign f_u_dadda_cla32_fa244_xor1 = f_u_dadda_cla32_fa244_xor0 ^ f_u_dadda_cla32_fa235_xor1;
  assign f_u_dadda_cla32_fa244_and1 = f_u_dadda_cla32_fa244_xor0 & f_u_dadda_cla32_fa235_xor1;
  assign f_u_dadda_cla32_fa244_or0 = f_u_dadda_cla32_fa244_and0 | f_u_dadda_cla32_fa244_and1;
  assign f_u_dadda_cla32_fa245_xor0 = f_u_dadda_cla32_fa236_xor1 ^ f_u_dadda_cla32_fa237_xor1;
  assign f_u_dadda_cla32_fa245_and0 = f_u_dadda_cla32_fa236_xor1 & f_u_dadda_cla32_fa237_xor1;
  assign f_u_dadda_cla32_fa245_xor1 = f_u_dadda_cla32_fa245_xor0 ^ f_u_dadda_cla32_fa238_xor1;
  assign f_u_dadda_cla32_fa245_and1 = f_u_dadda_cla32_fa245_xor0 & f_u_dadda_cla32_fa238_xor1;
  assign f_u_dadda_cla32_fa245_or0 = f_u_dadda_cla32_fa245_and0 | f_u_dadda_cla32_fa245_and1;
  assign f_u_dadda_cla32_ha26_xor0 = f_u_dadda_cla32_fa239_xor1 ^ f_u_dadda_cla32_fa240_xor1;
  assign f_u_dadda_cla32_ha26_and0 = f_u_dadda_cla32_fa239_xor1 & f_u_dadda_cla32_fa240_xor1;
  assign f_u_dadda_cla32_fa246_xor0 = f_u_dadda_cla32_ha26_and0 ^ f_u_dadda_cla32_fa245_or0;
  assign f_u_dadda_cla32_fa246_and0 = f_u_dadda_cla32_ha26_and0 & f_u_dadda_cla32_fa245_or0;
  assign f_u_dadda_cla32_fa246_xor1 = f_u_dadda_cla32_fa246_xor0 ^ f_u_dadda_cla32_fa244_or0;
  assign f_u_dadda_cla32_fa246_and1 = f_u_dadda_cla32_fa246_xor0 & f_u_dadda_cla32_fa244_or0;
  assign f_u_dadda_cla32_fa246_or0 = f_u_dadda_cla32_fa246_and0 | f_u_dadda_cla32_fa246_and1;
  assign f_u_dadda_cla32_fa247_xor0 = f_u_dadda_cla32_fa243_or0 ^ f_u_dadda_cla32_fa242_or0;
  assign f_u_dadda_cla32_fa247_and0 = f_u_dadda_cla32_fa243_or0 & f_u_dadda_cla32_fa242_or0;
  assign f_u_dadda_cla32_fa247_xor1 = f_u_dadda_cla32_fa247_xor0 ^ f_u_dadda_cla32_fa241_or0;
  assign f_u_dadda_cla32_fa247_and1 = f_u_dadda_cla32_fa247_xor0 & f_u_dadda_cla32_fa241_or0;
  assign f_u_dadda_cla32_fa247_or0 = f_u_dadda_cla32_fa247_and0 | f_u_dadda_cla32_fa247_and1;
  assign f_u_dadda_cla32_fa248_xor0 = f_u_dadda_cla32_fa240_or0 ^ f_u_dadda_cla32_fa239_or0;
  assign f_u_dadda_cla32_fa248_and0 = f_u_dadda_cla32_fa240_or0 & f_u_dadda_cla32_fa239_or0;
  assign f_u_dadda_cla32_fa248_xor1 = f_u_dadda_cla32_fa248_xor0 ^ f_u_dadda_cla32_fa238_or0;
  assign f_u_dadda_cla32_fa248_and1 = f_u_dadda_cla32_fa248_xor0 & f_u_dadda_cla32_fa238_or0;
  assign f_u_dadda_cla32_fa248_or0 = f_u_dadda_cla32_fa248_and0 | f_u_dadda_cla32_fa248_and1;
  assign f_u_dadda_cla32_fa249_xor0 = f_u_dadda_cla32_fa237_or0 ^ f_u_dadda_cla32_fa236_or0;
  assign f_u_dadda_cla32_fa249_and0 = f_u_dadda_cla32_fa237_or0 & f_u_dadda_cla32_fa236_or0;
  assign f_u_dadda_cla32_fa249_xor1 = f_u_dadda_cla32_fa249_xor0 ^ f_u_dadda_cla32_fa235_or0;
  assign f_u_dadda_cla32_fa249_and1 = f_u_dadda_cla32_fa249_xor0 & f_u_dadda_cla32_fa235_or0;
  assign f_u_dadda_cla32_fa249_or0 = f_u_dadda_cla32_fa249_and0 | f_u_dadda_cla32_fa249_and1;
  assign f_u_dadda_cla32_fa250_xor0 = f_u_dadda_cla32_fa234_or0 ^ f_u_dadda_cla32_fa233_or0;
  assign f_u_dadda_cla32_fa250_and0 = f_u_dadda_cla32_fa234_or0 & f_u_dadda_cla32_fa233_or0;
  assign f_u_dadda_cla32_fa250_xor1 = f_u_dadda_cla32_fa250_xor0 ^ f_u_dadda_cla32_fa232_or0;
  assign f_u_dadda_cla32_fa250_and1 = f_u_dadda_cla32_fa250_xor0 & f_u_dadda_cla32_fa232_or0;
  assign f_u_dadda_cla32_fa250_or0 = f_u_dadda_cla32_fa250_and0 | f_u_dadda_cla32_fa250_and1;
  assign f_u_dadda_cla32_fa251_xor0 = f_u_dadda_cla32_fa231_or0 ^ f_u_dadda_cla32_fa230_or0;
  assign f_u_dadda_cla32_fa251_and0 = f_u_dadda_cla32_fa231_or0 & f_u_dadda_cla32_fa230_or0;
  assign f_u_dadda_cla32_fa251_xor1 = f_u_dadda_cla32_fa251_xor0 ^ f_u_dadda_cla32_fa229_or0;
  assign f_u_dadda_cla32_fa251_and1 = f_u_dadda_cla32_fa251_xor0 & f_u_dadda_cla32_fa229_or0;
  assign f_u_dadda_cla32_fa251_or0 = f_u_dadda_cla32_fa251_and0 | f_u_dadda_cla32_fa251_and1;
  assign f_u_dadda_cla32_fa252_xor0 = f_u_dadda_cla32_fa228_or0 ^ f_u_dadda_cla32_fa227_or0;
  assign f_u_dadda_cla32_fa252_and0 = f_u_dadda_cla32_fa228_or0 & f_u_dadda_cla32_fa227_or0;
  assign f_u_dadda_cla32_fa252_xor1 = f_u_dadda_cla32_fa252_xor0 ^ f_u_dadda_cla32_fa226_or0;
  assign f_u_dadda_cla32_fa252_and1 = f_u_dadda_cla32_fa252_xor0 & f_u_dadda_cla32_fa226_or0;
  assign f_u_dadda_cla32_fa252_or0 = f_u_dadda_cla32_fa252_and0 | f_u_dadda_cla32_fa252_and1;
  assign f_u_dadda_cla32_and_26_2 = a[26] & b[2];
  assign f_u_dadda_cla32_and_25_3 = a[25] & b[3];
  assign f_u_dadda_cla32_fa253_xor0 = f_u_dadda_cla32_fa225_or0 ^ f_u_dadda_cla32_and_26_2;
  assign f_u_dadda_cla32_fa253_and0 = f_u_dadda_cla32_fa225_or0 & f_u_dadda_cla32_and_26_2;
  assign f_u_dadda_cla32_fa253_xor1 = f_u_dadda_cla32_fa253_xor0 ^ f_u_dadda_cla32_and_25_3;
  assign f_u_dadda_cla32_fa253_and1 = f_u_dadda_cla32_fa253_xor0 & f_u_dadda_cla32_and_25_3;
  assign f_u_dadda_cla32_fa253_or0 = f_u_dadda_cla32_fa253_and0 | f_u_dadda_cla32_fa253_and1;
  assign f_u_dadda_cla32_and_24_4 = a[24] & b[4];
  assign f_u_dadda_cla32_and_23_5 = a[23] & b[5];
  assign f_u_dadda_cla32_and_22_6 = a[22] & b[6];
  assign f_u_dadda_cla32_fa254_xor0 = f_u_dadda_cla32_and_24_4 ^ f_u_dadda_cla32_and_23_5;
  assign f_u_dadda_cla32_fa254_and0 = f_u_dadda_cla32_and_24_4 & f_u_dadda_cla32_and_23_5;
  assign f_u_dadda_cla32_fa254_xor1 = f_u_dadda_cla32_fa254_xor0 ^ f_u_dadda_cla32_and_22_6;
  assign f_u_dadda_cla32_fa254_and1 = f_u_dadda_cla32_fa254_xor0 & f_u_dadda_cla32_and_22_6;
  assign f_u_dadda_cla32_fa254_or0 = f_u_dadda_cla32_fa254_and0 | f_u_dadda_cla32_fa254_and1;
  assign f_u_dadda_cla32_and_21_7 = a[21] & b[7];
  assign f_u_dadda_cla32_and_20_8 = a[20] & b[8];
  assign f_u_dadda_cla32_and_19_9 = a[19] & b[9];
  assign f_u_dadda_cla32_fa255_xor0 = f_u_dadda_cla32_and_21_7 ^ f_u_dadda_cla32_and_20_8;
  assign f_u_dadda_cla32_fa255_and0 = f_u_dadda_cla32_and_21_7 & f_u_dadda_cla32_and_20_8;
  assign f_u_dadda_cla32_fa255_xor1 = f_u_dadda_cla32_fa255_xor0 ^ f_u_dadda_cla32_and_19_9;
  assign f_u_dadda_cla32_fa255_and1 = f_u_dadda_cla32_fa255_xor0 & f_u_dadda_cla32_and_19_9;
  assign f_u_dadda_cla32_fa255_or0 = f_u_dadda_cla32_fa255_and0 | f_u_dadda_cla32_fa255_and1;
  assign f_u_dadda_cla32_and_18_10 = a[18] & b[10];
  assign f_u_dadda_cla32_and_17_11 = a[17] & b[11];
  assign f_u_dadda_cla32_and_16_12 = a[16] & b[12];
  assign f_u_dadda_cla32_fa256_xor0 = f_u_dadda_cla32_and_18_10 ^ f_u_dadda_cla32_and_17_11;
  assign f_u_dadda_cla32_fa256_and0 = f_u_dadda_cla32_and_18_10 & f_u_dadda_cla32_and_17_11;
  assign f_u_dadda_cla32_fa256_xor1 = f_u_dadda_cla32_fa256_xor0 ^ f_u_dadda_cla32_and_16_12;
  assign f_u_dadda_cla32_fa256_and1 = f_u_dadda_cla32_fa256_xor0 & f_u_dadda_cla32_and_16_12;
  assign f_u_dadda_cla32_fa256_or0 = f_u_dadda_cla32_fa256_and0 | f_u_dadda_cla32_fa256_and1;
  assign f_u_dadda_cla32_and_15_13 = a[15] & b[13];
  assign f_u_dadda_cla32_and_14_14 = a[14] & b[14];
  assign f_u_dadda_cla32_and_13_15 = a[13] & b[15];
  assign f_u_dadda_cla32_fa257_xor0 = f_u_dadda_cla32_and_15_13 ^ f_u_dadda_cla32_and_14_14;
  assign f_u_dadda_cla32_fa257_and0 = f_u_dadda_cla32_and_15_13 & f_u_dadda_cla32_and_14_14;
  assign f_u_dadda_cla32_fa257_xor1 = f_u_dadda_cla32_fa257_xor0 ^ f_u_dadda_cla32_and_13_15;
  assign f_u_dadda_cla32_fa257_and1 = f_u_dadda_cla32_fa257_xor0 & f_u_dadda_cla32_and_13_15;
  assign f_u_dadda_cla32_fa257_or0 = f_u_dadda_cla32_fa257_and0 | f_u_dadda_cla32_fa257_and1;
  assign f_u_dadda_cla32_and_12_16 = a[12] & b[16];
  assign f_u_dadda_cla32_and_11_17 = a[11] & b[17];
  assign f_u_dadda_cla32_and_10_18 = a[10] & b[18];
  assign f_u_dadda_cla32_fa258_xor0 = f_u_dadda_cla32_and_12_16 ^ f_u_dadda_cla32_and_11_17;
  assign f_u_dadda_cla32_fa258_and0 = f_u_dadda_cla32_and_12_16 & f_u_dadda_cla32_and_11_17;
  assign f_u_dadda_cla32_fa258_xor1 = f_u_dadda_cla32_fa258_xor0 ^ f_u_dadda_cla32_and_10_18;
  assign f_u_dadda_cla32_fa258_and1 = f_u_dadda_cla32_fa258_xor0 & f_u_dadda_cla32_and_10_18;
  assign f_u_dadda_cla32_fa258_or0 = f_u_dadda_cla32_fa258_and0 | f_u_dadda_cla32_fa258_and1;
  assign f_u_dadda_cla32_and_9_19 = a[9] & b[19];
  assign f_u_dadda_cla32_and_8_20 = a[8] & b[20];
  assign f_u_dadda_cla32_and_7_21 = a[7] & b[21];
  assign f_u_dadda_cla32_fa259_xor0 = f_u_dadda_cla32_and_9_19 ^ f_u_dadda_cla32_and_8_20;
  assign f_u_dadda_cla32_fa259_and0 = f_u_dadda_cla32_and_9_19 & f_u_dadda_cla32_and_8_20;
  assign f_u_dadda_cla32_fa259_xor1 = f_u_dadda_cla32_fa259_xor0 ^ f_u_dadda_cla32_and_7_21;
  assign f_u_dadda_cla32_fa259_and1 = f_u_dadda_cla32_fa259_xor0 & f_u_dadda_cla32_and_7_21;
  assign f_u_dadda_cla32_fa259_or0 = f_u_dadda_cla32_fa259_and0 | f_u_dadda_cla32_fa259_and1;
  assign f_u_dadda_cla32_and_6_22 = a[6] & b[22];
  assign f_u_dadda_cla32_and_5_23 = a[5] & b[23];
  assign f_u_dadda_cla32_and_4_24 = a[4] & b[24];
  assign f_u_dadda_cla32_fa260_xor0 = f_u_dadda_cla32_and_6_22 ^ f_u_dadda_cla32_and_5_23;
  assign f_u_dadda_cla32_fa260_and0 = f_u_dadda_cla32_and_6_22 & f_u_dadda_cla32_and_5_23;
  assign f_u_dadda_cla32_fa260_xor1 = f_u_dadda_cla32_fa260_xor0 ^ f_u_dadda_cla32_and_4_24;
  assign f_u_dadda_cla32_fa260_and1 = f_u_dadda_cla32_fa260_xor0 & f_u_dadda_cla32_and_4_24;
  assign f_u_dadda_cla32_fa260_or0 = f_u_dadda_cla32_fa260_and0 | f_u_dadda_cla32_fa260_and1;
  assign f_u_dadda_cla32_and_3_25 = a[3] & b[25];
  assign f_u_dadda_cla32_and_2_26 = a[2] & b[26];
  assign f_u_dadda_cla32_and_1_27 = a[1] & b[27];
  assign f_u_dadda_cla32_fa261_xor0 = f_u_dadda_cla32_and_3_25 ^ f_u_dadda_cla32_and_2_26;
  assign f_u_dadda_cla32_fa261_and0 = f_u_dadda_cla32_and_3_25 & f_u_dadda_cla32_and_2_26;
  assign f_u_dadda_cla32_fa261_xor1 = f_u_dadda_cla32_fa261_xor0 ^ f_u_dadda_cla32_and_1_27;
  assign f_u_dadda_cla32_fa261_and1 = f_u_dadda_cla32_fa261_xor0 & f_u_dadda_cla32_and_1_27;
  assign f_u_dadda_cla32_fa261_or0 = f_u_dadda_cla32_fa261_and0 | f_u_dadda_cla32_fa261_and1;
  assign f_u_dadda_cla32_and_0_28 = a[0] & b[28];
  assign f_u_dadda_cla32_fa262_xor0 = f_u_dadda_cla32_and_0_28 ^ f_u_dadda_cla32_ha0_xor0;
  assign f_u_dadda_cla32_fa262_and0 = f_u_dadda_cla32_and_0_28 & f_u_dadda_cla32_ha0_xor0;
  assign f_u_dadda_cla32_fa262_xor1 = f_u_dadda_cla32_fa262_xor0 ^ f_u_dadda_cla32_fa246_xor1;
  assign f_u_dadda_cla32_fa262_and1 = f_u_dadda_cla32_fa262_xor0 & f_u_dadda_cla32_fa246_xor1;
  assign f_u_dadda_cla32_fa262_or0 = f_u_dadda_cla32_fa262_and0 | f_u_dadda_cla32_fa262_and1;
  assign f_u_dadda_cla32_fa263_xor0 = f_u_dadda_cla32_fa247_xor1 ^ f_u_dadda_cla32_fa248_xor1;
  assign f_u_dadda_cla32_fa263_and0 = f_u_dadda_cla32_fa247_xor1 & f_u_dadda_cla32_fa248_xor1;
  assign f_u_dadda_cla32_fa263_xor1 = f_u_dadda_cla32_fa263_xor0 ^ f_u_dadda_cla32_fa249_xor1;
  assign f_u_dadda_cla32_fa263_and1 = f_u_dadda_cla32_fa263_xor0 & f_u_dadda_cla32_fa249_xor1;
  assign f_u_dadda_cla32_fa263_or0 = f_u_dadda_cla32_fa263_and0 | f_u_dadda_cla32_fa263_and1;
  assign f_u_dadda_cla32_fa264_xor0 = f_u_dadda_cla32_fa250_xor1 ^ f_u_dadda_cla32_fa251_xor1;
  assign f_u_dadda_cla32_fa264_and0 = f_u_dadda_cla32_fa250_xor1 & f_u_dadda_cla32_fa251_xor1;
  assign f_u_dadda_cla32_fa264_xor1 = f_u_dadda_cla32_fa264_xor0 ^ f_u_dadda_cla32_fa252_xor1;
  assign f_u_dadda_cla32_fa264_and1 = f_u_dadda_cla32_fa264_xor0 & f_u_dadda_cla32_fa252_xor1;
  assign f_u_dadda_cla32_fa264_or0 = f_u_dadda_cla32_fa264_and0 | f_u_dadda_cla32_fa264_and1;
  assign f_u_dadda_cla32_fa265_xor0 = f_u_dadda_cla32_fa253_xor1 ^ f_u_dadda_cla32_fa254_xor1;
  assign f_u_dadda_cla32_fa265_and0 = f_u_dadda_cla32_fa253_xor1 & f_u_dadda_cla32_fa254_xor1;
  assign f_u_dadda_cla32_fa265_xor1 = f_u_dadda_cla32_fa265_xor0 ^ f_u_dadda_cla32_fa255_xor1;
  assign f_u_dadda_cla32_fa265_and1 = f_u_dadda_cla32_fa265_xor0 & f_u_dadda_cla32_fa255_xor1;
  assign f_u_dadda_cla32_fa265_or0 = f_u_dadda_cla32_fa265_and0 | f_u_dadda_cla32_fa265_and1;
  assign f_u_dadda_cla32_fa266_xor0 = f_u_dadda_cla32_fa256_xor1 ^ f_u_dadda_cla32_fa257_xor1;
  assign f_u_dadda_cla32_fa266_and0 = f_u_dadda_cla32_fa256_xor1 & f_u_dadda_cla32_fa257_xor1;
  assign f_u_dadda_cla32_fa266_xor1 = f_u_dadda_cla32_fa266_xor0 ^ f_u_dadda_cla32_fa258_xor1;
  assign f_u_dadda_cla32_fa266_and1 = f_u_dadda_cla32_fa266_xor0 & f_u_dadda_cla32_fa258_xor1;
  assign f_u_dadda_cla32_fa266_or0 = f_u_dadda_cla32_fa266_and0 | f_u_dadda_cla32_fa266_and1;
  assign f_u_dadda_cla32_fa267_xor0 = f_u_dadda_cla32_fa259_xor1 ^ f_u_dadda_cla32_fa260_xor1;
  assign f_u_dadda_cla32_fa267_and0 = f_u_dadda_cla32_fa259_xor1 & f_u_dadda_cla32_fa260_xor1;
  assign f_u_dadda_cla32_fa267_xor1 = f_u_dadda_cla32_fa267_xor0 ^ f_u_dadda_cla32_fa261_xor1;
  assign f_u_dadda_cla32_fa267_and1 = f_u_dadda_cla32_fa267_xor0 & f_u_dadda_cla32_fa261_xor1;
  assign f_u_dadda_cla32_fa267_or0 = f_u_dadda_cla32_fa267_and0 | f_u_dadda_cla32_fa267_and1;
  assign f_u_dadda_cla32_fa268_xor0 = f_u_dadda_cla32_fa267_or0 ^ f_u_dadda_cla32_fa266_or0;
  assign f_u_dadda_cla32_fa268_and0 = f_u_dadda_cla32_fa267_or0 & f_u_dadda_cla32_fa266_or0;
  assign f_u_dadda_cla32_fa268_xor1 = f_u_dadda_cla32_fa268_xor0 ^ f_u_dadda_cla32_fa265_or0;
  assign f_u_dadda_cla32_fa268_and1 = f_u_dadda_cla32_fa268_xor0 & f_u_dadda_cla32_fa265_or0;
  assign f_u_dadda_cla32_fa268_or0 = f_u_dadda_cla32_fa268_and0 | f_u_dadda_cla32_fa268_and1;
  assign f_u_dadda_cla32_fa269_xor0 = f_u_dadda_cla32_fa264_or0 ^ f_u_dadda_cla32_fa263_or0;
  assign f_u_dadda_cla32_fa269_and0 = f_u_dadda_cla32_fa264_or0 & f_u_dadda_cla32_fa263_or0;
  assign f_u_dadda_cla32_fa269_xor1 = f_u_dadda_cla32_fa269_xor0 ^ f_u_dadda_cla32_fa262_or0;
  assign f_u_dadda_cla32_fa269_and1 = f_u_dadda_cla32_fa269_xor0 & f_u_dadda_cla32_fa262_or0;
  assign f_u_dadda_cla32_fa269_or0 = f_u_dadda_cla32_fa269_and0 | f_u_dadda_cla32_fa269_and1;
  assign f_u_dadda_cla32_fa270_xor0 = f_u_dadda_cla32_fa261_or0 ^ f_u_dadda_cla32_fa260_or0;
  assign f_u_dadda_cla32_fa270_and0 = f_u_dadda_cla32_fa261_or0 & f_u_dadda_cla32_fa260_or0;
  assign f_u_dadda_cla32_fa270_xor1 = f_u_dadda_cla32_fa270_xor0 ^ f_u_dadda_cla32_fa259_or0;
  assign f_u_dadda_cla32_fa270_and1 = f_u_dadda_cla32_fa270_xor0 & f_u_dadda_cla32_fa259_or0;
  assign f_u_dadda_cla32_fa270_or0 = f_u_dadda_cla32_fa270_and0 | f_u_dadda_cla32_fa270_and1;
  assign f_u_dadda_cla32_fa271_xor0 = f_u_dadda_cla32_fa258_or0 ^ f_u_dadda_cla32_fa257_or0;
  assign f_u_dadda_cla32_fa271_and0 = f_u_dadda_cla32_fa258_or0 & f_u_dadda_cla32_fa257_or0;
  assign f_u_dadda_cla32_fa271_xor1 = f_u_dadda_cla32_fa271_xor0 ^ f_u_dadda_cla32_fa256_or0;
  assign f_u_dadda_cla32_fa271_and1 = f_u_dadda_cla32_fa271_xor0 & f_u_dadda_cla32_fa256_or0;
  assign f_u_dadda_cla32_fa271_or0 = f_u_dadda_cla32_fa271_and0 | f_u_dadda_cla32_fa271_and1;
  assign f_u_dadda_cla32_fa272_xor0 = f_u_dadda_cla32_fa255_or0 ^ f_u_dadda_cla32_fa254_or0;
  assign f_u_dadda_cla32_fa272_and0 = f_u_dadda_cla32_fa255_or0 & f_u_dadda_cla32_fa254_or0;
  assign f_u_dadda_cla32_fa272_xor1 = f_u_dadda_cla32_fa272_xor0 ^ f_u_dadda_cla32_fa253_or0;
  assign f_u_dadda_cla32_fa272_and1 = f_u_dadda_cla32_fa272_xor0 & f_u_dadda_cla32_fa253_or0;
  assign f_u_dadda_cla32_fa272_or0 = f_u_dadda_cla32_fa272_and0 | f_u_dadda_cla32_fa272_and1;
  assign f_u_dadda_cla32_fa273_xor0 = f_u_dadda_cla32_fa252_or0 ^ f_u_dadda_cla32_fa251_or0;
  assign f_u_dadda_cla32_fa273_and0 = f_u_dadda_cla32_fa252_or0 & f_u_dadda_cla32_fa251_or0;
  assign f_u_dadda_cla32_fa273_xor1 = f_u_dadda_cla32_fa273_xor0 ^ f_u_dadda_cla32_fa250_or0;
  assign f_u_dadda_cla32_fa273_and1 = f_u_dadda_cla32_fa273_xor0 & f_u_dadda_cla32_fa250_or0;
  assign f_u_dadda_cla32_fa273_or0 = f_u_dadda_cla32_fa273_and0 | f_u_dadda_cla32_fa273_and1;
  assign f_u_dadda_cla32_fa274_xor0 = f_u_dadda_cla32_fa249_or0 ^ f_u_dadda_cla32_fa248_or0;
  assign f_u_dadda_cla32_fa274_and0 = f_u_dadda_cla32_fa249_or0 & f_u_dadda_cla32_fa248_or0;
  assign f_u_dadda_cla32_fa274_xor1 = f_u_dadda_cla32_fa274_xor0 ^ f_u_dadda_cla32_fa247_or0;
  assign f_u_dadda_cla32_fa274_and1 = f_u_dadda_cla32_fa274_xor0 & f_u_dadda_cla32_fa247_or0;
  assign f_u_dadda_cla32_fa274_or0 = f_u_dadda_cla32_fa274_and0 | f_u_dadda_cla32_fa274_and1;
  assign f_u_dadda_cla32_and_25_4 = a[25] & b[4];
  assign f_u_dadda_cla32_and_24_5 = a[24] & b[5];
  assign f_u_dadda_cla32_fa275_xor0 = f_u_dadda_cla32_fa246_or0 ^ f_u_dadda_cla32_and_25_4;
  assign f_u_dadda_cla32_fa275_and0 = f_u_dadda_cla32_fa246_or0 & f_u_dadda_cla32_and_25_4;
  assign f_u_dadda_cla32_fa275_xor1 = f_u_dadda_cla32_fa275_xor0 ^ f_u_dadda_cla32_and_24_5;
  assign f_u_dadda_cla32_fa275_and1 = f_u_dadda_cla32_fa275_xor0 & f_u_dadda_cla32_and_24_5;
  assign f_u_dadda_cla32_fa275_or0 = f_u_dadda_cla32_fa275_and0 | f_u_dadda_cla32_fa275_and1;
  assign f_u_dadda_cla32_and_23_6 = a[23] & b[6];
  assign f_u_dadda_cla32_and_22_7 = a[22] & b[7];
  assign f_u_dadda_cla32_and_21_8 = a[21] & b[8];
  assign f_u_dadda_cla32_fa276_xor0 = f_u_dadda_cla32_and_23_6 ^ f_u_dadda_cla32_and_22_7;
  assign f_u_dadda_cla32_fa276_and0 = f_u_dadda_cla32_and_23_6 & f_u_dadda_cla32_and_22_7;
  assign f_u_dadda_cla32_fa276_xor1 = f_u_dadda_cla32_fa276_xor0 ^ f_u_dadda_cla32_and_21_8;
  assign f_u_dadda_cla32_fa276_and1 = f_u_dadda_cla32_fa276_xor0 & f_u_dadda_cla32_and_21_8;
  assign f_u_dadda_cla32_fa276_or0 = f_u_dadda_cla32_fa276_and0 | f_u_dadda_cla32_fa276_and1;
  assign f_u_dadda_cla32_and_20_9 = a[20] & b[9];
  assign f_u_dadda_cla32_and_19_10 = a[19] & b[10];
  assign f_u_dadda_cla32_and_18_11 = a[18] & b[11];
  assign f_u_dadda_cla32_fa277_xor0 = f_u_dadda_cla32_and_20_9 ^ f_u_dadda_cla32_and_19_10;
  assign f_u_dadda_cla32_fa277_and0 = f_u_dadda_cla32_and_20_9 & f_u_dadda_cla32_and_19_10;
  assign f_u_dadda_cla32_fa277_xor1 = f_u_dadda_cla32_fa277_xor0 ^ f_u_dadda_cla32_and_18_11;
  assign f_u_dadda_cla32_fa277_and1 = f_u_dadda_cla32_fa277_xor0 & f_u_dadda_cla32_and_18_11;
  assign f_u_dadda_cla32_fa277_or0 = f_u_dadda_cla32_fa277_and0 | f_u_dadda_cla32_fa277_and1;
  assign f_u_dadda_cla32_and_17_12 = a[17] & b[12];
  assign f_u_dadda_cla32_and_16_13 = a[16] & b[13];
  assign f_u_dadda_cla32_and_15_14 = a[15] & b[14];
  assign f_u_dadda_cla32_fa278_xor0 = f_u_dadda_cla32_and_17_12 ^ f_u_dadda_cla32_and_16_13;
  assign f_u_dadda_cla32_fa278_and0 = f_u_dadda_cla32_and_17_12 & f_u_dadda_cla32_and_16_13;
  assign f_u_dadda_cla32_fa278_xor1 = f_u_dadda_cla32_fa278_xor0 ^ f_u_dadda_cla32_and_15_14;
  assign f_u_dadda_cla32_fa278_and1 = f_u_dadda_cla32_fa278_xor0 & f_u_dadda_cla32_and_15_14;
  assign f_u_dadda_cla32_fa278_or0 = f_u_dadda_cla32_fa278_and0 | f_u_dadda_cla32_fa278_and1;
  assign f_u_dadda_cla32_and_14_15 = a[14] & b[15];
  assign f_u_dadda_cla32_and_13_16 = a[13] & b[16];
  assign f_u_dadda_cla32_and_12_17 = a[12] & b[17];
  assign f_u_dadda_cla32_fa279_xor0 = f_u_dadda_cla32_and_14_15 ^ f_u_dadda_cla32_and_13_16;
  assign f_u_dadda_cla32_fa279_and0 = f_u_dadda_cla32_and_14_15 & f_u_dadda_cla32_and_13_16;
  assign f_u_dadda_cla32_fa279_xor1 = f_u_dadda_cla32_fa279_xor0 ^ f_u_dadda_cla32_and_12_17;
  assign f_u_dadda_cla32_fa279_and1 = f_u_dadda_cla32_fa279_xor0 & f_u_dadda_cla32_and_12_17;
  assign f_u_dadda_cla32_fa279_or0 = f_u_dadda_cla32_fa279_and0 | f_u_dadda_cla32_fa279_and1;
  assign f_u_dadda_cla32_and_11_18 = a[11] & b[18];
  assign f_u_dadda_cla32_and_10_19 = a[10] & b[19];
  assign f_u_dadda_cla32_and_9_20 = a[9] & b[20];
  assign f_u_dadda_cla32_fa280_xor0 = f_u_dadda_cla32_and_11_18 ^ f_u_dadda_cla32_and_10_19;
  assign f_u_dadda_cla32_fa280_and0 = f_u_dadda_cla32_and_11_18 & f_u_dadda_cla32_and_10_19;
  assign f_u_dadda_cla32_fa280_xor1 = f_u_dadda_cla32_fa280_xor0 ^ f_u_dadda_cla32_and_9_20;
  assign f_u_dadda_cla32_fa280_and1 = f_u_dadda_cla32_fa280_xor0 & f_u_dadda_cla32_and_9_20;
  assign f_u_dadda_cla32_fa280_or0 = f_u_dadda_cla32_fa280_and0 | f_u_dadda_cla32_fa280_and1;
  assign f_u_dadda_cla32_and_8_21 = a[8] & b[21];
  assign f_u_dadda_cla32_and_7_22 = a[7] & b[22];
  assign f_u_dadda_cla32_and_6_23 = a[6] & b[23];
  assign f_u_dadda_cla32_fa281_xor0 = f_u_dadda_cla32_and_8_21 ^ f_u_dadda_cla32_and_7_22;
  assign f_u_dadda_cla32_fa281_and0 = f_u_dadda_cla32_and_8_21 & f_u_dadda_cla32_and_7_22;
  assign f_u_dadda_cla32_fa281_xor1 = f_u_dadda_cla32_fa281_xor0 ^ f_u_dadda_cla32_and_6_23;
  assign f_u_dadda_cla32_fa281_and1 = f_u_dadda_cla32_fa281_xor0 & f_u_dadda_cla32_and_6_23;
  assign f_u_dadda_cla32_fa281_or0 = f_u_dadda_cla32_fa281_and0 | f_u_dadda_cla32_fa281_and1;
  assign f_u_dadda_cla32_and_5_24 = a[5] & b[24];
  assign f_u_dadda_cla32_and_4_25 = a[4] & b[25];
  assign f_u_dadda_cla32_and_3_26 = a[3] & b[26];
  assign f_u_dadda_cla32_fa282_xor0 = f_u_dadda_cla32_and_5_24 ^ f_u_dadda_cla32_and_4_25;
  assign f_u_dadda_cla32_fa282_and0 = f_u_dadda_cla32_and_5_24 & f_u_dadda_cla32_and_4_25;
  assign f_u_dadda_cla32_fa282_xor1 = f_u_dadda_cla32_fa282_xor0 ^ f_u_dadda_cla32_and_3_26;
  assign f_u_dadda_cla32_fa282_and1 = f_u_dadda_cla32_fa282_xor0 & f_u_dadda_cla32_and_3_26;
  assign f_u_dadda_cla32_fa282_or0 = f_u_dadda_cla32_fa282_and0 | f_u_dadda_cla32_fa282_and1;
  assign f_u_dadda_cla32_and_2_27 = a[2] & b[27];
  assign f_u_dadda_cla32_and_1_28 = a[1] & b[28];
  assign f_u_dadda_cla32_and_0_29 = a[0] & b[29];
  assign f_u_dadda_cla32_fa283_xor0 = f_u_dadda_cla32_and_2_27 ^ f_u_dadda_cla32_and_1_28;
  assign f_u_dadda_cla32_fa283_and0 = f_u_dadda_cla32_and_2_27 & f_u_dadda_cla32_and_1_28;
  assign f_u_dadda_cla32_fa283_xor1 = f_u_dadda_cla32_fa283_xor0 ^ f_u_dadda_cla32_and_0_29;
  assign f_u_dadda_cla32_fa283_and1 = f_u_dadda_cla32_fa283_xor0 & f_u_dadda_cla32_and_0_29;
  assign f_u_dadda_cla32_fa283_or0 = f_u_dadda_cla32_fa283_and0 | f_u_dadda_cla32_fa283_and1;
  assign f_u_dadda_cla32_fa284_xor0 = f_u_dadda_cla32_fa0_xor1 ^ f_u_dadda_cla32_ha1_xor0;
  assign f_u_dadda_cla32_fa284_and0 = f_u_dadda_cla32_fa0_xor1 & f_u_dadda_cla32_ha1_xor0;
  assign f_u_dadda_cla32_fa284_xor1 = f_u_dadda_cla32_fa284_xor0 ^ f_u_dadda_cla32_fa268_xor1;
  assign f_u_dadda_cla32_fa284_and1 = f_u_dadda_cla32_fa284_xor0 & f_u_dadda_cla32_fa268_xor1;
  assign f_u_dadda_cla32_fa284_or0 = f_u_dadda_cla32_fa284_and0 | f_u_dadda_cla32_fa284_and1;
  assign f_u_dadda_cla32_fa285_xor0 = f_u_dadda_cla32_fa269_xor1 ^ f_u_dadda_cla32_fa270_xor1;
  assign f_u_dadda_cla32_fa285_and0 = f_u_dadda_cla32_fa269_xor1 & f_u_dadda_cla32_fa270_xor1;
  assign f_u_dadda_cla32_fa285_xor1 = f_u_dadda_cla32_fa285_xor0 ^ f_u_dadda_cla32_fa271_xor1;
  assign f_u_dadda_cla32_fa285_and1 = f_u_dadda_cla32_fa285_xor0 & f_u_dadda_cla32_fa271_xor1;
  assign f_u_dadda_cla32_fa285_or0 = f_u_dadda_cla32_fa285_and0 | f_u_dadda_cla32_fa285_and1;
  assign f_u_dadda_cla32_fa286_xor0 = f_u_dadda_cla32_fa272_xor1 ^ f_u_dadda_cla32_fa273_xor1;
  assign f_u_dadda_cla32_fa286_and0 = f_u_dadda_cla32_fa272_xor1 & f_u_dadda_cla32_fa273_xor1;
  assign f_u_dadda_cla32_fa286_xor1 = f_u_dadda_cla32_fa286_xor0 ^ f_u_dadda_cla32_fa274_xor1;
  assign f_u_dadda_cla32_fa286_and1 = f_u_dadda_cla32_fa286_xor0 & f_u_dadda_cla32_fa274_xor1;
  assign f_u_dadda_cla32_fa286_or0 = f_u_dadda_cla32_fa286_and0 | f_u_dadda_cla32_fa286_and1;
  assign f_u_dadda_cla32_fa287_xor0 = f_u_dadda_cla32_fa275_xor1 ^ f_u_dadda_cla32_fa276_xor1;
  assign f_u_dadda_cla32_fa287_and0 = f_u_dadda_cla32_fa275_xor1 & f_u_dadda_cla32_fa276_xor1;
  assign f_u_dadda_cla32_fa287_xor1 = f_u_dadda_cla32_fa287_xor0 ^ f_u_dadda_cla32_fa277_xor1;
  assign f_u_dadda_cla32_fa287_and1 = f_u_dadda_cla32_fa287_xor0 & f_u_dadda_cla32_fa277_xor1;
  assign f_u_dadda_cla32_fa287_or0 = f_u_dadda_cla32_fa287_and0 | f_u_dadda_cla32_fa287_and1;
  assign f_u_dadda_cla32_fa288_xor0 = f_u_dadda_cla32_fa278_xor1 ^ f_u_dadda_cla32_fa279_xor1;
  assign f_u_dadda_cla32_fa288_and0 = f_u_dadda_cla32_fa278_xor1 & f_u_dadda_cla32_fa279_xor1;
  assign f_u_dadda_cla32_fa288_xor1 = f_u_dadda_cla32_fa288_xor0 ^ f_u_dadda_cla32_fa280_xor1;
  assign f_u_dadda_cla32_fa288_and1 = f_u_dadda_cla32_fa288_xor0 & f_u_dadda_cla32_fa280_xor1;
  assign f_u_dadda_cla32_fa288_or0 = f_u_dadda_cla32_fa288_and0 | f_u_dadda_cla32_fa288_and1;
  assign f_u_dadda_cla32_fa289_xor0 = f_u_dadda_cla32_fa281_xor1 ^ f_u_dadda_cla32_fa282_xor1;
  assign f_u_dadda_cla32_fa289_and0 = f_u_dadda_cla32_fa281_xor1 & f_u_dadda_cla32_fa282_xor1;
  assign f_u_dadda_cla32_fa289_xor1 = f_u_dadda_cla32_fa289_xor0 ^ f_u_dadda_cla32_fa283_xor1;
  assign f_u_dadda_cla32_fa289_and1 = f_u_dadda_cla32_fa289_xor0 & f_u_dadda_cla32_fa283_xor1;
  assign f_u_dadda_cla32_fa289_or0 = f_u_dadda_cla32_fa289_and0 | f_u_dadda_cla32_fa289_and1;
  assign f_u_dadda_cla32_fa290_xor0 = f_u_dadda_cla32_fa289_or0 ^ f_u_dadda_cla32_fa288_or0;
  assign f_u_dadda_cla32_fa290_and0 = f_u_dadda_cla32_fa289_or0 & f_u_dadda_cla32_fa288_or0;
  assign f_u_dadda_cla32_fa290_xor1 = f_u_dadda_cla32_fa290_xor0 ^ f_u_dadda_cla32_fa287_or0;
  assign f_u_dadda_cla32_fa290_and1 = f_u_dadda_cla32_fa290_xor0 & f_u_dadda_cla32_fa287_or0;
  assign f_u_dadda_cla32_fa290_or0 = f_u_dadda_cla32_fa290_and0 | f_u_dadda_cla32_fa290_and1;
  assign f_u_dadda_cla32_fa291_xor0 = f_u_dadda_cla32_fa286_or0 ^ f_u_dadda_cla32_fa285_or0;
  assign f_u_dadda_cla32_fa291_and0 = f_u_dadda_cla32_fa286_or0 & f_u_dadda_cla32_fa285_or0;
  assign f_u_dadda_cla32_fa291_xor1 = f_u_dadda_cla32_fa291_xor0 ^ f_u_dadda_cla32_fa284_or0;
  assign f_u_dadda_cla32_fa291_and1 = f_u_dadda_cla32_fa291_xor0 & f_u_dadda_cla32_fa284_or0;
  assign f_u_dadda_cla32_fa291_or0 = f_u_dadda_cla32_fa291_and0 | f_u_dadda_cla32_fa291_and1;
  assign f_u_dadda_cla32_fa292_xor0 = f_u_dadda_cla32_fa283_or0 ^ f_u_dadda_cla32_fa282_or0;
  assign f_u_dadda_cla32_fa292_and0 = f_u_dadda_cla32_fa283_or0 & f_u_dadda_cla32_fa282_or0;
  assign f_u_dadda_cla32_fa292_xor1 = f_u_dadda_cla32_fa292_xor0 ^ f_u_dadda_cla32_fa281_or0;
  assign f_u_dadda_cla32_fa292_and1 = f_u_dadda_cla32_fa292_xor0 & f_u_dadda_cla32_fa281_or0;
  assign f_u_dadda_cla32_fa292_or0 = f_u_dadda_cla32_fa292_and0 | f_u_dadda_cla32_fa292_and1;
  assign f_u_dadda_cla32_fa293_xor0 = f_u_dadda_cla32_fa280_or0 ^ f_u_dadda_cla32_fa279_or0;
  assign f_u_dadda_cla32_fa293_and0 = f_u_dadda_cla32_fa280_or0 & f_u_dadda_cla32_fa279_or0;
  assign f_u_dadda_cla32_fa293_xor1 = f_u_dadda_cla32_fa293_xor0 ^ f_u_dadda_cla32_fa278_or0;
  assign f_u_dadda_cla32_fa293_and1 = f_u_dadda_cla32_fa293_xor0 & f_u_dadda_cla32_fa278_or0;
  assign f_u_dadda_cla32_fa293_or0 = f_u_dadda_cla32_fa293_and0 | f_u_dadda_cla32_fa293_and1;
  assign f_u_dadda_cla32_fa294_xor0 = f_u_dadda_cla32_fa277_or0 ^ f_u_dadda_cla32_fa276_or0;
  assign f_u_dadda_cla32_fa294_and0 = f_u_dadda_cla32_fa277_or0 & f_u_dadda_cla32_fa276_or0;
  assign f_u_dadda_cla32_fa294_xor1 = f_u_dadda_cla32_fa294_xor0 ^ f_u_dadda_cla32_fa275_or0;
  assign f_u_dadda_cla32_fa294_and1 = f_u_dadda_cla32_fa294_xor0 & f_u_dadda_cla32_fa275_or0;
  assign f_u_dadda_cla32_fa294_or0 = f_u_dadda_cla32_fa294_and0 | f_u_dadda_cla32_fa294_and1;
  assign f_u_dadda_cla32_fa295_xor0 = f_u_dadda_cla32_fa274_or0 ^ f_u_dadda_cla32_fa273_or0;
  assign f_u_dadda_cla32_fa295_and0 = f_u_dadda_cla32_fa274_or0 & f_u_dadda_cla32_fa273_or0;
  assign f_u_dadda_cla32_fa295_xor1 = f_u_dadda_cla32_fa295_xor0 ^ f_u_dadda_cla32_fa272_or0;
  assign f_u_dadda_cla32_fa295_and1 = f_u_dadda_cla32_fa295_xor0 & f_u_dadda_cla32_fa272_or0;
  assign f_u_dadda_cla32_fa295_or0 = f_u_dadda_cla32_fa295_and0 | f_u_dadda_cla32_fa295_and1;
  assign f_u_dadda_cla32_fa296_xor0 = f_u_dadda_cla32_fa271_or0 ^ f_u_dadda_cla32_fa270_or0;
  assign f_u_dadda_cla32_fa296_and0 = f_u_dadda_cla32_fa271_or0 & f_u_dadda_cla32_fa270_or0;
  assign f_u_dadda_cla32_fa296_xor1 = f_u_dadda_cla32_fa296_xor0 ^ f_u_dadda_cla32_fa269_or0;
  assign f_u_dadda_cla32_fa296_and1 = f_u_dadda_cla32_fa296_xor0 & f_u_dadda_cla32_fa269_or0;
  assign f_u_dadda_cla32_fa296_or0 = f_u_dadda_cla32_fa296_and0 | f_u_dadda_cla32_fa296_and1;
  assign f_u_dadda_cla32_and_24_6 = a[24] & b[6];
  assign f_u_dadda_cla32_and_23_7 = a[23] & b[7];
  assign f_u_dadda_cla32_fa297_xor0 = f_u_dadda_cla32_fa268_or0 ^ f_u_dadda_cla32_and_24_6;
  assign f_u_dadda_cla32_fa297_and0 = f_u_dadda_cla32_fa268_or0 & f_u_dadda_cla32_and_24_6;
  assign f_u_dadda_cla32_fa297_xor1 = f_u_dadda_cla32_fa297_xor0 ^ f_u_dadda_cla32_and_23_7;
  assign f_u_dadda_cla32_fa297_and1 = f_u_dadda_cla32_fa297_xor0 & f_u_dadda_cla32_and_23_7;
  assign f_u_dadda_cla32_fa297_or0 = f_u_dadda_cla32_fa297_and0 | f_u_dadda_cla32_fa297_and1;
  assign f_u_dadda_cla32_and_22_8 = a[22] & b[8];
  assign f_u_dadda_cla32_and_21_9 = a[21] & b[9];
  assign f_u_dadda_cla32_and_20_10 = a[20] & b[10];
  assign f_u_dadda_cla32_fa298_xor0 = f_u_dadda_cla32_and_22_8 ^ f_u_dadda_cla32_and_21_9;
  assign f_u_dadda_cla32_fa298_and0 = f_u_dadda_cla32_and_22_8 & f_u_dadda_cla32_and_21_9;
  assign f_u_dadda_cla32_fa298_xor1 = f_u_dadda_cla32_fa298_xor0 ^ f_u_dadda_cla32_and_20_10;
  assign f_u_dadda_cla32_fa298_and1 = f_u_dadda_cla32_fa298_xor0 & f_u_dadda_cla32_and_20_10;
  assign f_u_dadda_cla32_fa298_or0 = f_u_dadda_cla32_fa298_and0 | f_u_dadda_cla32_fa298_and1;
  assign f_u_dadda_cla32_and_19_11 = a[19] & b[11];
  assign f_u_dadda_cla32_and_18_12 = a[18] & b[12];
  assign f_u_dadda_cla32_and_17_13 = a[17] & b[13];
  assign f_u_dadda_cla32_fa299_xor0 = f_u_dadda_cla32_and_19_11 ^ f_u_dadda_cla32_and_18_12;
  assign f_u_dadda_cla32_fa299_and0 = f_u_dadda_cla32_and_19_11 & f_u_dadda_cla32_and_18_12;
  assign f_u_dadda_cla32_fa299_xor1 = f_u_dadda_cla32_fa299_xor0 ^ f_u_dadda_cla32_and_17_13;
  assign f_u_dadda_cla32_fa299_and1 = f_u_dadda_cla32_fa299_xor0 & f_u_dadda_cla32_and_17_13;
  assign f_u_dadda_cla32_fa299_or0 = f_u_dadda_cla32_fa299_and0 | f_u_dadda_cla32_fa299_and1;
  assign f_u_dadda_cla32_and_16_14 = a[16] & b[14];
  assign f_u_dadda_cla32_and_15_15 = a[15] & b[15];
  assign f_u_dadda_cla32_and_14_16 = a[14] & b[16];
  assign f_u_dadda_cla32_fa300_xor0 = f_u_dadda_cla32_and_16_14 ^ f_u_dadda_cla32_and_15_15;
  assign f_u_dadda_cla32_fa300_and0 = f_u_dadda_cla32_and_16_14 & f_u_dadda_cla32_and_15_15;
  assign f_u_dadda_cla32_fa300_xor1 = f_u_dadda_cla32_fa300_xor0 ^ f_u_dadda_cla32_and_14_16;
  assign f_u_dadda_cla32_fa300_and1 = f_u_dadda_cla32_fa300_xor0 & f_u_dadda_cla32_and_14_16;
  assign f_u_dadda_cla32_fa300_or0 = f_u_dadda_cla32_fa300_and0 | f_u_dadda_cla32_fa300_and1;
  assign f_u_dadda_cla32_and_13_17 = a[13] & b[17];
  assign f_u_dadda_cla32_and_12_18 = a[12] & b[18];
  assign f_u_dadda_cla32_and_11_19 = a[11] & b[19];
  assign f_u_dadda_cla32_fa301_xor0 = f_u_dadda_cla32_and_13_17 ^ f_u_dadda_cla32_and_12_18;
  assign f_u_dadda_cla32_fa301_and0 = f_u_dadda_cla32_and_13_17 & f_u_dadda_cla32_and_12_18;
  assign f_u_dadda_cla32_fa301_xor1 = f_u_dadda_cla32_fa301_xor0 ^ f_u_dadda_cla32_and_11_19;
  assign f_u_dadda_cla32_fa301_and1 = f_u_dadda_cla32_fa301_xor0 & f_u_dadda_cla32_and_11_19;
  assign f_u_dadda_cla32_fa301_or0 = f_u_dadda_cla32_fa301_and0 | f_u_dadda_cla32_fa301_and1;
  assign f_u_dadda_cla32_and_10_20 = a[10] & b[20];
  assign f_u_dadda_cla32_and_9_21 = a[9] & b[21];
  assign f_u_dadda_cla32_and_8_22 = a[8] & b[22];
  assign f_u_dadda_cla32_fa302_xor0 = f_u_dadda_cla32_and_10_20 ^ f_u_dadda_cla32_and_9_21;
  assign f_u_dadda_cla32_fa302_and0 = f_u_dadda_cla32_and_10_20 & f_u_dadda_cla32_and_9_21;
  assign f_u_dadda_cla32_fa302_xor1 = f_u_dadda_cla32_fa302_xor0 ^ f_u_dadda_cla32_and_8_22;
  assign f_u_dadda_cla32_fa302_and1 = f_u_dadda_cla32_fa302_xor0 & f_u_dadda_cla32_and_8_22;
  assign f_u_dadda_cla32_fa302_or0 = f_u_dadda_cla32_fa302_and0 | f_u_dadda_cla32_fa302_and1;
  assign f_u_dadda_cla32_and_7_23 = a[7] & b[23];
  assign f_u_dadda_cla32_and_6_24 = a[6] & b[24];
  assign f_u_dadda_cla32_and_5_25 = a[5] & b[25];
  assign f_u_dadda_cla32_fa303_xor0 = f_u_dadda_cla32_and_7_23 ^ f_u_dadda_cla32_and_6_24;
  assign f_u_dadda_cla32_fa303_and0 = f_u_dadda_cla32_and_7_23 & f_u_dadda_cla32_and_6_24;
  assign f_u_dadda_cla32_fa303_xor1 = f_u_dadda_cla32_fa303_xor0 ^ f_u_dadda_cla32_and_5_25;
  assign f_u_dadda_cla32_fa303_and1 = f_u_dadda_cla32_fa303_xor0 & f_u_dadda_cla32_and_5_25;
  assign f_u_dadda_cla32_fa303_or0 = f_u_dadda_cla32_fa303_and0 | f_u_dadda_cla32_fa303_and1;
  assign f_u_dadda_cla32_and_4_26 = a[4] & b[26];
  assign f_u_dadda_cla32_and_3_27 = a[3] & b[27];
  assign f_u_dadda_cla32_and_2_28 = a[2] & b[28];
  assign f_u_dadda_cla32_fa304_xor0 = f_u_dadda_cla32_and_4_26 ^ f_u_dadda_cla32_and_3_27;
  assign f_u_dadda_cla32_fa304_and0 = f_u_dadda_cla32_and_4_26 & f_u_dadda_cla32_and_3_27;
  assign f_u_dadda_cla32_fa304_xor1 = f_u_dadda_cla32_fa304_xor0 ^ f_u_dadda_cla32_and_2_28;
  assign f_u_dadda_cla32_fa304_and1 = f_u_dadda_cla32_fa304_xor0 & f_u_dadda_cla32_and_2_28;
  assign f_u_dadda_cla32_fa304_or0 = f_u_dadda_cla32_fa304_and0 | f_u_dadda_cla32_fa304_and1;
  assign f_u_dadda_cla32_and_1_29 = a[1] & b[29];
  assign f_u_dadda_cla32_and_0_30 = a[0] & b[30];
  assign f_u_dadda_cla32_fa305_xor0 = f_u_dadda_cla32_and_1_29 ^ f_u_dadda_cla32_and_0_30;
  assign f_u_dadda_cla32_fa305_and0 = f_u_dadda_cla32_and_1_29 & f_u_dadda_cla32_and_0_30;
  assign f_u_dadda_cla32_fa305_xor1 = f_u_dadda_cla32_fa305_xor0 ^ f_u_dadda_cla32_fa1_xor1;
  assign f_u_dadda_cla32_fa305_and1 = f_u_dadda_cla32_fa305_xor0 & f_u_dadda_cla32_fa1_xor1;
  assign f_u_dadda_cla32_fa305_or0 = f_u_dadda_cla32_fa305_and0 | f_u_dadda_cla32_fa305_and1;
  assign f_u_dadda_cla32_fa306_xor0 = f_u_dadda_cla32_fa2_xor1 ^ f_u_dadda_cla32_ha2_xor0;
  assign f_u_dadda_cla32_fa306_and0 = f_u_dadda_cla32_fa2_xor1 & f_u_dadda_cla32_ha2_xor0;
  assign f_u_dadda_cla32_fa306_xor1 = f_u_dadda_cla32_fa306_xor0 ^ f_u_dadda_cla32_fa290_xor1;
  assign f_u_dadda_cla32_fa306_and1 = f_u_dadda_cla32_fa306_xor0 & f_u_dadda_cla32_fa290_xor1;
  assign f_u_dadda_cla32_fa306_or0 = f_u_dadda_cla32_fa306_and0 | f_u_dadda_cla32_fa306_and1;
  assign f_u_dadda_cla32_fa307_xor0 = f_u_dadda_cla32_fa291_xor1 ^ f_u_dadda_cla32_fa292_xor1;
  assign f_u_dadda_cla32_fa307_and0 = f_u_dadda_cla32_fa291_xor1 & f_u_dadda_cla32_fa292_xor1;
  assign f_u_dadda_cla32_fa307_xor1 = f_u_dadda_cla32_fa307_xor0 ^ f_u_dadda_cla32_fa293_xor1;
  assign f_u_dadda_cla32_fa307_and1 = f_u_dadda_cla32_fa307_xor0 & f_u_dadda_cla32_fa293_xor1;
  assign f_u_dadda_cla32_fa307_or0 = f_u_dadda_cla32_fa307_and0 | f_u_dadda_cla32_fa307_and1;
  assign f_u_dadda_cla32_fa308_xor0 = f_u_dadda_cla32_fa294_xor1 ^ f_u_dadda_cla32_fa295_xor1;
  assign f_u_dadda_cla32_fa308_and0 = f_u_dadda_cla32_fa294_xor1 & f_u_dadda_cla32_fa295_xor1;
  assign f_u_dadda_cla32_fa308_xor1 = f_u_dadda_cla32_fa308_xor0 ^ f_u_dadda_cla32_fa296_xor1;
  assign f_u_dadda_cla32_fa308_and1 = f_u_dadda_cla32_fa308_xor0 & f_u_dadda_cla32_fa296_xor1;
  assign f_u_dadda_cla32_fa308_or0 = f_u_dadda_cla32_fa308_and0 | f_u_dadda_cla32_fa308_and1;
  assign f_u_dadda_cla32_fa309_xor0 = f_u_dadda_cla32_fa297_xor1 ^ f_u_dadda_cla32_fa298_xor1;
  assign f_u_dadda_cla32_fa309_and0 = f_u_dadda_cla32_fa297_xor1 & f_u_dadda_cla32_fa298_xor1;
  assign f_u_dadda_cla32_fa309_xor1 = f_u_dadda_cla32_fa309_xor0 ^ f_u_dadda_cla32_fa299_xor1;
  assign f_u_dadda_cla32_fa309_and1 = f_u_dadda_cla32_fa309_xor0 & f_u_dadda_cla32_fa299_xor1;
  assign f_u_dadda_cla32_fa309_or0 = f_u_dadda_cla32_fa309_and0 | f_u_dadda_cla32_fa309_and1;
  assign f_u_dadda_cla32_fa310_xor0 = f_u_dadda_cla32_fa300_xor1 ^ f_u_dadda_cla32_fa301_xor1;
  assign f_u_dadda_cla32_fa310_and0 = f_u_dadda_cla32_fa300_xor1 & f_u_dadda_cla32_fa301_xor1;
  assign f_u_dadda_cla32_fa310_xor1 = f_u_dadda_cla32_fa310_xor0 ^ f_u_dadda_cla32_fa302_xor1;
  assign f_u_dadda_cla32_fa310_and1 = f_u_dadda_cla32_fa310_xor0 & f_u_dadda_cla32_fa302_xor1;
  assign f_u_dadda_cla32_fa310_or0 = f_u_dadda_cla32_fa310_and0 | f_u_dadda_cla32_fa310_and1;
  assign f_u_dadda_cla32_fa311_xor0 = f_u_dadda_cla32_fa303_xor1 ^ f_u_dadda_cla32_fa304_xor1;
  assign f_u_dadda_cla32_fa311_and0 = f_u_dadda_cla32_fa303_xor1 & f_u_dadda_cla32_fa304_xor1;
  assign f_u_dadda_cla32_fa311_xor1 = f_u_dadda_cla32_fa311_xor0 ^ f_u_dadda_cla32_fa305_xor1;
  assign f_u_dadda_cla32_fa311_and1 = f_u_dadda_cla32_fa311_xor0 & f_u_dadda_cla32_fa305_xor1;
  assign f_u_dadda_cla32_fa311_or0 = f_u_dadda_cla32_fa311_and0 | f_u_dadda_cla32_fa311_and1;
  assign f_u_dadda_cla32_fa312_xor0 = f_u_dadda_cla32_fa311_or0 ^ f_u_dadda_cla32_fa310_or0;
  assign f_u_dadda_cla32_fa312_and0 = f_u_dadda_cla32_fa311_or0 & f_u_dadda_cla32_fa310_or0;
  assign f_u_dadda_cla32_fa312_xor1 = f_u_dadda_cla32_fa312_xor0 ^ f_u_dadda_cla32_fa309_or0;
  assign f_u_dadda_cla32_fa312_and1 = f_u_dadda_cla32_fa312_xor0 & f_u_dadda_cla32_fa309_or0;
  assign f_u_dadda_cla32_fa312_or0 = f_u_dadda_cla32_fa312_and0 | f_u_dadda_cla32_fa312_and1;
  assign f_u_dadda_cla32_fa313_xor0 = f_u_dadda_cla32_fa308_or0 ^ f_u_dadda_cla32_fa307_or0;
  assign f_u_dadda_cla32_fa313_and0 = f_u_dadda_cla32_fa308_or0 & f_u_dadda_cla32_fa307_or0;
  assign f_u_dadda_cla32_fa313_xor1 = f_u_dadda_cla32_fa313_xor0 ^ f_u_dadda_cla32_fa306_or0;
  assign f_u_dadda_cla32_fa313_and1 = f_u_dadda_cla32_fa313_xor0 & f_u_dadda_cla32_fa306_or0;
  assign f_u_dadda_cla32_fa313_or0 = f_u_dadda_cla32_fa313_and0 | f_u_dadda_cla32_fa313_and1;
  assign f_u_dadda_cla32_fa314_xor0 = f_u_dadda_cla32_fa305_or0 ^ f_u_dadda_cla32_fa304_or0;
  assign f_u_dadda_cla32_fa314_and0 = f_u_dadda_cla32_fa305_or0 & f_u_dadda_cla32_fa304_or0;
  assign f_u_dadda_cla32_fa314_xor1 = f_u_dadda_cla32_fa314_xor0 ^ f_u_dadda_cla32_fa303_or0;
  assign f_u_dadda_cla32_fa314_and1 = f_u_dadda_cla32_fa314_xor0 & f_u_dadda_cla32_fa303_or0;
  assign f_u_dadda_cla32_fa314_or0 = f_u_dadda_cla32_fa314_and0 | f_u_dadda_cla32_fa314_and1;
  assign f_u_dadda_cla32_fa315_xor0 = f_u_dadda_cla32_fa302_or0 ^ f_u_dadda_cla32_fa301_or0;
  assign f_u_dadda_cla32_fa315_and0 = f_u_dadda_cla32_fa302_or0 & f_u_dadda_cla32_fa301_or0;
  assign f_u_dadda_cla32_fa315_xor1 = f_u_dadda_cla32_fa315_xor0 ^ f_u_dadda_cla32_fa300_or0;
  assign f_u_dadda_cla32_fa315_and1 = f_u_dadda_cla32_fa315_xor0 & f_u_dadda_cla32_fa300_or0;
  assign f_u_dadda_cla32_fa315_or0 = f_u_dadda_cla32_fa315_and0 | f_u_dadda_cla32_fa315_and1;
  assign f_u_dadda_cla32_fa316_xor0 = f_u_dadda_cla32_fa299_or0 ^ f_u_dadda_cla32_fa298_or0;
  assign f_u_dadda_cla32_fa316_and0 = f_u_dadda_cla32_fa299_or0 & f_u_dadda_cla32_fa298_or0;
  assign f_u_dadda_cla32_fa316_xor1 = f_u_dadda_cla32_fa316_xor0 ^ f_u_dadda_cla32_fa297_or0;
  assign f_u_dadda_cla32_fa316_and1 = f_u_dadda_cla32_fa316_xor0 & f_u_dadda_cla32_fa297_or0;
  assign f_u_dadda_cla32_fa316_or0 = f_u_dadda_cla32_fa316_and0 | f_u_dadda_cla32_fa316_and1;
  assign f_u_dadda_cla32_fa317_xor0 = f_u_dadda_cla32_fa296_or0 ^ f_u_dadda_cla32_fa295_or0;
  assign f_u_dadda_cla32_fa317_and0 = f_u_dadda_cla32_fa296_or0 & f_u_dadda_cla32_fa295_or0;
  assign f_u_dadda_cla32_fa317_xor1 = f_u_dadda_cla32_fa317_xor0 ^ f_u_dadda_cla32_fa294_or0;
  assign f_u_dadda_cla32_fa317_and1 = f_u_dadda_cla32_fa317_xor0 & f_u_dadda_cla32_fa294_or0;
  assign f_u_dadda_cla32_fa317_or0 = f_u_dadda_cla32_fa317_and0 | f_u_dadda_cla32_fa317_and1;
  assign f_u_dadda_cla32_fa318_xor0 = f_u_dadda_cla32_fa293_or0 ^ f_u_dadda_cla32_fa292_or0;
  assign f_u_dadda_cla32_fa318_and0 = f_u_dadda_cla32_fa293_or0 & f_u_dadda_cla32_fa292_or0;
  assign f_u_dadda_cla32_fa318_xor1 = f_u_dadda_cla32_fa318_xor0 ^ f_u_dadda_cla32_fa291_or0;
  assign f_u_dadda_cla32_fa318_and1 = f_u_dadda_cla32_fa318_xor0 & f_u_dadda_cla32_fa291_or0;
  assign f_u_dadda_cla32_fa318_or0 = f_u_dadda_cla32_fa318_and0 | f_u_dadda_cla32_fa318_and1;
  assign f_u_dadda_cla32_and_23_8 = a[23] & b[8];
  assign f_u_dadda_cla32_and_22_9 = a[22] & b[9];
  assign f_u_dadda_cla32_fa319_xor0 = f_u_dadda_cla32_fa290_or0 ^ f_u_dadda_cla32_and_23_8;
  assign f_u_dadda_cla32_fa319_and0 = f_u_dadda_cla32_fa290_or0 & f_u_dadda_cla32_and_23_8;
  assign f_u_dadda_cla32_fa319_xor1 = f_u_dadda_cla32_fa319_xor0 ^ f_u_dadda_cla32_and_22_9;
  assign f_u_dadda_cla32_fa319_and1 = f_u_dadda_cla32_fa319_xor0 & f_u_dadda_cla32_and_22_9;
  assign f_u_dadda_cla32_fa319_or0 = f_u_dadda_cla32_fa319_and0 | f_u_dadda_cla32_fa319_and1;
  assign f_u_dadda_cla32_and_21_10 = a[21] & b[10];
  assign f_u_dadda_cla32_and_20_11 = a[20] & b[11];
  assign f_u_dadda_cla32_and_19_12 = a[19] & b[12];
  assign f_u_dadda_cla32_fa320_xor0 = f_u_dadda_cla32_and_21_10 ^ f_u_dadda_cla32_and_20_11;
  assign f_u_dadda_cla32_fa320_and0 = f_u_dadda_cla32_and_21_10 & f_u_dadda_cla32_and_20_11;
  assign f_u_dadda_cla32_fa320_xor1 = f_u_dadda_cla32_fa320_xor0 ^ f_u_dadda_cla32_and_19_12;
  assign f_u_dadda_cla32_fa320_and1 = f_u_dadda_cla32_fa320_xor0 & f_u_dadda_cla32_and_19_12;
  assign f_u_dadda_cla32_fa320_or0 = f_u_dadda_cla32_fa320_and0 | f_u_dadda_cla32_fa320_and1;
  assign f_u_dadda_cla32_and_18_13 = a[18] & b[13];
  assign f_u_dadda_cla32_and_17_14 = a[17] & b[14];
  assign f_u_dadda_cla32_and_16_15 = a[16] & b[15];
  assign f_u_dadda_cla32_fa321_xor0 = f_u_dadda_cla32_and_18_13 ^ f_u_dadda_cla32_and_17_14;
  assign f_u_dadda_cla32_fa321_and0 = f_u_dadda_cla32_and_18_13 & f_u_dadda_cla32_and_17_14;
  assign f_u_dadda_cla32_fa321_xor1 = f_u_dadda_cla32_fa321_xor0 ^ f_u_dadda_cla32_and_16_15;
  assign f_u_dadda_cla32_fa321_and1 = f_u_dadda_cla32_fa321_xor0 & f_u_dadda_cla32_and_16_15;
  assign f_u_dadda_cla32_fa321_or0 = f_u_dadda_cla32_fa321_and0 | f_u_dadda_cla32_fa321_and1;
  assign f_u_dadda_cla32_and_15_16 = a[15] & b[16];
  assign f_u_dadda_cla32_and_14_17 = a[14] & b[17];
  assign f_u_dadda_cla32_and_13_18 = a[13] & b[18];
  assign f_u_dadda_cla32_fa322_xor0 = f_u_dadda_cla32_and_15_16 ^ f_u_dadda_cla32_and_14_17;
  assign f_u_dadda_cla32_fa322_and0 = f_u_dadda_cla32_and_15_16 & f_u_dadda_cla32_and_14_17;
  assign f_u_dadda_cla32_fa322_xor1 = f_u_dadda_cla32_fa322_xor0 ^ f_u_dadda_cla32_and_13_18;
  assign f_u_dadda_cla32_fa322_and1 = f_u_dadda_cla32_fa322_xor0 & f_u_dadda_cla32_and_13_18;
  assign f_u_dadda_cla32_fa322_or0 = f_u_dadda_cla32_fa322_and0 | f_u_dadda_cla32_fa322_and1;
  assign f_u_dadda_cla32_and_12_19 = a[12] & b[19];
  assign f_u_dadda_cla32_and_11_20 = a[11] & b[20];
  assign f_u_dadda_cla32_and_10_21 = a[10] & b[21];
  assign f_u_dadda_cla32_fa323_xor0 = f_u_dadda_cla32_and_12_19 ^ f_u_dadda_cla32_and_11_20;
  assign f_u_dadda_cla32_fa323_and0 = f_u_dadda_cla32_and_12_19 & f_u_dadda_cla32_and_11_20;
  assign f_u_dadda_cla32_fa323_xor1 = f_u_dadda_cla32_fa323_xor0 ^ f_u_dadda_cla32_and_10_21;
  assign f_u_dadda_cla32_fa323_and1 = f_u_dadda_cla32_fa323_xor0 & f_u_dadda_cla32_and_10_21;
  assign f_u_dadda_cla32_fa323_or0 = f_u_dadda_cla32_fa323_and0 | f_u_dadda_cla32_fa323_and1;
  assign f_u_dadda_cla32_and_9_22 = a[9] & b[22];
  assign f_u_dadda_cla32_and_8_23 = a[8] & b[23];
  assign f_u_dadda_cla32_and_7_24 = a[7] & b[24];
  assign f_u_dadda_cla32_fa324_xor0 = f_u_dadda_cla32_and_9_22 ^ f_u_dadda_cla32_and_8_23;
  assign f_u_dadda_cla32_fa324_and0 = f_u_dadda_cla32_and_9_22 & f_u_dadda_cla32_and_8_23;
  assign f_u_dadda_cla32_fa324_xor1 = f_u_dadda_cla32_fa324_xor0 ^ f_u_dadda_cla32_and_7_24;
  assign f_u_dadda_cla32_fa324_and1 = f_u_dadda_cla32_fa324_xor0 & f_u_dadda_cla32_and_7_24;
  assign f_u_dadda_cla32_fa324_or0 = f_u_dadda_cla32_fa324_and0 | f_u_dadda_cla32_fa324_and1;
  assign f_u_dadda_cla32_and_6_25 = a[6] & b[25];
  assign f_u_dadda_cla32_and_5_26 = a[5] & b[26];
  assign f_u_dadda_cla32_and_4_27 = a[4] & b[27];
  assign f_u_dadda_cla32_fa325_xor0 = f_u_dadda_cla32_and_6_25 ^ f_u_dadda_cla32_and_5_26;
  assign f_u_dadda_cla32_fa325_and0 = f_u_dadda_cla32_and_6_25 & f_u_dadda_cla32_and_5_26;
  assign f_u_dadda_cla32_fa325_xor1 = f_u_dadda_cla32_fa325_xor0 ^ f_u_dadda_cla32_and_4_27;
  assign f_u_dadda_cla32_fa325_and1 = f_u_dadda_cla32_fa325_xor0 & f_u_dadda_cla32_and_4_27;
  assign f_u_dadda_cla32_fa325_or0 = f_u_dadda_cla32_fa325_and0 | f_u_dadda_cla32_fa325_and1;
  assign f_u_dadda_cla32_and_3_28 = a[3] & b[28];
  assign f_u_dadda_cla32_and_2_29 = a[2] & b[29];
  assign f_u_dadda_cla32_and_1_30 = a[1] & b[30];
  assign f_u_dadda_cla32_fa326_xor0 = f_u_dadda_cla32_and_3_28 ^ f_u_dadda_cla32_and_2_29;
  assign f_u_dadda_cla32_fa326_and0 = f_u_dadda_cla32_and_3_28 & f_u_dadda_cla32_and_2_29;
  assign f_u_dadda_cla32_fa326_xor1 = f_u_dadda_cla32_fa326_xor0 ^ f_u_dadda_cla32_and_1_30;
  assign f_u_dadda_cla32_fa326_and1 = f_u_dadda_cla32_fa326_xor0 & f_u_dadda_cla32_and_1_30;
  assign f_u_dadda_cla32_fa326_or0 = f_u_dadda_cla32_fa326_and0 | f_u_dadda_cla32_fa326_and1;
  assign f_u_dadda_cla32_and_0_31 = a[0] & b[31];
  assign f_u_dadda_cla32_fa327_xor0 = f_u_dadda_cla32_and_0_31 ^ f_u_dadda_cla32_fa3_xor1;
  assign f_u_dadda_cla32_fa327_and0 = f_u_dadda_cla32_and_0_31 & f_u_dadda_cla32_fa3_xor1;
  assign f_u_dadda_cla32_fa327_xor1 = f_u_dadda_cla32_fa327_xor0 ^ f_u_dadda_cla32_fa4_xor1;
  assign f_u_dadda_cla32_fa327_and1 = f_u_dadda_cla32_fa327_xor0 & f_u_dadda_cla32_fa4_xor1;
  assign f_u_dadda_cla32_fa327_or0 = f_u_dadda_cla32_fa327_and0 | f_u_dadda_cla32_fa327_and1;
  assign f_u_dadda_cla32_fa328_xor0 = f_u_dadda_cla32_fa5_xor1 ^ f_u_dadda_cla32_ha3_xor0;
  assign f_u_dadda_cla32_fa328_and0 = f_u_dadda_cla32_fa5_xor1 & f_u_dadda_cla32_ha3_xor0;
  assign f_u_dadda_cla32_fa328_xor1 = f_u_dadda_cla32_fa328_xor0 ^ f_u_dadda_cla32_fa312_xor1;
  assign f_u_dadda_cla32_fa328_and1 = f_u_dadda_cla32_fa328_xor0 & f_u_dadda_cla32_fa312_xor1;
  assign f_u_dadda_cla32_fa328_or0 = f_u_dadda_cla32_fa328_and0 | f_u_dadda_cla32_fa328_and1;
  assign f_u_dadda_cla32_fa329_xor0 = f_u_dadda_cla32_fa313_xor1 ^ f_u_dadda_cla32_fa314_xor1;
  assign f_u_dadda_cla32_fa329_and0 = f_u_dadda_cla32_fa313_xor1 & f_u_dadda_cla32_fa314_xor1;
  assign f_u_dadda_cla32_fa329_xor1 = f_u_dadda_cla32_fa329_xor0 ^ f_u_dadda_cla32_fa315_xor1;
  assign f_u_dadda_cla32_fa329_and1 = f_u_dadda_cla32_fa329_xor0 & f_u_dadda_cla32_fa315_xor1;
  assign f_u_dadda_cla32_fa329_or0 = f_u_dadda_cla32_fa329_and0 | f_u_dadda_cla32_fa329_and1;
  assign f_u_dadda_cla32_fa330_xor0 = f_u_dadda_cla32_fa316_xor1 ^ f_u_dadda_cla32_fa317_xor1;
  assign f_u_dadda_cla32_fa330_and0 = f_u_dadda_cla32_fa316_xor1 & f_u_dadda_cla32_fa317_xor1;
  assign f_u_dadda_cla32_fa330_xor1 = f_u_dadda_cla32_fa330_xor0 ^ f_u_dadda_cla32_fa318_xor1;
  assign f_u_dadda_cla32_fa330_and1 = f_u_dadda_cla32_fa330_xor0 & f_u_dadda_cla32_fa318_xor1;
  assign f_u_dadda_cla32_fa330_or0 = f_u_dadda_cla32_fa330_and0 | f_u_dadda_cla32_fa330_and1;
  assign f_u_dadda_cla32_fa331_xor0 = f_u_dadda_cla32_fa319_xor1 ^ f_u_dadda_cla32_fa320_xor1;
  assign f_u_dadda_cla32_fa331_and0 = f_u_dadda_cla32_fa319_xor1 & f_u_dadda_cla32_fa320_xor1;
  assign f_u_dadda_cla32_fa331_xor1 = f_u_dadda_cla32_fa331_xor0 ^ f_u_dadda_cla32_fa321_xor1;
  assign f_u_dadda_cla32_fa331_and1 = f_u_dadda_cla32_fa331_xor0 & f_u_dadda_cla32_fa321_xor1;
  assign f_u_dadda_cla32_fa331_or0 = f_u_dadda_cla32_fa331_and0 | f_u_dadda_cla32_fa331_and1;
  assign f_u_dadda_cla32_fa332_xor0 = f_u_dadda_cla32_fa322_xor1 ^ f_u_dadda_cla32_fa323_xor1;
  assign f_u_dadda_cla32_fa332_and0 = f_u_dadda_cla32_fa322_xor1 & f_u_dadda_cla32_fa323_xor1;
  assign f_u_dadda_cla32_fa332_xor1 = f_u_dadda_cla32_fa332_xor0 ^ f_u_dadda_cla32_fa324_xor1;
  assign f_u_dadda_cla32_fa332_and1 = f_u_dadda_cla32_fa332_xor0 & f_u_dadda_cla32_fa324_xor1;
  assign f_u_dadda_cla32_fa332_or0 = f_u_dadda_cla32_fa332_and0 | f_u_dadda_cla32_fa332_and1;
  assign f_u_dadda_cla32_fa333_xor0 = f_u_dadda_cla32_fa325_xor1 ^ f_u_dadda_cla32_fa326_xor1;
  assign f_u_dadda_cla32_fa333_and0 = f_u_dadda_cla32_fa325_xor1 & f_u_dadda_cla32_fa326_xor1;
  assign f_u_dadda_cla32_fa333_xor1 = f_u_dadda_cla32_fa333_xor0 ^ f_u_dadda_cla32_fa327_xor1;
  assign f_u_dadda_cla32_fa333_and1 = f_u_dadda_cla32_fa333_xor0 & f_u_dadda_cla32_fa327_xor1;
  assign f_u_dadda_cla32_fa333_or0 = f_u_dadda_cla32_fa333_and0 | f_u_dadda_cla32_fa333_and1;
  assign f_u_dadda_cla32_fa334_xor0 = f_u_dadda_cla32_fa333_or0 ^ f_u_dadda_cla32_fa332_or0;
  assign f_u_dadda_cla32_fa334_and0 = f_u_dadda_cla32_fa333_or0 & f_u_dadda_cla32_fa332_or0;
  assign f_u_dadda_cla32_fa334_xor1 = f_u_dadda_cla32_fa334_xor0 ^ f_u_dadda_cla32_fa331_or0;
  assign f_u_dadda_cla32_fa334_and1 = f_u_dadda_cla32_fa334_xor0 & f_u_dadda_cla32_fa331_or0;
  assign f_u_dadda_cla32_fa334_or0 = f_u_dadda_cla32_fa334_and0 | f_u_dadda_cla32_fa334_and1;
  assign f_u_dadda_cla32_fa335_xor0 = f_u_dadda_cla32_fa330_or0 ^ f_u_dadda_cla32_fa329_or0;
  assign f_u_dadda_cla32_fa335_and0 = f_u_dadda_cla32_fa330_or0 & f_u_dadda_cla32_fa329_or0;
  assign f_u_dadda_cla32_fa335_xor1 = f_u_dadda_cla32_fa335_xor0 ^ f_u_dadda_cla32_fa328_or0;
  assign f_u_dadda_cla32_fa335_and1 = f_u_dadda_cla32_fa335_xor0 & f_u_dadda_cla32_fa328_or0;
  assign f_u_dadda_cla32_fa335_or0 = f_u_dadda_cla32_fa335_and0 | f_u_dadda_cla32_fa335_and1;
  assign f_u_dadda_cla32_fa336_xor0 = f_u_dadda_cla32_fa327_or0 ^ f_u_dadda_cla32_fa326_or0;
  assign f_u_dadda_cla32_fa336_and0 = f_u_dadda_cla32_fa327_or0 & f_u_dadda_cla32_fa326_or0;
  assign f_u_dadda_cla32_fa336_xor1 = f_u_dadda_cla32_fa336_xor0 ^ f_u_dadda_cla32_fa325_or0;
  assign f_u_dadda_cla32_fa336_and1 = f_u_dadda_cla32_fa336_xor0 & f_u_dadda_cla32_fa325_or0;
  assign f_u_dadda_cla32_fa336_or0 = f_u_dadda_cla32_fa336_and0 | f_u_dadda_cla32_fa336_and1;
  assign f_u_dadda_cla32_fa337_xor0 = f_u_dadda_cla32_fa324_or0 ^ f_u_dadda_cla32_fa323_or0;
  assign f_u_dadda_cla32_fa337_and0 = f_u_dadda_cla32_fa324_or0 & f_u_dadda_cla32_fa323_or0;
  assign f_u_dadda_cla32_fa337_xor1 = f_u_dadda_cla32_fa337_xor0 ^ f_u_dadda_cla32_fa322_or0;
  assign f_u_dadda_cla32_fa337_and1 = f_u_dadda_cla32_fa337_xor0 & f_u_dadda_cla32_fa322_or0;
  assign f_u_dadda_cla32_fa337_or0 = f_u_dadda_cla32_fa337_and0 | f_u_dadda_cla32_fa337_and1;
  assign f_u_dadda_cla32_fa338_xor0 = f_u_dadda_cla32_fa321_or0 ^ f_u_dadda_cla32_fa320_or0;
  assign f_u_dadda_cla32_fa338_and0 = f_u_dadda_cla32_fa321_or0 & f_u_dadda_cla32_fa320_or0;
  assign f_u_dadda_cla32_fa338_xor1 = f_u_dadda_cla32_fa338_xor0 ^ f_u_dadda_cla32_fa319_or0;
  assign f_u_dadda_cla32_fa338_and1 = f_u_dadda_cla32_fa338_xor0 & f_u_dadda_cla32_fa319_or0;
  assign f_u_dadda_cla32_fa338_or0 = f_u_dadda_cla32_fa338_and0 | f_u_dadda_cla32_fa338_and1;
  assign f_u_dadda_cla32_fa339_xor0 = f_u_dadda_cla32_fa318_or0 ^ f_u_dadda_cla32_fa317_or0;
  assign f_u_dadda_cla32_fa339_and0 = f_u_dadda_cla32_fa318_or0 & f_u_dadda_cla32_fa317_or0;
  assign f_u_dadda_cla32_fa339_xor1 = f_u_dadda_cla32_fa339_xor0 ^ f_u_dadda_cla32_fa316_or0;
  assign f_u_dadda_cla32_fa339_and1 = f_u_dadda_cla32_fa339_xor0 & f_u_dadda_cla32_fa316_or0;
  assign f_u_dadda_cla32_fa339_or0 = f_u_dadda_cla32_fa339_and0 | f_u_dadda_cla32_fa339_and1;
  assign f_u_dadda_cla32_fa340_xor0 = f_u_dadda_cla32_fa315_or0 ^ f_u_dadda_cla32_fa314_or0;
  assign f_u_dadda_cla32_fa340_and0 = f_u_dadda_cla32_fa315_or0 & f_u_dadda_cla32_fa314_or0;
  assign f_u_dadda_cla32_fa340_xor1 = f_u_dadda_cla32_fa340_xor0 ^ f_u_dadda_cla32_fa313_or0;
  assign f_u_dadda_cla32_fa340_and1 = f_u_dadda_cla32_fa340_xor0 & f_u_dadda_cla32_fa313_or0;
  assign f_u_dadda_cla32_fa340_or0 = f_u_dadda_cla32_fa340_and0 | f_u_dadda_cla32_fa340_and1;
  assign f_u_dadda_cla32_and_24_8 = a[24] & b[8];
  assign f_u_dadda_cla32_and_23_9 = a[23] & b[9];
  assign f_u_dadda_cla32_fa341_xor0 = f_u_dadda_cla32_fa312_or0 ^ f_u_dadda_cla32_and_24_8;
  assign f_u_dadda_cla32_fa341_and0 = f_u_dadda_cla32_fa312_or0 & f_u_dadda_cla32_and_24_8;
  assign f_u_dadda_cla32_fa341_xor1 = f_u_dadda_cla32_fa341_xor0 ^ f_u_dadda_cla32_and_23_9;
  assign f_u_dadda_cla32_fa341_and1 = f_u_dadda_cla32_fa341_xor0 & f_u_dadda_cla32_and_23_9;
  assign f_u_dadda_cla32_fa341_or0 = f_u_dadda_cla32_fa341_and0 | f_u_dadda_cla32_fa341_and1;
  assign f_u_dadda_cla32_and_22_10 = a[22] & b[10];
  assign f_u_dadda_cla32_and_21_11 = a[21] & b[11];
  assign f_u_dadda_cla32_and_20_12 = a[20] & b[12];
  assign f_u_dadda_cla32_fa342_xor0 = f_u_dadda_cla32_and_22_10 ^ f_u_dadda_cla32_and_21_11;
  assign f_u_dadda_cla32_fa342_and0 = f_u_dadda_cla32_and_22_10 & f_u_dadda_cla32_and_21_11;
  assign f_u_dadda_cla32_fa342_xor1 = f_u_dadda_cla32_fa342_xor0 ^ f_u_dadda_cla32_and_20_12;
  assign f_u_dadda_cla32_fa342_and1 = f_u_dadda_cla32_fa342_xor0 & f_u_dadda_cla32_and_20_12;
  assign f_u_dadda_cla32_fa342_or0 = f_u_dadda_cla32_fa342_and0 | f_u_dadda_cla32_fa342_and1;
  assign f_u_dadda_cla32_and_19_13 = a[19] & b[13];
  assign f_u_dadda_cla32_and_18_14 = a[18] & b[14];
  assign f_u_dadda_cla32_and_17_15 = a[17] & b[15];
  assign f_u_dadda_cla32_fa343_xor0 = f_u_dadda_cla32_and_19_13 ^ f_u_dadda_cla32_and_18_14;
  assign f_u_dadda_cla32_fa343_and0 = f_u_dadda_cla32_and_19_13 & f_u_dadda_cla32_and_18_14;
  assign f_u_dadda_cla32_fa343_xor1 = f_u_dadda_cla32_fa343_xor0 ^ f_u_dadda_cla32_and_17_15;
  assign f_u_dadda_cla32_fa343_and1 = f_u_dadda_cla32_fa343_xor0 & f_u_dadda_cla32_and_17_15;
  assign f_u_dadda_cla32_fa343_or0 = f_u_dadda_cla32_fa343_and0 | f_u_dadda_cla32_fa343_and1;
  assign f_u_dadda_cla32_and_16_16 = a[16] & b[16];
  assign f_u_dadda_cla32_and_15_17 = a[15] & b[17];
  assign f_u_dadda_cla32_and_14_18 = a[14] & b[18];
  assign f_u_dadda_cla32_fa344_xor0 = f_u_dadda_cla32_and_16_16 ^ f_u_dadda_cla32_and_15_17;
  assign f_u_dadda_cla32_fa344_and0 = f_u_dadda_cla32_and_16_16 & f_u_dadda_cla32_and_15_17;
  assign f_u_dadda_cla32_fa344_xor1 = f_u_dadda_cla32_fa344_xor0 ^ f_u_dadda_cla32_and_14_18;
  assign f_u_dadda_cla32_fa344_and1 = f_u_dadda_cla32_fa344_xor0 & f_u_dadda_cla32_and_14_18;
  assign f_u_dadda_cla32_fa344_or0 = f_u_dadda_cla32_fa344_and0 | f_u_dadda_cla32_fa344_and1;
  assign f_u_dadda_cla32_and_13_19 = a[13] & b[19];
  assign f_u_dadda_cla32_and_12_20 = a[12] & b[20];
  assign f_u_dadda_cla32_and_11_21 = a[11] & b[21];
  assign f_u_dadda_cla32_fa345_xor0 = f_u_dadda_cla32_and_13_19 ^ f_u_dadda_cla32_and_12_20;
  assign f_u_dadda_cla32_fa345_and0 = f_u_dadda_cla32_and_13_19 & f_u_dadda_cla32_and_12_20;
  assign f_u_dadda_cla32_fa345_xor1 = f_u_dadda_cla32_fa345_xor0 ^ f_u_dadda_cla32_and_11_21;
  assign f_u_dadda_cla32_fa345_and1 = f_u_dadda_cla32_fa345_xor0 & f_u_dadda_cla32_and_11_21;
  assign f_u_dadda_cla32_fa345_or0 = f_u_dadda_cla32_fa345_and0 | f_u_dadda_cla32_fa345_and1;
  assign f_u_dadda_cla32_and_10_22 = a[10] & b[22];
  assign f_u_dadda_cla32_and_9_23 = a[9] & b[23];
  assign f_u_dadda_cla32_and_8_24 = a[8] & b[24];
  assign f_u_dadda_cla32_fa346_xor0 = f_u_dadda_cla32_and_10_22 ^ f_u_dadda_cla32_and_9_23;
  assign f_u_dadda_cla32_fa346_and0 = f_u_dadda_cla32_and_10_22 & f_u_dadda_cla32_and_9_23;
  assign f_u_dadda_cla32_fa346_xor1 = f_u_dadda_cla32_fa346_xor0 ^ f_u_dadda_cla32_and_8_24;
  assign f_u_dadda_cla32_fa346_and1 = f_u_dadda_cla32_fa346_xor0 & f_u_dadda_cla32_and_8_24;
  assign f_u_dadda_cla32_fa346_or0 = f_u_dadda_cla32_fa346_and0 | f_u_dadda_cla32_fa346_and1;
  assign f_u_dadda_cla32_and_7_25 = a[7] & b[25];
  assign f_u_dadda_cla32_and_6_26 = a[6] & b[26];
  assign f_u_dadda_cla32_and_5_27 = a[5] & b[27];
  assign f_u_dadda_cla32_fa347_xor0 = f_u_dadda_cla32_and_7_25 ^ f_u_dadda_cla32_and_6_26;
  assign f_u_dadda_cla32_fa347_and0 = f_u_dadda_cla32_and_7_25 & f_u_dadda_cla32_and_6_26;
  assign f_u_dadda_cla32_fa347_xor1 = f_u_dadda_cla32_fa347_xor0 ^ f_u_dadda_cla32_and_5_27;
  assign f_u_dadda_cla32_fa347_and1 = f_u_dadda_cla32_fa347_xor0 & f_u_dadda_cla32_and_5_27;
  assign f_u_dadda_cla32_fa347_or0 = f_u_dadda_cla32_fa347_and0 | f_u_dadda_cla32_fa347_and1;
  assign f_u_dadda_cla32_and_4_28 = a[4] & b[28];
  assign f_u_dadda_cla32_and_3_29 = a[3] & b[29];
  assign f_u_dadda_cla32_and_2_30 = a[2] & b[30];
  assign f_u_dadda_cla32_fa348_xor0 = f_u_dadda_cla32_and_4_28 ^ f_u_dadda_cla32_and_3_29;
  assign f_u_dadda_cla32_fa348_and0 = f_u_dadda_cla32_and_4_28 & f_u_dadda_cla32_and_3_29;
  assign f_u_dadda_cla32_fa348_xor1 = f_u_dadda_cla32_fa348_xor0 ^ f_u_dadda_cla32_and_2_30;
  assign f_u_dadda_cla32_fa348_and1 = f_u_dadda_cla32_fa348_xor0 & f_u_dadda_cla32_and_2_30;
  assign f_u_dadda_cla32_fa348_or0 = f_u_dadda_cla32_fa348_and0 | f_u_dadda_cla32_fa348_and1;
  assign f_u_dadda_cla32_and_1_31 = a[1] & b[31];
  assign f_u_dadda_cla32_fa349_xor0 = f_u_dadda_cla32_and_1_31 ^ f_u_dadda_cla32_fa6_xor1;
  assign f_u_dadda_cla32_fa349_and0 = f_u_dadda_cla32_and_1_31 & f_u_dadda_cla32_fa6_xor1;
  assign f_u_dadda_cla32_fa349_xor1 = f_u_dadda_cla32_fa349_xor0 ^ f_u_dadda_cla32_fa7_xor1;
  assign f_u_dadda_cla32_fa349_and1 = f_u_dadda_cla32_fa349_xor0 & f_u_dadda_cla32_fa7_xor1;
  assign f_u_dadda_cla32_fa349_or0 = f_u_dadda_cla32_fa349_and0 | f_u_dadda_cla32_fa349_and1;
  assign f_u_dadda_cla32_fa350_xor0 = f_u_dadda_cla32_fa8_xor1 ^ f_u_dadda_cla32_ha4_xor0;
  assign f_u_dadda_cla32_fa350_and0 = f_u_dadda_cla32_fa8_xor1 & f_u_dadda_cla32_ha4_xor0;
  assign f_u_dadda_cla32_fa350_xor1 = f_u_dadda_cla32_fa350_xor0 ^ f_u_dadda_cla32_fa334_xor1;
  assign f_u_dadda_cla32_fa350_and1 = f_u_dadda_cla32_fa350_xor0 & f_u_dadda_cla32_fa334_xor1;
  assign f_u_dadda_cla32_fa350_or0 = f_u_dadda_cla32_fa350_and0 | f_u_dadda_cla32_fa350_and1;
  assign f_u_dadda_cla32_fa351_xor0 = f_u_dadda_cla32_fa335_xor1 ^ f_u_dadda_cla32_fa336_xor1;
  assign f_u_dadda_cla32_fa351_and0 = f_u_dadda_cla32_fa335_xor1 & f_u_dadda_cla32_fa336_xor1;
  assign f_u_dadda_cla32_fa351_xor1 = f_u_dadda_cla32_fa351_xor0 ^ f_u_dadda_cla32_fa337_xor1;
  assign f_u_dadda_cla32_fa351_and1 = f_u_dadda_cla32_fa351_xor0 & f_u_dadda_cla32_fa337_xor1;
  assign f_u_dadda_cla32_fa351_or0 = f_u_dadda_cla32_fa351_and0 | f_u_dadda_cla32_fa351_and1;
  assign f_u_dadda_cla32_fa352_xor0 = f_u_dadda_cla32_fa338_xor1 ^ f_u_dadda_cla32_fa339_xor1;
  assign f_u_dadda_cla32_fa352_and0 = f_u_dadda_cla32_fa338_xor1 & f_u_dadda_cla32_fa339_xor1;
  assign f_u_dadda_cla32_fa352_xor1 = f_u_dadda_cla32_fa352_xor0 ^ f_u_dadda_cla32_fa340_xor1;
  assign f_u_dadda_cla32_fa352_and1 = f_u_dadda_cla32_fa352_xor0 & f_u_dadda_cla32_fa340_xor1;
  assign f_u_dadda_cla32_fa352_or0 = f_u_dadda_cla32_fa352_and0 | f_u_dadda_cla32_fa352_and1;
  assign f_u_dadda_cla32_fa353_xor0 = f_u_dadda_cla32_fa341_xor1 ^ f_u_dadda_cla32_fa342_xor1;
  assign f_u_dadda_cla32_fa353_and0 = f_u_dadda_cla32_fa341_xor1 & f_u_dadda_cla32_fa342_xor1;
  assign f_u_dadda_cla32_fa353_xor1 = f_u_dadda_cla32_fa353_xor0 ^ f_u_dadda_cla32_fa343_xor1;
  assign f_u_dadda_cla32_fa353_and1 = f_u_dadda_cla32_fa353_xor0 & f_u_dadda_cla32_fa343_xor1;
  assign f_u_dadda_cla32_fa353_or0 = f_u_dadda_cla32_fa353_and0 | f_u_dadda_cla32_fa353_and1;
  assign f_u_dadda_cla32_fa354_xor0 = f_u_dadda_cla32_fa344_xor1 ^ f_u_dadda_cla32_fa345_xor1;
  assign f_u_dadda_cla32_fa354_and0 = f_u_dadda_cla32_fa344_xor1 & f_u_dadda_cla32_fa345_xor1;
  assign f_u_dadda_cla32_fa354_xor1 = f_u_dadda_cla32_fa354_xor0 ^ f_u_dadda_cla32_fa346_xor1;
  assign f_u_dadda_cla32_fa354_and1 = f_u_dadda_cla32_fa354_xor0 & f_u_dadda_cla32_fa346_xor1;
  assign f_u_dadda_cla32_fa354_or0 = f_u_dadda_cla32_fa354_and0 | f_u_dadda_cla32_fa354_and1;
  assign f_u_dadda_cla32_fa355_xor0 = f_u_dadda_cla32_fa347_xor1 ^ f_u_dadda_cla32_fa348_xor1;
  assign f_u_dadda_cla32_fa355_and0 = f_u_dadda_cla32_fa347_xor1 & f_u_dadda_cla32_fa348_xor1;
  assign f_u_dadda_cla32_fa355_xor1 = f_u_dadda_cla32_fa355_xor0 ^ f_u_dadda_cla32_fa349_xor1;
  assign f_u_dadda_cla32_fa355_and1 = f_u_dadda_cla32_fa355_xor0 & f_u_dadda_cla32_fa349_xor1;
  assign f_u_dadda_cla32_fa355_or0 = f_u_dadda_cla32_fa355_and0 | f_u_dadda_cla32_fa355_and1;
  assign f_u_dadda_cla32_fa356_xor0 = f_u_dadda_cla32_fa355_or0 ^ f_u_dadda_cla32_fa354_or0;
  assign f_u_dadda_cla32_fa356_and0 = f_u_dadda_cla32_fa355_or0 & f_u_dadda_cla32_fa354_or0;
  assign f_u_dadda_cla32_fa356_xor1 = f_u_dadda_cla32_fa356_xor0 ^ f_u_dadda_cla32_fa353_or0;
  assign f_u_dadda_cla32_fa356_and1 = f_u_dadda_cla32_fa356_xor0 & f_u_dadda_cla32_fa353_or0;
  assign f_u_dadda_cla32_fa356_or0 = f_u_dadda_cla32_fa356_and0 | f_u_dadda_cla32_fa356_and1;
  assign f_u_dadda_cla32_fa357_xor0 = f_u_dadda_cla32_fa352_or0 ^ f_u_dadda_cla32_fa351_or0;
  assign f_u_dadda_cla32_fa357_and0 = f_u_dadda_cla32_fa352_or0 & f_u_dadda_cla32_fa351_or0;
  assign f_u_dadda_cla32_fa357_xor1 = f_u_dadda_cla32_fa357_xor0 ^ f_u_dadda_cla32_fa350_or0;
  assign f_u_dadda_cla32_fa357_and1 = f_u_dadda_cla32_fa357_xor0 & f_u_dadda_cla32_fa350_or0;
  assign f_u_dadda_cla32_fa357_or0 = f_u_dadda_cla32_fa357_and0 | f_u_dadda_cla32_fa357_and1;
  assign f_u_dadda_cla32_fa358_xor0 = f_u_dadda_cla32_fa349_or0 ^ f_u_dadda_cla32_fa348_or0;
  assign f_u_dadda_cla32_fa358_and0 = f_u_dadda_cla32_fa349_or0 & f_u_dadda_cla32_fa348_or0;
  assign f_u_dadda_cla32_fa358_xor1 = f_u_dadda_cla32_fa358_xor0 ^ f_u_dadda_cla32_fa347_or0;
  assign f_u_dadda_cla32_fa358_and1 = f_u_dadda_cla32_fa358_xor0 & f_u_dadda_cla32_fa347_or0;
  assign f_u_dadda_cla32_fa358_or0 = f_u_dadda_cla32_fa358_and0 | f_u_dadda_cla32_fa358_and1;
  assign f_u_dadda_cla32_fa359_xor0 = f_u_dadda_cla32_fa346_or0 ^ f_u_dadda_cla32_fa345_or0;
  assign f_u_dadda_cla32_fa359_and0 = f_u_dadda_cla32_fa346_or0 & f_u_dadda_cla32_fa345_or0;
  assign f_u_dadda_cla32_fa359_xor1 = f_u_dadda_cla32_fa359_xor0 ^ f_u_dadda_cla32_fa344_or0;
  assign f_u_dadda_cla32_fa359_and1 = f_u_dadda_cla32_fa359_xor0 & f_u_dadda_cla32_fa344_or0;
  assign f_u_dadda_cla32_fa359_or0 = f_u_dadda_cla32_fa359_and0 | f_u_dadda_cla32_fa359_and1;
  assign f_u_dadda_cla32_fa360_xor0 = f_u_dadda_cla32_fa343_or0 ^ f_u_dadda_cla32_fa342_or0;
  assign f_u_dadda_cla32_fa360_and0 = f_u_dadda_cla32_fa343_or0 & f_u_dadda_cla32_fa342_or0;
  assign f_u_dadda_cla32_fa360_xor1 = f_u_dadda_cla32_fa360_xor0 ^ f_u_dadda_cla32_fa341_or0;
  assign f_u_dadda_cla32_fa360_and1 = f_u_dadda_cla32_fa360_xor0 & f_u_dadda_cla32_fa341_or0;
  assign f_u_dadda_cla32_fa360_or0 = f_u_dadda_cla32_fa360_and0 | f_u_dadda_cla32_fa360_and1;
  assign f_u_dadda_cla32_fa361_xor0 = f_u_dadda_cla32_fa340_or0 ^ f_u_dadda_cla32_fa339_or0;
  assign f_u_dadda_cla32_fa361_and0 = f_u_dadda_cla32_fa340_or0 & f_u_dadda_cla32_fa339_or0;
  assign f_u_dadda_cla32_fa361_xor1 = f_u_dadda_cla32_fa361_xor0 ^ f_u_dadda_cla32_fa338_or0;
  assign f_u_dadda_cla32_fa361_and1 = f_u_dadda_cla32_fa361_xor0 & f_u_dadda_cla32_fa338_or0;
  assign f_u_dadda_cla32_fa361_or0 = f_u_dadda_cla32_fa361_and0 | f_u_dadda_cla32_fa361_and1;
  assign f_u_dadda_cla32_fa362_xor0 = f_u_dadda_cla32_fa337_or0 ^ f_u_dadda_cla32_fa336_or0;
  assign f_u_dadda_cla32_fa362_and0 = f_u_dadda_cla32_fa337_or0 & f_u_dadda_cla32_fa336_or0;
  assign f_u_dadda_cla32_fa362_xor1 = f_u_dadda_cla32_fa362_xor0 ^ f_u_dadda_cla32_fa335_or0;
  assign f_u_dadda_cla32_fa362_and1 = f_u_dadda_cla32_fa362_xor0 & f_u_dadda_cla32_fa335_or0;
  assign f_u_dadda_cla32_fa362_or0 = f_u_dadda_cla32_fa362_and0 | f_u_dadda_cla32_fa362_and1;
  assign f_u_dadda_cla32_and_26_7 = a[26] & b[7];
  assign f_u_dadda_cla32_and_25_8 = a[25] & b[8];
  assign f_u_dadda_cla32_fa363_xor0 = f_u_dadda_cla32_fa334_or0 ^ f_u_dadda_cla32_and_26_7;
  assign f_u_dadda_cla32_fa363_and0 = f_u_dadda_cla32_fa334_or0 & f_u_dadda_cla32_and_26_7;
  assign f_u_dadda_cla32_fa363_xor1 = f_u_dadda_cla32_fa363_xor0 ^ f_u_dadda_cla32_and_25_8;
  assign f_u_dadda_cla32_fa363_and1 = f_u_dadda_cla32_fa363_xor0 & f_u_dadda_cla32_and_25_8;
  assign f_u_dadda_cla32_fa363_or0 = f_u_dadda_cla32_fa363_and0 | f_u_dadda_cla32_fa363_and1;
  assign f_u_dadda_cla32_and_24_9 = a[24] & b[9];
  assign f_u_dadda_cla32_and_23_10 = a[23] & b[10];
  assign f_u_dadda_cla32_and_22_11 = a[22] & b[11];
  assign f_u_dadda_cla32_fa364_xor0 = f_u_dadda_cla32_and_24_9 ^ f_u_dadda_cla32_and_23_10;
  assign f_u_dadda_cla32_fa364_and0 = f_u_dadda_cla32_and_24_9 & f_u_dadda_cla32_and_23_10;
  assign f_u_dadda_cla32_fa364_xor1 = f_u_dadda_cla32_fa364_xor0 ^ f_u_dadda_cla32_and_22_11;
  assign f_u_dadda_cla32_fa364_and1 = f_u_dadda_cla32_fa364_xor0 & f_u_dadda_cla32_and_22_11;
  assign f_u_dadda_cla32_fa364_or0 = f_u_dadda_cla32_fa364_and0 | f_u_dadda_cla32_fa364_and1;
  assign f_u_dadda_cla32_and_21_12 = a[21] & b[12];
  assign f_u_dadda_cla32_and_20_13 = a[20] & b[13];
  assign f_u_dadda_cla32_and_19_14 = a[19] & b[14];
  assign f_u_dadda_cla32_fa365_xor0 = f_u_dadda_cla32_and_21_12 ^ f_u_dadda_cla32_and_20_13;
  assign f_u_dadda_cla32_fa365_and0 = f_u_dadda_cla32_and_21_12 & f_u_dadda_cla32_and_20_13;
  assign f_u_dadda_cla32_fa365_xor1 = f_u_dadda_cla32_fa365_xor0 ^ f_u_dadda_cla32_and_19_14;
  assign f_u_dadda_cla32_fa365_and1 = f_u_dadda_cla32_fa365_xor0 & f_u_dadda_cla32_and_19_14;
  assign f_u_dadda_cla32_fa365_or0 = f_u_dadda_cla32_fa365_and0 | f_u_dadda_cla32_fa365_and1;
  assign f_u_dadda_cla32_and_18_15 = a[18] & b[15];
  assign f_u_dadda_cla32_and_17_16 = a[17] & b[16];
  assign f_u_dadda_cla32_and_16_17 = a[16] & b[17];
  assign f_u_dadda_cla32_fa366_xor0 = f_u_dadda_cla32_and_18_15 ^ f_u_dadda_cla32_and_17_16;
  assign f_u_dadda_cla32_fa366_and0 = f_u_dadda_cla32_and_18_15 & f_u_dadda_cla32_and_17_16;
  assign f_u_dadda_cla32_fa366_xor1 = f_u_dadda_cla32_fa366_xor0 ^ f_u_dadda_cla32_and_16_17;
  assign f_u_dadda_cla32_fa366_and1 = f_u_dadda_cla32_fa366_xor0 & f_u_dadda_cla32_and_16_17;
  assign f_u_dadda_cla32_fa366_or0 = f_u_dadda_cla32_fa366_and0 | f_u_dadda_cla32_fa366_and1;
  assign f_u_dadda_cla32_and_15_18 = a[15] & b[18];
  assign f_u_dadda_cla32_and_14_19 = a[14] & b[19];
  assign f_u_dadda_cla32_and_13_20 = a[13] & b[20];
  assign f_u_dadda_cla32_fa367_xor0 = f_u_dadda_cla32_and_15_18 ^ f_u_dadda_cla32_and_14_19;
  assign f_u_dadda_cla32_fa367_and0 = f_u_dadda_cla32_and_15_18 & f_u_dadda_cla32_and_14_19;
  assign f_u_dadda_cla32_fa367_xor1 = f_u_dadda_cla32_fa367_xor0 ^ f_u_dadda_cla32_and_13_20;
  assign f_u_dadda_cla32_fa367_and1 = f_u_dadda_cla32_fa367_xor0 & f_u_dadda_cla32_and_13_20;
  assign f_u_dadda_cla32_fa367_or0 = f_u_dadda_cla32_fa367_and0 | f_u_dadda_cla32_fa367_and1;
  assign f_u_dadda_cla32_and_12_21 = a[12] & b[21];
  assign f_u_dadda_cla32_and_11_22 = a[11] & b[22];
  assign f_u_dadda_cla32_and_10_23 = a[10] & b[23];
  assign f_u_dadda_cla32_fa368_xor0 = f_u_dadda_cla32_and_12_21 ^ f_u_dadda_cla32_and_11_22;
  assign f_u_dadda_cla32_fa368_and0 = f_u_dadda_cla32_and_12_21 & f_u_dadda_cla32_and_11_22;
  assign f_u_dadda_cla32_fa368_xor1 = f_u_dadda_cla32_fa368_xor0 ^ f_u_dadda_cla32_and_10_23;
  assign f_u_dadda_cla32_fa368_and1 = f_u_dadda_cla32_fa368_xor0 & f_u_dadda_cla32_and_10_23;
  assign f_u_dadda_cla32_fa368_or0 = f_u_dadda_cla32_fa368_and0 | f_u_dadda_cla32_fa368_and1;
  assign f_u_dadda_cla32_and_9_24 = a[9] & b[24];
  assign f_u_dadda_cla32_and_8_25 = a[8] & b[25];
  assign f_u_dadda_cla32_and_7_26 = a[7] & b[26];
  assign f_u_dadda_cla32_fa369_xor0 = f_u_dadda_cla32_and_9_24 ^ f_u_dadda_cla32_and_8_25;
  assign f_u_dadda_cla32_fa369_and0 = f_u_dadda_cla32_and_9_24 & f_u_dadda_cla32_and_8_25;
  assign f_u_dadda_cla32_fa369_xor1 = f_u_dadda_cla32_fa369_xor0 ^ f_u_dadda_cla32_and_7_26;
  assign f_u_dadda_cla32_fa369_and1 = f_u_dadda_cla32_fa369_xor0 & f_u_dadda_cla32_and_7_26;
  assign f_u_dadda_cla32_fa369_or0 = f_u_dadda_cla32_fa369_and0 | f_u_dadda_cla32_fa369_and1;
  assign f_u_dadda_cla32_and_6_27 = a[6] & b[27];
  assign f_u_dadda_cla32_and_5_28 = a[5] & b[28];
  assign f_u_dadda_cla32_and_4_29 = a[4] & b[29];
  assign f_u_dadda_cla32_fa370_xor0 = f_u_dadda_cla32_and_6_27 ^ f_u_dadda_cla32_and_5_28;
  assign f_u_dadda_cla32_fa370_and0 = f_u_dadda_cla32_and_6_27 & f_u_dadda_cla32_and_5_28;
  assign f_u_dadda_cla32_fa370_xor1 = f_u_dadda_cla32_fa370_xor0 ^ f_u_dadda_cla32_and_4_29;
  assign f_u_dadda_cla32_fa370_and1 = f_u_dadda_cla32_fa370_xor0 & f_u_dadda_cla32_and_4_29;
  assign f_u_dadda_cla32_fa370_or0 = f_u_dadda_cla32_fa370_and0 | f_u_dadda_cla32_fa370_and1;
  assign f_u_dadda_cla32_and_3_30 = a[3] & b[30];
  assign f_u_dadda_cla32_and_2_31 = a[2] & b[31];
  assign f_u_dadda_cla32_fa371_xor0 = f_u_dadda_cla32_and_3_30 ^ f_u_dadda_cla32_and_2_31;
  assign f_u_dadda_cla32_fa371_and0 = f_u_dadda_cla32_and_3_30 & f_u_dadda_cla32_and_2_31;
  assign f_u_dadda_cla32_fa371_xor1 = f_u_dadda_cla32_fa371_xor0 ^ f_u_dadda_cla32_fa9_xor1;
  assign f_u_dadda_cla32_fa371_and1 = f_u_dadda_cla32_fa371_xor0 & f_u_dadda_cla32_fa9_xor1;
  assign f_u_dadda_cla32_fa371_or0 = f_u_dadda_cla32_fa371_and0 | f_u_dadda_cla32_fa371_and1;
  assign f_u_dadda_cla32_fa372_xor0 = f_u_dadda_cla32_fa10_xor1 ^ f_u_dadda_cla32_fa11_xor1;
  assign f_u_dadda_cla32_fa372_and0 = f_u_dadda_cla32_fa10_xor1 & f_u_dadda_cla32_fa11_xor1;
  assign f_u_dadda_cla32_fa372_xor1 = f_u_dadda_cla32_fa372_xor0 ^ f_u_dadda_cla32_fa356_xor1;
  assign f_u_dadda_cla32_fa372_and1 = f_u_dadda_cla32_fa372_xor0 & f_u_dadda_cla32_fa356_xor1;
  assign f_u_dadda_cla32_fa372_or0 = f_u_dadda_cla32_fa372_and0 | f_u_dadda_cla32_fa372_and1;
  assign f_u_dadda_cla32_fa373_xor0 = f_u_dadda_cla32_fa357_xor1 ^ f_u_dadda_cla32_fa358_xor1;
  assign f_u_dadda_cla32_fa373_and0 = f_u_dadda_cla32_fa357_xor1 & f_u_dadda_cla32_fa358_xor1;
  assign f_u_dadda_cla32_fa373_xor1 = f_u_dadda_cla32_fa373_xor0 ^ f_u_dadda_cla32_fa359_xor1;
  assign f_u_dadda_cla32_fa373_and1 = f_u_dadda_cla32_fa373_xor0 & f_u_dadda_cla32_fa359_xor1;
  assign f_u_dadda_cla32_fa373_or0 = f_u_dadda_cla32_fa373_and0 | f_u_dadda_cla32_fa373_and1;
  assign f_u_dadda_cla32_fa374_xor0 = f_u_dadda_cla32_fa360_xor1 ^ f_u_dadda_cla32_fa361_xor1;
  assign f_u_dadda_cla32_fa374_and0 = f_u_dadda_cla32_fa360_xor1 & f_u_dadda_cla32_fa361_xor1;
  assign f_u_dadda_cla32_fa374_xor1 = f_u_dadda_cla32_fa374_xor0 ^ f_u_dadda_cla32_fa362_xor1;
  assign f_u_dadda_cla32_fa374_and1 = f_u_dadda_cla32_fa374_xor0 & f_u_dadda_cla32_fa362_xor1;
  assign f_u_dadda_cla32_fa374_or0 = f_u_dadda_cla32_fa374_and0 | f_u_dadda_cla32_fa374_and1;
  assign f_u_dadda_cla32_fa375_xor0 = f_u_dadda_cla32_fa363_xor1 ^ f_u_dadda_cla32_fa364_xor1;
  assign f_u_dadda_cla32_fa375_and0 = f_u_dadda_cla32_fa363_xor1 & f_u_dadda_cla32_fa364_xor1;
  assign f_u_dadda_cla32_fa375_xor1 = f_u_dadda_cla32_fa375_xor0 ^ f_u_dadda_cla32_fa365_xor1;
  assign f_u_dadda_cla32_fa375_and1 = f_u_dadda_cla32_fa375_xor0 & f_u_dadda_cla32_fa365_xor1;
  assign f_u_dadda_cla32_fa375_or0 = f_u_dadda_cla32_fa375_and0 | f_u_dadda_cla32_fa375_and1;
  assign f_u_dadda_cla32_fa376_xor0 = f_u_dadda_cla32_fa366_xor1 ^ f_u_dadda_cla32_fa367_xor1;
  assign f_u_dadda_cla32_fa376_and0 = f_u_dadda_cla32_fa366_xor1 & f_u_dadda_cla32_fa367_xor1;
  assign f_u_dadda_cla32_fa376_xor1 = f_u_dadda_cla32_fa376_xor0 ^ f_u_dadda_cla32_fa368_xor1;
  assign f_u_dadda_cla32_fa376_and1 = f_u_dadda_cla32_fa376_xor0 & f_u_dadda_cla32_fa368_xor1;
  assign f_u_dadda_cla32_fa376_or0 = f_u_dadda_cla32_fa376_and0 | f_u_dadda_cla32_fa376_and1;
  assign f_u_dadda_cla32_fa377_xor0 = f_u_dadda_cla32_fa369_xor1 ^ f_u_dadda_cla32_fa370_xor1;
  assign f_u_dadda_cla32_fa377_and0 = f_u_dadda_cla32_fa369_xor1 & f_u_dadda_cla32_fa370_xor1;
  assign f_u_dadda_cla32_fa377_xor1 = f_u_dadda_cla32_fa377_xor0 ^ f_u_dadda_cla32_fa371_xor1;
  assign f_u_dadda_cla32_fa377_and1 = f_u_dadda_cla32_fa377_xor0 & f_u_dadda_cla32_fa371_xor1;
  assign f_u_dadda_cla32_fa377_or0 = f_u_dadda_cla32_fa377_and0 | f_u_dadda_cla32_fa377_and1;
  assign f_u_dadda_cla32_fa378_xor0 = f_u_dadda_cla32_fa377_or0 ^ f_u_dadda_cla32_fa376_or0;
  assign f_u_dadda_cla32_fa378_and0 = f_u_dadda_cla32_fa377_or0 & f_u_dadda_cla32_fa376_or0;
  assign f_u_dadda_cla32_fa378_xor1 = f_u_dadda_cla32_fa378_xor0 ^ f_u_dadda_cla32_fa375_or0;
  assign f_u_dadda_cla32_fa378_and1 = f_u_dadda_cla32_fa378_xor0 & f_u_dadda_cla32_fa375_or0;
  assign f_u_dadda_cla32_fa378_or0 = f_u_dadda_cla32_fa378_and0 | f_u_dadda_cla32_fa378_and1;
  assign f_u_dadda_cla32_fa379_xor0 = f_u_dadda_cla32_fa374_or0 ^ f_u_dadda_cla32_fa373_or0;
  assign f_u_dadda_cla32_fa379_and0 = f_u_dadda_cla32_fa374_or0 & f_u_dadda_cla32_fa373_or0;
  assign f_u_dadda_cla32_fa379_xor1 = f_u_dadda_cla32_fa379_xor0 ^ f_u_dadda_cla32_fa372_or0;
  assign f_u_dadda_cla32_fa379_and1 = f_u_dadda_cla32_fa379_xor0 & f_u_dadda_cla32_fa372_or0;
  assign f_u_dadda_cla32_fa379_or0 = f_u_dadda_cla32_fa379_and0 | f_u_dadda_cla32_fa379_and1;
  assign f_u_dadda_cla32_fa380_xor0 = f_u_dadda_cla32_fa371_or0 ^ f_u_dadda_cla32_fa370_or0;
  assign f_u_dadda_cla32_fa380_and0 = f_u_dadda_cla32_fa371_or0 & f_u_dadda_cla32_fa370_or0;
  assign f_u_dadda_cla32_fa380_xor1 = f_u_dadda_cla32_fa380_xor0 ^ f_u_dadda_cla32_fa369_or0;
  assign f_u_dadda_cla32_fa380_and1 = f_u_dadda_cla32_fa380_xor0 & f_u_dadda_cla32_fa369_or0;
  assign f_u_dadda_cla32_fa380_or0 = f_u_dadda_cla32_fa380_and0 | f_u_dadda_cla32_fa380_and1;
  assign f_u_dadda_cla32_fa381_xor0 = f_u_dadda_cla32_fa368_or0 ^ f_u_dadda_cla32_fa367_or0;
  assign f_u_dadda_cla32_fa381_and0 = f_u_dadda_cla32_fa368_or0 & f_u_dadda_cla32_fa367_or0;
  assign f_u_dadda_cla32_fa381_xor1 = f_u_dadda_cla32_fa381_xor0 ^ f_u_dadda_cla32_fa366_or0;
  assign f_u_dadda_cla32_fa381_and1 = f_u_dadda_cla32_fa381_xor0 & f_u_dadda_cla32_fa366_or0;
  assign f_u_dadda_cla32_fa381_or0 = f_u_dadda_cla32_fa381_and0 | f_u_dadda_cla32_fa381_and1;
  assign f_u_dadda_cla32_fa382_xor0 = f_u_dadda_cla32_fa365_or0 ^ f_u_dadda_cla32_fa364_or0;
  assign f_u_dadda_cla32_fa382_and0 = f_u_dadda_cla32_fa365_or0 & f_u_dadda_cla32_fa364_or0;
  assign f_u_dadda_cla32_fa382_xor1 = f_u_dadda_cla32_fa382_xor0 ^ f_u_dadda_cla32_fa363_or0;
  assign f_u_dadda_cla32_fa382_and1 = f_u_dadda_cla32_fa382_xor0 & f_u_dadda_cla32_fa363_or0;
  assign f_u_dadda_cla32_fa382_or0 = f_u_dadda_cla32_fa382_and0 | f_u_dadda_cla32_fa382_and1;
  assign f_u_dadda_cla32_fa383_xor0 = f_u_dadda_cla32_fa362_or0 ^ f_u_dadda_cla32_fa361_or0;
  assign f_u_dadda_cla32_fa383_and0 = f_u_dadda_cla32_fa362_or0 & f_u_dadda_cla32_fa361_or0;
  assign f_u_dadda_cla32_fa383_xor1 = f_u_dadda_cla32_fa383_xor0 ^ f_u_dadda_cla32_fa360_or0;
  assign f_u_dadda_cla32_fa383_and1 = f_u_dadda_cla32_fa383_xor0 & f_u_dadda_cla32_fa360_or0;
  assign f_u_dadda_cla32_fa383_or0 = f_u_dadda_cla32_fa383_and0 | f_u_dadda_cla32_fa383_and1;
  assign f_u_dadda_cla32_fa384_xor0 = f_u_dadda_cla32_fa359_or0 ^ f_u_dadda_cla32_fa358_or0;
  assign f_u_dadda_cla32_fa384_and0 = f_u_dadda_cla32_fa359_or0 & f_u_dadda_cla32_fa358_or0;
  assign f_u_dadda_cla32_fa384_xor1 = f_u_dadda_cla32_fa384_xor0 ^ f_u_dadda_cla32_fa357_or0;
  assign f_u_dadda_cla32_fa384_and1 = f_u_dadda_cla32_fa384_xor0 & f_u_dadda_cla32_fa357_or0;
  assign f_u_dadda_cla32_fa384_or0 = f_u_dadda_cla32_fa384_and0 | f_u_dadda_cla32_fa384_and1;
  assign f_u_dadda_cla32_and_28_6 = a[28] & b[6];
  assign f_u_dadda_cla32_and_27_7 = a[27] & b[7];
  assign f_u_dadda_cla32_fa385_xor0 = f_u_dadda_cla32_fa356_or0 ^ f_u_dadda_cla32_and_28_6;
  assign f_u_dadda_cla32_fa385_and0 = f_u_dadda_cla32_fa356_or0 & f_u_dadda_cla32_and_28_6;
  assign f_u_dadda_cla32_fa385_xor1 = f_u_dadda_cla32_fa385_xor0 ^ f_u_dadda_cla32_and_27_7;
  assign f_u_dadda_cla32_fa385_and1 = f_u_dadda_cla32_fa385_xor0 & f_u_dadda_cla32_and_27_7;
  assign f_u_dadda_cla32_fa385_or0 = f_u_dadda_cla32_fa385_and0 | f_u_dadda_cla32_fa385_and1;
  assign f_u_dadda_cla32_and_26_8 = a[26] & b[8];
  assign f_u_dadda_cla32_and_25_9 = a[25] & b[9];
  assign f_u_dadda_cla32_and_24_10 = a[24] & b[10];
  assign f_u_dadda_cla32_fa386_xor0 = f_u_dadda_cla32_and_26_8 ^ f_u_dadda_cla32_and_25_9;
  assign f_u_dadda_cla32_fa386_and0 = f_u_dadda_cla32_and_26_8 & f_u_dadda_cla32_and_25_9;
  assign f_u_dadda_cla32_fa386_xor1 = f_u_dadda_cla32_fa386_xor0 ^ f_u_dadda_cla32_and_24_10;
  assign f_u_dadda_cla32_fa386_and1 = f_u_dadda_cla32_fa386_xor0 & f_u_dadda_cla32_and_24_10;
  assign f_u_dadda_cla32_fa386_or0 = f_u_dadda_cla32_fa386_and0 | f_u_dadda_cla32_fa386_and1;
  assign f_u_dadda_cla32_and_23_11 = a[23] & b[11];
  assign f_u_dadda_cla32_and_22_12 = a[22] & b[12];
  assign f_u_dadda_cla32_and_21_13 = a[21] & b[13];
  assign f_u_dadda_cla32_fa387_xor0 = f_u_dadda_cla32_and_23_11 ^ f_u_dadda_cla32_and_22_12;
  assign f_u_dadda_cla32_fa387_and0 = f_u_dadda_cla32_and_23_11 & f_u_dadda_cla32_and_22_12;
  assign f_u_dadda_cla32_fa387_xor1 = f_u_dadda_cla32_fa387_xor0 ^ f_u_dadda_cla32_and_21_13;
  assign f_u_dadda_cla32_fa387_and1 = f_u_dadda_cla32_fa387_xor0 & f_u_dadda_cla32_and_21_13;
  assign f_u_dadda_cla32_fa387_or0 = f_u_dadda_cla32_fa387_and0 | f_u_dadda_cla32_fa387_and1;
  assign f_u_dadda_cla32_and_20_14 = a[20] & b[14];
  assign f_u_dadda_cla32_and_19_15 = a[19] & b[15];
  assign f_u_dadda_cla32_and_18_16 = a[18] & b[16];
  assign f_u_dadda_cla32_fa388_xor0 = f_u_dadda_cla32_and_20_14 ^ f_u_dadda_cla32_and_19_15;
  assign f_u_dadda_cla32_fa388_and0 = f_u_dadda_cla32_and_20_14 & f_u_dadda_cla32_and_19_15;
  assign f_u_dadda_cla32_fa388_xor1 = f_u_dadda_cla32_fa388_xor0 ^ f_u_dadda_cla32_and_18_16;
  assign f_u_dadda_cla32_fa388_and1 = f_u_dadda_cla32_fa388_xor0 & f_u_dadda_cla32_and_18_16;
  assign f_u_dadda_cla32_fa388_or0 = f_u_dadda_cla32_fa388_and0 | f_u_dadda_cla32_fa388_and1;
  assign f_u_dadda_cla32_and_17_17 = a[17] & b[17];
  assign f_u_dadda_cla32_and_16_18 = a[16] & b[18];
  assign f_u_dadda_cla32_and_15_19 = a[15] & b[19];
  assign f_u_dadda_cla32_fa389_xor0 = f_u_dadda_cla32_and_17_17 ^ f_u_dadda_cla32_and_16_18;
  assign f_u_dadda_cla32_fa389_and0 = f_u_dadda_cla32_and_17_17 & f_u_dadda_cla32_and_16_18;
  assign f_u_dadda_cla32_fa389_xor1 = f_u_dadda_cla32_fa389_xor0 ^ f_u_dadda_cla32_and_15_19;
  assign f_u_dadda_cla32_fa389_and1 = f_u_dadda_cla32_fa389_xor0 & f_u_dadda_cla32_and_15_19;
  assign f_u_dadda_cla32_fa389_or0 = f_u_dadda_cla32_fa389_and0 | f_u_dadda_cla32_fa389_and1;
  assign f_u_dadda_cla32_and_14_20 = a[14] & b[20];
  assign f_u_dadda_cla32_and_13_21 = a[13] & b[21];
  assign f_u_dadda_cla32_and_12_22 = a[12] & b[22];
  assign f_u_dadda_cla32_fa390_xor0 = f_u_dadda_cla32_and_14_20 ^ f_u_dadda_cla32_and_13_21;
  assign f_u_dadda_cla32_fa390_and0 = f_u_dadda_cla32_and_14_20 & f_u_dadda_cla32_and_13_21;
  assign f_u_dadda_cla32_fa390_xor1 = f_u_dadda_cla32_fa390_xor0 ^ f_u_dadda_cla32_and_12_22;
  assign f_u_dadda_cla32_fa390_and1 = f_u_dadda_cla32_fa390_xor0 & f_u_dadda_cla32_and_12_22;
  assign f_u_dadda_cla32_fa390_or0 = f_u_dadda_cla32_fa390_and0 | f_u_dadda_cla32_fa390_and1;
  assign f_u_dadda_cla32_and_11_23 = a[11] & b[23];
  assign f_u_dadda_cla32_and_10_24 = a[10] & b[24];
  assign f_u_dadda_cla32_and_9_25 = a[9] & b[25];
  assign f_u_dadda_cla32_fa391_xor0 = f_u_dadda_cla32_and_11_23 ^ f_u_dadda_cla32_and_10_24;
  assign f_u_dadda_cla32_fa391_and0 = f_u_dadda_cla32_and_11_23 & f_u_dadda_cla32_and_10_24;
  assign f_u_dadda_cla32_fa391_xor1 = f_u_dadda_cla32_fa391_xor0 ^ f_u_dadda_cla32_and_9_25;
  assign f_u_dadda_cla32_fa391_and1 = f_u_dadda_cla32_fa391_xor0 & f_u_dadda_cla32_and_9_25;
  assign f_u_dadda_cla32_fa391_or0 = f_u_dadda_cla32_fa391_and0 | f_u_dadda_cla32_fa391_and1;
  assign f_u_dadda_cla32_and_8_26 = a[8] & b[26];
  assign f_u_dadda_cla32_and_7_27 = a[7] & b[27];
  assign f_u_dadda_cla32_and_6_28 = a[6] & b[28];
  assign f_u_dadda_cla32_fa392_xor0 = f_u_dadda_cla32_and_8_26 ^ f_u_dadda_cla32_and_7_27;
  assign f_u_dadda_cla32_fa392_and0 = f_u_dadda_cla32_and_8_26 & f_u_dadda_cla32_and_7_27;
  assign f_u_dadda_cla32_fa392_xor1 = f_u_dadda_cla32_fa392_xor0 ^ f_u_dadda_cla32_and_6_28;
  assign f_u_dadda_cla32_fa392_and1 = f_u_dadda_cla32_fa392_xor0 & f_u_dadda_cla32_and_6_28;
  assign f_u_dadda_cla32_fa392_or0 = f_u_dadda_cla32_fa392_and0 | f_u_dadda_cla32_fa392_and1;
  assign f_u_dadda_cla32_and_5_29 = a[5] & b[29];
  assign f_u_dadda_cla32_and_4_30 = a[4] & b[30];
  assign f_u_dadda_cla32_and_3_31 = a[3] & b[31];
  assign f_u_dadda_cla32_fa393_xor0 = f_u_dadda_cla32_and_5_29 ^ f_u_dadda_cla32_and_4_30;
  assign f_u_dadda_cla32_fa393_and0 = f_u_dadda_cla32_and_5_29 & f_u_dadda_cla32_and_4_30;
  assign f_u_dadda_cla32_fa393_xor1 = f_u_dadda_cla32_fa393_xor0 ^ f_u_dadda_cla32_and_3_31;
  assign f_u_dadda_cla32_fa393_and1 = f_u_dadda_cla32_fa393_xor0 & f_u_dadda_cla32_and_3_31;
  assign f_u_dadda_cla32_fa393_or0 = f_u_dadda_cla32_fa393_and0 | f_u_dadda_cla32_fa393_and1;
  assign f_u_dadda_cla32_fa394_xor0 = f_u_dadda_cla32_fa12_xor1 ^ f_u_dadda_cla32_fa13_xor1;
  assign f_u_dadda_cla32_fa394_and0 = f_u_dadda_cla32_fa12_xor1 & f_u_dadda_cla32_fa13_xor1;
  assign f_u_dadda_cla32_fa394_xor1 = f_u_dadda_cla32_fa394_xor0 ^ f_u_dadda_cla32_fa378_xor1;
  assign f_u_dadda_cla32_fa394_and1 = f_u_dadda_cla32_fa394_xor0 & f_u_dadda_cla32_fa378_xor1;
  assign f_u_dadda_cla32_fa394_or0 = f_u_dadda_cla32_fa394_and0 | f_u_dadda_cla32_fa394_and1;
  assign f_u_dadda_cla32_fa395_xor0 = f_u_dadda_cla32_fa379_xor1 ^ f_u_dadda_cla32_fa380_xor1;
  assign f_u_dadda_cla32_fa395_and0 = f_u_dadda_cla32_fa379_xor1 & f_u_dadda_cla32_fa380_xor1;
  assign f_u_dadda_cla32_fa395_xor1 = f_u_dadda_cla32_fa395_xor0 ^ f_u_dadda_cla32_fa381_xor1;
  assign f_u_dadda_cla32_fa395_and1 = f_u_dadda_cla32_fa395_xor0 & f_u_dadda_cla32_fa381_xor1;
  assign f_u_dadda_cla32_fa395_or0 = f_u_dadda_cla32_fa395_and0 | f_u_dadda_cla32_fa395_and1;
  assign f_u_dadda_cla32_fa396_xor0 = f_u_dadda_cla32_fa382_xor1 ^ f_u_dadda_cla32_fa383_xor1;
  assign f_u_dadda_cla32_fa396_and0 = f_u_dadda_cla32_fa382_xor1 & f_u_dadda_cla32_fa383_xor1;
  assign f_u_dadda_cla32_fa396_xor1 = f_u_dadda_cla32_fa396_xor0 ^ f_u_dadda_cla32_fa384_xor1;
  assign f_u_dadda_cla32_fa396_and1 = f_u_dadda_cla32_fa396_xor0 & f_u_dadda_cla32_fa384_xor1;
  assign f_u_dadda_cla32_fa396_or0 = f_u_dadda_cla32_fa396_and0 | f_u_dadda_cla32_fa396_and1;
  assign f_u_dadda_cla32_fa397_xor0 = f_u_dadda_cla32_fa385_xor1 ^ f_u_dadda_cla32_fa386_xor1;
  assign f_u_dadda_cla32_fa397_and0 = f_u_dadda_cla32_fa385_xor1 & f_u_dadda_cla32_fa386_xor1;
  assign f_u_dadda_cla32_fa397_xor1 = f_u_dadda_cla32_fa397_xor0 ^ f_u_dadda_cla32_fa387_xor1;
  assign f_u_dadda_cla32_fa397_and1 = f_u_dadda_cla32_fa397_xor0 & f_u_dadda_cla32_fa387_xor1;
  assign f_u_dadda_cla32_fa397_or0 = f_u_dadda_cla32_fa397_and0 | f_u_dadda_cla32_fa397_and1;
  assign f_u_dadda_cla32_fa398_xor0 = f_u_dadda_cla32_fa388_xor1 ^ f_u_dadda_cla32_fa389_xor1;
  assign f_u_dadda_cla32_fa398_and0 = f_u_dadda_cla32_fa388_xor1 & f_u_dadda_cla32_fa389_xor1;
  assign f_u_dadda_cla32_fa398_xor1 = f_u_dadda_cla32_fa398_xor0 ^ f_u_dadda_cla32_fa390_xor1;
  assign f_u_dadda_cla32_fa398_and1 = f_u_dadda_cla32_fa398_xor0 & f_u_dadda_cla32_fa390_xor1;
  assign f_u_dadda_cla32_fa398_or0 = f_u_dadda_cla32_fa398_and0 | f_u_dadda_cla32_fa398_and1;
  assign f_u_dadda_cla32_fa399_xor0 = f_u_dadda_cla32_fa391_xor1 ^ f_u_dadda_cla32_fa392_xor1;
  assign f_u_dadda_cla32_fa399_and0 = f_u_dadda_cla32_fa391_xor1 & f_u_dadda_cla32_fa392_xor1;
  assign f_u_dadda_cla32_fa399_xor1 = f_u_dadda_cla32_fa399_xor0 ^ f_u_dadda_cla32_fa393_xor1;
  assign f_u_dadda_cla32_fa399_and1 = f_u_dadda_cla32_fa399_xor0 & f_u_dadda_cla32_fa393_xor1;
  assign f_u_dadda_cla32_fa399_or0 = f_u_dadda_cla32_fa399_and0 | f_u_dadda_cla32_fa399_and1;
  assign f_u_dadda_cla32_fa400_xor0 = f_u_dadda_cla32_fa399_or0 ^ f_u_dadda_cla32_fa398_or0;
  assign f_u_dadda_cla32_fa400_and0 = f_u_dadda_cla32_fa399_or0 & f_u_dadda_cla32_fa398_or0;
  assign f_u_dadda_cla32_fa400_xor1 = f_u_dadda_cla32_fa400_xor0 ^ f_u_dadda_cla32_fa397_or0;
  assign f_u_dadda_cla32_fa400_and1 = f_u_dadda_cla32_fa400_xor0 & f_u_dadda_cla32_fa397_or0;
  assign f_u_dadda_cla32_fa400_or0 = f_u_dadda_cla32_fa400_and0 | f_u_dadda_cla32_fa400_and1;
  assign f_u_dadda_cla32_fa401_xor0 = f_u_dadda_cla32_fa396_or0 ^ f_u_dadda_cla32_fa395_or0;
  assign f_u_dadda_cla32_fa401_and0 = f_u_dadda_cla32_fa396_or0 & f_u_dadda_cla32_fa395_or0;
  assign f_u_dadda_cla32_fa401_xor1 = f_u_dadda_cla32_fa401_xor0 ^ f_u_dadda_cla32_fa394_or0;
  assign f_u_dadda_cla32_fa401_and1 = f_u_dadda_cla32_fa401_xor0 & f_u_dadda_cla32_fa394_or0;
  assign f_u_dadda_cla32_fa401_or0 = f_u_dadda_cla32_fa401_and0 | f_u_dadda_cla32_fa401_and1;
  assign f_u_dadda_cla32_fa402_xor0 = f_u_dadda_cla32_fa393_or0 ^ f_u_dadda_cla32_fa392_or0;
  assign f_u_dadda_cla32_fa402_and0 = f_u_dadda_cla32_fa393_or0 & f_u_dadda_cla32_fa392_or0;
  assign f_u_dadda_cla32_fa402_xor1 = f_u_dadda_cla32_fa402_xor0 ^ f_u_dadda_cla32_fa391_or0;
  assign f_u_dadda_cla32_fa402_and1 = f_u_dadda_cla32_fa402_xor0 & f_u_dadda_cla32_fa391_or0;
  assign f_u_dadda_cla32_fa402_or0 = f_u_dadda_cla32_fa402_and0 | f_u_dadda_cla32_fa402_and1;
  assign f_u_dadda_cla32_fa403_xor0 = f_u_dadda_cla32_fa390_or0 ^ f_u_dadda_cla32_fa389_or0;
  assign f_u_dadda_cla32_fa403_and0 = f_u_dadda_cla32_fa390_or0 & f_u_dadda_cla32_fa389_or0;
  assign f_u_dadda_cla32_fa403_xor1 = f_u_dadda_cla32_fa403_xor0 ^ f_u_dadda_cla32_fa388_or0;
  assign f_u_dadda_cla32_fa403_and1 = f_u_dadda_cla32_fa403_xor0 & f_u_dadda_cla32_fa388_or0;
  assign f_u_dadda_cla32_fa403_or0 = f_u_dadda_cla32_fa403_and0 | f_u_dadda_cla32_fa403_and1;
  assign f_u_dadda_cla32_fa404_xor0 = f_u_dadda_cla32_fa387_or0 ^ f_u_dadda_cla32_fa386_or0;
  assign f_u_dadda_cla32_fa404_and0 = f_u_dadda_cla32_fa387_or0 & f_u_dadda_cla32_fa386_or0;
  assign f_u_dadda_cla32_fa404_xor1 = f_u_dadda_cla32_fa404_xor0 ^ f_u_dadda_cla32_fa385_or0;
  assign f_u_dadda_cla32_fa404_and1 = f_u_dadda_cla32_fa404_xor0 & f_u_dadda_cla32_fa385_or0;
  assign f_u_dadda_cla32_fa404_or0 = f_u_dadda_cla32_fa404_and0 | f_u_dadda_cla32_fa404_and1;
  assign f_u_dadda_cla32_fa405_xor0 = f_u_dadda_cla32_fa384_or0 ^ f_u_dadda_cla32_fa383_or0;
  assign f_u_dadda_cla32_fa405_and0 = f_u_dadda_cla32_fa384_or0 & f_u_dadda_cla32_fa383_or0;
  assign f_u_dadda_cla32_fa405_xor1 = f_u_dadda_cla32_fa405_xor0 ^ f_u_dadda_cla32_fa382_or0;
  assign f_u_dadda_cla32_fa405_and1 = f_u_dadda_cla32_fa405_xor0 & f_u_dadda_cla32_fa382_or0;
  assign f_u_dadda_cla32_fa405_or0 = f_u_dadda_cla32_fa405_and0 | f_u_dadda_cla32_fa405_and1;
  assign f_u_dadda_cla32_fa406_xor0 = f_u_dadda_cla32_fa381_or0 ^ f_u_dadda_cla32_fa380_or0;
  assign f_u_dadda_cla32_fa406_and0 = f_u_dadda_cla32_fa381_or0 & f_u_dadda_cla32_fa380_or0;
  assign f_u_dadda_cla32_fa406_xor1 = f_u_dadda_cla32_fa406_xor0 ^ f_u_dadda_cla32_fa379_or0;
  assign f_u_dadda_cla32_fa406_and1 = f_u_dadda_cla32_fa406_xor0 & f_u_dadda_cla32_fa379_or0;
  assign f_u_dadda_cla32_fa406_or0 = f_u_dadda_cla32_fa406_and0 | f_u_dadda_cla32_fa406_and1;
  assign f_u_dadda_cla32_and_30_5 = a[30] & b[5];
  assign f_u_dadda_cla32_and_29_6 = a[29] & b[6];
  assign f_u_dadda_cla32_fa407_xor0 = f_u_dadda_cla32_fa378_or0 ^ f_u_dadda_cla32_and_30_5;
  assign f_u_dadda_cla32_fa407_and0 = f_u_dadda_cla32_fa378_or0 & f_u_dadda_cla32_and_30_5;
  assign f_u_dadda_cla32_fa407_xor1 = f_u_dadda_cla32_fa407_xor0 ^ f_u_dadda_cla32_and_29_6;
  assign f_u_dadda_cla32_fa407_and1 = f_u_dadda_cla32_fa407_xor0 & f_u_dadda_cla32_and_29_6;
  assign f_u_dadda_cla32_fa407_or0 = f_u_dadda_cla32_fa407_and0 | f_u_dadda_cla32_fa407_and1;
  assign f_u_dadda_cla32_and_28_7 = a[28] & b[7];
  assign f_u_dadda_cla32_and_27_8 = a[27] & b[8];
  assign f_u_dadda_cla32_and_26_9 = a[26] & b[9];
  assign f_u_dadda_cla32_fa408_xor0 = f_u_dadda_cla32_and_28_7 ^ f_u_dadda_cla32_and_27_8;
  assign f_u_dadda_cla32_fa408_and0 = f_u_dadda_cla32_and_28_7 & f_u_dadda_cla32_and_27_8;
  assign f_u_dadda_cla32_fa408_xor1 = f_u_dadda_cla32_fa408_xor0 ^ f_u_dadda_cla32_and_26_9;
  assign f_u_dadda_cla32_fa408_and1 = f_u_dadda_cla32_fa408_xor0 & f_u_dadda_cla32_and_26_9;
  assign f_u_dadda_cla32_fa408_or0 = f_u_dadda_cla32_fa408_and0 | f_u_dadda_cla32_fa408_and1;
  assign f_u_dadda_cla32_and_25_10 = a[25] & b[10];
  assign f_u_dadda_cla32_and_24_11 = a[24] & b[11];
  assign f_u_dadda_cla32_and_23_12 = a[23] & b[12];
  assign f_u_dadda_cla32_fa409_xor0 = f_u_dadda_cla32_and_25_10 ^ f_u_dadda_cla32_and_24_11;
  assign f_u_dadda_cla32_fa409_and0 = f_u_dadda_cla32_and_25_10 & f_u_dadda_cla32_and_24_11;
  assign f_u_dadda_cla32_fa409_xor1 = f_u_dadda_cla32_fa409_xor0 ^ f_u_dadda_cla32_and_23_12;
  assign f_u_dadda_cla32_fa409_and1 = f_u_dadda_cla32_fa409_xor0 & f_u_dadda_cla32_and_23_12;
  assign f_u_dadda_cla32_fa409_or0 = f_u_dadda_cla32_fa409_and0 | f_u_dadda_cla32_fa409_and1;
  assign f_u_dadda_cla32_and_22_13 = a[22] & b[13];
  assign f_u_dadda_cla32_and_21_14 = a[21] & b[14];
  assign f_u_dadda_cla32_and_20_15 = a[20] & b[15];
  assign f_u_dadda_cla32_fa410_xor0 = f_u_dadda_cla32_and_22_13 ^ f_u_dadda_cla32_and_21_14;
  assign f_u_dadda_cla32_fa410_and0 = f_u_dadda_cla32_and_22_13 & f_u_dadda_cla32_and_21_14;
  assign f_u_dadda_cla32_fa410_xor1 = f_u_dadda_cla32_fa410_xor0 ^ f_u_dadda_cla32_and_20_15;
  assign f_u_dadda_cla32_fa410_and1 = f_u_dadda_cla32_fa410_xor0 & f_u_dadda_cla32_and_20_15;
  assign f_u_dadda_cla32_fa410_or0 = f_u_dadda_cla32_fa410_and0 | f_u_dadda_cla32_fa410_and1;
  assign f_u_dadda_cla32_and_19_16 = a[19] & b[16];
  assign f_u_dadda_cla32_and_18_17 = a[18] & b[17];
  assign f_u_dadda_cla32_and_17_18 = a[17] & b[18];
  assign f_u_dadda_cla32_fa411_xor0 = f_u_dadda_cla32_and_19_16 ^ f_u_dadda_cla32_and_18_17;
  assign f_u_dadda_cla32_fa411_and0 = f_u_dadda_cla32_and_19_16 & f_u_dadda_cla32_and_18_17;
  assign f_u_dadda_cla32_fa411_xor1 = f_u_dadda_cla32_fa411_xor0 ^ f_u_dadda_cla32_and_17_18;
  assign f_u_dadda_cla32_fa411_and1 = f_u_dadda_cla32_fa411_xor0 & f_u_dadda_cla32_and_17_18;
  assign f_u_dadda_cla32_fa411_or0 = f_u_dadda_cla32_fa411_and0 | f_u_dadda_cla32_fa411_and1;
  assign f_u_dadda_cla32_and_16_19 = a[16] & b[19];
  assign f_u_dadda_cla32_and_15_20 = a[15] & b[20];
  assign f_u_dadda_cla32_and_14_21 = a[14] & b[21];
  assign f_u_dadda_cla32_fa412_xor0 = f_u_dadda_cla32_and_16_19 ^ f_u_dadda_cla32_and_15_20;
  assign f_u_dadda_cla32_fa412_and0 = f_u_dadda_cla32_and_16_19 & f_u_dadda_cla32_and_15_20;
  assign f_u_dadda_cla32_fa412_xor1 = f_u_dadda_cla32_fa412_xor0 ^ f_u_dadda_cla32_and_14_21;
  assign f_u_dadda_cla32_fa412_and1 = f_u_dadda_cla32_fa412_xor0 & f_u_dadda_cla32_and_14_21;
  assign f_u_dadda_cla32_fa412_or0 = f_u_dadda_cla32_fa412_and0 | f_u_dadda_cla32_fa412_and1;
  assign f_u_dadda_cla32_and_13_22 = a[13] & b[22];
  assign f_u_dadda_cla32_and_12_23 = a[12] & b[23];
  assign f_u_dadda_cla32_and_11_24 = a[11] & b[24];
  assign f_u_dadda_cla32_fa413_xor0 = f_u_dadda_cla32_and_13_22 ^ f_u_dadda_cla32_and_12_23;
  assign f_u_dadda_cla32_fa413_and0 = f_u_dadda_cla32_and_13_22 & f_u_dadda_cla32_and_12_23;
  assign f_u_dadda_cla32_fa413_xor1 = f_u_dadda_cla32_fa413_xor0 ^ f_u_dadda_cla32_and_11_24;
  assign f_u_dadda_cla32_fa413_and1 = f_u_dadda_cla32_fa413_xor0 & f_u_dadda_cla32_and_11_24;
  assign f_u_dadda_cla32_fa413_or0 = f_u_dadda_cla32_fa413_and0 | f_u_dadda_cla32_fa413_and1;
  assign f_u_dadda_cla32_and_10_25 = a[10] & b[25];
  assign f_u_dadda_cla32_and_9_26 = a[9] & b[26];
  assign f_u_dadda_cla32_and_8_27 = a[8] & b[27];
  assign f_u_dadda_cla32_fa414_xor0 = f_u_dadda_cla32_and_10_25 ^ f_u_dadda_cla32_and_9_26;
  assign f_u_dadda_cla32_fa414_and0 = f_u_dadda_cla32_and_10_25 & f_u_dadda_cla32_and_9_26;
  assign f_u_dadda_cla32_fa414_xor1 = f_u_dadda_cla32_fa414_xor0 ^ f_u_dadda_cla32_and_8_27;
  assign f_u_dadda_cla32_fa414_and1 = f_u_dadda_cla32_fa414_xor0 & f_u_dadda_cla32_and_8_27;
  assign f_u_dadda_cla32_fa414_or0 = f_u_dadda_cla32_fa414_and0 | f_u_dadda_cla32_fa414_and1;
  assign f_u_dadda_cla32_and_7_28 = a[7] & b[28];
  assign f_u_dadda_cla32_and_6_29 = a[6] & b[29];
  assign f_u_dadda_cla32_and_5_30 = a[5] & b[30];
  assign f_u_dadda_cla32_fa415_xor0 = f_u_dadda_cla32_and_7_28 ^ f_u_dadda_cla32_and_6_29;
  assign f_u_dadda_cla32_fa415_and0 = f_u_dadda_cla32_and_7_28 & f_u_dadda_cla32_and_6_29;
  assign f_u_dadda_cla32_fa415_xor1 = f_u_dadda_cla32_fa415_xor0 ^ f_u_dadda_cla32_and_5_30;
  assign f_u_dadda_cla32_fa415_and1 = f_u_dadda_cla32_fa415_xor0 & f_u_dadda_cla32_and_5_30;
  assign f_u_dadda_cla32_fa415_or0 = f_u_dadda_cla32_fa415_and0 | f_u_dadda_cla32_fa415_and1;
  assign f_u_dadda_cla32_and_4_31 = a[4] & b[31];
  assign f_u_dadda_cla32_fa416_xor0 = f_u_dadda_cla32_and_4_31 ^ f_u_dadda_cla32_fa14_xor1;
  assign f_u_dadda_cla32_fa416_and0 = f_u_dadda_cla32_and_4_31 & f_u_dadda_cla32_fa14_xor1;
  assign f_u_dadda_cla32_fa416_xor1 = f_u_dadda_cla32_fa416_xor0 ^ f_u_dadda_cla32_fa400_xor1;
  assign f_u_dadda_cla32_fa416_and1 = f_u_dadda_cla32_fa416_xor0 & f_u_dadda_cla32_fa400_xor1;
  assign f_u_dadda_cla32_fa416_or0 = f_u_dadda_cla32_fa416_and0 | f_u_dadda_cla32_fa416_and1;
  assign f_u_dadda_cla32_fa417_xor0 = f_u_dadda_cla32_fa401_xor1 ^ f_u_dadda_cla32_fa402_xor1;
  assign f_u_dadda_cla32_fa417_and0 = f_u_dadda_cla32_fa401_xor1 & f_u_dadda_cla32_fa402_xor1;
  assign f_u_dadda_cla32_fa417_xor1 = f_u_dadda_cla32_fa417_xor0 ^ f_u_dadda_cla32_fa403_xor1;
  assign f_u_dadda_cla32_fa417_and1 = f_u_dadda_cla32_fa417_xor0 & f_u_dadda_cla32_fa403_xor1;
  assign f_u_dadda_cla32_fa417_or0 = f_u_dadda_cla32_fa417_and0 | f_u_dadda_cla32_fa417_and1;
  assign f_u_dadda_cla32_fa418_xor0 = f_u_dadda_cla32_fa404_xor1 ^ f_u_dadda_cla32_fa405_xor1;
  assign f_u_dadda_cla32_fa418_and0 = f_u_dadda_cla32_fa404_xor1 & f_u_dadda_cla32_fa405_xor1;
  assign f_u_dadda_cla32_fa418_xor1 = f_u_dadda_cla32_fa418_xor0 ^ f_u_dadda_cla32_fa406_xor1;
  assign f_u_dadda_cla32_fa418_and1 = f_u_dadda_cla32_fa418_xor0 & f_u_dadda_cla32_fa406_xor1;
  assign f_u_dadda_cla32_fa418_or0 = f_u_dadda_cla32_fa418_and0 | f_u_dadda_cla32_fa418_and1;
  assign f_u_dadda_cla32_fa419_xor0 = f_u_dadda_cla32_fa407_xor1 ^ f_u_dadda_cla32_fa408_xor1;
  assign f_u_dadda_cla32_fa419_and0 = f_u_dadda_cla32_fa407_xor1 & f_u_dadda_cla32_fa408_xor1;
  assign f_u_dadda_cla32_fa419_xor1 = f_u_dadda_cla32_fa419_xor0 ^ f_u_dadda_cla32_fa409_xor1;
  assign f_u_dadda_cla32_fa419_and1 = f_u_dadda_cla32_fa419_xor0 & f_u_dadda_cla32_fa409_xor1;
  assign f_u_dadda_cla32_fa419_or0 = f_u_dadda_cla32_fa419_and0 | f_u_dadda_cla32_fa419_and1;
  assign f_u_dadda_cla32_fa420_xor0 = f_u_dadda_cla32_fa410_xor1 ^ f_u_dadda_cla32_fa411_xor1;
  assign f_u_dadda_cla32_fa420_and0 = f_u_dadda_cla32_fa410_xor1 & f_u_dadda_cla32_fa411_xor1;
  assign f_u_dadda_cla32_fa420_xor1 = f_u_dadda_cla32_fa420_xor0 ^ f_u_dadda_cla32_fa412_xor1;
  assign f_u_dadda_cla32_fa420_and1 = f_u_dadda_cla32_fa420_xor0 & f_u_dadda_cla32_fa412_xor1;
  assign f_u_dadda_cla32_fa420_or0 = f_u_dadda_cla32_fa420_and0 | f_u_dadda_cla32_fa420_and1;
  assign f_u_dadda_cla32_fa421_xor0 = f_u_dadda_cla32_fa413_xor1 ^ f_u_dadda_cla32_fa414_xor1;
  assign f_u_dadda_cla32_fa421_and0 = f_u_dadda_cla32_fa413_xor1 & f_u_dadda_cla32_fa414_xor1;
  assign f_u_dadda_cla32_fa421_xor1 = f_u_dadda_cla32_fa421_xor0 ^ f_u_dadda_cla32_fa415_xor1;
  assign f_u_dadda_cla32_fa421_and1 = f_u_dadda_cla32_fa421_xor0 & f_u_dadda_cla32_fa415_xor1;
  assign f_u_dadda_cla32_fa421_or0 = f_u_dadda_cla32_fa421_and0 | f_u_dadda_cla32_fa421_and1;
  assign f_u_dadda_cla32_fa422_xor0 = f_u_dadda_cla32_fa421_or0 ^ f_u_dadda_cla32_fa420_or0;
  assign f_u_dadda_cla32_fa422_and0 = f_u_dadda_cla32_fa421_or0 & f_u_dadda_cla32_fa420_or0;
  assign f_u_dadda_cla32_fa422_xor1 = f_u_dadda_cla32_fa422_xor0 ^ f_u_dadda_cla32_fa419_or0;
  assign f_u_dadda_cla32_fa422_and1 = f_u_dadda_cla32_fa422_xor0 & f_u_dadda_cla32_fa419_or0;
  assign f_u_dadda_cla32_fa422_or0 = f_u_dadda_cla32_fa422_and0 | f_u_dadda_cla32_fa422_and1;
  assign f_u_dadda_cla32_fa423_xor0 = f_u_dadda_cla32_fa418_or0 ^ f_u_dadda_cla32_fa417_or0;
  assign f_u_dadda_cla32_fa423_and0 = f_u_dadda_cla32_fa418_or0 & f_u_dadda_cla32_fa417_or0;
  assign f_u_dadda_cla32_fa423_xor1 = f_u_dadda_cla32_fa423_xor0 ^ f_u_dadda_cla32_fa416_or0;
  assign f_u_dadda_cla32_fa423_and1 = f_u_dadda_cla32_fa423_xor0 & f_u_dadda_cla32_fa416_or0;
  assign f_u_dadda_cla32_fa423_or0 = f_u_dadda_cla32_fa423_and0 | f_u_dadda_cla32_fa423_and1;
  assign f_u_dadda_cla32_fa424_xor0 = f_u_dadda_cla32_fa415_or0 ^ f_u_dadda_cla32_fa414_or0;
  assign f_u_dadda_cla32_fa424_and0 = f_u_dadda_cla32_fa415_or0 & f_u_dadda_cla32_fa414_or0;
  assign f_u_dadda_cla32_fa424_xor1 = f_u_dadda_cla32_fa424_xor0 ^ f_u_dadda_cla32_fa413_or0;
  assign f_u_dadda_cla32_fa424_and1 = f_u_dadda_cla32_fa424_xor0 & f_u_dadda_cla32_fa413_or0;
  assign f_u_dadda_cla32_fa424_or0 = f_u_dadda_cla32_fa424_and0 | f_u_dadda_cla32_fa424_and1;
  assign f_u_dadda_cla32_fa425_xor0 = f_u_dadda_cla32_fa412_or0 ^ f_u_dadda_cla32_fa411_or0;
  assign f_u_dadda_cla32_fa425_and0 = f_u_dadda_cla32_fa412_or0 & f_u_dadda_cla32_fa411_or0;
  assign f_u_dadda_cla32_fa425_xor1 = f_u_dadda_cla32_fa425_xor0 ^ f_u_dadda_cla32_fa410_or0;
  assign f_u_dadda_cla32_fa425_and1 = f_u_dadda_cla32_fa425_xor0 & f_u_dadda_cla32_fa410_or0;
  assign f_u_dadda_cla32_fa425_or0 = f_u_dadda_cla32_fa425_and0 | f_u_dadda_cla32_fa425_and1;
  assign f_u_dadda_cla32_fa426_xor0 = f_u_dadda_cla32_fa409_or0 ^ f_u_dadda_cla32_fa408_or0;
  assign f_u_dadda_cla32_fa426_and0 = f_u_dadda_cla32_fa409_or0 & f_u_dadda_cla32_fa408_or0;
  assign f_u_dadda_cla32_fa426_xor1 = f_u_dadda_cla32_fa426_xor0 ^ f_u_dadda_cla32_fa407_or0;
  assign f_u_dadda_cla32_fa426_and1 = f_u_dadda_cla32_fa426_xor0 & f_u_dadda_cla32_fa407_or0;
  assign f_u_dadda_cla32_fa426_or0 = f_u_dadda_cla32_fa426_and0 | f_u_dadda_cla32_fa426_and1;
  assign f_u_dadda_cla32_fa427_xor0 = f_u_dadda_cla32_fa406_or0 ^ f_u_dadda_cla32_fa405_or0;
  assign f_u_dadda_cla32_fa427_and0 = f_u_dadda_cla32_fa406_or0 & f_u_dadda_cla32_fa405_or0;
  assign f_u_dadda_cla32_fa427_xor1 = f_u_dadda_cla32_fa427_xor0 ^ f_u_dadda_cla32_fa404_or0;
  assign f_u_dadda_cla32_fa427_and1 = f_u_dadda_cla32_fa427_xor0 & f_u_dadda_cla32_fa404_or0;
  assign f_u_dadda_cla32_fa427_or0 = f_u_dadda_cla32_fa427_and0 | f_u_dadda_cla32_fa427_and1;
  assign f_u_dadda_cla32_fa428_xor0 = f_u_dadda_cla32_fa403_or0 ^ f_u_dadda_cla32_fa402_or0;
  assign f_u_dadda_cla32_fa428_and0 = f_u_dadda_cla32_fa403_or0 & f_u_dadda_cla32_fa402_or0;
  assign f_u_dadda_cla32_fa428_xor1 = f_u_dadda_cla32_fa428_xor0 ^ f_u_dadda_cla32_fa401_or0;
  assign f_u_dadda_cla32_fa428_and1 = f_u_dadda_cla32_fa428_xor0 & f_u_dadda_cla32_fa401_or0;
  assign f_u_dadda_cla32_fa428_or0 = f_u_dadda_cla32_fa428_and0 | f_u_dadda_cla32_fa428_and1;
  assign f_u_dadda_cla32_and_31_5 = a[31] & b[5];
  assign f_u_dadda_cla32_fa429_xor0 = f_u_dadda_cla32_fa400_or0 ^ f_u_dadda_cla32_fa14_or0;
  assign f_u_dadda_cla32_fa429_and0 = f_u_dadda_cla32_fa400_or0 & f_u_dadda_cla32_fa14_or0;
  assign f_u_dadda_cla32_fa429_xor1 = f_u_dadda_cla32_fa429_xor0 ^ f_u_dadda_cla32_and_31_5;
  assign f_u_dadda_cla32_fa429_and1 = f_u_dadda_cla32_fa429_xor0 & f_u_dadda_cla32_and_31_5;
  assign f_u_dadda_cla32_fa429_or0 = f_u_dadda_cla32_fa429_and0 | f_u_dadda_cla32_fa429_and1;
  assign f_u_dadda_cla32_and_30_6 = a[30] & b[6];
  assign f_u_dadda_cla32_and_29_7 = a[29] & b[7];
  assign f_u_dadda_cla32_and_28_8 = a[28] & b[8];
  assign f_u_dadda_cla32_fa430_xor0 = f_u_dadda_cla32_and_30_6 ^ f_u_dadda_cla32_and_29_7;
  assign f_u_dadda_cla32_fa430_and0 = f_u_dadda_cla32_and_30_6 & f_u_dadda_cla32_and_29_7;
  assign f_u_dadda_cla32_fa430_xor1 = f_u_dadda_cla32_fa430_xor0 ^ f_u_dadda_cla32_and_28_8;
  assign f_u_dadda_cla32_fa430_and1 = f_u_dadda_cla32_fa430_xor0 & f_u_dadda_cla32_and_28_8;
  assign f_u_dadda_cla32_fa430_or0 = f_u_dadda_cla32_fa430_and0 | f_u_dadda_cla32_fa430_and1;
  assign f_u_dadda_cla32_and_27_9 = a[27] & b[9];
  assign f_u_dadda_cla32_and_26_10 = a[26] & b[10];
  assign f_u_dadda_cla32_and_25_11 = a[25] & b[11];
  assign f_u_dadda_cla32_fa431_xor0 = f_u_dadda_cla32_and_27_9 ^ f_u_dadda_cla32_and_26_10;
  assign f_u_dadda_cla32_fa431_and0 = f_u_dadda_cla32_and_27_9 & f_u_dadda_cla32_and_26_10;
  assign f_u_dadda_cla32_fa431_xor1 = f_u_dadda_cla32_fa431_xor0 ^ f_u_dadda_cla32_and_25_11;
  assign f_u_dadda_cla32_fa431_and1 = f_u_dadda_cla32_fa431_xor0 & f_u_dadda_cla32_and_25_11;
  assign f_u_dadda_cla32_fa431_or0 = f_u_dadda_cla32_fa431_and0 | f_u_dadda_cla32_fa431_and1;
  assign f_u_dadda_cla32_and_24_12 = a[24] & b[12];
  assign f_u_dadda_cla32_and_23_13 = a[23] & b[13];
  assign f_u_dadda_cla32_and_22_14 = a[22] & b[14];
  assign f_u_dadda_cla32_fa432_xor0 = f_u_dadda_cla32_and_24_12 ^ f_u_dadda_cla32_and_23_13;
  assign f_u_dadda_cla32_fa432_and0 = f_u_dadda_cla32_and_24_12 & f_u_dadda_cla32_and_23_13;
  assign f_u_dadda_cla32_fa432_xor1 = f_u_dadda_cla32_fa432_xor0 ^ f_u_dadda_cla32_and_22_14;
  assign f_u_dadda_cla32_fa432_and1 = f_u_dadda_cla32_fa432_xor0 & f_u_dadda_cla32_and_22_14;
  assign f_u_dadda_cla32_fa432_or0 = f_u_dadda_cla32_fa432_and0 | f_u_dadda_cla32_fa432_and1;
  assign f_u_dadda_cla32_and_21_15 = a[21] & b[15];
  assign f_u_dadda_cla32_and_20_16 = a[20] & b[16];
  assign f_u_dadda_cla32_and_19_17 = a[19] & b[17];
  assign f_u_dadda_cla32_fa433_xor0 = f_u_dadda_cla32_and_21_15 ^ f_u_dadda_cla32_and_20_16;
  assign f_u_dadda_cla32_fa433_and0 = f_u_dadda_cla32_and_21_15 & f_u_dadda_cla32_and_20_16;
  assign f_u_dadda_cla32_fa433_xor1 = f_u_dadda_cla32_fa433_xor0 ^ f_u_dadda_cla32_and_19_17;
  assign f_u_dadda_cla32_fa433_and1 = f_u_dadda_cla32_fa433_xor0 & f_u_dadda_cla32_and_19_17;
  assign f_u_dadda_cla32_fa433_or0 = f_u_dadda_cla32_fa433_and0 | f_u_dadda_cla32_fa433_and1;
  assign f_u_dadda_cla32_and_18_18 = a[18] & b[18];
  assign f_u_dadda_cla32_and_17_19 = a[17] & b[19];
  assign f_u_dadda_cla32_and_16_20 = a[16] & b[20];
  assign f_u_dadda_cla32_fa434_xor0 = f_u_dadda_cla32_and_18_18 ^ f_u_dadda_cla32_and_17_19;
  assign f_u_dadda_cla32_fa434_and0 = f_u_dadda_cla32_and_18_18 & f_u_dadda_cla32_and_17_19;
  assign f_u_dadda_cla32_fa434_xor1 = f_u_dadda_cla32_fa434_xor0 ^ f_u_dadda_cla32_and_16_20;
  assign f_u_dadda_cla32_fa434_and1 = f_u_dadda_cla32_fa434_xor0 & f_u_dadda_cla32_and_16_20;
  assign f_u_dadda_cla32_fa434_or0 = f_u_dadda_cla32_fa434_and0 | f_u_dadda_cla32_fa434_and1;
  assign f_u_dadda_cla32_and_15_21 = a[15] & b[21];
  assign f_u_dadda_cla32_and_14_22 = a[14] & b[22];
  assign f_u_dadda_cla32_and_13_23 = a[13] & b[23];
  assign f_u_dadda_cla32_fa435_xor0 = f_u_dadda_cla32_and_15_21 ^ f_u_dadda_cla32_and_14_22;
  assign f_u_dadda_cla32_fa435_and0 = f_u_dadda_cla32_and_15_21 & f_u_dadda_cla32_and_14_22;
  assign f_u_dadda_cla32_fa435_xor1 = f_u_dadda_cla32_fa435_xor0 ^ f_u_dadda_cla32_and_13_23;
  assign f_u_dadda_cla32_fa435_and1 = f_u_dadda_cla32_fa435_xor0 & f_u_dadda_cla32_and_13_23;
  assign f_u_dadda_cla32_fa435_or0 = f_u_dadda_cla32_fa435_and0 | f_u_dadda_cla32_fa435_and1;
  assign f_u_dadda_cla32_and_12_24 = a[12] & b[24];
  assign f_u_dadda_cla32_and_11_25 = a[11] & b[25];
  assign f_u_dadda_cla32_and_10_26 = a[10] & b[26];
  assign f_u_dadda_cla32_fa436_xor0 = f_u_dadda_cla32_and_12_24 ^ f_u_dadda_cla32_and_11_25;
  assign f_u_dadda_cla32_fa436_and0 = f_u_dadda_cla32_and_12_24 & f_u_dadda_cla32_and_11_25;
  assign f_u_dadda_cla32_fa436_xor1 = f_u_dadda_cla32_fa436_xor0 ^ f_u_dadda_cla32_and_10_26;
  assign f_u_dadda_cla32_fa436_and1 = f_u_dadda_cla32_fa436_xor0 & f_u_dadda_cla32_and_10_26;
  assign f_u_dadda_cla32_fa436_or0 = f_u_dadda_cla32_fa436_and0 | f_u_dadda_cla32_fa436_and1;
  assign f_u_dadda_cla32_and_9_27 = a[9] & b[27];
  assign f_u_dadda_cla32_and_8_28 = a[8] & b[28];
  assign f_u_dadda_cla32_and_7_29 = a[7] & b[29];
  assign f_u_dadda_cla32_fa437_xor0 = f_u_dadda_cla32_and_9_27 ^ f_u_dadda_cla32_and_8_28;
  assign f_u_dadda_cla32_fa437_and0 = f_u_dadda_cla32_and_9_27 & f_u_dadda_cla32_and_8_28;
  assign f_u_dadda_cla32_fa437_xor1 = f_u_dadda_cla32_fa437_xor0 ^ f_u_dadda_cla32_and_7_29;
  assign f_u_dadda_cla32_fa437_and1 = f_u_dadda_cla32_fa437_xor0 & f_u_dadda_cla32_and_7_29;
  assign f_u_dadda_cla32_fa437_or0 = f_u_dadda_cla32_fa437_and0 | f_u_dadda_cla32_fa437_and1;
  assign f_u_dadda_cla32_and_6_30 = a[6] & b[30];
  assign f_u_dadda_cla32_and_5_31 = a[5] & b[31];
  assign f_u_dadda_cla32_fa438_xor0 = f_u_dadda_cla32_and_6_30 ^ f_u_dadda_cla32_and_5_31;
  assign f_u_dadda_cla32_fa438_and0 = f_u_dadda_cla32_and_6_30 & f_u_dadda_cla32_and_5_31;
  assign f_u_dadda_cla32_fa438_xor1 = f_u_dadda_cla32_fa438_xor0 ^ f_u_dadda_cla32_fa422_xor1;
  assign f_u_dadda_cla32_fa438_and1 = f_u_dadda_cla32_fa438_xor0 & f_u_dadda_cla32_fa422_xor1;
  assign f_u_dadda_cla32_fa438_or0 = f_u_dadda_cla32_fa438_and0 | f_u_dadda_cla32_fa438_and1;
  assign f_u_dadda_cla32_fa439_xor0 = f_u_dadda_cla32_fa423_xor1 ^ f_u_dadda_cla32_fa424_xor1;
  assign f_u_dadda_cla32_fa439_and0 = f_u_dadda_cla32_fa423_xor1 & f_u_dadda_cla32_fa424_xor1;
  assign f_u_dadda_cla32_fa439_xor1 = f_u_dadda_cla32_fa439_xor0 ^ f_u_dadda_cla32_fa425_xor1;
  assign f_u_dadda_cla32_fa439_and1 = f_u_dadda_cla32_fa439_xor0 & f_u_dadda_cla32_fa425_xor1;
  assign f_u_dadda_cla32_fa439_or0 = f_u_dadda_cla32_fa439_and0 | f_u_dadda_cla32_fa439_and1;
  assign f_u_dadda_cla32_fa440_xor0 = f_u_dadda_cla32_fa426_xor1 ^ f_u_dadda_cla32_fa427_xor1;
  assign f_u_dadda_cla32_fa440_and0 = f_u_dadda_cla32_fa426_xor1 & f_u_dadda_cla32_fa427_xor1;
  assign f_u_dadda_cla32_fa440_xor1 = f_u_dadda_cla32_fa440_xor0 ^ f_u_dadda_cla32_fa428_xor1;
  assign f_u_dadda_cla32_fa440_and1 = f_u_dadda_cla32_fa440_xor0 & f_u_dadda_cla32_fa428_xor1;
  assign f_u_dadda_cla32_fa440_or0 = f_u_dadda_cla32_fa440_and0 | f_u_dadda_cla32_fa440_and1;
  assign f_u_dadda_cla32_fa441_xor0 = f_u_dadda_cla32_fa429_xor1 ^ f_u_dadda_cla32_fa430_xor1;
  assign f_u_dadda_cla32_fa441_and0 = f_u_dadda_cla32_fa429_xor1 & f_u_dadda_cla32_fa430_xor1;
  assign f_u_dadda_cla32_fa441_xor1 = f_u_dadda_cla32_fa441_xor0 ^ f_u_dadda_cla32_fa431_xor1;
  assign f_u_dadda_cla32_fa441_and1 = f_u_dadda_cla32_fa441_xor0 & f_u_dadda_cla32_fa431_xor1;
  assign f_u_dadda_cla32_fa441_or0 = f_u_dadda_cla32_fa441_and0 | f_u_dadda_cla32_fa441_and1;
  assign f_u_dadda_cla32_fa442_xor0 = f_u_dadda_cla32_fa432_xor1 ^ f_u_dadda_cla32_fa433_xor1;
  assign f_u_dadda_cla32_fa442_and0 = f_u_dadda_cla32_fa432_xor1 & f_u_dadda_cla32_fa433_xor1;
  assign f_u_dadda_cla32_fa442_xor1 = f_u_dadda_cla32_fa442_xor0 ^ f_u_dadda_cla32_fa434_xor1;
  assign f_u_dadda_cla32_fa442_and1 = f_u_dadda_cla32_fa442_xor0 & f_u_dadda_cla32_fa434_xor1;
  assign f_u_dadda_cla32_fa442_or0 = f_u_dadda_cla32_fa442_and0 | f_u_dadda_cla32_fa442_and1;
  assign f_u_dadda_cla32_fa443_xor0 = f_u_dadda_cla32_fa435_xor1 ^ f_u_dadda_cla32_fa436_xor1;
  assign f_u_dadda_cla32_fa443_and0 = f_u_dadda_cla32_fa435_xor1 & f_u_dadda_cla32_fa436_xor1;
  assign f_u_dadda_cla32_fa443_xor1 = f_u_dadda_cla32_fa443_xor0 ^ f_u_dadda_cla32_fa437_xor1;
  assign f_u_dadda_cla32_fa443_and1 = f_u_dadda_cla32_fa443_xor0 & f_u_dadda_cla32_fa437_xor1;
  assign f_u_dadda_cla32_fa443_or0 = f_u_dadda_cla32_fa443_and0 | f_u_dadda_cla32_fa443_and1;
  assign f_u_dadda_cla32_fa444_xor0 = f_u_dadda_cla32_fa443_or0 ^ f_u_dadda_cla32_fa442_or0;
  assign f_u_dadda_cla32_fa444_and0 = f_u_dadda_cla32_fa443_or0 & f_u_dadda_cla32_fa442_or0;
  assign f_u_dadda_cla32_fa444_xor1 = f_u_dadda_cla32_fa444_xor0 ^ f_u_dadda_cla32_fa441_or0;
  assign f_u_dadda_cla32_fa444_and1 = f_u_dadda_cla32_fa444_xor0 & f_u_dadda_cla32_fa441_or0;
  assign f_u_dadda_cla32_fa444_or0 = f_u_dadda_cla32_fa444_and0 | f_u_dadda_cla32_fa444_and1;
  assign f_u_dadda_cla32_fa445_xor0 = f_u_dadda_cla32_fa440_or0 ^ f_u_dadda_cla32_fa439_or0;
  assign f_u_dadda_cla32_fa445_and0 = f_u_dadda_cla32_fa440_or0 & f_u_dadda_cla32_fa439_or0;
  assign f_u_dadda_cla32_fa445_xor1 = f_u_dadda_cla32_fa445_xor0 ^ f_u_dadda_cla32_fa438_or0;
  assign f_u_dadda_cla32_fa445_and1 = f_u_dadda_cla32_fa445_xor0 & f_u_dadda_cla32_fa438_or0;
  assign f_u_dadda_cla32_fa445_or0 = f_u_dadda_cla32_fa445_and0 | f_u_dadda_cla32_fa445_and1;
  assign f_u_dadda_cla32_fa446_xor0 = f_u_dadda_cla32_fa437_or0 ^ f_u_dadda_cla32_fa436_or0;
  assign f_u_dadda_cla32_fa446_and0 = f_u_dadda_cla32_fa437_or0 & f_u_dadda_cla32_fa436_or0;
  assign f_u_dadda_cla32_fa446_xor1 = f_u_dadda_cla32_fa446_xor0 ^ f_u_dadda_cla32_fa435_or0;
  assign f_u_dadda_cla32_fa446_and1 = f_u_dadda_cla32_fa446_xor0 & f_u_dadda_cla32_fa435_or0;
  assign f_u_dadda_cla32_fa446_or0 = f_u_dadda_cla32_fa446_and0 | f_u_dadda_cla32_fa446_and1;
  assign f_u_dadda_cla32_fa447_xor0 = f_u_dadda_cla32_fa434_or0 ^ f_u_dadda_cla32_fa433_or0;
  assign f_u_dadda_cla32_fa447_and0 = f_u_dadda_cla32_fa434_or0 & f_u_dadda_cla32_fa433_or0;
  assign f_u_dadda_cla32_fa447_xor1 = f_u_dadda_cla32_fa447_xor0 ^ f_u_dadda_cla32_fa432_or0;
  assign f_u_dadda_cla32_fa447_and1 = f_u_dadda_cla32_fa447_xor0 & f_u_dadda_cla32_fa432_or0;
  assign f_u_dadda_cla32_fa447_or0 = f_u_dadda_cla32_fa447_and0 | f_u_dadda_cla32_fa447_and1;
  assign f_u_dadda_cla32_fa448_xor0 = f_u_dadda_cla32_fa431_or0 ^ f_u_dadda_cla32_fa430_or0;
  assign f_u_dadda_cla32_fa448_and0 = f_u_dadda_cla32_fa431_or0 & f_u_dadda_cla32_fa430_or0;
  assign f_u_dadda_cla32_fa448_xor1 = f_u_dadda_cla32_fa448_xor0 ^ f_u_dadda_cla32_fa429_or0;
  assign f_u_dadda_cla32_fa448_and1 = f_u_dadda_cla32_fa448_xor0 & f_u_dadda_cla32_fa429_or0;
  assign f_u_dadda_cla32_fa448_or0 = f_u_dadda_cla32_fa448_and0 | f_u_dadda_cla32_fa448_and1;
  assign f_u_dadda_cla32_fa449_xor0 = f_u_dadda_cla32_fa428_or0 ^ f_u_dadda_cla32_fa427_or0;
  assign f_u_dadda_cla32_fa449_and0 = f_u_dadda_cla32_fa428_or0 & f_u_dadda_cla32_fa427_or0;
  assign f_u_dadda_cla32_fa449_xor1 = f_u_dadda_cla32_fa449_xor0 ^ f_u_dadda_cla32_fa426_or0;
  assign f_u_dadda_cla32_fa449_and1 = f_u_dadda_cla32_fa449_xor0 & f_u_dadda_cla32_fa426_or0;
  assign f_u_dadda_cla32_fa449_or0 = f_u_dadda_cla32_fa449_and0 | f_u_dadda_cla32_fa449_and1;
  assign f_u_dadda_cla32_fa450_xor0 = f_u_dadda_cla32_fa425_or0 ^ f_u_dadda_cla32_fa424_or0;
  assign f_u_dadda_cla32_fa450_and0 = f_u_dadda_cla32_fa425_or0 & f_u_dadda_cla32_fa424_or0;
  assign f_u_dadda_cla32_fa450_xor1 = f_u_dadda_cla32_fa450_xor0 ^ f_u_dadda_cla32_fa423_or0;
  assign f_u_dadda_cla32_fa450_and1 = f_u_dadda_cla32_fa450_xor0 & f_u_dadda_cla32_fa423_or0;
  assign f_u_dadda_cla32_fa450_or0 = f_u_dadda_cla32_fa450_and0 | f_u_dadda_cla32_fa450_and1;
  assign f_u_dadda_cla32_and_31_6 = a[31] & b[6];
  assign f_u_dadda_cla32_and_30_7 = a[30] & b[7];
  assign f_u_dadda_cla32_fa451_xor0 = f_u_dadda_cla32_fa422_or0 ^ f_u_dadda_cla32_and_31_6;
  assign f_u_dadda_cla32_fa451_and0 = f_u_dadda_cla32_fa422_or0 & f_u_dadda_cla32_and_31_6;
  assign f_u_dadda_cla32_fa451_xor1 = f_u_dadda_cla32_fa451_xor0 ^ f_u_dadda_cla32_and_30_7;
  assign f_u_dadda_cla32_fa451_and1 = f_u_dadda_cla32_fa451_xor0 & f_u_dadda_cla32_and_30_7;
  assign f_u_dadda_cla32_fa451_or0 = f_u_dadda_cla32_fa451_and0 | f_u_dadda_cla32_fa451_and1;
  assign f_u_dadda_cla32_and_29_8 = a[29] & b[8];
  assign f_u_dadda_cla32_and_28_9 = a[28] & b[9];
  assign f_u_dadda_cla32_and_27_10 = a[27] & b[10];
  assign f_u_dadda_cla32_fa452_xor0 = f_u_dadda_cla32_and_29_8 ^ f_u_dadda_cla32_and_28_9;
  assign f_u_dadda_cla32_fa452_and0 = f_u_dadda_cla32_and_29_8 & f_u_dadda_cla32_and_28_9;
  assign f_u_dadda_cla32_fa452_xor1 = f_u_dadda_cla32_fa452_xor0 ^ f_u_dadda_cla32_and_27_10;
  assign f_u_dadda_cla32_fa452_and1 = f_u_dadda_cla32_fa452_xor0 & f_u_dadda_cla32_and_27_10;
  assign f_u_dadda_cla32_fa452_or0 = f_u_dadda_cla32_fa452_and0 | f_u_dadda_cla32_fa452_and1;
  assign f_u_dadda_cla32_and_26_11 = a[26] & b[11];
  assign f_u_dadda_cla32_and_25_12 = a[25] & b[12];
  assign f_u_dadda_cla32_and_24_13 = a[24] & b[13];
  assign f_u_dadda_cla32_fa453_xor0 = f_u_dadda_cla32_and_26_11 ^ f_u_dadda_cla32_and_25_12;
  assign f_u_dadda_cla32_fa453_and0 = f_u_dadda_cla32_and_26_11 & f_u_dadda_cla32_and_25_12;
  assign f_u_dadda_cla32_fa453_xor1 = f_u_dadda_cla32_fa453_xor0 ^ f_u_dadda_cla32_and_24_13;
  assign f_u_dadda_cla32_fa453_and1 = f_u_dadda_cla32_fa453_xor0 & f_u_dadda_cla32_and_24_13;
  assign f_u_dadda_cla32_fa453_or0 = f_u_dadda_cla32_fa453_and0 | f_u_dadda_cla32_fa453_and1;
  assign f_u_dadda_cla32_and_23_14 = a[23] & b[14];
  assign f_u_dadda_cla32_and_22_15 = a[22] & b[15];
  assign f_u_dadda_cla32_and_21_16 = a[21] & b[16];
  assign f_u_dadda_cla32_fa454_xor0 = f_u_dadda_cla32_and_23_14 ^ f_u_dadda_cla32_and_22_15;
  assign f_u_dadda_cla32_fa454_and0 = f_u_dadda_cla32_and_23_14 & f_u_dadda_cla32_and_22_15;
  assign f_u_dadda_cla32_fa454_xor1 = f_u_dadda_cla32_fa454_xor0 ^ f_u_dadda_cla32_and_21_16;
  assign f_u_dadda_cla32_fa454_and1 = f_u_dadda_cla32_fa454_xor0 & f_u_dadda_cla32_and_21_16;
  assign f_u_dadda_cla32_fa454_or0 = f_u_dadda_cla32_fa454_and0 | f_u_dadda_cla32_fa454_and1;
  assign f_u_dadda_cla32_and_20_17 = a[20] & b[17];
  assign f_u_dadda_cla32_and_19_18 = a[19] & b[18];
  assign f_u_dadda_cla32_and_18_19 = a[18] & b[19];
  assign f_u_dadda_cla32_fa455_xor0 = f_u_dadda_cla32_and_20_17 ^ f_u_dadda_cla32_and_19_18;
  assign f_u_dadda_cla32_fa455_and0 = f_u_dadda_cla32_and_20_17 & f_u_dadda_cla32_and_19_18;
  assign f_u_dadda_cla32_fa455_xor1 = f_u_dadda_cla32_fa455_xor0 ^ f_u_dadda_cla32_and_18_19;
  assign f_u_dadda_cla32_fa455_and1 = f_u_dadda_cla32_fa455_xor0 & f_u_dadda_cla32_and_18_19;
  assign f_u_dadda_cla32_fa455_or0 = f_u_dadda_cla32_fa455_and0 | f_u_dadda_cla32_fa455_and1;
  assign f_u_dadda_cla32_and_17_20 = a[17] & b[20];
  assign f_u_dadda_cla32_and_16_21 = a[16] & b[21];
  assign f_u_dadda_cla32_and_15_22 = a[15] & b[22];
  assign f_u_dadda_cla32_fa456_xor0 = f_u_dadda_cla32_and_17_20 ^ f_u_dadda_cla32_and_16_21;
  assign f_u_dadda_cla32_fa456_and0 = f_u_dadda_cla32_and_17_20 & f_u_dadda_cla32_and_16_21;
  assign f_u_dadda_cla32_fa456_xor1 = f_u_dadda_cla32_fa456_xor0 ^ f_u_dadda_cla32_and_15_22;
  assign f_u_dadda_cla32_fa456_and1 = f_u_dadda_cla32_fa456_xor0 & f_u_dadda_cla32_and_15_22;
  assign f_u_dadda_cla32_fa456_or0 = f_u_dadda_cla32_fa456_and0 | f_u_dadda_cla32_fa456_and1;
  assign f_u_dadda_cla32_and_14_23 = a[14] & b[23];
  assign f_u_dadda_cla32_and_13_24 = a[13] & b[24];
  assign f_u_dadda_cla32_and_12_25 = a[12] & b[25];
  assign f_u_dadda_cla32_fa457_xor0 = f_u_dadda_cla32_and_14_23 ^ f_u_dadda_cla32_and_13_24;
  assign f_u_dadda_cla32_fa457_and0 = f_u_dadda_cla32_and_14_23 & f_u_dadda_cla32_and_13_24;
  assign f_u_dadda_cla32_fa457_xor1 = f_u_dadda_cla32_fa457_xor0 ^ f_u_dadda_cla32_and_12_25;
  assign f_u_dadda_cla32_fa457_and1 = f_u_dadda_cla32_fa457_xor0 & f_u_dadda_cla32_and_12_25;
  assign f_u_dadda_cla32_fa457_or0 = f_u_dadda_cla32_fa457_and0 | f_u_dadda_cla32_fa457_and1;
  assign f_u_dadda_cla32_and_11_26 = a[11] & b[26];
  assign f_u_dadda_cla32_and_10_27 = a[10] & b[27];
  assign f_u_dadda_cla32_and_9_28 = a[9] & b[28];
  assign f_u_dadda_cla32_fa458_xor0 = f_u_dadda_cla32_and_11_26 ^ f_u_dadda_cla32_and_10_27;
  assign f_u_dadda_cla32_fa458_and0 = f_u_dadda_cla32_and_11_26 & f_u_dadda_cla32_and_10_27;
  assign f_u_dadda_cla32_fa458_xor1 = f_u_dadda_cla32_fa458_xor0 ^ f_u_dadda_cla32_and_9_28;
  assign f_u_dadda_cla32_fa458_and1 = f_u_dadda_cla32_fa458_xor0 & f_u_dadda_cla32_and_9_28;
  assign f_u_dadda_cla32_fa458_or0 = f_u_dadda_cla32_fa458_and0 | f_u_dadda_cla32_fa458_and1;
  assign f_u_dadda_cla32_and_8_29 = a[8] & b[29];
  assign f_u_dadda_cla32_and_7_30 = a[7] & b[30];
  assign f_u_dadda_cla32_and_6_31 = a[6] & b[31];
  assign f_u_dadda_cla32_fa459_xor0 = f_u_dadda_cla32_and_8_29 ^ f_u_dadda_cla32_and_7_30;
  assign f_u_dadda_cla32_fa459_and0 = f_u_dadda_cla32_and_8_29 & f_u_dadda_cla32_and_7_30;
  assign f_u_dadda_cla32_fa459_xor1 = f_u_dadda_cla32_fa459_xor0 ^ f_u_dadda_cla32_and_6_31;
  assign f_u_dadda_cla32_fa459_and1 = f_u_dadda_cla32_fa459_xor0 & f_u_dadda_cla32_and_6_31;
  assign f_u_dadda_cla32_fa459_or0 = f_u_dadda_cla32_fa459_and0 | f_u_dadda_cla32_fa459_and1;
  assign f_u_dadda_cla32_fa460_xor0 = f_u_dadda_cla32_fa444_xor1 ^ f_u_dadda_cla32_fa445_xor1;
  assign f_u_dadda_cla32_fa460_and0 = f_u_dadda_cla32_fa444_xor1 & f_u_dadda_cla32_fa445_xor1;
  assign f_u_dadda_cla32_fa460_xor1 = f_u_dadda_cla32_fa460_xor0 ^ f_u_dadda_cla32_fa446_xor1;
  assign f_u_dadda_cla32_fa460_and1 = f_u_dadda_cla32_fa460_xor0 & f_u_dadda_cla32_fa446_xor1;
  assign f_u_dadda_cla32_fa460_or0 = f_u_dadda_cla32_fa460_and0 | f_u_dadda_cla32_fa460_and1;
  assign f_u_dadda_cla32_fa461_xor0 = f_u_dadda_cla32_fa447_xor1 ^ f_u_dadda_cla32_fa448_xor1;
  assign f_u_dadda_cla32_fa461_and0 = f_u_dadda_cla32_fa447_xor1 & f_u_dadda_cla32_fa448_xor1;
  assign f_u_dadda_cla32_fa461_xor1 = f_u_dadda_cla32_fa461_xor0 ^ f_u_dadda_cla32_fa449_xor1;
  assign f_u_dadda_cla32_fa461_and1 = f_u_dadda_cla32_fa461_xor0 & f_u_dadda_cla32_fa449_xor1;
  assign f_u_dadda_cla32_fa461_or0 = f_u_dadda_cla32_fa461_and0 | f_u_dadda_cla32_fa461_and1;
  assign f_u_dadda_cla32_fa462_xor0 = f_u_dadda_cla32_fa450_xor1 ^ f_u_dadda_cla32_fa451_xor1;
  assign f_u_dadda_cla32_fa462_and0 = f_u_dadda_cla32_fa450_xor1 & f_u_dadda_cla32_fa451_xor1;
  assign f_u_dadda_cla32_fa462_xor1 = f_u_dadda_cla32_fa462_xor0 ^ f_u_dadda_cla32_fa452_xor1;
  assign f_u_dadda_cla32_fa462_and1 = f_u_dadda_cla32_fa462_xor0 & f_u_dadda_cla32_fa452_xor1;
  assign f_u_dadda_cla32_fa462_or0 = f_u_dadda_cla32_fa462_and0 | f_u_dadda_cla32_fa462_and1;
  assign f_u_dadda_cla32_fa463_xor0 = f_u_dadda_cla32_fa453_xor1 ^ f_u_dadda_cla32_fa454_xor1;
  assign f_u_dadda_cla32_fa463_and0 = f_u_dadda_cla32_fa453_xor1 & f_u_dadda_cla32_fa454_xor1;
  assign f_u_dadda_cla32_fa463_xor1 = f_u_dadda_cla32_fa463_xor0 ^ f_u_dadda_cla32_fa455_xor1;
  assign f_u_dadda_cla32_fa463_and1 = f_u_dadda_cla32_fa463_xor0 & f_u_dadda_cla32_fa455_xor1;
  assign f_u_dadda_cla32_fa463_or0 = f_u_dadda_cla32_fa463_and0 | f_u_dadda_cla32_fa463_and1;
  assign f_u_dadda_cla32_fa464_xor0 = f_u_dadda_cla32_fa456_xor1 ^ f_u_dadda_cla32_fa457_xor1;
  assign f_u_dadda_cla32_fa464_and0 = f_u_dadda_cla32_fa456_xor1 & f_u_dadda_cla32_fa457_xor1;
  assign f_u_dadda_cla32_fa464_xor1 = f_u_dadda_cla32_fa464_xor0 ^ f_u_dadda_cla32_fa458_xor1;
  assign f_u_dadda_cla32_fa464_and1 = f_u_dadda_cla32_fa464_xor0 & f_u_dadda_cla32_fa458_xor1;
  assign f_u_dadda_cla32_fa464_or0 = f_u_dadda_cla32_fa464_and0 | f_u_dadda_cla32_fa464_and1;
  assign f_u_dadda_cla32_fa465_xor0 = f_u_dadda_cla32_fa464_or0 ^ f_u_dadda_cla32_fa463_or0;
  assign f_u_dadda_cla32_fa465_and0 = f_u_dadda_cla32_fa464_or0 & f_u_dadda_cla32_fa463_or0;
  assign f_u_dadda_cla32_fa465_xor1 = f_u_dadda_cla32_fa465_xor0 ^ f_u_dadda_cla32_fa462_or0;
  assign f_u_dadda_cla32_fa465_and1 = f_u_dadda_cla32_fa465_xor0 & f_u_dadda_cla32_fa462_or0;
  assign f_u_dadda_cla32_fa465_or0 = f_u_dadda_cla32_fa465_and0 | f_u_dadda_cla32_fa465_and1;
  assign f_u_dadda_cla32_fa466_xor0 = f_u_dadda_cla32_fa461_or0 ^ f_u_dadda_cla32_fa460_or0;
  assign f_u_dadda_cla32_fa466_and0 = f_u_dadda_cla32_fa461_or0 & f_u_dadda_cla32_fa460_or0;
  assign f_u_dadda_cla32_fa466_xor1 = f_u_dadda_cla32_fa466_xor0 ^ f_u_dadda_cla32_fa459_or0;
  assign f_u_dadda_cla32_fa466_and1 = f_u_dadda_cla32_fa466_xor0 & f_u_dadda_cla32_fa459_or0;
  assign f_u_dadda_cla32_fa466_or0 = f_u_dadda_cla32_fa466_and0 | f_u_dadda_cla32_fa466_and1;
  assign f_u_dadda_cla32_fa467_xor0 = f_u_dadda_cla32_fa458_or0 ^ f_u_dadda_cla32_fa457_or0;
  assign f_u_dadda_cla32_fa467_and0 = f_u_dadda_cla32_fa458_or0 & f_u_dadda_cla32_fa457_or0;
  assign f_u_dadda_cla32_fa467_xor1 = f_u_dadda_cla32_fa467_xor0 ^ f_u_dadda_cla32_fa456_or0;
  assign f_u_dadda_cla32_fa467_and1 = f_u_dadda_cla32_fa467_xor0 & f_u_dadda_cla32_fa456_or0;
  assign f_u_dadda_cla32_fa467_or0 = f_u_dadda_cla32_fa467_and0 | f_u_dadda_cla32_fa467_and1;
  assign f_u_dadda_cla32_fa468_xor0 = f_u_dadda_cla32_fa455_or0 ^ f_u_dadda_cla32_fa454_or0;
  assign f_u_dadda_cla32_fa468_and0 = f_u_dadda_cla32_fa455_or0 & f_u_dadda_cla32_fa454_or0;
  assign f_u_dadda_cla32_fa468_xor1 = f_u_dadda_cla32_fa468_xor0 ^ f_u_dadda_cla32_fa453_or0;
  assign f_u_dadda_cla32_fa468_and1 = f_u_dadda_cla32_fa468_xor0 & f_u_dadda_cla32_fa453_or0;
  assign f_u_dadda_cla32_fa468_or0 = f_u_dadda_cla32_fa468_and0 | f_u_dadda_cla32_fa468_and1;
  assign f_u_dadda_cla32_fa469_xor0 = f_u_dadda_cla32_fa452_or0 ^ f_u_dadda_cla32_fa451_or0;
  assign f_u_dadda_cla32_fa469_and0 = f_u_dadda_cla32_fa452_or0 & f_u_dadda_cla32_fa451_or0;
  assign f_u_dadda_cla32_fa469_xor1 = f_u_dadda_cla32_fa469_xor0 ^ f_u_dadda_cla32_fa450_or0;
  assign f_u_dadda_cla32_fa469_and1 = f_u_dadda_cla32_fa469_xor0 & f_u_dadda_cla32_fa450_or0;
  assign f_u_dadda_cla32_fa469_or0 = f_u_dadda_cla32_fa469_and0 | f_u_dadda_cla32_fa469_and1;
  assign f_u_dadda_cla32_fa470_xor0 = f_u_dadda_cla32_fa449_or0 ^ f_u_dadda_cla32_fa448_or0;
  assign f_u_dadda_cla32_fa470_and0 = f_u_dadda_cla32_fa449_or0 & f_u_dadda_cla32_fa448_or0;
  assign f_u_dadda_cla32_fa470_xor1 = f_u_dadda_cla32_fa470_xor0 ^ f_u_dadda_cla32_fa447_or0;
  assign f_u_dadda_cla32_fa470_and1 = f_u_dadda_cla32_fa470_xor0 & f_u_dadda_cla32_fa447_or0;
  assign f_u_dadda_cla32_fa470_or0 = f_u_dadda_cla32_fa470_and0 | f_u_dadda_cla32_fa470_and1;
  assign f_u_dadda_cla32_fa471_xor0 = f_u_dadda_cla32_fa446_or0 ^ f_u_dadda_cla32_fa445_or0;
  assign f_u_dadda_cla32_fa471_and0 = f_u_dadda_cla32_fa446_or0 & f_u_dadda_cla32_fa445_or0;
  assign f_u_dadda_cla32_fa471_xor1 = f_u_dadda_cla32_fa471_xor0 ^ f_u_dadda_cla32_fa444_or0;
  assign f_u_dadda_cla32_fa471_and1 = f_u_dadda_cla32_fa471_xor0 & f_u_dadda_cla32_fa444_or0;
  assign f_u_dadda_cla32_fa471_or0 = f_u_dadda_cla32_fa471_and0 | f_u_dadda_cla32_fa471_and1;
  assign f_u_dadda_cla32_and_31_7 = a[31] & b[7];
  assign f_u_dadda_cla32_and_30_8 = a[30] & b[8];
  assign f_u_dadda_cla32_and_29_9 = a[29] & b[9];
  assign f_u_dadda_cla32_fa472_xor0 = f_u_dadda_cla32_and_31_7 ^ f_u_dadda_cla32_and_30_8;
  assign f_u_dadda_cla32_fa472_and0 = f_u_dadda_cla32_and_31_7 & f_u_dadda_cla32_and_30_8;
  assign f_u_dadda_cla32_fa472_xor1 = f_u_dadda_cla32_fa472_xor0 ^ f_u_dadda_cla32_and_29_9;
  assign f_u_dadda_cla32_fa472_and1 = f_u_dadda_cla32_fa472_xor0 & f_u_dadda_cla32_and_29_9;
  assign f_u_dadda_cla32_fa472_or0 = f_u_dadda_cla32_fa472_and0 | f_u_dadda_cla32_fa472_and1;
  assign f_u_dadda_cla32_and_28_10 = a[28] & b[10];
  assign f_u_dadda_cla32_and_27_11 = a[27] & b[11];
  assign f_u_dadda_cla32_and_26_12 = a[26] & b[12];
  assign f_u_dadda_cla32_fa473_xor0 = f_u_dadda_cla32_and_28_10 ^ f_u_dadda_cla32_and_27_11;
  assign f_u_dadda_cla32_fa473_and0 = f_u_dadda_cla32_and_28_10 & f_u_dadda_cla32_and_27_11;
  assign f_u_dadda_cla32_fa473_xor1 = f_u_dadda_cla32_fa473_xor0 ^ f_u_dadda_cla32_and_26_12;
  assign f_u_dadda_cla32_fa473_and1 = f_u_dadda_cla32_fa473_xor0 & f_u_dadda_cla32_and_26_12;
  assign f_u_dadda_cla32_fa473_or0 = f_u_dadda_cla32_fa473_and0 | f_u_dadda_cla32_fa473_and1;
  assign f_u_dadda_cla32_and_25_13 = a[25] & b[13];
  assign f_u_dadda_cla32_and_24_14 = a[24] & b[14];
  assign f_u_dadda_cla32_and_23_15 = a[23] & b[15];
  assign f_u_dadda_cla32_fa474_xor0 = f_u_dadda_cla32_and_25_13 ^ f_u_dadda_cla32_and_24_14;
  assign f_u_dadda_cla32_fa474_and0 = f_u_dadda_cla32_and_25_13 & f_u_dadda_cla32_and_24_14;
  assign f_u_dadda_cla32_fa474_xor1 = f_u_dadda_cla32_fa474_xor0 ^ f_u_dadda_cla32_and_23_15;
  assign f_u_dadda_cla32_fa474_and1 = f_u_dadda_cla32_fa474_xor0 & f_u_dadda_cla32_and_23_15;
  assign f_u_dadda_cla32_fa474_or0 = f_u_dadda_cla32_fa474_and0 | f_u_dadda_cla32_fa474_and1;
  assign f_u_dadda_cla32_and_22_16 = a[22] & b[16];
  assign f_u_dadda_cla32_and_21_17 = a[21] & b[17];
  assign f_u_dadda_cla32_and_20_18 = a[20] & b[18];
  assign f_u_dadda_cla32_fa475_xor0 = f_u_dadda_cla32_and_22_16 ^ f_u_dadda_cla32_and_21_17;
  assign f_u_dadda_cla32_fa475_and0 = f_u_dadda_cla32_and_22_16 & f_u_dadda_cla32_and_21_17;
  assign f_u_dadda_cla32_fa475_xor1 = f_u_dadda_cla32_fa475_xor0 ^ f_u_dadda_cla32_and_20_18;
  assign f_u_dadda_cla32_fa475_and1 = f_u_dadda_cla32_fa475_xor0 & f_u_dadda_cla32_and_20_18;
  assign f_u_dadda_cla32_fa475_or0 = f_u_dadda_cla32_fa475_and0 | f_u_dadda_cla32_fa475_and1;
  assign f_u_dadda_cla32_and_19_19 = a[19] & b[19];
  assign f_u_dadda_cla32_and_18_20 = a[18] & b[20];
  assign f_u_dadda_cla32_and_17_21 = a[17] & b[21];
  assign f_u_dadda_cla32_fa476_xor0 = f_u_dadda_cla32_and_19_19 ^ f_u_dadda_cla32_and_18_20;
  assign f_u_dadda_cla32_fa476_and0 = f_u_dadda_cla32_and_19_19 & f_u_dadda_cla32_and_18_20;
  assign f_u_dadda_cla32_fa476_xor1 = f_u_dadda_cla32_fa476_xor0 ^ f_u_dadda_cla32_and_17_21;
  assign f_u_dadda_cla32_fa476_and1 = f_u_dadda_cla32_fa476_xor0 & f_u_dadda_cla32_and_17_21;
  assign f_u_dadda_cla32_fa476_or0 = f_u_dadda_cla32_fa476_and0 | f_u_dadda_cla32_fa476_and1;
  assign f_u_dadda_cla32_and_16_22 = a[16] & b[22];
  assign f_u_dadda_cla32_and_15_23 = a[15] & b[23];
  assign f_u_dadda_cla32_and_14_24 = a[14] & b[24];
  assign f_u_dadda_cla32_fa477_xor0 = f_u_dadda_cla32_and_16_22 ^ f_u_dadda_cla32_and_15_23;
  assign f_u_dadda_cla32_fa477_and0 = f_u_dadda_cla32_and_16_22 & f_u_dadda_cla32_and_15_23;
  assign f_u_dadda_cla32_fa477_xor1 = f_u_dadda_cla32_fa477_xor0 ^ f_u_dadda_cla32_and_14_24;
  assign f_u_dadda_cla32_fa477_and1 = f_u_dadda_cla32_fa477_xor0 & f_u_dadda_cla32_and_14_24;
  assign f_u_dadda_cla32_fa477_or0 = f_u_dadda_cla32_fa477_and0 | f_u_dadda_cla32_fa477_and1;
  assign f_u_dadda_cla32_and_13_25 = a[13] & b[25];
  assign f_u_dadda_cla32_and_12_26 = a[12] & b[26];
  assign f_u_dadda_cla32_and_11_27 = a[11] & b[27];
  assign f_u_dadda_cla32_fa478_xor0 = f_u_dadda_cla32_and_13_25 ^ f_u_dadda_cla32_and_12_26;
  assign f_u_dadda_cla32_fa478_and0 = f_u_dadda_cla32_and_13_25 & f_u_dadda_cla32_and_12_26;
  assign f_u_dadda_cla32_fa478_xor1 = f_u_dadda_cla32_fa478_xor0 ^ f_u_dadda_cla32_and_11_27;
  assign f_u_dadda_cla32_fa478_and1 = f_u_dadda_cla32_fa478_xor0 & f_u_dadda_cla32_and_11_27;
  assign f_u_dadda_cla32_fa478_or0 = f_u_dadda_cla32_fa478_and0 | f_u_dadda_cla32_fa478_and1;
  assign f_u_dadda_cla32_and_10_28 = a[10] & b[28];
  assign f_u_dadda_cla32_and_9_29 = a[9] & b[29];
  assign f_u_dadda_cla32_and_8_30 = a[8] & b[30];
  assign f_u_dadda_cla32_fa479_xor0 = f_u_dadda_cla32_and_10_28 ^ f_u_dadda_cla32_and_9_29;
  assign f_u_dadda_cla32_fa479_and0 = f_u_dadda_cla32_and_10_28 & f_u_dadda_cla32_and_9_29;
  assign f_u_dadda_cla32_fa479_xor1 = f_u_dadda_cla32_fa479_xor0 ^ f_u_dadda_cla32_and_8_30;
  assign f_u_dadda_cla32_fa479_and1 = f_u_dadda_cla32_fa479_xor0 & f_u_dadda_cla32_and_8_30;
  assign f_u_dadda_cla32_fa479_or0 = f_u_dadda_cla32_fa479_and0 | f_u_dadda_cla32_fa479_and1;
  assign f_u_dadda_cla32_and_7_31 = a[7] & b[31];
  assign f_u_dadda_cla32_fa480_xor0 = f_u_dadda_cla32_and_7_31 ^ f_u_dadda_cla32_fa465_xor1;
  assign f_u_dadda_cla32_fa480_and0 = f_u_dadda_cla32_and_7_31 & f_u_dadda_cla32_fa465_xor1;
  assign f_u_dadda_cla32_fa480_xor1 = f_u_dadda_cla32_fa480_xor0 ^ f_u_dadda_cla32_fa466_xor1;
  assign f_u_dadda_cla32_fa480_and1 = f_u_dadda_cla32_fa480_xor0 & f_u_dadda_cla32_fa466_xor1;
  assign f_u_dadda_cla32_fa480_or0 = f_u_dadda_cla32_fa480_and0 | f_u_dadda_cla32_fa480_and1;
  assign f_u_dadda_cla32_fa481_xor0 = f_u_dadda_cla32_fa467_xor1 ^ f_u_dadda_cla32_fa468_xor1;
  assign f_u_dadda_cla32_fa481_and0 = f_u_dadda_cla32_fa467_xor1 & f_u_dadda_cla32_fa468_xor1;
  assign f_u_dadda_cla32_fa481_xor1 = f_u_dadda_cla32_fa481_xor0 ^ f_u_dadda_cla32_fa469_xor1;
  assign f_u_dadda_cla32_fa481_and1 = f_u_dadda_cla32_fa481_xor0 & f_u_dadda_cla32_fa469_xor1;
  assign f_u_dadda_cla32_fa481_or0 = f_u_dadda_cla32_fa481_and0 | f_u_dadda_cla32_fa481_and1;
  assign f_u_dadda_cla32_fa482_xor0 = f_u_dadda_cla32_fa470_xor1 ^ f_u_dadda_cla32_fa471_xor1;
  assign f_u_dadda_cla32_fa482_and0 = f_u_dadda_cla32_fa470_xor1 & f_u_dadda_cla32_fa471_xor1;
  assign f_u_dadda_cla32_fa482_xor1 = f_u_dadda_cla32_fa482_xor0 ^ f_u_dadda_cla32_fa472_xor1;
  assign f_u_dadda_cla32_fa482_and1 = f_u_dadda_cla32_fa482_xor0 & f_u_dadda_cla32_fa472_xor1;
  assign f_u_dadda_cla32_fa482_or0 = f_u_dadda_cla32_fa482_and0 | f_u_dadda_cla32_fa482_and1;
  assign f_u_dadda_cla32_fa483_xor0 = f_u_dadda_cla32_fa473_xor1 ^ f_u_dadda_cla32_fa474_xor1;
  assign f_u_dadda_cla32_fa483_and0 = f_u_dadda_cla32_fa473_xor1 & f_u_dadda_cla32_fa474_xor1;
  assign f_u_dadda_cla32_fa483_xor1 = f_u_dadda_cla32_fa483_xor0 ^ f_u_dadda_cla32_fa475_xor1;
  assign f_u_dadda_cla32_fa483_and1 = f_u_dadda_cla32_fa483_xor0 & f_u_dadda_cla32_fa475_xor1;
  assign f_u_dadda_cla32_fa483_or0 = f_u_dadda_cla32_fa483_and0 | f_u_dadda_cla32_fa483_and1;
  assign f_u_dadda_cla32_fa484_xor0 = f_u_dadda_cla32_fa476_xor1 ^ f_u_dadda_cla32_fa477_xor1;
  assign f_u_dadda_cla32_fa484_and0 = f_u_dadda_cla32_fa476_xor1 & f_u_dadda_cla32_fa477_xor1;
  assign f_u_dadda_cla32_fa484_xor1 = f_u_dadda_cla32_fa484_xor0 ^ f_u_dadda_cla32_fa478_xor1;
  assign f_u_dadda_cla32_fa484_and1 = f_u_dadda_cla32_fa484_xor0 & f_u_dadda_cla32_fa478_xor1;
  assign f_u_dadda_cla32_fa484_or0 = f_u_dadda_cla32_fa484_and0 | f_u_dadda_cla32_fa484_and1;
  assign f_u_dadda_cla32_fa485_xor0 = f_u_dadda_cla32_fa484_or0 ^ f_u_dadda_cla32_fa483_or0;
  assign f_u_dadda_cla32_fa485_and0 = f_u_dadda_cla32_fa484_or0 & f_u_dadda_cla32_fa483_or0;
  assign f_u_dadda_cla32_fa485_xor1 = f_u_dadda_cla32_fa485_xor0 ^ f_u_dadda_cla32_fa482_or0;
  assign f_u_dadda_cla32_fa485_and1 = f_u_dadda_cla32_fa485_xor0 & f_u_dadda_cla32_fa482_or0;
  assign f_u_dadda_cla32_fa485_or0 = f_u_dadda_cla32_fa485_and0 | f_u_dadda_cla32_fa485_and1;
  assign f_u_dadda_cla32_fa486_xor0 = f_u_dadda_cla32_fa481_or0 ^ f_u_dadda_cla32_fa480_or0;
  assign f_u_dadda_cla32_fa486_and0 = f_u_dadda_cla32_fa481_or0 & f_u_dadda_cla32_fa480_or0;
  assign f_u_dadda_cla32_fa486_xor1 = f_u_dadda_cla32_fa486_xor0 ^ f_u_dadda_cla32_fa479_or0;
  assign f_u_dadda_cla32_fa486_and1 = f_u_dadda_cla32_fa486_xor0 & f_u_dadda_cla32_fa479_or0;
  assign f_u_dadda_cla32_fa486_or0 = f_u_dadda_cla32_fa486_and0 | f_u_dadda_cla32_fa486_and1;
  assign f_u_dadda_cla32_fa487_xor0 = f_u_dadda_cla32_fa478_or0 ^ f_u_dadda_cla32_fa477_or0;
  assign f_u_dadda_cla32_fa487_and0 = f_u_dadda_cla32_fa478_or0 & f_u_dadda_cla32_fa477_or0;
  assign f_u_dadda_cla32_fa487_xor1 = f_u_dadda_cla32_fa487_xor0 ^ f_u_dadda_cla32_fa476_or0;
  assign f_u_dadda_cla32_fa487_and1 = f_u_dadda_cla32_fa487_xor0 & f_u_dadda_cla32_fa476_or0;
  assign f_u_dadda_cla32_fa487_or0 = f_u_dadda_cla32_fa487_and0 | f_u_dadda_cla32_fa487_and1;
  assign f_u_dadda_cla32_fa488_xor0 = f_u_dadda_cla32_fa475_or0 ^ f_u_dadda_cla32_fa474_or0;
  assign f_u_dadda_cla32_fa488_and0 = f_u_dadda_cla32_fa475_or0 & f_u_dadda_cla32_fa474_or0;
  assign f_u_dadda_cla32_fa488_xor1 = f_u_dadda_cla32_fa488_xor0 ^ f_u_dadda_cla32_fa473_or0;
  assign f_u_dadda_cla32_fa488_and1 = f_u_dadda_cla32_fa488_xor0 & f_u_dadda_cla32_fa473_or0;
  assign f_u_dadda_cla32_fa488_or0 = f_u_dadda_cla32_fa488_and0 | f_u_dadda_cla32_fa488_and1;
  assign f_u_dadda_cla32_fa489_xor0 = f_u_dadda_cla32_fa472_or0 ^ f_u_dadda_cla32_fa471_or0;
  assign f_u_dadda_cla32_fa489_and0 = f_u_dadda_cla32_fa472_or0 & f_u_dadda_cla32_fa471_or0;
  assign f_u_dadda_cla32_fa489_xor1 = f_u_dadda_cla32_fa489_xor0 ^ f_u_dadda_cla32_fa470_or0;
  assign f_u_dadda_cla32_fa489_and1 = f_u_dadda_cla32_fa489_xor0 & f_u_dadda_cla32_fa470_or0;
  assign f_u_dadda_cla32_fa489_or0 = f_u_dadda_cla32_fa489_and0 | f_u_dadda_cla32_fa489_and1;
  assign f_u_dadda_cla32_fa490_xor0 = f_u_dadda_cla32_fa469_or0 ^ f_u_dadda_cla32_fa468_or0;
  assign f_u_dadda_cla32_fa490_and0 = f_u_dadda_cla32_fa469_or0 & f_u_dadda_cla32_fa468_or0;
  assign f_u_dadda_cla32_fa490_xor1 = f_u_dadda_cla32_fa490_xor0 ^ f_u_dadda_cla32_fa467_or0;
  assign f_u_dadda_cla32_fa490_and1 = f_u_dadda_cla32_fa490_xor0 & f_u_dadda_cla32_fa467_or0;
  assign f_u_dadda_cla32_fa490_or0 = f_u_dadda_cla32_fa490_and0 | f_u_dadda_cla32_fa490_and1;
  assign f_u_dadda_cla32_and_31_8 = a[31] & b[8];
  assign f_u_dadda_cla32_fa491_xor0 = f_u_dadda_cla32_fa466_or0 ^ f_u_dadda_cla32_fa465_or0;
  assign f_u_dadda_cla32_fa491_and0 = f_u_dadda_cla32_fa466_or0 & f_u_dadda_cla32_fa465_or0;
  assign f_u_dadda_cla32_fa491_xor1 = f_u_dadda_cla32_fa491_xor0 ^ f_u_dadda_cla32_and_31_8;
  assign f_u_dadda_cla32_fa491_and1 = f_u_dadda_cla32_fa491_xor0 & f_u_dadda_cla32_and_31_8;
  assign f_u_dadda_cla32_fa491_or0 = f_u_dadda_cla32_fa491_and0 | f_u_dadda_cla32_fa491_and1;
  assign f_u_dadda_cla32_and_30_9 = a[30] & b[9];
  assign f_u_dadda_cla32_and_29_10 = a[29] & b[10];
  assign f_u_dadda_cla32_and_28_11 = a[28] & b[11];
  assign f_u_dadda_cla32_fa492_xor0 = f_u_dadda_cla32_and_30_9 ^ f_u_dadda_cla32_and_29_10;
  assign f_u_dadda_cla32_fa492_and0 = f_u_dadda_cla32_and_30_9 & f_u_dadda_cla32_and_29_10;
  assign f_u_dadda_cla32_fa492_xor1 = f_u_dadda_cla32_fa492_xor0 ^ f_u_dadda_cla32_and_28_11;
  assign f_u_dadda_cla32_fa492_and1 = f_u_dadda_cla32_fa492_xor0 & f_u_dadda_cla32_and_28_11;
  assign f_u_dadda_cla32_fa492_or0 = f_u_dadda_cla32_fa492_and0 | f_u_dadda_cla32_fa492_and1;
  assign f_u_dadda_cla32_and_27_12 = a[27] & b[12];
  assign f_u_dadda_cla32_and_26_13 = a[26] & b[13];
  assign f_u_dadda_cla32_and_25_14 = a[25] & b[14];
  assign f_u_dadda_cla32_fa493_xor0 = f_u_dadda_cla32_and_27_12 ^ f_u_dadda_cla32_and_26_13;
  assign f_u_dadda_cla32_fa493_and0 = f_u_dadda_cla32_and_27_12 & f_u_dadda_cla32_and_26_13;
  assign f_u_dadda_cla32_fa493_xor1 = f_u_dadda_cla32_fa493_xor0 ^ f_u_dadda_cla32_and_25_14;
  assign f_u_dadda_cla32_fa493_and1 = f_u_dadda_cla32_fa493_xor0 & f_u_dadda_cla32_and_25_14;
  assign f_u_dadda_cla32_fa493_or0 = f_u_dadda_cla32_fa493_and0 | f_u_dadda_cla32_fa493_and1;
  assign f_u_dadda_cla32_and_24_15 = a[24] & b[15];
  assign f_u_dadda_cla32_and_23_16 = a[23] & b[16];
  assign f_u_dadda_cla32_and_22_17 = a[22] & b[17];
  assign f_u_dadda_cla32_fa494_xor0 = f_u_dadda_cla32_and_24_15 ^ f_u_dadda_cla32_and_23_16;
  assign f_u_dadda_cla32_fa494_and0 = f_u_dadda_cla32_and_24_15 & f_u_dadda_cla32_and_23_16;
  assign f_u_dadda_cla32_fa494_xor1 = f_u_dadda_cla32_fa494_xor0 ^ f_u_dadda_cla32_and_22_17;
  assign f_u_dadda_cla32_fa494_and1 = f_u_dadda_cla32_fa494_xor0 & f_u_dadda_cla32_and_22_17;
  assign f_u_dadda_cla32_fa494_or0 = f_u_dadda_cla32_fa494_and0 | f_u_dadda_cla32_fa494_and1;
  assign f_u_dadda_cla32_and_21_18 = a[21] & b[18];
  assign f_u_dadda_cla32_and_20_19 = a[20] & b[19];
  assign f_u_dadda_cla32_and_19_20 = a[19] & b[20];
  assign f_u_dadda_cla32_fa495_xor0 = f_u_dadda_cla32_and_21_18 ^ f_u_dadda_cla32_and_20_19;
  assign f_u_dadda_cla32_fa495_and0 = f_u_dadda_cla32_and_21_18 & f_u_dadda_cla32_and_20_19;
  assign f_u_dadda_cla32_fa495_xor1 = f_u_dadda_cla32_fa495_xor0 ^ f_u_dadda_cla32_and_19_20;
  assign f_u_dadda_cla32_fa495_and1 = f_u_dadda_cla32_fa495_xor0 & f_u_dadda_cla32_and_19_20;
  assign f_u_dadda_cla32_fa495_or0 = f_u_dadda_cla32_fa495_and0 | f_u_dadda_cla32_fa495_and1;
  assign f_u_dadda_cla32_and_18_21 = a[18] & b[21];
  assign f_u_dadda_cla32_and_17_22 = a[17] & b[22];
  assign f_u_dadda_cla32_and_16_23 = a[16] & b[23];
  assign f_u_dadda_cla32_fa496_xor0 = f_u_dadda_cla32_and_18_21 ^ f_u_dadda_cla32_and_17_22;
  assign f_u_dadda_cla32_fa496_and0 = f_u_dadda_cla32_and_18_21 & f_u_dadda_cla32_and_17_22;
  assign f_u_dadda_cla32_fa496_xor1 = f_u_dadda_cla32_fa496_xor0 ^ f_u_dadda_cla32_and_16_23;
  assign f_u_dadda_cla32_fa496_and1 = f_u_dadda_cla32_fa496_xor0 & f_u_dadda_cla32_and_16_23;
  assign f_u_dadda_cla32_fa496_or0 = f_u_dadda_cla32_fa496_and0 | f_u_dadda_cla32_fa496_and1;
  assign f_u_dadda_cla32_and_15_24 = a[15] & b[24];
  assign f_u_dadda_cla32_and_14_25 = a[14] & b[25];
  assign f_u_dadda_cla32_and_13_26 = a[13] & b[26];
  assign f_u_dadda_cla32_fa497_xor0 = f_u_dadda_cla32_and_15_24 ^ f_u_dadda_cla32_and_14_25;
  assign f_u_dadda_cla32_fa497_and0 = f_u_dadda_cla32_and_15_24 & f_u_dadda_cla32_and_14_25;
  assign f_u_dadda_cla32_fa497_xor1 = f_u_dadda_cla32_fa497_xor0 ^ f_u_dadda_cla32_and_13_26;
  assign f_u_dadda_cla32_fa497_and1 = f_u_dadda_cla32_fa497_xor0 & f_u_dadda_cla32_and_13_26;
  assign f_u_dadda_cla32_fa497_or0 = f_u_dadda_cla32_fa497_and0 | f_u_dadda_cla32_fa497_and1;
  assign f_u_dadda_cla32_and_12_27 = a[12] & b[27];
  assign f_u_dadda_cla32_and_11_28 = a[11] & b[28];
  assign f_u_dadda_cla32_and_10_29 = a[10] & b[29];
  assign f_u_dadda_cla32_fa498_xor0 = f_u_dadda_cla32_and_12_27 ^ f_u_dadda_cla32_and_11_28;
  assign f_u_dadda_cla32_fa498_and0 = f_u_dadda_cla32_and_12_27 & f_u_dadda_cla32_and_11_28;
  assign f_u_dadda_cla32_fa498_xor1 = f_u_dadda_cla32_fa498_xor0 ^ f_u_dadda_cla32_and_10_29;
  assign f_u_dadda_cla32_fa498_and1 = f_u_dadda_cla32_fa498_xor0 & f_u_dadda_cla32_and_10_29;
  assign f_u_dadda_cla32_fa498_or0 = f_u_dadda_cla32_fa498_and0 | f_u_dadda_cla32_fa498_and1;
  assign f_u_dadda_cla32_and_9_30 = a[9] & b[30];
  assign f_u_dadda_cla32_and_8_31 = a[8] & b[31];
  assign f_u_dadda_cla32_fa499_xor0 = f_u_dadda_cla32_and_9_30 ^ f_u_dadda_cla32_and_8_31;
  assign f_u_dadda_cla32_fa499_and0 = f_u_dadda_cla32_and_9_30 & f_u_dadda_cla32_and_8_31;
  assign f_u_dadda_cla32_fa499_xor1 = f_u_dadda_cla32_fa499_xor0 ^ f_u_dadda_cla32_fa485_xor1;
  assign f_u_dadda_cla32_fa499_and1 = f_u_dadda_cla32_fa499_xor0 & f_u_dadda_cla32_fa485_xor1;
  assign f_u_dadda_cla32_fa499_or0 = f_u_dadda_cla32_fa499_and0 | f_u_dadda_cla32_fa499_and1;
  assign f_u_dadda_cla32_fa500_xor0 = f_u_dadda_cla32_fa486_xor1 ^ f_u_dadda_cla32_fa487_xor1;
  assign f_u_dadda_cla32_fa500_and0 = f_u_dadda_cla32_fa486_xor1 & f_u_dadda_cla32_fa487_xor1;
  assign f_u_dadda_cla32_fa500_xor1 = f_u_dadda_cla32_fa500_xor0 ^ f_u_dadda_cla32_fa488_xor1;
  assign f_u_dadda_cla32_fa500_and1 = f_u_dadda_cla32_fa500_xor0 & f_u_dadda_cla32_fa488_xor1;
  assign f_u_dadda_cla32_fa500_or0 = f_u_dadda_cla32_fa500_and0 | f_u_dadda_cla32_fa500_and1;
  assign f_u_dadda_cla32_fa501_xor0 = f_u_dadda_cla32_fa489_xor1 ^ f_u_dadda_cla32_fa490_xor1;
  assign f_u_dadda_cla32_fa501_and0 = f_u_dadda_cla32_fa489_xor1 & f_u_dadda_cla32_fa490_xor1;
  assign f_u_dadda_cla32_fa501_xor1 = f_u_dadda_cla32_fa501_xor0 ^ f_u_dadda_cla32_fa491_xor1;
  assign f_u_dadda_cla32_fa501_and1 = f_u_dadda_cla32_fa501_xor0 & f_u_dadda_cla32_fa491_xor1;
  assign f_u_dadda_cla32_fa501_or0 = f_u_dadda_cla32_fa501_and0 | f_u_dadda_cla32_fa501_and1;
  assign f_u_dadda_cla32_fa502_xor0 = f_u_dadda_cla32_fa492_xor1 ^ f_u_dadda_cla32_fa493_xor1;
  assign f_u_dadda_cla32_fa502_and0 = f_u_dadda_cla32_fa492_xor1 & f_u_dadda_cla32_fa493_xor1;
  assign f_u_dadda_cla32_fa502_xor1 = f_u_dadda_cla32_fa502_xor0 ^ f_u_dadda_cla32_fa494_xor1;
  assign f_u_dadda_cla32_fa502_and1 = f_u_dadda_cla32_fa502_xor0 & f_u_dadda_cla32_fa494_xor1;
  assign f_u_dadda_cla32_fa502_or0 = f_u_dadda_cla32_fa502_and0 | f_u_dadda_cla32_fa502_and1;
  assign f_u_dadda_cla32_fa503_xor0 = f_u_dadda_cla32_fa495_xor1 ^ f_u_dadda_cla32_fa496_xor1;
  assign f_u_dadda_cla32_fa503_and0 = f_u_dadda_cla32_fa495_xor1 & f_u_dadda_cla32_fa496_xor1;
  assign f_u_dadda_cla32_fa503_xor1 = f_u_dadda_cla32_fa503_xor0 ^ f_u_dadda_cla32_fa497_xor1;
  assign f_u_dadda_cla32_fa503_and1 = f_u_dadda_cla32_fa503_xor0 & f_u_dadda_cla32_fa497_xor1;
  assign f_u_dadda_cla32_fa503_or0 = f_u_dadda_cla32_fa503_and0 | f_u_dadda_cla32_fa503_and1;
  assign f_u_dadda_cla32_fa504_xor0 = f_u_dadda_cla32_fa503_or0 ^ f_u_dadda_cla32_fa502_or0;
  assign f_u_dadda_cla32_fa504_and0 = f_u_dadda_cla32_fa503_or0 & f_u_dadda_cla32_fa502_or0;
  assign f_u_dadda_cla32_fa504_xor1 = f_u_dadda_cla32_fa504_xor0 ^ f_u_dadda_cla32_fa501_or0;
  assign f_u_dadda_cla32_fa504_and1 = f_u_dadda_cla32_fa504_xor0 & f_u_dadda_cla32_fa501_or0;
  assign f_u_dadda_cla32_fa504_or0 = f_u_dadda_cla32_fa504_and0 | f_u_dadda_cla32_fa504_and1;
  assign f_u_dadda_cla32_fa505_xor0 = f_u_dadda_cla32_fa500_or0 ^ f_u_dadda_cla32_fa499_or0;
  assign f_u_dadda_cla32_fa505_and0 = f_u_dadda_cla32_fa500_or0 & f_u_dadda_cla32_fa499_or0;
  assign f_u_dadda_cla32_fa505_xor1 = f_u_dadda_cla32_fa505_xor0 ^ f_u_dadda_cla32_fa498_or0;
  assign f_u_dadda_cla32_fa505_and1 = f_u_dadda_cla32_fa505_xor0 & f_u_dadda_cla32_fa498_or0;
  assign f_u_dadda_cla32_fa505_or0 = f_u_dadda_cla32_fa505_and0 | f_u_dadda_cla32_fa505_and1;
  assign f_u_dadda_cla32_fa506_xor0 = f_u_dadda_cla32_fa497_or0 ^ f_u_dadda_cla32_fa496_or0;
  assign f_u_dadda_cla32_fa506_and0 = f_u_dadda_cla32_fa497_or0 & f_u_dadda_cla32_fa496_or0;
  assign f_u_dadda_cla32_fa506_xor1 = f_u_dadda_cla32_fa506_xor0 ^ f_u_dadda_cla32_fa495_or0;
  assign f_u_dadda_cla32_fa506_and1 = f_u_dadda_cla32_fa506_xor0 & f_u_dadda_cla32_fa495_or0;
  assign f_u_dadda_cla32_fa506_or0 = f_u_dadda_cla32_fa506_and0 | f_u_dadda_cla32_fa506_and1;
  assign f_u_dadda_cla32_fa507_xor0 = f_u_dadda_cla32_fa494_or0 ^ f_u_dadda_cla32_fa493_or0;
  assign f_u_dadda_cla32_fa507_and0 = f_u_dadda_cla32_fa494_or0 & f_u_dadda_cla32_fa493_or0;
  assign f_u_dadda_cla32_fa507_xor1 = f_u_dadda_cla32_fa507_xor0 ^ f_u_dadda_cla32_fa492_or0;
  assign f_u_dadda_cla32_fa507_and1 = f_u_dadda_cla32_fa507_xor0 & f_u_dadda_cla32_fa492_or0;
  assign f_u_dadda_cla32_fa507_or0 = f_u_dadda_cla32_fa507_and0 | f_u_dadda_cla32_fa507_and1;
  assign f_u_dadda_cla32_fa508_xor0 = f_u_dadda_cla32_fa491_or0 ^ f_u_dadda_cla32_fa490_or0;
  assign f_u_dadda_cla32_fa508_and0 = f_u_dadda_cla32_fa491_or0 & f_u_dadda_cla32_fa490_or0;
  assign f_u_dadda_cla32_fa508_xor1 = f_u_dadda_cla32_fa508_xor0 ^ f_u_dadda_cla32_fa489_or0;
  assign f_u_dadda_cla32_fa508_and1 = f_u_dadda_cla32_fa508_xor0 & f_u_dadda_cla32_fa489_or0;
  assign f_u_dadda_cla32_fa508_or0 = f_u_dadda_cla32_fa508_and0 | f_u_dadda_cla32_fa508_and1;
  assign f_u_dadda_cla32_fa509_xor0 = f_u_dadda_cla32_fa488_or0 ^ f_u_dadda_cla32_fa487_or0;
  assign f_u_dadda_cla32_fa509_and0 = f_u_dadda_cla32_fa488_or0 & f_u_dadda_cla32_fa487_or0;
  assign f_u_dadda_cla32_fa509_xor1 = f_u_dadda_cla32_fa509_xor0 ^ f_u_dadda_cla32_fa486_or0;
  assign f_u_dadda_cla32_fa509_and1 = f_u_dadda_cla32_fa509_xor0 & f_u_dadda_cla32_fa486_or0;
  assign f_u_dadda_cla32_fa509_or0 = f_u_dadda_cla32_fa509_and0 | f_u_dadda_cla32_fa509_and1;
  assign f_u_dadda_cla32_and_31_9 = a[31] & b[9];
  assign f_u_dadda_cla32_and_30_10 = a[30] & b[10];
  assign f_u_dadda_cla32_fa510_xor0 = f_u_dadda_cla32_fa485_or0 ^ f_u_dadda_cla32_and_31_9;
  assign f_u_dadda_cla32_fa510_and0 = f_u_dadda_cla32_fa485_or0 & f_u_dadda_cla32_and_31_9;
  assign f_u_dadda_cla32_fa510_xor1 = f_u_dadda_cla32_fa510_xor0 ^ f_u_dadda_cla32_and_30_10;
  assign f_u_dadda_cla32_fa510_and1 = f_u_dadda_cla32_fa510_xor0 & f_u_dadda_cla32_and_30_10;
  assign f_u_dadda_cla32_fa510_or0 = f_u_dadda_cla32_fa510_and0 | f_u_dadda_cla32_fa510_and1;
  assign f_u_dadda_cla32_and_29_11 = a[29] & b[11];
  assign f_u_dadda_cla32_and_28_12 = a[28] & b[12];
  assign f_u_dadda_cla32_and_27_13 = a[27] & b[13];
  assign f_u_dadda_cla32_fa511_xor0 = f_u_dadda_cla32_and_29_11 ^ f_u_dadda_cla32_and_28_12;
  assign f_u_dadda_cla32_fa511_and0 = f_u_dadda_cla32_and_29_11 & f_u_dadda_cla32_and_28_12;
  assign f_u_dadda_cla32_fa511_xor1 = f_u_dadda_cla32_fa511_xor0 ^ f_u_dadda_cla32_and_27_13;
  assign f_u_dadda_cla32_fa511_and1 = f_u_dadda_cla32_fa511_xor0 & f_u_dadda_cla32_and_27_13;
  assign f_u_dadda_cla32_fa511_or0 = f_u_dadda_cla32_fa511_and0 | f_u_dadda_cla32_fa511_and1;
  assign f_u_dadda_cla32_and_26_14 = a[26] & b[14];
  assign f_u_dadda_cla32_and_25_15 = a[25] & b[15];
  assign f_u_dadda_cla32_and_24_16 = a[24] & b[16];
  assign f_u_dadda_cla32_fa512_xor0 = f_u_dadda_cla32_and_26_14 ^ f_u_dadda_cla32_and_25_15;
  assign f_u_dadda_cla32_fa512_and0 = f_u_dadda_cla32_and_26_14 & f_u_dadda_cla32_and_25_15;
  assign f_u_dadda_cla32_fa512_xor1 = f_u_dadda_cla32_fa512_xor0 ^ f_u_dadda_cla32_and_24_16;
  assign f_u_dadda_cla32_fa512_and1 = f_u_dadda_cla32_fa512_xor0 & f_u_dadda_cla32_and_24_16;
  assign f_u_dadda_cla32_fa512_or0 = f_u_dadda_cla32_fa512_and0 | f_u_dadda_cla32_fa512_and1;
  assign f_u_dadda_cla32_and_23_17 = a[23] & b[17];
  assign f_u_dadda_cla32_and_22_18 = a[22] & b[18];
  assign f_u_dadda_cla32_and_21_19 = a[21] & b[19];
  assign f_u_dadda_cla32_fa513_xor0 = f_u_dadda_cla32_and_23_17 ^ f_u_dadda_cla32_and_22_18;
  assign f_u_dadda_cla32_fa513_and0 = f_u_dadda_cla32_and_23_17 & f_u_dadda_cla32_and_22_18;
  assign f_u_dadda_cla32_fa513_xor1 = f_u_dadda_cla32_fa513_xor0 ^ f_u_dadda_cla32_and_21_19;
  assign f_u_dadda_cla32_fa513_and1 = f_u_dadda_cla32_fa513_xor0 & f_u_dadda_cla32_and_21_19;
  assign f_u_dadda_cla32_fa513_or0 = f_u_dadda_cla32_fa513_and0 | f_u_dadda_cla32_fa513_and1;
  assign f_u_dadda_cla32_and_20_20 = a[20] & b[20];
  assign f_u_dadda_cla32_and_19_21 = a[19] & b[21];
  assign f_u_dadda_cla32_and_18_22 = a[18] & b[22];
  assign f_u_dadda_cla32_fa514_xor0 = f_u_dadda_cla32_and_20_20 ^ f_u_dadda_cla32_and_19_21;
  assign f_u_dadda_cla32_fa514_and0 = f_u_dadda_cla32_and_20_20 & f_u_dadda_cla32_and_19_21;
  assign f_u_dadda_cla32_fa514_xor1 = f_u_dadda_cla32_fa514_xor0 ^ f_u_dadda_cla32_and_18_22;
  assign f_u_dadda_cla32_fa514_and1 = f_u_dadda_cla32_fa514_xor0 & f_u_dadda_cla32_and_18_22;
  assign f_u_dadda_cla32_fa514_or0 = f_u_dadda_cla32_fa514_and0 | f_u_dadda_cla32_fa514_and1;
  assign f_u_dadda_cla32_and_17_23 = a[17] & b[23];
  assign f_u_dadda_cla32_and_16_24 = a[16] & b[24];
  assign f_u_dadda_cla32_and_15_25 = a[15] & b[25];
  assign f_u_dadda_cla32_fa515_xor0 = f_u_dadda_cla32_and_17_23 ^ f_u_dadda_cla32_and_16_24;
  assign f_u_dadda_cla32_fa515_and0 = f_u_dadda_cla32_and_17_23 & f_u_dadda_cla32_and_16_24;
  assign f_u_dadda_cla32_fa515_xor1 = f_u_dadda_cla32_fa515_xor0 ^ f_u_dadda_cla32_and_15_25;
  assign f_u_dadda_cla32_fa515_and1 = f_u_dadda_cla32_fa515_xor0 & f_u_dadda_cla32_and_15_25;
  assign f_u_dadda_cla32_fa515_or0 = f_u_dadda_cla32_fa515_and0 | f_u_dadda_cla32_fa515_and1;
  assign f_u_dadda_cla32_and_14_26 = a[14] & b[26];
  assign f_u_dadda_cla32_and_13_27 = a[13] & b[27];
  assign f_u_dadda_cla32_and_12_28 = a[12] & b[28];
  assign f_u_dadda_cla32_fa516_xor0 = f_u_dadda_cla32_and_14_26 ^ f_u_dadda_cla32_and_13_27;
  assign f_u_dadda_cla32_fa516_and0 = f_u_dadda_cla32_and_14_26 & f_u_dadda_cla32_and_13_27;
  assign f_u_dadda_cla32_fa516_xor1 = f_u_dadda_cla32_fa516_xor0 ^ f_u_dadda_cla32_and_12_28;
  assign f_u_dadda_cla32_fa516_and1 = f_u_dadda_cla32_fa516_xor0 & f_u_dadda_cla32_and_12_28;
  assign f_u_dadda_cla32_fa516_or0 = f_u_dadda_cla32_fa516_and0 | f_u_dadda_cla32_fa516_and1;
  assign f_u_dadda_cla32_and_11_29 = a[11] & b[29];
  assign f_u_dadda_cla32_and_10_30 = a[10] & b[30];
  assign f_u_dadda_cla32_and_9_31 = a[9] & b[31];
  assign f_u_dadda_cla32_fa517_xor0 = f_u_dadda_cla32_and_11_29 ^ f_u_dadda_cla32_and_10_30;
  assign f_u_dadda_cla32_fa517_and0 = f_u_dadda_cla32_and_11_29 & f_u_dadda_cla32_and_10_30;
  assign f_u_dadda_cla32_fa517_xor1 = f_u_dadda_cla32_fa517_xor0 ^ f_u_dadda_cla32_and_9_31;
  assign f_u_dadda_cla32_fa517_and1 = f_u_dadda_cla32_fa517_xor0 & f_u_dadda_cla32_and_9_31;
  assign f_u_dadda_cla32_fa517_or0 = f_u_dadda_cla32_fa517_and0 | f_u_dadda_cla32_fa517_and1;
  assign f_u_dadda_cla32_fa518_xor0 = f_u_dadda_cla32_fa504_xor1 ^ f_u_dadda_cla32_fa505_xor1;
  assign f_u_dadda_cla32_fa518_and0 = f_u_dadda_cla32_fa504_xor1 & f_u_dadda_cla32_fa505_xor1;
  assign f_u_dadda_cla32_fa518_xor1 = f_u_dadda_cla32_fa518_xor0 ^ f_u_dadda_cla32_fa506_xor1;
  assign f_u_dadda_cla32_fa518_and1 = f_u_dadda_cla32_fa518_xor0 & f_u_dadda_cla32_fa506_xor1;
  assign f_u_dadda_cla32_fa518_or0 = f_u_dadda_cla32_fa518_and0 | f_u_dadda_cla32_fa518_and1;
  assign f_u_dadda_cla32_fa519_xor0 = f_u_dadda_cla32_fa507_xor1 ^ f_u_dadda_cla32_fa508_xor1;
  assign f_u_dadda_cla32_fa519_and0 = f_u_dadda_cla32_fa507_xor1 & f_u_dadda_cla32_fa508_xor1;
  assign f_u_dadda_cla32_fa519_xor1 = f_u_dadda_cla32_fa519_xor0 ^ f_u_dadda_cla32_fa509_xor1;
  assign f_u_dadda_cla32_fa519_and1 = f_u_dadda_cla32_fa519_xor0 & f_u_dadda_cla32_fa509_xor1;
  assign f_u_dadda_cla32_fa519_or0 = f_u_dadda_cla32_fa519_and0 | f_u_dadda_cla32_fa519_and1;
  assign f_u_dadda_cla32_fa520_xor0 = f_u_dadda_cla32_fa510_xor1 ^ f_u_dadda_cla32_fa511_xor1;
  assign f_u_dadda_cla32_fa520_and0 = f_u_dadda_cla32_fa510_xor1 & f_u_dadda_cla32_fa511_xor1;
  assign f_u_dadda_cla32_fa520_xor1 = f_u_dadda_cla32_fa520_xor0 ^ f_u_dadda_cla32_fa512_xor1;
  assign f_u_dadda_cla32_fa520_and1 = f_u_dadda_cla32_fa520_xor0 & f_u_dadda_cla32_fa512_xor1;
  assign f_u_dadda_cla32_fa520_or0 = f_u_dadda_cla32_fa520_and0 | f_u_dadda_cla32_fa520_and1;
  assign f_u_dadda_cla32_fa521_xor0 = f_u_dadda_cla32_fa513_xor1 ^ f_u_dadda_cla32_fa514_xor1;
  assign f_u_dadda_cla32_fa521_and0 = f_u_dadda_cla32_fa513_xor1 & f_u_dadda_cla32_fa514_xor1;
  assign f_u_dadda_cla32_fa521_xor1 = f_u_dadda_cla32_fa521_xor0 ^ f_u_dadda_cla32_fa515_xor1;
  assign f_u_dadda_cla32_fa521_and1 = f_u_dadda_cla32_fa521_xor0 & f_u_dadda_cla32_fa515_xor1;
  assign f_u_dadda_cla32_fa521_or0 = f_u_dadda_cla32_fa521_and0 | f_u_dadda_cla32_fa521_and1;
  assign f_u_dadda_cla32_fa522_xor0 = f_u_dadda_cla32_fa521_or0 ^ f_u_dadda_cla32_fa520_or0;
  assign f_u_dadda_cla32_fa522_and0 = f_u_dadda_cla32_fa521_or0 & f_u_dadda_cla32_fa520_or0;
  assign f_u_dadda_cla32_fa522_xor1 = f_u_dadda_cla32_fa522_xor0 ^ f_u_dadda_cla32_fa519_or0;
  assign f_u_dadda_cla32_fa522_and1 = f_u_dadda_cla32_fa522_xor0 & f_u_dadda_cla32_fa519_or0;
  assign f_u_dadda_cla32_fa522_or0 = f_u_dadda_cla32_fa522_and0 | f_u_dadda_cla32_fa522_and1;
  assign f_u_dadda_cla32_fa523_xor0 = f_u_dadda_cla32_fa518_or0 ^ f_u_dadda_cla32_fa517_or0;
  assign f_u_dadda_cla32_fa523_and0 = f_u_dadda_cla32_fa518_or0 & f_u_dadda_cla32_fa517_or0;
  assign f_u_dadda_cla32_fa523_xor1 = f_u_dadda_cla32_fa523_xor0 ^ f_u_dadda_cla32_fa516_or0;
  assign f_u_dadda_cla32_fa523_and1 = f_u_dadda_cla32_fa523_xor0 & f_u_dadda_cla32_fa516_or0;
  assign f_u_dadda_cla32_fa523_or0 = f_u_dadda_cla32_fa523_and0 | f_u_dadda_cla32_fa523_and1;
  assign f_u_dadda_cla32_fa524_xor0 = f_u_dadda_cla32_fa515_or0 ^ f_u_dadda_cla32_fa514_or0;
  assign f_u_dadda_cla32_fa524_and0 = f_u_dadda_cla32_fa515_or0 & f_u_dadda_cla32_fa514_or0;
  assign f_u_dadda_cla32_fa524_xor1 = f_u_dadda_cla32_fa524_xor0 ^ f_u_dadda_cla32_fa513_or0;
  assign f_u_dadda_cla32_fa524_and1 = f_u_dadda_cla32_fa524_xor0 & f_u_dadda_cla32_fa513_or0;
  assign f_u_dadda_cla32_fa524_or0 = f_u_dadda_cla32_fa524_and0 | f_u_dadda_cla32_fa524_and1;
  assign f_u_dadda_cla32_fa525_xor0 = f_u_dadda_cla32_fa512_or0 ^ f_u_dadda_cla32_fa511_or0;
  assign f_u_dadda_cla32_fa525_and0 = f_u_dadda_cla32_fa512_or0 & f_u_dadda_cla32_fa511_or0;
  assign f_u_dadda_cla32_fa525_xor1 = f_u_dadda_cla32_fa525_xor0 ^ f_u_dadda_cla32_fa510_or0;
  assign f_u_dadda_cla32_fa525_and1 = f_u_dadda_cla32_fa525_xor0 & f_u_dadda_cla32_fa510_or0;
  assign f_u_dadda_cla32_fa525_or0 = f_u_dadda_cla32_fa525_and0 | f_u_dadda_cla32_fa525_and1;
  assign f_u_dadda_cla32_fa526_xor0 = f_u_dadda_cla32_fa509_or0 ^ f_u_dadda_cla32_fa508_or0;
  assign f_u_dadda_cla32_fa526_and0 = f_u_dadda_cla32_fa509_or0 & f_u_dadda_cla32_fa508_or0;
  assign f_u_dadda_cla32_fa526_xor1 = f_u_dadda_cla32_fa526_xor0 ^ f_u_dadda_cla32_fa507_or0;
  assign f_u_dadda_cla32_fa526_and1 = f_u_dadda_cla32_fa526_xor0 & f_u_dadda_cla32_fa507_or0;
  assign f_u_dadda_cla32_fa526_or0 = f_u_dadda_cla32_fa526_and0 | f_u_dadda_cla32_fa526_and1;
  assign f_u_dadda_cla32_fa527_xor0 = f_u_dadda_cla32_fa506_or0 ^ f_u_dadda_cla32_fa505_or0;
  assign f_u_dadda_cla32_fa527_and0 = f_u_dadda_cla32_fa506_or0 & f_u_dadda_cla32_fa505_or0;
  assign f_u_dadda_cla32_fa527_xor1 = f_u_dadda_cla32_fa527_xor0 ^ f_u_dadda_cla32_fa504_or0;
  assign f_u_dadda_cla32_fa527_and1 = f_u_dadda_cla32_fa527_xor0 & f_u_dadda_cla32_fa504_or0;
  assign f_u_dadda_cla32_fa527_or0 = f_u_dadda_cla32_fa527_and0 | f_u_dadda_cla32_fa527_and1;
  assign f_u_dadda_cla32_and_31_10 = a[31] & b[10];
  assign f_u_dadda_cla32_and_30_11 = a[30] & b[11];
  assign f_u_dadda_cla32_and_29_12 = a[29] & b[12];
  assign f_u_dadda_cla32_fa528_xor0 = f_u_dadda_cla32_and_31_10 ^ f_u_dadda_cla32_and_30_11;
  assign f_u_dadda_cla32_fa528_and0 = f_u_dadda_cla32_and_31_10 & f_u_dadda_cla32_and_30_11;
  assign f_u_dadda_cla32_fa528_xor1 = f_u_dadda_cla32_fa528_xor0 ^ f_u_dadda_cla32_and_29_12;
  assign f_u_dadda_cla32_fa528_and1 = f_u_dadda_cla32_fa528_xor0 & f_u_dadda_cla32_and_29_12;
  assign f_u_dadda_cla32_fa528_or0 = f_u_dadda_cla32_fa528_and0 | f_u_dadda_cla32_fa528_and1;
  assign f_u_dadda_cla32_and_28_13 = a[28] & b[13];
  assign f_u_dadda_cla32_and_27_14 = a[27] & b[14];
  assign f_u_dadda_cla32_and_26_15 = a[26] & b[15];
  assign f_u_dadda_cla32_fa529_xor0 = f_u_dadda_cla32_and_28_13 ^ f_u_dadda_cla32_and_27_14;
  assign f_u_dadda_cla32_fa529_and0 = f_u_dadda_cla32_and_28_13 & f_u_dadda_cla32_and_27_14;
  assign f_u_dadda_cla32_fa529_xor1 = f_u_dadda_cla32_fa529_xor0 ^ f_u_dadda_cla32_and_26_15;
  assign f_u_dadda_cla32_fa529_and1 = f_u_dadda_cla32_fa529_xor0 & f_u_dadda_cla32_and_26_15;
  assign f_u_dadda_cla32_fa529_or0 = f_u_dadda_cla32_fa529_and0 | f_u_dadda_cla32_fa529_and1;
  assign f_u_dadda_cla32_and_25_16 = a[25] & b[16];
  assign f_u_dadda_cla32_and_24_17 = a[24] & b[17];
  assign f_u_dadda_cla32_and_23_18 = a[23] & b[18];
  assign f_u_dadda_cla32_fa530_xor0 = f_u_dadda_cla32_and_25_16 ^ f_u_dadda_cla32_and_24_17;
  assign f_u_dadda_cla32_fa530_and0 = f_u_dadda_cla32_and_25_16 & f_u_dadda_cla32_and_24_17;
  assign f_u_dadda_cla32_fa530_xor1 = f_u_dadda_cla32_fa530_xor0 ^ f_u_dadda_cla32_and_23_18;
  assign f_u_dadda_cla32_fa530_and1 = f_u_dadda_cla32_fa530_xor0 & f_u_dadda_cla32_and_23_18;
  assign f_u_dadda_cla32_fa530_or0 = f_u_dadda_cla32_fa530_and0 | f_u_dadda_cla32_fa530_and1;
  assign f_u_dadda_cla32_and_22_19 = a[22] & b[19];
  assign f_u_dadda_cla32_and_21_20 = a[21] & b[20];
  assign f_u_dadda_cla32_and_20_21 = a[20] & b[21];
  assign f_u_dadda_cla32_fa531_xor0 = f_u_dadda_cla32_and_22_19 ^ f_u_dadda_cla32_and_21_20;
  assign f_u_dadda_cla32_fa531_and0 = f_u_dadda_cla32_and_22_19 & f_u_dadda_cla32_and_21_20;
  assign f_u_dadda_cla32_fa531_xor1 = f_u_dadda_cla32_fa531_xor0 ^ f_u_dadda_cla32_and_20_21;
  assign f_u_dadda_cla32_fa531_and1 = f_u_dadda_cla32_fa531_xor0 & f_u_dadda_cla32_and_20_21;
  assign f_u_dadda_cla32_fa531_or0 = f_u_dadda_cla32_fa531_and0 | f_u_dadda_cla32_fa531_and1;
  assign f_u_dadda_cla32_and_19_22 = a[19] & b[22];
  assign f_u_dadda_cla32_and_18_23 = a[18] & b[23];
  assign f_u_dadda_cla32_and_17_24 = a[17] & b[24];
  assign f_u_dadda_cla32_fa532_xor0 = f_u_dadda_cla32_and_19_22 ^ f_u_dadda_cla32_and_18_23;
  assign f_u_dadda_cla32_fa532_and0 = f_u_dadda_cla32_and_19_22 & f_u_dadda_cla32_and_18_23;
  assign f_u_dadda_cla32_fa532_xor1 = f_u_dadda_cla32_fa532_xor0 ^ f_u_dadda_cla32_and_17_24;
  assign f_u_dadda_cla32_fa532_and1 = f_u_dadda_cla32_fa532_xor0 & f_u_dadda_cla32_and_17_24;
  assign f_u_dadda_cla32_fa532_or0 = f_u_dadda_cla32_fa532_and0 | f_u_dadda_cla32_fa532_and1;
  assign f_u_dadda_cla32_and_16_25 = a[16] & b[25];
  assign f_u_dadda_cla32_and_15_26 = a[15] & b[26];
  assign f_u_dadda_cla32_and_14_27 = a[14] & b[27];
  assign f_u_dadda_cla32_fa533_xor0 = f_u_dadda_cla32_and_16_25 ^ f_u_dadda_cla32_and_15_26;
  assign f_u_dadda_cla32_fa533_and0 = f_u_dadda_cla32_and_16_25 & f_u_dadda_cla32_and_15_26;
  assign f_u_dadda_cla32_fa533_xor1 = f_u_dadda_cla32_fa533_xor0 ^ f_u_dadda_cla32_and_14_27;
  assign f_u_dadda_cla32_fa533_and1 = f_u_dadda_cla32_fa533_xor0 & f_u_dadda_cla32_and_14_27;
  assign f_u_dadda_cla32_fa533_or0 = f_u_dadda_cla32_fa533_and0 | f_u_dadda_cla32_fa533_and1;
  assign f_u_dadda_cla32_and_13_28 = a[13] & b[28];
  assign f_u_dadda_cla32_and_12_29 = a[12] & b[29];
  assign f_u_dadda_cla32_and_11_30 = a[11] & b[30];
  assign f_u_dadda_cla32_fa534_xor0 = f_u_dadda_cla32_and_13_28 ^ f_u_dadda_cla32_and_12_29;
  assign f_u_dadda_cla32_fa534_and0 = f_u_dadda_cla32_and_13_28 & f_u_dadda_cla32_and_12_29;
  assign f_u_dadda_cla32_fa534_xor1 = f_u_dadda_cla32_fa534_xor0 ^ f_u_dadda_cla32_and_11_30;
  assign f_u_dadda_cla32_fa534_and1 = f_u_dadda_cla32_fa534_xor0 & f_u_dadda_cla32_and_11_30;
  assign f_u_dadda_cla32_fa534_or0 = f_u_dadda_cla32_fa534_and0 | f_u_dadda_cla32_fa534_and1;
  assign f_u_dadda_cla32_and_10_31 = a[10] & b[31];
  assign f_u_dadda_cla32_fa535_xor0 = f_u_dadda_cla32_and_10_31 ^ f_u_dadda_cla32_fa522_xor1;
  assign f_u_dadda_cla32_fa535_and0 = f_u_dadda_cla32_and_10_31 & f_u_dadda_cla32_fa522_xor1;
  assign f_u_dadda_cla32_fa535_xor1 = f_u_dadda_cla32_fa535_xor0 ^ f_u_dadda_cla32_fa523_xor1;
  assign f_u_dadda_cla32_fa535_and1 = f_u_dadda_cla32_fa535_xor0 & f_u_dadda_cla32_fa523_xor1;
  assign f_u_dadda_cla32_fa535_or0 = f_u_dadda_cla32_fa535_and0 | f_u_dadda_cla32_fa535_and1;
  assign f_u_dadda_cla32_fa536_xor0 = f_u_dadda_cla32_fa524_xor1 ^ f_u_dadda_cla32_fa525_xor1;
  assign f_u_dadda_cla32_fa536_and0 = f_u_dadda_cla32_fa524_xor1 & f_u_dadda_cla32_fa525_xor1;
  assign f_u_dadda_cla32_fa536_xor1 = f_u_dadda_cla32_fa536_xor0 ^ f_u_dadda_cla32_fa526_xor1;
  assign f_u_dadda_cla32_fa536_and1 = f_u_dadda_cla32_fa536_xor0 & f_u_dadda_cla32_fa526_xor1;
  assign f_u_dadda_cla32_fa536_or0 = f_u_dadda_cla32_fa536_and0 | f_u_dadda_cla32_fa536_and1;
  assign f_u_dadda_cla32_fa537_xor0 = f_u_dadda_cla32_fa527_xor1 ^ f_u_dadda_cla32_fa528_xor1;
  assign f_u_dadda_cla32_fa537_and0 = f_u_dadda_cla32_fa527_xor1 & f_u_dadda_cla32_fa528_xor1;
  assign f_u_dadda_cla32_fa537_xor1 = f_u_dadda_cla32_fa537_xor0 ^ f_u_dadda_cla32_fa529_xor1;
  assign f_u_dadda_cla32_fa537_and1 = f_u_dadda_cla32_fa537_xor0 & f_u_dadda_cla32_fa529_xor1;
  assign f_u_dadda_cla32_fa537_or0 = f_u_dadda_cla32_fa537_and0 | f_u_dadda_cla32_fa537_and1;
  assign f_u_dadda_cla32_fa538_xor0 = f_u_dadda_cla32_fa530_xor1 ^ f_u_dadda_cla32_fa531_xor1;
  assign f_u_dadda_cla32_fa538_and0 = f_u_dadda_cla32_fa530_xor1 & f_u_dadda_cla32_fa531_xor1;
  assign f_u_dadda_cla32_fa538_xor1 = f_u_dadda_cla32_fa538_xor0 ^ f_u_dadda_cla32_fa532_xor1;
  assign f_u_dadda_cla32_fa538_and1 = f_u_dadda_cla32_fa538_xor0 & f_u_dadda_cla32_fa532_xor1;
  assign f_u_dadda_cla32_fa538_or0 = f_u_dadda_cla32_fa538_and0 | f_u_dadda_cla32_fa538_and1;
  assign f_u_dadda_cla32_fa539_xor0 = f_u_dadda_cla32_fa538_or0 ^ f_u_dadda_cla32_fa537_or0;
  assign f_u_dadda_cla32_fa539_and0 = f_u_dadda_cla32_fa538_or0 & f_u_dadda_cla32_fa537_or0;
  assign f_u_dadda_cla32_fa539_xor1 = f_u_dadda_cla32_fa539_xor0 ^ f_u_dadda_cla32_fa536_or0;
  assign f_u_dadda_cla32_fa539_and1 = f_u_dadda_cla32_fa539_xor0 & f_u_dadda_cla32_fa536_or0;
  assign f_u_dadda_cla32_fa539_or0 = f_u_dadda_cla32_fa539_and0 | f_u_dadda_cla32_fa539_and1;
  assign f_u_dadda_cla32_fa540_xor0 = f_u_dadda_cla32_fa535_or0 ^ f_u_dadda_cla32_fa534_or0;
  assign f_u_dadda_cla32_fa540_and0 = f_u_dadda_cla32_fa535_or0 & f_u_dadda_cla32_fa534_or0;
  assign f_u_dadda_cla32_fa540_xor1 = f_u_dadda_cla32_fa540_xor0 ^ f_u_dadda_cla32_fa533_or0;
  assign f_u_dadda_cla32_fa540_and1 = f_u_dadda_cla32_fa540_xor0 & f_u_dadda_cla32_fa533_or0;
  assign f_u_dadda_cla32_fa540_or0 = f_u_dadda_cla32_fa540_and0 | f_u_dadda_cla32_fa540_and1;
  assign f_u_dadda_cla32_fa541_xor0 = f_u_dadda_cla32_fa532_or0 ^ f_u_dadda_cla32_fa531_or0;
  assign f_u_dadda_cla32_fa541_and0 = f_u_dadda_cla32_fa532_or0 & f_u_dadda_cla32_fa531_or0;
  assign f_u_dadda_cla32_fa541_xor1 = f_u_dadda_cla32_fa541_xor0 ^ f_u_dadda_cla32_fa530_or0;
  assign f_u_dadda_cla32_fa541_and1 = f_u_dadda_cla32_fa541_xor0 & f_u_dadda_cla32_fa530_or0;
  assign f_u_dadda_cla32_fa541_or0 = f_u_dadda_cla32_fa541_and0 | f_u_dadda_cla32_fa541_and1;
  assign f_u_dadda_cla32_fa542_xor0 = f_u_dadda_cla32_fa529_or0 ^ f_u_dadda_cla32_fa528_or0;
  assign f_u_dadda_cla32_fa542_and0 = f_u_dadda_cla32_fa529_or0 & f_u_dadda_cla32_fa528_or0;
  assign f_u_dadda_cla32_fa542_xor1 = f_u_dadda_cla32_fa542_xor0 ^ f_u_dadda_cla32_fa527_or0;
  assign f_u_dadda_cla32_fa542_and1 = f_u_dadda_cla32_fa542_xor0 & f_u_dadda_cla32_fa527_or0;
  assign f_u_dadda_cla32_fa542_or0 = f_u_dadda_cla32_fa542_and0 | f_u_dadda_cla32_fa542_and1;
  assign f_u_dadda_cla32_fa543_xor0 = f_u_dadda_cla32_fa526_or0 ^ f_u_dadda_cla32_fa525_or0;
  assign f_u_dadda_cla32_fa543_and0 = f_u_dadda_cla32_fa526_or0 & f_u_dadda_cla32_fa525_or0;
  assign f_u_dadda_cla32_fa543_xor1 = f_u_dadda_cla32_fa543_xor0 ^ f_u_dadda_cla32_fa524_or0;
  assign f_u_dadda_cla32_fa543_and1 = f_u_dadda_cla32_fa543_xor0 & f_u_dadda_cla32_fa524_or0;
  assign f_u_dadda_cla32_fa543_or0 = f_u_dadda_cla32_fa543_and0 | f_u_dadda_cla32_fa543_and1;
  assign f_u_dadda_cla32_and_31_11 = a[31] & b[11];
  assign f_u_dadda_cla32_fa544_xor0 = f_u_dadda_cla32_fa523_or0 ^ f_u_dadda_cla32_fa522_or0;
  assign f_u_dadda_cla32_fa544_and0 = f_u_dadda_cla32_fa523_or0 & f_u_dadda_cla32_fa522_or0;
  assign f_u_dadda_cla32_fa544_xor1 = f_u_dadda_cla32_fa544_xor0 ^ f_u_dadda_cla32_and_31_11;
  assign f_u_dadda_cla32_fa544_and1 = f_u_dadda_cla32_fa544_xor0 & f_u_dadda_cla32_and_31_11;
  assign f_u_dadda_cla32_fa544_or0 = f_u_dadda_cla32_fa544_and0 | f_u_dadda_cla32_fa544_and1;
  assign f_u_dadda_cla32_and_30_12 = a[30] & b[12];
  assign f_u_dadda_cla32_and_29_13 = a[29] & b[13];
  assign f_u_dadda_cla32_and_28_14 = a[28] & b[14];
  assign f_u_dadda_cla32_fa545_xor0 = f_u_dadda_cla32_and_30_12 ^ f_u_dadda_cla32_and_29_13;
  assign f_u_dadda_cla32_fa545_and0 = f_u_dadda_cla32_and_30_12 & f_u_dadda_cla32_and_29_13;
  assign f_u_dadda_cla32_fa545_xor1 = f_u_dadda_cla32_fa545_xor0 ^ f_u_dadda_cla32_and_28_14;
  assign f_u_dadda_cla32_fa545_and1 = f_u_dadda_cla32_fa545_xor0 & f_u_dadda_cla32_and_28_14;
  assign f_u_dadda_cla32_fa545_or0 = f_u_dadda_cla32_fa545_and0 | f_u_dadda_cla32_fa545_and1;
  assign f_u_dadda_cla32_and_27_15 = a[27] & b[15];
  assign f_u_dadda_cla32_and_26_16 = a[26] & b[16];
  assign f_u_dadda_cla32_and_25_17 = a[25] & b[17];
  assign f_u_dadda_cla32_fa546_xor0 = f_u_dadda_cla32_and_27_15 ^ f_u_dadda_cla32_and_26_16;
  assign f_u_dadda_cla32_fa546_and0 = f_u_dadda_cla32_and_27_15 & f_u_dadda_cla32_and_26_16;
  assign f_u_dadda_cla32_fa546_xor1 = f_u_dadda_cla32_fa546_xor0 ^ f_u_dadda_cla32_and_25_17;
  assign f_u_dadda_cla32_fa546_and1 = f_u_dadda_cla32_fa546_xor0 & f_u_dadda_cla32_and_25_17;
  assign f_u_dadda_cla32_fa546_or0 = f_u_dadda_cla32_fa546_and0 | f_u_dadda_cla32_fa546_and1;
  assign f_u_dadda_cla32_and_24_18 = a[24] & b[18];
  assign f_u_dadda_cla32_and_23_19 = a[23] & b[19];
  assign f_u_dadda_cla32_and_22_20 = a[22] & b[20];
  assign f_u_dadda_cla32_fa547_xor0 = f_u_dadda_cla32_and_24_18 ^ f_u_dadda_cla32_and_23_19;
  assign f_u_dadda_cla32_fa547_and0 = f_u_dadda_cla32_and_24_18 & f_u_dadda_cla32_and_23_19;
  assign f_u_dadda_cla32_fa547_xor1 = f_u_dadda_cla32_fa547_xor0 ^ f_u_dadda_cla32_and_22_20;
  assign f_u_dadda_cla32_fa547_and1 = f_u_dadda_cla32_fa547_xor0 & f_u_dadda_cla32_and_22_20;
  assign f_u_dadda_cla32_fa547_or0 = f_u_dadda_cla32_fa547_and0 | f_u_dadda_cla32_fa547_and1;
  assign f_u_dadda_cla32_and_21_21 = a[21] & b[21];
  assign f_u_dadda_cla32_and_20_22 = a[20] & b[22];
  assign f_u_dadda_cla32_and_19_23 = a[19] & b[23];
  assign f_u_dadda_cla32_fa548_xor0 = f_u_dadda_cla32_and_21_21 ^ f_u_dadda_cla32_and_20_22;
  assign f_u_dadda_cla32_fa548_and0 = f_u_dadda_cla32_and_21_21 & f_u_dadda_cla32_and_20_22;
  assign f_u_dadda_cla32_fa548_xor1 = f_u_dadda_cla32_fa548_xor0 ^ f_u_dadda_cla32_and_19_23;
  assign f_u_dadda_cla32_fa548_and1 = f_u_dadda_cla32_fa548_xor0 & f_u_dadda_cla32_and_19_23;
  assign f_u_dadda_cla32_fa548_or0 = f_u_dadda_cla32_fa548_and0 | f_u_dadda_cla32_fa548_and1;
  assign f_u_dadda_cla32_and_18_24 = a[18] & b[24];
  assign f_u_dadda_cla32_and_17_25 = a[17] & b[25];
  assign f_u_dadda_cla32_and_16_26 = a[16] & b[26];
  assign f_u_dadda_cla32_fa549_xor0 = f_u_dadda_cla32_and_18_24 ^ f_u_dadda_cla32_and_17_25;
  assign f_u_dadda_cla32_fa549_and0 = f_u_dadda_cla32_and_18_24 & f_u_dadda_cla32_and_17_25;
  assign f_u_dadda_cla32_fa549_xor1 = f_u_dadda_cla32_fa549_xor0 ^ f_u_dadda_cla32_and_16_26;
  assign f_u_dadda_cla32_fa549_and1 = f_u_dadda_cla32_fa549_xor0 & f_u_dadda_cla32_and_16_26;
  assign f_u_dadda_cla32_fa549_or0 = f_u_dadda_cla32_fa549_and0 | f_u_dadda_cla32_fa549_and1;
  assign f_u_dadda_cla32_and_15_27 = a[15] & b[27];
  assign f_u_dadda_cla32_and_14_28 = a[14] & b[28];
  assign f_u_dadda_cla32_and_13_29 = a[13] & b[29];
  assign f_u_dadda_cla32_fa550_xor0 = f_u_dadda_cla32_and_15_27 ^ f_u_dadda_cla32_and_14_28;
  assign f_u_dadda_cla32_fa550_and0 = f_u_dadda_cla32_and_15_27 & f_u_dadda_cla32_and_14_28;
  assign f_u_dadda_cla32_fa550_xor1 = f_u_dadda_cla32_fa550_xor0 ^ f_u_dadda_cla32_and_13_29;
  assign f_u_dadda_cla32_fa550_and1 = f_u_dadda_cla32_fa550_xor0 & f_u_dadda_cla32_and_13_29;
  assign f_u_dadda_cla32_fa550_or0 = f_u_dadda_cla32_fa550_and0 | f_u_dadda_cla32_fa550_and1;
  assign f_u_dadda_cla32_and_12_30 = a[12] & b[30];
  assign f_u_dadda_cla32_and_11_31 = a[11] & b[31];
  assign f_u_dadda_cla32_fa551_xor0 = f_u_dadda_cla32_and_12_30 ^ f_u_dadda_cla32_and_11_31;
  assign f_u_dadda_cla32_fa551_and0 = f_u_dadda_cla32_and_12_30 & f_u_dadda_cla32_and_11_31;
  assign f_u_dadda_cla32_fa551_xor1 = f_u_dadda_cla32_fa551_xor0 ^ f_u_dadda_cla32_fa539_xor1;
  assign f_u_dadda_cla32_fa551_and1 = f_u_dadda_cla32_fa551_xor0 & f_u_dadda_cla32_fa539_xor1;
  assign f_u_dadda_cla32_fa551_or0 = f_u_dadda_cla32_fa551_and0 | f_u_dadda_cla32_fa551_and1;
  assign f_u_dadda_cla32_fa552_xor0 = f_u_dadda_cla32_fa540_xor1 ^ f_u_dadda_cla32_fa541_xor1;
  assign f_u_dadda_cla32_fa552_and0 = f_u_dadda_cla32_fa540_xor1 & f_u_dadda_cla32_fa541_xor1;
  assign f_u_dadda_cla32_fa552_xor1 = f_u_dadda_cla32_fa552_xor0 ^ f_u_dadda_cla32_fa542_xor1;
  assign f_u_dadda_cla32_fa552_and1 = f_u_dadda_cla32_fa552_xor0 & f_u_dadda_cla32_fa542_xor1;
  assign f_u_dadda_cla32_fa552_or0 = f_u_dadda_cla32_fa552_and0 | f_u_dadda_cla32_fa552_and1;
  assign f_u_dadda_cla32_fa553_xor0 = f_u_dadda_cla32_fa543_xor1 ^ f_u_dadda_cla32_fa544_xor1;
  assign f_u_dadda_cla32_fa553_and0 = f_u_dadda_cla32_fa543_xor1 & f_u_dadda_cla32_fa544_xor1;
  assign f_u_dadda_cla32_fa553_xor1 = f_u_dadda_cla32_fa553_xor0 ^ f_u_dadda_cla32_fa545_xor1;
  assign f_u_dadda_cla32_fa553_and1 = f_u_dadda_cla32_fa553_xor0 & f_u_dadda_cla32_fa545_xor1;
  assign f_u_dadda_cla32_fa553_or0 = f_u_dadda_cla32_fa553_and0 | f_u_dadda_cla32_fa553_and1;
  assign f_u_dadda_cla32_fa554_xor0 = f_u_dadda_cla32_fa546_xor1 ^ f_u_dadda_cla32_fa547_xor1;
  assign f_u_dadda_cla32_fa554_and0 = f_u_dadda_cla32_fa546_xor1 & f_u_dadda_cla32_fa547_xor1;
  assign f_u_dadda_cla32_fa554_xor1 = f_u_dadda_cla32_fa554_xor0 ^ f_u_dadda_cla32_fa548_xor1;
  assign f_u_dadda_cla32_fa554_and1 = f_u_dadda_cla32_fa554_xor0 & f_u_dadda_cla32_fa548_xor1;
  assign f_u_dadda_cla32_fa554_or0 = f_u_dadda_cla32_fa554_and0 | f_u_dadda_cla32_fa554_and1;
  assign f_u_dadda_cla32_fa555_xor0 = f_u_dadda_cla32_fa554_or0 ^ f_u_dadda_cla32_fa553_or0;
  assign f_u_dadda_cla32_fa555_and0 = f_u_dadda_cla32_fa554_or0 & f_u_dadda_cla32_fa553_or0;
  assign f_u_dadda_cla32_fa555_xor1 = f_u_dadda_cla32_fa555_xor0 ^ f_u_dadda_cla32_fa552_or0;
  assign f_u_dadda_cla32_fa555_and1 = f_u_dadda_cla32_fa555_xor0 & f_u_dadda_cla32_fa552_or0;
  assign f_u_dadda_cla32_fa555_or0 = f_u_dadda_cla32_fa555_and0 | f_u_dadda_cla32_fa555_and1;
  assign f_u_dadda_cla32_fa556_xor0 = f_u_dadda_cla32_fa551_or0 ^ f_u_dadda_cla32_fa550_or0;
  assign f_u_dadda_cla32_fa556_and0 = f_u_dadda_cla32_fa551_or0 & f_u_dadda_cla32_fa550_or0;
  assign f_u_dadda_cla32_fa556_xor1 = f_u_dadda_cla32_fa556_xor0 ^ f_u_dadda_cla32_fa549_or0;
  assign f_u_dadda_cla32_fa556_and1 = f_u_dadda_cla32_fa556_xor0 & f_u_dadda_cla32_fa549_or0;
  assign f_u_dadda_cla32_fa556_or0 = f_u_dadda_cla32_fa556_and0 | f_u_dadda_cla32_fa556_and1;
  assign f_u_dadda_cla32_fa557_xor0 = f_u_dadda_cla32_fa548_or0 ^ f_u_dadda_cla32_fa547_or0;
  assign f_u_dadda_cla32_fa557_and0 = f_u_dadda_cla32_fa548_or0 & f_u_dadda_cla32_fa547_or0;
  assign f_u_dadda_cla32_fa557_xor1 = f_u_dadda_cla32_fa557_xor0 ^ f_u_dadda_cla32_fa546_or0;
  assign f_u_dadda_cla32_fa557_and1 = f_u_dadda_cla32_fa557_xor0 & f_u_dadda_cla32_fa546_or0;
  assign f_u_dadda_cla32_fa557_or0 = f_u_dadda_cla32_fa557_and0 | f_u_dadda_cla32_fa557_and1;
  assign f_u_dadda_cla32_fa558_xor0 = f_u_dadda_cla32_fa545_or0 ^ f_u_dadda_cla32_fa544_or0;
  assign f_u_dadda_cla32_fa558_and0 = f_u_dadda_cla32_fa545_or0 & f_u_dadda_cla32_fa544_or0;
  assign f_u_dadda_cla32_fa558_xor1 = f_u_dadda_cla32_fa558_xor0 ^ f_u_dadda_cla32_fa543_or0;
  assign f_u_dadda_cla32_fa558_and1 = f_u_dadda_cla32_fa558_xor0 & f_u_dadda_cla32_fa543_or0;
  assign f_u_dadda_cla32_fa558_or0 = f_u_dadda_cla32_fa558_and0 | f_u_dadda_cla32_fa558_and1;
  assign f_u_dadda_cla32_fa559_xor0 = f_u_dadda_cla32_fa542_or0 ^ f_u_dadda_cla32_fa541_or0;
  assign f_u_dadda_cla32_fa559_and0 = f_u_dadda_cla32_fa542_or0 & f_u_dadda_cla32_fa541_or0;
  assign f_u_dadda_cla32_fa559_xor1 = f_u_dadda_cla32_fa559_xor0 ^ f_u_dadda_cla32_fa540_or0;
  assign f_u_dadda_cla32_fa559_and1 = f_u_dadda_cla32_fa559_xor0 & f_u_dadda_cla32_fa540_or0;
  assign f_u_dadda_cla32_fa559_or0 = f_u_dadda_cla32_fa559_and0 | f_u_dadda_cla32_fa559_and1;
  assign f_u_dadda_cla32_and_31_12 = a[31] & b[12];
  assign f_u_dadda_cla32_and_30_13 = a[30] & b[13];
  assign f_u_dadda_cla32_fa560_xor0 = f_u_dadda_cla32_fa539_or0 ^ f_u_dadda_cla32_and_31_12;
  assign f_u_dadda_cla32_fa560_and0 = f_u_dadda_cla32_fa539_or0 & f_u_dadda_cla32_and_31_12;
  assign f_u_dadda_cla32_fa560_xor1 = f_u_dadda_cla32_fa560_xor0 ^ f_u_dadda_cla32_and_30_13;
  assign f_u_dadda_cla32_fa560_and1 = f_u_dadda_cla32_fa560_xor0 & f_u_dadda_cla32_and_30_13;
  assign f_u_dadda_cla32_fa560_or0 = f_u_dadda_cla32_fa560_and0 | f_u_dadda_cla32_fa560_and1;
  assign f_u_dadda_cla32_and_29_14 = a[29] & b[14];
  assign f_u_dadda_cla32_and_28_15 = a[28] & b[15];
  assign f_u_dadda_cla32_and_27_16 = a[27] & b[16];
  assign f_u_dadda_cla32_fa561_xor0 = f_u_dadda_cla32_and_29_14 ^ f_u_dadda_cla32_and_28_15;
  assign f_u_dadda_cla32_fa561_and0 = f_u_dadda_cla32_and_29_14 & f_u_dadda_cla32_and_28_15;
  assign f_u_dadda_cla32_fa561_xor1 = f_u_dadda_cla32_fa561_xor0 ^ f_u_dadda_cla32_and_27_16;
  assign f_u_dadda_cla32_fa561_and1 = f_u_dadda_cla32_fa561_xor0 & f_u_dadda_cla32_and_27_16;
  assign f_u_dadda_cla32_fa561_or0 = f_u_dadda_cla32_fa561_and0 | f_u_dadda_cla32_fa561_and1;
  assign f_u_dadda_cla32_and_26_17 = a[26] & b[17];
  assign f_u_dadda_cla32_and_25_18 = a[25] & b[18];
  assign f_u_dadda_cla32_and_24_19 = a[24] & b[19];
  assign f_u_dadda_cla32_fa562_xor0 = f_u_dadda_cla32_and_26_17 ^ f_u_dadda_cla32_and_25_18;
  assign f_u_dadda_cla32_fa562_and0 = f_u_dadda_cla32_and_26_17 & f_u_dadda_cla32_and_25_18;
  assign f_u_dadda_cla32_fa562_xor1 = f_u_dadda_cla32_fa562_xor0 ^ f_u_dadda_cla32_and_24_19;
  assign f_u_dadda_cla32_fa562_and1 = f_u_dadda_cla32_fa562_xor0 & f_u_dadda_cla32_and_24_19;
  assign f_u_dadda_cla32_fa562_or0 = f_u_dadda_cla32_fa562_and0 | f_u_dadda_cla32_fa562_and1;
  assign f_u_dadda_cla32_and_23_20 = a[23] & b[20];
  assign f_u_dadda_cla32_and_22_21 = a[22] & b[21];
  assign f_u_dadda_cla32_and_21_22 = a[21] & b[22];
  assign f_u_dadda_cla32_fa563_xor0 = f_u_dadda_cla32_and_23_20 ^ f_u_dadda_cla32_and_22_21;
  assign f_u_dadda_cla32_fa563_and0 = f_u_dadda_cla32_and_23_20 & f_u_dadda_cla32_and_22_21;
  assign f_u_dadda_cla32_fa563_xor1 = f_u_dadda_cla32_fa563_xor0 ^ f_u_dadda_cla32_and_21_22;
  assign f_u_dadda_cla32_fa563_and1 = f_u_dadda_cla32_fa563_xor0 & f_u_dadda_cla32_and_21_22;
  assign f_u_dadda_cla32_fa563_or0 = f_u_dadda_cla32_fa563_and0 | f_u_dadda_cla32_fa563_and1;
  assign f_u_dadda_cla32_and_20_23 = a[20] & b[23];
  assign f_u_dadda_cla32_and_19_24 = a[19] & b[24];
  assign f_u_dadda_cla32_and_18_25 = a[18] & b[25];
  assign f_u_dadda_cla32_fa564_xor0 = f_u_dadda_cla32_and_20_23 ^ f_u_dadda_cla32_and_19_24;
  assign f_u_dadda_cla32_fa564_and0 = f_u_dadda_cla32_and_20_23 & f_u_dadda_cla32_and_19_24;
  assign f_u_dadda_cla32_fa564_xor1 = f_u_dadda_cla32_fa564_xor0 ^ f_u_dadda_cla32_and_18_25;
  assign f_u_dadda_cla32_fa564_and1 = f_u_dadda_cla32_fa564_xor0 & f_u_dadda_cla32_and_18_25;
  assign f_u_dadda_cla32_fa564_or0 = f_u_dadda_cla32_fa564_and0 | f_u_dadda_cla32_fa564_and1;
  assign f_u_dadda_cla32_and_17_26 = a[17] & b[26];
  assign f_u_dadda_cla32_and_16_27 = a[16] & b[27];
  assign f_u_dadda_cla32_and_15_28 = a[15] & b[28];
  assign f_u_dadda_cla32_fa565_xor0 = f_u_dadda_cla32_and_17_26 ^ f_u_dadda_cla32_and_16_27;
  assign f_u_dadda_cla32_fa565_and0 = f_u_dadda_cla32_and_17_26 & f_u_dadda_cla32_and_16_27;
  assign f_u_dadda_cla32_fa565_xor1 = f_u_dadda_cla32_fa565_xor0 ^ f_u_dadda_cla32_and_15_28;
  assign f_u_dadda_cla32_fa565_and1 = f_u_dadda_cla32_fa565_xor0 & f_u_dadda_cla32_and_15_28;
  assign f_u_dadda_cla32_fa565_or0 = f_u_dadda_cla32_fa565_and0 | f_u_dadda_cla32_fa565_and1;
  assign f_u_dadda_cla32_and_14_29 = a[14] & b[29];
  assign f_u_dadda_cla32_and_13_30 = a[13] & b[30];
  assign f_u_dadda_cla32_and_12_31 = a[12] & b[31];
  assign f_u_dadda_cla32_fa566_xor0 = f_u_dadda_cla32_and_14_29 ^ f_u_dadda_cla32_and_13_30;
  assign f_u_dadda_cla32_fa566_and0 = f_u_dadda_cla32_and_14_29 & f_u_dadda_cla32_and_13_30;
  assign f_u_dadda_cla32_fa566_xor1 = f_u_dadda_cla32_fa566_xor0 ^ f_u_dadda_cla32_and_12_31;
  assign f_u_dadda_cla32_fa566_and1 = f_u_dadda_cla32_fa566_xor0 & f_u_dadda_cla32_and_12_31;
  assign f_u_dadda_cla32_fa566_or0 = f_u_dadda_cla32_fa566_and0 | f_u_dadda_cla32_fa566_and1;
  assign f_u_dadda_cla32_fa567_xor0 = f_u_dadda_cla32_fa555_xor1 ^ f_u_dadda_cla32_fa556_xor1;
  assign f_u_dadda_cla32_fa567_and0 = f_u_dadda_cla32_fa555_xor1 & f_u_dadda_cla32_fa556_xor1;
  assign f_u_dadda_cla32_fa567_xor1 = f_u_dadda_cla32_fa567_xor0 ^ f_u_dadda_cla32_fa557_xor1;
  assign f_u_dadda_cla32_fa567_and1 = f_u_dadda_cla32_fa567_xor0 & f_u_dadda_cla32_fa557_xor1;
  assign f_u_dadda_cla32_fa567_or0 = f_u_dadda_cla32_fa567_and0 | f_u_dadda_cla32_fa567_and1;
  assign f_u_dadda_cla32_fa568_xor0 = f_u_dadda_cla32_fa558_xor1 ^ f_u_dadda_cla32_fa559_xor1;
  assign f_u_dadda_cla32_fa568_and0 = f_u_dadda_cla32_fa558_xor1 & f_u_dadda_cla32_fa559_xor1;
  assign f_u_dadda_cla32_fa568_xor1 = f_u_dadda_cla32_fa568_xor0 ^ f_u_dadda_cla32_fa560_xor1;
  assign f_u_dadda_cla32_fa568_and1 = f_u_dadda_cla32_fa568_xor0 & f_u_dadda_cla32_fa560_xor1;
  assign f_u_dadda_cla32_fa568_or0 = f_u_dadda_cla32_fa568_and0 | f_u_dadda_cla32_fa568_and1;
  assign f_u_dadda_cla32_fa569_xor0 = f_u_dadda_cla32_fa561_xor1 ^ f_u_dadda_cla32_fa562_xor1;
  assign f_u_dadda_cla32_fa569_and0 = f_u_dadda_cla32_fa561_xor1 & f_u_dadda_cla32_fa562_xor1;
  assign f_u_dadda_cla32_fa569_xor1 = f_u_dadda_cla32_fa569_xor0 ^ f_u_dadda_cla32_fa563_xor1;
  assign f_u_dadda_cla32_fa569_and1 = f_u_dadda_cla32_fa569_xor0 & f_u_dadda_cla32_fa563_xor1;
  assign f_u_dadda_cla32_fa569_or0 = f_u_dadda_cla32_fa569_and0 | f_u_dadda_cla32_fa569_and1;
  assign f_u_dadda_cla32_fa570_xor0 = f_u_dadda_cla32_fa569_or0 ^ f_u_dadda_cla32_fa568_or0;
  assign f_u_dadda_cla32_fa570_and0 = f_u_dadda_cla32_fa569_or0 & f_u_dadda_cla32_fa568_or0;
  assign f_u_dadda_cla32_fa570_xor1 = f_u_dadda_cla32_fa570_xor0 ^ f_u_dadda_cla32_fa567_or0;
  assign f_u_dadda_cla32_fa570_and1 = f_u_dadda_cla32_fa570_xor0 & f_u_dadda_cla32_fa567_or0;
  assign f_u_dadda_cla32_fa570_or0 = f_u_dadda_cla32_fa570_and0 | f_u_dadda_cla32_fa570_and1;
  assign f_u_dadda_cla32_fa571_xor0 = f_u_dadda_cla32_fa566_or0 ^ f_u_dadda_cla32_fa565_or0;
  assign f_u_dadda_cla32_fa571_and0 = f_u_dadda_cla32_fa566_or0 & f_u_dadda_cla32_fa565_or0;
  assign f_u_dadda_cla32_fa571_xor1 = f_u_dadda_cla32_fa571_xor0 ^ f_u_dadda_cla32_fa564_or0;
  assign f_u_dadda_cla32_fa571_and1 = f_u_dadda_cla32_fa571_xor0 & f_u_dadda_cla32_fa564_or0;
  assign f_u_dadda_cla32_fa571_or0 = f_u_dadda_cla32_fa571_and0 | f_u_dadda_cla32_fa571_and1;
  assign f_u_dadda_cla32_fa572_xor0 = f_u_dadda_cla32_fa563_or0 ^ f_u_dadda_cla32_fa562_or0;
  assign f_u_dadda_cla32_fa572_and0 = f_u_dadda_cla32_fa563_or0 & f_u_dadda_cla32_fa562_or0;
  assign f_u_dadda_cla32_fa572_xor1 = f_u_dadda_cla32_fa572_xor0 ^ f_u_dadda_cla32_fa561_or0;
  assign f_u_dadda_cla32_fa572_and1 = f_u_dadda_cla32_fa572_xor0 & f_u_dadda_cla32_fa561_or0;
  assign f_u_dadda_cla32_fa572_or0 = f_u_dadda_cla32_fa572_and0 | f_u_dadda_cla32_fa572_and1;
  assign f_u_dadda_cla32_fa573_xor0 = f_u_dadda_cla32_fa560_or0 ^ f_u_dadda_cla32_fa559_or0;
  assign f_u_dadda_cla32_fa573_and0 = f_u_dadda_cla32_fa560_or0 & f_u_dadda_cla32_fa559_or0;
  assign f_u_dadda_cla32_fa573_xor1 = f_u_dadda_cla32_fa573_xor0 ^ f_u_dadda_cla32_fa558_or0;
  assign f_u_dadda_cla32_fa573_and1 = f_u_dadda_cla32_fa573_xor0 & f_u_dadda_cla32_fa558_or0;
  assign f_u_dadda_cla32_fa573_or0 = f_u_dadda_cla32_fa573_and0 | f_u_dadda_cla32_fa573_and1;
  assign f_u_dadda_cla32_fa574_xor0 = f_u_dadda_cla32_fa557_or0 ^ f_u_dadda_cla32_fa556_or0;
  assign f_u_dadda_cla32_fa574_and0 = f_u_dadda_cla32_fa557_or0 & f_u_dadda_cla32_fa556_or0;
  assign f_u_dadda_cla32_fa574_xor1 = f_u_dadda_cla32_fa574_xor0 ^ f_u_dadda_cla32_fa555_or0;
  assign f_u_dadda_cla32_fa574_and1 = f_u_dadda_cla32_fa574_xor0 & f_u_dadda_cla32_fa555_or0;
  assign f_u_dadda_cla32_fa574_or0 = f_u_dadda_cla32_fa574_and0 | f_u_dadda_cla32_fa574_and1;
  assign f_u_dadda_cla32_and_31_13 = a[31] & b[13];
  assign f_u_dadda_cla32_and_30_14 = a[30] & b[14];
  assign f_u_dadda_cla32_and_29_15 = a[29] & b[15];
  assign f_u_dadda_cla32_fa575_xor0 = f_u_dadda_cla32_and_31_13 ^ f_u_dadda_cla32_and_30_14;
  assign f_u_dadda_cla32_fa575_and0 = f_u_dadda_cla32_and_31_13 & f_u_dadda_cla32_and_30_14;
  assign f_u_dadda_cla32_fa575_xor1 = f_u_dadda_cla32_fa575_xor0 ^ f_u_dadda_cla32_and_29_15;
  assign f_u_dadda_cla32_fa575_and1 = f_u_dadda_cla32_fa575_xor0 & f_u_dadda_cla32_and_29_15;
  assign f_u_dadda_cla32_fa575_or0 = f_u_dadda_cla32_fa575_and0 | f_u_dadda_cla32_fa575_and1;
  assign f_u_dadda_cla32_and_28_16 = a[28] & b[16];
  assign f_u_dadda_cla32_and_27_17 = a[27] & b[17];
  assign f_u_dadda_cla32_and_26_18 = a[26] & b[18];
  assign f_u_dadda_cla32_fa576_xor0 = f_u_dadda_cla32_and_28_16 ^ f_u_dadda_cla32_and_27_17;
  assign f_u_dadda_cla32_fa576_and0 = f_u_dadda_cla32_and_28_16 & f_u_dadda_cla32_and_27_17;
  assign f_u_dadda_cla32_fa576_xor1 = f_u_dadda_cla32_fa576_xor0 ^ f_u_dadda_cla32_and_26_18;
  assign f_u_dadda_cla32_fa576_and1 = f_u_dadda_cla32_fa576_xor0 & f_u_dadda_cla32_and_26_18;
  assign f_u_dadda_cla32_fa576_or0 = f_u_dadda_cla32_fa576_and0 | f_u_dadda_cla32_fa576_and1;
  assign f_u_dadda_cla32_and_25_19 = a[25] & b[19];
  assign f_u_dadda_cla32_and_24_20 = a[24] & b[20];
  assign f_u_dadda_cla32_and_23_21 = a[23] & b[21];
  assign f_u_dadda_cla32_fa577_xor0 = f_u_dadda_cla32_and_25_19 ^ f_u_dadda_cla32_and_24_20;
  assign f_u_dadda_cla32_fa577_and0 = f_u_dadda_cla32_and_25_19 & f_u_dadda_cla32_and_24_20;
  assign f_u_dadda_cla32_fa577_xor1 = f_u_dadda_cla32_fa577_xor0 ^ f_u_dadda_cla32_and_23_21;
  assign f_u_dadda_cla32_fa577_and1 = f_u_dadda_cla32_fa577_xor0 & f_u_dadda_cla32_and_23_21;
  assign f_u_dadda_cla32_fa577_or0 = f_u_dadda_cla32_fa577_and0 | f_u_dadda_cla32_fa577_and1;
  assign f_u_dadda_cla32_and_22_22 = a[22] & b[22];
  assign f_u_dadda_cla32_and_21_23 = a[21] & b[23];
  assign f_u_dadda_cla32_and_20_24 = a[20] & b[24];
  assign f_u_dadda_cla32_fa578_xor0 = f_u_dadda_cla32_and_22_22 ^ f_u_dadda_cla32_and_21_23;
  assign f_u_dadda_cla32_fa578_and0 = f_u_dadda_cla32_and_22_22 & f_u_dadda_cla32_and_21_23;
  assign f_u_dadda_cla32_fa578_xor1 = f_u_dadda_cla32_fa578_xor0 ^ f_u_dadda_cla32_and_20_24;
  assign f_u_dadda_cla32_fa578_and1 = f_u_dadda_cla32_fa578_xor0 & f_u_dadda_cla32_and_20_24;
  assign f_u_dadda_cla32_fa578_or0 = f_u_dadda_cla32_fa578_and0 | f_u_dadda_cla32_fa578_and1;
  assign f_u_dadda_cla32_and_19_25 = a[19] & b[25];
  assign f_u_dadda_cla32_and_18_26 = a[18] & b[26];
  assign f_u_dadda_cla32_and_17_27 = a[17] & b[27];
  assign f_u_dadda_cla32_fa579_xor0 = f_u_dadda_cla32_and_19_25 ^ f_u_dadda_cla32_and_18_26;
  assign f_u_dadda_cla32_fa579_and0 = f_u_dadda_cla32_and_19_25 & f_u_dadda_cla32_and_18_26;
  assign f_u_dadda_cla32_fa579_xor1 = f_u_dadda_cla32_fa579_xor0 ^ f_u_dadda_cla32_and_17_27;
  assign f_u_dadda_cla32_fa579_and1 = f_u_dadda_cla32_fa579_xor0 & f_u_dadda_cla32_and_17_27;
  assign f_u_dadda_cla32_fa579_or0 = f_u_dadda_cla32_fa579_and0 | f_u_dadda_cla32_fa579_and1;
  assign f_u_dadda_cla32_and_16_28 = a[16] & b[28];
  assign f_u_dadda_cla32_and_15_29 = a[15] & b[29];
  assign f_u_dadda_cla32_and_14_30 = a[14] & b[30];
  assign f_u_dadda_cla32_fa580_xor0 = f_u_dadda_cla32_and_16_28 ^ f_u_dadda_cla32_and_15_29;
  assign f_u_dadda_cla32_fa580_and0 = f_u_dadda_cla32_and_16_28 & f_u_dadda_cla32_and_15_29;
  assign f_u_dadda_cla32_fa580_xor1 = f_u_dadda_cla32_fa580_xor0 ^ f_u_dadda_cla32_and_14_30;
  assign f_u_dadda_cla32_fa580_and1 = f_u_dadda_cla32_fa580_xor0 & f_u_dadda_cla32_and_14_30;
  assign f_u_dadda_cla32_fa580_or0 = f_u_dadda_cla32_fa580_and0 | f_u_dadda_cla32_fa580_and1;
  assign f_u_dadda_cla32_and_13_31 = a[13] & b[31];
  assign f_u_dadda_cla32_fa581_xor0 = f_u_dadda_cla32_and_13_31 ^ f_u_dadda_cla32_fa570_xor1;
  assign f_u_dadda_cla32_fa581_and0 = f_u_dadda_cla32_and_13_31 & f_u_dadda_cla32_fa570_xor1;
  assign f_u_dadda_cla32_fa581_xor1 = f_u_dadda_cla32_fa581_xor0 ^ f_u_dadda_cla32_fa571_xor1;
  assign f_u_dadda_cla32_fa581_and1 = f_u_dadda_cla32_fa581_xor0 & f_u_dadda_cla32_fa571_xor1;
  assign f_u_dadda_cla32_fa581_or0 = f_u_dadda_cla32_fa581_and0 | f_u_dadda_cla32_fa581_and1;
  assign f_u_dadda_cla32_fa582_xor0 = f_u_dadda_cla32_fa572_xor1 ^ f_u_dadda_cla32_fa573_xor1;
  assign f_u_dadda_cla32_fa582_and0 = f_u_dadda_cla32_fa572_xor1 & f_u_dadda_cla32_fa573_xor1;
  assign f_u_dadda_cla32_fa582_xor1 = f_u_dadda_cla32_fa582_xor0 ^ f_u_dadda_cla32_fa574_xor1;
  assign f_u_dadda_cla32_fa582_and1 = f_u_dadda_cla32_fa582_xor0 & f_u_dadda_cla32_fa574_xor1;
  assign f_u_dadda_cla32_fa582_or0 = f_u_dadda_cla32_fa582_and0 | f_u_dadda_cla32_fa582_and1;
  assign f_u_dadda_cla32_fa583_xor0 = f_u_dadda_cla32_fa575_xor1 ^ f_u_dadda_cla32_fa576_xor1;
  assign f_u_dadda_cla32_fa583_and0 = f_u_dadda_cla32_fa575_xor1 & f_u_dadda_cla32_fa576_xor1;
  assign f_u_dadda_cla32_fa583_xor1 = f_u_dadda_cla32_fa583_xor0 ^ f_u_dadda_cla32_fa577_xor1;
  assign f_u_dadda_cla32_fa583_and1 = f_u_dadda_cla32_fa583_xor0 & f_u_dadda_cla32_fa577_xor1;
  assign f_u_dadda_cla32_fa583_or0 = f_u_dadda_cla32_fa583_and0 | f_u_dadda_cla32_fa583_and1;
  assign f_u_dadda_cla32_fa584_xor0 = f_u_dadda_cla32_fa583_or0 ^ f_u_dadda_cla32_fa582_or0;
  assign f_u_dadda_cla32_fa584_and0 = f_u_dadda_cla32_fa583_or0 & f_u_dadda_cla32_fa582_or0;
  assign f_u_dadda_cla32_fa584_xor1 = f_u_dadda_cla32_fa584_xor0 ^ f_u_dadda_cla32_fa581_or0;
  assign f_u_dadda_cla32_fa584_and1 = f_u_dadda_cla32_fa584_xor0 & f_u_dadda_cla32_fa581_or0;
  assign f_u_dadda_cla32_fa584_or0 = f_u_dadda_cla32_fa584_and0 | f_u_dadda_cla32_fa584_and1;
  assign f_u_dadda_cla32_fa585_xor0 = f_u_dadda_cla32_fa580_or0 ^ f_u_dadda_cla32_fa579_or0;
  assign f_u_dadda_cla32_fa585_and0 = f_u_dadda_cla32_fa580_or0 & f_u_dadda_cla32_fa579_or0;
  assign f_u_dadda_cla32_fa585_xor1 = f_u_dadda_cla32_fa585_xor0 ^ f_u_dadda_cla32_fa578_or0;
  assign f_u_dadda_cla32_fa585_and1 = f_u_dadda_cla32_fa585_xor0 & f_u_dadda_cla32_fa578_or0;
  assign f_u_dadda_cla32_fa585_or0 = f_u_dadda_cla32_fa585_and0 | f_u_dadda_cla32_fa585_and1;
  assign f_u_dadda_cla32_fa586_xor0 = f_u_dadda_cla32_fa577_or0 ^ f_u_dadda_cla32_fa576_or0;
  assign f_u_dadda_cla32_fa586_and0 = f_u_dadda_cla32_fa577_or0 & f_u_dadda_cla32_fa576_or0;
  assign f_u_dadda_cla32_fa586_xor1 = f_u_dadda_cla32_fa586_xor0 ^ f_u_dadda_cla32_fa575_or0;
  assign f_u_dadda_cla32_fa586_and1 = f_u_dadda_cla32_fa586_xor0 & f_u_dadda_cla32_fa575_or0;
  assign f_u_dadda_cla32_fa586_or0 = f_u_dadda_cla32_fa586_and0 | f_u_dadda_cla32_fa586_and1;
  assign f_u_dadda_cla32_fa587_xor0 = f_u_dadda_cla32_fa574_or0 ^ f_u_dadda_cla32_fa573_or0;
  assign f_u_dadda_cla32_fa587_and0 = f_u_dadda_cla32_fa574_or0 & f_u_dadda_cla32_fa573_or0;
  assign f_u_dadda_cla32_fa587_xor1 = f_u_dadda_cla32_fa587_xor0 ^ f_u_dadda_cla32_fa572_or0;
  assign f_u_dadda_cla32_fa587_and1 = f_u_dadda_cla32_fa587_xor0 & f_u_dadda_cla32_fa572_or0;
  assign f_u_dadda_cla32_fa587_or0 = f_u_dadda_cla32_fa587_and0 | f_u_dadda_cla32_fa587_and1;
  assign f_u_dadda_cla32_and_31_14 = a[31] & b[14];
  assign f_u_dadda_cla32_fa588_xor0 = f_u_dadda_cla32_fa571_or0 ^ f_u_dadda_cla32_fa570_or0;
  assign f_u_dadda_cla32_fa588_and0 = f_u_dadda_cla32_fa571_or0 & f_u_dadda_cla32_fa570_or0;
  assign f_u_dadda_cla32_fa588_xor1 = f_u_dadda_cla32_fa588_xor0 ^ f_u_dadda_cla32_and_31_14;
  assign f_u_dadda_cla32_fa588_and1 = f_u_dadda_cla32_fa588_xor0 & f_u_dadda_cla32_and_31_14;
  assign f_u_dadda_cla32_fa588_or0 = f_u_dadda_cla32_fa588_and0 | f_u_dadda_cla32_fa588_and1;
  assign f_u_dadda_cla32_and_30_15 = a[30] & b[15];
  assign f_u_dadda_cla32_and_29_16 = a[29] & b[16];
  assign f_u_dadda_cla32_and_28_17 = a[28] & b[17];
  assign f_u_dadda_cla32_fa589_xor0 = f_u_dadda_cla32_and_30_15 ^ f_u_dadda_cla32_and_29_16;
  assign f_u_dadda_cla32_fa589_and0 = f_u_dadda_cla32_and_30_15 & f_u_dadda_cla32_and_29_16;
  assign f_u_dadda_cla32_fa589_xor1 = f_u_dadda_cla32_fa589_xor0 ^ f_u_dadda_cla32_and_28_17;
  assign f_u_dadda_cla32_fa589_and1 = f_u_dadda_cla32_fa589_xor0 & f_u_dadda_cla32_and_28_17;
  assign f_u_dadda_cla32_fa589_or0 = f_u_dadda_cla32_fa589_and0 | f_u_dadda_cla32_fa589_and1;
  assign f_u_dadda_cla32_and_27_18 = a[27] & b[18];
  assign f_u_dadda_cla32_and_26_19 = a[26] & b[19];
  assign f_u_dadda_cla32_and_25_20 = a[25] & b[20];
  assign f_u_dadda_cla32_fa590_xor0 = f_u_dadda_cla32_and_27_18 ^ f_u_dadda_cla32_and_26_19;
  assign f_u_dadda_cla32_fa590_and0 = f_u_dadda_cla32_and_27_18 & f_u_dadda_cla32_and_26_19;
  assign f_u_dadda_cla32_fa590_xor1 = f_u_dadda_cla32_fa590_xor0 ^ f_u_dadda_cla32_and_25_20;
  assign f_u_dadda_cla32_fa590_and1 = f_u_dadda_cla32_fa590_xor0 & f_u_dadda_cla32_and_25_20;
  assign f_u_dadda_cla32_fa590_or0 = f_u_dadda_cla32_fa590_and0 | f_u_dadda_cla32_fa590_and1;
  assign f_u_dadda_cla32_and_24_21 = a[24] & b[21];
  assign f_u_dadda_cla32_and_23_22 = a[23] & b[22];
  assign f_u_dadda_cla32_and_22_23 = a[22] & b[23];
  assign f_u_dadda_cla32_fa591_xor0 = f_u_dadda_cla32_and_24_21 ^ f_u_dadda_cla32_and_23_22;
  assign f_u_dadda_cla32_fa591_and0 = f_u_dadda_cla32_and_24_21 & f_u_dadda_cla32_and_23_22;
  assign f_u_dadda_cla32_fa591_xor1 = f_u_dadda_cla32_fa591_xor0 ^ f_u_dadda_cla32_and_22_23;
  assign f_u_dadda_cla32_fa591_and1 = f_u_dadda_cla32_fa591_xor0 & f_u_dadda_cla32_and_22_23;
  assign f_u_dadda_cla32_fa591_or0 = f_u_dadda_cla32_fa591_and0 | f_u_dadda_cla32_fa591_and1;
  assign f_u_dadda_cla32_and_21_24 = a[21] & b[24];
  assign f_u_dadda_cla32_and_20_25 = a[20] & b[25];
  assign f_u_dadda_cla32_and_19_26 = a[19] & b[26];
  assign f_u_dadda_cla32_fa592_xor0 = f_u_dadda_cla32_and_21_24 ^ f_u_dadda_cla32_and_20_25;
  assign f_u_dadda_cla32_fa592_and0 = f_u_dadda_cla32_and_21_24 & f_u_dadda_cla32_and_20_25;
  assign f_u_dadda_cla32_fa592_xor1 = f_u_dadda_cla32_fa592_xor0 ^ f_u_dadda_cla32_and_19_26;
  assign f_u_dadda_cla32_fa592_and1 = f_u_dadda_cla32_fa592_xor0 & f_u_dadda_cla32_and_19_26;
  assign f_u_dadda_cla32_fa592_or0 = f_u_dadda_cla32_fa592_and0 | f_u_dadda_cla32_fa592_and1;
  assign f_u_dadda_cla32_and_18_27 = a[18] & b[27];
  assign f_u_dadda_cla32_and_17_28 = a[17] & b[28];
  assign f_u_dadda_cla32_and_16_29 = a[16] & b[29];
  assign f_u_dadda_cla32_fa593_xor0 = f_u_dadda_cla32_and_18_27 ^ f_u_dadda_cla32_and_17_28;
  assign f_u_dadda_cla32_fa593_and0 = f_u_dadda_cla32_and_18_27 & f_u_dadda_cla32_and_17_28;
  assign f_u_dadda_cla32_fa593_xor1 = f_u_dadda_cla32_fa593_xor0 ^ f_u_dadda_cla32_and_16_29;
  assign f_u_dadda_cla32_fa593_and1 = f_u_dadda_cla32_fa593_xor0 & f_u_dadda_cla32_and_16_29;
  assign f_u_dadda_cla32_fa593_or0 = f_u_dadda_cla32_fa593_and0 | f_u_dadda_cla32_fa593_and1;
  assign f_u_dadda_cla32_and_15_30 = a[15] & b[30];
  assign f_u_dadda_cla32_and_14_31 = a[14] & b[31];
  assign f_u_dadda_cla32_fa594_xor0 = f_u_dadda_cla32_and_15_30 ^ f_u_dadda_cla32_and_14_31;
  assign f_u_dadda_cla32_fa594_and0 = f_u_dadda_cla32_and_15_30 & f_u_dadda_cla32_and_14_31;
  assign f_u_dadda_cla32_fa594_xor1 = f_u_dadda_cla32_fa594_xor0 ^ f_u_dadda_cla32_fa584_xor1;
  assign f_u_dadda_cla32_fa594_and1 = f_u_dadda_cla32_fa594_xor0 & f_u_dadda_cla32_fa584_xor1;
  assign f_u_dadda_cla32_fa594_or0 = f_u_dadda_cla32_fa594_and0 | f_u_dadda_cla32_fa594_and1;
  assign f_u_dadda_cla32_fa595_xor0 = f_u_dadda_cla32_fa585_xor1 ^ f_u_dadda_cla32_fa586_xor1;
  assign f_u_dadda_cla32_fa595_and0 = f_u_dadda_cla32_fa585_xor1 & f_u_dadda_cla32_fa586_xor1;
  assign f_u_dadda_cla32_fa595_xor1 = f_u_dadda_cla32_fa595_xor0 ^ f_u_dadda_cla32_fa587_xor1;
  assign f_u_dadda_cla32_fa595_and1 = f_u_dadda_cla32_fa595_xor0 & f_u_dadda_cla32_fa587_xor1;
  assign f_u_dadda_cla32_fa595_or0 = f_u_dadda_cla32_fa595_and0 | f_u_dadda_cla32_fa595_and1;
  assign f_u_dadda_cla32_fa596_xor0 = f_u_dadda_cla32_fa588_xor1 ^ f_u_dadda_cla32_fa589_xor1;
  assign f_u_dadda_cla32_fa596_and0 = f_u_dadda_cla32_fa588_xor1 & f_u_dadda_cla32_fa589_xor1;
  assign f_u_dadda_cla32_fa596_xor1 = f_u_dadda_cla32_fa596_xor0 ^ f_u_dadda_cla32_fa590_xor1;
  assign f_u_dadda_cla32_fa596_and1 = f_u_dadda_cla32_fa596_xor0 & f_u_dadda_cla32_fa590_xor1;
  assign f_u_dadda_cla32_fa596_or0 = f_u_dadda_cla32_fa596_and0 | f_u_dadda_cla32_fa596_and1;
  assign f_u_dadda_cla32_fa597_xor0 = f_u_dadda_cla32_fa596_or0 ^ f_u_dadda_cla32_fa595_or0;
  assign f_u_dadda_cla32_fa597_and0 = f_u_dadda_cla32_fa596_or0 & f_u_dadda_cla32_fa595_or0;
  assign f_u_dadda_cla32_fa597_xor1 = f_u_dadda_cla32_fa597_xor0 ^ f_u_dadda_cla32_fa594_or0;
  assign f_u_dadda_cla32_fa597_and1 = f_u_dadda_cla32_fa597_xor0 & f_u_dadda_cla32_fa594_or0;
  assign f_u_dadda_cla32_fa597_or0 = f_u_dadda_cla32_fa597_and0 | f_u_dadda_cla32_fa597_and1;
  assign f_u_dadda_cla32_fa598_xor0 = f_u_dadda_cla32_fa593_or0 ^ f_u_dadda_cla32_fa592_or0;
  assign f_u_dadda_cla32_fa598_and0 = f_u_dadda_cla32_fa593_or0 & f_u_dadda_cla32_fa592_or0;
  assign f_u_dadda_cla32_fa598_xor1 = f_u_dadda_cla32_fa598_xor0 ^ f_u_dadda_cla32_fa591_or0;
  assign f_u_dadda_cla32_fa598_and1 = f_u_dadda_cla32_fa598_xor0 & f_u_dadda_cla32_fa591_or0;
  assign f_u_dadda_cla32_fa598_or0 = f_u_dadda_cla32_fa598_and0 | f_u_dadda_cla32_fa598_and1;
  assign f_u_dadda_cla32_fa599_xor0 = f_u_dadda_cla32_fa590_or0 ^ f_u_dadda_cla32_fa589_or0;
  assign f_u_dadda_cla32_fa599_and0 = f_u_dadda_cla32_fa590_or0 & f_u_dadda_cla32_fa589_or0;
  assign f_u_dadda_cla32_fa599_xor1 = f_u_dadda_cla32_fa599_xor0 ^ f_u_dadda_cla32_fa588_or0;
  assign f_u_dadda_cla32_fa599_and1 = f_u_dadda_cla32_fa599_xor0 & f_u_dadda_cla32_fa588_or0;
  assign f_u_dadda_cla32_fa599_or0 = f_u_dadda_cla32_fa599_and0 | f_u_dadda_cla32_fa599_and1;
  assign f_u_dadda_cla32_fa600_xor0 = f_u_dadda_cla32_fa587_or0 ^ f_u_dadda_cla32_fa586_or0;
  assign f_u_dadda_cla32_fa600_and0 = f_u_dadda_cla32_fa587_or0 & f_u_dadda_cla32_fa586_or0;
  assign f_u_dadda_cla32_fa600_xor1 = f_u_dadda_cla32_fa600_xor0 ^ f_u_dadda_cla32_fa585_or0;
  assign f_u_dadda_cla32_fa600_and1 = f_u_dadda_cla32_fa600_xor0 & f_u_dadda_cla32_fa585_or0;
  assign f_u_dadda_cla32_fa600_or0 = f_u_dadda_cla32_fa600_and0 | f_u_dadda_cla32_fa600_and1;
  assign f_u_dadda_cla32_and_31_15 = a[31] & b[15];
  assign f_u_dadda_cla32_and_30_16 = a[30] & b[16];
  assign f_u_dadda_cla32_fa601_xor0 = f_u_dadda_cla32_fa584_or0 ^ f_u_dadda_cla32_and_31_15;
  assign f_u_dadda_cla32_fa601_and0 = f_u_dadda_cla32_fa584_or0 & f_u_dadda_cla32_and_31_15;
  assign f_u_dadda_cla32_fa601_xor1 = f_u_dadda_cla32_fa601_xor0 ^ f_u_dadda_cla32_and_30_16;
  assign f_u_dadda_cla32_fa601_and1 = f_u_dadda_cla32_fa601_xor0 & f_u_dadda_cla32_and_30_16;
  assign f_u_dadda_cla32_fa601_or0 = f_u_dadda_cla32_fa601_and0 | f_u_dadda_cla32_fa601_and1;
  assign f_u_dadda_cla32_and_29_17 = a[29] & b[17];
  assign f_u_dadda_cla32_and_28_18 = a[28] & b[18];
  assign f_u_dadda_cla32_and_27_19 = a[27] & b[19];
  assign f_u_dadda_cla32_fa602_xor0 = f_u_dadda_cla32_and_29_17 ^ f_u_dadda_cla32_and_28_18;
  assign f_u_dadda_cla32_fa602_and0 = f_u_dadda_cla32_and_29_17 & f_u_dadda_cla32_and_28_18;
  assign f_u_dadda_cla32_fa602_xor1 = f_u_dadda_cla32_fa602_xor0 ^ f_u_dadda_cla32_and_27_19;
  assign f_u_dadda_cla32_fa602_and1 = f_u_dadda_cla32_fa602_xor0 & f_u_dadda_cla32_and_27_19;
  assign f_u_dadda_cla32_fa602_or0 = f_u_dadda_cla32_fa602_and0 | f_u_dadda_cla32_fa602_and1;
  assign f_u_dadda_cla32_and_26_20 = a[26] & b[20];
  assign f_u_dadda_cla32_and_25_21 = a[25] & b[21];
  assign f_u_dadda_cla32_and_24_22 = a[24] & b[22];
  assign f_u_dadda_cla32_fa603_xor0 = f_u_dadda_cla32_and_26_20 ^ f_u_dadda_cla32_and_25_21;
  assign f_u_dadda_cla32_fa603_and0 = f_u_dadda_cla32_and_26_20 & f_u_dadda_cla32_and_25_21;
  assign f_u_dadda_cla32_fa603_xor1 = f_u_dadda_cla32_fa603_xor0 ^ f_u_dadda_cla32_and_24_22;
  assign f_u_dadda_cla32_fa603_and1 = f_u_dadda_cla32_fa603_xor0 & f_u_dadda_cla32_and_24_22;
  assign f_u_dadda_cla32_fa603_or0 = f_u_dadda_cla32_fa603_and0 | f_u_dadda_cla32_fa603_and1;
  assign f_u_dadda_cla32_and_23_23 = a[23] & b[23];
  assign f_u_dadda_cla32_and_22_24 = a[22] & b[24];
  assign f_u_dadda_cla32_and_21_25 = a[21] & b[25];
  assign f_u_dadda_cla32_fa604_xor0 = f_u_dadda_cla32_and_23_23 ^ f_u_dadda_cla32_and_22_24;
  assign f_u_dadda_cla32_fa604_and0 = f_u_dadda_cla32_and_23_23 & f_u_dadda_cla32_and_22_24;
  assign f_u_dadda_cla32_fa604_xor1 = f_u_dadda_cla32_fa604_xor0 ^ f_u_dadda_cla32_and_21_25;
  assign f_u_dadda_cla32_fa604_and1 = f_u_dadda_cla32_fa604_xor0 & f_u_dadda_cla32_and_21_25;
  assign f_u_dadda_cla32_fa604_or0 = f_u_dadda_cla32_fa604_and0 | f_u_dadda_cla32_fa604_and1;
  assign f_u_dadda_cla32_and_20_26 = a[20] & b[26];
  assign f_u_dadda_cla32_and_19_27 = a[19] & b[27];
  assign f_u_dadda_cla32_and_18_28 = a[18] & b[28];
  assign f_u_dadda_cla32_fa605_xor0 = f_u_dadda_cla32_and_20_26 ^ f_u_dadda_cla32_and_19_27;
  assign f_u_dadda_cla32_fa605_and0 = f_u_dadda_cla32_and_20_26 & f_u_dadda_cla32_and_19_27;
  assign f_u_dadda_cla32_fa605_xor1 = f_u_dadda_cla32_fa605_xor0 ^ f_u_dadda_cla32_and_18_28;
  assign f_u_dadda_cla32_fa605_and1 = f_u_dadda_cla32_fa605_xor0 & f_u_dadda_cla32_and_18_28;
  assign f_u_dadda_cla32_fa605_or0 = f_u_dadda_cla32_fa605_and0 | f_u_dadda_cla32_fa605_and1;
  assign f_u_dadda_cla32_and_17_29 = a[17] & b[29];
  assign f_u_dadda_cla32_and_16_30 = a[16] & b[30];
  assign f_u_dadda_cla32_and_15_31 = a[15] & b[31];
  assign f_u_dadda_cla32_fa606_xor0 = f_u_dadda_cla32_and_17_29 ^ f_u_dadda_cla32_and_16_30;
  assign f_u_dadda_cla32_fa606_and0 = f_u_dadda_cla32_and_17_29 & f_u_dadda_cla32_and_16_30;
  assign f_u_dadda_cla32_fa606_xor1 = f_u_dadda_cla32_fa606_xor0 ^ f_u_dadda_cla32_and_15_31;
  assign f_u_dadda_cla32_fa606_and1 = f_u_dadda_cla32_fa606_xor0 & f_u_dadda_cla32_and_15_31;
  assign f_u_dadda_cla32_fa606_or0 = f_u_dadda_cla32_fa606_and0 | f_u_dadda_cla32_fa606_and1;
  assign f_u_dadda_cla32_fa607_xor0 = f_u_dadda_cla32_fa597_xor1 ^ f_u_dadda_cla32_fa598_xor1;
  assign f_u_dadda_cla32_fa607_and0 = f_u_dadda_cla32_fa597_xor1 & f_u_dadda_cla32_fa598_xor1;
  assign f_u_dadda_cla32_fa607_xor1 = f_u_dadda_cla32_fa607_xor0 ^ f_u_dadda_cla32_fa599_xor1;
  assign f_u_dadda_cla32_fa607_and1 = f_u_dadda_cla32_fa607_xor0 & f_u_dadda_cla32_fa599_xor1;
  assign f_u_dadda_cla32_fa607_or0 = f_u_dadda_cla32_fa607_and0 | f_u_dadda_cla32_fa607_and1;
  assign f_u_dadda_cla32_fa608_xor0 = f_u_dadda_cla32_fa600_xor1 ^ f_u_dadda_cla32_fa601_xor1;
  assign f_u_dadda_cla32_fa608_and0 = f_u_dadda_cla32_fa600_xor1 & f_u_dadda_cla32_fa601_xor1;
  assign f_u_dadda_cla32_fa608_xor1 = f_u_dadda_cla32_fa608_xor0 ^ f_u_dadda_cla32_fa602_xor1;
  assign f_u_dadda_cla32_fa608_and1 = f_u_dadda_cla32_fa608_xor0 & f_u_dadda_cla32_fa602_xor1;
  assign f_u_dadda_cla32_fa608_or0 = f_u_dadda_cla32_fa608_and0 | f_u_dadda_cla32_fa608_and1;
  assign f_u_dadda_cla32_fa609_xor0 = f_u_dadda_cla32_fa608_or0 ^ f_u_dadda_cla32_fa607_or0;
  assign f_u_dadda_cla32_fa609_and0 = f_u_dadda_cla32_fa608_or0 & f_u_dadda_cla32_fa607_or0;
  assign f_u_dadda_cla32_fa609_xor1 = f_u_dadda_cla32_fa609_xor0 ^ f_u_dadda_cla32_fa606_or0;
  assign f_u_dadda_cla32_fa609_and1 = f_u_dadda_cla32_fa609_xor0 & f_u_dadda_cla32_fa606_or0;
  assign f_u_dadda_cla32_fa609_or0 = f_u_dadda_cla32_fa609_and0 | f_u_dadda_cla32_fa609_and1;
  assign f_u_dadda_cla32_fa610_xor0 = f_u_dadda_cla32_fa605_or0 ^ f_u_dadda_cla32_fa604_or0;
  assign f_u_dadda_cla32_fa610_and0 = f_u_dadda_cla32_fa605_or0 & f_u_dadda_cla32_fa604_or0;
  assign f_u_dadda_cla32_fa610_xor1 = f_u_dadda_cla32_fa610_xor0 ^ f_u_dadda_cla32_fa603_or0;
  assign f_u_dadda_cla32_fa610_and1 = f_u_dadda_cla32_fa610_xor0 & f_u_dadda_cla32_fa603_or0;
  assign f_u_dadda_cla32_fa610_or0 = f_u_dadda_cla32_fa610_and0 | f_u_dadda_cla32_fa610_and1;
  assign f_u_dadda_cla32_fa611_xor0 = f_u_dadda_cla32_fa602_or0 ^ f_u_dadda_cla32_fa601_or0;
  assign f_u_dadda_cla32_fa611_and0 = f_u_dadda_cla32_fa602_or0 & f_u_dadda_cla32_fa601_or0;
  assign f_u_dadda_cla32_fa611_xor1 = f_u_dadda_cla32_fa611_xor0 ^ f_u_dadda_cla32_fa600_or0;
  assign f_u_dadda_cla32_fa611_and1 = f_u_dadda_cla32_fa611_xor0 & f_u_dadda_cla32_fa600_or0;
  assign f_u_dadda_cla32_fa611_or0 = f_u_dadda_cla32_fa611_and0 | f_u_dadda_cla32_fa611_and1;
  assign f_u_dadda_cla32_fa612_xor0 = f_u_dadda_cla32_fa599_or0 ^ f_u_dadda_cla32_fa598_or0;
  assign f_u_dadda_cla32_fa612_and0 = f_u_dadda_cla32_fa599_or0 & f_u_dadda_cla32_fa598_or0;
  assign f_u_dadda_cla32_fa612_xor1 = f_u_dadda_cla32_fa612_xor0 ^ f_u_dadda_cla32_fa597_or0;
  assign f_u_dadda_cla32_fa612_and1 = f_u_dadda_cla32_fa612_xor0 & f_u_dadda_cla32_fa597_or0;
  assign f_u_dadda_cla32_fa612_or0 = f_u_dadda_cla32_fa612_and0 | f_u_dadda_cla32_fa612_and1;
  assign f_u_dadda_cla32_and_31_16 = a[31] & b[16];
  assign f_u_dadda_cla32_and_30_17 = a[30] & b[17];
  assign f_u_dadda_cla32_and_29_18 = a[29] & b[18];
  assign f_u_dadda_cla32_fa613_xor0 = f_u_dadda_cla32_and_31_16 ^ f_u_dadda_cla32_and_30_17;
  assign f_u_dadda_cla32_fa613_and0 = f_u_dadda_cla32_and_31_16 & f_u_dadda_cla32_and_30_17;
  assign f_u_dadda_cla32_fa613_xor1 = f_u_dadda_cla32_fa613_xor0 ^ f_u_dadda_cla32_and_29_18;
  assign f_u_dadda_cla32_fa613_and1 = f_u_dadda_cla32_fa613_xor0 & f_u_dadda_cla32_and_29_18;
  assign f_u_dadda_cla32_fa613_or0 = f_u_dadda_cla32_fa613_and0 | f_u_dadda_cla32_fa613_and1;
  assign f_u_dadda_cla32_and_28_19 = a[28] & b[19];
  assign f_u_dadda_cla32_and_27_20 = a[27] & b[20];
  assign f_u_dadda_cla32_and_26_21 = a[26] & b[21];
  assign f_u_dadda_cla32_fa614_xor0 = f_u_dadda_cla32_and_28_19 ^ f_u_dadda_cla32_and_27_20;
  assign f_u_dadda_cla32_fa614_and0 = f_u_dadda_cla32_and_28_19 & f_u_dadda_cla32_and_27_20;
  assign f_u_dadda_cla32_fa614_xor1 = f_u_dadda_cla32_fa614_xor0 ^ f_u_dadda_cla32_and_26_21;
  assign f_u_dadda_cla32_fa614_and1 = f_u_dadda_cla32_fa614_xor0 & f_u_dadda_cla32_and_26_21;
  assign f_u_dadda_cla32_fa614_or0 = f_u_dadda_cla32_fa614_and0 | f_u_dadda_cla32_fa614_and1;
  assign f_u_dadda_cla32_and_25_22 = a[25] & b[22];
  assign f_u_dadda_cla32_and_24_23 = a[24] & b[23];
  assign f_u_dadda_cla32_and_23_24 = a[23] & b[24];
  assign f_u_dadda_cla32_fa615_xor0 = f_u_dadda_cla32_and_25_22 ^ f_u_dadda_cla32_and_24_23;
  assign f_u_dadda_cla32_fa615_and0 = f_u_dadda_cla32_and_25_22 & f_u_dadda_cla32_and_24_23;
  assign f_u_dadda_cla32_fa615_xor1 = f_u_dadda_cla32_fa615_xor0 ^ f_u_dadda_cla32_and_23_24;
  assign f_u_dadda_cla32_fa615_and1 = f_u_dadda_cla32_fa615_xor0 & f_u_dadda_cla32_and_23_24;
  assign f_u_dadda_cla32_fa615_or0 = f_u_dadda_cla32_fa615_and0 | f_u_dadda_cla32_fa615_and1;
  assign f_u_dadda_cla32_and_22_25 = a[22] & b[25];
  assign f_u_dadda_cla32_and_21_26 = a[21] & b[26];
  assign f_u_dadda_cla32_and_20_27 = a[20] & b[27];
  assign f_u_dadda_cla32_fa616_xor0 = f_u_dadda_cla32_and_22_25 ^ f_u_dadda_cla32_and_21_26;
  assign f_u_dadda_cla32_fa616_and0 = f_u_dadda_cla32_and_22_25 & f_u_dadda_cla32_and_21_26;
  assign f_u_dadda_cla32_fa616_xor1 = f_u_dadda_cla32_fa616_xor0 ^ f_u_dadda_cla32_and_20_27;
  assign f_u_dadda_cla32_fa616_and1 = f_u_dadda_cla32_fa616_xor0 & f_u_dadda_cla32_and_20_27;
  assign f_u_dadda_cla32_fa616_or0 = f_u_dadda_cla32_fa616_and0 | f_u_dadda_cla32_fa616_and1;
  assign f_u_dadda_cla32_and_19_28 = a[19] & b[28];
  assign f_u_dadda_cla32_and_18_29 = a[18] & b[29];
  assign f_u_dadda_cla32_and_17_30 = a[17] & b[30];
  assign f_u_dadda_cla32_fa617_xor0 = f_u_dadda_cla32_and_19_28 ^ f_u_dadda_cla32_and_18_29;
  assign f_u_dadda_cla32_fa617_and0 = f_u_dadda_cla32_and_19_28 & f_u_dadda_cla32_and_18_29;
  assign f_u_dadda_cla32_fa617_xor1 = f_u_dadda_cla32_fa617_xor0 ^ f_u_dadda_cla32_and_17_30;
  assign f_u_dadda_cla32_fa617_and1 = f_u_dadda_cla32_fa617_xor0 & f_u_dadda_cla32_and_17_30;
  assign f_u_dadda_cla32_fa617_or0 = f_u_dadda_cla32_fa617_and0 | f_u_dadda_cla32_fa617_and1;
  assign f_u_dadda_cla32_and_16_31 = a[16] & b[31];
  assign f_u_dadda_cla32_fa618_xor0 = f_u_dadda_cla32_and_16_31 ^ f_u_dadda_cla32_fa609_xor1;
  assign f_u_dadda_cla32_fa618_and0 = f_u_dadda_cla32_and_16_31 & f_u_dadda_cla32_fa609_xor1;
  assign f_u_dadda_cla32_fa618_xor1 = f_u_dadda_cla32_fa618_xor0 ^ f_u_dadda_cla32_fa610_xor1;
  assign f_u_dadda_cla32_fa618_and1 = f_u_dadda_cla32_fa618_xor0 & f_u_dadda_cla32_fa610_xor1;
  assign f_u_dadda_cla32_fa618_or0 = f_u_dadda_cla32_fa618_and0 | f_u_dadda_cla32_fa618_and1;
  assign f_u_dadda_cla32_fa619_xor0 = f_u_dadda_cla32_fa611_xor1 ^ f_u_dadda_cla32_fa612_xor1;
  assign f_u_dadda_cla32_fa619_and0 = f_u_dadda_cla32_fa611_xor1 & f_u_dadda_cla32_fa612_xor1;
  assign f_u_dadda_cla32_fa619_xor1 = f_u_dadda_cla32_fa619_xor0 ^ f_u_dadda_cla32_fa613_xor1;
  assign f_u_dadda_cla32_fa619_and1 = f_u_dadda_cla32_fa619_xor0 & f_u_dadda_cla32_fa613_xor1;
  assign f_u_dadda_cla32_fa619_or0 = f_u_dadda_cla32_fa619_and0 | f_u_dadda_cla32_fa619_and1;
  assign f_u_dadda_cla32_fa620_xor0 = f_u_dadda_cla32_fa619_or0 ^ f_u_dadda_cla32_fa618_or0;
  assign f_u_dadda_cla32_fa620_and0 = f_u_dadda_cla32_fa619_or0 & f_u_dadda_cla32_fa618_or0;
  assign f_u_dadda_cla32_fa620_xor1 = f_u_dadda_cla32_fa620_xor0 ^ f_u_dadda_cla32_fa617_or0;
  assign f_u_dadda_cla32_fa620_and1 = f_u_dadda_cla32_fa620_xor0 & f_u_dadda_cla32_fa617_or0;
  assign f_u_dadda_cla32_fa620_or0 = f_u_dadda_cla32_fa620_and0 | f_u_dadda_cla32_fa620_and1;
  assign f_u_dadda_cla32_fa621_xor0 = f_u_dadda_cla32_fa616_or0 ^ f_u_dadda_cla32_fa615_or0;
  assign f_u_dadda_cla32_fa621_and0 = f_u_dadda_cla32_fa616_or0 & f_u_dadda_cla32_fa615_or0;
  assign f_u_dadda_cla32_fa621_xor1 = f_u_dadda_cla32_fa621_xor0 ^ f_u_dadda_cla32_fa614_or0;
  assign f_u_dadda_cla32_fa621_and1 = f_u_dadda_cla32_fa621_xor0 & f_u_dadda_cla32_fa614_or0;
  assign f_u_dadda_cla32_fa621_or0 = f_u_dadda_cla32_fa621_and0 | f_u_dadda_cla32_fa621_and1;
  assign f_u_dadda_cla32_fa622_xor0 = f_u_dadda_cla32_fa613_or0 ^ f_u_dadda_cla32_fa612_or0;
  assign f_u_dadda_cla32_fa622_and0 = f_u_dadda_cla32_fa613_or0 & f_u_dadda_cla32_fa612_or0;
  assign f_u_dadda_cla32_fa622_xor1 = f_u_dadda_cla32_fa622_xor0 ^ f_u_dadda_cla32_fa611_or0;
  assign f_u_dadda_cla32_fa622_and1 = f_u_dadda_cla32_fa622_xor0 & f_u_dadda_cla32_fa611_or0;
  assign f_u_dadda_cla32_fa622_or0 = f_u_dadda_cla32_fa622_and0 | f_u_dadda_cla32_fa622_and1;
  assign f_u_dadda_cla32_and_31_17 = a[31] & b[17];
  assign f_u_dadda_cla32_fa623_xor0 = f_u_dadda_cla32_fa610_or0 ^ f_u_dadda_cla32_fa609_or0;
  assign f_u_dadda_cla32_fa623_and0 = f_u_dadda_cla32_fa610_or0 & f_u_dadda_cla32_fa609_or0;
  assign f_u_dadda_cla32_fa623_xor1 = f_u_dadda_cla32_fa623_xor0 ^ f_u_dadda_cla32_and_31_17;
  assign f_u_dadda_cla32_fa623_and1 = f_u_dadda_cla32_fa623_xor0 & f_u_dadda_cla32_and_31_17;
  assign f_u_dadda_cla32_fa623_or0 = f_u_dadda_cla32_fa623_and0 | f_u_dadda_cla32_fa623_and1;
  assign f_u_dadda_cla32_and_30_18 = a[30] & b[18];
  assign f_u_dadda_cla32_and_29_19 = a[29] & b[19];
  assign f_u_dadda_cla32_and_28_20 = a[28] & b[20];
  assign f_u_dadda_cla32_fa624_xor0 = f_u_dadda_cla32_and_30_18 ^ f_u_dadda_cla32_and_29_19;
  assign f_u_dadda_cla32_fa624_and0 = f_u_dadda_cla32_and_30_18 & f_u_dadda_cla32_and_29_19;
  assign f_u_dadda_cla32_fa624_xor1 = f_u_dadda_cla32_fa624_xor0 ^ f_u_dadda_cla32_and_28_20;
  assign f_u_dadda_cla32_fa624_and1 = f_u_dadda_cla32_fa624_xor0 & f_u_dadda_cla32_and_28_20;
  assign f_u_dadda_cla32_fa624_or0 = f_u_dadda_cla32_fa624_and0 | f_u_dadda_cla32_fa624_and1;
  assign f_u_dadda_cla32_and_27_21 = a[27] & b[21];
  assign f_u_dadda_cla32_and_26_22 = a[26] & b[22];
  assign f_u_dadda_cla32_and_25_23 = a[25] & b[23];
  assign f_u_dadda_cla32_fa625_xor0 = f_u_dadda_cla32_and_27_21 ^ f_u_dadda_cla32_and_26_22;
  assign f_u_dadda_cla32_fa625_and0 = f_u_dadda_cla32_and_27_21 & f_u_dadda_cla32_and_26_22;
  assign f_u_dadda_cla32_fa625_xor1 = f_u_dadda_cla32_fa625_xor0 ^ f_u_dadda_cla32_and_25_23;
  assign f_u_dadda_cla32_fa625_and1 = f_u_dadda_cla32_fa625_xor0 & f_u_dadda_cla32_and_25_23;
  assign f_u_dadda_cla32_fa625_or0 = f_u_dadda_cla32_fa625_and0 | f_u_dadda_cla32_fa625_and1;
  assign f_u_dadda_cla32_and_24_24 = a[24] & b[24];
  assign f_u_dadda_cla32_and_23_25 = a[23] & b[25];
  assign f_u_dadda_cla32_and_22_26 = a[22] & b[26];
  assign f_u_dadda_cla32_fa626_xor0 = f_u_dadda_cla32_and_24_24 ^ f_u_dadda_cla32_and_23_25;
  assign f_u_dadda_cla32_fa626_and0 = f_u_dadda_cla32_and_24_24 & f_u_dadda_cla32_and_23_25;
  assign f_u_dadda_cla32_fa626_xor1 = f_u_dadda_cla32_fa626_xor0 ^ f_u_dadda_cla32_and_22_26;
  assign f_u_dadda_cla32_fa626_and1 = f_u_dadda_cla32_fa626_xor0 & f_u_dadda_cla32_and_22_26;
  assign f_u_dadda_cla32_fa626_or0 = f_u_dadda_cla32_fa626_and0 | f_u_dadda_cla32_fa626_and1;
  assign f_u_dadda_cla32_and_21_27 = a[21] & b[27];
  assign f_u_dadda_cla32_and_20_28 = a[20] & b[28];
  assign f_u_dadda_cla32_and_19_29 = a[19] & b[29];
  assign f_u_dadda_cla32_fa627_xor0 = f_u_dadda_cla32_and_21_27 ^ f_u_dadda_cla32_and_20_28;
  assign f_u_dadda_cla32_fa627_and0 = f_u_dadda_cla32_and_21_27 & f_u_dadda_cla32_and_20_28;
  assign f_u_dadda_cla32_fa627_xor1 = f_u_dadda_cla32_fa627_xor0 ^ f_u_dadda_cla32_and_19_29;
  assign f_u_dadda_cla32_fa627_and1 = f_u_dadda_cla32_fa627_xor0 & f_u_dadda_cla32_and_19_29;
  assign f_u_dadda_cla32_fa627_or0 = f_u_dadda_cla32_fa627_and0 | f_u_dadda_cla32_fa627_and1;
  assign f_u_dadda_cla32_and_18_30 = a[18] & b[30];
  assign f_u_dadda_cla32_and_17_31 = a[17] & b[31];
  assign f_u_dadda_cla32_fa628_xor0 = f_u_dadda_cla32_and_18_30 ^ f_u_dadda_cla32_and_17_31;
  assign f_u_dadda_cla32_fa628_and0 = f_u_dadda_cla32_and_18_30 & f_u_dadda_cla32_and_17_31;
  assign f_u_dadda_cla32_fa628_xor1 = f_u_dadda_cla32_fa628_xor0 ^ f_u_dadda_cla32_fa620_xor1;
  assign f_u_dadda_cla32_fa628_and1 = f_u_dadda_cla32_fa628_xor0 & f_u_dadda_cla32_fa620_xor1;
  assign f_u_dadda_cla32_fa628_or0 = f_u_dadda_cla32_fa628_and0 | f_u_dadda_cla32_fa628_and1;
  assign f_u_dadda_cla32_fa629_xor0 = f_u_dadda_cla32_fa621_xor1 ^ f_u_dadda_cla32_fa622_xor1;
  assign f_u_dadda_cla32_fa629_and0 = f_u_dadda_cla32_fa621_xor1 & f_u_dadda_cla32_fa622_xor1;
  assign f_u_dadda_cla32_fa629_xor1 = f_u_dadda_cla32_fa629_xor0 ^ f_u_dadda_cla32_fa623_xor1;
  assign f_u_dadda_cla32_fa629_and1 = f_u_dadda_cla32_fa629_xor0 & f_u_dadda_cla32_fa623_xor1;
  assign f_u_dadda_cla32_fa629_or0 = f_u_dadda_cla32_fa629_and0 | f_u_dadda_cla32_fa629_and1;
  assign f_u_dadda_cla32_fa630_xor0 = f_u_dadda_cla32_fa629_or0 ^ f_u_dadda_cla32_fa628_or0;
  assign f_u_dadda_cla32_fa630_and0 = f_u_dadda_cla32_fa629_or0 & f_u_dadda_cla32_fa628_or0;
  assign f_u_dadda_cla32_fa630_xor1 = f_u_dadda_cla32_fa630_xor0 ^ f_u_dadda_cla32_fa627_or0;
  assign f_u_dadda_cla32_fa630_and1 = f_u_dadda_cla32_fa630_xor0 & f_u_dadda_cla32_fa627_or0;
  assign f_u_dadda_cla32_fa630_or0 = f_u_dadda_cla32_fa630_and0 | f_u_dadda_cla32_fa630_and1;
  assign f_u_dadda_cla32_fa631_xor0 = f_u_dadda_cla32_fa626_or0 ^ f_u_dadda_cla32_fa625_or0;
  assign f_u_dadda_cla32_fa631_and0 = f_u_dadda_cla32_fa626_or0 & f_u_dadda_cla32_fa625_or0;
  assign f_u_dadda_cla32_fa631_xor1 = f_u_dadda_cla32_fa631_xor0 ^ f_u_dadda_cla32_fa624_or0;
  assign f_u_dadda_cla32_fa631_and1 = f_u_dadda_cla32_fa631_xor0 & f_u_dadda_cla32_fa624_or0;
  assign f_u_dadda_cla32_fa631_or0 = f_u_dadda_cla32_fa631_and0 | f_u_dadda_cla32_fa631_and1;
  assign f_u_dadda_cla32_fa632_xor0 = f_u_dadda_cla32_fa623_or0 ^ f_u_dadda_cla32_fa622_or0;
  assign f_u_dadda_cla32_fa632_and0 = f_u_dadda_cla32_fa623_or0 & f_u_dadda_cla32_fa622_or0;
  assign f_u_dadda_cla32_fa632_xor1 = f_u_dadda_cla32_fa632_xor0 ^ f_u_dadda_cla32_fa621_or0;
  assign f_u_dadda_cla32_fa632_and1 = f_u_dadda_cla32_fa632_xor0 & f_u_dadda_cla32_fa621_or0;
  assign f_u_dadda_cla32_fa632_or0 = f_u_dadda_cla32_fa632_and0 | f_u_dadda_cla32_fa632_and1;
  assign f_u_dadda_cla32_and_31_18 = a[31] & b[18];
  assign f_u_dadda_cla32_and_30_19 = a[30] & b[19];
  assign f_u_dadda_cla32_fa633_xor0 = f_u_dadda_cla32_fa620_or0 ^ f_u_dadda_cla32_and_31_18;
  assign f_u_dadda_cla32_fa633_and0 = f_u_dadda_cla32_fa620_or0 & f_u_dadda_cla32_and_31_18;
  assign f_u_dadda_cla32_fa633_xor1 = f_u_dadda_cla32_fa633_xor0 ^ f_u_dadda_cla32_and_30_19;
  assign f_u_dadda_cla32_fa633_and1 = f_u_dadda_cla32_fa633_xor0 & f_u_dadda_cla32_and_30_19;
  assign f_u_dadda_cla32_fa633_or0 = f_u_dadda_cla32_fa633_and0 | f_u_dadda_cla32_fa633_and1;
  assign f_u_dadda_cla32_and_29_20 = a[29] & b[20];
  assign f_u_dadda_cla32_and_28_21 = a[28] & b[21];
  assign f_u_dadda_cla32_and_27_22 = a[27] & b[22];
  assign f_u_dadda_cla32_fa634_xor0 = f_u_dadda_cla32_and_29_20 ^ f_u_dadda_cla32_and_28_21;
  assign f_u_dadda_cla32_fa634_and0 = f_u_dadda_cla32_and_29_20 & f_u_dadda_cla32_and_28_21;
  assign f_u_dadda_cla32_fa634_xor1 = f_u_dadda_cla32_fa634_xor0 ^ f_u_dadda_cla32_and_27_22;
  assign f_u_dadda_cla32_fa634_and1 = f_u_dadda_cla32_fa634_xor0 & f_u_dadda_cla32_and_27_22;
  assign f_u_dadda_cla32_fa634_or0 = f_u_dadda_cla32_fa634_and0 | f_u_dadda_cla32_fa634_and1;
  assign f_u_dadda_cla32_and_26_23 = a[26] & b[23];
  assign f_u_dadda_cla32_and_25_24 = a[25] & b[24];
  assign f_u_dadda_cla32_and_24_25 = a[24] & b[25];
  assign f_u_dadda_cla32_fa635_xor0 = f_u_dadda_cla32_and_26_23 ^ f_u_dadda_cla32_and_25_24;
  assign f_u_dadda_cla32_fa635_and0 = f_u_dadda_cla32_and_26_23 & f_u_dadda_cla32_and_25_24;
  assign f_u_dadda_cla32_fa635_xor1 = f_u_dadda_cla32_fa635_xor0 ^ f_u_dadda_cla32_and_24_25;
  assign f_u_dadda_cla32_fa635_and1 = f_u_dadda_cla32_fa635_xor0 & f_u_dadda_cla32_and_24_25;
  assign f_u_dadda_cla32_fa635_or0 = f_u_dadda_cla32_fa635_and0 | f_u_dadda_cla32_fa635_and1;
  assign f_u_dadda_cla32_and_23_26 = a[23] & b[26];
  assign f_u_dadda_cla32_and_22_27 = a[22] & b[27];
  assign f_u_dadda_cla32_and_21_28 = a[21] & b[28];
  assign f_u_dadda_cla32_fa636_xor0 = f_u_dadda_cla32_and_23_26 ^ f_u_dadda_cla32_and_22_27;
  assign f_u_dadda_cla32_fa636_and0 = f_u_dadda_cla32_and_23_26 & f_u_dadda_cla32_and_22_27;
  assign f_u_dadda_cla32_fa636_xor1 = f_u_dadda_cla32_fa636_xor0 ^ f_u_dadda_cla32_and_21_28;
  assign f_u_dadda_cla32_fa636_and1 = f_u_dadda_cla32_fa636_xor0 & f_u_dadda_cla32_and_21_28;
  assign f_u_dadda_cla32_fa636_or0 = f_u_dadda_cla32_fa636_and0 | f_u_dadda_cla32_fa636_and1;
  assign f_u_dadda_cla32_and_20_29 = a[20] & b[29];
  assign f_u_dadda_cla32_and_19_30 = a[19] & b[30];
  assign f_u_dadda_cla32_and_18_31 = a[18] & b[31];
  assign f_u_dadda_cla32_fa637_xor0 = f_u_dadda_cla32_and_20_29 ^ f_u_dadda_cla32_and_19_30;
  assign f_u_dadda_cla32_fa637_and0 = f_u_dadda_cla32_and_20_29 & f_u_dadda_cla32_and_19_30;
  assign f_u_dadda_cla32_fa637_xor1 = f_u_dadda_cla32_fa637_xor0 ^ f_u_dadda_cla32_and_18_31;
  assign f_u_dadda_cla32_fa637_and1 = f_u_dadda_cla32_fa637_xor0 & f_u_dadda_cla32_and_18_31;
  assign f_u_dadda_cla32_fa637_or0 = f_u_dadda_cla32_fa637_and0 | f_u_dadda_cla32_fa637_and1;
  assign f_u_dadda_cla32_fa638_xor0 = f_u_dadda_cla32_fa630_xor1 ^ f_u_dadda_cla32_fa631_xor1;
  assign f_u_dadda_cla32_fa638_and0 = f_u_dadda_cla32_fa630_xor1 & f_u_dadda_cla32_fa631_xor1;
  assign f_u_dadda_cla32_fa638_xor1 = f_u_dadda_cla32_fa638_xor0 ^ f_u_dadda_cla32_fa632_xor1;
  assign f_u_dadda_cla32_fa638_and1 = f_u_dadda_cla32_fa638_xor0 & f_u_dadda_cla32_fa632_xor1;
  assign f_u_dadda_cla32_fa638_or0 = f_u_dadda_cla32_fa638_and0 | f_u_dadda_cla32_fa638_and1;
  assign f_u_dadda_cla32_fa639_xor0 = f_u_dadda_cla32_fa638_or0 ^ f_u_dadda_cla32_fa637_or0;
  assign f_u_dadda_cla32_fa639_and0 = f_u_dadda_cla32_fa638_or0 & f_u_dadda_cla32_fa637_or0;
  assign f_u_dadda_cla32_fa639_xor1 = f_u_dadda_cla32_fa639_xor0 ^ f_u_dadda_cla32_fa636_or0;
  assign f_u_dadda_cla32_fa639_and1 = f_u_dadda_cla32_fa639_xor0 & f_u_dadda_cla32_fa636_or0;
  assign f_u_dadda_cla32_fa639_or0 = f_u_dadda_cla32_fa639_and0 | f_u_dadda_cla32_fa639_and1;
  assign f_u_dadda_cla32_fa640_xor0 = f_u_dadda_cla32_fa635_or0 ^ f_u_dadda_cla32_fa634_or0;
  assign f_u_dadda_cla32_fa640_and0 = f_u_dadda_cla32_fa635_or0 & f_u_dadda_cla32_fa634_or0;
  assign f_u_dadda_cla32_fa640_xor1 = f_u_dadda_cla32_fa640_xor0 ^ f_u_dadda_cla32_fa633_or0;
  assign f_u_dadda_cla32_fa640_and1 = f_u_dadda_cla32_fa640_xor0 & f_u_dadda_cla32_fa633_or0;
  assign f_u_dadda_cla32_fa640_or0 = f_u_dadda_cla32_fa640_and0 | f_u_dadda_cla32_fa640_and1;
  assign f_u_dadda_cla32_fa641_xor0 = f_u_dadda_cla32_fa632_or0 ^ f_u_dadda_cla32_fa631_or0;
  assign f_u_dadda_cla32_fa641_and0 = f_u_dadda_cla32_fa632_or0 & f_u_dadda_cla32_fa631_or0;
  assign f_u_dadda_cla32_fa641_xor1 = f_u_dadda_cla32_fa641_xor0 ^ f_u_dadda_cla32_fa630_or0;
  assign f_u_dadda_cla32_fa641_and1 = f_u_dadda_cla32_fa641_xor0 & f_u_dadda_cla32_fa630_or0;
  assign f_u_dadda_cla32_fa641_or0 = f_u_dadda_cla32_fa641_and0 | f_u_dadda_cla32_fa641_and1;
  assign f_u_dadda_cla32_and_31_19 = a[31] & b[19];
  assign f_u_dadda_cla32_and_30_20 = a[30] & b[20];
  assign f_u_dadda_cla32_and_29_21 = a[29] & b[21];
  assign f_u_dadda_cla32_fa642_xor0 = f_u_dadda_cla32_and_31_19 ^ f_u_dadda_cla32_and_30_20;
  assign f_u_dadda_cla32_fa642_and0 = f_u_dadda_cla32_and_31_19 & f_u_dadda_cla32_and_30_20;
  assign f_u_dadda_cla32_fa642_xor1 = f_u_dadda_cla32_fa642_xor0 ^ f_u_dadda_cla32_and_29_21;
  assign f_u_dadda_cla32_fa642_and1 = f_u_dadda_cla32_fa642_xor0 & f_u_dadda_cla32_and_29_21;
  assign f_u_dadda_cla32_fa642_or0 = f_u_dadda_cla32_fa642_and0 | f_u_dadda_cla32_fa642_and1;
  assign f_u_dadda_cla32_and_28_22 = a[28] & b[22];
  assign f_u_dadda_cla32_and_27_23 = a[27] & b[23];
  assign f_u_dadda_cla32_and_26_24 = a[26] & b[24];
  assign f_u_dadda_cla32_fa643_xor0 = f_u_dadda_cla32_and_28_22 ^ f_u_dadda_cla32_and_27_23;
  assign f_u_dadda_cla32_fa643_and0 = f_u_dadda_cla32_and_28_22 & f_u_dadda_cla32_and_27_23;
  assign f_u_dadda_cla32_fa643_xor1 = f_u_dadda_cla32_fa643_xor0 ^ f_u_dadda_cla32_and_26_24;
  assign f_u_dadda_cla32_fa643_and1 = f_u_dadda_cla32_fa643_xor0 & f_u_dadda_cla32_and_26_24;
  assign f_u_dadda_cla32_fa643_or0 = f_u_dadda_cla32_fa643_and0 | f_u_dadda_cla32_fa643_and1;
  assign f_u_dadda_cla32_and_25_25 = a[25] & b[25];
  assign f_u_dadda_cla32_and_24_26 = a[24] & b[26];
  assign f_u_dadda_cla32_and_23_27 = a[23] & b[27];
  assign f_u_dadda_cla32_fa644_xor0 = f_u_dadda_cla32_and_25_25 ^ f_u_dadda_cla32_and_24_26;
  assign f_u_dadda_cla32_fa644_and0 = f_u_dadda_cla32_and_25_25 & f_u_dadda_cla32_and_24_26;
  assign f_u_dadda_cla32_fa644_xor1 = f_u_dadda_cla32_fa644_xor0 ^ f_u_dadda_cla32_and_23_27;
  assign f_u_dadda_cla32_fa644_and1 = f_u_dadda_cla32_fa644_xor0 & f_u_dadda_cla32_and_23_27;
  assign f_u_dadda_cla32_fa644_or0 = f_u_dadda_cla32_fa644_and0 | f_u_dadda_cla32_fa644_and1;
  assign f_u_dadda_cla32_and_22_28 = a[22] & b[28];
  assign f_u_dadda_cla32_and_21_29 = a[21] & b[29];
  assign f_u_dadda_cla32_and_20_30 = a[20] & b[30];
  assign f_u_dadda_cla32_fa645_xor0 = f_u_dadda_cla32_and_22_28 ^ f_u_dadda_cla32_and_21_29;
  assign f_u_dadda_cla32_fa645_and0 = f_u_dadda_cla32_and_22_28 & f_u_dadda_cla32_and_21_29;
  assign f_u_dadda_cla32_fa645_xor1 = f_u_dadda_cla32_fa645_xor0 ^ f_u_dadda_cla32_and_20_30;
  assign f_u_dadda_cla32_fa645_and1 = f_u_dadda_cla32_fa645_xor0 & f_u_dadda_cla32_and_20_30;
  assign f_u_dadda_cla32_fa645_or0 = f_u_dadda_cla32_fa645_and0 | f_u_dadda_cla32_fa645_and1;
  assign f_u_dadda_cla32_and_19_31 = a[19] & b[31];
  assign f_u_dadda_cla32_fa646_xor0 = f_u_dadda_cla32_and_19_31 ^ f_u_dadda_cla32_fa639_xor1;
  assign f_u_dadda_cla32_fa646_and0 = f_u_dadda_cla32_and_19_31 & f_u_dadda_cla32_fa639_xor1;
  assign f_u_dadda_cla32_fa646_xor1 = f_u_dadda_cla32_fa646_xor0 ^ f_u_dadda_cla32_fa640_xor1;
  assign f_u_dadda_cla32_fa646_and1 = f_u_dadda_cla32_fa646_xor0 & f_u_dadda_cla32_fa640_xor1;
  assign f_u_dadda_cla32_fa646_or0 = f_u_dadda_cla32_fa646_and0 | f_u_dadda_cla32_fa646_and1;
  assign f_u_dadda_cla32_fa647_xor0 = f_u_dadda_cla32_fa646_or0 ^ f_u_dadda_cla32_fa645_or0;
  assign f_u_dadda_cla32_fa647_and0 = f_u_dadda_cla32_fa646_or0 & f_u_dadda_cla32_fa645_or0;
  assign f_u_dadda_cla32_fa647_xor1 = f_u_dadda_cla32_fa647_xor0 ^ f_u_dadda_cla32_fa644_or0;
  assign f_u_dadda_cla32_fa647_and1 = f_u_dadda_cla32_fa647_xor0 & f_u_dadda_cla32_fa644_or0;
  assign f_u_dadda_cla32_fa647_or0 = f_u_dadda_cla32_fa647_and0 | f_u_dadda_cla32_fa647_and1;
  assign f_u_dadda_cla32_fa648_xor0 = f_u_dadda_cla32_fa643_or0 ^ f_u_dadda_cla32_fa642_or0;
  assign f_u_dadda_cla32_fa648_and0 = f_u_dadda_cla32_fa643_or0 & f_u_dadda_cla32_fa642_or0;
  assign f_u_dadda_cla32_fa648_xor1 = f_u_dadda_cla32_fa648_xor0 ^ f_u_dadda_cla32_fa641_or0;
  assign f_u_dadda_cla32_fa648_and1 = f_u_dadda_cla32_fa648_xor0 & f_u_dadda_cla32_fa641_or0;
  assign f_u_dadda_cla32_fa648_or0 = f_u_dadda_cla32_fa648_and0 | f_u_dadda_cla32_fa648_and1;
  assign f_u_dadda_cla32_and_31_20 = a[31] & b[20];
  assign f_u_dadda_cla32_fa649_xor0 = f_u_dadda_cla32_fa640_or0 ^ f_u_dadda_cla32_fa639_or0;
  assign f_u_dadda_cla32_fa649_and0 = f_u_dadda_cla32_fa640_or0 & f_u_dadda_cla32_fa639_or0;
  assign f_u_dadda_cla32_fa649_xor1 = f_u_dadda_cla32_fa649_xor0 ^ f_u_dadda_cla32_and_31_20;
  assign f_u_dadda_cla32_fa649_and1 = f_u_dadda_cla32_fa649_xor0 & f_u_dadda_cla32_and_31_20;
  assign f_u_dadda_cla32_fa649_or0 = f_u_dadda_cla32_fa649_and0 | f_u_dadda_cla32_fa649_and1;
  assign f_u_dadda_cla32_and_30_21 = a[30] & b[21];
  assign f_u_dadda_cla32_and_29_22 = a[29] & b[22];
  assign f_u_dadda_cla32_and_28_23 = a[28] & b[23];
  assign f_u_dadda_cla32_fa650_xor0 = f_u_dadda_cla32_and_30_21 ^ f_u_dadda_cla32_and_29_22;
  assign f_u_dadda_cla32_fa650_and0 = f_u_dadda_cla32_and_30_21 & f_u_dadda_cla32_and_29_22;
  assign f_u_dadda_cla32_fa650_xor1 = f_u_dadda_cla32_fa650_xor0 ^ f_u_dadda_cla32_and_28_23;
  assign f_u_dadda_cla32_fa650_and1 = f_u_dadda_cla32_fa650_xor0 & f_u_dadda_cla32_and_28_23;
  assign f_u_dadda_cla32_fa650_or0 = f_u_dadda_cla32_fa650_and0 | f_u_dadda_cla32_fa650_and1;
  assign f_u_dadda_cla32_and_27_24 = a[27] & b[24];
  assign f_u_dadda_cla32_and_26_25 = a[26] & b[25];
  assign f_u_dadda_cla32_and_25_26 = a[25] & b[26];
  assign f_u_dadda_cla32_fa651_xor0 = f_u_dadda_cla32_and_27_24 ^ f_u_dadda_cla32_and_26_25;
  assign f_u_dadda_cla32_fa651_and0 = f_u_dadda_cla32_and_27_24 & f_u_dadda_cla32_and_26_25;
  assign f_u_dadda_cla32_fa651_xor1 = f_u_dadda_cla32_fa651_xor0 ^ f_u_dadda_cla32_and_25_26;
  assign f_u_dadda_cla32_fa651_and1 = f_u_dadda_cla32_fa651_xor0 & f_u_dadda_cla32_and_25_26;
  assign f_u_dadda_cla32_fa651_or0 = f_u_dadda_cla32_fa651_and0 | f_u_dadda_cla32_fa651_and1;
  assign f_u_dadda_cla32_and_24_27 = a[24] & b[27];
  assign f_u_dadda_cla32_and_23_28 = a[23] & b[28];
  assign f_u_dadda_cla32_and_22_29 = a[22] & b[29];
  assign f_u_dadda_cla32_fa652_xor0 = f_u_dadda_cla32_and_24_27 ^ f_u_dadda_cla32_and_23_28;
  assign f_u_dadda_cla32_fa652_and0 = f_u_dadda_cla32_and_24_27 & f_u_dadda_cla32_and_23_28;
  assign f_u_dadda_cla32_fa652_xor1 = f_u_dadda_cla32_fa652_xor0 ^ f_u_dadda_cla32_and_22_29;
  assign f_u_dadda_cla32_fa652_and1 = f_u_dadda_cla32_fa652_xor0 & f_u_dadda_cla32_and_22_29;
  assign f_u_dadda_cla32_fa652_or0 = f_u_dadda_cla32_fa652_and0 | f_u_dadda_cla32_fa652_and1;
  assign f_u_dadda_cla32_and_21_30 = a[21] & b[30];
  assign f_u_dadda_cla32_and_20_31 = a[20] & b[31];
  assign f_u_dadda_cla32_fa653_xor0 = f_u_dadda_cla32_and_21_30 ^ f_u_dadda_cla32_and_20_31;
  assign f_u_dadda_cla32_fa653_and0 = f_u_dadda_cla32_and_21_30 & f_u_dadda_cla32_and_20_31;
  assign f_u_dadda_cla32_fa653_xor1 = f_u_dadda_cla32_fa653_xor0 ^ f_u_dadda_cla32_fa647_xor1;
  assign f_u_dadda_cla32_fa653_and1 = f_u_dadda_cla32_fa653_xor0 & f_u_dadda_cla32_fa647_xor1;
  assign f_u_dadda_cla32_fa653_or0 = f_u_dadda_cla32_fa653_and0 | f_u_dadda_cla32_fa653_and1;
  assign f_u_dadda_cla32_fa654_xor0 = f_u_dadda_cla32_fa653_or0 ^ f_u_dadda_cla32_fa652_or0;
  assign f_u_dadda_cla32_fa654_and0 = f_u_dadda_cla32_fa653_or0 & f_u_dadda_cla32_fa652_or0;
  assign f_u_dadda_cla32_fa654_xor1 = f_u_dadda_cla32_fa654_xor0 ^ f_u_dadda_cla32_fa651_or0;
  assign f_u_dadda_cla32_fa654_and1 = f_u_dadda_cla32_fa654_xor0 & f_u_dadda_cla32_fa651_or0;
  assign f_u_dadda_cla32_fa654_or0 = f_u_dadda_cla32_fa654_and0 | f_u_dadda_cla32_fa654_and1;
  assign f_u_dadda_cla32_fa655_xor0 = f_u_dadda_cla32_fa650_or0 ^ f_u_dadda_cla32_fa649_or0;
  assign f_u_dadda_cla32_fa655_and0 = f_u_dadda_cla32_fa650_or0 & f_u_dadda_cla32_fa649_or0;
  assign f_u_dadda_cla32_fa655_xor1 = f_u_dadda_cla32_fa655_xor0 ^ f_u_dadda_cla32_fa648_or0;
  assign f_u_dadda_cla32_fa655_and1 = f_u_dadda_cla32_fa655_xor0 & f_u_dadda_cla32_fa648_or0;
  assign f_u_dadda_cla32_fa655_or0 = f_u_dadda_cla32_fa655_and0 | f_u_dadda_cla32_fa655_and1;
  assign f_u_dadda_cla32_and_31_21 = a[31] & b[21];
  assign f_u_dadda_cla32_and_30_22 = a[30] & b[22];
  assign f_u_dadda_cla32_fa656_xor0 = f_u_dadda_cla32_fa647_or0 ^ f_u_dadda_cla32_and_31_21;
  assign f_u_dadda_cla32_fa656_and0 = f_u_dadda_cla32_fa647_or0 & f_u_dadda_cla32_and_31_21;
  assign f_u_dadda_cla32_fa656_xor1 = f_u_dadda_cla32_fa656_xor0 ^ f_u_dadda_cla32_and_30_22;
  assign f_u_dadda_cla32_fa656_and1 = f_u_dadda_cla32_fa656_xor0 & f_u_dadda_cla32_and_30_22;
  assign f_u_dadda_cla32_fa656_or0 = f_u_dadda_cla32_fa656_and0 | f_u_dadda_cla32_fa656_and1;
  assign f_u_dadda_cla32_and_29_23 = a[29] & b[23];
  assign f_u_dadda_cla32_and_28_24 = a[28] & b[24];
  assign f_u_dadda_cla32_and_27_25 = a[27] & b[25];
  assign f_u_dadda_cla32_fa657_xor0 = f_u_dadda_cla32_and_29_23 ^ f_u_dadda_cla32_and_28_24;
  assign f_u_dadda_cla32_fa657_and0 = f_u_dadda_cla32_and_29_23 & f_u_dadda_cla32_and_28_24;
  assign f_u_dadda_cla32_fa657_xor1 = f_u_dadda_cla32_fa657_xor0 ^ f_u_dadda_cla32_and_27_25;
  assign f_u_dadda_cla32_fa657_and1 = f_u_dadda_cla32_fa657_xor0 & f_u_dadda_cla32_and_27_25;
  assign f_u_dadda_cla32_fa657_or0 = f_u_dadda_cla32_fa657_and0 | f_u_dadda_cla32_fa657_and1;
  assign f_u_dadda_cla32_and_26_26 = a[26] & b[26];
  assign f_u_dadda_cla32_and_25_27 = a[25] & b[27];
  assign f_u_dadda_cla32_and_24_28 = a[24] & b[28];
  assign f_u_dadda_cla32_fa658_xor0 = f_u_dadda_cla32_and_26_26 ^ f_u_dadda_cla32_and_25_27;
  assign f_u_dadda_cla32_fa658_and0 = f_u_dadda_cla32_and_26_26 & f_u_dadda_cla32_and_25_27;
  assign f_u_dadda_cla32_fa658_xor1 = f_u_dadda_cla32_fa658_xor0 ^ f_u_dadda_cla32_and_24_28;
  assign f_u_dadda_cla32_fa658_and1 = f_u_dadda_cla32_fa658_xor0 & f_u_dadda_cla32_and_24_28;
  assign f_u_dadda_cla32_fa658_or0 = f_u_dadda_cla32_fa658_and0 | f_u_dadda_cla32_fa658_and1;
  assign f_u_dadda_cla32_and_23_29 = a[23] & b[29];
  assign f_u_dadda_cla32_and_22_30 = a[22] & b[30];
  assign f_u_dadda_cla32_and_21_31 = a[21] & b[31];
  assign f_u_dadda_cla32_fa659_xor0 = f_u_dadda_cla32_and_23_29 ^ f_u_dadda_cla32_and_22_30;
  assign f_u_dadda_cla32_fa659_and0 = f_u_dadda_cla32_and_23_29 & f_u_dadda_cla32_and_22_30;
  assign f_u_dadda_cla32_fa659_xor1 = f_u_dadda_cla32_fa659_xor0 ^ f_u_dadda_cla32_and_21_31;
  assign f_u_dadda_cla32_fa659_and1 = f_u_dadda_cla32_fa659_xor0 & f_u_dadda_cla32_and_21_31;
  assign f_u_dadda_cla32_fa659_or0 = f_u_dadda_cla32_fa659_and0 | f_u_dadda_cla32_fa659_and1;
  assign f_u_dadda_cla32_fa660_xor0 = f_u_dadda_cla32_fa659_or0 ^ f_u_dadda_cla32_fa658_or0;
  assign f_u_dadda_cla32_fa660_and0 = f_u_dadda_cla32_fa659_or0 & f_u_dadda_cla32_fa658_or0;
  assign f_u_dadda_cla32_fa660_xor1 = f_u_dadda_cla32_fa660_xor0 ^ f_u_dadda_cla32_fa657_or0;
  assign f_u_dadda_cla32_fa660_and1 = f_u_dadda_cla32_fa660_xor0 & f_u_dadda_cla32_fa657_or0;
  assign f_u_dadda_cla32_fa660_or0 = f_u_dadda_cla32_fa660_and0 | f_u_dadda_cla32_fa660_and1;
  assign f_u_dadda_cla32_fa661_xor0 = f_u_dadda_cla32_fa656_or0 ^ f_u_dadda_cla32_fa655_or0;
  assign f_u_dadda_cla32_fa661_and0 = f_u_dadda_cla32_fa656_or0 & f_u_dadda_cla32_fa655_or0;
  assign f_u_dadda_cla32_fa661_xor1 = f_u_dadda_cla32_fa661_xor0 ^ f_u_dadda_cla32_fa654_or0;
  assign f_u_dadda_cla32_fa661_and1 = f_u_dadda_cla32_fa661_xor0 & f_u_dadda_cla32_fa654_or0;
  assign f_u_dadda_cla32_fa661_or0 = f_u_dadda_cla32_fa661_and0 | f_u_dadda_cla32_fa661_and1;
  assign f_u_dadda_cla32_and_31_22 = a[31] & b[22];
  assign f_u_dadda_cla32_and_30_23 = a[30] & b[23];
  assign f_u_dadda_cla32_and_29_24 = a[29] & b[24];
  assign f_u_dadda_cla32_fa662_xor0 = f_u_dadda_cla32_and_31_22 ^ f_u_dadda_cla32_and_30_23;
  assign f_u_dadda_cla32_fa662_and0 = f_u_dadda_cla32_and_31_22 & f_u_dadda_cla32_and_30_23;
  assign f_u_dadda_cla32_fa662_xor1 = f_u_dadda_cla32_fa662_xor0 ^ f_u_dadda_cla32_and_29_24;
  assign f_u_dadda_cla32_fa662_and1 = f_u_dadda_cla32_fa662_xor0 & f_u_dadda_cla32_and_29_24;
  assign f_u_dadda_cla32_fa662_or0 = f_u_dadda_cla32_fa662_and0 | f_u_dadda_cla32_fa662_and1;
  assign f_u_dadda_cla32_and_28_25 = a[28] & b[25];
  assign f_u_dadda_cla32_and_27_26 = a[27] & b[26];
  assign f_u_dadda_cla32_and_26_27 = a[26] & b[27];
  assign f_u_dadda_cla32_fa663_xor0 = f_u_dadda_cla32_and_28_25 ^ f_u_dadda_cla32_and_27_26;
  assign f_u_dadda_cla32_fa663_and0 = f_u_dadda_cla32_and_28_25 & f_u_dadda_cla32_and_27_26;
  assign f_u_dadda_cla32_fa663_xor1 = f_u_dadda_cla32_fa663_xor0 ^ f_u_dadda_cla32_and_26_27;
  assign f_u_dadda_cla32_fa663_and1 = f_u_dadda_cla32_fa663_xor0 & f_u_dadda_cla32_and_26_27;
  assign f_u_dadda_cla32_fa663_or0 = f_u_dadda_cla32_fa663_and0 | f_u_dadda_cla32_fa663_and1;
  assign f_u_dadda_cla32_and_25_28 = a[25] & b[28];
  assign f_u_dadda_cla32_and_24_29 = a[24] & b[29];
  assign f_u_dadda_cla32_and_23_30 = a[23] & b[30];
  assign f_u_dadda_cla32_fa664_xor0 = f_u_dadda_cla32_and_25_28 ^ f_u_dadda_cla32_and_24_29;
  assign f_u_dadda_cla32_fa664_and0 = f_u_dadda_cla32_and_25_28 & f_u_dadda_cla32_and_24_29;
  assign f_u_dadda_cla32_fa664_xor1 = f_u_dadda_cla32_fa664_xor0 ^ f_u_dadda_cla32_and_23_30;
  assign f_u_dadda_cla32_fa664_and1 = f_u_dadda_cla32_fa664_xor0 & f_u_dadda_cla32_and_23_30;
  assign f_u_dadda_cla32_fa664_or0 = f_u_dadda_cla32_fa664_and0 | f_u_dadda_cla32_fa664_and1;
  assign f_u_dadda_cla32_fa665_xor0 = f_u_dadda_cla32_fa664_or0 ^ f_u_dadda_cla32_fa663_or0;
  assign f_u_dadda_cla32_fa665_and0 = f_u_dadda_cla32_fa664_or0 & f_u_dadda_cla32_fa663_or0;
  assign f_u_dadda_cla32_fa665_xor1 = f_u_dadda_cla32_fa665_xor0 ^ f_u_dadda_cla32_fa662_or0;
  assign f_u_dadda_cla32_fa665_and1 = f_u_dadda_cla32_fa665_xor0 & f_u_dadda_cla32_fa662_or0;
  assign f_u_dadda_cla32_fa665_or0 = f_u_dadda_cla32_fa665_and0 | f_u_dadda_cla32_fa665_and1;
  assign f_u_dadda_cla32_and_31_23 = a[31] & b[23];
  assign f_u_dadda_cla32_fa666_xor0 = f_u_dadda_cla32_fa661_or0 ^ f_u_dadda_cla32_fa660_or0;
  assign f_u_dadda_cla32_fa666_and0 = f_u_dadda_cla32_fa661_or0 & f_u_dadda_cla32_fa660_or0;
  assign f_u_dadda_cla32_fa666_xor1 = f_u_dadda_cla32_fa666_xor0 ^ f_u_dadda_cla32_and_31_23;
  assign f_u_dadda_cla32_fa666_and1 = f_u_dadda_cla32_fa666_xor0 & f_u_dadda_cla32_and_31_23;
  assign f_u_dadda_cla32_fa666_or0 = f_u_dadda_cla32_fa666_and0 | f_u_dadda_cla32_fa666_and1;
  assign f_u_dadda_cla32_and_30_24 = a[30] & b[24];
  assign f_u_dadda_cla32_and_29_25 = a[29] & b[25];
  assign f_u_dadda_cla32_and_28_26 = a[28] & b[26];
  assign f_u_dadda_cla32_fa667_xor0 = f_u_dadda_cla32_and_30_24 ^ f_u_dadda_cla32_and_29_25;
  assign f_u_dadda_cla32_fa667_and0 = f_u_dadda_cla32_and_30_24 & f_u_dadda_cla32_and_29_25;
  assign f_u_dadda_cla32_fa667_xor1 = f_u_dadda_cla32_fa667_xor0 ^ f_u_dadda_cla32_and_28_26;
  assign f_u_dadda_cla32_fa667_and1 = f_u_dadda_cla32_fa667_xor0 & f_u_dadda_cla32_and_28_26;
  assign f_u_dadda_cla32_fa667_or0 = f_u_dadda_cla32_fa667_and0 | f_u_dadda_cla32_fa667_and1;
  assign f_u_dadda_cla32_and_27_27 = a[27] & b[27];
  assign f_u_dadda_cla32_and_26_28 = a[26] & b[28];
  assign f_u_dadda_cla32_and_25_29 = a[25] & b[29];
  assign f_u_dadda_cla32_fa668_xor0 = f_u_dadda_cla32_and_27_27 ^ f_u_dadda_cla32_and_26_28;
  assign f_u_dadda_cla32_fa668_and0 = f_u_dadda_cla32_and_27_27 & f_u_dadda_cla32_and_26_28;
  assign f_u_dadda_cla32_fa668_xor1 = f_u_dadda_cla32_fa668_xor0 ^ f_u_dadda_cla32_and_25_29;
  assign f_u_dadda_cla32_fa668_and1 = f_u_dadda_cla32_fa668_xor0 & f_u_dadda_cla32_and_25_29;
  assign f_u_dadda_cla32_fa668_or0 = f_u_dadda_cla32_fa668_and0 | f_u_dadda_cla32_fa668_and1;
  assign f_u_dadda_cla32_fa669_xor0 = f_u_dadda_cla32_fa668_or0 ^ f_u_dadda_cla32_fa667_or0;
  assign f_u_dadda_cla32_fa669_and0 = f_u_dadda_cla32_fa668_or0 & f_u_dadda_cla32_fa667_or0;
  assign f_u_dadda_cla32_fa669_xor1 = f_u_dadda_cla32_fa669_xor0 ^ f_u_dadda_cla32_fa666_or0;
  assign f_u_dadda_cla32_fa669_and1 = f_u_dadda_cla32_fa669_xor0 & f_u_dadda_cla32_fa666_or0;
  assign f_u_dadda_cla32_fa669_or0 = f_u_dadda_cla32_fa669_and0 | f_u_dadda_cla32_fa669_and1;
  assign f_u_dadda_cla32_and_31_24 = a[31] & b[24];
  assign f_u_dadda_cla32_and_30_25 = a[30] & b[25];
  assign f_u_dadda_cla32_fa670_xor0 = f_u_dadda_cla32_fa665_or0 ^ f_u_dadda_cla32_and_31_24;
  assign f_u_dadda_cla32_fa670_and0 = f_u_dadda_cla32_fa665_or0 & f_u_dadda_cla32_and_31_24;
  assign f_u_dadda_cla32_fa670_xor1 = f_u_dadda_cla32_fa670_xor0 ^ f_u_dadda_cla32_and_30_25;
  assign f_u_dadda_cla32_fa670_and1 = f_u_dadda_cla32_fa670_xor0 & f_u_dadda_cla32_and_30_25;
  assign f_u_dadda_cla32_fa670_or0 = f_u_dadda_cla32_fa670_and0 | f_u_dadda_cla32_fa670_and1;
  assign f_u_dadda_cla32_and_29_26 = a[29] & b[26];
  assign f_u_dadda_cla32_and_28_27 = a[28] & b[27];
  assign f_u_dadda_cla32_and_27_28 = a[27] & b[28];
  assign f_u_dadda_cla32_fa671_xor0 = f_u_dadda_cla32_and_29_26 ^ f_u_dadda_cla32_and_28_27;
  assign f_u_dadda_cla32_fa671_and0 = f_u_dadda_cla32_and_29_26 & f_u_dadda_cla32_and_28_27;
  assign f_u_dadda_cla32_fa671_xor1 = f_u_dadda_cla32_fa671_xor0 ^ f_u_dadda_cla32_and_27_28;
  assign f_u_dadda_cla32_fa671_and1 = f_u_dadda_cla32_fa671_xor0 & f_u_dadda_cla32_and_27_28;
  assign f_u_dadda_cla32_fa671_or0 = f_u_dadda_cla32_fa671_and0 | f_u_dadda_cla32_fa671_and1;
  assign f_u_dadda_cla32_fa672_xor0 = f_u_dadda_cla32_fa671_or0 ^ f_u_dadda_cla32_fa670_or0;
  assign f_u_dadda_cla32_fa672_and0 = f_u_dadda_cla32_fa671_or0 & f_u_dadda_cla32_fa670_or0;
  assign f_u_dadda_cla32_fa672_xor1 = f_u_dadda_cla32_fa672_xor0 ^ f_u_dadda_cla32_fa669_or0;
  assign f_u_dadda_cla32_fa672_and1 = f_u_dadda_cla32_fa672_xor0 & f_u_dadda_cla32_fa669_or0;
  assign f_u_dadda_cla32_fa672_or0 = f_u_dadda_cla32_fa672_and0 | f_u_dadda_cla32_fa672_and1;
  assign f_u_dadda_cla32_and_31_25 = a[31] & b[25];
  assign f_u_dadda_cla32_and_30_26 = a[30] & b[26];
  assign f_u_dadda_cla32_and_29_27 = a[29] & b[27];
  assign f_u_dadda_cla32_fa673_xor0 = f_u_dadda_cla32_and_31_25 ^ f_u_dadda_cla32_and_30_26;
  assign f_u_dadda_cla32_fa673_and0 = f_u_dadda_cla32_and_31_25 & f_u_dadda_cla32_and_30_26;
  assign f_u_dadda_cla32_fa673_xor1 = f_u_dadda_cla32_fa673_xor0 ^ f_u_dadda_cla32_and_29_27;
  assign f_u_dadda_cla32_fa673_and1 = f_u_dadda_cla32_fa673_xor0 & f_u_dadda_cla32_and_29_27;
  assign f_u_dadda_cla32_fa673_or0 = f_u_dadda_cla32_fa673_and0 | f_u_dadda_cla32_fa673_and1;
  assign f_u_dadda_cla32_and_31_26 = a[31] & b[26];
  assign f_u_dadda_cla32_fa674_xor0 = f_u_dadda_cla32_fa673_or0 ^ f_u_dadda_cla32_fa672_or0;
  assign f_u_dadda_cla32_fa674_and0 = f_u_dadda_cla32_fa673_or0 & f_u_dadda_cla32_fa672_or0;
  assign f_u_dadda_cla32_fa674_xor1 = f_u_dadda_cla32_fa674_xor0 ^ f_u_dadda_cla32_and_31_26;
  assign f_u_dadda_cla32_fa674_and1 = f_u_dadda_cla32_fa674_xor0 & f_u_dadda_cla32_and_31_26;
  assign f_u_dadda_cla32_fa674_or0 = f_u_dadda_cla32_fa674_and0 | f_u_dadda_cla32_fa674_and1;
  assign f_u_dadda_cla32_and_4_0 = a[4] & b[0];
  assign f_u_dadda_cla32_and_3_1 = a[3] & b[1];
  assign f_u_dadda_cla32_ha27_xor0 = f_u_dadda_cla32_and_4_0 ^ f_u_dadda_cla32_and_3_1;
  assign f_u_dadda_cla32_ha27_and0 = f_u_dadda_cla32_and_4_0 & f_u_dadda_cla32_and_3_1;
  assign f_u_dadda_cla32_and_5_0 = a[5] & b[0];
  assign f_u_dadda_cla32_and_4_1 = a[4] & b[1];
  assign f_u_dadda_cla32_fa675_xor0 = f_u_dadda_cla32_ha27_and0 ^ f_u_dadda_cla32_and_5_0;
  assign f_u_dadda_cla32_fa675_and0 = f_u_dadda_cla32_ha27_and0 & f_u_dadda_cla32_and_5_0;
  assign f_u_dadda_cla32_fa675_xor1 = f_u_dadda_cla32_fa675_xor0 ^ f_u_dadda_cla32_and_4_1;
  assign f_u_dadda_cla32_fa675_and1 = f_u_dadda_cla32_fa675_xor0 & f_u_dadda_cla32_and_4_1;
  assign f_u_dadda_cla32_fa675_or0 = f_u_dadda_cla32_fa675_and0 | f_u_dadda_cla32_fa675_and1;
  assign f_u_dadda_cla32_and_3_2 = a[3] & b[2];
  assign f_u_dadda_cla32_and_2_3 = a[2] & b[3];
  assign f_u_dadda_cla32_ha28_xor0 = f_u_dadda_cla32_and_3_2 ^ f_u_dadda_cla32_and_2_3;
  assign f_u_dadda_cla32_ha28_and0 = f_u_dadda_cla32_and_3_2 & f_u_dadda_cla32_and_2_3;
  assign f_u_dadda_cla32_and_4_2 = a[4] & b[2];
  assign f_u_dadda_cla32_fa676_xor0 = f_u_dadda_cla32_ha28_and0 ^ f_u_dadda_cla32_fa675_or0;
  assign f_u_dadda_cla32_fa676_and0 = f_u_dadda_cla32_ha28_and0 & f_u_dadda_cla32_fa675_or0;
  assign f_u_dadda_cla32_fa676_xor1 = f_u_dadda_cla32_fa676_xor0 ^ f_u_dadda_cla32_and_4_2;
  assign f_u_dadda_cla32_fa676_and1 = f_u_dadda_cla32_fa676_xor0 & f_u_dadda_cla32_and_4_2;
  assign f_u_dadda_cla32_fa676_or0 = f_u_dadda_cla32_fa676_and0 | f_u_dadda_cla32_fa676_and1;
  assign f_u_dadda_cla32_and_3_3 = a[3] & b[3];
  assign f_u_dadda_cla32_and_2_4 = a[2] & b[4];
  assign f_u_dadda_cla32_and_1_5 = a[1] & b[5];
  assign f_u_dadda_cla32_fa677_xor0 = f_u_dadda_cla32_and_3_3 ^ f_u_dadda_cla32_and_2_4;
  assign f_u_dadda_cla32_fa677_and0 = f_u_dadda_cla32_and_3_3 & f_u_dadda_cla32_and_2_4;
  assign f_u_dadda_cla32_fa677_xor1 = f_u_dadda_cla32_fa677_xor0 ^ f_u_dadda_cla32_and_1_5;
  assign f_u_dadda_cla32_fa677_and1 = f_u_dadda_cla32_fa677_xor0 & f_u_dadda_cla32_and_1_5;
  assign f_u_dadda_cla32_fa677_or0 = f_u_dadda_cla32_fa677_and0 | f_u_dadda_cla32_fa677_and1;
  assign f_u_dadda_cla32_and_3_4 = a[3] & b[4];
  assign f_u_dadda_cla32_fa678_xor0 = f_u_dadda_cla32_fa677_or0 ^ f_u_dadda_cla32_fa676_or0;
  assign f_u_dadda_cla32_fa678_and0 = f_u_dadda_cla32_fa677_or0 & f_u_dadda_cla32_fa676_or0;
  assign f_u_dadda_cla32_fa678_xor1 = f_u_dadda_cla32_fa678_xor0 ^ f_u_dadda_cla32_and_3_4;
  assign f_u_dadda_cla32_fa678_and1 = f_u_dadda_cla32_fa678_xor0 & f_u_dadda_cla32_and_3_4;
  assign f_u_dadda_cla32_fa678_or0 = f_u_dadda_cla32_fa678_and0 | f_u_dadda_cla32_fa678_and1;
  assign f_u_dadda_cla32_and_2_5 = a[2] & b[5];
  assign f_u_dadda_cla32_and_1_6 = a[1] & b[6];
  assign f_u_dadda_cla32_and_0_7 = a[0] & b[7];
  assign f_u_dadda_cla32_fa679_xor0 = f_u_dadda_cla32_and_2_5 ^ f_u_dadda_cla32_and_1_6;
  assign f_u_dadda_cla32_fa679_and0 = f_u_dadda_cla32_and_2_5 & f_u_dadda_cla32_and_1_6;
  assign f_u_dadda_cla32_fa679_xor1 = f_u_dadda_cla32_fa679_xor0 ^ f_u_dadda_cla32_and_0_7;
  assign f_u_dadda_cla32_fa679_and1 = f_u_dadda_cla32_fa679_xor0 & f_u_dadda_cla32_and_0_7;
  assign f_u_dadda_cla32_fa679_or0 = f_u_dadda_cla32_fa679_and0 | f_u_dadda_cla32_fa679_and1;
  assign f_u_dadda_cla32_and_2_6 = a[2] & b[6];
  assign f_u_dadda_cla32_fa680_xor0 = f_u_dadda_cla32_fa679_or0 ^ f_u_dadda_cla32_fa678_or0;
  assign f_u_dadda_cla32_fa680_and0 = f_u_dadda_cla32_fa679_or0 & f_u_dadda_cla32_fa678_or0;
  assign f_u_dadda_cla32_fa680_xor1 = f_u_dadda_cla32_fa680_xor0 ^ f_u_dadda_cla32_and_2_6;
  assign f_u_dadda_cla32_fa680_and1 = f_u_dadda_cla32_fa680_xor0 & f_u_dadda_cla32_and_2_6;
  assign f_u_dadda_cla32_fa680_or0 = f_u_dadda_cla32_fa680_and0 | f_u_dadda_cla32_fa680_and1;
  assign f_u_dadda_cla32_and_1_7 = a[1] & b[7];
  assign f_u_dadda_cla32_and_0_8 = a[0] & b[8];
  assign f_u_dadda_cla32_fa681_xor0 = f_u_dadda_cla32_and_1_7 ^ f_u_dadda_cla32_and_0_8;
  assign f_u_dadda_cla32_fa681_and0 = f_u_dadda_cla32_and_1_7 & f_u_dadda_cla32_and_0_8;
  assign f_u_dadda_cla32_fa681_xor1 = f_u_dadda_cla32_fa681_xor0 ^ f_u_dadda_cla32_fa16_xor1;
  assign f_u_dadda_cla32_fa681_and1 = f_u_dadda_cla32_fa681_xor0 & f_u_dadda_cla32_fa16_xor1;
  assign f_u_dadda_cla32_fa681_or0 = f_u_dadda_cla32_fa681_and0 | f_u_dadda_cla32_fa681_and1;
  assign f_u_dadda_cla32_and_1_8 = a[1] & b[8];
  assign f_u_dadda_cla32_fa682_xor0 = f_u_dadda_cla32_fa681_or0 ^ f_u_dadda_cla32_fa680_or0;
  assign f_u_dadda_cla32_fa682_and0 = f_u_dadda_cla32_fa681_or0 & f_u_dadda_cla32_fa680_or0;
  assign f_u_dadda_cla32_fa682_xor1 = f_u_dadda_cla32_fa682_xor0 ^ f_u_dadda_cla32_and_1_8;
  assign f_u_dadda_cla32_fa682_and1 = f_u_dadda_cla32_fa682_xor0 & f_u_dadda_cla32_and_1_8;
  assign f_u_dadda_cla32_fa682_or0 = f_u_dadda_cla32_fa682_and0 | f_u_dadda_cla32_fa682_and1;
  assign f_u_dadda_cla32_and_0_9 = a[0] & b[9];
  assign f_u_dadda_cla32_fa683_xor0 = f_u_dadda_cla32_and_0_9 ^ f_u_dadda_cla32_fa18_xor1;
  assign f_u_dadda_cla32_fa683_and0 = f_u_dadda_cla32_and_0_9 & f_u_dadda_cla32_fa18_xor1;
  assign f_u_dadda_cla32_fa683_xor1 = f_u_dadda_cla32_fa683_xor0 ^ f_u_dadda_cla32_fa19_xor1;
  assign f_u_dadda_cla32_fa683_and1 = f_u_dadda_cla32_fa683_xor0 & f_u_dadda_cla32_fa19_xor1;
  assign f_u_dadda_cla32_fa683_or0 = f_u_dadda_cla32_fa683_and0 | f_u_dadda_cla32_fa683_and1;
  assign f_u_dadda_cla32_and_0_10 = a[0] & b[10];
  assign f_u_dadda_cla32_fa684_xor0 = f_u_dadda_cla32_fa683_or0 ^ f_u_dadda_cla32_fa682_or0;
  assign f_u_dadda_cla32_fa684_and0 = f_u_dadda_cla32_fa683_or0 & f_u_dadda_cla32_fa682_or0;
  assign f_u_dadda_cla32_fa684_xor1 = f_u_dadda_cla32_fa684_xor0 ^ f_u_dadda_cla32_and_0_10;
  assign f_u_dadda_cla32_fa684_and1 = f_u_dadda_cla32_fa684_xor0 & f_u_dadda_cla32_and_0_10;
  assign f_u_dadda_cla32_fa684_or0 = f_u_dadda_cla32_fa684_and0 | f_u_dadda_cla32_fa684_and1;
  assign f_u_dadda_cla32_fa685_xor0 = f_u_dadda_cla32_fa21_xor1 ^ f_u_dadda_cla32_fa22_xor1;
  assign f_u_dadda_cla32_fa685_and0 = f_u_dadda_cla32_fa21_xor1 & f_u_dadda_cla32_fa22_xor1;
  assign f_u_dadda_cla32_fa685_xor1 = f_u_dadda_cla32_fa685_xor0 ^ f_u_dadda_cla32_fa23_xor1;
  assign f_u_dadda_cla32_fa685_and1 = f_u_dadda_cla32_fa685_xor0 & f_u_dadda_cla32_fa23_xor1;
  assign f_u_dadda_cla32_fa685_or0 = f_u_dadda_cla32_fa685_and0 | f_u_dadda_cla32_fa685_and1;
  assign f_u_dadda_cla32_fa686_xor0 = f_u_dadda_cla32_fa685_or0 ^ f_u_dadda_cla32_fa684_or0;
  assign f_u_dadda_cla32_fa686_and0 = f_u_dadda_cla32_fa685_or0 & f_u_dadda_cla32_fa684_or0;
  assign f_u_dadda_cla32_fa686_xor1 = f_u_dadda_cla32_fa686_xor0 ^ f_u_dadda_cla32_fa25_xor1;
  assign f_u_dadda_cla32_fa686_and1 = f_u_dadda_cla32_fa686_xor0 & f_u_dadda_cla32_fa25_xor1;
  assign f_u_dadda_cla32_fa686_or0 = f_u_dadda_cla32_fa686_and0 | f_u_dadda_cla32_fa686_and1;
  assign f_u_dadda_cla32_fa687_xor0 = f_u_dadda_cla32_fa26_xor1 ^ f_u_dadda_cla32_fa27_xor1;
  assign f_u_dadda_cla32_fa687_and0 = f_u_dadda_cla32_fa26_xor1 & f_u_dadda_cla32_fa27_xor1;
  assign f_u_dadda_cla32_fa687_xor1 = f_u_dadda_cla32_fa687_xor0 ^ f_u_dadda_cla32_fa28_xor1;
  assign f_u_dadda_cla32_fa687_and1 = f_u_dadda_cla32_fa687_xor0 & f_u_dadda_cla32_fa28_xor1;
  assign f_u_dadda_cla32_fa687_or0 = f_u_dadda_cla32_fa687_and0 | f_u_dadda_cla32_fa687_and1;
  assign f_u_dadda_cla32_fa688_xor0 = f_u_dadda_cla32_fa687_or0 ^ f_u_dadda_cla32_fa686_or0;
  assign f_u_dadda_cla32_fa688_and0 = f_u_dadda_cla32_fa687_or0 & f_u_dadda_cla32_fa686_or0;
  assign f_u_dadda_cla32_fa688_xor1 = f_u_dadda_cla32_fa688_xor0 ^ f_u_dadda_cla32_fa31_xor1;
  assign f_u_dadda_cla32_fa688_and1 = f_u_dadda_cla32_fa688_xor0 & f_u_dadda_cla32_fa31_xor1;
  assign f_u_dadda_cla32_fa688_or0 = f_u_dadda_cla32_fa688_and0 | f_u_dadda_cla32_fa688_and1;
  assign f_u_dadda_cla32_fa689_xor0 = f_u_dadda_cla32_fa32_xor1 ^ f_u_dadda_cla32_fa33_xor1;
  assign f_u_dadda_cla32_fa689_and0 = f_u_dadda_cla32_fa32_xor1 & f_u_dadda_cla32_fa33_xor1;
  assign f_u_dadda_cla32_fa689_xor1 = f_u_dadda_cla32_fa689_xor0 ^ f_u_dadda_cla32_fa34_xor1;
  assign f_u_dadda_cla32_fa689_and1 = f_u_dadda_cla32_fa689_xor0 & f_u_dadda_cla32_fa34_xor1;
  assign f_u_dadda_cla32_fa689_or0 = f_u_dadda_cla32_fa689_and0 | f_u_dadda_cla32_fa689_and1;
  assign f_u_dadda_cla32_fa690_xor0 = f_u_dadda_cla32_fa689_or0 ^ f_u_dadda_cla32_fa688_or0;
  assign f_u_dadda_cla32_fa690_and0 = f_u_dadda_cla32_fa689_or0 & f_u_dadda_cla32_fa688_or0;
  assign f_u_dadda_cla32_fa690_xor1 = f_u_dadda_cla32_fa690_xor0 ^ f_u_dadda_cla32_fa38_xor1;
  assign f_u_dadda_cla32_fa690_and1 = f_u_dadda_cla32_fa690_xor0 & f_u_dadda_cla32_fa38_xor1;
  assign f_u_dadda_cla32_fa690_or0 = f_u_dadda_cla32_fa690_and0 | f_u_dadda_cla32_fa690_and1;
  assign f_u_dadda_cla32_fa691_xor0 = f_u_dadda_cla32_fa39_xor1 ^ f_u_dadda_cla32_fa40_xor1;
  assign f_u_dadda_cla32_fa691_and0 = f_u_dadda_cla32_fa39_xor1 & f_u_dadda_cla32_fa40_xor1;
  assign f_u_dadda_cla32_fa691_xor1 = f_u_dadda_cla32_fa691_xor0 ^ f_u_dadda_cla32_fa41_xor1;
  assign f_u_dadda_cla32_fa691_and1 = f_u_dadda_cla32_fa691_xor0 & f_u_dadda_cla32_fa41_xor1;
  assign f_u_dadda_cla32_fa691_or0 = f_u_dadda_cla32_fa691_and0 | f_u_dadda_cla32_fa691_and1;
  assign f_u_dadda_cla32_fa692_xor0 = f_u_dadda_cla32_fa691_or0 ^ f_u_dadda_cla32_fa690_or0;
  assign f_u_dadda_cla32_fa692_and0 = f_u_dadda_cla32_fa691_or0 & f_u_dadda_cla32_fa690_or0;
  assign f_u_dadda_cla32_fa692_xor1 = f_u_dadda_cla32_fa692_xor0 ^ f_u_dadda_cla32_fa46_xor1;
  assign f_u_dadda_cla32_fa692_and1 = f_u_dadda_cla32_fa692_xor0 & f_u_dadda_cla32_fa46_xor1;
  assign f_u_dadda_cla32_fa692_or0 = f_u_dadda_cla32_fa692_and0 | f_u_dadda_cla32_fa692_and1;
  assign f_u_dadda_cla32_fa693_xor0 = f_u_dadda_cla32_fa47_xor1 ^ f_u_dadda_cla32_fa48_xor1;
  assign f_u_dadda_cla32_fa693_and0 = f_u_dadda_cla32_fa47_xor1 & f_u_dadda_cla32_fa48_xor1;
  assign f_u_dadda_cla32_fa693_xor1 = f_u_dadda_cla32_fa693_xor0 ^ f_u_dadda_cla32_fa49_xor1;
  assign f_u_dadda_cla32_fa693_and1 = f_u_dadda_cla32_fa693_xor0 & f_u_dadda_cla32_fa49_xor1;
  assign f_u_dadda_cla32_fa693_or0 = f_u_dadda_cla32_fa693_and0 | f_u_dadda_cla32_fa693_and1;
  assign f_u_dadda_cla32_fa694_xor0 = f_u_dadda_cla32_fa693_or0 ^ f_u_dadda_cla32_fa692_or0;
  assign f_u_dadda_cla32_fa694_and0 = f_u_dadda_cla32_fa693_or0 & f_u_dadda_cla32_fa692_or0;
  assign f_u_dadda_cla32_fa694_xor1 = f_u_dadda_cla32_fa694_xor0 ^ f_u_dadda_cla32_fa55_xor1;
  assign f_u_dadda_cla32_fa694_and1 = f_u_dadda_cla32_fa694_xor0 & f_u_dadda_cla32_fa55_xor1;
  assign f_u_dadda_cla32_fa694_or0 = f_u_dadda_cla32_fa694_and0 | f_u_dadda_cla32_fa694_and1;
  assign f_u_dadda_cla32_fa695_xor0 = f_u_dadda_cla32_fa56_xor1 ^ f_u_dadda_cla32_fa57_xor1;
  assign f_u_dadda_cla32_fa695_and0 = f_u_dadda_cla32_fa56_xor1 & f_u_dadda_cla32_fa57_xor1;
  assign f_u_dadda_cla32_fa695_xor1 = f_u_dadda_cla32_fa695_xor0 ^ f_u_dadda_cla32_fa58_xor1;
  assign f_u_dadda_cla32_fa695_and1 = f_u_dadda_cla32_fa695_xor0 & f_u_dadda_cla32_fa58_xor1;
  assign f_u_dadda_cla32_fa695_or0 = f_u_dadda_cla32_fa695_and0 | f_u_dadda_cla32_fa695_and1;
  assign f_u_dadda_cla32_fa696_xor0 = f_u_dadda_cla32_fa695_or0 ^ f_u_dadda_cla32_fa694_or0;
  assign f_u_dadda_cla32_fa696_and0 = f_u_dadda_cla32_fa695_or0 & f_u_dadda_cla32_fa694_or0;
  assign f_u_dadda_cla32_fa696_xor1 = f_u_dadda_cla32_fa696_xor0 ^ f_u_dadda_cla32_fa65_xor1;
  assign f_u_dadda_cla32_fa696_and1 = f_u_dadda_cla32_fa696_xor0 & f_u_dadda_cla32_fa65_xor1;
  assign f_u_dadda_cla32_fa696_or0 = f_u_dadda_cla32_fa696_and0 | f_u_dadda_cla32_fa696_and1;
  assign f_u_dadda_cla32_fa697_xor0 = f_u_dadda_cla32_fa66_xor1 ^ f_u_dadda_cla32_fa67_xor1;
  assign f_u_dadda_cla32_fa697_and0 = f_u_dadda_cla32_fa66_xor1 & f_u_dadda_cla32_fa67_xor1;
  assign f_u_dadda_cla32_fa697_xor1 = f_u_dadda_cla32_fa697_xor0 ^ f_u_dadda_cla32_fa68_xor1;
  assign f_u_dadda_cla32_fa697_and1 = f_u_dadda_cla32_fa697_xor0 & f_u_dadda_cla32_fa68_xor1;
  assign f_u_dadda_cla32_fa697_or0 = f_u_dadda_cla32_fa697_and0 | f_u_dadda_cla32_fa697_and1;
  assign f_u_dadda_cla32_fa698_xor0 = f_u_dadda_cla32_fa697_or0 ^ f_u_dadda_cla32_fa696_or0;
  assign f_u_dadda_cla32_fa698_and0 = f_u_dadda_cla32_fa697_or0 & f_u_dadda_cla32_fa696_or0;
  assign f_u_dadda_cla32_fa698_xor1 = f_u_dadda_cla32_fa698_xor0 ^ f_u_dadda_cla32_fa76_xor1;
  assign f_u_dadda_cla32_fa698_and1 = f_u_dadda_cla32_fa698_xor0 & f_u_dadda_cla32_fa76_xor1;
  assign f_u_dadda_cla32_fa698_or0 = f_u_dadda_cla32_fa698_and0 | f_u_dadda_cla32_fa698_and1;
  assign f_u_dadda_cla32_fa699_xor0 = f_u_dadda_cla32_fa77_xor1 ^ f_u_dadda_cla32_fa78_xor1;
  assign f_u_dadda_cla32_fa699_and0 = f_u_dadda_cla32_fa77_xor1 & f_u_dadda_cla32_fa78_xor1;
  assign f_u_dadda_cla32_fa699_xor1 = f_u_dadda_cla32_fa699_xor0 ^ f_u_dadda_cla32_fa79_xor1;
  assign f_u_dadda_cla32_fa699_and1 = f_u_dadda_cla32_fa699_xor0 & f_u_dadda_cla32_fa79_xor1;
  assign f_u_dadda_cla32_fa699_or0 = f_u_dadda_cla32_fa699_and0 | f_u_dadda_cla32_fa699_and1;
  assign f_u_dadda_cla32_fa700_xor0 = f_u_dadda_cla32_fa699_or0 ^ f_u_dadda_cla32_fa698_or0;
  assign f_u_dadda_cla32_fa700_and0 = f_u_dadda_cla32_fa699_or0 & f_u_dadda_cla32_fa698_or0;
  assign f_u_dadda_cla32_fa700_xor1 = f_u_dadda_cla32_fa700_xor0 ^ f_u_dadda_cla32_fa88_xor1;
  assign f_u_dadda_cla32_fa700_and1 = f_u_dadda_cla32_fa700_xor0 & f_u_dadda_cla32_fa88_xor1;
  assign f_u_dadda_cla32_fa700_or0 = f_u_dadda_cla32_fa700_and0 | f_u_dadda_cla32_fa700_and1;
  assign f_u_dadda_cla32_fa701_xor0 = f_u_dadda_cla32_fa89_xor1 ^ f_u_dadda_cla32_fa90_xor1;
  assign f_u_dadda_cla32_fa701_and0 = f_u_dadda_cla32_fa89_xor1 & f_u_dadda_cla32_fa90_xor1;
  assign f_u_dadda_cla32_fa701_xor1 = f_u_dadda_cla32_fa701_xor0 ^ f_u_dadda_cla32_fa91_xor1;
  assign f_u_dadda_cla32_fa701_and1 = f_u_dadda_cla32_fa701_xor0 & f_u_dadda_cla32_fa91_xor1;
  assign f_u_dadda_cla32_fa701_or0 = f_u_dadda_cla32_fa701_and0 | f_u_dadda_cla32_fa701_and1;
  assign f_u_dadda_cla32_fa702_xor0 = f_u_dadda_cla32_fa701_or0 ^ f_u_dadda_cla32_fa700_or0;
  assign f_u_dadda_cla32_fa702_and0 = f_u_dadda_cla32_fa701_or0 & f_u_dadda_cla32_fa700_or0;
  assign f_u_dadda_cla32_fa702_xor1 = f_u_dadda_cla32_fa702_xor0 ^ f_u_dadda_cla32_fa101_xor1;
  assign f_u_dadda_cla32_fa702_and1 = f_u_dadda_cla32_fa702_xor0 & f_u_dadda_cla32_fa101_xor1;
  assign f_u_dadda_cla32_fa702_or0 = f_u_dadda_cla32_fa702_and0 | f_u_dadda_cla32_fa702_and1;
  assign f_u_dadda_cla32_fa703_xor0 = f_u_dadda_cla32_fa102_xor1 ^ f_u_dadda_cla32_fa103_xor1;
  assign f_u_dadda_cla32_fa703_and0 = f_u_dadda_cla32_fa102_xor1 & f_u_dadda_cla32_fa103_xor1;
  assign f_u_dadda_cla32_fa703_xor1 = f_u_dadda_cla32_fa703_xor0 ^ f_u_dadda_cla32_fa104_xor1;
  assign f_u_dadda_cla32_fa703_and1 = f_u_dadda_cla32_fa703_xor0 & f_u_dadda_cla32_fa104_xor1;
  assign f_u_dadda_cla32_fa703_or0 = f_u_dadda_cla32_fa703_and0 | f_u_dadda_cla32_fa703_and1;
  assign f_u_dadda_cla32_fa704_xor0 = f_u_dadda_cla32_fa703_or0 ^ f_u_dadda_cla32_fa702_or0;
  assign f_u_dadda_cla32_fa704_and0 = f_u_dadda_cla32_fa703_or0 & f_u_dadda_cla32_fa702_or0;
  assign f_u_dadda_cla32_fa704_xor1 = f_u_dadda_cla32_fa704_xor0 ^ f_u_dadda_cla32_fa115_xor1;
  assign f_u_dadda_cla32_fa704_and1 = f_u_dadda_cla32_fa704_xor0 & f_u_dadda_cla32_fa115_xor1;
  assign f_u_dadda_cla32_fa704_or0 = f_u_dadda_cla32_fa704_and0 | f_u_dadda_cla32_fa704_and1;
  assign f_u_dadda_cla32_fa705_xor0 = f_u_dadda_cla32_fa116_xor1 ^ f_u_dadda_cla32_fa117_xor1;
  assign f_u_dadda_cla32_fa705_and0 = f_u_dadda_cla32_fa116_xor1 & f_u_dadda_cla32_fa117_xor1;
  assign f_u_dadda_cla32_fa705_xor1 = f_u_dadda_cla32_fa705_xor0 ^ f_u_dadda_cla32_fa118_xor1;
  assign f_u_dadda_cla32_fa705_and1 = f_u_dadda_cla32_fa705_xor0 & f_u_dadda_cla32_fa118_xor1;
  assign f_u_dadda_cla32_fa705_or0 = f_u_dadda_cla32_fa705_and0 | f_u_dadda_cla32_fa705_and1;
  assign f_u_dadda_cla32_fa706_xor0 = f_u_dadda_cla32_fa705_or0 ^ f_u_dadda_cla32_fa704_or0;
  assign f_u_dadda_cla32_fa706_and0 = f_u_dadda_cla32_fa705_or0 & f_u_dadda_cla32_fa704_or0;
  assign f_u_dadda_cla32_fa706_xor1 = f_u_dadda_cla32_fa706_xor0 ^ f_u_dadda_cla32_fa130_xor1;
  assign f_u_dadda_cla32_fa706_and1 = f_u_dadda_cla32_fa706_xor0 & f_u_dadda_cla32_fa130_xor1;
  assign f_u_dadda_cla32_fa706_or0 = f_u_dadda_cla32_fa706_and0 | f_u_dadda_cla32_fa706_and1;
  assign f_u_dadda_cla32_fa707_xor0 = f_u_dadda_cla32_fa131_xor1 ^ f_u_dadda_cla32_fa132_xor1;
  assign f_u_dadda_cla32_fa707_and0 = f_u_dadda_cla32_fa131_xor1 & f_u_dadda_cla32_fa132_xor1;
  assign f_u_dadda_cla32_fa707_xor1 = f_u_dadda_cla32_fa707_xor0 ^ f_u_dadda_cla32_fa133_xor1;
  assign f_u_dadda_cla32_fa707_and1 = f_u_dadda_cla32_fa707_xor0 & f_u_dadda_cla32_fa133_xor1;
  assign f_u_dadda_cla32_fa707_or0 = f_u_dadda_cla32_fa707_and0 | f_u_dadda_cla32_fa707_and1;
  assign f_u_dadda_cla32_fa708_xor0 = f_u_dadda_cla32_fa707_or0 ^ f_u_dadda_cla32_fa706_or0;
  assign f_u_dadda_cla32_fa708_and0 = f_u_dadda_cla32_fa707_or0 & f_u_dadda_cla32_fa706_or0;
  assign f_u_dadda_cla32_fa708_xor1 = f_u_dadda_cla32_fa708_xor0 ^ f_u_dadda_cla32_fa146_xor1;
  assign f_u_dadda_cla32_fa708_and1 = f_u_dadda_cla32_fa708_xor0 & f_u_dadda_cla32_fa146_xor1;
  assign f_u_dadda_cla32_fa708_or0 = f_u_dadda_cla32_fa708_and0 | f_u_dadda_cla32_fa708_and1;
  assign f_u_dadda_cla32_fa709_xor0 = f_u_dadda_cla32_fa147_xor1 ^ f_u_dadda_cla32_fa148_xor1;
  assign f_u_dadda_cla32_fa709_and0 = f_u_dadda_cla32_fa147_xor1 & f_u_dadda_cla32_fa148_xor1;
  assign f_u_dadda_cla32_fa709_xor1 = f_u_dadda_cla32_fa709_xor0 ^ f_u_dadda_cla32_fa149_xor1;
  assign f_u_dadda_cla32_fa709_and1 = f_u_dadda_cla32_fa709_xor0 & f_u_dadda_cla32_fa149_xor1;
  assign f_u_dadda_cla32_fa709_or0 = f_u_dadda_cla32_fa709_and0 | f_u_dadda_cla32_fa709_and1;
  assign f_u_dadda_cla32_fa710_xor0 = f_u_dadda_cla32_fa709_or0 ^ f_u_dadda_cla32_fa708_or0;
  assign f_u_dadda_cla32_fa710_and0 = f_u_dadda_cla32_fa709_or0 & f_u_dadda_cla32_fa708_or0;
  assign f_u_dadda_cla32_fa710_xor1 = f_u_dadda_cla32_fa710_xor0 ^ f_u_dadda_cla32_fa163_xor1;
  assign f_u_dadda_cla32_fa710_and1 = f_u_dadda_cla32_fa710_xor0 & f_u_dadda_cla32_fa163_xor1;
  assign f_u_dadda_cla32_fa710_or0 = f_u_dadda_cla32_fa710_and0 | f_u_dadda_cla32_fa710_and1;
  assign f_u_dadda_cla32_fa711_xor0 = f_u_dadda_cla32_fa164_xor1 ^ f_u_dadda_cla32_fa165_xor1;
  assign f_u_dadda_cla32_fa711_and0 = f_u_dadda_cla32_fa164_xor1 & f_u_dadda_cla32_fa165_xor1;
  assign f_u_dadda_cla32_fa711_xor1 = f_u_dadda_cla32_fa711_xor0 ^ f_u_dadda_cla32_fa166_xor1;
  assign f_u_dadda_cla32_fa711_and1 = f_u_dadda_cla32_fa711_xor0 & f_u_dadda_cla32_fa166_xor1;
  assign f_u_dadda_cla32_fa711_or0 = f_u_dadda_cla32_fa711_and0 | f_u_dadda_cla32_fa711_and1;
  assign f_u_dadda_cla32_fa712_xor0 = f_u_dadda_cla32_fa711_or0 ^ f_u_dadda_cla32_fa710_or0;
  assign f_u_dadda_cla32_fa712_and0 = f_u_dadda_cla32_fa711_or0 & f_u_dadda_cla32_fa710_or0;
  assign f_u_dadda_cla32_fa712_xor1 = f_u_dadda_cla32_fa712_xor0 ^ f_u_dadda_cla32_fa181_xor1;
  assign f_u_dadda_cla32_fa712_and1 = f_u_dadda_cla32_fa712_xor0 & f_u_dadda_cla32_fa181_xor1;
  assign f_u_dadda_cla32_fa712_or0 = f_u_dadda_cla32_fa712_and0 | f_u_dadda_cla32_fa712_and1;
  assign f_u_dadda_cla32_fa713_xor0 = f_u_dadda_cla32_fa182_xor1 ^ f_u_dadda_cla32_fa183_xor1;
  assign f_u_dadda_cla32_fa713_and0 = f_u_dadda_cla32_fa182_xor1 & f_u_dadda_cla32_fa183_xor1;
  assign f_u_dadda_cla32_fa713_xor1 = f_u_dadda_cla32_fa713_xor0 ^ f_u_dadda_cla32_fa184_xor1;
  assign f_u_dadda_cla32_fa713_and1 = f_u_dadda_cla32_fa713_xor0 & f_u_dadda_cla32_fa184_xor1;
  assign f_u_dadda_cla32_fa713_or0 = f_u_dadda_cla32_fa713_and0 | f_u_dadda_cla32_fa713_and1;
  assign f_u_dadda_cla32_fa714_xor0 = f_u_dadda_cla32_fa713_or0 ^ f_u_dadda_cla32_fa712_or0;
  assign f_u_dadda_cla32_fa714_and0 = f_u_dadda_cla32_fa713_or0 & f_u_dadda_cla32_fa712_or0;
  assign f_u_dadda_cla32_fa714_xor1 = f_u_dadda_cla32_fa714_xor0 ^ f_u_dadda_cla32_fa200_xor1;
  assign f_u_dadda_cla32_fa714_and1 = f_u_dadda_cla32_fa714_xor0 & f_u_dadda_cla32_fa200_xor1;
  assign f_u_dadda_cla32_fa714_or0 = f_u_dadda_cla32_fa714_and0 | f_u_dadda_cla32_fa714_and1;
  assign f_u_dadda_cla32_fa715_xor0 = f_u_dadda_cla32_fa201_xor1 ^ f_u_dadda_cla32_fa202_xor1;
  assign f_u_dadda_cla32_fa715_and0 = f_u_dadda_cla32_fa201_xor1 & f_u_dadda_cla32_fa202_xor1;
  assign f_u_dadda_cla32_fa715_xor1 = f_u_dadda_cla32_fa715_xor0 ^ f_u_dadda_cla32_fa203_xor1;
  assign f_u_dadda_cla32_fa715_and1 = f_u_dadda_cla32_fa715_xor0 & f_u_dadda_cla32_fa203_xor1;
  assign f_u_dadda_cla32_fa715_or0 = f_u_dadda_cla32_fa715_and0 | f_u_dadda_cla32_fa715_and1;
  assign f_u_dadda_cla32_fa716_xor0 = f_u_dadda_cla32_fa715_or0 ^ f_u_dadda_cla32_fa714_or0;
  assign f_u_dadda_cla32_fa716_and0 = f_u_dadda_cla32_fa715_or0 & f_u_dadda_cla32_fa714_or0;
  assign f_u_dadda_cla32_fa716_xor1 = f_u_dadda_cla32_fa716_xor0 ^ f_u_dadda_cla32_fa220_xor1;
  assign f_u_dadda_cla32_fa716_and1 = f_u_dadda_cla32_fa716_xor0 & f_u_dadda_cla32_fa220_xor1;
  assign f_u_dadda_cla32_fa716_or0 = f_u_dadda_cla32_fa716_and0 | f_u_dadda_cla32_fa716_and1;
  assign f_u_dadda_cla32_fa717_xor0 = f_u_dadda_cla32_fa221_xor1 ^ f_u_dadda_cla32_fa222_xor1;
  assign f_u_dadda_cla32_fa717_and0 = f_u_dadda_cla32_fa221_xor1 & f_u_dadda_cla32_fa222_xor1;
  assign f_u_dadda_cla32_fa717_xor1 = f_u_dadda_cla32_fa717_xor0 ^ f_u_dadda_cla32_fa223_xor1;
  assign f_u_dadda_cla32_fa717_and1 = f_u_dadda_cla32_fa717_xor0 & f_u_dadda_cla32_fa223_xor1;
  assign f_u_dadda_cla32_fa717_or0 = f_u_dadda_cla32_fa717_and0 | f_u_dadda_cla32_fa717_and1;
  assign f_u_dadda_cla32_fa718_xor0 = f_u_dadda_cla32_fa717_or0 ^ f_u_dadda_cla32_fa716_or0;
  assign f_u_dadda_cla32_fa718_and0 = f_u_dadda_cla32_fa717_or0 & f_u_dadda_cla32_fa716_or0;
  assign f_u_dadda_cla32_fa718_xor1 = f_u_dadda_cla32_fa718_xor0 ^ f_u_dadda_cla32_fa241_xor1;
  assign f_u_dadda_cla32_fa718_and1 = f_u_dadda_cla32_fa718_xor0 & f_u_dadda_cla32_fa241_xor1;
  assign f_u_dadda_cla32_fa718_or0 = f_u_dadda_cla32_fa718_and0 | f_u_dadda_cla32_fa718_and1;
  assign f_u_dadda_cla32_fa719_xor0 = f_u_dadda_cla32_fa242_xor1 ^ f_u_dadda_cla32_fa243_xor1;
  assign f_u_dadda_cla32_fa719_and0 = f_u_dadda_cla32_fa242_xor1 & f_u_dadda_cla32_fa243_xor1;
  assign f_u_dadda_cla32_fa719_xor1 = f_u_dadda_cla32_fa719_xor0 ^ f_u_dadda_cla32_fa244_xor1;
  assign f_u_dadda_cla32_fa719_and1 = f_u_dadda_cla32_fa719_xor0 & f_u_dadda_cla32_fa244_xor1;
  assign f_u_dadda_cla32_fa719_or0 = f_u_dadda_cla32_fa719_and0 | f_u_dadda_cla32_fa719_and1;
  assign f_u_dadda_cla32_fa720_xor0 = f_u_dadda_cla32_fa719_or0 ^ f_u_dadda_cla32_fa718_or0;
  assign f_u_dadda_cla32_fa720_and0 = f_u_dadda_cla32_fa719_or0 & f_u_dadda_cla32_fa718_or0;
  assign f_u_dadda_cla32_fa720_xor1 = f_u_dadda_cla32_fa720_xor0 ^ f_u_dadda_cla32_fa262_xor1;
  assign f_u_dadda_cla32_fa720_and1 = f_u_dadda_cla32_fa720_xor0 & f_u_dadda_cla32_fa262_xor1;
  assign f_u_dadda_cla32_fa720_or0 = f_u_dadda_cla32_fa720_and0 | f_u_dadda_cla32_fa720_and1;
  assign f_u_dadda_cla32_fa721_xor0 = f_u_dadda_cla32_fa263_xor1 ^ f_u_dadda_cla32_fa264_xor1;
  assign f_u_dadda_cla32_fa721_and0 = f_u_dadda_cla32_fa263_xor1 & f_u_dadda_cla32_fa264_xor1;
  assign f_u_dadda_cla32_fa721_xor1 = f_u_dadda_cla32_fa721_xor0 ^ f_u_dadda_cla32_fa265_xor1;
  assign f_u_dadda_cla32_fa721_and1 = f_u_dadda_cla32_fa721_xor0 & f_u_dadda_cla32_fa265_xor1;
  assign f_u_dadda_cla32_fa721_or0 = f_u_dadda_cla32_fa721_and0 | f_u_dadda_cla32_fa721_and1;
  assign f_u_dadda_cla32_fa722_xor0 = f_u_dadda_cla32_fa721_or0 ^ f_u_dadda_cla32_fa720_or0;
  assign f_u_dadda_cla32_fa722_and0 = f_u_dadda_cla32_fa721_or0 & f_u_dadda_cla32_fa720_or0;
  assign f_u_dadda_cla32_fa722_xor1 = f_u_dadda_cla32_fa722_xor0 ^ f_u_dadda_cla32_fa284_xor1;
  assign f_u_dadda_cla32_fa722_and1 = f_u_dadda_cla32_fa722_xor0 & f_u_dadda_cla32_fa284_xor1;
  assign f_u_dadda_cla32_fa722_or0 = f_u_dadda_cla32_fa722_and0 | f_u_dadda_cla32_fa722_and1;
  assign f_u_dadda_cla32_fa723_xor0 = f_u_dadda_cla32_fa285_xor1 ^ f_u_dadda_cla32_fa286_xor1;
  assign f_u_dadda_cla32_fa723_and0 = f_u_dadda_cla32_fa285_xor1 & f_u_dadda_cla32_fa286_xor1;
  assign f_u_dadda_cla32_fa723_xor1 = f_u_dadda_cla32_fa723_xor0 ^ f_u_dadda_cla32_fa287_xor1;
  assign f_u_dadda_cla32_fa723_and1 = f_u_dadda_cla32_fa723_xor0 & f_u_dadda_cla32_fa287_xor1;
  assign f_u_dadda_cla32_fa723_or0 = f_u_dadda_cla32_fa723_and0 | f_u_dadda_cla32_fa723_and1;
  assign f_u_dadda_cla32_fa724_xor0 = f_u_dadda_cla32_fa723_or0 ^ f_u_dadda_cla32_fa722_or0;
  assign f_u_dadda_cla32_fa724_and0 = f_u_dadda_cla32_fa723_or0 & f_u_dadda_cla32_fa722_or0;
  assign f_u_dadda_cla32_fa724_xor1 = f_u_dadda_cla32_fa724_xor0 ^ f_u_dadda_cla32_fa306_xor1;
  assign f_u_dadda_cla32_fa724_and1 = f_u_dadda_cla32_fa724_xor0 & f_u_dadda_cla32_fa306_xor1;
  assign f_u_dadda_cla32_fa724_or0 = f_u_dadda_cla32_fa724_and0 | f_u_dadda_cla32_fa724_and1;
  assign f_u_dadda_cla32_fa725_xor0 = f_u_dadda_cla32_fa307_xor1 ^ f_u_dadda_cla32_fa308_xor1;
  assign f_u_dadda_cla32_fa725_and0 = f_u_dadda_cla32_fa307_xor1 & f_u_dadda_cla32_fa308_xor1;
  assign f_u_dadda_cla32_fa725_xor1 = f_u_dadda_cla32_fa725_xor0 ^ f_u_dadda_cla32_fa309_xor1;
  assign f_u_dadda_cla32_fa725_and1 = f_u_dadda_cla32_fa725_xor0 & f_u_dadda_cla32_fa309_xor1;
  assign f_u_dadda_cla32_fa725_or0 = f_u_dadda_cla32_fa725_and0 | f_u_dadda_cla32_fa725_and1;
  assign f_u_dadda_cla32_fa726_xor0 = f_u_dadda_cla32_fa725_or0 ^ f_u_dadda_cla32_fa724_or0;
  assign f_u_dadda_cla32_fa726_and0 = f_u_dadda_cla32_fa725_or0 & f_u_dadda_cla32_fa724_or0;
  assign f_u_dadda_cla32_fa726_xor1 = f_u_dadda_cla32_fa726_xor0 ^ f_u_dadda_cla32_fa328_xor1;
  assign f_u_dadda_cla32_fa726_and1 = f_u_dadda_cla32_fa726_xor0 & f_u_dadda_cla32_fa328_xor1;
  assign f_u_dadda_cla32_fa726_or0 = f_u_dadda_cla32_fa726_and0 | f_u_dadda_cla32_fa726_and1;
  assign f_u_dadda_cla32_fa727_xor0 = f_u_dadda_cla32_fa329_xor1 ^ f_u_dadda_cla32_fa330_xor1;
  assign f_u_dadda_cla32_fa727_and0 = f_u_dadda_cla32_fa329_xor1 & f_u_dadda_cla32_fa330_xor1;
  assign f_u_dadda_cla32_fa727_xor1 = f_u_dadda_cla32_fa727_xor0 ^ f_u_dadda_cla32_fa331_xor1;
  assign f_u_dadda_cla32_fa727_and1 = f_u_dadda_cla32_fa727_xor0 & f_u_dadda_cla32_fa331_xor1;
  assign f_u_dadda_cla32_fa727_or0 = f_u_dadda_cla32_fa727_and0 | f_u_dadda_cla32_fa727_and1;
  assign f_u_dadda_cla32_fa728_xor0 = f_u_dadda_cla32_fa727_or0 ^ f_u_dadda_cla32_fa726_or0;
  assign f_u_dadda_cla32_fa728_and0 = f_u_dadda_cla32_fa727_or0 & f_u_dadda_cla32_fa726_or0;
  assign f_u_dadda_cla32_fa728_xor1 = f_u_dadda_cla32_fa728_xor0 ^ f_u_dadda_cla32_fa350_xor1;
  assign f_u_dadda_cla32_fa728_and1 = f_u_dadda_cla32_fa728_xor0 & f_u_dadda_cla32_fa350_xor1;
  assign f_u_dadda_cla32_fa728_or0 = f_u_dadda_cla32_fa728_and0 | f_u_dadda_cla32_fa728_and1;
  assign f_u_dadda_cla32_fa729_xor0 = f_u_dadda_cla32_fa351_xor1 ^ f_u_dadda_cla32_fa352_xor1;
  assign f_u_dadda_cla32_fa729_and0 = f_u_dadda_cla32_fa351_xor1 & f_u_dadda_cla32_fa352_xor1;
  assign f_u_dadda_cla32_fa729_xor1 = f_u_dadda_cla32_fa729_xor0 ^ f_u_dadda_cla32_fa353_xor1;
  assign f_u_dadda_cla32_fa729_and1 = f_u_dadda_cla32_fa729_xor0 & f_u_dadda_cla32_fa353_xor1;
  assign f_u_dadda_cla32_fa729_or0 = f_u_dadda_cla32_fa729_and0 | f_u_dadda_cla32_fa729_and1;
  assign f_u_dadda_cla32_fa730_xor0 = f_u_dadda_cla32_fa729_or0 ^ f_u_dadda_cla32_fa728_or0;
  assign f_u_dadda_cla32_fa730_and0 = f_u_dadda_cla32_fa729_or0 & f_u_dadda_cla32_fa728_or0;
  assign f_u_dadda_cla32_fa730_xor1 = f_u_dadda_cla32_fa730_xor0 ^ f_u_dadda_cla32_fa372_xor1;
  assign f_u_dadda_cla32_fa730_and1 = f_u_dadda_cla32_fa730_xor0 & f_u_dadda_cla32_fa372_xor1;
  assign f_u_dadda_cla32_fa730_or0 = f_u_dadda_cla32_fa730_and0 | f_u_dadda_cla32_fa730_and1;
  assign f_u_dadda_cla32_fa731_xor0 = f_u_dadda_cla32_fa373_xor1 ^ f_u_dadda_cla32_fa374_xor1;
  assign f_u_dadda_cla32_fa731_and0 = f_u_dadda_cla32_fa373_xor1 & f_u_dadda_cla32_fa374_xor1;
  assign f_u_dadda_cla32_fa731_xor1 = f_u_dadda_cla32_fa731_xor0 ^ f_u_dadda_cla32_fa375_xor1;
  assign f_u_dadda_cla32_fa731_and1 = f_u_dadda_cla32_fa731_xor0 & f_u_dadda_cla32_fa375_xor1;
  assign f_u_dadda_cla32_fa731_or0 = f_u_dadda_cla32_fa731_and0 | f_u_dadda_cla32_fa731_and1;
  assign f_u_dadda_cla32_fa732_xor0 = f_u_dadda_cla32_fa731_or0 ^ f_u_dadda_cla32_fa730_or0;
  assign f_u_dadda_cla32_fa732_and0 = f_u_dadda_cla32_fa731_or0 & f_u_dadda_cla32_fa730_or0;
  assign f_u_dadda_cla32_fa732_xor1 = f_u_dadda_cla32_fa732_xor0 ^ f_u_dadda_cla32_fa394_xor1;
  assign f_u_dadda_cla32_fa732_and1 = f_u_dadda_cla32_fa732_xor0 & f_u_dadda_cla32_fa394_xor1;
  assign f_u_dadda_cla32_fa732_or0 = f_u_dadda_cla32_fa732_and0 | f_u_dadda_cla32_fa732_and1;
  assign f_u_dadda_cla32_fa733_xor0 = f_u_dadda_cla32_fa395_xor1 ^ f_u_dadda_cla32_fa396_xor1;
  assign f_u_dadda_cla32_fa733_and0 = f_u_dadda_cla32_fa395_xor1 & f_u_dadda_cla32_fa396_xor1;
  assign f_u_dadda_cla32_fa733_xor1 = f_u_dadda_cla32_fa733_xor0 ^ f_u_dadda_cla32_fa397_xor1;
  assign f_u_dadda_cla32_fa733_and1 = f_u_dadda_cla32_fa733_xor0 & f_u_dadda_cla32_fa397_xor1;
  assign f_u_dadda_cla32_fa733_or0 = f_u_dadda_cla32_fa733_and0 | f_u_dadda_cla32_fa733_and1;
  assign f_u_dadda_cla32_fa734_xor0 = f_u_dadda_cla32_fa733_or0 ^ f_u_dadda_cla32_fa732_or0;
  assign f_u_dadda_cla32_fa734_and0 = f_u_dadda_cla32_fa733_or0 & f_u_dadda_cla32_fa732_or0;
  assign f_u_dadda_cla32_fa734_xor1 = f_u_dadda_cla32_fa734_xor0 ^ f_u_dadda_cla32_fa416_xor1;
  assign f_u_dadda_cla32_fa734_and1 = f_u_dadda_cla32_fa734_xor0 & f_u_dadda_cla32_fa416_xor1;
  assign f_u_dadda_cla32_fa734_or0 = f_u_dadda_cla32_fa734_and0 | f_u_dadda_cla32_fa734_and1;
  assign f_u_dadda_cla32_fa735_xor0 = f_u_dadda_cla32_fa417_xor1 ^ f_u_dadda_cla32_fa418_xor1;
  assign f_u_dadda_cla32_fa735_and0 = f_u_dadda_cla32_fa417_xor1 & f_u_dadda_cla32_fa418_xor1;
  assign f_u_dadda_cla32_fa735_xor1 = f_u_dadda_cla32_fa735_xor0 ^ f_u_dadda_cla32_fa419_xor1;
  assign f_u_dadda_cla32_fa735_and1 = f_u_dadda_cla32_fa735_xor0 & f_u_dadda_cla32_fa419_xor1;
  assign f_u_dadda_cla32_fa735_or0 = f_u_dadda_cla32_fa735_and0 | f_u_dadda_cla32_fa735_and1;
  assign f_u_dadda_cla32_fa736_xor0 = f_u_dadda_cla32_fa735_or0 ^ f_u_dadda_cla32_fa734_or0;
  assign f_u_dadda_cla32_fa736_and0 = f_u_dadda_cla32_fa735_or0 & f_u_dadda_cla32_fa734_or0;
  assign f_u_dadda_cla32_fa736_xor1 = f_u_dadda_cla32_fa736_xor0 ^ f_u_dadda_cla32_fa438_xor1;
  assign f_u_dadda_cla32_fa736_and1 = f_u_dadda_cla32_fa736_xor0 & f_u_dadda_cla32_fa438_xor1;
  assign f_u_dadda_cla32_fa736_or0 = f_u_dadda_cla32_fa736_and0 | f_u_dadda_cla32_fa736_and1;
  assign f_u_dadda_cla32_fa737_xor0 = f_u_dadda_cla32_fa439_xor1 ^ f_u_dadda_cla32_fa440_xor1;
  assign f_u_dadda_cla32_fa737_and0 = f_u_dadda_cla32_fa439_xor1 & f_u_dadda_cla32_fa440_xor1;
  assign f_u_dadda_cla32_fa737_xor1 = f_u_dadda_cla32_fa737_xor0 ^ f_u_dadda_cla32_fa441_xor1;
  assign f_u_dadda_cla32_fa737_and1 = f_u_dadda_cla32_fa737_xor0 & f_u_dadda_cla32_fa441_xor1;
  assign f_u_dadda_cla32_fa737_or0 = f_u_dadda_cla32_fa737_and0 | f_u_dadda_cla32_fa737_and1;
  assign f_u_dadda_cla32_fa738_xor0 = f_u_dadda_cla32_fa737_or0 ^ f_u_dadda_cla32_fa736_or0;
  assign f_u_dadda_cla32_fa738_and0 = f_u_dadda_cla32_fa737_or0 & f_u_dadda_cla32_fa736_or0;
  assign f_u_dadda_cla32_fa738_xor1 = f_u_dadda_cla32_fa738_xor0 ^ f_u_dadda_cla32_fa459_xor1;
  assign f_u_dadda_cla32_fa738_and1 = f_u_dadda_cla32_fa738_xor0 & f_u_dadda_cla32_fa459_xor1;
  assign f_u_dadda_cla32_fa738_or0 = f_u_dadda_cla32_fa738_and0 | f_u_dadda_cla32_fa738_and1;
  assign f_u_dadda_cla32_fa739_xor0 = f_u_dadda_cla32_fa460_xor1 ^ f_u_dadda_cla32_fa461_xor1;
  assign f_u_dadda_cla32_fa739_and0 = f_u_dadda_cla32_fa460_xor1 & f_u_dadda_cla32_fa461_xor1;
  assign f_u_dadda_cla32_fa739_xor1 = f_u_dadda_cla32_fa739_xor0 ^ f_u_dadda_cla32_fa462_xor1;
  assign f_u_dadda_cla32_fa739_and1 = f_u_dadda_cla32_fa739_xor0 & f_u_dadda_cla32_fa462_xor1;
  assign f_u_dadda_cla32_fa739_or0 = f_u_dadda_cla32_fa739_and0 | f_u_dadda_cla32_fa739_and1;
  assign f_u_dadda_cla32_fa740_xor0 = f_u_dadda_cla32_fa739_or0 ^ f_u_dadda_cla32_fa738_or0;
  assign f_u_dadda_cla32_fa740_and0 = f_u_dadda_cla32_fa739_or0 & f_u_dadda_cla32_fa738_or0;
  assign f_u_dadda_cla32_fa740_xor1 = f_u_dadda_cla32_fa740_xor0 ^ f_u_dadda_cla32_fa479_xor1;
  assign f_u_dadda_cla32_fa740_and1 = f_u_dadda_cla32_fa740_xor0 & f_u_dadda_cla32_fa479_xor1;
  assign f_u_dadda_cla32_fa740_or0 = f_u_dadda_cla32_fa740_and0 | f_u_dadda_cla32_fa740_and1;
  assign f_u_dadda_cla32_fa741_xor0 = f_u_dadda_cla32_fa480_xor1 ^ f_u_dadda_cla32_fa481_xor1;
  assign f_u_dadda_cla32_fa741_and0 = f_u_dadda_cla32_fa480_xor1 & f_u_dadda_cla32_fa481_xor1;
  assign f_u_dadda_cla32_fa741_xor1 = f_u_dadda_cla32_fa741_xor0 ^ f_u_dadda_cla32_fa482_xor1;
  assign f_u_dadda_cla32_fa741_and1 = f_u_dadda_cla32_fa741_xor0 & f_u_dadda_cla32_fa482_xor1;
  assign f_u_dadda_cla32_fa741_or0 = f_u_dadda_cla32_fa741_and0 | f_u_dadda_cla32_fa741_and1;
  assign f_u_dadda_cla32_fa742_xor0 = f_u_dadda_cla32_fa741_or0 ^ f_u_dadda_cla32_fa740_or0;
  assign f_u_dadda_cla32_fa742_and0 = f_u_dadda_cla32_fa741_or0 & f_u_dadda_cla32_fa740_or0;
  assign f_u_dadda_cla32_fa742_xor1 = f_u_dadda_cla32_fa742_xor0 ^ f_u_dadda_cla32_fa498_xor1;
  assign f_u_dadda_cla32_fa742_and1 = f_u_dadda_cla32_fa742_xor0 & f_u_dadda_cla32_fa498_xor1;
  assign f_u_dadda_cla32_fa742_or0 = f_u_dadda_cla32_fa742_and0 | f_u_dadda_cla32_fa742_and1;
  assign f_u_dadda_cla32_fa743_xor0 = f_u_dadda_cla32_fa499_xor1 ^ f_u_dadda_cla32_fa500_xor1;
  assign f_u_dadda_cla32_fa743_and0 = f_u_dadda_cla32_fa499_xor1 & f_u_dadda_cla32_fa500_xor1;
  assign f_u_dadda_cla32_fa743_xor1 = f_u_dadda_cla32_fa743_xor0 ^ f_u_dadda_cla32_fa501_xor1;
  assign f_u_dadda_cla32_fa743_and1 = f_u_dadda_cla32_fa743_xor0 & f_u_dadda_cla32_fa501_xor1;
  assign f_u_dadda_cla32_fa743_or0 = f_u_dadda_cla32_fa743_and0 | f_u_dadda_cla32_fa743_and1;
  assign f_u_dadda_cla32_fa744_xor0 = f_u_dadda_cla32_fa743_or0 ^ f_u_dadda_cla32_fa742_or0;
  assign f_u_dadda_cla32_fa744_and0 = f_u_dadda_cla32_fa743_or0 & f_u_dadda_cla32_fa742_or0;
  assign f_u_dadda_cla32_fa744_xor1 = f_u_dadda_cla32_fa744_xor0 ^ f_u_dadda_cla32_fa516_xor1;
  assign f_u_dadda_cla32_fa744_and1 = f_u_dadda_cla32_fa744_xor0 & f_u_dadda_cla32_fa516_xor1;
  assign f_u_dadda_cla32_fa744_or0 = f_u_dadda_cla32_fa744_and0 | f_u_dadda_cla32_fa744_and1;
  assign f_u_dadda_cla32_fa745_xor0 = f_u_dadda_cla32_fa517_xor1 ^ f_u_dadda_cla32_fa518_xor1;
  assign f_u_dadda_cla32_fa745_and0 = f_u_dadda_cla32_fa517_xor1 & f_u_dadda_cla32_fa518_xor1;
  assign f_u_dadda_cla32_fa745_xor1 = f_u_dadda_cla32_fa745_xor0 ^ f_u_dadda_cla32_fa519_xor1;
  assign f_u_dadda_cla32_fa745_and1 = f_u_dadda_cla32_fa745_xor0 & f_u_dadda_cla32_fa519_xor1;
  assign f_u_dadda_cla32_fa745_or0 = f_u_dadda_cla32_fa745_and0 | f_u_dadda_cla32_fa745_and1;
  assign f_u_dadda_cla32_fa746_xor0 = f_u_dadda_cla32_fa745_or0 ^ f_u_dadda_cla32_fa744_or0;
  assign f_u_dadda_cla32_fa746_and0 = f_u_dadda_cla32_fa745_or0 & f_u_dadda_cla32_fa744_or0;
  assign f_u_dadda_cla32_fa746_xor1 = f_u_dadda_cla32_fa746_xor0 ^ f_u_dadda_cla32_fa533_xor1;
  assign f_u_dadda_cla32_fa746_and1 = f_u_dadda_cla32_fa746_xor0 & f_u_dadda_cla32_fa533_xor1;
  assign f_u_dadda_cla32_fa746_or0 = f_u_dadda_cla32_fa746_and0 | f_u_dadda_cla32_fa746_and1;
  assign f_u_dadda_cla32_fa747_xor0 = f_u_dadda_cla32_fa534_xor1 ^ f_u_dadda_cla32_fa535_xor1;
  assign f_u_dadda_cla32_fa747_and0 = f_u_dadda_cla32_fa534_xor1 & f_u_dadda_cla32_fa535_xor1;
  assign f_u_dadda_cla32_fa747_xor1 = f_u_dadda_cla32_fa747_xor0 ^ f_u_dadda_cla32_fa536_xor1;
  assign f_u_dadda_cla32_fa747_and1 = f_u_dadda_cla32_fa747_xor0 & f_u_dadda_cla32_fa536_xor1;
  assign f_u_dadda_cla32_fa747_or0 = f_u_dadda_cla32_fa747_and0 | f_u_dadda_cla32_fa747_and1;
  assign f_u_dadda_cla32_fa748_xor0 = f_u_dadda_cla32_fa747_or0 ^ f_u_dadda_cla32_fa746_or0;
  assign f_u_dadda_cla32_fa748_and0 = f_u_dadda_cla32_fa747_or0 & f_u_dadda_cla32_fa746_or0;
  assign f_u_dadda_cla32_fa748_xor1 = f_u_dadda_cla32_fa748_xor0 ^ f_u_dadda_cla32_fa549_xor1;
  assign f_u_dadda_cla32_fa748_and1 = f_u_dadda_cla32_fa748_xor0 & f_u_dadda_cla32_fa549_xor1;
  assign f_u_dadda_cla32_fa748_or0 = f_u_dadda_cla32_fa748_and0 | f_u_dadda_cla32_fa748_and1;
  assign f_u_dadda_cla32_fa749_xor0 = f_u_dadda_cla32_fa550_xor1 ^ f_u_dadda_cla32_fa551_xor1;
  assign f_u_dadda_cla32_fa749_and0 = f_u_dadda_cla32_fa550_xor1 & f_u_dadda_cla32_fa551_xor1;
  assign f_u_dadda_cla32_fa749_xor1 = f_u_dadda_cla32_fa749_xor0 ^ f_u_dadda_cla32_fa552_xor1;
  assign f_u_dadda_cla32_fa749_and1 = f_u_dadda_cla32_fa749_xor0 & f_u_dadda_cla32_fa552_xor1;
  assign f_u_dadda_cla32_fa749_or0 = f_u_dadda_cla32_fa749_and0 | f_u_dadda_cla32_fa749_and1;
  assign f_u_dadda_cla32_fa750_xor0 = f_u_dadda_cla32_fa749_or0 ^ f_u_dadda_cla32_fa748_or0;
  assign f_u_dadda_cla32_fa750_and0 = f_u_dadda_cla32_fa749_or0 & f_u_dadda_cla32_fa748_or0;
  assign f_u_dadda_cla32_fa750_xor1 = f_u_dadda_cla32_fa750_xor0 ^ f_u_dadda_cla32_fa564_xor1;
  assign f_u_dadda_cla32_fa750_and1 = f_u_dadda_cla32_fa750_xor0 & f_u_dadda_cla32_fa564_xor1;
  assign f_u_dadda_cla32_fa750_or0 = f_u_dadda_cla32_fa750_and0 | f_u_dadda_cla32_fa750_and1;
  assign f_u_dadda_cla32_fa751_xor0 = f_u_dadda_cla32_fa565_xor1 ^ f_u_dadda_cla32_fa566_xor1;
  assign f_u_dadda_cla32_fa751_and0 = f_u_dadda_cla32_fa565_xor1 & f_u_dadda_cla32_fa566_xor1;
  assign f_u_dadda_cla32_fa751_xor1 = f_u_dadda_cla32_fa751_xor0 ^ f_u_dadda_cla32_fa567_xor1;
  assign f_u_dadda_cla32_fa751_and1 = f_u_dadda_cla32_fa751_xor0 & f_u_dadda_cla32_fa567_xor1;
  assign f_u_dadda_cla32_fa751_or0 = f_u_dadda_cla32_fa751_and0 | f_u_dadda_cla32_fa751_and1;
  assign f_u_dadda_cla32_fa752_xor0 = f_u_dadda_cla32_fa751_or0 ^ f_u_dadda_cla32_fa750_or0;
  assign f_u_dadda_cla32_fa752_and0 = f_u_dadda_cla32_fa751_or0 & f_u_dadda_cla32_fa750_or0;
  assign f_u_dadda_cla32_fa752_xor1 = f_u_dadda_cla32_fa752_xor0 ^ f_u_dadda_cla32_fa578_xor1;
  assign f_u_dadda_cla32_fa752_and1 = f_u_dadda_cla32_fa752_xor0 & f_u_dadda_cla32_fa578_xor1;
  assign f_u_dadda_cla32_fa752_or0 = f_u_dadda_cla32_fa752_and0 | f_u_dadda_cla32_fa752_and1;
  assign f_u_dadda_cla32_fa753_xor0 = f_u_dadda_cla32_fa579_xor1 ^ f_u_dadda_cla32_fa580_xor1;
  assign f_u_dadda_cla32_fa753_and0 = f_u_dadda_cla32_fa579_xor1 & f_u_dadda_cla32_fa580_xor1;
  assign f_u_dadda_cla32_fa753_xor1 = f_u_dadda_cla32_fa753_xor0 ^ f_u_dadda_cla32_fa581_xor1;
  assign f_u_dadda_cla32_fa753_and1 = f_u_dadda_cla32_fa753_xor0 & f_u_dadda_cla32_fa581_xor1;
  assign f_u_dadda_cla32_fa753_or0 = f_u_dadda_cla32_fa753_and0 | f_u_dadda_cla32_fa753_and1;
  assign f_u_dadda_cla32_fa754_xor0 = f_u_dadda_cla32_fa753_or0 ^ f_u_dadda_cla32_fa752_or0;
  assign f_u_dadda_cla32_fa754_and0 = f_u_dadda_cla32_fa753_or0 & f_u_dadda_cla32_fa752_or0;
  assign f_u_dadda_cla32_fa754_xor1 = f_u_dadda_cla32_fa754_xor0 ^ f_u_dadda_cla32_fa591_xor1;
  assign f_u_dadda_cla32_fa754_and1 = f_u_dadda_cla32_fa754_xor0 & f_u_dadda_cla32_fa591_xor1;
  assign f_u_dadda_cla32_fa754_or0 = f_u_dadda_cla32_fa754_and0 | f_u_dadda_cla32_fa754_and1;
  assign f_u_dadda_cla32_fa755_xor0 = f_u_dadda_cla32_fa592_xor1 ^ f_u_dadda_cla32_fa593_xor1;
  assign f_u_dadda_cla32_fa755_and0 = f_u_dadda_cla32_fa592_xor1 & f_u_dadda_cla32_fa593_xor1;
  assign f_u_dadda_cla32_fa755_xor1 = f_u_dadda_cla32_fa755_xor0 ^ f_u_dadda_cla32_fa594_xor1;
  assign f_u_dadda_cla32_fa755_and1 = f_u_dadda_cla32_fa755_xor0 & f_u_dadda_cla32_fa594_xor1;
  assign f_u_dadda_cla32_fa755_or0 = f_u_dadda_cla32_fa755_and0 | f_u_dadda_cla32_fa755_and1;
  assign f_u_dadda_cla32_fa756_xor0 = f_u_dadda_cla32_fa755_or0 ^ f_u_dadda_cla32_fa754_or0;
  assign f_u_dadda_cla32_fa756_and0 = f_u_dadda_cla32_fa755_or0 & f_u_dadda_cla32_fa754_or0;
  assign f_u_dadda_cla32_fa756_xor1 = f_u_dadda_cla32_fa756_xor0 ^ f_u_dadda_cla32_fa603_xor1;
  assign f_u_dadda_cla32_fa756_and1 = f_u_dadda_cla32_fa756_xor0 & f_u_dadda_cla32_fa603_xor1;
  assign f_u_dadda_cla32_fa756_or0 = f_u_dadda_cla32_fa756_and0 | f_u_dadda_cla32_fa756_and1;
  assign f_u_dadda_cla32_fa757_xor0 = f_u_dadda_cla32_fa604_xor1 ^ f_u_dadda_cla32_fa605_xor1;
  assign f_u_dadda_cla32_fa757_and0 = f_u_dadda_cla32_fa604_xor1 & f_u_dadda_cla32_fa605_xor1;
  assign f_u_dadda_cla32_fa757_xor1 = f_u_dadda_cla32_fa757_xor0 ^ f_u_dadda_cla32_fa606_xor1;
  assign f_u_dadda_cla32_fa757_and1 = f_u_dadda_cla32_fa757_xor0 & f_u_dadda_cla32_fa606_xor1;
  assign f_u_dadda_cla32_fa757_or0 = f_u_dadda_cla32_fa757_and0 | f_u_dadda_cla32_fa757_and1;
  assign f_u_dadda_cla32_fa758_xor0 = f_u_dadda_cla32_fa757_or0 ^ f_u_dadda_cla32_fa756_or0;
  assign f_u_dadda_cla32_fa758_and0 = f_u_dadda_cla32_fa757_or0 & f_u_dadda_cla32_fa756_or0;
  assign f_u_dadda_cla32_fa758_xor1 = f_u_dadda_cla32_fa758_xor0 ^ f_u_dadda_cla32_fa614_xor1;
  assign f_u_dadda_cla32_fa758_and1 = f_u_dadda_cla32_fa758_xor0 & f_u_dadda_cla32_fa614_xor1;
  assign f_u_dadda_cla32_fa758_or0 = f_u_dadda_cla32_fa758_and0 | f_u_dadda_cla32_fa758_and1;
  assign f_u_dadda_cla32_fa759_xor0 = f_u_dadda_cla32_fa615_xor1 ^ f_u_dadda_cla32_fa616_xor1;
  assign f_u_dadda_cla32_fa759_and0 = f_u_dadda_cla32_fa615_xor1 & f_u_dadda_cla32_fa616_xor1;
  assign f_u_dadda_cla32_fa759_xor1 = f_u_dadda_cla32_fa759_xor0 ^ f_u_dadda_cla32_fa617_xor1;
  assign f_u_dadda_cla32_fa759_and1 = f_u_dadda_cla32_fa759_xor0 & f_u_dadda_cla32_fa617_xor1;
  assign f_u_dadda_cla32_fa759_or0 = f_u_dadda_cla32_fa759_and0 | f_u_dadda_cla32_fa759_and1;
  assign f_u_dadda_cla32_fa760_xor0 = f_u_dadda_cla32_fa759_or0 ^ f_u_dadda_cla32_fa758_or0;
  assign f_u_dadda_cla32_fa760_and0 = f_u_dadda_cla32_fa759_or0 & f_u_dadda_cla32_fa758_or0;
  assign f_u_dadda_cla32_fa760_xor1 = f_u_dadda_cla32_fa760_xor0 ^ f_u_dadda_cla32_fa624_xor1;
  assign f_u_dadda_cla32_fa760_and1 = f_u_dadda_cla32_fa760_xor0 & f_u_dadda_cla32_fa624_xor1;
  assign f_u_dadda_cla32_fa760_or0 = f_u_dadda_cla32_fa760_and0 | f_u_dadda_cla32_fa760_and1;
  assign f_u_dadda_cla32_fa761_xor0 = f_u_dadda_cla32_fa625_xor1 ^ f_u_dadda_cla32_fa626_xor1;
  assign f_u_dadda_cla32_fa761_and0 = f_u_dadda_cla32_fa625_xor1 & f_u_dadda_cla32_fa626_xor1;
  assign f_u_dadda_cla32_fa761_xor1 = f_u_dadda_cla32_fa761_xor0 ^ f_u_dadda_cla32_fa627_xor1;
  assign f_u_dadda_cla32_fa761_and1 = f_u_dadda_cla32_fa761_xor0 & f_u_dadda_cla32_fa627_xor1;
  assign f_u_dadda_cla32_fa761_or0 = f_u_dadda_cla32_fa761_and0 | f_u_dadda_cla32_fa761_and1;
  assign f_u_dadda_cla32_fa762_xor0 = f_u_dadda_cla32_fa761_or0 ^ f_u_dadda_cla32_fa760_or0;
  assign f_u_dadda_cla32_fa762_and0 = f_u_dadda_cla32_fa761_or0 & f_u_dadda_cla32_fa760_or0;
  assign f_u_dadda_cla32_fa762_xor1 = f_u_dadda_cla32_fa762_xor0 ^ f_u_dadda_cla32_fa633_xor1;
  assign f_u_dadda_cla32_fa762_and1 = f_u_dadda_cla32_fa762_xor0 & f_u_dadda_cla32_fa633_xor1;
  assign f_u_dadda_cla32_fa762_or0 = f_u_dadda_cla32_fa762_and0 | f_u_dadda_cla32_fa762_and1;
  assign f_u_dadda_cla32_fa763_xor0 = f_u_dadda_cla32_fa634_xor1 ^ f_u_dadda_cla32_fa635_xor1;
  assign f_u_dadda_cla32_fa763_and0 = f_u_dadda_cla32_fa634_xor1 & f_u_dadda_cla32_fa635_xor1;
  assign f_u_dadda_cla32_fa763_xor1 = f_u_dadda_cla32_fa763_xor0 ^ f_u_dadda_cla32_fa636_xor1;
  assign f_u_dadda_cla32_fa763_and1 = f_u_dadda_cla32_fa763_xor0 & f_u_dadda_cla32_fa636_xor1;
  assign f_u_dadda_cla32_fa763_or0 = f_u_dadda_cla32_fa763_and0 | f_u_dadda_cla32_fa763_and1;
  assign f_u_dadda_cla32_fa764_xor0 = f_u_dadda_cla32_fa763_or0 ^ f_u_dadda_cla32_fa762_or0;
  assign f_u_dadda_cla32_fa764_and0 = f_u_dadda_cla32_fa763_or0 & f_u_dadda_cla32_fa762_or0;
  assign f_u_dadda_cla32_fa764_xor1 = f_u_dadda_cla32_fa764_xor0 ^ f_u_dadda_cla32_fa641_xor1;
  assign f_u_dadda_cla32_fa764_and1 = f_u_dadda_cla32_fa764_xor0 & f_u_dadda_cla32_fa641_xor1;
  assign f_u_dadda_cla32_fa764_or0 = f_u_dadda_cla32_fa764_and0 | f_u_dadda_cla32_fa764_and1;
  assign f_u_dadda_cla32_fa765_xor0 = f_u_dadda_cla32_fa642_xor1 ^ f_u_dadda_cla32_fa643_xor1;
  assign f_u_dadda_cla32_fa765_and0 = f_u_dadda_cla32_fa642_xor1 & f_u_dadda_cla32_fa643_xor1;
  assign f_u_dadda_cla32_fa765_xor1 = f_u_dadda_cla32_fa765_xor0 ^ f_u_dadda_cla32_fa644_xor1;
  assign f_u_dadda_cla32_fa765_and1 = f_u_dadda_cla32_fa765_xor0 & f_u_dadda_cla32_fa644_xor1;
  assign f_u_dadda_cla32_fa765_or0 = f_u_dadda_cla32_fa765_and0 | f_u_dadda_cla32_fa765_and1;
  assign f_u_dadda_cla32_fa766_xor0 = f_u_dadda_cla32_fa765_or0 ^ f_u_dadda_cla32_fa764_or0;
  assign f_u_dadda_cla32_fa766_and0 = f_u_dadda_cla32_fa765_or0 & f_u_dadda_cla32_fa764_or0;
  assign f_u_dadda_cla32_fa766_xor1 = f_u_dadda_cla32_fa766_xor0 ^ f_u_dadda_cla32_fa648_xor1;
  assign f_u_dadda_cla32_fa766_and1 = f_u_dadda_cla32_fa766_xor0 & f_u_dadda_cla32_fa648_xor1;
  assign f_u_dadda_cla32_fa766_or0 = f_u_dadda_cla32_fa766_and0 | f_u_dadda_cla32_fa766_and1;
  assign f_u_dadda_cla32_fa767_xor0 = f_u_dadda_cla32_fa649_xor1 ^ f_u_dadda_cla32_fa650_xor1;
  assign f_u_dadda_cla32_fa767_and0 = f_u_dadda_cla32_fa649_xor1 & f_u_dadda_cla32_fa650_xor1;
  assign f_u_dadda_cla32_fa767_xor1 = f_u_dadda_cla32_fa767_xor0 ^ f_u_dadda_cla32_fa651_xor1;
  assign f_u_dadda_cla32_fa767_and1 = f_u_dadda_cla32_fa767_xor0 & f_u_dadda_cla32_fa651_xor1;
  assign f_u_dadda_cla32_fa767_or0 = f_u_dadda_cla32_fa767_and0 | f_u_dadda_cla32_fa767_and1;
  assign f_u_dadda_cla32_fa768_xor0 = f_u_dadda_cla32_fa767_or0 ^ f_u_dadda_cla32_fa766_or0;
  assign f_u_dadda_cla32_fa768_and0 = f_u_dadda_cla32_fa767_or0 & f_u_dadda_cla32_fa766_or0;
  assign f_u_dadda_cla32_fa768_xor1 = f_u_dadda_cla32_fa768_xor0 ^ f_u_dadda_cla32_fa654_xor1;
  assign f_u_dadda_cla32_fa768_and1 = f_u_dadda_cla32_fa768_xor0 & f_u_dadda_cla32_fa654_xor1;
  assign f_u_dadda_cla32_fa768_or0 = f_u_dadda_cla32_fa768_and0 | f_u_dadda_cla32_fa768_and1;
  assign f_u_dadda_cla32_fa769_xor0 = f_u_dadda_cla32_fa655_xor1 ^ f_u_dadda_cla32_fa656_xor1;
  assign f_u_dadda_cla32_fa769_and0 = f_u_dadda_cla32_fa655_xor1 & f_u_dadda_cla32_fa656_xor1;
  assign f_u_dadda_cla32_fa769_xor1 = f_u_dadda_cla32_fa769_xor0 ^ f_u_dadda_cla32_fa657_xor1;
  assign f_u_dadda_cla32_fa769_and1 = f_u_dadda_cla32_fa769_xor0 & f_u_dadda_cla32_fa657_xor1;
  assign f_u_dadda_cla32_fa769_or0 = f_u_dadda_cla32_fa769_and0 | f_u_dadda_cla32_fa769_and1;
  assign f_u_dadda_cla32_and_22_31 = a[22] & b[31];
  assign f_u_dadda_cla32_fa770_xor0 = f_u_dadda_cla32_fa769_or0 ^ f_u_dadda_cla32_fa768_or0;
  assign f_u_dadda_cla32_fa770_and0 = f_u_dadda_cla32_fa769_or0 & f_u_dadda_cla32_fa768_or0;
  assign f_u_dadda_cla32_fa770_xor1 = f_u_dadda_cla32_fa770_xor0 ^ f_u_dadda_cla32_and_22_31;
  assign f_u_dadda_cla32_fa770_and1 = f_u_dadda_cla32_fa770_xor0 & f_u_dadda_cla32_and_22_31;
  assign f_u_dadda_cla32_fa770_or0 = f_u_dadda_cla32_fa770_and0 | f_u_dadda_cla32_fa770_and1;
  assign f_u_dadda_cla32_fa771_xor0 = f_u_dadda_cla32_fa660_xor1 ^ f_u_dadda_cla32_fa661_xor1;
  assign f_u_dadda_cla32_fa771_and0 = f_u_dadda_cla32_fa660_xor1 & f_u_dadda_cla32_fa661_xor1;
  assign f_u_dadda_cla32_fa771_xor1 = f_u_dadda_cla32_fa771_xor0 ^ f_u_dadda_cla32_fa662_xor1;
  assign f_u_dadda_cla32_fa771_and1 = f_u_dadda_cla32_fa771_xor0 & f_u_dadda_cla32_fa662_xor1;
  assign f_u_dadda_cla32_fa771_or0 = f_u_dadda_cla32_fa771_and0 | f_u_dadda_cla32_fa771_and1;
  assign f_u_dadda_cla32_and_24_30 = a[24] & b[30];
  assign f_u_dadda_cla32_fa772_xor0 = f_u_dadda_cla32_fa771_or0 ^ f_u_dadda_cla32_fa770_or0;
  assign f_u_dadda_cla32_fa772_and0 = f_u_dadda_cla32_fa771_or0 & f_u_dadda_cla32_fa770_or0;
  assign f_u_dadda_cla32_fa772_xor1 = f_u_dadda_cla32_fa772_xor0 ^ f_u_dadda_cla32_and_24_30;
  assign f_u_dadda_cla32_fa772_and1 = f_u_dadda_cla32_fa772_xor0 & f_u_dadda_cla32_and_24_30;
  assign f_u_dadda_cla32_fa772_or0 = f_u_dadda_cla32_fa772_and0 | f_u_dadda_cla32_fa772_and1;
  assign f_u_dadda_cla32_and_23_31 = a[23] & b[31];
  assign f_u_dadda_cla32_fa773_xor0 = f_u_dadda_cla32_and_23_31 ^ f_u_dadda_cla32_fa665_xor1;
  assign f_u_dadda_cla32_fa773_and0 = f_u_dadda_cla32_and_23_31 & f_u_dadda_cla32_fa665_xor1;
  assign f_u_dadda_cla32_fa773_xor1 = f_u_dadda_cla32_fa773_xor0 ^ f_u_dadda_cla32_fa666_xor1;
  assign f_u_dadda_cla32_fa773_and1 = f_u_dadda_cla32_fa773_xor0 & f_u_dadda_cla32_fa666_xor1;
  assign f_u_dadda_cla32_fa773_or0 = f_u_dadda_cla32_fa773_and0 | f_u_dadda_cla32_fa773_and1;
  assign f_u_dadda_cla32_and_26_29 = a[26] & b[29];
  assign f_u_dadda_cla32_fa774_xor0 = f_u_dadda_cla32_fa773_or0 ^ f_u_dadda_cla32_fa772_or0;
  assign f_u_dadda_cla32_fa774_and0 = f_u_dadda_cla32_fa773_or0 & f_u_dadda_cla32_fa772_or0;
  assign f_u_dadda_cla32_fa774_xor1 = f_u_dadda_cla32_fa774_xor0 ^ f_u_dadda_cla32_and_26_29;
  assign f_u_dadda_cla32_fa774_and1 = f_u_dadda_cla32_fa774_xor0 & f_u_dadda_cla32_and_26_29;
  assign f_u_dadda_cla32_fa774_or0 = f_u_dadda_cla32_fa774_and0 | f_u_dadda_cla32_fa774_and1;
  assign f_u_dadda_cla32_and_25_30 = a[25] & b[30];
  assign f_u_dadda_cla32_and_24_31 = a[24] & b[31];
  assign f_u_dadda_cla32_fa775_xor0 = f_u_dadda_cla32_and_25_30 ^ f_u_dadda_cla32_and_24_31;
  assign f_u_dadda_cla32_fa775_and0 = f_u_dadda_cla32_and_25_30 & f_u_dadda_cla32_and_24_31;
  assign f_u_dadda_cla32_fa775_xor1 = f_u_dadda_cla32_fa775_xor0 ^ f_u_dadda_cla32_fa669_xor1;
  assign f_u_dadda_cla32_fa775_and1 = f_u_dadda_cla32_fa775_xor0 & f_u_dadda_cla32_fa669_xor1;
  assign f_u_dadda_cla32_fa775_or0 = f_u_dadda_cla32_fa775_and0 | f_u_dadda_cla32_fa775_and1;
  assign f_u_dadda_cla32_and_28_28 = a[28] & b[28];
  assign f_u_dadda_cla32_fa776_xor0 = f_u_dadda_cla32_fa775_or0 ^ f_u_dadda_cla32_fa774_or0;
  assign f_u_dadda_cla32_fa776_and0 = f_u_dadda_cla32_fa775_or0 & f_u_dadda_cla32_fa774_or0;
  assign f_u_dadda_cla32_fa776_xor1 = f_u_dadda_cla32_fa776_xor0 ^ f_u_dadda_cla32_and_28_28;
  assign f_u_dadda_cla32_fa776_and1 = f_u_dadda_cla32_fa776_xor0 & f_u_dadda_cla32_and_28_28;
  assign f_u_dadda_cla32_fa776_or0 = f_u_dadda_cla32_fa776_and0 | f_u_dadda_cla32_fa776_and1;
  assign f_u_dadda_cla32_and_27_29 = a[27] & b[29];
  assign f_u_dadda_cla32_and_26_30 = a[26] & b[30];
  assign f_u_dadda_cla32_and_25_31 = a[25] & b[31];
  assign f_u_dadda_cla32_fa777_xor0 = f_u_dadda_cla32_and_27_29 ^ f_u_dadda_cla32_and_26_30;
  assign f_u_dadda_cla32_fa777_and0 = f_u_dadda_cla32_and_27_29 & f_u_dadda_cla32_and_26_30;
  assign f_u_dadda_cla32_fa777_xor1 = f_u_dadda_cla32_fa777_xor0 ^ f_u_dadda_cla32_and_25_31;
  assign f_u_dadda_cla32_fa777_and1 = f_u_dadda_cla32_fa777_xor0 & f_u_dadda_cla32_and_25_31;
  assign f_u_dadda_cla32_fa777_or0 = f_u_dadda_cla32_fa777_and0 | f_u_dadda_cla32_fa777_and1;
  assign f_u_dadda_cla32_and_30_27 = a[30] & b[27];
  assign f_u_dadda_cla32_fa778_xor0 = f_u_dadda_cla32_fa777_or0 ^ f_u_dadda_cla32_fa776_or0;
  assign f_u_dadda_cla32_fa778_and0 = f_u_dadda_cla32_fa777_or0 & f_u_dadda_cla32_fa776_or0;
  assign f_u_dadda_cla32_fa778_xor1 = f_u_dadda_cla32_fa778_xor0 ^ f_u_dadda_cla32_and_30_27;
  assign f_u_dadda_cla32_fa778_and1 = f_u_dadda_cla32_fa778_xor0 & f_u_dadda_cla32_and_30_27;
  assign f_u_dadda_cla32_fa778_or0 = f_u_dadda_cla32_fa778_and0 | f_u_dadda_cla32_fa778_and1;
  assign f_u_dadda_cla32_and_29_28 = a[29] & b[28];
  assign f_u_dadda_cla32_and_28_29 = a[28] & b[29];
  assign f_u_dadda_cla32_and_27_30 = a[27] & b[30];
  assign f_u_dadda_cla32_fa779_xor0 = f_u_dadda_cla32_and_29_28 ^ f_u_dadda_cla32_and_28_29;
  assign f_u_dadda_cla32_fa779_and0 = f_u_dadda_cla32_and_29_28 & f_u_dadda_cla32_and_28_29;
  assign f_u_dadda_cla32_fa779_xor1 = f_u_dadda_cla32_fa779_xor0 ^ f_u_dadda_cla32_and_27_30;
  assign f_u_dadda_cla32_fa779_and1 = f_u_dadda_cla32_fa779_xor0 & f_u_dadda_cla32_and_27_30;
  assign f_u_dadda_cla32_fa779_or0 = f_u_dadda_cla32_fa779_and0 | f_u_dadda_cla32_fa779_and1;
  assign f_u_dadda_cla32_fa780_xor0 = f_u_dadda_cla32_fa779_or0 ^ f_u_dadda_cla32_fa778_or0;
  assign f_u_dadda_cla32_fa780_and0 = f_u_dadda_cla32_fa779_or0 & f_u_dadda_cla32_fa778_or0;
  assign f_u_dadda_cla32_fa780_xor1 = f_u_dadda_cla32_fa780_xor0 ^ f_u_dadda_cla32_fa674_or0;
  assign f_u_dadda_cla32_fa780_and1 = f_u_dadda_cla32_fa780_xor0 & f_u_dadda_cla32_fa674_or0;
  assign f_u_dadda_cla32_fa780_or0 = f_u_dadda_cla32_fa780_and0 | f_u_dadda_cla32_fa780_and1;
  assign f_u_dadda_cla32_and_31_27 = a[31] & b[27];
  assign f_u_dadda_cla32_and_30_28 = a[30] & b[28];
  assign f_u_dadda_cla32_and_29_29 = a[29] & b[29];
  assign f_u_dadda_cla32_fa781_xor0 = f_u_dadda_cla32_and_31_27 ^ f_u_dadda_cla32_and_30_28;
  assign f_u_dadda_cla32_fa781_and0 = f_u_dadda_cla32_and_31_27 & f_u_dadda_cla32_and_30_28;
  assign f_u_dadda_cla32_fa781_xor1 = f_u_dadda_cla32_fa781_xor0 ^ f_u_dadda_cla32_and_29_29;
  assign f_u_dadda_cla32_fa781_and1 = f_u_dadda_cla32_fa781_xor0 & f_u_dadda_cla32_and_29_29;
  assign f_u_dadda_cla32_fa781_or0 = f_u_dadda_cla32_fa781_and0 | f_u_dadda_cla32_fa781_and1;
  assign f_u_dadda_cla32_and_31_28 = a[31] & b[28];
  assign f_u_dadda_cla32_fa782_xor0 = f_u_dadda_cla32_fa781_or0 ^ f_u_dadda_cla32_fa780_or0;
  assign f_u_dadda_cla32_fa782_and0 = f_u_dadda_cla32_fa781_or0 & f_u_dadda_cla32_fa780_or0;
  assign f_u_dadda_cla32_fa782_xor1 = f_u_dadda_cla32_fa782_xor0 ^ f_u_dadda_cla32_and_31_28;
  assign f_u_dadda_cla32_fa782_and1 = f_u_dadda_cla32_fa782_xor0 & f_u_dadda_cla32_and_31_28;
  assign f_u_dadda_cla32_fa782_or0 = f_u_dadda_cla32_fa782_and0 | f_u_dadda_cla32_fa782_and1;
  assign f_u_dadda_cla32_and_3_0 = a[3] & b[0];
  assign f_u_dadda_cla32_and_2_1 = a[2] & b[1];
  assign f_u_dadda_cla32_ha29_xor0 = f_u_dadda_cla32_and_3_0 ^ f_u_dadda_cla32_and_2_1;
  assign f_u_dadda_cla32_ha29_and0 = f_u_dadda_cla32_and_3_0 & f_u_dadda_cla32_and_2_1;
  assign f_u_dadda_cla32_and_2_2 = a[2] & b[2];
  assign f_u_dadda_cla32_and_1_3 = a[1] & b[3];
  assign f_u_dadda_cla32_fa783_xor0 = f_u_dadda_cla32_ha29_and0 ^ f_u_dadda_cla32_and_2_2;
  assign f_u_dadda_cla32_fa783_and0 = f_u_dadda_cla32_ha29_and0 & f_u_dadda_cla32_and_2_2;
  assign f_u_dadda_cla32_fa783_xor1 = f_u_dadda_cla32_fa783_xor0 ^ f_u_dadda_cla32_and_1_3;
  assign f_u_dadda_cla32_fa783_and1 = f_u_dadda_cla32_fa783_xor0 & f_u_dadda_cla32_and_1_3;
  assign f_u_dadda_cla32_fa783_or0 = f_u_dadda_cla32_fa783_and0 | f_u_dadda_cla32_fa783_and1;
  assign f_u_dadda_cla32_and_1_4 = a[1] & b[4];
  assign f_u_dadda_cla32_and_0_5 = a[0] & b[5];
  assign f_u_dadda_cla32_fa784_xor0 = f_u_dadda_cla32_fa783_or0 ^ f_u_dadda_cla32_and_1_4;
  assign f_u_dadda_cla32_fa784_and0 = f_u_dadda_cla32_fa783_or0 & f_u_dadda_cla32_and_1_4;
  assign f_u_dadda_cla32_fa784_xor1 = f_u_dadda_cla32_fa784_xor0 ^ f_u_dadda_cla32_and_0_5;
  assign f_u_dadda_cla32_fa784_and1 = f_u_dadda_cla32_fa784_xor0 & f_u_dadda_cla32_and_0_5;
  assign f_u_dadda_cla32_fa784_or0 = f_u_dadda_cla32_fa784_and0 | f_u_dadda_cla32_fa784_and1;
  assign f_u_dadda_cla32_and_0_6 = a[0] & b[6];
  assign f_u_dadda_cla32_fa785_xor0 = f_u_dadda_cla32_fa784_or0 ^ f_u_dadda_cla32_and_0_6;
  assign f_u_dadda_cla32_fa785_and0 = f_u_dadda_cla32_fa784_or0 & f_u_dadda_cla32_and_0_6;
  assign f_u_dadda_cla32_fa785_xor1 = f_u_dadda_cla32_fa785_xor0 ^ f_u_dadda_cla32_ha5_xor0;
  assign f_u_dadda_cla32_fa785_and1 = f_u_dadda_cla32_fa785_xor0 & f_u_dadda_cla32_ha5_xor0;
  assign f_u_dadda_cla32_fa785_or0 = f_u_dadda_cla32_fa785_and0 | f_u_dadda_cla32_fa785_and1;
  assign f_u_dadda_cla32_fa786_xor0 = f_u_dadda_cla32_fa785_or0 ^ f_u_dadda_cla32_fa15_xor1;
  assign f_u_dadda_cla32_fa786_and0 = f_u_dadda_cla32_fa785_or0 & f_u_dadda_cla32_fa15_xor1;
  assign f_u_dadda_cla32_fa786_xor1 = f_u_dadda_cla32_fa786_xor0 ^ f_u_dadda_cla32_ha6_xor0;
  assign f_u_dadda_cla32_fa786_and1 = f_u_dadda_cla32_fa786_xor0 & f_u_dadda_cla32_ha6_xor0;
  assign f_u_dadda_cla32_fa786_or0 = f_u_dadda_cla32_fa786_and0 | f_u_dadda_cla32_fa786_and1;
  assign f_u_dadda_cla32_fa787_xor0 = f_u_dadda_cla32_fa786_or0 ^ f_u_dadda_cla32_fa17_xor1;
  assign f_u_dadda_cla32_fa787_and0 = f_u_dadda_cla32_fa786_or0 & f_u_dadda_cla32_fa17_xor1;
  assign f_u_dadda_cla32_fa787_xor1 = f_u_dadda_cla32_fa787_xor0 ^ f_u_dadda_cla32_ha7_xor0;
  assign f_u_dadda_cla32_fa787_and1 = f_u_dadda_cla32_fa787_xor0 & f_u_dadda_cla32_ha7_xor0;
  assign f_u_dadda_cla32_fa787_or0 = f_u_dadda_cla32_fa787_and0 | f_u_dadda_cla32_fa787_and1;
  assign f_u_dadda_cla32_fa788_xor0 = f_u_dadda_cla32_fa787_or0 ^ f_u_dadda_cla32_fa20_xor1;
  assign f_u_dadda_cla32_fa788_and0 = f_u_dadda_cla32_fa787_or0 & f_u_dadda_cla32_fa20_xor1;
  assign f_u_dadda_cla32_fa788_xor1 = f_u_dadda_cla32_fa788_xor0 ^ f_u_dadda_cla32_ha8_xor0;
  assign f_u_dadda_cla32_fa788_and1 = f_u_dadda_cla32_fa788_xor0 & f_u_dadda_cla32_ha8_xor0;
  assign f_u_dadda_cla32_fa788_or0 = f_u_dadda_cla32_fa788_and0 | f_u_dadda_cla32_fa788_and1;
  assign f_u_dadda_cla32_fa789_xor0 = f_u_dadda_cla32_fa788_or0 ^ f_u_dadda_cla32_fa24_xor1;
  assign f_u_dadda_cla32_fa789_and0 = f_u_dadda_cla32_fa788_or0 & f_u_dadda_cla32_fa24_xor1;
  assign f_u_dadda_cla32_fa789_xor1 = f_u_dadda_cla32_fa789_xor0 ^ f_u_dadda_cla32_ha9_xor0;
  assign f_u_dadda_cla32_fa789_and1 = f_u_dadda_cla32_fa789_xor0 & f_u_dadda_cla32_ha9_xor0;
  assign f_u_dadda_cla32_fa789_or0 = f_u_dadda_cla32_fa789_and0 | f_u_dadda_cla32_fa789_and1;
  assign f_u_dadda_cla32_fa790_xor0 = f_u_dadda_cla32_fa789_or0 ^ f_u_dadda_cla32_fa29_xor1;
  assign f_u_dadda_cla32_fa790_and0 = f_u_dadda_cla32_fa789_or0 & f_u_dadda_cla32_fa29_xor1;
  assign f_u_dadda_cla32_fa790_xor1 = f_u_dadda_cla32_fa790_xor0 ^ f_u_dadda_cla32_ha10_xor0;
  assign f_u_dadda_cla32_fa790_and1 = f_u_dadda_cla32_fa790_xor0 & f_u_dadda_cla32_ha10_xor0;
  assign f_u_dadda_cla32_fa790_or0 = f_u_dadda_cla32_fa790_and0 | f_u_dadda_cla32_fa790_and1;
  assign f_u_dadda_cla32_fa791_xor0 = f_u_dadda_cla32_fa790_or0 ^ f_u_dadda_cla32_fa35_xor1;
  assign f_u_dadda_cla32_fa791_and0 = f_u_dadda_cla32_fa790_or0 & f_u_dadda_cla32_fa35_xor1;
  assign f_u_dadda_cla32_fa791_xor1 = f_u_dadda_cla32_fa791_xor0 ^ f_u_dadda_cla32_ha11_xor0;
  assign f_u_dadda_cla32_fa791_and1 = f_u_dadda_cla32_fa791_xor0 & f_u_dadda_cla32_ha11_xor0;
  assign f_u_dadda_cla32_fa791_or0 = f_u_dadda_cla32_fa791_and0 | f_u_dadda_cla32_fa791_and1;
  assign f_u_dadda_cla32_fa792_xor0 = f_u_dadda_cla32_fa791_or0 ^ f_u_dadda_cla32_fa42_xor1;
  assign f_u_dadda_cla32_fa792_and0 = f_u_dadda_cla32_fa791_or0 & f_u_dadda_cla32_fa42_xor1;
  assign f_u_dadda_cla32_fa792_xor1 = f_u_dadda_cla32_fa792_xor0 ^ f_u_dadda_cla32_ha12_xor0;
  assign f_u_dadda_cla32_fa792_and1 = f_u_dadda_cla32_fa792_xor0 & f_u_dadda_cla32_ha12_xor0;
  assign f_u_dadda_cla32_fa792_or0 = f_u_dadda_cla32_fa792_and0 | f_u_dadda_cla32_fa792_and1;
  assign f_u_dadda_cla32_fa793_xor0 = f_u_dadda_cla32_fa792_or0 ^ f_u_dadda_cla32_fa50_xor1;
  assign f_u_dadda_cla32_fa793_and0 = f_u_dadda_cla32_fa792_or0 & f_u_dadda_cla32_fa50_xor1;
  assign f_u_dadda_cla32_fa793_xor1 = f_u_dadda_cla32_fa793_xor0 ^ f_u_dadda_cla32_ha13_xor0;
  assign f_u_dadda_cla32_fa793_and1 = f_u_dadda_cla32_fa793_xor0 & f_u_dadda_cla32_ha13_xor0;
  assign f_u_dadda_cla32_fa793_or0 = f_u_dadda_cla32_fa793_and0 | f_u_dadda_cla32_fa793_and1;
  assign f_u_dadda_cla32_fa794_xor0 = f_u_dadda_cla32_fa793_or0 ^ f_u_dadda_cla32_fa59_xor1;
  assign f_u_dadda_cla32_fa794_and0 = f_u_dadda_cla32_fa793_or0 & f_u_dadda_cla32_fa59_xor1;
  assign f_u_dadda_cla32_fa794_xor1 = f_u_dadda_cla32_fa794_xor0 ^ f_u_dadda_cla32_ha14_xor0;
  assign f_u_dadda_cla32_fa794_and1 = f_u_dadda_cla32_fa794_xor0 & f_u_dadda_cla32_ha14_xor0;
  assign f_u_dadda_cla32_fa794_or0 = f_u_dadda_cla32_fa794_and0 | f_u_dadda_cla32_fa794_and1;
  assign f_u_dadda_cla32_fa795_xor0 = f_u_dadda_cla32_fa794_or0 ^ f_u_dadda_cla32_fa69_xor1;
  assign f_u_dadda_cla32_fa795_and0 = f_u_dadda_cla32_fa794_or0 & f_u_dadda_cla32_fa69_xor1;
  assign f_u_dadda_cla32_fa795_xor1 = f_u_dadda_cla32_fa795_xor0 ^ f_u_dadda_cla32_ha15_xor0;
  assign f_u_dadda_cla32_fa795_and1 = f_u_dadda_cla32_fa795_xor0 & f_u_dadda_cla32_ha15_xor0;
  assign f_u_dadda_cla32_fa795_or0 = f_u_dadda_cla32_fa795_and0 | f_u_dadda_cla32_fa795_and1;
  assign f_u_dadda_cla32_fa796_xor0 = f_u_dadda_cla32_fa795_or0 ^ f_u_dadda_cla32_fa80_xor1;
  assign f_u_dadda_cla32_fa796_and0 = f_u_dadda_cla32_fa795_or0 & f_u_dadda_cla32_fa80_xor1;
  assign f_u_dadda_cla32_fa796_xor1 = f_u_dadda_cla32_fa796_xor0 ^ f_u_dadda_cla32_ha16_xor0;
  assign f_u_dadda_cla32_fa796_and1 = f_u_dadda_cla32_fa796_xor0 & f_u_dadda_cla32_ha16_xor0;
  assign f_u_dadda_cla32_fa796_or0 = f_u_dadda_cla32_fa796_and0 | f_u_dadda_cla32_fa796_and1;
  assign f_u_dadda_cla32_fa797_xor0 = f_u_dadda_cla32_fa796_or0 ^ f_u_dadda_cla32_fa92_xor1;
  assign f_u_dadda_cla32_fa797_and0 = f_u_dadda_cla32_fa796_or0 & f_u_dadda_cla32_fa92_xor1;
  assign f_u_dadda_cla32_fa797_xor1 = f_u_dadda_cla32_fa797_xor0 ^ f_u_dadda_cla32_ha17_xor0;
  assign f_u_dadda_cla32_fa797_and1 = f_u_dadda_cla32_fa797_xor0 & f_u_dadda_cla32_ha17_xor0;
  assign f_u_dadda_cla32_fa797_or0 = f_u_dadda_cla32_fa797_and0 | f_u_dadda_cla32_fa797_and1;
  assign f_u_dadda_cla32_fa798_xor0 = f_u_dadda_cla32_fa797_or0 ^ f_u_dadda_cla32_fa105_xor1;
  assign f_u_dadda_cla32_fa798_and0 = f_u_dadda_cla32_fa797_or0 & f_u_dadda_cla32_fa105_xor1;
  assign f_u_dadda_cla32_fa798_xor1 = f_u_dadda_cla32_fa798_xor0 ^ f_u_dadda_cla32_ha18_xor0;
  assign f_u_dadda_cla32_fa798_and1 = f_u_dadda_cla32_fa798_xor0 & f_u_dadda_cla32_ha18_xor0;
  assign f_u_dadda_cla32_fa798_or0 = f_u_dadda_cla32_fa798_and0 | f_u_dadda_cla32_fa798_and1;
  assign f_u_dadda_cla32_fa799_xor0 = f_u_dadda_cla32_fa798_or0 ^ f_u_dadda_cla32_fa119_xor1;
  assign f_u_dadda_cla32_fa799_and0 = f_u_dadda_cla32_fa798_or0 & f_u_dadda_cla32_fa119_xor1;
  assign f_u_dadda_cla32_fa799_xor1 = f_u_dadda_cla32_fa799_xor0 ^ f_u_dadda_cla32_ha19_xor0;
  assign f_u_dadda_cla32_fa799_and1 = f_u_dadda_cla32_fa799_xor0 & f_u_dadda_cla32_ha19_xor0;
  assign f_u_dadda_cla32_fa799_or0 = f_u_dadda_cla32_fa799_and0 | f_u_dadda_cla32_fa799_and1;
  assign f_u_dadda_cla32_fa800_xor0 = f_u_dadda_cla32_fa799_or0 ^ f_u_dadda_cla32_fa134_xor1;
  assign f_u_dadda_cla32_fa800_and0 = f_u_dadda_cla32_fa799_or0 & f_u_dadda_cla32_fa134_xor1;
  assign f_u_dadda_cla32_fa800_xor1 = f_u_dadda_cla32_fa800_xor0 ^ f_u_dadda_cla32_ha20_xor0;
  assign f_u_dadda_cla32_fa800_and1 = f_u_dadda_cla32_fa800_xor0 & f_u_dadda_cla32_ha20_xor0;
  assign f_u_dadda_cla32_fa800_or0 = f_u_dadda_cla32_fa800_and0 | f_u_dadda_cla32_fa800_and1;
  assign f_u_dadda_cla32_fa801_xor0 = f_u_dadda_cla32_fa800_or0 ^ f_u_dadda_cla32_fa150_xor1;
  assign f_u_dadda_cla32_fa801_and0 = f_u_dadda_cla32_fa800_or0 & f_u_dadda_cla32_fa150_xor1;
  assign f_u_dadda_cla32_fa801_xor1 = f_u_dadda_cla32_fa801_xor0 ^ f_u_dadda_cla32_ha21_xor0;
  assign f_u_dadda_cla32_fa801_and1 = f_u_dadda_cla32_fa801_xor0 & f_u_dadda_cla32_ha21_xor0;
  assign f_u_dadda_cla32_fa801_or0 = f_u_dadda_cla32_fa801_and0 | f_u_dadda_cla32_fa801_and1;
  assign f_u_dadda_cla32_fa802_xor0 = f_u_dadda_cla32_fa801_or0 ^ f_u_dadda_cla32_fa167_xor1;
  assign f_u_dadda_cla32_fa802_and0 = f_u_dadda_cla32_fa801_or0 & f_u_dadda_cla32_fa167_xor1;
  assign f_u_dadda_cla32_fa802_xor1 = f_u_dadda_cla32_fa802_xor0 ^ f_u_dadda_cla32_ha22_xor0;
  assign f_u_dadda_cla32_fa802_and1 = f_u_dadda_cla32_fa802_xor0 & f_u_dadda_cla32_ha22_xor0;
  assign f_u_dadda_cla32_fa802_or0 = f_u_dadda_cla32_fa802_and0 | f_u_dadda_cla32_fa802_and1;
  assign f_u_dadda_cla32_fa803_xor0 = f_u_dadda_cla32_fa802_or0 ^ f_u_dadda_cla32_fa185_xor1;
  assign f_u_dadda_cla32_fa803_and0 = f_u_dadda_cla32_fa802_or0 & f_u_dadda_cla32_fa185_xor1;
  assign f_u_dadda_cla32_fa803_xor1 = f_u_dadda_cla32_fa803_xor0 ^ f_u_dadda_cla32_ha23_xor0;
  assign f_u_dadda_cla32_fa803_and1 = f_u_dadda_cla32_fa803_xor0 & f_u_dadda_cla32_ha23_xor0;
  assign f_u_dadda_cla32_fa803_or0 = f_u_dadda_cla32_fa803_and0 | f_u_dadda_cla32_fa803_and1;
  assign f_u_dadda_cla32_fa804_xor0 = f_u_dadda_cla32_fa803_or0 ^ f_u_dadda_cla32_fa204_xor1;
  assign f_u_dadda_cla32_fa804_and0 = f_u_dadda_cla32_fa803_or0 & f_u_dadda_cla32_fa204_xor1;
  assign f_u_dadda_cla32_fa804_xor1 = f_u_dadda_cla32_fa804_xor0 ^ f_u_dadda_cla32_ha24_xor0;
  assign f_u_dadda_cla32_fa804_and1 = f_u_dadda_cla32_fa804_xor0 & f_u_dadda_cla32_ha24_xor0;
  assign f_u_dadda_cla32_fa804_or0 = f_u_dadda_cla32_fa804_and0 | f_u_dadda_cla32_fa804_and1;
  assign f_u_dadda_cla32_fa805_xor0 = f_u_dadda_cla32_fa804_or0 ^ f_u_dadda_cla32_fa224_xor1;
  assign f_u_dadda_cla32_fa805_and0 = f_u_dadda_cla32_fa804_or0 & f_u_dadda_cla32_fa224_xor1;
  assign f_u_dadda_cla32_fa805_xor1 = f_u_dadda_cla32_fa805_xor0 ^ f_u_dadda_cla32_ha25_xor0;
  assign f_u_dadda_cla32_fa805_and1 = f_u_dadda_cla32_fa805_xor0 & f_u_dadda_cla32_ha25_xor0;
  assign f_u_dadda_cla32_fa805_or0 = f_u_dadda_cla32_fa805_and0 | f_u_dadda_cla32_fa805_and1;
  assign f_u_dadda_cla32_fa806_xor0 = f_u_dadda_cla32_fa805_or0 ^ f_u_dadda_cla32_fa245_xor1;
  assign f_u_dadda_cla32_fa806_and0 = f_u_dadda_cla32_fa805_or0 & f_u_dadda_cla32_fa245_xor1;
  assign f_u_dadda_cla32_fa806_xor1 = f_u_dadda_cla32_fa806_xor0 ^ f_u_dadda_cla32_ha26_xor0;
  assign f_u_dadda_cla32_fa806_and1 = f_u_dadda_cla32_fa806_xor0 & f_u_dadda_cla32_ha26_xor0;
  assign f_u_dadda_cla32_fa806_or0 = f_u_dadda_cla32_fa806_and0 | f_u_dadda_cla32_fa806_and1;
  assign f_u_dadda_cla32_fa807_xor0 = f_u_dadda_cla32_fa806_or0 ^ f_u_dadda_cla32_fa266_xor1;
  assign f_u_dadda_cla32_fa807_and0 = f_u_dadda_cla32_fa806_or0 & f_u_dadda_cla32_fa266_xor1;
  assign f_u_dadda_cla32_fa807_xor1 = f_u_dadda_cla32_fa807_xor0 ^ f_u_dadda_cla32_fa267_xor1;
  assign f_u_dadda_cla32_fa807_and1 = f_u_dadda_cla32_fa807_xor0 & f_u_dadda_cla32_fa267_xor1;
  assign f_u_dadda_cla32_fa807_or0 = f_u_dadda_cla32_fa807_and0 | f_u_dadda_cla32_fa807_and1;
  assign f_u_dadda_cla32_fa808_xor0 = f_u_dadda_cla32_fa807_or0 ^ f_u_dadda_cla32_fa288_xor1;
  assign f_u_dadda_cla32_fa808_and0 = f_u_dadda_cla32_fa807_or0 & f_u_dadda_cla32_fa288_xor1;
  assign f_u_dadda_cla32_fa808_xor1 = f_u_dadda_cla32_fa808_xor0 ^ f_u_dadda_cla32_fa289_xor1;
  assign f_u_dadda_cla32_fa808_and1 = f_u_dadda_cla32_fa808_xor0 & f_u_dadda_cla32_fa289_xor1;
  assign f_u_dadda_cla32_fa808_or0 = f_u_dadda_cla32_fa808_and0 | f_u_dadda_cla32_fa808_and1;
  assign f_u_dadda_cla32_fa809_xor0 = f_u_dadda_cla32_fa808_or0 ^ f_u_dadda_cla32_fa310_xor1;
  assign f_u_dadda_cla32_fa809_and0 = f_u_dadda_cla32_fa808_or0 & f_u_dadda_cla32_fa310_xor1;
  assign f_u_dadda_cla32_fa809_xor1 = f_u_dadda_cla32_fa809_xor0 ^ f_u_dadda_cla32_fa311_xor1;
  assign f_u_dadda_cla32_fa809_and1 = f_u_dadda_cla32_fa809_xor0 & f_u_dadda_cla32_fa311_xor1;
  assign f_u_dadda_cla32_fa809_or0 = f_u_dadda_cla32_fa809_and0 | f_u_dadda_cla32_fa809_and1;
  assign f_u_dadda_cla32_fa810_xor0 = f_u_dadda_cla32_fa809_or0 ^ f_u_dadda_cla32_fa332_xor1;
  assign f_u_dadda_cla32_fa810_and0 = f_u_dadda_cla32_fa809_or0 & f_u_dadda_cla32_fa332_xor1;
  assign f_u_dadda_cla32_fa810_xor1 = f_u_dadda_cla32_fa810_xor0 ^ f_u_dadda_cla32_fa333_xor1;
  assign f_u_dadda_cla32_fa810_and1 = f_u_dadda_cla32_fa810_xor0 & f_u_dadda_cla32_fa333_xor1;
  assign f_u_dadda_cla32_fa810_or0 = f_u_dadda_cla32_fa810_and0 | f_u_dadda_cla32_fa810_and1;
  assign f_u_dadda_cla32_fa811_xor0 = f_u_dadda_cla32_fa810_or0 ^ f_u_dadda_cla32_fa354_xor1;
  assign f_u_dadda_cla32_fa811_and0 = f_u_dadda_cla32_fa810_or0 & f_u_dadda_cla32_fa354_xor1;
  assign f_u_dadda_cla32_fa811_xor1 = f_u_dadda_cla32_fa811_xor0 ^ f_u_dadda_cla32_fa355_xor1;
  assign f_u_dadda_cla32_fa811_and1 = f_u_dadda_cla32_fa811_xor0 & f_u_dadda_cla32_fa355_xor1;
  assign f_u_dadda_cla32_fa811_or0 = f_u_dadda_cla32_fa811_and0 | f_u_dadda_cla32_fa811_and1;
  assign f_u_dadda_cla32_fa812_xor0 = f_u_dadda_cla32_fa811_or0 ^ f_u_dadda_cla32_fa376_xor1;
  assign f_u_dadda_cla32_fa812_and0 = f_u_dadda_cla32_fa811_or0 & f_u_dadda_cla32_fa376_xor1;
  assign f_u_dadda_cla32_fa812_xor1 = f_u_dadda_cla32_fa812_xor0 ^ f_u_dadda_cla32_fa377_xor1;
  assign f_u_dadda_cla32_fa812_and1 = f_u_dadda_cla32_fa812_xor0 & f_u_dadda_cla32_fa377_xor1;
  assign f_u_dadda_cla32_fa812_or0 = f_u_dadda_cla32_fa812_and0 | f_u_dadda_cla32_fa812_and1;
  assign f_u_dadda_cla32_fa813_xor0 = f_u_dadda_cla32_fa812_or0 ^ f_u_dadda_cla32_fa398_xor1;
  assign f_u_dadda_cla32_fa813_and0 = f_u_dadda_cla32_fa812_or0 & f_u_dadda_cla32_fa398_xor1;
  assign f_u_dadda_cla32_fa813_xor1 = f_u_dadda_cla32_fa813_xor0 ^ f_u_dadda_cla32_fa399_xor1;
  assign f_u_dadda_cla32_fa813_and1 = f_u_dadda_cla32_fa813_xor0 & f_u_dadda_cla32_fa399_xor1;
  assign f_u_dadda_cla32_fa813_or0 = f_u_dadda_cla32_fa813_and0 | f_u_dadda_cla32_fa813_and1;
  assign f_u_dadda_cla32_fa814_xor0 = f_u_dadda_cla32_fa813_or0 ^ f_u_dadda_cla32_fa420_xor1;
  assign f_u_dadda_cla32_fa814_and0 = f_u_dadda_cla32_fa813_or0 & f_u_dadda_cla32_fa420_xor1;
  assign f_u_dadda_cla32_fa814_xor1 = f_u_dadda_cla32_fa814_xor0 ^ f_u_dadda_cla32_fa421_xor1;
  assign f_u_dadda_cla32_fa814_and1 = f_u_dadda_cla32_fa814_xor0 & f_u_dadda_cla32_fa421_xor1;
  assign f_u_dadda_cla32_fa814_or0 = f_u_dadda_cla32_fa814_and0 | f_u_dadda_cla32_fa814_and1;
  assign f_u_dadda_cla32_fa815_xor0 = f_u_dadda_cla32_fa814_or0 ^ f_u_dadda_cla32_fa442_xor1;
  assign f_u_dadda_cla32_fa815_and0 = f_u_dadda_cla32_fa814_or0 & f_u_dadda_cla32_fa442_xor1;
  assign f_u_dadda_cla32_fa815_xor1 = f_u_dadda_cla32_fa815_xor0 ^ f_u_dadda_cla32_fa443_xor1;
  assign f_u_dadda_cla32_fa815_and1 = f_u_dadda_cla32_fa815_xor0 & f_u_dadda_cla32_fa443_xor1;
  assign f_u_dadda_cla32_fa815_or0 = f_u_dadda_cla32_fa815_and0 | f_u_dadda_cla32_fa815_and1;
  assign f_u_dadda_cla32_fa816_xor0 = f_u_dadda_cla32_fa815_or0 ^ f_u_dadda_cla32_fa463_xor1;
  assign f_u_dadda_cla32_fa816_and0 = f_u_dadda_cla32_fa815_or0 & f_u_dadda_cla32_fa463_xor1;
  assign f_u_dadda_cla32_fa816_xor1 = f_u_dadda_cla32_fa816_xor0 ^ f_u_dadda_cla32_fa464_xor1;
  assign f_u_dadda_cla32_fa816_and1 = f_u_dadda_cla32_fa816_xor0 & f_u_dadda_cla32_fa464_xor1;
  assign f_u_dadda_cla32_fa816_or0 = f_u_dadda_cla32_fa816_and0 | f_u_dadda_cla32_fa816_and1;
  assign f_u_dadda_cla32_fa817_xor0 = f_u_dadda_cla32_fa816_or0 ^ f_u_dadda_cla32_fa483_xor1;
  assign f_u_dadda_cla32_fa817_and0 = f_u_dadda_cla32_fa816_or0 & f_u_dadda_cla32_fa483_xor1;
  assign f_u_dadda_cla32_fa817_xor1 = f_u_dadda_cla32_fa817_xor0 ^ f_u_dadda_cla32_fa484_xor1;
  assign f_u_dadda_cla32_fa817_and1 = f_u_dadda_cla32_fa817_xor0 & f_u_dadda_cla32_fa484_xor1;
  assign f_u_dadda_cla32_fa817_or0 = f_u_dadda_cla32_fa817_and0 | f_u_dadda_cla32_fa817_and1;
  assign f_u_dadda_cla32_fa818_xor0 = f_u_dadda_cla32_fa817_or0 ^ f_u_dadda_cla32_fa502_xor1;
  assign f_u_dadda_cla32_fa818_and0 = f_u_dadda_cla32_fa817_or0 & f_u_dadda_cla32_fa502_xor1;
  assign f_u_dadda_cla32_fa818_xor1 = f_u_dadda_cla32_fa818_xor0 ^ f_u_dadda_cla32_fa503_xor1;
  assign f_u_dadda_cla32_fa818_and1 = f_u_dadda_cla32_fa818_xor0 & f_u_dadda_cla32_fa503_xor1;
  assign f_u_dadda_cla32_fa818_or0 = f_u_dadda_cla32_fa818_and0 | f_u_dadda_cla32_fa818_and1;
  assign f_u_dadda_cla32_fa819_xor0 = f_u_dadda_cla32_fa818_or0 ^ f_u_dadda_cla32_fa520_xor1;
  assign f_u_dadda_cla32_fa819_and0 = f_u_dadda_cla32_fa818_or0 & f_u_dadda_cla32_fa520_xor1;
  assign f_u_dadda_cla32_fa819_xor1 = f_u_dadda_cla32_fa819_xor0 ^ f_u_dadda_cla32_fa521_xor1;
  assign f_u_dadda_cla32_fa819_and1 = f_u_dadda_cla32_fa819_xor0 & f_u_dadda_cla32_fa521_xor1;
  assign f_u_dadda_cla32_fa819_or0 = f_u_dadda_cla32_fa819_and0 | f_u_dadda_cla32_fa819_and1;
  assign f_u_dadda_cla32_fa820_xor0 = f_u_dadda_cla32_fa819_or0 ^ f_u_dadda_cla32_fa537_xor1;
  assign f_u_dadda_cla32_fa820_and0 = f_u_dadda_cla32_fa819_or0 & f_u_dadda_cla32_fa537_xor1;
  assign f_u_dadda_cla32_fa820_xor1 = f_u_dadda_cla32_fa820_xor0 ^ f_u_dadda_cla32_fa538_xor1;
  assign f_u_dadda_cla32_fa820_and1 = f_u_dadda_cla32_fa820_xor0 & f_u_dadda_cla32_fa538_xor1;
  assign f_u_dadda_cla32_fa820_or0 = f_u_dadda_cla32_fa820_and0 | f_u_dadda_cla32_fa820_and1;
  assign f_u_dadda_cla32_fa821_xor0 = f_u_dadda_cla32_fa820_or0 ^ f_u_dadda_cla32_fa553_xor1;
  assign f_u_dadda_cla32_fa821_and0 = f_u_dadda_cla32_fa820_or0 & f_u_dadda_cla32_fa553_xor1;
  assign f_u_dadda_cla32_fa821_xor1 = f_u_dadda_cla32_fa821_xor0 ^ f_u_dadda_cla32_fa554_xor1;
  assign f_u_dadda_cla32_fa821_and1 = f_u_dadda_cla32_fa821_xor0 & f_u_dadda_cla32_fa554_xor1;
  assign f_u_dadda_cla32_fa821_or0 = f_u_dadda_cla32_fa821_and0 | f_u_dadda_cla32_fa821_and1;
  assign f_u_dadda_cla32_fa822_xor0 = f_u_dadda_cla32_fa821_or0 ^ f_u_dadda_cla32_fa568_xor1;
  assign f_u_dadda_cla32_fa822_and0 = f_u_dadda_cla32_fa821_or0 & f_u_dadda_cla32_fa568_xor1;
  assign f_u_dadda_cla32_fa822_xor1 = f_u_dadda_cla32_fa822_xor0 ^ f_u_dadda_cla32_fa569_xor1;
  assign f_u_dadda_cla32_fa822_and1 = f_u_dadda_cla32_fa822_xor0 & f_u_dadda_cla32_fa569_xor1;
  assign f_u_dadda_cla32_fa822_or0 = f_u_dadda_cla32_fa822_and0 | f_u_dadda_cla32_fa822_and1;
  assign f_u_dadda_cla32_fa823_xor0 = f_u_dadda_cla32_fa822_or0 ^ f_u_dadda_cla32_fa582_xor1;
  assign f_u_dadda_cla32_fa823_and0 = f_u_dadda_cla32_fa822_or0 & f_u_dadda_cla32_fa582_xor1;
  assign f_u_dadda_cla32_fa823_xor1 = f_u_dadda_cla32_fa823_xor0 ^ f_u_dadda_cla32_fa583_xor1;
  assign f_u_dadda_cla32_fa823_and1 = f_u_dadda_cla32_fa823_xor0 & f_u_dadda_cla32_fa583_xor1;
  assign f_u_dadda_cla32_fa823_or0 = f_u_dadda_cla32_fa823_and0 | f_u_dadda_cla32_fa823_and1;
  assign f_u_dadda_cla32_fa824_xor0 = f_u_dadda_cla32_fa823_or0 ^ f_u_dadda_cla32_fa595_xor1;
  assign f_u_dadda_cla32_fa824_and0 = f_u_dadda_cla32_fa823_or0 & f_u_dadda_cla32_fa595_xor1;
  assign f_u_dadda_cla32_fa824_xor1 = f_u_dadda_cla32_fa824_xor0 ^ f_u_dadda_cla32_fa596_xor1;
  assign f_u_dadda_cla32_fa824_and1 = f_u_dadda_cla32_fa824_xor0 & f_u_dadda_cla32_fa596_xor1;
  assign f_u_dadda_cla32_fa824_or0 = f_u_dadda_cla32_fa824_and0 | f_u_dadda_cla32_fa824_and1;
  assign f_u_dadda_cla32_fa825_xor0 = f_u_dadda_cla32_fa824_or0 ^ f_u_dadda_cla32_fa607_xor1;
  assign f_u_dadda_cla32_fa825_and0 = f_u_dadda_cla32_fa824_or0 & f_u_dadda_cla32_fa607_xor1;
  assign f_u_dadda_cla32_fa825_xor1 = f_u_dadda_cla32_fa825_xor0 ^ f_u_dadda_cla32_fa608_xor1;
  assign f_u_dadda_cla32_fa825_and1 = f_u_dadda_cla32_fa825_xor0 & f_u_dadda_cla32_fa608_xor1;
  assign f_u_dadda_cla32_fa825_or0 = f_u_dadda_cla32_fa825_and0 | f_u_dadda_cla32_fa825_and1;
  assign f_u_dadda_cla32_fa826_xor0 = f_u_dadda_cla32_fa825_or0 ^ f_u_dadda_cla32_fa618_xor1;
  assign f_u_dadda_cla32_fa826_and0 = f_u_dadda_cla32_fa825_or0 & f_u_dadda_cla32_fa618_xor1;
  assign f_u_dadda_cla32_fa826_xor1 = f_u_dadda_cla32_fa826_xor0 ^ f_u_dadda_cla32_fa619_xor1;
  assign f_u_dadda_cla32_fa826_and1 = f_u_dadda_cla32_fa826_xor0 & f_u_dadda_cla32_fa619_xor1;
  assign f_u_dadda_cla32_fa826_or0 = f_u_dadda_cla32_fa826_and0 | f_u_dadda_cla32_fa826_and1;
  assign f_u_dadda_cla32_fa827_xor0 = f_u_dadda_cla32_fa826_or0 ^ f_u_dadda_cla32_fa628_xor1;
  assign f_u_dadda_cla32_fa827_and0 = f_u_dadda_cla32_fa826_or0 & f_u_dadda_cla32_fa628_xor1;
  assign f_u_dadda_cla32_fa827_xor1 = f_u_dadda_cla32_fa827_xor0 ^ f_u_dadda_cla32_fa629_xor1;
  assign f_u_dadda_cla32_fa827_and1 = f_u_dadda_cla32_fa827_xor0 & f_u_dadda_cla32_fa629_xor1;
  assign f_u_dadda_cla32_fa827_or0 = f_u_dadda_cla32_fa827_and0 | f_u_dadda_cla32_fa827_and1;
  assign f_u_dadda_cla32_fa828_xor0 = f_u_dadda_cla32_fa827_or0 ^ f_u_dadda_cla32_fa637_xor1;
  assign f_u_dadda_cla32_fa828_and0 = f_u_dadda_cla32_fa827_or0 & f_u_dadda_cla32_fa637_xor1;
  assign f_u_dadda_cla32_fa828_xor1 = f_u_dadda_cla32_fa828_xor0 ^ f_u_dadda_cla32_fa638_xor1;
  assign f_u_dadda_cla32_fa828_and1 = f_u_dadda_cla32_fa828_xor0 & f_u_dadda_cla32_fa638_xor1;
  assign f_u_dadda_cla32_fa828_or0 = f_u_dadda_cla32_fa828_and0 | f_u_dadda_cla32_fa828_and1;
  assign f_u_dadda_cla32_fa829_xor0 = f_u_dadda_cla32_fa828_or0 ^ f_u_dadda_cla32_fa645_xor1;
  assign f_u_dadda_cla32_fa829_and0 = f_u_dadda_cla32_fa828_or0 & f_u_dadda_cla32_fa645_xor1;
  assign f_u_dadda_cla32_fa829_xor1 = f_u_dadda_cla32_fa829_xor0 ^ f_u_dadda_cla32_fa646_xor1;
  assign f_u_dadda_cla32_fa829_and1 = f_u_dadda_cla32_fa829_xor0 & f_u_dadda_cla32_fa646_xor1;
  assign f_u_dadda_cla32_fa829_or0 = f_u_dadda_cla32_fa829_and0 | f_u_dadda_cla32_fa829_and1;
  assign f_u_dadda_cla32_fa830_xor0 = f_u_dadda_cla32_fa829_or0 ^ f_u_dadda_cla32_fa652_xor1;
  assign f_u_dadda_cla32_fa830_and0 = f_u_dadda_cla32_fa829_or0 & f_u_dadda_cla32_fa652_xor1;
  assign f_u_dadda_cla32_fa830_xor1 = f_u_dadda_cla32_fa830_xor0 ^ f_u_dadda_cla32_fa653_xor1;
  assign f_u_dadda_cla32_fa830_and1 = f_u_dadda_cla32_fa830_xor0 & f_u_dadda_cla32_fa653_xor1;
  assign f_u_dadda_cla32_fa830_or0 = f_u_dadda_cla32_fa830_and0 | f_u_dadda_cla32_fa830_and1;
  assign f_u_dadda_cla32_fa831_xor0 = f_u_dadda_cla32_fa830_or0 ^ f_u_dadda_cla32_fa658_xor1;
  assign f_u_dadda_cla32_fa831_and0 = f_u_dadda_cla32_fa830_or0 & f_u_dadda_cla32_fa658_xor1;
  assign f_u_dadda_cla32_fa831_xor1 = f_u_dadda_cla32_fa831_xor0 ^ f_u_dadda_cla32_fa659_xor1;
  assign f_u_dadda_cla32_fa831_and1 = f_u_dadda_cla32_fa831_xor0 & f_u_dadda_cla32_fa659_xor1;
  assign f_u_dadda_cla32_fa831_or0 = f_u_dadda_cla32_fa831_and0 | f_u_dadda_cla32_fa831_and1;
  assign f_u_dadda_cla32_fa832_xor0 = f_u_dadda_cla32_fa831_or0 ^ f_u_dadda_cla32_fa663_xor1;
  assign f_u_dadda_cla32_fa832_and0 = f_u_dadda_cla32_fa831_or0 & f_u_dadda_cla32_fa663_xor1;
  assign f_u_dadda_cla32_fa832_xor1 = f_u_dadda_cla32_fa832_xor0 ^ f_u_dadda_cla32_fa664_xor1;
  assign f_u_dadda_cla32_fa832_and1 = f_u_dadda_cla32_fa832_xor0 & f_u_dadda_cla32_fa664_xor1;
  assign f_u_dadda_cla32_fa832_or0 = f_u_dadda_cla32_fa832_and0 | f_u_dadda_cla32_fa832_and1;
  assign f_u_dadda_cla32_fa833_xor0 = f_u_dadda_cla32_fa832_or0 ^ f_u_dadda_cla32_fa667_xor1;
  assign f_u_dadda_cla32_fa833_and0 = f_u_dadda_cla32_fa832_or0 & f_u_dadda_cla32_fa667_xor1;
  assign f_u_dadda_cla32_fa833_xor1 = f_u_dadda_cla32_fa833_xor0 ^ f_u_dadda_cla32_fa668_xor1;
  assign f_u_dadda_cla32_fa833_and1 = f_u_dadda_cla32_fa833_xor0 & f_u_dadda_cla32_fa668_xor1;
  assign f_u_dadda_cla32_fa833_or0 = f_u_dadda_cla32_fa833_and0 | f_u_dadda_cla32_fa833_and1;
  assign f_u_dadda_cla32_fa834_xor0 = f_u_dadda_cla32_fa833_or0 ^ f_u_dadda_cla32_fa670_xor1;
  assign f_u_dadda_cla32_fa834_and0 = f_u_dadda_cla32_fa833_or0 & f_u_dadda_cla32_fa670_xor1;
  assign f_u_dadda_cla32_fa834_xor1 = f_u_dadda_cla32_fa834_xor0 ^ f_u_dadda_cla32_fa671_xor1;
  assign f_u_dadda_cla32_fa834_and1 = f_u_dadda_cla32_fa834_xor0 & f_u_dadda_cla32_fa671_xor1;
  assign f_u_dadda_cla32_fa834_or0 = f_u_dadda_cla32_fa834_and0 | f_u_dadda_cla32_fa834_and1;
  assign f_u_dadda_cla32_fa835_xor0 = f_u_dadda_cla32_fa834_or0 ^ f_u_dadda_cla32_fa672_xor1;
  assign f_u_dadda_cla32_fa835_and0 = f_u_dadda_cla32_fa834_or0 & f_u_dadda_cla32_fa672_xor1;
  assign f_u_dadda_cla32_fa835_xor1 = f_u_dadda_cla32_fa835_xor0 ^ f_u_dadda_cla32_fa673_xor1;
  assign f_u_dadda_cla32_fa835_and1 = f_u_dadda_cla32_fa835_xor0 & f_u_dadda_cla32_fa673_xor1;
  assign f_u_dadda_cla32_fa835_or0 = f_u_dadda_cla32_fa835_and0 | f_u_dadda_cla32_fa835_and1;
  assign f_u_dadda_cla32_and_26_31 = a[26] & b[31];
  assign f_u_dadda_cla32_fa836_xor0 = f_u_dadda_cla32_fa835_or0 ^ f_u_dadda_cla32_and_26_31;
  assign f_u_dadda_cla32_fa836_and0 = f_u_dadda_cla32_fa835_or0 & f_u_dadda_cla32_and_26_31;
  assign f_u_dadda_cla32_fa836_xor1 = f_u_dadda_cla32_fa836_xor0 ^ f_u_dadda_cla32_fa674_xor1;
  assign f_u_dadda_cla32_fa836_and1 = f_u_dadda_cla32_fa836_xor0 & f_u_dadda_cla32_fa674_xor1;
  assign f_u_dadda_cla32_fa836_or0 = f_u_dadda_cla32_fa836_and0 | f_u_dadda_cla32_fa836_and1;
  assign f_u_dadda_cla32_and_28_30 = a[28] & b[30];
  assign f_u_dadda_cla32_and_27_31 = a[27] & b[31];
  assign f_u_dadda_cla32_fa837_xor0 = f_u_dadda_cla32_fa836_or0 ^ f_u_dadda_cla32_and_28_30;
  assign f_u_dadda_cla32_fa837_and0 = f_u_dadda_cla32_fa836_or0 & f_u_dadda_cla32_and_28_30;
  assign f_u_dadda_cla32_fa837_xor1 = f_u_dadda_cla32_fa837_xor0 ^ f_u_dadda_cla32_and_27_31;
  assign f_u_dadda_cla32_fa837_and1 = f_u_dadda_cla32_fa837_xor0 & f_u_dadda_cla32_and_27_31;
  assign f_u_dadda_cla32_fa837_or0 = f_u_dadda_cla32_fa837_and0 | f_u_dadda_cla32_fa837_and1;
  assign f_u_dadda_cla32_and_30_29 = a[30] & b[29];
  assign f_u_dadda_cla32_and_29_30 = a[29] & b[30];
  assign f_u_dadda_cla32_fa838_xor0 = f_u_dadda_cla32_fa837_or0 ^ f_u_dadda_cla32_and_30_29;
  assign f_u_dadda_cla32_fa838_and0 = f_u_dadda_cla32_fa837_or0 & f_u_dadda_cla32_and_30_29;
  assign f_u_dadda_cla32_fa838_xor1 = f_u_dadda_cla32_fa838_xor0 ^ f_u_dadda_cla32_and_29_30;
  assign f_u_dadda_cla32_fa838_and1 = f_u_dadda_cla32_fa838_xor0 & f_u_dadda_cla32_and_29_30;
  assign f_u_dadda_cla32_fa838_or0 = f_u_dadda_cla32_fa838_and0 | f_u_dadda_cla32_fa838_and1;
  assign f_u_dadda_cla32_and_31_29 = a[31] & b[29];
  assign f_u_dadda_cla32_fa839_xor0 = f_u_dadda_cla32_fa838_or0 ^ f_u_dadda_cla32_fa782_or0;
  assign f_u_dadda_cla32_fa839_and0 = f_u_dadda_cla32_fa838_or0 & f_u_dadda_cla32_fa782_or0;
  assign f_u_dadda_cla32_fa839_xor1 = f_u_dadda_cla32_fa839_xor0 ^ f_u_dadda_cla32_and_31_29;
  assign f_u_dadda_cla32_fa839_and1 = f_u_dadda_cla32_fa839_xor0 & f_u_dadda_cla32_and_31_29;
  assign f_u_dadda_cla32_fa839_or0 = f_u_dadda_cla32_fa839_and0 | f_u_dadda_cla32_fa839_and1;
  assign f_u_dadda_cla32_and_2_0 = a[2] & b[0];
  assign f_u_dadda_cla32_and_1_1 = a[1] & b[1];
  assign f_u_dadda_cla32_ha30_xor0 = f_u_dadda_cla32_and_2_0 ^ f_u_dadda_cla32_and_1_1;
  assign f_u_dadda_cla32_ha30_and0 = f_u_dadda_cla32_and_2_0 & f_u_dadda_cla32_and_1_1;
  assign f_u_dadda_cla32_and_1_2 = a[1] & b[2];
  assign f_u_dadda_cla32_and_0_3 = a[0] & b[3];
  assign f_u_dadda_cla32_fa840_xor0 = f_u_dadda_cla32_ha30_and0 ^ f_u_dadda_cla32_and_1_2;
  assign f_u_dadda_cla32_fa840_and0 = f_u_dadda_cla32_ha30_and0 & f_u_dadda_cla32_and_1_2;
  assign f_u_dadda_cla32_fa840_xor1 = f_u_dadda_cla32_fa840_xor0 ^ f_u_dadda_cla32_and_0_3;
  assign f_u_dadda_cla32_fa840_and1 = f_u_dadda_cla32_fa840_xor0 & f_u_dadda_cla32_and_0_3;
  assign f_u_dadda_cla32_fa840_or0 = f_u_dadda_cla32_fa840_and0 | f_u_dadda_cla32_fa840_and1;
  assign f_u_dadda_cla32_and_0_4 = a[0] & b[4];
  assign f_u_dadda_cla32_fa841_xor0 = f_u_dadda_cla32_fa840_or0 ^ f_u_dadda_cla32_and_0_4;
  assign f_u_dadda_cla32_fa841_and0 = f_u_dadda_cla32_fa840_or0 & f_u_dadda_cla32_and_0_4;
  assign f_u_dadda_cla32_fa841_xor1 = f_u_dadda_cla32_fa841_xor0 ^ f_u_dadda_cla32_ha27_xor0;
  assign f_u_dadda_cla32_fa841_and1 = f_u_dadda_cla32_fa841_xor0 & f_u_dadda_cla32_ha27_xor0;
  assign f_u_dadda_cla32_fa841_or0 = f_u_dadda_cla32_fa841_and0 | f_u_dadda_cla32_fa841_and1;
  assign f_u_dadda_cla32_fa842_xor0 = f_u_dadda_cla32_fa841_or0 ^ f_u_dadda_cla32_fa675_xor1;
  assign f_u_dadda_cla32_fa842_and0 = f_u_dadda_cla32_fa841_or0 & f_u_dadda_cla32_fa675_xor1;
  assign f_u_dadda_cla32_fa842_xor1 = f_u_dadda_cla32_fa842_xor0 ^ f_u_dadda_cla32_ha28_xor0;
  assign f_u_dadda_cla32_fa842_and1 = f_u_dadda_cla32_fa842_xor0 & f_u_dadda_cla32_ha28_xor0;
  assign f_u_dadda_cla32_fa842_or0 = f_u_dadda_cla32_fa842_and0 | f_u_dadda_cla32_fa842_and1;
  assign f_u_dadda_cla32_fa843_xor0 = f_u_dadda_cla32_fa842_or0 ^ f_u_dadda_cla32_fa676_xor1;
  assign f_u_dadda_cla32_fa843_and0 = f_u_dadda_cla32_fa842_or0 & f_u_dadda_cla32_fa676_xor1;
  assign f_u_dadda_cla32_fa843_xor1 = f_u_dadda_cla32_fa843_xor0 ^ f_u_dadda_cla32_fa677_xor1;
  assign f_u_dadda_cla32_fa843_and1 = f_u_dadda_cla32_fa843_xor0 & f_u_dadda_cla32_fa677_xor1;
  assign f_u_dadda_cla32_fa843_or0 = f_u_dadda_cla32_fa843_and0 | f_u_dadda_cla32_fa843_and1;
  assign f_u_dadda_cla32_fa844_xor0 = f_u_dadda_cla32_fa843_or0 ^ f_u_dadda_cla32_fa678_xor1;
  assign f_u_dadda_cla32_fa844_and0 = f_u_dadda_cla32_fa843_or0 & f_u_dadda_cla32_fa678_xor1;
  assign f_u_dadda_cla32_fa844_xor1 = f_u_dadda_cla32_fa844_xor0 ^ f_u_dadda_cla32_fa679_xor1;
  assign f_u_dadda_cla32_fa844_and1 = f_u_dadda_cla32_fa844_xor0 & f_u_dadda_cla32_fa679_xor1;
  assign f_u_dadda_cla32_fa844_or0 = f_u_dadda_cla32_fa844_and0 | f_u_dadda_cla32_fa844_and1;
  assign f_u_dadda_cla32_fa845_xor0 = f_u_dadda_cla32_fa844_or0 ^ f_u_dadda_cla32_fa680_xor1;
  assign f_u_dadda_cla32_fa845_and0 = f_u_dadda_cla32_fa844_or0 & f_u_dadda_cla32_fa680_xor1;
  assign f_u_dadda_cla32_fa845_xor1 = f_u_dadda_cla32_fa845_xor0 ^ f_u_dadda_cla32_fa681_xor1;
  assign f_u_dadda_cla32_fa845_and1 = f_u_dadda_cla32_fa845_xor0 & f_u_dadda_cla32_fa681_xor1;
  assign f_u_dadda_cla32_fa845_or0 = f_u_dadda_cla32_fa845_and0 | f_u_dadda_cla32_fa845_and1;
  assign f_u_dadda_cla32_fa846_xor0 = f_u_dadda_cla32_fa845_or0 ^ f_u_dadda_cla32_fa682_xor1;
  assign f_u_dadda_cla32_fa846_and0 = f_u_dadda_cla32_fa845_or0 & f_u_dadda_cla32_fa682_xor1;
  assign f_u_dadda_cla32_fa846_xor1 = f_u_dadda_cla32_fa846_xor0 ^ f_u_dadda_cla32_fa683_xor1;
  assign f_u_dadda_cla32_fa846_and1 = f_u_dadda_cla32_fa846_xor0 & f_u_dadda_cla32_fa683_xor1;
  assign f_u_dadda_cla32_fa846_or0 = f_u_dadda_cla32_fa846_and0 | f_u_dadda_cla32_fa846_and1;
  assign f_u_dadda_cla32_fa847_xor0 = f_u_dadda_cla32_fa846_or0 ^ f_u_dadda_cla32_fa684_xor1;
  assign f_u_dadda_cla32_fa847_and0 = f_u_dadda_cla32_fa846_or0 & f_u_dadda_cla32_fa684_xor1;
  assign f_u_dadda_cla32_fa847_xor1 = f_u_dadda_cla32_fa847_xor0 ^ f_u_dadda_cla32_fa685_xor1;
  assign f_u_dadda_cla32_fa847_and1 = f_u_dadda_cla32_fa847_xor0 & f_u_dadda_cla32_fa685_xor1;
  assign f_u_dadda_cla32_fa847_or0 = f_u_dadda_cla32_fa847_and0 | f_u_dadda_cla32_fa847_and1;
  assign f_u_dadda_cla32_fa848_xor0 = f_u_dadda_cla32_fa847_or0 ^ f_u_dadda_cla32_fa686_xor1;
  assign f_u_dadda_cla32_fa848_and0 = f_u_dadda_cla32_fa847_or0 & f_u_dadda_cla32_fa686_xor1;
  assign f_u_dadda_cla32_fa848_xor1 = f_u_dadda_cla32_fa848_xor0 ^ f_u_dadda_cla32_fa687_xor1;
  assign f_u_dadda_cla32_fa848_and1 = f_u_dadda_cla32_fa848_xor0 & f_u_dadda_cla32_fa687_xor1;
  assign f_u_dadda_cla32_fa848_or0 = f_u_dadda_cla32_fa848_and0 | f_u_dadda_cla32_fa848_and1;
  assign f_u_dadda_cla32_fa849_xor0 = f_u_dadda_cla32_fa848_or0 ^ f_u_dadda_cla32_fa688_xor1;
  assign f_u_dadda_cla32_fa849_and0 = f_u_dadda_cla32_fa848_or0 & f_u_dadda_cla32_fa688_xor1;
  assign f_u_dadda_cla32_fa849_xor1 = f_u_dadda_cla32_fa849_xor0 ^ f_u_dadda_cla32_fa689_xor1;
  assign f_u_dadda_cla32_fa849_and1 = f_u_dadda_cla32_fa849_xor0 & f_u_dadda_cla32_fa689_xor1;
  assign f_u_dadda_cla32_fa849_or0 = f_u_dadda_cla32_fa849_and0 | f_u_dadda_cla32_fa849_and1;
  assign f_u_dadda_cla32_fa850_xor0 = f_u_dadda_cla32_fa849_or0 ^ f_u_dadda_cla32_fa690_xor1;
  assign f_u_dadda_cla32_fa850_and0 = f_u_dadda_cla32_fa849_or0 & f_u_dadda_cla32_fa690_xor1;
  assign f_u_dadda_cla32_fa850_xor1 = f_u_dadda_cla32_fa850_xor0 ^ f_u_dadda_cla32_fa691_xor1;
  assign f_u_dadda_cla32_fa850_and1 = f_u_dadda_cla32_fa850_xor0 & f_u_dadda_cla32_fa691_xor1;
  assign f_u_dadda_cla32_fa850_or0 = f_u_dadda_cla32_fa850_and0 | f_u_dadda_cla32_fa850_and1;
  assign f_u_dadda_cla32_fa851_xor0 = f_u_dadda_cla32_fa850_or0 ^ f_u_dadda_cla32_fa692_xor1;
  assign f_u_dadda_cla32_fa851_and0 = f_u_dadda_cla32_fa850_or0 & f_u_dadda_cla32_fa692_xor1;
  assign f_u_dadda_cla32_fa851_xor1 = f_u_dadda_cla32_fa851_xor0 ^ f_u_dadda_cla32_fa693_xor1;
  assign f_u_dadda_cla32_fa851_and1 = f_u_dadda_cla32_fa851_xor0 & f_u_dadda_cla32_fa693_xor1;
  assign f_u_dadda_cla32_fa851_or0 = f_u_dadda_cla32_fa851_and0 | f_u_dadda_cla32_fa851_and1;
  assign f_u_dadda_cla32_fa852_xor0 = f_u_dadda_cla32_fa851_or0 ^ f_u_dadda_cla32_fa694_xor1;
  assign f_u_dadda_cla32_fa852_and0 = f_u_dadda_cla32_fa851_or0 & f_u_dadda_cla32_fa694_xor1;
  assign f_u_dadda_cla32_fa852_xor1 = f_u_dadda_cla32_fa852_xor0 ^ f_u_dadda_cla32_fa695_xor1;
  assign f_u_dadda_cla32_fa852_and1 = f_u_dadda_cla32_fa852_xor0 & f_u_dadda_cla32_fa695_xor1;
  assign f_u_dadda_cla32_fa852_or0 = f_u_dadda_cla32_fa852_and0 | f_u_dadda_cla32_fa852_and1;
  assign f_u_dadda_cla32_fa853_xor0 = f_u_dadda_cla32_fa852_or0 ^ f_u_dadda_cla32_fa696_xor1;
  assign f_u_dadda_cla32_fa853_and0 = f_u_dadda_cla32_fa852_or0 & f_u_dadda_cla32_fa696_xor1;
  assign f_u_dadda_cla32_fa853_xor1 = f_u_dadda_cla32_fa853_xor0 ^ f_u_dadda_cla32_fa697_xor1;
  assign f_u_dadda_cla32_fa853_and1 = f_u_dadda_cla32_fa853_xor0 & f_u_dadda_cla32_fa697_xor1;
  assign f_u_dadda_cla32_fa853_or0 = f_u_dadda_cla32_fa853_and0 | f_u_dadda_cla32_fa853_and1;
  assign f_u_dadda_cla32_fa854_xor0 = f_u_dadda_cla32_fa853_or0 ^ f_u_dadda_cla32_fa698_xor1;
  assign f_u_dadda_cla32_fa854_and0 = f_u_dadda_cla32_fa853_or0 & f_u_dadda_cla32_fa698_xor1;
  assign f_u_dadda_cla32_fa854_xor1 = f_u_dadda_cla32_fa854_xor0 ^ f_u_dadda_cla32_fa699_xor1;
  assign f_u_dadda_cla32_fa854_and1 = f_u_dadda_cla32_fa854_xor0 & f_u_dadda_cla32_fa699_xor1;
  assign f_u_dadda_cla32_fa854_or0 = f_u_dadda_cla32_fa854_and0 | f_u_dadda_cla32_fa854_and1;
  assign f_u_dadda_cla32_fa855_xor0 = f_u_dadda_cla32_fa854_or0 ^ f_u_dadda_cla32_fa700_xor1;
  assign f_u_dadda_cla32_fa855_and0 = f_u_dadda_cla32_fa854_or0 & f_u_dadda_cla32_fa700_xor1;
  assign f_u_dadda_cla32_fa855_xor1 = f_u_dadda_cla32_fa855_xor0 ^ f_u_dadda_cla32_fa701_xor1;
  assign f_u_dadda_cla32_fa855_and1 = f_u_dadda_cla32_fa855_xor0 & f_u_dadda_cla32_fa701_xor1;
  assign f_u_dadda_cla32_fa855_or0 = f_u_dadda_cla32_fa855_and0 | f_u_dadda_cla32_fa855_and1;
  assign f_u_dadda_cla32_fa856_xor0 = f_u_dadda_cla32_fa855_or0 ^ f_u_dadda_cla32_fa702_xor1;
  assign f_u_dadda_cla32_fa856_and0 = f_u_dadda_cla32_fa855_or0 & f_u_dadda_cla32_fa702_xor1;
  assign f_u_dadda_cla32_fa856_xor1 = f_u_dadda_cla32_fa856_xor0 ^ f_u_dadda_cla32_fa703_xor1;
  assign f_u_dadda_cla32_fa856_and1 = f_u_dadda_cla32_fa856_xor0 & f_u_dadda_cla32_fa703_xor1;
  assign f_u_dadda_cla32_fa856_or0 = f_u_dadda_cla32_fa856_and0 | f_u_dadda_cla32_fa856_and1;
  assign f_u_dadda_cla32_fa857_xor0 = f_u_dadda_cla32_fa856_or0 ^ f_u_dadda_cla32_fa704_xor1;
  assign f_u_dadda_cla32_fa857_and0 = f_u_dadda_cla32_fa856_or0 & f_u_dadda_cla32_fa704_xor1;
  assign f_u_dadda_cla32_fa857_xor1 = f_u_dadda_cla32_fa857_xor0 ^ f_u_dadda_cla32_fa705_xor1;
  assign f_u_dadda_cla32_fa857_and1 = f_u_dadda_cla32_fa857_xor0 & f_u_dadda_cla32_fa705_xor1;
  assign f_u_dadda_cla32_fa857_or0 = f_u_dadda_cla32_fa857_and0 | f_u_dadda_cla32_fa857_and1;
  assign f_u_dadda_cla32_fa858_xor0 = f_u_dadda_cla32_fa857_or0 ^ f_u_dadda_cla32_fa706_xor1;
  assign f_u_dadda_cla32_fa858_and0 = f_u_dadda_cla32_fa857_or0 & f_u_dadda_cla32_fa706_xor1;
  assign f_u_dadda_cla32_fa858_xor1 = f_u_dadda_cla32_fa858_xor0 ^ f_u_dadda_cla32_fa707_xor1;
  assign f_u_dadda_cla32_fa858_and1 = f_u_dadda_cla32_fa858_xor0 & f_u_dadda_cla32_fa707_xor1;
  assign f_u_dadda_cla32_fa858_or0 = f_u_dadda_cla32_fa858_and0 | f_u_dadda_cla32_fa858_and1;
  assign f_u_dadda_cla32_fa859_xor0 = f_u_dadda_cla32_fa858_or0 ^ f_u_dadda_cla32_fa708_xor1;
  assign f_u_dadda_cla32_fa859_and0 = f_u_dadda_cla32_fa858_or0 & f_u_dadda_cla32_fa708_xor1;
  assign f_u_dadda_cla32_fa859_xor1 = f_u_dadda_cla32_fa859_xor0 ^ f_u_dadda_cla32_fa709_xor1;
  assign f_u_dadda_cla32_fa859_and1 = f_u_dadda_cla32_fa859_xor0 & f_u_dadda_cla32_fa709_xor1;
  assign f_u_dadda_cla32_fa859_or0 = f_u_dadda_cla32_fa859_and0 | f_u_dadda_cla32_fa859_and1;
  assign f_u_dadda_cla32_fa860_xor0 = f_u_dadda_cla32_fa859_or0 ^ f_u_dadda_cla32_fa710_xor1;
  assign f_u_dadda_cla32_fa860_and0 = f_u_dadda_cla32_fa859_or0 & f_u_dadda_cla32_fa710_xor1;
  assign f_u_dadda_cla32_fa860_xor1 = f_u_dadda_cla32_fa860_xor0 ^ f_u_dadda_cla32_fa711_xor1;
  assign f_u_dadda_cla32_fa860_and1 = f_u_dadda_cla32_fa860_xor0 & f_u_dadda_cla32_fa711_xor1;
  assign f_u_dadda_cla32_fa860_or0 = f_u_dadda_cla32_fa860_and0 | f_u_dadda_cla32_fa860_and1;
  assign f_u_dadda_cla32_fa861_xor0 = f_u_dadda_cla32_fa860_or0 ^ f_u_dadda_cla32_fa712_xor1;
  assign f_u_dadda_cla32_fa861_and0 = f_u_dadda_cla32_fa860_or0 & f_u_dadda_cla32_fa712_xor1;
  assign f_u_dadda_cla32_fa861_xor1 = f_u_dadda_cla32_fa861_xor0 ^ f_u_dadda_cla32_fa713_xor1;
  assign f_u_dadda_cla32_fa861_and1 = f_u_dadda_cla32_fa861_xor0 & f_u_dadda_cla32_fa713_xor1;
  assign f_u_dadda_cla32_fa861_or0 = f_u_dadda_cla32_fa861_and0 | f_u_dadda_cla32_fa861_and1;
  assign f_u_dadda_cla32_fa862_xor0 = f_u_dadda_cla32_fa861_or0 ^ f_u_dadda_cla32_fa714_xor1;
  assign f_u_dadda_cla32_fa862_and0 = f_u_dadda_cla32_fa861_or0 & f_u_dadda_cla32_fa714_xor1;
  assign f_u_dadda_cla32_fa862_xor1 = f_u_dadda_cla32_fa862_xor0 ^ f_u_dadda_cla32_fa715_xor1;
  assign f_u_dadda_cla32_fa862_and1 = f_u_dadda_cla32_fa862_xor0 & f_u_dadda_cla32_fa715_xor1;
  assign f_u_dadda_cla32_fa862_or0 = f_u_dadda_cla32_fa862_and0 | f_u_dadda_cla32_fa862_and1;
  assign f_u_dadda_cla32_fa863_xor0 = f_u_dadda_cla32_fa862_or0 ^ f_u_dadda_cla32_fa716_xor1;
  assign f_u_dadda_cla32_fa863_and0 = f_u_dadda_cla32_fa862_or0 & f_u_dadda_cla32_fa716_xor1;
  assign f_u_dadda_cla32_fa863_xor1 = f_u_dadda_cla32_fa863_xor0 ^ f_u_dadda_cla32_fa717_xor1;
  assign f_u_dadda_cla32_fa863_and1 = f_u_dadda_cla32_fa863_xor0 & f_u_dadda_cla32_fa717_xor1;
  assign f_u_dadda_cla32_fa863_or0 = f_u_dadda_cla32_fa863_and0 | f_u_dadda_cla32_fa863_and1;
  assign f_u_dadda_cla32_fa864_xor0 = f_u_dadda_cla32_fa863_or0 ^ f_u_dadda_cla32_fa718_xor1;
  assign f_u_dadda_cla32_fa864_and0 = f_u_dadda_cla32_fa863_or0 & f_u_dadda_cla32_fa718_xor1;
  assign f_u_dadda_cla32_fa864_xor1 = f_u_dadda_cla32_fa864_xor0 ^ f_u_dadda_cla32_fa719_xor1;
  assign f_u_dadda_cla32_fa864_and1 = f_u_dadda_cla32_fa864_xor0 & f_u_dadda_cla32_fa719_xor1;
  assign f_u_dadda_cla32_fa864_or0 = f_u_dadda_cla32_fa864_and0 | f_u_dadda_cla32_fa864_and1;
  assign f_u_dadda_cla32_fa865_xor0 = f_u_dadda_cla32_fa864_or0 ^ f_u_dadda_cla32_fa720_xor1;
  assign f_u_dadda_cla32_fa865_and0 = f_u_dadda_cla32_fa864_or0 & f_u_dadda_cla32_fa720_xor1;
  assign f_u_dadda_cla32_fa865_xor1 = f_u_dadda_cla32_fa865_xor0 ^ f_u_dadda_cla32_fa721_xor1;
  assign f_u_dadda_cla32_fa865_and1 = f_u_dadda_cla32_fa865_xor0 & f_u_dadda_cla32_fa721_xor1;
  assign f_u_dadda_cla32_fa865_or0 = f_u_dadda_cla32_fa865_and0 | f_u_dadda_cla32_fa865_and1;
  assign f_u_dadda_cla32_fa866_xor0 = f_u_dadda_cla32_fa865_or0 ^ f_u_dadda_cla32_fa722_xor1;
  assign f_u_dadda_cla32_fa866_and0 = f_u_dadda_cla32_fa865_or0 & f_u_dadda_cla32_fa722_xor1;
  assign f_u_dadda_cla32_fa866_xor1 = f_u_dadda_cla32_fa866_xor0 ^ f_u_dadda_cla32_fa723_xor1;
  assign f_u_dadda_cla32_fa866_and1 = f_u_dadda_cla32_fa866_xor0 & f_u_dadda_cla32_fa723_xor1;
  assign f_u_dadda_cla32_fa866_or0 = f_u_dadda_cla32_fa866_and0 | f_u_dadda_cla32_fa866_and1;
  assign f_u_dadda_cla32_fa867_xor0 = f_u_dadda_cla32_fa866_or0 ^ f_u_dadda_cla32_fa724_xor1;
  assign f_u_dadda_cla32_fa867_and0 = f_u_dadda_cla32_fa866_or0 & f_u_dadda_cla32_fa724_xor1;
  assign f_u_dadda_cla32_fa867_xor1 = f_u_dadda_cla32_fa867_xor0 ^ f_u_dadda_cla32_fa725_xor1;
  assign f_u_dadda_cla32_fa867_and1 = f_u_dadda_cla32_fa867_xor0 & f_u_dadda_cla32_fa725_xor1;
  assign f_u_dadda_cla32_fa867_or0 = f_u_dadda_cla32_fa867_and0 | f_u_dadda_cla32_fa867_and1;
  assign f_u_dadda_cla32_fa868_xor0 = f_u_dadda_cla32_fa867_or0 ^ f_u_dadda_cla32_fa726_xor1;
  assign f_u_dadda_cla32_fa868_and0 = f_u_dadda_cla32_fa867_or0 & f_u_dadda_cla32_fa726_xor1;
  assign f_u_dadda_cla32_fa868_xor1 = f_u_dadda_cla32_fa868_xor0 ^ f_u_dadda_cla32_fa727_xor1;
  assign f_u_dadda_cla32_fa868_and1 = f_u_dadda_cla32_fa868_xor0 & f_u_dadda_cla32_fa727_xor1;
  assign f_u_dadda_cla32_fa868_or0 = f_u_dadda_cla32_fa868_and0 | f_u_dadda_cla32_fa868_and1;
  assign f_u_dadda_cla32_fa869_xor0 = f_u_dadda_cla32_fa868_or0 ^ f_u_dadda_cla32_fa728_xor1;
  assign f_u_dadda_cla32_fa869_and0 = f_u_dadda_cla32_fa868_or0 & f_u_dadda_cla32_fa728_xor1;
  assign f_u_dadda_cla32_fa869_xor1 = f_u_dadda_cla32_fa869_xor0 ^ f_u_dadda_cla32_fa729_xor1;
  assign f_u_dadda_cla32_fa869_and1 = f_u_dadda_cla32_fa869_xor0 & f_u_dadda_cla32_fa729_xor1;
  assign f_u_dadda_cla32_fa869_or0 = f_u_dadda_cla32_fa869_and0 | f_u_dadda_cla32_fa869_and1;
  assign f_u_dadda_cla32_fa870_xor0 = f_u_dadda_cla32_fa869_or0 ^ f_u_dadda_cla32_fa730_xor1;
  assign f_u_dadda_cla32_fa870_and0 = f_u_dadda_cla32_fa869_or0 & f_u_dadda_cla32_fa730_xor1;
  assign f_u_dadda_cla32_fa870_xor1 = f_u_dadda_cla32_fa870_xor0 ^ f_u_dadda_cla32_fa731_xor1;
  assign f_u_dadda_cla32_fa870_and1 = f_u_dadda_cla32_fa870_xor0 & f_u_dadda_cla32_fa731_xor1;
  assign f_u_dadda_cla32_fa870_or0 = f_u_dadda_cla32_fa870_and0 | f_u_dadda_cla32_fa870_and1;
  assign f_u_dadda_cla32_fa871_xor0 = f_u_dadda_cla32_fa870_or0 ^ f_u_dadda_cla32_fa732_xor1;
  assign f_u_dadda_cla32_fa871_and0 = f_u_dadda_cla32_fa870_or0 & f_u_dadda_cla32_fa732_xor1;
  assign f_u_dadda_cla32_fa871_xor1 = f_u_dadda_cla32_fa871_xor0 ^ f_u_dadda_cla32_fa733_xor1;
  assign f_u_dadda_cla32_fa871_and1 = f_u_dadda_cla32_fa871_xor0 & f_u_dadda_cla32_fa733_xor1;
  assign f_u_dadda_cla32_fa871_or0 = f_u_dadda_cla32_fa871_and0 | f_u_dadda_cla32_fa871_and1;
  assign f_u_dadda_cla32_fa872_xor0 = f_u_dadda_cla32_fa871_or0 ^ f_u_dadda_cla32_fa734_xor1;
  assign f_u_dadda_cla32_fa872_and0 = f_u_dadda_cla32_fa871_or0 & f_u_dadda_cla32_fa734_xor1;
  assign f_u_dadda_cla32_fa872_xor1 = f_u_dadda_cla32_fa872_xor0 ^ f_u_dadda_cla32_fa735_xor1;
  assign f_u_dadda_cla32_fa872_and1 = f_u_dadda_cla32_fa872_xor0 & f_u_dadda_cla32_fa735_xor1;
  assign f_u_dadda_cla32_fa872_or0 = f_u_dadda_cla32_fa872_and0 | f_u_dadda_cla32_fa872_and1;
  assign f_u_dadda_cla32_fa873_xor0 = f_u_dadda_cla32_fa872_or0 ^ f_u_dadda_cla32_fa736_xor1;
  assign f_u_dadda_cla32_fa873_and0 = f_u_dadda_cla32_fa872_or0 & f_u_dadda_cla32_fa736_xor1;
  assign f_u_dadda_cla32_fa873_xor1 = f_u_dadda_cla32_fa873_xor0 ^ f_u_dadda_cla32_fa737_xor1;
  assign f_u_dadda_cla32_fa873_and1 = f_u_dadda_cla32_fa873_xor0 & f_u_dadda_cla32_fa737_xor1;
  assign f_u_dadda_cla32_fa873_or0 = f_u_dadda_cla32_fa873_and0 | f_u_dadda_cla32_fa873_and1;
  assign f_u_dadda_cla32_fa874_xor0 = f_u_dadda_cla32_fa873_or0 ^ f_u_dadda_cla32_fa738_xor1;
  assign f_u_dadda_cla32_fa874_and0 = f_u_dadda_cla32_fa873_or0 & f_u_dadda_cla32_fa738_xor1;
  assign f_u_dadda_cla32_fa874_xor1 = f_u_dadda_cla32_fa874_xor0 ^ f_u_dadda_cla32_fa739_xor1;
  assign f_u_dadda_cla32_fa874_and1 = f_u_dadda_cla32_fa874_xor0 & f_u_dadda_cla32_fa739_xor1;
  assign f_u_dadda_cla32_fa874_or0 = f_u_dadda_cla32_fa874_and0 | f_u_dadda_cla32_fa874_and1;
  assign f_u_dadda_cla32_fa875_xor0 = f_u_dadda_cla32_fa874_or0 ^ f_u_dadda_cla32_fa740_xor1;
  assign f_u_dadda_cla32_fa875_and0 = f_u_dadda_cla32_fa874_or0 & f_u_dadda_cla32_fa740_xor1;
  assign f_u_dadda_cla32_fa875_xor1 = f_u_dadda_cla32_fa875_xor0 ^ f_u_dadda_cla32_fa741_xor1;
  assign f_u_dadda_cla32_fa875_and1 = f_u_dadda_cla32_fa875_xor0 & f_u_dadda_cla32_fa741_xor1;
  assign f_u_dadda_cla32_fa875_or0 = f_u_dadda_cla32_fa875_and0 | f_u_dadda_cla32_fa875_and1;
  assign f_u_dadda_cla32_fa876_xor0 = f_u_dadda_cla32_fa875_or0 ^ f_u_dadda_cla32_fa742_xor1;
  assign f_u_dadda_cla32_fa876_and0 = f_u_dadda_cla32_fa875_or0 & f_u_dadda_cla32_fa742_xor1;
  assign f_u_dadda_cla32_fa876_xor1 = f_u_dadda_cla32_fa876_xor0 ^ f_u_dadda_cla32_fa743_xor1;
  assign f_u_dadda_cla32_fa876_and1 = f_u_dadda_cla32_fa876_xor0 & f_u_dadda_cla32_fa743_xor1;
  assign f_u_dadda_cla32_fa876_or0 = f_u_dadda_cla32_fa876_and0 | f_u_dadda_cla32_fa876_and1;
  assign f_u_dadda_cla32_fa877_xor0 = f_u_dadda_cla32_fa876_or0 ^ f_u_dadda_cla32_fa744_xor1;
  assign f_u_dadda_cla32_fa877_and0 = f_u_dadda_cla32_fa876_or0 & f_u_dadda_cla32_fa744_xor1;
  assign f_u_dadda_cla32_fa877_xor1 = f_u_dadda_cla32_fa877_xor0 ^ f_u_dadda_cla32_fa745_xor1;
  assign f_u_dadda_cla32_fa877_and1 = f_u_dadda_cla32_fa877_xor0 & f_u_dadda_cla32_fa745_xor1;
  assign f_u_dadda_cla32_fa877_or0 = f_u_dadda_cla32_fa877_and0 | f_u_dadda_cla32_fa877_and1;
  assign f_u_dadda_cla32_fa878_xor0 = f_u_dadda_cla32_fa877_or0 ^ f_u_dadda_cla32_fa746_xor1;
  assign f_u_dadda_cla32_fa878_and0 = f_u_dadda_cla32_fa877_or0 & f_u_dadda_cla32_fa746_xor1;
  assign f_u_dadda_cla32_fa878_xor1 = f_u_dadda_cla32_fa878_xor0 ^ f_u_dadda_cla32_fa747_xor1;
  assign f_u_dadda_cla32_fa878_and1 = f_u_dadda_cla32_fa878_xor0 & f_u_dadda_cla32_fa747_xor1;
  assign f_u_dadda_cla32_fa878_or0 = f_u_dadda_cla32_fa878_and0 | f_u_dadda_cla32_fa878_and1;
  assign f_u_dadda_cla32_fa879_xor0 = f_u_dadda_cla32_fa878_or0 ^ f_u_dadda_cla32_fa748_xor1;
  assign f_u_dadda_cla32_fa879_and0 = f_u_dadda_cla32_fa878_or0 & f_u_dadda_cla32_fa748_xor1;
  assign f_u_dadda_cla32_fa879_xor1 = f_u_dadda_cla32_fa879_xor0 ^ f_u_dadda_cla32_fa749_xor1;
  assign f_u_dadda_cla32_fa879_and1 = f_u_dadda_cla32_fa879_xor0 & f_u_dadda_cla32_fa749_xor1;
  assign f_u_dadda_cla32_fa879_or0 = f_u_dadda_cla32_fa879_and0 | f_u_dadda_cla32_fa879_and1;
  assign f_u_dadda_cla32_fa880_xor0 = f_u_dadda_cla32_fa879_or0 ^ f_u_dadda_cla32_fa750_xor1;
  assign f_u_dadda_cla32_fa880_and0 = f_u_dadda_cla32_fa879_or0 & f_u_dadda_cla32_fa750_xor1;
  assign f_u_dadda_cla32_fa880_xor1 = f_u_dadda_cla32_fa880_xor0 ^ f_u_dadda_cla32_fa751_xor1;
  assign f_u_dadda_cla32_fa880_and1 = f_u_dadda_cla32_fa880_xor0 & f_u_dadda_cla32_fa751_xor1;
  assign f_u_dadda_cla32_fa880_or0 = f_u_dadda_cla32_fa880_and0 | f_u_dadda_cla32_fa880_and1;
  assign f_u_dadda_cla32_fa881_xor0 = f_u_dadda_cla32_fa880_or0 ^ f_u_dadda_cla32_fa752_xor1;
  assign f_u_dadda_cla32_fa881_and0 = f_u_dadda_cla32_fa880_or0 & f_u_dadda_cla32_fa752_xor1;
  assign f_u_dadda_cla32_fa881_xor1 = f_u_dadda_cla32_fa881_xor0 ^ f_u_dadda_cla32_fa753_xor1;
  assign f_u_dadda_cla32_fa881_and1 = f_u_dadda_cla32_fa881_xor0 & f_u_dadda_cla32_fa753_xor1;
  assign f_u_dadda_cla32_fa881_or0 = f_u_dadda_cla32_fa881_and0 | f_u_dadda_cla32_fa881_and1;
  assign f_u_dadda_cla32_fa882_xor0 = f_u_dadda_cla32_fa881_or0 ^ f_u_dadda_cla32_fa754_xor1;
  assign f_u_dadda_cla32_fa882_and0 = f_u_dadda_cla32_fa881_or0 & f_u_dadda_cla32_fa754_xor1;
  assign f_u_dadda_cla32_fa882_xor1 = f_u_dadda_cla32_fa882_xor0 ^ f_u_dadda_cla32_fa755_xor1;
  assign f_u_dadda_cla32_fa882_and1 = f_u_dadda_cla32_fa882_xor0 & f_u_dadda_cla32_fa755_xor1;
  assign f_u_dadda_cla32_fa882_or0 = f_u_dadda_cla32_fa882_and0 | f_u_dadda_cla32_fa882_and1;
  assign f_u_dadda_cla32_fa883_xor0 = f_u_dadda_cla32_fa882_or0 ^ f_u_dadda_cla32_fa756_xor1;
  assign f_u_dadda_cla32_fa883_and0 = f_u_dadda_cla32_fa882_or0 & f_u_dadda_cla32_fa756_xor1;
  assign f_u_dadda_cla32_fa883_xor1 = f_u_dadda_cla32_fa883_xor0 ^ f_u_dadda_cla32_fa757_xor1;
  assign f_u_dadda_cla32_fa883_and1 = f_u_dadda_cla32_fa883_xor0 & f_u_dadda_cla32_fa757_xor1;
  assign f_u_dadda_cla32_fa883_or0 = f_u_dadda_cla32_fa883_and0 | f_u_dadda_cla32_fa883_and1;
  assign f_u_dadda_cla32_fa884_xor0 = f_u_dadda_cla32_fa883_or0 ^ f_u_dadda_cla32_fa758_xor1;
  assign f_u_dadda_cla32_fa884_and0 = f_u_dadda_cla32_fa883_or0 & f_u_dadda_cla32_fa758_xor1;
  assign f_u_dadda_cla32_fa884_xor1 = f_u_dadda_cla32_fa884_xor0 ^ f_u_dadda_cla32_fa759_xor1;
  assign f_u_dadda_cla32_fa884_and1 = f_u_dadda_cla32_fa884_xor0 & f_u_dadda_cla32_fa759_xor1;
  assign f_u_dadda_cla32_fa884_or0 = f_u_dadda_cla32_fa884_and0 | f_u_dadda_cla32_fa884_and1;
  assign f_u_dadda_cla32_fa885_xor0 = f_u_dadda_cla32_fa884_or0 ^ f_u_dadda_cla32_fa760_xor1;
  assign f_u_dadda_cla32_fa885_and0 = f_u_dadda_cla32_fa884_or0 & f_u_dadda_cla32_fa760_xor1;
  assign f_u_dadda_cla32_fa885_xor1 = f_u_dadda_cla32_fa885_xor0 ^ f_u_dadda_cla32_fa761_xor1;
  assign f_u_dadda_cla32_fa885_and1 = f_u_dadda_cla32_fa885_xor0 & f_u_dadda_cla32_fa761_xor1;
  assign f_u_dadda_cla32_fa885_or0 = f_u_dadda_cla32_fa885_and0 | f_u_dadda_cla32_fa885_and1;
  assign f_u_dadda_cla32_fa886_xor0 = f_u_dadda_cla32_fa885_or0 ^ f_u_dadda_cla32_fa762_xor1;
  assign f_u_dadda_cla32_fa886_and0 = f_u_dadda_cla32_fa885_or0 & f_u_dadda_cla32_fa762_xor1;
  assign f_u_dadda_cla32_fa886_xor1 = f_u_dadda_cla32_fa886_xor0 ^ f_u_dadda_cla32_fa763_xor1;
  assign f_u_dadda_cla32_fa886_and1 = f_u_dadda_cla32_fa886_xor0 & f_u_dadda_cla32_fa763_xor1;
  assign f_u_dadda_cla32_fa886_or0 = f_u_dadda_cla32_fa886_and0 | f_u_dadda_cla32_fa886_and1;
  assign f_u_dadda_cla32_fa887_xor0 = f_u_dadda_cla32_fa886_or0 ^ f_u_dadda_cla32_fa764_xor1;
  assign f_u_dadda_cla32_fa887_and0 = f_u_dadda_cla32_fa886_or0 & f_u_dadda_cla32_fa764_xor1;
  assign f_u_dadda_cla32_fa887_xor1 = f_u_dadda_cla32_fa887_xor0 ^ f_u_dadda_cla32_fa765_xor1;
  assign f_u_dadda_cla32_fa887_and1 = f_u_dadda_cla32_fa887_xor0 & f_u_dadda_cla32_fa765_xor1;
  assign f_u_dadda_cla32_fa887_or0 = f_u_dadda_cla32_fa887_and0 | f_u_dadda_cla32_fa887_and1;
  assign f_u_dadda_cla32_fa888_xor0 = f_u_dadda_cla32_fa887_or0 ^ f_u_dadda_cla32_fa766_xor1;
  assign f_u_dadda_cla32_fa888_and0 = f_u_dadda_cla32_fa887_or0 & f_u_dadda_cla32_fa766_xor1;
  assign f_u_dadda_cla32_fa888_xor1 = f_u_dadda_cla32_fa888_xor0 ^ f_u_dadda_cla32_fa767_xor1;
  assign f_u_dadda_cla32_fa888_and1 = f_u_dadda_cla32_fa888_xor0 & f_u_dadda_cla32_fa767_xor1;
  assign f_u_dadda_cla32_fa888_or0 = f_u_dadda_cla32_fa888_and0 | f_u_dadda_cla32_fa888_and1;
  assign f_u_dadda_cla32_fa889_xor0 = f_u_dadda_cla32_fa888_or0 ^ f_u_dadda_cla32_fa768_xor1;
  assign f_u_dadda_cla32_fa889_and0 = f_u_dadda_cla32_fa888_or0 & f_u_dadda_cla32_fa768_xor1;
  assign f_u_dadda_cla32_fa889_xor1 = f_u_dadda_cla32_fa889_xor0 ^ f_u_dadda_cla32_fa769_xor1;
  assign f_u_dadda_cla32_fa889_and1 = f_u_dadda_cla32_fa889_xor0 & f_u_dadda_cla32_fa769_xor1;
  assign f_u_dadda_cla32_fa889_or0 = f_u_dadda_cla32_fa889_and0 | f_u_dadda_cla32_fa889_and1;
  assign f_u_dadda_cla32_fa890_xor0 = f_u_dadda_cla32_fa889_or0 ^ f_u_dadda_cla32_fa770_xor1;
  assign f_u_dadda_cla32_fa890_and0 = f_u_dadda_cla32_fa889_or0 & f_u_dadda_cla32_fa770_xor1;
  assign f_u_dadda_cla32_fa890_xor1 = f_u_dadda_cla32_fa890_xor0 ^ f_u_dadda_cla32_fa771_xor1;
  assign f_u_dadda_cla32_fa890_and1 = f_u_dadda_cla32_fa890_xor0 & f_u_dadda_cla32_fa771_xor1;
  assign f_u_dadda_cla32_fa890_or0 = f_u_dadda_cla32_fa890_and0 | f_u_dadda_cla32_fa890_and1;
  assign f_u_dadda_cla32_fa891_xor0 = f_u_dadda_cla32_fa890_or0 ^ f_u_dadda_cla32_fa772_xor1;
  assign f_u_dadda_cla32_fa891_and0 = f_u_dadda_cla32_fa890_or0 & f_u_dadda_cla32_fa772_xor1;
  assign f_u_dadda_cla32_fa891_xor1 = f_u_dadda_cla32_fa891_xor0 ^ f_u_dadda_cla32_fa773_xor1;
  assign f_u_dadda_cla32_fa891_and1 = f_u_dadda_cla32_fa891_xor0 & f_u_dadda_cla32_fa773_xor1;
  assign f_u_dadda_cla32_fa891_or0 = f_u_dadda_cla32_fa891_and0 | f_u_dadda_cla32_fa891_and1;
  assign f_u_dadda_cla32_fa892_xor0 = f_u_dadda_cla32_fa891_or0 ^ f_u_dadda_cla32_fa774_xor1;
  assign f_u_dadda_cla32_fa892_and0 = f_u_dadda_cla32_fa891_or0 & f_u_dadda_cla32_fa774_xor1;
  assign f_u_dadda_cla32_fa892_xor1 = f_u_dadda_cla32_fa892_xor0 ^ f_u_dadda_cla32_fa775_xor1;
  assign f_u_dadda_cla32_fa892_and1 = f_u_dadda_cla32_fa892_xor0 & f_u_dadda_cla32_fa775_xor1;
  assign f_u_dadda_cla32_fa892_or0 = f_u_dadda_cla32_fa892_and0 | f_u_dadda_cla32_fa892_and1;
  assign f_u_dadda_cla32_fa893_xor0 = f_u_dadda_cla32_fa892_or0 ^ f_u_dadda_cla32_fa776_xor1;
  assign f_u_dadda_cla32_fa893_and0 = f_u_dadda_cla32_fa892_or0 & f_u_dadda_cla32_fa776_xor1;
  assign f_u_dadda_cla32_fa893_xor1 = f_u_dadda_cla32_fa893_xor0 ^ f_u_dadda_cla32_fa777_xor1;
  assign f_u_dadda_cla32_fa893_and1 = f_u_dadda_cla32_fa893_xor0 & f_u_dadda_cla32_fa777_xor1;
  assign f_u_dadda_cla32_fa893_or0 = f_u_dadda_cla32_fa893_and0 | f_u_dadda_cla32_fa893_and1;
  assign f_u_dadda_cla32_fa894_xor0 = f_u_dadda_cla32_fa893_or0 ^ f_u_dadda_cla32_fa778_xor1;
  assign f_u_dadda_cla32_fa894_and0 = f_u_dadda_cla32_fa893_or0 & f_u_dadda_cla32_fa778_xor1;
  assign f_u_dadda_cla32_fa894_xor1 = f_u_dadda_cla32_fa894_xor0 ^ f_u_dadda_cla32_fa779_xor1;
  assign f_u_dadda_cla32_fa894_and1 = f_u_dadda_cla32_fa894_xor0 & f_u_dadda_cla32_fa779_xor1;
  assign f_u_dadda_cla32_fa894_or0 = f_u_dadda_cla32_fa894_and0 | f_u_dadda_cla32_fa894_and1;
  assign f_u_dadda_cla32_fa895_xor0 = f_u_dadda_cla32_fa894_or0 ^ f_u_dadda_cla32_fa780_xor1;
  assign f_u_dadda_cla32_fa895_and0 = f_u_dadda_cla32_fa894_or0 & f_u_dadda_cla32_fa780_xor1;
  assign f_u_dadda_cla32_fa895_xor1 = f_u_dadda_cla32_fa895_xor0 ^ f_u_dadda_cla32_fa781_xor1;
  assign f_u_dadda_cla32_fa895_and1 = f_u_dadda_cla32_fa895_xor0 & f_u_dadda_cla32_fa781_xor1;
  assign f_u_dadda_cla32_fa895_or0 = f_u_dadda_cla32_fa895_and0 | f_u_dadda_cla32_fa895_and1;
  assign f_u_dadda_cla32_and_28_31 = a[28] & b[31];
  assign f_u_dadda_cla32_fa896_xor0 = f_u_dadda_cla32_fa895_or0 ^ f_u_dadda_cla32_and_28_31;
  assign f_u_dadda_cla32_fa896_and0 = f_u_dadda_cla32_fa895_or0 & f_u_dadda_cla32_and_28_31;
  assign f_u_dadda_cla32_fa896_xor1 = f_u_dadda_cla32_fa896_xor0 ^ f_u_dadda_cla32_fa782_xor1;
  assign f_u_dadda_cla32_fa896_and1 = f_u_dadda_cla32_fa896_xor0 & f_u_dadda_cla32_fa782_xor1;
  assign f_u_dadda_cla32_fa896_or0 = f_u_dadda_cla32_fa896_and0 | f_u_dadda_cla32_fa896_and1;
  assign f_u_dadda_cla32_and_30_30 = a[30] & b[30];
  assign f_u_dadda_cla32_and_29_31 = a[29] & b[31];
  assign f_u_dadda_cla32_fa897_xor0 = f_u_dadda_cla32_fa896_or0 ^ f_u_dadda_cla32_and_30_30;
  assign f_u_dadda_cla32_fa897_and0 = f_u_dadda_cla32_fa896_or0 & f_u_dadda_cla32_and_30_30;
  assign f_u_dadda_cla32_fa897_xor1 = f_u_dadda_cla32_fa897_xor0 ^ f_u_dadda_cla32_and_29_31;
  assign f_u_dadda_cla32_fa897_and1 = f_u_dadda_cla32_fa897_xor0 & f_u_dadda_cla32_and_29_31;
  assign f_u_dadda_cla32_fa897_or0 = f_u_dadda_cla32_fa897_and0 | f_u_dadda_cla32_fa897_and1;
  assign f_u_dadda_cla32_and_31_30 = a[31] & b[30];
  assign f_u_dadda_cla32_fa898_xor0 = f_u_dadda_cla32_fa897_or0 ^ f_u_dadda_cla32_fa839_or0;
  assign f_u_dadda_cla32_fa898_and0 = f_u_dadda_cla32_fa897_or0 & f_u_dadda_cla32_fa839_or0;
  assign f_u_dadda_cla32_fa898_xor1 = f_u_dadda_cla32_fa898_xor0 ^ f_u_dadda_cla32_and_31_30;
  assign f_u_dadda_cla32_fa898_and1 = f_u_dadda_cla32_fa898_xor0 & f_u_dadda_cla32_and_31_30;
  assign f_u_dadda_cla32_fa898_or0 = f_u_dadda_cla32_fa898_and0 | f_u_dadda_cla32_fa898_and1;
  assign f_u_dadda_cla32_and_0_0 = a[0] & b[0];
  assign f_u_dadda_cla32_and_1_0 = a[1] & b[0];
  assign f_u_dadda_cla32_and_0_2 = a[0] & b[2];
  assign f_u_dadda_cla32_and_30_31 = a[30] & b[31];
  assign f_u_dadda_cla32_and_0_1 = a[0] & b[1];
  assign f_u_dadda_cla32_and_31_31 = a[31] & b[31];
  assign f_u_dadda_cla32_u_cla62_pg_logic0_or0 = f_u_dadda_cla32_and_1_0 | f_u_dadda_cla32_and_0_1;
  assign f_u_dadda_cla32_u_cla62_pg_logic0_and0 = f_u_dadda_cla32_and_1_0 & f_u_dadda_cla32_and_0_1;
  assign f_u_dadda_cla32_u_cla62_pg_logic0_xor0 = f_u_dadda_cla32_and_1_0 ^ f_u_dadda_cla32_and_0_1;
  assign f_u_dadda_cla32_u_cla62_pg_logic1_or0 = f_u_dadda_cla32_and_0_2 | f_u_dadda_cla32_ha30_xor0;
  assign f_u_dadda_cla32_u_cla62_pg_logic1_and0 = f_u_dadda_cla32_and_0_2 & f_u_dadda_cla32_ha30_xor0;
  assign f_u_dadda_cla32_u_cla62_pg_logic1_xor0 = f_u_dadda_cla32_and_0_2 ^ f_u_dadda_cla32_ha30_xor0;
  assign f_u_dadda_cla32_u_cla62_xor1 = f_u_dadda_cla32_u_cla62_pg_logic1_xor0 ^ f_u_dadda_cla32_u_cla62_pg_logic0_and0;
  assign f_u_dadda_cla32_u_cla62_and0 = f_u_dadda_cla32_u_cla62_pg_logic0_and0 & f_u_dadda_cla32_u_cla62_pg_logic1_or0;
  assign f_u_dadda_cla32_u_cla62_or0 = f_u_dadda_cla32_u_cla62_pg_logic1_and0 | f_u_dadda_cla32_u_cla62_and0;
  assign f_u_dadda_cla32_u_cla62_pg_logic2_or0 = f_u_dadda_cla32_ha29_xor0 | f_u_dadda_cla32_fa840_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic2_and0 = f_u_dadda_cla32_ha29_xor0 & f_u_dadda_cla32_fa840_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic2_xor0 = f_u_dadda_cla32_ha29_xor0 ^ f_u_dadda_cla32_fa840_xor1;
  assign f_u_dadda_cla32_u_cla62_xor2 = f_u_dadda_cla32_u_cla62_pg_logic2_xor0 ^ f_u_dadda_cla32_u_cla62_or0;
  assign f_u_dadda_cla32_u_cla62_and1 = f_u_dadda_cla32_u_cla62_pg_logic2_or0 & f_u_dadda_cla32_u_cla62_pg_logic0_or0;
  assign f_u_dadda_cla32_u_cla62_and2 = f_u_dadda_cla32_u_cla62_pg_logic0_and0 & f_u_dadda_cla32_u_cla62_pg_logic2_or0;
  assign f_u_dadda_cla32_u_cla62_and3 = f_u_dadda_cla32_u_cla62_and2 & f_u_dadda_cla32_u_cla62_pg_logic1_or0;
  assign f_u_dadda_cla32_u_cla62_and4 = f_u_dadda_cla32_u_cla62_pg_logic1_and0 & f_u_dadda_cla32_u_cla62_pg_logic2_or0;
  assign f_u_dadda_cla32_u_cla62_or1 = f_u_dadda_cla32_u_cla62_and3 | f_u_dadda_cla32_u_cla62_and4;
  assign f_u_dadda_cla32_u_cla62_or2 = f_u_dadda_cla32_u_cla62_pg_logic2_and0 | f_u_dadda_cla32_u_cla62_or1;
  assign f_u_dadda_cla32_u_cla62_pg_logic3_or0 = f_u_dadda_cla32_fa783_xor1 | f_u_dadda_cla32_fa841_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic3_and0 = f_u_dadda_cla32_fa783_xor1 & f_u_dadda_cla32_fa841_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic3_xor0 = f_u_dadda_cla32_fa783_xor1 ^ f_u_dadda_cla32_fa841_xor1;
  assign f_u_dadda_cla32_u_cla62_xor3 = f_u_dadda_cla32_u_cla62_pg_logic3_xor0 ^ f_u_dadda_cla32_u_cla62_or2;
  assign f_u_dadda_cla32_u_cla62_and5 = f_u_dadda_cla32_u_cla62_pg_logic3_or0 & f_u_dadda_cla32_u_cla62_pg_logic1_or0;
  assign f_u_dadda_cla32_u_cla62_and6 = f_u_dadda_cla32_u_cla62_pg_logic0_and0 & f_u_dadda_cla32_u_cla62_pg_logic2_or0;
  assign f_u_dadda_cla32_u_cla62_and7 = f_u_dadda_cla32_u_cla62_pg_logic3_or0 & f_u_dadda_cla32_u_cla62_pg_logic1_or0;
  assign f_u_dadda_cla32_u_cla62_and8 = f_u_dadda_cla32_u_cla62_and6 & f_u_dadda_cla32_u_cla62_and7;
  assign f_u_dadda_cla32_u_cla62_and9 = f_u_dadda_cla32_u_cla62_pg_logic1_and0 & f_u_dadda_cla32_u_cla62_pg_logic3_or0;
  assign f_u_dadda_cla32_u_cla62_and10 = f_u_dadda_cla32_u_cla62_and9 & f_u_dadda_cla32_u_cla62_pg_logic2_or0;
  assign f_u_dadda_cla32_u_cla62_and11 = f_u_dadda_cla32_u_cla62_pg_logic2_and0 & f_u_dadda_cla32_u_cla62_pg_logic3_or0;
  assign f_u_dadda_cla32_u_cla62_or3 = f_u_dadda_cla32_u_cla62_and8 | f_u_dadda_cla32_u_cla62_and11;
  assign f_u_dadda_cla32_u_cla62_or4 = f_u_dadda_cla32_u_cla62_and10 | f_u_dadda_cla32_u_cla62_or3;
  assign f_u_dadda_cla32_u_cla62_or5 = f_u_dadda_cla32_u_cla62_pg_logic3_and0 | f_u_dadda_cla32_u_cla62_or4;
  assign f_u_dadda_cla32_u_cla62_pg_logic4_or0 = f_u_dadda_cla32_fa784_xor1 | f_u_dadda_cla32_fa842_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic4_and0 = f_u_dadda_cla32_fa784_xor1 & f_u_dadda_cla32_fa842_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic4_xor0 = f_u_dadda_cla32_fa784_xor1 ^ f_u_dadda_cla32_fa842_xor1;
  assign f_u_dadda_cla32_u_cla62_xor4 = f_u_dadda_cla32_u_cla62_pg_logic4_xor0 ^ f_u_dadda_cla32_u_cla62_or5;
  assign f_u_dadda_cla32_u_cla62_and12 = f_u_dadda_cla32_u_cla62_or5 & f_u_dadda_cla32_u_cla62_pg_logic4_or0;
  assign f_u_dadda_cla32_u_cla62_or6 = f_u_dadda_cla32_u_cla62_pg_logic4_and0 | f_u_dadda_cla32_u_cla62_and12;
  assign f_u_dadda_cla32_u_cla62_pg_logic5_or0 = f_u_dadda_cla32_fa785_xor1 | f_u_dadda_cla32_fa843_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic5_and0 = f_u_dadda_cla32_fa785_xor1 & f_u_dadda_cla32_fa843_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic5_xor0 = f_u_dadda_cla32_fa785_xor1 ^ f_u_dadda_cla32_fa843_xor1;
  assign f_u_dadda_cla32_u_cla62_xor5 = f_u_dadda_cla32_u_cla62_pg_logic5_xor0 ^ f_u_dadda_cla32_u_cla62_or6;
  assign f_u_dadda_cla32_u_cla62_and13 = f_u_dadda_cla32_u_cla62_or5 & f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  assign f_u_dadda_cla32_u_cla62_and14 = f_u_dadda_cla32_u_cla62_and13 & f_u_dadda_cla32_u_cla62_pg_logic4_or0;
  assign f_u_dadda_cla32_u_cla62_and15 = f_u_dadda_cla32_u_cla62_pg_logic4_and0 & f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  assign f_u_dadda_cla32_u_cla62_or7 = f_u_dadda_cla32_u_cla62_and14 | f_u_dadda_cla32_u_cla62_and15;
  assign f_u_dadda_cla32_u_cla62_or8 = f_u_dadda_cla32_u_cla62_pg_logic5_and0 | f_u_dadda_cla32_u_cla62_or7;
  assign f_u_dadda_cla32_u_cla62_pg_logic6_or0 = f_u_dadda_cla32_fa786_xor1 | f_u_dadda_cla32_fa844_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic6_and0 = f_u_dadda_cla32_fa786_xor1 & f_u_dadda_cla32_fa844_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic6_xor0 = f_u_dadda_cla32_fa786_xor1 ^ f_u_dadda_cla32_fa844_xor1;
  assign f_u_dadda_cla32_u_cla62_xor6 = f_u_dadda_cla32_u_cla62_pg_logic6_xor0 ^ f_u_dadda_cla32_u_cla62_or8;
  assign f_u_dadda_cla32_u_cla62_and16 = f_u_dadda_cla32_u_cla62_or5 & f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  assign f_u_dadda_cla32_u_cla62_and17 = f_u_dadda_cla32_u_cla62_pg_logic6_or0 & f_u_dadda_cla32_u_cla62_pg_logic4_or0;
  assign f_u_dadda_cla32_u_cla62_and18 = f_u_dadda_cla32_u_cla62_and16 & f_u_dadda_cla32_u_cla62_and17;
  assign f_u_dadda_cla32_u_cla62_and19 = f_u_dadda_cla32_u_cla62_pg_logic4_and0 & f_u_dadda_cla32_u_cla62_pg_logic6_or0;
  assign f_u_dadda_cla32_u_cla62_and20 = f_u_dadda_cla32_u_cla62_and19 & f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  assign f_u_dadda_cla32_u_cla62_and21 = f_u_dadda_cla32_u_cla62_pg_logic5_and0 & f_u_dadda_cla32_u_cla62_pg_logic6_or0;
  assign f_u_dadda_cla32_u_cla62_or9 = f_u_dadda_cla32_u_cla62_and18 | f_u_dadda_cla32_u_cla62_and20;
  assign f_u_dadda_cla32_u_cla62_or10 = f_u_dadda_cla32_u_cla62_or9 | f_u_dadda_cla32_u_cla62_and21;
  assign f_u_dadda_cla32_u_cla62_or11 = f_u_dadda_cla32_u_cla62_pg_logic6_and0 | f_u_dadda_cla32_u_cla62_or10;
  assign f_u_dadda_cla32_u_cla62_pg_logic7_or0 = f_u_dadda_cla32_fa787_xor1 | f_u_dadda_cla32_fa845_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic7_and0 = f_u_dadda_cla32_fa787_xor1 & f_u_dadda_cla32_fa845_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic7_xor0 = f_u_dadda_cla32_fa787_xor1 ^ f_u_dadda_cla32_fa845_xor1;
  assign f_u_dadda_cla32_u_cla62_xor7 = f_u_dadda_cla32_u_cla62_pg_logic7_xor0 ^ f_u_dadda_cla32_u_cla62_or11;
  assign f_u_dadda_cla32_u_cla62_and22 = f_u_dadda_cla32_u_cla62_or5 & f_u_dadda_cla32_u_cla62_pg_logic6_or0;
  assign f_u_dadda_cla32_u_cla62_and23 = f_u_dadda_cla32_u_cla62_pg_logic7_or0 & f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  assign f_u_dadda_cla32_u_cla62_and24 = f_u_dadda_cla32_u_cla62_and22 & f_u_dadda_cla32_u_cla62_and23;
  assign f_u_dadda_cla32_u_cla62_and25 = f_u_dadda_cla32_u_cla62_and24 & f_u_dadda_cla32_u_cla62_pg_logic4_or0;
  assign f_u_dadda_cla32_u_cla62_and26 = f_u_dadda_cla32_u_cla62_pg_logic4_and0 & f_u_dadda_cla32_u_cla62_pg_logic6_or0;
  assign f_u_dadda_cla32_u_cla62_and27 = f_u_dadda_cla32_u_cla62_pg_logic7_or0 & f_u_dadda_cla32_u_cla62_pg_logic5_or0;
  assign f_u_dadda_cla32_u_cla62_and28 = f_u_dadda_cla32_u_cla62_and26 & f_u_dadda_cla32_u_cla62_and27;
  assign f_u_dadda_cla32_u_cla62_and29 = f_u_dadda_cla32_u_cla62_pg_logic5_and0 & f_u_dadda_cla32_u_cla62_pg_logic7_or0;
  assign f_u_dadda_cla32_u_cla62_and30 = f_u_dadda_cla32_u_cla62_and29 & f_u_dadda_cla32_u_cla62_pg_logic6_or0;
  assign f_u_dadda_cla32_u_cla62_and31 = f_u_dadda_cla32_u_cla62_pg_logic6_and0 & f_u_dadda_cla32_u_cla62_pg_logic7_or0;
  assign f_u_dadda_cla32_u_cla62_or12 = f_u_dadda_cla32_u_cla62_and25 | f_u_dadda_cla32_u_cla62_and30;
  assign f_u_dadda_cla32_u_cla62_or13 = f_u_dadda_cla32_u_cla62_and28 | f_u_dadda_cla32_u_cla62_and31;
  assign f_u_dadda_cla32_u_cla62_or14 = f_u_dadda_cla32_u_cla62_or12 | f_u_dadda_cla32_u_cla62_or13;
  assign f_u_dadda_cla32_u_cla62_or15 = f_u_dadda_cla32_u_cla62_pg_logic7_and0 | f_u_dadda_cla32_u_cla62_or14;
  assign f_u_dadda_cla32_u_cla62_pg_logic8_or0 = f_u_dadda_cla32_fa788_xor1 | f_u_dadda_cla32_fa846_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic8_and0 = f_u_dadda_cla32_fa788_xor1 & f_u_dadda_cla32_fa846_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic8_xor0 = f_u_dadda_cla32_fa788_xor1 ^ f_u_dadda_cla32_fa846_xor1;
  assign f_u_dadda_cla32_u_cla62_xor8 = f_u_dadda_cla32_u_cla62_pg_logic8_xor0 ^ f_u_dadda_cla32_u_cla62_or15;
  assign f_u_dadda_cla32_u_cla62_and32 = f_u_dadda_cla32_u_cla62_or15 & f_u_dadda_cla32_u_cla62_pg_logic8_or0;
  assign f_u_dadda_cla32_u_cla62_or16 = f_u_dadda_cla32_u_cla62_pg_logic8_and0 | f_u_dadda_cla32_u_cla62_and32;
  assign f_u_dadda_cla32_u_cla62_pg_logic9_or0 = f_u_dadda_cla32_fa789_xor1 | f_u_dadda_cla32_fa847_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic9_and0 = f_u_dadda_cla32_fa789_xor1 & f_u_dadda_cla32_fa847_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic9_xor0 = f_u_dadda_cla32_fa789_xor1 ^ f_u_dadda_cla32_fa847_xor1;
  assign f_u_dadda_cla32_u_cla62_xor9 = f_u_dadda_cla32_u_cla62_pg_logic9_xor0 ^ f_u_dadda_cla32_u_cla62_or16;
  assign f_u_dadda_cla32_u_cla62_and33 = f_u_dadda_cla32_u_cla62_or15 & f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  assign f_u_dadda_cla32_u_cla62_and34 = f_u_dadda_cla32_u_cla62_and33 & f_u_dadda_cla32_u_cla62_pg_logic8_or0;
  assign f_u_dadda_cla32_u_cla62_and35 = f_u_dadda_cla32_u_cla62_pg_logic8_and0 & f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  assign f_u_dadda_cla32_u_cla62_or17 = f_u_dadda_cla32_u_cla62_and34 | f_u_dadda_cla32_u_cla62_and35;
  assign f_u_dadda_cla32_u_cla62_or18 = f_u_dadda_cla32_u_cla62_pg_logic9_and0 | f_u_dadda_cla32_u_cla62_or17;
  assign f_u_dadda_cla32_u_cla62_pg_logic10_or0 = f_u_dadda_cla32_fa790_xor1 | f_u_dadda_cla32_fa848_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic10_and0 = f_u_dadda_cla32_fa790_xor1 & f_u_dadda_cla32_fa848_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic10_xor0 = f_u_dadda_cla32_fa790_xor1 ^ f_u_dadda_cla32_fa848_xor1;
  assign f_u_dadda_cla32_u_cla62_xor10 = f_u_dadda_cla32_u_cla62_pg_logic10_xor0 ^ f_u_dadda_cla32_u_cla62_or18;
  assign f_u_dadda_cla32_u_cla62_and36 = f_u_dadda_cla32_u_cla62_or15 & f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  assign f_u_dadda_cla32_u_cla62_and37 = f_u_dadda_cla32_u_cla62_pg_logic10_or0 & f_u_dadda_cla32_u_cla62_pg_logic8_or0;
  assign f_u_dadda_cla32_u_cla62_and38 = f_u_dadda_cla32_u_cla62_and36 & f_u_dadda_cla32_u_cla62_and37;
  assign f_u_dadda_cla32_u_cla62_and39 = f_u_dadda_cla32_u_cla62_pg_logic8_and0 & f_u_dadda_cla32_u_cla62_pg_logic10_or0;
  assign f_u_dadda_cla32_u_cla62_and40 = f_u_dadda_cla32_u_cla62_and39 & f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  assign f_u_dadda_cla32_u_cla62_and41 = f_u_dadda_cla32_u_cla62_pg_logic9_and0 & f_u_dadda_cla32_u_cla62_pg_logic10_or0;
  assign f_u_dadda_cla32_u_cla62_or19 = f_u_dadda_cla32_u_cla62_and38 | f_u_dadda_cla32_u_cla62_and40;
  assign f_u_dadda_cla32_u_cla62_or20 = f_u_dadda_cla32_u_cla62_or19 | f_u_dadda_cla32_u_cla62_and41;
  assign f_u_dadda_cla32_u_cla62_or21 = f_u_dadda_cla32_u_cla62_pg_logic10_and0 | f_u_dadda_cla32_u_cla62_or20;
  assign f_u_dadda_cla32_u_cla62_pg_logic11_or0 = f_u_dadda_cla32_fa791_xor1 | f_u_dadda_cla32_fa849_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic11_and0 = f_u_dadda_cla32_fa791_xor1 & f_u_dadda_cla32_fa849_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic11_xor0 = f_u_dadda_cla32_fa791_xor1 ^ f_u_dadda_cla32_fa849_xor1;
  assign f_u_dadda_cla32_u_cla62_xor11 = f_u_dadda_cla32_u_cla62_pg_logic11_xor0 ^ f_u_dadda_cla32_u_cla62_or21;
  assign f_u_dadda_cla32_u_cla62_and42 = f_u_dadda_cla32_u_cla62_or15 & f_u_dadda_cla32_u_cla62_pg_logic10_or0;
  assign f_u_dadda_cla32_u_cla62_and43 = f_u_dadda_cla32_u_cla62_pg_logic11_or0 & f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  assign f_u_dadda_cla32_u_cla62_and44 = f_u_dadda_cla32_u_cla62_and42 & f_u_dadda_cla32_u_cla62_and43;
  assign f_u_dadda_cla32_u_cla62_and45 = f_u_dadda_cla32_u_cla62_and44 & f_u_dadda_cla32_u_cla62_pg_logic8_or0;
  assign f_u_dadda_cla32_u_cla62_and46 = f_u_dadda_cla32_u_cla62_pg_logic8_and0 & f_u_dadda_cla32_u_cla62_pg_logic10_or0;
  assign f_u_dadda_cla32_u_cla62_and47 = f_u_dadda_cla32_u_cla62_pg_logic11_or0 & f_u_dadda_cla32_u_cla62_pg_logic9_or0;
  assign f_u_dadda_cla32_u_cla62_and48 = f_u_dadda_cla32_u_cla62_and46 & f_u_dadda_cla32_u_cla62_and47;
  assign f_u_dadda_cla32_u_cla62_and49 = f_u_dadda_cla32_u_cla62_pg_logic9_and0 & f_u_dadda_cla32_u_cla62_pg_logic11_or0;
  assign f_u_dadda_cla32_u_cla62_and50 = f_u_dadda_cla32_u_cla62_and49 & f_u_dadda_cla32_u_cla62_pg_logic10_or0;
  assign f_u_dadda_cla32_u_cla62_and51 = f_u_dadda_cla32_u_cla62_pg_logic10_and0 & f_u_dadda_cla32_u_cla62_pg_logic11_or0;
  assign f_u_dadda_cla32_u_cla62_or22 = f_u_dadda_cla32_u_cla62_and45 | f_u_dadda_cla32_u_cla62_and50;
  assign f_u_dadda_cla32_u_cla62_or23 = f_u_dadda_cla32_u_cla62_and48 | f_u_dadda_cla32_u_cla62_and51;
  assign f_u_dadda_cla32_u_cla62_or24 = f_u_dadda_cla32_u_cla62_or22 | f_u_dadda_cla32_u_cla62_or23;
  assign f_u_dadda_cla32_u_cla62_or25 = f_u_dadda_cla32_u_cla62_pg_logic11_and0 | f_u_dadda_cla32_u_cla62_or24;
  assign f_u_dadda_cla32_u_cla62_pg_logic12_or0 = f_u_dadda_cla32_fa792_xor1 | f_u_dadda_cla32_fa850_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic12_and0 = f_u_dadda_cla32_fa792_xor1 & f_u_dadda_cla32_fa850_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic12_xor0 = f_u_dadda_cla32_fa792_xor1 ^ f_u_dadda_cla32_fa850_xor1;
  assign f_u_dadda_cla32_u_cla62_xor12 = f_u_dadda_cla32_u_cla62_pg_logic12_xor0 ^ f_u_dadda_cla32_u_cla62_or25;
  assign f_u_dadda_cla32_u_cla62_and52 = f_u_dadda_cla32_u_cla62_or25 & f_u_dadda_cla32_u_cla62_pg_logic12_or0;
  assign f_u_dadda_cla32_u_cla62_or26 = f_u_dadda_cla32_u_cla62_pg_logic12_and0 | f_u_dadda_cla32_u_cla62_and52;
  assign f_u_dadda_cla32_u_cla62_pg_logic13_or0 = f_u_dadda_cla32_fa793_xor1 | f_u_dadda_cla32_fa851_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic13_and0 = f_u_dadda_cla32_fa793_xor1 & f_u_dadda_cla32_fa851_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic13_xor0 = f_u_dadda_cla32_fa793_xor1 ^ f_u_dadda_cla32_fa851_xor1;
  assign f_u_dadda_cla32_u_cla62_xor13 = f_u_dadda_cla32_u_cla62_pg_logic13_xor0 ^ f_u_dadda_cla32_u_cla62_or26;
  assign f_u_dadda_cla32_u_cla62_and53 = f_u_dadda_cla32_u_cla62_or25 & f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  assign f_u_dadda_cla32_u_cla62_and54 = f_u_dadda_cla32_u_cla62_and53 & f_u_dadda_cla32_u_cla62_pg_logic12_or0;
  assign f_u_dadda_cla32_u_cla62_and55 = f_u_dadda_cla32_u_cla62_pg_logic12_and0 & f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  assign f_u_dadda_cla32_u_cla62_or27 = f_u_dadda_cla32_u_cla62_and54 | f_u_dadda_cla32_u_cla62_and55;
  assign f_u_dadda_cla32_u_cla62_or28 = f_u_dadda_cla32_u_cla62_pg_logic13_and0 | f_u_dadda_cla32_u_cla62_or27;
  assign f_u_dadda_cla32_u_cla62_pg_logic14_or0 = f_u_dadda_cla32_fa794_xor1 | f_u_dadda_cla32_fa852_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic14_and0 = f_u_dadda_cla32_fa794_xor1 & f_u_dadda_cla32_fa852_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic14_xor0 = f_u_dadda_cla32_fa794_xor1 ^ f_u_dadda_cla32_fa852_xor1;
  assign f_u_dadda_cla32_u_cla62_xor14 = f_u_dadda_cla32_u_cla62_pg_logic14_xor0 ^ f_u_dadda_cla32_u_cla62_or28;
  assign f_u_dadda_cla32_u_cla62_and56 = f_u_dadda_cla32_u_cla62_or25 & f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  assign f_u_dadda_cla32_u_cla62_and57 = f_u_dadda_cla32_u_cla62_pg_logic14_or0 & f_u_dadda_cla32_u_cla62_pg_logic12_or0;
  assign f_u_dadda_cla32_u_cla62_and58 = f_u_dadda_cla32_u_cla62_and56 & f_u_dadda_cla32_u_cla62_and57;
  assign f_u_dadda_cla32_u_cla62_and59 = f_u_dadda_cla32_u_cla62_pg_logic12_and0 & f_u_dadda_cla32_u_cla62_pg_logic14_or0;
  assign f_u_dadda_cla32_u_cla62_and60 = f_u_dadda_cla32_u_cla62_and59 & f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  assign f_u_dadda_cla32_u_cla62_and61 = f_u_dadda_cla32_u_cla62_pg_logic13_and0 & f_u_dadda_cla32_u_cla62_pg_logic14_or0;
  assign f_u_dadda_cla32_u_cla62_or29 = f_u_dadda_cla32_u_cla62_and58 | f_u_dadda_cla32_u_cla62_and60;
  assign f_u_dadda_cla32_u_cla62_or30 = f_u_dadda_cla32_u_cla62_or29 | f_u_dadda_cla32_u_cla62_and61;
  assign f_u_dadda_cla32_u_cla62_or31 = f_u_dadda_cla32_u_cla62_pg_logic14_and0 | f_u_dadda_cla32_u_cla62_or30;
  assign f_u_dadda_cla32_u_cla62_pg_logic15_or0 = f_u_dadda_cla32_fa795_xor1 | f_u_dadda_cla32_fa853_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic15_and0 = f_u_dadda_cla32_fa795_xor1 & f_u_dadda_cla32_fa853_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic15_xor0 = f_u_dadda_cla32_fa795_xor1 ^ f_u_dadda_cla32_fa853_xor1;
  assign f_u_dadda_cla32_u_cla62_xor15 = f_u_dadda_cla32_u_cla62_pg_logic15_xor0 ^ f_u_dadda_cla32_u_cla62_or31;
  assign f_u_dadda_cla32_u_cla62_and62 = f_u_dadda_cla32_u_cla62_or25 & f_u_dadda_cla32_u_cla62_pg_logic14_or0;
  assign f_u_dadda_cla32_u_cla62_and63 = f_u_dadda_cla32_u_cla62_pg_logic15_or0 & f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  assign f_u_dadda_cla32_u_cla62_and64 = f_u_dadda_cla32_u_cla62_and62 & f_u_dadda_cla32_u_cla62_and63;
  assign f_u_dadda_cla32_u_cla62_and65 = f_u_dadda_cla32_u_cla62_and64 & f_u_dadda_cla32_u_cla62_pg_logic12_or0;
  assign f_u_dadda_cla32_u_cla62_and66 = f_u_dadda_cla32_u_cla62_pg_logic12_and0 & f_u_dadda_cla32_u_cla62_pg_logic14_or0;
  assign f_u_dadda_cla32_u_cla62_and67 = f_u_dadda_cla32_u_cla62_pg_logic15_or0 & f_u_dadda_cla32_u_cla62_pg_logic13_or0;
  assign f_u_dadda_cla32_u_cla62_and68 = f_u_dadda_cla32_u_cla62_and66 & f_u_dadda_cla32_u_cla62_and67;
  assign f_u_dadda_cla32_u_cla62_and69 = f_u_dadda_cla32_u_cla62_pg_logic13_and0 & f_u_dadda_cla32_u_cla62_pg_logic15_or0;
  assign f_u_dadda_cla32_u_cla62_and70 = f_u_dadda_cla32_u_cla62_and69 & f_u_dadda_cla32_u_cla62_pg_logic14_or0;
  assign f_u_dadda_cla32_u_cla62_and71 = f_u_dadda_cla32_u_cla62_pg_logic14_and0 & f_u_dadda_cla32_u_cla62_pg_logic15_or0;
  assign f_u_dadda_cla32_u_cla62_or32 = f_u_dadda_cla32_u_cla62_and65 | f_u_dadda_cla32_u_cla62_and70;
  assign f_u_dadda_cla32_u_cla62_or33 = f_u_dadda_cla32_u_cla62_and68 | f_u_dadda_cla32_u_cla62_and71;
  assign f_u_dadda_cla32_u_cla62_or34 = f_u_dadda_cla32_u_cla62_or32 | f_u_dadda_cla32_u_cla62_or33;
  assign f_u_dadda_cla32_u_cla62_or35 = f_u_dadda_cla32_u_cla62_pg_logic15_and0 | f_u_dadda_cla32_u_cla62_or34;
  assign f_u_dadda_cla32_u_cla62_pg_logic16_or0 = f_u_dadda_cla32_fa796_xor1 | f_u_dadda_cla32_fa854_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic16_and0 = f_u_dadda_cla32_fa796_xor1 & f_u_dadda_cla32_fa854_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic16_xor0 = f_u_dadda_cla32_fa796_xor1 ^ f_u_dadda_cla32_fa854_xor1;
  assign f_u_dadda_cla32_u_cla62_xor16 = f_u_dadda_cla32_u_cla62_pg_logic16_xor0 ^ f_u_dadda_cla32_u_cla62_or35;
  assign f_u_dadda_cla32_u_cla62_and72 = f_u_dadda_cla32_u_cla62_or35 & f_u_dadda_cla32_u_cla62_pg_logic16_or0;
  assign f_u_dadda_cla32_u_cla62_or36 = f_u_dadda_cla32_u_cla62_pg_logic16_and0 | f_u_dadda_cla32_u_cla62_and72;
  assign f_u_dadda_cla32_u_cla62_pg_logic17_or0 = f_u_dadda_cla32_fa797_xor1 | f_u_dadda_cla32_fa855_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic17_and0 = f_u_dadda_cla32_fa797_xor1 & f_u_dadda_cla32_fa855_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic17_xor0 = f_u_dadda_cla32_fa797_xor1 ^ f_u_dadda_cla32_fa855_xor1;
  assign f_u_dadda_cla32_u_cla62_xor17 = f_u_dadda_cla32_u_cla62_pg_logic17_xor0 ^ f_u_dadda_cla32_u_cla62_or36;
  assign f_u_dadda_cla32_u_cla62_and73 = f_u_dadda_cla32_u_cla62_or35 & f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  assign f_u_dadda_cla32_u_cla62_and74 = f_u_dadda_cla32_u_cla62_and73 & f_u_dadda_cla32_u_cla62_pg_logic16_or0;
  assign f_u_dadda_cla32_u_cla62_and75 = f_u_dadda_cla32_u_cla62_pg_logic16_and0 & f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  assign f_u_dadda_cla32_u_cla62_or37 = f_u_dadda_cla32_u_cla62_and74 | f_u_dadda_cla32_u_cla62_and75;
  assign f_u_dadda_cla32_u_cla62_or38 = f_u_dadda_cla32_u_cla62_pg_logic17_and0 | f_u_dadda_cla32_u_cla62_or37;
  assign f_u_dadda_cla32_u_cla62_pg_logic18_or0 = f_u_dadda_cla32_fa798_xor1 | f_u_dadda_cla32_fa856_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic18_and0 = f_u_dadda_cla32_fa798_xor1 & f_u_dadda_cla32_fa856_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic18_xor0 = f_u_dadda_cla32_fa798_xor1 ^ f_u_dadda_cla32_fa856_xor1;
  assign f_u_dadda_cla32_u_cla62_xor18 = f_u_dadda_cla32_u_cla62_pg_logic18_xor0 ^ f_u_dadda_cla32_u_cla62_or38;
  assign f_u_dadda_cla32_u_cla62_and76 = f_u_dadda_cla32_u_cla62_or35 & f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  assign f_u_dadda_cla32_u_cla62_and77 = f_u_dadda_cla32_u_cla62_pg_logic18_or0 & f_u_dadda_cla32_u_cla62_pg_logic16_or0;
  assign f_u_dadda_cla32_u_cla62_and78 = f_u_dadda_cla32_u_cla62_and76 & f_u_dadda_cla32_u_cla62_and77;
  assign f_u_dadda_cla32_u_cla62_and79 = f_u_dadda_cla32_u_cla62_pg_logic16_and0 & f_u_dadda_cla32_u_cla62_pg_logic18_or0;
  assign f_u_dadda_cla32_u_cla62_and80 = f_u_dadda_cla32_u_cla62_and79 & f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  assign f_u_dadda_cla32_u_cla62_and81 = f_u_dadda_cla32_u_cla62_pg_logic17_and0 & f_u_dadda_cla32_u_cla62_pg_logic18_or0;
  assign f_u_dadda_cla32_u_cla62_or39 = f_u_dadda_cla32_u_cla62_and78 | f_u_dadda_cla32_u_cla62_and80;
  assign f_u_dadda_cla32_u_cla62_or40 = f_u_dadda_cla32_u_cla62_or39 | f_u_dadda_cla32_u_cla62_and81;
  assign f_u_dadda_cla32_u_cla62_or41 = f_u_dadda_cla32_u_cla62_pg_logic18_and0 | f_u_dadda_cla32_u_cla62_or40;
  assign f_u_dadda_cla32_u_cla62_pg_logic19_or0 = f_u_dadda_cla32_fa799_xor1 | f_u_dadda_cla32_fa857_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic19_and0 = f_u_dadda_cla32_fa799_xor1 & f_u_dadda_cla32_fa857_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic19_xor0 = f_u_dadda_cla32_fa799_xor1 ^ f_u_dadda_cla32_fa857_xor1;
  assign f_u_dadda_cla32_u_cla62_xor19 = f_u_dadda_cla32_u_cla62_pg_logic19_xor0 ^ f_u_dadda_cla32_u_cla62_or41;
  assign f_u_dadda_cla32_u_cla62_and82 = f_u_dadda_cla32_u_cla62_or35 & f_u_dadda_cla32_u_cla62_pg_logic18_or0;
  assign f_u_dadda_cla32_u_cla62_and83 = f_u_dadda_cla32_u_cla62_pg_logic19_or0 & f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  assign f_u_dadda_cla32_u_cla62_and84 = f_u_dadda_cla32_u_cla62_and82 & f_u_dadda_cla32_u_cla62_and83;
  assign f_u_dadda_cla32_u_cla62_and85 = f_u_dadda_cla32_u_cla62_and84 & f_u_dadda_cla32_u_cla62_pg_logic16_or0;
  assign f_u_dadda_cla32_u_cla62_and86 = f_u_dadda_cla32_u_cla62_pg_logic16_and0 & f_u_dadda_cla32_u_cla62_pg_logic18_or0;
  assign f_u_dadda_cla32_u_cla62_and87 = f_u_dadda_cla32_u_cla62_pg_logic19_or0 & f_u_dadda_cla32_u_cla62_pg_logic17_or0;
  assign f_u_dadda_cla32_u_cla62_and88 = f_u_dadda_cla32_u_cla62_and86 & f_u_dadda_cla32_u_cla62_and87;
  assign f_u_dadda_cla32_u_cla62_and89 = f_u_dadda_cla32_u_cla62_pg_logic17_and0 & f_u_dadda_cla32_u_cla62_pg_logic19_or0;
  assign f_u_dadda_cla32_u_cla62_and90 = f_u_dadda_cla32_u_cla62_and89 & f_u_dadda_cla32_u_cla62_pg_logic18_or0;
  assign f_u_dadda_cla32_u_cla62_and91 = f_u_dadda_cla32_u_cla62_pg_logic18_and0 & f_u_dadda_cla32_u_cla62_pg_logic19_or0;
  assign f_u_dadda_cla32_u_cla62_or42 = f_u_dadda_cla32_u_cla62_and85 | f_u_dadda_cla32_u_cla62_and90;
  assign f_u_dadda_cla32_u_cla62_or43 = f_u_dadda_cla32_u_cla62_and88 | f_u_dadda_cla32_u_cla62_and91;
  assign f_u_dadda_cla32_u_cla62_or44 = f_u_dadda_cla32_u_cla62_or42 | f_u_dadda_cla32_u_cla62_or43;
  assign f_u_dadda_cla32_u_cla62_or45 = f_u_dadda_cla32_u_cla62_pg_logic19_and0 | f_u_dadda_cla32_u_cla62_or44;
  assign f_u_dadda_cla32_u_cla62_pg_logic20_or0 = f_u_dadda_cla32_fa800_xor1 | f_u_dadda_cla32_fa858_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic20_and0 = f_u_dadda_cla32_fa800_xor1 & f_u_dadda_cla32_fa858_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic20_xor0 = f_u_dadda_cla32_fa800_xor1 ^ f_u_dadda_cla32_fa858_xor1;
  assign f_u_dadda_cla32_u_cla62_xor20 = f_u_dadda_cla32_u_cla62_pg_logic20_xor0 ^ f_u_dadda_cla32_u_cla62_or45;
  assign f_u_dadda_cla32_u_cla62_and92 = f_u_dadda_cla32_u_cla62_or45 & f_u_dadda_cla32_u_cla62_pg_logic20_or0;
  assign f_u_dadda_cla32_u_cla62_or46 = f_u_dadda_cla32_u_cla62_pg_logic20_and0 | f_u_dadda_cla32_u_cla62_and92;
  assign f_u_dadda_cla32_u_cla62_pg_logic21_or0 = f_u_dadda_cla32_fa801_xor1 | f_u_dadda_cla32_fa859_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic21_and0 = f_u_dadda_cla32_fa801_xor1 & f_u_dadda_cla32_fa859_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic21_xor0 = f_u_dadda_cla32_fa801_xor1 ^ f_u_dadda_cla32_fa859_xor1;
  assign f_u_dadda_cla32_u_cla62_xor21 = f_u_dadda_cla32_u_cla62_pg_logic21_xor0 ^ f_u_dadda_cla32_u_cla62_or46;
  assign f_u_dadda_cla32_u_cla62_and93 = f_u_dadda_cla32_u_cla62_or45 & f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  assign f_u_dadda_cla32_u_cla62_and94 = f_u_dadda_cla32_u_cla62_and93 & f_u_dadda_cla32_u_cla62_pg_logic20_or0;
  assign f_u_dadda_cla32_u_cla62_and95 = f_u_dadda_cla32_u_cla62_pg_logic20_and0 & f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  assign f_u_dadda_cla32_u_cla62_or47 = f_u_dadda_cla32_u_cla62_and94 | f_u_dadda_cla32_u_cla62_and95;
  assign f_u_dadda_cla32_u_cla62_or48 = f_u_dadda_cla32_u_cla62_pg_logic21_and0 | f_u_dadda_cla32_u_cla62_or47;
  assign f_u_dadda_cla32_u_cla62_pg_logic22_or0 = f_u_dadda_cla32_fa802_xor1 | f_u_dadda_cla32_fa860_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic22_and0 = f_u_dadda_cla32_fa802_xor1 & f_u_dadda_cla32_fa860_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic22_xor0 = f_u_dadda_cla32_fa802_xor1 ^ f_u_dadda_cla32_fa860_xor1;
  assign f_u_dadda_cla32_u_cla62_xor22 = f_u_dadda_cla32_u_cla62_pg_logic22_xor0 ^ f_u_dadda_cla32_u_cla62_or48;
  assign f_u_dadda_cla32_u_cla62_and96 = f_u_dadda_cla32_u_cla62_or45 & f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  assign f_u_dadda_cla32_u_cla62_and97 = f_u_dadda_cla32_u_cla62_pg_logic22_or0 & f_u_dadda_cla32_u_cla62_pg_logic20_or0;
  assign f_u_dadda_cla32_u_cla62_and98 = f_u_dadda_cla32_u_cla62_and96 & f_u_dadda_cla32_u_cla62_and97;
  assign f_u_dadda_cla32_u_cla62_and99 = f_u_dadda_cla32_u_cla62_pg_logic20_and0 & f_u_dadda_cla32_u_cla62_pg_logic22_or0;
  assign f_u_dadda_cla32_u_cla62_and100 = f_u_dadda_cla32_u_cla62_and99 & f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  assign f_u_dadda_cla32_u_cla62_and101 = f_u_dadda_cla32_u_cla62_pg_logic21_and0 & f_u_dadda_cla32_u_cla62_pg_logic22_or0;
  assign f_u_dadda_cla32_u_cla62_or49 = f_u_dadda_cla32_u_cla62_and98 | f_u_dadda_cla32_u_cla62_and100;
  assign f_u_dadda_cla32_u_cla62_or50 = f_u_dadda_cla32_u_cla62_or49 | f_u_dadda_cla32_u_cla62_and101;
  assign f_u_dadda_cla32_u_cla62_or51 = f_u_dadda_cla32_u_cla62_pg_logic22_and0 | f_u_dadda_cla32_u_cla62_or50;
  assign f_u_dadda_cla32_u_cla62_pg_logic23_or0 = f_u_dadda_cla32_fa803_xor1 | f_u_dadda_cla32_fa861_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic23_and0 = f_u_dadda_cla32_fa803_xor1 & f_u_dadda_cla32_fa861_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic23_xor0 = f_u_dadda_cla32_fa803_xor1 ^ f_u_dadda_cla32_fa861_xor1;
  assign f_u_dadda_cla32_u_cla62_xor23 = f_u_dadda_cla32_u_cla62_pg_logic23_xor0 ^ f_u_dadda_cla32_u_cla62_or51;
  assign f_u_dadda_cla32_u_cla62_and102 = f_u_dadda_cla32_u_cla62_or45 & f_u_dadda_cla32_u_cla62_pg_logic22_or0;
  assign f_u_dadda_cla32_u_cla62_and103 = f_u_dadda_cla32_u_cla62_pg_logic23_or0 & f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  assign f_u_dadda_cla32_u_cla62_and104 = f_u_dadda_cla32_u_cla62_and102 & f_u_dadda_cla32_u_cla62_and103;
  assign f_u_dadda_cla32_u_cla62_and105 = f_u_dadda_cla32_u_cla62_and104 & f_u_dadda_cla32_u_cla62_pg_logic20_or0;
  assign f_u_dadda_cla32_u_cla62_and106 = f_u_dadda_cla32_u_cla62_pg_logic20_and0 & f_u_dadda_cla32_u_cla62_pg_logic22_or0;
  assign f_u_dadda_cla32_u_cla62_and107 = f_u_dadda_cla32_u_cla62_pg_logic23_or0 & f_u_dadda_cla32_u_cla62_pg_logic21_or0;
  assign f_u_dadda_cla32_u_cla62_and108 = f_u_dadda_cla32_u_cla62_and106 & f_u_dadda_cla32_u_cla62_and107;
  assign f_u_dadda_cla32_u_cla62_and109 = f_u_dadda_cla32_u_cla62_pg_logic21_and0 & f_u_dadda_cla32_u_cla62_pg_logic23_or0;
  assign f_u_dadda_cla32_u_cla62_and110 = f_u_dadda_cla32_u_cla62_and109 & f_u_dadda_cla32_u_cla62_pg_logic22_or0;
  assign f_u_dadda_cla32_u_cla62_and111 = f_u_dadda_cla32_u_cla62_pg_logic22_and0 & f_u_dadda_cla32_u_cla62_pg_logic23_or0;
  assign f_u_dadda_cla32_u_cla62_or52 = f_u_dadda_cla32_u_cla62_and105 | f_u_dadda_cla32_u_cla62_and110;
  assign f_u_dadda_cla32_u_cla62_or53 = f_u_dadda_cla32_u_cla62_and108 | f_u_dadda_cla32_u_cla62_and111;
  assign f_u_dadda_cla32_u_cla62_or54 = f_u_dadda_cla32_u_cla62_or52 | f_u_dadda_cla32_u_cla62_or53;
  assign f_u_dadda_cla32_u_cla62_or55 = f_u_dadda_cla32_u_cla62_pg_logic23_and0 | f_u_dadda_cla32_u_cla62_or54;
  assign f_u_dadda_cla32_u_cla62_pg_logic24_or0 = f_u_dadda_cla32_fa804_xor1 | f_u_dadda_cla32_fa862_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic24_and0 = f_u_dadda_cla32_fa804_xor1 & f_u_dadda_cla32_fa862_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic24_xor0 = f_u_dadda_cla32_fa804_xor1 ^ f_u_dadda_cla32_fa862_xor1;
  assign f_u_dadda_cla32_u_cla62_xor24 = f_u_dadda_cla32_u_cla62_pg_logic24_xor0 ^ f_u_dadda_cla32_u_cla62_or55;
  assign f_u_dadda_cla32_u_cla62_and112 = f_u_dadda_cla32_u_cla62_or55 & f_u_dadda_cla32_u_cla62_pg_logic24_or0;
  assign f_u_dadda_cla32_u_cla62_or56 = f_u_dadda_cla32_u_cla62_pg_logic24_and0 | f_u_dadda_cla32_u_cla62_and112;
  assign f_u_dadda_cla32_u_cla62_pg_logic25_or0 = f_u_dadda_cla32_fa805_xor1 | f_u_dadda_cla32_fa863_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic25_and0 = f_u_dadda_cla32_fa805_xor1 & f_u_dadda_cla32_fa863_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic25_xor0 = f_u_dadda_cla32_fa805_xor1 ^ f_u_dadda_cla32_fa863_xor1;
  assign f_u_dadda_cla32_u_cla62_xor25 = f_u_dadda_cla32_u_cla62_pg_logic25_xor0 ^ f_u_dadda_cla32_u_cla62_or56;
  assign f_u_dadda_cla32_u_cla62_and113 = f_u_dadda_cla32_u_cla62_or55 & f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  assign f_u_dadda_cla32_u_cla62_and114 = f_u_dadda_cla32_u_cla62_and113 & f_u_dadda_cla32_u_cla62_pg_logic24_or0;
  assign f_u_dadda_cla32_u_cla62_and115 = f_u_dadda_cla32_u_cla62_pg_logic24_and0 & f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  assign f_u_dadda_cla32_u_cla62_or57 = f_u_dadda_cla32_u_cla62_and114 | f_u_dadda_cla32_u_cla62_and115;
  assign f_u_dadda_cla32_u_cla62_or58 = f_u_dadda_cla32_u_cla62_pg_logic25_and0 | f_u_dadda_cla32_u_cla62_or57;
  assign f_u_dadda_cla32_u_cla62_pg_logic26_or0 = f_u_dadda_cla32_fa806_xor1 | f_u_dadda_cla32_fa864_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic26_and0 = f_u_dadda_cla32_fa806_xor1 & f_u_dadda_cla32_fa864_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic26_xor0 = f_u_dadda_cla32_fa806_xor1 ^ f_u_dadda_cla32_fa864_xor1;
  assign f_u_dadda_cla32_u_cla62_xor26 = f_u_dadda_cla32_u_cla62_pg_logic26_xor0 ^ f_u_dadda_cla32_u_cla62_or58;
  assign f_u_dadda_cla32_u_cla62_and116 = f_u_dadda_cla32_u_cla62_or55 & f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  assign f_u_dadda_cla32_u_cla62_and117 = f_u_dadda_cla32_u_cla62_pg_logic26_or0 & f_u_dadda_cla32_u_cla62_pg_logic24_or0;
  assign f_u_dadda_cla32_u_cla62_and118 = f_u_dadda_cla32_u_cla62_and116 & f_u_dadda_cla32_u_cla62_and117;
  assign f_u_dadda_cla32_u_cla62_and119 = f_u_dadda_cla32_u_cla62_pg_logic24_and0 & f_u_dadda_cla32_u_cla62_pg_logic26_or0;
  assign f_u_dadda_cla32_u_cla62_and120 = f_u_dadda_cla32_u_cla62_and119 & f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  assign f_u_dadda_cla32_u_cla62_and121 = f_u_dadda_cla32_u_cla62_pg_logic25_and0 & f_u_dadda_cla32_u_cla62_pg_logic26_or0;
  assign f_u_dadda_cla32_u_cla62_or59 = f_u_dadda_cla32_u_cla62_and118 | f_u_dadda_cla32_u_cla62_and120;
  assign f_u_dadda_cla32_u_cla62_or60 = f_u_dadda_cla32_u_cla62_or59 | f_u_dadda_cla32_u_cla62_and121;
  assign f_u_dadda_cla32_u_cla62_or61 = f_u_dadda_cla32_u_cla62_pg_logic26_and0 | f_u_dadda_cla32_u_cla62_or60;
  assign f_u_dadda_cla32_u_cla62_pg_logic27_or0 = f_u_dadda_cla32_fa807_xor1 | f_u_dadda_cla32_fa865_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic27_and0 = f_u_dadda_cla32_fa807_xor1 & f_u_dadda_cla32_fa865_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic27_xor0 = f_u_dadda_cla32_fa807_xor1 ^ f_u_dadda_cla32_fa865_xor1;
  assign f_u_dadda_cla32_u_cla62_xor27 = f_u_dadda_cla32_u_cla62_pg_logic27_xor0 ^ f_u_dadda_cla32_u_cla62_or61;
  assign f_u_dadda_cla32_u_cla62_and122 = f_u_dadda_cla32_u_cla62_or55 & f_u_dadda_cla32_u_cla62_pg_logic26_or0;
  assign f_u_dadda_cla32_u_cla62_and123 = f_u_dadda_cla32_u_cla62_pg_logic27_or0 & f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  assign f_u_dadda_cla32_u_cla62_and124 = f_u_dadda_cla32_u_cla62_and122 & f_u_dadda_cla32_u_cla62_and123;
  assign f_u_dadda_cla32_u_cla62_and125 = f_u_dadda_cla32_u_cla62_and124 & f_u_dadda_cla32_u_cla62_pg_logic24_or0;
  assign f_u_dadda_cla32_u_cla62_and126 = f_u_dadda_cla32_u_cla62_pg_logic24_and0 & f_u_dadda_cla32_u_cla62_pg_logic26_or0;
  assign f_u_dadda_cla32_u_cla62_and127 = f_u_dadda_cla32_u_cla62_pg_logic27_or0 & f_u_dadda_cla32_u_cla62_pg_logic25_or0;
  assign f_u_dadda_cla32_u_cla62_and128 = f_u_dadda_cla32_u_cla62_and126 & f_u_dadda_cla32_u_cla62_and127;
  assign f_u_dadda_cla32_u_cla62_and129 = f_u_dadda_cla32_u_cla62_pg_logic25_and0 & f_u_dadda_cla32_u_cla62_pg_logic27_or0;
  assign f_u_dadda_cla32_u_cla62_and130 = f_u_dadda_cla32_u_cla62_and129 & f_u_dadda_cla32_u_cla62_pg_logic26_or0;
  assign f_u_dadda_cla32_u_cla62_and131 = f_u_dadda_cla32_u_cla62_pg_logic26_and0 & f_u_dadda_cla32_u_cla62_pg_logic27_or0;
  assign f_u_dadda_cla32_u_cla62_or62 = f_u_dadda_cla32_u_cla62_and125 | f_u_dadda_cla32_u_cla62_and130;
  assign f_u_dadda_cla32_u_cla62_or63 = f_u_dadda_cla32_u_cla62_and128 | f_u_dadda_cla32_u_cla62_and131;
  assign f_u_dadda_cla32_u_cla62_or64 = f_u_dadda_cla32_u_cla62_or62 | f_u_dadda_cla32_u_cla62_or63;
  assign f_u_dadda_cla32_u_cla62_or65 = f_u_dadda_cla32_u_cla62_pg_logic27_and0 | f_u_dadda_cla32_u_cla62_or64;
  assign f_u_dadda_cla32_u_cla62_pg_logic28_or0 = f_u_dadda_cla32_fa808_xor1 | f_u_dadda_cla32_fa866_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic28_and0 = f_u_dadda_cla32_fa808_xor1 & f_u_dadda_cla32_fa866_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic28_xor0 = f_u_dadda_cla32_fa808_xor1 ^ f_u_dadda_cla32_fa866_xor1;
  assign f_u_dadda_cla32_u_cla62_xor28 = f_u_dadda_cla32_u_cla62_pg_logic28_xor0 ^ f_u_dadda_cla32_u_cla62_or65;
  assign f_u_dadda_cla32_u_cla62_and132 = f_u_dadda_cla32_u_cla62_or65 & f_u_dadda_cla32_u_cla62_pg_logic28_or0;
  assign f_u_dadda_cla32_u_cla62_or66 = f_u_dadda_cla32_u_cla62_pg_logic28_and0 | f_u_dadda_cla32_u_cla62_and132;
  assign f_u_dadda_cla32_u_cla62_pg_logic29_or0 = f_u_dadda_cla32_fa809_xor1 | f_u_dadda_cla32_fa867_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic29_and0 = f_u_dadda_cla32_fa809_xor1 & f_u_dadda_cla32_fa867_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic29_xor0 = f_u_dadda_cla32_fa809_xor1 ^ f_u_dadda_cla32_fa867_xor1;
  assign f_u_dadda_cla32_u_cla62_xor29 = f_u_dadda_cla32_u_cla62_pg_logic29_xor0 ^ f_u_dadda_cla32_u_cla62_or66;
  assign f_u_dadda_cla32_u_cla62_and133 = f_u_dadda_cla32_u_cla62_or65 & f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  assign f_u_dadda_cla32_u_cla62_and134 = f_u_dadda_cla32_u_cla62_and133 & f_u_dadda_cla32_u_cla62_pg_logic28_or0;
  assign f_u_dadda_cla32_u_cla62_and135 = f_u_dadda_cla32_u_cla62_pg_logic28_and0 & f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  assign f_u_dadda_cla32_u_cla62_or67 = f_u_dadda_cla32_u_cla62_and134 | f_u_dadda_cla32_u_cla62_and135;
  assign f_u_dadda_cla32_u_cla62_or68 = f_u_dadda_cla32_u_cla62_pg_logic29_and0 | f_u_dadda_cla32_u_cla62_or67;
  assign f_u_dadda_cla32_u_cla62_pg_logic30_or0 = f_u_dadda_cla32_fa810_xor1 | f_u_dadda_cla32_fa868_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic30_and0 = f_u_dadda_cla32_fa810_xor1 & f_u_dadda_cla32_fa868_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic30_xor0 = f_u_dadda_cla32_fa810_xor1 ^ f_u_dadda_cla32_fa868_xor1;
  assign f_u_dadda_cla32_u_cla62_xor30 = f_u_dadda_cla32_u_cla62_pg_logic30_xor0 ^ f_u_dadda_cla32_u_cla62_or68;
  assign f_u_dadda_cla32_u_cla62_and136 = f_u_dadda_cla32_u_cla62_or65 & f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  assign f_u_dadda_cla32_u_cla62_and137 = f_u_dadda_cla32_u_cla62_pg_logic30_or0 & f_u_dadda_cla32_u_cla62_pg_logic28_or0;
  assign f_u_dadda_cla32_u_cla62_and138 = f_u_dadda_cla32_u_cla62_and136 & f_u_dadda_cla32_u_cla62_and137;
  assign f_u_dadda_cla32_u_cla62_and139 = f_u_dadda_cla32_u_cla62_pg_logic28_and0 & f_u_dadda_cla32_u_cla62_pg_logic30_or0;
  assign f_u_dadda_cla32_u_cla62_and140 = f_u_dadda_cla32_u_cla62_and139 & f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  assign f_u_dadda_cla32_u_cla62_and141 = f_u_dadda_cla32_u_cla62_pg_logic29_and0 & f_u_dadda_cla32_u_cla62_pg_logic30_or0;
  assign f_u_dadda_cla32_u_cla62_or69 = f_u_dadda_cla32_u_cla62_and138 | f_u_dadda_cla32_u_cla62_and140;
  assign f_u_dadda_cla32_u_cla62_or70 = f_u_dadda_cla32_u_cla62_or69 | f_u_dadda_cla32_u_cla62_and141;
  assign f_u_dadda_cla32_u_cla62_or71 = f_u_dadda_cla32_u_cla62_pg_logic30_and0 | f_u_dadda_cla32_u_cla62_or70;
  assign f_u_dadda_cla32_u_cla62_pg_logic31_or0 = f_u_dadda_cla32_fa811_xor1 | f_u_dadda_cla32_fa869_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic31_and0 = f_u_dadda_cla32_fa811_xor1 & f_u_dadda_cla32_fa869_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic31_xor0 = f_u_dadda_cla32_fa811_xor1 ^ f_u_dadda_cla32_fa869_xor1;
  assign f_u_dadda_cla32_u_cla62_xor31 = f_u_dadda_cla32_u_cla62_pg_logic31_xor0 ^ f_u_dadda_cla32_u_cla62_or71;
  assign f_u_dadda_cla32_u_cla62_and142 = f_u_dadda_cla32_u_cla62_or65 & f_u_dadda_cla32_u_cla62_pg_logic30_or0;
  assign f_u_dadda_cla32_u_cla62_and143 = f_u_dadda_cla32_u_cla62_pg_logic31_or0 & f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  assign f_u_dadda_cla32_u_cla62_and144 = f_u_dadda_cla32_u_cla62_and142 & f_u_dadda_cla32_u_cla62_and143;
  assign f_u_dadda_cla32_u_cla62_and145 = f_u_dadda_cla32_u_cla62_and144 & f_u_dadda_cla32_u_cla62_pg_logic28_or0;
  assign f_u_dadda_cla32_u_cla62_and146 = f_u_dadda_cla32_u_cla62_pg_logic28_and0 & f_u_dadda_cla32_u_cla62_pg_logic30_or0;
  assign f_u_dadda_cla32_u_cla62_and147 = f_u_dadda_cla32_u_cla62_pg_logic31_or0 & f_u_dadda_cla32_u_cla62_pg_logic29_or0;
  assign f_u_dadda_cla32_u_cla62_and148 = f_u_dadda_cla32_u_cla62_and146 & f_u_dadda_cla32_u_cla62_and147;
  assign f_u_dadda_cla32_u_cla62_and149 = f_u_dadda_cla32_u_cla62_pg_logic29_and0 & f_u_dadda_cla32_u_cla62_pg_logic31_or0;
  assign f_u_dadda_cla32_u_cla62_and150 = f_u_dadda_cla32_u_cla62_and149 & f_u_dadda_cla32_u_cla62_pg_logic30_or0;
  assign f_u_dadda_cla32_u_cla62_and151 = f_u_dadda_cla32_u_cla62_pg_logic30_and0 & f_u_dadda_cla32_u_cla62_pg_logic31_or0;
  assign f_u_dadda_cla32_u_cla62_or72 = f_u_dadda_cla32_u_cla62_and145 | f_u_dadda_cla32_u_cla62_and150;
  assign f_u_dadda_cla32_u_cla62_or73 = f_u_dadda_cla32_u_cla62_and148 | f_u_dadda_cla32_u_cla62_and151;
  assign f_u_dadda_cla32_u_cla62_or74 = f_u_dadda_cla32_u_cla62_or72 | f_u_dadda_cla32_u_cla62_or73;
  assign f_u_dadda_cla32_u_cla62_or75 = f_u_dadda_cla32_u_cla62_pg_logic31_and0 | f_u_dadda_cla32_u_cla62_or74;
  assign f_u_dadda_cla32_u_cla62_pg_logic32_or0 = f_u_dadda_cla32_fa812_xor1 | f_u_dadda_cla32_fa870_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic32_and0 = f_u_dadda_cla32_fa812_xor1 & f_u_dadda_cla32_fa870_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic32_xor0 = f_u_dadda_cla32_fa812_xor1 ^ f_u_dadda_cla32_fa870_xor1;
  assign f_u_dadda_cla32_u_cla62_xor32 = f_u_dadda_cla32_u_cla62_pg_logic32_xor0 ^ f_u_dadda_cla32_u_cla62_or75;
  assign f_u_dadda_cla32_u_cla62_and152 = f_u_dadda_cla32_u_cla62_or75 & f_u_dadda_cla32_u_cla62_pg_logic32_or0;
  assign f_u_dadda_cla32_u_cla62_or76 = f_u_dadda_cla32_u_cla62_pg_logic32_and0 | f_u_dadda_cla32_u_cla62_and152;
  assign f_u_dadda_cla32_u_cla62_pg_logic33_or0 = f_u_dadda_cla32_fa813_xor1 | f_u_dadda_cla32_fa871_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic33_and0 = f_u_dadda_cla32_fa813_xor1 & f_u_dadda_cla32_fa871_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic33_xor0 = f_u_dadda_cla32_fa813_xor1 ^ f_u_dadda_cla32_fa871_xor1;
  assign f_u_dadda_cla32_u_cla62_xor33 = f_u_dadda_cla32_u_cla62_pg_logic33_xor0 ^ f_u_dadda_cla32_u_cla62_or76;
  assign f_u_dadda_cla32_u_cla62_and153 = f_u_dadda_cla32_u_cla62_or75 & f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  assign f_u_dadda_cla32_u_cla62_and154 = f_u_dadda_cla32_u_cla62_and153 & f_u_dadda_cla32_u_cla62_pg_logic32_or0;
  assign f_u_dadda_cla32_u_cla62_and155 = f_u_dadda_cla32_u_cla62_pg_logic32_and0 & f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  assign f_u_dadda_cla32_u_cla62_or77 = f_u_dadda_cla32_u_cla62_and154 | f_u_dadda_cla32_u_cla62_and155;
  assign f_u_dadda_cla32_u_cla62_or78 = f_u_dadda_cla32_u_cla62_pg_logic33_and0 | f_u_dadda_cla32_u_cla62_or77;
  assign f_u_dadda_cla32_u_cla62_pg_logic34_or0 = f_u_dadda_cla32_fa814_xor1 | f_u_dadda_cla32_fa872_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic34_and0 = f_u_dadda_cla32_fa814_xor1 & f_u_dadda_cla32_fa872_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic34_xor0 = f_u_dadda_cla32_fa814_xor1 ^ f_u_dadda_cla32_fa872_xor1;
  assign f_u_dadda_cla32_u_cla62_xor34 = f_u_dadda_cla32_u_cla62_pg_logic34_xor0 ^ f_u_dadda_cla32_u_cla62_or78;
  assign f_u_dadda_cla32_u_cla62_and156 = f_u_dadda_cla32_u_cla62_or75 & f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  assign f_u_dadda_cla32_u_cla62_and157 = f_u_dadda_cla32_u_cla62_pg_logic34_or0 & f_u_dadda_cla32_u_cla62_pg_logic32_or0;
  assign f_u_dadda_cla32_u_cla62_and158 = f_u_dadda_cla32_u_cla62_and156 & f_u_dadda_cla32_u_cla62_and157;
  assign f_u_dadda_cla32_u_cla62_and159 = f_u_dadda_cla32_u_cla62_pg_logic32_and0 & f_u_dadda_cla32_u_cla62_pg_logic34_or0;
  assign f_u_dadda_cla32_u_cla62_and160 = f_u_dadda_cla32_u_cla62_and159 & f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  assign f_u_dadda_cla32_u_cla62_and161 = f_u_dadda_cla32_u_cla62_pg_logic33_and0 & f_u_dadda_cla32_u_cla62_pg_logic34_or0;
  assign f_u_dadda_cla32_u_cla62_or79 = f_u_dadda_cla32_u_cla62_and158 | f_u_dadda_cla32_u_cla62_and160;
  assign f_u_dadda_cla32_u_cla62_or80 = f_u_dadda_cla32_u_cla62_or79 | f_u_dadda_cla32_u_cla62_and161;
  assign f_u_dadda_cla32_u_cla62_or81 = f_u_dadda_cla32_u_cla62_pg_logic34_and0 | f_u_dadda_cla32_u_cla62_or80;
  assign f_u_dadda_cla32_u_cla62_pg_logic35_or0 = f_u_dadda_cla32_fa815_xor1 | f_u_dadda_cla32_fa873_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic35_and0 = f_u_dadda_cla32_fa815_xor1 & f_u_dadda_cla32_fa873_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic35_xor0 = f_u_dadda_cla32_fa815_xor1 ^ f_u_dadda_cla32_fa873_xor1;
  assign f_u_dadda_cla32_u_cla62_xor35 = f_u_dadda_cla32_u_cla62_pg_logic35_xor0 ^ f_u_dadda_cla32_u_cla62_or81;
  assign f_u_dadda_cla32_u_cla62_and162 = f_u_dadda_cla32_u_cla62_or75 & f_u_dadda_cla32_u_cla62_pg_logic34_or0;
  assign f_u_dadda_cla32_u_cla62_and163 = f_u_dadda_cla32_u_cla62_pg_logic35_or0 & f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  assign f_u_dadda_cla32_u_cla62_and164 = f_u_dadda_cla32_u_cla62_and162 & f_u_dadda_cla32_u_cla62_and163;
  assign f_u_dadda_cla32_u_cla62_and165 = f_u_dadda_cla32_u_cla62_and164 & f_u_dadda_cla32_u_cla62_pg_logic32_or0;
  assign f_u_dadda_cla32_u_cla62_and166 = f_u_dadda_cla32_u_cla62_pg_logic32_and0 & f_u_dadda_cla32_u_cla62_pg_logic34_or0;
  assign f_u_dadda_cla32_u_cla62_and167 = f_u_dadda_cla32_u_cla62_pg_logic35_or0 & f_u_dadda_cla32_u_cla62_pg_logic33_or0;
  assign f_u_dadda_cla32_u_cla62_and168 = f_u_dadda_cla32_u_cla62_and166 & f_u_dadda_cla32_u_cla62_and167;
  assign f_u_dadda_cla32_u_cla62_and169 = f_u_dadda_cla32_u_cla62_pg_logic33_and0 & f_u_dadda_cla32_u_cla62_pg_logic35_or0;
  assign f_u_dadda_cla32_u_cla62_and170 = f_u_dadda_cla32_u_cla62_and169 & f_u_dadda_cla32_u_cla62_pg_logic34_or0;
  assign f_u_dadda_cla32_u_cla62_and171 = f_u_dadda_cla32_u_cla62_pg_logic34_and0 & f_u_dadda_cla32_u_cla62_pg_logic35_or0;
  assign f_u_dadda_cla32_u_cla62_or82 = f_u_dadda_cla32_u_cla62_and165 | f_u_dadda_cla32_u_cla62_and170;
  assign f_u_dadda_cla32_u_cla62_or83 = f_u_dadda_cla32_u_cla62_and168 | f_u_dadda_cla32_u_cla62_and171;
  assign f_u_dadda_cla32_u_cla62_or84 = f_u_dadda_cla32_u_cla62_or82 | f_u_dadda_cla32_u_cla62_or83;
  assign f_u_dadda_cla32_u_cla62_or85 = f_u_dadda_cla32_u_cla62_pg_logic35_and0 | f_u_dadda_cla32_u_cla62_or84;
  assign f_u_dadda_cla32_u_cla62_pg_logic36_or0 = f_u_dadda_cla32_fa816_xor1 | f_u_dadda_cla32_fa874_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic36_and0 = f_u_dadda_cla32_fa816_xor1 & f_u_dadda_cla32_fa874_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic36_xor0 = f_u_dadda_cla32_fa816_xor1 ^ f_u_dadda_cla32_fa874_xor1;
  assign f_u_dadda_cla32_u_cla62_xor36 = f_u_dadda_cla32_u_cla62_pg_logic36_xor0 ^ f_u_dadda_cla32_u_cla62_or85;
  assign f_u_dadda_cla32_u_cla62_and172 = f_u_dadda_cla32_u_cla62_or85 & f_u_dadda_cla32_u_cla62_pg_logic36_or0;
  assign f_u_dadda_cla32_u_cla62_or86 = f_u_dadda_cla32_u_cla62_pg_logic36_and0 | f_u_dadda_cla32_u_cla62_and172;
  assign f_u_dadda_cla32_u_cla62_pg_logic37_or0 = f_u_dadda_cla32_fa817_xor1 | f_u_dadda_cla32_fa875_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic37_and0 = f_u_dadda_cla32_fa817_xor1 & f_u_dadda_cla32_fa875_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic37_xor0 = f_u_dadda_cla32_fa817_xor1 ^ f_u_dadda_cla32_fa875_xor1;
  assign f_u_dadda_cla32_u_cla62_xor37 = f_u_dadda_cla32_u_cla62_pg_logic37_xor0 ^ f_u_dadda_cla32_u_cla62_or86;
  assign f_u_dadda_cla32_u_cla62_and173 = f_u_dadda_cla32_u_cla62_or85 & f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  assign f_u_dadda_cla32_u_cla62_and174 = f_u_dadda_cla32_u_cla62_and173 & f_u_dadda_cla32_u_cla62_pg_logic36_or0;
  assign f_u_dadda_cla32_u_cla62_and175 = f_u_dadda_cla32_u_cla62_pg_logic36_and0 & f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  assign f_u_dadda_cla32_u_cla62_or87 = f_u_dadda_cla32_u_cla62_and174 | f_u_dadda_cla32_u_cla62_and175;
  assign f_u_dadda_cla32_u_cla62_or88 = f_u_dadda_cla32_u_cla62_pg_logic37_and0 | f_u_dadda_cla32_u_cla62_or87;
  assign f_u_dadda_cla32_u_cla62_pg_logic38_or0 = f_u_dadda_cla32_fa818_xor1 | f_u_dadda_cla32_fa876_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic38_and0 = f_u_dadda_cla32_fa818_xor1 & f_u_dadda_cla32_fa876_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic38_xor0 = f_u_dadda_cla32_fa818_xor1 ^ f_u_dadda_cla32_fa876_xor1;
  assign f_u_dadda_cla32_u_cla62_xor38 = f_u_dadda_cla32_u_cla62_pg_logic38_xor0 ^ f_u_dadda_cla32_u_cla62_or88;
  assign f_u_dadda_cla32_u_cla62_and176 = f_u_dadda_cla32_u_cla62_or85 & f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  assign f_u_dadda_cla32_u_cla62_and177 = f_u_dadda_cla32_u_cla62_pg_logic38_or0 & f_u_dadda_cla32_u_cla62_pg_logic36_or0;
  assign f_u_dadda_cla32_u_cla62_and178 = f_u_dadda_cla32_u_cla62_and176 & f_u_dadda_cla32_u_cla62_and177;
  assign f_u_dadda_cla32_u_cla62_and179 = f_u_dadda_cla32_u_cla62_pg_logic36_and0 & f_u_dadda_cla32_u_cla62_pg_logic38_or0;
  assign f_u_dadda_cla32_u_cla62_and180 = f_u_dadda_cla32_u_cla62_and179 & f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  assign f_u_dadda_cla32_u_cla62_and181 = f_u_dadda_cla32_u_cla62_pg_logic37_and0 & f_u_dadda_cla32_u_cla62_pg_logic38_or0;
  assign f_u_dadda_cla32_u_cla62_or89 = f_u_dadda_cla32_u_cla62_and178 | f_u_dadda_cla32_u_cla62_and180;
  assign f_u_dadda_cla32_u_cla62_or90 = f_u_dadda_cla32_u_cla62_or89 | f_u_dadda_cla32_u_cla62_and181;
  assign f_u_dadda_cla32_u_cla62_or91 = f_u_dadda_cla32_u_cla62_pg_logic38_and0 | f_u_dadda_cla32_u_cla62_or90;
  assign f_u_dadda_cla32_u_cla62_pg_logic39_or0 = f_u_dadda_cla32_fa819_xor1 | f_u_dadda_cla32_fa877_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic39_and0 = f_u_dadda_cla32_fa819_xor1 & f_u_dadda_cla32_fa877_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic39_xor0 = f_u_dadda_cla32_fa819_xor1 ^ f_u_dadda_cla32_fa877_xor1;
  assign f_u_dadda_cla32_u_cla62_xor39 = f_u_dadda_cla32_u_cla62_pg_logic39_xor0 ^ f_u_dadda_cla32_u_cla62_or91;
  assign f_u_dadda_cla32_u_cla62_and182 = f_u_dadda_cla32_u_cla62_or85 & f_u_dadda_cla32_u_cla62_pg_logic38_or0;
  assign f_u_dadda_cla32_u_cla62_and183 = f_u_dadda_cla32_u_cla62_pg_logic39_or0 & f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  assign f_u_dadda_cla32_u_cla62_and184 = f_u_dadda_cla32_u_cla62_and182 & f_u_dadda_cla32_u_cla62_and183;
  assign f_u_dadda_cla32_u_cla62_and185 = f_u_dadda_cla32_u_cla62_and184 & f_u_dadda_cla32_u_cla62_pg_logic36_or0;
  assign f_u_dadda_cla32_u_cla62_and186 = f_u_dadda_cla32_u_cla62_pg_logic36_and0 & f_u_dadda_cla32_u_cla62_pg_logic38_or0;
  assign f_u_dadda_cla32_u_cla62_and187 = f_u_dadda_cla32_u_cla62_pg_logic39_or0 & f_u_dadda_cla32_u_cla62_pg_logic37_or0;
  assign f_u_dadda_cla32_u_cla62_and188 = f_u_dadda_cla32_u_cla62_and186 & f_u_dadda_cla32_u_cla62_and187;
  assign f_u_dadda_cla32_u_cla62_and189 = f_u_dadda_cla32_u_cla62_pg_logic37_and0 & f_u_dadda_cla32_u_cla62_pg_logic39_or0;
  assign f_u_dadda_cla32_u_cla62_and190 = f_u_dadda_cla32_u_cla62_and189 & f_u_dadda_cla32_u_cla62_pg_logic38_or0;
  assign f_u_dadda_cla32_u_cla62_and191 = f_u_dadda_cla32_u_cla62_pg_logic38_and0 & f_u_dadda_cla32_u_cla62_pg_logic39_or0;
  assign f_u_dadda_cla32_u_cla62_or92 = f_u_dadda_cla32_u_cla62_and185 | f_u_dadda_cla32_u_cla62_and190;
  assign f_u_dadda_cla32_u_cla62_or93 = f_u_dadda_cla32_u_cla62_and188 | f_u_dadda_cla32_u_cla62_and191;
  assign f_u_dadda_cla32_u_cla62_or94 = f_u_dadda_cla32_u_cla62_or92 | f_u_dadda_cla32_u_cla62_or93;
  assign f_u_dadda_cla32_u_cla62_or95 = f_u_dadda_cla32_u_cla62_pg_logic39_and0 | f_u_dadda_cla32_u_cla62_or94;
  assign f_u_dadda_cla32_u_cla62_pg_logic40_or0 = f_u_dadda_cla32_fa820_xor1 | f_u_dadda_cla32_fa878_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic40_and0 = f_u_dadda_cla32_fa820_xor1 & f_u_dadda_cla32_fa878_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic40_xor0 = f_u_dadda_cla32_fa820_xor1 ^ f_u_dadda_cla32_fa878_xor1;
  assign f_u_dadda_cla32_u_cla62_xor40 = f_u_dadda_cla32_u_cla62_pg_logic40_xor0 ^ f_u_dadda_cla32_u_cla62_or95;
  assign f_u_dadda_cla32_u_cla62_and192 = f_u_dadda_cla32_u_cla62_or95 & f_u_dadda_cla32_u_cla62_pg_logic40_or0;
  assign f_u_dadda_cla32_u_cla62_or96 = f_u_dadda_cla32_u_cla62_pg_logic40_and0 | f_u_dadda_cla32_u_cla62_and192;
  assign f_u_dadda_cla32_u_cla62_pg_logic41_or0 = f_u_dadda_cla32_fa821_xor1 | f_u_dadda_cla32_fa879_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic41_and0 = f_u_dadda_cla32_fa821_xor1 & f_u_dadda_cla32_fa879_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic41_xor0 = f_u_dadda_cla32_fa821_xor1 ^ f_u_dadda_cla32_fa879_xor1;
  assign f_u_dadda_cla32_u_cla62_xor41 = f_u_dadda_cla32_u_cla62_pg_logic41_xor0 ^ f_u_dadda_cla32_u_cla62_or96;
  assign f_u_dadda_cla32_u_cla62_and193 = f_u_dadda_cla32_u_cla62_or95 & f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  assign f_u_dadda_cla32_u_cla62_and194 = f_u_dadda_cla32_u_cla62_and193 & f_u_dadda_cla32_u_cla62_pg_logic40_or0;
  assign f_u_dadda_cla32_u_cla62_and195 = f_u_dadda_cla32_u_cla62_pg_logic40_and0 & f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  assign f_u_dadda_cla32_u_cla62_or97 = f_u_dadda_cla32_u_cla62_and194 | f_u_dadda_cla32_u_cla62_and195;
  assign f_u_dadda_cla32_u_cla62_or98 = f_u_dadda_cla32_u_cla62_pg_logic41_and0 | f_u_dadda_cla32_u_cla62_or97;
  assign f_u_dadda_cla32_u_cla62_pg_logic42_or0 = f_u_dadda_cla32_fa822_xor1 | f_u_dadda_cla32_fa880_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic42_and0 = f_u_dadda_cla32_fa822_xor1 & f_u_dadda_cla32_fa880_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic42_xor0 = f_u_dadda_cla32_fa822_xor1 ^ f_u_dadda_cla32_fa880_xor1;
  assign f_u_dadda_cla32_u_cla62_xor42 = f_u_dadda_cla32_u_cla62_pg_logic42_xor0 ^ f_u_dadda_cla32_u_cla62_or98;
  assign f_u_dadda_cla32_u_cla62_and196 = f_u_dadda_cla32_u_cla62_or95 & f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  assign f_u_dadda_cla32_u_cla62_and197 = f_u_dadda_cla32_u_cla62_pg_logic42_or0 & f_u_dadda_cla32_u_cla62_pg_logic40_or0;
  assign f_u_dadda_cla32_u_cla62_and198 = f_u_dadda_cla32_u_cla62_and196 & f_u_dadda_cla32_u_cla62_and197;
  assign f_u_dadda_cla32_u_cla62_and199 = f_u_dadda_cla32_u_cla62_pg_logic40_and0 & f_u_dadda_cla32_u_cla62_pg_logic42_or0;
  assign f_u_dadda_cla32_u_cla62_and200 = f_u_dadda_cla32_u_cla62_and199 & f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  assign f_u_dadda_cla32_u_cla62_and201 = f_u_dadda_cla32_u_cla62_pg_logic41_and0 & f_u_dadda_cla32_u_cla62_pg_logic42_or0;
  assign f_u_dadda_cla32_u_cla62_or99 = f_u_dadda_cla32_u_cla62_and198 | f_u_dadda_cla32_u_cla62_and200;
  assign f_u_dadda_cla32_u_cla62_or100 = f_u_dadda_cla32_u_cla62_or99 | f_u_dadda_cla32_u_cla62_and201;
  assign f_u_dadda_cla32_u_cla62_or101 = f_u_dadda_cla32_u_cla62_pg_logic42_and0 | f_u_dadda_cla32_u_cla62_or100;
  assign f_u_dadda_cla32_u_cla62_pg_logic43_or0 = f_u_dadda_cla32_fa823_xor1 | f_u_dadda_cla32_fa881_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic43_and0 = f_u_dadda_cla32_fa823_xor1 & f_u_dadda_cla32_fa881_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic43_xor0 = f_u_dadda_cla32_fa823_xor1 ^ f_u_dadda_cla32_fa881_xor1;
  assign f_u_dadda_cla32_u_cla62_xor43 = f_u_dadda_cla32_u_cla62_pg_logic43_xor0 ^ f_u_dadda_cla32_u_cla62_or101;
  assign f_u_dadda_cla32_u_cla62_and202 = f_u_dadda_cla32_u_cla62_or95 & f_u_dadda_cla32_u_cla62_pg_logic42_or0;
  assign f_u_dadda_cla32_u_cla62_and203 = f_u_dadda_cla32_u_cla62_pg_logic43_or0 & f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  assign f_u_dadda_cla32_u_cla62_and204 = f_u_dadda_cla32_u_cla62_and202 & f_u_dadda_cla32_u_cla62_and203;
  assign f_u_dadda_cla32_u_cla62_and205 = f_u_dadda_cla32_u_cla62_and204 & f_u_dadda_cla32_u_cla62_pg_logic40_or0;
  assign f_u_dadda_cla32_u_cla62_and206 = f_u_dadda_cla32_u_cla62_pg_logic40_and0 & f_u_dadda_cla32_u_cla62_pg_logic42_or0;
  assign f_u_dadda_cla32_u_cla62_and207 = f_u_dadda_cla32_u_cla62_pg_logic43_or0 & f_u_dadda_cla32_u_cla62_pg_logic41_or0;
  assign f_u_dadda_cla32_u_cla62_and208 = f_u_dadda_cla32_u_cla62_and206 & f_u_dadda_cla32_u_cla62_and207;
  assign f_u_dadda_cla32_u_cla62_and209 = f_u_dadda_cla32_u_cla62_pg_logic41_and0 & f_u_dadda_cla32_u_cla62_pg_logic43_or0;
  assign f_u_dadda_cla32_u_cla62_and210 = f_u_dadda_cla32_u_cla62_and209 & f_u_dadda_cla32_u_cla62_pg_logic42_or0;
  assign f_u_dadda_cla32_u_cla62_and211 = f_u_dadda_cla32_u_cla62_pg_logic42_and0 & f_u_dadda_cla32_u_cla62_pg_logic43_or0;
  assign f_u_dadda_cla32_u_cla62_or102 = f_u_dadda_cla32_u_cla62_and205 | f_u_dadda_cla32_u_cla62_and210;
  assign f_u_dadda_cla32_u_cla62_or103 = f_u_dadda_cla32_u_cla62_and208 | f_u_dadda_cla32_u_cla62_and211;
  assign f_u_dadda_cla32_u_cla62_or104 = f_u_dadda_cla32_u_cla62_or102 | f_u_dadda_cla32_u_cla62_or103;
  assign f_u_dadda_cla32_u_cla62_or105 = f_u_dadda_cla32_u_cla62_pg_logic43_and0 | f_u_dadda_cla32_u_cla62_or104;
  assign f_u_dadda_cla32_u_cla62_pg_logic44_or0 = f_u_dadda_cla32_fa824_xor1 | f_u_dadda_cla32_fa882_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic44_and0 = f_u_dadda_cla32_fa824_xor1 & f_u_dadda_cla32_fa882_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic44_xor0 = f_u_dadda_cla32_fa824_xor1 ^ f_u_dadda_cla32_fa882_xor1;
  assign f_u_dadda_cla32_u_cla62_xor44 = f_u_dadda_cla32_u_cla62_pg_logic44_xor0 ^ f_u_dadda_cla32_u_cla62_or105;
  assign f_u_dadda_cla32_u_cla62_and212 = f_u_dadda_cla32_u_cla62_or105 & f_u_dadda_cla32_u_cla62_pg_logic44_or0;
  assign f_u_dadda_cla32_u_cla62_or106 = f_u_dadda_cla32_u_cla62_pg_logic44_and0 | f_u_dadda_cla32_u_cla62_and212;
  assign f_u_dadda_cla32_u_cla62_pg_logic45_or0 = f_u_dadda_cla32_fa825_xor1 | f_u_dadda_cla32_fa883_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic45_and0 = f_u_dadda_cla32_fa825_xor1 & f_u_dadda_cla32_fa883_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic45_xor0 = f_u_dadda_cla32_fa825_xor1 ^ f_u_dadda_cla32_fa883_xor1;
  assign f_u_dadda_cla32_u_cla62_xor45 = f_u_dadda_cla32_u_cla62_pg_logic45_xor0 ^ f_u_dadda_cla32_u_cla62_or106;
  assign f_u_dadda_cla32_u_cla62_and213 = f_u_dadda_cla32_u_cla62_or105 & f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  assign f_u_dadda_cla32_u_cla62_and214 = f_u_dadda_cla32_u_cla62_and213 & f_u_dadda_cla32_u_cla62_pg_logic44_or0;
  assign f_u_dadda_cla32_u_cla62_and215 = f_u_dadda_cla32_u_cla62_pg_logic44_and0 & f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  assign f_u_dadda_cla32_u_cla62_or107 = f_u_dadda_cla32_u_cla62_and214 | f_u_dadda_cla32_u_cla62_and215;
  assign f_u_dadda_cla32_u_cla62_or108 = f_u_dadda_cla32_u_cla62_pg_logic45_and0 | f_u_dadda_cla32_u_cla62_or107;
  assign f_u_dadda_cla32_u_cla62_pg_logic46_or0 = f_u_dadda_cla32_fa826_xor1 | f_u_dadda_cla32_fa884_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic46_and0 = f_u_dadda_cla32_fa826_xor1 & f_u_dadda_cla32_fa884_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic46_xor0 = f_u_dadda_cla32_fa826_xor1 ^ f_u_dadda_cla32_fa884_xor1;
  assign f_u_dadda_cla32_u_cla62_xor46 = f_u_dadda_cla32_u_cla62_pg_logic46_xor0 ^ f_u_dadda_cla32_u_cla62_or108;
  assign f_u_dadda_cla32_u_cla62_and216 = f_u_dadda_cla32_u_cla62_or105 & f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  assign f_u_dadda_cla32_u_cla62_and217 = f_u_dadda_cla32_u_cla62_pg_logic46_or0 & f_u_dadda_cla32_u_cla62_pg_logic44_or0;
  assign f_u_dadda_cla32_u_cla62_and218 = f_u_dadda_cla32_u_cla62_and216 & f_u_dadda_cla32_u_cla62_and217;
  assign f_u_dadda_cla32_u_cla62_and219 = f_u_dadda_cla32_u_cla62_pg_logic44_and0 & f_u_dadda_cla32_u_cla62_pg_logic46_or0;
  assign f_u_dadda_cla32_u_cla62_and220 = f_u_dadda_cla32_u_cla62_and219 & f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  assign f_u_dadda_cla32_u_cla62_and221 = f_u_dadda_cla32_u_cla62_pg_logic45_and0 & f_u_dadda_cla32_u_cla62_pg_logic46_or0;
  assign f_u_dadda_cla32_u_cla62_or109 = f_u_dadda_cla32_u_cla62_and218 | f_u_dadda_cla32_u_cla62_and220;
  assign f_u_dadda_cla32_u_cla62_or110 = f_u_dadda_cla32_u_cla62_or109 | f_u_dadda_cla32_u_cla62_and221;
  assign f_u_dadda_cla32_u_cla62_or111 = f_u_dadda_cla32_u_cla62_pg_logic46_and0 | f_u_dadda_cla32_u_cla62_or110;
  assign f_u_dadda_cla32_u_cla62_pg_logic47_or0 = f_u_dadda_cla32_fa827_xor1 | f_u_dadda_cla32_fa885_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic47_and0 = f_u_dadda_cla32_fa827_xor1 & f_u_dadda_cla32_fa885_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic47_xor0 = f_u_dadda_cla32_fa827_xor1 ^ f_u_dadda_cla32_fa885_xor1;
  assign f_u_dadda_cla32_u_cla62_xor47 = f_u_dadda_cla32_u_cla62_pg_logic47_xor0 ^ f_u_dadda_cla32_u_cla62_or111;
  assign f_u_dadda_cla32_u_cla62_and222 = f_u_dadda_cla32_u_cla62_or105 & f_u_dadda_cla32_u_cla62_pg_logic46_or0;
  assign f_u_dadda_cla32_u_cla62_and223 = f_u_dadda_cla32_u_cla62_pg_logic47_or0 & f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  assign f_u_dadda_cla32_u_cla62_and224 = f_u_dadda_cla32_u_cla62_and222 & f_u_dadda_cla32_u_cla62_and223;
  assign f_u_dadda_cla32_u_cla62_and225 = f_u_dadda_cla32_u_cla62_and224 & f_u_dadda_cla32_u_cla62_pg_logic44_or0;
  assign f_u_dadda_cla32_u_cla62_and226 = f_u_dadda_cla32_u_cla62_pg_logic44_and0 & f_u_dadda_cla32_u_cla62_pg_logic46_or0;
  assign f_u_dadda_cla32_u_cla62_and227 = f_u_dadda_cla32_u_cla62_pg_logic47_or0 & f_u_dadda_cla32_u_cla62_pg_logic45_or0;
  assign f_u_dadda_cla32_u_cla62_and228 = f_u_dadda_cla32_u_cla62_and226 & f_u_dadda_cla32_u_cla62_and227;
  assign f_u_dadda_cla32_u_cla62_and229 = f_u_dadda_cla32_u_cla62_pg_logic45_and0 & f_u_dadda_cla32_u_cla62_pg_logic47_or0;
  assign f_u_dadda_cla32_u_cla62_and230 = f_u_dadda_cla32_u_cla62_and229 & f_u_dadda_cla32_u_cla62_pg_logic46_or0;
  assign f_u_dadda_cla32_u_cla62_and231 = f_u_dadda_cla32_u_cla62_pg_logic46_and0 & f_u_dadda_cla32_u_cla62_pg_logic47_or0;
  assign f_u_dadda_cla32_u_cla62_or112 = f_u_dadda_cla32_u_cla62_and225 | f_u_dadda_cla32_u_cla62_and230;
  assign f_u_dadda_cla32_u_cla62_or113 = f_u_dadda_cla32_u_cla62_and228 | f_u_dadda_cla32_u_cla62_and231;
  assign f_u_dadda_cla32_u_cla62_or114 = f_u_dadda_cla32_u_cla62_or112 | f_u_dadda_cla32_u_cla62_or113;
  assign f_u_dadda_cla32_u_cla62_or115 = f_u_dadda_cla32_u_cla62_pg_logic47_and0 | f_u_dadda_cla32_u_cla62_or114;
  assign f_u_dadda_cla32_u_cla62_pg_logic48_or0 = f_u_dadda_cla32_fa828_xor1 | f_u_dadda_cla32_fa886_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic48_and0 = f_u_dadda_cla32_fa828_xor1 & f_u_dadda_cla32_fa886_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic48_xor0 = f_u_dadda_cla32_fa828_xor1 ^ f_u_dadda_cla32_fa886_xor1;
  assign f_u_dadda_cla32_u_cla62_xor48 = f_u_dadda_cla32_u_cla62_pg_logic48_xor0 ^ f_u_dadda_cla32_u_cla62_or115;
  assign f_u_dadda_cla32_u_cla62_and232 = f_u_dadda_cla32_u_cla62_or115 & f_u_dadda_cla32_u_cla62_pg_logic48_or0;
  assign f_u_dadda_cla32_u_cla62_or116 = f_u_dadda_cla32_u_cla62_pg_logic48_and0 | f_u_dadda_cla32_u_cla62_and232;
  assign f_u_dadda_cla32_u_cla62_pg_logic49_or0 = f_u_dadda_cla32_fa829_xor1 | f_u_dadda_cla32_fa887_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic49_and0 = f_u_dadda_cla32_fa829_xor1 & f_u_dadda_cla32_fa887_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic49_xor0 = f_u_dadda_cla32_fa829_xor1 ^ f_u_dadda_cla32_fa887_xor1;
  assign f_u_dadda_cla32_u_cla62_xor49 = f_u_dadda_cla32_u_cla62_pg_logic49_xor0 ^ f_u_dadda_cla32_u_cla62_or116;
  assign f_u_dadda_cla32_u_cla62_and233 = f_u_dadda_cla32_u_cla62_or115 & f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  assign f_u_dadda_cla32_u_cla62_and234 = f_u_dadda_cla32_u_cla62_and233 & f_u_dadda_cla32_u_cla62_pg_logic48_or0;
  assign f_u_dadda_cla32_u_cla62_and235 = f_u_dadda_cla32_u_cla62_pg_logic48_and0 & f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  assign f_u_dadda_cla32_u_cla62_or117 = f_u_dadda_cla32_u_cla62_and234 | f_u_dadda_cla32_u_cla62_and235;
  assign f_u_dadda_cla32_u_cla62_or118 = f_u_dadda_cla32_u_cla62_pg_logic49_and0 | f_u_dadda_cla32_u_cla62_or117;
  assign f_u_dadda_cla32_u_cla62_pg_logic50_or0 = f_u_dadda_cla32_fa830_xor1 | f_u_dadda_cla32_fa888_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic50_and0 = f_u_dadda_cla32_fa830_xor1 & f_u_dadda_cla32_fa888_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic50_xor0 = f_u_dadda_cla32_fa830_xor1 ^ f_u_dadda_cla32_fa888_xor1;
  assign f_u_dadda_cla32_u_cla62_xor50 = f_u_dadda_cla32_u_cla62_pg_logic50_xor0 ^ f_u_dadda_cla32_u_cla62_or118;
  assign f_u_dadda_cla32_u_cla62_and236 = f_u_dadda_cla32_u_cla62_or115 & f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  assign f_u_dadda_cla32_u_cla62_and237 = f_u_dadda_cla32_u_cla62_pg_logic50_or0 & f_u_dadda_cla32_u_cla62_pg_logic48_or0;
  assign f_u_dadda_cla32_u_cla62_and238 = f_u_dadda_cla32_u_cla62_and236 & f_u_dadda_cla32_u_cla62_and237;
  assign f_u_dadda_cla32_u_cla62_and239 = f_u_dadda_cla32_u_cla62_pg_logic48_and0 & f_u_dadda_cla32_u_cla62_pg_logic50_or0;
  assign f_u_dadda_cla32_u_cla62_and240 = f_u_dadda_cla32_u_cla62_and239 & f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  assign f_u_dadda_cla32_u_cla62_and241 = f_u_dadda_cla32_u_cla62_pg_logic49_and0 & f_u_dadda_cla32_u_cla62_pg_logic50_or0;
  assign f_u_dadda_cla32_u_cla62_or119 = f_u_dadda_cla32_u_cla62_and238 | f_u_dadda_cla32_u_cla62_and240;
  assign f_u_dadda_cla32_u_cla62_or120 = f_u_dadda_cla32_u_cla62_or119 | f_u_dadda_cla32_u_cla62_and241;
  assign f_u_dadda_cla32_u_cla62_or121 = f_u_dadda_cla32_u_cla62_pg_logic50_and0 | f_u_dadda_cla32_u_cla62_or120;
  assign f_u_dadda_cla32_u_cla62_pg_logic51_or0 = f_u_dadda_cla32_fa831_xor1 | f_u_dadda_cla32_fa889_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic51_and0 = f_u_dadda_cla32_fa831_xor1 & f_u_dadda_cla32_fa889_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic51_xor0 = f_u_dadda_cla32_fa831_xor1 ^ f_u_dadda_cla32_fa889_xor1;
  assign f_u_dadda_cla32_u_cla62_xor51 = f_u_dadda_cla32_u_cla62_pg_logic51_xor0 ^ f_u_dadda_cla32_u_cla62_or121;
  assign f_u_dadda_cla32_u_cla62_and242 = f_u_dadda_cla32_u_cla62_or115 & f_u_dadda_cla32_u_cla62_pg_logic50_or0;
  assign f_u_dadda_cla32_u_cla62_and243 = f_u_dadda_cla32_u_cla62_pg_logic51_or0 & f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  assign f_u_dadda_cla32_u_cla62_and244 = f_u_dadda_cla32_u_cla62_and242 & f_u_dadda_cla32_u_cla62_and243;
  assign f_u_dadda_cla32_u_cla62_and245 = f_u_dadda_cla32_u_cla62_and244 & f_u_dadda_cla32_u_cla62_pg_logic48_or0;
  assign f_u_dadda_cla32_u_cla62_and246 = f_u_dadda_cla32_u_cla62_pg_logic48_and0 & f_u_dadda_cla32_u_cla62_pg_logic50_or0;
  assign f_u_dadda_cla32_u_cla62_and247 = f_u_dadda_cla32_u_cla62_pg_logic51_or0 & f_u_dadda_cla32_u_cla62_pg_logic49_or0;
  assign f_u_dadda_cla32_u_cla62_and248 = f_u_dadda_cla32_u_cla62_and246 & f_u_dadda_cla32_u_cla62_and247;
  assign f_u_dadda_cla32_u_cla62_and249 = f_u_dadda_cla32_u_cla62_pg_logic49_and0 & f_u_dadda_cla32_u_cla62_pg_logic51_or0;
  assign f_u_dadda_cla32_u_cla62_and250 = f_u_dadda_cla32_u_cla62_and249 & f_u_dadda_cla32_u_cla62_pg_logic50_or0;
  assign f_u_dadda_cla32_u_cla62_and251 = f_u_dadda_cla32_u_cla62_pg_logic50_and0 & f_u_dadda_cla32_u_cla62_pg_logic51_or0;
  assign f_u_dadda_cla32_u_cla62_or122 = f_u_dadda_cla32_u_cla62_and245 | f_u_dadda_cla32_u_cla62_and250;
  assign f_u_dadda_cla32_u_cla62_or123 = f_u_dadda_cla32_u_cla62_and248 | f_u_dadda_cla32_u_cla62_and251;
  assign f_u_dadda_cla32_u_cla62_or124 = f_u_dadda_cla32_u_cla62_or122 | f_u_dadda_cla32_u_cla62_or123;
  assign f_u_dadda_cla32_u_cla62_or125 = f_u_dadda_cla32_u_cla62_pg_logic51_and0 | f_u_dadda_cla32_u_cla62_or124;
  assign f_u_dadda_cla32_u_cla62_pg_logic52_or0 = f_u_dadda_cla32_fa832_xor1 | f_u_dadda_cla32_fa890_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic52_and0 = f_u_dadda_cla32_fa832_xor1 & f_u_dadda_cla32_fa890_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic52_xor0 = f_u_dadda_cla32_fa832_xor1 ^ f_u_dadda_cla32_fa890_xor1;
  assign f_u_dadda_cla32_u_cla62_xor52 = f_u_dadda_cla32_u_cla62_pg_logic52_xor0 ^ f_u_dadda_cla32_u_cla62_or125;
  assign f_u_dadda_cla32_u_cla62_and252 = f_u_dadda_cla32_u_cla62_or125 & f_u_dadda_cla32_u_cla62_pg_logic52_or0;
  assign f_u_dadda_cla32_u_cla62_or126 = f_u_dadda_cla32_u_cla62_pg_logic52_and0 | f_u_dadda_cla32_u_cla62_and252;
  assign f_u_dadda_cla32_u_cla62_pg_logic53_or0 = f_u_dadda_cla32_fa833_xor1 | f_u_dadda_cla32_fa891_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic53_and0 = f_u_dadda_cla32_fa833_xor1 & f_u_dadda_cla32_fa891_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic53_xor0 = f_u_dadda_cla32_fa833_xor1 ^ f_u_dadda_cla32_fa891_xor1;
  assign f_u_dadda_cla32_u_cla62_xor53 = f_u_dadda_cla32_u_cla62_pg_logic53_xor0 ^ f_u_dadda_cla32_u_cla62_or126;
  assign f_u_dadda_cla32_u_cla62_and253 = f_u_dadda_cla32_u_cla62_or125 & f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  assign f_u_dadda_cla32_u_cla62_and254 = f_u_dadda_cla32_u_cla62_and253 & f_u_dadda_cla32_u_cla62_pg_logic52_or0;
  assign f_u_dadda_cla32_u_cla62_and255 = f_u_dadda_cla32_u_cla62_pg_logic52_and0 & f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  assign f_u_dadda_cla32_u_cla62_or127 = f_u_dadda_cla32_u_cla62_and254 | f_u_dadda_cla32_u_cla62_and255;
  assign f_u_dadda_cla32_u_cla62_or128 = f_u_dadda_cla32_u_cla62_pg_logic53_and0 | f_u_dadda_cla32_u_cla62_or127;
  assign f_u_dadda_cla32_u_cla62_pg_logic54_or0 = f_u_dadda_cla32_fa834_xor1 | f_u_dadda_cla32_fa892_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic54_and0 = f_u_dadda_cla32_fa834_xor1 & f_u_dadda_cla32_fa892_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic54_xor0 = f_u_dadda_cla32_fa834_xor1 ^ f_u_dadda_cla32_fa892_xor1;
  assign f_u_dadda_cla32_u_cla62_xor54 = f_u_dadda_cla32_u_cla62_pg_logic54_xor0 ^ f_u_dadda_cla32_u_cla62_or128;
  assign f_u_dadda_cla32_u_cla62_and256 = f_u_dadda_cla32_u_cla62_or125 & f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  assign f_u_dadda_cla32_u_cla62_and257 = f_u_dadda_cla32_u_cla62_pg_logic54_or0 & f_u_dadda_cla32_u_cla62_pg_logic52_or0;
  assign f_u_dadda_cla32_u_cla62_and258 = f_u_dadda_cla32_u_cla62_and256 & f_u_dadda_cla32_u_cla62_and257;
  assign f_u_dadda_cla32_u_cla62_and259 = f_u_dadda_cla32_u_cla62_pg_logic52_and0 & f_u_dadda_cla32_u_cla62_pg_logic54_or0;
  assign f_u_dadda_cla32_u_cla62_and260 = f_u_dadda_cla32_u_cla62_and259 & f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  assign f_u_dadda_cla32_u_cla62_and261 = f_u_dadda_cla32_u_cla62_pg_logic53_and0 & f_u_dadda_cla32_u_cla62_pg_logic54_or0;
  assign f_u_dadda_cla32_u_cla62_or129 = f_u_dadda_cla32_u_cla62_and258 | f_u_dadda_cla32_u_cla62_and260;
  assign f_u_dadda_cla32_u_cla62_or130 = f_u_dadda_cla32_u_cla62_or129 | f_u_dadda_cla32_u_cla62_and261;
  assign f_u_dadda_cla32_u_cla62_or131 = f_u_dadda_cla32_u_cla62_pg_logic54_and0 | f_u_dadda_cla32_u_cla62_or130;
  assign f_u_dadda_cla32_u_cla62_pg_logic55_or0 = f_u_dadda_cla32_fa835_xor1 | f_u_dadda_cla32_fa893_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic55_and0 = f_u_dadda_cla32_fa835_xor1 & f_u_dadda_cla32_fa893_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic55_xor0 = f_u_dadda_cla32_fa835_xor1 ^ f_u_dadda_cla32_fa893_xor1;
  assign f_u_dadda_cla32_u_cla62_xor55 = f_u_dadda_cla32_u_cla62_pg_logic55_xor0 ^ f_u_dadda_cla32_u_cla62_or131;
  assign f_u_dadda_cla32_u_cla62_and262 = f_u_dadda_cla32_u_cla62_or125 & f_u_dadda_cla32_u_cla62_pg_logic54_or0;
  assign f_u_dadda_cla32_u_cla62_and263 = f_u_dadda_cla32_u_cla62_pg_logic55_or0 & f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  assign f_u_dadda_cla32_u_cla62_and264 = f_u_dadda_cla32_u_cla62_and262 & f_u_dadda_cla32_u_cla62_and263;
  assign f_u_dadda_cla32_u_cla62_and265 = f_u_dadda_cla32_u_cla62_and264 & f_u_dadda_cla32_u_cla62_pg_logic52_or0;
  assign f_u_dadda_cla32_u_cla62_and266 = f_u_dadda_cla32_u_cla62_pg_logic52_and0 & f_u_dadda_cla32_u_cla62_pg_logic54_or0;
  assign f_u_dadda_cla32_u_cla62_and267 = f_u_dadda_cla32_u_cla62_pg_logic55_or0 & f_u_dadda_cla32_u_cla62_pg_logic53_or0;
  assign f_u_dadda_cla32_u_cla62_and268 = f_u_dadda_cla32_u_cla62_and266 & f_u_dadda_cla32_u_cla62_and267;
  assign f_u_dadda_cla32_u_cla62_and269 = f_u_dadda_cla32_u_cla62_pg_logic53_and0 & f_u_dadda_cla32_u_cla62_pg_logic55_or0;
  assign f_u_dadda_cla32_u_cla62_and270 = f_u_dadda_cla32_u_cla62_and269 & f_u_dadda_cla32_u_cla62_pg_logic54_or0;
  assign f_u_dadda_cla32_u_cla62_and271 = f_u_dadda_cla32_u_cla62_pg_logic54_and0 & f_u_dadda_cla32_u_cla62_pg_logic55_or0;
  assign f_u_dadda_cla32_u_cla62_or132 = f_u_dadda_cla32_u_cla62_and265 | f_u_dadda_cla32_u_cla62_and270;
  assign f_u_dadda_cla32_u_cla62_or133 = f_u_dadda_cla32_u_cla62_and268 | f_u_dadda_cla32_u_cla62_and271;
  assign f_u_dadda_cla32_u_cla62_or134 = f_u_dadda_cla32_u_cla62_or132 | f_u_dadda_cla32_u_cla62_or133;
  assign f_u_dadda_cla32_u_cla62_or135 = f_u_dadda_cla32_u_cla62_pg_logic55_and0 | f_u_dadda_cla32_u_cla62_or134;
  assign f_u_dadda_cla32_u_cla62_pg_logic56_or0 = f_u_dadda_cla32_fa836_xor1 | f_u_dadda_cla32_fa894_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic56_and0 = f_u_dadda_cla32_fa836_xor1 & f_u_dadda_cla32_fa894_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic56_xor0 = f_u_dadda_cla32_fa836_xor1 ^ f_u_dadda_cla32_fa894_xor1;
  assign f_u_dadda_cla32_u_cla62_xor56 = f_u_dadda_cla32_u_cla62_pg_logic56_xor0 ^ f_u_dadda_cla32_u_cla62_or135;
  assign f_u_dadda_cla32_u_cla62_and272 = f_u_dadda_cla32_u_cla62_or135 & f_u_dadda_cla32_u_cla62_pg_logic56_or0;
  assign f_u_dadda_cla32_u_cla62_or136 = f_u_dadda_cla32_u_cla62_pg_logic56_and0 | f_u_dadda_cla32_u_cla62_and272;
  assign f_u_dadda_cla32_u_cla62_pg_logic57_or0 = f_u_dadda_cla32_fa837_xor1 | f_u_dadda_cla32_fa895_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic57_and0 = f_u_dadda_cla32_fa837_xor1 & f_u_dadda_cla32_fa895_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic57_xor0 = f_u_dadda_cla32_fa837_xor1 ^ f_u_dadda_cla32_fa895_xor1;
  assign f_u_dadda_cla32_u_cla62_xor57 = f_u_dadda_cla32_u_cla62_pg_logic57_xor0 ^ f_u_dadda_cla32_u_cla62_or136;
  assign f_u_dadda_cla32_u_cla62_and273 = f_u_dadda_cla32_u_cla62_or135 & f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  assign f_u_dadda_cla32_u_cla62_and274 = f_u_dadda_cla32_u_cla62_and273 & f_u_dadda_cla32_u_cla62_pg_logic56_or0;
  assign f_u_dadda_cla32_u_cla62_and275 = f_u_dadda_cla32_u_cla62_pg_logic56_and0 & f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  assign f_u_dadda_cla32_u_cla62_or137 = f_u_dadda_cla32_u_cla62_and274 | f_u_dadda_cla32_u_cla62_and275;
  assign f_u_dadda_cla32_u_cla62_or138 = f_u_dadda_cla32_u_cla62_pg_logic57_and0 | f_u_dadda_cla32_u_cla62_or137;
  assign f_u_dadda_cla32_u_cla62_pg_logic58_or0 = f_u_dadda_cla32_fa838_xor1 | f_u_dadda_cla32_fa896_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic58_and0 = f_u_dadda_cla32_fa838_xor1 & f_u_dadda_cla32_fa896_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic58_xor0 = f_u_dadda_cla32_fa838_xor1 ^ f_u_dadda_cla32_fa896_xor1;
  assign f_u_dadda_cla32_u_cla62_xor58 = f_u_dadda_cla32_u_cla62_pg_logic58_xor0 ^ f_u_dadda_cla32_u_cla62_or138;
  assign f_u_dadda_cla32_u_cla62_and276 = f_u_dadda_cla32_u_cla62_or135 & f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  assign f_u_dadda_cla32_u_cla62_and277 = f_u_dadda_cla32_u_cla62_pg_logic58_or0 & f_u_dadda_cla32_u_cla62_pg_logic56_or0;
  assign f_u_dadda_cla32_u_cla62_and278 = f_u_dadda_cla32_u_cla62_and276 & f_u_dadda_cla32_u_cla62_and277;
  assign f_u_dadda_cla32_u_cla62_and279 = f_u_dadda_cla32_u_cla62_pg_logic56_and0 & f_u_dadda_cla32_u_cla62_pg_logic58_or0;
  assign f_u_dadda_cla32_u_cla62_and280 = f_u_dadda_cla32_u_cla62_and279 & f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  assign f_u_dadda_cla32_u_cla62_and281 = f_u_dadda_cla32_u_cla62_pg_logic57_and0 & f_u_dadda_cla32_u_cla62_pg_logic58_or0;
  assign f_u_dadda_cla32_u_cla62_or139 = f_u_dadda_cla32_u_cla62_and278 | f_u_dadda_cla32_u_cla62_and280;
  assign f_u_dadda_cla32_u_cla62_or140 = f_u_dadda_cla32_u_cla62_or139 | f_u_dadda_cla32_u_cla62_and281;
  assign f_u_dadda_cla32_u_cla62_or141 = f_u_dadda_cla32_u_cla62_pg_logic58_and0 | f_u_dadda_cla32_u_cla62_or140;
  assign f_u_dadda_cla32_u_cla62_pg_logic59_or0 = f_u_dadda_cla32_fa839_xor1 | f_u_dadda_cla32_fa897_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic59_and0 = f_u_dadda_cla32_fa839_xor1 & f_u_dadda_cla32_fa897_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic59_xor0 = f_u_dadda_cla32_fa839_xor1 ^ f_u_dadda_cla32_fa897_xor1;
  assign f_u_dadda_cla32_u_cla62_xor59 = f_u_dadda_cla32_u_cla62_pg_logic59_xor0 ^ f_u_dadda_cla32_u_cla62_or141;
  assign f_u_dadda_cla32_u_cla62_and282 = f_u_dadda_cla32_u_cla62_or135 & f_u_dadda_cla32_u_cla62_pg_logic58_or0;
  assign f_u_dadda_cla32_u_cla62_and283 = f_u_dadda_cla32_u_cla62_pg_logic59_or0 & f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  assign f_u_dadda_cla32_u_cla62_and284 = f_u_dadda_cla32_u_cla62_and282 & f_u_dadda_cla32_u_cla62_and283;
  assign f_u_dadda_cla32_u_cla62_and285 = f_u_dadda_cla32_u_cla62_and284 & f_u_dadda_cla32_u_cla62_pg_logic56_or0;
  assign f_u_dadda_cla32_u_cla62_and286 = f_u_dadda_cla32_u_cla62_pg_logic56_and0 & f_u_dadda_cla32_u_cla62_pg_logic58_or0;
  assign f_u_dadda_cla32_u_cla62_and287 = f_u_dadda_cla32_u_cla62_pg_logic59_or0 & f_u_dadda_cla32_u_cla62_pg_logic57_or0;
  assign f_u_dadda_cla32_u_cla62_and288 = f_u_dadda_cla32_u_cla62_and286 & f_u_dadda_cla32_u_cla62_and287;
  assign f_u_dadda_cla32_u_cla62_and289 = f_u_dadda_cla32_u_cla62_pg_logic57_and0 & f_u_dadda_cla32_u_cla62_pg_logic59_or0;
  assign f_u_dadda_cla32_u_cla62_and290 = f_u_dadda_cla32_u_cla62_and289 & f_u_dadda_cla32_u_cla62_pg_logic58_or0;
  assign f_u_dadda_cla32_u_cla62_and291 = f_u_dadda_cla32_u_cla62_pg_logic58_and0 & f_u_dadda_cla32_u_cla62_pg_logic59_or0;
  assign f_u_dadda_cla32_u_cla62_or142 = f_u_dadda_cla32_u_cla62_and285 | f_u_dadda_cla32_u_cla62_and290;
  assign f_u_dadda_cla32_u_cla62_or143 = f_u_dadda_cla32_u_cla62_and288 | f_u_dadda_cla32_u_cla62_and291;
  assign f_u_dadda_cla32_u_cla62_or144 = f_u_dadda_cla32_u_cla62_or142 | f_u_dadda_cla32_u_cla62_or143;
  assign f_u_dadda_cla32_u_cla62_or145 = f_u_dadda_cla32_u_cla62_pg_logic59_and0 | f_u_dadda_cla32_u_cla62_or144;
  assign f_u_dadda_cla32_u_cla62_pg_logic60_or0 = f_u_dadda_cla32_and_30_31 | f_u_dadda_cla32_fa898_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic60_and0 = f_u_dadda_cla32_and_30_31 & f_u_dadda_cla32_fa898_xor1;
  assign f_u_dadda_cla32_u_cla62_pg_logic60_xor0 = f_u_dadda_cla32_and_30_31 ^ f_u_dadda_cla32_fa898_xor1;
  assign f_u_dadda_cla32_u_cla62_xor60 = f_u_dadda_cla32_u_cla62_pg_logic60_xor0 ^ f_u_dadda_cla32_u_cla62_or145;
  assign f_u_dadda_cla32_u_cla62_and292 = f_u_dadda_cla32_u_cla62_or145 & f_u_dadda_cla32_u_cla62_pg_logic60_or0;
  assign f_u_dadda_cla32_u_cla62_or146 = f_u_dadda_cla32_u_cla62_pg_logic60_and0 | f_u_dadda_cla32_u_cla62_and292;
  assign f_u_dadda_cla32_u_cla62_pg_logic61_or0 = f_u_dadda_cla32_fa898_or0 | f_u_dadda_cla32_and_31_31;
  assign f_u_dadda_cla32_u_cla62_pg_logic61_and0 = f_u_dadda_cla32_fa898_or0 & f_u_dadda_cla32_and_31_31;
  assign f_u_dadda_cla32_u_cla62_pg_logic61_xor0 = f_u_dadda_cla32_fa898_or0 ^ f_u_dadda_cla32_and_31_31;
  assign f_u_dadda_cla32_u_cla62_xor61 = f_u_dadda_cla32_u_cla62_pg_logic61_xor0 ^ f_u_dadda_cla32_u_cla62_or146;
  assign f_u_dadda_cla32_u_cla62_and293 = f_u_dadda_cla32_u_cla62_or145 & f_u_dadda_cla32_u_cla62_pg_logic61_or0;
  assign f_u_dadda_cla32_u_cla62_and294 = f_u_dadda_cla32_u_cla62_and293 & f_u_dadda_cla32_u_cla62_pg_logic60_or0;
  assign f_u_dadda_cla32_u_cla62_and295 = f_u_dadda_cla32_u_cla62_pg_logic60_and0 & f_u_dadda_cla32_u_cla62_pg_logic61_or0;
  assign f_u_dadda_cla32_u_cla62_or147 = f_u_dadda_cla32_u_cla62_and294 | f_u_dadda_cla32_u_cla62_and295;
  assign f_u_dadda_cla32_u_cla62_or148 = f_u_dadda_cla32_u_cla62_pg_logic61_and0 | f_u_dadda_cla32_u_cla62_or147;

  assign f_u_dadda_cla32_out[0] = f_u_dadda_cla32_and_0_0;
  assign f_u_dadda_cla32_out[1] = f_u_dadda_cla32_u_cla62_pg_logic0_xor0;
  assign f_u_dadda_cla32_out[2] = f_u_dadda_cla32_u_cla62_xor1;
  assign f_u_dadda_cla32_out[3] = f_u_dadda_cla32_u_cla62_xor2;
  assign f_u_dadda_cla32_out[4] = f_u_dadda_cla32_u_cla62_xor3;
  assign f_u_dadda_cla32_out[5] = f_u_dadda_cla32_u_cla62_xor4;
  assign f_u_dadda_cla32_out[6] = f_u_dadda_cla32_u_cla62_xor5;
  assign f_u_dadda_cla32_out[7] = f_u_dadda_cla32_u_cla62_xor6;
  assign f_u_dadda_cla32_out[8] = f_u_dadda_cla32_u_cla62_xor7;
  assign f_u_dadda_cla32_out[9] = f_u_dadda_cla32_u_cla62_xor8;
  assign f_u_dadda_cla32_out[10] = f_u_dadda_cla32_u_cla62_xor9;
  assign f_u_dadda_cla32_out[11] = f_u_dadda_cla32_u_cla62_xor10;
  assign f_u_dadda_cla32_out[12] = f_u_dadda_cla32_u_cla62_xor11;
  assign f_u_dadda_cla32_out[13] = f_u_dadda_cla32_u_cla62_xor12;
  assign f_u_dadda_cla32_out[14] = f_u_dadda_cla32_u_cla62_xor13;
  assign f_u_dadda_cla32_out[15] = f_u_dadda_cla32_u_cla62_xor14;
  assign f_u_dadda_cla32_out[16] = f_u_dadda_cla32_u_cla62_xor15;
  assign f_u_dadda_cla32_out[17] = f_u_dadda_cla32_u_cla62_xor16;
  assign f_u_dadda_cla32_out[18] = f_u_dadda_cla32_u_cla62_xor17;
  assign f_u_dadda_cla32_out[19] = f_u_dadda_cla32_u_cla62_xor18;
  assign f_u_dadda_cla32_out[20] = f_u_dadda_cla32_u_cla62_xor19;
  assign f_u_dadda_cla32_out[21] = f_u_dadda_cla32_u_cla62_xor20;
  assign f_u_dadda_cla32_out[22] = f_u_dadda_cla32_u_cla62_xor21;
  assign f_u_dadda_cla32_out[23] = f_u_dadda_cla32_u_cla62_xor22;
  assign f_u_dadda_cla32_out[24] = f_u_dadda_cla32_u_cla62_xor23;
  assign f_u_dadda_cla32_out[25] = f_u_dadda_cla32_u_cla62_xor24;
  assign f_u_dadda_cla32_out[26] = f_u_dadda_cla32_u_cla62_xor25;
  assign f_u_dadda_cla32_out[27] = f_u_dadda_cla32_u_cla62_xor26;
  assign f_u_dadda_cla32_out[28] = f_u_dadda_cla32_u_cla62_xor27;
  assign f_u_dadda_cla32_out[29] = f_u_dadda_cla32_u_cla62_xor28;
  assign f_u_dadda_cla32_out[30] = f_u_dadda_cla32_u_cla62_xor29;
  assign f_u_dadda_cla32_out[31] = f_u_dadda_cla32_u_cla62_xor30;
  assign f_u_dadda_cla32_out[32] = f_u_dadda_cla32_u_cla62_xor31;
  assign f_u_dadda_cla32_out[33] = f_u_dadda_cla32_u_cla62_xor32;
  assign f_u_dadda_cla32_out[34] = f_u_dadda_cla32_u_cla62_xor33;
  assign f_u_dadda_cla32_out[35] = f_u_dadda_cla32_u_cla62_xor34;
  assign f_u_dadda_cla32_out[36] = f_u_dadda_cla32_u_cla62_xor35;
  assign f_u_dadda_cla32_out[37] = f_u_dadda_cla32_u_cla62_xor36;
  assign f_u_dadda_cla32_out[38] = f_u_dadda_cla32_u_cla62_xor37;
  assign f_u_dadda_cla32_out[39] = f_u_dadda_cla32_u_cla62_xor38;
  assign f_u_dadda_cla32_out[40] = f_u_dadda_cla32_u_cla62_xor39;
  assign f_u_dadda_cla32_out[41] = f_u_dadda_cla32_u_cla62_xor40;
  assign f_u_dadda_cla32_out[42] = f_u_dadda_cla32_u_cla62_xor41;
  assign f_u_dadda_cla32_out[43] = f_u_dadda_cla32_u_cla62_xor42;
  assign f_u_dadda_cla32_out[44] = f_u_dadda_cla32_u_cla62_xor43;
  assign f_u_dadda_cla32_out[45] = f_u_dadda_cla32_u_cla62_xor44;
  assign f_u_dadda_cla32_out[46] = f_u_dadda_cla32_u_cla62_xor45;
  assign f_u_dadda_cla32_out[47] = f_u_dadda_cla32_u_cla62_xor46;
  assign f_u_dadda_cla32_out[48] = f_u_dadda_cla32_u_cla62_xor47;
  assign f_u_dadda_cla32_out[49] = f_u_dadda_cla32_u_cla62_xor48;
  assign f_u_dadda_cla32_out[50] = f_u_dadda_cla32_u_cla62_xor49;
  assign f_u_dadda_cla32_out[51] = f_u_dadda_cla32_u_cla62_xor50;
  assign f_u_dadda_cla32_out[52] = f_u_dadda_cla32_u_cla62_xor51;
  assign f_u_dadda_cla32_out[53] = f_u_dadda_cla32_u_cla62_xor52;
  assign f_u_dadda_cla32_out[54] = f_u_dadda_cla32_u_cla62_xor53;
  assign f_u_dadda_cla32_out[55] = f_u_dadda_cla32_u_cla62_xor54;
  assign f_u_dadda_cla32_out[56] = f_u_dadda_cla32_u_cla62_xor55;
  assign f_u_dadda_cla32_out[57] = f_u_dadda_cla32_u_cla62_xor56;
  assign f_u_dadda_cla32_out[58] = f_u_dadda_cla32_u_cla62_xor57;
  assign f_u_dadda_cla32_out[59] = f_u_dadda_cla32_u_cla62_xor58;
  assign f_u_dadda_cla32_out[60] = f_u_dadda_cla32_u_cla62_xor59;
  assign f_u_dadda_cla32_out[61] = f_u_dadda_cla32_u_cla62_xor60;
  assign f_u_dadda_cla32_out[62] = f_u_dadda_cla32_u_cla62_xor61;
  assign f_u_dadda_cla32_out[63] = f_u_dadda_cla32_u_cla62_or148;
endmodule