module u_rca12(input [11:0] a, input [11:0] b, output [12:0] u_rca12_out);
  wire u_rca12_ha_xor0;
  wire u_rca12_ha_and0;
  wire u_rca12_fa1_xor0;
  wire u_rca12_fa1_and0;
  wire u_rca12_fa1_xor1;
  wire u_rca12_fa1_and1;
  wire u_rca12_fa1_or0;
  wire u_rca12_fa2_xor0;
  wire u_rca12_fa2_and0;
  wire u_rca12_fa2_xor1;
  wire u_rca12_fa2_and1;
  wire u_rca12_fa2_or0;
  wire u_rca12_fa3_xor0;
  wire u_rca12_fa3_and0;
  wire u_rca12_fa3_xor1;
  wire u_rca12_fa3_and1;
  wire u_rca12_fa3_or0;
  wire u_rca12_fa4_xor0;
  wire u_rca12_fa4_and0;
  wire u_rca12_fa4_xor1;
  wire u_rca12_fa4_and1;
  wire u_rca12_fa4_or0;
  wire u_rca12_fa5_xor0;
  wire u_rca12_fa5_and0;
  wire u_rca12_fa5_xor1;
  wire u_rca12_fa5_and1;
  wire u_rca12_fa5_or0;
  wire u_rca12_fa6_xor0;
  wire u_rca12_fa6_and0;
  wire u_rca12_fa6_xor1;
  wire u_rca12_fa6_and1;
  wire u_rca12_fa6_or0;
  wire u_rca12_fa7_xor0;
  wire u_rca12_fa7_and0;
  wire u_rca12_fa7_xor1;
  wire u_rca12_fa7_and1;
  wire u_rca12_fa7_or0;
  wire u_rca12_fa8_xor0;
  wire u_rca12_fa8_and0;
  wire u_rca12_fa8_xor1;
  wire u_rca12_fa8_and1;
  wire u_rca12_fa8_or0;
  wire u_rca12_fa9_xor0;
  wire u_rca12_fa9_and0;
  wire u_rca12_fa9_xor1;
  wire u_rca12_fa9_and1;
  wire u_rca12_fa9_or0;
  wire u_rca12_fa10_xor0;
  wire u_rca12_fa10_and0;
  wire u_rca12_fa10_xor1;
  wire u_rca12_fa10_and1;
  wire u_rca12_fa10_or0;
  wire u_rca12_fa11_xor0;
  wire u_rca12_fa11_and0;
  wire u_rca12_fa11_xor1;
  wire u_rca12_fa11_and1;
  wire u_rca12_fa11_or0;

  assign u_rca12_ha_xor0 = a[0] ^ b[0];
  assign u_rca12_ha_and0 = a[0] & b[0];
  assign u_rca12_fa1_xor0 = a[1] ^ b[1];
  assign u_rca12_fa1_and0 = a[1] & b[1];
  assign u_rca12_fa1_xor1 = u_rca12_fa1_xor0 ^ u_rca12_ha_and0;
  assign u_rca12_fa1_and1 = u_rca12_fa1_xor0 & u_rca12_ha_and0;
  assign u_rca12_fa1_or0 = u_rca12_fa1_and0 | u_rca12_fa1_and1;
  assign u_rca12_fa2_xor0 = a[2] ^ b[2];
  assign u_rca12_fa2_and0 = a[2] & b[2];
  assign u_rca12_fa2_xor1 = u_rca12_fa2_xor0 ^ u_rca12_fa1_or0;
  assign u_rca12_fa2_and1 = u_rca12_fa2_xor0 & u_rca12_fa1_or0;
  assign u_rca12_fa2_or0 = u_rca12_fa2_and0 | u_rca12_fa2_and1;
  assign u_rca12_fa3_xor0 = a[3] ^ b[3];
  assign u_rca12_fa3_and0 = a[3] & b[3];
  assign u_rca12_fa3_xor1 = u_rca12_fa3_xor0 ^ u_rca12_fa2_or0;
  assign u_rca12_fa3_and1 = u_rca12_fa3_xor0 & u_rca12_fa2_or0;
  assign u_rca12_fa3_or0 = u_rca12_fa3_and0 | u_rca12_fa3_and1;
  assign u_rca12_fa4_xor0 = a[4] ^ b[4];
  assign u_rca12_fa4_and0 = a[4] & b[4];
  assign u_rca12_fa4_xor1 = u_rca12_fa4_xor0 ^ u_rca12_fa3_or0;
  assign u_rca12_fa4_and1 = u_rca12_fa4_xor0 & u_rca12_fa3_or0;
  assign u_rca12_fa4_or0 = u_rca12_fa4_and0 | u_rca12_fa4_and1;
  assign u_rca12_fa5_xor0 = a[5] ^ b[5];
  assign u_rca12_fa5_and0 = a[5] & b[5];
  assign u_rca12_fa5_xor1 = u_rca12_fa5_xor0 ^ u_rca12_fa4_or0;
  assign u_rca12_fa5_and1 = u_rca12_fa5_xor0 & u_rca12_fa4_or0;
  assign u_rca12_fa5_or0 = u_rca12_fa5_and0 | u_rca12_fa5_and1;
  assign u_rca12_fa6_xor0 = a[6] ^ b[6];
  assign u_rca12_fa6_and0 = a[6] & b[6];
  assign u_rca12_fa6_xor1 = u_rca12_fa6_xor0 ^ u_rca12_fa5_or0;
  assign u_rca12_fa6_and1 = u_rca12_fa6_xor0 & u_rca12_fa5_or0;
  assign u_rca12_fa6_or0 = u_rca12_fa6_and0 | u_rca12_fa6_and1;
  assign u_rca12_fa7_xor0 = a[7] ^ b[7];
  assign u_rca12_fa7_and0 = a[7] & b[7];
  assign u_rca12_fa7_xor1 = u_rca12_fa7_xor0 ^ u_rca12_fa6_or0;
  assign u_rca12_fa7_and1 = u_rca12_fa7_xor0 & u_rca12_fa6_or0;
  assign u_rca12_fa7_or0 = u_rca12_fa7_and0 | u_rca12_fa7_and1;
  assign u_rca12_fa8_xor0 = a[8] ^ b[8];
  assign u_rca12_fa8_and0 = a[8] & b[8];
  assign u_rca12_fa8_xor1 = u_rca12_fa8_xor0 ^ u_rca12_fa7_or0;
  assign u_rca12_fa8_and1 = u_rca12_fa8_xor0 & u_rca12_fa7_or0;
  assign u_rca12_fa8_or0 = u_rca12_fa8_and0 | u_rca12_fa8_and1;
  assign u_rca12_fa9_xor0 = a[9] ^ b[9];
  assign u_rca12_fa9_and0 = a[9] & b[9];
  assign u_rca12_fa9_xor1 = u_rca12_fa9_xor0 ^ u_rca12_fa8_or0;
  assign u_rca12_fa9_and1 = u_rca12_fa9_xor0 & u_rca12_fa8_or0;
  assign u_rca12_fa9_or0 = u_rca12_fa9_and0 | u_rca12_fa9_and1;
  assign u_rca12_fa10_xor0 = a[10] ^ b[10];
  assign u_rca12_fa10_and0 = a[10] & b[10];
  assign u_rca12_fa10_xor1 = u_rca12_fa10_xor0 ^ u_rca12_fa9_or0;
  assign u_rca12_fa10_and1 = u_rca12_fa10_xor0 & u_rca12_fa9_or0;
  assign u_rca12_fa10_or0 = u_rca12_fa10_and0 | u_rca12_fa10_and1;
  assign u_rca12_fa11_xor0 = a[11] ^ b[11];
  assign u_rca12_fa11_and0 = a[11] & b[11];
  assign u_rca12_fa11_xor1 = u_rca12_fa11_xor0 ^ u_rca12_fa10_or0;
  assign u_rca12_fa11_and1 = u_rca12_fa11_xor0 & u_rca12_fa10_or0;
  assign u_rca12_fa11_or0 = u_rca12_fa11_and0 | u_rca12_fa11_and1;

  assign u_rca12_out[0] = u_rca12_ha_xor0;
  assign u_rca12_out[1] = u_rca12_fa1_xor1;
  assign u_rca12_out[2] = u_rca12_fa2_xor1;
  assign u_rca12_out[3] = u_rca12_fa3_xor1;
  assign u_rca12_out[4] = u_rca12_fa4_xor1;
  assign u_rca12_out[5] = u_rca12_fa5_xor1;
  assign u_rca12_out[6] = u_rca12_fa6_xor1;
  assign u_rca12_out[7] = u_rca12_fa7_xor1;
  assign u_rca12_out[8] = u_rca12_fa8_xor1;
  assign u_rca12_out[9] = u_rca12_fa9_xor1;
  assign u_rca12_out[10] = u_rca12_fa10_xor1;
  assign u_rca12_out[11] = u_rca12_fa11_xor1;
  assign u_rca12_out[12] = u_rca12_fa11_or0;
endmodule