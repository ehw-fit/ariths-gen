module f_arrdiv32(input [31:0] a, input [31:0] b, output [31:0] f_arrdiv32_out);
  wire f_arrdiv32_fs0_xor0;
  wire f_arrdiv32_fs0_not0;
  wire f_arrdiv32_fs0_and0;
  wire f_arrdiv32_fs0_not1;
  wire f_arrdiv32_fs1_xor1;
  wire f_arrdiv32_fs1_not1;
  wire f_arrdiv32_fs1_and1;
  wire f_arrdiv32_fs1_or0;
  wire f_arrdiv32_fs2_xor1;
  wire f_arrdiv32_fs2_not1;
  wire f_arrdiv32_fs2_and1;
  wire f_arrdiv32_fs2_or0;
  wire f_arrdiv32_fs3_xor1;
  wire f_arrdiv32_fs3_not1;
  wire f_arrdiv32_fs3_and1;
  wire f_arrdiv32_fs3_or0;
  wire f_arrdiv32_fs4_xor1;
  wire f_arrdiv32_fs4_not1;
  wire f_arrdiv32_fs4_and1;
  wire f_arrdiv32_fs4_or0;
  wire f_arrdiv32_fs5_xor1;
  wire f_arrdiv32_fs5_not1;
  wire f_arrdiv32_fs5_and1;
  wire f_arrdiv32_fs5_or0;
  wire f_arrdiv32_fs6_xor1;
  wire f_arrdiv32_fs6_not1;
  wire f_arrdiv32_fs6_and1;
  wire f_arrdiv32_fs6_or0;
  wire f_arrdiv32_fs7_xor1;
  wire f_arrdiv32_fs7_not1;
  wire f_arrdiv32_fs7_and1;
  wire f_arrdiv32_fs7_or0;
  wire f_arrdiv32_fs8_xor1;
  wire f_arrdiv32_fs8_not1;
  wire f_arrdiv32_fs8_and1;
  wire f_arrdiv32_fs8_or0;
  wire f_arrdiv32_fs9_xor1;
  wire f_arrdiv32_fs9_not1;
  wire f_arrdiv32_fs9_and1;
  wire f_arrdiv32_fs9_or0;
  wire f_arrdiv32_fs10_xor1;
  wire f_arrdiv32_fs10_not1;
  wire f_arrdiv32_fs10_and1;
  wire f_arrdiv32_fs10_or0;
  wire f_arrdiv32_fs11_xor1;
  wire f_arrdiv32_fs11_not1;
  wire f_arrdiv32_fs11_and1;
  wire f_arrdiv32_fs11_or0;
  wire f_arrdiv32_fs12_xor1;
  wire f_arrdiv32_fs12_not1;
  wire f_arrdiv32_fs12_and1;
  wire f_arrdiv32_fs12_or0;
  wire f_arrdiv32_fs13_xor1;
  wire f_arrdiv32_fs13_not1;
  wire f_arrdiv32_fs13_and1;
  wire f_arrdiv32_fs13_or0;
  wire f_arrdiv32_fs14_xor1;
  wire f_arrdiv32_fs14_not1;
  wire f_arrdiv32_fs14_and1;
  wire f_arrdiv32_fs14_or0;
  wire f_arrdiv32_fs15_xor1;
  wire f_arrdiv32_fs15_not1;
  wire f_arrdiv32_fs15_and1;
  wire f_arrdiv32_fs15_or0;
  wire f_arrdiv32_fs16_xor1;
  wire f_arrdiv32_fs16_not1;
  wire f_arrdiv32_fs16_and1;
  wire f_arrdiv32_fs16_or0;
  wire f_arrdiv32_fs17_xor1;
  wire f_arrdiv32_fs17_not1;
  wire f_arrdiv32_fs17_and1;
  wire f_arrdiv32_fs17_or0;
  wire f_arrdiv32_fs18_xor1;
  wire f_arrdiv32_fs18_not1;
  wire f_arrdiv32_fs18_and1;
  wire f_arrdiv32_fs18_or0;
  wire f_arrdiv32_fs19_xor1;
  wire f_arrdiv32_fs19_not1;
  wire f_arrdiv32_fs19_and1;
  wire f_arrdiv32_fs19_or0;
  wire f_arrdiv32_fs20_xor1;
  wire f_arrdiv32_fs20_not1;
  wire f_arrdiv32_fs20_and1;
  wire f_arrdiv32_fs20_or0;
  wire f_arrdiv32_fs21_xor1;
  wire f_arrdiv32_fs21_not1;
  wire f_arrdiv32_fs21_and1;
  wire f_arrdiv32_fs21_or0;
  wire f_arrdiv32_fs22_xor1;
  wire f_arrdiv32_fs22_not1;
  wire f_arrdiv32_fs22_and1;
  wire f_arrdiv32_fs22_or0;
  wire f_arrdiv32_fs23_xor1;
  wire f_arrdiv32_fs23_not1;
  wire f_arrdiv32_fs23_and1;
  wire f_arrdiv32_fs23_or0;
  wire f_arrdiv32_fs24_xor1;
  wire f_arrdiv32_fs24_not1;
  wire f_arrdiv32_fs24_and1;
  wire f_arrdiv32_fs24_or0;
  wire f_arrdiv32_fs25_xor1;
  wire f_arrdiv32_fs25_not1;
  wire f_arrdiv32_fs25_and1;
  wire f_arrdiv32_fs25_or0;
  wire f_arrdiv32_fs26_xor1;
  wire f_arrdiv32_fs26_not1;
  wire f_arrdiv32_fs26_and1;
  wire f_arrdiv32_fs26_or0;
  wire f_arrdiv32_fs27_xor1;
  wire f_arrdiv32_fs27_not1;
  wire f_arrdiv32_fs27_and1;
  wire f_arrdiv32_fs27_or0;
  wire f_arrdiv32_fs28_xor1;
  wire f_arrdiv32_fs28_not1;
  wire f_arrdiv32_fs28_and1;
  wire f_arrdiv32_fs28_or0;
  wire f_arrdiv32_fs29_xor1;
  wire f_arrdiv32_fs29_not1;
  wire f_arrdiv32_fs29_and1;
  wire f_arrdiv32_fs29_or0;
  wire f_arrdiv32_fs30_xor1;
  wire f_arrdiv32_fs30_not1;
  wire f_arrdiv32_fs30_and1;
  wire f_arrdiv32_fs30_or0;
  wire f_arrdiv32_fs31_xor1;
  wire f_arrdiv32_fs31_not1;
  wire f_arrdiv32_fs31_and1;
  wire f_arrdiv32_fs31_or0;
  wire f_arrdiv32_mux2to10_and0;
  wire f_arrdiv32_mux2to10_not0;
  wire f_arrdiv32_mux2to10_and1;
  wire f_arrdiv32_mux2to10_xor0;
  wire f_arrdiv32_mux2to11_not0;
  wire f_arrdiv32_mux2to11_and1;
  wire f_arrdiv32_mux2to12_not0;
  wire f_arrdiv32_mux2to12_and1;
  wire f_arrdiv32_mux2to13_not0;
  wire f_arrdiv32_mux2to13_and1;
  wire f_arrdiv32_mux2to14_not0;
  wire f_arrdiv32_mux2to14_and1;
  wire f_arrdiv32_mux2to15_not0;
  wire f_arrdiv32_mux2to15_and1;
  wire f_arrdiv32_mux2to16_not0;
  wire f_arrdiv32_mux2to16_and1;
  wire f_arrdiv32_mux2to17_not0;
  wire f_arrdiv32_mux2to17_and1;
  wire f_arrdiv32_mux2to18_not0;
  wire f_arrdiv32_mux2to18_and1;
  wire f_arrdiv32_mux2to19_not0;
  wire f_arrdiv32_mux2to19_and1;
  wire f_arrdiv32_mux2to110_not0;
  wire f_arrdiv32_mux2to110_and1;
  wire f_arrdiv32_mux2to111_not0;
  wire f_arrdiv32_mux2to111_and1;
  wire f_arrdiv32_mux2to112_not0;
  wire f_arrdiv32_mux2to112_and1;
  wire f_arrdiv32_mux2to113_not0;
  wire f_arrdiv32_mux2to113_and1;
  wire f_arrdiv32_mux2to114_not0;
  wire f_arrdiv32_mux2to114_and1;
  wire f_arrdiv32_mux2to115_not0;
  wire f_arrdiv32_mux2to115_and1;
  wire f_arrdiv32_mux2to116_not0;
  wire f_arrdiv32_mux2to116_and1;
  wire f_arrdiv32_mux2to117_not0;
  wire f_arrdiv32_mux2to117_and1;
  wire f_arrdiv32_mux2to118_not0;
  wire f_arrdiv32_mux2to118_and1;
  wire f_arrdiv32_mux2to119_not0;
  wire f_arrdiv32_mux2to119_and1;
  wire f_arrdiv32_mux2to120_not0;
  wire f_arrdiv32_mux2to120_and1;
  wire f_arrdiv32_mux2to121_not0;
  wire f_arrdiv32_mux2to121_and1;
  wire f_arrdiv32_mux2to122_not0;
  wire f_arrdiv32_mux2to122_and1;
  wire f_arrdiv32_mux2to123_not0;
  wire f_arrdiv32_mux2to123_and1;
  wire f_arrdiv32_mux2to124_not0;
  wire f_arrdiv32_mux2to124_and1;
  wire f_arrdiv32_mux2to125_not0;
  wire f_arrdiv32_mux2to125_and1;
  wire f_arrdiv32_mux2to126_not0;
  wire f_arrdiv32_mux2to126_and1;
  wire f_arrdiv32_mux2to127_not0;
  wire f_arrdiv32_mux2to127_and1;
  wire f_arrdiv32_mux2to128_not0;
  wire f_arrdiv32_mux2to128_and1;
  wire f_arrdiv32_mux2to129_not0;
  wire f_arrdiv32_mux2to129_and1;
  wire f_arrdiv32_mux2to130_not0;
  wire f_arrdiv32_mux2to130_and1;
  wire f_arrdiv32_not0;
  wire f_arrdiv32_fs32_xor0;
  wire f_arrdiv32_fs32_not0;
  wire f_arrdiv32_fs32_and0;
  wire f_arrdiv32_fs32_not1;
  wire f_arrdiv32_fs33_xor0;
  wire f_arrdiv32_fs33_not0;
  wire f_arrdiv32_fs33_and0;
  wire f_arrdiv32_fs33_xor1;
  wire f_arrdiv32_fs33_not1;
  wire f_arrdiv32_fs33_and1;
  wire f_arrdiv32_fs33_or0;
  wire f_arrdiv32_fs34_xor0;
  wire f_arrdiv32_fs34_not0;
  wire f_arrdiv32_fs34_and0;
  wire f_arrdiv32_fs34_xor1;
  wire f_arrdiv32_fs34_not1;
  wire f_arrdiv32_fs34_and1;
  wire f_arrdiv32_fs34_or0;
  wire f_arrdiv32_fs35_xor0;
  wire f_arrdiv32_fs35_not0;
  wire f_arrdiv32_fs35_and0;
  wire f_arrdiv32_fs35_xor1;
  wire f_arrdiv32_fs35_not1;
  wire f_arrdiv32_fs35_and1;
  wire f_arrdiv32_fs35_or0;
  wire f_arrdiv32_fs36_xor0;
  wire f_arrdiv32_fs36_not0;
  wire f_arrdiv32_fs36_and0;
  wire f_arrdiv32_fs36_xor1;
  wire f_arrdiv32_fs36_not1;
  wire f_arrdiv32_fs36_and1;
  wire f_arrdiv32_fs36_or0;
  wire f_arrdiv32_fs37_xor0;
  wire f_arrdiv32_fs37_not0;
  wire f_arrdiv32_fs37_and0;
  wire f_arrdiv32_fs37_xor1;
  wire f_arrdiv32_fs37_not1;
  wire f_arrdiv32_fs37_and1;
  wire f_arrdiv32_fs37_or0;
  wire f_arrdiv32_fs38_xor0;
  wire f_arrdiv32_fs38_not0;
  wire f_arrdiv32_fs38_and0;
  wire f_arrdiv32_fs38_xor1;
  wire f_arrdiv32_fs38_not1;
  wire f_arrdiv32_fs38_and1;
  wire f_arrdiv32_fs38_or0;
  wire f_arrdiv32_fs39_xor0;
  wire f_arrdiv32_fs39_not0;
  wire f_arrdiv32_fs39_and0;
  wire f_arrdiv32_fs39_xor1;
  wire f_arrdiv32_fs39_not1;
  wire f_arrdiv32_fs39_and1;
  wire f_arrdiv32_fs39_or0;
  wire f_arrdiv32_fs40_xor0;
  wire f_arrdiv32_fs40_not0;
  wire f_arrdiv32_fs40_and0;
  wire f_arrdiv32_fs40_xor1;
  wire f_arrdiv32_fs40_not1;
  wire f_arrdiv32_fs40_and1;
  wire f_arrdiv32_fs40_or0;
  wire f_arrdiv32_fs41_xor0;
  wire f_arrdiv32_fs41_not0;
  wire f_arrdiv32_fs41_and0;
  wire f_arrdiv32_fs41_xor1;
  wire f_arrdiv32_fs41_not1;
  wire f_arrdiv32_fs41_and1;
  wire f_arrdiv32_fs41_or0;
  wire f_arrdiv32_fs42_xor0;
  wire f_arrdiv32_fs42_not0;
  wire f_arrdiv32_fs42_and0;
  wire f_arrdiv32_fs42_xor1;
  wire f_arrdiv32_fs42_not1;
  wire f_arrdiv32_fs42_and1;
  wire f_arrdiv32_fs42_or0;
  wire f_arrdiv32_fs43_xor0;
  wire f_arrdiv32_fs43_not0;
  wire f_arrdiv32_fs43_and0;
  wire f_arrdiv32_fs43_xor1;
  wire f_arrdiv32_fs43_not1;
  wire f_arrdiv32_fs43_and1;
  wire f_arrdiv32_fs43_or0;
  wire f_arrdiv32_fs44_xor0;
  wire f_arrdiv32_fs44_not0;
  wire f_arrdiv32_fs44_and0;
  wire f_arrdiv32_fs44_xor1;
  wire f_arrdiv32_fs44_not1;
  wire f_arrdiv32_fs44_and1;
  wire f_arrdiv32_fs44_or0;
  wire f_arrdiv32_fs45_xor0;
  wire f_arrdiv32_fs45_not0;
  wire f_arrdiv32_fs45_and0;
  wire f_arrdiv32_fs45_xor1;
  wire f_arrdiv32_fs45_not1;
  wire f_arrdiv32_fs45_and1;
  wire f_arrdiv32_fs45_or0;
  wire f_arrdiv32_fs46_xor0;
  wire f_arrdiv32_fs46_not0;
  wire f_arrdiv32_fs46_and0;
  wire f_arrdiv32_fs46_xor1;
  wire f_arrdiv32_fs46_not1;
  wire f_arrdiv32_fs46_and1;
  wire f_arrdiv32_fs46_or0;
  wire f_arrdiv32_fs47_xor0;
  wire f_arrdiv32_fs47_not0;
  wire f_arrdiv32_fs47_and0;
  wire f_arrdiv32_fs47_xor1;
  wire f_arrdiv32_fs47_not1;
  wire f_arrdiv32_fs47_and1;
  wire f_arrdiv32_fs47_or0;
  wire f_arrdiv32_fs48_xor0;
  wire f_arrdiv32_fs48_not0;
  wire f_arrdiv32_fs48_and0;
  wire f_arrdiv32_fs48_xor1;
  wire f_arrdiv32_fs48_not1;
  wire f_arrdiv32_fs48_and1;
  wire f_arrdiv32_fs48_or0;
  wire f_arrdiv32_fs49_xor0;
  wire f_arrdiv32_fs49_not0;
  wire f_arrdiv32_fs49_and0;
  wire f_arrdiv32_fs49_xor1;
  wire f_arrdiv32_fs49_not1;
  wire f_arrdiv32_fs49_and1;
  wire f_arrdiv32_fs49_or0;
  wire f_arrdiv32_fs50_xor0;
  wire f_arrdiv32_fs50_not0;
  wire f_arrdiv32_fs50_and0;
  wire f_arrdiv32_fs50_xor1;
  wire f_arrdiv32_fs50_not1;
  wire f_arrdiv32_fs50_and1;
  wire f_arrdiv32_fs50_or0;
  wire f_arrdiv32_fs51_xor0;
  wire f_arrdiv32_fs51_not0;
  wire f_arrdiv32_fs51_and0;
  wire f_arrdiv32_fs51_xor1;
  wire f_arrdiv32_fs51_not1;
  wire f_arrdiv32_fs51_and1;
  wire f_arrdiv32_fs51_or0;
  wire f_arrdiv32_fs52_xor0;
  wire f_arrdiv32_fs52_not0;
  wire f_arrdiv32_fs52_and0;
  wire f_arrdiv32_fs52_xor1;
  wire f_arrdiv32_fs52_not1;
  wire f_arrdiv32_fs52_and1;
  wire f_arrdiv32_fs52_or0;
  wire f_arrdiv32_fs53_xor0;
  wire f_arrdiv32_fs53_not0;
  wire f_arrdiv32_fs53_and0;
  wire f_arrdiv32_fs53_xor1;
  wire f_arrdiv32_fs53_not1;
  wire f_arrdiv32_fs53_and1;
  wire f_arrdiv32_fs53_or0;
  wire f_arrdiv32_fs54_xor0;
  wire f_arrdiv32_fs54_not0;
  wire f_arrdiv32_fs54_and0;
  wire f_arrdiv32_fs54_xor1;
  wire f_arrdiv32_fs54_not1;
  wire f_arrdiv32_fs54_and1;
  wire f_arrdiv32_fs54_or0;
  wire f_arrdiv32_fs55_xor0;
  wire f_arrdiv32_fs55_not0;
  wire f_arrdiv32_fs55_and0;
  wire f_arrdiv32_fs55_xor1;
  wire f_arrdiv32_fs55_not1;
  wire f_arrdiv32_fs55_and1;
  wire f_arrdiv32_fs55_or0;
  wire f_arrdiv32_fs56_xor0;
  wire f_arrdiv32_fs56_not0;
  wire f_arrdiv32_fs56_and0;
  wire f_arrdiv32_fs56_xor1;
  wire f_arrdiv32_fs56_not1;
  wire f_arrdiv32_fs56_and1;
  wire f_arrdiv32_fs56_or0;
  wire f_arrdiv32_fs57_xor0;
  wire f_arrdiv32_fs57_not0;
  wire f_arrdiv32_fs57_and0;
  wire f_arrdiv32_fs57_xor1;
  wire f_arrdiv32_fs57_not1;
  wire f_arrdiv32_fs57_and1;
  wire f_arrdiv32_fs57_or0;
  wire f_arrdiv32_fs58_xor0;
  wire f_arrdiv32_fs58_not0;
  wire f_arrdiv32_fs58_and0;
  wire f_arrdiv32_fs58_xor1;
  wire f_arrdiv32_fs58_not1;
  wire f_arrdiv32_fs58_and1;
  wire f_arrdiv32_fs58_or0;
  wire f_arrdiv32_fs59_xor0;
  wire f_arrdiv32_fs59_not0;
  wire f_arrdiv32_fs59_and0;
  wire f_arrdiv32_fs59_xor1;
  wire f_arrdiv32_fs59_not1;
  wire f_arrdiv32_fs59_and1;
  wire f_arrdiv32_fs59_or0;
  wire f_arrdiv32_fs60_xor0;
  wire f_arrdiv32_fs60_not0;
  wire f_arrdiv32_fs60_and0;
  wire f_arrdiv32_fs60_xor1;
  wire f_arrdiv32_fs60_not1;
  wire f_arrdiv32_fs60_and1;
  wire f_arrdiv32_fs60_or0;
  wire f_arrdiv32_fs61_xor0;
  wire f_arrdiv32_fs61_not0;
  wire f_arrdiv32_fs61_and0;
  wire f_arrdiv32_fs61_xor1;
  wire f_arrdiv32_fs61_not1;
  wire f_arrdiv32_fs61_and1;
  wire f_arrdiv32_fs61_or0;
  wire f_arrdiv32_fs62_xor0;
  wire f_arrdiv32_fs62_not0;
  wire f_arrdiv32_fs62_and0;
  wire f_arrdiv32_fs62_xor1;
  wire f_arrdiv32_fs62_not1;
  wire f_arrdiv32_fs62_and1;
  wire f_arrdiv32_fs62_or0;
  wire f_arrdiv32_fs63_xor0;
  wire f_arrdiv32_fs63_not0;
  wire f_arrdiv32_fs63_and0;
  wire f_arrdiv32_fs63_xor1;
  wire f_arrdiv32_fs63_not1;
  wire f_arrdiv32_fs63_and1;
  wire f_arrdiv32_fs63_or0;
  wire f_arrdiv32_mux2to131_and0;
  wire f_arrdiv32_mux2to131_not0;
  wire f_arrdiv32_mux2to131_and1;
  wire f_arrdiv32_mux2to131_xor0;
  wire f_arrdiv32_mux2to132_and0;
  wire f_arrdiv32_mux2to132_not0;
  wire f_arrdiv32_mux2to132_and1;
  wire f_arrdiv32_mux2to132_xor0;
  wire f_arrdiv32_mux2to133_and0;
  wire f_arrdiv32_mux2to133_not0;
  wire f_arrdiv32_mux2to133_and1;
  wire f_arrdiv32_mux2to133_xor0;
  wire f_arrdiv32_mux2to134_and0;
  wire f_arrdiv32_mux2to134_not0;
  wire f_arrdiv32_mux2to134_and1;
  wire f_arrdiv32_mux2to134_xor0;
  wire f_arrdiv32_mux2to135_and0;
  wire f_arrdiv32_mux2to135_not0;
  wire f_arrdiv32_mux2to135_and1;
  wire f_arrdiv32_mux2to135_xor0;
  wire f_arrdiv32_mux2to136_and0;
  wire f_arrdiv32_mux2to136_not0;
  wire f_arrdiv32_mux2to136_and1;
  wire f_arrdiv32_mux2to136_xor0;
  wire f_arrdiv32_mux2to137_and0;
  wire f_arrdiv32_mux2to137_not0;
  wire f_arrdiv32_mux2to137_and1;
  wire f_arrdiv32_mux2to137_xor0;
  wire f_arrdiv32_mux2to138_and0;
  wire f_arrdiv32_mux2to138_not0;
  wire f_arrdiv32_mux2to138_and1;
  wire f_arrdiv32_mux2to138_xor0;
  wire f_arrdiv32_mux2to139_and0;
  wire f_arrdiv32_mux2to139_not0;
  wire f_arrdiv32_mux2to139_and1;
  wire f_arrdiv32_mux2to139_xor0;
  wire f_arrdiv32_mux2to140_and0;
  wire f_arrdiv32_mux2to140_not0;
  wire f_arrdiv32_mux2to140_and1;
  wire f_arrdiv32_mux2to140_xor0;
  wire f_arrdiv32_mux2to141_and0;
  wire f_arrdiv32_mux2to141_not0;
  wire f_arrdiv32_mux2to141_and1;
  wire f_arrdiv32_mux2to141_xor0;
  wire f_arrdiv32_mux2to142_and0;
  wire f_arrdiv32_mux2to142_not0;
  wire f_arrdiv32_mux2to142_and1;
  wire f_arrdiv32_mux2to142_xor0;
  wire f_arrdiv32_mux2to143_and0;
  wire f_arrdiv32_mux2to143_not0;
  wire f_arrdiv32_mux2to143_and1;
  wire f_arrdiv32_mux2to143_xor0;
  wire f_arrdiv32_mux2to144_and0;
  wire f_arrdiv32_mux2to144_not0;
  wire f_arrdiv32_mux2to144_and1;
  wire f_arrdiv32_mux2to144_xor0;
  wire f_arrdiv32_mux2to145_and0;
  wire f_arrdiv32_mux2to145_not0;
  wire f_arrdiv32_mux2to145_and1;
  wire f_arrdiv32_mux2to145_xor0;
  wire f_arrdiv32_mux2to146_and0;
  wire f_arrdiv32_mux2to146_not0;
  wire f_arrdiv32_mux2to146_and1;
  wire f_arrdiv32_mux2to146_xor0;
  wire f_arrdiv32_mux2to147_and0;
  wire f_arrdiv32_mux2to147_not0;
  wire f_arrdiv32_mux2to147_and1;
  wire f_arrdiv32_mux2to147_xor0;
  wire f_arrdiv32_mux2to148_and0;
  wire f_arrdiv32_mux2to148_not0;
  wire f_arrdiv32_mux2to148_and1;
  wire f_arrdiv32_mux2to148_xor0;
  wire f_arrdiv32_mux2to149_and0;
  wire f_arrdiv32_mux2to149_not0;
  wire f_arrdiv32_mux2to149_and1;
  wire f_arrdiv32_mux2to149_xor0;
  wire f_arrdiv32_mux2to150_and0;
  wire f_arrdiv32_mux2to150_not0;
  wire f_arrdiv32_mux2to150_and1;
  wire f_arrdiv32_mux2to150_xor0;
  wire f_arrdiv32_mux2to151_and0;
  wire f_arrdiv32_mux2to151_not0;
  wire f_arrdiv32_mux2to151_and1;
  wire f_arrdiv32_mux2to151_xor0;
  wire f_arrdiv32_mux2to152_and0;
  wire f_arrdiv32_mux2to152_not0;
  wire f_arrdiv32_mux2to152_and1;
  wire f_arrdiv32_mux2to152_xor0;
  wire f_arrdiv32_mux2to153_and0;
  wire f_arrdiv32_mux2to153_not0;
  wire f_arrdiv32_mux2to153_and1;
  wire f_arrdiv32_mux2to153_xor0;
  wire f_arrdiv32_mux2to154_and0;
  wire f_arrdiv32_mux2to154_not0;
  wire f_arrdiv32_mux2to154_and1;
  wire f_arrdiv32_mux2to154_xor0;
  wire f_arrdiv32_mux2to155_and0;
  wire f_arrdiv32_mux2to155_not0;
  wire f_arrdiv32_mux2to155_and1;
  wire f_arrdiv32_mux2to155_xor0;
  wire f_arrdiv32_mux2to156_and0;
  wire f_arrdiv32_mux2to156_not0;
  wire f_arrdiv32_mux2to156_and1;
  wire f_arrdiv32_mux2to156_xor0;
  wire f_arrdiv32_mux2to157_and0;
  wire f_arrdiv32_mux2to157_not0;
  wire f_arrdiv32_mux2to157_and1;
  wire f_arrdiv32_mux2to157_xor0;
  wire f_arrdiv32_mux2to158_and0;
  wire f_arrdiv32_mux2to158_not0;
  wire f_arrdiv32_mux2to158_and1;
  wire f_arrdiv32_mux2to158_xor0;
  wire f_arrdiv32_mux2to159_and0;
  wire f_arrdiv32_mux2to159_not0;
  wire f_arrdiv32_mux2to159_and1;
  wire f_arrdiv32_mux2to159_xor0;
  wire f_arrdiv32_mux2to160_and0;
  wire f_arrdiv32_mux2to160_not0;
  wire f_arrdiv32_mux2to160_and1;
  wire f_arrdiv32_mux2to160_xor0;
  wire f_arrdiv32_mux2to161_and0;
  wire f_arrdiv32_mux2to161_not0;
  wire f_arrdiv32_mux2to161_and1;
  wire f_arrdiv32_mux2to161_xor0;
  wire f_arrdiv32_not1;
  wire f_arrdiv32_fs64_xor0;
  wire f_arrdiv32_fs64_not0;
  wire f_arrdiv32_fs64_and0;
  wire f_arrdiv32_fs64_not1;
  wire f_arrdiv32_fs65_xor0;
  wire f_arrdiv32_fs65_not0;
  wire f_arrdiv32_fs65_and0;
  wire f_arrdiv32_fs65_xor1;
  wire f_arrdiv32_fs65_not1;
  wire f_arrdiv32_fs65_and1;
  wire f_arrdiv32_fs65_or0;
  wire f_arrdiv32_fs66_xor0;
  wire f_arrdiv32_fs66_not0;
  wire f_arrdiv32_fs66_and0;
  wire f_arrdiv32_fs66_xor1;
  wire f_arrdiv32_fs66_not1;
  wire f_arrdiv32_fs66_and1;
  wire f_arrdiv32_fs66_or0;
  wire f_arrdiv32_fs67_xor0;
  wire f_arrdiv32_fs67_not0;
  wire f_arrdiv32_fs67_and0;
  wire f_arrdiv32_fs67_xor1;
  wire f_arrdiv32_fs67_not1;
  wire f_arrdiv32_fs67_and1;
  wire f_arrdiv32_fs67_or0;
  wire f_arrdiv32_fs68_xor0;
  wire f_arrdiv32_fs68_not0;
  wire f_arrdiv32_fs68_and0;
  wire f_arrdiv32_fs68_xor1;
  wire f_arrdiv32_fs68_not1;
  wire f_arrdiv32_fs68_and1;
  wire f_arrdiv32_fs68_or0;
  wire f_arrdiv32_fs69_xor0;
  wire f_arrdiv32_fs69_not0;
  wire f_arrdiv32_fs69_and0;
  wire f_arrdiv32_fs69_xor1;
  wire f_arrdiv32_fs69_not1;
  wire f_arrdiv32_fs69_and1;
  wire f_arrdiv32_fs69_or0;
  wire f_arrdiv32_fs70_xor0;
  wire f_arrdiv32_fs70_not0;
  wire f_arrdiv32_fs70_and0;
  wire f_arrdiv32_fs70_xor1;
  wire f_arrdiv32_fs70_not1;
  wire f_arrdiv32_fs70_and1;
  wire f_arrdiv32_fs70_or0;
  wire f_arrdiv32_fs71_xor0;
  wire f_arrdiv32_fs71_not0;
  wire f_arrdiv32_fs71_and0;
  wire f_arrdiv32_fs71_xor1;
  wire f_arrdiv32_fs71_not1;
  wire f_arrdiv32_fs71_and1;
  wire f_arrdiv32_fs71_or0;
  wire f_arrdiv32_fs72_xor0;
  wire f_arrdiv32_fs72_not0;
  wire f_arrdiv32_fs72_and0;
  wire f_arrdiv32_fs72_xor1;
  wire f_arrdiv32_fs72_not1;
  wire f_arrdiv32_fs72_and1;
  wire f_arrdiv32_fs72_or0;
  wire f_arrdiv32_fs73_xor0;
  wire f_arrdiv32_fs73_not0;
  wire f_arrdiv32_fs73_and0;
  wire f_arrdiv32_fs73_xor1;
  wire f_arrdiv32_fs73_not1;
  wire f_arrdiv32_fs73_and1;
  wire f_arrdiv32_fs73_or0;
  wire f_arrdiv32_fs74_xor0;
  wire f_arrdiv32_fs74_not0;
  wire f_arrdiv32_fs74_and0;
  wire f_arrdiv32_fs74_xor1;
  wire f_arrdiv32_fs74_not1;
  wire f_arrdiv32_fs74_and1;
  wire f_arrdiv32_fs74_or0;
  wire f_arrdiv32_fs75_xor0;
  wire f_arrdiv32_fs75_not0;
  wire f_arrdiv32_fs75_and0;
  wire f_arrdiv32_fs75_xor1;
  wire f_arrdiv32_fs75_not1;
  wire f_arrdiv32_fs75_and1;
  wire f_arrdiv32_fs75_or0;
  wire f_arrdiv32_fs76_xor0;
  wire f_arrdiv32_fs76_not0;
  wire f_arrdiv32_fs76_and0;
  wire f_arrdiv32_fs76_xor1;
  wire f_arrdiv32_fs76_not1;
  wire f_arrdiv32_fs76_and1;
  wire f_arrdiv32_fs76_or0;
  wire f_arrdiv32_fs77_xor0;
  wire f_arrdiv32_fs77_not0;
  wire f_arrdiv32_fs77_and0;
  wire f_arrdiv32_fs77_xor1;
  wire f_arrdiv32_fs77_not1;
  wire f_arrdiv32_fs77_and1;
  wire f_arrdiv32_fs77_or0;
  wire f_arrdiv32_fs78_xor0;
  wire f_arrdiv32_fs78_not0;
  wire f_arrdiv32_fs78_and0;
  wire f_arrdiv32_fs78_xor1;
  wire f_arrdiv32_fs78_not1;
  wire f_arrdiv32_fs78_and1;
  wire f_arrdiv32_fs78_or0;
  wire f_arrdiv32_fs79_xor0;
  wire f_arrdiv32_fs79_not0;
  wire f_arrdiv32_fs79_and0;
  wire f_arrdiv32_fs79_xor1;
  wire f_arrdiv32_fs79_not1;
  wire f_arrdiv32_fs79_and1;
  wire f_arrdiv32_fs79_or0;
  wire f_arrdiv32_fs80_xor0;
  wire f_arrdiv32_fs80_not0;
  wire f_arrdiv32_fs80_and0;
  wire f_arrdiv32_fs80_xor1;
  wire f_arrdiv32_fs80_not1;
  wire f_arrdiv32_fs80_and1;
  wire f_arrdiv32_fs80_or0;
  wire f_arrdiv32_fs81_xor0;
  wire f_arrdiv32_fs81_not0;
  wire f_arrdiv32_fs81_and0;
  wire f_arrdiv32_fs81_xor1;
  wire f_arrdiv32_fs81_not1;
  wire f_arrdiv32_fs81_and1;
  wire f_arrdiv32_fs81_or0;
  wire f_arrdiv32_fs82_xor0;
  wire f_arrdiv32_fs82_not0;
  wire f_arrdiv32_fs82_and0;
  wire f_arrdiv32_fs82_xor1;
  wire f_arrdiv32_fs82_not1;
  wire f_arrdiv32_fs82_and1;
  wire f_arrdiv32_fs82_or0;
  wire f_arrdiv32_fs83_xor0;
  wire f_arrdiv32_fs83_not0;
  wire f_arrdiv32_fs83_and0;
  wire f_arrdiv32_fs83_xor1;
  wire f_arrdiv32_fs83_not1;
  wire f_arrdiv32_fs83_and1;
  wire f_arrdiv32_fs83_or0;
  wire f_arrdiv32_fs84_xor0;
  wire f_arrdiv32_fs84_not0;
  wire f_arrdiv32_fs84_and0;
  wire f_arrdiv32_fs84_xor1;
  wire f_arrdiv32_fs84_not1;
  wire f_arrdiv32_fs84_and1;
  wire f_arrdiv32_fs84_or0;
  wire f_arrdiv32_fs85_xor0;
  wire f_arrdiv32_fs85_not0;
  wire f_arrdiv32_fs85_and0;
  wire f_arrdiv32_fs85_xor1;
  wire f_arrdiv32_fs85_not1;
  wire f_arrdiv32_fs85_and1;
  wire f_arrdiv32_fs85_or0;
  wire f_arrdiv32_fs86_xor0;
  wire f_arrdiv32_fs86_not0;
  wire f_arrdiv32_fs86_and0;
  wire f_arrdiv32_fs86_xor1;
  wire f_arrdiv32_fs86_not1;
  wire f_arrdiv32_fs86_and1;
  wire f_arrdiv32_fs86_or0;
  wire f_arrdiv32_fs87_xor0;
  wire f_arrdiv32_fs87_not0;
  wire f_arrdiv32_fs87_and0;
  wire f_arrdiv32_fs87_xor1;
  wire f_arrdiv32_fs87_not1;
  wire f_arrdiv32_fs87_and1;
  wire f_arrdiv32_fs87_or0;
  wire f_arrdiv32_fs88_xor0;
  wire f_arrdiv32_fs88_not0;
  wire f_arrdiv32_fs88_and0;
  wire f_arrdiv32_fs88_xor1;
  wire f_arrdiv32_fs88_not1;
  wire f_arrdiv32_fs88_and1;
  wire f_arrdiv32_fs88_or0;
  wire f_arrdiv32_fs89_xor0;
  wire f_arrdiv32_fs89_not0;
  wire f_arrdiv32_fs89_and0;
  wire f_arrdiv32_fs89_xor1;
  wire f_arrdiv32_fs89_not1;
  wire f_arrdiv32_fs89_and1;
  wire f_arrdiv32_fs89_or0;
  wire f_arrdiv32_fs90_xor0;
  wire f_arrdiv32_fs90_not0;
  wire f_arrdiv32_fs90_and0;
  wire f_arrdiv32_fs90_xor1;
  wire f_arrdiv32_fs90_not1;
  wire f_arrdiv32_fs90_and1;
  wire f_arrdiv32_fs90_or0;
  wire f_arrdiv32_fs91_xor0;
  wire f_arrdiv32_fs91_not0;
  wire f_arrdiv32_fs91_and0;
  wire f_arrdiv32_fs91_xor1;
  wire f_arrdiv32_fs91_not1;
  wire f_arrdiv32_fs91_and1;
  wire f_arrdiv32_fs91_or0;
  wire f_arrdiv32_fs92_xor0;
  wire f_arrdiv32_fs92_not0;
  wire f_arrdiv32_fs92_and0;
  wire f_arrdiv32_fs92_xor1;
  wire f_arrdiv32_fs92_not1;
  wire f_arrdiv32_fs92_and1;
  wire f_arrdiv32_fs92_or0;
  wire f_arrdiv32_fs93_xor0;
  wire f_arrdiv32_fs93_not0;
  wire f_arrdiv32_fs93_and0;
  wire f_arrdiv32_fs93_xor1;
  wire f_arrdiv32_fs93_not1;
  wire f_arrdiv32_fs93_and1;
  wire f_arrdiv32_fs93_or0;
  wire f_arrdiv32_fs94_xor0;
  wire f_arrdiv32_fs94_not0;
  wire f_arrdiv32_fs94_and0;
  wire f_arrdiv32_fs94_xor1;
  wire f_arrdiv32_fs94_not1;
  wire f_arrdiv32_fs94_and1;
  wire f_arrdiv32_fs94_or0;
  wire f_arrdiv32_fs95_xor0;
  wire f_arrdiv32_fs95_not0;
  wire f_arrdiv32_fs95_and0;
  wire f_arrdiv32_fs95_xor1;
  wire f_arrdiv32_fs95_not1;
  wire f_arrdiv32_fs95_and1;
  wire f_arrdiv32_fs95_or0;
  wire f_arrdiv32_mux2to162_and0;
  wire f_arrdiv32_mux2to162_not0;
  wire f_arrdiv32_mux2to162_and1;
  wire f_arrdiv32_mux2to162_xor0;
  wire f_arrdiv32_mux2to163_and0;
  wire f_arrdiv32_mux2to163_not0;
  wire f_arrdiv32_mux2to163_and1;
  wire f_arrdiv32_mux2to163_xor0;
  wire f_arrdiv32_mux2to164_and0;
  wire f_arrdiv32_mux2to164_not0;
  wire f_arrdiv32_mux2to164_and1;
  wire f_arrdiv32_mux2to164_xor0;
  wire f_arrdiv32_mux2to165_and0;
  wire f_arrdiv32_mux2to165_not0;
  wire f_arrdiv32_mux2to165_and1;
  wire f_arrdiv32_mux2to165_xor0;
  wire f_arrdiv32_mux2to166_and0;
  wire f_arrdiv32_mux2to166_not0;
  wire f_arrdiv32_mux2to166_and1;
  wire f_arrdiv32_mux2to166_xor0;
  wire f_arrdiv32_mux2to167_and0;
  wire f_arrdiv32_mux2to167_not0;
  wire f_arrdiv32_mux2to167_and1;
  wire f_arrdiv32_mux2to167_xor0;
  wire f_arrdiv32_mux2to168_and0;
  wire f_arrdiv32_mux2to168_not0;
  wire f_arrdiv32_mux2to168_and1;
  wire f_arrdiv32_mux2to168_xor0;
  wire f_arrdiv32_mux2to169_and0;
  wire f_arrdiv32_mux2to169_not0;
  wire f_arrdiv32_mux2to169_and1;
  wire f_arrdiv32_mux2to169_xor0;
  wire f_arrdiv32_mux2to170_and0;
  wire f_arrdiv32_mux2to170_not0;
  wire f_arrdiv32_mux2to170_and1;
  wire f_arrdiv32_mux2to170_xor0;
  wire f_arrdiv32_mux2to171_and0;
  wire f_arrdiv32_mux2to171_not0;
  wire f_arrdiv32_mux2to171_and1;
  wire f_arrdiv32_mux2to171_xor0;
  wire f_arrdiv32_mux2to172_and0;
  wire f_arrdiv32_mux2to172_not0;
  wire f_arrdiv32_mux2to172_and1;
  wire f_arrdiv32_mux2to172_xor0;
  wire f_arrdiv32_mux2to173_and0;
  wire f_arrdiv32_mux2to173_not0;
  wire f_arrdiv32_mux2to173_and1;
  wire f_arrdiv32_mux2to173_xor0;
  wire f_arrdiv32_mux2to174_and0;
  wire f_arrdiv32_mux2to174_not0;
  wire f_arrdiv32_mux2to174_and1;
  wire f_arrdiv32_mux2to174_xor0;
  wire f_arrdiv32_mux2to175_and0;
  wire f_arrdiv32_mux2to175_not0;
  wire f_arrdiv32_mux2to175_and1;
  wire f_arrdiv32_mux2to175_xor0;
  wire f_arrdiv32_mux2to176_and0;
  wire f_arrdiv32_mux2to176_not0;
  wire f_arrdiv32_mux2to176_and1;
  wire f_arrdiv32_mux2to176_xor0;
  wire f_arrdiv32_mux2to177_and0;
  wire f_arrdiv32_mux2to177_not0;
  wire f_arrdiv32_mux2to177_and1;
  wire f_arrdiv32_mux2to177_xor0;
  wire f_arrdiv32_mux2to178_and0;
  wire f_arrdiv32_mux2to178_not0;
  wire f_arrdiv32_mux2to178_and1;
  wire f_arrdiv32_mux2to178_xor0;
  wire f_arrdiv32_mux2to179_and0;
  wire f_arrdiv32_mux2to179_not0;
  wire f_arrdiv32_mux2to179_and1;
  wire f_arrdiv32_mux2to179_xor0;
  wire f_arrdiv32_mux2to180_and0;
  wire f_arrdiv32_mux2to180_not0;
  wire f_arrdiv32_mux2to180_and1;
  wire f_arrdiv32_mux2to180_xor0;
  wire f_arrdiv32_mux2to181_and0;
  wire f_arrdiv32_mux2to181_not0;
  wire f_arrdiv32_mux2to181_and1;
  wire f_arrdiv32_mux2to181_xor0;
  wire f_arrdiv32_mux2to182_and0;
  wire f_arrdiv32_mux2to182_not0;
  wire f_arrdiv32_mux2to182_and1;
  wire f_arrdiv32_mux2to182_xor0;
  wire f_arrdiv32_mux2to183_and0;
  wire f_arrdiv32_mux2to183_not0;
  wire f_arrdiv32_mux2to183_and1;
  wire f_arrdiv32_mux2to183_xor0;
  wire f_arrdiv32_mux2to184_and0;
  wire f_arrdiv32_mux2to184_not0;
  wire f_arrdiv32_mux2to184_and1;
  wire f_arrdiv32_mux2to184_xor0;
  wire f_arrdiv32_mux2to185_and0;
  wire f_arrdiv32_mux2to185_not0;
  wire f_arrdiv32_mux2to185_and1;
  wire f_arrdiv32_mux2to185_xor0;
  wire f_arrdiv32_mux2to186_and0;
  wire f_arrdiv32_mux2to186_not0;
  wire f_arrdiv32_mux2to186_and1;
  wire f_arrdiv32_mux2to186_xor0;
  wire f_arrdiv32_mux2to187_and0;
  wire f_arrdiv32_mux2to187_not0;
  wire f_arrdiv32_mux2to187_and1;
  wire f_arrdiv32_mux2to187_xor0;
  wire f_arrdiv32_mux2to188_and0;
  wire f_arrdiv32_mux2to188_not0;
  wire f_arrdiv32_mux2to188_and1;
  wire f_arrdiv32_mux2to188_xor0;
  wire f_arrdiv32_mux2to189_and0;
  wire f_arrdiv32_mux2to189_not0;
  wire f_arrdiv32_mux2to189_and1;
  wire f_arrdiv32_mux2to189_xor0;
  wire f_arrdiv32_mux2to190_and0;
  wire f_arrdiv32_mux2to190_not0;
  wire f_arrdiv32_mux2to190_and1;
  wire f_arrdiv32_mux2to190_xor0;
  wire f_arrdiv32_mux2to191_and0;
  wire f_arrdiv32_mux2to191_not0;
  wire f_arrdiv32_mux2to191_and1;
  wire f_arrdiv32_mux2to191_xor0;
  wire f_arrdiv32_mux2to192_and0;
  wire f_arrdiv32_mux2to192_not0;
  wire f_arrdiv32_mux2to192_and1;
  wire f_arrdiv32_mux2to192_xor0;
  wire f_arrdiv32_not2;
  wire f_arrdiv32_fs96_xor0;
  wire f_arrdiv32_fs96_not0;
  wire f_arrdiv32_fs96_and0;
  wire f_arrdiv32_fs96_not1;
  wire f_arrdiv32_fs97_xor0;
  wire f_arrdiv32_fs97_not0;
  wire f_arrdiv32_fs97_and0;
  wire f_arrdiv32_fs97_xor1;
  wire f_arrdiv32_fs97_not1;
  wire f_arrdiv32_fs97_and1;
  wire f_arrdiv32_fs97_or0;
  wire f_arrdiv32_fs98_xor0;
  wire f_arrdiv32_fs98_not0;
  wire f_arrdiv32_fs98_and0;
  wire f_arrdiv32_fs98_xor1;
  wire f_arrdiv32_fs98_not1;
  wire f_arrdiv32_fs98_and1;
  wire f_arrdiv32_fs98_or0;
  wire f_arrdiv32_fs99_xor0;
  wire f_arrdiv32_fs99_not0;
  wire f_arrdiv32_fs99_and0;
  wire f_arrdiv32_fs99_xor1;
  wire f_arrdiv32_fs99_not1;
  wire f_arrdiv32_fs99_and1;
  wire f_arrdiv32_fs99_or0;
  wire f_arrdiv32_fs100_xor0;
  wire f_arrdiv32_fs100_not0;
  wire f_arrdiv32_fs100_and0;
  wire f_arrdiv32_fs100_xor1;
  wire f_arrdiv32_fs100_not1;
  wire f_arrdiv32_fs100_and1;
  wire f_arrdiv32_fs100_or0;
  wire f_arrdiv32_fs101_xor0;
  wire f_arrdiv32_fs101_not0;
  wire f_arrdiv32_fs101_and0;
  wire f_arrdiv32_fs101_xor1;
  wire f_arrdiv32_fs101_not1;
  wire f_arrdiv32_fs101_and1;
  wire f_arrdiv32_fs101_or0;
  wire f_arrdiv32_fs102_xor0;
  wire f_arrdiv32_fs102_not0;
  wire f_arrdiv32_fs102_and0;
  wire f_arrdiv32_fs102_xor1;
  wire f_arrdiv32_fs102_not1;
  wire f_arrdiv32_fs102_and1;
  wire f_arrdiv32_fs102_or0;
  wire f_arrdiv32_fs103_xor0;
  wire f_arrdiv32_fs103_not0;
  wire f_arrdiv32_fs103_and0;
  wire f_arrdiv32_fs103_xor1;
  wire f_arrdiv32_fs103_not1;
  wire f_arrdiv32_fs103_and1;
  wire f_arrdiv32_fs103_or0;
  wire f_arrdiv32_fs104_xor0;
  wire f_arrdiv32_fs104_not0;
  wire f_arrdiv32_fs104_and0;
  wire f_arrdiv32_fs104_xor1;
  wire f_arrdiv32_fs104_not1;
  wire f_arrdiv32_fs104_and1;
  wire f_arrdiv32_fs104_or0;
  wire f_arrdiv32_fs105_xor0;
  wire f_arrdiv32_fs105_not0;
  wire f_arrdiv32_fs105_and0;
  wire f_arrdiv32_fs105_xor1;
  wire f_arrdiv32_fs105_not1;
  wire f_arrdiv32_fs105_and1;
  wire f_arrdiv32_fs105_or0;
  wire f_arrdiv32_fs106_xor0;
  wire f_arrdiv32_fs106_not0;
  wire f_arrdiv32_fs106_and0;
  wire f_arrdiv32_fs106_xor1;
  wire f_arrdiv32_fs106_not1;
  wire f_arrdiv32_fs106_and1;
  wire f_arrdiv32_fs106_or0;
  wire f_arrdiv32_fs107_xor0;
  wire f_arrdiv32_fs107_not0;
  wire f_arrdiv32_fs107_and0;
  wire f_arrdiv32_fs107_xor1;
  wire f_arrdiv32_fs107_not1;
  wire f_arrdiv32_fs107_and1;
  wire f_arrdiv32_fs107_or0;
  wire f_arrdiv32_fs108_xor0;
  wire f_arrdiv32_fs108_not0;
  wire f_arrdiv32_fs108_and0;
  wire f_arrdiv32_fs108_xor1;
  wire f_arrdiv32_fs108_not1;
  wire f_arrdiv32_fs108_and1;
  wire f_arrdiv32_fs108_or0;
  wire f_arrdiv32_fs109_xor0;
  wire f_arrdiv32_fs109_not0;
  wire f_arrdiv32_fs109_and0;
  wire f_arrdiv32_fs109_xor1;
  wire f_arrdiv32_fs109_not1;
  wire f_arrdiv32_fs109_and1;
  wire f_arrdiv32_fs109_or0;
  wire f_arrdiv32_fs110_xor0;
  wire f_arrdiv32_fs110_not0;
  wire f_arrdiv32_fs110_and0;
  wire f_arrdiv32_fs110_xor1;
  wire f_arrdiv32_fs110_not1;
  wire f_arrdiv32_fs110_and1;
  wire f_arrdiv32_fs110_or0;
  wire f_arrdiv32_fs111_xor0;
  wire f_arrdiv32_fs111_not0;
  wire f_arrdiv32_fs111_and0;
  wire f_arrdiv32_fs111_xor1;
  wire f_arrdiv32_fs111_not1;
  wire f_arrdiv32_fs111_and1;
  wire f_arrdiv32_fs111_or0;
  wire f_arrdiv32_fs112_xor0;
  wire f_arrdiv32_fs112_not0;
  wire f_arrdiv32_fs112_and0;
  wire f_arrdiv32_fs112_xor1;
  wire f_arrdiv32_fs112_not1;
  wire f_arrdiv32_fs112_and1;
  wire f_arrdiv32_fs112_or0;
  wire f_arrdiv32_fs113_xor0;
  wire f_arrdiv32_fs113_not0;
  wire f_arrdiv32_fs113_and0;
  wire f_arrdiv32_fs113_xor1;
  wire f_arrdiv32_fs113_not1;
  wire f_arrdiv32_fs113_and1;
  wire f_arrdiv32_fs113_or0;
  wire f_arrdiv32_fs114_xor0;
  wire f_arrdiv32_fs114_not0;
  wire f_arrdiv32_fs114_and0;
  wire f_arrdiv32_fs114_xor1;
  wire f_arrdiv32_fs114_not1;
  wire f_arrdiv32_fs114_and1;
  wire f_arrdiv32_fs114_or0;
  wire f_arrdiv32_fs115_xor0;
  wire f_arrdiv32_fs115_not0;
  wire f_arrdiv32_fs115_and0;
  wire f_arrdiv32_fs115_xor1;
  wire f_arrdiv32_fs115_not1;
  wire f_arrdiv32_fs115_and1;
  wire f_arrdiv32_fs115_or0;
  wire f_arrdiv32_fs116_xor0;
  wire f_arrdiv32_fs116_not0;
  wire f_arrdiv32_fs116_and0;
  wire f_arrdiv32_fs116_xor1;
  wire f_arrdiv32_fs116_not1;
  wire f_arrdiv32_fs116_and1;
  wire f_arrdiv32_fs116_or0;
  wire f_arrdiv32_fs117_xor0;
  wire f_arrdiv32_fs117_not0;
  wire f_arrdiv32_fs117_and0;
  wire f_arrdiv32_fs117_xor1;
  wire f_arrdiv32_fs117_not1;
  wire f_arrdiv32_fs117_and1;
  wire f_arrdiv32_fs117_or0;
  wire f_arrdiv32_fs118_xor0;
  wire f_arrdiv32_fs118_not0;
  wire f_arrdiv32_fs118_and0;
  wire f_arrdiv32_fs118_xor1;
  wire f_arrdiv32_fs118_not1;
  wire f_arrdiv32_fs118_and1;
  wire f_arrdiv32_fs118_or0;
  wire f_arrdiv32_fs119_xor0;
  wire f_arrdiv32_fs119_not0;
  wire f_arrdiv32_fs119_and0;
  wire f_arrdiv32_fs119_xor1;
  wire f_arrdiv32_fs119_not1;
  wire f_arrdiv32_fs119_and1;
  wire f_arrdiv32_fs119_or0;
  wire f_arrdiv32_fs120_xor0;
  wire f_arrdiv32_fs120_not0;
  wire f_arrdiv32_fs120_and0;
  wire f_arrdiv32_fs120_xor1;
  wire f_arrdiv32_fs120_not1;
  wire f_arrdiv32_fs120_and1;
  wire f_arrdiv32_fs120_or0;
  wire f_arrdiv32_fs121_xor0;
  wire f_arrdiv32_fs121_not0;
  wire f_arrdiv32_fs121_and0;
  wire f_arrdiv32_fs121_xor1;
  wire f_arrdiv32_fs121_not1;
  wire f_arrdiv32_fs121_and1;
  wire f_arrdiv32_fs121_or0;
  wire f_arrdiv32_fs122_xor0;
  wire f_arrdiv32_fs122_not0;
  wire f_arrdiv32_fs122_and0;
  wire f_arrdiv32_fs122_xor1;
  wire f_arrdiv32_fs122_not1;
  wire f_arrdiv32_fs122_and1;
  wire f_arrdiv32_fs122_or0;
  wire f_arrdiv32_fs123_xor0;
  wire f_arrdiv32_fs123_not0;
  wire f_arrdiv32_fs123_and0;
  wire f_arrdiv32_fs123_xor1;
  wire f_arrdiv32_fs123_not1;
  wire f_arrdiv32_fs123_and1;
  wire f_arrdiv32_fs123_or0;
  wire f_arrdiv32_fs124_xor0;
  wire f_arrdiv32_fs124_not0;
  wire f_arrdiv32_fs124_and0;
  wire f_arrdiv32_fs124_xor1;
  wire f_arrdiv32_fs124_not1;
  wire f_arrdiv32_fs124_and1;
  wire f_arrdiv32_fs124_or0;
  wire f_arrdiv32_fs125_xor0;
  wire f_arrdiv32_fs125_not0;
  wire f_arrdiv32_fs125_and0;
  wire f_arrdiv32_fs125_xor1;
  wire f_arrdiv32_fs125_not1;
  wire f_arrdiv32_fs125_and1;
  wire f_arrdiv32_fs125_or0;
  wire f_arrdiv32_fs126_xor0;
  wire f_arrdiv32_fs126_not0;
  wire f_arrdiv32_fs126_and0;
  wire f_arrdiv32_fs126_xor1;
  wire f_arrdiv32_fs126_not1;
  wire f_arrdiv32_fs126_and1;
  wire f_arrdiv32_fs126_or0;
  wire f_arrdiv32_fs127_xor0;
  wire f_arrdiv32_fs127_not0;
  wire f_arrdiv32_fs127_and0;
  wire f_arrdiv32_fs127_xor1;
  wire f_arrdiv32_fs127_not1;
  wire f_arrdiv32_fs127_and1;
  wire f_arrdiv32_fs127_or0;
  wire f_arrdiv32_mux2to193_and0;
  wire f_arrdiv32_mux2to193_not0;
  wire f_arrdiv32_mux2to193_and1;
  wire f_arrdiv32_mux2to193_xor0;
  wire f_arrdiv32_mux2to194_and0;
  wire f_arrdiv32_mux2to194_not0;
  wire f_arrdiv32_mux2to194_and1;
  wire f_arrdiv32_mux2to194_xor0;
  wire f_arrdiv32_mux2to195_and0;
  wire f_arrdiv32_mux2to195_not0;
  wire f_arrdiv32_mux2to195_and1;
  wire f_arrdiv32_mux2to195_xor0;
  wire f_arrdiv32_mux2to196_and0;
  wire f_arrdiv32_mux2to196_not0;
  wire f_arrdiv32_mux2to196_and1;
  wire f_arrdiv32_mux2to196_xor0;
  wire f_arrdiv32_mux2to197_and0;
  wire f_arrdiv32_mux2to197_not0;
  wire f_arrdiv32_mux2to197_and1;
  wire f_arrdiv32_mux2to197_xor0;
  wire f_arrdiv32_mux2to198_and0;
  wire f_arrdiv32_mux2to198_not0;
  wire f_arrdiv32_mux2to198_and1;
  wire f_arrdiv32_mux2to198_xor0;
  wire f_arrdiv32_mux2to199_and0;
  wire f_arrdiv32_mux2to199_not0;
  wire f_arrdiv32_mux2to199_and1;
  wire f_arrdiv32_mux2to199_xor0;
  wire f_arrdiv32_mux2to1100_and0;
  wire f_arrdiv32_mux2to1100_not0;
  wire f_arrdiv32_mux2to1100_and1;
  wire f_arrdiv32_mux2to1100_xor0;
  wire f_arrdiv32_mux2to1101_and0;
  wire f_arrdiv32_mux2to1101_not0;
  wire f_arrdiv32_mux2to1101_and1;
  wire f_arrdiv32_mux2to1101_xor0;
  wire f_arrdiv32_mux2to1102_and0;
  wire f_arrdiv32_mux2to1102_not0;
  wire f_arrdiv32_mux2to1102_and1;
  wire f_arrdiv32_mux2to1102_xor0;
  wire f_arrdiv32_mux2to1103_and0;
  wire f_arrdiv32_mux2to1103_not0;
  wire f_arrdiv32_mux2to1103_and1;
  wire f_arrdiv32_mux2to1103_xor0;
  wire f_arrdiv32_mux2to1104_and0;
  wire f_arrdiv32_mux2to1104_not0;
  wire f_arrdiv32_mux2to1104_and1;
  wire f_arrdiv32_mux2to1104_xor0;
  wire f_arrdiv32_mux2to1105_and0;
  wire f_arrdiv32_mux2to1105_not0;
  wire f_arrdiv32_mux2to1105_and1;
  wire f_arrdiv32_mux2to1105_xor0;
  wire f_arrdiv32_mux2to1106_and0;
  wire f_arrdiv32_mux2to1106_not0;
  wire f_arrdiv32_mux2to1106_and1;
  wire f_arrdiv32_mux2to1106_xor0;
  wire f_arrdiv32_mux2to1107_and0;
  wire f_arrdiv32_mux2to1107_not0;
  wire f_arrdiv32_mux2to1107_and1;
  wire f_arrdiv32_mux2to1107_xor0;
  wire f_arrdiv32_mux2to1108_and0;
  wire f_arrdiv32_mux2to1108_not0;
  wire f_arrdiv32_mux2to1108_and1;
  wire f_arrdiv32_mux2to1108_xor0;
  wire f_arrdiv32_mux2to1109_and0;
  wire f_arrdiv32_mux2to1109_not0;
  wire f_arrdiv32_mux2to1109_and1;
  wire f_arrdiv32_mux2to1109_xor0;
  wire f_arrdiv32_mux2to1110_and0;
  wire f_arrdiv32_mux2to1110_not0;
  wire f_arrdiv32_mux2to1110_and1;
  wire f_arrdiv32_mux2to1110_xor0;
  wire f_arrdiv32_mux2to1111_and0;
  wire f_arrdiv32_mux2to1111_not0;
  wire f_arrdiv32_mux2to1111_and1;
  wire f_arrdiv32_mux2to1111_xor0;
  wire f_arrdiv32_mux2to1112_and0;
  wire f_arrdiv32_mux2to1112_not0;
  wire f_arrdiv32_mux2to1112_and1;
  wire f_arrdiv32_mux2to1112_xor0;
  wire f_arrdiv32_mux2to1113_and0;
  wire f_arrdiv32_mux2to1113_not0;
  wire f_arrdiv32_mux2to1113_and1;
  wire f_arrdiv32_mux2to1113_xor0;
  wire f_arrdiv32_mux2to1114_and0;
  wire f_arrdiv32_mux2to1114_not0;
  wire f_arrdiv32_mux2to1114_and1;
  wire f_arrdiv32_mux2to1114_xor0;
  wire f_arrdiv32_mux2to1115_and0;
  wire f_arrdiv32_mux2to1115_not0;
  wire f_arrdiv32_mux2to1115_and1;
  wire f_arrdiv32_mux2to1115_xor0;
  wire f_arrdiv32_mux2to1116_and0;
  wire f_arrdiv32_mux2to1116_not0;
  wire f_arrdiv32_mux2to1116_and1;
  wire f_arrdiv32_mux2to1116_xor0;
  wire f_arrdiv32_mux2to1117_and0;
  wire f_arrdiv32_mux2to1117_not0;
  wire f_arrdiv32_mux2to1117_and1;
  wire f_arrdiv32_mux2to1117_xor0;
  wire f_arrdiv32_mux2to1118_and0;
  wire f_arrdiv32_mux2to1118_not0;
  wire f_arrdiv32_mux2to1118_and1;
  wire f_arrdiv32_mux2to1118_xor0;
  wire f_arrdiv32_mux2to1119_and0;
  wire f_arrdiv32_mux2to1119_not0;
  wire f_arrdiv32_mux2to1119_and1;
  wire f_arrdiv32_mux2to1119_xor0;
  wire f_arrdiv32_mux2to1120_and0;
  wire f_arrdiv32_mux2to1120_not0;
  wire f_arrdiv32_mux2to1120_and1;
  wire f_arrdiv32_mux2to1120_xor0;
  wire f_arrdiv32_mux2to1121_and0;
  wire f_arrdiv32_mux2to1121_not0;
  wire f_arrdiv32_mux2to1121_and1;
  wire f_arrdiv32_mux2to1121_xor0;
  wire f_arrdiv32_mux2to1122_and0;
  wire f_arrdiv32_mux2to1122_not0;
  wire f_arrdiv32_mux2to1122_and1;
  wire f_arrdiv32_mux2to1122_xor0;
  wire f_arrdiv32_mux2to1123_and0;
  wire f_arrdiv32_mux2to1123_not0;
  wire f_arrdiv32_mux2to1123_and1;
  wire f_arrdiv32_mux2to1123_xor0;
  wire f_arrdiv32_not3;
  wire f_arrdiv32_fs128_xor0;
  wire f_arrdiv32_fs128_not0;
  wire f_arrdiv32_fs128_and0;
  wire f_arrdiv32_fs128_not1;
  wire f_arrdiv32_fs129_xor0;
  wire f_arrdiv32_fs129_not0;
  wire f_arrdiv32_fs129_and0;
  wire f_arrdiv32_fs129_xor1;
  wire f_arrdiv32_fs129_not1;
  wire f_arrdiv32_fs129_and1;
  wire f_arrdiv32_fs129_or0;
  wire f_arrdiv32_fs130_xor0;
  wire f_arrdiv32_fs130_not0;
  wire f_arrdiv32_fs130_and0;
  wire f_arrdiv32_fs130_xor1;
  wire f_arrdiv32_fs130_not1;
  wire f_arrdiv32_fs130_and1;
  wire f_arrdiv32_fs130_or0;
  wire f_arrdiv32_fs131_xor0;
  wire f_arrdiv32_fs131_not0;
  wire f_arrdiv32_fs131_and0;
  wire f_arrdiv32_fs131_xor1;
  wire f_arrdiv32_fs131_not1;
  wire f_arrdiv32_fs131_and1;
  wire f_arrdiv32_fs131_or0;
  wire f_arrdiv32_fs132_xor0;
  wire f_arrdiv32_fs132_not0;
  wire f_arrdiv32_fs132_and0;
  wire f_arrdiv32_fs132_xor1;
  wire f_arrdiv32_fs132_not1;
  wire f_arrdiv32_fs132_and1;
  wire f_arrdiv32_fs132_or0;
  wire f_arrdiv32_fs133_xor0;
  wire f_arrdiv32_fs133_not0;
  wire f_arrdiv32_fs133_and0;
  wire f_arrdiv32_fs133_xor1;
  wire f_arrdiv32_fs133_not1;
  wire f_arrdiv32_fs133_and1;
  wire f_arrdiv32_fs133_or0;
  wire f_arrdiv32_fs134_xor0;
  wire f_arrdiv32_fs134_not0;
  wire f_arrdiv32_fs134_and0;
  wire f_arrdiv32_fs134_xor1;
  wire f_arrdiv32_fs134_not1;
  wire f_arrdiv32_fs134_and1;
  wire f_arrdiv32_fs134_or0;
  wire f_arrdiv32_fs135_xor0;
  wire f_arrdiv32_fs135_not0;
  wire f_arrdiv32_fs135_and0;
  wire f_arrdiv32_fs135_xor1;
  wire f_arrdiv32_fs135_not1;
  wire f_arrdiv32_fs135_and1;
  wire f_arrdiv32_fs135_or0;
  wire f_arrdiv32_fs136_xor0;
  wire f_arrdiv32_fs136_not0;
  wire f_arrdiv32_fs136_and0;
  wire f_arrdiv32_fs136_xor1;
  wire f_arrdiv32_fs136_not1;
  wire f_arrdiv32_fs136_and1;
  wire f_arrdiv32_fs136_or0;
  wire f_arrdiv32_fs137_xor0;
  wire f_arrdiv32_fs137_not0;
  wire f_arrdiv32_fs137_and0;
  wire f_arrdiv32_fs137_xor1;
  wire f_arrdiv32_fs137_not1;
  wire f_arrdiv32_fs137_and1;
  wire f_arrdiv32_fs137_or0;
  wire f_arrdiv32_fs138_xor0;
  wire f_arrdiv32_fs138_not0;
  wire f_arrdiv32_fs138_and0;
  wire f_arrdiv32_fs138_xor1;
  wire f_arrdiv32_fs138_not1;
  wire f_arrdiv32_fs138_and1;
  wire f_arrdiv32_fs138_or0;
  wire f_arrdiv32_fs139_xor0;
  wire f_arrdiv32_fs139_not0;
  wire f_arrdiv32_fs139_and0;
  wire f_arrdiv32_fs139_xor1;
  wire f_arrdiv32_fs139_not1;
  wire f_arrdiv32_fs139_and1;
  wire f_arrdiv32_fs139_or0;
  wire f_arrdiv32_fs140_xor0;
  wire f_arrdiv32_fs140_not0;
  wire f_arrdiv32_fs140_and0;
  wire f_arrdiv32_fs140_xor1;
  wire f_arrdiv32_fs140_not1;
  wire f_arrdiv32_fs140_and1;
  wire f_arrdiv32_fs140_or0;
  wire f_arrdiv32_fs141_xor0;
  wire f_arrdiv32_fs141_not0;
  wire f_arrdiv32_fs141_and0;
  wire f_arrdiv32_fs141_xor1;
  wire f_arrdiv32_fs141_not1;
  wire f_arrdiv32_fs141_and1;
  wire f_arrdiv32_fs141_or0;
  wire f_arrdiv32_fs142_xor0;
  wire f_arrdiv32_fs142_not0;
  wire f_arrdiv32_fs142_and0;
  wire f_arrdiv32_fs142_xor1;
  wire f_arrdiv32_fs142_not1;
  wire f_arrdiv32_fs142_and1;
  wire f_arrdiv32_fs142_or0;
  wire f_arrdiv32_fs143_xor0;
  wire f_arrdiv32_fs143_not0;
  wire f_arrdiv32_fs143_and0;
  wire f_arrdiv32_fs143_xor1;
  wire f_arrdiv32_fs143_not1;
  wire f_arrdiv32_fs143_and1;
  wire f_arrdiv32_fs143_or0;
  wire f_arrdiv32_fs144_xor0;
  wire f_arrdiv32_fs144_not0;
  wire f_arrdiv32_fs144_and0;
  wire f_arrdiv32_fs144_xor1;
  wire f_arrdiv32_fs144_not1;
  wire f_arrdiv32_fs144_and1;
  wire f_arrdiv32_fs144_or0;
  wire f_arrdiv32_fs145_xor0;
  wire f_arrdiv32_fs145_not0;
  wire f_arrdiv32_fs145_and0;
  wire f_arrdiv32_fs145_xor1;
  wire f_arrdiv32_fs145_not1;
  wire f_arrdiv32_fs145_and1;
  wire f_arrdiv32_fs145_or0;
  wire f_arrdiv32_fs146_xor0;
  wire f_arrdiv32_fs146_not0;
  wire f_arrdiv32_fs146_and0;
  wire f_arrdiv32_fs146_xor1;
  wire f_arrdiv32_fs146_not1;
  wire f_arrdiv32_fs146_and1;
  wire f_arrdiv32_fs146_or0;
  wire f_arrdiv32_fs147_xor0;
  wire f_arrdiv32_fs147_not0;
  wire f_arrdiv32_fs147_and0;
  wire f_arrdiv32_fs147_xor1;
  wire f_arrdiv32_fs147_not1;
  wire f_arrdiv32_fs147_and1;
  wire f_arrdiv32_fs147_or0;
  wire f_arrdiv32_fs148_xor0;
  wire f_arrdiv32_fs148_not0;
  wire f_arrdiv32_fs148_and0;
  wire f_arrdiv32_fs148_xor1;
  wire f_arrdiv32_fs148_not1;
  wire f_arrdiv32_fs148_and1;
  wire f_arrdiv32_fs148_or0;
  wire f_arrdiv32_fs149_xor0;
  wire f_arrdiv32_fs149_not0;
  wire f_arrdiv32_fs149_and0;
  wire f_arrdiv32_fs149_xor1;
  wire f_arrdiv32_fs149_not1;
  wire f_arrdiv32_fs149_and1;
  wire f_arrdiv32_fs149_or0;
  wire f_arrdiv32_fs150_xor0;
  wire f_arrdiv32_fs150_not0;
  wire f_arrdiv32_fs150_and0;
  wire f_arrdiv32_fs150_xor1;
  wire f_arrdiv32_fs150_not1;
  wire f_arrdiv32_fs150_and1;
  wire f_arrdiv32_fs150_or0;
  wire f_arrdiv32_fs151_xor0;
  wire f_arrdiv32_fs151_not0;
  wire f_arrdiv32_fs151_and0;
  wire f_arrdiv32_fs151_xor1;
  wire f_arrdiv32_fs151_not1;
  wire f_arrdiv32_fs151_and1;
  wire f_arrdiv32_fs151_or0;
  wire f_arrdiv32_fs152_xor0;
  wire f_arrdiv32_fs152_not0;
  wire f_arrdiv32_fs152_and0;
  wire f_arrdiv32_fs152_xor1;
  wire f_arrdiv32_fs152_not1;
  wire f_arrdiv32_fs152_and1;
  wire f_arrdiv32_fs152_or0;
  wire f_arrdiv32_fs153_xor0;
  wire f_arrdiv32_fs153_not0;
  wire f_arrdiv32_fs153_and0;
  wire f_arrdiv32_fs153_xor1;
  wire f_arrdiv32_fs153_not1;
  wire f_arrdiv32_fs153_and1;
  wire f_arrdiv32_fs153_or0;
  wire f_arrdiv32_fs154_xor0;
  wire f_arrdiv32_fs154_not0;
  wire f_arrdiv32_fs154_and0;
  wire f_arrdiv32_fs154_xor1;
  wire f_arrdiv32_fs154_not1;
  wire f_arrdiv32_fs154_and1;
  wire f_arrdiv32_fs154_or0;
  wire f_arrdiv32_fs155_xor0;
  wire f_arrdiv32_fs155_not0;
  wire f_arrdiv32_fs155_and0;
  wire f_arrdiv32_fs155_xor1;
  wire f_arrdiv32_fs155_not1;
  wire f_arrdiv32_fs155_and1;
  wire f_arrdiv32_fs155_or0;
  wire f_arrdiv32_fs156_xor0;
  wire f_arrdiv32_fs156_not0;
  wire f_arrdiv32_fs156_and0;
  wire f_arrdiv32_fs156_xor1;
  wire f_arrdiv32_fs156_not1;
  wire f_arrdiv32_fs156_and1;
  wire f_arrdiv32_fs156_or0;
  wire f_arrdiv32_fs157_xor0;
  wire f_arrdiv32_fs157_not0;
  wire f_arrdiv32_fs157_and0;
  wire f_arrdiv32_fs157_xor1;
  wire f_arrdiv32_fs157_not1;
  wire f_arrdiv32_fs157_and1;
  wire f_arrdiv32_fs157_or0;
  wire f_arrdiv32_fs158_xor0;
  wire f_arrdiv32_fs158_not0;
  wire f_arrdiv32_fs158_and0;
  wire f_arrdiv32_fs158_xor1;
  wire f_arrdiv32_fs158_not1;
  wire f_arrdiv32_fs158_and1;
  wire f_arrdiv32_fs158_or0;
  wire f_arrdiv32_fs159_xor0;
  wire f_arrdiv32_fs159_not0;
  wire f_arrdiv32_fs159_and0;
  wire f_arrdiv32_fs159_xor1;
  wire f_arrdiv32_fs159_not1;
  wire f_arrdiv32_fs159_and1;
  wire f_arrdiv32_fs159_or0;
  wire f_arrdiv32_mux2to1124_and0;
  wire f_arrdiv32_mux2to1124_not0;
  wire f_arrdiv32_mux2to1124_and1;
  wire f_arrdiv32_mux2to1124_xor0;
  wire f_arrdiv32_mux2to1125_and0;
  wire f_arrdiv32_mux2to1125_not0;
  wire f_arrdiv32_mux2to1125_and1;
  wire f_arrdiv32_mux2to1125_xor0;
  wire f_arrdiv32_mux2to1126_and0;
  wire f_arrdiv32_mux2to1126_not0;
  wire f_arrdiv32_mux2to1126_and1;
  wire f_arrdiv32_mux2to1126_xor0;
  wire f_arrdiv32_mux2to1127_and0;
  wire f_arrdiv32_mux2to1127_not0;
  wire f_arrdiv32_mux2to1127_and1;
  wire f_arrdiv32_mux2to1127_xor0;
  wire f_arrdiv32_mux2to1128_and0;
  wire f_arrdiv32_mux2to1128_not0;
  wire f_arrdiv32_mux2to1128_and1;
  wire f_arrdiv32_mux2to1128_xor0;
  wire f_arrdiv32_mux2to1129_and0;
  wire f_arrdiv32_mux2to1129_not0;
  wire f_arrdiv32_mux2to1129_and1;
  wire f_arrdiv32_mux2to1129_xor0;
  wire f_arrdiv32_mux2to1130_and0;
  wire f_arrdiv32_mux2to1130_not0;
  wire f_arrdiv32_mux2to1130_and1;
  wire f_arrdiv32_mux2to1130_xor0;
  wire f_arrdiv32_mux2to1131_and0;
  wire f_arrdiv32_mux2to1131_not0;
  wire f_arrdiv32_mux2to1131_and1;
  wire f_arrdiv32_mux2to1131_xor0;
  wire f_arrdiv32_mux2to1132_and0;
  wire f_arrdiv32_mux2to1132_not0;
  wire f_arrdiv32_mux2to1132_and1;
  wire f_arrdiv32_mux2to1132_xor0;
  wire f_arrdiv32_mux2to1133_and0;
  wire f_arrdiv32_mux2to1133_not0;
  wire f_arrdiv32_mux2to1133_and1;
  wire f_arrdiv32_mux2to1133_xor0;
  wire f_arrdiv32_mux2to1134_and0;
  wire f_arrdiv32_mux2to1134_not0;
  wire f_arrdiv32_mux2to1134_and1;
  wire f_arrdiv32_mux2to1134_xor0;
  wire f_arrdiv32_mux2to1135_and0;
  wire f_arrdiv32_mux2to1135_not0;
  wire f_arrdiv32_mux2to1135_and1;
  wire f_arrdiv32_mux2to1135_xor0;
  wire f_arrdiv32_mux2to1136_and0;
  wire f_arrdiv32_mux2to1136_not0;
  wire f_arrdiv32_mux2to1136_and1;
  wire f_arrdiv32_mux2to1136_xor0;
  wire f_arrdiv32_mux2to1137_and0;
  wire f_arrdiv32_mux2to1137_not0;
  wire f_arrdiv32_mux2to1137_and1;
  wire f_arrdiv32_mux2to1137_xor0;
  wire f_arrdiv32_mux2to1138_and0;
  wire f_arrdiv32_mux2to1138_not0;
  wire f_arrdiv32_mux2to1138_and1;
  wire f_arrdiv32_mux2to1138_xor0;
  wire f_arrdiv32_mux2to1139_and0;
  wire f_arrdiv32_mux2to1139_not0;
  wire f_arrdiv32_mux2to1139_and1;
  wire f_arrdiv32_mux2to1139_xor0;
  wire f_arrdiv32_mux2to1140_and0;
  wire f_arrdiv32_mux2to1140_not0;
  wire f_arrdiv32_mux2to1140_and1;
  wire f_arrdiv32_mux2to1140_xor0;
  wire f_arrdiv32_mux2to1141_and0;
  wire f_arrdiv32_mux2to1141_not0;
  wire f_arrdiv32_mux2to1141_and1;
  wire f_arrdiv32_mux2to1141_xor0;
  wire f_arrdiv32_mux2to1142_and0;
  wire f_arrdiv32_mux2to1142_not0;
  wire f_arrdiv32_mux2to1142_and1;
  wire f_arrdiv32_mux2to1142_xor0;
  wire f_arrdiv32_mux2to1143_and0;
  wire f_arrdiv32_mux2to1143_not0;
  wire f_arrdiv32_mux2to1143_and1;
  wire f_arrdiv32_mux2to1143_xor0;
  wire f_arrdiv32_mux2to1144_and0;
  wire f_arrdiv32_mux2to1144_not0;
  wire f_arrdiv32_mux2to1144_and1;
  wire f_arrdiv32_mux2to1144_xor0;
  wire f_arrdiv32_mux2to1145_and0;
  wire f_arrdiv32_mux2to1145_not0;
  wire f_arrdiv32_mux2to1145_and1;
  wire f_arrdiv32_mux2to1145_xor0;
  wire f_arrdiv32_mux2to1146_and0;
  wire f_arrdiv32_mux2to1146_not0;
  wire f_arrdiv32_mux2to1146_and1;
  wire f_arrdiv32_mux2to1146_xor0;
  wire f_arrdiv32_mux2to1147_and0;
  wire f_arrdiv32_mux2to1147_not0;
  wire f_arrdiv32_mux2to1147_and1;
  wire f_arrdiv32_mux2to1147_xor0;
  wire f_arrdiv32_mux2to1148_and0;
  wire f_arrdiv32_mux2to1148_not0;
  wire f_arrdiv32_mux2to1148_and1;
  wire f_arrdiv32_mux2to1148_xor0;
  wire f_arrdiv32_mux2to1149_and0;
  wire f_arrdiv32_mux2to1149_not0;
  wire f_arrdiv32_mux2to1149_and1;
  wire f_arrdiv32_mux2to1149_xor0;
  wire f_arrdiv32_mux2to1150_and0;
  wire f_arrdiv32_mux2to1150_not0;
  wire f_arrdiv32_mux2to1150_and1;
  wire f_arrdiv32_mux2to1150_xor0;
  wire f_arrdiv32_mux2to1151_and0;
  wire f_arrdiv32_mux2to1151_not0;
  wire f_arrdiv32_mux2to1151_and1;
  wire f_arrdiv32_mux2to1151_xor0;
  wire f_arrdiv32_mux2to1152_and0;
  wire f_arrdiv32_mux2to1152_not0;
  wire f_arrdiv32_mux2to1152_and1;
  wire f_arrdiv32_mux2to1152_xor0;
  wire f_arrdiv32_mux2to1153_and0;
  wire f_arrdiv32_mux2to1153_not0;
  wire f_arrdiv32_mux2to1153_and1;
  wire f_arrdiv32_mux2to1153_xor0;
  wire f_arrdiv32_mux2to1154_and0;
  wire f_arrdiv32_mux2to1154_not0;
  wire f_arrdiv32_mux2to1154_and1;
  wire f_arrdiv32_mux2to1154_xor0;
  wire f_arrdiv32_not4;
  wire f_arrdiv32_fs160_xor0;
  wire f_arrdiv32_fs160_not0;
  wire f_arrdiv32_fs160_and0;
  wire f_arrdiv32_fs160_not1;
  wire f_arrdiv32_fs161_xor0;
  wire f_arrdiv32_fs161_not0;
  wire f_arrdiv32_fs161_and0;
  wire f_arrdiv32_fs161_xor1;
  wire f_arrdiv32_fs161_not1;
  wire f_arrdiv32_fs161_and1;
  wire f_arrdiv32_fs161_or0;
  wire f_arrdiv32_fs162_xor0;
  wire f_arrdiv32_fs162_not0;
  wire f_arrdiv32_fs162_and0;
  wire f_arrdiv32_fs162_xor1;
  wire f_arrdiv32_fs162_not1;
  wire f_arrdiv32_fs162_and1;
  wire f_arrdiv32_fs162_or0;
  wire f_arrdiv32_fs163_xor0;
  wire f_arrdiv32_fs163_not0;
  wire f_arrdiv32_fs163_and0;
  wire f_arrdiv32_fs163_xor1;
  wire f_arrdiv32_fs163_not1;
  wire f_arrdiv32_fs163_and1;
  wire f_arrdiv32_fs163_or0;
  wire f_arrdiv32_fs164_xor0;
  wire f_arrdiv32_fs164_not0;
  wire f_arrdiv32_fs164_and0;
  wire f_arrdiv32_fs164_xor1;
  wire f_arrdiv32_fs164_not1;
  wire f_arrdiv32_fs164_and1;
  wire f_arrdiv32_fs164_or0;
  wire f_arrdiv32_fs165_xor0;
  wire f_arrdiv32_fs165_not0;
  wire f_arrdiv32_fs165_and0;
  wire f_arrdiv32_fs165_xor1;
  wire f_arrdiv32_fs165_not1;
  wire f_arrdiv32_fs165_and1;
  wire f_arrdiv32_fs165_or0;
  wire f_arrdiv32_fs166_xor0;
  wire f_arrdiv32_fs166_not0;
  wire f_arrdiv32_fs166_and0;
  wire f_arrdiv32_fs166_xor1;
  wire f_arrdiv32_fs166_not1;
  wire f_arrdiv32_fs166_and1;
  wire f_arrdiv32_fs166_or0;
  wire f_arrdiv32_fs167_xor0;
  wire f_arrdiv32_fs167_not0;
  wire f_arrdiv32_fs167_and0;
  wire f_arrdiv32_fs167_xor1;
  wire f_arrdiv32_fs167_not1;
  wire f_arrdiv32_fs167_and1;
  wire f_arrdiv32_fs167_or0;
  wire f_arrdiv32_fs168_xor0;
  wire f_arrdiv32_fs168_not0;
  wire f_arrdiv32_fs168_and0;
  wire f_arrdiv32_fs168_xor1;
  wire f_arrdiv32_fs168_not1;
  wire f_arrdiv32_fs168_and1;
  wire f_arrdiv32_fs168_or0;
  wire f_arrdiv32_fs169_xor0;
  wire f_arrdiv32_fs169_not0;
  wire f_arrdiv32_fs169_and0;
  wire f_arrdiv32_fs169_xor1;
  wire f_arrdiv32_fs169_not1;
  wire f_arrdiv32_fs169_and1;
  wire f_arrdiv32_fs169_or0;
  wire f_arrdiv32_fs170_xor0;
  wire f_arrdiv32_fs170_not0;
  wire f_arrdiv32_fs170_and0;
  wire f_arrdiv32_fs170_xor1;
  wire f_arrdiv32_fs170_not1;
  wire f_arrdiv32_fs170_and1;
  wire f_arrdiv32_fs170_or0;
  wire f_arrdiv32_fs171_xor0;
  wire f_arrdiv32_fs171_not0;
  wire f_arrdiv32_fs171_and0;
  wire f_arrdiv32_fs171_xor1;
  wire f_arrdiv32_fs171_not1;
  wire f_arrdiv32_fs171_and1;
  wire f_arrdiv32_fs171_or0;
  wire f_arrdiv32_fs172_xor0;
  wire f_arrdiv32_fs172_not0;
  wire f_arrdiv32_fs172_and0;
  wire f_arrdiv32_fs172_xor1;
  wire f_arrdiv32_fs172_not1;
  wire f_arrdiv32_fs172_and1;
  wire f_arrdiv32_fs172_or0;
  wire f_arrdiv32_fs173_xor0;
  wire f_arrdiv32_fs173_not0;
  wire f_arrdiv32_fs173_and0;
  wire f_arrdiv32_fs173_xor1;
  wire f_arrdiv32_fs173_not1;
  wire f_arrdiv32_fs173_and1;
  wire f_arrdiv32_fs173_or0;
  wire f_arrdiv32_fs174_xor0;
  wire f_arrdiv32_fs174_not0;
  wire f_arrdiv32_fs174_and0;
  wire f_arrdiv32_fs174_xor1;
  wire f_arrdiv32_fs174_not1;
  wire f_arrdiv32_fs174_and1;
  wire f_arrdiv32_fs174_or0;
  wire f_arrdiv32_fs175_xor0;
  wire f_arrdiv32_fs175_not0;
  wire f_arrdiv32_fs175_and0;
  wire f_arrdiv32_fs175_xor1;
  wire f_arrdiv32_fs175_not1;
  wire f_arrdiv32_fs175_and1;
  wire f_arrdiv32_fs175_or0;
  wire f_arrdiv32_fs176_xor0;
  wire f_arrdiv32_fs176_not0;
  wire f_arrdiv32_fs176_and0;
  wire f_arrdiv32_fs176_xor1;
  wire f_arrdiv32_fs176_not1;
  wire f_arrdiv32_fs176_and1;
  wire f_arrdiv32_fs176_or0;
  wire f_arrdiv32_fs177_xor0;
  wire f_arrdiv32_fs177_not0;
  wire f_arrdiv32_fs177_and0;
  wire f_arrdiv32_fs177_xor1;
  wire f_arrdiv32_fs177_not1;
  wire f_arrdiv32_fs177_and1;
  wire f_arrdiv32_fs177_or0;
  wire f_arrdiv32_fs178_xor0;
  wire f_arrdiv32_fs178_not0;
  wire f_arrdiv32_fs178_and0;
  wire f_arrdiv32_fs178_xor1;
  wire f_arrdiv32_fs178_not1;
  wire f_arrdiv32_fs178_and1;
  wire f_arrdiv32_fs178_or0;
  wire f_arrdiv32_fs179_xor0;
  wire f_arrdiv32_fs179_not0;
  wire f_arrdiv32_fs179_and0;
  wire f_arrdiv32_fs179_xor1;
  wire f_arrdiv32_fs179_not1;
  wire f_arrdiv32_fs179_and1;
  wire f_arrdiv32_fs179_or0;
  wire f_arrdiv32_fs180_xor0;
  wire f_arrdiv32_fs180_not0;
  wire f_arrdiv32_fs180_and0;
  wire f_arrdiv32_fs180_xor1;
  wire f_arrdiv32_fs180_not1;
  wire f_arrdiv32_fs180_and1;
  wire f_arrdiv32_fs180_or0;
  wire f_arrdiv32_fs181_xor0;
  wire f_arrdiv32_fs181_not0;
  wire f_arrdiv32_fs181_and0;
  wire f_arrdiv32_fs181_xor1;
  wire f_arrdiv32_fs181_not1;
  wire f_arrdiv32_fs181_and1;
  wire f_arrdiv32_fs181_or0;
  wire f_arrdiv32_fs182_xor0;
  wire f_arrdiv32_fs182_not0;
  wire f_arrdiv32_fs182_and0;
  wire f_arrdiv32_fs182_xor1;
  wire f_arrdiv32_fs182_not1;
  wire f_arrdiv32_fs182_and1;
  wire f_arrdiv32_fs182_or0;
  wire f_arrdiv32_fs183_xor0;
  wire f_arrdiv32_fs183_not0;
  wire f_arrdiv32_fs183_and0;
  wire f_arrdiv32_fs183_xor1;
  wire f_arrdiv32_fs183_not1;
  wire f_arrdiv32_fs183_and1;
  wire f_arrdiv32_fs183_or0;
  wire f_arrdiv32_fs184_xor0;
  wire f_arrdiv32_fs184_not0;
  wire f_arrdiv32_fs184_and0;
  wire f_arrdiv32_fs184_xor1;
  wire f_arrdiv32_fs184_not1;
  wire f_arrdiv32_fs184_and1;
  wire f_arrdiv32_fs184_or0;
  wire f_arrdiv32_fs185_xor0;
  wire f_arrdiv32_fs185_not0;
  wire f_arrdiv32_fs185_and0;
  wire f_arrdiv32_fs185_xor1;
  wire f_arrdiv32_fs185_not1;
  wire f_arrdiv32_fs185_and1;
  wire f_arrdiv32_fs185_or0;
  wire f_arrdiv32_fs186_xor0;
  wire f_arrdiv32_fs186_not0;
  wire f_arrdiv32_fs186_and0;
  wire f_arrdiv32_fs186_xor1;
  wire f_arrdiv32_fs186_not1;
  wire f_arrdiv32_fs186_and1;
  wire f_arrdiv32_fs186_or0;
  wire f_arrdiv32_fs187_xor0;
  wire f_arrdiv32_fs187_not0;
  wire f_arrdiv32_fs187_and0;
  wire f_arrdiv32_fs187_xor1;
  wire f_arrdiv32_fs187_not1;
  wire f_arrdiv32_fs187_and1;
  wire f_arrdiv32_fs187_or0;
  wire f_arrdiv32_fs188_xor0;
  wire f_arrdiv32_fs188_not0;
  wire f_arrdiv32_fs188_and0;
  wire f_arrdiv32_fs188_xor1;
  wire f_arrdiv32_fs188_not1;
  wire f_arrdiv32_fs188_and1;
  wire f_arrdiv32_fs188_or0;
  wire f_arrdiv32_fs189_xor0;
  wire f_arrdiv32_fs189_not0;
  wire f_arrdiv32_fs189_and0;
  wire f_arrdiv32_fs189_xor1;
  wire f_arrdiv32_fs189_not1;
  wire f_arrdiv32_fs189_and1;
  wire f_arrdiv32_fs189_or0;
  wire f_arrdiv32_fs190_xor0;
  wire f_arrdiv32_fs190_not0;
  wire f_arrdiv32_fs190_and0;
  wire f_arrdiv32_fs190_xor1;
  wire f_arrdiv32_fs190_not1;
  wire f_arrdiv32_fs190_and1;
  wire f_arrdiv32_fs190_or0;
  wire f_arrdiv32_fs191_xor0;
  wire f_arrdiv32_fs191_not0;
  wire f_arrdiv32_fs191_and0;
  wire f_arrdiv32_fs191_xor1;
  wire f_arrdiv32_fs191_not1;
  wire f_arrdiv32_fs191_and1;
  wire f_arrdiv32_fs191_or0;
  wire f_arrdiv32_mux2to1155_and0;
  wire f_arrdiv32_mux2to1155_not0;
  wire f_arrdiv32_mux2to1155_and1;
  wire f_arrdiv32_mux2to1155_xor0;
  wire f_arrdiv32_mux2to1156_and0;
  wire f_arrdiv32_mux2to1156_not0;
  wire f_arrdiv32_mux2to1156_and1;
  wire f_arrdiv32_mux2to1156_xor0;
  wire f_arrdiv32_mux2to1157_and0;
  wire f_arrdiv32_mux2to1157_not0;
  wire f_arrdiv32_mux2to1157_and1;
  wire f_arrdiv32_mux2to1157_xor0;
  wire f_arrdiv32_mux2to1158_and0;
  wire f_arrdiv32_mux2to1158_not0;
  wire f_arrdiv32_mux2to1158_and1;
  wire f_arrdiv32_mux2to1158_xor0;
  wire f_arrdiv32_mux2to1159_and0;
  wire f_arrdiv32_mux2to1159_not0;
  wire f_arrdiv32_mux2to1159_and1;
  wire f_arrdiv32_mux2to1159_xor0;
  wire f_arrdiv32_mux2to1160_and0;
  wire f_arrdiv32_mux2to1160_not0;
  wire f_arrdiv32_mux2to1160_and1;
  wire f_arrdiv32_mux2to1160_xor0;
  wire f_arrdiv32_mux2to1161_and0;
  wire f_arrdiv32_mux2to1161_not0;
  wire f_arrdiv32_mux2to1161_and1;
  wire f_arrdiv32_mux2to1161_xor0;
  wire f_arrdiv32_mux2to1162_and0;
  wire f_arrdiv32_mux2to1162_not0;
  wire f_arrdiv32_mux2to1162_and1;
  wire f_arrdiv32_mux2to1162_xor0;
  wire f_arrdiv32_mux2to1163_and0;
  wire f_arrdiv32_mux2to1163_not0;
  wire f_arrdiv32_mux2to1163_and1;
  wire f_arrdiv32_mux2to1163_xor0;
  wire f_arrdiv32_mux2to1164_and0;
  wire f_arrdiv32_mux2to1164_not0;
  wire f_arrdiv32_mux2to1164_and1;
  wire f_arrdiv32_mux2to1164_xor0;
  wire f_arrdiv32_mux2to1165_and0;
  wire f_arrdiv32_mux2to1165_not0;
  wire f_arrdiv32_mux2to1165_and1;
  wire f_arrdiv32_mux2to1165_xor0;
  wire f_arrdiv32_mux2to1166_and0;
  wire f_arrdiv32_mux2to1166_not0;
  wire f_arrdiv32_mux2to1166_and1;
  wire f_arrdiv32_mux2to1166_xor0;
  wire f_arrdiv32_mux2to1167_and0;
  wire f_arrdiv32_mux2to1167_not0;
  wire f_arrdiv32_mux2to1167_and1;
  wire f_arrdiv32_mux2to1167_xor0;
  wire f_arrdiv32_mux2to1168_and0;
  wire f_arrdiv32_mux2to1168_not0;
  wire f_arrdiv32_mux2to1168_and1;
  wire f_arrdiv32_mux2to1168_xor0;
  wire f_arrdiv32_mux2to1169_and0;
  wire f_arrdiv32_mux2to1169_not0;
  wire f_arrdiv32_mux2to1169_and1;
  wire f_arrdiv32_mux2to1169_xor0;
  wire f_arrdiv32_mux2to1170_and0;
  wire f_arrdiv32_mux2to1170_not0;
  wire f_arrdiv32_mux2to1170_and1;
  wire f_arrdiv32_mux2to1170_xor0;
  wire f_arrdiv32_mux2to1171_and0;
  wire f_arrdiv32_mux2to1171_not0;
  wire f_arrdiv32_mux2to1171_and1;
  wire f_arrdiv32_mux2to1171_xor0;
  wire f_arrdiv32_mux2to1172_and0;
  wire f_arrdiv32_mux2to1172_not0;
  wire f_arrdiv32_mux2to1172_and1;
  wire f_arrdiv32_mux2to1172_xor0;
  wire f_arrdiv32_mux2to1173_and0;
  wire f_arrdiv32_mux2to1173_not0;
  wire f_arrdiv32_mux2to1173_and1;
  wire f_arrdiv32_mux2to1173_xor0;
  wire f_arrdiv32_mux2to1174_and0;
  wire f_arrdiv32_mux2to1174_not0;
  wire f_arrdiv32_mux2to1174_and1;
  wire f_arrdiv32_mux2to1174_xor0;
  wire f_arrdiv32_mux2to1175_and0;
  wire f_arrdiv32_mux2to1175_not0;
  wire f_arrdiv32_mux2to1175_and1;
  wire f_arrdiv32_mux2to1175_xor0;
  wire f_arrdiv32_mux2to1176_and0;
  wire f_arrdiv32_mux2to1176_not0;
  wire f_arrdiv32_mux2to1176_and1;
  wire f_arrdiv32_mux2to1176_xor0;
  wire f_arrdiv32_mux2to1177_and0;
  wire f_arrdiv32_mux2to1177_not0;
  wire f_arrdiv32_mux2to1177_and1;
  wire f_arrdiv32_mux2to1177_xor0;
  wire f_arrdiv32_mux2to1178_and0;
  wire f_arrdiv32_mux2to1178_not0;
  wire f_arrdiv32_mux2to1178_and1;
  wire f_arrdiv32_mux2to1178_xor0;
  wire f_arrdiv32_mux2to1179_and0;
  wire f_arrdiv32_mux2to1179_not0;
  wire f_arrdiv32_mux2to1179_and1;
  wire f_arrdiv32_mux2to1179_xor0;
  wire f_arrdiv32_mux2to1180_and0;
  wire f_arrdiv32_mux2to1180_not0;
  wire f_arrdiv32_mux2to1180_and1;
  wire f_arrdiv32_mux2to1180_xor0;
  wire f_arrdiv32_mux2to1181_and0;
  wire f_arrdiv32_mux2to1181_not0;
  wire f_arrdiv32_mux2to1181_and1;
  wire f_arrdiv32_mux2to1181_xor0;
  wire f_arrdiv32_mux2to1182_and0;
  wire f_arrdiv32_mux2to1182_not0;
  wire f_arrdiv32_mux2to1182_and1;
  wire f_arrdiv32_mux2to1182_xor0;
  wire f_arrdiv32_mux2to1183_and0;
  wire f_arrdiv32_mux2to1183_not0;
  wire f_arrdiv32_mux2to1183_and1;
  wire f_arrdiv32_mux2to1183_xor0;
  wire f_arrdiv32_mux2to1184_and0;
  wire f_arrdiv32_mux2to1184_not0;
  wire f_arrdiv32_mux2to1184_and1;
  wire f_arrdiv32_mux2to1184_xor0;
  wire f_arrdiv32_mux2to1185_and0;
  wire f_arrdiv32_mux2to1185_not0;
  wire f_arrdiv32_mux2to1185_and1;
  wire f_arrdiv32_mux2to1185_xor0;
  wire f_arrdiv32_not5;
  wire f_arrdiv32_fs192_xor0;
  wire f_arrdiv32_fs192_not0;
  wire f_arrdiv32_fs192_and0;
  wire f_arrdiv32_fs192_not1;
  wire f_arrdiv32_fs193_xor0;
  wire f_arrdiv32_fs193_not0;
  wire f_arrdiv32_fs193_and0;
  wire f_arrdiv32_fs193_xor1;
  wire f_arrdiv32_fs193_not1;
  wire f_arrdiv32_fs193_and1;
  wire f_arrdiv32_fs193_or0;
  wire f_arrdiv32_fs194_xor0;
  wire f_arrdiv32_fs194_not0;
  wire f_arrdiv32_fs194_and0;
  wire f_arrdiv32_fs194_xor1;
  wire f_arrdiv32_fs194_not1;
  wire f_arrdiv32_fs194_and1;
  wire f_arrdiv32_fs194_or0;
  wire f_arrdiv32_fs195_xor0;
  wire f_arrdiv32_fs195_not0;
  wire f_arrdiv32_fs195_and0;
  wire f_arrdiv32_fs195_xor1;
  wire f_arrdiv32_fs195_not1;
  wire f_arrdiv32_fs195_and1;
  wire f_arrdiv32_fs195_or0;
  wire f_arrdiv32_fs196_xor0;
  wire f_arrdiv32_fs196_not0;
  wire f_arrdiv32_fs196_and0;
  wire f_arrdiv32_fs196_xor1;
  wire f_arrdiv32_fs196_not1;
  wire f_arrdiv32_fs196_and1;
  wire f_arrdiv32_fs196_or0;
  wire f_arrdiv32_fs197_xor0;
  wire f_arrdiv32_fs197_not0;
  wire f_arrdiv32_fs197_and0;
  wire f_arrdiv32_fs197_xor1;
  wire f_arrdiv32_fs197_not1;
  wire f_arrdiv32_fs197_and1;
  wire f_arrdiv32_fs197_or0;
  wire f_arrdiv32_fs198_xor0;
  wire f_arrdiv32_fs198_not0;
  wire f_arrdiv32_fs198_and0;
  wire f_arrdiv32_fs198_xor1;
  wire f_arrdiv32_fs198_not1;
  wire f_arrdiv32_fs198_and1;
  wire f_arrdiv32_fs198_or0;
  wire f_arrdiv32_fs199_xor0;
  wire f_arrdiv32_fs199_not0;
  wire f_arrdiv32_fs199_and0;
  wire f_arrdiv32_fs199_xor1;
  wire f_arrdiv32_fs199_not1;
  wire f_arrdiv32_fs199_and1;
  wire f_arrdiv32_fs199_or0;
  wire f_arrdiv32_fs200_xor0;
  wire f_arrdiv32_fs200_not0;
  wire f_arrdiv32_fs200_and0;
  wire f_arrdiv32_fs200_xor1;
  wire f_arrdiv32_fs200_not1;
  wire f_arrdiv32_fs200_and1;
  wire f_arrdiv32_fs200_or0;
  wire f_arrdiv32_fs201_xor0;
  wire f_arrdiv32_fs201_not0;
  wire f_arrdiv32_fs201_and0;
  wire f_arrdiv32_fs201_xor1;
  wire f_arrdiv32_fs201_not1;
  wire f_arrdiv32_fs201_and1;
  wire f_arrdiv32_fs201_or0;
  wire f_arrdiv32_fs202_xor0;
  wire f_arrdiv32_fs202_not0;
  wire f_arrdiv32_fs202_and0;
  wire f_arrdiv32_fs202_xor1;
  wire f_arrdiv32_fs202_not1;
  wire f_arrdiv32_fs202_and1;
  wire f_arrdiv32_fs202_or0;
  wire f_arrdiv32_fs203_xor0;
  wire f_arrdiv32_fs203_not0;
  wire f_arrdiv32_fs203_and0;
  wire f_arrdiv32_fs203_xor1;
  wire f_arrdiv32_fs203_not1;
  wire f_arrdiv32_fs203_and1;
  wire f_arrdiv32_fs203_or0;
  wire f_arrdiv32_fs204_xor0;
  wire f_arrdiv32_fs204_not0;
  wire f_arrdiv32_fs204_and0;
  wire f_arrdiv32_fs204_xor1;
  wire f_arrdiv32_fs204_not1;
  wire f_arrdiv32_fs204_and1;
  wire f_arrdiv32_fs204_or0;
  wire f_arrdiv32_fs205_xor0;
  wire f_arrdiv32_fs205_not0;
  wire f_arrdiv32_fs205_and0;
  wire f_arrdiv32_fs205_xor1;
  wire f_arrdiv32_fs205_not1;
  wire f_arrdiv32_fs205_and1;
  wire f_arrdiv32_fs205_or0;
  wire f_arrdiv32_fs206_xor0;
  wire f_arrdiv32_fs206_not0;
  wire f_arrdiv32_fs206_and0;
  wire f_arrdiv32_fs206_xor1;
  wire f_arrdiv32_fs206_not1;
  wire f_arrdiv32_fs206_and1;
  wire f_arrdiv32_fs206_or0;
  wire f_arrdiv32_fs207_xor0;
  wire f_arrdiv32_fs207_not0;
  wire f_arrdiv32_fs207_and0;
  wire f_arrdiv32_fs207_xor1;
  wire f_arrdiv32_fs207_not1;
  wire f_arrdiv32_fs207_and1;
  wire f_arrdiv32_fs207_or0;
  wire f_arrdiv32_fs208_xor0;
  wire f_arrdiv32_fs208_not0;
  wire f_arrdiv32_fs208_and0;
  wire f_arrdiv32_fs208_xor1;
  wire f_arrdiv32_fs208_not1;
  wire f_arrdiv32_fs208_and1;
  wire f_arrdiv32_fs208_or0;
  wire f_arrdiv32_fs209_xor0;
  wire f_arrdiv32_fs209_not0;
  wire f_arrdiv32_fs209_and0;
  wire f_arrdiv32_fs209_xor1;
  wire f_arrdiv32_fs209_not1;
  wire f_arrdiv32_fs209_and1;
  wire f_arrdiv32_fs209_or0;
  wire f_arrdiv32_fs210_xor0;
  wire f_arrdiv32_fs210_not0;
  wire f_arrdiv32_fs210_and0;
  wire f_arrdiv32_fs210_xor1;
  wire f_arrdiv32_fs210_not1;
  wire f_arrdiv32_fs210_and1;
  wire f_arrdiv32_fs210_or0;
  wire f_arrdiv32_fs211_xor0;
  wire f_arrdiv32_fs211_not0;
  wire f_arrdiv32_fs211_and0;
  wire f_arrdiv32_fs211_xor1;
  wire f_arrdiv32_fs211_not1;
  wire f_arrdiv32_fs211_and1;
  wire f_arrdiv32_fs211_or0;
  wire f_arrdiv32_fs212_xor0;
  wire f_arrdiv32_fs212_not0;
  wire f_arrdiv32_fs212_and0;
  wire f_arrdiv32_fs212_xor1;
  wire f_arrdiv32_fs212_not1;
  wire f_arrdiv32_fs212_and1;
  wire f_arrdiv32_fs212_or0;
  wire f_arrdiv32_fs213_xor0;
  wire f_arrdiv32_fs213_not0;
  wire f_arrdiv32_fs213_and0;
  wire f_arrdiv32_fs213_xor1;
  wire f_arrdiv32_fs213_not1;
  wire f_arrdiv32_fs213_and1;
  wire f_arrdiv32_fs213_or0;
  wire f_arrdiv32_fs214_xor0;
  wire f_arrdiv32_fs214_not0;
  wire f_arrdiv32_fs214_and0;
  wire f_arrdiv32_fs214_xor1;
  wire f_arrdiv32_fs214_not1;
  wire f_arrdiv32_fs214_and1;
  wire f_arrdiv32_fs214_or0;
  wire f_arrdiv32_fs215_xor0;
  wire f_arrdiv32_fs215_not0;
  wire f_arrdiv32_fs215_and0;
  wire f_arrdiv32_fs215_xor1;
  wire f_arrdiv32_fs215_not1;
  wire f_arrdiv32_fs215_and1;
  wire f_arrdiv32_fs215_or0;
  wire f_arrdiv32_fs216_xor0;
  wire f_arrdiv32_fs216_not0;
  wire f_arrdiv32_fs216_and0;
  wire f_arrdiv32_fs216_xor1;
  wire f_arrdiv32_fs216_not1;
  wire f_arrdiv32_fs216_and1;
  wire f_arrdiv32_fs216_or0;
  wire f_arrdiv32_fs217_xor0;
  wire f_arrdiv32_fs217_not0;
  wire f_arrdiv32_fs217_and0;
  wire f_arrdiv32_fs217_xor1;
  wire f_arrdiv32_fs217_not1;
  wire f_arrdiv32_fs217_and1;
  wire f_arrdiv32_fs217_or0;
  wire f_arrdiv32_fs218_xor0;
  wire f_arrdiv32_fs218_not0;
  wire f_arrdiv32_fs218_and0;
  wire f_arrdiv32_fs218_xor1;
  wire f_arrdiv32_fs218_not1;
  wire f_arrdiv32_fs218_and1;
  wire f_arrdiv32_fs218_or0;
  wire f_arrdiv32_fs219_xor0;
  wire f_arrdiv32_fs219_not0;
  wire f_arrdiv32_fs219_and0;
  wire f_arrdiv32_fs219_xor1;
  wire f_arrdiv32_fs219_not1;
  wire f_arrdiv32_fs219_and1;
  wire f_arrdiv32_fs219_or0;
  wire f_arrdiv32_fs220_xor0;
  wire f_arrdiv32_fs220_not0;
  wire f_arrdiv32_fs220_and0;
  wire f_arrdiv32_fs220_xor1;
  wire f_arrdiv32_fs220_not1;
  wire f_arrdiv32_fs220_and1;
  wire f_arrdiv32_fs220_or0;
  wire f_arrdiv32_fs221_xor0;
  wire f_arrdiv32_fs221_not0;
  wire f_arrdiv32_fs221_and0;
  wire f_arrdiv32_fs221_xor1;
  wire f_arrdiv32_fs221_not1;
  wire f_arrdiv32_fs221_and1;
  wire f_arrdiv32_fs221_or0;
  wire f_arrdiv32_fs222_xor0;
  wire f_arrdiv32_fs222_not0;
  wire f_arrdiv32_fs222_and0;
  wire f_arrdiv32_fs222_xor1;
  wire f_arrdiv32_fs222_not1;
  wire f_arrdiv32_fs222_and1;
  wire f_arrdiv32_fs222_or0;
  wire f_arrdiv32_fs223_xor0;
  wire f_arrdiv32_fs223_not0;
  wire f_arrdiv32_fs223_and0;
  wire f_arrdiv32_fs223_xor1;
  wire f_arrdiv32_fs223_not1;
  wire f_arrdiv32_fs223_and1;
  wire f_arrdiv32_fs223_or0;
  wire f_arrdiv32_mux2to1186_and0;
  wire f_arrdiv32_mux2to1186_not0;
  wire f_arrdiv32_mux2to1186_and1;
  wire f_arrdiv32_mux2to1186_xor0;
  wire f_arrdiv32_mux2to1187_and0;
  wire f_arrdiv32_mux2to1187_not0;
  wire f_arrdiv32_mux2to1187_and1;
  wire f_arrdiv32_mux2to1187_xor0;
  wire f_arrdiv32_mux2to1188_and0;
  wire f_arrdiv32_mux2to1188_not0;
  wire f_arrdiv32_mux2to1188_and1;
  wire f_arrdiv32_mux2to1188_xor0;
  wire f_arrdiv32_mux2to1189_and0;
  wire f_arrdiv32_mux2to1189_not0;
  wire f_arrdiv32_mux2to1189_and1;
  wire f_arrdiv32_mux2to1189_xor0;
  wire f_arrdiv32_mux2to1190_and0;
  wire f_arrdiv32_mux2to1190_not0;
  wire f_arrdiv32_mux2to1190_and1;
  wire f_arrdiv32_mux2to1190_xor0;
  wire f_arrdiv32_mux2to1191_and0;
  wire f_arrdiv32_mux2to1191_not0;
  wire f_arrdiv32_mux2to1191_and1;
  wire f_arrdiv32_mux2to1191_xor0;
  wire f_arrdiv32_mux2to1192_and0;
  wire f_arrdiv32_mux2to1192_not0;
  wire f_arrdiv32_mux2to1192_and1;
  wire f_arrdiv32_mux2to1192_xor0;
  wire f_arrdiv32_mux2to1193_and0;
  wire f_arrdiv32_mux2to1193_not0;
  wire f_arrdiv32_mux2to1193_and1;
  wire f_arrdiv32_mux2to1193_xor0;
  wire f_arrdiv32_mux2to1194_and0;
  wire f_arrdiv32_mux2to1194_not0;
  wire f_arrdiv32_mux2to1194_and1;
  wire f_arrdiv32_mux2to1194_xor0;
  wire f_arrdiv32_mux2to1195_and0;
  wire f_arrdiv32_mux2to1195_not0;
  wire f_arrdiv32_mux2to1195_and1;
  wire f_arrdiv32_mux2to1195_xor0;
  wire f_arrdiv32_mux2to1196_and0;
  wire f_arrdiv32_mux2to1196_not0;
  wire f_arrdiv32_mux2to1196_and1;
  wire f_arrdiv32_mux2to1196_xor0;
  wire f_arrdiv32_mux2to1197_and0;
  wire f_arrdiv32_mux2to1197_not0;
  wire f_arrdiv32_mux2to1197_and1;
  wire f_arrdiv32_mux2to1197_xor0;
  wire f_arrdiv32_mux2to1198_and0;
  wire f_arrdiv32_mux2to1198_not0;
  wire f_arrdiv32_mux2to1198_and1;
  wire f_arrdiv32_mux2to1198_xor0;
  wire f_arrdiv32_mux2to1199_and0;
  wire f_arrdiv32_mux2to1199_not0;
  wire f_arrdiv32_mux2to1199_and1;
  wire f_arrdiv32_mux2to1199_xor0;
  wire f_arrdiv32_mux2to1200_and0;
  wire f_arrdiv32_mux2to1200_not0;
  wire f_arrdiv32_mux2to1200_and1;
  wire f_arrdiv32_mux2to1200_xor0;
  wire f_arrdiv32_mux2to1201_and0;
  wire f_arrdiv32_mux2to1201_not0;
  wire f_arrdiv32_mux2to1201_and1;
  wire f_arrdiv32_mux2to1201_xor0;
  wire f_arrdiv32_mux2to1202_and0;
  wire f_arrdiv32_mux2to1202_not0;
  wire f_arrdiv32_mux2to1202_and1;
  wire f_arrdiv32_mux2to1202_xor0;
  wire f_arrdiv32_mux2to1203_and0;
  wire f_arrdiv32_mux2to1203_not0;
  wire f_arrdiv32_mux2to1203_and1;
  wire f_arrdiv32_mux2to1203_xor0;
  wire f_arrdiv32_mux2to1204_and0;
  wire f_arrdiv32_mux2to1204_not0;
  wire f_arrdiv32_mux2to1204_and1;
  wire f_arrdiv32_mux2to1204_xor0;
  wire f_arrdiv32_mux2to1205_and0;
  wire f_arrdiv32_mux2to1205_not0;
  wire f_arrdiv32_mux2to1205_and1;
  wire f_arrdiv32_mux2to1205_xor0;
  wire f_arrdiv32_mux2to1206_and0;
  wire f_arrdiv32_mux2to1206_not0;
  wire f_arrdiv32_mux2to1206_and1;
  wire f_arrdiv32_mux2to1206_xor0;
  wire f_arrdiv32_mux2to1207_and0;
  wire f_arrdiv32_mux2to1207_not0;
  wire f_arrdiv32_mux2to1207_and1;
  wire f_arrdiv32_mux2to1207_xor0;
  wire f_arrdiv32_mux2to1208_and0;
  wire f_arrdiv32_mux2to1208_not0;
  wire f_arrdiv32_mux2to1208_and1;
  wire f_arrdiv32_mux2to1208_xor0;
  wire f_arrdiv32_mux2to1209_and0;
  wire f_arrdiv32_mux2to1209_not0;
  wire f_arrdiv32_mux2to1209_and1;
  wire f_arrdiv32_mux2to1209_xor0;
  wire f_arrdiv32_mux2to1210_and0;
  wire f_arrdiv32_mux2to1210_not0;
  wire f_arrdiv32_mux2to1210_and1;
  wire f_arrdiv32_mux2to1210_xor0;
  wire f_arrdiv32_mux2to1211_and0;
  wire f_arrdiv32_mux2to1211_not0;
  wire f_arrdiv32_mux2to1211_and1;
  wire f_arrdiv32_mux2to1211_xor0;
  wire f_arrdiv32_mux2to1212_and0;
  wire f_arrdiv32_mux2to1212_not0;
  wire f_arrdiv32_mux2to1212_and1;
  wire f_arrdiv32_mux2to1212_xor0;
  wire f_arrdiv32_mux2to1213_and0;
  wire f_arrdiv32_mux2to1213_not0;
  wire f_arrdiv32_mux2to1213_and1;
  wire f_arrdiv32_mux2to1213_xor0;
  wire f_arrdiv32_mux2to1214_and0;
  wire f_arrdiv32_mux2to1214_not0;
  wire f_arrdiv32_mux2to1214_and1;
  wire f_arrdiv32_mux2to1214_xor0;
  wire f_arrdiv32_mux2to1215_and0;
  wire f_arrdiv32_mux2to1215_not0;
  wire f_arrdiv32_mux2to1215_and1;
  wire f_arrdiv32_mux2to1215_xor0;
  wire f_arrdiv32_mux2to1216_and0;
  wire f_arrdiv32_mux2to1216_not0;
  wire f_arrdiv32_mux2to1216_and1;
  wire f_arrdiv32_mux2to1216_xor0;
  wire f_arrdiv32_not6;
  wire f_arrdiv32_fs224_xor0;
  wire f_arrdiv32_fs224_not0;
  wire f_arrdiv32_fs224_and0;
  wire f_arrdiv32_fs224_not1;
  wire f_arrdiv32_fs225_xor0;
  wire f_arrdiv32_fs225_not0;
  wire f_arrdiv32_fs225_and0;
  wire f_arrdiv32_fs225_xor1;
  wire f_arrdiv32_fs225_not1;
  wire f_arrdiv32_fs225_and1;
  wire f_arrdiv32_fs225_or0;
  wire f_arrdiv32_fs226_xor0;
  wire f_arrdiv32_fs226_not0;
  wire f_arrdiv32_fs226_and0;
  wire f_arrdiv32_fs226_xor1;
  wire f_arrdiv32_fs226_not1;
  wire f_arrdiv32_fs226_and1;
  wire f_arrdiv32_fs226_or0;
  wire f_arrdiv32_fs227_xor0;
  wire f_arrdiv32_fs227_not0;
  wire f_arrdiv32_fs227_and0;
  wire f_arrdiv32_fs227_xor1;
  wire f_arrdiv32_fs227_not1;
  wire f_arrdiv32_fs227_and1;
  wire f_arrdiv32_fs227_or0;
  wire f_arrdiv32_fs228_xor0;
  wire f_arrdiv32_fs228_not0;
  wire f_arrdiv32_fs228_and0;
  wire f_arrdiv32_fs228_xor1;
  wire f_arrdiv32_fs228_not1;
  wire f_arrdiv32_fs228_and1;
  wire f_arrdiv32_fs228_or0;
  wire f_arrdiv32_fs229_xor0;
  wire f_arrdiv32_fs229_not0;
  wire f_arrdiv32_fs229_and0;
  wire f_arrdiv32_fs229_xor1;
  wire f_arrdiv32_fs229_not1;
  wire f_arrdiv32_fs229_and1;
  wire f_arrdiv32_fs229_or0;
  wire f_arrdiv32_fs230_xor0;
  wire f_arrdiv32_fs230_not0;
  wire f_arrdiv32_fs230_and0;
  wire f_arrdiv32_fs230_xor1;
  wire f_arrdiv32_fs230_not1;
  wire f_arrdiv32_fs230_and1;
  wire f_arrdiv32_fs230_or0;
  wire f_arrdiv32_fs231_xor0;
  wire f_arrdiv32_fs231_not0;
  wire f_arrdiv32_fs231_and0;
  wire f_arrdiv32_fs231_xor1;
  wire f_arrdiv32_fs231_not1;
  wire f_arrdiv32_fs231_and1;
  wire f_arrdiv32_fs231_or0;
  wire f_arrdiv32_fs232_xor0;
  wire f_arrdiv32_fs232_not0;
  wire f_arrdiv32_fs232_and0;
  wire f_arrdiv32_fs232_xor1;
  wire f_arrdiv32_fs232_not1;
  wire f_arrdiv32_fs232_and1;
  wire f_arrdiv32_fs232_or0;
  wire f_arrdiv32_fs233_xor0;
  wire f_arrdiv32_fs233_not0;
  wire f_arrdiv32_fs233_and0;
  wire f_arrdiv32_fs233_xor1;
  wire f_arrdiv32_fs233_not1;
  wire f_arrdiv32_fs233_and1;
  wire f_arrdiv32_fs233_or0;
  wire f_arrdiv32_fs234_xor0;
  wire f_arrdiv32_fs234_not0;
  wire f_arrdiv32_fs234_and0;
  wire f_arrdiv32_fs234_xor1;
  wire f_arrdiv32_fs234_not1;
  wire f_arrdiv32_fs234_and1;
  wire f_arrdiv32_fs234_or0;
  wire f_arrdiv32_fs235_xor0;
  wire f_arrdiv32_fs235_not0;
  wire f_arrdiv32_fs235_and0;
  wire f_arrdiv32_fs235_xor1;
  wire f_arrdiv32_fs235_not1;
  wire f_arrdiv32_fs235_and1;
  wire f_arrdiv32_fs235_or0;
  wire f_arrdiv32_fs236_xor0;
  wire f_arrdiv32_fs236_not0;
  wire f_arrdiv32_fs236_and0;
  wire f_arrdiv32_fs236_xor1;
  wire f_arrdiv32_fs236_not1;
  wire f_arrdiv32_fs236_and1;
  wire f_arrdiv32_fs236_or0;
  wire f_arrdiv32_fs237_xor0;
  wire f_arrdiv32_fs237_not0;
  wire f_arrdiv32_fs237_and0;
  wire f_arrdiv32_fs237_xor1;
  wire f_arrdiv32_fs237_not1;
  wire f_arrdiv32_fs237_and1;
  wire f_arrdiv32_fs237_or0;
  wire f_arrdiv32_fs238_xor0;
  wire f_arrdiv32_fs238_not0;
  wire f_arrdiv32_fs238_and0;
  wire f_arrdiv32_fs238_xor1;
  wire f_arrdiv32_fs238_not1;
  wire f_arrdiv32_fs238_and1;
  wire f_arrdiv32_fs238_or0;
  wire f_arrdiv32_fs239_xor0;
  wire f_arrdiv32_fs239_not0;
  wire f_arrdiv32_fs239_and0;
  wire f_arrdiv32_fs239_xor1;
  wire f_arrdiv32_fs239_not1;
  wire f_arrdiv32_fs239_and1;
  wire f_arrdiv32_fs239_or0;
  wire f_arrdiv32_fs240_xor0;
  wire f_arrdiv32_fs240_not0;
  wire f_arrdiv32_fs240_and0;
  wire f_arrdiv32_fs240_xor1;
  wire f_arrdiv32_fs240_not1;
  wire f_arrdiv32_fs240_and1;
  wire f_arrdiv32_fs240_or0;
  wire f_arrdiv32_fs241_xor0;
  wire f_arrdiv32_fs241_not0;
  wire f_arrdiv32_fs241_and0;
  wire f_arrdiv32_fs241_xor1;
  wire f_arrdiv32_fs241_not1;
  wire f_arrdiv32_fs241_and1;
  wire f_arrdiv32_fs241_or0;
  wire f_arrdiv32_fs242_xor0;
  wire f_arrdiv32_fs242_not0;
  wire f_arrdiv32_fs242_and0;
  wire f_arrdiv32_fs242_xor1;
  wire f_arrdiv32_fs242_not1;
  wire f_arrdiv32_fs242_and1;
  wire f_arrdiv32_fs242_or0;
  wire f_arrdiv32_fs243_xor0;
  wire f_arrdiv32_fs243_not0;
  wire f_arrdiv32_fs243_and0;
  wire f_arrdiv32_fs243_xor1;
  wire f_arrdiv32_fs243_not1;
  wire f_arrdiv32_fs243_and1;
  wire f_arrdiv32_fs243_or0;
  wire f_arrdiv32_fs244_xor0;
  wire f_arrdiv32_fs244_not0;
  wire f_arrdiv32_fs244_and0;
  wire f_arrdiv32_fs244_xor1;
  wire f_arrdiv32_fs244_not1;
  wire f_arrdiv32_fs244_and1;
  wire f_arrdiv32_fs244_or0;
  wire f_arrdiv32_fs245_xor0;
  wire f_arrdiv32_fs245_not0;
  wire f_arrdiv32_fs245_and0;
  wire f_arrdiv32_fs245_xor1;
  wire f_arrdiv32_fs245_not1;
  wire f_arrdiv32_fs245_and1;
  wire f_arrdiv32_fs245_or0;
  wire f_arrdiv32_fs246_xor0;
  wire f_arrdiv32_fs246_not0;
  wire f_arrdiv32_fs246_and0;
  wire f_arrdiv32_fs246_xor1;
  wire f_arrdiv32_fs246_not1;
  wire f_arrdiv32_fs246_and1;
  wire f_arrdiv32_fs246_or0;
  wire f_arrdiv32_fs247_xor0;
  wire f_arrdiv32_fs247_not0;
  wire f_arrdiv32_fs247_and0;
  wire f_arrdiv32_fs247_xor1;
  wire f_arrdiv32_fs247_not1;
  wire f_arrdiv32_fs247_and1;
  wire f_arrdiv32_fs247_or0;
  wire f_arrdiv32_fs248_xor0;
  wire f_arrdiv32_fs248_not0;
  wire f_arrdiv32_fs248_and0;
  wire f_arrdiv32_fs248_xor1;
  wire f_arrdiv32_fs248_not1;
  wire f_arrdiv32_fs248_and1;
  wire f_arrdiv32_fs248_or0;
  wire f_arrdiv32_fs249_xor0;
  wire f_arrdiv32_fs249_not0;
  wire f_arrdiv32_fs249_and0;
  wire f_arrdiv32_fs249_xor1;
  wire f_arrdiv32_fs249_not1;
  wire f_arrdiv32_fs249_and1;
  wire f_arrdiv32_fs249_or0;
  wire f_arrdiv32_fs250_xor0;
  wire f_arrdiv32_fs250_not0;
  wire f_arrdiv32_fs250_and0;
  wire f_arrdiv32_fs250_xor1;
  wire f_arrdiv32_fs250_not1;
  wire f_arrdiv32_fs250_and1;
  wire f_arrdiv32_fs250_or0;
  wire f_arrdiv32_fs251_xor0;
  wire f_arrdiv32_fs251_not0;
  wire f_arrdiv32_fs251_and0;
  wire f_arrdiv32_fs251_xor1;
  wire f_arrdiv32_fs251_not1;
  wire f_arrdiv32_fs251_and1;
  wire f_arrdiv32_fs251_or0;
  wire f_arrdiv32_fs252_xor0;
  wire f_arrdiv32_fs252_not0;
  wire f_arrdiv32_fs252_and0;
  wire f_arrdiv32_fs252_xor1;
  wire f_arrdiv32_fs252_not1;
  wire f_arrdiv32_fs252_and1;
  wire f_arrdiv32_fs252_or0;
  wire f_arrdiv32_fs253_xor0;
  wire f_arrdiv32_fs253_not0;
  wire f_arrdiv32_fs253_and0;
  wire f_arrdiv32_fs253_xor1;
  wire f_arrdiv32_fs253_not1;
  wire f_arrdiv32_fs253_and1;
  wire f_arrdiv32_fs253_or0;
  wire f_arrdiv32_fs254_xor0;
  wire f_arrdiv32_fs254_not0;
  wire f_arrdiv32_fs254_and0;
  wire f_arrdiv32_fs254_xor1;
  wire f_arrdiv32_fs254_not1;
  wire f_arrdiv32_fs254_and1;
  wire f_arrdiv32_fs254_or0;
  wire f_arrdiv32_fs255_xor0;
  wire f_arrdiv32_fs255_not0;
  wire f_arrdiv32_fs255_and0;
  wire f_arrdiv32_fs255_xor1;
  wire f_arrdiv32_fs255_not1;
  wire f_arrdiv32_fs255_and1;
  wire f_arrdiv32_fs255_or0;
  wire f_arrdiv32_mux2to1217_and0;
  wire f_arrdiv32_mux2to1217_not0;
  wire f_arrdiv32_mux2to1217_and1;
  wire f_arrdiv32_mux2to1217_xor0;
  wire f_arrdiv32_mux2to1218_and0;
  wire f_arrdiv32_mux2to1218_not0;
  wire f_arrdiv32_mux2to1218_and1;
  wire f_arrdiv32_mux2to1218_xor0;
  wire f_arrdiv32_mux2to1219_and0;
  wire f_arrdiv32_mux2to1219_not0;
  wire f_arrdiv32_mux2to1219_and1;
  wire f_arrdiv32_mux2to1219_xor0;
  wire f_arrdiv32_mux2to1220_and0;
  wire f_arrdiv32_mux2to1220_not0;
  wire f_arrdiv32_mux2to1220_and1;
  wire f_arrdiv32_mux2to1220_xor0;
  wire f_arrdiv32_mux2to1221_and0;
  wire f_arrdiv32_mux2to1221_not0;
  wire f_arrdiv32_mux2to1221_and1;
  wire f_arrdiv32_mux2to1221_xor0;
  wire f_arrdiv32_mux2to1222_and0;
  wire f_arrdiv32_mux2to1222_not0;
  wire f_arrdiv32_mux2to1222_and1;
  wire f_arrdiv32_mux2to1222_xor0;
  wire f_arrdiv32_mux2to1223_and0;
  wire f_arrdiv32_mux2to1223_not0;
  wire f_arrdiv32_mux2to1223_and1;
  wire f_arrdiv32_mux2to1223_xor0;
  wire f_arrdiv32_mux2to1224_and0;
  wire f_arrdiv32_mux2to1224_not0;
  wire f_arrdiv32_mux2to1224_and1;
  wire f_arrdiv32_mux2to1224_xor0;
  wire f_arrdiv32_mux2to1225_and0;
  wire f_arrdiv32_mux2to1225_not0;
  wire f_arrdiv32_mux2to1225_and1;
  wire f_arrdiv32_mux2to1225_xor0;
  wire f_arrdiv32_mux2to1226_and0;
  wire f_arrdiv32_mux2to1226_not0;
  wire f_arrdiv32_mux2to1226_and1;
  wire f_arrdiv32_mux2to1226_xor0;
  wire f_arrdiv32_mux2to1227_and0;
  wire f_arrdiv32_mux2to1227_not0;
  wire f_arrdiv32_mux2to1227_and1;
  wire f_arrdiv32_mux2to1227_xor0;
  wire f_arrdiv32_mux2to1228_and0;
  wire f_arrdiv32_mux2to1228_not0;
  wire f_arrdiv32_mux2to1228_and1;
  wire f_arrdiv32_mux2to1228_xor0;
  wire f_arrdiv32_mux2to1229_and0;
  wire f_arrdiv32_mux2to1229_not0;
  wire f_arrdiv32_mux2to1229_and1;
  wire f_arrdiv32_mux2to1229_xor0;
  wire f_arrdiv32_mux2to1230_and0;
  wire f_arrdiv32_mux2to1230_not0;
  wire f_arrdiv32_mux2to1230_and1;
  wire f_arrdiv32_mux2to1230_xor0;
  wire f_arrdiv32_mux2to1231_and0;
  wire f_arrdiv32_mux2to1231_not0;
  wire f_arrdiv32_mux2to1231_and1;
  wire f_arrdiv32_mux2to1231_xor0;
  wire f_arrdiv32_mux2to1232_and0;
  wire f_arrdiv32_mux2to1232_not0;
  wire f_arrdiv32_mux2to1232_and1;
  wire f_arrdiv32_mux2to1232_xor0;
  wire f_arrdiv32_mux2to1233_and0;
  wire f_arrdiv32_mux2to1233_not0;
  wire f_arrdiv32_mux2to1233_and1;
  wire f_arrdiv32_mux2to1233_xor0;
  wire f_arrdiv32_mux2to1234_and0;
  wire f_arrdiv32_mux2to1234_not0;
  wire f_arrdiv32_mux2to1234_and1;
  wire f_arrdiv32_mux2to1234_xor0;
  wire f_arrdiv32_mux2to1235_and0;
  wire f_arrdiv32_mux2to1235_not0;
  wire f_arrdiv32_mux2to1235_and1;
  wire f_arrdiv32_mux2to1235_xor0;
  wire f_arrdiv32_mux2to1236_and0;
  wire f_arrdiv32_mux2to1236_not0;
  wire f_arrdiv32_mux2to1236_and1;
  wire f_arrdiv32_mux2to1236_xor0;
  wire f_arrdiv32_mux2to1237_and0;
  wire f_arrdiv32_mux2to1237_not0;
  wire f_arrdiv32_mux2to1237_and1;
  wire f_arrdiv32_mux2to1237_xor0;
  wire f_arrdiv32_mux2to1238_and0;
  wire f_arrdiv32_mux2to1238_not0;
  wire f_arrdiv32_mux2to1238_and1;
  wire f_arrdiv32_mux2to1238_xor0;
  wire f_arrdiv32_mux2to1239_and0;
  wire f_arrdiv32_mux2to1239_not0;
  wire f_arrdiv32_mux2to1239_and1;
  wire f_arrdiv32_mux2to1239_xor0;
  wire f_arrdiv32_mux2to1240_and0;
  wire f_arrdiv32_mux2to1240_not0;
  wire f_arrdiv32_mux2to1240_and1;
  wire f_arrdiv32_mux2to1240_xor0;
  wire f_arrdiv32_mux2to1241_and0;
  wire f_arrdiv32_mux2to1241_not0;
  wire f_arrdiv32_mux2to1241_and1;
  wire f_arrdiv32_mux2to1241_xor0;
  wire f_arrdiv32_mux2to1242_and0;
  wire f_arrdiv32_mux2to1242_not0;
  wire f_arrdiv32_mux2to1242_and1;
  wire f_arrdiv32_mux2to1242_xor0;
  wire f_arrdiv32_mux2to1243_and0;
  wire f_arrdiv32_mux2to1243_not0;
  wire f_arrdiv32_mux2to1243_and1;
  wire f_arrdiv32_mux2to1243_xor0;
  wire f_arrdiv32_mux2to1244_and0;
  wire f_arrdiv32_mux2to1244_not0;
  wire f_arrdiv32_mux2to1244_and1;
  wire f_arrdiv32_mux2to1244_xor0;
  wire f_arrdiv32_mux2to1245_and0;
  wire f_arrdiv32_mux2to1245_not0;
  wire f_arrdiv32_mux2to1245_and1;
  wire f_arrdiv32_mux2to1245_xor0;
  wire f_arrdiv32_mux2to1246_and0;
  wire f_arrdiv32_mux2to1246_not0;
  wire f_arrdiv32_mux2to1246_and1;
  wire f_arrdiv32_mux2to1246_xor0;
  wire f_arrdiv32_mux2to1247_and0;
  wire f_arrdiv32_mux2to1247_not0;
  wire f_arrdiv32_mux2to1247_and1;
  wire f_arrdiv32_mux2to1247_xor0;
  wire f_arrdiv32_not7;
  wire f_arrdiv32_fs256_xor0;
  wire f_arrdiv32_fs256_not0;
  wire f_arrdiv32_fs256_and0;
  wire f_arrdiv32_fs256_not1;
  wire f_arrdiv32_fs257_xor0;
  wire f_arrdiv32_fs257_not0;
  wire f_arrdiv32_fs257_and0;
  wire f_arrdiv32_fs257_xor1;
  wire f_arrdiv32_fs257_not1;
  wire f_arrdiv32_fs257_and1;
  wire f_arrdiv32_fs257_or0;
  wire f_arrdiv32_fs258_xor0;
  wire f_arrdiv32_fs258_not0;
  wire f_arrdiv32_fs258_and0;
  wire f_arrdiv32_fs258_xor1;
  wire f_arrdiv32_fs258_not1;
  wire f_arrdiv32_fs258_and1;
  wire f_arrdiv32_fs258_or0;
  wire f_arrdiv32_fs259_xor0;
  wire f_arrdiv32_fs259_not0;
  wire f_arrdiv32_fs259_and0;
  wire f_arrdiv32_fs259_xor1;
  wire f_arrdiv32_fs259_not1;
  wire f_arrdiv32_fs259_and1;
  wire f_arrdiv32_fs259_or0;
  wire f_arrdiv32_fs260_xor0;
  wire f_arrdiv32_fs260_not0;
  wire f_arrdiv32_fs260_and0;
  wire f_arrdiv32_fs260_xor1;
  wire f_arrdiv32_fs260_not1;
  wire f_arrdiv32_fs260_and1;
  wire f_arrdiv32_fs260_or0;
  wire f_arrdiv32_fs261_xor0;
  wire f_arrdiv32_fs261_not0;
  wire f_arrdiv32_fs261_and0;
  wire f_arrdiv32_fs261_xor1;
  wire f_arrdiv32_fs261_not1;
  wire f_arrdiv32_fs261_and1;
  wire f_arrdiv32_fs261_or0;
  wire f_arrdiv32_fs262_xor0;
  wire f_arrdiv32_fs262_not0;
  wire f_arrdiv32_fs262_and0;
  wire f_arrdiv32_fs262_xor1;
  wire f_arrdiv32_fs262_not1;
  wire f_arrdiv32_fs262_and1;
  wire f_arrdiv32_fs262_or0;
  wire f_arrdiv32_fs263_xor0;
  wire f_arrdiv32_fs263_not0;
  wire f_arrdiv32_fs263_and0;
  wire f_arrdiv32_fs263_xor1;
  wire f_arrdiv32_fs263_not1;
  wire f_arrdiv32_fs263_and1;
  wire f_arrdiv32_fs263_or0;
  wire f_arrdiv32_fs264_xor0;
  wire f_arrdiv32_fs264_not0;
  wire f_arrdiv32_fs264_and0;
  wire f_arrdiv32_fs264_xor1;
  wire f_arrdiv32_fs264_not1;
  wire f_arrdiv32_fs264_and1;
  wire f_arrdiv32_fs264_or0;
  wire f_arrdiv32_fs265_xor0;
  wire f_arrdiv32_fs265_not0;
  wire f_arrdiv32_fs265_and0;
  wire f_arrdiv32_fs265_xor1;
  wire f_arrdiv32_fs265_not1;
  wire f_arrdiv32_fs265_and1;
  wire f_arrdiv32_fs265_or0;
  wire f_arrdiv32_fs266_xor0;
  wire f_arrdiv32_fs266_not0;
  wire f_arrdiv32_fs266_and0;
  wire f_arrdiv32_fs266_xor1;
  wire f_arrdiv32_fs266_not1;
  wire f_arrdiv32_fs266_and1;
  wire f_arrdiv32_fs266_or0;
  wire f_arrdiv32_fs267_xor0;
  wire f_arrdiv32_fs267_not0;
  wire f_arrdiv32_fs267_and0;
  wire f_arrdiv32_fs267_xor1;
  wire f_arrdiv32_fs267_not1;
  wire f_arrdiv32_fs267_and1;
  wire f_arrdiv32_fs267_or0;
  wire f_arrdiv32_fs268_xor0;
  wire f_arrdiv32_fs268_not0;
  wire f_arrdiv32_fs268_and0;
  wire f_arrdiv32_fs268_xor1;
  wire f_arrdiv32_fs268_not1;
  wire f_arrdiv32_fs268_and1;
  wire f_arrdiv32_fs268_or0;
  wire f_arrdiv32_fs269_xor0;
  wire f_arrdiv32_fs269_not0;
  wire f_arrdiv32_fs269_and0;
  wire f_arrdiv32_fs269_xor1;
  wire f_arrdiv32_fs269_not1;
  wire f_arrdiv32_fs269_and1;
  wire f_arrdiv32_fs269_or0;
  wire f_arrdiv32_fs270_xor0;
  wire f_arrdiv32_fs270_not0;
  wire f_arrdiv32_fs270_and0;
  wire f_arrdiv32_fs270_xor1;
  wire f_arrdiv32_fs270_not1;
  wire f_arrdiv32_fs270_and1;
  wire f_arrdiv32_fs270_or0;
  wire f_arrdiv32_fs271_xor0;
  wire f_arrdiv32_fs271_not0;
  wire f_arrdiv32_fs271_and0;
  wire f_arrdiv32_fs271_xor1;
  wire f_arrdiv32_fs271_not1;
  wire f_arrdiv32_fs271_and1;
  wire f_arrdiv32_fs271_or0;
  wire f_arrdiv32_fs272_xor0;
  wire f_arrdiv32_fs272_not0;
  wire f_arrdiv32_fs272_and0;
  wire f_arrdiv32_fs272_xor1;
  wire f_arrdiv32_fs272_not1;
  wire f_arrdiv32_fs272_and1;
  wire f_arrdiv32_fs272_or0;
  wire f_arrdiv32_fs273_xor0;
  wire f_arrdiv32_fs273_not0;
  wire f_arrdiv32_fs273_and0;
  wire f_arrdiv32_fs273_xor1;
  wire f_arrdiv32_fs273_not1;
  wire f_arrdiv32_fs273_and1;
  wire f_arrdiv32_fs273_or0;
  wire f_arrdiv32_fs274_xor0;
  wire f_arrdiv32_fs274_not0;
  wire f_arrdiv32_fs274_and0;
  wire f_arrdiv32_fs274_xor1;
  wire f_arrdiv32_fs274_not1;
  wire f_arrdiv32_fs274_and1;
  wire f_arrdiv32_fs274_or0;
  wire f_arrdiv32_fs275_xor0;
  wire f_arrdiv32_fs275_not0;
  wire f_arrdiv32_fs275_and0;
  wire f_arrdiv32_fs275_xor1;
  wire f_arrdiv32_fs275_not1;
  wire f_arrdiv32_fs275_and1;
  wire f_arrdiv32_fs275_or0;
  wire f_arrdiv32_fs276_xor0;
  wire f_arrdiv32_fs276_not0;
  wire f_arrdiv32_fs276_and0;
  wire f_arrdiv32_fs276_xor1;
  wire f_arrdiv32_fs276_not1;
  wire f_arrdiv32_fs276_and1;
  wire f_arrdiv32_fs276_or0;
  wire f_arrdiv32_fs277_xor0;
  wire f_arrdiv32_fs277_not0;
  wire f_arrdiv32_fs277_and0;
  wire f_arrdiv32_fs277_xor1;
  wire f_arrdiv32_fs277_not1;
  wire f_arrdiv32_fs277_and1;
  wire f_arrdiv32_fs277_or0;
  wire f_arrdiv32_fs278_xor0;
  wire f_arrdiv32_fs278_not0;
  wire f_arrdiv32_fs278_and0;
  wire f_arrdiv32_fs278_xor1;
  wire f_arrdiv32_fs278_not1;
  wire f_arrdiv32_fs278_and1;
  wire f_arrdiv32_fs278_or0;
  wire f_arrdiv32_fs279_xor0;
  wire f_arrdiv32_fs279_not0;
  wire f_arrdiv32_fs279_and0;
  wire f_arrdiv32_fs279_xor1;
  wire f_arrdiv32_fs279_not1;
  wire f_arrdiv32_fs279_and1;
  wire f_arrdiv32_fs279_or0;
  wire f_arrdiv32_fs280_xor0;
  wire f_arrdiv32_fs280_not0;
  wire f_arrdiv32_fs280_and0;
  wire f_arrdiv32_fs280_xor1;
  wire f_arrdiv32_fs280_not1;
  wire f_arrdiv32_fs280_and1;
  wire f_arrdiv32_fs280_or0;
  wire f_arrdiv32_fs281_xor0;
  wire f_arrdiv32_fs281_not0;
  wire f_arrdiv32_fs281_and0;
  wire f_arrdiv32_fs281_xor1;
  wire f_arrdiv32_fs281_not1;
  wire f_arrdiv32_fs281_and1;
  wire f_arrdiv32_fs281_or0;
  wire f_arrdiv32_fs282_xor0;
  wire f_arrdiv32_fs282_not0;
  wire f_arrdiv32_fs282_and0;
  wire f_arrdiv32_fs282_xor1;
  wire f_arrdiv32_fs282_not1;
  wire f_arrdiv32_fs282_and1;
  wire f_arrdiv32_fs282_or0;
  wire f_arrdiv32_fs283_xor0;
  wire f_arrdiv32_fs283_not0;
  wire f_arrdiv32_fs283_and0;
  wire f_arrdiv32_fs283_xor1;
  wire f_arrdiv32_fs283_not1;
  wire f_arrdiv32_fs283_and1;
  wire f_arrdiv32_fs283_or0;
  wire f_arrdiv32_fs284_xor0;
  wire f_arrdiv32_fs284_not0;
  wire f_arrdiv32_fs284_and0;
  wire f_arrdiv32_fs284_xor1;
  wire f_arrdiv32_fs284_not1;
  wire f_arrdiv32_fs284_and1;
  wire f_arrdiv32_fs284_or0;
  wire f_arrdiv32_fs285_xor0;
  wire f_arrdiv32_fs285_not0;
  wire f_arrdiv32_fs285_and0;
  wire f_arrdiv32_fs285_xor1;
  wire f_arrdiv32_fs285_not1;
  wire f_arrdiv32_fs285_and1;
  wire f_arrdiv32_fs285_or0;
  wire f_arrdiv32_fs286_xor0;
  wire f_arrdiv32_fs286_not0;
  wire f_arrdiv32_fs286_and0;
  wire f_arrdiv32_fs286_xor1;
  wire f_arrdiv32_fs286_not1;
  wire f_arrdiv32_fs286_and1;
  wire f_arrdiv32_fs286_or0;
  wire f_arrdiv32_fs287_xor0;
  wire f_arrdiv32_fs287_not0;
  wire f_arrdiv32_fs287_and0;
  wire f_arrdiv32_fs287_xor1;
  wire f_arrdiv32_fs287_not1;
  wire f_arrdiv32_fs287_and1;
  wire f_arrdiv32_fs287_or0;
  wire f_arrdiv32_mux2to1248_and0;
  wire f_arrdiv32_mux2to1248_not0;
  wire f_arrdiv32_mux2to1248_and1;
  wire f_arrdiv32_mux2to1248_xor0;
  wire f_arrdiv32_mux2to1249_and0;
  wire f_arrdiv32_mux2to1249_not0;
  wire f_arrdiv32_mux2to1249_and1;
  wire f_arrdiv32_mux2to1249_xor0;
  wire f_arrdiv32_mux2to1250_and0;
  wire f_arrdiv32_mux2to1250_not0;
  wire f_arrdiv32_mux2to1250_and1;
  wire f_arrdiv32_mux2to1250_xor0;
  wire f_arrdiv32_mux2to1251_and0;
  wire f_arrdiv32_mux2to1251_not0;
  wire f_arrdiv32_mux2to1251_and1;
  wire f_arrdiv32_mux2to1251_xor0;
  wire f_arrdiv32_mux2to1252_and0;
  wire f_arrdiv32_mux2to1252_not0;
  wire f_arrdiv32_mux2to1252_and1;
  wire f_arrdiv32_mux2to1252_xor0;
  wire f_arrdiv32_mux2to1253_and0;
  wire f_arrdiv32_mux2to1253_not0;
  wire f_arrdiv32_mux2to1253_and1;
  wire f_arrdiv32_mux2to1253_xor0;
  wire f_arrdiv32_mux2to1254_and0;
  wire f_arrdiv32_mux2to1254_not0;
  wire f_arrdiv32_mux2to1254_and1;
  wire f_arrdiv32_mux2to1254_xor0;
  wire f_arrdiv32_mux2to1255_and0;
  wire f_arrdiv32_mux2to1255_not0;
  wire f_arrdiv32_mux2to1255_and1;
  wire f_arrdiv32_mux2to1255_xor0;
  wire f_arrdiv32_mux2to1256_and0;
  wire f_arrdiv32_mux2to1256_not0;
  wire f_arrdiv32_mux2to1256_and1;
  wire f_arrdiv32_mux2to1256_xor0;
  wire f_arrdiv32_mux2to1257_and0;
  wire f_arrdiv32_mux2to1257_not0;
  wire f_arrdiv32_mux2to1257_and1;
  wire f_arrdiv32_mux2to1257_xor0;
  wire f_arrdiv32_mux2to1258_and0;
  wire f_arrdiv32_mux2to1258_not0;
  wire f_arrdiv32_mux2to1258_and1;
  wire f_arrdiv32_mux2to1258_xor0;
  wire f_arrdiv32_mux2to1259_and0;
  wire f_arrdiv32_mux2to1259_not0;
  wire f_arrdiv32_mux2to1259_and1;
  wire f_arrdiv32_mux2to1259_xor0;
  wire f_arrdiv32_mux2to1260_and0;
  wire f_arrdiv32_mux2to1260_not0;
  wire f_arrdiv32_mux2to1260_and1;
  wire f_arrdiv32_mux2to1260_xor0;
  wire f_arrdiv32_mux2to1261_and0;
  wire f_arrdiv32_mux2to1261_not0;
  wire f_arrdiv32_mux2to1261_and1;
  wire f_arrdiv32_mux2to1261_xor0;
  wire f_arrdiv32_mux2to1262_and0;
  wire f_arrdiv32_mux2to1262_not0;
  wire f_arrdiv32_mux2to1262_and1;
  wire f_arrdiv32_mux2to1262_xor0;
  wire f_arrdiv32_mux2to1263_and0;
  wire f_arrdiv32_mux2to1263_not0;
  wire f_arrdiv32_mux2to1263_and1;
  wire f_arrdiv32_mux2to1263_xor0;
  wire f_arrdiv32_mux2to1264_and0;
  wire f_arrdiv32_mux2to1264_not0;
  wire f_arrdiv32_mux2to1264_and1;
  wire f_arrdiv32_mux2to1264_xor0;
  wire f_arrdiv32_mux2to1265_and0;
  wire f_arrdiv32_mux2to1265_not0;
  wire f_arrdiv32_mux2to1265_and1;
  wire f_arrdiv32_mux2to1265_xor0;
  wire f_arrdiv32_mux2to1266_and0;
  wire f_arrdiv32_mux2to1266_not0;
  wire f_arrdiv32_mux2to1266_and1;
  wire f_arrdiv32_mux2to1266_xor0;
  wire f_arrdiv32_mux2to1267_and0;
  wire f_arrdiv32_mux2to1267_not0;
  wire f_arrdiv32_mux2to1267_and1;
  wire f_arrdiv32_mux2to1267_xor0;
  wire f_arrdiv32_mux2to1268_and0;
  wire f_arrdiv32_mux2to1268_not0;
  wire f_arrdiv32_mux2to1268_and1;
  wire f_arrdiv32_mux2to1268_xor0;
  wire f_arrdiv32_mux2to1269_and0;
  wire f_arrdiv32_mux2to1269_not0;
  wire f_arrdiv32_mux2to1269_and1;
  wire f_arrdiv32_mux2to1269_xor0;
  wire f_arrdiv32_mux2to1270_and0;
  wire f_arrdiv32_mux2to1270_not0;
  wire f_arrdiv32_mux2to1270_and1;
  wire f_arrdiv32_mux2to1270_xor0;
  wire f_arrdiv32_mux2to1271_and0;
  wire f_arrdiv32_mux2to1271_not0;
  wire f_arrdiv32_mux2to1271_and1;
  wire f_arrdiv32_mux2to1271_xor0;
  wire f_arrdiv32_mux2to1272_and0;
  wire f_arrdiv32_mux2to1272_not0;
  wire f_arrdiv32_mux2to1272_and1;
  wire f_arrdiv32_mux2to1272_xor0;
  wire f_arrdiv32_mux2to1273_and0;
  wire f_arrdiv32_mux2to1273_not0;
  wire f_arrdiv32_mux2to1273_and1;
  wire f_arrdiv32_mux2to1273_xor0;
  wire f_arrdiv32_mux2to1274_and0;
  wire f_arrdiv32_mux2to1274_not0;
  wire f_arrdiv32_mux2to1274_and1;
  wire f_arrdiv32_mux2to1274_xor0;
  wire f_arrdiv32_mux2to1275_and0;
  wire f_arrdiv32_mux2to1275_not0;
  wire f_arrdiv32_mux2to1275_and1;
  wire f_arrdiv32_mux2to1275_xor0;
  wire f_arrdiv32_mux2to1276_and0;
  wire f_arrdiv32_mux2to1276_not0;
  wire f_arrdiv32_mux2to1276_and1;
  wire f_arrdiv32_mux2to1276_xor0;
  wire f_arrdiv32_mux2to1277_and0;
  wire f_arrdiv32_mux2to1277_not0;
  wire f_arrdiv32_mux2to1277_and1;
  wire f_arrdiv32_mux2to1277_xor0;
  wire f_arrdiv32_mux2to1278_and0;
  wire f_arrdiv32_mux2to1278_not0;
  wire f_arrdiv32_mux2to1278_and1;
  wire f_arrdiv32_mux2to1278_xor0;
  wire f_arrdiv32_not8;
  wire f_arrdiv32_fs288_xor0;
  wire f_arrdiv32_fs288_not0;
  wire f_arrdiv32_fs288_and0;
  wire f_arrdiv32_fs288_not1;
  wire f_arrdiv32_fs289_xor0;
  wire f_arrdiv32_fs289_not0;
  wire f_arrdiv32_fs289_and0;
  wire f_arrdiv32_fs289_xor1;
  wire f_arrdiv32_fs289_not1;
  wire f_arrdiv32_fs289_and1;
  wire f_arrdiv32_fs289_or0;
  wire f_arrdiv32_fs290_xor0;
  wire f_arrdiv32_fs290_not0;
  wire f_arrdiv32_fs290_and0;
  wire f_arrdiv32_fs290_xor1;
  wire f_arrdiv32_fs290_not1;
  wire f_arrdiv32_fs290_and1;
  wire f_arrdiv32_fs290_or0;
  wire f_arrdiv32_fs291_xor0;
  wire f_arrdiv32_fs291_not0;
  wire f_arrdiv32_fs291_and0;
  wire f_arrdiv32_fs291_xor1;
  wire f_arrdiv32_fs291_not1;
  wire f_arrdiv32_fs291_and1;
  wire f_arrdiv32_fs291_or0;
  wire f_arrdiv32_fs292_xor0;
  wire f_arrdiv32_fs292_not0;
  wire f_arrdiv32_fs292_and0;
  wire f_arrdiv32_fs292_xor1;
  wire f_arrdiv32_fs292_not1;
  wire f_arrdiv32_fs292_and1;
  wire f_arrdiv32_fs292_or0;
  wire f_arrdiv32_fs293_xor0;
  wire f_arrdiv32_fs293_not0;
  wire f_arrdiv32_fs293_and0;
  wire f_arrdiv32_fs293_xor1;
  wire f_arrdiv32_fs293_not1;
  wire f_arrdiv32_fs293_and1;
  wire f_arrdiv32_fs293_or0;
  wire f_arrdiv32_fs294_xor0;
  wire f_arrdiv32_fs294_not0;
  wire f_arrdiv32_fs294_and0;
  wire f_arrdiv32_fs294_xor1;
  wire f_arrdiv32_fs294_not1;
  wire f_arrdiv32_fs294_and1;
  wire f_arrdiv32_fs294_or0;
  wire f_arrdiv32_fs295_xor0;
  wire f_arrdiv32_fs295_not0;
  wire f_arrdiv32_fs295_and0;
  wire f_arrdiv32_fs295_xor1;
  wire f_arrdiv32_fs295_not1;
  wire f_arrdiv32_fs295_and1;
  wire f_arrdiv32_fs295_or0;
  wire f_arrdiv32_fs296_xor0;
  wire f_arrdiv32_fs296_not0;
  wire f_arrdiv32_fs296_and0;
  wire f_arrdiv32_fs296_xor1;
  wire f_arrdiv32_fs296_not1;
  wire f_arrdiv32_fs296_and1;
  wire f_arrdiv32_fs296_or0;
  wire f_arrdiv32_fs297_xor0;
  wire f_arrdiv32_fs297_not0;
  wire f_arrdiv32_fs297_and0;
  wire f_arrdiv32_fs297_xor1;
  wire f_arrdiv32_fs297_not1;
  wire f_arrdiv32_fs297_and1;
  wire f_arrdiv32_fs297_or0;
  wire f_arrdiv32_fs298_xor0;
  wire f_arrdiv32_fs298_not0;
  wire f_arrdiv32_fs298_and0;
  wire f_arrdiv32_fs298_xor1;
  wire f_arrdiv32_fs298_not1;
  wire f_arrdiv32_fs298_and1;
  wire f_arrdiv32_fs298_or0;
  wire f_arrdiv32_fs299_xor0;
  wire f_arrdiv32_fs299_not0;
  wire f_arrdiv32_fs299_and0;
  wire f_arrdiv32_fs299_xor1;
  wire f_arrdiv32_fs299_not1;
  wire f_arrdiv32_fs299_and1;
  wire f_arrdiv32_fs299_or0;
  wire f_arrdiv32_fs300_xor0;
  wire f_arrdiv32_fs300_not0;
  wire f_arrdiv32_fs300_and0;
  wire f_arrdiv32_fs300_xor1;
  wire f_arrdiv32_fs300_not1;
  wire f_arrdiv32_fs300_and1;
  wire f_arrdiv32_fs300_or0;
  wire f_arrdiv32_fs301_xor0;
  wire f_arrdiv32_fs301_not0;
  wire f_arrdiv32_fs301_and0;
  wire f_arrdiv32_fs301_xor1;
  wire f_arrdiv32_fs301_not1;
  wire f_arrdiv32_fs301_and1;
  wire f_arrdiv32_fs301_or0;
  wire f_arrdiv32_fs302_xor0;
  wire f_arrdiv32_fs302_not0;
  wire f_arrdiv32_fs302_and0;
  wire f_arrdiv32_fs302_xor1;
  wire f_arrdiv32_fs302_not1;
  wire f_arrdiv32_fs302_and1;
  wire f_arrdiv32_fs302_or0;
  wire f_arrdiv32_fs303_xor0;
  wire f_arrdiv32_fs303_not0;
  wire f_arrdiv32_fs303_and0;
  wire f_arrdiv32_fs303_xor1;
  wire f_arrdiv32_fs303_not1;
  wire f_arrdiv32_fs303_and1;
  wire f_arrdiv32_fs303_or0;
  wire f_arrdiv32_fs304_xor0;
  wire f_arrdiv32_fs304_not0;
  wire f_arrdiv32_fs304_and0;
  wire f_arrdiv32_fs304_xor1;
  wire f_arrdiv32_fs304_not1;
  wire f_arrdiv32_fs304_and1;
  wire f_arrdiv32_fs304_or0;
  wire f_arrdiv32_fs305_xor0;
  wire f_arrdiv32_fs305_not0;
  wire f_arrdiv32_fs305_and0;
  wire f_arrdiv32_fs305_xor1;
  wire f_arrdiv32_fs305_not1;
  wire f_arrdiv32_fs305_and1;
  wire f_arrdiv32_fs305_or0;
  wire f_arrdiv32_fs306_xor0;
  wire f_arrdiv32_fs306_not0;
  wire f_arrdiv32_fs306_and0;
  wire f_arrdiv32_fs306_xor1;
  wire f_arrdiv32_fs306_not1;
  wire f_arrdiv32_fs306_and1;
  wire f_arrdiv32_fs306_or0;
  wire f_arrdiv32_fs307_xor0;
  wire f_arrdiv32_fs307_not0;
  wire f_arrdiv32_fs307_and0;
  wire f_arrdiv32_fs307_xor1;
  wire f_arrdiv32_fs307_not1;
  wire f_arrdiv32_fs307_and1;
  wire f_arrdiv32_fs307_or0;
  wire f_arrdiv32_fs308_xor0;
  wire f_arrdiv32_fs308_not0;
  wire f_arrdiv32_fs308_and0;
  wire f_arrdiv32_fs308_xor1;
  wire f_arrdiv32_fs308_not1;
  wire f_arrdiv32_fs308_and1;
  wire f_arrdiv32_fs308_or0;
  wire f_arrdiv32_fs309_xor0;
  wire f_arrdiv32_fs309_not0;
  wire f_arrdiv32_fs309_and0;
  wire f_arrdiv32_fs309_xor1;
  wire f_arrdiv32_fs309_not1;
  wire f_arrdiv32_fs309_and1;
  wire f_arrdiv32_fs309_or0;
  wire f_arrdiv32_fs310_xor0;
  wire f_arrdiv32_fs310_not0;
  wire f_arrdiv32_fs310_and0;
  wire f_arrdiv32_fs310_xor1;
  wire f_arrdiv32_fs310_not1;
  wire f_arrdiv32_fs310_and1;
  wire f_arrdiv32_fs310_or0;
  wire f_arrdiv32_fs311_xor0;
  wire f_arrdiv32_fs311_not0;
  wire f_arrdiv32_fs311_and0;
  wire f_arrdiv32_fs311_xor1;
  wire f_arrdiv32_fs311_not1;
  wire f_arrdiv32_fs311_and1;
  wire f_arrdiv32_fs311_or0;
  wire f_arrdiv32_fs312_xor0;
  wire f_arrdiv32_fs312_not0;
  wire f_arrdiv32_fs312_and0;
  wire f_arrdiv32_fs312_xor1;
  wire f_arrdiv32_fs312_not1;
  wire f_arrdiv32_fs312_and1;
  wire f_arrdiv32_fs312_or0;
  wire f_arrdiv32_fs313_xor0;
  wire f_arrdiv32_fs313_not0;
  wire f_arrdiv32_fs313_and0;
  wire f_arrdiv32_fs313_xor1;
  wire f_arrdiv32_fs313_not1;
  wire f_arrdiv32_fs313_and1;
  wire f_arrdiv32_fs313_or0;
  wire f_arrdiv32_fs314_xor0;
  wire f_arrdiv32_fs314_not0;
  wire f_arrdiv32_fs314_and0;
  wire f_arrdiv32_fs314_xor1;
  wire f_arrdiv32_fs314_not1;
  wire f_arrdiv32_fs314_and1;
  wire f_arrdiv32_fs314_or0;
  wire f_arrdiv32_fs315_xor0;
  wire f_arrdiv32_fs315_not0;
  wire f_arrdiv32_fs315_and0;
  wire f_arrdiv32_fs315_xor1;
  wire f_arrdiv32_fs315_not1;
  wire f_arrdiv32_fs315_and1;
  wire f_arrdiv32_fs315_or0;
  wire f_arrdiv32_fs316_xor0;
  wire f_arrdiv32_fs316_not0;
  wire f_arrdiv32_fs316_and0;
  wire f_arrdiv32_fs316_xor1;
  wire f_arrdiv32_fs316_not1;
  wire f_arrdiv32_fs316_and1;
  wire f_arrdiv32_fs316_or0;
  wire f_arrdiv32_fs317_xor0;
  wire f_arrdiv32_fs317_not0;
  wire f_arrdiv32_fs317_and0;
  wire f_arrdiv32_fs317_xor1;
  wire f_arrdiv32_fs317_not1;
  wire f_arrdiv32_fs317_and1;
  wire f_arrdiv32_fs317_or0;
  wire f_arrdiv32_fs318_xor0;
  wire f_arrdiv32_fs318_not0;
  wire f_arrdiv32_fs318_and0;
  wire f_arrdiv32_fs318_xor1;
  wire f_arrdiv32_fs318_not1;
  wire f_arrdiv32_fs318_and1;
  wire f_arrdiv32_fs318_or0;
  wire f_arrdiv32_fs319_xor0;
  wire f_arrdiv32_fs319_not0;
  wire f_arrdiv32_fs319_and0;
  wire f_arrdiv32_fs319_xor1;
  wire f_arrdiv32_fs319_not1;
  wire f_arrdiv32_fs319_and1;
  wire f_arrdiv32_fs319_or0;
  wire f_arrdiv32_mux2to1279_and0;
  wire f_arrdiv32_mux2to1279_not0;
  wire f_arrdiv32_mux2to1279_and1;
  wire f_arrdiv32_mux2to1279_xor0;
  wire f_arrdiv32_mux2to1280_and0;
  wire f_arrdiv32_mux2to1280_not0;
  wire f_arrdiv32_mux2to1280_and1;
  wire f_arrdiv32_mux2to1280_xor0;
  wire f_arrdiv32_mux2to1281_and0;
  wire f_arrdiv32_mux2to1281_not0;
  wire f_arrdiv32_mux2to1281_and1;
  wire f_arrdiv32_mux2to1281_xor0;
  wire f_arrdiv32_mux2to1282_and0;
  wire f_arrdiv32_mux2to1282_not0;
  wire f_arrdiv32_mux2to1282_and1;
  wire f_arrdiv32_mux2to1282_xor0;
  wire f_arrdiv32_mux2to1283_and0;
  wire f_arrdiv32_mux2to1283_not0;
  wire f_arrdiv32_mux2to1283_and1;
  wire f_arrdiv32_mux2to1283_xor0;
  wire f_arrdiv32_mux2to1284_and0;
  wire f_arrdiv32_mux2to1284_not0;
  wire f_arrdiv32_mux2to1284_and1;
  wire f_arrdiv32_mux2to1284_xor0;
  wire f_arrdiv32_mux2to1285_and0;
  wire f_arrdiv32_mux2to1285_not0;
  wire f_arrdiv32_mux2to1285_and1;
  wire f_arrdiv32_mux2to1285_xor0;
  wire f_arrdiv32_mux2to1286_and0;
  wire f_arrdiv32_mux2to1286_not0;
  wire f_arrdiv32_mux2to1286_and1;
  wire f_arrdiv32_mux2to1286_xor0;
  wire f_arrdiv32_mux2to1287_and0;
  wire f_arrdiv32_mux2to1287_not0;
  wire f_arrdiv32_mux2to1287_and1;
  wire f_arrdiv32_mux2to1287_xor0;
  wire f_arrdiv32_mux2to1288_and0;
  wire f_arrdiv32_mux2to1288_not0;
  wire f_arrdiv32_mux2to1288_and1;
  wire f_arrdiv32_mux2to1288_xor0;
  wire f_arrdiv32_mux2to1289_and0;
  wire f_arrdiv32_mux2to1289_not0;
  wire f_arrdiv32_mux2to1289_and1;
  wire f_arrdiv32_mux2to1289_xor0;
  wire f_arrdiv32_mux2to1290_and0;
  wire f_arrdiv32_mux2to1290_not0;
  wire f_arrdiv32_mux2to1290_and1;
  wire f_arrdiv32_mux2to1290_xor0;
  wire f_arrdiv32_mux2to1291_and0;
  wire f_arrdiv32_mux2to1291_not0;
  wire f_arrdiv32_mux2to1291_and1;
  wire f_arrdiv32_mux2to1291_xor0;
  wire f_arrdiv32_mux2to1292_and0;
  wire f_arrdiv32_mux2to1292_not0;
  wire f_arrdiv32_mux2to1292_and1;
  wire f_arrdiv32_mux2to1292_xor0;
  wire f_arrdiv32_mux2to1293_and0;
  wire f_arrdiv32_mux2to1293_not0;
  wire f_arrdiv32_mux2to1293_and1;
  wire f_arrdiv32_mux2to1293_xor0;
  wire f_arrdiv32_mux2to1294_and0;
  wire f_arrdiv32_mux2to1294_not0;
  wire f_arrdiv32_mux2to1294_and1;
  wire f_arrdiv32_mux2to1294_xor0;
  wire f_arrdiv32_mux2to1295_and0;
  wire f_arrdiv32_mux2to1295_not0;
  wire f_arrdiv32_mux2to1295_and1;
  wire f_arrdiv32_mux2to1295_xor0;
  wire f_arrdiv32_mux2to1296_and0;
  wire f_arrdiv32_mux2to1296_not0;
  wire f_arrdiv32_mux2to1296_and1;
  wire f_arrdiv32_mux2to1296_xor0;
  wire f_arrdiv32_mux2to1297_and0;
  wire f_arrdiv32_mux2to1297_not0;
  wire f_arrdiv32_mux2to1297_and1;
  wire f_arrdiv32_mux2to1297_xor0;
  wire f_arrdiv32_mux2to1298_and0;
  wire f_arrdiv32_mux2to1298_not0;
  wire f_arrdiv32_mux2to1298_and1;
  wire f_arrdiv32_mux2to1298_xor0;
  wire f_arrdiv32_mux2to1299_and0;
  wire f_arrdiv32_mux2to1299_not0;
  wire f_arrdiv32_mux2to1299_and1;
  wire f_arrdiv32_mux2to1299_xor0;
  wire f_arrdiv32_mux2to1300_and0;
  wire f_arrdiv32_mux2to1300_not0;
  wire f_arrdiv32_mux2to1300_and1;
  wire f_arrdiv32_mux2to1300_xor0;
  wire f_arrdiv32_mux2to1301_and0;
  wire f_arrdiv32_mux2to1301_not0;
  wire f_arrdiv32_mux2to1301_and1;
  wire f_arrdiv32_mux2to1301_xor0;
  wire f_arrdiv32_mux2to1302_and0;
  wire f_arrdiv32_mux2to1302_not0;
  wire f_arrdiv32_mux2to1302_and1;
  wire f_arrdiv32_mux2to1302_xor0;
  wire f_arrdiv32_mux2to1303_and0;
  wire f_arrdiv32_mux2to1303_not0;
  wire f_arrdiv32_mux2to1303_and1;
  wire f_arrdiv32_mux2to1303_xor0;
  wire f_arrdiv32_mux2to1304_and0;
  wire f_arrdiv32_mux2to1304_not0;
  wire f_arrdiv32_mux2to1304_and1;
  wire f_arrdiv32_mux2to1304_xor0;
  wire f_arrdiv32_mux2to1305_and0;
  wire f_arrdiv32_mux2to1305_not0;
  wire f_arrdiv32_mux2to1305_and1;
  wire f_arrdiv32_mux2to1305_xor0;
  wire f_arrdiv32_mux2to1306_and0;
  wire f_arrdiv32_mux2to1306_not0;
  wire f_arrdiv32_mux2to1306_and1;
  wire f_arrdiv32_mux2to1306_xor0;
  wire f_arrdiv32_mux2to1307_and0;
  wire f_arrdiv32_mux2to1307_not0;
  wire f_arrdiv32_mux2to1307_and1;
  wire f_arrdiv32_mux2to1307_xor0;
  wire f_arrdiv32_mux2to1308_and0;
  wire f_arrdiv32_mux2to1308_not0;
  wire f_arrdiv32_mux2to1308_and1;
  wire f_arrdiv32_mux2to1308_xor0;
  wire f_arrdiv32_mux2to1309_and0;
  wire f_arrdiv32_mux2to1309_not0;
  wire f_arrdiv32_mux2to1309_and1;
  wire f_arrdiv32_mux2to1309_xor0;
  wire f_arrdiv32_not9;
  wire f_arrdiv32_fs320_xor0;
  wire f_arrdiv32_fs320_not0;
  wire f_arrdiv32_fs320_and0;
  wire f_arrdiv32_fs320_not1;
  wire f_arrdiv32_fs321_xor0;
  wire f_arrdiv32_fs321_not0;
  wire f_arrdiv32_fs321_and0;
  wire f_arrdiv32_fs321_xor1;
  wire f_arrdiv32_fs321_not1;
  wire f_arrdiv32_fs321_and1;
  wire f_arrdiv32_fs321_or0;
  wire f_arrdiv32_fs322_xor0;
  wire f_arrdiv32_fs322_not0;
  wire f_arrdiv32_fs322_and0;
  wire f_arrdiv32_fs322_xor1;
  wire f_arrdiv32_fs322_not1;
  wire f_arrdiv32_fs322_and1;
  wire f_arrdiv32_fs322_or0;
  wire f_arrdiv32_fs323_xor0;
  wire f_arrdiv32_fs323_not0;
  wire f_arrdiv32_fs323_and0;
  wire f_arrdiv32_fs323_xor1;
  wire f_arrdiv32_fs323_not1;
  wire f_arrdiv32_fs323_and1;
  wire f_arrdiv32_fs323_or0;
  wire f_arrdiv32_fs324_xor0;
  wire f_arrdiv32_fs324_not0;
  wire f_arrdiv32_fs324_and0;
  wire f_arrdiv32_fs324_xor1;
  wire f_arrdiv32_fs324_not1;
  wire f_arrdiv32_fs324_and1;
  wire f_arrdiv32_fs324_or0;
  wire f_arrdiv32_fs325_xor0;
  wire f_arrdiv32_fs325_not0;
  wire f_arrdiv32_fs325_and0;
  wire f_arrdiv32_fs325_xor1;
  wire f_arrdiv32_fs325_not1;
  wire f_arrdiv32_fs325_and1;
  wire f_arrdiv32_fs325_or0;
  wire f_arrdiv32_fs326_xor0;
  wire f_arrdiv32_fs326_not0;
  wire f_arrdiv32_fs326_and0;
  wire f_arrdiv32_fs326_xor1;
  wire f_arrdiv32_fs326_not1;
  wire f_arrdiv32_fs326_and1;
  wire f_arrdiv32_fs326_or0;
  wire f_arrdiv32_fs327_xor0;
  wire f_arrdiv32_fs327_not0;
  wire f_arrdiv32_fs327_and0;
  wire f_arrdiv32_fs327_xor1;
  wire f_arrdiv32_fs327_not1;
  wire f_arrdiv32_fs327_and1;
  wire f_arrdiv32_fs327_or0;
  wire f_arrdiv32_fs328_xor0;
  wire f_arrdiv32_fs328_not0;
  wire f_arrdiv32_fs328_and0;
  wire f_arrdiv32_fs328_xor1;
  wire f_arrdiv32_fs328_not1;
  wire f_arrdiv32_fs328_and1;
  wire f_arrdiv32_fs328_or0;
  wire f_arrdiv32_fs329_xor0;
  wire f_arrdiv32_fs329_not0;
  wire f_arrdiv32_fs329_and0;
  wire f_arrdiv32_fs329_xor1;
  wire f_arrdiv32_fs329_not1;
  wire f_arrdiv32_fs329_and1;
  wire f_arrdiv32_fs329_or0;
  wire f_arrdiv32_fs330_xor0;
  wire f_arrdiv32_fs330_not0;
  wire f_arrdiv32_fs330_and0;
  wire f_arrdiv32_fs330_xor1;
  wire f_arrdiv32_fs330_not1;
  wire f_arrdiv32_fs330_and1;
  wire f_arrdiv32_fs330_or0;
  wire f_arrdiv32_fs331_xor0;
  wire f_arrdiv32_fs331_not0;
  wire f_arrdiv32_fs331_and0;
  wire f_arrdiv32_fs331_xor1;
  wire f_arrdiv32_fs331_not1;
  wire f_arrdiv32_fs331_and1;
  wire f_arrdiv32_fs331_or0;
  wire f_arrdiv32_fs332_xor0;
  wire f_arrdiv32_fs332_not0;
  wire f_arrdiv32_fs332_and0;
  wire f_arrdiv32_fs332_xor1;
  wire f_arrdiv32_fs332_not1;
  wire f_arrdiv32_fs332_and1;
  wire f_arrdiv32_fs332_or0;
  wire f_arrdiv32_fs333_xor0;
  wire f_arrdiv32_fs333_not0;
  wire f_arrdiv32_fs333_and0;
  wire f_arrdiv32_fs333_xor1;
  wire f_arrdiv32_fs333_not1;
  wire f_arrdiv32_fs333_and1;
  wire f_arrdiv32_fs333_or0;
  wire f_arrdiv32_fs334_xor0;
  wire f_arrdiv32_fs334_not0;
  wire f_arrdiv32_fs334_and0;
  wire f_arrdiv32_fs334_xor1;
  wire f_arrdiv32_fs334_not1;
  wire f_arrdiv32_fs334_and1;
  wire f_arrdiv32_fs334_or0;
  wire f_arrdiv32_fs335_xor0;
  wire f_arrdiv32_fs335_not0;
  wire f_arrdiv32_fs335_and0;
  wire f_arrdiv32_fs335_xor1;
  wire f_arrdiv32_fs335_not1;
  wire f_arrdiv32_fs335_and1;
  wire f_arrdiv32_fs335_or0;
  wire f_arrdiv32_fs336_xor0;
  wire f_arrdiv32_fs336_not0;
  wire f_arrdiv32_fs336_and0;
  wire f_arrdiv32_fs336_xor1;
  wire f_arrdiv32_fs336_not1;
  wire f_arrdiv32_fs336_and1;
  wire f_arrdiv32_fs336_or0;
  wire f_arrdiv32_fs337_xor0;
  wire f_arrdiv32_fs337_not0;
  wire f_arrdiv32_fs337_and0;
  wire f_arrdiv32_fs337_xor1;
  wire f_arrdiv32_fs337_not1;
  wire f_arrdiv32_fs337_and1;
  wire f_arrdiv32_fs337_or0;
  wire f_arrdiv32_fs338_xor0;
  wire f_arrdiv32_fs338_not0;
  wire f_arrdiv32_fs338_and0;
  wire f_arrdiv32_fs338_xor1;
  wire f_arrdiv32_fs338_not1;
  wire f_arrdiv32_fs338_and1;
  wire f_arrdiv32_fs338_or0;
  wire f_arrdiv32_fs339_xor0;
  wire f_arrdiv32_fs339_not0;
  wire f_arrdiv32_fs339_and0;
  wire f_arrdiv32_fs339_xor1;
  wire f_arrdiv32_fs339_not1;
  wire f_arrdiv32_fs339_and1;
  wire f_arrdiv32_fs339_or0;
  wire f_arrdiv32_fs340_xor0;
  wire f_arrdiv32_fs340_not0;
  wire f_arrdiv32_fs340_and0;
  wire f_arrdiv32_fs340_xor1;
  wire f_arrdiv32_fs340_not1;
  wire f_arrdiv32_fs340_and1;
  wire f_arrdiv32_fs340_or0;
  wire f_arrdiv32_fs341_xor0;
  wire f_arrdiv32_fs341_not0;
  wire f_arrdiv32_fs341_and0;
  wire f_arrdiv32_fs341_xor1;
  wire f_arrdiv32_fs341_not1;
  wire f_arrdiv32_fs341_and1;
  wire f_arrdiv32_fs341_or0;
  wire f_arrdiv32_fs342_xor0;
  wire f_arrdiv32_fs342_not0;
  wire f_arrdiv32_fs342_and0;
  wire f_arrdiv32_fs342_xor1;
  wire f_arrdiv32_fs342_not1;
  wire f_arrdiv32_fs342_and1;
  wire f_arrdiv32_fs342_or0;
  wire f_arrdiv32_fs343_xor0;
  wire f_arrdiv32_fs343_not0;
  wire f_arrdiv32_fs343_and0;
  wire f_arrdiv32_fs343_xor1;
  wire f_arrdiv32_fs343_not1;
  wire f_arrdiv32_fs343_and1;
  wire f_arrdiv32_fs343_or0;
  wire f_arrdiv32_fs344_xor0;
  wire f_arrdiv32_fs344_not0;
  wire f_arrdiv32_fs344_and0;
  wire f_arrdiv32_fs344_xor1;
  wire f_arrdiv32_fs344_not1;
  wire f_arrdiv32_fs344_and1;
  wire f_arrdiv32_fs344_or0;
  wire f_arrdiv32_fs345_xor0;
  wire f_arrdiv32_fs345_not0;
  wire f_arrdiv32_fs345_and0;
  wire f_arrdiv32_fs345_xor1;
  wire f_arrdiv32_fs345_not1;
  wire f_arrdiv32_fs345_and1;
  wire f_arrdiv32_fs345_or0;
  wire f_arrdiv32_fs346_xor0;
  wire f_arrdiv32_fs346_not0;
  wire f_arrdiv32_fs346_and0;
  wire f_arrdiv32_fs346_xor1;
  wire f_arrdiv32_fs346_not1;
  wire f_arrdiv32_fs346_and1;
  wire f_arrdiv32_fs346_or0;
  wire f_arrdiv32_fs347_xor0;
  wire f_arrdiv32_fs347_not0;
  wire f_arrdiv32_fs347_and0;
  wire f_arrdiv32_fs347_xor1;
  wire f_arrdiv32_fs347_not1;
  wire f_arrdiv32_fs347_and1;
  wire f_arrdiv32_fs347_or0;
  wire f_arrdiv32_fs348_xor0;
  wire f_arrdiv32_fs348_not0;
  wire f_arrdiv32_fs348_and0;
  wire f_arrdiv32_fs348_xor1;
  wire f_arrdiv32_fs348_not1;
  wire f_arrdiv32_fs348_and1;
  wire f_arrdiv32_fs348_or0;
  wire f_arrdiv32_fs349_xor0;
  wire f_arrdiv32_fs349_not0;
  wire f_arrdiv32_fs349_and0;
  wire f_arrdiv32_fs349_xor1;
  wire f_arrdiv32_fs349_not1;
  wire f_arrdiv32_fs349_and1;
  wire f_arrdiv32_fs349_or0;
  wire f_arrdiv32_fs350_xor0;
  wire f_arrdiv32_fs350_not0;
  wire f_arrdiv32_fs350_and0;
  wire f_arrdiv32_fs350_xor1;
  wire f_arrdiv32_fs350_not1;
  wire f_arrdiv32_fs350_and1;
  wire f_arrdiv32_fs350_or0;
  wire f_arrdiv32_fs351_xor0;
  wire f_arrdiv32_fs351_not0;
  wire f_arrdiv32_fs351_and0;
  wire f_arrdiv32_fs351_xor1;
  wire f_arrdiv32_fs351_not1;
  wire f_arrdiv32_fs351_and1;
  wire f_arrdiv32_fs351_or0;
  wire f_arrdiv32_mux2to1310_and0;
  wire f_arrdiv32_mux2to1310_not0;
  wire f_arrdiv32_mux2to1310_and1;
  wire f_arrdiv32_mux2to1310_xor0;
  wire f_arrdiv32_mux2to1311_and0;
  wire f_arrdiv32_mux2to1311_not0;
  wire f_arrdiv32_mux2to1311_and1;
  wire f_arrdiv32_mux2to1311_xor0;
  wire f_arrdiv32_mux2to1312_and0;
  wire f_arrdiv32_mux2to1312_not0;
  wire f_arrdiv32_mux2to1312_and1;
  wire f_arrdiv32_mux2to1312_xor0;
  wire f_arrdiv32_mux2to1313_and0;
  wire f_arrdiv32_mux2to1313_not0;
  wire f_arrdiv32_mux2to1313_and1;
  wire f_arrdiv32_mux2to1313_xor0;
  wire f_arrdiv32_mux2to1314_and0;
  wire f_arrdiv32_mux2to1314_not0;
  wire f_arrdiv32_mux2to1314_and1;
  wire f_arrdiv32_mux2to1314_xor0;
  wire f_arrdiv32_mux2to1315_and0;
  wire f_arrdiv32_mux2to1315_not0;
  wire f_arrdiv32_mux2to1315_and1;
  wire f_arrdiv32_mux2to1315_xor0;
  wire f_arrdiv32_mux2to1316_and0;
  wire f_arrdiv32_mux2to1316_not0;
  wire f_arrdiv32_mux2to1316_and1;
  wire f_arrdiv32_mux2to1316_xor0;
  wire f_arrdiv32_mux2to1317_and0;
  wire f_arrdiv32_mux2to1317_not0;
  wire f_arrdiv32_mux2to1317_and1;
  wire f_arrdiv32_mux2to1317_xor0;
  wire f_arrdiv32_mux2to1318_and0;
  wire f_arrdiv32_mux2to1318_not0;
  wire f_arrdiv32_mux2to1318_and1;
  wire f_arrdiv32_mux2to1318_xor0;
  wire f_arrdiv32_mux2to1319_and0;
  wire f_arrdiv32_mux2to1319_not0;
  wire f_arrdiv32_mux2to1319_and1;
  wire f_arrdiv32_mux2to1319_xor0;
  wire f_arrdiv32_mux2to1320_and0;
  wire f_arrdiv32_mux2to1320_not0;
  wire f_arrdiv32_mux2to1320_and1;
  wire f_arrdiv32_mux2to1320_xor0;
  wire f_arrdiv32_mux2to1321_and0;
  wire f_arrdiv32_mux2to1321_not0;
  wire f_arrdiv32_mux2to1321_and1;
  wire f_arrdiv32_mux2to1321_xor0;
  wire f_arrdiv32_mux2to1322_and0;
  wire f_arrdiv32_mux2to1322_not0;
  wire f_arrdiv32_mux2to1322_and1;
  wire f_arrdiv32_mux2to1322_xor0;
  wire f_arrdiv32_mux2to1323_and0;
  wire f_arrdiv32_mux2to1323_not0;
  wire f_arrdiv32_mux2to1323_and1;
  wire f_arrdiv32_mux2to1323_xor0;
  wire f_arrdiv32_mux2to1324_and0;
  wire f_arrdiv32_mux2to1324_not0;
  wire f_arrdiv32_mux2to1324_and1;
  wire f_arrdiv32_mux2to1324_xor0;
  wire f_arrdiv32_mux2to1325_and0;
  wire f_arrdiv32_mux2to1325_not0;
  wire f_arrdiv32_mux2to1325_and1;
  wire f_arrdiv32_mux2to1325_xor0;
  wire f_arrdiv32_mux2to1326_and0;
  wire f_arrdiv32_mux2to1326_not0;
  wire f_arrdiv32_mux2to1326_and1;
  wire f_arrdiv32_mux2to1326_xor0;
  wire f_arrdiv32_mux2to1327_and0;
  wire f_arrdiv32_mux2to1327_not0;
  wire f_arrdiv32_mux2to1327_and1;
  wire f_arrdiv32_mux2to1327_xor0;
  wire f_arrdiv32_mux2to1328_and0;
  wire f_arrdiv32_mux2to1328_not0;
  wire f_arrdiv32_mux2to1328_and1;
  wire f_arrdiv32_mux2to1328_xor0;
  wire f_arrdiv32_mux2to1329_and0;
  wire f_arrdiv32_mux2to1329_not0;
  wire f_arrdiv32_mux2to1329_and1;
  wire f_arrdiv32_mux2to1329_xor0;
  wire f_arrdiv32_mux2to1330_and0;
  wire f_arrdiv32_mux2to1330_not0;
  wire f_arrdiv32_mux2to1330_and1;
  wire f_arrdiv32_mux2to1330_xor0;
  wire f_arrdiv32_mux2to1331_and0;
  wire f_arrdiv32_mux2to1331_not0;
  wire f_arrdiv32_mux2to1331_and1;
  wire f_arrdiv32_mux2to1331_xor0;
  wire f_arrdiv32_mux2to1332_and0;
  wire f_arrdiv32_mux2to1332_not0;
  wire f_arrdiv32_mux2to1332_and1;
  wire f_arrdiv32_mux2to1332_xor0;
  wire f_arrdiv32_mux2to1333_and0;
  wire f_arrdiv32_mux2to1333_not0;
  wire f_arrdiv32_mux2to1333_and1;
  wire f_arrdiv32_mux2to1333_xor0;
  wire f_arrdiv32_mux2to1334_and0;
  wire f_arrdiv32_mux2to1334_not0;
  wire f_arrdiv32_mux2to1334_and1;
  wire f_arrdiv32_mux2to1334_xor0;
  wire f_arrdiv32_mux2to1335_and0;
  wire f_arrdiv32_mux2to1335_not0;
  wire f_arrdiv32_mux2to1335_and1;
  wire f_arrdiv32_mux2to1335_xor0;
  wire f_arrdiv32_mux2to1336_and0;
  wire f_arrdiv32_mux2to1336_not0;
  wire f_arrdiv32_mux2to1336_and1;
  wire f_arrdiv32_mux2to1336_xor0;
  wire f_arrdiv32_mux2to1337_and0;
  wire f_arrdiv32_mux2to1337_not0;
  wire f_arrdiv32_mux2to1337_and1;
  wire f_arrdiv32_mux2to1337_xor0;
  wire f_arrdiv32_mux2to1338_and0;
  wire f_arrdiv32_mux2to1338_not0;
  wire f_arrdiv32_mux2to1338_and1;
  wire f_arrdiv32_mux2to1338_xor0;
  wire f_arrdiv32_mux2to1339_and0;
  wire f_arrdiv32_mux2to1339_not0;
  wire f_arrdiv32_mux2to1339_and1;
  wire f_arrdiv32_mux2to1339_xor0;
  wire f_arrdiv32_mux2to1340_and0;
  wire f_arrdiv32_mux2to1340_not0;
  wire f_arrdiv32_mux2to1340_and1;
  wire f_arrdiv32_mux2to1340_xor0;
  wire f_arrdiv32_not10;
  wire f_arrdiv32_fs352_xor0;
  wire f_arrdiv32_fs352_not0;
  wire f_arrdiv32_fs352_and0;
  wire f_arrdiv32_fs352_not1;
  wire f_arrdiv32_fs353_xor0;
  wire f_arrdiv32_fs353_not0;
  wire f_arrdiv32_fs353_and0;
  wire f_arrdiv32_fs353_xor1;
  wire f_arrdiv32_fs353_not1;
  wire f_arrdiv32_fs353_and1;
  wire f_arrdiv32_fs353_or0;
  wire f_arrdiv32_fs354_xor0;
  wire f_arrdiv32_fs354_not0;
  wire f_arrdiv32_fs354_and0;
  wire f_arrdiv32_fs354_xor1;
  wire f_arrdiv32_fs354_not1;
  wire f_arrdiv32_fs354_and1;
  wire f_arrdiv32_fs354_or0;
  wire f_arrdiv32_fs355_xor0;
  wire f_arrdiv32_fs355_not0;
  wire f_arrdiv32_fs355_and0;
  wire f_arrdiv32_fs355_xor1;
  wire f_arrdiv32_fs355_not1;
  wire f_arrdiv32_fs355_and1;
  wire f_arrdiv32_fs355_or0;
  wire f_arrdiv32_fs356_xor0;
  wire f_arrdiv32_fs356_not0;
  wire f_arrdiv32_fs356_and0;
  wire f_arrdiv32_fs356_xor1;
  wire f_arrdiv32_fs356_not1;
  wire f_arrdiv32_fs356_and1;
  wire f_arrdiv32_fs356_or0;
  wire f_arrdiv32_fs357_xor0;
  wire f_arrdiv32_fs357_not0;
  wire f_arrdiv32_fs357_and0;
  wire f_arrdiv32_fs357_xor1;
  wire f_arrdiv32_fs357_not1;
  wire f_arrdiv32_fs357_and1;
  wire f_arrdiv32_fs357_or0;
  wire f_arrdiv32_fs358_xor0;
  wire f_arrdiv32_fs358_not0;
  wire f_arrdiv32_fs358_and0;
  wire f_arrdiv32_fs358_xor1;
  wire f_arrdiv32_fs358_not1;
  wire f_arrdiv32_fs358_and1;
  wire f_arrdiv32_fs358_or0;
  wire f_arrdiv32_fs359_xor0;
  wire f_arrdiv32_fs359_not0;
  wire f_arrdiv32_fs359_and0;
  wire f_arrdiv32_fs359_xor1;
  wire f_arrdiv32_fs359_not1;
  wire f_arrdiv32_fs359_and1;
  wire f_arrdiv32_fs359_or0;
  wire f_arrdiv32_fs360_xor0;
  wire f_arrdiv32_fs360_not0;
  wire f_arrdiv32_fs360_and0;
  wire f_arrdiv32_fs360_xor1;
  wire f_arrdiv32_fs360_not1;
  wire f_arrdiv32_fs360_and1;
  wire f_arrdiv32_fs360_or0;
  wire f_arrdiv32_fs361_xor0;
  wire f_arrdiv32_fs361_not0;
  wire f_arrdiv32_fs361_and0;
  wire f_arrdiv32_fs361_xor1;
  wire f_arrdiv32_fs361_not1;
  wire f_arrdiv32_fs361_and1;
  wire f_arrdiv32_fs361_or0;
  wire f_arrdiv32_fs362_xor0;
  wire f_arrdiv32_fs362_not0;
  wire f_arrdiv32_fs362_and0;
  wire f_arrdiv32_fs362_xor1;
  wire f_arrdiv32_fs362_not1;
  wire f_arrdiv32_fs362_and1;
  wire f_arrdiv32_fs362_or0;
  wire f_arrdiv32_fs363_xor0;
  wire f_arrdiv32_fs363_not0;
  wire f_arrdiv32_fs363_and0;
  wire f_arrdiv32_fs363_xor1;
  wire f_arrdiv32_fs363_not1;
  wire f_arrdiv32_fs363_and1;
  wire f_arrdiv32_fs363_or0;
  wire f_arrdiv32_fs364_xor0;
  wire f_arrdiv32_fs364_not0;
  wire f_arrdiv32_fs364_and0;
  wire f_arrdiv32_fs364_xor1;
  wire f_arrdiv32_fs364_not1;
  wire f_arrdiv32_fs364_and1;
  wire f_arrdiv32_fs364_or0;
  wire f_arrdiv32_fs365_xor0;
  wire f_arrdiv32_fs365_not0;
  wire f_arrdiv32_fs365_and0;
  wire f_arrdiv32_fs365_xor1;
  wire f_arrdiv32_fs365_not1;
  wire f_arrdiv32_fs365_and1;
  wire f_arrdiv32_fs365_or0;
  wire f_arrdiv32_fs366_xor0;
  wire f_arrdiv32_fs366_not0;
  wire f_arrdiv32_fs366_and0;
  wire f_arrdiv32_fs366_xor1;
  wire f_arrdiv32_fs366_not1;
  wire f_arrdiv32_fs366_and1;
  wire f_arrdiv32_fs366_or0;
  wire f_arrdiv32_fs367_xor0;
  wire f_arrdiv32_fs367_not0;
  wire f_arrdiv32_fs367_and0;
  wire f_arrdiv32_fs367_xor1;
  wire f_arrdiv32_fs367_not1;
  wire f_arrdiv32_fs367_and1;
  wire f_arrdiv32_fs367_or0;
  wire f_arrdiv32_fs368_xor0;
  wire f_arrdiv32_fs368_not0;
  wire f_arrdiv32_fs368_and0;
  wire f_arrdiv32_fs368_xor1;
  wire f_arrdiv32_fs368_not1;
  wire f_arrdiv32_fs368_and1;
  wire f_arrdiv32_fs368_or0;
  wire f_arrdiv32_fs369_xor0;
  wire f_arrdiv32_fs369_not0;
  wire f_arrdiv32_fs369_and0;
  wire f_arrdiv32_fs369_xor1;
  wire f_arrdiv32_fs369_not1;
  wire f_arrdiv32_fs369_and1;
  wire f_arrdiv32_fs369_or0;
  wire f_arrdiv32_fs370_xor0;
  wire f_arrdiv32_fs370_not0;
  wire f_arrdiv32_fs370_and0;
  wire f_arrdiv32_fs370_xor1;
  wire f_arrdiv32_fs370_not1;
  wire f_arrdiv32_fs370_and1;
  wire f_arrdiv32_fs370_or0;
  wire f_arrdiv32_fs371_xor0;
  wire f_arrdiv32_fs371_not0;
  wire f_arrdiv32_fs371_and0;
  wire f_arrdiv32_fs371_xor1;
  wire f_arrdiv32_fs371_not1;
  wire f_arrdiv32_fs371_and1;
  wire f_arrdiv32_fs371_or0;
  wire f_arrdiv32_fs372_xor0;
  wire f_arrdiv32_fs372_not0;
  wire f_arrdiv32_fs372_and0;
  wire f_arrdiv32_fs372_xor1;
  wire f_arrdiv32_fs372_not1;
  wire f_arrdiv32_fs372_and1;
  wire f_arrdiv32_fs372_or0;
  wire f_arrdiv32_fs373_xor0;
  wire f_arrdiv32_fs373_not0;
  wire f_arrdiv32_fs373_and0;
  wire f_arrdiv32_fs373_xor1;
  wire f_arrdiv32_fs373_not1;
  wire f_arrdiv32_fs373_and1;
  wire f_arrdiv32_fs373_or0;
  wire f_arrdiv32_fs374_xor0;
  wire f_arrdiv32_fs374_not0;
  wire f_arrdiv32_fs374_and0;
  wire f_arrdiv32_fs374_xor1;
  wire f_arrdiv32_fs374_not1;
  wire f_arrdiv32_fs374_and1;
  wire f_arrdiv32_fs374_or0;
  wire f_arrdiv32_fs375_xor0;
  wire f_arrdiv32_fs375_not0;
  wire f_arrdiv32_fs375_and0;
  wire f_arrdiv32_fs375_xor1;
  wire f_arrdiv32_fs375_not1;
  wire f_arrdiv32_fs375_and1;
  wire f_arrdiv32_fs375_or0;
  wire f_arrdiv32_fs376_xor0;
  wire f_arrdiv32_fs376_not0;
  wire f_arrdiv32_fs376_and0;
  wire f_arrdiv32_fs376_xor1;
  wire f_arrdiv32_fs376_not1;
  wire f_arrdiv32_fs376_and1;
  wire f_arrdiv32_fs376_or0;
  wire f_arrdiv32_fs377_xor0;
  wire f_arrdiv32_fs377_not0;
  wire f_arrdiv32_fs377_and0;
  wire f_arrdiv32_fs377_xor1;
  wire f_arrdiv32_fs377_not1;
  wire f_arrdiv32_fs377_and1;
  wire f_arrdiv32_fs377_or0;
  wire f_arrdiv32_fs378_xor0;
  wire f_arrdiv32_fs378_not0;
  wire f_arrdiv32_fs378_and0;
  wire f_arrdiv32_fs378_xor1;
  wire f_arrdiv32_fs378_not1;
  wire f_arrdiv32_fs378_and1;
  wire f_arrdiv32_fs378_or0;
  wire f_arrdiv32_fs379_xor0;
  wire f_arrdiv32_fs379_not0;
  wire f_arrdiv32_fs379_and0;
  wire f_arrdiv32_fs379_xor1;
  wire f_arrdiv32_fs379_not1;
  wire f_arrdiv32_fs379_and1;
  wire f_arrdiv32_fs379_or0;
  wire f_arrdiv32_fs380_xor0;
  wire f_arrdiv32_fs380_not0;
  wire f_arrdiv32_fs380_and0;
  wire f_arrdiv32_fs380_xor1;
  wire f_arrdiv32_fs380_not1;
  wire f_arrdiv32_fs380_and1;
  wire f_arrdiv32_fs380_or0;
  wire f_arrdiv32_fs381_xor0;
  wire f_arrdiv32_fs381_not0;
  wire f_arrdiv32_fs381_and0;
  wire f_arrdiv32_fs381_xor1;
  wire f_arrdiv32_fs381_not1;
  wire f_arrdiv32_fs381_and1;
  wire f_arrdiv32_fs381_or0;
  wire f_arrdiv32_fs382_xor0;
  wire f_arrdiv32_fs382_not0;
  wire f_arrdiv32_fs382_and0;
  wire f_arrdiv32_fs382_xor1;
  wire f_arrdiv32_fs382_not1;
  wire f_arrdiv32_fs382_and1;
  wire f_arrdiv32_fs382_or0;
  wire f_arrdiv32_fs383_xor0;
  wire f_arrdiv32_fs383_not0;
  wire f_arrdiv32_fs383_and0;
  wire f_arrdiv32_fs383_xor1;
  wire f_arrdiv32_fs383_not1;
  wire f_arrdiv32_fs383_and1;
  wire f_arrdiv32_fs383_or0;
  wire f_arrdiv32_mux2to1341_and0;
  wire f_arrdiv32_mux2to1341_not0;
  wire f_arrdiv32_mux2to1341_and1;
  wire f_arrdiv32_mux2to1341_xor0;
  wire f_arrdiv32_mux2to1342_and0;
  wire f_arrdiv32_mux2to1342_not0;
  wire f_arrdiv32_mux2to1342_and1;
  wire f_arrdiv32_mux2to1342_xor0;
  wire f_arrdiv32_mux2to1343_and0;
  wire f_arrdiv32_mux2to1343_not0;
  wire f_arrdiv32_mux2to1343_and1;
  wire f_arrdiv32_mux2to1343_xor0;
  wire f_arrdiv32_mux2to1344_and0;
  wire f_arrdiv32_mux2to1344_not0;
  wire f_arrdiv32_mux2to1344_and1;
  wire f_arrdiv32_mux2to1344_xor0;
  wire f_arrdiv32_mux2to1345_and0;
  wire f_arrdiv32_mux2to1345_not0;
  wire f_arrdiv32_mux2to1345_and1;
  wire f_arrdiv32_mux2to1345_xor0;
  wire f_arrdiv32_mux2to1346_and0;
  wire f_arrdiv32_mux2to1346_not0;
  wire f_arrdiv32_mux2to1346_and1;
  wire f_arrdiv32_mux2to1346_xor0;
  wire f_arrdiv32_mux2to1347_and0;
  wire f_arrdiv32_mux2to1347_not0;
  wire f_arrdiv32_mux2to1347_and1;
  wire f_arrdiv32_mux2to1347_xor0;
  wire f_arrdiv32_mux2to1348_and0;
  wire f_arrdiv32_mux2to1348_not0;
  wire f_arrdiv32_mux2to1348_and1;
  wire f_arrdiv32_mux2to1348_xor0;
  wire f_arrdiv32_mux2to1349_and0;
  wire f_arrdiv32_mux2to1349_not0;
  wire f_arrdiv32_mux2to1349_and1;
  wire f_arrdiv32_mux2to1349_xor0;
  wire f_arrdiv32_mux2to1350_and0;
  wire f_arrdiv32_mux2to1350_not0;
  wire f_arrdiv32_mux2to1350_and1;
  wire f_arrdiv32_mux2to1350_xor0;
  wire f_arrdiv32_mux2to1351_and0;
  wire f_arrdiv32_mux2to1351_not0;
  wire f_arrdiv32_mux2to1351_and1;
  wire f_arrdiv32_mux2to1351_xor0;
  wire f_arrdiv32_mux2to1352_and0;
  wire f_arrdiv32_mux2to1352_not0;
  wire f_arrdiv32_mux2to1352_and1;
  wire f_arrdiv32_mux2to1352_xor0;
  wire f_arrdiv32_mux2to1353_and0;
  wire f_arrdiv32_mux2to1353_not0;
  wire f_arrdiv32_mux2to1353_and1;
  wire f_arrdiv32_mux2to1353_xor0;
  wire f_arrdiv32_mux2to1354_and0;
  wire f_arrdiv32_mux2to1354_not0;
  wire f_arrdiv32_mux2to1354_and1;
  wire f_arrdiv32_mux2to1354_xor0;
  wire f_arrdiv32_mux2to1355_and0;
  wire f_arrdiv32_mux2to1355_not0;
  wire f_arrdiv32_mux2to1355_and1;
  wire f_arrdiv32_mux2to1355_xor0;
  wire f_arrdiv32_mux2to1356_and0;
  wire f_arrdiv32_mux2to1356_not0;
  wire f_arrdiv32_mux2to1356_and1;
  wire f_arrdiv32_mux2to1356_xor0;
  wire f_arrdiv32_mux2to1357_and0;
  wire f_arrdiv32_mux2to1357_not0;
  wire f_arrdiv32_mux2to1357_and1;
  wire f_arrdiv32_mux2to1357_xor0;
  wire f_arrdiv32_mux2to1358_and0;
  wire f_arrdiv32_mux2to1358_not0;
  wire f_arrdiv32_mux2to1358_and1;
  wire f_arrdiv32_mux2to1358_xor0;
  wire f_arrdiv32_mux2to1359_and0;
  wire f_arrdiv32_mux2to1359_not0;
  wire f_arrdiv32_mux2to1359_and1;
  wire f_arrdiv32_mux2to1359_xor0;
  wire f_arrdiv32_mux2to1360_and0;
  wire f_arrdiv32_mux2to1360_not0;
  wire f_arrdiv32_mux2to1360_and1;
  wire f_arrdiv32_mux2to1360_xor0;
  wire f_arrdiv32_mux2to1361_and0;
  wire f_arrdiv32_mux2to1361_not0;
  wire f_arrdiv32_mux2to1361_and1;
  wire f_arrdiv32_mux2to1361_xor0;
  wire f_arrdiv32_mux2to1362_and0;
  wire f_arrdiv32_mux2to1362_not0;
  wire f_arrdiv32_mux2to1362_and1;
  wire f_arrdiv32_mux2to1362_xor0;
  wire f_arrdiv32_mux2to1363_and0;
  wire f_arrdiv32_mux2to1363_not0;
  wire f_arrdiv32_mux2to1363_and1;
  wire f_arrdiv32_mux2to1363_xor0;
  wire f_arrdiv32_mux2to1364_and0;
  wire f_arrdiv32_mux2to1364_not0;
  wire f_arrdiv32_mux2to1364_and1;
  wire f_arrdiv32_mux2to1364_xor0;
  wire f_arrdiv32_mux2to1365_and0;
  wire f_arrdiv32_mux2to1365_not0;
  wire f_arrdiv32_mux2to1365_and1;
  wire f_arrdiv32_mux2to1365_xor0;
  wire f_arrdiv32_mux2to1366_and0;
  wire f_arrdiv32_mux2to1366_not0;
  wire f_arrdiv32_mux2to1366_and1;
  wire f_arrdiv32_mux2to1366_xor0;
  wire f_arrdiv32_mux2to1367_and0;
  wire f_arrdiv32_mux2to1367_not0;
  wire f_arrdiv32_mux2to1367_and1;
  wire f_arrdiv32_mux2to1367_xor0;
  wire f_arrdiv32_mux2to1368_and0;
  wire f_arrdiv32_mux2to1368_not0;
  wire f_arrdiv32_mux2to1368_and1;
  wire f_arrdiv32_mux2to1368_xor0;
  wire f_arrdiv32_mux2to1369_and0;
  wire f_arrdiv32_mux2to1369_not0;
  wire f_arrdiv32_mux2to1369_and1;
  wire f_arrdiv32_mux2to1369_xor0;
  wire f_arrdiv32_mux2to1370_and0;
  wire f_arrdiv32_mux2to1370_not0;
  wire f_arrdiv32_mux2to1370_and1;
  wire f_arrdiv32_mux2to1370_xor0;
  wire f_arrdiv32_mux2to1371_and0;
  wire f_arrdiv32_mux2to1371_not0;
  wire f_arrdiv32_mux2to1371_and1;
  wire f_arrdiv32_mux2to1371_xor0;
  wire f_arrdiv32_not11;
  wire f_arrdiv32_fs384_xor0;
  wire f_arrdiv32_fs384_not0;
  wire f_arrdiv32_fs384_and0;
  wire f_arrdiv32_fs384_not1;
  wire f_arrdiv32_fs385_xor0;
  wire f_arrdiv32_fs385_not0;
  wire f_arrdiv32_fs385_and0;
  wire f_arrdiv32_fs385_xor1;
  wire f_arrdiv32_fs385_not1;
  wire f_arrdiv32_fs385_and1;
  wire f_arrdiv32_fs385_or0;
  wire f_arrdiv32_fs386_xor0;
  wire f_arrdiv32_fs386_not0;
  wire f_arrdiv32_fs386_and0;
  wire f_arrdiv32_fs386_xor1;
  wire f_arrdiv32_fs386_not1;
  wire f_arrdiv32_fs386_and1;
  wire f_arrdiv32_fs386_or0;
  wire f_arrdiv32_fs387_xor0;
  wire f_arrdiv32_fs387_not0;
  wire f_arrdiv32_fs387_and0;
  wire f_arrdiv32_fs387_xor1;
  wire f_arrdiv32_fs387_not1;
  wire f_arrdiv32_fs387_and1;
  wire f_arrdiv32_fs387_or0;
  wire f_arrdiv32_fs388_xor0;
  wire f_arrdiv32_fs388_not0;
  wire f_arrdiv32_fs388_and0;
  wire f_arrdiv32_fs388_xor1;
  wire f_arrdiv32_fs388_not1;
  wire f_arrdiv32_fs388_and1;
  wire f_arrdiv32_fs388_or0;
  wire f_arrdiv32_fs389_xor0;
  wire f_arrdiv32_fs389_not0;
  wire f_arrdiv32_fs389_and0;
  wire f_arrdiv32_fs389_xor1;
  wire f_arrdiv32_fs389_not1;
  wire f_arrdiv32_fs389_and1;
  wire f_arrdiv32_fs389_or0;
  wire f_arrdiv32_fs390_xor0;
  wire f_arrdiv32_fs390_not0;
  wire f_arrdiv32_fs390_and0;
  wire f_arrdiv32_fs390_xor1;
  wire f_arrdiv32_fs390_not1;
  wire f_arrdiv32_fs390_and1;
  wire f_arrdiv32_fs390_or0;
  wire f_arrdiv32_fs391_xor0;
  wire f_arrdiv32_fs391_not0;
  wire f_arrdiv32_fs391_and0;
  wire f_arrdiv32_fs391_xor1;
  wire f_arrdiv32_fs391_not1;
  wire f_arrdiv32_fs391_and1;
  wire f_arrdiv32_fs391_or0;
  wire f_arrdiv32_fs392_xor0;
  wire f_arrdiv32_fs392_not0;
  wire f_arrdiv32_fs392_and0;
  wire f_arrdiv32_fs392_xor1;
  wire f_arrdiv32_fs392_not1;
  wire f_arrdiv32_fs392_and1;
  wire f_arrdiv32_fs392_or0;
  wire f_arrdiv32_fs393_xor0;
  wire f_arrdiv32_fs393_not0;
  wire f_arrdiv32_fs393_and0;
  wire f_arrdiv32_fs393_xor1;
  wire f_arrdiv32_fs393_not1;
  wire f_arrdiv32_fs393_and1;
  wire f_arrdiv32_fs393_or0;
  wire f_arrdiv32_fs394_xor0;
  wire f_arrdiv32_fs394_not0;
  wire f_arrdiv32_fs394_and0;
  wire f_arrdiv32_fs394_xor1;
  wire f_arrdiv32_fs394_not1;
  wire f_arrdiv32_fs394_and1;
  wire f_arrdiv32_fs394_or0;
  wire f_arrdiv32_fs395_xor0;
  wire f_arrdiv32_fs395_not0;
  wire f_arrdiv32_fs395_and0;
  wire f_arrdiv32_fs395_xor1;
  wire f_arrdiv32_fs395_not1;
  wire f_arrdiv32_fs395_and1;
  wire f_arrdiv32_fs395_or0;
  wire f_arrdiv32_fs396_xor0;
  wire f_arrdiv32_fs396_not0;
  wire f_arrdiv32_fs396_and0;
  wire f_arrdiv32_fs396_xor1;
  wire f_arrdiv32_fs396_not1;
  wire f_arrdiv32_fs396_and1;
  wire f_arrdiv32_fs396_or0;
  wire f_arrdiv32_fs397_xor0;
  wire f_arrdiv32_fs397_not0;
  wire f_arrdiv32_fs397_and0;
  wire f_arrdiv32_fs397_xor1;
  wire f_arrdiv32_fs397_not1;
  wire f_arrdiv32_fs397_and1;
  wire f_arrdiv32_fs397_or0;
  wire f_arrdiv32_fs398_xor0;
  wire f_arrdiv32_fs398_not0;
  wire f_arrdiv32_fs398_and0;
  wire f_arrdiv32_fs398_xor1;
  wire f_arrdiv32_fs398_not1;
  wire f_arrdiv32_fs398_and1;
  wire f_arrdiv32_fs398_or0;
  wire f_arrdiv32_fs399_xor0;
  wire f_arrdiv32_fs399_not0;
  wire f_arrdiv32_fs399_and0;
  wire f_arrdiv32_fs399_xor1;
  wire f_arrdiv32_fs399_not1;
  wire f_arrdiv32_fs399_and1;
  wire f_arrdiv32_fs399_or0;
  wire f_arrdiv32_fs400_xor0;
  wire f_arrdiv32_fs400_not0;
  wire f_arrdiv32_fs400_and0;
  wire f_arrdiv32_fs400_xor1;
  wire f_arrdiv32_fs400_not1;
  wire f_arrdiv32_fs400_and1;
  wire f_arrdiv32_fs400_or0;
  wire f_arrdiv32_fs401_xor0;
  wire f_arrdiv32_fs401_not0;
  wire f_arrdiv32_fs401_and0;
  wire f_arrdiv32_fs401_xor1;
  wire f_arrdiv32_fs401_not1;
  wire f_arrdiv32_fs401_and1;
  wire f_arrdiv32_fs401_or0;
  wire f_arrdiv32_fs402_xor0;
  wire f_arrdiv32_fs402_not0;
  wire f_arrdiv32_fs402_and0;
  wire f_arrdiv32_fs402_xor1;
  wire f_arrdiv32_fs402_not1;
  wire f_arrdiv32_fs402_and1;
  wire f_arrdiv32_fs402_or0;
  wire f_arrdiv32_fs403_xor0;
  wire f_arrdiv32_fs403_not0;
  wire f_arrdiv32_fs403_and0;
  wire f_arrdiv32_fs403_xor1;
  wire f_arrdiv32_fs403_not1;
  wire f_arrdiv32_fs403_and1;
  wire f_arrdiv32_fs403_or0;
  wire f_arrdiv32_fs404_xor0;
  wire f_arrdiv32_fs404_not0;
  wire f_arrdiv32_fs404_and0;
  wire f_arrdiv32_fs404_xor1;
  wire f_arrdiv32_fs404_not1;
  wire f_arrdiv32_fs404_and1;
  wire f_arrdiv32_fs404_or0;
  wire f_arrdiv32_fs405_xor0;
  wire f_arrdiv32_fs405_not0;
  wire f_arrdiv32_fs405_and0;
  wire f_arrdiv32_fs405_xor1;
  wire f_arrdiv32_fs405_not1;
  wire f_arrdiv32_fs405_and1;
  wire f_arrdiv32_fs405_or0;
  wire f_arrdiv32_fs406_xor0;
  wire f_arrdiv32_fs406_not0;
  wire f_arrdiv32_fs406_and0;
  wire f_arrdiv32_fs406_xor1;
  wire f_arrdiv32_fs406_not1;
  wire f_arrdiv32_fs406_and1;
  wire f_arrdiv32_fs406_or0;
  wire f_arrdiv32_fs407_xor0;
  wire f_arrdiv32_fs407_not0;
  wire f_arrdiv32_fs407_and0;
  wire f_arrdiv32_fs407_xor1;
  wire f_arrdiv32_fs407_not1;
  wire f_arrdiv32_fs407_and1;
  wire f_arrdiv32_fs407_or0;
  wire f_arrdiv32_fs408_xor0;
  wire f_arrdiv32_fs408_not0;
  wire f_arrdiv32_fs408_and0;
  wire f_arrdiv32_fs408_xor1;
  wire f_arrdiv32_fs408_not1;
  wire f_arrdiv32_fs408_and1;
  wire f_arrdiv32_fs408_or0;
  wire f_arrdiv32_fs409_xor0;
  wire f_arrdiv32_fs409_not0;
  wire f_arrdiv32_fs409_and0;
  wire f_arrdiv32_fs409_xor1;
  wire f_arrdiv32_fs409_not1;
  wire f_arrdiv32_fs409_and1;
  wire f_arrdiv32_fs409_or0;
  wire f_arrdiv32_fs410_xor0;
  wire f_arrdiv32_fs410_not0;
  wire f_arrdiv32_fs410_and0;
  wire f_arrdiv32_fs410_xor1;
  wire f_arrdiv32_fs410_not1;
  wire f_arrdiv32_fs410_and1;
  wire f_arrdiv32_fs410_or0;
  wire f_arrdiv32_fs411_xor0;
  wire f_arrdiv32_fs411_not0;
  wire f_arrdiv32_fs411_and0;
  wire f_arrdiv32_fs411_xor1;
  wire f_arrdiv32_fs411_not1;
  wire f_arrdiv32_fs411_and1;
  wire f_arrdiv32_fs411_or0;
  wire f_arrdiv32_fs412_xor0;
  wire f_arrdiv32_fs412_not0;
  wire f_arrdiv32_fs412_and0;
  wire f_arrdiv32_fs412_xor1;
  wire f_arrdiv32_fs412_not1;
  wire f_arrdiv32_fs412_and1;
  wire f_arrdiv32_fs412_or0;
  wire f_arrdiv32_fs413_xor0;
  wire f_arrdiv32_fs413_not0;
  wire f_arrdiv32_fs413_and0;
  wire f_arrdiv32_fs413_xor1;
  wire f_arrdiv32_fs413_not1;
  wire f_arrdiv32_fs413_and1;
  wire f_arrdiv32_fs413_or0;
  wire f_arrdiv32_fs414_xor0;
  wire f_arrdiv32_fs414_not0;
  wire f_arrdiv32_fs414_and0;
  wire f_arrdiv32_fs414_xor1;
  wire f_arrdiv32_fs414_not1;
  wire f_arrdiv32_fs414_and1;
  wire f_arrdiv32_fs414_or0;
  wire f_arrdiv32_fs415_xor0;
  wire f_arrdiv32_fs415_not0;
  wire f_arrdiv32_fs415_and0;
  wire f_arrdiv32_fs415_xor1;
  wire f_arrdiv32_fs415_not1;
  wire f_arrdiv32_fs415_and1;
  wire f_arrdiv32_fs415_or0;
  wire f_arrdiv32_mux2to1372_and0;
  wire f_arrdiv32_mux2to1372_not0;
  wire f_arrdiv32_mux2to1372_and1;
  wire f_arrdiv32_mux2to1372_xor0;
  wire f_arrdiv32_mux2to1373_and0;
  wire f_arrdiv32_mux2to1373_not0;
  wire f_arrdiv32_mux2to1373_and1;
  wire f_arrdiv32_mux2to1373_xor0;
  wire f_arrdiv32_mux2to1374_and0;
  wire f_arrdiv32_mux2to1374_not0;
  wire f_arrdiv32_mux2to1374_and1;
  wire f_arrdiv32_mux2to1374_xor0;
  wire f_arrdiv32_mux2to1375_and0;
  wire f_arrdiv32_mux2to1375_not0;
  wire f_arrdiv32_mux2to1375_and1;
  wire f_arrdiv32_mux2to1375_xor0;
  wire f_arrdiv32_mux2to1376_and0;
  wire f_arrdiv32_mux2to1376_not0;
  wire f_arrdiv32_mux2to1376_and1;
  wire f_arrdiv32_mux2to1376_xor0;
  wire f_arrdiv32_mux2to1377_and0;
  wire f_arrdiv32_mux2to1377_not0;
  wire f_arrdiv32_mux2to1377_and1;
  wire f_arrdiv32_mux2to1377_xor0;
  wire f_arrdiv32_mux2to1378_and0;
  wire f_arrdiv32_mux2to1378_not0;
  wire f_arrdiv32_mux2to1378_and1;
  wire f_arrdiv32_mux2to1378_xor0;
  wire f_arrdiv32_mux2to1379_and0;
  wire f_arrdiv32_mux2to1379_not0;
  wire f_arrdiv32_mux2to1379_and1;
  wire f_arrdiv32_mux2to1379_xor0;
  wire f_arrdiv32_mux2to1380_and0;
  wire f_arrdiv32_mux2to1380_not0;
  wire f_arrdiv32_mux2to1380_and1;
  wire f_arrdiv32_mux2to1380_xor0;
  wire f_arrdiv32_mux2to1381_and0;
  wire f_arrdiv32_mux2to1381_not0;
  wire f_arrdiv32_mux2to1381_and1;
  wire f_arrdiv32_mux2to1381_xor0;
  wire f_arrdiv32_mux2to1382_and0;
  wire f_arrdiv32_mux2to1382_not0;
  wire f_arrdiv32_mux2to1382_and1;
  wire f_arrdiv32_mux2to1382_xor0;
  wire f_arrdiv32_mux2to1383_and0;
  wire f_arrdiv32_mux2to1383_not0;
  wire f_arrdiv32_mux2to1383_and1;
  wire f_arrdiv32_mux2to1383_xor0;
  wire f_arrdiv32_mux2to1384_and0;
  wire f_arrdiv32_mux2to1384_not0;
  wire f_arrdiv32_mux2to1384_and1;
  wire f_arrdiv32_mux2to1384_xor0;
  wire f_arrdiv32_mux2to1385_and0;
  wire f_arrdiv32_mux2to1385_not0;
  wire f_arrdiv32_mux2to1385_and1;
  wire f_arrdiv32_mux2to1385_xor0;
  wire f_arrdiv32_mux2to1386_and0;
  wire f_arrdiv32_mux2to1386_not0;
  wire f_arrdiv32_mux2to1386_and1;
  wire f_arrdiv32_mux2to1386_xor0;
  wire f_arrdiv32_mux2to1387_and0;
  wire f_arrdiv32_mux2to1387_not0;
  wire f_arrdiv32_mux2to1387_and1;
  wire f_arrdiv32_mux2to1387_xor0;
  wire f_arrdiv32_mux2to1388_and0;
  wire f_arrdiv32_mux2to1388_not0;
  wire f_arrdiv32_mux2to1388_and1;
  wire f_arrdiv32_mux2to1388_xor0;
  wire f_arrdiv32_mux2to1389_and0;
  wire f_arrdiv32_mux2to1389_not0;
  wire f_arrdiv32_mux2to1389_and1;
  wire f_arrdiv32_mux2to1389_xor0;
  wire f_arrdiv32_mux2to1390_and0;
  wire f_arrdiv32_mux2to1390_not0;
  wire f_arrdiv32_mux2to1390_and1;
  wire f_arrdiv32_mux2to1390_xor0;
  wire f_arrdiv32_mux2to1391_and0;
  wire f_arrdiv32_mux2to1391_not0;
  wire f_arrdiv32_mux2to1391_and1;
  wire f_arrdiv32_mux2to1391_xor0;
  wire f_arrdiv32_mux2to1392_and0;
  wire f_arrdiv32_mux2to1392_not0;
  wire f_arrdiv32_mux2to1392_and1;
  wire f_arrdiv32_mux2to1392_xor0;
  wire f_arrdiv32_mux2to1393_and0;
  wire f_arrdiv32_mux2to1393_not0;
  wire f_arrdiv32_mux2to1393_and1;
  wire f_arrdiv32_mux2to1393_xor0;
  wire f_arrdiv32_mux2to1394_and0;
  wire f_arrdiv32_mux2to1394_not0;
  wire f_arrdiv32_mux2to1394_and1;
  wire f_arrdiv32_mux2to1394_xor0;
  wire f_arrdiv32_mux2to1395_and0;
  wire f_arrdiv32_mux2to1395_not0;
  wire f_arrdiv32_mux2to1395_and1;
  wire f_arrdiv32_mux2to1395_xor0;
  wire f_arrdiv32_mux2to1396_and0;
  wire f_arrdiv32_mux2to1396_not0;
  wire f_arrdiv32_mux2to1396_and1;
  wire f_arrdiv32_mux2to1396_xor0;
  wire f_arrdiv32_mux2to1397_and0;
  wire f_arrdiv32_mux2to1397_not0;
  wire f_arrdiv32_mux2to1397_and1;
  wire f_arrdiv32_mux2to1397_xor0;
  wire f_arrdiv32_mux2to1398_and0;
  wire f_arrdiv32_mux2to1398_not0;
  wire f_arrdiv32_mux2to1398_and1;
  wire f_arrdiv32_mux2to1398_xor0;
  wire f_arrdiv32_mux2to1399_and0;
  wire f_arrdiv32_mux2to1399_not0;
  wire f_arrdiv32_mux2to1399_and1;
  wire f_arrdiv32_mux2to1399_xor0;
  wire f_arrdiv32_mux2to1400_and0;
  wire f_arrdiv32_mux2to1400_not0;
  wire f_arrdiv32_mux2to1400_and1;
  wire f_arrdiv32_mux2to1400_xor0;
  wire f_arrdiv32_mux2to1401_and0;
  wire f_arrdiv32_mux2to1401_not0;
  wire f_arrdiv32_mux2to1401_and1;
  wire f_arrdiv32_mux2to1401_xor0;
  wire f_arrdiv32_mux2to1402_and0;
  wire f_arrdiv32_mux2to1402_not0;
  wire f_arrdiv32_mux2to1402_and1;
  wire f_arrdiv32_mux2to1402_xor0;
  wire f_arrdiv32_not12;
  wire f_arrdiv32_fs416_xor0;
  wire f_arrdiv32_fs416_not0;
  wire f_arrdiv32_fs416_and0;
  wire f_arrdiv32_fs416_not1;
  wire f_arrdiv32_fs417_xor0;
  wire f_arrdiv32_fs417_not0;
  wire f_arrdiv32_fs417_and0;
  wire f_arrdiv32_fs417_xor1;
  wire f_arrdiv32_fs417_not1;
  wire f_arrdiv32_fs417_and1;
  wire f_arrdiv32_fs417_or0;
  wire f_arrdiv32_fs418_xor0;
  wire f_arrdiv32_fs418_not0;
  wire f_arrdiv32_fs418_and0;
  wire f_arrdiv32_fs418_xor1;
  wire f_arrdiv32_fs418_not1;
  wire f_arrdiv32_fs418_and1;
  wire f_arrdiv32_fs418_or0;
  wire f_arrdiv32_fs419_xor0;
  wire f_arrdiv32_fs419_not0;
  wire f_arrdiv32_fs419_and0;
  wire f_arrdiv32_fs419_xor1;
  wire f_arrdiv32_fs419_not1;
  wire f_arrdiv32_fs419_and1;
  wire f_arrdiv32_fs419_or0;
  wire f_arrdiv32_fs420_xor0;
  wire f_arrdiv32_fs420_not0;
  wire f_arrdiv32_fs420_and0;
  wire f_arrdiv32_fs420_xor1;
  wire f_arrdiv32_fs420_not1;
  wire f_arrdiv32_fs420_and1;
  wire f_arrdiv32_fs420_or0;
  wire f_arrdiv32_fs421_xor0;
  wire f_arrdiv32_fs421_not0;
  wire f_arrdiv32_fs421_and0;
  wire f_arrdiv32_fs421_xor1;
  wire f_arrdiv32_fs421_not1;
  wire f_arrdiv32_fs421_and1;
  wire f_arrdiv32_fs421_or0;
  wire f_arrdiv32_fs422_xor0;
  wire f_arrdiv32_fs422_not0;
  wire f_arrdiv32_fs422_and0;
  wire f_arrdiv32_fs422_xor1;
  wire f_arrdiv32_fs422_not1;
  wire f_arrdiv32_fs422_and1;
  wire f_arrdiv32_fs422_or0;
  wire f_arrdiv32_fs423_xor0;
  wire f_arrdiv32_fs423_not0;
  wire f_arrdiv32_fs423_and0;
  wire f_arrdiv32_fs423_xor1;
  wire f_arrdiv32_fs423_not1;
  wire f_arrdiv32_fs423_and1;
  wire f_arrdiv32_fs423_or0;
  wire f_arrdiv32_fs424_xor0;
  wire f_arrdiv32_fs424_not0;
  wire f_arrdiv32_fs424_and0;
  wire f_arrdiv32_fs424_xor1;
  wire f_arrdiv32_fs424_not1;
  wire f_arrdiv32_fs424_and1;
  wire f_arrdiv32_fs424_or0;
  wire f_arrdiv32_fs425_xor0;
  wire f_arrdiv32_fs425_not0;
  wire f_arrdiv32_fs425_and0;
  wire f_arrdiv32_fs425_xor1;
  wire f_arrdiv32_fs425_not1;
  wire f_arrdiv32_fs425_and1;
  wire f_arrdiv32_fs425_or0;
  wire f_arrdiv32_fs426_xor0;
  wire f_arrdiv32_fs426_not0;
  wire f_arrdiv32_fs426_and0;
  wire f_arrdiv32_fs426_xor1;
  wire f_arrdiv32_fs426_not1;
  wire f_arrdiv32_fs426_and1;
  wire f_arrdiv32_fs426_or0;
  wire f_arrdiv32_fs427_xor0;
  wire f_arrdiv32_fs427_not0;
  wire f_arrdiv32_fs427_and0;
  wire f_arrdiv32_fs427_xor1;
  wire f_arrdiv32_fs427_not1;
  wire f_arrdiv32_fs427_and1;
  wire f_arrdiv32_fs427_or0;
  wire f_arrdiv32_fs428_xor0;
  wire f_arrdiv32_fs428_not0;
  wire f_arrdiv32_fs428_and0;
  wire f_arrdiv32_fs428_xor1;
  wire f_arrdiv32_fs428_not1;
  wire f_arrdiv32_fs428_and1;
  wire f_arrdiv32_fs428_or0;
  wire f_arrdiv32_fs429_xor0;
  wire f_arrdiv32_fs429_not0;
  wire f_arrdiv32_fs429_and0;
  wire f_arrdiv32_fs429_xor1;
  wire f_arrdiv32_fs429_not1;
  wire f_arrdiv32_fs429_and1;
  wire f_arrdiv32_fs429_or0;
  wire f_arrdiv32_fs430_xor0;
  wire f_arrdiv32_fs430_not0;
  wire f_arrdiv32_fs430_and0;
  wire f_arrdiv32_fs430_xor1;
  wire f_arrdiv32_fs430_not1;
  wire f_arrdiv32_fs430_and1;
  wire f_arrdiv32_fs430_or0;
  wire f_arrdiv32_fs431_xor0;
  wire f_arrdiv32_fs431_not0;
  wire f_arrdiv32_fs431_and0;
  wire f_arrdiv32_fs431_xor1;
  wire f_arrdiv32_fs431_not1;
  wire f_arrdiv32_fs431_and1;
  wire f_arrdiv32_fs431_or0;
  wire f_arrdiv32_fs432_xor0;
  wire f_arrdiv32_fs432_not0;
  wire f_arrdiv32_fs432_and0;
  wire f_arrdiv32_fs432_xor1;
  wire f_arrdiv32_fs432_not1;
  wire f_arrdiv32_fs432_and1;
  wire f_arrdiv32_fs432_or0;
  wire f_arrdiv32_fs433_xor0;
  wire f_arrdiv32_fs433_not0;
  wire f_arrdiv32_fs433_and0;
  wire f_arrdiv32_fs433_xor1;
  wire f_arrdiv32_fs433_not1;
  wire f_arrdiv32_fs433_and1;
  wire f_arrdiv32_fs433_or0;
  wire f_arrdiv32_fs434_xor0;
  wire f_arrdiv32_fs434_not0;
  wire f_arrdiv32_fs434_and0;
  wire f_arrdiv32_fs434_xor1;
  wire f_arrdiv32_fs434_not1;
  wire f_arrdiv32_fs434_and1;
  wire f_arrdiv32_fs434_or0;
  wire f_arrdiv32_fs435_xor0;
  wire f_arrdiv32_fs435_not0;
  wire f_arrdiv32_fs435_and0;
  wire f_arrdiv32_fs435_xor1;
  wire f_arrdiv32_fs435_not1;
  wire f_arrdiv32_fs435_and1;
  wire f_arrdiv32_fs435_or0;
  wire f_arrdiv32_fs436_xor0;
  wire f_arrdiv32_fs436_not0;
  wire f_arrdiv32_fs436_and0;
  wire f_arrdiv32_fs436_xor1;
  wire f_arrdiv32_fs436_not1;
  wire f_arrdiv32_fs436_and1;
  wire f_arrdiv32_fs436_or0;
  wire f_arrdiv32_fs437_xor0;
  wire f_arrdiv32_fs437_not0;
  wire f_arrdiv32_fs437_and0;
  wire f_arrdiv32_fs437_xor1;
  wire f_arrdiv32_fs437_not1;
  wire f_arrdiv32_fs437_and1;
  wire f_arrdiv32_fs437_or0;
  wire f_arrdiv32_fs438_xor0;
  wire f_arrdiv32_fs438_not0;
  wire f_arrdiv32_fs438_and0;
  wire f_arrdiv32_fs438_xor1;
  wire f_arrdiv32_fs438_not1;
  wire f_arrdiv32_fs438_and1;
  wire f_arrdiv32_fs438_or0;
  wire f_arrdiv32_fs439_xor0;
  wire f_arrdiv32_fs439_not0;
  wire f_arrdiv32_fs439_and0;
  wire f_arrdiv32_fs439_xor1;
  wire f_arrdiv32_fs439_not1;
  wire f_arrdiv32_fs439_and1;
  wire f_arrdiv32_fs439_or0;
  wire f_arrdiv32_fs440_xor0;
  wire f_arrdiv32_fs440_not0;
  wire f_arrdiv32_fs440_and0;
  wire f_arrdiv32_fs440_xor1;
  wire f_arrdiv32_fs440_not1;
  wire f_arrdiv32_fs440_and1;
  wire f_arrdiv32_fs440_or0;
  wire f_arrdiv32_fs441_xor0;
  wire f_arrdiv32_fs441_not0;
  wire f_arrdiv32_fs441_and0;
  wire f_arrdiv32_fs441_xor1;
  wire f_arrdiv32_fs441_not1;
  wire f_arrdiv32_fs441_and1;
  wire f_arrdiv32_fs441_or0;
  wire f_arrdiv32_fs442_xor0;
  wire f_arrdiv32_fs442_not0;
  wire f_arrdiv32_fs442_and0;
  wire f_arrdiv32_fs442_xor1;
  wire f_arrdiv32_fs442_not1;
  wire f_arrdiv32_fs442_and1;
  wire f_arrdiv32_fs442_or0;
  wire f_arrdiv32_fs443_xor0;
  wire f_arrdiv32_fs443_not0;
  wire f_arrdiv32_fs443_and0;
  wire f_arrdiv32_fs443_xor1;
  wire f_arrdiv32_fs443_not1;
  wire f_arrdiv32_fs443_and1;
  wire f_arrdiv32_fs443_or0;
  wire f_arrdiv32_fs444_xor0;
  wire f_arrdiv32_fs444_not0;
  wire f_arrdiv32_fs444_and0;
  wire f_arrdiv32_fs444_xor1;
  wire f_arrdiv32_fs444_not1;
  wire f_arrdiv32_fs444_and1;
  wire f_arrdiv32_fs444_or0;
  wire f_arrdiv32_fs445_xor0;
  wire f_arrdiv32_fs445_not0;
  wire f_arrdiv32_fs445_and0;
  wire f_arrdiv32_fs445_xor1;
  wire f_arrdiv32_fs445_not1;
  wire f_arrdiv32_fs445_and1;
  wire f_arrdiv32_fs445_or0;
  wire f_arrdiv32_fs446_xor0;
  wire f_arrdiv32_fs446_not0;
  wire f_arrdiv32_fs446_and0;
  wire f_arrdiv32_fs446_xor1;
  wire f_arrdiv32_fs446_not1;
  wire f_arrdiv32_fs446_and1;
  wire f_arrdiv32_fs446_or0;
  wire f_arrdiv32_fs447_xor0;
  wire f_arrdiv32_fs447_not0;
  wire f_arrdiv32_fs447_and0;
  wire f_arrdiv32_fs447_xor1;
  wire f_arrdiv32_fs447_not1;
  wire f_arrdiv32_fs447_and1;
  wire f_arrdiv32_fs447_or0;
  wire f_arrdiv32_mux2to1403_and0;
  wire f_arrdiv32_mux2to1403_not0;
  wire f_arrdiv32_mux2to1403_and1;
  wire f_arrdiv32_mux2to1403_xor0;
  wire f_arrdiv32_mux2to1404_and0;
  wire f_arrdiv32_mux2to1404_not0;
  wire f_arrdiv32_mux2to1404_and1;
  wire f_arrdiv32_mux2to1404_xor0;
  wire f_arrdiv32_mux2to1405_and0;
  wire f_arrdiv32_mux2to1405_not0;
  wire f_arrdiv32_mux2to1405_and1;
  wire f_arrdiv32_mux2to1405_xor0;
  wire f_arrdiv32_mux2to1406_and0;
  wire f_arrdiv32_mux2to1406_not0;
  wire f_arrdiv32_mux2to1406_and1;
  wire f_arrdiv32_mux2to1406_xor0;
  wire f_arrdiv32_mux2to1407_and0;
  wire f_arrdiv32_mux2to1407_not0;
  wire f_arrdiv32_mux2to1407_and1;
  wire f_arrdiv32_mux2to1407_xor0;
  wire f_arrdiv32_mux2to1408_and0;
  wire f_arrdiv32_mux2to1408_not0;
  wire f_arrdiv32_mux2to1408_and1;
  wire f_arrdiv32_mux2to1408_xor0;
  wire f_arrdiv32_mux2to1409_and0;
  wire f_arrdiv32_mux2to1409_not0;
  wire f_arrdiv32_mux2to1409_and1;
  wire f_arrdiv32_mux2to1409_xor0;
  wire f_arrdiv32_mux2to1410_and0;
  wire f_arrdiv32_mux2to1410_not0;
  wire f_arrdiv32_mux2to1410_and1;
  wire f_arrdiv32_mux2to1410_xor0;
  wire f_arrdiv32_mux2to1411_and0;
  wire f_arrdiv32_mux2to1411_not0;
  wire f_arrdiv32_mux2to1411_and1;
  wire f_arrdiv32_mux2to1411_xor0;
  wire f_arrdiv32_mux2to1412_and0;
  wire f_arrdiv32_mux2to1412_not0;
  wire f_arrdiv32_mux2to1412_and1;
  wire f_arrdiv32_mux2to1412_xor0;
  wire f_arrdiv32_mux2to1413_and0;
  wire f_arrdiv32_mux2to1413_not0;
  wire f_arrdiv32_mux2to1413_and1;
  wire f_arrdiv32_mux2to1413_xor0;
  wire f_arrdiv32_mux2to1414_and0;
  wire f_arrdiv32_mux2to1414_not0;
  wire f_arrdiv32_mux2to1414_and1;
  wire f_arrdiv32_mux2to1414_xor0;
  wire f_arrdiv32_mux2to1415_and0;
  wire f_arrdiv32_mux2to1415_not0;
  wire f_arrdiv32_mux2to1415_and1;
  wire f_arrdiv32_mux2to1415_xor0;
  wire f_arrdiv32_mux2to1416_and0;
  wire f_arrdiv32_mux2to1416_not0;
  wire f_arrdiv32_mux2to1416_and1;
  wire f_arrdiv32_mux2to1416_xor0;
  wire f_arrdiv32_mux2to1417_and0;
  wire f_arrdiv32_mux2to1417_not0;
  wire f_arrdiv32_mux2to1417_and1;
  wire f_arrdiv32_mux2to1417_xor0;
  wire f_arrdiv32_mux2to1418_and0;
  wire f_arrdiv32_mux2to1418_not0;
  wire f_arrdiv32_mux2to1418_and1;
  wire f_arrdiv32_mux2to1418_xor0;
  wire f_arrdiv32_mux2to1419_and0;
  wire f_arrdiv32_mux2to1419_not0;
  wire f_arrdiv32_mux2to1419_and1;
  wire f_arrdiv32_mux2to1419_xor0;
  wire f_arrdiv32_mux2to1420_and0;
  wire f_arrdiv32_mux2to1420_not0;
  wire f_arrdiv32_mux2to1420_and1;
  wire f_arrdiv32_mux2to1420_xor0;
  wire f_arrdiv32_mux2to1421_and0;
  wire f_arrdiv32_mux2to1421_not0;
  wire f_arrdiv32_mux2to1421_and1;
  wire f_arrdiv32_mux2to1421_xor0;
  wire f_arrdiv32_mux2to1422_and0;
  wire f_arrdiv32_mux2to1422_not0;
  wire f_arrdiv32_mux2to1422_and1;
  wire f_arrdiv32_mux2to1422_xor0;
  wire f_arrdiv32_mux2to1423_and0;
  wire f_arrdiv32_mux2to1423_not0;
  wire f_arrdiv32_mux2to1423_and1;
  wire f_arrdiv32_mux2to1423_xor0;
  wire f_arrdiv32_mux2to1424_and0;
  wire f_arrdiv32_mux2to1424_not0;
  wire f_arrdiv32_mux2to1424_and1;
  wire f_arrdiv32_mux2to1424_xor0;
  wire f_arrdiv32_mux2to1425_and0;
  wire f_arrdiv32_mux2to1425_not0;
  wire f_arrdiv32_mux2to1425_and1;
  wire f_arrdiv32_mux2to1425_xor0;
  wire f_arrdiv32_mux2to1426_and0;
  wire f_arrdiv32_mux2to1426_not0;
  wire f_arrdiv32_mux2to1426_and1;
  wire f_arrdiv32_mux2to1426_xor0;
  wire f_arrdiv32_mux2to1427_and0;
  wire f_arrdiv32_mux2to1427_not0;
  wire f_arrdiv32_mux2to1427_and1;
  wire f_arrdiv32_mux2to1427_xor0;
  wire f_arrdiv32_mux2to1428_and0;
  wire f_arrdiv32_mux2to1428_not0;
  wire f_arrdiv32_mux2to1428_and1;
  wire f_arrdiv32_mux2to1428_xor0;
  wire f_arrdiv32_mux2to1429_and0;
  wire f_arrdiv32_mux2to1429_not0;
  wire f_arrdiv32_mux2to1429_and1;
  wire f_arrdiv32_mux2to1429_xor0;
  wire f_arrdiv32_mux2to1430_and0;
  wire f_arrdiv32_mux2to1430_not0;
  wire f_arrdiv32_mux2to1430_and1;
  wire f_arrdiv32_mux2to1430_xor0;
  wire f_arrdiv32_mux2to1431_and0;
  wire f_arrdiv32_mux2to1431_not0;
  wire f_arrdiv32_mux2to1431_and1;
  wire f_arrdiv32_mux2to1431_xor0;
  wire f_arrdiv32_mux2to1432_and0;
  wire f_arrdiv32_mux2to1432_not0;
  wire f_arrdiv32_mux2to1432_and1;
  wire f_arrdiv32_mux2to1432_xor0;
  wire f_arrdiv32_mux2to1433_and0;
  wire f_arrdiv32_mux2to1433_not0;
  wire f_arrdiv32_mux2to1433_and1;
  wire f_arrdiv32_mux2to1433_xor0;
  wire f_arrdiv32_not13;
  wire f_arrdiv32_fs448_xor0;
  wire f_arrdiv32_fs448_not0;
  wire f_arrdiv32_fs448_and0;
  wire f_arrdiv32_fs448_not1;
  wire f_arrdiv32_fs449_xor0;
  wire f_arrdiv32_fs449_not0;
  wire f_arrdiv32_fs449_and0;
  wire f_arrdiv32_fs449_xor1;
  wire f_arrdiv32_fs449_not1;
  wire f_arrdiv32_fs449_and1;
  wire f_arrdiv32_fs449_or0;
  wire f_arrdiv32_fs450_xor0;
  wire f_arrdiv32_fs450_not0;
  wire f_arrdiv32_fs450_and0;
  wire f_arrdiv32_fs450_xor1;
  wire f_arrdiv32_fs450_not1;
  wire f_arrdiv32_fs450_and1;
  wire f_arrdiv32_fs450_or0;
  wire f_arrdiv32_fs451_xor0;
  wire f_arrdiv32_fs451_not0;
  wire f_arrdiv32_fs451_and0;
  wire f_arrdiv32_fs451_xor1;
  wire f_arrdiv32_fs451_not1;
  wire f_arrdiv32_fs451_and1;
  wire f_arrdiv32_fs451_or0;
  wire f_arrdiv32_fs452_xor0;
  wire f_arrdiv32_fs452_not0;
  wire f_arrdiv32_fs452_and0;
  wire f_arrdiv32_fs452_xor1;
  wire f_arrdiv32_fs452_not1;
  wire f_arrdiv32_fs452_and1;
  wire f_arrdiv32_fs452_or0;
  wire f_arrdiv32_fs453_xor0;
  wire f_arrdiv32_fs453_not0;
  wire f_arrdiv32_fs453_and0;
  wire f_arrdiv32_fs453_xor1;
  wire f_arrdiv32_fs453_not1;
  wire f_arrdiv32_fs453_and1;
  wire f_arrdiv32_fs453_or0;
  wire f_arrdiv32_fs454_xor0;
  wire f_arrdiv32_fs454_not0;
  wire f_arrdiv32_fs454_and0;
  wire f_arrdiv32_fs454_xor1;
  wire f_arrdiv32_fs454_not1;
  wire f_arrdiv32_fs454_and1;
  wire f_arrdiv32_fs454_or0;
  wire f_arrdiv32_fs455_xor0;
  wire f_arrdiv32_fs455_not0;
  wire f_arrdiv32_fs455_and0;
  wire f_arrdiv32_fs455_xor1;
  wire f_arrdiv32_fs455_not1;
  wire f_arrdiv32_fs455_and1;
  wire f_arrdiv32_fs455_or0;
  wire f_arrdiv32_fs456_xor0;
  wire f_arrdiv32_fs456_not0;
  wire f_arrdiv32_fs456_and0;
  wire f_arrdiv32_fs456_xor1;
  wire f_arrdiv32_fs456_not1;
  wire f_arrdiv32_fs456_and1;
  wire f_arrdiv32_fs456_or0;
  wire f_arrdiv32_fs457_xor0;
  wire f_arrdiv32_fs457_not0;
  wire f_arrdiv32_fs457_and0;
  wire f_arrdiv32_fs457_xor1;
  wire f_arrdiv32_fs457_not1;
  wire f_arrdiv32_fs457_and1;
  wire f_arrdiv32_fs457_or0;
  wire f_arrdiv32_fs458_xor0;
  wire f_arrdiv32_fs458_not0;
  wire f_arrdiv32_fs458_and0;
  wire f_arrdiv32_fs458_xor1;
  wire f_arrdiv32_fs458_not1;
  wire f_arrdiv32_fs458_and1;
  wire f_arrdiv32_fs458_or0;
  wire f_arrdiv32_fs459_xor0;
  wire f_arrdiv32_fs459_not0;
  wire f_arrdiv32_fs459_and0;
  wire f_arrdiv32_fs459_xor1;
  wire f_arrdiv32_fs459_not1;
  wire f_arrdiv32_fs459_and1;
  wire f_arrdiv32_fs459_or0;
  wire f_arrdiv32_fs460_xor0;
  wire f_arrdiv32_fs460_not0;
  wire f_arrdiv32_fs460_and0;
  wire f_arrdiv32_fs460_xor1;
  wire f_arrdiv32_fs460_not1;
  wire f_arrdiv32_fs460_and1;
  wire f_arrdiv32_fs460_or0;
  wire f_arrdiv32_fs461_xor0;
  wire f_arrdiv32_fs461_not0;
  wire f_arrdiv32_fs461_and0;
  wire f_arrdiv32_fs461_xor1;
  wire f_arrdiv32_fs461_not1;
  wire f_arrdiv32_fs461_and1;
  wire f_arrdiv32_fs461_or0;
  wire f_arrdiv32_fs462_xor0;
  wire f_arrdiv32_fs462_not0;
  wire f_arrdiv32_fs462_and0;
  wire f_arrdiv32_fs462_xor1;
  wire f_arrdiv32_fs462_not1;
  wire f_arrdiv32_fs462_and1;
  wire f_arrdiv32_fs462_or0;
  wire f_arrdiv32_fs463_xor0;
  wire f_arrdiv32_fs463_not0;
  wire f_arrdiv32_fs463_and0;
  wire f_arrdiv32_fs463_xor1;
  wire f_arrdiv32_fs463_not1;
  wire f_arrdiv32_fs463_and1;
  wire f_arrdiv32_fs463_or0;
  wire f_arrdiv32_fs464_xor0;
  wire f_arrdiv32_fs464_not0;
  wire f_arrdiv32_fs464_and0;
  wire f_arrdiv32_fs464_xor1;
  wire f_arrdiv32_fs464_not1;
  wire f_arrdiv32_fs464_and1;
  wire f_arrdiv32_fs464_or0;
  wire f_arrdiv32_fs465_xor0;
  wire f_arrdiv32_fs465_not0;
  wire f_arrdiv32_fs465_and0;
  wire f_arrdiv32_fs465_xor1;
  wire f_arrdiv32_fs465_not1;
  wire f_arrdiv32_fs465_and1;
  wire f_arrdiv32_fs465_or0;
  wire f_arrdiv32_fs466_xor0;
  wire f_arrdiv32_fs466_not0;
  wire f_arrdiv32_fs466_and0;
  wire f_arrdiv32_fs466_xor1;
  wire f_arrdiv32_fs466_not1;
  wire f_arrdiv32_fs466_and1;
  wire f_arrdiv32_fs466_or0;
  wire f_arrdiv32_fs467_xor0;
  wire f_arrdiv32_fs467_not0;
  wire f_arrdiv32_fs467_and0;
  wire f_arrdiv32_fs467_xor1;
  wire f_arrdiv32_fs467_not1;
  wire f_arrdiv32_fs467_and1;
  wire f_arrdiv32_fs467_or0;
  wire f_arrdiv32_fs468_xor0;
  wire f_arrdiv32_fs468_not0;
  wire f_arrdiv32_fs468_and0;
  wire f_arrdiv32_fs468_xor1;
  wire f_arrdiv32_fs468_not1;
  wire f_arrdiv32_fs468_and1;
  wire f_arrdiv32_fs468_or0;
  wire f_arrdiv32_fs469_xor0;
  wire f_arrdiv32_fs469_not0;
  wire f_arrdiv32_fs469_and0;
  wire f_arrdiv32_fs469_xor1;
  wire f_arrdiv32_fs469_not1;
  wire f_arrdiv32_fs469_and1;
  wire f_arrdiv32_fs469_or0;
  wire f_arrdiv32_fs470_xor0;
  wire f_arrdiv32_fs470_not0;
  wire f_arrdiv32_fs470_and0;
  wire f_arrdiv32_fs470_xor1;
  wire f_arrdiv32_fs470_not1;
  wire f_arrdiv32_fs470_and1;
  wire f_arrdiv32_fs470_or0;
  wire f_arrdiv32_fs471_xor0;
  wire f_arrdiv32_fs471_not0;
  wire f_arrdiv32_fs471_and0;
  wire f_arrdiv32_fs471_xor1;
  wire f_arrdiv32_fs471_not1;
  wire f_arrdiv32_fs471_and1;
  wire f_arrdiv32_fs471_or0;
  wire f_arrdiv32_fs472_xor0;
  wire f_arrdiv32_fs472_not0;
  wire f_arrdiv32_fs472_and0;
  wire f_arrdiv32_fs472_xor1;
  wire f_arrdiv32_fs472_not1;
  wire f_arrdiv32_fs472_and1;
  wire f_arrdiv32_fs472_or0;
  wire f_arrdiv32_fs473_xor0;
  wire f_arrdiv32_fs473_not0;
  wire f_arrdiv32_fs473_and0;
  wire f_arrdiv32_fs473_xor1;
  wire f_arrdiv32_fs473_not1;
  wire f_arrdiv32_fs473_and1;
  wire f_arrdiv32_fs473_or0;
  wire f_arrdiv32_fs474_xor0;
  wire f_arrdiv32_fs474_not0;
  wire f_arrdiv32_fs474_and0;
  wire f_arrdiv32_fs474_xor1;
  wire f_arrdiv32_fs474_not1;
  wire f_arrdiv32_fs474_and1;
  wire f_arrdiv32_fs474_or0;
  wire f_arrdiv32_fs475_xor0;
  wire f_arrdiv32_fs475_not0;
  wire f_arrdiv32_fs475_and0;
  wire f_arrdiv32_fs475_xor1;
  wire f_arrdiv32_fs475_not1;
  wire f_arrdiv32_fs475_and1;
  wire f_arrdiv32_fs475_or0;
  wire f_arrdiv32_fs476_xor0;
  wire f_arrdiv32_fs476_not0;
  wire f_arrdiv32_fs476_and0;
  wire f_arrdiv32_fs476_xor1;
  wire f_arrdiv32_fs476_not1;
  wire f_arrdiv32_fs476_and1;
  wire f_arrdiv32_fs476_or0;
  wire f_arrdiv32_fs477_xor0;
  wire f_arrdiv32_fs477_not0;
  wire f_arrdiv32_fs477_and0;
  wire f_arrdiv32_fs477_xor1;
  wire f_arrdiv32_fs477_not1;
  wire f_arrdiv32_fs477_and1;
  wire f_arrdiv32_fs477_or0;
  wire f_arrdiv32_fs478_xor0;
  wire f_arrdiv32_fs478_not0;
  wire f_arrdiv32_fs478_and0;
  wire f_arrdiv32_fs478_xor1;
  wire f_arrdiv32_fs478_not1;
  wire f_arrdiv32_fs478_and1;
  wire f_arrdiv32_fs478_or0;
  wire f_arrdiv32_fs479_xor0;
  wire f_arrdiv32_fs479_not0;
  wire f_arrdiv32_fs479_and0;
  wire f_arrdiv32_fs479_xor1;
  wire f_arrdiv32_fs479_not1;
  wire f_arrdiv32_fs479_and1;
  wire f_arrdiv32_fs479_or0;
  wire f_arrdiv32_mux2to1434_and0;
  wire f_arrdiv32_mux2to1434_not0;
  wire f_arrdiv32_mux2to1434_and1;
  wire f_arrdiv32_mux2to1434_xor0;
  wire f_arrdiv32_mux2to1435_and0;
  wire f_arrdiv32_mux2to1435_not0;
  wire f_arrdiv32_mux2to1435_and1;
  wire f_arrdiv32_mux2to1435_xor0;
  wire f_arrdiv32_mux2to1436_and0;
  wire f_arrdiv32_mux2to1436_not0;
  wire f_arrdiv32_mux2to1436_and1;
  wire f_arrdiv32_mux2to1436_xor0;
  wire f_arrdiv32_mux2to1437_and0;
  wire f_arrdiv32_mux2to1437_not0;
  wire f_arrdiv32_mux2to1437_and1;
  wire f_arrdiv32_mux2to1437_xor0;
  wire f_arrdiv32_mux2to1438_and0;
  wire f_arrdiv32_mux2to1438_not0;
  wire f_arrdiv32_mux2to1438_and1;
  wire f_arrdiv32_mux2to1438_xor0;
  wire f_arrdiv32_mux2to1439_and0;
  wire f_arrdiv32_mux2to1439_not0;
  wire f_arrdiv32_mux2to1439_and1;
  wire f_arrdiv32_mux2to1439_xor0;
  wire f_arrdiv32_mux2to1440_and0;
  wire f_arrdiv32_mux2to1440_not0;
  wire f_arrdiv32_mux2to1440_and1;
  wire f_arrdiv32_mux2to1440_xor0;
  wire f_arrdiv32_mux2to1441_and0;
  wire f_arrdiv32_mux2to1441_not0;
  wire f_arrdiv32_mux2to1441_and1;
  wire f_arrdiv32_mux2to1441_xor0;
  wire f_arrdiv32_mux2to1442_and0;
  wire f_arrdiv32_mux2to1442_not0;
  wire f_arrdiv32_mux2to1442_and1;
  wire f_arrdiv32_mux2to1442_xor0;
  wire f_arrdiv32_mux2to1443_and0;
  wire f_arrdiv32_mux2to1443_not0;
  wire f_arrdiv32_mux2to1443_and1;
  wire f_arrdiv32_mux2to1443_xor0;
  wire f_arrdiv32_mux2to1444_and0;
  wire f_arrdiv32_mux2to1444_not0;
  wire f_arrdiv32_mux2to1444_and1;
  wire f_arrdiv32_mux2to1444_xor0;
  wire f_arrdiv32_mux2to1445_and0;
  wire f_arrdiv32_mux2to1445_not0;
  wire f_arrdiv32_mux2to1445_and1;
  wire f_arrdiv32_mux2to1445_xor0;
  wire f_arrdiv32_mux2to1446_and0;
  wire f_arrdiv32_mux2to1446_not0;
  wire f_arrdiv32_mux2to1446_and1;
  wire f_arrdiv32_mux2to1446_xor0;
  wire f_arrdiv32_mux2to1447_and0;
  wire f_arrdiv32_mux2to1447_not0;
  wire f_arrdiv32_mux2to1447_and1;
  wire f_arrdiv32_mux2to1447_xor0;
  wire f_arrdiv32_mux2to1448_and0;
  wire f_arrdiv32_mux2to1448_not0;
  wire f_arrdiv32_mux2to1448_and1;
  wire f_arrdiv32_mux2to1448_xor0;
  wire f_arrdiv32_mux2to1449_and0;
  wire f_arrdiv32_mux2to1449_not0;
  wire f_arrdiv32_mux2to1449_and1;
  wire f_arrdiv32_mux2to1449_xor0;
  wire f_arrdiv32_mux2to1450_and0;
  wire f_arrdiv32_mux2to1450_not0;
  wire f_arrdiv32_mux2to1450_and1;
  wire f_arrdiv32_mux2to1450_xor0;
  wire f_arrdiv32_mux2to1451_and0;
  wire f_arrdiv32_mux2to1451_not0;
  wire f_arrdiv32_mux2to1451_and1;
  wire f_arrdiv32_mux2to1451_xor0;
  wire f_arrdiv32_mux2to1452_and0;
  wire f_arrdiv32_mux2to1452_not0;
  wire f_arrdiv32_mux2to1452_and1;
  wire f_arrdiv32_mux2to1452_xor0;
  wire f_arrdiv32_mux2to1453_and0;
  wire f_arrdiv32_mux2to1453_not0;
  wire f_arrdiv32_mux2to1453_and1;
  wire f_arrdiv32_mux2to1453_xor0;
  wire f_arrdiv32_mux2to1454_and0;
  wire f_arrdiv32_mux2to1454_not0;
  wire f_arrdiv32_mux2to1454_and1;
  wire f_arrdiv32_mux2to1454_xor0;
  wire f_arrdiv32_mux2to1455_and0;
  wire f_arrdiv32_mux2to1455_not0;
  wire f_arrdiv32_mux2to1455_and1;
  wire f_arrdiv32_mux2to1455_xor0;
  wire f_arrdiv32_mux2to1456_and0;
  wire f_arrdiv32_mux2to1456_not0;
  wire f_arrdiv32_mux2to1456_and1;
  wire f_arrdiv32_mux2to1456_xor0;
  wire f_arrdiv32_mux2to1457_and0;
  wire f_arrdiv32_mux2to1457_not0;
  wire f_arrdiv32_mux2to1457_and1;
  wire f_arrdiv32_mux2to1457_xor0;
  wire f_arrdiv32_mux2to1458_and0;
  wire f_arrdiv32_mux2to1458_not0;
  wire f_arrdiv32_mux2to1458_and1;
  wire f_arrdiv32_mux2to1458_xor0;
  wire f_arrdiv32_mux2to1459_and0;
  wire f_arrdiv32_mux2to1459_not0;
  wire f_arrdiv32_mux2to1459_and1;
  wire f_arrdiv32_mux2to1459_xor0;
  wire f_arrdiv32_mux2to1460_and0;
  wire f_arrdiv32_mux2to1460_not0;
  wire f_arrdiv32_mux2to1460_and1;
  wire f_arrdiv32_mux2to1460_xor0;
  wire f_arrdiv32_mux2to1461_and0;
  wire f_arrdiv32_mux2to1461_not0;
  wire f_arrdiv32_mux2to1461_and1;
  wire f_arrdiv32_mux2to1461_xor0;
  wire f_arrdiv32_mux2to1462_and0;
  wire f_arrdiv32_mux2to1462_not0;
  wire f_arrdiv32_mux2to1462_and1;
  wire f_arrdiv32_mux2to1462_xor0;
  wire f_arrdiv32_mux2to1463_and0;
  wire f_arrdiv32_mux2to1463_not0;
  wire f_arrdiv32_mux2to1463_and1;
  wire f_arrdiv32_mux2to1463_xor0;
  wire f_arrdiv32_mux2to1464_and0;
  wire f_arrdiv32_mux2to1464_not0;
  wire f_arrdiv32_mux2to1464_and1;
  wire f_arrdiv32_mux2to1464_xor0;
  wire f_arrdiv32_not14;
  wire f_arrdiv32_fs480_xor0;
  wire f_arrdiv32_fs480_not0;
  wire f_arrdiv32_fs480_and0;
  wire f_arrdiv32_fs480_not1;
  wire f_arrdiv32_fs481_xor0;
  wire f_arrdiv32_fs481_not0;
  wire f_arrdiv32_fs481_and0;
  wire f_arrdiv32_fs481_xor1;
  wire f_arrdiv32_fs481_not1;
  wire f_arrdiv32_fs481_and1;
  wire f_arrdiv32_fs481_or0;
  wire f_arrdiv32_fs482_xor0;
  wire f_arrdiv32_fs482_not0;
  wire f_arrdiv32_fs482_and0;
  wire f_arrdiv32_fs482_xor1;
  wire f_arrdiv32_fs482_not1;
  wire f_arrdiv32_fs482_and1;
  wire f_arrdiv32_fs482_or0;
  wire f_arrdiv32_fs483_xor0;
  wire f_arrdiv32_fs483_not0;
  wire f_arrdiv32_fs483_and0;
  wire f_arrdiv32_fs483_xor1;
  wire f_arrdiv32_fs483_not1;
  wire f_arrdiv32_fs483_and1;
  wire f_arrdiv32_fs483_or0;
  wire f_arrdiv32_fs484_xor0;
  wire f_arrdiv32_fs484_not0;
  wire f_arrdiv32_fs484_and0;
  wire f_arrdiv32_fs484_xor1;
  wire f_arrdiv32_fs484_not1;
  wire f_arrdiv32_fs484_and1;
  wire f_arrdiv32_fs484_or0;
  wire f_arrdiv32_fs485_xor0;
  wire f_arrdiv32_fs485_not0;
  wire f_arrdiv32_fs485_and0;
  wire f_arrdiv32_fs485_xor1;
  wire f_arrdiv32_fs485_not1;
  wire f_arrdiv32_fs485_and1;
  wire f_arrdiv32_fs485_or0;
  wire f_arrdiv32_fs486_xor0;
  wire f_arrdiv32_fs486_not0;
  wire f_arrdiv32_fs486_and0;
  wire f_arrdiv32_fs486_xor1;
  wire f_arrdiv32_fs486_not1;
  wire f_arrdiv32_fs486_and1;
  wire f_arrdiv32_fs486_or0;
  wire f_arrdiv32_fs487_xor0;
  wire f_arrdiv32_fs487_not0;
  wire f_arrdiv32_fs487_and0;
  wire f_arrdiv32_fs487_xor1;
  wire f_arrdiv32_fs487_not1;
  wire f_arrdiv32_fs487_and1;
  wire f_arrdiv32_fs487_or0;
  wire f_arrdiv32_fs488_xor0;
  wire f_arrdiv32_fs488_not0;
  wire f_arrdiv32_fs488_and0;
  wire f_arrdiv32_fs488_xor1;
  wire f_arrdiv32_fs488_not1;
  wire f_arrdiv32_fs488_and1;
  wire f_arrdiv32_fs488_or0;
  wire f_arrdiv32_fs489_xor0;
  wire f_arrdiv32_fs489_not0;
  wire f_arrdiv32_fs489_and0;
  wire f_arrdiv32_fs489_xor1;
  wire f_arrdiv32_fs489_not1;
  wire f_arrdiv32_fs489_and1;
  wire f_arrdiv32_fs489_or0;
  wire f_arrdiv32_fs490_xor0;
  wire f_arrdiv32_fs490_not0;
  wire f_arrdiv32_fs490_and0;
  wire f_arrdiv32_fs490_xor1;
  wire f_arrdiv32_fs490_not1;
  wire f_arrdiv32_fs490_and1;
  wire f_arrdiv32_fs490_or0;
  wire f_arrdiv32_fs491_xor0;
  wire f_arrdiv32_fs491_not0;
  wire f_arrdiv32_fs491_and0;
  wire f_arrdiv32_fs491_xor1;
  wire f_arrdiv32_fs491_not1;
  wire f_arrdiv32_fs491_and1;
  wire f_arrdiv32_fs491_or0;
  wire f_arrdiv32_fs492_xor0;
  wire f_arrdiv32_fs492_not0;
  wire f_arrdiv32_fs492_and0;
  wire f_arrdiv32_fs492_xor1;
  wire f_arrdiv32_fs492_not1;
  wire f_arrdiv32_fs492_and1;
  wire f_arrdiv32_fs492_or0;
  wire f_arrdiv32_fs493_xor0;
  wire f_arrdiv32_fs493_not0;
  wire f_arrdiv32_fs493_and0;
  wire f_arrdiv32_fs493_xor1;
  wire f_arrdiv32_fs493_not1;
  wire f_arrdiv32_fs493_and1;
  wire f_arrdiv32_fs493_or0;
  wire f_arrdiv32_fs494_xor0;
  wire f_arrdiv32_fs494_not0;
  wire f_arrdiv32_fs494_and0;
  wire f_arrdiv32_fs494_xor1;
  wire f_arrdiv32_fs494_not1;
  wire f_arrdiv32_fs494_and1;
  wire f_arrdiv32_fs494_or0;
  wire f_arrdiv32_fs495_xor0;
  wire f_arrdiv32_fs495_not0;
  wire f_arrdiv32_fs495_and0;
  wire f_arrdiv32_fs495_xor1;
  wire f_arrdiv32_fs495_not1;
  wire f_arrdiv32_fs495_and1;
  wire f_arrdiv32_fs495_or0;
  wire f_arrdiv32_fs496_xor0;
  wire f_arrdiv32_fs496_not0;
  wire f_arrdiv32_fs496_and0;
  wire f_arrdiv32_fs496_xor1;
  wire f_arrdiv32_fs496_not1;
  wire f_arrdiv32_fs496_and1;
  wire f_arrdiv32_fs496_or0;
  wire f_arrdiv32_fs497_xor0;
  wire f_arrdiv32_fs497_not0;
  wire f_arrdiv32_fs497_and0;
  wire f_arrdiv32_fs497_xor1;
  wire f_arrdiv32_fs497_not1;
  wire f_arrdiv32_fs497_and1;
  wire f_arrdiv32_fs497_or0;
  wire f_arrdiv32_fs498_xor0;
  wire f_arrdiv32_fs498_not0;
  wire f_arrdiv32_fs498_and0;
  wire f_arrdiv32_fs498_xor1;
  wire f_arrdiv32_fs498_not1;
  wire f_arrdiv32_fs498_and1;
  wire f_arrdiv32_fs498_or0;
  wire f_arrdiv32_fs499_xor0;
  wire f_arrdiv32_fs499_not0;
  wire f_arrdiv32_fs499_and0;
  wire f_arrdiv32_fs499_xor1;
  wire f_arrdiv32_fs499_not1;
  wire f_arrdiv32_fs499_and1;
  wire f_arrdiv32_fs499_or0;
  wire f_arrdiv32_fs500_xor0;
  wire f_arrdiv32_fs500_not0;
  wire f_arrdiv32_fs500_and0;
  wire f_arrdiv32_fs500_xor1;
  wire f_arrdiv32_fs500_not1;
  wire f_arrdiv32_fs500_and1;
  wire f_arrdiv32_fs500_or0;
  wire f_arrdiv32_fs501_xor0;
  wire f_arrdiv32_fs501_not0;
  wire f_arrdiv32_fs501_and0;
  wire f_arrdiv32_fs501_xor1;
  wire f_arrdiv32_fs501_not1;
  wire f_arrdiv32_fs501_and1;
  wire f_arrdiv32_fs501_or0;
  wire f_arrdiv32_fs502_xor0;
  wire f_arrdiv32_fs502_not0;
  wire f_arrdiv32_fs502_and0;
  wire f_arrdiv32_fs502_xor1;
  wire f_arrdiv32_fs502_not1;
  wire f_arrdiv32_fs502_and1;
  wire f_arrdiv32_fs502_or0;
  wire f_arrdiv32_fs503_xor0;
  wire f_arrdiv32_fs503_not0;
  wire f_arrdiv32_fs503_and0;
  wire f_arrdiv32_fs503_xor1;
  wire f_arrdiv32_fs503_not1;
  wire f_arrdiv32_fs503_and1;
  wire f_arrdiv32_fs503_or0;
  wire f_arrdiv32_fs504_xor0;
  wire f_arrdiv32_fs504_not0;
  wire f_arrdiv32_fs504_and0;
  wire f_arrdiv32_fs504_xor1;
  wire f_arrdiv32_fs504_not1;
  wire f_arrdiv32_fs504_and1;
  wire f_arrdiv32_fs504_or0;
  wire f_arrdiv32_fs505_xor0;
  wire f_arrdiv32_fs505_not0;
  wire f_arrdiv32_fs505_and0;
  wire f_arrdiv32_fs505_xor1;
  wire f_arrdiv32_fs505_not1;
  wire f_arrdiv32_fs505_and1;
  wire f_arrdiv32_fs505_or0;
  wire f_arrdiv32_fs506_xor0;
  wire f_arrdiv32_fs506_not0;
  wire f_arrdiv32_fs506_and0;
  wire f_arrdiv32_fs506_xor1;
  wire f_arrdiv32_fs506_not1;
  wire f_arrdiv32_fs506_and1;
  wire f_arrdiv32_fs506_or0;
  wire f_arrdiv32_fs507_xor0;
  wire f_arrdiv32_fs507_not0;
  wire f_arrdiv32_fs507_and0;
  wire f_arrdiv32_fs507_xor1;
  wire f_arrdiv32_fs507_not1;
  wire f_arrdiv32_fs507_and1;
  wire f_arrdiv32_fs507_or0;
  wire f_arrdiv32_fs508_xor0;
  wire f_arrdiv32_fs508_not0;
  wire f_arrdiv32_fs508_and0;
  wire f_arrdiv32_fs508_xor1;
  wire f_arrdiv32_fs508_not1;
  wire f_arrdiv32_fs508_and1;
  wire f_arrdiv32_fs508_or0;
  wire f_arrdiv32_fs509_xor0;
  wire f_arrdiv32_fs509_not0;
  wire f_arrdiv32_fs509_and0;
  wire f_arrdiv32_fs509_xor1;
  wire f_arrdiv32_fs509_not1;
  wire f_arrdiv32_fs509_and1;
  wire f_arrdiv32_fs509_or0;
  wire f_arrdiv32_fs510_xor0;
  wire f_arrdiv32_fs510_not0;
  wire f_arrdiv32_fs510_and0;
  wire f_arrdiv32_fs510_xor1;
  wire f_arrdiv32_fs510_not1;
  wire f_arrdiv32_fs510_and1;
  wire f_arrdiv32_fs510_or0;
  wire f_arrdiv32_fs511_xor0;
  wire f_arrdiv32_fs511_not0;
  wire f_arrdiv32_fs511_and0;
  wire f_arrdiv32_fs511_xor1;
  wire f_arrdiv32_fs511_not1;
  wire f_arrdiv32_fs511_and1;
  wire f_arrdiv32_fs511_or0;
  wire f_arrdiv32_mux2to1465_and0;
  wire f_arrdiv32_mux2to1465_not0;
  wire f_arrdiv32_mux2to1465_and1;
  wire f_arrdiv32_mux2to1465_xor0;
  wire f_arrdiv32_mux2to1466_and0;
  wire f_arrdiv32_mux2to1466_not0;
  wire f_arrdiv32_mux2to1466_and1;
  wire f_arrdiv32_mux2to1466_xor0;
  wire f_arrdiv32_mux2to1467_and0;
  wire f_arrdiv32_mux2to1467_not0;
  wire f_arrdiv32_mux2to1467_and1;
  wire f_arrdiv32_mux2to1467_xor0;
  wire f_arrdiv32_mux2to1468_and0;
  wire f_arrdiv32_mux2to1468_not0;
  wire f_arrdiv32_mux2to1468_and1;
  wire f_arrdiv32_mux2to1468_xor0;
  wire f_arrdiv32_mux2to1469_and0;
  wire f_arrdiv32_mux2to1469_not0;
  wire f_arrdiv32_mux2to1469_and1;
  wire f_arrdiv32_mux2to1469_xor0;
  wire f_arrdiv32_mux2to1470_and0;
  wire f_arrdiv32_mux2to1470_not0;
  wire f_arrdiv32_mux2to1470_and1;
  wire f_arrdiv32_mux2to1470_xor0;
  wire f_arrdiv32_mux2to1471_and0;
  wire f_arrdiv32_mux2to1471_not0;
  wire f_arrdiv32_mux2to1471_and1;
  wire f_arrdiv32_mux2to1471_xor0;
  wire f_arrdiv32_mux2to1472_and0;
  wire f_arrdiv32_mux2to1472_not0;
  wire f_arrdiv32_mux2to1472_and1;
  wire f_arrdiv32_mux2to1472_xor0;
  wire f_arrdiv32_mux2to1473_and0;
  wire f_arrdiv32_mux2to1473_not0;
  wire f_arrdiv32_mux2to1473_and1;
  wire f_arrdiv32_mux2to1473_xor0;
  wire f_arrdiv32_mux2to1474_and0;
  wire f_arrdiv32_mux2to1474_not0;
  wire f_arrdiv32_mux2to1474_and1;
  wire f_arrdiv32_mux2to1474_xor0;
  wire f_arrdiv32_mux2to1475_and0;
  wire f_arrdiv32_mux2to1475_not0;
  wire f_arrdiv32_mux2to1475_and1;
  wire f_arrdiv32_mux2to1475_xor0;
  wire f_arrdiv32_mux2to1476_and0;
  wire f_arrdiv32_mux2to1476_not0;
  wire f_arrdiv32_mux2to1476_and1;
  wire f_arrdiv32_mux2to1476_xor0;
  wire f_arrdiv32_mux2to1477_and0;
  wire f_arrdiv32_mux2to1477_not0;
  wire f_arrdiv32_mux2to1477_and1;
  wire f_arrdiv32_mux2to1477_xor0;
  wire f_arrdiv32_mux2to1478_and0;
  wire f_arrdiv32_mux2to1478_not0;
  wire f_arrdiv32_mux2to1478_and1;
  wire f_arrdiv32_mux2to1478_xor0;
  wire f_arrdiv32_mux2to1479_and0;
  wire f_arrdiv32_mux2to1479_not0;
  wire f_arrdiv32_mux2to1479_and1;
  wire f_arrdiv32_mux2to1479_xor0;
  wire f_arrdiv32_mux2to1480_and0;
  wire f_arrdiv32_mux2to1480_not0;
  wire f_arrdiv32_mux2to1480_and1;
  wire f_arrdiv32_mux2to1480_xor0;
  wire f_arrdiv32_mux2to1481_and0;
  wire f_arrdiv32_mux2to1481_not0;
  wire f_arrdiv32_mux2to1481_and1;
  wire f_arrdiv32_mux2to1481_xor0;
  wire f_arrdiv32_mux2to1482_and0;
  wire f_arrdiv32_mux2to1482_not0;
  wire f_arrdiv32_mux2to1482_and1;
  wire f_arrdiv32_mux2to1482_xor0;
  wire f_arrdiv32_mux2to1483_and0;
  wire f_arrdiv32_mux2to1483_not0;
  wire f_arrdiv32_mux2to1483_and1;
  wire f_arrdiv32_mux2to1483_xor0;
  wire f_arrdiv32_mux2to1484_and0;
  wire f_arrdiv32_mux2to1484_not0;
  wire f_arrdiv32_mux2to1484_and1;
  wire f_arrdiv32_mux2to1484_xor0;
  wire f_arrdiv32_mux2to1485_and0;
  wire f_arrdiv32_mux2to1485_not0;
  wire f_arrdiv32_mux2to1485_and1;
  wire f_arrdiv32_mux2to1485_xor0;
  wire f_arrdiv32_mux2to1486_and0;
  wire f_arrdiv32_mux2to1486_not0;
  wire f_arrdiv32_mux2to1486_and1;
  wire f_arrdiv32_mux2to1486_xor0;
  wire f_arrdiv32_mux2to1487_and0;
  wire f_arrdiv32_mux2to1487_not0;
  wire f_arrdiv32_mux2to1487_and1;
  wire f_arrdiv32_mux2to1487_xor0;
  wire f_arrdiv32_mux2to1488_and0;
  wire f_arrdiv32_mux2to1488_not0;
  wire f_arrdiv32_mux2to1488_and1;
  wire f_arrdiv32_mux2to1488_xor0;
  wire f_arrdiv32_mux2to1489_and0;
  wire f_arrdiv32_mux2to1489_not0;
  wire f_arrdiv32_mux2to1489_and1;
  wire f_arrdiv32_mux2to1489_xor0;
  wire f_arrdiv32_mux2to1490_and0;
  wire f_arrdiv32_mux2to1490_not0;
  wire f_arrdiv32_mux2to1490_and1;
  wire f_arrdiv32_mux2to1490_xor0;
  wire f_arrdiv32_mux2to1491_and0;
  wire f_arrdiv32_mux2to1491_not0;
  wire f_arrdiv32_mux2to1491_and1;
  wire f_arrdiv32_mux2to1491_xor0;
  wire f_arrdiv32_mux2to1492_and0;
  wire f_arrdiv32_mux2to1492_not0;
  wire f_arrdiv32_mux2to1492_and1;
  wire f_arrdiv32_mux2to1492_xor0;
  wire f_arrdiv32_mux2to1493_and0;
  wire f_arrdiv32_mux2to1493_not0;
  wire f_arrdiv32_mux2to1493_and1;
  wire f_arrdiv32_mux2to1493_xor0;
  wire f_arrdiv32_mux2to1494_and0;
  wire f_arrdiv32_mux2to1494_not0;
  wire f_arrdiv32_mux2to1494_and1;
  wire f_arrdiv32_mux2to1494_xor0;
  wire f_arrdiv32_mux2to1495_and0;
  wire f_arrdiv32_mux2to1495_not0;
  wire f_arrdiv32_mux2to1495_and1;
  wire f_arrdiv32_mux2to1495_xor0;
  wire f_arrdiv32_not15;
  wire f_arrdiv32_fs512_xor0;
  wire f_arrdiv32_fs512_not0;
  wire f_arrdiv32_fs512_and0;
  wire f_arrdiv32_fs512_not1;
  wire f_arrdiv32_fs513_xor0;
  wire f_arrdiv32_fs513_not0;
  wire f_arrdiv32_fs513_and0;
  wire f_arrdiv32_fs513_xor1;
  wire f_arrdiv32_fs513_not1;
  wire f_arrdiv32_fs513_and1;
  wire f_arrdiv32_fs513_or0;
  wire f_arrdiv32_fs514_xor0;
  wire f_arrdiv32_fs514_not0;
  wire f_arrdiv32_fs514_and0;
  wire f_arrdiv32_fs514_xor1;
  wire f_arrdiv32_fs514_not1;
  wire f_arrdiv32_fs514_and1;
  wire f_arrdiv32_fs514_or0;
  wire f_arrdiv32_fs515_xor0;
  wire f_arrdiv32_fs515_not0;
  wire f_arrdiv32_fs515_and0;
  wire f_arrdiv32_fs515_xor1;
  wire f_arrdiv32_fs515_not1;
  wire f_arrdiv32_fs515_and1;
  wire f_arrdiv32_fs515_or0;
  wire f_arrdiv32_fs516_xor0;
  wire f_arrdiv32_fs516_not0;
  wire f_arrdiv32_fs516_and0;
  wire f_arrdiv32_fs516_xor1;
  wire f_arrdiv32_fs516_not1;
  wire f_arrdiv32_fs516_and1;
  wire f_arrdiv32_fs516_or0;
  wire f_arrdiv32_fs517_xor0;
  wire f_arrdiv32_fs517_not0;
  wire f_arrdiv32_fs517_and0;
  wire f_arrdiv32_fs517_xor1;
  wire f_arrdiv32_fs517_not1;
  wire f_arrdiv32_fs517_and1;
  wire f_arrdiv32_fs517_or0;
  wire f_arrdiv32_fs518_xor0;
  wire f_arrdiv32_fs518_not0;
  wire f_arrdiv32_fs518_and0;
  wire f_arrdiv32_fs518_xor1;
  wire f_arrdiv32_fs518_not1;
  wire f_arrdiv32_fs518_and1;
  wire f_arrdiv32_fs518_or0;
  wire f_arrdiv32_fs519_xor0;
  wire f_arrdiv32_fs519_not0;
  wire f_arrdiv32_fs519_and0;
  wire f_arrdiv32_fs519_xor1;
  wire f_arrdiv32_fs519_not1;
  wire f_arrdiv32_fs519_and1;
  wire f_arrdiv32_fs519_or0;
  wire f_arrdiv32_fs520_xor0;
  wire f_arrdiv32_fs520_not0;
  wire f_arrdiv32_fs520_and0;
  wire f_arrdiv32_fs520_xor1;
  wire f_arrdiv32_fs520_not1;
  wire f_arrdiv32_fs520_and1;
  wire f_arrdiv32_fs520_or0;
  wire f_arrdiv32_fs521_xor0;
  wire f_arrdiv32_fs521_not0;
  wire f_arrdiv32_fs521_and0;
  wire f_arrdiv32_fs521_xor1;
  wire f_arrdiv32_fs521_not1;
  wire f_arrdiv32_fs521_and1;
  wire f_arrdiv32_fs521_or0;
  wire f_arrdiv32_fs522_xor0;
  wire f_arrdiv32_fs522_not0;
  wire f_arrdiv32_fs522_and0;
  wire f_arrdiv32_fs522_xor1;
  wire f_arrdiv32_fs522_not1;
  wire f_arrdiv32_fs522_and1;
  wire f_arrdiv32_fs522_or0;
  wire f_arrdiv32_fs523_xor0;
  wire f_arrdiv32_fs523_not0;
  wire f_arrdiv32_fs523_and0;
  wire f_arrdiv32_fs523_xor1;
  wire f_arrdiv32_fs523_not1;
  wire f_arrdiv32_fs523_and1;
  wire f_arrdiv32_fs523_or0;
  wire f_arrdiv32_fs524_xor0;
  wire f_arrdiv32_fs524_not0;
  wire f_arrdiv32_fs524_and0;
  wire f_arrdiv32_fs524_xor1;
  wire f_arrdiv32_fs524_not1;
  wire f_arrdiv32_fs524_and1;
  wire f_arrdiv32_fs524_or0;
  wire f_arrdiv32_fs525_xor0;
  wire f_arrdiv32_fs525_not0;
  wire f_arrdiv32_fs525_and0;
  wire f_arrdiv32_fs525_xor1;
  wire f_arrdiv32_fs525_not1;
  wire f_arrdiv32_fs525_and1;
  wire f_arrdiv32_fs525_or0;
  wire f_arrdiv32_fs526_xor0;
  wire f_arrdiv32_fs526_not0;
  wire f_arrdiv32_fs526_and0;
  wire f_arrdiv32_fs526_xor1;
  wire f_arrdiv32_fs526_not1;
  wire f_arrdiv32_fs526_and1;
  wire f_arrdiv32_fs526_or0;
  wire f_arrdiv32_fs527_xor0;
  wire f_arrdiv32_fs527_not0;
  wire f_arrdiv32_fs527_and0;
  wire f_arrdiv32_fs527_xor1;
  wire f_arrdiv32_fs527_not1;
  wire f_arrdiv32_fs527_and1;
  wire f_arrdiv32_fs527_or0;
  wire f_arrdiv32_fs528_xor0;
  wire f_arrdiv32_fs528_not0;
  wire f_arrdiv32_fs528_and0;
  wire f_arrdiv32_fs528_xor1;
  wire f_arrdiv32_fs528_not1;
  wire f_arrdiv32_fs528_and1;
  wire f_arrdiv32_fs528_or0;
  wire f_arrdiv32_fs529_xor0;
  wire f_arrdiv32_fs529_not0;
  wire f_arrdiv32_fs529_and0;
  wire f_arrdiv32_fs529_xor1;
  wire f_arrdiv32_fs529_not1;
  wire f_arrdiv32_fs529_and1;
  wire f_arrdiv32_fs529_or0;
  wire f_arrdiv32_fs530_xor0;
  wire f_arrdiv32_fs530_not0;
  wire f_arrdiv32_fs530_and0;
  wire f_arrdiv32_fs530_xor1;
  wire f_arrdiv32_fs530_not1;
  wire f_arrdiv32_fs530_and1;
  wire f_arrdiv32_fs530_or0;
  wire f_arrdiv32_fs531_xor0;
  wire f_arrdiv32_fs531_not0;
  wire f_arrdiv32_fs531_and0;
  wire f_arrdiv32_fs531_xor1;
  wire f_arrdiv32_fs531_not1;
  wire f_arrdiv32_fs531_and1;
  wire f_arrdiv32_fs531_or0;
  wire f_arrdiv32_fs532_xor0;
  wire f_arrdiv32_fs532_not0;
  wire f_arrdiv32_fs532_and0;
  wire f_arrdiv32_fs532_xor1;
  wire f_arrdiv32_fs532_not1;
  wire f_arrdiv32_fs532_and1;
  wire f_arrdiv32_fs532_or0;
  wire f_arrdiv32_fs533_xor0;
  wire f_arrdiv32_fs533_not0;
  wire f_arrdiv32_fs533_and0;
  wire f_arrdiv32_fs533_xor1;
  wire f_arrdiv32_fs533_not1;
  wire f_arrdiv32_fs533_and1;
  wire f_arrdiv32_fs533_or0;
  wire f_arrdiv32_fs534_xor0;
  wire f_arrdiv32_fs534_not0;
  wire f_arrdiv32_fs534_and0;
  wire f_arrdiv32_fs534_xor1;
  wire f_arrdiv32_fs534_not1;
  wire f_arrdiv32_fs534_and1;
  wire f_arrdiv32_fs534_or0;
  wire f_arrdiv32_fs535_xor0;
  wire f_arrdiv32_fs535_not0;
  wire f_arrdiv32_fs535_and0;
  wire f_arrdiv32_fs535_xor1;
  wire f_arrdiv32_fs535_not1;
  wire f_arrdiv32_fs535_and1;
  wire f_arrdiv32_fs535_or0;
  wire f_arrdiv32_fs536_xor0;
  wire f_arrdiv32_fs536_not0;
  wire f_arrdiv32_fs536_and0;
  wire f_arrdiv32_fs536_xor1;
  wire f_arrdiv32_fs536_not1;
  wire f_arrdiv32_fs536_and1;
  wire f_arrdiv32_fs536_or0;
  wire f_arrdiv32_fs537_xor0;
  wire f_arrdiv32_fs537_not0;
  wire f_arrdiv32_fs537_and0;
  wire f_arrdiv32_fs537_xor1;
  wire f_arrdiv32_fs537_not1;
  wire f_arrdiv32_fs537_and1;
  wire f_arrdiv32_fs537_or0;
  wire f_arrdiv32_fs538_xor0;
  wire f_arrdiv32_fs538_not0;
  wire f_arrdiv32_fs538_and0;
  wire f_arrdiv32_fs538_xor1;
  wire f_arrdiv32_fs538_not1;
  wire f_arrdiv32_fs538_and1;
  wire f_arrdiv32_fs538_or0;
  wire f_arrdiv32_fs539_xor0;
  wire f_arrdiv32_fs539_not0;
  wire f_arrdiv32_fs539_and0;
  wire f_arrdiv32_fs539_xor1;
  wire f_arrdiv32_fs539_not1;
  wire f_arrdiv32_fs539_and1;
  wire f_arrdiv32_fs539_or0;
  wire f_arrdiv32_fs540_xor0;
  wire f_arrdiv32_fs540_not0;
  wire f_arrdiv32_fs540_and0;
  wire f_arrdiv32_fs540_xor1;
  wire f_arrdiv32_fs540_not1;
  wire f_arrdiv32_fs540_and1;
  wire f_arrdiv32_fs540_or0;
  wire f_arrdiv32_fs541_xor0;
  wire f_arrdiv32_fs541_not0;
  wire f_arrdiv32_fs541_and0;
  wire f_arrdiv32_fs541_xor1;
  wire f_arrdiv32_fs541_not1;
  wire f_arrdiv32_fs541_and1;
  wire f_arrdiv32_fs541_or0;
  wire f_arrdiv32_fs542_xor0;
  wire f_arrdiv32_fs542_not0;
  wire f_arrdiv32_fs542_and0;
  wire f_arrdiv32_fs542_xor1;
  wire f_arrdiv32_fs542_not1;
  wire f_arrdiv32_fs542_and1;
  wire f_arrdiv32_fs542_or0;
  wire f_arrdiv32_fs543_xor0;
  wire f_arrdiv32_fs543_not0;
  wire f_arrdiv32_fs543_and0;
  wire f_arrdiv32_fs543_xor1;
  wire f_arrdiv32_fs543_not1;
  wire f_arrdiv32_fs543_and1;
  wire f_arrdiv32_fs543_or0;
  wire f_arrdiv32_mux2to1496_and0;
  wire f_arrdiv32_mux2to1496_not0;
  wire f_arrdiv32_mux2to1496_and1;
  wire f_arrdiv32_mux2to1496_xor0;
  wire f_arrdiv32_mux2to1497_and0;
  wire f_arrdiv32_mux2to1497_not0;
  wire f_arrdiv32_mux2to1497_and1;
  wire f_arrdiv32_mux2to1497_xor0;
  wire f_arrdiv32_mux2to1498_and0;
  wire f_arrdiv32_mux2to1498_not0;
  wire f_arrdiv32_mux2to1498_and1;
  wire f_arrdiv32_mux2to1498_xor0;
  wire f_arrdiv32_mux2to1499_and0;
  wire f_arrdiv32_mux2to1499_not0;
  wire f_arrdiv32_mux2to1499_and1;
  wire f_arrdiv32_mux2to1499_xor0;
  wire f_arrdiv32_mux2to1500_and0;
  wire f_arrdiv32_mux2to1500_not0;
  wire f_arrdiv32_mux2to1500_and1;
  wire f_arrdiv32_mux2to1500_xor0;
  wire f_arrdiv32_mux2to1501_and0;
  wire f_arrdiv32_mux2to1501_not0;
  wire f_arrdiv32_mux2to1501_and1;
  wire f_arrdiv32_mux2to1501_xor0;
  wire f_arrdiv32_mux2to1502_and0;
  wire f_arrdiv32_mux2to1502_not0;
  wire f_arrdiv32_mux2to1502_and1;
  wire f_arrdiv32_mux2to1502_xor0;
  wire f_arrdiv32_mux2to1503_and0;
  wire f_arrdiv32_mux2to1503_not0;
  wire f_arrdiv32_mux2to1503_and1;
  wire f_arrdiv32_mux2to1503_xor0;
  wire f_arrdiv32_mux2to1504_and0;
  wire f_arrdiv32_mux2to1504_not0;
  wire f_arrdiv32_mux2to1504_and1;
  wire f_arrdiv32_mux2to1504_xor0;
  wire f_arrdiv32_mux2to1505_and0;
  wire f_arrdiv32_mux2to1505_not0;
  wire f_arrdiv32_mux2to1505_and1;
  wire f_arrdiv32_mux2to1505_xor0;
  wire f_arrdiv32_mux2to1506_and0;
  wire f_arrdiv32_mux2to1506_not0;
  wire f_arrdiv32_mux2to1506_and1;
  wire f_arrdiv32_mux2to1506_xor0;
  wire f_arrdiv32_mux2to1507_and0;
  wire f_arrdiv32_mux2to1507_not0;
  wire f_arrdiv32_mux2to1507_and1;
  wire f_arrdiv32_mux2to1507_xor0;
  wire f_arrdiv32_mux2to1508_and0;
  wire f_arrdiv32_mux2to1508_not0;
  wire f_arrdiv32_mux2to1508_and1;
  wire f_arrdiv32_mux2to1508_xor0;
  wire f_arrdiv32_mux2to1509_and0;
  wire f_arrdiv32_mux2to1509_not0;
  wire f_arrdiv32_mux2to1509_and1;
  wire f_arrdiv32_mux2to1509_xor0;
  wire f_arrdiv32_mux2to1510_and0;
  wire f_arrdiv32_mux2to1510_not0;
  wire f_arrdiv32_mux2to1510_and1;
  wire f_arrdiv32_mux2to1510_xor0;
  wire f_arrdiv32_mux2to1511_and0;
  wire f_arrdiv32_mux2to1511_not0;
  wire f_arrdiv32_mux2to1511_and1;
  wire f_arrdiv32_mux2to1511_xor0;
  wire f_arrdiv32_mux2to1512_and0;
  wire f_arrdiv32_mux2to1512_not0;
  wire f_arrdiv32_mux2to1512_and1;
  wire f_arrdiv32_mux2to1512_xor0;
  wire f_arrdiv32_mux2to1513_and0;
  wire f_arrdiv32_mux2to1513_not0;
  wire f_arrdiv32_mux2to1513_and1;
  wire f_arrdiv32_mux2to1513_xor0;
  wire f_arrdiv32_mux2to1514_and0;
  wire f_arrdiv32_mux2to1514_not0;
  wire f_arrdiv32_mux2to1514_and1;
  wire f_arrdiv32_mux2to1514_xor0;
  wire f_arrdiv32_mux2to1515_and0;
  wire f_arrdiv32_mux2to1515_not0;
  wire f_arrdiv32_mux2to1515_and1;
  wire f_arrdiv32_mux2to1515_xor0;
  wire f_arrdiv32_mux2to1516_and0;
  wire f_arrdiv32_mux2to1516_not0;
  wire f_arrdiv32_mux2to1516_and1;
  wire f_arrdiv32_mux2to1516_xor0;
  wire f_arrdiv32_mux2to1517_and0;
  wire f_arrdiv32_mux2to1517_not0;
  wire f_arrdiv32_mux2to1517_and1;
  wire f_arrdiv32_mux2to1517_xor0;
  wire f_arrdiv32_mux2to1518_and0;
  wire f_arrdiv32_mux2to1518_not0;
  wire f_arrdiv32_mux2to1518_and1;
  wire f_arrdiv32_mux2to1518_xor0;
  wire f_arrdiv32_mux2to1519_and0;
  wire f_arrdiv32_mux2to1519_not0;
  wire f_arrdiv32_mux2to1519_and1;
  wire f_arrdiv32_mux2to1519_xor0;
  wire f_arrdiv32_mux2to1520_and0;
  wire f_arrdiv32_mux2to1520_not0;
  wire f_arrdiv32_mux2to1520_and1;
  wire f_arrdiv32_mux2to1520_xor0;
  wire f_arrdiv32_mux2to1521_and0;
  wire f_arrdiv32_mux2to1521_not0;
  wire f_arrdiv32_mux2to1521_and1;
  wire f_arrdiv32_mux2to1521_xor0;
  wire f_arrdiv32_mux2to1522_and0;
  wire f_arrdiv32_mux2to1522_not0;
  wire f_arrdiv32_mux2to1522_and1;
  wire f_arrdiv32_mux2to1522_xor0;
  wire f_arrdiv32_mux2to1523_and0;
  wire f_arrdiv32_mux2to1523_not0;
  wire f_arrdiv32_mux2to1523_and1;
  wire f_arrdiv32_mux2to1523_xor0;
  wire f_arrdiv32_mux2to1524_and0;
  wire f_arrdiv32_mux2to1524_not0;
  wire f_arrdiv32_mux2to1524_and1;
  wire f_arrdiv32_mux2to1524_xor0;
  wire f_arrdiv32_mux2to1525_and0;
  wire f_arrdiv32_mux2to1525_not0;
  wire f_arrdiv32_mux2to1525_and1;
  wire f_arrdiv32_mux2to1525_xor0;
  wire f_arrdiv32_mux2to1526_and0;
  wire f_arrdiv32_mux2to1526_not0;
  wire f_arrdiv32_mux2to1526_and1;
  wire f_arrdiv32_mux2to1526_xor0;
  wire f_arrdiv32_not16;
  wire f_arrdiv32_fs544_xor0;
  wire f_arrdiv32_fs544_not0;
  wire f_arrdiv32_fs544_and0;
  wire f_arrdiv32_fs544_not1;
  wire f_arrdiv32_fs545_xor0;
  wire f_arrdiv32_fs545_not0;
  wire f_arrdiv32_fs545_and0;
  wire f_arrdiv32_fs545_xor1;
  wire f_arrdiv32_fs545_not1;
  wire f_arrdiv32_fs545_and1;
  wire f_arrdiv32_fs545_or0;
  wire f_arrdiv32_fs546_xor0;
  wire f_arrdiv32_fs546_not0;
  wire f_arrdiv32_fs546_and0;
  wire f_arrdiv32_fs546_xor1;
  wire f_arrdiv32_fs546_not1;
  wire f_arrdiv32_fs546_and1;
  wire f_arrdiv32_fs546_or0;
  wire f_arrdiv32_fs547_xor0;
  wire f_arrdiv32_fs547_not0;
  wire f_arrdiv32_fs547_and0;
  wire f_arrdiv32_fs547_xor1;
  wire f_arrdiv32_fs547_not1;
  wire f_arrdiv32_fs547_and1;
  wire f_arrdiv32_fs547_or0;
  wire f_arrdiv32_fs548_xor0;
  wire f_arrdiv32_fs548_not0;
  wire f_arrdiv32_fs548_and0;
  wire f_arrdiv32_fs548_xor1;
  wire f_arrdiv32_fs548_not1;
  wire f_arrdiv32_fs548_and1;
  wire f_arrdiv32_fs548_or0;
  wire f_arrdiv32_fs549_xor0;
  wire f_arrdiv32_fs549_not0;
  wire f_arrdiv32_fs549_and0;
  wire f_arrdiv32_fs549_xor1;
  wire f_arrdiv32_fs549_not1;
  wire f_arrdiv32_fs549_and1;
  wire f_arrdiv32_fs549_or0;
  wire f_arrdiv32_fs550_xor0;
  wire f_arrdiv32_fs550_not0;
  wire f_arrdiv32_fs550_and0;
  wire f_arrdiv32_fs550_xor1;
  wire f_arrdiv32_fs550_not1;
  wire f_arrdiv32_fs550_and1;
  wire f_arrdiv32_fs550_or0;
  wire f_arrdiv32_fs551_xor0;
  wire f_arrdiv32_fs551_not0;
  wire f_arrdiv32_fs551_and0;
  wire f_arrdiv32_fs551_xor1;
  wire f_arrdiv32_fs551_not1;
  wire f_arrdiv32_fs551_and1;
  wire f_arrdiv32_fs551_or0;
  wire f_arrdiv32_fs552_xor0;
  wire f_arrdiv32_fs552_not0;
  wire f_arrdiv32_fs552_and0;
  wire f_arrdiv32_fs552_xor1;
  wire f_arrdiv32_fs552_not1;
  wire f_arrdiv32_fs552_and1;
  wire f_arrdiv32_fs552_or0;
  wire f_arrdiv32_fs553_xor0;
  wire f_arrdiv32_fs553_not0;
  wire f_arrdiv32_fs553_and0;
  wire f_arrdiv32_fs553_xor1;
  wire f_arrdiv32_fs553_not1;
  wire f_arrdiv32_fs553_and1;
  wire f_arrdiv32_fs553_or0;
  wire f_arrdiv32_fs554_xor0;
  wire f_arrdiv32_fs554_not0;
  wire f_arrdiv32_fs554_and0;
  wire f_arrdiv32_fs554_xor1;
  wire f_arrdiv32_fs554_not1;
  wire f_arrdiv32_fs554_and1;
  wire f_arrdiv32_fs554_or0;
  wire f_arrdiv32_fs555_xor0;
  wire f_arrdiv32_fs555_not0;
  wire f_arrdiv32_fs555_and0;
  wire f_arrdiv32_fs555_xor1;
  wire f_arrdiv32_fs555_not1;
  wire f_arrdiv32_fs555_and1;
  wire f_arrdiv32_fs555_or0;
  wire f_arrdiv32_fs556_xor0;
  wire f_arrdiv32_fs556_not0;
  wire f_arrdiv32_fs556_and0;
  wire f_arrdiv32_fs556_xor1;
  wire f_arrdiv32_fs556_not1;
  wire f_arrdiv32_fs556_and1;
  wire f_arrdiv32_fs556_or0;
  wire f_arrdiv32_fs557_xor0;
  wire f_arrdiv32_fs557_not0;
  wire f_arrdiv32_fs557_and0;
  wire f_arrdiv32_fs557_xor1;
  wire f_arrdiv32_fs557_not1;
  wire f_arrdiv32_fs557_and1;
  wire f_arrdiv32_fs557_or0;
  wire f_arrdiv32_fs558_xor0;
  wire f_arrdiv32_fs558_not0;
  wire f_arrdiv32_fs558_and0;
  wire f_arrdiv32_fs558_xor1;
  wire f_arrdiv32_fs558_not1;
  wire f_arrdiv32_fs558_and1;
  wire f_arrdiv32_fs558_or0;
  wire f_arrdiv32_fs559_xor0;
  wire f_arrdiv32_fs559_not0;
  wire f_arrdiv32_fs559_and0;
  wire f_arrdiv32_fs559_xor1;
  wire f_arrdiv32_fs559_not1;
  wire f_arrdiv32_fs559_and1;
  wire f_arrdiv32_fs559_or0;
  wire f_arrdiv32_fs560_xor0;
  wire f_arrdiv32_fs560_not0;
  wire f_arrdiv32_fs560_and0;
  wire f_arrdiv32_fs560_xor1;
  wire f_arrdiv32_fs560_not1;
  wire f_arrdiv32_fs560_and1;
  wire f_arrdiv32_fs560_or0;
  wire f_arrdiv32_fs561_xor0;
  wire f_arrdiv32_fs561_not0;
  wire f_arrdiv32_fs561_and0;
  wire f_arrdiv32_fs561_xor1;
  wire f_arrdiv32_fs561_not1;
  wire f_arrdiv32_fs561_and1;
  wire f_arrdiv32_fs561_or0;
  wire f_arrdiv32_fs562_xor0;
  wire f_arrdiv32_fs562_not0;
  wire f_arrdiv32_fs562_and0;
  wire f_arrdiv32_fs562_xor1;
  wire f_arrdiv32_fs562_not1;
  wire f_arrdiv32_fs562_and1;
  wire f_arrdiv32_fs562_or0;
  wire f_arrdiv32_fs563_xor0;
  wire f_arrdiv32_fs563_not0;
  wire f_arrdiv32_fs563_and0;
  wire f_arrdiv32_fs563_xor1;
  wire f_arrdiv32_fs563_not1;
  wire f_arrdiv32_fs563_and1;
  wire f_arrdiv32_fs563_or0;
  wire f_arrdiv32_fs564_xor0;
  wire f_arrdiv32_fs564_not0;
  wire f_arrdiv32_fs564_and0;
  wire f_arrdiv32_fs564_xor1;
  wire f_arrdiv32_fs564_not1;
  wire f_arrdiv32_fs564_and1;
  wire f_arrdiv32_fs564_or0;
  wire f_arrdiv32_fs565_xor0;
  wire f_arrdiv32_fs565_not0;
  wire f_arrdiv32_fs565_and0;
  wire f_arrdiv32_fs565_xor1;
  wire f_arrdiv32_fs565_not1;
  wire f_arrdiv32_fs565_and1;
  wire f_arrdiv32_fs565_or0;
  wire f_arrdiv32_fs566_xor0;
  wire f_arrdiv32_fs566_not0;
  wire f_arrdiv32_fs566_and0;
  wire f_arrdiv32_fs566_xor1;
  wire f_arrdiv32_fs566_not1;
  wire f_arrdiv32_fs566_and1;
  wire f_arrdiv32_fs566_or0;
  wire f_arrdiv32_fs567_xor0;
  wire f_arrdiv32_fs567_not0;
  wire f_arrdiv32_fs567_and0;
  wire f_arrdiv32_fs567_xor1;
  wire f_arrdiv32_fs567_not1;
  wire f_arrdiv32_fs567_and1;
  wire f_arrdiv32_fs567_or0;
  wire f_arrdiv32_fs568_xor0;
  wire f_arrdiv32_fs568_not0;
  wire f_arrdiv32_fs568_and0;
  wire f_arrdiv32_fs568_xor1;
  wire f_arrdiv32_fs568_not1;
  wire f_arrdiv32_fs568_and1;
  wire f_arrdiv32_fs568_or0;
  wire f_arrdiv32_fs569_xor0;
  wire f_arrdiv32_fs569_not0;
  wire f_arrdiv32_fs569_and0;
  wire f_arrdiv32_fs569_xor1;
  wire f_arrdiv32_fs569_not1;
  wire f_arrdiv32_fs569_and1;
  wire f_arrdiv32_fs569_or0;
  wire f_arrdiv32_fs570_xor0;
  wire f_arrdiv32_fs570_not0;
  wire f_arrdiv32_fs570_and0;
  wire f_arrdiv32_fs570_xor1;
  wire f_arrdiv32_fs570_not1;
  wire f_arrdiv32_fs570_and1;
  wire f_arrdiv32_fs570_or0;
  wire f_arrdiv32_fs571_xor0;
  wire f_arrdiv32_fs571_not0;
  wire f_arrdiv32_fs571_and0;
  wire f_arrdiv32_fs571_xor1;
  wire f_arrdiv32_fs571_not1;
  wire f_arrdiv32_fs571_and1;
  wire f_arrdiv32_fs571_or0;
  wire f_arrdiv32_fs572_xor0;
  wire f_arrdiv32_fs572_not0;
  wire f_arrdiv32_fs572_and0;
  wire f_arrdiv32_fs572_xor1;
  wire f_arrdiv32_fs572_not1;
  wire f_arrdiv32_fs572_and1;
  wire f_arrdiv32_fs572_or0;
  wire f_arrdiv32_fs573_xor0;
  wire f_arrdiv32_fs573_not0;
  wire f_arrdiv32_fs573_and0;
  wire f_arrdiv32_fs573_xor1;
  wire f_arrdiv32_fs573_not1;
  wire f_arrdiv32_fs573_and1;
  wire f_arrdiv32_fs573_or0;
  wire f_arrdiv32_fs574_xor0;
  wire f_arrdiv32_fs574_not0;
  wire f_arrdiv32_fs574_and0;
  wire f_arrdiv32_fs574_xor1;
  wire f_arrdiv32_fs574_not1;
  wire f_arrdiv32_fs574_and1;
  wire f_arrdiv32_fs574_or0;
  wire f_arrdiv32_fs575_xor0;
  wire f_arrdiv32_fs575_not0;
  wire f_arrdiv32_fs575_and0;
  wire f_arrdiv32_fs575_xor1;
  wire f_arrdiv32_fs575_not1;
  wire f_arrdiv32_fs575_and1;
  wire f_arrdiv32_fs575_or0;
  wire f_arrdiv32_mux2to1527_and0;
  wire f_arrdiv32_mux2to1527_not0;
  wire f_arrdiv32_mux2to1527_and1;
  wire f_arrdiv32_mux2to1527_xor0;
  wire f_arrdiv32_mux2to1528_and0;
  wire f_arrdiv32_mux2to1528_not0;
  wire f_arrdiv32_mux2to1528_and1;
  wire f_arrdiv32_mux2to1528_xor0;
  wire f_arrdiv32_mux2to1529_and0;
  wire f_arrdiv32_mux2to1529_not0;
  wire f_arrdiv32_mux2to1529_and1;
  wire f_arrdiv32_mux2to1529_xor0;
  wire f_arrdiv32_mux2to1530_and0;
  wire f_arrdiv32_mux2to1530_not0;
  wire f_arrdiv32_mux2to1530_and1;
  wire f_arrdiv32_mux2to1530_xor0;
  wire f_arrdiv32_mux2to1531_and0;
  wire f_arrdiv32_mux2to1531_not0;
  wire f_arrdiv32_mux2to1531_and1;
  wire f_arrdiv32_mux2to1531_xor0;
  wire f_arrdiv32_mux2to1532_and0;
  wire f_arrdiv32_mux2to1532_not0;
  wire f_arrdiv32_mux2to1532_and1;
  wire f_arrdiv32_mux2to1532_xor0;
  wire f_arrdiv32_mux2to1533_and0;
  wire f_arrdiv32_mux2to1533_not0;
  wire f_arrdiv32_mux2to1533_and1;
  wire f_arrdiv32_mux2to1533_xor0;
  wire f_arrdiv32_mux2to1534_and0;
  wire f_arrdiv32_mux2to1534_not0;
  wire f_arrdiv32_mux2to1534_and1;
  wire f_arrdiv32_mux2to1534_xor0;
  wire f_arrdiv32_mux2to1535_and0;
  wire f_arrdiv32_mux2to1535_not0;
  wire f_arrdiv32_mux2to1535_and1;
  wire f_arrdiv32_mux2to1535_xor0;
  wire f_arrdiv32_mux2to1536_and0;
  wire f_arrdiv32_mux2to1536_not0;
  wire f_arrdiv32_mux2to1536_and1;
  wire f_arrdiv32_mux2to1536_xor0;
  wire f_arrdiv32_mux2to1537_and0;
  wire f_arrdiv32_mux2to1537_not0;
  wire f_arrdiv32_mux2to1537_and1;
  wire f_arrdiv32_mux2to1537_xor0;
  wire f_arrdiv32_mux2to1538_and0;
  wire f_arrdiv32_mux2to1538_not0;
  wire f_arrdiv32_mux2to1538_and1;
  wire f_arrdiv32_mux2to1538_xor0;
  wire f_arrdiv32_mux2to1539_and0;
  wire f_arrdiv32_mux2to1539_not0;
  wire f_arrdiv32_mux2to1539_and1;
  wire f_arrdiv32_mux2to1539_xor0;
  wire f_arrdiv32_mux2to1540_and0;
  wire f_arrdiv32_mux2to1540_not0;
  wire f_arrdiv32_mux2to1540_and1;
  wire f_arrdiv32_mux2to1540_xor0;
  wire f_arrdiv32_mux2to1541_and0;
  wire f_arrdiv32_mux2to1541_not0;
  wire f_arrdiv32_mux2to1541_and1;
  wire f_arrdiv32_mux2to1541_xor0;
  wire f_arrdiv32_mux2to1542_and0;
  wire f_arrdiv32_mux2to1542_not0;
  wire f_arrdiv32_mux2to1542_and1;
  wire f_arrdiv32_mux2to1542_xor0;
  wire f_arrdiv32_mux2to1543_and0;
  wire f_arrdiv32_mux2to1543_not0;
  wire f_arrdiv32_mux2to1543_and1;
  wire f_arrdiv32_mux2to1543_xor0;
  wire f_arrdiv32_mux2to1544_and0;
  wire f_arrdiv32_mux2to1544_not0;
  wire f_arrdiv32_mux2to1544_and1;
  wire f_arrdiv32_mux2to1544_xor0;
  wire f_arrdiv32_mux2to1545_and0;
  wire f_arrdiv32_mux2to1545_not0;
  wire f_arrdiv32_mux2to1545_and1;
  wire f_arrdiv32_mux2to1545_xor0;
  wire f_arrdiv32_mux2to1546_and0;
  wire f_arrdiv32_mux2to1546_not0;
  wire f_arrdiv32_mux2to1546_and1;
  wire f_arrdiv32_mux2to1546_xor0;
  wire f_arrdiv32_mux2to1547_and0;
  wire f_arrdiv32_mux2to1547_not0;
  wire f_arrdiv32_mux2to1547_and1;
  wire f_arrdiv32_mux2to1547_xor0;
  wire f_arrdiv32_mux2to1548_and0;
  wire f_arrdiv32_mux2to1548_not0;
  wire f_arrdiv32_mux2to1548_and1;
  wire f_arrdiv32_mux2to1548_xor0;
  wire f_arrdiv32_mux2to1549_and0;
  wire f_arrdiv32_mux2to1549_not0;
  wire f_arrdiv32_mux2to1549_and1;
  wire f_arrdiv32_mux2to1549_xor0;
  wire f_arrdiv32_mux2to1550_and0;
  wire f_arrdiv32_mux2to1550_not0;
  wire f_arrdiv32_mux2to1550_and1;
  wire f_arrdiv32_mux2to1550_xor0;
  wire f_arrdiv32_mux2to1551_and0;
  wire f_arrdiv32_mux2to1551_not0;
  wire f_arrdiv32_mux2to1551_and1;
  wire f_arrdiv32_mux2to1551_xor0;
  wire f_arrdiv32_mux2to1552_and0;
  wire f_arrdiv32_mux2to1552_not0;
  wire f_arrdiv32_mux2to1552_and1;
  wire f_arrdiv32_mux2to1552_xor0;
  wire f_arrdiv32_mux2to1553_and0;
  wire f_arrdiv32_mux2to1553_not0;
  wire f_arrdiv32_mux2to1553_and1;
  wire f_arrdiv32_mux2to1553_xor0;
  wire f_arrdiv32_mux2to1554_and0;
  wire f_arrdiv32_mux2to1554_not0;
  wire f_arrdiv32_mux2to1554_and1;
  wire f_arrdiv32_mux2to1554_xor0;
  wire f_arrdiv32_mux2to1555_and0;
  wire f_arrdiv32_mux2to1555_not0;
  wire f_arrdiv32_mux2to1555_and1;
  wire f_arrdiv32_mux2to1555_xor0;
  wire f_arrdiv32_mux2to1556_and0;
  wire f_arrdiv32_mux2to1556_not0;
  wire f_arrdiv32_mux2to1556_and1;
  wire f_arrdiv32_mux2to1556_xor0;
  wire f_arrdiv32_mux2to1557_and0;
  wire f_arrdiv32_mux2to1557_not0;
  wire f_arrdiv32_mux2to1557_and1;
  wire f_arrdiv32_mux2to1557_xor0;
  wire f_arrdiv32_not17;
  wire f_arrdiv32_fs576_xor0;
  wire f_arrdiv32_fs576_not0;
  wire f_arrdiv32_fs576_and0;
  wire f_arrdiv32_fs576_not1;
  wire f_arrdiv32_fs577_xor0;
  wire f_arrdiv32_fs577_not0;
  wire f_arrdiv32_fs577_and0;
  wire f_arrdiv32_fs577_xor1;
  wire f_arrdiv32_fs577_not1;
  wire f_arrdiv32_fs577_and1;
  wire f_arrdiv32_fs577_or0;
  wire f_arrdiv32_fs578_xor0;
  wire f_arrdiv32_fs578_not0;
  wire f_arrdiv32_fs578_and0;
  wire f_arrdiv32_fs578_xor1;
  wire f_arrdiv32_fs578_not1;
  wire f_arrdiv32_fs578_and1;
  wire f_arrdiv32_fs578_or0;
  wire f_arrdiv32_fs579_xor0;
  wire f_arrdiv32_fs579_not0;
  wire f_arrdiv32_fs579_and0;
  wire f_arrdiv32_fs579_xor1;
  wire f_arrdiv32_fs579_not1;
  wire f_arrdiv32_fs579_and1;
  wire f_arrdiv32_fs579_or0;
  wire f_arrdiv32_fs580_xor0;
  wire f_arrdiv32_fs580_not0;
  wire f_arrdiv32_fs580_and0;
  wire f_arrdiv32_fs580_xor1;
  wire f_arrdiv32_fs580_not1;
  wire f_arrdiv32_fs580_and1;
  wire f_arrdiv32_fs580_or0;
  wire f_arrdiv32_fs581_xor0;
  wire f_arrdiv32_fs581_not0;
  wire f_arrdiv32_fs581_and0;
  wire f_arrdiv32_fs581_xor1;
  wire f_arrdiv32_fs581_not1;
  wire f_arrdiv32_fs581_and1;
  wire f_arrdiv32_fs581_or0;
  wire f_arrdiv32_fs582_xor0;
  wire f_arrdiv32_fs582_not0;
  wire f_arrdiv32_fs582_and0;
  wire f_arrdiv32_fs582_xor1;
  wire f_arrdiv32_fs582_not1;
  wire f_arrdiv32_fs582_and1;
  wire f_arrdiv32_fs582_or0;
  wire f_arrdiv32_fs583_xor0;
  wire f_arrdiv32_fs583_not0;
  wire f_arrdiv32_fs583_and0;
  wire f_arrdiv32_fs583_xor1;
  wire f_arrdiv32_fs583_not1;
  wire f_arrdiv32_fs583_and1;
  wire f_arrdiv32_fs583_or0;
  wire f_arrdiv32_fs584_xor0;
  wire f_arrdiv32_fs584_not0;
  wire f_arrdiv32_fs584_and0;
  wire f_arrdiv32_fs584_xor1;
  wire f_arrdiv32_fs584_not1;
  wire f_arrdiv32_fs584_and1;
  wire f_arrdiv32_fs584_or0;
  wire f_arrdiv32_fs585_xor0;
  wire f_arrdiv32_fs585_not0;
  wire f_arrdiv32_fs585_and0;
  wire f_arrdiv32_fs585_xor1;
  wire f_arrdiv32_fs585_not1;
  wire f_arrdiv32_fs585_and1;
  wire f_arrdiv32_fs585_or0;
  wire f_arrdiv32_fs586_xor0;
  wire f_arrdiv32_fs586_not0;
  wire f_arrdiv32_fs586_and0;
  wire f_arrdiv32_fs586_xor1;
  wire f_arrdiv32_fs586_not1;
  wire f_arrdiv32_fs586_and1;
  wire f_arrdiv32_fs586_or0;
  wire f_arrdiv32_fs587_xor0;
  wire f_arrdiv32_fs587_not0;
  wire f_arrdiv32_fs587_and0;
  wire f_arrdiv32_fs587_xor1;
  wire f_arrdiv32_fs587_not1;
  wire f_arrdiv32_fs587_and1;
  wire f_arrdiv32_fs587_or0;
  wire f_arrdiv32_fs588_xor0;
  wire f_arrdiv32_fs588_not0;
  wire f_arrdiv32_fs588_and0;
  wire f_arrdiv32_fs588_xor1;
  wire f_arrdiv32_fs588_not1;
  wire f_arrdiv32_fs588_and1;
  wire f_arrdiv32_fs588_or0;
  wire f_arrdiv32_fs589_xor0;
  wire f_arrdiv32_fs589_not0;
  wire f_arrdiv32_fs589_and0;
  wire f_arrdiv32_fs589_xor1;
  wire f_arrdiv32_fs589_not1;
  wire f_arrdiv32_fs589_and1;
  wire f_arrdiv32_fs589_or0;
  wire f_arrdiv32_fs590_xor0;
  wire f_arrdiv32_fs590_not0;
  wire f_arrdiv32_fs590_and0;
  wire f_arrdiv32_fs590_xor1;
  wire f_arrdiv32_fs590_not1;
  wire f_arrdiv32_fs590_and1;
  wire f_arrdiv32_fs590_or0;
  wire f_arrdiv32_fs591_xor0;
  wire f_arrdiv32_fs591_not0;
  wire f_arrdiv32_fs591_and0;
  wire f_arrdiv32_fs591_xor1;
  wire f_arrdiv32_fs591_not1;
  wire f_arrdiv32_fs591_and1;
  wire f_arrdiv32_fs591_or0;
  wire f_arrdiv32_fs592_xor0;
  wire f_arrdiv32_fs592_not0;
  wire f_arrdiv32_fs592_and0;
  wire f_arrdiv32_fs592_xor1;
  wire f_arrdiv32_fs592_not1;
  wire f_arrdiv32_fs592_and1;
  wire f_arrdiv32_fs592_or0;
  wire f_arrdiv32_fs593_xor0;
  wire f_arrdiv32_fs593_not0;
  wire f_arrdiv32_fs593_and0;
  wire f_arrdiv32_fs593_xor1;
  wire f_arrdiv32_fs593_not1;
  wire f_arrdiv32_fs593_and1;
  wire f_arrdiv32_fs593_or0;
  wire f_arrdiv32_fs594_xor0;
  wire f_arrdiv32_fs594_not0;
  wire f_arrdiv32_fs594_and0;
  wire f_arrdiv32_fs594_xor1;
  wire f_arrdiv32_fs594_not1;
  wire f_arrdiv32_fs594_and1;
  wire f_arrdiv32_fs594_or0;
  wire f_arrdiv32_fs595_xor0;
  wire f_arrdiv32_fs595_not0;
  wire f_arrdiv32_fs595_and0;
  wire f_arrdiv32_fs595_xor1;
  wire f_arrdiv32_fs595_not1;
  wire f_arrdiv32_fs595_and1;
  wire f_arrdiv32_fs595_or0;
  wire f_arrdiv32_fs596_xor0;
  wire f_arrdiv32_fs596_not0;
  wire f_arrdiv32_fs596_and0;
  wire f_arrdiv32_fs596_xor1;
  wire f_arrdiv32_fs596_not1;
  wire f_arrdiv32_fs596_and1;
  wire f_arrdiv32_fs596_or0;
  wire f_arrdiv32_fs597_xor0;
  wire f_arrdiv32_fs597_not0;
  wire f_arrdiv32_fs597_and0;
  wire f_arrdiv32_fs597_xor1;
  wire f_arrdiv32_fs597_not1;
  wire f_arrdiv32_fs597_and1;
  wire f_arrdiv32_fs597_or0;
  wire f_arrdiv32_fs598_xor0;
  wire f_arrdiv32_fs598_not0;
  wire f_arrdiv32_fs598_and0;
  wire f_arrdiv32_fs598_xor1;
  wire f_arrdiv32_fs598_not1;
  wire f_arrdiv32_fs598_and1;
  wire f_arrdiv32_fs598_or0;
  wire f_arrdiv32_fs599_xor0;
  wire f_arrdiv32_fs599_not0;
  wire f_arrdiv32_fs599_and0;
  wire f_arrdiv32_fs599_xor1;
  wire f_arrdiv32_fs599_not1;
  wire f_arrdiv32_fs599_and1;
  wire f_arrdiv32_fs599_or0;
  wire f_arrdiv32_fs600_xor0;
  wire f_arrdiv32_fs600_not0;
  wire f_arrdiv32_fs600_and0;
  wire f_arrdiv32_fs600_xor1;
  wire f_arrdiv32_fs600_not1;
  wire f_arrdiv32_fs600_and1;
  wire f_arrdiv32_fs600_or0;
  wire f_arrdiv32_fs601_xor0;
  wire f_arrdiv32_fs601_not0;
  wire f_arrdiv32_fs601_and0;
  wire f_arrdiv32_fs601_xor1;
  wire f_arrdiv32_fs601_not1;
  wire f_arrdiv32_fs601_and1;
  wire f_arrdiv32_fs601_or0;
  wire f_arrdiv32_fs602_xor0;
  wire f_arrdiv32_fs602_not0;
  wire f_arrdiv32_fs602_and0;
  wire f_arrdiv32_fs602_xor1;
  wire f_arrdiv32_fs602_not1;
  wire f_arrdiv32_fs602_and1;
  wire f_arrdiv32_fs602_or0;
  wire f_arrdiv32_fs603_xor0;
  wire f_arrdiv32_fs603_not0;
  wire f_arrdiv32_fs603_and0;
  wire f_arrdiv32_fs603_xor1;
  wire f_arrdiv32_fs603_not1;
  wire f_arrdiv32_fs603_and1;
  wire f_arrdiv32_fs603_or0;
  wire f_arrdiv32_fs604_xor0;
  wire f_arrdiv32_fs604_not0;
  wire f_arrdiv32_fs604_and0;
  wire f_arrdiv32_fs604_xor1;
  wire f_arrdiv32_fs604_not1;
  wire f_arrdiv32_fs604_and1;
  wire f_arrdiv32_fs604_or0;
  wire f_arrdiv32_fs605_xor0;
  wire f_arrdiv32_fs605_not0;
  wire f_arrdiv32_fs605_and0;
  wire f_arrdiv32_fs605_xor1;
  wire f_arrdiv32_fs605_not1;
  wire f_arrdiv32_fs605_and1;
  wire f_arrdiv32_fs605_or0;
  wire f_arrdiv32_fs606_xor0;
  wire f_arrdiv32_fs606_not0;
  wire f_arrdiv32_fs606_and0;
  wire f_arrdiv32_fs606_xor1;
  wire f_arrdiv32_fs606_not1;
  wire f_arrdiv32_fs606_and1;
  wire f_arrdiv32_fs606_or0;
  wire f_arrdiv32_fs607_xor0;
  wire f_arrdiv32_fs607_not0;
  wire f_arrdiv32_fs607_and0;
  wire f_arrdiv32_fs607_xor1;
  wire f_arrdiv32_fs607_not1;
  wire f_arrdiv32_fs607_and1;
  wire f_arrdiv32_fs607_or0;
  wire f_arrdiv32_mux2to1558_and0;
  wire f_arrdiv32_mux2to1558_not0;
  wire f_arrdiv32_mux2to1558_and1;
  wire f_arrdiv32_mux2to1558_xor0;
  wire f_arrdiv32_mux2to1559_and0;
  wire f_arrdiv32_mux2to1559_not0;
  wire f_arrdiv32_mux2to1559_and1;
  wire f_arrdiv32_mux2to1559_xor0;
  wire f_arrdiv32_mux2to1560_and0;
  wire f_arrdiv32_mux2to1560_not0;
  wire f_arrdiv32_mux2to1560_and1;
  wire f_arrdiv32_mux2to1560_xor0;
  wire f_arrdiv32_mux2to1561_and0;
  wire f_arrdiv32_mux2to1561_not0;
  wire f_arrdiv32_mux2to1561_and1;
  wire f_arrdiv32_mux2to1561_xor0;
  wire f_arrdiv32_mux2to1562_and0;
  wire f_arrdiv32_mux2to1562_not0;
  wire f_arrdiv32_mux2to1562_and1;
  wire f_arrdiv32_mux2to1562_xor0;
  wire f_arrdiv32_mux2to1563_and0;
  wire f_arrdiv32_mux2to1563_not0;
  wire f_arrdiv32_mux2to1563_and1;
  wire f_arrdiv32_mux2to1563_xor0;
  wire f_arrdiv32_mux2to1564_and0;
  wire f_arrdiv32_mux2to1564_not0;
  wire f_arrdiv32_mux2to1564_and1;
  wire f_arrdiv32_mux2to1564_xor0;
  wire f_arrdiv32_mux2to1565_and0;
  wire f_arrdiv32_mux2to1565_not0;
  wire f_arrdiv32_mux2to1565_and1;
  wire f_arrdiv32_mux2to1565_xor0;
  wire f_arrdiv32_mux2to1566_and0;
  wire f_arrdiv32_mux2to1566_not0;
  wire f_arrdiv32_mux2to1566_and1;
  wire f_arrdiv32_mux2to1566_xor0;
  wire f_arrdiv32_mux2to1567_and0;
  wire f_arrdiv32_mux2to1567_not0;
  wire f_arrdiv32_mux2to1567_and1;
  wire f_arrdiv32_mux2to1567_xor0;
  wire f_arrdiv32_mux2to1568_and0;
  wire f_arrdiv32_mux2to1568_not0;
  wire f_arrdiv32_mux2to1568_and1;
  wire f_arrdiv32_mux2to1568_xor0;
  wire f_arrdiv32_mux2to1569_and0;
  wire f_arrdiv32_mux2to1569_not0;
  wire f_arrdiv32_mux2to1569_and1;
  wire f_arrdiv32_mux2to1569_xor0;
  wire f_arrdiv32_mux2to1570_and0;
  wire f_arrdiv32_mux2to1570_not0;
  wire f_arrdiv32_mux2to1570_and1;
  wire f_arrdiv32_mux2to1570_xor0;
  wire f_arrdiv32_mux2to1571_and0;
  wire f_arrdiv32_mux2to1571_not0;
  wire f_arrdiv32_mux2to1571_and1;
  wire f_arrdiv32_mux2to1571_xor0;
  wire f_arrdiv32_mux2to1572_and0;
  wire f_arrdiv32_mux2to1572_not0;
  wire f_arrdiv32_mux2to1572_and1;
  wire f_arrdiv32_mux2to1572_xor0;
  wire f_arrdiv32_mux2to1573_and0;
  wire f_arrdiv32_mux2to1573_not0;
  wire f_arrdiv32_mux2to1573_and1;
  wire f_arrdiv32_mux2to1573_xor0;
  wire f_arrdiv32_mux2to1574_and0;
  wire f_arrdiv32_mux2to1574_not0;
  wire f_arrdiv32_mux2to1574_and1;
  wire f_arrdiv32_mux2to1574_xor0;
  wire f_arrdiv32_mux2to1575_and0;
  wire f_arrdiv32_mux2to1575_not0;
  wire f_arrdiv32_mux2to1575_and1;
  wire f_arrdiv32_mux2to1575_xor0;
  wire f_arrdiv32_mux2to1576_and0;
  wire f_arrdiv32_mux2to1576_not0;
  wire f_arrdiv32_mux2to1576_and1;
  wire f_arrdiv32_mux2to1576_xor0;
  wire f_arrdiv32_mux2to1577_and0;
  wire f_arrdiv32_mux2to1577_not0;
  wire f_arrdiv32_mux2to1577_and1;
  wire f_arrdiv32_mux2to1577_xor0;
  wire f_arrdiv32_mux2to1578_and0;
  wire f_arrdiv32_mux2to1578_not0;
  wire f_arrdiv32_mux2to1578_and1;
  wire f_arrdiv32_mux2to1578_xor0;
  wire f_arrdiv32_mux2to1579_and0;
  wire f_arrdiv32_mux2to1579_not0;
  wire f_arrdiv32_mux2to1579_and1;
  wire f_arrdiv32_mux2to1579_xor0;
  wire f_arrdiv32_mux2to1580_and0;
  wire f_arrdiv32_mux2to1580_not0;
  wire f_arrdiv32_mux2to1580_and1;
  wire f_arrdiv32_mux2to1580_xor0;
  wire f_arrdiv32_mux2to1581_and0;
  wire f_arrdiv32_mux2to1581_not0;
  wire f_arrdiv32_mux2to1581_and1;
  wire f_arrdiv32_mux2to1581_xor0;
  wire f_arrdiv32_mux2to1582_and0;
  wire f_arrdiv32_mux2to1582_not0;
  wire f_arrdiv32_mux2to1582_and1;
  wire f_arrdiv32_mux2to1582_xor0;
  wire f_arrdiv32_mux2to1583_and0;
  wire f_arrdiv32_mux2to1583_not0;
  wire f_arrdiv32_mux2to1583_and1;
  wire f_arrdiv32_mux2to1583_xor0;
  wire f_arrdiv32_mux2to1584_and0;
  wire f_arrdiv32_mux2to1584_not0;
  wire f_arrdiv32_mux2to1584_and1;
  wire f_arrdiv32_mux2to1584_xor0;
  wire f_arrdiv32_mux2to1585_and0;
  wire f_arrdiv32_mux2to1585_not0;
  wire f_arrdiv32_mux2to1585_and1;
  wire f_arrdiv32_mux2to1585_xor0;
  wire f_arrdiv32_mux2to1586_and0;
  wire f_arrdiv32_mux2to1586_not0;
  wire f_arrdiv32_mux2to1586_and1;
  wire f_arrdiv32_mux2to1586_xor0;
  wire f_arrdiv32_mux2to1587_and0;
  wire f_arrdiv32_mux2to1587_not0;
  wire f_arrdiv32_mux2to1587_and1;
  wire f_arrdiv32_mux2to1587_xor0;
  wire f_arrdiv32_mux2to1588_and0;
  wire f_arrdiv32_mux2to1588_not0;
  wire f_arrdiv32_mux2to1588_and1;
  wire f_arrdiv32_mux2to1588_xor0;
  wire f_arrdiv32_not18;
  wire f_arrdiv32_fs608_xor0;
  wire f_arrdiv32_fs608_not0;
  wire f_arrdiv32_fs608_and0;
  wire f_arrdiv32_fs608_not1;
  wire f_arrdiv32_fs609_xor0;
  wire f_arrdiv32_fs609_not0;
  wire f_arrdiv32_fs609_and0;
  wire f_arrdiv32_fs609_xor1;
  wire f_arrdiv32_fs609_not1;
  wire f_arrdiv32_fs609_and1;
  wire f_arrdiv32_fs609_or0;
  wire f_arrdiv32_fs610_xor0;
  wire f_arrdiv32_fs610_not0;
  wire f_arrdiv32_fs610_and0;
  wire f_arrdiv32_fs610_xor1;
  wire f_arrdiv32_fs610_not1;
  wire f_arrdiv32_fs610_and1;
  wire f_arrdiv32_fs610_or0;
  wire f_arrdiv32_fs611_xor0;
  wire f_arrdiv32_fs611_not0;
  wire f_arrdiv32_fs611_and0;
  wire f_arrdiv32_fs611_xor1;
  wire f_arrdiv32_fs611_not1;
  wire f_arrdiv32_fs611_and1;
  wire f_arrdiv32_fs611_or0;
  wire f_arrdiv32_fs612_xor0;
  wire f_arrdiv32_fs612_not0;
  wire f_arrdiv32_fs612_and0;
  wire f_arrdiv32_fs612_xor1;
  wire f_arrdiv32_fs612_not1;
  wire f_arrdiv32_fs612_and1;
  wire f_arrdiv32_fs612_or0;
  wire f_arrdiv32_fs613_xor0;
  wire f_arrdiv32_fs613_not0;
  wire f_arrdiv32_fs613_and0;
  wire f_arrdiv32_fs613_xor1;
  wire f_arrdiv32_fs613_not1;
  wire f_arrdiv32_fs613_and1;
  wire f_arrdiv32_fs613_or0;
  wire f_arrdiv32_fs614_xor0;
  wire f_arrdiv32_fs614_not0;
  wire f_arrdiv32_fs614_and0;
  wire f_arrdiv32_fs614_xor1;
  wire f_arrdiv32_fs614_not1;
  wire f_arrdiv32_fs614_and1;
  wire f_arrdiv32_fs614_or0;
  wire f_arrdiv32_fs615_xor0;
  wire f_arrdiv32_fs615_not0;
  wire f_arrdiv32_fs615_and0;
  wire f_arrdiv32_fs615_xor1;
  wire f_arrdiv32_fs615_not1;
  wire f_arrdiv32_fs615_and1;
  wire f_arrdiv32_fs615_or0;
  wire f_arrdiv32_fs616_xor0;
  wire f_arrdiv32_fs616_not0;
  wire f_arrdiv32_fs616_and0;
  wire f_arrdiv32_fs616_xor1;
  wire f_arrdiv32_fs616_not1;
  wire f_arrdiv32_fs616_and1;
  wire f_arrdiv32_fs616_or0;
  wire f_arrdiv32_fs617_xor0;
  wire f_arrdiv32_fs617_not0;
  wire f_arrdiv32_fs617_and0;
  wire f_arrdiv32_fs617_xor1;
  wire f_arrdiv32_fs617_not1;
  wire f_arrdiv32_fs617_and1;
  wire f_arrdiv32_fs617_or0;
  wire f_arrdiv32_fs618_xor0;
  wire f_arrdiv32_fs618_not0;
  wire f_arrdiv32_fs618_and0;
  wire f_arrdiv32_fs618_xor1;
  wire f_arrdiv32_fs618_not1;
  wire f_arrdiv32_fs618_and1;
  wire f_arrdiv32_fs618_or0;
  wire f_arrdiv32_fs619_xor0;
  wire f_arrdiv32_fs619_not0;
  wire f_arrdiv32_fs619_and0;
  wire f_arrdiv32_fs619_xor1;
  wire f_arrdiv32_fs619_not1;
  wire f_arrdiv32_fs619_and1;
  wire f_arrdiv32_fs619_or0;
  wire f_arrdiv32_fs620_xor0;
  wire f_arrdiv32_fs620_not0;
  wire f_arrdiv32_fs620_and0;
  wire f_arrdiv32_fs620_xor1;
  wire f_arrdiv32_fs620_not1;
  wire f_arrdiv32_fs620_and1;
  wire f_arrdiv32_fs620_or0;
  wire f_arrdiv32_fs621_xor0;
  wire f_arrdiv32_fs621_not0;
  wire f_arrdiv32_fs621_and0;
  wire f_arrdiv32_fs621_xor1;
  wire f_arrdiv32_fs621_not1;
  wire f_arrdiv32_fs621_and1;
  wire f_arrdiv32_fs621_or0;
  wire f_arrdiv32_fs622_xor0;
  wire f_arrdiv32_fs622_not0;
  wire f_arrdiv32_fs622_and0;
  wire f_arrdiv32_fs622_xor1;
  wire f_arrdiv32_fs622_not1;
  wire f_arrdiv32_fs622_and1;
  wire f_arrdiv32_fs622_or0;
  wire f_arrdiv32_fs623_xor0;
  wire f_arrdiv32_fs623_not0;
  wire f_arrdiv32_fs623_and0;
  wire f_arrdiv32_fs623_xor1;
  wire f_arrdiv32_fs623_not1;
  wire f_arrdiv32_fs623_and1;
  wire f_arrdiv32_fs623_or0;
  wire f_arrdiv32_fs624_xor0;
  wire f_arrdiv32_fs624_not0;
  wire f_arrdiv32_fs624_and0;
  wire f_arrdiv32_fs624_xor1;
  wire f_arrdiv32_fs624_not1;
  wire f_arrdiv32_fs624_and1;
  wire f_arrdiv32_fs624_or0;
  wire f_arrdiv32_fs625_xor0;
  wire f_arrdiv32_fs625_not0;
  wire f_arrdiv32_fs625_and0;
  wire f_arrdiv32_fs625_xor1;
  wire f_arrdiv32_fs625_not1;
  wire f_arrdiv32_fs625_and1;
  wire f_arrdiv32_fs625_or0;
  wire f_arrdiv32_fs626_xor0;
  wire f_arrdiv32_fs626_not0;
  wire f_arrdiv32_fs626_and0;
  wire f_arrdiv32_fs626_xor1;
  wire f_arrdiv32_fs626_not1;
  wire f_arrdiv32_fs626_and1;
  wire f_arrdiv32_fs626_or0;
  wire f_arrdiv32_fs627_xor0;
  wire f_arrdiv32_fs627_not0;
  wire f_arrdiv32_fs627_and0;
  wire f_arrdiv32_fs627_xor1;
  wire f_arrdiv32_fs627_not1;
  wire f_arrdiv32_fs627_and1;
  wire f_arrdiv32_fs627_or0;
  wire f_arrdiv32_fs628_xor0;
  wire f_arrdiv32_fs628_not0;
  wire f_arrdiv32_fs628_and0;
  wire f_arrdiv32_fs628_xor1;
  wire f_arrdiv32_fs628_not1;
  wire f_arrdiv32_fs628_and1;
  wire f_arrdiv32_fs628_or0;
  wire f_arrdiv32_fs629_xor0;
  wire f_arrdiv32_fs629_not0;
  wire f_arrdiv32_fs629_and0;
  wire f_arrdiv32_fs629_xor1;
  wire f_arrdiv32_fs629_not1;
  wire f_arrdiv32_fs629_and1;
  wire f_arrdiv32_fs629_or0;
  wire f_arrdiv32_fs630_xor0;
  wire f_arrdiv32_fs630_not0;
  wire f_arrdiv32_fs630_and0;
  wire f_arrdiv32_fs630_xor1;
  wire f_arrdiv32_fs630_not1;
  wire f_arrdiv32_fs630_and1;
  wire f_arrdiv32_fs630_or0;
  wire f_arrdiv32_fs631_xor0;
  wire f_arrdiv32_fs631_not0;
  wire f_arrdiv32_fs631_and0;
  wire f_arrdiv32_fs631_xor1;
  wire f_arrdiv32_fs631_not1;
  wire f_arrdiv32_fs631_and1;
  wire f_arrdiv32_fs631_or0;
  wire f_arrdiv32_fs632_xor0;
  wire f_arrdiv32_fs632_not0;
  wire f_arrdiv32_fs632_and0;
  wire f_arrdiv32_fs632_xor1;
  wire f_arrdiv32_fs632_not1;
  wire f_arrdiv32_fs632_and1;
  wire f_arrdiv32_fs632_or0;
  wire f_arrdiv32_fs633_xor0;
  wire f_arrdiv32_fs633_not0;
  wire f_arrdiv32_fs633_and0;
  wire f_arrdiv32_fs633_xor1;
  wire f_arrdiv32_fs633_not1;
  wire f_arrdiv32_fs633_and1;
  wire f_arrdiv32_fs633_or0;
  wire f_arrdiv32_fs634_xor0;
  wire f_arrdiv32_fs634_not0;
  wire f_arrdiv32_fs634_and0;
  wire f_arrdiv32_fs634_xor1;
  wire f_arrdiv32_fs634_not1;
  wire f_arrdiv32_fs634_and1;
  wire f_arrdiv32_fs634_or0;
  wire f_arrdiv32_fs635_xor0;
  wire f_arrdiv32_fs635_not0;
  wire f_arrdiv32_fs635_and0;
  wire f_arrdiv32_fs635_xor1;
  wire f_arrdiv32_fs635_not1;
  wire f_arrdiv32_fs635_and1;
  wire f_arrdiv32_fs635_or0;
  wire f_arrdiv32_fs636_xor0;
  wire f_arrdiv32_fs636_not0;
  wire f_arrdiv32_fs636_and0;
  wire f_arrdiv32_fs636_xor1;
  wire f_arrdiv32_fs636_not1;
  wire f_arrdiv32_fs636_and1;
  wire f_arrdiv32_fs636_or0;
  wire f_arrdiv32_fs637_xor0;
  wire f_arrdiv32_fs637_not0;
  wire f_arrdiv32_fs637_and0;
  wire f_arrdiv32_fs637_xor1;
  wire f_arrdiv32_fs637_not1;
  wire f_arrdiv32_fs637_and1;
  wire f_arrdiv32_fs637_or0;
  wire f_arrdiv32_fs638_xor0;
  wire f_arrdiv32_fs638_not0;
  wire f_arrdiv32_fs638_and0;
  wire f_arrdiv32_fs638_xor1;
  wire f_arrdiv32_fs638_not1;
  wire f_arrdiv32_fs638_and1;
  wire f_arrdiv32_fs638_or0;
  wire f_arrdiv32_fs639_xor0;
  wire f_arrdiv32_fs639_not0;
  wire f_arrdiv32_fs639_and0;
  wire f_arrdiv32_fs639_xor1;
  wire f_arrdiv32_fs639_not1;
  wire f_arrdiv32_fs639_and1;
  wire f_arrdiv32_fs639_or0;
  wire f_arrdiv32_mux2to1589_and0;
  wire f_arrdiv32_mux2to1589_not0;
  wire f_arrdiv32_mux2to1589_and1;
  wire f_arrdiv32_mux2to1589_xor0;
  wire f_arrdiv32_mux2to1590_and0;
  wire f_arrdiv32_mux2to1590_not0;
  wire f_arrdiv32_mux2to1590_and1;
  wire f_arrdiv32_mux2to1590_xor0;
  wire f_arrdiv32_mux2to1591_and0;
  wire f_arrdiv32_mux2to1591_not0;
  wire f_arrdiv32_mux2to1591_and1;
  wire f_arrdiv32_mux2to1591_xor0;
  wire f_arrdiv32_mux2to1592_and0;
  wire f_arrdiv32_mux2to1592_not0;
  wire f_arrdiv32_mux2to1592_and1;
  wire f_arrdiv32_mux2to1592_xor0;
  wire f_arrdiv32_mux2to1593_and0;
  wire f_arrdiv32_mux2to1593_not0;
  wire f_arrdiv32_mux2to1593_and1;
  wire f_arrdiv32_mux2to1593_xor0;
  wire f_arrdiv32_mux2to1594_and0;
  wire f_arrdiv32_mux2to1594_not0;
  wire f_arrdiv32_mux2to1594_and1;
  wire f_arrdiv32_mux2to1594_xor0;
  wire f_arrdiv32_mux2to1595_and0;
  wire f_arrdiv32_mux2to1595_not0;
  wire f_arrdiv32_mux2to1595_and1;
  wire f_arrdiv32_mux2to1595_xor0;
  wire f_arrdiv32_mux2to1596_and0;
  wire f_arrdiv32_mux2to1596_not0;
  wire f_arrdiv32_mux2to1596_and1;
  wire f_arrdiv32_mux2to1596_xor0;
  wire f_arrdiv32_mux2to1597_and0;
  wire f_arrdiv32_mux2to1597_not0;
  wire f_arrdiv32_mux2to1597_and1;
  wire f_arrdiv32_mux2to1597_xor0;
  wire f_arrdiv32_mux2to1598_and0;
  wire f_arrdiv32_mux2to1598_not0;
  wire f_arrdiv32_mux2to1598_and1;
  wire f_arrdiv32_mux2to1598_xor0;
  wire f_arrdiv32_mux2to1599_and0;
  wire f_arrdiv32_mux2to1599_not0;
  wire f_arrdiv32_mux2to1599_and1;
  wire f_arrdiv32_mux2to1599_xor0;
  wire f_arrdiv32_mux2to1600_and0;
  wire f_arrdiv32_mux2to1600_not0;
  wire f_arrdiv32_mux2to1600_and1;
  wire f_arrdiv32_mux2to1600_xor0;
  wire f_arrdiv32_mux2to1601_and0;
  wire f_arrdiv32_mux2to1601_not0;
  wire f_arrdiv32_mux2to1601_and1;
  wire f_arrdiv32_mux2to1601_xor0;
  wire f_arrdiv32_mux2to1602_and0;
  wire f_arrdiv32_mux2to1602_not0;
  wire f_arrdiv32_mux2to1602_and1;
  wire f_arrdiv32_mux2to1602_xor0;
  wire f_arrdiv32_mux2to1603_and0;
  wire f_arrdiv32_mux2to1603_not0;
  wire f_arrdiv32_mux2to1603_and1;
  wire f_arrdiv32_mux2to1603_xor0;
  wire f_arrdiv32_mux2to1604_and0;
  wire f_arrdiv32_mux2to1604_not0;
  wire f_arrdiv32_mux2to1604_and1;
  wire f_arrdiv32_mux2to1604_xor0;
  wire f_arrdiv32_mux2to1605_and0;
  wire f_arrdiv32_mux2to1605_not0;
  wire f_arrdiv32_mux2to1605_and1;
  wire f_arrdiv32_mux2to1605_xor0;
  wire f_arrdiv32_mux2to1606_and0;
  wire f_arrdiv32_mux2to1606_not0;
  wire f_arrdiv32_mux2to1606_and1;
  wire f_arrdiv32_mux2to1606_xor0;
  wire f_arrdiv32_mux2to1607_and0;
  wire f_arrdiv32_mux2to1607_not0;
  wire f_arrdiv32_mux2to1607_and1;
  wire f_arrdiv32_mux2to1607_xor0;
  wire f_arrdiv32_mux2to1608_and0;
  wire f_arrdiv32_mux2to1608_not0;
  wire f_arrdiv32_mux2to1608_and1;
  wire f_arrdiv32_mux2to1608_xor0;
  wire f_arrdiv32_mux2to1609_and0;
  wire f_arrdiv32_mux2to1609_not0;
  wire f_arrdiv32_mux2to1609_and1;
  wire f_arrdiv32_mux2to1609_xor0;
  wire f_arrdiv32_mux2to1610_and0;
  wire f_arrdiv32_mux2to1610_not0;
  wire f_arrdiv32_mux2to1610_and1;
  wire f_arrdiv32_mux2to1610_xor0;
  wire f_arrdiv32_mux2to1611_and0;
  wire f_arrdiv32_mux2to1611_not0;
  wire f_arrdiv32_mux2to1611_and1;
  wire f_arrdiv32_mux2to1611_xor0;
  wire f_arrdiv32_mux2to1612_and0;
  wire f_arrdiv32_mux2to1612_not0;
  wire f_arrdiv32_mux2to1612_and1;
  wire f_arrdiv32_mux2to1612_xor0;
  wire f_arrdiv32_mux2to1613_and0;
  wire f_arrdiv32_mux2to1613_not0;
  wire f_arrdiv32_mux2to1613_and1;
  wire f_arrdiv32_mux2to1613_xor0;
  wire f_arrdiv32_mux2to1614_and0;
  wire f_arrdiv32_mux2to1614_not0;
  wire f_arrdiv32_mux2to1614_and1;
  wire f_arrdiv32_mux2to1614_xor0;
  wire f_arrdiv32_mux2to1615_and0;
  wire f_arrdiv32_mux2to1615_not0;
  wire f_arrdiv32_mux2to1615_and1;
  wire f_arrdiv32_mux2to1615_xor0;
  wire f_arrdiv32_mux2to1616_and0;
  wire f_arrdiv32_mux2to1616_not0;
  wire f_arrdiv32_mux2to1616_and1;
  wire f_arrdiv32_mux2to1616_xor0;
  wire f_arrdiv32_mux2to1617_and0;
  wire f_arrdiv32_mux2to1617_not0;
  wire f_arrdiv32_mux2to1617_and1;
  wire f_arrdiv32_mux2to1617_xor0;
  wire f_arrdiv32_mux2to1618_and0;
  wire f_arrdiv32_mux2to1618_not0;
  wire f_arrdiv32_mux2to1618_and1;
  wire f_arrdiv32_mux2to1618_xor0;
  wire f_arrdiv32_mux2to1619_and0;
  wire f_arrdiv32_mux2to1619_not0;
  wire f_arrdiv32_mux2to1619_and1;
  wire f_arrdiv32_mux2to1619_xor0;
  wire f_arrdiv32_not19;
  wire f_arrdiv32_fs640_xor0;
  wire f_arrdiv32_fs640_not0;
  wire f_arrdiv32_fs640_and0;
  wire f_arrdiv32_fs640_not1;
  wire f_arrdiv32_fs641_xor0;
  wire f_arrdiv32_fs641_not0;
  wire f_arrdiv32_fs641_and0;
  wire f_arrdiv32_fs641_xor1;
  wire f_arrdiv32_fs641_not1;
  wire f_arrdiv32_fs641_and1;
  wire f_arrdiv32_fs641_or0;
  wire f_arrdiv32_fs642_xor0;
  wire f_arrdiv32_fs642_not0;
  wire f_arrdiv32_fs642_and0;
  wire f_arrdiv32_fs642_xor1;
  wire f_arrdiv32_fs642_not1;
  wire f_arrdiv32_fs642_and1;
  wire f_arrdiv32_fs642_or0;
  wire f_arrdiv32_fs643_xor0;
  wire f_arrdiv32_fs643_not0;
  wire f_arrdiv32_fs643_and0;
  wire f_arrdiv32_fs643_xor1;
  wire f_arrdiv32_fs643_not1;
  wire f_arrdiv32_fs643_and1;
  wire f_arrdiv32_fs643_or0;
  wire f_arrdiv32_fs644_xor0;
  wire f_arrdiv32_fs644_not0;
  wire f_arrdiv32_fs644_and0;
  wire f_arrdiv32_fs644_xor1;
  wire f_arrdiv32_fs644_not1;
  wire f_arrdiv32_fs644_and1;
  wire f_arrdiv32_fs644_or0;
  wire f_arrdiv32_fs645_xor0;
  wire f_arrdiv32_fs645_not0;
  wire f_arrdiv32_fs645_and0;
  wire f_arrdiv32_fs645_xor1;
  wire f_arrdiv32_fs645_not1;
  wire f_arrdiv32_fs645_and1;
  wire f_arrdiv32_fs645_or0;
  wire f_arrdiv32_fs646_xor0;
  wire f_arrdiv32_fs646_not0;
  wire f_arrdiv32_fs646_and0;
  wire f_arrdiv32_fs646_xor1;
  wire f_arrdiv32_fs646_not1;
  wire f_arrdiv32_fs646_and1;
  wire f_arrdiv32_fs646_or0;
  wire f_arrdiv32_fs647_xor0;
  wire f_arrdiv32_fs647_not0;
  wire f_arrdiv32_fs647_and0;
  wire f_arrdiv32_fs647_xor1;
  wire f_arrdiv32_fs647_not1;
  wire f_arrdiv32_fs647_and1;
  wire f_arrdiv32_fs647_or0;
  wire f_arrdiv32_fs648_xor0;
  wire f_arrdiv32_fs648_not0;
  wire f_arrdiv32_fs648_and0;
  wire f_arrdiv32_fs648_xor1;
  wire f_arrdiv32_fs648_not1;
  wire f_arrdiv32_fs648_and1;
  wire f_arrdiv32_fs648_or0;
  wire f_arrdiv32_fs649_xor0;
  wire f_arrdiv32_fs649_not0;
  wire f_arrdiv32_fs649_and0;
  wire f_arrdiv32_fs649_xor1;
  wire f_arrdiv32_fs649_not1;
  wire f_arrdiv32_fs649_and1;
  wire f_arrdiv32_fs649_or0;
  wire f_arrdiv32_fs650_xor0;
  wire f_arrdiv32_fs650_not0;
  wire f_arrdiv32_fs650_and0;
  wire f_arrdiv32_fs650_xor1;
  wire f_arrdiv32_fs650_not1;
  wire f_arrdiv32_fs650_and1;
  wire f_arrdiv32_fs650_or0;
  wire f_arrdiv32_fs651_xor0;
  wire f_arrdiv32_fs651_not0;
  wire f_arrdiv32_fs651_and0;
  wire f_arrdiv32_fs651_xor1;
  wire f_arrdiv32_fs651_not1;
  wire f_arrdiv32_fs651_and1;
  wire f_arrdiv32_fs651_or0;
  wire f_arrdiv32_fs652_xor0;
  wire f_arrdiv32_fs652_not0;
  wire f_arrdiv32_fs652_and0;
  wire f_arrdiv32_fs652_xor1;
  wire f_arrdiv32_fs652_not1;
  wire f_arrdiv32_fs652_and1;
  wire f_arrdiv32_fs652_or0;
  wire f_arrdiv32_fs653_xor0;
  wire f_arrdiv32_fs653_not0;
  wire f_arrdiv32_fs653_and0;
  wire f_arrdiv32_fs653_xor1;
  wire f_arrdiv32_fs653_not1;
  wire f_arrdiv32_fs653_and1;
  wire f_arrdiv32_fs653_or0;
  wire f_arrdiv32_fs654_xor0;
  wire f_arrdiv32_fs654_not0;
  wire f_arrdiv32_fs654_and0;
  wire f_arrdiv32_fs654_xor1;
  wire f_arrdiv32_fs654_not1;
  wire f_arrdiv32_fs654_and1;
  wire f_arrdiv32_fs654_or0;
  wire f_arrdiv32_fs655_xor0;
  wire f_arrdiv32_fs655_not0;
  wire f_arrdiv32_fs655_and0;
  wire f_arrdiv32_fs655_xor1;
  wire f_arrdiv32_fs655_not1;
  wire f_arrdiv32_fs655_and1;
  wire f_arrdiv32_fs655_or0;
  wire f_arrdiv32_fs656_xor0;
  wire f_arrdiv32_fs656_not0;
  wire f_arrdiv32_fs656_and0;
  wire f_arrdiv32_fs656_xor1;
  wire f_arrdiv32_fs656_not1;
  wire f_arrdiv32_fs656_and1;
  wire f_arrdiv32_fs656_or0;
  wire f_arrdiv32_fs657_xor0;
  wire f_arrdiv32_fs657_not0;
  wire f_arrdiv32_fs657_and0;
  wire f_arrdiv32_fs657_xor1;
  wire f_arrdiv32_fs657_not1;
  wire f_arrdiv32_fs657_and1;
  wire f_arrdiv32_fs657_or0;
  wire f_arrdiv32_fs658_xor0;
  wire f_arrdiv32_fs658_not0;
  wire f_arrdiv32_fs658_and0;
  wire f_arrdiv32_fs658_xor1;
  wire f_arrdiv32_fs658_not1;
  wire f_arrdiv32_fs658_and1;
  wire f_arrdiv32_fs658_or0;
  wire f_arrdiv32_fs659_xor0;
  wire f_arrdiv32_fs659_not0;
  wire f_arrdiv32_fs659_and0;
  wire f_arrdiv32_fs659_xor1;
  wire f_arrdiv32_fs659_not1;
  wire f_arrdiv32_fs659_and1;
  wire f_arrdiv32_fs659_or0;
  wire f_arrdiv32_fs660_xor0;
  wire f_arrdiv32_fs660_not0;
  wire f_arrdiv32_fs660_and0;
  wire f_arrdiv32_fs660_xor1;
  wire f_arrdiv32_fs660_not1;
  wire f_arrdiv32_fs660_and1;
  wire f_arrdiv32_fs660_or0;
  wire f_arrdiv32_fs661_xor0;
  wire f_arrdiv32_fs661_not0;
  wire f_arrdiv32_fs661_and0;
  wire f_arrdiv32_fs661_xor1;
  wire f_arrdiv32_fs661_not1;
  wire f_arrdiv32_fs661_and1;
  wire f_arrdiv32_fs661_or0;
  wire f_arrdiv32_fs662_xor0;
  wire f_arrdiv32_fs662_not0;
  wire f_arrdiv32_fs662_and0;
  wire f_arrdiv32_fs662_xor1;
  wire f_arrdiv32_fs662_not1;
  wire f_arrdiv32_fs662_and1;
  wire f_arrdiv32_fs662_or0;
  wire f_arrdiv32_fs663_xor0;
  wire f_arrdiv32_fs663_not0;
  wire f_arrdiv32_fs663_and0;
  wire f_arrdiv32_fs663_xor1;
  wire f_arrdiv32_fs663_not1;
  wire f_arrdiv32_fs663_and1;
  wire f_arrdiv32_fs663_or0;
  wire f_arrdiv32_fs664_xor0;
  wire f_arrdiv32_fs664_not0;
  wire f_arrdiv32_fs664_and0;
  wire f_arrdiv32_fs664_xor1;
  wire f_arrdiv32_fs664_not1;
  wire f_arrdiv32_fs664_and1;
  wire f_arrdiv32_fs664_or0;
  wire f_arrdiv32_fs665_xor0;
  wire f_arrdiv32_fs665_not0;
  wire f_arrdiv32_fs665_and0;
  wire f_arrdiv32_fs665_xor1;
  wire f_arrdiv32_fs665_not1;
  wire f_arrdiv32_fs665_and1;
  wire f_arrdiv32_fs665_or0;
  wire f_arrdiv32_fs666_xor0;
  wire f_arrdiv32_fs666_not0;
  wire f_arrdiv32_fs666_and0;
  wire f_arrdiv32_fs666_xor1;
  wire f_arrdiv32_fs666_not1;
  wire f_arrdiv32_fs666_and1;
  wire f_arrdiv32_fs666_or0;
  wire f_arrdiv32_fs667_xor0;
  wire f_arrdiv32_fs667_not0;
  wire f_arrdiv32_fs667_and0;
  wire f_arrdiv32_fs667_xor1;
  wire f_arrdiv32_fs667_not1;
  wire f_arrdiv32_fs667_and1;
  wire f_arrdiv32_fs667_or0;
  wire f_arrdiv32_fs668_xor0;
  wire f_arrdiv32_fs668_not0;
  wire f_arrdiv32_fs668_and0;
  wire f_arrdiv32_fs668_xor1;
  wire f_arrdiv32_fs668_not1;
  wire f_arrdiv32_fs668_and1;
  wire f_arrdiv32_fs668_or0;
  wire f_arrdiv32_fs669_xor0;
  wire f_arrdiv32_fs669_not0;
  wire f_arrdiv32_fs669_and0;
  wire f_arrdiv32_fs669_xor1;
  wire f_arrdiv32_fs669_not1;
  wire f_arrdiv32_fs669_and1;
  wire f_arrdiv32_fs669_or0;
  wire f_arrdiv32_fs670_xor0;
  wire f_arrdiv32_fs670_not0;
  wire f_arrdiv32_fs670_and0;
  wire f_arrdiv32_fs670_xor1;
  wire f_arrdiv32_fs670_not1;
  wire f_arrdiv32_fs670_and1;
  wire f_arrdiv32_fs670_or0;
  wire f_arrdiv32_fs671_xor0;
  wire f_arrdiv32_fs671_not0;
  wire f_arrdiv32_fs671_and0;
  wire f_arrdiv32_fs671_xor1;
  wire f_arrdiv32_fs671_not1;
  wire f_arrdiv32_fs671_and1;
  wire f_arrdiv32_fs671_or0;
  wire f_arrdiv32_mux2to1620_and0;
  wire f_arrdiv32_mux2to1620_not0;
  wire f_arrdiv32_mux2to1620_and1;
  wire f_arrdiv32_mux2to1620_xor0;
  wire f_arrdiv32_mux2to1621_and0;
  wire f_arrdiv32_mux2to1621_not0;
  wire f_arrdiv32_mux2to1621_and1;
  wire f_arrdiv32_mux2to1621_xor0;
  wire f_arrdiv32_mux2to1622_and0;
  wire f_arrdiv32_mux2to1622_not0;
  wire f_arrdiv32_mux2to1622_and1;
  wire f_arrdiv32_mux2to1622_xor0;
  wire f_arrdiv32_mux2to1623_and0;
  wire f_arrdiv32_mux2to1623_not0;
  wire f_arrdiv32_mux2to1623_and1;
  wire f_arrdiv32_mux2to1623_xor0;
  wire f_arrdiv32_mux2to1624_and0;
  wire f_arrdiv32_mux2to1624_not0;
  wire f_arrdiv32_mux2to1624_and1;
  wire f_arrdiv32_mux2to1624_xor0;
  wire f_arrdiv32_mux2to1625_and0;
  wire f_arrdiv32_mux2to1625_not0;
  wire f_arrdiv32_mux2to1625_and1;
  wire f_arrdiv32_mux2to1625_xor0;
  wire f_arrdiv32_mux2to1626_and0;
  wire f_arrdiv32_mux2to1626_not0;
  wire f_arrdiv32_mux2to1626_and1;
  wire f_arrdiv32_mux2to1626_xor0;
  wire f_arrdiv32_mux2to1627_and0;
  wire f_arrdiv32_mux2to1627_not0;
  wire f_arrdiv32_mux2to1627_and1;
  wire f_arrdiv32_mux2to1627_xor0;
  wire f_arrdiv32_mux2to1628_and0;
  wire f_arrdiv32_mux2to1628_not0;
  wire f_arrdiv32_mux2to1628_and1;
  wire f_arrdiv32_mux2to1628_xor0;
  wire f_arrdiv32_mux2to1629_and0;
  wire f_arrdiv32_mux2to1629_not0;
  wire f_arrdiv32_mux2to1629_and1;
  wire f_arrdiv32_mux2to1629_xor0;
  wire f_arrdiv32_mux2to1630_and0;
  wire f_arrdiv32_mux2to1630_not0;
  wire f_arrdiv32_mux2to1630_and1;
  wire f_arrdiv32_mux2to1630_xor0;
  wire f_arrdiv32_mux2to1631_and0;
  wire f_arrdiv32_mux2to1631_not0;
  wire f_arrdiv32_mux2to1631_and1;
  wire f_arrdiv32_mux2to1631_xor0;
  wire f_arrdiv32_mux2to1632_and0;
  wire f_arrdiv32_mux2to1632_not0;
  wire f_arrdiv32_mux2to1632_and1;
  wire f_arrdiv32_mux2to1632_xor0;
  wire f_arrdiv32_mux2to1633_and0;
  wire f_arrdiv32_mux2to1633_not0;
  wire f_arrdiv32_mux2to1633_and1;
  wire f_arrdiv32_mux2to1633_xor0;
  wire f_arrdiv32_mux2to1634_and0;
  wire f_arrdiv32_mux2to1634_not0;
  wire f_arrdiv32_mux2to1634_and1;
  wire f_arrdiv32_mux2to1634_xor0;
  wire f_arrdiv32_mux2to1635_and0;
  wire f_arrdiv32_mux2to1635_not0;
  wire f_arrdiv32_mux2to1635_and1;
  wire f_arrdiv32_mux2to1635_xor0;
  wire f_arrdiv32_mux2to1636_and0;
  wire f_arrdiv32_mux2to1636_not0;
  wire f_arrdiv32_mux2to1636_and1;
  wire f_arrdiv32_mux2to1636_xor0;
  wire f_arrdiv32_mux2to1637_and0;
  wire f_arrdiv32_mux2to1637_not0;
  wire f_arrdiv32_mux2to1637_and1;
  wire f_arrdiv32_mux2to1637_xor0;
  wire f_arrdiv32_mux2to1638_and0;
  wire f_arrdiv32_mux2to1638_not0;
  wire f_arrdiv32_mux2to1638_and1;
  wire f_arrdiv32_mux2to1638_xor0;
  wire f_arrdiv32_mux2to1639_and0;
  wire f_arrdiv32_mux2to1639_not0;
  wire f_arrdiv32_mux2to1639_and1;
  wire f_arrdiv32_mux2to1639_xor0;
  wire f_arrdiv32_mux2to1640_and0;
  wire f_arrdiv32_mux2to1640_not0;
  wire f_arrdiv32_mux2to1640_and1;
  wire f_arrdiv32_mux2to1640_xor0;
  wire f_arrdiv32_mux2to1641_and0;
  wire f_arrdiv32_mux2to1641_not0;
  wire f_arrdiv32_mux2to1641_and1;
  wire f_arrdiv32_mux2to1641_xor0;
  wire f_arrdiv32_mux2to1642_and0;
  wire f_arrdiv32_mux2to1642_not0;
  wire f_arrdiv32_mux2to1642_and1;
  wire f_arrdiv32_mux2to1642_xor0;
  wire f_arrdiv32_mux2to1643_and0;
  wire f_arrdiv32_mux2to1643_not0;
  wire f_arrdiv32_mux2to1643_and1;
  wire f_arrdiv32_mux2to1643_xor0;
  wire f_arrdiv32_mux2to1644_and0;
  wire f_arrdiv32_mux2to1644_not0;
  wire f_arrdiv32_mux2to1644_and1;
  wire f_arrdiv32_mux2to1644_xor0;
  wire f_arrdiv32_mux2to1645_and0;
  wire f_arrdiv32_mux2to1645_not0;
  wire f_arrdiv32_mux2to1645_and1;
  wire f_arrdiv32_mux2to1645_xor0;
  wire f_arrdiv32_mux2to1646_and0;
  wire f_arrdiv32_mux2to1646_not0;
  wire f_arrdiv32_mux2to1646_and1;
  wire f_arrdiv32_mux2to1646_xor0;
  wire f_arrdiv32_mux2to1647_and0;
  wire f_arrdiv32_mux2to1647_not0;
  wire f_arrdiv32_mux2to1647_and1;
  wire f_arrdiv32_mux2to1647_xor0;
  wire f_arrdiv32_mux2to1648_and0;
  wire f_arrdiv32_mux2to1648_not0;
  wire f_arrdiv32_mux2to1648_and1;
  wire f_arrdiv32_mux2to1648_xor0;
  wire f_arrdiv32_mux2to1649_and0;
  wire f_arrdiv32_mux2to1649_not0;
  wire f_arrdiv32_mux2to1649_and1;
  wire f_arrdiv32_mux2to1649_xor0;
  wire f_arrdiv32_mux2to1650_and0;
  wire f_arrdiv32_mux2to1650_not0;
  wire f_arrdiv32_mux2to1650_and1;
  wire f_arrdiv32_mux2to1650_xor0;
  wire f_arrdiv32_not20;
  wire f_arrdiv32_fs672_xor0;
  wire f_arrdiv32_fs672_not0;
  wire f_arrdiv32_fs672_and0;
  wire f_arrdiv32_fs672_not1;
  wire f_arrdiv32_fs673_xor0;
  wire f_arrdiv32_fs673_not0;
  wire f_arrdiv32_fs673_and0;
  wire f_arrdiv32_fs673_xor1;
  wire f_arrdiv32_fs673_not1;
  wire f_arrdiv32_fs673_and1;
  wire f_arrdiv32_fs673_or0;
  wire f_arrdiv32_fs674_xor0;
  wire f_arrdiv32_fs674_not0;
  wire f_arrdiv32_fs674_and0;
  wire f_arrdiv32_fs674_xor1;
  wire f_arrdiv32_fs674_not1;
  wire f_arrdiv32_fs674_and1;
  wire f_arrdiv32_fs674_or0;
  wire f_arrdiv32_fs675_xor0;
  wire f_arrdiv32_fs675_not0;
  wire f_arrdiv32_fs675_and0;
  wire f_arrdiv32_fs675_xor1;
  wire f_arrdiv32_fs675_not1;
  wire f_arrdiv32_fs675_and1;
  wire f_arrdiv32_fs675_or0;
  wire f_arrdiv32_fs676_xor0;
  wire f_arrdiv32_fs676_not0;
  wire f_arrdiv32_fs676_and0;
  wire f_arrdiv32_fs676_xor1;
  wire f_arrdiv32_fs676_not1;
  wire f_arrdiv32_fs676_and1;
  wire f_arrdiv32_fs676_or0;
  wire f_arrdiv32_fs677_xor0;
  wire f_arrdiv32_fs677_not0;
  wire f_arrdiv32_fs677_and0;
  wire f_arrdiv32_fs677_xor1;
  wire f_arrdiv32_fs677_not1;
  wire f_arrdiv32_fs677_and1;
  wire f_arrdiv32_fs677_or0;
  wire f_arrdiv32_fs678_xor0;
  wire f_arrdiv32_fs678_not0;
  wire f_arrdiv32_fs678_and0;
  wire f_arrdiv32_fs678_xor1;
  wire f_arrdiv32_fs678_not1;
  wire f_arrdiv32_fs678_and1;
  wire f_arrdiv32_fs678_or0;
  wire f_arrdiv32_fs679_xor0;
  wire f_arrdiv32_fs679_not0;
  wire f_arrdiv32_fs679_and0;
  wire f_arrdiv32_fs679_xor1;
  wire f_arrdiv32_fs679_not1;
  wire f_arrdiv32_fs679_and1;
  wire f_arrdiv32_fs679_or0;
  wire f_arrdiv32_fs680_xor0;
  wire f_arrdiv32_fs680_not0;
  wire f_arrdiv32_fs680_and0;
  wire f_arrdiv32_fs680_xor1;
  wire f_arrdiv32_fs680_not1;
  wire f_arrdiv32_fs680_and1;
  wire f_arrdiv32_fs680_or0;
  wire f_arrdiv32_fs681_xor0;
  wire f_arrdiv32_fs681_not0;
  wire f_arrdiv32_fs681_and0;
  wire f_arrdiv32_fs681_xor1;
  wire f_arrdiv32_fs681_not1;
  wire f_arrdiv32_fs681_and1;
  wire f_arrdiv32_fs681_or0;
  wire f_arrdiv32_fs682_xor0;
  wire f_arrdiv32_fs682_not0;
  wire f_arrdiv32_fs682_and0;
  wire f_arrdiv32_fs682_xor1;
  wire f_arrdiv32_fs682_not1;
  wire f_arrdiv32_fs682_and1;
  wire f_arrdiv32_fs682_or0;
  wire f_arrdiv32_fs683_xor0;
  wire f_arrdiv32_fs683_not0;
  wire f_arrdiv32_fs683_and0;
  wire f_arrdiv32_fs683_xor1;
  wire f_arrdiv32_fs683_not1;
  wire f_arrdiv32_fs683_and1;
  wire f_arrdiv32_fs683_or0;
  wire f_arrdiv32_fs684_xor0;
  wire f_arrdiv32_fs684_not0;
  wire f_arrdiv32_fs684_and0;
  wire f_arrdiv32_fs684_xor1;
  wire f_arrdiv32_fs684_not1;
  wire f_arrdiv32_fs684_and1;
  wire f_arrdiv32_fs684_or0;
  wire f_arrdiv32_fs685_xor0;
  wire f_arrdiv32_fs685_not0;
  wire f_arrdiv32_fs685_and0;
  wire f_arrdiv32_fs685_xor1;
  wire f_arrdiv32_fs685_not1;
  wire f_arrdiv32_fs685_and1;
  wire f_arrdiv32_fs685_or0;
  wire f_arrdiv32_fs686_xor0;
  wire f_arrdiv32_fs686_not0;
  wire f_arrdiv32_fs686_and0;
  wire f_arrdiv32_fs686_xor1;
  wire f_arrdiv32_fs686_not1;
  wire f_arrdiv32_fs686_and1;
  wire f_arrdiv32_fs686_or0;
  wire f_arrdiv32_fs687_xor0;
  wire f_arrdiv32_fs687_not0;
  wire f_arrdiv32_fs687_and0;
  wire f_arrdiv32_fs687_xor1;
  wire f_arrdiv32_fs687_not1;
  wire f_arrdiv32_fs687_and1;
  wire f_arrdiv32_fs687_or0;
  wire f_arrdiv32_fs688_xor0;
  wire f_arrdiv32_fs688_not0;
  wire f_arrdiv32_fs688_and0;
  wire f_arrdiv32_fs688_xor1;
  wire f_arrdiv32_fs688_not1;
  wire f_arrdiv32_fs688_and1;
  wire f_arrdiv32_fs688_or0;
  wire f_arrdiv32_fs689_xor0;
  wire f_arrdiv32_fs689_not0;
  wire f_arrdiv32_fs689_and0;
  wire f_arrdiv32_fs689_xor1;
  wire f_arrdiv32_fs689_not1;
  wire f_arrdiv32_fs689_and1;
  wire f_arrdiv32_fs689_or0;
  wire f_arrdiv32_fs690_xor0;
  wire f_arrdiv32_fs690_not0;
  wire f_arrdiv32_fs690_and0;
  wire f_arrdiv32_fs690_xor1;
  wire f_arrdiv32_fs690_not1;
  wire f_arrdiv32_fs690_and1;
  wire f_arrdiv32_fs690_or0;
  wire f_arrdiv32_fs691_xor0;
  wire f_arrdiv32_fs691_not0;
  wire f_arrdiv32_fs691_and0;
  wire f_arrdiv32_fs691_xor1;
  wire f_arrdiv32_fs691_not1;
  wire f_arrdiv32_fs691_and1;
  wire f_arrdiv32_fs691_or0;
  wire f_arrdiv32_fs692_xor0;
  wire f_arrdiv32_fs692_not0;
  wire f_arrdiv32_fs692_and0;
  wire f_arrdiv32_fs692_xor1;
  wire f_arrdiv32_fs692_not1;
  wire f_arrdiv32_fs692_and1;
  wire f_arrdiv32_fs692_or0;
  wire f_arrdiv32_fs693_xor0;
  wire f_arrdiv32_fs693_not0;
  wire f_arrdiv32_fs693_and0;
  wire f_arrdiv32_fs693_xor1;
  wire f_arrdiv32_fs693_not1;
  wire f_arrdiv32_fs693_and1;
  wire f_arrdiv32_fs693_or0;
  wire f_arrdiv32_fs694_xor0;
  wire f_arrdiv32_fs694_not0;
  wire f_arrdiv32_fs694_and0;
  wire f_arrdiv32_fs694_xor1;
  wire f_arrdiv32_fs694_not1;
  wire f_arrdiv32_fs694_and1;
  wire f_arrdiv32_fs694_or0;
  wire f_arrdiv32_fs695_xor0;
  wire f_arrdiv32_fs695_not0;
  wire f_arrdiv32_fs695_and0;
  wire f_arrdiv32_fs695_xor1;
  wire f_arrdiv32_fs695_not1;
  wire f_arrdiv32_fs695_and1;
  wire f_arrdiv32_fs695_or0;
  wire f_arrdiv32_fs696_xor0;
  wire f_arrdiv32_fs696_not0;
  wire f_arrdiv32_fs696_and0;
  wire f_arrdiv32_fs696_xor1;
  wire f_arrdiv32_fs696_not1;
  wire f_arrdiv32_fs696_and1;
  wire f_arrdiv32_fs696_or0;
  wire f_arrdiv32_fs697_xor0;
  wire f_arrdiv32_fs697_not0;
  wire f_arrdiv32_fs697_and0;
  wire f_arrdiv32_fs697_xor1;
  wire f_arrdiv32_fs697_not1;
  wire f_arrdiv32_fs697_and1;
  wire f_arrdiv32_fs697_or0;
  wire f_arrdiv32_fs698_xor0;
  wire f_arrdiv32_fs698_not0;
  wire f_arrdiv32_fs698_and0;
  wire f_arrdiv32_fs698_xor1;
  wire f_arrdiv32_fs698_not1;
  wire f_arrdiv32_fs698_and1;
  wire f_arrdiv32_fs698_or0;
  wire f_arrdiv32_fs699_xor0;
  wire f_arrdiv32_fs699_not0;
  wire f_arrdiv32_fs699_and0;
  wire f_arrdiv32_fs699_xor1;
  wire f_arrdiv32_fs699_not1;
  wire f_arrdiv32_fs699_and1;
  wire f_arrdiv32_fs699_or0;
  wire f_arrdiv32_fs700_xor0;
  wire f_arrdiv32_fs700_not0;
  wire f_arrdiv32_fs700_and0;
  wire f_arrdiv32_fs700_xor1;
  wire f_arrdiv32_fs700_not1;
  wire f_arrdiv32_fs700_and1;
  wire f_arrdiv32_fs700_or0;
  wire f_arrdiv32_fs701_xor0;
  wire f_arrdiv32_fs701_not0;
  wire f_arrdiv32_fs701_and0;
  wire f_arrdiv32_fs701_xor1;
  wire f_arrdiv32_fs701_not1;
  wire f_arrdiv32_fs701_and1;
  wire f_arrdiv32_fs701_or0;
  wire f_arrdiv32_fs702_xor0;
  wire f_arrdiv32_fs702_not0;
  wire f_arrdiv32_fs702_and0;
  wire f_arrdiv32_fs702_xor1;
  wire f_arrdiv32_fs702_not1;
  wire f_arrdiv32_fs702_and1;
  wire f_arrdiv32_fs702_or0;
  wire f_arrdiv32_fs703_xor0;
  wire f_arrdiv32_fs703_not0;
  wire f_arrdiv32_fs703_and0;
  wire f_arrdiv32_fs703_xor1;
  wire f_arrdiv32_fs703_not1;
  wire f_arrdiv32_fs703_and1;
  wire f_arrdiv32_fs703_or0;
  wire f_arrdiv32_mux2to1651_and0;
  wire f_arrdiv32_mux2to1651_not0;
  wire f_arrdiv32_mux2to1651_and1;
  wire f_arrdiv32_mux2to1651_xor0;
  wire f_arrdiv32_mux2to1652_and0;
  wire f_arrdiv32_mux2to1652_not0;
  wire f_arrdiv32_mux2to1652_and1;
  wire f_arrdiv32_mux2to1652_xor0;
  wire f_arrdiv32_mux2to1653_and0;
  wire f_arrdiv32_mux2to1653_not0;
  wire f_arrdiv32_mux2to1653_and1;
  wire f_arrdiv32_mux2to1653_xor0;
  wire f_arrdiv32_mux2to1654_and0;
  wire f_arrdiv32_mux2to1654_not0;
  wire f_arrdiv32_mux2to1654_and1;
  wire f_arrdiv32_mux2to1654_xor0;
  wire f_arrdiv32_mux2to1655_and0;
  wire f_arrdiv32_mux2to1655_not0;
  wire f_arrdiv32_mux2to1655_and1;
  wire f_arrdiv32_mux2to1655_xor0;
  wire f_arrdiv32_mux2to1656_and0;
  wire f_arrdiv32_mux2to1656_not0;
  wire f_arrdiv32_mux2to1656_and1;
  wire f_arrdiv32_mux2to1656_xor0;
  wire f_arrdiv32_mux2to1657_and0;
  wire f_arrdiv32_mux2to1657_not0;
  wire f_arrdiv32_mux2to1657_and1;
  wire f_arrdiv32_mux2to1657_xor0;
  wire f_arrdiv32_mux2to1658_and0;
  wire f_arrdiv32_mux2to1658_not0;
  wire f_arrdiv32_mux2to1658_and1;
  wire f_arrdiv32_mux2to1658_xor0;
  wire f_arrdiv32_mux2to1659_and0;
  wire f_arrdiv32_mux2to1659_not0;
  wire f_arrdiv32_mux2to1659_and1;
  wire f_arrdiv32_mux2to1659_xor0;
  wire f_arrdiv32_mux2to1660_and0;
  wire f_arrdiv32_mux2to1660_not0;
  wire f_arrdiv32_mux2to1660_and1;
  wire f_arrdiv32_mux2to1660_xor0;
  wire f_arrdiv32_mux2to1661_and0;
  wire f_arrdiv32_mux2to1661_not0;
  wire f_arrdiv32_mux2to1661_and1;
  wire f_arrdiv32_mux2to1661_xor0;
  wire f_arrdiv32_mux2to1662_and0;
  wire f_arrdiv32_mux2to1662_not0;
  wire f_arrdiv32_mux2to1662_and1;
  wire f_arrdiv32_mux2to1662_xor0;
  wire f_arrdiv32_mux2to1663_and0;
  wire f_arrdiv32_mux2to1663_not0;
  wire f_arrdiv32_mux2to1663_and1;
  wire f_arrdiv32_mux2to1663_xor0;
  wire f_arrdiv32_mux2to1664_and0;
  wire f_arrdiv32_mux2to1664_not0;
  wire f_arrdiv32_mux2to1664_and1;
  wire f_arrdiv32_mux2to1664_xor0;
  wire f_arrdiv32_mux2to1665_and0;
  wire f_arrdiv32_mux2to1665_not0;
  wire f_arrdiv32_mux2to1665_and1;
  wire f_arrdiv32_mux2to1665_xor0;
  wire f_arrdiv32_mux2to1666_and0;
  wire f_arrdiv32_mux2to1666_not0;
  wire f_arrdiv32_mux2to1666_and1;
  wire f_arrdiv32_mux2to1666_xor0;
  wire f_arrdiv32_mux2to1667_and0;
  wire f_arrdiv32_mux2to1667_not0;
  wire f_arrdiv32_mux2to1667_and1;
  wire f_arrdiv32_mux2to1667_xor0;
  wire f_arrdiv32_mux2to1668_and0;
  wire f_arrdiv32_mux2to1668_not0;
  wire f_arrdiv32_mux2to1668_and1;
  wire f_arrdiv32_mux2to1668_xor0;
  wire f_arrdiv32_mux2to1669_and0;
  wire f_arrdiv32_mux2to1669_not0;
  wire f_arrdiv32_mux2to1669_and1;
  wire f_arrdiv32_mux2to1669_xor0;
  wire f_arrdiv32_mux2to1670_and0;
  wire f_arrdiv32_mux2to1670_not0;
  wire f_arrdiv32_mux2to1670_and1;
  wire f_arrdiv32_mux2to1670_xor0;
  wire f_arrdiv32_mux2to1671_and0;
  wire f_arrdiv32_mux2to1671_not0;
  wire f_arrdiv32_mux2to1671_and1;
  wire f_arrdiv32_mux2to1671_xor0;
  wire f_arrdiv32_mux2to1672_and0;
  wire f_arrdiv32_mux2to1672_not0;
  wire f_arrdiv32_mux2to1672_and1;
  wire f_arrdiv32_mux2to1672_xor0;
  wire f_arrdiv32_mux2to1673_and0;
  wire f_arrdiv32_mux2to1673_not0;
  wire f_arrdiv32_mux2to1673_and1;
  wire f_arrdiv32_mux2to1673_xor0;
  wire f_arrdiv32_mux2to1674_and0;
  wire f_arrdiv32_mux2to1674_not0;
  wire f_arrdiv32_mux2to1674_and1;
  wire f_arrdiv32_mux2to1674_xor0;
  wire f_arrdiv32_mux2to1675_and0;
  wire f_arrdiv32_mux2to1675_not0;
  wire f_arrdiv32_mux2to1675_and1;
  wire f_arrdiv32_mux2to1675_xor0;
  wire f_arrdiv32_mux2to1676_and0;
  wire f_arrdiv32_mux2to1676_not0;
  wire f_arrdiv32_mux2to1676_and1;
  wire f_arrdiv32_mux2to1676_xor0;
  wire f_arrdiv32_mux2to1677_and0;
  wire f_arrdiv32_mux2to1677_not0;
  wire f_arrdiv32_mux2to1677_and1;
  wire f_arrdiv32_mux2to1677_xor0;
  wire f_arrdiv32_mux2to1678_and0;
  wire f_arrdiv32_mux2to1678_not0;
  wire f_arrdiv32_mux2to1678_and1;
  wire f_arrdiv32_mux2to1678_xor0;
  wire f_arrdiv32_mux2to1679_and0;
  wire f_arrdiv32_mux2to1679_not0;
  wire f_arrdiv32_mux2to1679_and1;
  wire f_arrdiv32_mux2to1679_xor0;
  wire f_arrdiv32_mux2to1680_and0;
  wire f_arrdiv32_mux2to1680_not0;
  wire f_arrdiv32_mux2to1680_and1;
  wire f_arrdiv32_mux2to1680_xor0;
  wire f_arrdiv32_mux2to1681_and0;
  wire f_arrdiv32_mux2to1681_not0;
  wire f_arrdiv32_mux2to1681_and1;
  wire f_arrdiv32_mux2to1681_xor0;
  wire f_arrdiv32_not21;
  wire f_arrdiv32_fs704_xor0;
  wire f_arrdiv32_fs704_not0;
  wire f_arrdiv32_fs704_and0;
  wire f_arrdiv32_fs704_not1;
  wire f_arrdiv32_fs705_xor0;
  wire f_arrdiv32_fs705_not0;
  wire f_arrdiv32_fs705_and0;
  wire f_arrdiv32_fs705_xor1;
  wire f_arrdiv32_fs705_not1;
  wire f_arrdiv32_fs705_and1;
  wire f_arrdiv32_fs705_or0;
  wire f_arrdiv32_fs706_xor0;
  wire f_arrdiv32_fs706_not0;
  wire f_arrdiv32_fs706_and0;
  wire f_arrdiv32_fs706_xor1;
  wire f_arrdiv32_fs706_not1;
  wire f_arrdiv32_fs706_and1;
  wire f_arrdiv32_fs706_or0;
  wire f_arrdiv32_fs707_xor0;
  wire f_arrdiv32_fs707_not0;
  wire f_arrdiv32_fs707_and0;
  wire f_arrdiv32_fs707_xor1;
  wire f_arrdiv32_fs707_not1;
  wire f_arrdiv32_fs707_and1;
  wire f_arrdiv32_fs707_or0;
  wire f_arrdiv32_fs708_xor0;
  wire f_arrdiv32_fs708_not0;
  wire f_arrdiv32_fs708_and0;
  wire f_arrdiv32_fs708_xor1;
  wire f_arrdiv32_fs708_not1;
  wire f_arrdiv32_fs708_and1;
  wire f_arrdiv32_fs708_or0;
  wire f_arrdiv32_fs709_xor0;
  wire f_arrdiv32_fs709_not0;
  wire f_arrdiv32_fs709_and0;
  wire f_arrdiv32_fs709_xor1;
  wire f_arrdiv32_fs709_not1;
  wire f_arrdiv32_fs709_and1;
  wire f_arrdiv32_fs709_or0;
  wire f_arrdiv32_fs710_xor0;
  wire f_arrdiv32_fs710_not0;
  wire f_arrdiv32_fs710_and0;
  wire f_arrdiv32_fs710_xor1;
  wire f_arrdiv32_fs710_not1;
  wire f_arrdiv32_fs710_and1;
  wire f_arrdiv32_fs710_or0;
  wire f_arrdiv32_fs711_xor0;
  wire f_arrdiv32_fs711_not0;
  wire f_arrdiv32_fs711_and0;
  wire f_arrdiv32_fs711_xor1;
  wire f_arrdiv32_fs711_not1;
  wire f_arrdiv32_fs711_and1;
  wire f_arrdiv32_fs711_or0;
  wire f_arrdiv32_fs712_xor0;
  wire f_arrdiv32_fs712_not0;
  wire f_arrdiv32_fs712_and0;
  wire f_arrdiv32_fs712_xor1;
  wire f_arrdiv32_fs712_not1;
  wire f_arrdiv32_fs712_and1;
  wire f_arrdiv32_fs712_or0;
  wire f_arrdiv32_fs713_xor0;
  wire f_arrdiv32_fs713_not0;
  wire f_arrdiv32_fs713_and0;
  wire f_arrdiv32_fs713_xor1;
  wire f_arrdiv32_fs713_not1;
  wire f_arrdiv32_fs713_and1;
  wire f_arrdiv32_fs713_or0;
  wire f_arrdiv32_fs714_xor0;
  wire f_arrdiv32_fs714_not0;
  wire f_arrdiv32_fs714_and0;
  wire f_arrdiv32_fs714_xor1;
  wire f_arrdiv32_fs714_not1;
  wire f_arrdiv32_fs714_and1;
  wire f_arrdiv32_fs714_or0;
  wire f_arrdiv32_fs715_xor0;
  wire f_arrdiv32_fs715_not0;
  wire f_arrdiv32_fs715_and0;
  wire f_arrdiv32_fs715_xor1;
  wire f_arrdiv32_fs715_not1;
  wire f_arrdiv32_fs715_and1;
  wire f_arrdiv32_fs715_or0;
  wire f_arrdiv32_fs716_xor0;
  wire f_arrdiv32_fs716_not0;
  wire f_arrdiv32_fs716_and0;
  wire f_arrdiv32_fs716_xor1;
  wire f_arrdiv32_fs716_not1;
  wire f_arrdiv32_fs716_and1;
  wire f_arrdiv32_fs716_or0;
  wire f_arrdiv32_fs717_xor0;
  wire f_arrdiv32_fs717_not0;
  wire f_arrdiv32_fs717_and0;
  wire f_arrdiv32_fs717_xor1;
  wire f_arrdiv32_fs717_not1;
  wire f_arrdiv32_fs717_and1;
  wire f_arrdiv32_fs717_or0;
  wire f_arrdiv32_fs718_xor0;
  wire f_arrdiv32_fs718_not0;
  wire f_arrdiv32_fs718_and0;
  wire f_arrdiv32_fs718_xor1;
  wire f_arrdiv32_fs718_not1;
  wire f_arrdiv32_fs718_and1;
  wire f_arrdiv32_fs718_or0;
  wire f_arrdiv32_fs719_xor0;
  wire f_arrdiv32_fs719_not0;
  wire f_arrdiv32_fs719_and0;
  wire f_arrdiv32_fs719_xor1;
  wire f_arrdiv32_fs719_not1;
  wire f_arrdiv32_fs719_and1;
  wire f_arrdiv32_fs719_or0;
  wire f_arrdiv32_fs720_xor0;
  wire f_arrdiv32_fs720_not0;
  wire f_arrdiv32_fs720_and0;
  wire f_arrdiv32_fs720_xor1;
  wire f_arrdiv32_fs720_not1;
  wire f_arrdiv32_fs720_and1;
  wire f_arrdiv32_fs720_or0;
  wire f_arrdiv32_fs721_xor0;
  wire f_arrdiv32_fs721_not0;
  wire f_arrdiv32_fs721_and0;
  wire f_arrdiv32_fs721_xor1;
  wire f_arrdiv32_fs721_not1;
  wire f_arrdiv32_fs721_and1;
  wire f_arrdiv32_fs721_or0;
  wire f_arrdiv32_fs722_xor0;
  wire f_arrdiv32_fs722_not0;
  wire f_arrdiv32_fs722_and0;
  wire f_arrdiv32_fs722_xor1;
  wire f_arrdiv32_fs722_not1;
  wire f_arrdiv32_fs722_and1;
  wire f_arrdiv32_fs722_or0;
  wire f_arrdiv32_fs723_xor0;
  wire f_arrdiv32_fs723_not0;
  wire f_arrdiv32_fs723_and0;
  wire f_arrdiv32_fs723_xor1;
  wire f_arrdiv32_fs723_not1;
  wire f_arrdiv32_fs723_and1;
  wire f_arrdiv32_fs723_or0;
  wire f_arrdiv32_fs724_xor0;
  wire f_arrdiv32_fs724_not0;
  wire f_arrdiv32_fs724_and0;
  wire f_arrdiv32_fs724_xor1;
  wire f_arrdiv32_fs724_not1;
  wire f_arrdiv32_fs724_and1;
  wire f_arrdiv32_fs724_or0;
  wire f_arrdiv32_fs725_xor0;
  wire f_arrdiv32_fs725_not0;
  wire f_arrdiv32_fs725_and0;
  wire f_arrdiv32_fs725_xor1;
  wire f_arrdiv32_fs725_not1;
  wire f_arrdiv32_fs725_and1;
  wire f_arrdiv32_fs725_or0;
  wire f_arrdiv32_fs726_xor0;
  wire f_arrdiv32_fs726_not0;
  wire f_arrdiv32_fs726_and0;
  wire f_arrdiv32_fs726_xor1;
  wire f_arrdiv32_fs726_not1;
  wire f_arrdiv32_fs726_and1;
  wire f_arrdiv32_fs726_or0;
  wire f_arrdiv32_fs727_xor0;
  wire f_arrdiv32_fs727_not0;
  wire f_arrdiv32_fs727_and0;
  wire f_arrdiv32_fs727_xor1;
  wire f_arrdiv32_fs727_not1;
  wire f_arrdiv32_fs727_and1;
  wire f_arrdiv32_fs727_or0;
  wire f_arrdiv32_fs728_xor0;
  wire f_arrdiv32_fs728_not0;
  wire f_arrdiv32_fs728_and0;
  wire f_arrdiv32_fs728_xor1;
  wire f_arrdiv32_fs728_not1;
  wire f_arrdiv32_fs728_and1;
  wire f_arrdiv32_fs728_or0;
  wire f_arrdiv32_fs729_xor0;
  wire f_arrdiv32_fs729_not0;
  wire f_arrdiv32_fs729_and0;
  wire f_arrdiv32_fs729_xor1;
  wire f_arrdiv32_fs729_not1;
  wire f_arrdiv32_fs729_and1;
  wire f_arrdiv32_fs729_or0;
  wire f_arrdiv32_fs730_xor0;
  wire f_arrdiv32_fs730_not0;
  wire f_arrdiv32_fs730_and0;
  wire f_arrdiv32_fs730_xor1;
  wire f_arrdiv32_fs730_not1;
  wire f_arrdiv32_fs730_and1;
  wire f_arrdiv32_fs730_or0;
  wire f_arrdiv32_fs731_xor0;
  wire f_arrdiv32_fs731_not0;
  wire f_arrdiv32_fs731_and0;
  wire f_arrdiv32_fs731_xor1;
  wire f_arrdiv32_fs731_not1;
  wire f_arrdiv32_fs731_and1;
  wire f_arrdiv32_fs731_or0;
  wire f_arrdiv32_fs732_xor0;
  wire f_arrdiv32_fs732_not0;
  wire f_arrdiv32_fs732_and0;
  wire f_arrdiv32_fs732_xor1;
  wire f_arrdiv32_fs732_not1;
  wire f_arrdiv32_fs732_and1;
  wire f_arrdiv32_fs732_or0;
  wire f_arrdiv32_fs733_xor0;
  wire f_arrdiv32_fs733_not0;
  wire f_arrdiv32_fs733_and0;
  wire f_arrdiv32_fs733_xor1;
  wire f_arrdiv32_fs733_not1;
  wire f_arrdiv32_fs733_and1;
  wire f_arrdiv32_fs733_or0;
  wire f_arrdiv32_fs734_xor0;
  wire f_arrdiv32_fs734_not0;
  wire f_arrdiv32_fs734_and0;
  wire f_arrdiv32_fs734_xor1;
  wire f_arrdiv32_fs734_not1;
  wire f_arrdiv32_fs734_and1;
  wire f_arrdiv32_fs734_or0;
  wire f_arrdiv32_fs735_xor0;
  wire f_arrdiv32_fs735_not0;
  wire f_arrdiv32_fs735_and0;
  wire f_arrdiv32_fs735_xor1;
  wire f_arrdiv32_fs735_not1;
  wire f_arrdiv32_fs735_and1;
  wire f_arrdiv32_fs735_or0;
  wire f_arrdiv32_mux2to1682_and0;
  wire f_arrdiv32_mux2to1682_not0;
  wire f_arrdiv32_mux2to1682_and1;
  wire f_arrdiv32_mux2to1682_xor0;
  wire f_arrdiv32_mux2to1683_and0;
  wire f_arrdiv32_mux2to1683_not0;
  wire f_arrdiv32_mux2to1683_and1;
  wire f_arrdiv32_mux2to1683_xor0;
  wire f_arrdiv32_mux2to1684_and0;
  wire f_arrdiv32_mux2to1684_not0;
  wire f_arrdiv32_mux2to1684_and1;
  wire f_arrdiv32_mux2to1684_xor0;
  wire f_arrdiv32_mux2to1685_and0;
  wire f_arrdiv32_mux2to1685_not0;
  wire f_arrdiv32_mux2to1685_and1;
  wire f_arrdiv32_mux2to1685_xor0;
  wire f_arrdiv32_mux2to1686_and0;
  wire f_arrdiv32_mux2to1686_not0;
  wire f_arrdiv32_mux2to1686_and1;
  wire f_arrdiv32_mux2to1686_xor0;
  wire f_arrdiv32_mux2to1687_and0;
  wire f_arrdiv32_mux2to1687_not0;
  wire f_arrdiv32_mux2to1687_and1;
  wire f_arrdiv32_mux2to1687_xor0;
  wire f_arrdiv32_mux2to1688_and0;
  wire f_arrdiv32_mux2to1688_not0;
  wire f_arrdiv32_mux2to1688_and1;
  wire f_arrdiv32_mux2to1688_xor0;
  wire f_arrdiv32_mux2to1689_and0;
  wire f_arrdiv32_mux2to1689_not0;
  wire f_arrdiv32_mux2to1689_and1;
  wire f_arrdiv32_mux2to1689_xor0;
  wire f_arrdiv32_mux2to1690_and0;
  wire f_arrdiv32_mux2to1690_not0;
  wire f_arrdiv32_mux2to1690_and1;
  wire f_arrdiv32_mux2to1690_xor0;
  wire f_arrdiv32_mux2to1691_and0;
  wire f_arrdiv32_mux2to1691_not0;
  wire f_arrdiv32_mux2to1691_and1;
  wire f_arrdiv32_mux2to1691_xor0;
  wire f_arrdiv32_mux2to1692_and0;
  wire f_arrdiv32_mux2to1692_not0;
  wire f_arrdiv32_mux2to1692_and1;
  wire f_arrdiv32_mux2to1692_xor0;
  wire f_arrdiv32_mux2to1693_and0;
  wire f_arrdiv32_mux2to1693_not0;
  wire f_arrdiv32_mux2to1693_and1;
  wire f_arrdiv32_mux2to1693_xor0;
  wire f_arrdiv32_mux2to1694_and0;
  wire f_arrdiv32_mux2to1694_not0;
  wire f_arrdiv32_mux2to1694_and1;
  wire f_arrdiv32_mux2to1694_xor0;
  wire f_arrdiv32_mux2to1695_and0;
  wire f_arrdiv32_mux2to1695_not0;
  wire f_arrdiv32_mux2to1695_and1;
  wire f_arrdiv32_mux2to1695_xor0;
  wire f_arrdiv32_mux2to1696_and0;
  wire f_arrdiv32_mux2to1696_not0;
  wire f_arrdiv32_mux2to1696_and1;
  wire f_arrdiv32_mux2to1696_xor0;
  wire f_arrdiv32_mux2to1697_and0;
  wire f_arrdiv32_mux2to1697_not0;
  wire f_arrdiv32_mux2to1697_and1;
  wire f_arrdiv32_mux2to1697_xor0;
  wire f_arrdiv32_mux2to1698_and0;
  wire f_arrdiv32_mux2to1698_not0;
  wire f_arrdiv32_mux2to1698_and1;
  wire f_arrdiv32_mux2to1698_xor0;
  wire f_arrdiv32_mux2to1699_and0;
  wire f_arrdiv32_mux2to1699_not0;
  wire f_arrdiv32_mux2to1699_and1;
  wire f_arrdiv32_mux2to1699_xor0;
  wire f_arrdiv32_mux2to1700_and0;
  wire f_arrdiv32_mux2to1700_not0;
  wire f_arrdiv32_mux2to1700_and1;
  wire f_arrdiv32_mux2to1700_xor0;
  wire f_arrdiv32_mux2to1701_and0;
  wire f_arrdiv32_mux2to1701_not0;
  wire f_arrdiv32_mux2to1701_and1;
  wire f_arrdiv32_mux2to1701_xor0;
  wire f_arrdiv32_mux2to1702_and0;
  wire f_arrdiv32_mux2to1702_not0;
  wire f_arrdiv32_mux2to1702_and1;
  wire f_arrdiv32_mux2to1702_xor0;
  wire f_arrdiv32_mux2to1703_and0;
  wire f_arrdiv32_mux2to1703_not0;
  wire f_arrdiv32_mux2to1703_and1;
  wire f_arrdiv32_mux2to1703_xor0;
  wire f_arrdiv32_mux2to1704_and0;
  wire f_arrdiv32_mux2to1704_not0;
  wire f_arrdiv32_mux2to1704_and1;
  wire f_arrdiv32_mux2to1704_xor0;
  wire f_arrdiv32_mux2to1705_and0;
  wire f_arrdiv32_mux2to1705_not0;
  wire f_arrdiv32_mux2to1705_and1;
  wire f_arrdiv32_mux2to1705_xor0;
  wire f_arrdiv32_mux2to1706_and0;
  wire f_arrdiv32_mux2to1706_not0;
  wire f_arrdiv32_mux2to1706_and1;
  wire f_arrdiv32_mux2to1706_xor0;
  wire f_arrdiv32_mux2to1707_and0;
  wire f_arrdiv32_mux2to1707_not0;
  wire f_arrdiv32_mux2to1707_and1;
  wire f_arrdiv32_mux2to1707_xor0;
  wire f_arrdiv32_mux2to1708_and0;
  wire f_arrdiv32_mux2to1708_not0;
  wire f_arrdiv32_mux2to1708_and1;
  wire f_arrdiv32_mux2to1708_xor0;
  wire f_arrdiv32_mux2to1709_and0;
  wire f_arrdiv32_mux2to1709_not0;
  wire f_arrdiv32_mux2to1709_and1;
  wire f_arrdiv32_mux2to1709_xor0;
  wire f_arrdiv32_mux2to1710_and0;
  wire f_arrdiv32_mux2to1710_not0;
  wire f_arrdiv32_mux2to1710_and1;
  wire f_arrdiv32_mux2to1710_xor0;
  wire f_arrdiv32_mux2to1711_and0;
  wire f_arrdiv32_mux2to1711_not0;
  wire f_arrdiv32_mux2to1711_and1;
  wire f_arrdiv32_mux2to1711_xor0;
  wire f_arrdiv32_mux2to1712_and0;
  wire f_arrdiv32_mux2to1712_not0;
  wire f_arrdiv32_mux2to1712_and1;
  wire f_arrdiv32_mux2to1712_xor0;
  wire f_arrdiv32_not22;
  wire f_arrdiv32_fs736_xor0;
  wire f_arrdiv32_fs736_not0;
  wire f_arrdiv32_fs736_and0;
  wire f_arrdiv32_fs736_not1;
  wire f_arrdiv32_fs737_xor0;
  wire f_arrdiv32_fs737_not0;
  wire f_arrdiv32_fs737_and0;
  wire f_arrdiv32_fs737_xor1;
  wire f_arrdiv32_fs737_not1;
  wire f_arrdiv32_fs737_and1;
  wire f_arrdiv32_fs737_or0;
  wire f_arrdiv32_fs738_xor0;
  wire f_arrdiv32_fs738_not0;
  wire f_arrdiv32_fs738_and0;
  wire f_arrdiv32_fs738_xor1;
  wire f_arrdiv32_fs738_not1;
  wire f_arrdiv32_fs738_and1;
  wire f_arrdiv32_fs738_or0;
  wire f_arrdiv32_fs739_xor0;
  wire f_arrdiv32_fs739_not0;
  wire f_arrdiv32_fs739_and0;
  wire f_arrdiv32_fs739_xor1;
  wire f_arrdiv32_fs739_not1;
  wire f_arrdiv32_fs739_and1;
  wire f_arrdiv32_fs739_or0;
  wire f_arrdiv32_fs740_xor0;
  wire f_arrdiv32_fs740_not0;
  wire f_arrdiv32_fs740_and0;
  wire f_arrdiv32_fs740_xor1;
  wire f_arrdiv32_fs740_not1;
  wire f_arrdiv32_fs740_and1;
  wire f_arrdiv32_fs740_or0;
  wire f_arrdiv32_fs741_xor0;
  wire f_arrdiv32_fs741_not0;
  wire f_arrdiv32_fs741_and0;
  wire f_arrdiv32_fs741_xor1;
  wire f_arrdiv32_fs741_not1;
  wire f_arrdiv32_fs741_and1;
  wire f_arrdiv32_fs741_or0;
  wire f_arrdiv32_fs742_xor0;
  wire f_arrdiv32_fs742_not0;
  wire f_arrdiv32_fs742_and0;
  wire f_arrdiv32_fs742_xor1;
  wire f_arrdiv32_fs742_not1;
  wire f_arrdiv32_fs742_and1;
  wire f_arrdiv32_fs742_or0;
  wire f_arrdiv32_fs743_xor0;
  wire f_arrdiv32_fs743_not0;
  wire f_arrdiv32_fs743_and0;
  wire f_arrdiv32_fs743_xor1;
  wire f_arrdiv32_fs743_not1;
  wire f_arrdiv32_fs743_and1;
  wire f_arrdiv32_fs743_or0;
  wire f_arrdiv32_fs744_xor0;
  wire f_arrdiv32_fs744_not0;
  wire f_arrdiv32_fs744_and0;
  wire f_arrdiv32_fs744_xor1;
  wire f_arrdiv32_fs744_not1;
  wire f_arrdiv32_fs744_and1;
  wire f_arrdiv32_fs744_or0;
  wire f_arrdiv32_fs745_xor0;
  wire f_arrdiv32_fs745_not0;
  wire f_arrdiv32_fs745_and0;
  wire f_arrdiv32_fs745_xor1;
  wire f_arrdiv32_fs745_not1;
  wire f_arrdiv32_fs745_and1;
  wire f_arrdiv32_fs745_or0;
  wire f_arrdiv32_fs746_xor0;
  wire f_arrdiv32_fs746_not0;
  wire f_arrdiv32_fs746_and0;
  wire f_arrdiv32_fs746_xor1;
  wire f_arrdiv32_fs746_not1;
  wire f_arrdiv32_fs746_and1;
  wire f_arrdiv32_fs746_or0;
  wire f_arrdiv32_fs747_xor0;
  wire f_arrdiv32_fs747_not0;
  wire f_arrdiv32_fs747_and0;
  wire f_arrdiv32_fs747_xor1;
  wire f_arrdiv32_fs747_not1;
  wire f_arrdiv32_fs747_and1;
  wire f_arrdiv32_fs747_or0;
  wire f_arrdiv32_fs748_xor0;
  wire f_arrdiv32_fs748_not0;
  wire f_arrdiv32_fs748_and0;
  wire f_arrdiv32_fs748_xor1;
  wire f_arrdiv32_fs748_not1;
  wire f_arrdiv32_fs748_and1;
  wire f_arrdiv32_fs748_or0;
  wire f_arrdiv32_fs749_xor0;
  wire f_arrdiv32_fs749_not0;
  wire f_arrdiv32_fs749_and0;
  wire f_arrdiv32_fs749_xor1;
  wire f_arrdiv32_fs749_not1;
  wire f_arrdiv32_fs749_and1;
  wire f_arrdiv32_fs749_or0;
  wire f_arrdiv32_fs750_xor0;
  wire f_arrdiv32_fs750_not0;
  wire f_arrdiv32_fs750_and0;
  wire f_arrdiv32_fs750_xor1;
  wire f_arrdiv32_fs750_not1;
  wire f_arrdiv32_fs750_and1;
  wire f_arrdiv32_fs750_or0;
  wire f_arrdiv32_fs751_xor0;
  wire f_arrdiv32_fs751_not0;
  wire f_arrdiv32_fs751_and0;
  wire f_arrdiv32_fs751_xor1;
  wire f_arrdiv32_fs751_not1;
  wire f_arrdiv32_fs751_and1;
  wire f_arrdiv32_fs751_or0;
  wire f_arrdiv32_fs752_xor0;
  wire f_arrdiv32_fs752_not0;
  wire f_arrdiv32_fs752_and0;
  wire f_arrdiv32_fs752_xor1;
  wire f_arrdiv32_fs752_not1;
  wire f_arrdiv32_fs752_and1;
  wire f_arrdiv32_fs752_or0;
  wire f_arrdiv32_fs753_xor0;
  wire f_arrdiv32_fs753_not0;
  wire f_arrdiv32_fs753_and0;
  wire f_arrdiv32_fs753_xor1;
  wire f_arrdiv32_fs753_not1;
  wire f_arrdiv32_fs753_and1;
  wire f_arrdiv32_fs753_or0;
  wire f_arrdiv32_fs754_xor0;
  wire f_arrdiv32_fs754_not0;
  wire f_arrdiv32_fs754_and0;
  wire f_arrdiv32_fs754_xor1;
  wire f_arrdiv32_fs754_not1;
  wire f_arrdiv32_fs754_and1;
  wire f_arrdiv32_fs754_or0;
  wire f_arrdiv32_fs755_xor0;
  wire f_arrdiv32_fs755_not0;
  wire f_arrdiv32_fs755_and0;
  wire f_arrdiv32_fs755_xor1;
  wire f_arrdiv32_fs755_not1;
  wire f_arrdiv32_fs755_and1;
  wire f_arrdiv32_fs755_or0;
  wire f_arrdiv32_fs756_xor0;
  wire f_arrdiv32_fs756_not0;
  wire f_arrdiv32_fs756_and0;
  wire f_arrdiv32_fs756_xor1;
  wire f_arrdiv32_fs756_not1;
  wire f_arrdiv32_fs756_and1;
  wire f_arrdiv32_fs756_or0;
  wire f_arrdiv32_fs757_xor0;
  wire f_arrdiv32_fs757_not0;
  wire f_arrdiv32_fs757_and0;
  wire f_arrdiv32_fs757_xor1;
  wire f_arrdiv32_fs757_not1;
  wire f_arrdiv32_fs757_and1;
  wire f_arrdiv32_fs757_or0;
  wire f_arrdiv32_fs758_xor0;
  wire f_arrdiv32_fs758_not0;
  wire f_arrdiv32_fs758_and0;
  wire f_arrdiv32_fs758_xor1;
  wire f_arrdiv32_fs758_not1;
  wire f_arrdiv32_fs758_and1;
  wire f_arrdiv32_fs758_or0;
  wire f_arrdiv32_fs759_xor0;
  wire f_arrdiv32_fs759_not0;
  wire f_arrdiv32_fs759_and0;
  wire f_arrdiv32_fs759_xor1;
  wire f_arrdiv32_fs759_not1;
  wire f_arrdiv32_fs759_and1;
  wire f_arrdiv32_fs759_or0;
  wire f_arrdiv32_fs760_xor0;
  wire f_arrdiv32_fs760_not0;
  wire f_arrdiv32_fs760_and0;
  wire f_arrdiv32_fs760_xor1;
  wire f_arrdiv32_fs760_not1;
  wire f_arrdiv32_fs760_and1;
  wire f_arrdiv32_fs760_or0;
  wire f_arrdiv32_fs761_xor0;
  wire f_arrdiv32_fs761_not0;
  wire f_arrdiv32_fs761_and0;
  wire f_arrdiv32_fs761_xor1;
  wire f_arrdiv32_fs761_not1;
  wire f_arrdiv32_fs761_and1;
  wire f_arrdiv32_fs761_or0;
  wire f_arrdiv32_fs762_xor0;
  wire f_arrdiv32_fs762_not0;
  wire f_arrdiv32_fs762_and0;
  wire f_arrdiv32_fs762_xor1;
  wire f_arrdiv32_fs762_not1;
  wire f_arrdiv32_fs762_and1;
  wire f_arrdiv32_fs762_or0;
  wire f_arrdiv32_fs763_xor0;
  wire f_arrdiv32_fs763_not0;
  wire f_arrdiv32_fs763_and0;
  wire f_arrdiv32_fs763_xor1;
  wire f_arrdiv32_fs763_not1;
  wire f_arrdiv32_fs763_and1;
  wire f_arrdiv32_fs763_or0;
  wire f_arrdiv32_fs764_xor0;
  wire f_arrdiv32_fs764_not0;
  wire f_arrdiv32_fs764_and0;
  wire f_arrdiv32_fs764_xor1;
  wire f_arrdiv32_fs764_not1;
  wire f_arrdiv32_fs764_and1;
  wire f_arrdiv32_fs764_or0;
  wire f_arrdiv32_fs765_xor0;
  wire f_arrdiv32_fs765_not0;
  wire f_arrdiv32_fs765_and0;
  wire f_arrdiv32_fs765_xor1;
  wire f_arrdiv32_fs765_not1;
  wire f_arrdiv32_fs765_and1;
  wire f_arrdiv32_fs765_or0;
  wire f_arrdiv32_fs766_xor0;
  wire f_arrdiv32_fs766_not0;
  wire f_arrdiv32_fs766_and0;
  wire f_arrdiv32_fs766_xor1;
  wire f_arrdiv32_fs766_not1;
  wire f_arrdiv32_fs766_and1;
  wire f_arrdiv32_fs766_or0;
  wire f_arrdiv32_fs767_xor0;
  wire f_arrdiv32_fs767_not0;
  wire f_arrdiv32_fs767_and0;
  wire f_arrdiv32_fs767_xor1;
  wire f_arrdiv32_fs767_not1;
  wire f_arrdiv32_fs767_and1;
  wire f_arrdiv32_fs767_or0;
  wire f_arrdiv32_mux2to1713_and0;
  wire f_arrdiv32_mux2to1713_not0;
  wire f_arrdiv32_mux2to1713_and1;
  wire f_arrdiv32_mux2to1713_xor0;
  wire f_arrdiv32_mux2to1714_and0;
  wire f_arrdiv32_mux2to1714_not0;
  wire f_arrdiv32_mux2to1714_and1;
  wire f_arrdiv32_mux2to1714_xor0;
  wire f_arrdiv32_mux2to1715_and0;
  wire f_arrdiv32_mux2to1715_not0;
  wire f_arrdiv32_mux2to1715_and1;
  wire f_arrdiv32_mux2to1715_xor0;
  wire f_arrdiv32_mux2to1716_and0;
  wire f_arrdiv32_mux2to1716_not0;
  wire f_arrdiv32_mux2to1716_and1;
  wire f_arrdiv32_mux2to1716_xor0;
  wire f_arrdiv32_mux2to1717_and0;
  wire f_arrdiv32_mux2to1717_not0;
  wire f_arrdiv32_mux2to1717_and1;
  wire f_arrdiv32_mux2to1717_xor0;
  wire f_arrdiv32_mux2to1718_and0;
  wire f_arrdiv32_mux2to1718_not0;
  wire f_arrdiv32_mux2to1718_and1;
  wire f_arrdiv32_mux2to1718_xor0;
  wire f_arrdiv32_mux2to1719_and0;
  wire f_arrdiv32_mux2to1719_not0;
  wire f_arrdiv32_mux2to1719_and1;
  wire f_arrdiv32_mux2to1719_xor0;
  wire f_arrdiv32_mux2to1720_and0;
  wire f_arrdiv32_mux2to1720_not0;
  wire f_arrdiv32_mux2to1720_and1;
  wire f_arrdiv32_mux2to1720_xor0;
  wire f_arrdiv32_mux2to1721_and0;
  wire f_arrdiv32_mux2to1721_not0;
  wire f_arrdiv32_mux2to1721_and1;
  wire f_arrdiv32_mux2to1721_xor0;
  wire f_arrdiv32_mux2to1722_and0;
  wire f_arrdiv32_mux2to1722_not0;
  wire f_arrdiv32_mux2to1722_and1;
  wire f_arrdiv32_mux2to1722_xor0;
  wire f_arrdiv32_mux2to1723_and0;
  wire f_arrdiv32_mux2to1723_not0;
  wire f_arrdiv32_mux2to1723_and1;
  wire f_arrdiv32_mux2to1723_xor0;
  wire f_arrdiv32_mux2to1724_and0;
  wire f_arrdiv32_mux2to1724_not0;
  wire f_arrdiv32_mux2to1724_and1;
  wire f_arrdiv32_mux2to1724_xor0;
  wire f_arrdiv32_mux2to1725_and0;
  wire f_arrdiv32_mux2to1725_not0;
  wire f_arrdiv32_mux2to1725_and1;
  wire f_arrdiv32_mux2to1725_xor0;
  wire f_arrdiv32_mux2to1726_and0;
  wire f_arrdiv32_mux2to1726_not0;
  wire f_arrdiv32_mux2to1726_and1;
  wire f_arrdiv32_mux2to1726_xor0;
  wire f_arrdiv32_mux2to1727_and0;
  wire f_arrdiv32_mux2to1727_not0;
  wire f_arrdiv32_mux2to1727_and1;
  wire f_arrdiv32_mux2to1727_xor0;
  wire f_arrdiv32_mux2to1728_and0;
  wire f_arrdiv32_mux2to1728_not0;
  wire f_arrdiv32_mux2to1728_and1;
  wire f_arrdiv32_mux2to1728_xor0;
  wire f_arrdiv32_mux2to1729_and0;
  wire f_arrdiv32_mux2to1729_not0;
  wire f_arrdiv32_mux2to1729_and1;
  wire f_arrdiv32_mux2to1729_xor0;
  wire f_arrdiv32_mux2to1730_and0;
  wire f_arrdiv32_mux2to1730_not0;
  wire f_arrdiv32_mux2to1730_and1;
  wire f_arrdiv32_mux2to1730_xor0;
  wire f_arrdiv32_mux2to1731_and0;
  wire f_arrdiv32_mux2to1731_not0;
  wire f_arrdiv32_mux2to1731_and1;
  wire f_arrdiv32_mux2to1731_xor0;
  wire f_arrdiv32_mux2to1732_and0;
  wire f_arrdiv32_mux2to1732_not0;
  wire f_arrdiv32_mux2to1732_and1;
  wire f_arrdiv32_mux2to1732_xor0;
  wire f_arrdiv32_mux2to1733_and0;
  wire f_arrdiv32_mux2to1733_not0;
  wire f_arrdiv32_mux2to1733_and1;
  wire f_arrdiv32_mux2to1733_xor0;
  wire f_arrdiv32_mux2to1734_and0;
  wire f_arrdiv32_mux2to1734_not0;
  wire f_arrdiv32_mux2to1734_and1;
  wire f_arrdiv32_mux2to1734_xor0;
  wire f_arrdiv32_mux2to1735_and0;
  wire f_arrdiv32_mux2to1735_not0;
  wire f_arrdiv32_mux2to1735_and1;
  wire f_arrdiv32_mux2to1735_xor0;
  wire f_arrdiv32_mux2to1736_and0;
  wire f_arrdiv32_mux2to1736_not0;
  wire f_arrdiv32_mux2to1736_and1;
  wire f_arrdiv32_mux2to1736_xor0;
  wire f_arrdiv32_mux2to1737_and0;
  wire f_arrdiv32_mux2to1737_not0;
  wire f_arrdiv32_mux2to1737_and1;
  wire f_arrdiv32_mux2to1737_xor0;
  wire f_arrdiv32_mux2to1738_and0;
  wire f_arrdiv32_mux2to1738_not0;
  wire f_arrdiv32_mux2to1738_and1;
  wire f_arrdiv32_mux2to1738_xor0;
  wire f_arrdiv32_mux2to1739_and0;
  wire f_arrdiv32_mux2to1739_not0;
  wire f_arrdiv32_mux2to1739_and1;
  wire f_arrdiv32_mux2to1739_xor0;
  wire f_arrdiv32_mux2to1740_and0;
  wire f_arrdiv32_mux2to1740_not0;
  wire f_arrdiv32_mux2to1740_and1;
  wire f_arrdiv32_mux2to1740_xor0;
  wire f_arrdiv32_mux2to1741_and0;
  wire f_arrdiv32_mux2to1741_not0;
  wire f_arrdiv32_mux2to1741_and1;
  wire f_arrdiv32_mux2to1741_xor0;
  wire f_arrdiv32_mux2to1742_and0;
  wire f_arrdiv32_mux2to1742_not0;
  wire f_arrdiv32_mux2to1742_and1;
  wire f_arrdiv32_mux2to1742_xor0;
  wire f_arrdiv32_mux2to1743_and0;
  wire f_arrdiv32_mux2to1743_not0;
  wire f_arrdiv32_mux2to1743_and1;
  wire f_arrdiv32_mux2to1743_xor0;
  wire f_arrdiv32_not23;
  wire f_arrdiv32_fs768_xor0;
  wire f_arrdiv32_fs768_not0;
  wire f_arrdiv32_fs768_and0;
  wire f_arrdiv32_fs768_not1;
  wire f_arrdiv32_fs769_xor0;
  wire f_arrdiv32_fs769_not0;
  wire f_arrdiv32_fs769_and0;
  wire f_arrdiv32_fs769_xor1;
  wire f_arrdiv32_fs769_not1;
  wire f_arrdiv32_fs769_and1;
  wire f_arrdiv32_fs769_or0;
  wire f_arrdiv32_fs770_xor0;
  wire f_arrdiv32_fs770_not0;
  wire f_arrdiv32_fs770_and0;
  wire f_arrdiv32_fs770_xor1;
  wire f_arrdiv32_fs770_not1;
  wire f_arrdiv32_fs770_and1;
  wire f_arrdiv32_fs770_or0;
  wire f_arrdiv32_fs771_xor0;
  wire f_arrdiv32_fs771_not0;
  wire f_arrdiv32_fs771_and0;
  wire f_arrdiv32_fs771_xor1;
  wire f_arrdiv32_fs771_not1;
  wire f_arrdiv32_fs771_and1;
  wire f_arrdiv32_fs771_or0;
  wire f_arrdiv32_fs772_xor0;
  wire f_arrdiv32_fs772_not0;
  wire f_arrdiv32_fs772_and0;
  wire f_arrdiv32_fs772_xor1;
  wire f_arrdiv32_fs772_not1;
  wire f_arrdiv32_fs772_and1;
  wire f_arrdiv32_fs772_or0;
  wire f_arrdiv32_fs773_xor0;
  wire f_arrdiv32_fs773_not0;
  wire f_arrdiv32_fs773_and0;
  wire f_arrdiv32_fs773_xor1;
  wire f_arrdiv32_fs773_not1;
  wire f_arrdiv32_fs773_and1;
  wire f_arrdiv32_fs773_or0;
  wire f_arrdiv32_fs774_xor0;
  wire f_arrdiv32_fs774_not0;
  wire f_arrdiv32_fs774_and0;
  wire f_arrdiv32_fs774_xor1;
  wire f_arrdiv32_fs774_not1;
  wire f_arrdiv32_fs774_and1;
  wire f_arrdiv32_fs774_or0;
  wire f_arrdiv32_fs775_xor0;
  wire f_arrdiv32_fs775_not0;
  wire f_arrdiv32_fs775_and0;
  wire f_arrdiv32_fs775_xor1;
  wire f_arrdiv32_fs775_not1;
  wire f_arrdiv32_fs775_and1;
  wire f_arrdiv32_fs775_or0;
  wire f_arrdiv32_fs776_xor0;
  wire f_arrdiv32_fs776_not0;
  wire f_arrdiv32_fs776_and0;
  wire f_arrdiv32_fs776_xor1;
  wire f_arrdiv32_fs776_not1;
  wire f_arrdiv32_fs776_and1;
  wire f_arrdiv32_fs776_or0;
  wire f_arrdiv32_fs777_xor0;
  wire f_arrdiv32_fs777_not0;
  wire f_arrdiv32_fs777_and0;
  wire f_arrdiv32_fs777_xor1;
  wire f_arrdiv32_fs777_not1;
  wire f_arrdiv32_fs777_and1;
  wire f_arrdiv32_fs777_or0;
  wire f_arrdiv32_fs778_xor0;
  wire f_arrdiv32_fs778_not0;
  wire f_arrdiv32_fs778_and0;
  wire f_arrdiv32_fs778_xor1;
  wire f_arrdiv32_fs778_not1;
  wire f_arrdiv32_fs778_and1;
  wire f_arrdiv32_fs778_or0;
  wire f_arrdiv32_fs779_xor0;
  wire f_arrdiv32_fs779_not0;
  wire f_arrdiv32_fs779_and0;
  wire f_arrdiv32_fs779_xor1;
  wire f_arrdiv32_fs779_not1;
  wire f_arrdiv32_fs779_and1;
  wire f_arrdiv32_fs779_or0;
  wire f_arrdiv32_fs780_xor0;
  wire f_arrdiv32_fs780_not0;
  wire f_arrdiv32_fs780_and0;
  wire f_arrdiv32_fs780_xor1;
  wire f_arrdiv32_fs780_not1;
  wire f_arrdiv32_fs780_and1;
  wire f_arrdiv32_fs780_or0;
  wire f_arrdiv32_fs781_xor0;
  wire f_arrdiv32_fs781_not0;
  wire f_arrdiv32_fs781_and0;
  wire f_arrdiv32_fs781_xor1;
  wire f_arrdiv32_fs781_not1;
  wire f_arrdiv32_fs781_and1;
  wire f_arrdiv32_fs781_or0;
  wire f_arrdiv32_fs782_xor0;
  wire f_arrdiv32_fs782_not0;
  wire f_arrdiv32_fs782_and0;
  wire f_arrdiv32_fs782_xor1;
  wire f_arrdiv32_fs782_not1;
  wire f_arrdiv32_fs782_and1;
  wire f_arrdiv32_fs782_or0;
  wire f_arrdiv32_fs783_xor0;
  wire f_arrdiv32_fs783_not0;
  wire f_arrdiv32_fs783_and0;
  wire f_arrdiv32_fs783_xor1;
  wire f_arrdiv32_fs783_not1;
  wire f_arrdiv32_fs783_and1;
  wire f_arrdiv32_fs783_or0;
  wire f_arrdiv32_fs784_xor0;
  wire f_arrdiv32_fs784_not0;
  wire f_arrdiv32_fs784_and0;
  wire f_arrdiv32_fs784_xor1;
  wire f_arrdiv32_fs784_not1;
  wire f_arrdiv32_fs784_and1;
  wire f_arrdiv32_fs784_or0;
  wire f_arrdiv32_fs785_xor0;
  wire f_arrdiv32_fs785_not0;
  wire f_arrdiv32_fs785_and0;
  wire f_arrdiv32_fs785_xor1;
  wire f_arrdiv32_fs785_not1;
  wire f_arrdiv32_fs785_and1;
  wire f_arrdiv32_fs785_or0;
  wire f_arrdiv32_fs786_xor0;
  wire f_arrdiv32_fs786_not0;
  wire f_arrdiv32_fs786_and0;
  wire f_arrdiv32_fs786_xor1;
  wire f_arrdiv32_fs786_not1;
  wire f_arrdiv32_fs786_and1;
  wire f_arrdiv32_fs786_or0;
  wire f_arrdiv32_fs787_xor0;
  wire f_arrdiv32_fs787_not0;
  wire f_arrdiv32_fs787_and0;
  wire f_arrdiv32_fs787_xor1;
  wire f_arrdiv32_fs787_not1;
  wire f_arrdiv32_fs787_and1;
  wire f_arrdiv32_fs787_or0;
  wire f_arrdiv32_fs788_xor0;
  wire f_arrdiv32_fs788_not0;
  wire f_arrdiv32_fs788_and0;
  wire f_arrdiv32_fs788_xor1;
  wire f_arrdiv32_fs788_not1;
  wire f_arrdiv32_fs788_and1;
  wire f_arrdiv32_fs788_or0;
  wire f_arrdiv32_fs789_xor0;
  wire f_arrdiv32_fs789_not0;
  wire f_arrdiv32_fs789_and0;
  wire f_arrdiv32_fs789_xor1;
  wire f_arrdiv32_fs789_not1;
  wire f_arrdiv32_fs789_and1;
  wire f_arrdiv32_fs789_or0;
  wire f_arrdiv32_fs790_xor0;
  wire f_arrdiv32_fs790_not0;
  wire f_arrdiv32_fs790_and0;
  wire f_arrdiv32_fs790_xor1;
  wire f_arrdiv32_fs790_not1;
  wire f_arrdiv32_fs790_and1;
  wire f_arrdiv32_fs790_or0;
  wire f_arrdiv32_fs791_xor0;
  wire f_arrdiv32_fs791_not0;
  wire f_arrdiv32_fs791_and0;
  wire f_arrdiv32_fs791_xor1;
  wire f_arrdiv32_fs791_not1;
  wire f_arrdiv32_fs791_and1;
  wire f_arrdiv32_fs791_or0;
  wire f_arrdiv32_fs792_xor0;
  wire f_arrdiv32_fs792_not0;
  wire f_arrdiv32_fs792_and0;
  wire f_arrdiv32_fs792_xor1;
  wire f_arrdiv32_fs792_not1;
  wire f_arrdiv32_fs792_and1;
  wire f_arrdiv32_fs792_or0;
  wire f_arrdiv32_fs793_xor0;
  wire f_arrdiv32_fs793_not0;
  wire f_arrdiv32_fs793_and0;
  wire f_arrdiv32_fs793_xor1;
  wire f_arrdiv32_fs793_not1;
  wire f_arrdiv32_fs793_and1;
  wire f_arrdiv32_fs793_or0;
  wire f_arrdiv32_fs794_xor0;
  wire f_arrdiv32_fs794_not0;
  wire f_arrdiv32_fs794_and0;
  wire f_arrdiv32_fs794_xor1;
  wire f_arrdiv32_fs794_not1;
  wire f_arrdiv32_fs794_and1;
  wire f_arrdiv32_fs794_or0;
  wire f_arrdiv32_fs795_xor0;
  wire f_arrdiv32_fs795_not0;
  wire f_arrdiv32_fs795_and0;
  wire f_arrdiv32_fs795_xor1;
  wire f_arrdiv32_fs795_not1;
  wire f_arrdiv32_fs795_and1;
  wire f_arrdiv32_fs795_or0;
  wire f_arrdiv32_fs796_xor0;
  wire f_arrdiv32_fs796_not0;
  wire f_arrdiv32_fs796_and0;
  wire f_arrdiv32_fs796_xor1;
  wire f_arrdiv32_fs796_not1;
  wire f_arrdiv32_fs796_and1;
  wire f_arrdiv32_fs796_or0;
  wire f_arrdiv32_fs797_xor0;
  wire f_arrdiv32_fs797_not0;
  wire f_arrdiv32_fs797_and0;
  wire f_arrdiv32_fs797_xor1;
  wire f_arrdiv32_fs797_not1;
  wire f_arrdiv32_fs797_and1;
  wire f_arrdiv32_fs797_or0;
  wire f_arrdiv32_fs798_xor0;
  wire f_arrdiv32_fs798_not0;
  wire f_arrdiv32_fs798_and0;
  wire f_arrdiv32_fs798_xor1;
  wire f_arrdiv32_fs798_not1;
  wire f_arrdiv32_fs798_and1;
  wire f_arrdiv32_fs798_or0;
  wire f_arrdiv32_fs799_xor0;
  wire f_arrdiv32_fs799_not0;
  wire f_arrdiv32_fs799_and0;
  wire f_arrdiv32_fs799_xor1;
  wire f_arrdiv32_fs799_not1;
  wire f_arrdiv32_fs799_and1;
  wire f_arrdiv32_fs799_or0;
  wire f_arrdiv32_mux2to1744_and0;
  wire f_arrdiv32_mux2to1744_not0;
  wire f_arrdiv32_mux2to1744_and1;
  wire f_arrdiv32_mux2to1744_xor0;
  wire f_arrdiv32_mux2to1745_and0;
  wire f_arrdiv32_mux2to1745_not0;
  wire f_arrdiv32_mux2to1745_and1;
  wire f_arrdiv32_mux2to1745_xor0;
  wire f_arrdiv32_mux2to1746_and0;
  wire f_arrdiv32_mux2to1746_not0;
  wire f_arrdiv32_mux2to1746_and1;
  wire f_arrdiv32_mux2to1746_xor0;
  wire f_arrdiv32_mux2to1747_and0;
  wire f_arrdiv32_mux2to1747_not0;
  wire f_arrdiv32_mux2to1747_and1;
  wire f_arrdiv32_mux2to1747_xor0;
  wire f_arrdiv32_mux2to1748_and0;
  wire f_arrdiv32_mux2to1748_not0;
  wire f_arrdiv32_mux2to1748_and1;
  wire f_arrdiv32_mux2to1748_xor0;
  wire f_arrdiv32_mux2to1749_and0;
  wire f_arrdiv32_mux2to1749_not0;
  wire f_arrdiv32_mux2to1749_and1;
  wire f_arrdiv32_mux2to1749_xor0;
  wire f_arrdiv32_mux2to1750_and0;
  wire f_arrdiv32_mux2to1750_not0;
  wire f_arrdiv32_mux2to1750_and1;
  wire f_arrdiv32_mux2to1750_xor0;
  wire f_arrdiv32_mux2to1751_and0;
  wire f_arrdiv32_mux2to1751_not0;
  wire f_arrdiv32_mux2to1751_and1;
  wire f_arrdiv32_mux2to1751_xor0;
  wire f_arrdiv32_mux2to1752_and0;
  wire f_arrdiv32_mux2to1752_not0;
  wire f_arrdiv32_mux2to1752_and1;
  wire f_arrdiv32_mux2to1752_xor0;
  wire f_arrdiv32_mux2to1753_and0;
  wire f_arrdiv32_mux2to1753_not0;
  wire f_arrdiv32_mux2to1753_and1;
  wire f_arrdiv32_mux2to1753_xor0;
  wire f_arrdiv32_mux2to1754_and0;
  wire f_arrdiv32_mux2to1754_not0;
  wire f_arrdiv32_mux2to1754_and1;
  wire f_arrdiv32_mux2to1754_xor0;
  wire f_arrdiv32_mux2to1755_and0;
  wire f_arrdiv32_mux2to1755_not0;
  wire f_arrdiv32_mux2to1755_and1;
  wire f_arrdiv32_mux2to1755_xor0;
  wire f_arrdiv32_mux2to1756_and0;
  wire f_arrdiv32_mux2to1756_not0;
  wire f_arrdiv32_mux2to1756_and1;
  wire f_arrdiv32_mux2to1756_xor0;
  wire f_arrdiv32_mux2to1757_and0;
  wire f_arrdiv32_mux2to1757_not0;
  wire f_arrdiv32_mux2to1757_and1;
  wire f_arrdiv32_mux2to1757_xor0;
  wire f_arrdiv32_mux2to1758_and0;
  wire f_arrdiv32_mux2to1758_not0;
  wire f_arrdiv32_mux2to1758_and1;
  wire f_arrdiv32_mux2to1758_xor0;
  wire f_arrdiv32_mux2to1759_and0;
  wire f_arrdiv32_mux2to1759_not0;
  wire f_arrdiv32_mux2to1759_and1;
  wire f_arrdiv32_mux2to1759_xor0;
  wire f_arrdiv32_mux2to1760_and0;
  wire f_arrdiv32_mux2to1760_not0;
  wire f_arrdiv32_mux2to1760_and1;
  wire f_arrdiv32_mux2to1760_xor0;
  wire f_arrdiv32_mux2to1761_and0;
  wire f_arrdiv32_mux2to1761_not0;
  wire f_arrdiv32_mux2to1761_and1;
  wire f_arrdiv32_mux2to1761_xor0;
  wire f_arrdiv32_mux2to1762_and0;
  wire f_arrdiv32_mux2to1762_not0;
  wire f_arrdiv32_mux2to1762_and1;
  wire f_arrdiv32_mux2to1762_xor0;
  wire f_arrdiv32_mux2to1763_and0;
  wire f_arrdiv32_mux2to1763_not0;
  wire f_arrdiv32_mux2to1763_and1;
  wire f_arrdiv32_mux2to1763_xor0;
  wire f_arrdiv32_mux2to1764_and0;
  wire f_arrdiv32_mux2to1764_not0;
  wire f_arrdiv32_mux2to1764_and1;
  wire f_arrdiv32_mux2to1764_xor0;
  wire f_arrdiv32_mux2to1765_and0;
  wire f_arrdiv32_mux2to1765_not0;
  wire f_arrdiv32_mux2to1765_and1;
  wire f_arrdiv32_mux2to1765_xor0;
  wire f_arrdiv32_mux2to1766_and0;
  wire f_arrdiv32_mux2to1766_not0;
  wire f_arrdiv32_mux2to1766_and1;
  wire f_arrdiv32_mux2to1766_xor0;
  wire f_arrdiv32_mux2to1767_and0;
  wire f_arrdiv32_mux2to1767_not0;
  wire f_arrdiv32_mux2to1767_and1;
  wire f_arrdiv32_mux2to1767_xor0;
  wire f_arrdiv32_mux2to1768_and0;
  wire f_arrdiv32_mux2to1768_not0;
  wire f_arrdiv32_mux2to1768_and1;
  wire f_arrdiv32_mux2to1768_xor0;
  wire f_arrdiv32_mux2to1769_and0;
  wire f_arrdiv32_mux2to1769_not0;
  wire f_arrdiv32_mux2to1769_and1;
  wire f_arrdiv32_mux2to1769_xor0;
  wire f_arrdiv32_mux2to1770_and0;
  wire f_arrdiv32_mux2to1770_not0;
  wire f_arrdiv32_mux2to1770_and1;
  wire f_arrdiv32_mux2to1770_xor0;
  wire f_arrdiv32_mux2to1771_and0;
  wire f_arrdiv32_mux2to1771_not0;
  wire f_arrdiv32_mux2to1771_and1;
  wire f_arrdiv32_mux2to1771_xor0;
  wire f_arrdiv32_mux2to1772_and0;
  wire f_arrdiv32_mux2to1772_not0;
  wire f_arrdiv32_mux2to1772_and1;
  wire f_arrdiv32_mux2to1772_xor0;
  wire f_arrdiv32_mux2to1773_and0;
  wire f_arrdiv32_mux2to1773_not0;
  wire f_arrdiv32_mux2to1773_and1;
  wire f_arrdiv32_mux2to1773_xor0;
  wire f_arrdiv32_mux2to1774_and0;
  wire f_arrdiv32_mux2to1774_not0;
  wire f_arrdiv32_mux2to1774_and1;
  wire f_arrdiv32_mux2to1774_xor0;
  wire f_arrdiv32_not24;
  wire f_arrdiv32_fs800_xor0;
  wire f_arrdiv32_fs800_not0;
  wire f_arrdiv32_fs800_and0;
  wire f_arrdiv32_fs800_not1;
  wire f_arrdiv32_fs801_xor0;
  wire f_arrdiv32_fs801_not0;
  wire f_arrdiv32_fs801_and0;
  wire f_arrdiv32_fs801_xor1;
  wire f_arrdiv32_fs801_not1;
  wire f_arrdiv32_fs801_and1;
  wire f_arrdiv32_fs801_or0;
  wire f_arrdiv32_fs802_xor0;
  wire f_arrdiv32_fs802_not0;
  wire f_arrdiv32_fs802_and0;
  wire f_arrdiv32_fs802_xor1;
  wire f_arrdiv32_fs802_not1;
  wire f_arrdiv32_fs802_and1;
  wire f_arrdiv32_fs802_or0;
  wire f_arrdiv32_fs803_xor0;
  wire f_arrdiv32_fs803_not0;
  wire f_arrdiv32_fs803_and0;
  wire f_arrdiv32_fs803_xor1;
  wire f_arrdiv32_fs803_not1;
  wire f_arrdiv32_fs803_and1;
  wire f_arrdiv32_fs803_or0;
  wire f_arrdiv32_fs804_xor0;
  wire f_arrdiv32_fs804_not0;
  wire f_arrdiv32_fs804_and0;
  wire f_arrdiv32_fs804_xor1;
  wire f_arrdiv32_fs804_not1;
  wire f_arrdiv32_fs804_and1;
  wire f_arrdiv32_fs804_or0;
  wire f_arrdiv32_fs805_xor0;
  wire f_arrdiv32_fs805_not0;
  wire f_arrdiv32_fs805_and0;
  wire f_arrdiv32_fs805_xor1;
  wire f_arrdiv32_fs805_not1;
  wire f_arrdiv32_fs805_and1;
  wire f_arrdiv32_fs805_or0;
  wire f_arrdiv32_fs806_xor0;
  wire f_arrdiv32_fs806_not0;
  wire f_arrdiv32_fs806_and0;
  wire f_arrdiv32_fs806_xor1;
  wire f_arrdiv32_fs806_not1;
  wire f_arrdiv32_fs806_and1;
  wire f_arrdiv32_fs806_or0;
  wire f_arrdiv32_fs807_xor0;
  wire f_arrdiv32_fs807_not0;
  wire f_arrdiv32_fs807_and0;
  wire f_arrdiv32_fs807_xor1;
  wire f_arrdiv32_fs807_not1;
  wire f_arrdiv32_fs807_and1;
  wire f_arrdiv32_fs807_or0;
  wire f_arrdiv32_fs808_xor0;
  wire f_arrdiv32_fs808_not0;
  wire f_arrdiv32_fs808_and0;
  wire f_arrdiv32_fs808_xor1;
  wire f_arrdiv32_fs808_not1;
  wire f_arrdiv32_fs808_and1;
  wire f_arrdiv32_fs808_or0;
  wire f_arrdiv32_fs809_xor0;
  wire f_arrdiv32_fs809_not0;
  wire f_arrdiv32_fs809_and0;
  wire f_arrdiv32_fs809_xor1;
  wire f_arrdiv32_fs809_not1;
  wire f_arrdiv32_fs809_and1;
  wire f_arrdiv32_fs809_or0;
  wire f_arrdiv32_fs810_xor0;
  wire f_arrdiv32_fs810_not0;
  wire f_arrdiv32_fs810_and0;
  wire f_arrdiv32_fs810_xor1;
  wire f_arrdiv32_fs810_not1;
  wire f_arrdiv32_fs810_and1;
  wire f_arrdiv32_fs810_or0;
  wire f_arrdiv32_fs811_xor0;
  wire f_arrdiv32_fs811_not0;
  wire f_arrdiv32_fs811_and0;
  wire f_arrdiv32_fs811_xor1;
  wire f_arrdiv32_fs811_not1;
  wire f_arrdiv32_fs811_and1;
  wire f_arrdiv32_fs811_or0;
  wire f_arrdiv32_fs812_xor0;
  wire f_arrdiv32_fs812_not0;
  wire f_arrdiv32_fs812_and0;
  wire f_arrdiv32_fs812_xor1;
  wire f_arrdiv32_fs812_not1;
  wire f_arrdiv32_fs812_and1;
  wire f_arrdiv32_fs812_or0;
  wire f_arrdiv32_fs813_xor0;
  wire f_arrdiv32_fs813_not0;
  wire f_arrdiv32_fs813_and0;
  wire f_arrdiv32_fs813_xor1;
  wire f_arrdiv32_fs813_not1;
  wire f_arrdiv32_fs813_and1;
  wire f_arrdiv32_fs813_or0;
  wire f_arrdiv32_fs814_xor0;
  wire f_arrdiv32_fs814_not0;
  wire f_arrdiv32_fs814_and0;
  wire f_arrdiv32_fs814_xor1;
  wire f_arrdiv32_fs814_not1;
  wire f_arrdiv32_fs814_and1;
  wire f_arrdiv32_fs814_or0;
  wire f_arrdiv32_fs815_xor0;
  wire f_arrdiv32_fs815_not0;
  wire f_arrdiv32_fs815_and0;
  wire f_arrdiv32_fs815_xor1;
  wire f_arrdiv32_fs815_not1;
  wire f_arrdiv32_fs815_and1;
  wire f_arrdiv32_fs815_or0;
  wire f_arrdiv32_fs816_xor0;
  wire f_arrdiv32_fs816_not0;
  wire f_arrdiv32_fs816_and0;
  wire f_arrdiv32_fs816_xor1;
  wire f_arrdiv32_fs816_not1;
  wire f_arrdiv32_fs816_and1;
  wire f_arrdiv32_fs816_or0;
  wire f_arrdiv32_fs817_xor0;
  wire f_arrdiv32_fs817_not0;
  wire f_arrdiv32_fs817_and0;
  wire f_arrdiv32_fs817_xor1;
  wire f_arrdiv32_fs817_not1;
  wire f_arrdiv32_fs817_and1;
  wire f_arrdiv32_fs817_or0;
  wire f_arrdiv32_fs818_xor0;
  wire f_arrdiv32_fs818_not0;
  wire f_arrdiv32_fs818_and0;
  wire f_arrdiv32_fs818_xor1;
  wire f_arrdiv32_fs818_not1;
  wire f_arrdiv32_fs818_and1;
  wire f_arrdiv32_fs818_or0;
  wire f_arrdiv32_fs819_xor0;
  wire f_arrdiv32_fs819_not0;
  wire f_arrdiv32_fs819_and0;
  wire f_arrdiv32_fs819_xor1;
  wire f_arrdiv32_fs819_not1;
  wire f_arrdiv32_fs819_and1;
  wire f_arrdiv32_fs819_or0;
  wire f_arrdiv32_fs820_xor0;
  wire f_arrdiv32_fs820_not0;
  wire f_arrdiv32_fs820_and0;
  wire f_arrdiv32_fs820_xor1;
  wire f_arrdiv32_fs820_not1;
  wire f_arrdiv32_fs820_and1;
  wire f_arrdiv32_fs820_or0;
  wire f_arrdiv32_fs821_xor0;
  wire f_arrdiv32_fs821_not0;
  wire f_arrdiv32_fs821_and0;
  wire f_arrdiv32_fs821_xor1;
  wire f_arrdiv32_fs821_not1;
  wire f_arrdiv32_fs821_and1;
  wire f_arrdiv32_fs821_or0;
  wire f_arrdiv32_fs822_xor0;
  wire f_arrdiv32_fs822_not0;
  wire f_arrdiv32_fs822_and0;
  wire f_arrdiv32_fs822_xor1;
  wire f_arrdiv32_fs822_not1;
  wire f_arrdiv32_fs822_and1;
  wire f_arrdiv32_fs822_or0;
  wire f_arrdiv32_fs823_xor0;
  wire f_arrdiv32_fs823_not0;
  wire f_arrdiv32_fs823_and0;
  wire f_arrdiv32_fs823_xor1;
  wire f_arrdiv32_fs823_not1;
  wire f_arrdiv32_fs823_and1;
  wire f_arrdiv32_fs823_or0;
  wire f_arrdiv32_fs824_xor0;
  wire f_arrdiv32_fs824_not0;
  wire f_arrdiv32_fs824_and0;
  wire f_arrdiv32_fs824_xor1;
  wire f_arrdiv32_fs824_not1;
  wire f_arrdiv32_fs824_and1;
  wire f_arrdiv32_fs824_or0;
  wire f_arrdiv32_fs825_xor0;
  wire f_arrdiv32_fs825_not0;
  wire f_arrdiv32_fs825_and0;
  wire f_arrdiv32_fs825_xor1;
  wire f_arrdiv32_fs825_not1;
  wire f_arrdiv32_fs825_and1;
  wire f_arrdiv32_fs825_or0;
  wire f_arrdiv32_fs826_xor0;
  wire f_arrdiv32_fs826_not0;
  wire f_arrdiv32_fs826_and0;
  wire f_arrdiv32_fs826_xor1;
  wire f_arrdiv32_fs826_not1;
  wire f_arrdiv32_fs826_and1;
  wire f_arrdiv32_fs826_or0;
  wire f_arrdiv32_fs827_xor0;
  wire f_arrdiv32_fs827_not0;
  wire f_arrdiv32_fs827_and0;
  wire f_arrdiv32_fs827_xor1;
  wire f_arrdiv32_fs827_not1;
  wire f_arrdiv32_fs827_and1;
  wire f_arrdiv32_fs827_or0;
  wire f_arrdiv32_fs828_xor0;
  wire f_arrdiv32_fs828_not0;
  wire f_arrdiv32_fs828_and0;
  wire f_arrdiv32_fs828_xor1;
  wire f_arrdiv32_fs828_not1;
  wire f_arrdiv32_fs828_and1;
  wire f_arrdiv32_fs828_or0;
  wire f_arrdiv32_fs829_xor0;
  wire f_arrdiv32_fs829_not0;
  wire f_arrdiv32_fs829_and0;
  wire f_arrdiv32_fs829_xor1;
  wire f_arrdiv32_fs829_not1;
  wire f_arrdiv32_fs829_and1;
  wire f_arrdiv32_fs829_or0;
  wire f_arrdiv32_fs830_xor0;
  wire f_arrdiv32_fs830_not0;
  wire f_arrdiv32_fs830_and0;
  wire f_arrdiv32_fs830_xor1;
  wire f_arrdiv32_fs830_not1;
  wire f_arrdiv32_fs830_and1;
  wire f_arrdiv32_fs830_or0;
  wire f_arrdiv32_fs831_xor0;
  wire f_arrdiv32_fs831_not0;
  wire f_arrdiv32_fs831_and0;
  wire f_arrdiv32_fs831_xor1;
  wire f_arrdiv32_fs831_not1;
  wire f_arrdiv32_fs831_and1;
  wire f_arrdiv32_fs831_or0;
  wire f_arrdiv32_mux2to1775_and0;
  wire f_arrdiv32_mux2to1775_not0;
  wire f_arrdiv32_mux2to1775_and1;
  wire f_arrdiv32_mux2to1775_xor0;
  wire f_arrdiv32_mux2to1776_and0;
  wire f_arrdiv32_mux2to1776_not0;
  wire f_arrdiv32_mux2to1776_and1;
  wire f_arrdiv32_mux2to1776_xor0;
  wire f_arrdiv32_mux2to1777_and0;
  wire f_arrdiv32_mux2to1777_not0;
  wire f_arrdiv32_mux2to1777_and1;
  wire f_arrdiv32_mux2to1777_xor0;
  wire f_arrdiv32_mux2to1778_and0;
  wire f_arrdiv32_mux2to1778_not0;
  wire f_arrdiv32_mux2to1778_and1;
  wire f_arrdiv32_mux2to1778_xor0;
  wire f_arrdiv32_mux2to1779_and0;
  wire f_arrdiv32_mux2to1779_not0;
  wire f_arrdiv32_mux2to1779_and1;
  wire f_arrdiv32_mux2to1779_xor0;
  wire f_arrdiv32_mux2to1780_and0;
  wire f_arrdiv32_mux2to1780_not0;
  wire f_arrdiv32_mux2to1780_and1;
  wire f_arrdiv32_mux2to1780_xor0;
  wire f_arrdiv32_mux2to1781_and0;
  wire f_arrdiv32_mux2to1781_not0;
  wire f_arrdiv32_mux2to1781_and1;
  wire f_arrdiv32_mux2to1781_xor0;
  wire f_arrdiv32_mux2to1782_and0;
  wire f_arrdiv32_mux2to1782_not0;
  wire f_arrdiv32_mux2to1782_and1;
  wire f_arrdiv32_mux2to1782_xor0;
  wire f_arrdiv32_mux2to1783_and0;
  wire f_arrdiv32_mux2to1783_not0;
  wire f_arrdiv32_mux2to1783_and1;
  wire f_arrdiv32_mux2to1783_xor0;
  wire f_arrdiv32_mux2to1784_and0;
  wire f_arrdiv32_mux2to1784_not0;
  wire f_arrdiv32_mux2to1784_and1;
  wire f_arrdiv32_mux2to1784_xor0;
  wire f_arrdiv32_mux2to1785_and0;
  wire f_arrdiv32_mux2to1785_not0;
  wire f_arrdiv32_mux2to1785_and1;
  wire f_arrdiv32_mux2to1785_xor0;
  wire f_arrdiv32_mux2to1786_and0;
  wire f_arrdiv32_mux2to1786_not0;
  wire f_arrdiv32_mux2to1786_and1;
  wire f_arrdiv32_mux2to1786_xor0;
  wire f_arrdiv32_mux2to1787_and0;
  wire f_arrdiv32_mux2to1787_not0;
  wire f_arrdiv32_mux2to1787_and1;
  wire f_arrdiv32_mux2to1787_xor0;
  wire f_arrdiv32_mux2to1788_and0;
  wire f_arrdiv32_mux2to1788_not0;
  wire f_arrdiv32_mux2to1788_and1;
  wire f_arrdiv32_mux2to1788_xor0;
  wire f_arrdiv32_mux2to1789_and0;
  wire f_arrdiv32_mux2to1789_not0;
  wire f_arrdiv32_mux2to1789_and1;
  wire f_arrdiv32_mux2to1789_xor0;
  wire f_arrdiv32_mux2to1790_and0;
  wire f_arrdiv32_mux2to1790_not0;
  wire f_arrdiv32_mux2to1790_and1;
  wire f_arrdiv32_mux2to1790_xor0;
  wire f_arrdiv32_mux2to1791_and0;
  wire f_arrdiv32_mux2to1791_not0;
  wire f_arrdiv32_mux2to1791_and1;
  wire f_arrdiv32_mux2to1791_xor0;
  wire f_arrdiv32_mux2to1792_and0;
  wire f_arrdiv32_mux2to1792_not0;
  wire f_arrdiv32_mux2to1792_and1;
  wire f_arrdiv32_mux2to1792_xor0;
  wire f_arrdiv32_mux2to1793_and0;
  wire f_arrdiv32_mux2to1793_not0;
  wire f_arrdiv32_mux2to1793_and1;
  wire f_arrdiv32_mux2to1793_xor0;
  wire f_arrdiv32_mux2to1794_and0;
  wire f_arrdiv32_mux2to1794_not0;
  wire f_arrdiv32_mux2to1794_and1;
  wire f_arrdiv32_mux2to1794_xor0;
  wire f_arrdiv32_mux2to1795_and0;
  wire f_arrdiv32_mux2to1795_not0;
  wire f_arrdiv32_mux2to1795_and1;
  wire f_arrdiv32_mux2to1795_xor0;
  wire f_arrdiv32_mux2to1796_and0;
  wire f_arrdiv32_mux2to1796_not0;
  wire f_arrdiv32_mux2to1796_and1;
  wire f_arrdiv32_mux2to1796_xor0;
  wire f_arrdiv32_mux2to1797_and0;
  wire f_arrdiv32_mux2to1797_not0;
  wire f_arrdiv32_mux2to1797_and1;
  wire f_arrdiv32_mux2to1797_xor0;
  wire f_arrdiv32_mux2to1798_and0;
  wire f_arrdiv32_mux2to1798_not0;
  wire f_arrdiv32_mux2to1798_and1;
  wire f_arrdiv32_mux2to1798_xor0;
  wire f_arrdiv32_mux2to1799_and0;
  wire f_arrdiv32_mux2to1799_not0;
  wire f_arrdiv32_mux2to1799_and1;
  wire f_arrdiv32_mux2to1799_xor0;
  wire f_arrdiv32_mux2to1800_and0;
  wire f_arrdiv32_mux2to1800_not0;
  wire f_arrdiv32_mux2to1800_and1;
  wire f_arrdiv32_mux2to1800_xor0;
  wire f_arrdiv32_mux2to1801_and0;
  wire f_arrdiv32_mux2to1801_not0;
  wire f_arrdiv32_mux2to1801_and1;
  wire f_arrdiv32_mux2to1801_xor0;
  wire f_arrdiv32_mux2to1802_and0;
  wire f_arrdiv32_mux2to1802_not0;
  wire f_arrdiv32_mux2to1802_and1;
  wire f_arrdiv32_mux2to1802_xor0;
  wire f_arrdiv32_mux2to1803_and0;
  wire f_arrdiv32_mux2to1803_not0;
  wire f_arrdiv32_mux2to1803_and1;
  wire f_arrdiv32_mux2to1803_xor0;
  wire f_arrdiv32_mux2to1804_and0;
  wire f_arrdiv32_mux2to1804_not0;
  wire f_arrdiv32_mux2to1804_and1;
  wire f_arrdiv32_mux2to1804_xor0;
  wire f_arrdiv32_mux2to1805_and0;
  wire f_arrdiv32_mux2to1805_not0;
  wire f_arrdiv32_mux2to1805_and1;
  wire f_arrdiv32_mux2to1805_xor0;
  wire f_arrdiv32_not25;
  wire f_arrdiv32_fs832_xor0;
  wire f_arrdiv32_fs832_not0;
  wire f_arrdiv32_fs832_and0;
  wire f_arrdiv32_fs832_not1;
  wire f_arrdiv32_fs833_xor0;
  wire f_arrdiv32_fs833_not0;
  wire f_arrdiv32_fs833_and0;
  wire f_arrdiv32_fs833_xor1;
  wire f_arrdiv32_fs833_not1;
  wire f_arrdiv32_fs833_and1;
  wire f_arrdiv32_fs833_or0;
  wire f_arrdiv32_fs834_xor0;
  wire f_arrdiv32_fs834_not0;
  wire f_arrdiv32_fs834_and0;
  wire f_arrdiv32_fs834_xor1;
  wire f_arrdiv32_fs834_not1;
  wire f_arrdiv32_fs834_and1;
  wire f_arrdiv32_fs834_or0;
  wire f_arrdiv32_fs835_xor0;
  wire f_arrdiv32_fs835_not0;
  wire f_arrdiv32_fs835_and0;
  wire f_arrdiv32_fs835_xor1;
  wire f_arrdiv32_fs835_not1;
  wire f_arrdiv32_fs835_and1;
  wire f_arrdiv32_fs835_or0;
  wire f_arrdiv32_fs836_xor0;
  wire f_arrdiv32_fs836_not0;
  wire f_arrdiv32_fs836_and0;
  wire f_arrdiv32_fs836_xor1;
  wire f_arrdiv32_fs836_not1;
  wire f_arrdiv32_fs836_and1;
  wire f_arrdiv32_fs836_or0;
  wire f_arrdiv32_fs837_xor0;
  wire f_arrdiv32_fs837_not0;
  wire f_arrdiv32_fs837_and0;
  wire f_arrdiv32_fs837_xor1;
  wire f_arrdiv32_fs837_not1;
  wire f_arrdiv32_fs837_and1;
  wire f_arrdiv32_fs837_or0;
  wire f_arrdiv32_fs838_xor0;
  wire f_arrdiv32_fs838_not0;
  wire f_arrdiv32_fs838_and0;
  wire f_arrdiv32_fs838_xor1;
  wire f_arrdiv32_fs838_not1;
  wire f_arrdiv32_fs838_and1;
  wire f_arrdiv32_fs838_or0;
  wire f_arrdiv32_fs839_xor0;
  wire f_arrdiv32_fs839_not0;
  wire f_arrdiv32_fs839_and0;
  wire f_arrdiv32_fs839_xor1;
  wire f_arrdiv32_fs839_not1;
  wire f_arrdiv32_fs839_and1;
  wire f_arrdiv32_fs839_or0;
  wire f_arrdiv32_fs840_xor0;
  wire f_arrdiv32_fs840_not0;
  wire f_arrdiv32_fs840_and0;
  wire f_arrdiv32_fs840_xor1;
  wire f_arrdiv32_fs840_not1;
  wire f_arrdiv32_fs840_and1;
  wire f_arrdiv32_fs840_or0;
  wire f_arrdiv32_fs841_xor0;
  wire f_arrdiv32_fs841_not0;
  wire f_arrdiv32_fs841_and0;
  wire f_arrdiv32_fs841_xor1;
  wire f_arrdiv32_fs841_not1;
  wire f_arrdiv32_fs841_and1;
  wire f_arrdiv32_fs841_or0;
  wire f_arrdiv32_fs842_xor0;
  wire f_arrdiv32_fs842_not0;
  wire f_arrdiv32_fs842_and0;
  wire f_arrdiv32_fs842_xor1;
  wire f_arrdiv32_fs842_not1;
  wire f_arrdiv32_fs842_and1;
  wire f_arrdiv32_fs842_or0;
  wire f_arrdiv32_fs843_xor0;
  wire f_arrdiv32_fs843_not0;
  wire f_arrdiv32_fs843_and0;
  wire f_arrdiv32_fs843_xor1;
  wire f_arrdiv32_fs843_not1;
  wire f_arrdiv32_fs843_and1;
  wire f_arrdiv32_fs843_or0;
  wire f_arrdiv32_fs844_xor0;
  wire f_arrdiv32_fs844_not0;
  wire f_arrdiv32_fs844_and0;
  wire f_arrdiv32_fs844_xor1;
  wire f_arrdiv32_fs844_not1;
  wire f_arrdiv32_fs844_and1;
  wire f_arrdiv32_fs844_or0;
  wire f_arrdiv32_fs845_xor0;
  wire f_arrdiv32_fs845_not0;
  wire f_arrdiv32_fs845_and0;
  wire f_arrdiv32_fs845_xor1;
  wire f_arrdiv32_fs845_not1;
  wire f_arrdiv32_fs845_and1;
  wire f_arrdiv32_fs845_or0;
  wire f_arrdiv32_fs846_xor0;
  wire f_arrdiv32_fs846_not0;
  wire f_arrdiv32_fs846_and0;
  wire f_arrdiv32_fs846_xor1;
  wire f_arrdiv32_fs846_not1;
  wire f_arrdiv32_fs846_and1;
  wire f_arrdiv32_fs846_or0;
  wire f_arrdiv32_fs847_xor0;
  wire f_arrdiv32_fs847_not0;
  wire f_arrdiv32_fs847_and0;
  wire f_arrdiv32_fs847_xor1;
  wire f_arrdiv32_fs847_not1;
  wire f_arrdiv32_fs847_and1;
  wire f_arrdiv32_fs847_or0;
  wire f_arrdiv32_fs848_xor0;
  wire f_arrdiv32_fs848_not0;
  wire f_arrdiv32_fs848_and0;
  wire f_arrdiv32_fs848_xor1;
  wire f_arrdiv32_fs848_not1;
  wire f_arrdiv32_fs848_and1;
  wire f_arrdiv32_fs848_or0;
  wire f_arrdiv32_fs849_xor0;
  wire f_arrdiv32_fs849_not0;
  wire f_arrdiv32_fs849_and0;
  wire f_arrdiv32_fs849_xor1;
  wire f_arrdiv32_fs849_not1;
  wire f_arrdiv32_fs849_and1;
  wire f_arrdiv32_fs849_or0;
  wire f_arrdiv32_fs850_xor0;
  wire f_arrdiv32_fs850_not0;
  wire f_arrdiv32_fs850_and0;
  wire f_arrdiv32_fs850_xor1;
  wire f_arrdiv32_fs850_not1;
  wire f_arrdiv32_fs850_and1;
  wire f_arrdiv32_fs850_or0;
  wire f_arrdiv32_fs851_xor0;
  wire f_arrdiv32_fs851_not0;
  wire f_arrdiv32_fs851_and0;
  wire f_arrdiv32_fs851_xor1;
  wire f_arrdiv32_fs851_not1;
  wire f_arrdiv32_fs851_and1;
  wire f_arrdiv32_fs851_or0;
  wire f_arrdiv32_fs852_xor0;
  wire f_arrdiv32_fs852_not0;
  wire f_arrdiv32_fs852_and0;
  wire f_arrdiv32_fs852_xor1;
  wire f_arrdiv32_fs852_not1;
  wire f_arrdiv32_fs852_and1;
  wire f_arrdiv32_fs852_or0;
  wire f_arrdiv32_fs853_xor0;
  wire f_arrdiv32_fs853_not0;
  wire f_arrdiv32_fs853_and0;
  wire f_arrdiv32_fs853_xor1;
  wire f_arrdiv32_fs853_not1;
  wire f_arrdiv32_fs853_and1;
  wire f_arrdiv32_fs853_or0;
  wire f_arrdiv32_fs854_xor0;
  wire f_arrdiv32_fs854_not0;
  wire f_arrdiv32_fs854_and0;
  wire f_arrdiv32_fs854_xor1;
  wire f_arrdiv32_fs854_not1;
  wire f_arrdiv32_fs854_and1;
  wire f_arrdiv32_fs854_or0;
  wire f_arrdiv32_fs855_xor0;
  wire f_arrdiv32_fs855_not0;
  wire f_arrdiv32_fs855_and0;
  wire f_arrdiv32_fs855_xor1;
  wire f_arrdiv32_fs855_not1;
  wire f_arrdiv32_fs855_and1;
  wire f_arrdiv32_fs855_or0;
  wire f_arrdiv32_fs856_xor0;
  wire f_arrdiv32_fs856_not0;
  wire f_arrdiv32_fs856_and0;
  wire f_arrdiv32_fs856_xor1;
  wire f_arrdiv32_fs856_not1;
  wire f_arrdiv32_fs856_and1;
  wire f_arrdiv32_fs856_or0;
  wire f_arrdiv32_fs857_xor0;
  wire f_arrdiv32_fs857_not0;
  wire f_arrdiv32_fs857_and0;
  wire f_arrdiv32_fs857_xor1;
  wire f_arrdiv32_fs857_not1;
  wire f_arrdiv32_fs857_and1;
  wire f_arrdiv32_fs857_or0;
  wire f_arrdiv32_fs858_xor0;
  wire f_arrdiv32_fs858_not0;
  wire f_arrdiv32_fs858_and0;
  wire f_arrdiv32_fs858_xor1;
  wire f_arrdiv32_fs858_not1;
  wire f_arrdiv32_fs858_and1;
  wire f_arrdiv32_fs858_or0;
  wire f_arrdiv32_fs859_xor0;
  wire f_arrdiv32_fs859_not0;
  wire f_arrdiv32_fs859_and0;
  wire f_arrdiv32_fs859_xor1;
  wire f_arrdiv32_fs859_not1;
  wire f_arrdiv32_fs859_and1;
  wire f_arrdiv32_fs859_or0;
  wire f_arrdiv32_fs860_xor0;
  wire f_arrdiv32_fs860_not0;
  wire f_arrdiv32_fs860_and0;
  wire f_arrdiv32_fs860_xor1;
  wire f_arrdiv32_fs860_not1;
  wire f_arrdiv32_fs860_and1;
  wire f_arrdiv32_fs860_or0;
  wire f_arrdiv32_fs861_xor0;
  wire f_arrdiv32_fs861_not0;
  wire f_arrdiv32_fs861_and0;
  wire f_arrdiv32_fs861_xor1;
  wire f_arrdiv32_fs861_not1;
  wire f_arrdiv32_fs861_and1;
  wire f_arrdiv32_fs861_or0;
  wire f_arrdiv32_fs862_xor0;
  wire f_arrdiv32_fs862_not0;
  wire f_arrdiv32_fs862_and0;
  wire f_arrdiv32_fs862_xor1;
  wire f_arrdiv32_fs862_not1;
  wire f_arrdiv32_fs862_and1;
  wire f_arrdiv32_fs862_or0;
  wire f_arrdiv32_fs863_xor0;
  wire f_arrdiv32_fs863_not0;
  wire f_arrdiv32_fs863_and0;
  wire f_arrdiv32_fs863_xor1;
  wire f_arrdiv32_fs863_not1;
  wire f_arrdiv32_fs863_and1;
  wire f_arrdiv32_fs863_or0;
  wire f_arrdiv32_mux2to1806_and0;
  wire f_arrdiv32_mux2to1806_not0;
  wire f_arrdiv32_mux2to1806_and1;
  wire f_arrdiv32_mux2to1806_xor0;
  wire f_arrdiv32_mux2to1807_and0;
  wire f_arrdiv32_mux2to1807_not0;
  wire f_arrdiv32_mux2to1807_and1;
  wire f_arrdiv32_mux2to1807_xor0;
  wire f_arrdiv32_mux2to1808_and0;
  wire f_arrdiv32_mux2to1808_not0;
  wire f_arrdiv32_mux2to1808_and1;
  wire f_arrdiv32_mux2to1808_xor0;
  wire f_arrdiv32_mux2to1809_and0;
  wire f_arrdiv32_mux2to1809_not0;
  wire f_arrdiv32_mux2to1809_and1;
  wire f_arrdiv32_mux2to1809_xor0;
  wire f_arrdiv32_mux2to1810_and0;
  wire f_arrdiv32_mux2to1810_not0;
  wire f_arrdiv32_mux2to1810_and1;
  wire f_arrdiv32_mux2to1810_xor0;
  wire f_arrdiv32_mux2to1811_and0;
  wire f_arrdiv32_mux2to1811_not0;
  wire f_arrdiv32_mux2to1811_and1;
  wire f_arrdiv32_mux2to1811_xor0;
  wire f_arrdiv32_mux2to1812_and0;
  wire f_arrdiv32_mux2to1812_not0;
  wire f_arrdiv32_mux2to1812_and1;
  wire f_arrdiv32_mux2to1812_xor0;
  wire f_arrdiv32_mux2to1813_and0;
  wire f_arrdiv32_mux2to1813_not0;
  wire f_arrdiv32_mux2to1813_and1;
  wire f_arrdiv32_mux2to1813_xor0;
  wire f_arrdiv32_mux2to1814_and0;
  wire f_arrdiv32_mux2to1814_not0;
  wire f_arrdiv32_mux2to1814_and1;
  wire f_arrdiv32_mux2to1814_xor0;
  wire f_arrdiv32_mux2to1815_and0;
  wire f_arrdiv32_mux2to1815_not0;
  wire f_arrdiv32_mux2to1815_and1;
  wire f_arrdiv32_mux2to1815_xor0;
  wire f_arrdiv32_mux2to1816_and0;
  wire f_arrdiv32_mux2to1816_not0;
  wire f_arrdiv32_mux2to1816_and1;
  wire f_arrdiv32_mux2to1816_xor0;
  wire f_arrdiv32_mux2to1817_and0;
  wire f_arrdiv32_mux2to1817_not0;
  wire f_arrdiv32_mux2to1817_and1;
  wire f_arrdiv32_mux2to1817_xor0;
  wire f_arrdiv32_mux2to1818_and0;
  wire f_arrdiv32_mux2to1818_not0;
  wire f_arrdiv32_mux2to1818_and1;
  wire f_arrdiv32_mux2to1818_xor0;
  wire f_arrdiv32_mux2to1819_and0;
  wire f_arrdiv32_mux2to1819_not0;
  wire f_arrdiv32_mux2to1819_and1;
  wire f_arrdiv32_mux2to1819_xor0;
  wire f_arrdiv32_mux2to1820_and0;
  wire f_arrdiv32_mux2to1820_not0;
  wire f_arrdiv32_mux2to1820_and1;
  wire f_arrdiv32_mux2to1820_xor0;
  wire f_arrdiv32_mux2to1821_and0;
  wire f_arrdiv32_mux2to1821_not0;
  wire f_arrdiv32_mux2to1821_and1;
  wire f_arrdiv32_mux2to1821_xor0;
  wire f_arrdiv32_mux2to1822_and0;
  wire f_arrdiv32_mux2to1822_not0;
  wire f_arrdiv32_mux2to1822_and1;
  wire f_arrdiv32_mux2to1822_xor0;
  wire f_arrdiv32_mux2to1823_and0;
  wire f_arrdiv32_mux2to1823_not0;
  wire f_arrdiv32_mux2to1823_and1;
  wire f_arrdiv32_mux2to1823_xor0;
  wire f_arrdiv32_mux2to1824_and0;
  wire f_arrdiv32_mux2to1824_not0;
  wire f_arrdiv32_mux2to1824_and1;
  wire f_arrdiv32_mux2to1824_xor0;
  wire f_arrdiv32_mux2to1825_and0;
  wire f_arrdiv32_mux2to1825_not0;
  wire f_arrdiv32_mux2to1825_and1;
  wire f_arrdiv32_mux2to1825_xor0;
  wire f_arrdiv32_mux2to1826_and0;
  wire f_arrdiv32_mux2to1826_not0;
  wire f_arrdiv32_mux2to1826_and1;
  wire f_arrdiv32_mux2to1826_xor0;
  wire f_arrdiv32_mux2to1827_and0;
  wire f_arrdiv32_mux2to1827_not0;
  wire f_arrdiv32_mux2to1827_and1;
  wire f_arrdiv32_mux2to1827_xor0;
  wire f_arrdiv32_mux2to1828_and0;
  wire f_arrdiv32_mux2to1828_not0;
  wire f_arrdiv32_mux2to1828_and1;
  wire f_arrdiv32_mux2to1828_xor0;
  wire f_arrdiv32_mux2to1829_and0;
  wire f_arrdiv32_mux2to1829_not0;
  wire f_arrdiv32_mux2to1829_and1;
  wire f_arrdiv32_mux2to1829_xor0;
  wire f_arrdiv32_mux2to1830_and0;
  wire f_arrdiv32_mux2to1830_not0;
  wire f_arrdiv32_mux2to1830_and1;
  wire f_arrdiv32_mux2to1830_xor0;
  wire f_arrdiv32_mux2to1831_and0;
  wire f_arrdiv32_mux2to1831_not0;
  wire f_arrdiv32_mux2to1831_and1;
  wire f_arrdiv32_mux2to1831_xor0;
  wire f_arrdiv32_mux2to1832_and0;
  wire f_arrdiv32_mux2to1832_not0;
  wire f_arrdiv32_mux2to1832_and1;
  wire f_arrdiv32_mux2to1832_xor0;
  wire f_arrdiv32_mux2to1833_and0;
  wire f_arrdiv32_mux2to1833_not0;
  wire f_arrdiv32_mux2to1833_and1;
  wire f_arrdiv32_mux2to1833_xor0;
  wire f_arrdiv32_mux2to1834_and0;
  wire f_arrdiv32_mux2to1834_not0;
  wire f_arrdiv32_mux2to1834_and1;
  wire f_arrdiv32_mux2to1834_xor0;
  wire f_arrdiv32_mux2to1835_and0;
  wire f_arrdiv32_mux2to1835_not0;
  wire f_arrdiv32_mux2to1835_and1;
  wire f_arrdiv32_mux2to1835_xor0;
  wire f_arrdiv32_mux2to1836_and0;
  wire f_arrdiv32_mux2to1836_not0;
  wire f_arrdiv32_mux2to1836_and1;
  wire f_arrdiv32_mux2to1836_xor0;
  wire f_arrdiv32_not26;
  wire f_arrdiv32_fs864_xor0;
  wire f_arrdiv32_fs864_not0;
  wire f_arrdiv32_fs864_and0;
  wire f_arrdiv32_fs864_not1;
  wire f_arrdiv32_fs865_xor0;
  wire f_arrdiv32_fs865_not0;
  wire f_arrdiv32_fs865_and0;
  wire f_arrdiv32_fs865_xor1;
  wire f_arrdiv32_fs865_not1;
  wire f_arrdiv32_fs865_and1;
  wire f_arrdiv32_fs865_or0;
  wire f_arrdiv32_fs866_xor0;
  wire f_arrdiv32_fs866_not0;
  wire f_arrdiv32_fs866_and0;
  wire f_arrdiv32_fs866_xor1;
  wire f_arrdiv32_fs866_not1;
  wire f_arrdiv32_fs866_and1;
  wire f_arrdiv32_fs866_or0;
  wire f_arrdiv32_fs867_xor0;
  wire f_arrdiv32_fs867_not0;
  wire f_arrdiv32_fs867_and0;
  wire f_arrdiv32_fs867_xor1;
  wire f_arrdiv32_fs867_not1;
  wire f_arrdiv32_fs867_and1;
  wire f_arrdiv32_fs867_or0;
  wire f_arrdiv32_fs868_xor0;
  wire f_arrdiv32_fs868_not0;
  wire f_arrdiv32_fs868_and0;
  wire f_arrdiv32_fs868_xor1;
  wire f_arrdiv32_fs868_not1;
  wire f_arrdiv32_fs868_and1;
  wire f_arrdiv32_fs868_or0;
  wire f_arrdiv32_fs869_xor0;
  wire f_arrdiv32_fs869_not0;
  wire f_arrdiv32_fs869_and0;
  wire f_arrdiv32_fs869_xor1;
  wire f_arrdiv32_fs869_not1;
  wire f_arrdiv32_fs869_and1;
  wire f_arrdiv32_fs869_or0;
  wire f_arrdiv32_fs870_xor0;
  wire f_arrdiv32_fs870_not0;
  wire f_arrdiv32_fs870_and0;
  wire f_arrdiv32_fs870_xor1;
  wire f_arrdiv32_fs870_not1;
  wire f_arrdiv32_fs870_and1;
  wire f_arrdiv32_fs870_or0;
  wire f_arrdiv32_fs871_xor0;
  wire f_arrdiv32_fs871_not0;
  wire f_arrdiv32_fs871_and0;
  wire f_arrdiv32_fs871_xor1;
  wire f_arrdiv32_fs871_not1;
  wire f_arrdiv32_fs871_and1;
  wire f_arrdiv32_fs871_or0;
  wire f_arrdiv32_fs872_xor0;
  wire f_arrdiv32_fs872_not0;
  wire f_arrdiv32_fs872_and0;
  wire f_arrdiv32_fs872_xor1;
  wire f_arrdiv32_fs872_not1;
  wire f_arrdiv32_fs872_and1;
  wire f_arrdiv32_fs872_or0;
  wire f_arrdiv32_fs873_xor0;
  wire f_arrdiv32_fs873_not0;
  wire f_arrdiv32_fs873_and0;
  wire f_arrdiv32_fs873_xor1;
  wire f_arrdiv32_fs873_not1;
  wire f_arrdiv32_fs873_and1;
  wire f_arrdiv32_fs873_or0;
  wire f_arrdiv32_fs874_xor0;
  wire f_arrdiv32_fs874_not0;
  wire f_arrdiv32_fs874_and0;
  wire f_arrdiv32_fs874_xor1;
  wire f_arrdiv32_fs874_not1;
  wire f_arrdiv32_fs874_and1;
  wire f_arrdiv32_fs874_or0;
  wire f_arrdiv32_fs875_xor0;
  wire f_arrdiv32_fs875_not0;
  wire f_arrdiv32_fs875_and0;
  wire f_arrdiv32_fs875_xor1;
  wire f_arrdiv32_fs875_not1;
  wire f_arrdiv32_fs875_and1;
  wire f_arrdiv32_fs875_or0;
  wire f_arrdiv32_fs876_xor0;
  wire f_arrdiv32_fs876_not0;
  wire f_arrdiv32_fs876_and0;
  wire f_arrdiv32_fs876_xor1;
  wire f_arrdiv32_fs876_not1;
  wire f_arrdiv32_fs876_and1;
  wire f_arrdiv32_fs876_or0;
  wire f_arrdiv32_fs877_xor0;
  wire f_arrdiv32_fs877_not0;
  wire f_arrdiv32_fs877_and0;
  wire f_arrdiv32_fs877_xor1;
  wire f_arrdiv32_fs877_not1;
  wire f_arrdiv32_fs877_and1;
  wire f_arrdiv32_fs877_or0;
  wire f_arrdiv32_fs878_xor0;
  wire f_arrdiv32_fs878_not0;
  wire f_arrdiv32_fs878_and0;
  wire f_arrdiv32_fs878_xor1;
  wire f_arrdiv32_fs878_not1;
  wire f_arrdiv32_fs878_and1;
  wire f_arrdiv32_fs878_or0;
  wire f_arrdiv32_fs879_xor0;
  wire f_arrdiv32_fs879_not0;
  wire f_arrdiv32_fs879_and0;
  wire f_arrdiv32_fs879_xor1;
  wire f_arrdiv32_fs879_not1;
  wire f_arrdiv32_fs879_and1;
  wire f_arrdiv32_fs879_or0;
  wire f_arrdiv32_fs880_xor0;
  wire f_arrdiv32_fs880_not0;
  wire f_arrdiv32_fs880_and0;
  wire f_arrdiv32_fs880_xor1;
  wire f_arrdiv32_fs880_not1;
  wire f_arrdiv32_fs880_and1;
  wire f_arrdiv32_fs880_or0;
  wire f_arrdiv32_fs881_xor0;
  wire f_arrdiv32_fs881_not0;
  wire f_arrdiv32_fs881_and0;
  wire f_arrdiv32_fs881_xor1;
  wire f_arrdiv32_fs881_not1;
  wire f_arrdiv32_fs881_and1;
  wire f_arrdiv32_fs881_or0;
  wire f_arrdiv32_fs882_xor0;
  wire f_arrdiv32_fs882_not0;
  wire f_arrdiv32_fs882_and0;
  wire f_arrdiv32_fs882_xor1;
  wire f_arrdiv32_fs882_not1;
  wire f_arrdiv32_fs882_and1;
  wire f_arrdiv32_fs882_or0;
  wire f_arrdiv32_fs883_xor0;
  wire f_arrdiv32_fs883_not0;
  wire f_arrdiv32_fs883_and0;
  wire f_arrdiv32_fs883_xor1;
  wire f_arrdiv32_fs883_not1;
  wire f_arrdiv32_fs883_and1;
  wire f_arrdiv32_fs883_or0;
  wire f_arrdiv32_fs884_xor0;
  wire f_arrdiv32_fs884_not0;
  wire f_arrdiv32_fs884_and0;
  wire f_arrdiv32_fs884_xor1;
  wire f_arrdiv32_fs884_not1;
  wire f_arrdiv32_fs884_and1;
  wire f_arrdiv32_fs884_or0;
  wire f_arrdiv32_fs885_xor0;
  wire f_arrdiv32_fs885_not0;
  wire f_arrdiv32_fs885_and0;
  wire f_arrdiv32_fs885_xor1;
  wire f_arrdiv32_fs885_not1;
  wire f_arrdiv32_fs885_and1;
  wire f_arrdiv32_fs885_or0;
  wire f_arrdiv32_fs886_xor0;
  wire f_arrdiv32_fs886_not0;
  wire f_arrdiv32_fs886_and0;
  wire f_arrdiv32_fs886_xor1;
  wire f_arrdiv32_fs886_not1;
  wire f_arrdiv32_fs886_and1;
  wire f_arrdiv32_fs886_or0;
  wire f_arrdiv32_fs887_xor0;
  wire f_arrdiv32_fs887_not0;
  wire f_arrdiv32_fs887_and0;
  wire f_arrdiv32_fs887_xor1;
  wire f_arrdiv32_fs887_not1;
  wire f_arrdiv32_fs887_and1;
  wire f_arrdiv32_fs887_or0;
  wire f_arrdiv32_fs888_xor0;
  wire f_arrdiv32_fs888_not0;
  wire f_arrdiv32_fs888_and0;
  wire f_arrdiv32_fs888_xor1;
  wire f_arrdiv32_fs888_not1;
  wire f_arrdiv32_fs888_and1;
  wire f_arrdiv32_fs888_or0;
  wire f_arrdiv32_fs889_xor0;
  wire f_arrdiv32_fs889_not0;
  wire f_arrdiv32_fs889_and0;
  wire f_arrdiv32_fs889_xor1;
  wire f_arrdiv32_fs889_not1;
  wire f_arrdiv32_fs889_and1;
  wire f_arrdiv32_fs889_or0;
  wire f_arrdiv32_fs890_xor0;
  wire f_arrdiv32_fs890_not0;
  wire f_arrdiv32_fs890_and0;
  wire f_arrdiv32_fs890_xor1;
  wire f_arrdiv32_fs890_not1;
  wire f_arrdiv32_fs890_and1;
  wire f_arrdiv32_fs890_or0;
  wire f_arrdiv32_fs891_xor0;
  wire f_arrdiv32_fs891_not0;
  wire f_arrdiv32_fs891_and0;
  wire f_arrdiv32_fs891_xor1;
  wire f_arrdiv32_fs891_not1;
  wire f_arrdiv32_fs891_and1;
  wire f_arrdiv32_fs891_or0;
  wire f_arrdiv32_fs892_xor0;
  wire f_arrdiv32_fs892_not0;
  wire f_arrdiv32_fs892_and0;
  wire f_arrdiv32_fs892_xor1;
  wire f_arrdiv32_fs892_not1;
  wire f_arrdiv32_fs892_and1;
  wire f_arrdiv32_fs892_or0;
  wire f_arrdiv32_fs893_xor0;
  wire f_arrdiv32_fs893_not0;
  wire f_arrdiv32_fs893_and0;
  wire f_arrdiv32_fs893_xor1;
  wire f_arrdiv32_fs893_not1;
  wire f_arrdiv32_fs893_and1;
  wire f_arrdiv32_fs893_or0;
  wire f_arrdiv32_fs894_xor0;
  wire f_arrdiv32_fs894_not0;
  wire f_arrdiv32_fs894_and0;
  wire f_arrdiv32_fs894_xor1;
  wire f_arrdiv32_fs894_not1;
  wire f_arrdiv32_fs894_and1;
  wire f_arrdiv32_fs894_or0;
  wire f_arrdiv32_fs895_xor0;
  wire f_arrdiv32_fs895_not0;
  wire f_arrdiv32_fs895_and0;
  wire f_arrdiv32_fs895_xor1;
  wire f_arrdiv32_fs895_not1;
  wire f_arrdiv32_fs895_and1;
  wire f_arrdiv32_fs895_or0;
  wire f_arrdiv32_mux2to1837_and0;
  wire f_arrdiv32_mux2to1837_not0;
  wire f_arrdiv32_mux2to1837_and1;
  wire f_arrdiv32_mux2to1837_xor0;
  wire f_arrdiv32_mux2to1838_and0;
  wire f_arrdiv32_mux2to1838_not0;
  wire f_arrdiv32_mux2to1838_and1;
  wire f_arrdiv32_mux2to1838_xor0;
  wire f_arrdiv32_mux2to1839_and0;
  wire f_arrdiv32_mux2to1839_not0;
  wire f_arrdiv32_mux2to1839_and1;
  wire f_arrdiv32_mux2to1839_xor0;
  wire f_arrdiv32_mux2to1840_and0;
  wire f_arrdiv32_mux2to1840_not0;
  wire f_arrdiv32_mux2to1840_and1;
  wire f_arrdiv32_mux2to1840_xor0;
  wire f_arrdiv32_mux2to1841_and0;
  wire f_arrdiv32_mux2to1841_not0;
  wire f_arrdiv32_mux2to1841_and1;
  wire f_arrdiv32_mux2to1841_xor0;
  wire f_arrdiv32_mux2to1842_and0;
  wire f_arrdiv32_mux2to1842_not0;
  wire f_arrdiv32_mux2to1842_and1;
  wire f_arrdiv32_mux2to1842_xor0;
  wire f_arrdiv32_mux2to1843_and0;
  wire f_arrdiv32_mux2to1843_not0;
  wire f_arrdiv32_mux2to1843_and1;
  wire f_arrdiv32_mux2to1843_xor0;
  wire f_arrdiv32_mux2to1844_and0;
  wire f_arrdiv32_mux2to1844_not0;
  wire f_arrdiv32_mux2to1844_and1;
  wire f_arrdiv32_mux2to1844_xor0;
  wire f_arrdiv32_mux2to1845_and0;
  wire f_arrdiv32_mux2to1845_not0;
  wire f_arrdiv32_mux2to1845_and1;
  wire f_arrdiv32_mux2to1845_xor0;
  wire f_arrdiv32_mux2to1846_and0;
  wire f_arrdiv32_mux2to1846_not0;
  wire f_arrdiv32_mux2to1846_and1;
  wire f_arrdiv32_mux2to1846_xor0;
  wire f_arrdiv32_mux2to1847_and0;
  wire f_arrdiv32_mux2to1847_not0;
  wire f_arrdiv32_mux2to1847_and1;
  wire f_arrdiv32_mux2to1847_xor0;
  wire f_arrdiv32_mux2to1848_and0;
  wire f_arrdiv32_mux2to1848_not0;
  wire f_arrdiv32_mux2to1848_and1;
  wire f_arrdiv32_mux2to1848_xor0;
  wire f_arrdiv32_mux2to1849_and0;
  wire f_arrdiv32_mux2to1849_not0;
  wire f_arrdiv32_mux2to1849_and1;
  wire f_arrdiv32_mux2to1849_xor0;
  wire f_arrdiv32_mux2to1850_and0;
  wire f_arrdiv32_mux2to1850_not0;
  wire f_arrdiv32_mux2to1850_and1;
  wire f_arrdiv32_mux2to1850_xor0;
  wire f_arrdiv32_mux2to1851_and0;
  wire f_arrdiv32_mux2to1851_not0;
  wire f_arrdiv32_mux2to1851_and1;
  wire f_arrdiv32_mux2to1851_xor0;
  wire f_arrdiv32_mux2to1852_and0;
  wire f_arrdiv32_mux2to1852_not0;
  wire f_arrdiv32_mux2to1852_and1;
  wire f_arrdiv32_mux2to1852_xor0;
  wire f_arrdiv32_mux2to1853_and0;
  wire f_arrdiv32_mux2to1853_not0;
  wire f_arrdiv32_mux2to1853_and1;
  wire f_arrdiv32_mux2to1853_xor0;
  wire f_arrdiv32_mux2to1854_and0;
  wire f_arrdiv32_mux2to1854_not0;
  wire f_arrdiv32_mux2to1854_and1;
  wire f_arrdiv32_mux2to1854_xor0;
  wire f_arrdiv32_mux2to1855_and0;
  wire f_arrdiv32_mux2to1855_not0;
  wire f_arrdiv32_mux2to1855_and1;
  wire f_arrdiv32_mux2to1855_xor0;
  wire f_arrdiv32_mux2to1856_and0;
  wire f_arrdiv32_mux2to1856_not0;
  wire f_arrdiv32_mux2to1856_and1;
  wire f_arrdiv32_mux2to1856_xor0;
  wire f_arrdiv32_mux2to1857_and0;
  wire f_arrdiv32_mux2to1857_not0;
  wire f_arrdiv32_mux2to1857_and1;
  wire f_arrdiv32_mux2to1857_xor0;
  wire f_arrdiv32_mux2to1858_and0;
  wire f_arrdiv32_mux2to1858_not0;
  wire f_arrdiv32_mux2to1858_and1;
  wire f_arrdiv32_mux2to1858_xor0;
  wire f_arrdiv32_mux2to1859_and0;
  wire f_arrdiv32_mux2to1859_not0;
  wire f_arrdiv32_mux2to1859_and1;
  wire f_arrdiv32_mux2to1859_xor0;
  wire f_arrdiv32_mux2to1860_and0;
  wire f_arrdiv32_mux2to1860_not0;
  wire f_arrdiv32_mux2to1860_and1;
  wire f_arrdiv32_mux2to1860_xor0;
  wire f_arrdiv32_mux2to1861_and0;
  wire f_arrdiv32_mux2to1861_not0;
  wire f_arrdiv32_mux2to1861_and1;
  wire f_arrdiv32_mux2to1861_xor0;
  wire f_arrdiv32_mux2to1862_and0;
  wire f_arrdiv32_mux2to1862_not0;
  wire f_arrdiv32_mux2to1862_and1;
  wire f_arrdiv32_mux2to1862_xor0;
  wire f_arrdiv32_mux2to1863_and0;
  wire f_arrdiv32_mux2to1863_not0;
  wire f_arrdiv32_mux2to1863_and1;
  wire f_arrdiv32_mux2to1863_xor0;
  wire f_arrdiv32_mux2to1864_and0;
  wire f_arrdiv32_mux2to1864_not0;
  wire f_arrdiv32_mux2to1864_and1;
  wire f_arrdiv32_mux2to1864_xor0;
  wire f_arrdiv32_mux2to1865_and0;
  wire f_arrdiv32_mux2to1865_not0;
  wire f_arrdiv32_mux2to1865_and1;
  wire f_arrdiv32_mux2to1865_xor0;
  wire f_arrdiv32_mux2to1866_and0;
  wire f_arrdiv32_mux2to1866_not0;
  wire f_arrdiv32_mux2to1866_and1;
  wire f_arrdiv32_mux2to1866_xor0;
  wire f_arrdiv32_mux2to1867_and0;
  wire f_arrdiv32_mux2to1867_not0;
  wire f_arrdiv32_mux2to1867_and1;
  wire f_arrdiv32_mux2to1867_xor0;
  wire f_arrdiv32_not27;
  wire f_arrdiv32_fs896_xor0;
  wire f_arrdiv32_fs896_not0;
  wire f_arrdiv32_fs896_and0;
  wire f_arrdiv32_fs896_not1;
  wire f_arrdiv32_fs897_xor0;
  wire f_arrdiv32_fs897_not0;
  wire f_arrdiv32_fs897_and0;
  wire f_arrdiv32_fs897_xor1;
  wire f_arrdiv32_fs897_not1;
  wire f_arrdiv32_fs897_and1;
  wire f_arrdiv32_fs897_or0;
  wire f_arrdiv32_fs898_xor0;
  wire f_arrdiv32_fs898_not0;
  wire f_arrdiv32_fs898_and0;
  wire f_arrdiv32_fs898_xor1;
  wire f_arrdiv32_fs898_not1;
  wire f_arrdiv32_fs898_and1;
  wire f_arrdiv32_fs898_or0;
  wire f_arrdiv32_fs899_xor0;
  wire f_arrdiv32_fs899_not0;
  wire f_arrdiv32_fs899_and0;
  wire f_arrdiv32_fs899_xor1;
  wire f_arrdiv32_fs899_not1;
  wire f_arrdiv32_fs899_and1;
  wire f_arrdiv32_fs899_or0;
  wire f_arrdiv32_fs900_xor0;
  wire f_arrdiv32_fs900_not0;
  wire f_arrdiv32_fs900_and0;
  wire f_arrdiv32_fs900_xor1;
  wire f_arrdiv32_fs900_not1;
  wire f_arrdiv32_fs900_and1;
  wire f_arrdiv32_fs900_or0;
  wire f_arrdiv32_fs901_xor0;
  wire f_arrdiv32_fs901_not0;
  wire f_arrdiv32_fs901_and0;
  wire f_arrdiv32_fs901_xor1;
  wire f_arrdiv32_fs901_not1;
  wire f_arrdiv32_fs901_and1;
  wire f_arrdiv32_fs901_or0;
  wire f_arrdiv32_fs902_xor0;
  wire f_arrdiv32_fs902_not0;
  wire f_arrdiv32_fs902_and0;
  wire f_arrdiv32_fs902_xor1;
  wire f_arrdiv32_fs902_not1;
  wire f_arrdiv32_fs902_and1;
  wire f_arrdiv32_fs902_or0;
  wire f_arrdiv32_fs903_xor0;
  wire f_arrdiv32_fs903_not0;
  wire f_arrdiv32_fs903_and0;
  wire f_arrdiv32_fs903_xor1;
  wire f_arrdiv32_fs903_not1;
  wire f_arrdiv32_fs903_and1;
  wire f_arrdiv32_fs903_or0;
  wire f_arrdiv32_fs904_xor0;
  wire f_arrdiv32_fs904_not0;
  wire f_arrdiv32_fs904_and0;
  wire f_arrdiv32_fs904_xor1;
  wire f_arrdiv32_fs904_not1;
  wire f_arrdiv32_fs904_and1;
  wire f_arrdiv32_fs904_or0;
  wire f_arrdiv32_fs905_xor0;
  wire f_arrdiv32_fs905_not0;
  wire f_arrdiv32_fs905_and0;
  wire f_arrdiv32_fs905_xor1;
  wire f_arrdiv32_fs905_not1;
  wire f_arrdiv32_fs905_and1;
  wire f_arrdiv32_fs905_or0;
  wire f_arrdiv32_fs906_xor0;
  wire f_arrdiv32_fs906_not0;
  wire f_arrdiv32_fs906_and0;
  wire f_arrdiv32_fs906_xor1;
  wire f_arrdiv32_fs906_not1;
  wire f_arrdiv32_fs906_and1;
  wire f_arrdiv32_fs906_or0;
  wire f_arrdiv32_fs907_xor0;
  wire f_arrdiv32_fs907_not0;
  wire f_arrdiv32_fs907_and0;
  wire f_arrdiv32_fs907_xor1;
  wire f_arrdiv32_fs907_not1;
  wire f_arrdiv32_fs907_and1;
  wire f_arrdiv32_fs907_or0;
  wire f_arrdiv32_fs908_xor0;
  wire f_arrdiv32_fs908_not0;
  wire f_arrdiv32_fs908_and0;
  wire f_arrdiv32_fs908_xor1;
  wire f_arrdiv32_fs908_not1;
  wire f_arrdiv32_fs908_and1;
  wire f_arrdiv32_fs908_or0;
  wire f_arrdiv32_fs909_xor0;
  wire f_arrdiv32_fs909_not0;
  wire f_arrdiv32_fs909_and0;
  wire f_arrdiv32_fs909_xor1;
  wire f_arrdiv32_fs909_not1;
  wire f_arrdiv32_fs909_and1;
  wire f_arrdiv32_fs909_or0;
  wire f_arrdiv32_fs910_xor0;
  wire f_arrdiv32_fs910_not0;
  wire f_arrdiv32_fs910_and0;
  wire f_arrdiv32_fs910_xor1;
  wire f_arrdiv32_fs910_not1;
  wire f_arrdiv32_fs910_and1;
  wire f_arrdiv32_fs910_or0;
  wire f_arrdiv32_fs911_xor0;
  wire f_arrdiv32_fs911_not0;
  wire f_arrdiv32_fs911_and0;
  wire f_arrdiv32_fs911_xor1;
  wire f_arrdiv32_fs911_not1;
  wire f_arrdiv32_fs911_and1;
  wire f_arrdiv32_fs911_or0;
  wire f_arrdiv32_fs912_xor0;
  wire f_arrdiv32_fs912_not0;
  wire f_arrdiv32_fs912_and0;
  wire f_arrdiv32_fs912_xor1;
  wire f_arrdiv32_fs912_not1;
  wire f_arrdiv32_fs912_and1;
  wire f_arrdiv32_fs912_or0;
  wire f_arrdiv32_fs913_xor0;
  wire f_arrdiv32_fs913_not0;
  wire f_arrdiv32_fs913_and0;
  wire f_arrdiv32_fs913_xor1;
  wire f_arrdiv32_fs913_not1;
  wire f_arrdiv32_fs913_and1;
  wire f_arrdiv32_fs913_or0;
  wire f_arrdiv32_fs914_xor0;
  wire f_arrdiv32_fs914_not0;
  wire f_arrdiv32_fs914_and0;
  wire f_arrdiv32_fs914_xor1;
  wire f_arrdiv32_fs914_not1;
  wire f_arrdiv32_fs914_and1;
  wire f_arrdiv32_fs914_or0;
  wire f_arrdiv32_fs915_xor0;
  wire f_arrdiv32_fs915_not0;
  wire f_arrdiv32_fs915_and0;
  wire f_arrdiv32_fs915_xor1;
  wire f_arrdiv32_fs915_not1;
  wire f_arrdiv32_fs915_and1;
  wire f_arrdiv32_fs915_or0;
  wire f_arrdiv32_fs916_xor0;
  wire f_arrdiv32_fs916_not0;
  wire f_arrdiv32_fs916_and0;
  wire f_arrdiv32_fs916_xor1;
  wire f_arrdiv32_fs916_not1;
  wire f_arrdiv32_fs916_and1;
  wire f_arrdiv32_fs916_or0;
  wire f_arrdiv32_fs917_xor0;
  wire f_arrdiv32_fs917_not0;
  wire f_arrdiv32_fs917_and0;
  wire f_arrdiv32_fs917_xor1;
  wire f_arrdiv32_fs917_not1;
  wire f_arrdiv32_fs917_and1;
  wire f_arrdiv32_fs917_or0;
  wire f_arrdiv32_fs918_xor0;
  wire f_arrdiv32_fs918_not0;
  wire f_arrdiv32_fs918_and0;
  wire f_arrdiv32_fs918_xor1;
  wire f_arrdiv32_fs918_not1;
  wire f_arrdiv32_fs918_and1;
  wire f_arrdiv32_fs918_or0;
  wire f_arrdiv32_fs919_xor0;
  wire f_arrdiv32_fs919_not0;
  wire f_arrdiv32_fs919_and0;
  wire f_arrdiv32_fs919_xor1;
  wire f_arrdiv32_fs919_not1;
  wire f_arrdiv32_fs919_and1;
  wire f_arrdiv32_fs919_or0;
  wire f_arrdiv32_fs920_xor0;
  wire f_arrdiv32_fs920_not0;
  wire f_arrdiv32_fs920_and0;
  wire f_arrdiv32_fs920_xor1;
  wire f_arrdiv32_fs920_not1;
  wire f_arrdiv32_fs920_and1;
  wire f_arrdiv32_fs920_or0;
  wire f_arrdiv32_fs921_xor0;
  wire f_arrdiv32_fs921_not0;
  wire f_arrdiv32_fs921_and0;
  wire f_arrdiv32_fs921_xor1;
  wire f_arrdiv32_fs921_not1;
  wire f_arrdiv32_fs921_and1;
  wire f_arrdiv32_fs921_or0;
  wire f_arrdiv32_fs922_xor0;
  wire f_arrdiv32_fs922_not0;
  wire f_arrdiv32_fs922_and0;
  wire f_arrdiv32_fs922_xor1;
  wire f_arrdiv32_fs922_not1;
  wire f_arrdiv32_fs922_and1;
  wire f_arrdiv32_fs922_or0;
  wire f_arrdiv32_fs923_xor0;
  wire f_arrdiv32_fs923_not0;
  wire f_arrdiv32_fs923_and0;
  wire f_arrdiv32_fs923_xor1;
  wire f_arrdiv32_fs923_not1;
  wire f_arrdiv32_fs923_and1;
  wire f_arrdiv32_fs923_or0;
  wire f_arrdiv32_fs924_xor0;
  wire f_arrdiv32_fs924_not0;
  wire f_arrdiv32_fs924_and0;
  wire f_arrdiv32_fs924_xor1;
  wire f_arrdiv32_fs924_not1;
  wire f_arrdiv32_fs924_and1;
  wire f_arrdiv32_fs924_or0;
  wire f_arrdiv32_fs925_xor0;
  wire f_arrdiv32_fs925_not0;
  wire f_arrdiv32_fs925_and0;
  wire f_arrdiv32_fs925_xor1;
  wire f_arrdiv32_fs925_not1;
  wire f_arrdiv32_fs925_and1;
  wire f_arrdiv32_fs925_or0;
  wire f_arrdiv32_fs926_xor0;
  wire f_arrdiv32_fs926_not0;
  wire f_arrdiv32_fs926_and0;
  wire f_arrdiv32_fs926_xor1;
  wire f_arrdiv32_fs926_not1;
  wire f_arrdiv32_fs926_and1;
  wire f_arrdiv32_fs926_or0;
  wire f_arrdiv32_fs927_xor0;
  wire f_arrdiv32_fs927_not0;
  wire f_arrdiv32_fs927_and0;
  wire f_arrdiv32_fs927_xor1;
  wire f_arrdiv32_fs927_not1;
  wire f_arrdiv32_fs927_and1;
  wire f_arrdiv32_fs927_or0;
  wire f_arrdiv32_mux2to1868_and0;
  wire f_arrdiv32_mux2to1868_not0;
  wire f_arrdiv32_mux2to1868_and1;
  wire f_arrdiv32_mux2to1868_xor0;
  wire f_arrdiv32_mux2to1869_and0;
  wire f_arrdiv32_mux2to1869_not0;
  wire f_arrdiv32_mux2to1869_and1;
  wire f_arrdiv32_mux2to1869_xor0;
  wire f_arrdiv32_mux2to1870_and0;
  wire f_arrdiv32_mux2to1870_not0;
  wire f_arrdiv32_mux2to1870_and1;
  wire f_arrdiv32_mux2to1870_xor0;
  wire f_arrdiv32_mux2to1871_and0;
  wire f_arrdiv32_mux2to1871_not0;
  wire f_arrdiv32_mux2to1871_and1;
  wire f_arrdiv32_mux2to1871_xor0;
  wire f_arrdiv32_mux2to1872_and0;
  wire f_arrdiv32_mux2to1872_not0;
  wire f_arrdiv32_mux2to1872_and1;
  wire f_arrdiv32_mux2to1872_xor0;
  wire f_arrdiv32_mux2to1873_and0;
  wire f_arrdiv32_mux2to1873_not0;
  wire f_arrdiv32_mux2to1873_and1;
  wire f_arrdiv32_mux2to1873_xor0;
  wire f_arrdiv32_mux2to1874_and0;
  wire f_arrdiv32_mux2to1874_not0;
  wire f_arrdiv32_mux2to1874_and1;
  wire f_arrdiv32_mux2to1874_xor0;
  wire f_arrdiv32_mux2to1875_and0;
  wire f_arrdiv32_mux2to1875_not0;
  wire f_arrdiv32_mux2to1875_and1;
  wire f_arrdiv32_mux2to1875_xor0;
  wire f_arrdiv32_mux2to1876_and0;
  wire f_arrdiv32_mux2to1876_not0;
  wire f_arrdiv32_mux2to1876_and1;
  wire f_arrdiv32_mux2to1876_xor0;
  wire f_arrdiv32_mux2to1877_and0;
  wire f_arrdiv32_mux2to1877_not0;
  wire f_arrdiv32_mux2to1877_and1;
  wire f_arrdiv32_mux2to1877_xor0;
  wire f_arrdiv32_mux2to1878_and0;
  wire f_arrdiv32_mux2to1878_not0;
  wire f_arrdiv32_mux2to1878_and1;
  wire f_arrdiv32_mux2to1878_xor0;
  wire f_arrdiv32_mux2to1879_and0;
  wire f_arrdiv32_mux2to1879_not0;
  wire f_arrdiv32_mux2to1879_and1;
  wire f_arrdiv32_mux2to1879_xor0;
  wire f_arrdiv32_mux2to1880_and0;
  wire f_arrdiv32_mux2to1880_not0;
  wire f_arrdiv32_mux2to1880_and1;
  wire f_arrdiv32_mux2to1880_xor0;
  wire f_arrdiv32_mux2to1881_and0;
  wire f_arrdiv32_mux2to1881_not0;
  wire f_arrdiv32_mux2to1881_and1;
  wire f_arrdiv32_mux2to1881_xor0;
  wire f_arrdiv32_mux2to1882_and0;
  wire f_arrdiv32_mux2to1882_not0;
  wire f_arrdiv32_mux2to1882_and1;
  wire f_arrdiv32_mux2to1882_xor0;
  wire f_arrdiv32_mux2to1883_and0;
  wire f_arrdiv32_mux2to1883_not0;
  wire f_arrdiv32_mux2to1883_and1;
  wire f_arrdiv32_mux2to1883_xor0;
  wire f_arrdiv32_mux2to1884_and0;
  wire f_arrdiv32_mux2to1884_not0;
  wire f_arrdiv32_mux2to1884_and1;
  wire f_arrdiv32_mux2to1884_xor0;
  wire f_arrdiv32_mux2to1885_and0;
  wire f_arrdiv32_mux2to1885_not0;
  wire f_arrdiv32_mux2to1885_and1;
  wire f_arrdiv32_mux2to1885_xor0;
  wire f_arrdiv32_mux2to1886_and0;
  wire f_arrdiv32_mux2to1886_not0;
  wire f_arrdiv32_mux2to1886_and1;
  wire f_arrdiv32_mux2to1886_xor0;
  wire f_arrdiv32_mux2to1887_and0;
  wire f_arrdiv32_mux2to1887_not0;
  wire f_arrdiv32_mux2to1887_and1;
  wire f_arrdiv32_mux2to1887_xor0;
  wire f_arrdiv32_mux2to1888_and0;
  wire f_arrdiv32_mux2to1888_not0;
  wire f_arrdiv32_mux2to1888_and1;
  wire f_arrdiv32_mux2to1888_xor0;
  wire f_arrdiv32_mux2to1889_and0;
  wire f_arrdiv32_mux2to1889_not0;
  wire f_arrdiv32_mux2to1889_and1;
  wire f_arrdiv32_mux2to1889_xor0;
  wire f_arrdiv32_mux2to1890_and0;
  wire f_arrdiv32_mux2to1890_not0;
  wire f_arrdiv32_mux2to1890_and1;
  wire f_arrdiv32_mux2to1890_xor0;
  wire f_arrdiv32_mux2to1891_and0;
  wire f_arrdiv32_mux2to1891_not0;
  wire f_arrdiv32_mux2to1891_and1;
  wire f_arrdiv32_mux2to1891_xor0;
  wire f_arrdiv32_mux2to1892_and0;
  wire f_arrdiv32_mux2to1892_not0;
  wire f_arrdiv32_mux2to1892_and1;
  wire f_arrdiv32_mux2to1892_xor0;
  wire f_arrdiv32_mux2to1893_and0;
  wire f_arrdiv32_mux2to1893_not0;
  wire f_arrdiv32_mux2to1893_and1;
  wire f_arrdiv32_mux2to1893_xor0;
  wire f_arrdiv32_mux2to1894_and0;
  wire f_arrdiv32_mux2to1894_not0;
  wire f_arrdiv32_mux2to1894_and1;
  wire f_arrdiv32_mux2to1894_xor0;
  wire f_arrdiv32_mux2to1895_and0;
  wire f_arrdiv32_mux2to1895_not0;
  wire f_arrdiv32_mux2to1895_and1;
  wire f_arrdiv32_mux2to1895_xor0;
  wire f_arrdiv32_mux2to1896_and0;
  wire f_arrdiv32_mux2to1896_not0;
  wire f_arrdiv32_mux2to1896_and1;
  wire f_arrdiv32_mux2to1896_xor0;
  wire f_arrdiv32_mux2to1897_and0;
  wire f_arrdiv32_mux2to1897_not0;
  wire f_arrdiv32_mux2to1897_and1;
  wire f_arrdiv32_mux2to1897_xor0;
  wire f_arrdiv32_mux2to1898_and0;
  wire f_arrdiv32_mux2to1898_not0;
  wire f_arrdiv32_mux2to1898_and1;
  wire f_arrdiv32_mux2to1898_xor0;
  wire f_arrdiv32_not28;
  wire f_arrdiv32_fs928_xor0;
  wire f_arrdiv32_fs928_not0;
  wire f_arrdiv32_fs928_and0;
  wire f_arrdiv32_fs928_not1;
  wire f_arrdiv32_fs929_xor0;
  wire f_arrdiv32_fs929_not0;
  wire f_arrdiv32_fs929_and0;
  wire f_arrdiv32_fs929_xor1;
  wire f_arrdiv32_fs929_not1;
  wire f_arrdiv32_fs929_and1;
  wire f_arrdiv32_fs929_or0;
  wire f_arrdiv32_fs930_xor0;
  wire f_arrdiv32_fs930_not0;
  wire f_arrdiv32_fs930_and0;
  wire f_arrdiv32_fs930_xor1;
  wire f_arrdiv32_fs930_not1;
  wire f_arrdiv32_fs930_and1;
  wire f_arrdiv32_fs930_or0;
  wire f_arrdiv32_fs931_xor0;
  wire f_arrdiv32_fs931_not0;
  wire f_arrdiv32_fs931_and0;
  wire f_arrdiv32_fs931_xor1;
  wire f_arrdiv32_fs931_not1;
  wire f_arrdiv32_fs931_and1;
  wire f_arrdiv32_fs931_or0;
  wire f_arrdiv32_fs932_xor0;
  wire f_arrdiv32_fs932_not0;
  wire f_arrdiv32_fs932_and0;
  wire f_arrdiv32_fs932_xor1;
  wire f_arrdiv32_fs932_not1;
  wire f_arrdiv32_fs932_and1;
  wire f_arrdiv32_fs932_or0;
  wire f_arrdiv32_fs933_xor0;
  wire f_arrdiv32_fs933_not0;
  wire f_arrdiv32_fs933_and0;
  wire f_arrdiv32_fs933_xor1;
  wire f_arrdiv32_fs933_not1;
  wire f_arrdiv32_fs933_and1;
  wire f_arrdiv32_fs933_or0;
  wire f_arrdiv32_fs934_xor0;
  wire f_arrdiv32_fs934_not0;
  wire f_arrdiv32_fs934_and0;
  wire f_arrdiv32_fs934_xor1;
  wire f_arrdiv32_fs934_not1;
  wire f_arrdiv32_fs934_and1;
  wire f_arrdiv32_fs934_or0;
  wire f_arrdiv32_fs935_xor0;
  wire f_arrdiv32_fs935_not0;
  wire f_arrdiv32_fs935_and0;
  wire f_arrdiv32_fs935_xor1;
  wire f_arrdiv32_fs935_not1;
  wire f_arrdiv32_fs935_and1;
  wire f_arrdiv32_fs935_or0;
  wire f_arrdiv32_fs936_xor0;
  wire f_arrdiv32_fs936_not0;
  wire f_arrdiv32_fs936_and0;
  wire f_arrdiv32_fs936_xor1;
  wire f_arrdiv32_fs936_not1;
  wire f_arrdiv32_fs936_and1;
  wire f_arrdiv32_fs936_or0;
  wire f_arrdiv32_fs937_xor0;
  wire f_arrdiv32_fs937_not0;
  wire f_arrdiv32_fs937_and0;
  wire f_arrdiv32_fs937_xor1;
  wire f_arrdiv32_fs937_not1;
  wire f_arrdiv32_fs937_and1;
  wire f_arrdiv32_fs937_or0;
  wire f_arrdiv32_fs938_xor0;
  wire f_arrdiv32_fs938_not0;
  wire f_arrdiv32_fs938_and0;
  wire f_arrdiv32_fs938_xor1;
  wire f_arrdiv32_fs938_not1;
  wire f_arrdiv32_fs938_and1;
  wire f_arrdiv32_fs938_or0;
  wire f_arrdiv32_fs939_xor0;
  wire f_arrdiv32_fs939_not0;
  wire f_arrdiv32_fs939_and0;
  wire f_arrdiv32_fs939_xor1;
  wire f_arrdiv32_fs939_not1;
  wire f_arrdiv32_fs939_and1;
  wire f_arrdiv32_fs939_or0;
  wire f_arrdiv32_fs940_xor0;
  wire f_arrdiv32_fs940_not0;
  wire f_arrdiv32_fs940_and0;
  wire f_arrdiv32_fs940_xor1;
  wire f_arrdiv32_fs940_not1;
  wire f_arrdiv32_fs940_and1;
  wire f_arrdiv32_fs940_or0;
  wire f_arrdiv32_fs941_xor0;
  wire f_arrdiv32_fs941_not0;
  wire f_arrdiv32_fs941_and0;
  wire f_arrdiv32_fs941_xor1;
  wire f_arrdiv32_fs941_not1;
  wire f_arrdiv32_fs941_and1;
  wire f_arrdiv32_fs941_or0;
  wire f_arrdiv32_fs942_xor0;
  wire f_arrdiv32_fs942_not0;
  wire f_arrdiv32_fs942_and0;
  wire f_arrdiv32_fs942_xor1;
  wire f_arrdiv32_fs942_not1;
  wire f_arrdiv32_fs942_and1;
  wire f_arrdiv32_fs942_or0;
  wire f_arrdiv32_fs943_xor0;
  wire f_arrdiv32_fs943_not0;
  wire f_arrdiv32_fs943_and0;
  wire f_arrdiv32_fs943_xor1;
  wire f_arrdiv32_fs943_not1;
  wire f_arrdiv32_fs943_and1;
  wire f_arrdiv32_fs943_or0;
  wire f_arrdiv32_fs944_xor0;
  wire f_arrdiv32_fs944_not0;
  wire f_arrdiv32_fs944_and0;
  wire f_arrdiv32_fs944_xor1;
  wire f_arrdiv32_fs944_not1;
  wire f_arrdiv32_fs944_and1;
  wire f_arrdiv32_fs944_or0;
  wire f_arrdiv32_fs945_xor0;
  wire f_arrdiv32_fs945_not0;
  wire f_arrdiv32_fs945_and0;
  wire f_arrdiv32_fs945_xor1;
  wire f_arrdiv32_fs945_not1;
  wire f_arrdiv32_fs945_and1;
  wire f_arrdiv32_fs945_or0;
  wire f_arrdiv32_fs946_xor0;
  wire f_arrdiv32_fs946_not0;
  wire f_arrdiv32_fs946_and0;
  wire f_arrdiv32_fs946_xor1;
  wire f_arrdiv32_fs946_not1;
  wire f_arrdiv32_fs946_and1;
  wire f_arrdiv32_fs946_or0;
  wire f_arrdiv32_fs947_xor0;
  wire f_arrdiv32_fs947_not0;
  wire f_arrdiv32_fs947_and0;
  wire f_arrdiv32_fs947_xor1;
  wire f_arrdiv32_fs947_not1;
  wire f_arrdiv32_fs947_and1;
  wire f_arrdiv32_fs947_or0;
  wire f_arrdiv32_fs948_xor0;
  wire f_arrdiv32_fs948_not0;
  wire f_arrdiv32_fs948_and0;
  wire f_arrdiv32_fs948_xor1;
  wire f_arrdiv32_fs948_not1;
  wire f_arrdiv32_fs948_and1;
  wire f_arrdiv32_fs948_or0;
  wire f_arrdiv32_fs949_xor0;
  wire f_arrdiv32_fs949_not0;
  wire f_arrdiv32_fs949_and0;
  wire f_arrdiv32_fs949_xor1;
  wire f_arrdiv32_fs949_not1;
  wire f_arrdiv32_fs949_and1;
  wire f_arrdiv32_fs949_or0;
  wire f_arrdiv32_fs950_xor0;
  wire f_arrdiv32_fs950_not0;
  wire f_arrdiv32_fs950_and0;
  wire f_arrdiv32_fs950_xor1;
  wire f_arrdiv32_fs950_not1;
  wire f_arrdiv32_fs950_and1;
  wire f_arrdiv32_fs950_or0;
  wire f_arrdiv32_fs951_xor0;
  wire f_arrdiv32_fs951_not0;
  wire f_arrdiv32_fs951_and0;
  wire f_arrdiv32_fs951_xor1;
  wire f_arrdiv32_fs951_not1;
  wire f_arrdiv32_fs951_and1;
  wire f_arrdiv32_fs951_or0;
  wire f_arrdiv32_fs952_xor0;
  wire f_arrdiv32_fs952_not0;
  wire f_arrdiv32_fs952_and0;
  wire f_arrdiv32_fs952_xor1;
  wire f_arrdiv32_fs952_not1;
  wire f_arrdiv32_fs952_and1;
  wire f_arrdiv32_fs952_or0;
  wire f_arrdiv32_fs953_xor0;
  wire f_arrdiv32_fs953_not0;
  wire f_arrdiv32_fs953_and0;
  wire f_arrdiv32_fs953_xor1;
  wire f_arrdiv32_fs953_not1;
  wire f_arrdiv32_fs953_and1;
  wire f_arrdiv32_fs953_or0;
  wire f_arrdiv32_fs954_xor0;
  wire f_arrdiv32_fs954_not0;
  wire f_arrdiv32_fs954_and0;
  wire f_arrdiv32_fs954_xor1;
  wire f_arrdiv32_fs954_not1;
  wire f_arrdiv32_fs954_and1;
  wire f_arrdiv32_fs954_or0;
  wire f_arrdiv32_fs955_xor0;
  wire f_arrdiv32_fs955_not0;
  wire f_arrdiv32_fs955_and0;
  wire f_arrdiv32_fs955_xor1;
  wire f_arrdiv32_fs955_not1;
  wire f_arrdiv32_fs955_and1;
  wire f_arrdiv32_fs955_or0;
  wire f_arrdiv32_fs956_xor0;
  wire f_arrdiv32_fs956_not0;
  wire f_arrdiv32_fs956_and0;
  wire f_arrdiv32_fs956_xor1;
  wire f_arrdiv32_fs956_not1;
  wire f_arrdiv32_fs956_and1;
  wire f_arrdiv32_fs956_or0;
  wire f_arrdiv32_fs957_xor0;
  wire f_arrdiv32_fs957_not0;
  wire f_arrdiv32_fs957_and0;
  wire f_arrdiv32_fs957_xor1;
  wire f_arrdiv32_fs957_not1;
  wire f_arrdiv32_fs957_and1;
  wire f_arrdiv32_fs957_or0;
  wire f_arrdiv32_fs958_xor0;
  wire f_arrdiv32_fs958_not0;
  wire f_arrdiv32_fs958_and0;
  wire f_arrdiv32_fs958_xor1;
  wire f_arrdiv32_fs958_not1;
  wire f_arrdiv32_fs958_and1;
  wire f_arrdiv32_fs958_or0;
  wire f_arrdiv32_fs959_xor0;
  wire f_arrdiv32_fs959_not0;
  wire f_arrdiv32_fs959_and0;
  wire f_arrdiv32_fs959_xor1;
  wire f_arrdiv32_fs959_not1;
  wire f_arrdiv32_fs959_and1;
  wire f_arrdiv32_fs959_or0;
  wire f_arrdiv32_mux2to1899_and0;
  wire f_arrdiv32_mux2to1899_not0;
  wire f_arrdiv32_mux2to1899_and1;
  wire f_arrdiv32_mux2to1899_xor0;
  wire f_arrdiv32_mux2to1900_and0;
  wire f_arrdiv32_mux2to1900_not0;
  wire f_arrdiv32_mux2to1900_and1;
  wire f_arrdiv32_mux2to1900_xor0;
  wire f_arrdiv32_mux2to1901_and0;
  wire f_arrdiv32_mux2to1901_not0;
  wire f_arrdiv32_mux2to1901_and1;
  wire f_arrdiv32_mux2to1901_xor0;
  wire f_arrdiv32_mux2to1902_and0;
  wire f_arrdiv32_mux2to1902_not0;
  wire f_arrdiv32_mux2to1902_and1;
  wire f_arrdiv32_mux2to1902_xor0;
  wire f_arrdiv32_mux2to1903_and0;
  wire f_arrdiv32_mux2to1903_not0;
  wire f_arrdiv32_mux2to1903_and1;
  wire f_arrdiv32_mux2to1903_xor0;
  wire f_arrdiv32_mux2to1904_and0;
  wire f_arrdiv32_mux2to1904_not0;
  wire f_arrdiv32_mux2to1904_and1;
  wire f_arrdiv32_mux2to1904_xor0;
  wire f_arrdiv32_mux2to1905_and0;
  wire f_arrdiv32_mux2to1905_not0;
  wire f_arrdiv32_mux2to1905_and1;
  wire f_arrdiv32_mux2to1905_xor0;
  wire f_arrdiv32_mux2to1906_and0;
  wire f_arrdiv32_mux2to1906_not0;
  wire f_arrdiv32_mux2to1906_and1;
  wire f_arrdiv32_mux2to1906_xor0;
  wire f_arrdiv32_mux2to1907_and0;
  wire f_arrdiv32_mux2to1907_not0;
  wire f_arrdiv32_mux2to1907_and1;
  wire f_arrdiv32_mux2to1907_xor0;
  wire f_arrdiv32_mux2to1908_and0;
  wire f_arrdiv32_mux2to1908_not0;
  wire f_arrdiv32_mux2to1908_and1;
  wire f_arrdiv32_mux2to1908_xor0;
  wire f_arrdiv32_mux2to1909_and0;
  wire f_arrdiv32_mux2to1909_not0;
  wire f_arrdiv32_mux2to1909_and1;
  wire f_arrdiv32_mux2to1909_xor0;
  wire f_arrdiv32_mux2to1910_and0;
  wire f_arrdiv32_mux2to1910_not0;
  wire f_arrdiv32_mux2to1910_and1;
  wire f_arrdiv32_mux2to1910_xor0;
  wire f_arrdiv32_mux2to1911_and0;
  wire f_arrdiv32_mux2to1911_not0;
  wire f_arrdiv32_mux2to1911_and1;
  wire f_arrdiv32_mux2to1911_xor0;
  wire f_arrdiv32_mux2to1912_and0;
  wire f_arrdiv32_mux2to1912_not0;
  wire f_arrdiv32_mux2to1912_and1;
  wire f_arrdiv32_mux2to1912_xor0;
  wire f_arrdiv32_mux2to1913_and0;
  wire f_arrdiv32_mux2to1913_not0;
  wire f_arrdiv32_mux2to1913_and1;
  wire f_arrdiv32_mux2to1913_xor0;
  wire f_arrdiv32_mux2to1914_and0;
  wire f_arrdiv32_mux2to1914_not0;
  wire f_arrdiv32_mux2to1914_and1;
  wire f_arrdiv32_mux2to1914_xor0;
  wire f_arrdiv32_mux2to1915_and0;
  wire f_arrdiv32_mux2to1915_not0;
  wire f_arrdiv32_mux2to1915_and1;
  wire f_arrdiv32_mux2to1915_xor0;
  wire f_arrdiv32_mux2to1916_and0;
  wire f_arrdiv32_mux2to1916_not0;
  wire f_arrdiv32_mux2to1916_and1;
  wire f_arrdiv32_mux2to1916_xor0;
  wire f_arrdiv32_mux2to1917_and0;
  wire f_arrdiv32_mux2to1917_not0;
  wire f_arrdiv32_mux2to1917_and1;
  wire f_arrdiv32_mux2to1917_xor0;
  wire f_arrdiv32_mux2to1918_and0;
  wire f_arrdiv32_mux2to1918_not0;
  wire f_arrdiv32_mux2to1918_and1;
  wire f_arrdiv32_mux2to1918_xor0;
  wire f_arrdiv32_mux2to1919_and0;
  wire f_arrdiv32_mux2to1919_not0;
  wire f_arrdiv32_mux2to1919_and1;
  wire f_arrdiv32_mux2to1919_xor0;
  wire f_arrdiv32_mux2to1920_and0;
  wire f_arrdiv32_mux2to1920_not0;
  wire f_arrdiv32_mux2to1920_and1;
  wire f_arrdiv32_mux2to1920_xor0;
  wire f_arrdiv32_mux2to1921_and0;
  wire f_arrdiv32_mux2to1921_not0;
  wire f_arrdiv32_mux2to1921_and1;
  wire f_arrdiv32_mux2to1921_xor0;
  wire f_arrdiv32_mux2to1922_and0;
  wire f_arrdiv32_mux2to1922_not0;
  wire f_arrdiv32_mux2to1922_and1;
  wire f_arrdiv32_mux2to1922_xor0;
  wire f_arrdiv32_mux2to1923_and0;
  wire f_arrdiv32_mux2to1923_not0;
  wire f_arrdiv32_mux2to1923_and1;
  wire f_arrdiv32_mux2to1923_xor0;
  wire f_arrdiv32_mux2to1924_and0;
  wire f_arrdiv32_mux2to1924_not0;
  wire f_arrdiv32_mux2to1924_and1;
  wire f_arrdiv32_mux2to1924_xor0;
  wire f_arrdiv32_mux2to1925_and0;
  wire f_arrdiv32_mux2to1925_not0;
  wire f_arrdiv32_mux2to1925_and1;
  wire f_arrdiv32_mux2to1925_xor0;
  wire f_arrdiv32_mux2to1926_and0;
  wire f_arrdiv32_mux2to1926_not0;
  wire f_arrdiv32_mux2to1926_and1;
  wire f_arrdiv32_mux2to1926_xor0;
  wire f_arrdiv32_mux2to1927_and0;
  wire f_arrdiv32_mux2to1927_not0;
  wire f_arrdiv32_mux2to1927_and1;
  wire f_arrdiv32_mux2to1927_xor0;
  wire f_arrdiv32_mux2to1928_and0;
  wire f_arrdiv32_mux2to1928_not0;
  wire f_arrdiv32_mux2to1928_and1;
  wire f_arrdiv32_mux2to1928_xor0;
  wire f_arrdiv32_mux2to1929_and0;
  wire f_arrdiv32_mux2to1929_not0;
  wire f_arrdiv32_mux2to1929_and1;
  wire f_arrdiv32_mux2to1929_xor0;
  wire f_arrdiv32_not29;
  wire f_arrdiv32_fs960_xor0;
  wire f_arrdiv32_fs960_not0;
  wire f_arrdiv32_fs960_and0;
  wire f_arrdiv32_fs960_not1;
  wire f_arrdiv32_fs961_xor0;
  wire f_arrdiv32_fs961_not0;
  wire f_arrdiv32_fs961_and0;
  wire f_arrdiv32_fs961_xor1;
  wire f_arrdiv32_fs961_not1;
  wire f_arrdiv32_fs961_and1;
  wire f_arrdiv32_fs961_or0;
  wire f_arrdiv32_fs962_xor0;
  wire f_arrdiv32_fs962_not0;
  wire f_arrdiv32_fs962_and0;
  wire f_arrdiv32_fs962_xor1;
  wire f_arrdiv32_fs962_not1;
  wire f_arrdiv32_fs962_and1;
  wire f_arrdiv32_fs962_or0;
  wire f_arrdiv32_fs963_xor0;
  wire f_arrdiv32_fs963_not0;
  wire f_arrdiv32_fs963_and0;
  wire f_arrdiv32_fs963_xor1;
  wire f_arrdiv32_fs963_not1;
  wire f_arrdiv32_fs963_and1;
  wire f_arrdiv32_fs963_or0;
  wire f_arrdiv32_fs964_xor0;
  wire f_arrdiv32_fs964_not0;
  wire f_arrdiv32_fs964_and0;
  wire f_arrdiv32_fs964_xor1;
  wire f_arrdiv32_fs964_not1;
  wire f_arrdiv32_fs964_and1;
  wire f_arrdiv32_fs964_or0;
  wire f_arrdiv32_fs965_xor0;
  wire f_arrdiv32_fs965_not0;
  wire f_arrdiv32_fs965_and0;
  wire f_arrdiv32_fs965_xor1;
  wire f_arrdiv32_fs965_not1;
  wire f_arrdiv32_fs965_and1;
  wire f_arrdiv32_fs965_or0;
  wire f_arrdiv32_fs966_xor0;
  wire f_arrdiv32_fs966_not0;
  wire f_arrdiv32_fs966_and0;
  wire f_arrdiv32_fs966_xor1;
  wire f_arrdiv32_fs966_not1;
  wire f_arrdiv32_fs966_and1;
  wire f_arrdiv32_fs966_or0;
  wire f_arrdiv32_fs967_xor0;
  wire f_arrdiv32_fs967_not0;
  wire f_arrdiv32_fs967_and0;
  wire f_arrdiv32_fs967_xor1;
  wire f_arrdiv32_fs967_not1;
  wire f_arrdiv32_fs967_and1;
  wire f_arrdiv32_fs967_or0;
  wire f_arrdiv32_fs968_xor0;
  wire f_arrdiv32_fs968_not0;
  wire f_arrdiv32_fs968_and0;
  wire f_arrdiv32_fs968_xor1;
  wire f_arrdiv32_fs968_not1;
  wire f_arrdiv32_fs968_and1;
  wire f_arrdiv32_fs968_or0;
  wire f_arrdiv32_fs969_xor0;
  wire f_arrdiv32_fs969_not0;
  wire f_arrdiv32_fs969_and0;
  wire f_arrdiv32_fs969_xor1;
  wire f_arrdiv32_fs969_not1;
  wire f_arrdiv32_fs969_and1;
  wire f_arrdiv32_fs969_or0;
  wire f_arrdiv32_fs970_xor0;
  wire f_arrdiv32_fs970_not0;
  wire f_arrdiv32_fs970_and0;
  wire f_arrdiv32_fs970_xor1;
  wire f_arrdiv32_fs970_not1;
  wire f_arrdiv32_fs970_and1;
  wire f_arrdiv32_fs970_or0;
  wire f_arrdiv32_fs971_xor0;
  wire f_arrdiv32_fs971_not0;
  wire f_arrdiv32_fs971_and0;
  wire f_arrdiv32_fs971_xor1;
  wire f_arrdiv32_fs971_not1;
  wire f_arrdiv32_fs971_and1;
  wire f_arrdiv32_fs971_or0;
  wire f_arrdiv32_fs972_xor0;
  wire f_arrdiv32_fs972_not0;
  wire f_arrdiv32_fs972_and0;
  wire f_arrdiv32_fs972_xor1;
  wire f_arrdiv32_fs972_not1;
  wire f_arrdiv32_fs972_and1;
  wire f_arrdiv32_fs972_or0;
  wire f_arrdiv32_fs973_xor0;
  wire f_arrdiv32_fs973_not0;
  wire f_arrdiv32_fs973_and0;
  wire f_arrdiv32_fs973_xor1;
  wire f_arrdiv32_fs973_not1;
  wire f_arrdiv32_fs973_and1;
  wire f_arrdiv32_fs973_or0;
  wire f_arrdiv32_fs974_xor0;
  wire f_arrdiv32_fs974_not0;
  wire f_arrdiv32_fs974_and0;
  wire f_arrdiv32_fs974_xor1;
  wire f_arrdiv32_fs974_not1;
  wire f_arrdiv32_fs974_and1;
  wire f_arrdiv32_fs974_or0;
  wire f_arrdiv32_fs975_xor0;
  wire f_arrdiv32_fs975_not0;
  wire f_arrdiv32_fs975_and0;
  wire f_arrdiv32_fs975_xor1;
  wire f_arrdiv32_fs975_not1;
  wire f_arrdiv32_fs975_and1;
  wire f_arrdiv32_fs975_or0;
  wire f_arrdiv32_fs976_xor0;
  wire f_arrdiv32_fs976_not0;
  wire f_arrdiv32_fs976_and0;
  wire f_arrdiv32_fs976_xor1;
  wire f_arrdiv32_fs976_not1;
  wire f_arrdiv32_fs976_and1;
  wire f_arrdiv32_fs976_or0;
  wire f_arrdiv32_fs977_xor0;
  wire f_arrdiv32_fs977_not0;
  wire f_arrdiv32_fs977_and0;
  wire f_arrdiv32_fs977_xor1;
  wire f_arrdiv32_fs977_not1;
  wire f_arrdiv32_fs977_and1;
  wire f_arrdiv32_fs977_or0;
  wire f_arrdiv32_fs978_xor0;
  wire f_arrdiv32_fs978_not0;
  wire f_arrdiv32_fs978_and0;
  wire f_arrdiv32_fs978_xor1;
  wire f_arrdiv32_fs978_not1;
  wire f_arrdiv32_fs978_and1;
  wire f_arrdiv32_fs978_or0;
  wire f_arrdiv32_fs979_xor0;
  wire f_arrdiv32_fs979_not0;
  wire f_arrdiv32_fs979_and0;
  wire f_arrdiv32_fs979_xor1;
  wire f_arrdiv32_fs979_not1;
  wire f_arrdiv32_fs979_and1;
  wire f_arrdiv32_fs979_or0;
  wire f_arrdiv32_fs980_xor0;
  wire f_arrdiv32_fs980_not0;
  wire f_arrdiv32_fs980_and0;
  wire f_arrdiv32_fs980_xor1;
  wire f_arrdiv32_fs980_not1;
  wire f_arrdiv32_fs980_and1;
  wire f_arrdiv32_fs980_or0;
  wire f_arrdiv32_fs981_xor0;
  wire f_arrdiv32_fs981_not0;
  wire f_arrdiv32_fs981_and0;
  wire f_arrdiv32_fs981_xor1;
  wire f_arrdiv32_fs981_not1;
  wire f_arrdiv32_fs981_and1;
  wire f_arrdiv32_fs981_or0;
  wire f_arrdiv32_fs982_xor0;
  wire f_arrdiv32_fs982_not0;
  wire f_arrdiv32_fs982_and0;
  wire f_arrdiv32_fs982_xor1;
  wire f_arrdiv32_fs982_not1;
  wire f_arrdiv32_fs982_and1;
  wire f_arrdiv32_fs982_or0;
  wire f_arrdiv32_fs983_xor0;
  wire f_arrdiv32_fs983_not0;
  wire f_arrdiv32_fs983_and0;
  wire f_arrdiv32_fs983_xor1;
  wire f_arrdiv32_fs983_not1;
  wire f_arrdiv32_fs983_and1;
  wire f_arrdiv32_fs983_or0;
  wire f_arrdiv32_fs984_xor0;
  wire f_arrdiv32_fs984_not0;
  wire f_arrdiv32_fs984_and0;
  wire f_arrdiv32_fs984_xor1;
  wire f_arrdiv32_fs984_not1;
  wire f_arrdiv32_fs984_and1;
  wire f_arrdiv32_fs984_or0;
  wire f_arrdiv32_fs985_xor0;
  wire f_arrdiv32_fs985_not0;
  wire f_arrdiv32_fs985_and0;
  wire f_arrdiv32_fs985_xor1;
  wire f_arrdiv32_fs985_not1;
  wire f_arrdiv32_fs985_and1;
  wire f_arrdiv32_fs985_or0;
  wire f_arrdiv32_fs986_xor0;
  wire f_arrdiv32_fs986_not0;
  wire f_arrdiv32_fs986_and0;
  wire f_arrdiv32_fs986_xor1;
  wire f_arrdiv32_fs986_not1;
  wire f_arrdiv32_fs986_and1;
  wire f_arrdiv32_fs986_or0;
  wire f_arrdiv32_fs987_xor0;
  wire f_arrdiv32_fs987_not0;
  wire f_arrdiv32_fs987_and0;
  wire f_arrdiv32_fs987_xor1;
  wire f_arrdiv32_fs987_not1;
  wire f_arrdiv32_fs987_and1;
  wire f_arrdiv32_fs987_or0;
  wire f_arrdiv32_fs988_xor0;
  wire f_arrdiv32_fs988_not0;
  wire f_arrdiv32_fs988_and0;
  wire f_arrdiv32_fs988_xor1;
  wire f_arrdiv32_fs988_not1;
  wire f_arrdiv32_fs988_and1;
  wire f_arrdiv32_fs988_or0;
  wire f_arrdiv32_fs989_xor0;
  wire f_arrdiv32_fs989_not0;
  wire f_arrdiv32_fs989_and0;
  wire f_arrdiv32_fs989_xor1;
  wire f_arrdiv32_fs989_not1;
  wire f_arrdiv32_fs989_and1;
  wire f_arrdiv32_fs989_or0;
  wire f_arrdiv32_fs990_xor0;
  wire f_arrdiv32_fs990_not0;
  wire f_arrdiv32_fs990_and0;
  wire f_arrdiv32_fs990_xor1;
  wire f_arrdiv32_fs990_not1;
  wire f_arrdiv32_fs990_and1;
  wire f_arrdiv32_fs990_or0;
  wire f_arrdiv32_fs991_xor0;
  wire f_arrdiv32_fs991_not0;
  wire f_arrdiv32_fs991_and0;
  wire f_arrdiv32_fs991_xor1;
  wire f_arrdiv32_fs991_not1;
  wire f_arrdiv32_fs991_and1;
  wire f_arrdiv32_fs991_or0;
  wire f_arrdiv32_mux2to1930_and0;
  wire f_arrdiv32_mux2to1930_not0;
  wire f_arrdiv32_mux2to1930_and1;
  wire f_arrdiv32_mux2to1930_xor0;
  wire f_arrdiv32_mux2to1931_and0;
  wire f_arrdiv32_mux2to1931_not0;
  wire f_arrdiv32_mux2to1931_and1;
  wire f_arrdiv32_mux2to1931_xor0;
  wire f_arrdiv32_mux2to1932_and0;
  wire f_arrdiv32_mux2to1932_not0;
  wire f_arrdiv32_mux2to1932_and1;
  wire f_arrdiv32_mux2to1932_xor0;
  wire f_arrdiv32_mux2to1933_and0;
  wire f_arrdiv32_mux2to1933_not0;
  wire f_arrdiv32_mux2to1933_and1;
  wire f_arrdiv32_mux2to1933_xor0;
  wire f_arrdiv32_mux2to1934_and0;
  wire f_arrdiv32_mux2to1934_not0;
  wire f_arrdiv32_mux2to1934_and1;
  wire f_arrdiv32_mux2to1934_xor0;
  wire f_arrdiv32_mux2to1935_and0;
  wire f_arrdiv32_mux2to1935_not0;
  wire f_arrdiv32_mux2to1935_and1;
  wire f_arrdiv32_mux2to1935_xor0;
  wire f_arrdiv32_mux2to1936_and0;
  wire f_arrdiv32_mux2to1936_not0;
  wire f_arrdiv32_mux2to1936_and1;
  wire f_arrdiv32_mux2to1936_xor0;
  wire f_arrdiv32_mux2to1937_and0;
  wire f_arrdiv32_mux2to1937_not0;
  wire f_arrdiv32_mux2to1937_and1;
  wire f_arrdiv32_mux2to1937_xor0;
  wire f_arrdiv32_mux2to1938_and0;
  wire f_arrdiv32_mux2to1938_not0;
  wire f_arrdiv32_mux2to1938_and1;
  wire f_arrdiv32_mux2to1938_xor0;
  wire f_arrdiv32_mux2to1939_and0;
  wire f_arrdiv32_mux2to1939_not0;
  wire f_arrdiv32_mux2to1939_and1;
  wire f_arrdiv32_mux2to1939_xor0;
  wire f_arrdiv32_mux2to1940_and0;
  wire f_arrdiv32_mux2to1940_not0;
  wire f_arrdiv32_mux2to1940_and1;
  wire f_arrdiv32_mux2to1940_xor0;
  wire f_arrdiv32_mux2to1941_and0;
  wire f_arrdiv32_mux2to1941_not0;
  wire f_arrdiv32_mux2to1941_and1;
  wire f_arrdiv32_mux2to1941_xor0;
  wire f_arrdiv32_mux2to1942_and0;
  wire f_arrdiv32_mux2to1942_not0;
  wire f_arrdiv32_mux2to1942_and1;
  wire f_arrdiv32_mux2to1942_xor0;
  wire f_arrdiv32_mux2to1943_and0;
  wire f_arrdiv32_mux2to1943_not0;
  wire f_arrdiv32_mux2to1943_and1;
  wire f_arrdiv32_mux2to1943_xor0;
  wire f_arrdiv32_mux2to1944_and0;
  wire f_arrdiv32_mux2to1944_not0;
  wire f_arrdiv32_mux2to1944_and1;
  wire f_arrdiv32_mux2to1944_xor0;
  wire f_arrdiv32_mux2to1945_and0;
  wire f_arrdiv32_mux2to1945_not0;
  wire f_arrdiv32_mux2to1945_and1;
  wire f_arrdiv32_mux2to1945_xor0;
  wire f_arrdiv32_mux2to1946_and0;
  wire f_arrdiv32_mux2to1946_not0;
  wire f_arrdiv32_mux2to1946_and1;
  wire f_arrdiv32_mux2to1946_xor0;
  wire f_arrdiv32_mux2to1947_and0;
  wire f_arrdiv32_mux2to1947_not0;
  wire f_arrdiv32_mux2to1947_and1;
  wire f_arrdiv32_mux2to1947_xor0;
  wire f_arrdiv32_mux2to1948_and0;
  wire f_arrdiv32_mux2to1948_not0;
  wire f_arrdiv32_mux2to1948_and1;
  wire f_arrdiv32_mux2to1948_xor0;
  wire f_arrdiv32_mux2to1949_and0;
  wire f_arrdiv32_mux2to1949_not0;
  wire f_arrdiv32_mux2to1949_and1;
  wire f_arrdiv32_mux2to1949_xor0;
  wire f_arrdiv32_mux2to1950_and0;
  wire f_arrdiv32_mux2to1950_not0;
  wire f_arrdiv32_mux2to1950_and1;
  wire f_arrdiv32_mux2to1950_xor0;
  wire f_arrdiv32_mux2to1951_and0;
  wire f_arrdiv32_mux2to1951_not0;
  wire f_arrdiv32_mux2to1951_and1;
  wire f_arrdiv32_mux2to1951_xor0;
  wire f_arrdiv32_mux2to1952_and0;
  wire f_arrdiv32_mux2to1952_not0;
  wire f_arrdiv32_mux2to1952_and1;
  wire f_arrdiv32_mux2to1952_xor0;
  wire f_arrdiv32_mux2to1953_and0;
  wire f_arrdiv32_mux2to1953_not0;
  wire f_arrdiv32_mux2to1953_and1;
  wire f_arrdiv32_mux2to1953_xor0;
  wire f_arrdiv32_mux2to1954_and0;
  wire f_arrdiv32_mux2to1954_not0;
  wire f_arrdiv32_mux2to1954_and1;
  wire f_arrdiv32_mux2to1954_xor0;
  wire f_arrdiv32_mux2to1955_and0;
  wire f_arrdiv32_mux2to1955_not0;
  wire f_arrdiv32_mux2to1955_and1;
  wire f_arrdiv32_mux2to1955_xor0;
  wire f_arrdiv32_mux2to1956_and0;
  wire f_arrdiv32_mux2to1956_not0;
  wire f_arrdiv32_mux2to1956_and1;
  wire f_arrdiv32_mux2to1956_xor0;
  wire f_arrdiv32_mux2to1957_and0;
  wire f_arrdiv32_mux2to1957_not0;
  wire f_arrdiv32_mux2to1957_and1;
  wire f_arrdiv32_mux2to1957_xor0;
  wire f_arrdiv32_mux2to1958_and0;
  wire f_arrdiv32_mux2to1958_not0;
  wire f_arrdiv32_mux2to1958_and1;
  wire f_arrdiv32_mux2to1958_xor0;
  wire f_arrdiv32_mux2to1959_and0;
  wire f_arrdiv32_mux2to1959_not0;
  wire f_arrdiv32_mux2to1959_and1;
  wire f_arrdiv32_mux2to1959_xor0;
  wire f_arrdiv32_mux2to1960_and0;
  wire f_arrdiv32_mux2to1960_not0;
  wire f_arrdiv32_mux2to1960_and1;
  wire f_arrdiv32_mux2to1960_xor0;
  wire f_arrdiv32_not30;
  wire f_arrdiv32_fs992_xor0;
  wire f_arrdiv32_fs992_not0;
  wire f_arrdiv32_fs992_and0;
  wire f_arrdiv32_fs992_not1;
  wire f_arrdiv32_fs993_xor0;
  wire f_arrdiv32_fs993_not0;
  wire f_arrdiv32_fs993_and0;
  wire f_arrdiv32_fs993_xor1;
  wire f_arrdiv32_fs993_not1;
  wire f_arrdiv32_fs993_and1;
  wire f_arrdiv32_fs993_or0;
  wire f_arrdiv32_fs994_xor0;
  wire f_arrdiv32_fs994_not0;
  wire f_arrdiv32_fs994_and0;
  wire f_arrdiv32_fs994_xor1;
  wire f_arrdiv32_fs994_not1;
  wire f_arrdiv32_fs994_and1;
  wire f_arrdiv32_fs994_or0;
  wire f_arrdiv32_fs995_xor0;
  wire f_arrdiv32_fs995_not0;
  wire f_arrdiv32_fs995_and0;
  wire f_arrdiv32_fs995_xor1;
  wire f_arrdiv32_fs995_not1;
  wire f_arrdiv32_fs995_and1;
  wire f_arrdiv32_fs995_or0;
  wire f_arrdiv32_fs996_xor0;
  wire f_arrdiv32_fs996_not0;
  wire f_arrdiv32_fs996_and0;
  wire f_arrdiv32_fs996_xor1;
  wire f_arrdiv32_fs996_not1;
  wire f_arrdiv32_fs996_and1;
  wire f_arrdiv32_fs996_or0;
  wire f_arrdiv32_fs997_xor0;
  wire f_arrdiv32_fs997_not0;
  wire f_arrdiv32_fs997_and0;
  wire f_arrdiv32_fs997_xor1;
  wire f_arrdiv32_fs997_not1;
  wire f_arrdiv32_fs997_and1;
  wire f_arrdiv32_fs997_or0;
  wire f_arrdiv32_fs998_xor0;
  wire f_arrdiv32_fs998_not0;
  wire f_arrdiv32_fs998_and0;
  wire f_arrdiv32_fs998_xor1;
  wire f_arrdiv32_fs998_not1;
  wire f_arrdiv32_fs998_and1;
  wire f_arrdiv32_fs998_or0;
  wire f_arrdiv32_fs999_xor0;
  wire f_arrdiv32_fs999_not0;
  wire f_arrdiv32_fs999_and0;
  wire f_arrdiv32_fs999_xor1;
  wire f_arrdiv32_fs999_not1;
  wire f_arrdiv32_fs999_and1;
  wire f_arrdiv32_fs999_or0;
  wire f_arrdiv32_fs1000_xor0;
  wire f_arrdiv32_fs1000_not0;
  wire f_arrdiv32_fs1000_and0;
  wire f_arrdiv32_fs1000_xor1;
  wire f_arrdiv32_fs1000_not1;
  wire f_arrdiv32_fs1000_and1;
  wire f_arrdiv32_fs1000_or0;
  wire f_arrdiv32_fs1001_xor0;
  wire f_arrdiv32_fs1001_not0;
  wire f_arrdiv32_fs1001_and0;
  wire f_arrdiv32_fs1001_xor1;
  wire f_arrdiv32_fs1001_not1;
  wire f_arrdiv32_fs1001_and1;
  wire f_arrdiv32_fs1001_or0;
  wire f_arrdiv32_fs1002_xor0;
  wire f_arrdiv32_fs1002_not0;
  wire f_arrdiv32_fs1002_and0;
  wire f_arrdiv32_fs1002_xor1;
  wire f_arrdiv32_fs1002_not1;
  wire f_arrdiv32_fs1002_and1;
  wire f_arrdiv32_fs1002_or0;
  wire f_arrdiv32_fs1003_xor0;
  wire f_arrdiv32_fs1003_not0;
  wire f_arrdiv32_fs1003_and0;
  wire f_arrdiv32_fs1003_xor1;
  wire f_arrdiv32_fs1003_not1;
  wire f_arrdiv32_fs1003_and1;
  wire f_arrdiv32_fs1003_or0;
  wire f_arrdiv32_fs1004_xor0;
  wire f_arrdiv32_fs1004_not0;
  wire f_arrdiv32_fs1004_and0;
  wire f_arrdiv32_fs1004_xor1;
  wire f_arrdiv32_fs1004_not1;
  wire f_arrdiv32_fs1004_and1;
  wire f_arrdiv32_fs1004_or0;
  wire f_arrdiv32_fs1005_xor0;
  wire f_arrdiv32_fs1005_not0;
  wire f_arrdiv32_fs1005_and0;
  wire f_arrdiv32_fs1005_xor1;
  wire f_arrdiv32_fs1005_not1;
  wire f_arrdiv32_fs1005_and1;
  wire f_arrdiv32_fs1005_or0;
  wire f_arrdiv32_fs1006_xor0;
  wire f_arrdiv32_fs1006_not0;
  wire f_arrdiv32_fs1006_and0;
  wire f_arrdiv32_fs1006_xor1;
  wire f_arrdiv32_fs1006_not1;
  wire f_arrdiv32_fs1006_and1;
  wire f_arrdiv32_fs1006_or0;
  wire f_arrdiv32_fs1007_xor0;
  wire f_arrdiv32_fs1007_not0;
  wire f_arrdiv32_fs1007_and0;
  wire f_arrdiv32_fs1007_xor1;
  wire f_arrdiv32_fs1007_not1;
  wire f_arrdiv32_fs1007_and1;
  wire f_arrdiv32_fs1007_or0;
  wire f_arrdiv32_fs1008_xor0;
  wire f_arrdiv32_fs1008_not0;
  wire f_arrdiv32_fs1008_and0;
  wire f_arrdiv32_fs1008_xor1;
  wire f_arrdiv32_fs1008_not1;
  wire f_arrdiv32_fs1008_and1;
  wire f_arrdiv32_fs1008_or0;
  wire f_arrdiv32_fs1009_xor0;
  wire f_arrdiv32_fs1009_not0;
  wire f_arrdiv32_fs1009_and0;
  wire f_arrdiv32_fs1009_xor1;
  wire f_arrdiv32_fs1009_not1;
  wire f_arrdiv32_fs1009_and1;
  wire f_arrdiv32_fs1009_or0;
  wire f_arrdiv32_fs1010_xor0;
  wire f_arrdiv32_fs1010_not0;
  wire f_arrdiv32_fs1010_and0;
  wire f_arrdiv32_fs1010_xor1;
  wire f_arrdiv32_fs1010_not1;
  wire f_arrdiv32_fs1010_and1;
  wire f_arrdiv32_fs1010_or0;
  wire f_arrdiv32_fs1011_xor0;
  wire f_arrdiv32_fs1011_not0;
  wire f_arrdiv32_fs1011_and0;
  wire f_arrdiv32_fs1011_xor1;
  wire f_arrdiv32_fs1011_not1;
  wire f_arrdiv32_fs1011_and1;
  wire f_arrdiv32_fs1011_or0;
  wire f_arrdiv32_fs1012_xor0;
  wire f_arrdiv32_fs1012_not0;
  wire f_arrdiv32_fs1012_and0;
  wire f_arrdiv32_fs1012_xor1;
  wire f_arrdiv32_fs1012_not1;
  wire f_arrdiv32_fs1012_and1;
  wire f_arrdiv32_fs1012_or0;
  wire f_arrdiv32_fs1013_xor0;
  wire f_arrdiv32_fs1013_not0;
  wire f_arrdiv32_fs1013_and0;
  wire f_arrdiv32_fs1013_xor1;
  wire f_arrdiv32_fs1013_not1;
  wire f_arrdiv32_fs1013_and1;
  wire f_arrdiv32_fs1013_or0;
  wire f_arrdiv32_fs1014_xor0;
  wire f_arrdiv32_fs1014_not0;
  wire f_arrdiv32_fs1014_and0;
  wire f_arrdiv32_fs1014_xor1;
  wire f_arrdiv32_fs1014_not1;
  wire f_arrdiv32_fs1014_and1;
  wire f_arrdiv32_fs1014_or0;
  wire f_arrdiv32_fs1015_xor0;
  wire f_arrdiv32_fs1015_not0;
  wire f_arrdiv32_fs1015_and0;
  wire f_arrdiv32_fs1015_xor1;
  wire f_arrdiv32_fs1015_not1;
  wire f_arrdiv32_fs1015_and1;
  wire f_arrdiv32_fs1015_or0;
  wire f_arrdiv32_fs1016_xor0;
  wire f_arrdiv32_fs1016_not0;
  wire f_arrdiv32_fs1016_and0;
  wire f_arrdiv32_fs1016_xor1;
  wire f_arrdiv32_fs1016_not1;
  wire f_arrdiv32_fs1016_and1;
  wire f_arrdiv32_fs1016_or0;
  wire f_arrdiv32_fs1017_xor0;
  wire f_arrdiv32_fs1017_not0;
  wire f_arrdiv32_fs1017_and0;
  wire f_arrdiv32_fs1017_xor1;
  wire f_arrdiv32_fs1017_not1;
  wire f_arrdiv32_fs1017_and1;
  wire f_arrdiv32_fs1017_or0;
  wire f_arrdiv32_fs1018_xor0;
  wire f_arrdiv32_fs1018_not0;
  wire f_arrdiv32_fs1018_and0;
  wire f_arrdiv32_fs1018_xor1;
  wire f_arrdiv32_fs1018_not1;
  wire f_arrdiv32_fs1018_and1;
  wire f_arrdiv32_fs1018_or0;
  wire f_arrdiv32_fs1019_xor0;
  wire f_arrdiv32_fs1019_not0;
  wire f_arrdiv32_fs1019_and0;
  wire f_arrdiv32_fs1019_xor1;
  wire f_arrdiv32_fs1019_not1;
  wire f_arrdiv32_fs1019_and1;
  wire f_arrdiv32_fs1019_or0;
  wire f_arrdiv32_fs1020_xor0;
  wire f_arrdiv32_fs1020_not0;
  wire f_arrdiv32_fs1020_and0;
  wire f_arrdiv32_fs1020_xor1;
  wire f_arrdiv32_fs1020_not1;
  wire f_arrdiv32_fs1020_and1;
  wire f_arrdiv32_fs1020_or0;
  wire f_arrdiv32_fs1021_xor0;
  wire f_arrdiv32_fs1021_not0;
  wire f_arrdiv32_fs1021_and0;
  wire f_arrdiv32_fs1021_xor1;
  wire f_arrdiv32_fs1021_not1;
  wire f_arrdiv32_fs1021_and1;
  wire f_arrdiv32_fs1021_or0;
  wire f_arrdiv32_fs1022_xor0;
  wire f_arrdiv32_fs1022_not0;
  wire f_arrdiv32_fs1022_and0;
  wire f_arrdiv32_fs1022_xor1;
  wire f_arrdiv32_fs1022_not1;
  wire f_arrdiv32_fs1022_and1;
  wire f_arrdiv32_fs1022_or0;
  wire f_arrdiv32_fs1023_xor0;
  wire f_arrdiv32_fs1023_not0;
  wire f_arrdiv32_fs1023_and0;
  wire f_arrdiv32_fs1023_xor1;
  wire f_arrdiv32_fs1023_not1;
  wire f_arrdiv32_fs1023_and1;
  wire f_arrdiv32_fs1023_or0;
  wire f_arrdiv32_not31;

  assign f_arrdiv32_fs0_xor0 = a[31] ^ b[0];
  assign f_arrdiv32_fs0_not0 = ~a[31];
  assign f_arrdiv32_fs0_and0 = f_arrdiv32_fs0_not0 & b[0];
  assign f_arrdiv32_fs0_not1 = ~f_arrdiv32_fs0_xor0;
  assign f_arrdiv32_fs1_xor1 = f_arrdiv32_fs0_and0 ^ b[1];
  assign f_arrdiv32_fs1_not1 = ~b[1];
  assign f_arrdiv32_fs1_and1 = f_arrdiv32_fs1_not1 & f_arrdiv32_fs0_and0;
  assign f_arrdiv32_fs1_or0 = f_arrdiv32_fs1_and1 | b[1];
  assign f_arrdiv32_fs2_xor1 = f_arrdiv32_fs1_or0 ^ b[2];
  assign f_arrdiv32_fs2_not1 = ~b[2];
  assign f_arrdiv32_fs2_and1 = f_arrdiv32_fs2_not1 & f_arrdiv32_fs1_or0;
  assign f_arrdiv32_fs2_or0 = f_arrdiv32_fs2_and1 | b[2];
  assign f_arrdiv32_fs3_xor1 = f_arrdiv32_fs2_or0 ^ b[3];
  assign f_arrdiv32_fs3_not1 = ~b[3];
  assign f_arrdiv32_fs3_and1 = f_arrdiv32_fs3_not1 & f_arrdiv32_fs2_or0;
  assign f_arrdiv32_fs3_or0 = f_arrdiv32_fs3_and1 | b[3];
  assign f_arrdiv32_fs4_xor1 = f_arrdiv32_fs3_or0 ^ b[4];
  assign f_arrdiv32_fs4_not1 = ~b[4];
  assign f_arrdiv32_fs4_and1 = f_arrdiv32_fs4_not1 & f_arrdiv32_fs3_or0;
  assign f_arrdiv32_fs4_or0 = f_arrdiv32_fs4_and1 | b[4];
  assign f_arrdiv32_fs5_xor1 = f_arrdiv32_fs4_or0 ^ b[5];
  assign f_arrdiv32_fs5_not1 = ~b[5];
  assign f_arrdiv32_fs5_and1 = f_arrdiv32_fs5_not1 & f_arrdiv32_fs4_or0;
  assign f_arrdiv32_fs5_or0 = f_arrdiv32_fs5_and1 | b[5];
  assign f_arrdiv32_fs6_xor1 = f_arrdiv32_fs5_or0 ^ b[6];
  assign f_arrdiv32_fs6_not1 = ~b[6];
  assign f_arrdiv32_fs6_and1 = f_arrdiv32_fs6_not1 & f_arrdiv32_fs5_or0;
  assign f_arrdiv32_fs6_or0 = f_arrdiv32_fs6_and1 | b[6];
  assign f_arrdiv32_fs7_xor1 = f_arrdiv32_fs6_or0 ^ b[7];
  assign f_arrdiv32_fs7_not1 = ~b[7];
  assign f_arrdiv32_fs7_and1 = f_arrdiv32_fs7_not1 & f_arrdiv32_fs6_or0;
  assign f_arrdiv32_fs7_or0 = f_arrdiv32_fs7_and1 | b[7];
  assign f_arrdiv32_fs8_xor1 = f_arrdiv32_fs7_or0 ^ b[8];
  assign f_arrdiv32_fs8_not1 = ~b[8];
  assign f_arrdiv32_fs8_and1 = f_arrdiv32_fs8_not1 & f_arrdiv32_fs7_or0;
  assign f_arrdiv32_fs8_or0 = f_arrdiv32_fs8_and1 | b[8];
  assign f_arrdiv32_fs9_xor1 = f_arrdiv32_fs8_or0 ^ b[9];
  assign f_arrdiv32_fs9_not1 = ~b[9];
  assign f_arrdiv32_fs9_and1 = f_arrdiv32_fs9_not1 & f_arrdiv32_fs8_or0;
  assign f_arrdiv32_fs9_or0 = f_arrdiv32_fs9_and1 | b[9];
  assign f_arrdiv32_fs10_xor1 = f_arrdiv32_fs9_or0 ^ b[10];
  assign f_arrdiv32_fs10_not1 = ~b[10];
  assign f_arrdiv32_fs10_and1 = f_arrdiv32_fs10_not1 & f_arrdiv32_fs9_or0;
  assign f_arrdiv32_fs10_or0 = f_arrdiv32_fs10_and1 | b[10];
  assign f_arrdiv32_fs11_xor1 = f_arrdiv32_fs10_or0 ^ b[11];
  assign f_arrdiv32_fs11_not1 = ~b[11];
  assign f_arrdiv32_fs11_and1 = f_arrdiv32_fs11_not1 & f_arrdiv32_fs10_or0;
  assign f_arrdiv32_fs11_or0 = f_arrdiv32_fs11_and1 | b[11];
  assign f_arrdiv32_fs12_xor1 = f_arrdiv32_fs11_or0 ^ b[12];
  assign f_arrdiv32_fs12_not1 = ~b[12];
  assign f_arrdiv32_fs12_and1 = f_arrdiv32_fs12_not1 & f_arrdiv32_fs11_or0;
  assign f_arrdiv32_fs12_or0 = f_arrdiv32_fs12_and1 | b[12];
  assign f_arrdiv32_fs13_xor1 = f_arrdiv32_fs12_or0 ^ b[13];
  assign f_arrdiv32_fs13_not1 = ~b[13];
  assign f_arrdiv32_fs13_and1 = f_arrdiv32_fs13_not1 & f_arrdiv32_fs12_or0;
  assign f_arrdiv32_fs13_or0 = f_arrdiv32_fs13_and1 | b[13];
  assign f_arrdiv32_fs14_xor1 = f_arrdiv32_fs13_or0 ^ b[14];
  assign f_arrdiv32_fs14_not1 = ~b[14];
  assign f_arrdiv32_fs14_and1 = f_arrdiv32_fs14_not1 & f_arrdiv32_fs13_or0;
  assign f_arrdiv32_fs14_or0 = f_arrdiv32_fs14_and1 | b[14];
  assign f_arrdiv32_fs15_xor1 = f_arrdiv32_fs14_or0 ^ b[15];
  assign f_arrdiv32_fs15_not1 = ~b[15];
  assign f_arrdiv32_fs15_and1 = f_arrdiv32_fs15_not1 & f_arrdiv32_fs14_or0;
  assign f_arrdiv32_fs15_or0 = f_arrdiv32_fs15_and1 | b[15];
  assign f_arrdiv32_fs16_xor1 = f_arrdiv32_fs15_or0 ^ b[16];
  assign f_arrdiv32_fs16_not1 = ~b[16];
  assign f_arrdiv32_fs16_and1 = f_arrdiv32_fs16_not1 & f_arrdiv32_fs15_or0;
  assign f_arrdiv32_fs16_or0 = f_arrdiv32_fs16_and1 | b[16];
  assign f_arrdiv32_fs17_xor1 = f_arrdiv32_fs16_or0 ^ b[17];
  assign f_arrdiv32_fs17_not1 = ~b[17];
  assign f_arrdiv32_fs17_and1 = f_arrdiv32_fs17_not1 & f_arrdiv32_fs16_or0;
  assign f_arrdiv32_fs17_or0 = f_arrdiv32_fs17_and1 | b[17];
  assign f_arrdiv32_fs18_xor1 = f_arrdiv32_fs17_or0 ^ b[18];
  assign f_arrdiv32_fs18_not1 = ~b[18];
  assign f_arrdiv32_fs18_and1 = f_arrdiv32_fs18_not1 & f_arrdiv32_fs17_or0;
  assign f_arrdiv32_fs18_or0 = f_arrdiv32_fs18_and1 | b[18];
  assign f_arrdiv32_fs19_xor1 = f_arrdiv32_fs18_or0 ^ b[19];
  assign f_arrdiv32_fs19_not1 = ~b[19];
  assign f_arrdiv32_fs19_and1 = f_arrdiv32_fs19_not1 & f_arrdiv32_fs18_or0;
  assign f_arrdiv32_fs19_or0 = f_arrdiv32_fs19_and1 | b[19];
  assign f_arrdiv32_fs20_xor1 = f_arrdiv32_fs19_or0 ^ b[20];
  assign f_arrdiv32_fs20_not1 = ~b[20];
  assign f_arrdiv32_fs20_and1 = f_arrdiv32_fs20_not1 & f_arrdiv32_fs19_or0;
  assign f_arrdiv32_fs20_or0 = f_arrdiv32_fs20_and1 | b[20];
  assign f_arrdiv32_fs21_xor1 = f_arrdiv32_fs20_or0 ^ b[21];
  assign f_arrdiv32_fs21_not1 = ~b[21];
  assign f_arrdiv32_fs21_and1 = f_arrdiv32_fs21_not1 & f_arrdiv32_fs20_or0;
  assign f_arrdiv32_fs21_or0 = f_arrdiv32_fs21_and1 | b[21];
  assign f_arrdiv32_fs22_xor1 = f_arrdiv32_fs21_or0 ^ b[22];
  assign f_arrdiv32_fs22_not1 = ~b[22];
  assign f_arrdiv32_fs22_and1 = f_arrdiv32_fs22_not1 & f_arrdiv32_fs21_or0;
  assign f_arrdiv32_fs22_or0 = f_arrdiv32_fs22_and1 | b[22];
  assign f_arrdiv32_fs23_xor1 = f_arrdiv32_fs22_or0 ^ b[23];
  assign f_arrdiv32_fs23_not1 = ~b[23];
  assign f_arrdiv32_fs23_and1 = f_arrdiv32_fs23_not1 & f_arrdiv32_fs22_or0;
  assign f_arrdiv32_fs23_or0 = f_arrdiv32_fs23_and1 | b[23];
  assign f_arrdiv32_fs24_xor1 = f_arrdiv32_fs23_or0 ^ b[24];
  assign f_arrdiv32_fs24_not1 = ~b[24];
  assign f_arrdiv32_fs24_and1 = f_arrdiv32_fs24_not1 & f_arrdiv32_fs23_or0;
  assign f_arrdiv32_fs24_or0 = f_arrdiv32_fs24_and1 | b[24];
  assign f_arrdiv32_fs25_xor1 = f_arrdiv32_fs24_or0 ^ b[25];
  assign f_arrdiv32_fs25_not1 = ~b[25];
  assign f_arrdiv32_fs25_and1 = f_arrdiv32_fs25_not1 & f_arrdiv32_fs24_or0;
  assign f_arrdiv32_fs25_or0 = f_arrdiv32_fs25_and1 | b[25];
  assign f_arrdiv32_fs26_xor1 = f_arrdiv32_fs25_or0 ^ b[26];
  assign f_arrdiv32_fs26_not1 = ~b[26];
  assign f_arrdiv32_fs26_and1 = f_arrdiv32_fs26_not1 & f_arrdiv32_fs25_or0;
  assign f_arrdiv32_fs26_or0 = f_arrdiv32_fs26_and1 | b[26];
  assign f_arrdiv32_fs27_xor1 = f_arrdiv32_fs26_or0 ^ b[27];
  assign f_arrdiv32_fs27_not1 = ~b[27];
  assign f_arrdiv32_fs27_and1 = f_arrdiv32_fs27_not1 & f_arrdiv32_fs26_or0;
  assign f_arrdiv32_fs27_or0 = f_arrdiv32_fs27_and1 | b[27];
  assign f_arrdiv32_fs28_xor1 = f_arrdiv32_fs27_or0 ^ b[28];
  assign f_arrdiv32_fs28_not1 = ~b[28];
  assign f_arrdiv32_fs28_and1 = f_arrdiv32_fs28_not1 & f_arrdiv32_fs27_or0;
  assign f_arrdiv32_fs28_or0 = f_arrdiv32_fs28_and1 | b[28];
  assign f_arrdiv32_fs29_xor1 = f_arrdiv32_fs28_or0 ^ b[29];
  assign f_arrdiv32_fs29_not1 = ~b[29];
  assign f_arrdiv32_fs29_and1 = f_arrdiv32_fs29_not1 & f_arrdiv32_fs28_or0;
  assign f_arrdiv32_fs29_or0 = f_arrdiv32_fs29_and1 | b[29];
  assign f_arrdiv32_fs30_xor1 = f_arrdiv32_fs29_or0 ^ b[30];
  assign f_arrdiv32_fs30_not1 = ~b[30];
  assign f_arrdiv32_fs30_and1 = f_arrdiv32_fs30_not1 & f_arrdiv32_fs29_or0;
  assign f_arrdiv32_fs30_or0 = f_arrdiv32_fs30_and1 | b[30];
  assign f_arrdiv32_fs31_xor1 = f_arrdiv32_fs30_or0 ^ b[31];
  assign f_arrdiv32_fs31_not1 = ~b[31];
  assign f_arrdiv32_fs31_and1 = f_arrdiv32_fs31_not1 & f_arrdiv32_fs30_or0;
  assign f_arrdiv32_fs31_or0 = f_arrdiv32_fs31_and1 | b[31];
  assign f_arrdiv32_mux2to10_and0 = a[31] & f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to10_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to10_and1 = f_arrdiv32_fs0_xor0 & f_arrdiv32_mux2to10_not0;
  assign f_arrdiv32_mux2to10_xor0 = f_arrdiv32_mux2to10_and0 ^ f_arrdiv32_mux2to10_and1;
  assign f_arrdiv32_mux2to11_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to11_and1 = f_arrdiv32_fs1_xor1 & f_arrdiv32_mux2to11_not0;
  assign f_arrdiv32_mux2to12_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to12_and1 = f_arrdiv32_fs2_xor1 & f_arrdiv32_mux2to12_not0;
  assign f_arrdiv32_mux2to13_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to13_and1 = f_arrdiv32_fs3_xor1 & f_arrdiv32_mux2to13_not0;
  assign f_arrdiv32_mux2to14_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to14_and1 = f_arrdiv32_fs4_xor1 & f_arrdiv32_mux2to14_not0;
  assign f_arrdiv32_mux2to15_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to15_and1 = f_arrdiv32_fs5_xor1 & f_arrdiv32_mux2to15_not0;
  assign f_arrdiv32_mux2to16_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to16_and1 = f_arrdiv32_fs6_xor1 & f_arrdiv32_mux2to16_not0;
  assign f_arrdiv32_mux2to17_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to17_and1 = f_arrdiv32_fs7_xor1 & f_arrdiv32_mux2to17_not0;
  assign f_arrdiv32_mux2to18_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to18_and1 = f_arrdiv32_fs8_xor1 & f_arrdiv32_mux2to18_not0;
  assign f_arrdiv32_mux2to19_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to19_and1 = f_arrdiv32_fs9_xor1 & f_arrdiv32_mux2to19_not0;
  assign f_arrdiv32_mux2to110_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to110_and1 = f_arrdiv32_fs10_xor1 & f_arrdiv32_mux2to110_not0;
  assign f_arrdiv32_mux2to111_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to111_and1 = f_arrdiv32_fs11_xor1 & f_arrdiv32_mux2to111_not0;
  assign f_arrdiv32_mux2to112_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to112_and1 = f_arrdiv32_fs12_xor1 & f_arrdiv32_mux2to112_not0;
  assign f_arrdiv32_mux2to113_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to113_and1 = f_arrdiv32_fs13_xor1 & f_arrdiv32_mux2to113_not0;
  assign f_arrdiv32_mux2to114_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to114_and1 = f_arrdiv32_fs14_xor1 & f_arrdiv32_mux2to114_not0;
  assign f_arrdiv32_mux2to115_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to115_and1 = f_arrdiv32_fs15_xor1 & f_arrdiv32_mux2to115_not0;
  assign f_arrdiv32_mux2to116_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to116_and1 = f_arrdiv32_fs16_xor1 & f_arrdiv32_mux2to116_not0;
  assign f_arrdiv32_mux2to117_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to117_and1 = f_arrdiv32_fs17_xor1 & f_arrdiv32_mux2to117_not0;
  assign f_arrdiv32_mux2to118_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to118_and1 = f_arrdiv32_fs18_xor1 & f_arrdiv32_mux2to118_not0;
  assign f_arrdiv32_mux2to119_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to119_and1 = f_arrdiv32_fs19_xor1 & f_arrdiv32_mux2to119_not0;
  assign f_arrdiv32_mux2to120_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to120_and1 = f_arrdiv32_fs20_xor1 & f_arrdiv32_mux2to120_not0;
  assign f_arrdiv32_mux2to121_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to121_and1 = f_arrdiv32_fs21_xor1 & f_arrdiv32_mux2to121_not0;
  assign f_arrdiv32_mux2to122_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to122_and1 = f_arrdiv32_fs22_xor1 & f_arrdiv32_mux2to122_not0;
  assign f_arrdiv32_mux2to123_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to123_and1 = f_arrdiv32_fs23_xor1 & f_arrdiv32_mux2to123_not0;
  assign f_arrdiv32_mux2to124_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to124_and1 = f_arrdiv32_fs24_xor1 & f_arrdiv32_mux2to124_not0;
  assign f_arrdiv32_mux2to125_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to125_and1 = f_arrdiv32_fs25_xor1 & f_arrdiv32_mux2to125_not0;
  assign f_arrdiv32_mux2to126_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to126_and1 = f_arrdiv32_fs26_xor1 & f_arrdiv32_mux2to126_not0;
  assign f_arrdiv32_mux2to127_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to127_and1 = f_arrdiv32_fs27_xor1 & f_arrdiv32_mux2to127_not0;
  assign f_arrdiv32_mux2to128_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to128_and1 = f_arrdiv32_fs28_xor1 & f_arrdiv32_mux2to128_not0;
  assign f_arrdiv32_mux2to129_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to129_and1 = f_arrdiv32_fs29_xor1 & f_arrdiv32_mux2to129_not0;
  assign f_arrdiv32_mux2to130_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_mux2to130_and1 = f_arrdiv32_fs30_xor1 & f_arrdiv32_mux2to130_not0;
  assign f_arrdiv32_not0 = ~f_arrdiv32_fs31_or0;
  assign f_arrdiv32_fs32_xor0 = a[30] ^ b[0];
  assign f_arrdiv32_fs32_not0 = ~a[30];
  assign f_arrdiv32_fs32_and0 = f_arrdiv32_fs32_not0 & b[0];
  assign f_arrdiv32_fs32_not1 = ~f_arrdiv32_fs32_xor0;
  assign f_arrdiv32_fs33_xor0 = f_arrdiv32_mux2to10_xor0 ^ b[1];
  assign f_arrdiv32_fs33_not0 = ~f_arrdiv32_mux2to10_xor0;
  assign f_arrdiv32_fs33_and0 = f_arrdiv32_fs33_not0 & b[1];
  assign f_arrdiv32_fs33_xor1 = f_arrdiv32_fs32_and0 ^ f_arrdiv32_fs33_xor0;
  assign f_arrdiv32_fs33_not1 = ~f_arrdiv32_fs33_xor0;
  assign f_arrdiv32_fs33_and1 = f_arrdiv32_fs33_not1 & f_arrdiv32_fs32_and0;
  assign f_arrdiv32_fs33_or0 = f_arrdiv32_fs33_and1 | f_arrdiv32_fs33_and0;
  assign f_arrdiv32_fs34_xor0 = f_arrdiv32_mux2to11_and1 ^ b[2];
  assign f_arrdiv32_fs34_not0 = ~f_arrdiv32_mux2to11_and1;
  assign f_arrdiv32_fs34_and0 = f_arrdiv32_fs34_not0 & b[2];
  assign f_arrdiv32_fs34_xor1 = f_arrdiv32_fs33_or0 ^ f_arrdiv32_fs34_xor0;
  assign f_arrdiv32_fs34_not1 = ~f_arrdiv32_fs34_xor0;
  assign f_arrdiv32_fs34_and1 = f_arrdiv32_fs34_not1 & f_arrdiv32_fs33_or0;
  assign f_arrdiv32_fs34_or0 = f_arrdiv32_fs34_and1 | f_arrdiv32_fs34_and0;
  assign f_arrdiv32_fs35_xor0 = f_arrdiv32_mux2to12_and1 ^ b[3];
  assign f_arrdiv32_fs35_not0 = ~f_arrdiv32_mux2to12_and1;
  assign f_arrdiv32_fs35_and0 = f_arrdiv32_fs35_not0 & b[3];
  assign f_arrdiv32_fs35_xor1 = f_arrdiv32_fs34_or0 ^ f_arrdiv32_fs35_xor0;
  assign f_arrdiv32_fs35_not1 = ~f_arrdiv32_fs35_xor0;
  assign f_arrdiv32_fs35_and1 = f_arrdiv32_fs35_not1 & f_arrdiv32_fs34_or0;
  assign f_arrdiv32_fs35_or0 = f_arrdiv32_fs35_and1 | f_arrdiv32_fs35_and0;
  assign f_arrdiv32_fs36_xor0 = f_arrdiv32_mux2to13_and1 ^ b[4];
  assign f_arrdiv32_fs36_not0 = ~f_arrdiv32_mux2to13_and1;
  assign f_arrdiv32_fs36_and0 = f_arrdiv32_fs36_not0 & b[4];
  assign f_arrdiv32_fs36_xor1 = f_arrdiv32_fs35_or0 ^ f_arrdiv32_fs36_xor0;
  assign f_arrdiv32_fs36_not1 = ~f_arrdiv32_fs36_xor0;
  assign f_arrdiv32_fs36_and1 = f_arrdiv32_fs36_not1 & f_arrdiv32_fs35_or0;
  assign f_arrdiv32_fs36_or0 = f_arrdiv32_fs36_and1 | f_arrdiv32_fs36_and0;
  assign f_arrdiv32_fs37_xor0 = f_arrdiv32_mux2to14_and1 ^ b[5];
  assign f_arrdiv32_fs37_not0 = ~f_arrdiv32_mux2to14_and1;
  assign f_arrdiv32_fs37_and0 = f_arrdiv32_fs37_not0 & b[5];
  assign f_arrdiv32_fs37_xor1 = f_arrdiv32_fs36_or0 ^ f_arrdiv32_fs37_xor0;
  assign f_arrdiv32_fs37_not1 = ~f_arrdiv32_fs37_xor0;
  assign f_arrdiv32_fs37_and1 = f_arrdiv32_fs37_not1 & f_arrdiv32_fs36_or0;
  assign f_arrdiv32_fs37_or0 = f_arrdiv32_fs37_and1 | f_arrdiv32_fs37_and0;
  assign f_arrdiv32_fs38_xor0 = f_arrdiv32_mux2to15_and1 ^ b[6];
  assign f_arrdiv32_fs38_not0 = ~f_arrdiv32_mux2to15_and1;
  assign f_arrdiv32_fs38_and0 = f_arrdiv32_fs38_not0 & b[6];
  assign f_arrdiv32_fs38_xor1 = f_arrdiv32_fs37_or0 ^ f_arrdiv32_fs38_xor0;
  assign f_arrdiv32_fs38_not1 = ~f_arrdiv32_fs38_xor0;
  assign f_arrdiv32_fs38_and1 = f_arrdiv32_fs38_not1 & f_arrdiv32_fs37_or0;
  assign f_arrdiv32_fs38_or0 = f_arrdiv32_fs38_and1 | f_arrdiv32_fs38_and0;
  assign f_arrdiv32_fs39_xor0 = f_arrdiv32_mux2to16_and1 ^ b[7];
  assign f_arrdiv32_fs39_not0 = ~f_arrdiv32_mux2to16_and1;
  assign f_arrdiv32_fs39_and0 = f_arrdiv32_fs39_not0 & b[7];
  assign f_arrdiv32_fs39_xor1 = f_arrdiv32_fs38_or0 ^ f_arrdiv32_fs39_xor0;
  assign f_arrdiv32_fs39_not1 = ~f_arrdiv32_fs39_xor0;
  assign f_arrdiv32_fs39_and1 = f_arrdiv32_fs39_not1 & f_arrdiv32_fs38_or0;
  assign f_arrdiv32_fs39_or0 = f_arrdiv32_fs39_and1 | f_arrdiv32_fs39_and0;
  assign f_arrdiv32_fs40_xor0 = f_arrdiv32_mux2to17_and1 ^ b[8];
  assign f_arrdiv32_fs40_not0 = ~f_arrdiv32_mux2to17_and1;
  assign f_arrdiv32_fs40_and0 = f_arrdiv32_fs40_not0 & b[8];
  assign f_arrdiv32_fs40_xor1 = f_arrdiv32_fs39_or0 ^ f_arrdiv32_fs40_xor0;
  assign f_arrdiv32_fs40_not1 = ~f_arrdiv32_fs40_xor0;
  assign f_arrdiv32_fs40_and1 = f_arrdiv32_fs40_not1 & f_arrdiv32_fs39_or0;
  assign f_arrdiv32_fs40_or0 = f_arrdiv32_fs40_and1 | f_arrdiv32_fs40_and0;
  assign f_arrdiv32_fs41_xor0 = f_arrdiv32_mux2to18_and1 ^ b[9];
  assign f_arrdiv32_fs41_not0 = ~f_arrdiv32_mux2to18_and1;
  assign f_arrdiv32_fs41_and0 = f_arrdiv32_fs41_not0 & b[9];
  assign f_arrdiv32_fs41_xor1 = f_arrdiv32_fs40_or0 ^ f_arrdiv32_fs41_xor0;
  assign f_arrdiv32_fs41_not1 = ~f_arrdiv32_fs41_xor0;
  assign f_arrdiv32_fs41_and1 = f_arrdiv32_fs41_not1 & f_arrdiv32_fs40_or0;
  assign f_arrdiv32_fs41_or0 = f_arrdiv32_fs41_and1 | f_arrdiv32_fs41_and0;
  assign f_arrdiv32_fs42_xor0 = f_arrdiv32_mux2to19_and1 ^ b[10];
  assign f_arrdiv32_fs42_not0 = ~f_arrdiv32_mux2to19_and1;
  assign f_arrdiv32_fs42_and0 = f_arrdiv32_fs42_not0 & b[10];
  assign f_arrdiv32_fs42_xor1 = f_arrdiv32_fs41_or0 ^ f_arrdiv32_fs42_xor0;
  assign f_arrdiv32_fs42_not1 = ~f_arrdiv32_fs42_xor0;
  assign f_arrdiv32_fs42_and1 = f_arrdiv32_fs42_not1 & f_arrdiv32_fs41_or0;
  assign f_arrdiv32_fs42_or0 = f_arrdiv32_fs42_and1 | f_arrdiv32_fs42_and0;
  assign f_arrdiv32_fs43_xor0 = f_arrdiv32_mux2to110_and1 ^ b[11];
  assign f_arrdiv32_fs43_not0 = ~f_arrdiv32_mux2to110_and1;
  assign f_arrdiv32_fs43_and0 = f_arrdiv32_fs43_not0 & b[11];
  assign f_arrdiv32_fs43_xor1 = f_arrdiv32_fs42_or0 ^ f_arrdiv32_fs43_xor0;
  assign f_arrdiv32_fs43_not1 = ~f_arrdiv32_fs43_xor0;
  assign f_arrdiv32_fs43_and1 = f_arrdiv32_fs43_not1 & f_arrdiv32_fs42_or0;
  assign f_arrdiv32_fs43_or0 = f_arrdiv32_fs43_and1 | f_arrdiv32_fs43_and0;
  assign f_arrdiv32_fs44_xor0 = f_arrdiv32_mux2to111_and1 ^ b[12];
  assign f_arrdiv32_fs44_not0 = ~f_arrdiv32_mux2to111_and1;
  assign f_arrdiv32_fs44_and0 = f_arrdiv32_fs44_not0 & b[12];
  assign f_arrdiv32_fs44_xor1 = f_arrdiv32_fs43_or0 ^ f_arrdiv32_fs44_xor0;
  assign f_arrdiv32_fs44_not1 = ~f_arrdiv32_fs44_xor0;
  assign f_arrdiv32_fs44_and1 = f_arrdiv32_fs44_not1 & f_arrdiv32_fs43_or0;
  assign f_arrdiv32_fs44_or0 = f_arrdiv32_fs44_and1 | f_arrdiv32_fs44_and0;
  assign f_arrdiv32_fs45_xor0 = f_arrdiv32_mux2to112_and1 ^ b[13];
  assign f_arrdiv32_fs45_not0 = ~f_arrdiv32_mux2to112_and1;
  assign f_arrdiv32_fs45_and0 = f_arrdiv32_fs45_not0 & b[13];
  assign f_arrdiv32_fs45_xor1 = f_arrdiv32_fs44_or0 ^ f_arrdiv32_fs45_xor0;
  assign f_arrdiv32_fs45_not1 = ~f_arrdiv32_fs45_xor0;
  assign f_arrdiv32_fs45_and1 = f_arrdiv32_fs45_not1 & f_arrdiv32_fs44_or0;
  assign f_arrdiv32_fs45_or0 = f_arrdiv32_fs45_and1 | f_arrdiv32_fs45_and0;
  assign f_arrdiv32_fs46_xor0 = f_arrdiv32_mux2to113_and1 ^ b[14];
  assign f_arrdiv32_fs46_not0 = ~f_arrdiv32_mux2to113_and1;
  assign f_arrdiv32_fs46_and0 = f_arrdiv32_fs46_not0 & b[14];
  assign f_arrdiv32_fs46_xor1 = f_arrdiv32_fs45_or0 ^ f_arrdiv32_fs46_xor0;
  assign f_arrdiv32_fs46_not1 = ~f_arrdiv32_fs46_xor0;
  assign f_arrdiv32_fs46_and1 = f_arrdiv32_fs46_not1 & f_arrdiv32_fs45_or0;
  assign f_arrdiv32_fs46_or0 = f_arrdiv32_fs46_and1 | f_arrdiv32_fs46_and0;
  assign f_arrdiv32_fs47_xor0 = f_arrdiv32_mux2to114_and1 ^ b[15];
  assign f_arrdiv32_fs47_not0 = ~f_arrdiv32_mux2to114_and1;
  assign f_arrdiv32_fs47_and0 = f_arrdiv32_fs47_not0 & b[15];
  assign f_arrdiv32_fs47_xor1 = f_arrdiv32_fs46_or0 ^ f_arrdiv32_fs47_xor0;
  assign f_arrdiv32_fs47_not1 = ~f_arrdiv32_fs47_xor0;
  assign f_arrdiv32_fs47_and1 = f_arrdiv32_fs47_not1 & f_arrdiv32_fs46_or0;
  assign f_arrdiv32_fs47_or0 = f_arrdiv32_fs47_and1 | f_arrdiv32_fs47_and0;
  assign f_arrdiv32_fs48_xor0 = f_arrdiv32_mux2to115_and1 ^ b[16];
  assign f_arrdiv32_fs48_not0 = ~f_arrdiv32_mux2to115_and1;
  assign f_arrdiv32_fs48_and0 = f_arrdiv32_fs48_not0 & b[16];
  assign f_arrdiv32_fs48_xor1 = f_arrdiv32_fs47_or0 ^ f_arrdiv32_fs48_xor0;
  assign f_arrdiv32_fs48_not1 = ~f_arrdiv32_fs48_xor0;
  assign f_arrdiv32_fs48_and1 = f_arrdiv32_fs48_not1 & f_arrdiv32_fs47_or0;
  assign f_arrdiv32_fs48_or0 = f_arrdiv32_fs48_and1 | f_arrdiv32_fs48_and0;
  assign f_arrdiv32_fs49_xor0 = f_arrdiv32_mux2to116_and1 ^ b[17];
  assign f_arrdiv32_fs49_not0 = ~f_arrdiv32_mux2to116_and1;
  assign f_arrdiv32_fs49_and0 = f_arrdiv32_fs49_not0 & b[17];
  assign f_arrdiv32_fs49_xor1 = f_arrdiv32_fs48_or0 ^ f_arrdiv32_fs49_xor0;
  assign f_arrdiv32_fs49_not1 = ~f_arrdiv32_fs49_xor0;
  assign f_arrdiv32_fs49_and1 = f_arrdiv32_fs49_not1 & f_arrdiv32_fs48_or0;
  assign f_arrdiv32_fs49_or0 = f_arrdiv32_fs49_and1 | f_arrdiv32_fs49_and0;
  assign f_arrdiv32_fs50_xor0 = f_arrdiv32_mux2to117_and1 ^ b[18];
  assign f_arrdiv32_fs50_not0 = ~f_arrdiv32_mux2to117_and1;
  assign f_arrdiv32_fs50_and0 = f_arrdiv32_fs50_not0 & b[18];
  assign f_arrdiv32_fs50_xor1 = f_arrdiv32_fs49_or0 ^ f_arrdiv32_fs50_xor0;
  assign f_arrdiv32_fs50_not1 = ~f_arrdiv32_fs50_xor0;
  assign f_arrdiv32_fs50_and1 = f_arrdiv32_fs50_not1 & f_arrdiv32_fs49_or0;
  assign f_arrdiv32_fs50_or0 = f_arrdiv32_fs50_and1 | f_arrdiv32_fs50_and0;
  assign f_arrdiv32_fs51_xor0 = f_arrdiv32_mux2to118_and1 ^ b[19];
  assign f_arrdiv32_fs51_not0 = ~f_arrdiv32_mux2to118_and1;
  assign f_arrdiv32_fs51_and0 = f_arrdiv32_fs51_not0 & b[19];
  assign f_arrdiv32_fs51_xor1 = f_arrdiv32_fs50_or0 ^ f_arrdiv32_fs51_xor0;
  assign f_arrdiv32_fs51_not1 = ~f_arrdiv32_fs51_xor0;
  assign f_arrdiv32_fs51_and1 = f_arrdiv32_fs51_not1 & f_arrdiv32_fs50_or0;
  assign f_arrdiv32_fs51_or0 = f_arrdiv32_fs51_and1 | f_arrdiv32_fs51_and0;
  assign f_arrdiv32_fs52_xor0 = f_arrdiv32_mux2to119_and1 ^ b[20];
  assign f_arrdiv32_fs52_not0 = ~f_arrdiv32_mux2to119_and1;
  assign f_arrdiv32_fs52_and0 = f_arrdiv32_fs52_not0 & b[20];
  assign f_arrdiv32_fs52_xor1 = f_arrdiv32_fs51_or0 ^ f_arrdiv32_fs52_xor0;
  assign f_arrdiv32_fs52_not1 = ~f_arrdiv32_fs52_xor0;
  assign f_arrdiv32_fs52_and1 = f_arrdiv32_fs52_not1 & f_arrdiv32_fs51_or0;
  assign f_arrdiv32_fs52_or0 = f_arrdiv32_fs52_and1 | f_arrdiv32_fs52_and0;
  assign f_arrdiv32_fs53_xor0 = f_arrdiv32_mux2to120_and1 ^ b[21];
  assign f_arrdiv32_fs53_not0 = ~f_arrdiv32_mux2to120_and1;
  assign f_arrdiv32_fs53_and0 = f_arrdiv32_fs53_not0 & b[21];
  assign f_arrdiv32_fs53_xor1 = f_arrdiv32_fs52_or0 ^ f_arrdiv32_fs53_xor0;
  assign f_arrdiv32_fs53_not1 = ~f_arrdiv32_fs53_xor0;
  assign f_arrdiv32_fs53_and1 = f_arrdiv32_fs53_not1 & f_arrdiv32_fs52_or0;
  assign f_arrdiv32_fs53_or0 = f_arrdiv32_fs53_and1 | f_arrdiv32_fs53_and0;
  assign f_arrdiv32_fs54_xor0 = f_arrdiv32_mux2to121_and1 ^ b[22];
  assign f_arrdiv32_fs54_not0 = ~f_arrdiv32_mux2to121_and1;
  assign f_arrdiv32_fs54_and0 = f_arrdiv32_fs54_not0 & b[22];
  assign f_arrdiv32_fs54_xor1 = f_arrdiv32_fs53_or0 ^ f_arrdiv32_fs54_xor0;
  assign f_arrdiv32_fs54_not1 = ~f_arrdiv32_fs54_xor0;
  assign f_arrdiv32_fs54_and1 = f_arrdiv32_fs54_not1 & f_arrdiv32_fs53_or0;
  assign f_arrdiv32_fs54_or0 = f_arrdiv32_fs54_and1 | f_arrdiv32_fs54_and0;
  assign f_arrdiv32_fs55_xor0 = f_arrdiv32_mux2to122_and1 ^ b[23];
  assign f_arrdiv32_fs55_not0 = ~f_arrdiv32_mux2to122_and1;
  assign f_arrdiv32_fs55_and0 = f_arrdiv32_fs55_not0 & b[23];
  assign f_arrdiv32_fs55_xor1 = f_arrdiv32_fs54_or0 ^ f_arrdiv32_fs55_xor0;
  assign f_arrdiv32_fs55_not1 = ~f_arrdiv32_fs55_xor0;
  assign f_arrdiv32_fs55_and1 = f_arrdiv32_fs55_not1 & f_arrdiv32_fs54_or0;
  assign f_arrdiv32_fs55_or0 = f_arrdiv32_fs55_and1 | f_arrdiv32_fs55_and0;
  assign f_arrdiv32_fs56_xor0 = f_arrdiv32_mux2to123_and1 ^ b[24];
  assign f_arrdiv32_fs56_not0 = ~f_arrdiv32_mux2to123_and1;
  assign f_arrdiv32_fs56_and0 = f_arrdiv32_fs56_not0 & b[24];
  assign f_arrdiv32_fs56_xor1 = f_arrdiv32_fs55_or0 ^ f_arrdiv32_fs56_xor0;
  assign f_arrdiv32_fs56_not1 = ~f_arrdiv32_fs56_xor0;
  assign f_arrdiv32_fs56_and1 = f_arrdiv32_fs56_not1 & f_arrdiv32_fs55_or0;
  assign f_arrdiv32_fs56_or0 = f_arrdiv32_fs56_and1 | f_arrdiv32_fs56_and0;
  assign f_arrdiv32_fs57_xor0 = f_arrdiv32_mux2to124_and1 ^ b[25];
  assign f_arrdiv32_fs57_not0 = ~f_arrdiv32_mux2to124_and1;
  assign f_arrdiv32_fs57_and0 = f_arrdiv32_fs57_not0 & b[25];
  assign f_arrdiv32_fs57_xor1 = f_arrdiv32_fs56_or0 ^ f_arrdiv32_fs57_xor0;
  assign f_arrdiv32_fs57_not1 = ~f_arrdiv32_fs57_xor0;
  assign f_arrdiv32_fs57_and1 = f_arrdiv32_fs57_not1 & f_arrdiv32_fs56_or0;
  assign f_arrdiv32_fs57_or0 = f_arrdiv32_fs57_and1 | f_arrdiv32_fs57_and0;
  assign f_arrdiv32_fs58_xor0 = f_arrdiv32_mux2to125_and1 ^ b[26];
  assign f_arrdiv32_fs58_not0 = ~f_arrdiv32_mux2to125_and1;
  assign f_arrdiv32_fs58_and0 = f_arrdiv32_fs58_not0 & b[26];
  assign f_arrdiv32_fs58_xor1 = f_arrdiv32_fs57_or0 ^ f_arrdiv32_fs58_xor0;
  assign f_arrdiv32_fs58_not1 = ~f_arrdiv32_fs58_xor0;
  assign f_arrdiv32_fs58_and1 = f_arrdiv32_fs58_not1 & f_arrdiv32_fs57_or0;
  assign f_arrdiv32_fs58_or0 = f_arrdiv32_fs58_and1 | f_arrdiv32_fs58_and0;
  assign f_arrdiv32_fs59_xor0 = f_arrdiv32_mux2to126_and1 ^ b[27];
  assign f_arrdiv32_fs59_not0 = ~f_arrdiv32_mux2to126_and1;
  assign f_arrdiv32_fs59_and0 = f_arrdiv32_fs59_not0 & b[27];
  assign f_arrdiv32_fs59_xor1 = f_arrdiv32_fs58_or0 ^ f_arrdiv32_fs59_xor0;
  assign f_arrdiv32_fs59_not1 = ~f_arrdiv32_fs59_xor0;
  assign f_arrdiv32_fs59_and1 = f_arrdiv32_fs59_not1 & f_arrdiv32_fs58_or0;
  assign f_arrdiv32_fs59_or0 = f_arrdiv32_fs59_and1 | f_arrdiv32_fs59_and0;
  assign f_arrdiv32_fs60_xor0 = f_arrdiv32_mux2to127_and1 ^ b[28];
  assign f_arrdiv32_fs60_not0 = ~f_arrdiv32_mux2to127_and1;
  assign f_arrdiv32_fs60_and0 = f_arrdiv32_fs60_not0 & b[28];
  assign f_arrdiv32_fs60_xor1 = f_arrdiv32_fs59_or0 ^ f_arrdiv32_fs60_xor0;
  assign f_arrdiv32_fs60_not1 = ~f_arrdiv32_fs60_xor0;
  assign f_arrdiv32_fs60_and1 = f_arrdiv32_fs60_not1 & f_arrdiv32_fs59_or0;
  assign f_arrdiv32_fs60_or0 = f_arrdiv32_fs60_and1 | f_arrdiv32_fs60_and0;
  assign f_arrdiv32_fs61_xor0 = f_arrdiv32_mux2to128_and1 ^ b[29];
  assign f_arrdiv32_fs61_not0 = ~f_arrdiv32_mux2to128_and1;
  assign f_arrdiv32_fs61_and0 = f_arrdiv32_fs61_not0 & b[29];
  assign f_arrdiv32_fs61_xor1 = f_arrdiv32_fs60_or0 ^ f_arrdiv32_fs61_xor0;
  assign f_arrdiv32_fs61_not1 = ~f_arrdiv32_fs61_xor0;
  assign f_arrdiv32_fs61_and1 = f_arrdiv32_fs61_not1 & f_arrdiv32_fs60_or0;
  assign f_arrdiv32_fs61_or0 = f_arrdiv32_fs61_and1 | f_arrdiv32_fs61_and0;
  assign f_arrdiv32_fs62_xor0 = f_arrdiv32_mux2to129_and1 ^ b[30];
  assign f_arrdiv32_fs62_not0 = ~f_arrdiv32_mux2to129_and1;
  assign f_arrdiv32_fs62_and0 = f_arrdiv32_fs62_not0 & b[30];
  assign f_arrdiv32_fs62_xor1 = f_arrdiv32_fs61_or0 ^ f_arrdiv32_fs62_xor0;
  assign f_arrdiv32_fs62_not1 = ~f_arrdiv32_fs62_xor0;
  assign f_arrdiv32_fs62_and1 = f_arrdiv32_fs62_not1 & f_arrdiv32_fs61_or0;
  assign f_arrdiv32_fs62_or0 = f_arrdiv32_fs62_and1 | f_arrdiv32_fs62_and0;
  assign f_arrdiv32_fs63_xor0 = f_arrdiv32_mux2to130_and1 ^ b[31];
  assign f_arrdiv32_fs63_not0 = ~f_arrdiv32_mux2to130_and1;
  assign f_arrdiv32_fs63_and0 = f_arrdiv32_fs63_not0 & b[31];
  assign f_arrdiv32_fs63_xor1 = f_arrdiv32_fs62_or0 ^ f_arrdiv32_fs63_xor0;
  assign f_arrdiv32_fs63_not1 = ~f_arrdiv32_fs63_xor0;
  assign f_arrdiv32_fs63_and1 = f_arrdiv32_fs63_not1 & f_arrdiv32_fs62_or0;
  assign f_arrdiv32_fs63_or0 = f_arrdiv32_fs63_and1 | f_arrdiv32_fs63_and0;
  assign f_arrdiv32_mux2to131_and0 = a[30] & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to131_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to131_and1 = f_arrdiv32_fs32_xor0 & f_arrdiv32_mux2to131_not0;
  assign f_arrdiv32_mux2to131_xor0 = f_arrdiv32_mux2to131_and0 ^ f_arrdiv32_mux2to131_and1;
  assign f_arrdiv32_mux2to132_and0 = f_arrdiv32_mux2to10_xor0 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to132_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to132_and1 = f_arrdiv32_fs33_xor1 & f_arrdiv32_mux2to132_not0;
  assign f_arrdiv32_mux2to132_xor0 = f_arrdiv32_mux2to132_and0 ^ f_arrdiv32_mux2to132_and1;
  assign f_arrdiv32_mux2to133_and0 = f_arrdiv32_mux2to11_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to133_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to133_and1 = f_arrdiv32_fs34_xor1 & f_arrdiv32_mux2to133_not0;
  assign f_arrdiv32_mux2to133_xor0 = f_arrdiv32_mux2to133_and0 ^ f_arrdiv32_mux2to133_and1;
  assign f_arrdiv32_mux2to134_and0 = f_arrdiv32_mux2to12_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to134_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to134_and1 = f_arrdiv32_fs35_xor1 & f_arrdiv32_mux2to134_not0;
  assign f_arrdiv32_mux2to134_xor0 = f_arrdiv32_mux2to134_and0 ^ f_arrdiv32_mux2to134_and1;
  assign f_arrdiv32_mux2to135_and0 = f_arrdiv32_mux2to13_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to135_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to135_and1 = f_arrdiv32_fs36_xor1 & f_arrdiv32_mux2to135_not0;
  assign f_arrdiv32_mux2to135_xor0 = f_arrdiv32_mux2to135_and0 ^ f_arrdiv32_mux2to135_and1;
  assign f_arrdiv32_mux2to136_and0 = f_arrdiv32_mux2to14_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to136_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to136_and1 = f_arrdiv32_fs37_xor1 & f_arrdiv32_mux2to136_not0;
  assign f_arrdiv32_mux2to136_xor0 = f_arrdiv32_mux2to136_and0 ^ f_arrdiv32_mux2to136_and1;
  assign f_arrdiv32_mux2to137_and0 = f_arrdiv32_mux2to15_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to137_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to137_and1 = f_arrdiv32_fs38_xor1 & f_arrdiv32_mux2to137_not0;
  assign f_arrdiv32_mux2to137_xor0 = f_arrdiv32_mux2to137_and0 ^ f_arrdiv32_mux2to137_and1;
  assign f_arrdiv32_mux2to138_and0 = f_arrdiv32_mux2to16_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to138_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to138_and1 = f_arrdiv32_fs39_xor1 & f_arrdiv32_mux2to138_not0;
  assign f_arrdiv32_mux2to138_xor0 = f_arrdiv32_mux2to138_and0 ^ f_arrdiv32_mux2to138_and1;
  assign f_arrdiv32_mux2to139_and0 = f_arrdiv32_mux2to17_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to139_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to139_and1 = f_arrdiv32_fs40_xor1 & f_arrdiv32_mux2to139_not0;
  assign f_arrdiv32_mux2to139_xor0 = f_arrdiv32_mux2to139_and0 ^ f_arrdiv32_mux2to139_and1;
  assign f_arrdiv32_mux2to140_and0 = f_arrdiv32_mux2to18_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to140_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to140_and1 = f_arrdiv32_fs41_xor1 & f_arrdiv32_mux2to140_not0;
  assign f_arrdiv32_mux2to140_xor0 = f_arrdiv32_mux2to140_and0 ^ f_arrdiv32_mux2to140_and1;
  assign f_arrdiv32_mux2to141_and0 = f_arrdiv32_mux2to19_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to141_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to141_and1 = f_arrdiv32_fs42_xor1 & f_arrdiv32_mux2to141_not0;
  assign f_arrdiv32_mux2to141_xor0 = f_arrdiv32_mux2to141_and0 ^ f_arrdiv32_mux2to141_and1;
  assign f_arrdiv32_mux2to142_and0 = f_arrdiv32_mux2to110_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to142_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to142_and1 = f_arrdiv32_fs43_xor1 & f_arrdiv32_mux2to142_not0;
  assign f_arrdiv32_mux2to142_xor0 = f_arrdiv32_mux2to142_and0 ^ f_arrdiv32_mux2to142_and1;
  assign f_arrdiv32_mux2to143_and0 = f_arrdiv32_mux2to111_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to143_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to143_and1 = f_arrdiv32_fs44_xor1 & f_arrdiv32_mux2to143_not0;
  assign f_arrdiv32_mux2to143_xor0 = f_arrdiv32_mux2to143_and0 ^ f_arrdiv32_mux2to143_and1;
  assign f_arrdiv32_mux2to144_and0 = f_arrdiv32_mux2to112_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to144_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to144_and1 = f_arrdiv32_fs45_xor1 & f_arrdiv32_mux2to144_not0;
  assign f_arrdiv32_mux2to144_xor0 = f_arrdiv32_mux2to144_and0 ^ f_arrdiv32_mux2to144_and1;
  assign f_arrdiv32_mux2to145_and0 = f_arrdiv32_mux2to113_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to145_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to145_and1 = f_arrdiv32_fs46_xor1 & f_arrdiv32_mux2to145_not0;
  assign f_arrdiv32_mux2to145_xor0 = f_arrdiv32_mux2to145_and0 ^ f_arrdiv32_mux2to145_and1;
  assign f_arrdiv32_mux2to146_and0 = f_arrdiv32_mux2to114_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to146_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to146_and1 = f_arrdiv32_fs47_xor1 & f_arrdiv32_mux2to146_not0;
  assign f_arrdiv32_mux2to146_xor0 = f_arrdiv32_mux2to146_and0 ^ f_arrdiv32_mux2to146_and1;
  assign f_arrdiv32_mux2to147_and0 = f_arrdiv32_mux2to115_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to147_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to147_and1 = f_arrdiv32_fs48_xor1 & f_arrdiv32_mux2to147_not0;
  assign f_arrdiv32_mux2to147_xor0 = f_arrdiv32_mux2to147_and0 ^ f_arrdiv32_mux2to147_and1;
  assign f_arrdiv32_mux2to148_and0 = f_arrdiv32_mux2to116_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to148_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to148_and1 = f_arrdiv32_fs49_xor1 & f_arrdiv32_mux2to148_not0;
  assign f_arrdiv32_mux2to148_xor0 = f_arrdiv32_mux2to148_and0 ^ f_arrdiv32_mux2to148_and1;
  assign f_arrdiv32_mux2to149_and0 = f_arrdiv32_mux2to117_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to149_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to149_and1 = f_arrdiv32_fs50_xor1 & f_arrdiv32_mux2to149_not0;
  assign f_arrdiv32_mux2to149_xor0 = f_arrdiv32_mux2to149_and0 ^ f_arrdiv32_mux2to149_and1;
  assign f_arrdiv32_mux2to150_and0 = f_arrdiv32_mux2to118_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to150_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to150_and1 = f_arrdiv32_fs51_xor1 & f_arrdiv32_mux2to150_not0;
  assign f_arrdiv32_mux2to150_xor0 = f_arrdiv32_mux2to150_and0 ^ f_arrdiv32_mux2to150_and1;
  assign f_arrdiv32_mux2to151_and0 = f_arrdiv32_mux2to119_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to151_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to151_and1 = f_arrdiv32_fs52_xor1 & f_arrdiv32_mux2to151_not0;
  assign f_arrdiv32_mux2to151_xor0 = f_arrdiv32_mux2to151_and0 ^ f_arrdiv32_mux2to151_and1;
  assign f_arrdiv32_mux2to152_and0 = f_arrdiv32_mux2to120_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to152_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to152_and1 = f_arrdiv32_fs53_xor1 & f_arrdiv32_mux2to152_not0;
  assign f_arrdiv32_mux2to152_xor0 = f_arrdiv32_mux2to152_and0 ^ f_arrdiv32_mux2to152_and1;
  assign f_arrdiv32_mux2to153_and0 = f_arrdiv32_mux2to121_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to153_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to153_and1 = f_arrdiv32_fs54_xor1 & f_arrdiv32_mux2to153_not0;
  assign f_arrdiv32_mux2to153_xor0 = f_arrdiv32_mux2to153_and0 ^ f_arrdiv32_mux2to153_and1;
  assign f_arrdiv32_mux2to154_and0 = f_arrdiv32_mux2to122_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to154_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to154_and1 = f_arrdiv32_fs55_xor1 & f_arrdiv32_mux2to154_not0;
  assign f_arrdiv32_mux2to154_xor0 = f_arrdiv32_mux2to154_and0 ^ f_arrdiv32_mux2to154_and1;
  assign f_arrdiv32_mux2to155_and0 = f_arrdiv32_mux2to123_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to155_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to155_and1 = f_arrdiv32_fs56_xor1 & f_arrdiv32_mux2to155_not0;
  assign f_arrdiv32_mux2to155_xor0 = f_arrdiv32_mux2to155_and0 ^ f_arrdiv32_mux2to155_and1;
  assign f_arrdiv32_mux2to156_and0 = f_arrdiv32_mux2to124_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to156_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to156_and1 = f_arrdiv32_fs57_xor1 & f_arrdiv32_mux2to156_not0;
  assign f_arrdiv32_mux2to156_xor0 = f_arrdiv32_mux2to156_and0 ^ f_arrdiv32_mux2to156_and1;
  assign f_arrdiv32_mux2to157_and0 = f_arrdiv32_mux2to125_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to157_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to157_and1 = f_arrdiv32_fs58_xor1 & f_arrdiv32_mux2to157_not0;
  assign f_arrdiv32_mux2to157_xor0 = f_arrdiv32_mux2to157_and0 ^ f_arrdiv32_mux2to157_and1;
  assign f_arrdiv32_mux2to158_and0 = f_arrdiv32_mux2to126_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to158_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to158_and1 = f_arrdiv32_fs59_xor1 & f_arrdiv32_mux2to158_not0;
  assign f_arrdiv32_mux2to158_xor0 = f_arrdiv32_mux2to158_and0 ^ f_arrdiv32_mux2to158_and1;
  assign f_arrdiv32_mux2to159_and0 = f_arrdiv32_mux2to127_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to159_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to159_and1 = f_arrdiv32_fs60_xor1 & f_arrdiv32_mux2to159_not0;
  assign f_arrdiv32_mux2to159_xor0 = f_arrdiv32_mux2to159_and0 ^ f_arrdiv32_mux2to159_and1;
  assign f_arrdiv32_mux2to160_and0 = f_arrdiv32_mux2to128_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to160_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to160_and1 = f_arrdiv32_fs61_xor1 & f_arrdiv32_mux2to160_not0;
  assign f_arrdiv32_mux2to160_xor0 = f_arrdiv32_mux2to160_and0 ^ f_arrdiv32_mux2to160_and1;
  assign f_arrdiv32_mux2to161_and0 = f_arrdiv32_mux2to129_and1 & f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to161_not0 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_mux2to161_and1 = f_arrdiv32_fs62_xor1 & f_arrdiv32_mux2to161_not0;
  assign f_arrdiv32_mux2to161_xor0 = f_arrdiv32_mux2to161_and0 ^ f_arrdiv32_mux2to161_and1;
  assign f_arrdiv32_not1 = ~f_arrdiv32_fs63_or0;
  assign f_arrdiv32_fs64_xor0 = a[29] ^ b[0];
  assign f_arrdiv32_fs64_not0 = ~a[29];
  assign f_arrdiv32_fs64_and0 = f_arrdiv32_fs64_not0 & b[0];
  assign f_arrdiv32_fs64_not1 = ~f_arrdiv32_fs64_xor0;
  assign f_arrdiv32_fs65_xor0 = f_arrdiv32_mux2to131_xor0 ^ b[1];
  assign f_arrdiv32_fs65_not0 = ~f_arrdiv32_mux2to131_xor0;
  assign f_arrdiv32_fs65_and0 = f_arrdiv32_fs65_not0 & b[1];
  assign f_arrdiv32_fs65_xor1 = f_arrdiv32_fs64_and0 ^ f_arrdiv32_fs65_xor0;
  assign f_arrdiv32_fs65_not1 = ~f_arrdiv32_fs65_xor0;
  assign f_arrdiv32_fs65_and1 = f_arrdiv32_fs65_not1 & f_arrdiv32_fs64_and0;
  assign f_arrdiv32_fs65_or0 = f_arrdiv32_fs65_and1 | f_arrdiv32_fs65_and0;
  assign f_arrdiv32_fs66_xor0 = f_arrdiv32_mux2to132_xor0 ^ b[2];
  assign f_arrdiv32_fs66_not0 = ~f_arrdiv32_mux2to132_xor0;
  assign f_arrdiv32_fs66_and0 = f_arrdiv32_fs66_not0 & b[2];
  assign f_arrdiv32_fs66_xor1 = f_arrdiv32_fs65_or0 ^ f_arrdiv32_fs66_xor0;
  assign f_arrdiv32_fs66_not1 = ~f_arrdiv32_fs66_xor0;
  assign f_arrdiv32_fs66_and1 = f_arrdiv32_fs66_not1 & f_arrdiv32_fs65_or0;
  assign f_arrdiv32_fs66_or0 = f_arrdiv32_fs66_and1 | f_arrdiv32_fs66_and0;
  assign f_arrdiv32_fs67_xor0 = f_arrdiv32_mux2to133_xor0 ^ b[3];
  assign f_arrdiv32_fs67_not0 = ~f_arrdiv32_mux2to133_xor0;
  assign f_arrdiv32_fs67_and0 = f_arrdiv32_fs67_not0 & b[3];
  assign f_arrdiv32_fs67_xor1 = f_arrdiv32_fs66_or0 ^ f_arrdiv32_fs67_xor0;
  assign f_arrdiv32_fs67_not1 = ~f_arrdiv32_fs67_xor0;
  assign f_arrdiv32_fs67_and1 = f_arrdiv32_fs67_not1 & f_arrdiv32_fs66_or0;
  assign f_arrdiv32_fs67_or0 = f_arrdiv32_fs67_and1 | f_arrdiv32_fs67_and0;
  assign f_arrdiv32_fs68_xor0 = f_arrdiv32_mux2to134_xor0 ^ b[4];
  assign f_arrdiv32_fs68_not0 = ~f_arrdiv32_mux2to134_xor0;
  assign f_arrdiv32_fs68_and0 = f_arrdiv32_fs68_not0 & b[4];
  assign f_arrdiv32_fs68_xor1 = f_arrdiv32_fs67_or0 ^ f_arrdiv32_fs68_xor0;
  assign f_arrdiv32_fs68_not1 = ~f_arrdiv32_fs68_xor0;
  assign f_arrdiv32_fs68_and1 = f_arrdiv32_fs68_not1 & f_arrdiv32_fs67_or0;
  assign f_arrdiv32_fs68_or0 = f_arrdiv32_fs68_and1 | f_arrdiv32_fs68_and0;
  assign f_arrdiv32_fs69_xor0 = f_arrdiv32_mux2to135_xor0 ^ b[5];
  assign f_arrdiv32_fs69_not0 = ~f_arrdiv32_mux2to135_xor0;
  assign f_arrdiv32_fs69_and0 = f_arrdiv32_fs69_not0 & b[5];
  assign f_arrdiv32_fs69_xor1 = f_arrdiv32_fs68_or0 ^ f_arrdiv32_fs69_xor0;
  assign f_arrdiv32_fs69_not1 = ~f_arrdiv32_fs69_xor0;
  assign f_arrdiv32_fs69_and1 = f_arrdiv32_fs69_not1 & f_arrdiv32_fs68_or0;
  assign f_arrdiv32_fs69_or0 = f_arrdiv32_fs69_and1 | f_arrdiv32_fs69_and0;
  assign f_arrdiv32_fs70_xor0 = f_arrdiv32_mux2to136_xor0 ^ b[6];
  assign f_arrdiv32_fs70_not0 = ~f_arrdiv32_mux2to136_xor0;
  assign f_arrdiv32_fs70_and0 = f_arrdiv32_fs70_not0 & b[6];
  assign f_arrdiv32_fs70_xor1 = f_arrdiv32_fs69_or0 ^ f_arrdiv32_fs70_xor0;
  assign f_arrdiv32_fs70_not1 = ~f_arrdiv32_fs70_xor0;
  assign f_arrdiv32_fs70_and1 = f_arrdiv32_fs70_not1 & f_arrdiv32_fs69_or0;
  assign f_arrdiv32_fs70_or0 = f_arrdiv32_fs70_and1 | f_arrdiv32_fs70_and0;
  assign f_arrdiv32_fs71_xor0 = f_arrdiv32_mux2to137_xor0 ^ b[7];
  assign f_arrdiv32_fs71_not0 = ~f_arrdiv32_mux2to137_xor0;
  assign f_arrdiv32_fs71_and0 = f_arrdiv32_fs71_not0 & b[7];
  assign f_arrdiv32_fs71_xor1 = f_arrdiv32_fs70_or0 ^ f_arrdiv32_fs71_xor0;
  assign f_arrdiv32_fs71_not1 = ~f_arrdiv32_fs71_xor0;
  assign f_arrdiv32_fs71_and1 = f_arrdiv32_fs71_not1 & f_arrdiv32_fs70_or0;
  assign f_arrdiv32_fs71_or0 = f_arrdiv32_fs71_and1 | f_arrdiv32_fs71_and0;
  assign f_arrdiv32_fs72_xor0 = f_arrdiv32_mux2to138_xor0 ^ b[8];
  assign f_arrdiv32_fs72_not0 = ~f_arrdiv32_mux2to138_xor0;
  assign f_arrdiv32_fs72_and0 = f_arrdiv32_fs72_not0 & b[8];
  assign f_arrdiv32_fs72_xor1 = f_arrdiv32_fs71_or0 ^ f_arrdiv32_fs72_xor0;
  assign f_arrdiv32_fs72_not1 = ~f_arrdiv32_fs72_xor0;
  assign f_arrdiv32_fs72_and1 = f_arrdiv32_fs72_not1 & f_arrdiv32_fs71_or0;
  assign f_arrdiv32_fs72_or0 = f_arrdiv32_fs72_and1 | f_arrdiv32_fs72_and0;
  assign f_arrdiv32_fs73_xor0 = f_arrdiv32_mux2to139_xor0 ^ b[9];
  assign f_arrdiv32_fs73_not0 = ~f_arrdiv32_mux2to139_xor0;
  assign f_arrdiv32_fs73_and0 = f_arrdiv32_fs73_not0 & b[9];
  assign f_arrdiv32_fs73_xor1 = f_arrdiv32_fs72_or0 ^ f_arrdiv32_fs73_xor0;
  assign f_arrdiv32_fs73_not1 = ~f_arrdiv32_fs73_xor0;
  assign f_arrdiv32_fs73_and1 = f_arrdiv32_fs73_not1 & f_arrdiv32_fs72_or0;
  assign f_arrdiv32_fs73_or0 = f_arrdiv32_fs73_and1 | f_arrdiv32_fs73_and0;
  assign f_arrdiv32_fs74_xor0 = f_arrdiv32_mux2to140_xor0 ^ b[10];
  assign f_arrdiv32_fs74_not0 = ~f_arrdiv32_mux2to140_xor0;
  assign f_arrdiv32_fs74_and0 = f_arrdiv32_fs74_not0 & b[10];
  assign f_arrdiv32_fs74_xor1 = f_arrdiv32_fs73_or0 ^ f_arrdiv32_fs74_xor0;
  assign f_arrdiv32_fs74_not1 = ~f_arrdiv32_fs74_xor0;
  assign f_arrdiv32_fs74_and1 = f_arrdiv32_fs74_not1 & f_arrdiv32_fs73_or0;
  assign f_arrdiv32_fs74_or0 = f_arrdiv32_fs74_and1 | f_arrdiv32_fs74_and0;
  assign f_arrdiv32_fs75_xor0 = f_arrdiv32_mux2to141_xor0 ^ b[11];
  assign f_arrdiv32_fs75_not0 = ~f_arrdiv32_mux2to141_xor0;
  assign f_arrdiv32_fs75_and0 = f_arrdiv32_fs75_not0 & b[11];
  assign f_arrdiv32_fs75_xor1 = f_arrdiv32_fs74_or0 ^ f_arrdiv32_fs75_xor0;
  assign f_arrdiv32_fs75_not1 = ~f_arrdiv32_fs75_xor0;
  assign f_arrdiv32_fs75_and1 = f_arrdiv32_fs75_not1 & f_arrdiv32_fs74_or0;
  assign f_arrdiv32_fs75_or0 = f_arrdiv32_fs75_and1 | f_arrdiv32_fs75_and0;
  assign f_arrdiv32_fs76_xor0 = f_arrdiv32_mux2to142_xor0 ^ b[12];
  assign f_arrdiv32_fs76_not0 = ~f_arrdiv32_mux2to142_xor0;
  assign f_arrdiv32_fs76_and0 = f_arrdiv32_fs76_not0 & b[12];
  assign f_arrdiv32_fs76_xor1 = f_arrdiv32_fs75_or0 ^ f_arrdiv32_fs76_xor0;
  assign f_arrdiv32_fs76_not1 = ~f_arrdiv32_fs76_xor0;
  assign f_arrdiv32_fs76_and1 = f_arrdiv32_fs76_not1 & f_arrdiv32_fs75_or0;
  assign f_arrdiv32_fs76_or0 = f_arrdiv32_fs76_and1 | f_arrdiv32_fs76_and0;
  assign f_arrdiv32_fs77_xor0 = f_arrdiv32_mux2to143_xor0 ^ b[13];
  assign f_arrdiv32_fs77_not0 = ~f_arrdiv32_mux2to143_xor0;
  assign f_arrdiv32_fs77_and0 = f_arrdiv32_fs77_not0 & b[13];
  assign f_arrdiv32_fs77_xor1 = f_arrdiv32_fs76_or0 ^ f_arrdiv32_fs77_xor0;
  assign f_arrdiv32_fs77_not1 = ~f_arrdiv32_fs77_xor0;
  assign f_arrdiv32_fs77_and1 = f_arrdiv32_fs77_not1 & f_arrdiv32_fs76_or0;
  assign f_arrdiv32_fs77_or0 = f_arrdiv32_fs77_and1 | f_arrdiv32_fs77_and0;
  assign f_arrdiv32_fs78_xor0 = f_arrdiv32_mux2to144_xor0 ^ b[14];
  assign f_arrdiv32_fs78_not0 = ~f_arrdiv32_mux2to144_xor0;
  assign f_arrdiv32_fs78_and0 = f_arrdiv32_fs78_not0 & b[14];
  assign f_arrdiv32_fs78_xor1 = f_arrdiv32_fs77_or0 ^ f_arrdiv32_fs78_xor0;
  assign f_arrdiv32_fs78_not1 = ~f_arrdiv32_fs78_xor0;
  assign f_arrdiv32_fs78_and1 = f_arrdiv32_fs78_not1 & f_arrdiv32_fs77_or0;
  assign f_arrdiv32_fs78_or0 = f_arrdiv32_fs78_and1 | f_arrdiv32_fs78_and0;
  assign f_arrdiv32_fs79_xor0 = f_arrdiv32_mux2to145_xor0 ^ b[15];
  assign f_arrdiv32_fs79_not0 = ~f_arrdiv32_mux2to145_xor0;
  assign f_arrdiv32_fs79_and0 = f_arrdiv32_fs79_not0 & b[15];
  assign f_arrdiv32_fs79_xor1 = f_arrdiv32_fs78_or0 ^ f_arrdiv32_fs79_xor0;
  assign f_arrdiv32_fs79_not1 = ~f_arrdiv32_fs79_xor0;
  assign f_arrdiv32_fs79_and1 = f_arrdiv32_fs79_not1 & f_arrdiv32_fs78_or0;
  assign f_arrdiv32_fs79_or0 = f_arrdiv32_fs79_and1 | f_arrdiv32_fs79_and0;
  assign f_arrdiv32_fs80_xor0 = f_arrdiv32_mux2to146_xor0 ^ b[16];
  assign f_arrdiv32_fs80_not0 = ~f_arrdiv32_mux2to146_xor0;
  assign f_arrdiv32_fs80_and0 = f_arrdiv32_fs80_not0 & b[16];
  assign f_arrdiv32_fs80_xor1 = f_arrdiv32_fs79_or0 ^ f_arrdiv32_fs80_xor0;
  assign f_arrdiv32_fs80_not1 = ~f_arrdiv32_fs80_xor0;
  assign f_arrdiv32_fs80_and1 = f_arrdiv32_fs80_not1 & f_arrdiv32_fs79_or0;
  assign f_arrdiv32_fs80_or0 = f_arrdiv32_fs80_and1 | f_arrdiv32_fs80_and0;
  assign f_arrdiv32_fs81_xor0 = f_arrdiv32_mux2to147_xor0 ^ b[17];
  assign f_arrdiv32_fs81_not0 = ~f_arrdiv32_mux2to147_xor0;
  assign f_arrdiv32_fs81_and0 = f_arrdiv32_fs81_not0 & b[17];
  assign f_arrdiv32_fs81_xor1 = f_arrdiv32_fs80_or0 ^ f_arrdiv32_fs81_xor0;
  assign f_arrdiv32_fs81_not1 = ~f_arrdiv32_fs81_xor0;
  assign f_arrdiv32_fs81_and1 = f_arrdiv32_fs81_not1 & f_arrdiv32_fs80_or0;
  assign f_arrdiv32_fs81_or0 = f_arrdiv32_fs81_and1 | f_arrdiv32_fs81_and0;
  assign f_arrdiv32_fs82_xor0 = f_arrdiv32_mux2to148_xor0 ^ b[18];
  assign f_arrdiv32_fs82_not0 = ~f_arrdiv32_mux2to148_xor0;
  assign f_arrdiv32_fs82_and0 = f_arrdiv32_fs82_not0 & b[18];
  assign f_arrdiv32_fs82_xor1 = f_arrdiv32_fs81_or0 ^ f_arrdiv32_fs82_xor0;
  assign f_arrdiv32_fs82_not1 = ~f_arrdiv32_fs82_xor0;
  assign f_arrdiv32_fs82_and1 = f_arrdiv32_fs82_not1 & f_arrdiv32_fs81_or0;
  assign f_arrdiv32_fs82_or0 = f_arrdiv32_fs82_and1 | f_arrdiv32_fs82_and0;
  assign f_arrdiv32_fs83_xor0 = f_arrdiv32_mux2to149_xor0 ^ b[19];
  assign f_arrdiv32_fs83_not0 = ~f_arrdiv32_mux2to149_xor0;
  assign f_arrdiv32_fs83_and0 = f_arrdiv32_fs83_not0 & b[19];
  assign f_arrdiv32_fs83_xor1 = f_arrdiv32_fs82_or0 ^ f_arrdiv32_fs83_xor0;
  assign f_arrdiv32_fs83_not1 = ~f_arrdiv32_fs83_xor0;
  assign f_arrdiv32_fs83_and1 = f_arrdiv32_fs83_not1 & f_arrdiv32_fs82_or0;
  assign f_arrdiv32_fs83_or0 = f_arrdiv32_fs83_and1 | f_arrdiv32_fs83_and0;
  assign f_arrdiv32_fs84_xor0 = f_arrdiv32_mux2to150_xor0 ^ b[20];
  assign f_arrdiv32_fs84_not0 = ~f_arrdiv32_mux2to150_xor0;
  assign f_arrdiv32_fs84_and0 = f_arrdiv32_fs84_not0 & b[20];
  assign f_arrdiv32_fs84_xor1 = f_arrdiv32_fs83_or0 ^ f_arrdiv32_fs84_xor0;
  assign f_arrdiv32_fs84_not1 = ~f_arrdiv32_fs84_xor0;
  assign f_arrdiv32_fs84_and1 = f_arrdiv32_fs84_not1 & f_arrdiv32_fs83_or0;
  assign f_arrdiv32_fs84_or0 = f_arrdiv32_fs84_and1 | f_arrdiv32_fs84_and0;
  assign f_arrdiv32_fs85_xor0 = f_arrdiv32_mux2to151_xor0 ^ b[21];
  assign f_arrdiv32_fs85_not0 = ~f_arrdiv32_mux2to151_xor0;
  assign f_arrdiv32_fs85_and0 = f_arrdiv32_fs85_not0 & b[21];
  assign f_arrdiv32_fs85_xor1 = f_arrdiv32_fs84_or0 ^ f_arrdiv32_fs85_xor0;
  assign f_arrdiv32_fs85_not1 = ~f_arrdiv32_fs85_xor0;
  assign f_arrdiv32_fs85_and1 = f_arrdiv32_fs85_not1 & f_arrdiv32_fs84_or0;
  assign f_arrdiv32_fs85_or0 = f_arrdiv32_fs85_and1 | f_arrdiv32_fs85_and0;
  assign f_arrdiv32_fs86_xor0 = f_arrdiv32_mux2to152_xor0 ^ b[22];
  assign f_arrdiv32_fs86_not0 = ~f_arrdiv32_mux2to152_xor0;
  assign f_arrdiv32_fs86_and0 = f_arrdiv32_fs86_not0 & b[22];
  assign f_arrdiv32_fs86_xor1 = f_arrdiv32_fs85_or0 ^ f_arrdiv32_fs86_xor0;
  assign f_arrdiv32_fs86_not1 = ~f_arrdiv32_fs86_xor0;
  assign f_arrdiv32_fs86_and1 = f_arrdiv32_fs86_not1 & f_arrdiv32_fs85_or0;
  assign f_arrdiv32_fs86_or0 = f_arrdiv32_fs86_and1 | f_arrdiv32_fs86_and0;
  assign f_arrdiv32_fs87_xor0 = f_arrdiv32_mux2to153_xor0 ^ b[23];
  assign f_arrdiv32_fs87_not0 = ~f_arrdiv32_mux2to153_xor0;
  assign f_arrdiv32_fs87_and0 = f_arrdiv32_fs87_not0 & b[23];
  assign f_arrdiv32_fs87_xor1 = f_arrdiv32_fs86_or0 ^ f_arrdiv32_fs87_xor0;
  assign f_arrdiv32_fs87_not1 = ~f_arrdiv32_fs87_xor0;
  assign f_arrdiv32_fs87_and1 = f_arrdiv32_fs87_not1 & f_arrdiv32_fs86_or0;
  assign f_arrdiv32_fs87_or0 = f_arrdiv32_fs87_and1 | f_arrdiv32_fs87_and0;
  assign f_arrdiv32_fs88_xor0 = f_arrdiv32_mux2to154_xor0 ^ b[24];
  assign f_arrdiv32_fs88_not0 = ~f_arrdiv32_mux2to154_xor0;
  assign f_arrdiv32_fs88_and0 = f_arrdiv32_fs88_not0 & b[24];
  assign f_arrdiv32_fs88_xor1 = f_arrdiv32_fs87_or0 ^ f_arrdiv32_fs88_xor0;
  assign f_arrdiv32_fs88_not1 = ~f_arrdiv32_fs88_xor0;
  assign f_arrdiv32_fs88_and1 = f_arrdiv32_fs88_not1 & f_arrdiv32_fs87_or0;
  assign f_arrdiv32_fs88_or0 = f_arrdiv32_fs88_and1 | f_arrdiv32_fs88_and0;
  assign f_arrdiv32_fs89_xor0 = f_arrdiv32_mux2to155_xor0 ^ b[25];
  assign f_arrdiv32_fs89_not0 = ~f_arrdiv32_mux2to155_xor0;
  assign f_arrdiv32_fs89_and0 = f_arrdiv32_fs89_not0 & b[25];
  assign f_arrdiv32_fs89_xor1 = f_arrdiv32_fs88_or0 ^ f_arrdiv32_fs89_xor0;
  assign f_arrdiv32_fs89_not1 = ~f_arrdiv32_fs89_xor0;
  assign f_arrdiv32_fs89_and1 = f_arrdiv32_fs89_not1 & f_arrdiv32_fs88_or0;
  assign f_arrdiv32_fs89_or0 = f_arrdiv32_fs89_and1 | f_arrdiv32_fs89_and0;
  assign f_arrdiv32_fs90_xor0 = f_arrdiv32_mux2to156_xor0 ^ b[26];
  assign f_arrdiv32_fs90_not0 = ~f_arrdiv32_mux2to156_xor0;
  assign f_arrdiv32_fs90_and0 = f_arrdiv32_fs90_not0 & b[26];
  assign f_arrdiv32_fs90_xor1 = f_arrdiv32_fs89_or0 ^ f_arrdiv32_fs90_xor0;
  assign f_arrdiv32_fs90_not1 = ~f_arrdiv32_fs90_xor0;
  assign f_arrdiv32_fs90_and1 = f_arrdiv32_fs90_not1 & f_arrdiv32_fs89_or0;
  assign f_arrdiv32_fs90_or0 = f_arrdiv32_fs90_and1 | f_arrdiv32_fs90_and0;
  assign f_arrdiv32_fs91_xor0 = f_arrdiv32_mux2to157_xor0 ^ b[27];
  assign f_arrdiv32_fs91_not0 = ~f_arrdiv32_mux2to157_xor0;
  assign f_arrdiv32_fs91_and0 = f_arrdiv32_fs91_not0 & b[27];
  assign f_arrdiv32_fs91_xor1 = f_arrdiv32_fs90_or0 ^ f_arrdiv32_fs91_xor0;
  assign f_arrdiv32_fs91_not1 = ~f_arrdiv32_fs91_xor0;
  assign f_arrdiv32_fs91_and1 = f_arrdiv32_fs91_not1 & f_arrdiv32_fs90_or0;
  assign f_arrdiv32_fs91_or0 = f_arrdiv32_fs91_and1 | f_arrdiv32_fs91_and0;
  assign f_arrdiv32_fs92_xor0 = f_arrdiv32_mux2to158_xor0 ^ b[28];
  assign f_arrdiv32_fs92_not0 = ~f_arrdiv32_mux2to158_xor0;
  assign f_arrdiv32_fs92_and0 = f_arrdiv32_fs92_not0 & b[28];
  assign f_arrdiv32_fs92_xor1 = f_arrdiv32_fs91_or0 ^ f_arrdiv32_fs92_xor0;
  assign f_arrdiv32_fs92_not1 = ~f_arrdiv32_fs92_xor0;
  assign f_arrdiv32_fs92_and1 = f_arrdiv32_fs92_not1 & f_arrdiv32_fs91_or0;
  assign f_arrdiv32_fs92_or0 = f_arrdiv32_fs92_and1 | f_arrdiv32_fs92_and0;
  assign f_arrdiv32_fs93_xor0 = f_arrdiv32_mux2to159_xor0 ^ b[29];
  assign f_arrdiv32_fs93_not0 = ~f_arrdiv32_mux2to159_xor0;
  assign f_arrdiv32_fs93_and0 = f_arrdiv32_fs93_not0 & b[29];
  assign f_arrdiv32_fs93_xor1 = f_arrdiv32_fs92_or0 ^ f_arrdiv32_fs93_xor0;
  assign f_arrdiv32_fs93_not1 = ~f_arrdiv32_fs93_xor0;
  assign f_arrdiv32_fs93_and1 = f_arrdiv32_fs93_not1 & f_arrdiv32_fs92_or0;
  assign f_arrdiv32_fs93_or0 = f_arrdiv32_fs93_and1 | f_arrdiv32_fs93_and0;
  assign f_arrdiv32_fs94_xor0 = f_arrdiv32_mux2to160_xor0 ^ b[30];
  assign f_arrdiv32_fs94_not0 = ~f_arrdiv32_mux2to160_xor0;
  assign f_arrdiv32_fs94_and0 = f_arrdiv32_fs94_not0 & b[30];
  assign f_arrdiv32_fs94_xor1 = f_arrdiv32_fs93_or0 ^ f_arrdiv32_fs94_xor0;
  assign f_arrdiv32_fs94_not1 = ~f_arrdiv32_fs94_xor0;
  assign f_arrdiv32_fs94_and1 = f_arrdiv32_fs94_not1 & f_arrdiv32_fs93_or0;
  assign f_arrdiv32_fs94_or0 = f_arrdiv32_fs94_and1 | f_arrdiv32_fs94_and0;
  assign f_arrdiv32_fs95_xor0 = f_arrdiv32_mux2to161_xor0 ^ b[31];
  assign f_arrdiv32_fs95_not0 = ~f_arrdiv32_mux2to161_xor0;
  assign f_arrdiv32_fs95_and0 = f_arrdiv32_fs95_not0 & b[31];
  assign f_arrdiv32_fs95_xor1 = f_arrdiv32_fs94_or0 ^ f_arrdiv32_fs95_xor0;
  assign f_arrdiv32_fs95_not1 = ~f_arrdiv32_fs95_xor0;
  assign f_arrdiv32_fs95_and1 = f_arrdiv32_fs95_not1 & f_arrdiv32_fs94_or0;
  assign f_arrdiv32_fs95_or0 = f_arrdiv32_fs95_and1 | f_arrdiv32_fs95_and0;
  assign f_arrdiv32_mux2to162_and0 = a[29] & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to162_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to162_and1 = f_arrdiv32_fs64_xor0 & f_arrdiv32_mux2to162_not0;
  assign f_arrdiv32_mux2to162_xor0 = f_arrdiv32_mux2to162_and0 ^ f_arrdiv32_mux2to162_and1;
  assign f_arrdiv32_mux2to163_and0 = f_arrdiv32_mux2to131_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to163_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to163_and1 = f_arrdiv32_fs65_xor1 & f_arrdiv32_mux2to163_not0;
  assign f_arrdiv32_mux2to163_xor0 = f_arrdiv32_mux2to163_and0 ^ f_arrdiv32_mux2to163_and1;
  assign f_arrdiv32_mux2to164_and0 = f_arrdiv32_mux2to132_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to164_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to164_and1 = f_arrdiv32_fs66_xor1 & f_arrdiv32_mux2to164_not0;
  assign f_arrdiv32_mux2to164_xor0 = f_arrdiv32_mux2to164_and0 ^ f_arrdiv32_mux2to164_and1;
  assign f_arrdiv32_mux2to165_and0 = f_arrdiv32_mux2to133_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to165_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to165_and1 = f_arrdiv32_fs67_xor1 & f_arrdiv32_mux2to165_not0;
  assign f_arrdiv32_mux2to165_xor0 = f_arrdiv32_mux2to165_and0 ^ f_arrdiv32_mux2to165_and1;
  assign f_arrdiv32_mux2to166_and0 = f_arrdiv32_mux2to134_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to166_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to166_and1 = f_arrdiv32_fs68_xor1 & f_arrdiv32_mux2to166_not0;
  assign f_arrdiv32_mux2to166_xor0 = f_arrdiv32_mux2to166_and0 ^ f_arrdiv32_mux2to166_and1;
  assign f_arrdiv32_mux2to167_and0 = f_arrdiv32_mux2to135_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to167_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to167_and1 = f_arrdiv32_fs69_xor1 & f_arrdiv32_mux2to167_not0;
  assign f_arrdiv32_mux2to167_xor0 = f_arrdiv32_mux2to167_and0 ^ f_arrdiv32_mux2to167_and1;
  assign f_arrdiv32_mux2to168_and0 = f_arrdiv32_mux2to136_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to168_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to168_and1 = f_arrdiv32_fs70_xor1 & f_arrdiv32_mux2to168_not0;
  assign f_arrdiv32_mux2to168_xor0 = f_arrdiv32_mux2to168_and0 ^ f_arrdiv32_mux2to168_and1;
  assign f_arrdiv32_mux2to169_and0 = f_arrdiv32_mux2to137_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to169_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to169_and1 = f_arrdiv32_fs71_xor1 & f_arrdiv32_mux2to169_not0;
  assign f_arrdiv32_mux2to169_xor0 = f_arrdiv32_mux2to169_and0 ^ f_arrdiv32_mux2to169_and1;
  assign f_arrdiv32_mux2to170_and0 = f_arrdiv32_mux2to138_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to170_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to170_and1 = f_arrdiv32_fs72_xor1 & f_arrdiv32_mux2to170_not0;
  assign f_arrdiv32_mux2to170_xor0 = f_arrdiv32_mux2to170_and0 ^ f_arrdiv32_mux2to170_and1;
  assign f_arrdiv32_mux2to171_and0 = f_arrdiv32_mux2to139_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to171_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to171_and1 = f_arrdiv32_fs73_xor1 & f_arrdiv32_mux2to171_not0;
  assign f_arrdiv32_mux2to171_xor0 = f_arrdiv32_mux2to171_and0 ^ f_arrdiv32_mux2to171_and1;
  assign f_arrdiv32_mux2to172_and0 = f_arrdiv32_mux2to140_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to172_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to172_and1 = f_arrdiv32_fs74_xor1 & f_arrdiv32_mux2to172_not0;
  assign f_arrdiv32_mux2to172_xor0 = f_arrdiv32_mux2to172_and0 ^ f_arrdiv32_mux2to172_and1;
  assign f_arrdiv32_mux2to173_and0 = f_arrdiv32_mux2to141_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to173_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to173_and1 = f_arrdiv32_fs75_xor1 & f_arrdiv32_mux2to173_not0;
  assign f_arrdiv32_mux2to173_xor0 = f_arrdiv32_mux2to173_and0 ^ f_arrdiv32_mux2to173_and1;
  assign f_arrdiv32_mux2to174_and0 = f_arrdiv32_mux2to142_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to174_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to174_and1 = f_arrdiv32_fs76_xor1 & f_arrdiv32_mux2to174_not0;
  assign f_arrdiv32_mux2to174_xor0 = f_arrdiv32_mux2to174_and0 ^ f_arrdiv32_mux2to174_and1;
  assign f_arrdiv32_mux2to175_and0 = f_arrdiv32_mux2to143_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to175_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to175_and1 = f_arrdiv32_fs77_xor1 & f_arrdiv32_mux2to175_not0;
  assign f_arrdiv32_mux2to175_xor0 = f_arrdiv32_mux2to175_and0 ^ f_arrdiv32_mux2to175_and1;
  assign f_arrdiv32_mux2to176_and0 = f_arrdiv32_mux2to144_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to176_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to176_and1 = f_arrdiv32_fs78_xor1 & f_arrdiv32_mux2to176_not0;
  assign f_arrdiv32_mux2to176_xor0 = f_arrdiv32_mux2to176_and0 ^ f_arrdiv32_mux2to176_and1;
  assign f_arrdiv32_mux2to177_and0 = f_arrdiv32_mux2to145_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to177_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to177_and1 = f_arrdiv32_fs79_xor1 & f_arrdiv32_mux2to177_not0;
  assign f_arrdiv32_mux2to177_xor0 = f_arrdiv32_mux2to177_and0 ^ f_arrdiv32_mux2to177_and1;
  assign f_arrdiv32_mux2to178_and0 = f_arrdiv32_mux2to146_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to178_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to178_and1 = f_arrdiv32_fs80_xor1 & f_arrdiv32_mux2to178_not0;
  assign f_arrdiv32_mux2to178_xor0 = f_arrdiv32_mux2to178_and0 ^ f_arrdiv32_mux2to178_and1;
  assign f_arrdiv32_mux2to179_and0 = f_arrdiv32_mux2to147_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to179_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to179_and1 = f_arrdiv32_fs81_xor1 & f_arrdiv32_mux2to179_not0;
  assign f_arrdiv32_mux2to179_xor0 = f_arrdiv32_mux2to179_and0 ^ f_arrdiv32_mux2to179_and1;
  assign f_arrdiv32_mux2to180_and0 = f_arrdiv32_mux2to148_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to180_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to180_and1 = f_arrdiv32_fs82_xor1 & f_arrdiv32_mux2to180_not0;
  assign f_arrdiv32_mux2to180_xor0 = f_arrdiv32_mux2to180_and0 ^ f_arrdiv32_mux2to180_and1;
  assign f_arrdiv32_mux2to181_and0 = f_arrdiv32_mux2to149_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to181_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to181_and1 = f_arrdiv32_fs83_xor1 & f_arrdiv32_mux2to181_not0;
  assign f_arrdiv32_mux2to181_xor0 = f_arrdiv32_mux2to181_and0 ^ f_arrdiv32_mux2to181_and1;
  assign f_arrdiv32_mux2to182_and0 = f_arrdiv32_mux2to150_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to182_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to182_and1 = f_arrdiv32_fs84_xor1 & f_arrdiv32_mux2to182_not0;
  assign f_arrdiv32_mux2to182_xor0 = f_arrdiv32_mux2to182_and0 ^ f_arrdiv32_mux2to182_and1;
  assign f_arrdiv32_mux2to183_and0 = f_arrdiv32_mux2to151_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to183_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to183_and1 = f_arrdiv32_fs85_xor1 & f_arrdiv32_mux2to183_not0;
  assign f_arrdiv32_mux2to183_xor0 = f_arrdiv32_mux2to183_and0 ^ f_arrdiv32_mux2to183_and1;
  assign f_arrdiv32_mux2to184_and0 = f_arrdiv32_mux2to152_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to184_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to184_and1 = f_arrdiv32_fs86_xor1 & f_arrdiv32_mux2to184_not0;
  assign f_arrdiv32_mux2to184_xor0 = f_arrdiv32_mux2to184_and0 ^ f_arrdiv32_mux2to184_and1;
  assign f_arrdiv32_mux2to185_and0 = f_arrdiv32_mux2to153_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to185_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to185_and1 = f_arrdiv32_fs87_xor1 & f_arrdiv32_mux2to185_not0;
  assign f_arrdiv32_mux2to185_xor0 = f_arrdiv32_mux2to185_and0 ^ f_arrdiv32_mux2to185_and1;
  assign f_arrdiv32_mux2to186_and0 = f_arrdiv32_mux2to154_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to186_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to186_and1 = f_arrdiv32_fs88_xor1 & f_arrdiv32_mux2to186_not0;
  assign f_arrdiv32_mux2to186_xor0 = f_arrdiv32_mux2to186_and0 ^ f_arrdiv32_mux2to186_and1;
  assign f_arrdiv32_mux2to187_and0 = f_arrdiv32_mux2to155_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to187_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to187_and1 = f_arrdiv32_fs89_xor1 & f_arrdiv32_mux2to187_not0;
  assign f_arrdiv32_mux2to187_xor0 = f_arrdiv32_mux2to187_and0 ^ f_arrdiv32_mux2to187_and1;
  assign f_arrdiv32_mux2to188_and0 = f_arrdiv32_mux2to156_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to188_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to188_and1 = f_arrdiv32_fs90_xor1 & f_arrdiv32_mux2to188_not0;
  assign f_arrdiv32_mux2to188_xor0 = f_arrdiv32_mux2to188_and0 ^ f_arrdiv32_mux2to188_and1;
  assign f_arrdiv32_mux2to189_and0 = f_arrdiv32_mux2to157_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to189_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to189_and1 = f_arrdiv32_fs91_xor1 & f_arrdiv32_mux2to189_not0;
  assign f_arrdiv32_mux2to189_xor0 = f_arrdiv32_mux2to189_and0 ^ f_arrdiv32_mux2to189_and1;
  assign f_arrdiv32_mux2to190_and0 = f_arrdiv32_mux2to158_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to190_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to190_and1 = f_arrdiv32_fs92_xor1 & f_arrdiv32_mux2to190_not0;
  assign f_arrdiv32_mux2to190_xor0 = f_arrdiv32_mux2to190_and0 ^ f_arrdiv32_mux2to190_and1;
  assign f_arrdiv32_mux2to191_and0 = f_arrdiv32_mux2to159_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to191_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to191_and1 = f_arrdiv32_fs93_xor1 & f_arrdiv32_mux2to191_not0;
  assign f_arrdiv32_mux2to191_xor0 = f_arrdiv32_mux2to191_and0 ^ f_arrdiv32_mux2to191_and1;
  assign f_arrdiv32_mux2to192_and0 = f_arrdiv32_mux2to160_xor0 & f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to192_not0 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_mux2to192_and1 = f_arrdiv32_fs94_xor1 & f_arrdiv32_mux2to192_not0;
  assign f_arrdiv32_mux2to192_xor0 = f_arrdiv32_mux2to192_and0 ^ f_arrdiv32_mux2to192_and1;
  assign f_arrdiv32_not2 = ~f_arrdiv32_fs95_or0;
  assign f_arrdiv32_fs96_xor0 = a[28] ^ b[0];
  assign f_arrdiv32_fs96_not0 = ~a[28];
  assign f_arrdiv32_fs96_and0 = f_arrdiv32_fs96_not0 & b[0];
  assign f_arrdiv32_fs96_not1 = ~f_arrdiv32_fs96_xor0;
  assign f_arrdiv32_fs97_xor0 = f_arrdiv32_mux2to162_xor0 ^ b[1];
  assign f_arrdiv32_fs97_not0 = ~f_arrdiv32_mux2to162_xor0;
  assign f_arrdiv32_fs97_and0 = f_arrdiv32_fs97_not0 & b[1];
  assign f_arrdiv32_fs97_xor1 = f_arrdiv32_fs96_and0 ^ f_arrdiv32_fs97_xor0;
  assign f_arrdiv32_fs97_not1 = ~f_arrdiv32_fs97_xor0;
  assign f_arrdiv32_fs97_and1 = f_arrdiv32_fs97_not1 & f_arrdiv32_fs96_and0;
  assign f_arrdiv32_fs97_or0 = f_arrdiv32_fs97_and1 | f_arrdiv32_fs97_and0;
  assign f_arrdiv32_fs98_xor0 = f_arrdiv32_mux2to163_xor0 ^ b[2];
  assign f_arrdiv32_fs98_not0 = ~f_arrdiv32_mux2to163_xor0;
  assign f_arrdiv32_fs98_and0 = f_arrdiv32_fs98_not0 & b[2];
  assign f_arrdiv32_fs98_xor1 = f_arrdiv32_fs97_or0 ^ f_arrdiv32_fs98_xor0;
  assign f_arrdiv32_fs98_not1 = ~f_arrdiv32_fs98_xor0;
  assign f_arrdiv32_fs98_and1 = f_arrdiv32_fs98_not1 & f_arrdiv32_fs97_or0;
  assign f_arrdiv32_fs98_or0 = f_arrdiv32_fs98_and1 | f_arrdiv32_fs98_and0;
  assign f_arrdiv32_fs99_xor0 = f_arrdiv32_mux2to164_xor0 ^ b[3];
  assign f_arrdiv32_fs99_not0 = ~f_arrdiv32_mux2to164_xor0;
  assign f_arrdiv32_fs99_and0 = f_arrdiv32_fs99_not0 & b[3];
  assign f_arrdiv32_fs99_xor1 = f_arrdiv32_fs98_or0 ^ f_arrdiv32_fs99_xor0;
  assign f_arrdiv32_fs99_not1 = ~f_arrdiv32_fs99_xor0;
  assign f_arrdiv32_fs99_and1 = f_arrdiv32_fs99_not1 & f_arrdiv32_fs98_or0;
  assign f_arrdiv32_fs99_or0 = f_arrdiv32_fs99_and1 | f_arrdiv32_fs99_and0;
  assign f_arrdiv32_fs100_xor0 = f_arrdiv32_mux2to165_xor0 ^ b[4];
  assign f_arrdiv32_fs100_not0 = ~f_arrdiv32_mux2to165_xor0;
  assign f_arrdiv32_fs100_and0 = f_arrdiv32_fs100_not0 & b[4];
  assign f_arrdiv32_fs100_xor1 = f_arrdiv32_fs99_or0 ^ f_arrdiv32_fs100_xor0;
  assign f_arrdiv32_fs100_not1 = ~f_arrdiv32_fs100_xor0;
  assign f_arrdiv32_fs100_and1 = f_arrdiv32_fs100_not1 & f_arrdiv32_fs99_or0;
  assign f_arrdiv32_fs100_or0 = f_arrdiv32_fs100_and1 | f_arrdiv32_fs100_and0;
  assign f_arrdiv32_fs101_xor0 = f_arrdiv32_mux2to166_xor0 ^ b[5];
  assign f_arrdiv32_fs101_not0 = ~f_arrdiv32_mux2to166_xor0;
  assign f_arrdiv32_fs101_and0 = f_arrdiv32_fs101_not0 & b[5];
  assign f_arrdiv32_fs101_xor1 = f_arrdiv32_fs100_or0 ^ f_arrdiv32_fs101_xor0;
  assign f_arrdiv32_fs101_not1 = ~f_arrdiv32_fs101_xor0;
  assign f_arrdiv32_fs101_and1 = f_arrdiv32_fs101_not1 & f_arrdiv32_fs100_or0;
  assign f_arrdiv32_fs101_or0 = f_arrdiv32_fs101_and1 | f_arrdiv32_fs101_and0;
  assign f_arrdiv32_fs102_xor0 = f_arrdiv32_mux2to167_xor0 ^ b[6];
  assign f_arrdiv32_fs102_not0 = ~f_arrdiv32_mux2to167_xor0;
  assign f_arrdiv32_fs102_and0 = f_arrdiv32_fs102_not0 & b[6];
  assign f_arrdiv32_fs102_xor1 = f_arrdiv32_fs101_or0 ^ f_arrdiv32_fs102_xor0;
  assign f_arrdiv32_fs102_not1 = ~f_arrdiv32_fs102_xor0;
  assign f_arrdiv32_fs102_and1 = f_arrdiv32_fs102_not1 & f_arrdiv32_fs101_or0;
  assign f_arrdiv32_fs102_or0 = f_arrdiv32_fs102_and1 | f_arrdiv32_fs102_and0;
  assign f_arrdiv32_fs103_xor0 = f_arrdiv32_mux2to168_xor0 ^ b[7];
  assign f_arrdiv32_fs103_not0 = ~f_arrdiv32_mux2to168_xor0;
  assign f_arrdiv32_fs103_and0 = f_arrdiv32_fs103_not0 & b[7];
  assign f_arrdiv32_fs103_xor1 = f_arrdiv32_fs102_or0 ^ f_arrdiv32_fs103_xor0;
  assign f_arrdiv32_fs103_not1 = ~f_arrdiv32_fs103_xor0;
  assign f_arrdiv32_fs103_and1 = f_arrdiv32_fs103_not1 & f_arrdiv32_fs102_or0;
  assign f_arrdiv32_fs103_or0 = f_arrdiv32_fs103_and1 | f_arrdiv32_fs103_and0;
  assign f_arrdiv32_fs104_xor0 = f_arrdiv32_mux2to169_xor0 ^ b[8];
  assign f_arrdiv32_fs104_not0 = ~f_arrdiv32_mux2to169_xor0;
  assign f_arrdiv32_fs104_and0 = f_arrdiv32_fs104_not0 & b[8];
  assign f_arrdiv32_fs104_xor1 = f_arrdiv32_fs103_or0 ^ f_arrdiv32_fs104_xor0;
  assign f_arrdiv32_fs104_not1 = ~f_arrdiv32_fs104_xor0;
  assign f_arrdiv32_fs104_and1 = f_arrdiv32_fs104_not1 & f_arrdiv32_fs103_or0;
  assign f_arrdiv32_fs104_or0 = f_arrdiv32_fs104_and1 | f_arrdiv32_fs104_and0;
  assign f_arrdiv32_fs105_xor0 = f_arrdiv32_mux2to170_xor0 ^ b[9];
  assign f_arrdiv32_fs105_not0 = ~f_arrdiv32_mux2to170_xor0;
  assign f_arrdiv32_fs105_and0 = f_arrdiv32_fs105_not0 & b[9];
  assign f_arrdiv32_fs105_xor1 = f_arrdiv32_fs104_or0 ^ f_arrdiv32_fs105_xor0;
  assign f_arrdiv32_fs105_not1 = ~f_arrdiv32_fs105_xor0;
  assign f_arrdiv32_fs105_and1 = f_arrdiv32_fs105_not1 & f_arrdiv32_fs104_or0;
  assign f_arrdiv32_fs105_or0 = f_arrdiv32_fs105_and1 | f_arrdiv32_fs105_and0;
  assign f_arrdiv32_fs106_xor0 = f_arrdiv32_mux2to171_xor0 ^ b[10];
  assign f_arrdiv32_fs106_not0 = ~f_arrdiv32_mux2to171_xor0;
  assign f_arrdiv32_fs106_and0 = f_arrdiv32_fs106_not0 & b[10];
  assign f_arrdiv32_fs106_xor1 = f_arrdiv32_fs105_or0 ^ f_arrdiv32_fs106_xor0;
  assign f_arrdiv32_fs106_not1 = ~f_arrdiv32_fs106_xor0;
  assign f_arrdiv32_fs106_and1 = f_arrdiv32_fs106_not1 & f_arrdiv32_fs105_or0;
  assign f_arrdiv32_fs106_or0 = f_arrdiv32_fs106_and1 | f_arrdiv32_fs106_and0;
  assign f_arrdiv32_fs107_xor0 = f_arrdiv32_mux2to172_xor0 ^ b[11];
  assign f_arrdiv32_fs107_not0 = ~f_arrdiv32_mux2to172_xor0;
  assign f_arrdiv32_fs107_and0 = f_arrdiv32_fs107_not0 & b[11];
  assign f_arrdiv32_fs107_xor1 = f_arrdiv32_fs106_or0 ^ f_arrdiv32_fs107_xor0;
  assign f_arrdiv32_fs107_not1 = ~f_arrdiv32_fs107_xor0;
  assign f_arrdiv32_fs107_and1 = f_arrdiv32_fs107_not1 & f_arrdiv32_fs106_or0;
  assign f_arrdiv32_fs107_or0 = f_arrdiv32_fs107_and1 | f_arrdiv32_fs107_and0;
  assign f_arrdiv32_fs108_xor0 = f_arrdiv32_mux2to173_xor0 ^ b[12];
  assign f_arrdiv32_fs108_not0 = ~f_arrdiv32_mux2to173_xor0;
  assign f_arrdiv32_fs108_and0 = f_arrdiv32_fs108_not0 & b[12];
  assign f_arrdiv32_fs108_xor1 = f_arrdiv32_fs107_or0 ^ f_arrdiv32_fs108_xor0;
  assign f_arrdiv32_fs108_not1 = ~f_arrdiv32_fs108_xor0;
  assign f_arrdiv32_fs108_and1 = f_arrdiv32_fs108_not1 & f_arrdiv32_fs107_or0;
  assign f_arrdiv32_fs108_or0 = f_arrdiv32_fs108_and1 | f_arrdiv32_fs108_and0;
  assign f_arrdiv32_fs109_xor0 = f_arrdiv32_mux2to174_xor0 ^ b[13];
  assign f_arrdiv32_fs109_not0 = ~f_arrdiv32_mux2to174_xor0;
  assign f_arrdiv32_fs109_and0 = f_arrdiv32_fs109_not0 & b[13];
  assign f_arrdiv32_fs109_xor1 = f_arrdiv32_fs108_or0 ^ f_arrdiv32_fs109_xor0;
  assign f_arrdiv32_fs109_not1 = ~f_arrdiv32_fs109_xor0;
  assign f_arrdiv32_fs109_and1 = f_arrdiv32_fs109_not1 & f_arrdiv32_fs108_or0;
  assign f_arrdiv32_fs109_or0 = f_arrdiv32_fs109_and1 | f_arrdiv32_fs109_and0;
  assign f_arrdiv32_fs110_xor0 = f_arrdiv32_mux2to175_xor0 ^ b[14];
  assign f_arrdiv32_fs110_not0 = ~f_arrdiv32_mux2to175_xor0;
  assign f_arrdiv32_fs110_and0 = f_arrdiv32_fs110_not0 & b[14];
  assign f_arrdiv32_fs110_xor1 = f_arrdiv32_fs109_or0 ^ f_arrdiv32_fs110_xor0;
  assign f_arrdiv32_fs110_not1 = ~f_arrdiv32_fs110_xor0;
  assign f_arrdiv32_fs110_and1 = f_arrdiv32_fs110_not1 & f_arrdiv32_fs109_or0;
  assign f_arrdiv32_fs110_or0 = f_arrdiv32_fs110_and1 | f_arrdiv32_fs110_and0;
  assign f_arrdiv32_fs111_xor0 = f_arrdiv32_mux2to176_xor0 ^ b[15];
  assign f_arrdiv32_fs111_not0 = ~f_arrdiv32_mux2to176_xor0;
  assign f_arrdiv32_fs111_and0 = f_arrdiv32_fs111_not0 & b[15];
  assign f_arrdiv32_fs111_xor1 = f_arrdiv32_fs110_or0 ^ f_arrdiv32_fs111_xor0;
  assign f_arrdiv32_fs111_not1 = ~f_arrdiv32_fs111_xor0;
  assign f_arrdiv32_fs111_and1 = f_arrdiv32_fs111_not1 & f_arrdiv32_fs110_or0;
  assign f_arrdiv32_fs111_or0 = f_arrdiv32_fs111_and1 | f_arrdiv32_fs111_and0;
  assign f_arrdiv32_fs112_xor0 = f_arrdiv32_mux2to177_xor0 ^ b[16];
  assign f_arrdiv32_fs112_not0 = ~f_arrdiv32_mux2to177_xor0;
  assign f_arrdiv32_fs112_and0 = f_arrdiv32_fs112_not0 & b[16];
  assign f_arrdiv32_fs112_xor1 = f_arrdiv32_fs111_or0 ^ f_arrdiv32_fs112_xor0;
  assign f_arrdiv32_fs112_not1 = ~f_arrdiv32_fs112_xor0;
  assign f_arrdiv32_fs112_and1 = f_arrdiv32_fs112_not1 & f_arrdiv32_fs111_or0;
  assign f_arrdiv32_fs112_or0 = f_arrdiv32_fs112_and1 | f_arrdiv32_fs112_and0;
  assign f_arrdiv32_fs113_xor0 = f_arrdiv32_mux2to178_xor0 ^ b[17];
  assign f_arrdiv32_fs113_not0 = ~f_arrdiv32_mux2to178_xor0;
  assign f_arrdiv32_fs113_and0 = f_arrdiv32_fs113_not0 & b[17];
  assign f_arrdiv32_fs113_xor1 = f_arrdiv32_fs112_or0 ^ f_arrdiv32_fs113_xor0;
  assign f_arrdiv32_fs113_not1 = ~f_arrdiv32_fs113_xor0;
  assign f_arrdiv32_fs113_and1 = f_arrdiv32_fs113_not1 & f_arrdiv32_fs112_or0;
  assign f_arrdiv32_fs113_or0 = f_arrdiv32_fs113_and1 | f_arrdiv32_fs113_and0;
  assign f_arrdiv32_fs114_xor0 = f_arrdiv32_mux2to179_xor0 ^ b[18];
  assign f_arrdiv32_fs114_not0 = ~f_arrdiv32_mux2to179_xor0;
  assign f_arrdiv32_fs114_and0 = f_arrdiv32_fs114_not0 & b[18];
  assign f_arrdiv32_fs114_xor1 = f_arrdiv32_fs113_or0 ^ f_arrdiv32_fs114_xor0;
  assign f_arrdiv32_fs114_not1 = ~f_arrdiv32_fs114_xor0;
  assign f_arrdiv32_fs114_and1 = f_arrdiv32_fs114_not1 & f_arrdiv32_fs113_or0;
  assign f_arrdiv32_fs114_or0 = f_arrdiv32_fs114_and1 | f_arrdiv32_fs114_and0;
  assign f_arrdiv32_fs115_xor0 = f_arrdiv32_mux2to180_xor0 ^ b[19];
  assign f_arrdiv32_fs115_not0 = ~f_arrdiv32_mux2to180_xor0;
  assign f_arrdiv32_fs115_and0 = f_arrdiv32_fs115_not0 & b[19];
  assign f_arrdiv32_fs115_xor1 = f_arrdiv32_fs114_or0 ^ f_arrdiv32_fs115_xor0;
  assign f_arrdiv32_fs115_not1 = ~f_arrdiv32_fs115_xor0;
  assign f_arrdiv32_fs115_and1 = f_arrdiv32_fs115_not1 & f_arrdiv32_fs114_or0;
  assign f_arrdiv32_fs115_or0 = f_arrdiv32_fs115_and1 | f_arrdiv32_fs115_and0;
  assign f_arrdiv32_fs116_xor0 = f_arrdiv32_mux2to181_xor0 ^ b[20];
  assign f_arrdiv32_fs116_not0 = ~f_arrdiv32_mux2to181_xor0;
  assign f_arrdiv32_fs116_and0 = f_arrdiv32_fs116_not0 & b[20];
  assign f_arrdiv32_fs116_xor1 = f_arrdiv32_fs115_or0 ^ f_arrdiv32_fs116_xor0;
  assign f_arrdiv32_fs116_not1 = ~f_arrdiv32_fs116_xor0;
  assign f_arrdiv32_fs116_and1 = f_arrdiv32_fs116_not1 & f_arrdiv32_fs115_or0;
  assign f_arrdiv32_fs116_or0 = f_arrdiv32_fs116_and1 | f_arrdiv32_fs116_and0;
  assign f_arrdiv32_fs117_xor0 = f_arrdiv32_mux2to182_xor0 ^ b[21];
  assign f_arrdiv32_fs117_not0 = ~f_arrdiv32_mux2to182_xor0;
  assign f_arrdiv32_fs117_and0 = f_arrdiv32_fs117_not0 & b[21];
  assign f_arrdiv32_fs117_xor1 = f_arrdiv32_fs116_or0 ^ f_arrdiv32_fs117_xor0;
  assign f_arrdiv32_fs117_not1 = ~f_arrdiv32_fs117_xor0;
  assign f_arrdiv32_fs117_and1 = f_arrdiv32_fs117_not1 & f_arrdiv32_fs116_or0;
  assign f_arrdiv32_fs117_or0 = f_arrdiv32_fs117_and1 | f_arrdiv32_fs117_and0;
  assign f_arrdiv32_fs118_xor0 = f_arrdiv32_mux2to183_xor0 ^ b[22];
  assign f_arrdiv32_fs118_not0 = ~f_arrdiv32_mux2to183_xor0;
  assign f_arrdiv32_fs118_and0 = f_arrdiv32_fs118_not0 & b[22];
  assign f_arrdiv32_fs118_xor1 = f_arrdiv32_fs117_or0 ^ f_arrdiv32_fs118_xor0;
  assign f_arrdiv32_fs118_not1 = ~f_arrdiv32_fs118_xor0;
  assign f_arrdiv32_fs118_and1 = f_arrdiv32_fs118_not1 & f_arrdiv32_fs117_or0;
  assign f_arrdiv32_fs118_or0 = f_arrdiv32_fs118_and1 | f_arrdiv32_fs118_and0;
  assign f_arrdiv32_fs119_xor0 = f_arrdiv32_mux2to184_xor0 ^ b[23];
  assign f_arrdiv32_fs119_not0 = ~f_arrdiv32_mux2to184_xor0;
  assign f_arrdiv32_fs119_and0 = f_arrdiv32_fs119_not0 & b[23];
  assign f_arrdiv32_fs119_xor1 = f_arrdiv32_fs118_or0 ^ f_arrdiv32_fs119_xor0;
  assign f_arrdiv32_fs119_not1 = ~f_arrdiv32_fs119_xor0;
  assign f_arrdiv32_fs119_and1 = f_arrdiv32_fs119_not1 & f_arrdiv32_fs118_or0;
  assign f_arrdiv32_fs119_or0 = f_arrdiv32_fs119_and1 | f_arrdiv32_fs119_and0;
  assign f_arrdiv32_fs120_xor0 = f_arrdiv32_mux2to185_xor0 ^ b[24];
  assign f_arrdiv32_fs120_not0 = ~f_arrdiv32_mux2to185_xor0;
  assign f_arrdiv32_fs120_and0 = f_arrdiv32_fs120_not0 & b[24];
  assign f_arrdiv32_fs120_xor1 = f_arrdiv32_fs119_or0 ^ f_arrdiv32_fs120_xor0;
  assign f_arrdiv32_fs120_not1 = ~f_arrdiv32_fs120_xor0;
  assign f_arrdiv32_fs120_and1 = f_arrdiv32_fs120_not1 & f_arrdiv32_fs119_or0;
  assign f_arrdiv32_fs120_or0 = f_arrdiv32_fs120_and1 | f_arrdiv32_fs120_and0;
  assign f_arrdiv32_fs121_xor0 = f_arrdiv32_mux2to186_xor0 ^ b[25];
  assign f_arrdiv32_fs121_not0 = ~f_arrdiv32_mux2to186_xor0;
  assign f_arrdiv32_fs121_and0 = f_arrdiv32_fs121_not0 & b[25];
  assign f_arrdiv32_fs121_xor1 = f_arrdiv32_fs120_or0 ^ f_arrdiv32_fs121_xor0;
  assign f_arrdiv32_fs121_not1 = ~f_arrdiv32_fs121_xor0;
  assign f_arrdiv32_fs121_and1 = f_arrdiv32_fs121_not1 & f_arrdiv32_fs120_or0;
  assign f_arrdiv32_fs121_or0 = f_arrdiv32_fs121_and1 | f_arrdiv32_fs121_and0;
  assign f_arrdiv32_fs122_xor0 = f_arrdiv32_mux2to187_xor0 ^ b[26];
  assign f_arrdiv32_fs122_not0 = ~f_arrdiv32_mux2to187_xor0;
  assign f_arrdiv32_fs122_and0 = f_arrdiv32_fs122_not0 & b[26];
  assign f_arrdiv32_fs122_xor1 = f_arrdiv32_fs121_or0 ^ f_arrdiv32_fs122_xor0;
  assign f_arrdiv32_fs122_not1 = ~f_arrdiv32_fs122_xor0;
  assign f_arrdiv32_fs122_and1 = f_arrdiv32_fs122_not1 & f_arrdiv32_fs121_or0;
  assign f_arrdiv32_fs122_or0 = f_arrdiv32_fs122_and1 | f_arrdiv32_fs122_and0;
  assign f_arrdiv32_fs123_xor0 = f_arrdiv32_mux2to188_xor0 ^ b[27];
  assign f_arrdiv32_fs123_not0 = ~f_arrdiv32_mux2to188_xor0;
  assign f_arrdiv32_fs123_and0 = f_arrdiv32_fs123_not0 & b[27];
  assign f_arrdiv32_fs123_xor1 = f_arrdiv32_fs122_or0 ^ f_arrdiv32_fs123_xor0;
  assign f_arrdiv32_fs123_not1 = ~f_arrdiv32_fs123_xor0;
  assign f_arrdiv32_fs123_and1 = f_arrdiv32_fs123_not1 & f_arrdiv32_fs122_or0;
  assign f_arrdiv32_fs123_or0 = f_arrdiv32_fs123_and1 | f_arrdiv32_fs123_and0;
  assign f_arrdiv32_fs124_xor0 = f_arrdiv32_mux2to189_xor0 ^ b[28];
  assign f_arrdiv32_fs124_not0 = ~f_arrdiv32_mux2to189_xor0;
  assign f_arrdiv32_fs124_and0 = f_arrdiv32_fs124_not0 & b[28];
  assign f_arrdiv32_fs124_xor1 = f_arrdiv32_fs123_or0 ^ f_arrdiv32_fs124_xor0;
  assign f_arrdiv32_fs124_not1 = ~f_arrdiv32_fs124_xor0;
  assign f_arrdiv32_fs124_and1 = f_arrdiv32_fs124_not1 & f_arrdiv32_fs123_or0;
  assign f_arrdiv32_fs124_or0 = f_arrdiv32_fs124_and1 | f_arrdiv32_fs124_and0;
  assign f_arrdiv32_fs125_xor0 = f_arrdiv32_mux2to190_xor0 ^ b[29];
  assign f_arrdiv32_fs125_not0 = ~f_arrdiv32_mux2to190_xor0;
  assign f_arrdiv32_fs125_and0 = f_arrdiv32_fs125_not0 & b[29];
  assign f_arrdiv32_fs125_xor1 = f_arrdiv32_fs124_or0 ^ f_arrdiv32_fs125_xor0;
  assign f_arrdiv32_fs125_not1 = ~f_arrdiv32_fs125_xor0;
  assign f_arrdiv32_fs125_and1 = f_arrdiv32_fs125_not1 & f_arrdiv32_fs124_or0;
  assign f_arrdiv32_fs125_or0 = f_arrdiv32_fs125_and1 | f_arrdiv32_fs125_and0;
  assign f_arrdiv32_fs126_xor0 = f_arrdiv32_mux2to191_xor0 ^ b[30];
  assign f_arrdiv32_fs126_not0 = ~f_arrdiv32_mux2to191_xor0;
  assign f_arrdiv32_fs126_and0 = f_arrdiv32_fs126_not0 & b[30];
  assign f_arrdiv32_fs126_xor1 = f_arrdiv32_fs125_or0 ^ f_arrdiv32_fs126_xor0;
  assign f_arrdiv32_fs126_not1 = ~f_arrdiv32_fs126_xor0;
  assign f_arrdiv32_fs126_and1 = f_arrdiv32_fs126_not1 & f_arrdiv32_fs125_or0;
  assign f_arrdiv32_fs126_or0 = f_arrdiv32_fs126_and1 | f_arrdiv32_fs126_and0;
  assign f_arrdiv32_fs127_xor0 = f_arrdiv32_mux2to192_xor0 ^ b[31];
  assign f_arrdiv32_fs127_not0 = ~f_arrdiv32_mux2to192_xor0;
  assign f_arrdiv32_fs127_and0 = f_arrdiv32_fs127_not0 & b[31];
  assign f_arrdiv32_fs127_xor1 = f_arrdiv32_fs126_or0 ^ f_arrdiv32_fs127_xor0;
  assign f_arrdiv32_fs127_not1 = ~f_arrdiv32_fs127_xor0;
  assign f_arrdiv32_fs127_and1 = f_arrdiv32_fs127_not1 & f_arrdiv32_fs126_or0;
  assign f_arrdiv32_fs127_or0 = f_arrdiv32_fs127_and1 | f_arrdiv32_fs127_and0;
  assign f_arrdiv32_mux2to193_and0 = a[28] & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to193_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to193_and1 = f_arrdiv32_fs96_xor0 & f_arrdiv32_mux2to193_not0;
  assign f_arrdiv32_mux2to193_xor0 = f_arrdiv32_mux2to193_and0 ^ f_arrdiv32_mux2to193_and1;
  assign f_arrdiv32_mux2to194_and0 = f_arrdiv32_mux2to162_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to194_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to194_and1 = f_arrdiv32_fs97_xor1 & f_arrdiv32_mux2to194_not0;
  assign f_arrdiv32_mux2to194_xor0 = f_arrdiv32_mux2to194_and0 ^ f_arrdiv32_mux2to194_and1;
  assign f_arrdiv32_mux2to195_and0 = f_arrdiv32_mux2to163_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to195_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to195_and1 = f_arrdiv32_fs98_xor1 & f_arrdiv32_mux2to195_not0;
  assign f_arrdiv32_mux2to195_xor0 = f_arrdiv32_mux2to195_and0 ^ f_arrdiv32_mux2to195_and1;
  assign f_arrdiv32_mux2to196_and0 = f_arrdiv32_mux2to164_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to196_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to196_and1 = f_arrdiv32_fs99_xor1 & f_arrdiv32_mux2to196_not0;
  assign f_arrdiv32_mux2to196_xor0 = f_arrdiv32_mux2to196_and0 ^ f_arrdiv32_mux2to196_and1;
  assign f_arrdiv32_mux2to197_and0 = f_arrdiv32_mux2to165_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to197_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to197_and1 = f_arrdiv32_fs100_xor1 & f_arrdiv32_mux2to197_not0;
  assign f_arrdiv32_mux2to197_xor0 = f_arrdiv32_mux2to197_and0 ^ f_arrdiv32_mux2to197_and1;
  assign f_arrdiv32_mux2to198_and0 = f_arrdiv32_mux2to166_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to198_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to198_and1 = f_arrdiv32_fs101_xor1 & f_arrdiv32_mux2to198_not0;
  assign f_arrdiv32_mux2to198_xor0 = f_arrdiv32_mux2to198_and0 ^ f_arrdiv32_mux2to198_and1;
  assign f_arrdiv32_mux2to199_and0 = f_arrdiv32_mux2to167_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to199_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to199_and1 = f_arrdiv32_fs102_xor1 & f_arrdiv32_mux2to199_not0;
  assign f_arrdiv32_mux2to199_xor0 = f_arrdiv32_mux2to199_and0 ^ f_arrdiv32_mux2to199_and1;
  assign f_arrdiv32_mux2to1100_and0 = f_arrdiv32_mux2to168_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1100_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1100_and1 = f_arrdiv32_fs103_xor1 & f_arrdiv32_mux2to1100_not0;
  assign f_arrdiv32_mux2to1100_xor0 = f_arrdiv32_mux2to1100_and0 ^ f_arrdiv32_mux2to1100_and1;
  assign f_arrdiv32_mux2to1101_and0 = f_arrdiv32_mux2to169_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1101_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1101_and1 = f_arrdiv32_fs104_xor1 & f_arrdiv32_mux2to1101_not0;
  assign f_arrdiv32_mux2to1101_xor0 = f_arrdiv32_mux2to1101_and0 ^ f_arrdiv32_mux2to1101_and1;
  assign f_arrdiv32_mux2to1102_and0 = f_arrdiv32_mux2to170_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1102_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1102_and1 = f_arrdiv32_fs105_xor1 & f_arrdiv32_mux2to1102_not0;
  assign f_arrdiv32_mux2to1102_xor0 = f_arrdiv32_mux2to1102_and0 ^ f_arrdiv32_mux2to1102_and1;
  assign f_arrdiv32_mux2to1103_and0 = f_arrdiv32_mux2to171_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1103_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1103_and1 = f_arrdiv32_fs106_xor1 & f_arrdiv32_mux2to1103_not0;
  assign f_arrdiv32_mux2to1103_xor0 = f_arrdiv32_mux2to1103_and0 ^ f_arrdiv32_mux2to1103_and1;
  assign f_arrdiv32_mux2to1104_and0 = f_arrdiv32_mux2to172_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1104_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1104_and1 = f_arrdiv32_fs107_xor1 & f_arrdiv32_mux2to1104_not0;
  assign f_arrdiv32_mux2to1104_xor0 = f_arrdiv32_mux2to1104_and0 ^ f_arrdiv32_mux2to1104_and1;
  assign f_arrdiv32_mux2to1105_and0 = f_arrdiv32_mux2to173_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1105_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1105_and1 = f_arrdiv32_fs108_xor1 & f_arrdiv32_mux2to1105_not0;
  assign f_arrdiv32_mux2to1105_xor0 = f_arrdiv32_mux2to1105_and0 ^ f_arrdiv32_mux2to1105_and1;
  assign f_arrdiv32_mux2to1106_and0 = f_arrdiv32_mux2to174_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1106_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1106_and1 = f_arrdiv32_fs109_xor1 & f_arrdiv32_mux2to1106_not0;
  assign f_arrdiv32_mux2to1106_xor0 = f_arrdiv32_mux2to1106_and0 ^ f_arrdiv32_mux2to1106_and1;
  assign f_arrdiv32_mux2to1107_and0 = f_arrdiv32_mux2to175_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1107_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1107_and1 = f_arrdiv32_fs110_xor1 & f_arrdiv32_mux2to1107_not0;
  assign f_arrdiv32_mux2to1107_xor0 = f_arrdiv32_mux2to1107_and0 ^ f_arrdiv32_mux2to1107_and1;
  assign f_arrdiv32_mux2to1108_and0 = f_arrdiv32_mux2to176_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1108_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1108_and1 = f_arrdiv32_fs111_xor1 & f_arrdiv32_mux2to1108_not0;
  assign f_arrdiv32_mux2to1108_xor0 = f_arrdiv32_mux2to1108_and0 ^ f_arrdiv32_mux2to1108_and1;
  assign f_arrdiv32_mux2to1109_and0 = f_arrdiv32_mux2to177_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1109_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1109_and1 = f_arrdiv32_fs112_xor1 & f_arrdiv32_mux2to1109_not0;
  assign f_arrdiv32_mux2to1109_xor0 = f_arrdiv32_mux2to1109_and0 ^ f_arrdiv32_mux2to1109_and1;
  assign f_arrdiv32_mux2to1110_and0 = f_arrdiv32_mux2to178_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1110_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1110_and1 = f_arrdiv32_fs113_xor1 & f_arrdiv32_mux2to1110_not0;
  assign f_arrdiv32_mux2to1110_xor0 = f_arrdiv32_mux2to1110_and0 ^ f_arrdiv32_mux2to1110_and1;
  assign f_arrdiv32_mux2to1111_and0 = f_arrdiv32_mux2to179_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1111_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1111_and1 = f_arrdiv32_fs114_xor1 & f_arrdiv32_mux2to1111_not0;
  assign f_arrdiv32_mux2to1111_xor0 = f_arrdiv32_mux2to1111_and0 ^ f_arrdiv32_mux2to1111_and1;
  assign f_arrdiv32_mux2to1112_and0 = f_arrdiv32_mux2to180_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1112_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1112_and1 = f_arrdiv32_fs115_xor1 & f_arrdiv32_mux2to1112_not0;
  assign f_arrdiv32_mux2to1112_xor0 = f_arrdiv32_mux2to1112_and0 ^ f_arrdiv32_mux2to1112_and1;
  assign f_arrdiv32_mux2to1113_and0 = f_arrdiv32_mux2to181_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1113_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1113_and1 = f_arrdiv32_fs116_xor1 & f_arrdiv32_mux2to1113_not0;
  assign f_arrdiv32_mux2to1113_xor0 = f_arrdiv32_mux2to1113_and0 ^ f_arrdiv32_mux2to1113_and1;
  assign f_arrdiv32_mux2to1114_and0 = f_arrdiv32_mux2to182_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1114_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1114_and1 = f_arrdiv32_fs117_xor1 & f_arrdiv32_mux2to1114_not0;
  assign f_arrdiv32_mux2to1114_xor0 = f_arrdiv32_mux2to1114_and0 ^ f_arrdiv32_mux2to1114_and1;
  assign f_arrdiv32_mux2to1115_and0 = f_arrdiv32_mux2to183_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1115_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1115_and1 = f_arrdiv32_fs118_xor1 & f_arrdiv32_mux2to1115_not0;
  assign f_arrdiv32_mux2to1115_xor0 = f_arrdiv32_mux2to1115_and0 ^ f_arrdiv32_mux2to1115_and1;
  assign f_arrdiv32_mux2to1116_and0 = f_arrdiv32_mux2to184_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1116_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1116_and1 = f_arrdiv32_fs119_xor1 & f_arrdiv32_mux2to1116_not0;
  assign f_arrdiv32_mux2to1116_xor0 = f_arrdiv32_mux2to1116_and0 ^ f_arrdiv32_mux2to1116_and1;
  assign f_arrdiv32_mux2to1117_and0 = f_arrdiv32_mux2to185_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1117_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1117_and1 = f_arrdiv32_fs120_xor1 & f_arrdiv32_mux2to1117_not0;
  assign f_arrdiv32_mux2to1117_xor0 = f_arrdiv32_mux2to1117_and0 ^ f_arrdiv32_mux2to1117_and1;
  assign f_arrdiv32_mux2to1118_and0 = f_arrdiv32_mux2to186_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1118_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1118_and1 = f_arrdiv32_fs121_xor1 & f_arrdiv32_mux2to1118_not0;
  assign f_arrdiv32_mux2to1118_xor0 = f_arrdiv32_mux2to1118_and0 ^ f_arrdiv32_mux2to1118_and1;
  assign f_arrdiv32_mux2to1119_and0 = f_arrdiv32_mux2to187_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1119_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1119_and1 = f_arrdiv32_fs122_xor1 & f_arrdiv32_mux2to1119_not0;
  assign f_arrdiv32_mux2to1119_xor0 = f_arrdiv32_mux2to1119_and0 ^ f_arrdiv32_mux2to1119_and1;
  assign f_arrdiv32_mux2to1120_and0 = f_arrdiv32_mux2to188_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1120_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1120_and1 = f_arrdiv32_fs123_xor1 & f_arrdiv32_mux2to1120_not0;
  assign f_arrdiv32_mux2to1120_xor0 = f_arrdiv32_mux2to1120_and0 ^ f_arrdiv32_mux2to1120_and1;
  assign f_arrdiv32_mux2to1121_and0 = f_arrdiv32_mux2to189_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1121_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1121_and1 = f_arrdiv32_fs124_xor1 & f_arrdiv32_mux2to1121_not0;
  assign f_arrdiv32_mux2to1121_xor0 = f_arrdiv32_mux2to1121_and0 ^ f_arrdiv32_mux2to1121_and1;
  assign f_arrdiv32_mux2to1122_and0 = f_arrdiv32_mux2to190_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1122_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1122_and1 = f_arrdiv32_fs125_xor1 & f_arrdiv32_mux2to1122_not0;
  assign f_arrdiv32_mux2to1122_xor0 = f_arrdiv32_mux2to1122_and0 ^ f_arrdiv32_mux2to1122_and1;
  assign f_arrdiv32_mux2to1123_and0 = f_arrdiv32_mux2to191_xor0 & f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1123_not0 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_mux2to1123_and1 = f_arrdiv32_fs126_xor1 & f_arrdiv32_mux2to1123_not0;
  assign f_arrdiv32_mux2to1123_xor0 = f_arrdiv32_mux2to1123_and0 ^ f_arrdiv32_mux2to1123_and1;
  assign f_arrdiv32_not3 = ~f_arrdiv32_fs127_or0;
  assign f_arrdiv32_fs128_xor0 = a[27] ^ b[0];
  assign f_arrdiv32_fs128_not0 = ~a[27];
  assign f_arrdiv32_fs128_and0 = f_arrdiv32_fs128_not0 & b[0];
  assign f_arrdiv32_fs128_not1 = ~f_arrdiv32_fs128_xor0;
  assign f_arrdiv32_fs129_xor0 = f_arrdiv32_mux2to193_xor0 ^ b[1];
  assign f_arrdiv32_fs129_not0 = ~f_arrdiv32_mux2to193_xor0;
  assign f_arrdiv32_fs129_and0 = f_arrdiv32_fs129_not0 & b[1];
  assign f_arrdiv32_fs129_xor1 = f_arrdiv32_fs128_and0 ^ f_arrdiv32_fs129_xor0;
  assign f_arrdiv32_fs129_not1 = ~f_arrdiv32_fs129_xor0;
  assign f_arrdiv32_fs129_and1 = f_arrdiv32_fs129_not1 & f_arrdiv32_fs128_and0;
  assign f_arrdiv32_fs129_or0 = f_arrdiv32_fs129_and1 | f_arrdiv32_fs129_and0;
  assign f_arrdiv32_fs130_xor0 = f_arrdiv32_mux2to194_xor0 ^ b[2];
  assign f_arrdiv32_fs130_not0 = ~f_arrdiv32_mux2to194_xor0;
  assign f_arrdiv32_fs130_and0 = f_arrdiv32_fs130_not0 & b[2];
  assign f_arrdiv32_fs130_xor1 = f_arrdiv32_fs129_or0 ^ f_arrdiv32_fs130_xor0;
  assign f_arrdiv32_fs130_not1 = ~f_arrdiv32_fs130_xor0;
  assign f_arrdiv32_fs130_and1 = f_arrdiv32_fs130_not1 & f_arrdiv32_fs129_or0;
  assign f_arrdiv32_fs130_or0 = f_arrdiv32_fs130_and1 | f_arrdiv32_fs130_and0;
  assign f_arrdiv32_fs131_xor0 = f_arrdiv32_mux2to195_xor0 ^ b[3];
  assign f_arrdiv32_fs131_not0 = ~f_arrdiv32_mux2to195_xor0;
  assign f_arrdiv32_fs131_and0 = f_arrdiv32_fs131_not0 & b[3];
  assign f_arrdiv32_fs131_xor1 = f_arrdiv32_fs130_or0 ^ f_arrdiv32_fs131_xor0;
  assign f_arrdiv32_fs131_not1 = ~f_arrdiv32_fs131_xor0;
  assign f_arrdiv32_fs131_and1 = f_arrdiv32_fs131_not1 & f_arrdiv32_fs130_or0;
  assign f_arrdiv32_fs131_or0 = f_arrdiv32_fs131_and1 | f_arrdiv32_fs131_and0;
  assign f_arrdiv32_fs132_xor0 = f_arrdiv32_mux2to196_xor0 ^ b[4];
  assign f_arrdiv32_fs132_not0 = ~f_arrdiv32_mux2to196_xor0;
  assign f_arrdiv32_fs132_and0 = f_arrdiv32_fs132_not0 & b[4];
  assign f_arrdiv32_fs132_xor1 = f_arrdiv32_fs131_or0 ^ f_arrdiv32_fs132_xor0;
  assign f_arrdiv32_fs132_not1 = ~f_arrdiv32_fs132_xor0;
  assign f_arrdiv32_fs132_and1 = f_arrdiv32_fs132_not1 & f_arrdiv32_fs131_or0;
  assign f_arrdiv32_fs132_or0 = f_arrdiv32_fs132_and1 | f_arrdiv32_fs132_and0;
  assign f_arrdiv32_fs133_xor0 = f_arrdiv32_mux2to197_xor0 ^ b[5];
  assign f_arrdiv32_fs133_not0 = ~f_arrdiv32_mux2to197_xor0;
  assign f_arrdiv32_fs133_and0 = f_arrdiv32_fs133_not0 & b[5];
  assign f_arrdiv32_fs133_xor1 = f_arrdiv32_fs132_or0 ^ f_arrdiv32_fs133_xor0;
  assign f_arrdiv32_fs133_not1 = ~f_arrdiv32_fs133_xor0;
  assign f_arrdiv32_fs133_and1 = f_arrdiv32_fs133_not1 & f_arrdiv32_fs132_or0;
  assign f_arrdiv32_fs133_or0 = f_arrdiv32_fs133_and1 | f_arrdiv32_fs133_and0;
  assign f_arrdiv32_fs134_xor0 = f_arrdiv32_mux2to198_xor0 ^ b[6];
  assign f_arrdiv32_fs134_not0 = ~f_arrdiv32_mux2to198_xor0;
  assign f_arrdiv32_fs134_and0 = f_arrdiv32_fs134_not0 & b[6];
  assign f_arrdiv32_fs134_xor1 = f_arrdiv32_fs133_or0 ^ f_arrdiv32_fs134_xor0;
  assign f_arrdiv32_fs134_not1 = ~f_arrdiv32_fs134_xor0;
  assign f_arrdiv32_fs134_and1 = f_arrdiv32_fs134_not1 & f_arrdiv32_fs133_or0;
  assign f_arrdiv32_fs134_or0 = f_arrdiv32_fs134_and1 | f_arrdiv32_fs134_and0;
  assign f_arrdiv32_fs135_xor0 = f_arrdiv32_mux2to199_xor0 ^ b[7];
  assign f_arrdiv32_fs135_not0 = ~f_arrdiv32_mux2to199_xor0;
  assign f_arrdiv32_fs135_and0 = f_arrdiv32_fs135_not0 & b[7];
  assign f_arrdiv32_fs135_xor1 = f_arrdiv32_fs134_or0 ^ f_arrdiv32_fs135_xor0;
  assign f_arrdiv32_fs135_not1 = ~f_arrdiv32_fs135_xor0;
  assign f_arrdiv32_fs135_and1 = f_arrdiv32_fs135_not1 & f_arrdiv32_fs134_or0;
  assign f_arrdiv32_fs135_or0 = f_arrdiv32_fs135_and1 | f_arrdiv32_fs135_and0;
  assign f_arrdiv32_fs136_xor0 = f_arrdiv32_mux2to1100_xor0 ^ b[8];
  assign f_arrdiv32_fs136_not0 = ~f_arrdiv32_mux2to1100_xor0;
  assign f_arrdiv32_fs136_and0 = f_arrdiv32_fs136_not0 & b[8];
  assign f_arrdiv32_fs136_xor1 = f_arrdiv32_fs135_or0 ^ f_arrdiv32_fs136_xor0;
  assign f_arrdiv32_fs136_not1 = ~f_arrdiv32_fs136_xor0;
  assign f_arrdiv32_fs136_and1 = f_arrdiv32_fs136_not1 & f_arrdiv32_fs135_or0;
  assign f_arrdiv32_fs136_or0 = f_arrdiv32_fs136_and1 | f_arrdiv32_fs136_and0;
  assign f_arrdiv32_fs137_xor0 = f_arrdiv32_mux2to1101_xor0 ^ b[9];
  assign f_arrdiv32_fs137_not0 = ~f_arrdiv32_mux2to1101_xor0;
  assign f_arrdiv32_fs137_and0 = f_arrdiv32_fs137_not0 & b[9];
  assign f_arrdiv32_fs137_xor1 = f_arrdiv32_fs136_or0 ^ f_arrdiv32_fs137_xor0;
  assign f_arrdiv32_fs137_not1 = ~f_arrdiv32_fs137_xor0;
  assign f_arrdiv32_fs137_and1 = f_arrdiv32_fs137_not1 & f_arrdiv32_fs136_or0;
  assign f_arrdiv32_fs137_or0 = f_arrdiv32_fs137_and1 | f_arrdiv32_fs137_and0;
  assign f_arrdiv32_fs138_xor0 = f_arrdiv32_mux2to1102_xor0 ^ b[10];
  assign f_arrdiv32_fs138_not0 = ~f_arrdiv32_mux2to1102_xor0;
  assign f_arrdiv32_fs138_and0 = f_arrdiv32_fs138_not0 & b[10];
  assign f_arrdiv32_fs138_xor1 = f_arrdiv32_fs137_or0 ^ f_arrdiv32_fs138_xor0;
  assign f_arrdiv32_fs138_not1 = ~f_arrdiv32_fs138_xor0;
  assign f_arrdiv32_fs138_and1 = f_arrdiv32_fs138_not1 & f_arrdiv32_fs137_or0;
  assign f_arrdiv32_fs138_or0 = f_arrdiv32_fs138_and1 | f_arrdiv32_fs138_and0;
  assign f_arrdiv32_fs139_xor0 = f_arrdiv32_mux2to1103_xor0 ^ b[11];
  assign f_arrdiv32_fs139_not0 = ~f_arrdiv32_mux2to1103_xor0;
  assign f_arrdiv32_fs139_and0 = f_arrdiv32_fs139_not0 & b[11];
  assign f_arrdiv32_fs139_xor1 = f_arrdiv32_fs138_or0 ^ f_arrdiv32_fs139_xor0;
  assign f_arrdiv32_fs139_not1 = ~f_arrdiv32_fs139_xor0;
  assign f_arrdiv32_fs139_and1 = f_arrdiv32_fs139_not1 & f_arrdiv32_fs138_or0;
  assign f_arrdiv32_fs139_or0 = f_arrdiv32_fs139_and1 | f_arrdiv32_fs139_and0;
  assign f_arrdiv32_fs140_xor0 = f_arrdiv32_mux2to1104_xor0 ^ b[12];
  assign f_arrdiv32_fs140_not0 = ~f_arrdiv32_mux2to1104_xor0;
  assign f_arrdiv32_fs140_and0 = f_arrdiv32_fs140_not0 & b[12];
  assign f_arrdiv32_fs140_xor1 = f_arrdiv32_fs139_or0 ^ f_arrdiv32_fs140_xor0;
  assign f_arrdiv32_fs140_not1 = ~f_arrdiv32_fs140_xor0;
  assign f_arrdiv32_fs140_and1 = f_arrdiv32_fs140_not1 & f_arrdiv32_fs139_or0;
  assign f_arrdiv32_fs140_or0 = f_arrdiv32_fs140_and1 | f_arrdiv32_fs140_and0;
  assign f_arrdiv32_fs141_xor0 = f_arrdiv32_mux2to1105_xor0 ^ b[13];
  assign f_arrdiv32_fs141_not0 = ~f_arrdiv32_mux2to1105_xor0;
  assign f_arrdiv32_fs141_and0 = f_arrdiv32_fs141_not0 & b[13];
  assign f_arrdiv32_fs141_xor1 = f_arrdiv32_fs140_or0 ^ f_arrdiv32_fs141_xor0;
  assign f_arrdiv32_fs141_not1 = ~f_arrdiv32_fs141_xor0;
  assign f_arrdiv32_fs141_and1 = f_arrdiv32_fs141_not1 & f_arrdiv32_fs140_or0;
  assign f_arrdiv32_fs141_or0 = f_arrdiv32_fs141_and1 | f_arrdiv32_fs141_and0;
  assign f_arrdiv32_fs142_xor0 = f_arrdiv32_mux2to1106_xor0 ^ b[14];
  assign f_arrdiv32_fs142_not0 = ~f_arrdiv32_mux2to1106_xor0;
  assign f_arrdiv32_fs142_and0 = f_arrdiv32_fs142_not0 & b[14];
  assign f_arrdiv32_fs142_xor1 = f_arrdiv32_fs141_or0 ^ f_arrdiv32_fs142_xor0;
  assign f_arrdiv32_fs142_not1 = ~f_arrdiv32_fs142_xor0;
  assign f_arrdiv32_fs142_and1 = f_arrdiv32_fs142_not1 & f_arrdiv32_fs141_or0;
  assign f_arrdiv32_fs142_or0 = f_arrdiv32_fs142_and1 | f_arrdiv32_fs142_and0;
  assign f_arrdiv32_fs143_xor0 = f_arrdiv32_mux2to1107_xor0 ^ b[15];
  assign f_arrdiv32_fs143_not0 = ~f_arrdiv32_mux2to1107_xor0;
  assign f_arrdiv32_fs143_and0 = f_arrdiv32_fs143_not0 & b[15];
  assign f_arrdiv32_fs143_xor1 = f_arrdiv32_fs142_or0 ^ f_arrdiv32_fs143_xor0;
  assign f_arrdiv32_fs143_not1 = ~f_arrdiv32_fs143_xor0;
  assign f_arrdiv32_fs143_and1 = f_arrdiv32_fs143_not1 & f_arrdiv32_fs142_or0;
  assign f_arrdiv32_fs143_or0 = f_arrdiv32_fs143_and1 | f_arrdiv32_fs143_and0;
  assign f_arrdiv32_fs144_xor0 = f_arrdiv32_mux2to1108_xor0 ^ b[16];
  assign f_arrdiv32_fs144_not0 = ~f_arrdiv32_mux2to1108_xor0;
  assign f_arrdiv32_fs144_and0 = f_arrdiv32_fs144_not0 & b[16];
  assign f_arrdiv32_fs144_xor1 = f_arrdiv32_fs143_or0 ^ f_arrdiv32_fs144_xor0;
  assign f_arrdiv32_fs144_not1 = ~f_arrdiv32_fs144_xor0;
  assign f_arrdiv32_fs144_and1 = f_arrdiv32_fs144_not1 & f_arrdiv32_fs143_or0;
  assign f_arrdiv32_fs144_or0 = f_arrdiv32_fs144_and1 | f_arrdiv32_fs144_and0;
  assign f_arrdiv32_fs145_xor0 = f_arrdiv32_mux2to1109_xor0 ^ b[17];
  assign f_arrdiv32_fs145_not0 = ~f_arrdiv32_mux2to1109_xor0;
  assign f_arrdiv32_fs145_and0 = f_arrdiv32_fs145_not0 & b[17];
  assign f_arrdiv32_fs145_xor1 = f_arrdiv32_fs144_or0 ^ f_arrdiv32_fs145_xor0;
  assign f_arrdiv32_fs145_not1 = ~f_arrdiv32_fs145_xor0;
  assign f_arrdiv32_fs145_and1 = f_arrdiv32_fs145_not1 & f_arrdiv32_fs144_or0;
  assign f_arrdiv32_fs145_or0 = f_arrdiv32_fs145_and1 | f_arrdiv32_fs145_and0;
  assign f_arrdiv32_fs146_xor0 = f_arrdiv32_mux2to1110_xor0 ^ b[18];
  assign f_arrdiv32_fs146_not0 = ~f_arrdiv32_mux2to1110_xor0;
  assign f_arrdiv32_fs146_and0 = f_arrdiv32_fs146_not0 & b[18];
  assign f_arrdiv32_fs146_xor1 = f_arrdiv32_fs145_or0 ^ f_arrdiv32_fs146_xor0;
  assign f_arrdiv32_fs146_not1 = ~f_arrdiv32_fs146_xor0;
  assign f_arrdiv32_fs146_and1 = f_arrdiv32_fs146_not1 & f_arrdiv32_fs145_or0;
  assign f_arrdiv32_fs146_or0 = f_arrdiv32_fs146_and1 | f_arrdiv32_fs146_and0;
  assign f_arrdiv32_fs147_xor0 = f_arrdiv32_mux2to1111_xor0 ^ b[19];
  assign f_arrdiv32_fs147_not0 = ~f_arrdiv32_mux2to1111_xor0;
  assign f_arrdiv32_fs147_and0 = f_arrdiv32_fs147_not0 & b[19];
  assign f_arrdiv32_fs147_xor1 = f_arrdiv32_fs146_or0 ^ f_arrdiv32_fs147_xor0;
  assign f_arrdiv32_fs147_not1 = ~f_arrdiv32_fs147_xor0;
  assign f_arrdiv32_fs147_and1 = f_arrdiv32_fs147_not1 & f_arrdiv32_fs146_or0;
  assign f_arrdiv32_fs147_or0 = f_arrdiv32_fs147_and1 | f_arrdiv32_fs147_and0;
  assign f_arrdiv32_fs148_xor0 = f_arrdiv32_mux2to1112_xor0 ^ b[20];
  assign f_arrdiv32_fs148_not0 = ~f_arrdiv32_mux2to1112_xor0;
  assign f_arrdiv32_fs148_and0 = f_arrdiv32_fs148_not0 & b[20];
  assign f_arrdiv32_fs148_xor1 = f_arrdiv32_fs147_or0 ^ f_arrdiv32_fs148_xor0;
  assign f_arrdiv32_fs148_not1 = ~f_arrdiv32_fs148_xor0;
  assign f_arrdiv32_fs148_and1 = f_arrdiv32_fs148_not1 & f_arrdiv32_fs147_or0;
  assign f_arrdiv32_fs148_or0 = f_arrdiv32_fs148_and1 | f_arrdiv32_fs148_and0;
  assign f_arrdiv32_fs149_xor0 = f_arrdiv32_mux2to1113_xor0 ^ b[21];
  assign f_arrdiv32_fs149_not0 = ~f_arrdiv32_mux2to1113_xor0;
  assign f_arrdiv32_fs149_and0 = f_arrdiv32_fs149_not0 & b[21];
  assign f_arrdiv32_fs149_xor1 = f_arrdiv32_fs148_or0 ^ f_arrdiv32_fs149_xor0;
  assign f_arrdiv32_fs149_not1 = ~f_arrdiv32_fs149_xor0;
  assign f_arrdiv32_fs149_and1 = f_arrdiv32_fs149_not1 & f_arrdiv32_fs148_or0;
  assign f_arrdiv32_fs149_or0 = f_arrdiv32_fs149_and1 | f_arrdiv32_fs149_and0;
  assign f_arrdiv32_fs150_xor0 = f_arrdiv32_mux2to1114_xor0 ^ b[22];
  assign f_arrdiv32_fs150_not0 = ~f_arrdiv32_mux2to1114_xor0;
  assign f_arrdiv32_fs150_and0 = f_arrdiv32_fs150_not0 & b[22];
  assign f_arrdiv32_fs150_xor1 = f_arrdiv32_fs149_or0 ^ f_arrdiv32_fs150_xor0;
  assign f_arrdiv32_fs150_not1 = ~f_arrdiv32_fs150_xor0;
  assign f_arrdiv32_fs150_and1 = f_arrdiv32_fs150_not1 & f_arrdiv32_fs149_or0;
  assign f_arrdiv32_fs150_or0 = f_arrdiv32_fs150_and1 | f_arrdiv32_fs150_and0;
  assign f_arrdiv32_fs151_xor0 = f_arrdiv32_mux2to1115_xor0 ^ b[23];
  assign f_arrdiv32_fs151_not0 = ~f_arrdiv32_mux2to1115_xor0;
  assign f_arrdiv32_fs151_and0 = f_arrdiv32_fs151_not0 & b[23];
  assign f_arrdiv32_fs151_xor1 = f_arrdiv32_fs150_or0 ^ f_arrdiv32_fs151_xor0;
  assign f_arrdiv32_fs151_not1 = ~f_arrdiv32_fs151_xor0;
  assign f_arrdiv32_fs151_and1 = f_arrdiv32_fs151_not1 & f_arrdiv32_fs150_or0;
  assign f_arrdiv32_fs151_or0 = f_arrdiv32_fs151_and1 | f_arrdiv32_fs151_and0;
  assign f_arrdiv32_fs152_xor0 = f_arrdiv32_mux2to1116_xor0 ^ b[24];
  assign f_arrdiv32_fs152_not0 = ~f_arrdiv32_mux2to1116_xor0;
  assign f_arrdiv32_fs152_and0 = f_arrdiv32_fs152_not0 & b[24];
  assign f_arrdiv32_fs152_xor1 = f_arrdiv32_fs151_or0 ^ f_arrdiv32_fs152_xor0;
  assign f_arrdiv32_fs152_not1 = ~f_arrdiv32_fs152_xor0;
  assign f_arrdiv32_fs152_and1 = f_arrdiv32_fs152_not1 & f_arrdiv32_fs151_or0;
  assign f_arrdiv32_fs152_or0 = f_arrdiv32_fs152_and1 | f_arrdiv32_fs152_and0;
  assign f_arrdiv32_fs153_xor0 = f_arrdiv32_mux2to1117_xor0 ^ b[25];
  assign f_arrdiv32_fs153_not0 = ~f_arrdiv32_mux2to1117_xor0;
  assign f_arrdiv32_fs153_and0 = f_arrdiv32_fs153_not0 & b[25];
  assign f_arrdiv32_fs153_xor1 = f_arrdiv32_fs152_or0 ^ f_arrdiv32_fs153_xor0;
  assign f_arrdiv32_fs153_not1 = ~f_arrdiv32_fs153_xor0;
  assign f_arrdiv32_fs153_and1 = f_arrdiv32_fs153_not1 & f_arrdiv32_fs152_or0;
  assign f_arrdiv32_fs153_or0 = f_arrdiv32_fs153_and1 | f_arrdiv32_fs153_and0;
  assign f_arrdiv32_fs154_xor0 = f_arrdiv32_mux2to1118_xor0 ^ b[26];
  assign f_arrdiv32_fs154_not0 = ~f_arrdiv32_mux2to1118_xor0;
  assign f_arrdiv32_fs154_and0 = f_arrdiv32_fs154_not0 & b[26];
  assign f_arrdiv32_fs154_xor1 = f_arrdiv32_fs153_or0 ^ f_arrdiv32_fs154_xor0;
  assign f_arrdiv32_fs154_not1 = ~f_arrdiv32_fs154_xor0;
  assign f_arrdiv32_fs154_and1 = f_arrdiv32_fs154_not1 & f_arrdiv32_fs153_or0;
  assign f_arrdiv32_fs154_or0 = f_arrdiv32_fs154_and1 | f_arrdiv32_fs154_and0;
  assign f_arrdiv32_fs155_xor0 = f_arrdiv32_mux2to1119_xor0 ^ b[27];
  assign f_arrdiv32_fs155_not0 = ~f_arrdiv32_mux2to1119_xor0;
  assign f_arrdiv32_fs155_and0 = f_arrdiv32_fs155_not0 & b[27];
  assign f_arrdiv32_fs155_xor1 = f_arrdiv32_fs154_or0 ^ f_arrdiv32_fs155_xor0;
  assign f_arrdiv32_fs155_not1 = ~f_arrdiv32_fs155_xor0;
  assign f_arrdiv32_fs155_and1 = f_arrdiv32_fs155_not1 & f_arrdiv32_fs154_or0;
  assign f_arrdiv32_fs155_or0 = f_arrdiv32_fs155_and1 | f_arrdiv32_fs155_and0;
  assign f_arrdiv32_fs156_xor0 = f_arrdiv32_mux2to1120_xor0 ^ b[28];
  assign f_arrdiv32_fs156_not0 = ~f_arrdiv32_mux2to1120_xor0;
  assign f_arrdiv32_fs156_and0 = f_arrdiv32_fs156_not0 & b[28];
  assign f_arrdiv32_fs156_xor1 = f_arrdiv32_fs155_or0 ^ f_arrdiv32_fs156_xor0;
  assign f_arrdiv32_fs156_not1 = ~f_arrdiv32_fs156_xor0;
  assign f_arrdiv32_fs156_and1 = f_arrdiv32_fs156_not1 & f_arrdiv32_fs155_or0;
  assign f_arrdiv32_fs156_or0 = f_arrdiv32_fs156_and1 | f_arrdiv32_fs156_and0;
  assign f_arrdiv32_fs157_xor0 = f_arrdiv32_mux2to1121_xor0 ^ b[29];
  assign f_arrdiv32_fs157_not0 = ~f_arrdiv32_mux2to1121_xor0;
  assign f_arrdiv32_fs157_and0 = f_arrdiv32_fs157_not0 & b[29];
  assign f_arrdiv32_fs157_xor1 = f_arrdiv32_fs156_or0 ^ f_arrdiv32_fs157_xor0;
  assign f_arrdiv32_fs157_not1 = ~f_arrdiv32_fs157_xor0;
  assign f_arrdiv32_fs157_and1 = f_arrdiv32_fs157_not1 & f_arrdiv32_fs156_or0;
  assign f_arrdiv32_fs157_or0 = f_arrdiv32_fs157_and1 | f_arrdiv32_fs157_and0;
  assign f_arrdiv32_fs158_xor0 = f_arrdiv32_mux2to1122_xor0 ^ b[30];
  assign f_arrdiv32_fs158_not0 = ~f_arrdiv32_mux2to1122_xor0;
  assign f_arrdiv32_fs158_and0 = f_arrdiv32_fs158_not0 & b[30];
  assign f_arrdiv32_fs158_xor1 = f_arrdiv32_fs157_or0 ^ f_arrdiv32_fs158_xor0;
  assign f_arrdiv32_fs158_not1 = ~f_arrdiv32_fs158_xor0;
  assign f_arrdiv32_fs158_and1 = f_arrdiv32_fs158_not1 & f_arrdiv32_fs157_or0;
  assign f_arrdiv32_fs158_or0 = f_arrdiv32_fs158_and1 | f_arrdiv32_fs158_and0;
  assign f_arrdiv32_fs159_xor0 = f_arrdiv32_mux2to1123_xor0 ^ b[31];
  assign f_arrdiv32_fs159_not0 = ~f_arrdiv32_mux2to1123_xor0;
  assign f_arrdiv32_fs159_and0 = f_arrdiv32_fs159_not0 & b[31];
  assign f_arrdiv32_fs159_xor1 = f_arrdiv32_fs158_or0 ^ f_arrdiv32_fs159_xor0;
  assign f_arrdiv32_fs159_not1 = ~f_arrdiv32_fs159_xor0;
  assign f_arrdiv32_fs159_and1 = f_arrdiv32_fs159_not1 & f_arrdiv32_fs158_or0;
  assign f_arrdiv32_fs159_or0 = f_arrdiv32_fs159_and1 | f_arrdiv32_fs159_and0;
  assign f_arrdiv32_mux2to1124_and0 = a[27] & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1124_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1124_and1 = f_arrdiv32_fs128_xor0 & f_arrdiv32_mux2to1124_not0;
  assign f_arrdiv32_mux2to1124_xor0 = f_arrdiv32_mux2to1124_and0 ^ f_arrdiv32_mux2to1124_and1;
  assign f_arrdiv32_mux2to1125_and0 = f_arrdiv32_mux2to193_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1125_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1125_and1 = f_arrdiv32_fs129_xor1 & f_arrdiv32_mux2to1125_not0;
  assign f_arrdiv32_mux2to1125_xor0 = f_arrdiv32_mux2to1125_and0 ^ f_arrdiv32_mux2to1125_and1;
  assign f_arrdiv32_mux2to1126_and0 = f_arrdiv32_mux2to194_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1126_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1126_and1 = f_arrdiv32_fs130_xor1 & f_arrdiv32_mux2to1126_not0;
  assign f_arrdiv32_mux2to1126_xor0 = f_arrdiv32_mux2to1126_and0 ^ f_arrdiv32_mux2to1126_and1;
  assign f_arrdiv32_mux2to1127_and0 = f_arrdiv32_mux2to195_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1127_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1127_and1 = f_arrdiv32_fs131_xor1 & f_arrdiv32_mux2to1127_not0;
  assign f_arrdiv32_mux2to1127_xor0 = f_arrdiv32_mux2to1127_and0 ^ f_arrdiv32_mux2to1127_and1;
  assign f_arrdiv32_mux2to1128_and0 = f_arrdiv32_mux2to196_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1128_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1128_and1 = f_arrdiv32_fs132_xor1 & f_arrdiv32_mux2to1128_not0;
  assign f_arrdiv32_mux2to1128_xor0 = f_arrdiv32_mux2to1128_and0 ^ f_arrdiv32_mux2to1128_and1;
  assign f_arrdiv32_mux2to1129_and0 = f_arrdiv32_mux2to197_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1129_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1129_and1 = f_arrdiv32_fs133_xor1 & f_arrdiv32_mux2to1129_not0;
  assign f_arrdiv32_mux2to1129_xor0 = f_arrdiv32_mux2to1129_and0 ^ f_arrdiv32_mux2to1129_and1;
  assign f_arrdiv32_mux2to1130_and0 = f_arrdiv32_mux2to198_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1130_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1130_and1 = f_arrdiv32_fs134_xor1 & f_arrdiv32_mux2to1130_not0;
  assign f_arrdiv32_mux2to1130_xor0 = f_arrdiv32_mux2to1130_and0 ^ f_arrdiv32_mux2to1130_and1;
  assign f_arrdiv32_mux2to1131_and0 = f_arrdiv32_mux2to199_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1131_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1131_and1 = f_arrdiv32_fs135_xor1 & f_arrdiv32_mux2to1131_not0;
  assign f_arrdiv32_mux2to1131_xor0 = f_arrdiv32_mux2to1131_and0 ^ f_arrdiv32_mux2to1131_and1;
  assign f_arrdiv32_mux2to1132_and0 = f_arrdiv32_mux2to1100_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1132_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1132_and1 = f_arrdiv32_fs136_xor1 & f_arrdiv32_mux2to1132_not0;
  assign f_arrdiv32_mux2to1132_xor0 = f_arrdiv32_mux2to1132_and0 ^ f_arrdiv32_mux2to1132_and1;
  assign f_arrdiv32_mux2to1133_and0 = f_arrdiv32_mux2to1101_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1133_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1133_and1 = f_arrdiv32_fs137_xor1 & f_arrdiv32_mux2to1133_not0;
  assign f_arrdiv32_mux2to1133_xor0 = f_arrdiv32_mux2to1133_and0 ^ f_arrdiv32_mux2to1133_and1;
  assign f_arrdiv32_mux2to1134_and0 = f_arrdiv32_mux2to1102_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1134_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1134_and1 = f_arrdiv32_fs138_xor1 & f_arrdiv32_mux2to1134_not0;
  assign f_arrdiv32_mux2to1134_xor0 = f_arrdiv32_mux2to1134_and0 ^ f_arrdiv32_mux2to1134_and1;
  assign f_arrdiv32_mux2to1135_and0 = f_arrdiv32_mux2to1103_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1135_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1135_and1 = f_arrdiv32_fs139_xor1 & f_arrdiv32_mux2to1135_not0;
  assign f_arrdiv32_mux2to1135_xor0 = f_arrdiv32_mux2to1135_and0 ^ f_arrdiv32_mux2to1135_and1;
  assign f_arrdiv32_mux2to1136_and0 = f_arrdiv32_mux2to1104_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1136_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1136_and1 = f_arrdiv32_fs140_xor1 & f_arrdiv32_mux2to1136_not0;
  assign f_arrdiv32_mux2to1136_xor0 = f_arrdiv32_mux2to1136_and0 ^ f_arrdiv32_mux2to1136_and1;
  assign f_arrdiv32_mux2to1137_and0 = f_arrdiv32_mux2to1105_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1137_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1137_and1 = f_arrdiv32_fs141_xor1 & f_arrdiv32_mux2to1137_not0;
  assign f_arrdiv32_mux2to1137_xor0 = f_arrdiv32_mux2to1137_and0 ^ f_arrdiv32_mux2to1137_and1;
  assign f_arrdiv32_mux2to1138_and0 = f_arrdiv32_mux2to1106_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1138_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1138_and1 = f_arrdiv32_fs142_xor1 & f_arrdiv32_mux2to1138_not0;
  assign f_arrdiv32_mux2to1138_xor0 = f_arrdiv32_mux2to1138_and0 ^ f_arrdiv32_mux2to1138_and1;
  assign f_arrdiv32_mux2to1139_and0 = f_arrdiv32_mux2to1107_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1139_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1139_and1 = f_arrdiv32_fs143_xor1 & f_arrdiv32_mux2to1139_not0;
  assign f_arrdiv32_mux2to1139_xor0 = f_arrdiv32_mux2to1139_and0 ^ f_arrdiv32_mux2to1139_and1;
  assign f_arrdiv32_mux2to1140_and0 = f_arrdiv32_mux2to1108_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1140_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1140_and1 = f_arrdiv32_fs144_xor1 & f_arrdiv32_mux2to1140_not0;
  assign f_arrdiv32_mux2to1140_xor0 = f_arrdiv32_mux2to1140_and0 ^ f_arrdiv32_mux2to1140_and1;
  assign f_arrdiv32_mux2to1141_and0 = f_arrdiv32_mux2to1109_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1141_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1141_and1 = f_arrdiv32_fs145_xor1 & f_arrdiv32_mux2to1141_not0;
  assign f_arrdiv32_mux2to1141_xor0 = f_arrdiv32_mux2to1141_and0 ^ f_arrdiv32_mux2to1141_and1;
  assign f_arrdiv32_mux2to1142_and0 = f_arrdiv32_mux2to1110_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1142_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1142_and1 = f_arrdiv32_fs146_xor1 & f_arrdiv32_mux2to1142_not0;
  assign f_arrdiv32_mux2to1142_xor0 = f_arrdiv32_mux2to1142_and0 ^ f_arrdiv32_mux2to1142_and1;
  assign f_arrdiv32_mux2to1143_and0 = f_arrdiv32_mux2to1111_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1143_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1143_and1 = f_arrdiv32_fs147_xor1 & f_arrdiv32_mux2to1143_not0;
  assign f_arrdiv32_mux2to1143_xor0 = f_arrdiv32_mux2to1143_and0 ^ f_arrdiv32_mux2to1143_and1;
  assign f_arrdiv32_mux2to1144_and0 = f_arrdiv32_mux2to1112_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1144_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1144_and1 = f_arrdiv32_fs148_xor1 & f_arrdiv32_mux2to1144_not0;
  assign f_arrdiv32_mux2to1144_xor0 = f_arrdiv32_mux2to1144_and0 ^ f_arrdiv32_mux2to1144_and1;
  assign f_arrdiv32_mux2to1145_and0 = f_arrdiv32_mux2to1113_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1145_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1145_and1 = f_arrdiv32_fs149_xor1 & f_arrdiv32_mux2to1145_not0;
  assign f_arrdiv32_mux2to1145_xor0 = f_arrdiv32_mux2to1145_and0 ^ f_arrdiv32_mux2to1145_and1;
  assign f_arrdiv32_mux2to1146_and0 = f_arrdiv32_mux2to1114_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1146_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1146_and1 = f_arrdiv32_fs150_xor1 & f_arrdiv32_mux2to1146_not0;
  assign f_arrdiv32_mux2to1146_xor0 = f_arrdiv32_mux2to1146_and0 ^ f_arrdiv32_mux2to1146_and1;
  assign f_arrdiv32_mux2to1147_and0 = f_arrdiv32_mux2to1115_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1147_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1147_and1 = f_arrdiv32_fs151_xor1 & f_arrdiv32_mux2to1147_not0;
  assign f_arrdiv32_mux2to1147_xor0 = f_arrdiv32_mux2to1147_and0 ^ f_arrdiv32_mux2to1147_and1;
  assign f_arrdiv32_mux2to1148_and0 = f_arrdiv32_mux2to1116_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1148_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1148_and1 = f_arrdiv32_fs152_xor1 & f_arrdiv32_mux2to1148_not0;
  assign f_arrdiv32_mux2to1148_xor0 = f_arrdiv32_mux2to1148_and0 ^ f_arrdiv32_mux2to1148_and1;
  assign f_arrdiv32_mux2to1149_and0 = f_arrdiv32_mux2to1117_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1149_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1149_and1 = f_arrdiv32_fs153_xor1 & f_arrdiv32_mux2to1149_not0;
  assign f_arrdiv32_mux2to1149_xor0 = f_arrdiv32_mux2to1149_and0 ^ f_arrdiv32_mux2to1149_and1;
  assign f_arrdiv32_mux2to1150_and0 = f_arrdiv32_mux2to1118_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1150_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1150_and1 = f_arrdiv32_fs154_xor1 & f_arrdiv32_mux2to1150_not0;
  assign f_arrdiv32_mux2to1150_xor0 = f_arrdiv32_mux2to1150_and0 ^ f_arrdiv32_mux2to1150_and1;
  assign f_arrdiv32_mux2to1151_and0 = f_arrdiv32_mux2to1119_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1151_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1151_and1 = f_arrdiv32_fs155_xor1 & f_arrdiv32_mux2to1151_not0;
  assign f_arrdiv32_mux2to1151_xor0 = f_arrdiv32_mux2to1151_and0 ^ f_arrdiv32_mux2to1151_and1;
  assign f_arrdiv32_mux2to1152_and0 = f_arrdiv32_mux2to1120_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1152_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1152_and1 = f_arrdiv32_fs156_xor1 & f_arrdiv32_mux2to1152_not0;
  assign f_arrdiv32_mux2to1152_xor0 = f_arrdiv32_mux2to1152_and0 ^ f_arrdiv32_mux2to1152_and1;
  assign f_arrdiv32_mux2to1153_and0 = f_arrdiv32_mux2to1121_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1153_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1153_and1 = f_arrdiv32_fs157_xor1 & f_arrdiv32_mux2to1153_not0;
  assign f_arrdiv32_mux2to1153_xor0 = f_arrdiv32_mux2to1153_and0 ^ f_arrdiv32_mux2to1153_and1;
  assign f_arrdiv32_mux2to1154_and0 = f_arrdiv32_mux2to1122_xor0 & f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1154_not0 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_mux2to1154_and1 = f_arrdiv32_fs158_xor1 & f_arrdiv32_mux2to1154_not0;
  assign f_arrdiv32_mux2to1154_xor0 = f_arrdiv32_mux2to1154_and0 ^ f_arrdiv32_mux2to1154_and1;
  assign f_arrdiv32_not4 = ~f_arrdiv32_fs159_or0;
  assign f_arrdiv32_fs160_xor0 = a[26] ^ b[0];
  assign f_arrdiv32_fs160_not0 = ~a[26];
  assign f_arrdiv32_fs160_and0 = f_arrdiv32_fs160_not0 & b[0];
  assign f_arrdiv32_fs160_not1 = ~f_arrdiv32_fs160_xor0;
  assign f_arrdiv32_fs161_xor0 = f_arrdiv32_mux2to1124_xor0 ^ b[1];
  assign f_arrdiv32_fs161_not0 = ~f_arrdiv32_mux2to1124_xor0;
  assign f_arrdiv32_fs161_and0 = f_arrdiv32_fs161_not0 & b[1];
  assign f_arrdiv32_fs161_xor1 = f_arrdiv32_fs160_and0 ^ f_arrdiv32_fs161_xor0;
  assign f_arrdiv32_fs161_not1 = ~f_arrdiv32_fs161_xor0;
  assign f_arrdiv32_fs161_and1 = f_arrdiv32_fs161_not1 & f_arrdiv32_fs160_and0;
  assign f_arrdiv32_fs161_or0 = f_arrdiv32_fs161_and1 | f_arrdiv32_fs161_and0;
  assign f_arrdiv32_fs162_xor0 = f_arrdiv32_mux2to1125_xor0 ^ b[2];
  assign f_arrdiv32_fs162_not0 = ~f_arrdiv32_mux2to1125_xor0;
  assign f_arrdiv32_fs162_and0 = f_arrdiv32_fs162_not0 & b[2];
  assign f_arrdiv32_fs162_xor1 = f_arrdiv32_fs161_or0 ^ f_arrdiv32_fs162_xor0;
  assign f_arrdiv32_fs162_not1 = ~f_arrdiv32_fs162_xor0;
  assign f_arrdiv32_fs162_and1 = f_arrdiv32_fs162_not1 & f_arrdiv32_fs161_or0;
  assign f_arrdiv32_fs162_or0 = f_arrdiv32_fs162_and1 | f_arrdiv32_fs162_and0;
  assign f_arrdiv32_fs163_xor0 = f_arrdiv32_mux2to1126_xor0 ^ b[3];
  assign f_arrdiv32_fs163_not0 = ~f_arrdiv32_mux2to1126_xor0;
  assign f_arrdiv32_fs163_and0 = f_arrdiv32_fs163_not0 & b[3];
  assign f_arrdiv32_fs163_xor1 = f_arrdiv32_fs162_or0 ^ f_arrdiv32_fs163_xor0;
  assign f_arrdiv32_fs163_not1 = ~f_arrdiv32_fs163_xor0;
  assign f_arrdiv32_fs163_and1 = f_arrdiv32_fs163_not1 & f_arrdiv32_fs162_or0;
  assign f_arrdiv32_fs163_or0 = f_arrdiv32_fs163_and1 | f_arrdiv32_fs163_and0;
  assign f_arrdiv32_fs164_xor0 = f_arrdiv32_mux2to1127_xor0 ^ b[4];
  assign f_arrdiv32_fs164_not0 = ~f_arrdiv32_mux2to1127_xor0;
  assign f_arrdiv32_fs164_and0 = f_arrdiv32_fs164_not0 & b[4];
  assign f_arrdiv32_fs164_xor1 = f_arrdiv32_fs163_or0 ^ f_arrdiv32_fs164_xor0;
  assign f_arrdiv32_fs164_not1 = ~f_arrdiv32_fs164_xor0;
  assign f_arrdiv32_fs164_and1 = f_arrdiv32_fs164_not1 & f_arrdiv32_fs163_or0;
  assign f_arrdiv32_fs164_or0 = f_arrdiv32_fs164_and1 | f_arrdiv32_fs164_and0;
  assign f_arrdiv32_fs165_xor0 = f_arrdiv32_mux2to1128_xor0 ^ b[5];
  assign f_arrdiv32_fs165_not0 = ~f_arrdiv32_mux2to1128_xor0;
  assign f_arrdiv32_fs165_and0 = f_arrdiv32_fs165_not0 & b[5];
  assign f_arrdiv32_fs165_xor1 = f_arrdiv32_fs164_or0 ^ f_arrdiv32_fs165_xor0;
  assign f_arrdiv32_fs165_not1 = ~f_arrdiv32_fs165_xor0;
  assign f_arrdiv32_fs165_and1 = f_arrdiv32_fs165_not1 & f_arrdiv32_fs164_or0;
  assign f_arrdiv32_fs165_or0 = f_arrdiv32_fs165_and1 | f_arrdiv32_fs165_and0;
  assign f_arrdiv32_fs166_xor0 = f_arrdiv32_mux2to1129_xor0 ^ b[6];
  assign f_arrdiv32_fs166_not0 = ~f_arrdiv32_mux2to1129_xor0;
  assign f_arrdiv32_fs166_and0 = f_arrdiv32_fs166_not0 & b[6];
  assign f_arrdiv32_fs166_xor1 = f_arrdiv32_fs165_or0 ^ f_arrdiv32_fs166_xor0;
  assign f_arrdiv32_fs166_not1 = ~f_arrdiv32_fs166_xor0;
  assign f_arrdiv32_fs166_and1 = f_arrdiv32_fs166_not1 & f_arrdiv32_fs165_or0;
  assign f_arrdiv32_fs166_or0 = f_arrdiv32_fs166_and1 | f_arrdiv32_fs166_and0;
  assign f_arrdiv32_fs167_xor0 = f_arrdiv32_mux2to1130_xor0 ^ b[7];
  assign f_arrdiv32_fs167_not0 = ~f_arrdiv32_mux2to1130_xor0;
  assign f_arrdiv32_fs167_and0 = f_arrdiv32_fs167_not0 & b[7];
  assign f_arrdiv32_fs167_xor1 = f_arrdiv32_fs166_or0 ^ f_arrdiv32_fs167_xor0;
  assign f_arrdiv32_fs167_not1 = ~f_arrdiv32_fs167_xor0;
  assign f_arrdiv32_fs167_and1 = f_arrdiv32_fs167_not1 & f_arrdiv32_fs166_or0;
  assign f_arrdiv32_fs167_or0 = f_arrdiv32_fs167_and1 | f_arrdiv32_fs167_and0;
  assign f_arrdiv32_fs168_xor0 = f_arrdiv32_mux2to1131_xor0 ^ b[8];
  assign f_arrdiv32_fs168_not0 = ~f_arrdiv32_mux2to1131_xor0;
  assign f_arrdiv32_fs168_and0 = f_arrdiv32_fs168_not0 & b[8];
  assign f_arrdiv32_fs168_xor1 = f_arrdiv32_fs167_or0 ^ f_arrdiv32_fs168_xor0;
  assign f_arrdiv32_fs168_not1 = ~f_arrdiv32_fs168_xor0;
  assign f_arrdiv32_fs168_and1 = f_arrdiv32_fs168_not1 & f_arrdiv32_fs167_or0;
  assign f_arrdiv32_fs168_or0 = f_arrdiv32_fs168_and1 | f_arrdiv32_fs168_and0;
  assign f_arrdiv32_fs169_xor0 = f_arrdiv32_mux2to1132_xor0 ^ b[9];
  assign f_arrdiv32_fs169_not0 = ~f_arrdiv32_mux2to1132_xor0;
  assign f_arrdiv32_fs169_and0 = f_arrdiv32_fs169_not0 & b[9];
  assign f_arrdiv32_fs169_xor1 = f_arrdiv32_fs168_or0 ^ f_arrdiv32_fs169_xor0;
  assign f_arrdiv32_fs169_not1 = ~f_arrdiv32_fs169_xor0;
  assign f_arrdiv32_fs169_and1 = f_arrdiv32_fs169_not1 & f_arrdiv32_fs168_or0;
  assign f_arrdiv32_fs169_or0 = f_arrdiv32_fs169_and1 | f_arrdiv32_fs169_and0;
  assign f_arrdiv32_fs170_xor0 = f_arrdiv32_mux2to1133_xor0 ^ b[10];
  assign f_arrdiv32_fs170_not0 = ~f_arrdiv32_mux2to1133_xor0;
  assign f_arrdiv32_fs170_and0 = f_arrdiv32_fs170_not0 & b[10];
  assign f_arrdiv32_fs170_xor1 = f_arrdiv32_fs169_or0 ^ f_arrdiv32_fs170_xor0;
  assign f_arrdiv32_fs170_not1 = ~f_arrdiv32_fs170_xor0;
  assign f_arrdiv32_fs170_and1 = f_arrdiv32_fs170_not1 & f_arrdiv32_fs169_or0;
  assign f_arrdiv32_fs170_or0 = f_arrdiv32_fs170_and1 | f_arrdiv32_fs170_and0;
  assign f_arrdiv32_fs171_xor0 = f_arrdiv32_mux2to1134_xor0 ^ b[11];
  assign f_arrdiv32_fs171_not0 = ~f_arrdiv32_mux2to1134_xor0;
  assign f_arrdiv32_fs171_and0 = f_arrdiv32_fs171_not0 & b[11];
  assign f_arrdiv32_fs171_xor1 = f_arrdiv32_fs170_or0 ^ f_arrdiv32_fs171_xor0;
  assign f_arrdiv32_fs171_not1 = ~f_arrdiv32_fs171_xor0;
  assign f_arrdiv32_fs171_and1 = f_arrdiv32_fs171_not1 & f_arrdiv32_fs170_or0;
  assign f_arrdiv32_fs171_or0 = f_arrdiv32_fs171_and1 | f_arrdiv32_fs171_and0;
  assign f_arrdiv32_fs172_xor0 = f_arrdiv32_mux2to1135_xor0 ^ b[12];
  assign f_arrdiv32_fs172_not0 = ~f_arrdiv32_mux2to1135_xor0;
  assign f_arrdiv32_fs172_and0 = f_arrdiv32_fs172_not0 & b[12];
  assign f_arrdiv32_fs172_xor1 = f_arrdiv32_fs171_or0 ^ f_arrdiv32_fs172_xor0;
  assign f_arrdiv32_fs172_not1 = ~f_arrdiv32_fs172_xor0;
  assign f_arrdiv32_fs172_and1 = f_arrdiv32_fs172_not1 & f_arrdiv32_fs171_or0;
  assign f_arrdiv32_fs172_or0 = f_arrdiv32_fs172_and1 | f_arrdiv32_fs172_and0;
  assign f_arrdiv32_fs173_xor0 = f_arrdiv32_mux2to1136_xor0 ^ b[13];
  assign f_arrdiv32_fs173_not0 = ~f_arrdiv32_mux2to1136_xor0;
  assign f_arrdiv32_fs173_and0 = f_arrdiv32_fs173_not0 & b[13];
  assign f_arrdiv32_fs173_xor1 = f_arrdiv32_fs172_or0 ^ f_arrdiv32_fs173_xor0;
  assign f_arrdiv32_fs173_not1 = ~f_arrdiv32_fs173_xor0;
  assign f_arrdiv32_fs173_and1 = f_arrdiv32_fs173_not1 & f_arrdiv32_fs172_or0;
  assign f_arrdiv32_fs173_or0 = f_arrdiv32_fs173_and1 | f_arrdiv32_fs173_and0;
  assign f_arrdiv32_fs174_xor0 = f_arrdiv32_mux2to1137_xor0 ^ b[14];
  assign f_arrdiv32_fs174_not0 = ~f_arrdiv32_mux2to1137_xor0;
  assign f_arrdiv32_fs174_and0 = f_arrdiv32_fs174_not0 & b[14];
  assign f_arrdiv32_fs174_xor1 = f_arrdiv32_fs173_or0 ^ f_arrdiv32_fs174_xor0;
  assign f_arrdiv32_fs174_not1 = ~f_arrdiv32_fs174_xor0;
  assign f_arrdiv32_fs174_and1 = f_arrdiv32_fs174_not1 & f_arrdiv32_fs173_or0;
  assign f_arrdiv32_fs174_or0 = f_arrdiv32_fs174_and1 | f_arrdiv32_fs174_and0;
  assign f_arrdiv32_fs175_xor0 = f_arrdiv32_mux2to1138_xor0 ^ b[15];
  assign f_arrdiv32_fs175_not0 = ~f_arrdiv32_mux2to1138_xor0;
  assign f_arrdiv32_fs175_and0 = f_arrdiv32_fs175_not0 & b[15];
  assign f_arrdiv32_fs175_xor1 = f_arrdiv32_fs174_or0 ^ f_arrdiv32_fs175_xor0;
  assign f_arrdiv32_fs175_not1 = ~f_arrdiv32_fs175_xor0;
  assign f_arrdiv32_fs175_and1 = f_arrdiv32_fs175_not1 & f_arrdiv32_fs174_or0;
  assign f_arrdiv32_fs175_or0 = f_arrdiv32_fs175_and1 | f_arrdiv32_fs175_and0;
  assign f_arrdiv32_fs176_xor0 = f_arrdiv32_mux2to1139_xor0 ^ b[16];
  assign f_arrdiv32_fs176_not0 = ~f_arrdiv32_mux2to1139_xor0;
  assign f_arrdiv32_fs176_and0 = f_arrdiv32_fs176_not0 & b[16];
  assign f_arrdiv32_fs176_xor1 = f_arrdiv32_fs175_or0 ^ f_arrdiv32_fs176_xor0;
  assign f_arrdiv32_fs176_not1 = ~f_arrdiv32_fs176_xor0;
  assign f_arrdiv32_fs176_and1 = f_arrdiv32_fs176_not1 & f_arrdiv32_fs175_or0;
  assign f_arrdiv32_fs176_or0 = f_arrdiv32_fs176_and1 | f_arrdiv32_fs176_and0;
  assign f_arrdiv32_fs177_xor0 = f_arrdiv32_mux2to1140_xor0 ^ b[17];
  assign f_arrdiv32_fs177_not0 = ~f_arrdiv32_mux2to1140_xor0;
  assign f_arrdiv32_fs177_and0 = f_arrdiv32_fs177_not0 & b[17];
  assign f_arrdiv32_fs177_xor1 = f_arrdiv32_fs176_or0 ^ f_arrdiv32_fs177_xor0;
  assign f_arrdiv32_fs177_not1 = ~f_arrdiv32_fs177_xor0;
  assign f_arrdiv32_fs177_and1 = f_arrdiv32_fs177_not1 & f_arrdiv32_fs176_or0;
  assign f_arrdiv32_fs177_or0 = f_arrdiv32_fs177_and1 | f_arrdiv32_fs177_and0;
  assign f_arrdiv32_fs178_xor0 = f_arrdiv32_mux2to1141_xor0 ^ b[18];
  assign f_arrdiv32_fs178_not0 = ~f_arrdiv32_mux2to1141_xor0;
  assign f_arrdiv32_fs178_and0 = f_arrdiv32_fs178_not0 & b[18];
  assign f_arrdiv32_fs178_xor1 = f_arrdiv32_fs177_or0 ^ f_arrdiv32_fs178_xor0;
  assign f_arrdiv32_fs178_not1 = ~f_arrdiv32_fs178_xor0;
  assign f_arrdiv32_fs178_and1 = f_arrdiv32_fs178_not1 & f_arrdiv32_fs177_or0;
  assign f_arrdiv32_fs178_or0 = f_arrdiv32_fs178_and1 | f_arrdiv32_fs178_and0;
  assign f_arrdiv32_fs179_xor0 = f_arrdiv32_mux2to1142_xor0 ^ b[19];
  assign f_arrdiv32_fs179_not0 = ~f_arrdiv32_mux2to1142_xor0;
  assign f_arrdiv32_fs179_and0 = f_arrdiv32_fs179_not0 & b[19];
  assign f_arrdiv32_fs179_xor1 = f_arrdiv32_fs178_or0 ^ f_arrdiv32_fs179_xor0;
  assign f_arrdiv32_fs179_not1 = ~f_arrdiv32_fs179_xor0;
  assign f_arrdiv32_fs179_and1 = f_arrdiv32_fs179_not1 & f_arrdiv32_fs178_or0;
  assign f_arrdiv32_fs179_or0 = f_arrdiv32_fs179_and1 | f_arrdiv32_fs179_and0;
  assign f_arrdiv32_fs180_xor0 = f_arrdiv32_mux2to1143_xor0 ^ b[20];
  assign f_arrdiv32_fs180_not0 = ~f_arrdiv32_mux2to1143_xor0;
  assign f_arrdiv32_fs180_and0 = f_arrdiv32_fs180_not0 & b[20];
  assign f_arrdiv32_fs180_xor1 = f_arrdiv32_fs179_or0 ^ f_arrdiv32_fs180_xor0;
  assign f_arrdiv32_fs180_not1 = ~f_arrdiv32_fs180_xor0;
  assign f_arrdiv32_fs180_and1 = f_arrdiv32_fs180_not1 & f_arrdiv32_fs179_or0;
  assign f_arrdiv32_fs180_or0 = f_arrdiv32_fs180_and1 | f_arrdiv32_fs180_and0;
  assign f_arrdiv32_fs181_xor0 = f_arrdiv32_mux2to1144_xor0 ^ b[21];
  assign f_arrdiv32_fs181_not0 = ~f_arrdiv32_mux2to1144_xor0;
  assign f_arrdiv32_fs181_and0 = f_arrdiv32_fs181_not0 & b[21];
  assign f_arrdiv32_fs181_xor1 = f_arrdiv32_fs180_or0 ^ f_arrdiv32_fs181_xor0;
  assign f_arrdiv32_fs181_not1 = ~f_arrdiv32_fs181_xor0;
  assign f_arrdiv32_fs181_and1 = f_arrdiv32_fs181_not1 & f_arrdiv32_fs180_or0;
  assign f_arrdiv32_fs181_or0 = f_arrdiv32_fs181_and1 | f_arrdiv32_fs181_and0;
  assign f_arrdiv32_fs182_xor0 = f_arrdiv32_mux2to1145_xor0 ^ b[22];
  assign f_arrdiv32_fs182_not0 = ~f_arrdiv32_mux2to1145_xor0;
  assign f_arrdiv32_fs182_and0 = f_arrdiv32_fs182_not0 & b[22];
  assign f_arrdiv32_fs182_xor1 = f_arrdiv32_fs181_or0 ^ f_arrdiv32_fs182_xor0;
  assign f_arrdiv32_fs182_not1 = ~f_arrdiv32_fs182_xor0;
  assign f_arrdiv32_fs182_and1 = f_arrdiv32_fs182_not1 & f_arrdiv32_fs181_or0;
  assign f_arrdiv32_fs182_or0 = f_arrdiv32_fs182_and1 | f_arrdiv32_fs182_and0;
  assign f_arrdiv32_fs183_xor0 = f_arrdiv32_mux2to1146_xor0 ^ b[23];
  assign f_arrdiv32_fs183_not0 = ~f_arrdiv32_mux2to1146_xor0;
  assign f_arrdiv32_fs183_and0 = f_arrdiv32_fs183_not0 & b[23];
  assign f_arrdiv32_fs183_xor1 = f_arrdiv32_fs182_or0 ^ f_arrdiv32_fs183_xor0;
  assign f_arrdiv32_fs183_not1 = ~f_arrdiv32_fs183_xor0;
  assign f_arrdiv32_fs183_and1 = f_arrdiv32_fs183_not1 & f_arrdiv32_fs182_or0;
  assign f_arrdiv32_fs183_or0 = f_arrdiv32_fs183_and1 | f_arrdiv32_fs183_and0;
  assign f_arrdiv32_fs184_xor0 = f_arrdiv32_mux2to1147_xor0 ^ b[24];
  assign f_arrdiv32_fs184_not0 = ~f_arrdiv32_mux2to1147_xor0;
  assign f_arrdiv32_fs184_and0 = f_arrdiv32_fs184_not0 & b[24];
  assign f_arrdiv32_fs184_xor1 = f_arrdiv32_fs183_or0 ^ f_arrdiv32_fs184_xor0;
  assign f_arrdiv32_fs184_not1 = ~f_arrdiv32_fs184_xor0;
  assign f_arrdiv32_fs184_and1 = f_arrdiv32_fs184_not1 & f_arrdiv32_fs183_or0;
  assign f_arrdiv32_fs184_or0 = f_arrdiv32_fs184_and1 | f_arrdiv32_fs184_and0;
  assign f_arrdiv32_fs185_xor0 = f_arrdiv32_mux2to1148_xor0 ^ b[25];
  assign f_arrdiv32_fs185_not0 = ~f_arrdiv32_mux2to1148_xor0;
  assign f_arrdiv32_fs185_and0 = f_arrdiv32_fs185_not0 & b[25];
  assign f_arrdiv32_fs185_xor1 = f_arrdiv32_fs184_or0 ^ f_arrdiv32_fs185_xor0;
  assign f_arrdiv32_fs185_not1 = ~f_arrdiv32_fs185_xor0;
  assign f_arrdiv32_fs185_and1 = f_arrdiv32_fs185_not1 & f_arrdiv32_fs184_or0;
  assign f_arrdiv32_fs185_or0 = f_arrdiv32_fs185_and1 | f_arrdiv32_fs185_and0;
  assign f_arrdiv32_fs186_xor0 = f_arrdiv32_mux2to1149_xor0 ^ b[26];
  assign f_arrdiv32_fs186_not0 = ~f_arrdiv32_mux2to1149_xor0;
  assign f_arrdiv32_fs186_and0 = f_arrdiv32_fs186_not0 & b[26];
  assign f_arrdiv32_fs186_xor1 = f_arrdiv32_fs185_or0 ^ f_arrdiv32_fs186_xor0;
  assign f_arrdiv32_fs186_not1 = ~f_arrdiv32_fs186_xor0;
  assign f_arrdiv32_fs186_and1 = f_arrdiv32_fs186_not1 & f_arrdiv32_fs185_or0;
  assign f_arrdiv32_fs186_or0 = f_arrdiv32_fs186_and1 | f_arrdiv32_fs186_and0;
  assign f_arrdiv32_fs187_xor0 = f_arrdiv32_mux2to1150_xor0 ^ b[27];
  assign f_arrdiv32_fs187_not0 = ~f_arrdiv32_mux2to1150_xor0;
  assign f_arrdiv32_fs187_and0 = f_arrdiv32_fs187_not0 & b[27];
  assign f_arrdiv32_fs187_xor1 = f_arrdiv32_fs186_or0 ^ f_arrdiv32_fs187_xor0;
  assign f_arrdiv32_fs187_not1 = ~f_arrdiv32_fs187_xor0;
  assign f_arrdiv32_fs187_and1 = f_arrdiv32_fs187_not1 & f_arrdiv32_fs186_or0;
  assign f_arrdiv32_fs187_or0 = f_arrdiv32_fs187_and1 | f_arrdiv32_fs187_and0;
  assign f_arrdiv32_fs188_xor0 = f_arrdiv32_mux2to1151_xor0 ^ b[28];
  assign f_arrdiv32_fs188_not0 = ~f_arrdiv32_mux2to1151_xor0;
  assign f_arrdiv32_fs188_and0 = f_arrdiv32_fs188_not0 & b[28];
  assign f_arrdiv32_fs188_xor1 = f_arrdiv32_fs187_or0 ^ f_arrdiv32_fs188_xor0;
  assign f_arrdiv32_fs188_not1 = ~f_arrdiv32_fs188_xor0;
  assign f_arrdiv32_fs188_and1 = f_arrdiv32_fs188_not1 & f_arrdiv32_fs187_or0;
  assign f_arrdiv32_fs188_or0 = f_arrdiv32_fs188_and1 | f_arrdiv32_fs188_and0;
  assign f_arrdiv32_fs189_xor0 = f_arrdiv32_mux2to1152_xor0 ^ b[29];
  assign f_arrdiv32_fs189_not0 = ~f_arrdiv32_mux2to1152_xor0;
  assign f_arrdiv32_fs189_and0 = f_arrdiv32_fs189_not0 & b[29];
  assign f_arrdiv32_fs189_xor1 = f_arrdiv32_fs188_or0 ^ f_arrdiv32_fs189_xor0;
  assign f_arrdiv32_fs189_not1 = ~f_arrdiv32_fs189_xor0;
  assign f_arrdiv32_fs189_and1 = f_arrdiv32_fs189_not1 & f_arrdiv32_fs188_or0;
  assign f_arrdiv32_fs189_or0 = f_arrdiv32_fs189_and1 | f_arrdiv32_fs189_and0;
  assign f_arrdiv32_fs190_xor0 = f_arrdiv32_mux2to1153_xor0 ^ b[30];
  assign f_arrdiv32_fs190_not0 = ~f_arrdiv32_mux2to1153_xor0;
  assign f_arrdiv32_fs190_and0 = f_arrdiv32_fs190_not0 & b[30];
  assign f_arrdiv32_fs190_xor1 = f_arrdiv32_fs189_or0 ^ f_arrdiv32_fs190_xor0;
  assign f_arrdiv32_fs190_not1 = ~f_arrdiv32_fs190_xor0;
  assign f_arrdiv32_fs190_and1 = f_arrdiv32_fs190_not1 & f_arrdiv32_fs189_or0;
  assign f_arrdiv32_fs190_or0 = f_arrdiv32_fs190_and1 | f_arrdiv32_fs190_and0;
  assign f_arrdiv32_fs191_xor0 = f_arrdiv32_mux2to1154_xor0 ^ b[31];
  assign f_arrdiv32_fs191_not0 = ~f_arrdiv32_mux2to1154_xor0;
  assign f_arrdiv32_fs191_and0 = f_arrdiv32_fs191_not0 & b[31];
  assign f_arrdiv32_fs191_xor1 = f_arrdiv32_fs190_or0 ^ f_arrdiv32_fs191_xor0;
  assign f_arrdiv32_fs191_not1 = ~f_arrdiv32_fs191_xor0;
  assign f_arrdiv32_fs191_and1 = f_arrdiv32_fs191_not1 & f_arrdiv32_fs190_or0;
  assign f_arrdiv32_fs191_or0 = f_arrdiv32_fs191_and1 | f_arrdiv32_fs191_and0;
  assign f_arrdiv32_mux2to1155_and0 = a[26] & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1155_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1155_and1 = f_arrdiv32_fs160_xor0 & f_arrdiv32_mux2to1155_not0;
  assign f_arrdiv32_mux2to1155_xor0 = f_arrdiv32_mux2to1155_and0 ^ f_arrdiv32_mux2to1155_and1;
  assign f_arrdiv32_mux2to1156_and0 = f_arrdiv32_mux2to1124_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1156_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1156_and1 = f_arrdiv32_fs161_xor1 & f_arrdiv32_mux2to1156_not0;
  assign f_arrdiv32_mux2to1156_xor0 = f_arrdiv32_mux2to1156_and0 ^ f_arrdiv32_mux2to1156_and1;
  assign f_arrdiv32_mux2to1157_and0 = f_arrdiv32_mux2to1125_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1157_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1157_and1 = f_arrdiv32_fs162_xor1 & f_arrdiv32_mux2to1157_not0;
  assign f_arrdiv32_mux2to1157_xor0 = f_arrdiv32_mux2to1157_and0 ^ f_arrdiv32_mux2to1157_and1;
  assign f_arrdiv32_mux2to1158_and0 = f_arrdiv32_mux2to1126_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1158_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1158_and1 = f_arrdiv32_fs163_xor1 & f_arrdiv32_mux2to1158_not0;
  assign f_arrdiv32_mux2to1158_xor0 = f_arrdiv32_mux2to1158_and0 ^ f_arrdiv32_mux2to1158_and1;
  assign f_arrdiv32_mux2to1159_and0 = f_arrdiv32_mux2to1127_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1159_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1159_and1 = f_arrdiv32_fs164_xor1 & f_arrdiv32_mux2to1159_not0;
  assign f_arrdiv32_mux2to1159_xor0 = f_arrdiv32_mux2to1159_and0 ^ f_arrdiv32_mux2to1159_and1;
  assign f_arrdiv32_mux2to1160_and0 = f_arrdiv32_mux2to1128_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1160_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1160_and1 = f_arrdiv32_fs165_xor1 & f_arrdiv32_mux2to1160_not0;
  assign f_arrdiv32_mux2to1160_xor0 = f_arrdiv32_mux2to1160_and0 ^ f_arrdiv32_mux2to1160_and1;
  assign f_arrdiv32_mux2to1161_and0 = f_arrdiv32_mux2to1129_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1161_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1161_and1 = f_arrdiv32_fs166_xor1 & f_arrdiv32_mux2to1161_not0;
  assign f_arrdiv32_mux2to1161_xor0 = f_arrdiv32_mux2to1161_and0 ^ f_arrdiv32_mux2to1161_and1;
  assign f_arrdiv32_mux2to1162_and0 = f_arrdiv32_mux2to1130_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1162_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1162_and1 = f_arrdiv32_fs167_xor1 & f_arrdiv32_mux2to1162_not0;
  assign f_arrdiv32_mux2to1162_xor0 = f_arrdiv32_mux2to1162_and0 ^ f_arrdiv32_mux2to1162_and1;
  assign f_arrdiv32_mux2to1163_and0 = f_arrdiv32_mux2to1131_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1163_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1163_and1 = f_arrdiv32_fs168_xor1 & f_arrdiv32_mux2to1163_not0;
  assign f_arrdiv32_mux2to1163_xor0 = f_arrdiv32_mux2to1163_and0 ^ f_arrdiv32_mux2to1163_and1;
  assign f_arrdiv32_mux2to1164_and0 = f_arrdiv32_mux2to1132_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1164_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1164_and1 = f_arrdiv32_fs169_xor1 & f_arrdiv32_mux2to1164_not0;
  assign f_arrdiv32_mux2to1164_xor0 = f_arrdiv32_mux2to1164_and0 ^ f_arrdiv32_mux2to1164_and1;
  assign f_arrdiv32_mux2to1165_and0 = f_arrdiv32_mux2to1133_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1165_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1165_and1 = f_arrdiv32_fs170_xor1 & f_arrdiv32_mux2to1165_not0;
  assign f_arrdiv32_mux2to1165_xor0 = f_arrdiv32_mux2to1165_and0 ^ f_arrdiv32_mux2to1165_and1;
  assign f_arrdiv32_mux2to1166_and0 = f_arrdiv32_mux2to1134_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1166_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1166_and1 = f_arrdiv32_fs171_xor1 & f_arrdiv32_mux2to1166_not0;
  assign f_arrdiv32_mux2to1166_xor0 = f_arrdiv32_mux2to1166_and0 ^ f_arrdiv32_mux2to1166_and1;
  assign f_arrdiv32_mux2to1167_and0 = f_arrdiv32_mux2to1135_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1167_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1167_and1 = f_arrdiv32_fs172_xor1 & f_arrdiv32_mux2to1167_not0;
  assign f_arrdiv32_mux2to1167_xor0 = f_arrdiv32_mux2to1167_and0 ^ f_arrdiv32_mux2to1167_and1;
  assign f_arrdiv32_mux2to1168_and0 = f_arrdiv32_mux2to1136_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1168_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1168_and1 = f_arrdiv32_fs173_xor1 & f_arrdiv32_mux2to1168_not0;
  assign f_arrdiv32_mux2to1168_xor0 = f_arrdiv32_mux2to1168_and0 ^ f_arrdiv32_mux2to1168_and1;
  assign f_arrdiv32_mux2to1169_and0 = f_arrdiv32_mux2to1137_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1169_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1169_and1 = f_arrdiv32_fs174_xor1 & f_arrdiv32_mux2to1169_not0;
  assign f_arrdiv32_mux2to1169_xor0 = f_arrdiv32_mux2to1169_and0 ^ f_arrdiv32_mux2to1169_and1;
  assign f_arrdiv32_mux2to1170_and0 = f_arrdiv32_mux2to1138_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1170_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1170_and1 = f_arrdiv32_fs175_xor1 & f_arrdiv32_mux2to1170_not0;
  assign f_arrdiv32_mux2to1170_xor0 = f_arrdiv32_mux2to1170_and0 ^ f_arrdiv32_mux2to1170_and1;
  assign f_arrdiv32_mux2to1171_and0 = f_arrdiv32_mux2to1139_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1171_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1171_and1 = f_arrdiv32_fs176_xor1 & f_arrdiv32_mux2to1171_not0;
  assign f_arrdiv32_mux2to1171_xor0 = f_arrdiv32_mux2to1171_and0 ^ f_arrdiv32_mux2to1171_and1;
  assign f_arrdiv32_mux2to1172_and0 = f_arrdiv32_mux2to1140_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1172_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1172_and1 = f_arrdiv32_fs177_xor1 & f_arrdiv32_mux2to1172_not0;
  assign f_arrdiv32_mux2to1172_xor0 = f_arrdiv32_mux2to1172_and0 ^ f_arrdiv32_mux2to1172_and1;
  assign f_arrdiv32_mux2to1173_and0 = f_arrdiv32_mux2to1141_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1173_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1173_and1 = f_arrdiv32_fs178_xor1 & f_arrdiv32_mux2to1173_not0;
  assign f_arrdiv32_mux2to1173_xor0 = f_arrdiv32_mux2to1173_and0 ^ f_arrdiv32_mux2to1173_and1;
  assign f_arrdiv32_mux2to1174_and0 = f_arrdiv32_mux2to1142_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1174_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1174_and1 = f_arrdiv32_fs179_xor1 & f_arrdiv32_mux2to1174_not0;
  assign f_arrdiv32_mux2to1174_xor0 = f_arrdiv32_mux2to1174_and0 ^ f_arrdiv32_mux2to1174_and1;
  assign f_arrdiv32_mux2to1175_and0 = f_arrdiv32_mux2to1143_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1175_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1175_and1 = f_arrdiv32_fs180_xor1 & f_arrdiv32_mux2to1175_not0;
  assign f_arrdiv32_mux2to1175_xor0 = f_arrdiv32_mux2to1175_and0 ^ f_arrdiv32_mux2to1175_and1;
  assign f_arrdiv32_mux2to1176_and0 = f_arrdiv32_mux2to1144_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1176_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1176_and1 = f_arrdiv32_fs181_xor1 & f_arrdiv32_mux2to1176_not0;
  assign f_arrdiv32_mux2to1176_xor0 = f_arrdiv32_mux2to1176_and0 ^ f_arrdiv32_mux2to1176_and1;
  assign f_arrdiv32_mux2to1177_and0 = f_arrdiv32_mux2to1145_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1177_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1177_and1 = f_arrdiv32_fs182_xor1 & f_arrdiv32_mux2to1177_not0;
  assign f_arrdiv32_mux2to1177_xor0 = f_arrdiv32_mux2to1177_and0 ^ f_arrdiv32_mux2to1177_and1;
  assign f_arrdiv32_mux2to1178_and0 = f_arrdiv32_mux2to1146_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1178_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1178_and1 = f_arrdiv32_fs183_xor1 & f_arrdiv32_mux2to1178_not0;
  assign f_arrdiv32_mux2to1178_xor0 = f_arrdiv32_mux2to1178_and0 ^ f_arrdiv32_mux2to1178_and1;
  assign f_arrdiv32_mux2to1179_and0 = f_arrdiv32_mux2to1147_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1179_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1179_and1 = f_arrdiv32_fs184_xor1 & f_arrdiv32_mux2to1179_not0;
  assign f_arrdiv32_mux2to1179_xor0 = f_arrdiv32_mux2to1179_and0 ^ f_arrdiv32_mux2to1179_and1;
  assign f_arrdiv32_mux2to1180_and0 = f_arrdiv32_mux2to1148_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1180_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1180_and1 = f_arrdiv32_fs185_xor1 & f_arrdiv32_mux2to1180_not0;
  assign f_arrdiv32_mux2to1180_xor0 = f_arrdiv32_mux2to1180_and0 ^ f_arrdiv32_mux2to1180_and1;
  assign f_arrdiv32_mux2to1181_and0 = f_arrdiv32_mux2to1149_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1181_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1181_and1 = f_arrdiv32_fs186_xor1 & f_arrdiv32_mux2to1181_not0;
  assign f_arrdiv32_mux2to1181_xor0 = f_arrdiv32_mux2to1181_and0 ^ f_arrdiv32_mux2to1181_and1;
  assign f_arrdiv32_mux2to1182_and0 = f_arrdiv32_mux2to1150_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1182_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1182_and1 = f_arrdiv32_fs187_xor1 & f_arrdiv32_mux2to1182_not0;
  assign f_arrdiv32_mux2to1182_xor0 = f_arrdiv32_mux2to1182_and0 ^ f_arrdiv32_mux2to1182_and1;
  assign f_arrdiv32_mux2to1183_and0 = f_arrdiv32_mux2to1151_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1183_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1183_and1 = f_arrdiv32_fs188_xor1 & f_arrdiv32_mux2to1183_not0;
  assign f_arrdiv32_mux2to1183_xor0 = f_arrdiv32_mux2to1183_and0 ^ f_arrdiv32_mux2to1183_and1;
  assign f_arrdiv32_mux2to1184_and0 = f_arrdiv32_mux2to1152_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1184_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1184_and1 = f_arrdiv32_fs189_xor1 & f_arrdiv32_mux2to1184_not0;
  assign f_arrdiv32_mux2to1184_xor0 = f_arrdiv32_mux2to1184_and0 ^ f_arrdiv32_mux2to1184_and1;
  assign f_arrdiv32_mux2to1185_and0 = f_arrdiv32_mux2to1153_xor0 & f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1185_not0 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_mux2to1185_and1 = f_arrdiv32_fs190_xor1 & f_arrdiv32_mux2to1185_not0;
  assign f_arrdiv32_mux2to1185_xor0 = f_arrdiv32_mux2to1185_and0 ^ f_arrdiv32_mux2to1185_and1;
  assign f_arrdiv32_not5 = ~f_arrdiv32_fs191_or0;
  assign f_arrdiv32_fs192_xor0 = a[25] ^ b[0];
  assign f_arrdiv32_fs192_not0 = ~a[25];
  assign f_arrdiv32_fs192_and0 = f_arrdiv32_fs192_not0 & b[0];
  assign f_arrdiv32_fs192_not1 = ~f_arrdiv32_fs192_xor0;
  assign f_arrdiv32_fs193_xor0 = f_arrdiv32_mux2to1155_xor0 ^ b[1];
  assign f_arrdiv32_fs193_not0 = ~f_arrdiv32_mux2to1155_xor0;
  assign f_arrdiv32_fs193_and0 = f_arrdiv32_fs193_not0 & b[1];
  assign f_arrdiv32_fs193_xor1 = f_arrdiv32_fs192_and0 ^ f_arrdiv32_fs193_xor0;
  assign f_arrdiv32_fs193_not1 = ~f_arrdiv32_fs193_xor0;
  assign f_arrdiv32_fs193_and1 = f_arrdiv32_fs193_not1 & f_arrdiv32_fs192_and0;
  assign f_arrdiv32_fs193_or0 = f_arrdiv32_fs193_and1 | f_arrdiv32_fs193_and0;
  assign f_arrdiv32_fs194_xor0 = f_arrdiv32_mux2to1156_xor0 ^ b[2];
  assign f_arrdiv32_fs194_not0 = ~f_arrdiv32_mux2to1156_xor0;
  assign f_arrdiv32_fs194_and0 = f_arrdiv32_fs194_not0 & b[2];
  assign f_arrdiv32_fs194_xor1 = f_arrdiv32_fs193_or0 ^ f_arrdiv32_fs194_xor0;
  assign f_arrdiv32_fs194_not1 = ~f_arrdiv32_fs194_xor0;
  assign f_arrdiv32_fs194_and1 = f_arrdiv32_fs194_not1 & f_arrdiv32_fs193_or0;
  assign f_arrdiv32_fs194_or0 = f_arrdiv32_fs194_and1 | f_arrdiv32_fs194_and0;
  assign f_arrdiv32_fs195_xor0 = f_arrdiv32_mux2to1157_xor0 ^ b[3];
  assign f_arrdiv32_fs195_not0 = ~f_arrdiv32_mux2to1157_xor0;
  assign f_arrdiv32_fs195_and0 = f_arrdiv32_fs195_not0 & b[3];
  assign f_arrdiv32_fs195_xor1 = f_arrdiv32_fs194_or0 ^ f_arrdiv32_fs195_xor0;
  assign f_arrdiv32_fs195_not1 = ~f_arrdiv32_fs195_xor0;
  assign f_arrdiv32_fs195_and1 = f_arrdiv32_fs195_not1 & f_arrdiv32_fs194_or0;
  assign f_arrdiv32_fs195_or0 = f_arrdiv32_fs195_and1 | f_arrdiv32_fs195_and0;
  assign f_arrdiv32_fs196_xor0 = f_arrdiv32_mux2to1158_xor0 ^ b[4];
  assign f_arrdiv32_fs196_not0 = ~f_arrdiv32_mux2to1158_xor0;
  assign f_arrdiv32_fs196_and0 = f_arrdiv32_fs196_not0 & b[4];
  assign f_arrdiv32_fs196_xor1 = f_arrdiv32_fs195_or0 ^ f_arrdiv32_fs196_xor0;
  assign f_arrdiv32_fs196_not1 = ~f_arrdiv32_fs196_xor0;
  assign f_arrdiv32_fs196_and1 = f_arrdiv32_fs196_not1 & f_arrdiv32_fs195_or0;
  assign f_arrdiv32_fs196_or0 = f_arrdiv32_fs196_and1 | f_arrdiv32_fs196_and0;
  assign f_arrdiv32_fs197_xor0 = f_arrdiv32_mux2to1159_xor0 ^ b[5];
  assign f_arrdiv32_fs197_not0 = ~f_arrdiv32_mux2to1159_xor0;
  assign f_arrdiv32_fs197_and0 = f_arrdiv32_fs197_not0 & b[5];
  assign f_arrdiv32_fs197_xor1 = f_arrdiv32_fs196_or0 ^ f_arrdiv32_fs197_xor0;
  assign f_arrdiv32_fs197_not1 = ~f_arrdiv32_fs197_xor0;
  assign f_arrdiv32_fs197_and1 = f_arrdiv32_fs197_not1 & f_arrdiv32_fs196_or0;
  assign f_arrdiv32_fs197_or0 = f_arrdiv32_fs197_and1 | f_arrdiv32_fs197_and0;
  assign f_arrdiv32_fs198_xor0 = f_arrdiv32_mux2to1160_xor0 ^ b[6];
  assign f_arrdiv32_fs198_not0 = ~f_arrdiv32_mux2to1160_xor0;
  assign f_arrdiv32_fs198_and0 = f_arrdiv32_fs198_not0 & b[6];
  assign f_arrdiv32_fs198_xor1 = f_arrdiv32_fs197_or0 ^ f_arrdiv32_fs198_xor0;
  assign f_arrdiv32_fs198_not1 = ~f_arrdiv32_fs198_xor0;
  assign f_arrdiv32_fs198_and1 = f_arrdiv32_fs198_not1 & f_arrdiv32_fs197_or0;
  assign f_arrdiv32_fs198_or0 = f_arrdiv32_fs198_and1 | f_arrdiv32_fs198_and0;
  assign f_arrdiv32_fs199_xor0 = f_arrdiv32_mux2to1161_xor0 ^ b[7];
  assign f_arrdiv32_fs199_not0 = ~f_arrdiv32_mux2to1161_xor0;
  assign f_arrdiv32_fs199_and0 = f_arrdiv32_fs199_not0 & b[7];
  assign f_arrdiv32_fs199_xor1 = f_arrdiv32_fs198_or0 ^ f_arrdiv32_fs199_xor0;
  assign f_arrdiv32_fs199_not1 = ~f_arrdiv32_fs199_xor0;
  assign f_arrdiv32_fs199_and1 = f_arrdiv32_fs199_not1 & f_arrdiv32_fs198_or0;
  assign f_arrdiv32_fs199_or0 = f_arrdiv32_fs199_and1 | f_arrdiv32_fs199_and0;
  assign f_arrdiv32_fs200_xor0 = f_arrdiv32_mux2to1162_xor0 ^ b[8];
  assign f_arrdiv32_fs200_not0 = ~f_arrdiv32_mux2to1162_xor0;
  assign f_arrdiv32_fs200_and0 = f_arrdiv32_fs200_not0 & b[8];
  assign f_arrdiv32_fs200_xor1 = f_arrdiv32_fs199_or0 ^ f_arrdiv32_fs200_xor0;
  assign f_arrdiv32_fs200_not1 = ~f_arrdiv32_fs200_xor0;
  assign f_arrdiv32_fs200_and1 = f_arrdiv32_fs200_not1 & f_arrdiv32_fs199_or0;
  assign f_arrdiv32_fs200_or0 = f_arrdiv32_fs200_and1 | f_arrdiv32_fs200_and0;
  assign f_arrdiv32_fs201_xor0 = f_arrdiv32_mux2to1163_xor0 ^ b[9];
  assign f_arrdiv32_fs201_not0 = ~f_arrdiv32_mux2to1163_xor0;
  assign f_arrdiv32_fs201_and0 = f_arrdiv32_fs201_not0 & b[9];
  assign f_arrdiv32_fs201_xor1 = f_arrdiv32_fs200_or0 ^ f_arrdiv32_fs201_xor0;
  assign f_arrdiv32_fs201_not1 = ~f_arrdiv32_fs201_xor0;
  assign f_arrdiv32_fs201_and1 = f_arrdiv32_fs201_not1 & f_arrdiv32_fs200_or0;
  assign f_arrdiv32_fs201_or0 = f_arrdiv32_fs201_and1 | f_arrdiv32_fs201_and0;
  assign f_arrdiv32_fs202_xor0 = f_arrdiv32_mux2to1164_xor0 ^ b[10];
  assign f_arrdiv32_fs202_not0 = ~f_arrdiv32_mux2to1164_xor0;
  assign f_arrdiv32_fs202_and0 = f_arrdiv32_fs202_not0 & b[10];
  assign f_arrdiv32_fs202_xor1 = f_arrdiv32_fs201_or0 ^ f_arrdiv32_fs202_xor0;
  assign f_arrdiv32_fs202_not1 = ~f_arrdiv32_fs202_xor0;
  assign f_arrdiv32_fs202_and1 = f_arrdiv32_fs202_not1 & f_arrdiv32_fs201_or0;
  assign f_arrdiv32_fs202_or0 = f_arrdiv32_fs202_and1 | f_arrdiv32_fs202_and0;
  assign f_arrdiv32_fs203_xor0 = f_arrdiv32_mux2to1165_xor0 ^ b[11];
  assign f_arrdiv32_fs203_not0 = ~f_arrdiv32_mux2to1165_xor0;
  assign f_arrdiv32_fs203_and0 = f_arrdiv32_fs203_not0 & b[11];
  assign f_arrdiv32_fs203_xor1 = f_arrdiv32_fs202_or0 ^ f_arrdiv32_fs203_xor0;
  assign f_arrdiv32_fs203_not1 = ~f_arrdiv32_fs203_xor0;
  assign f_arrdiv32_fs203_and1 = f_arrdiv32_fs203_not1 & f_arrdiv32_fs202_or0;
  assign f_arrdiv32_fs203_or0 = f_arrdiv32_fs203_and1 | f_arrdiv32_fs203_and0;
  assign f_arrdiv32_fs204_xor0 = f_arrdiv32_mux2to1166_xor0 ^ b[12];
  assign f_arrdiv32_fs204_not0 = ~f_arrdiv32_mux2to1166_xor0;
  assign f_arrdiv32_fs204_and0 = f_arrdiv32_fs204_not0 & b[12];
  assign f_arrdiv32_fs204_xor1 = f_arrdiv32_fs203_or0 ^ f_arrdiv32_fs204_xor0;
  assign f_arrdiv32_fs204_not1 = ~f_arrdiv32_fs204_xor0;
  assign f_arrdiv32_fs204_and1 = f_arrdiv32_fs204_not1 & f_arrdiv32_fs203_or0;
  assign f_arrdiv32_fs204_or0 = f_arrdiv32_fs204_and1 | f_arrdiv32_fs204_and0;
  assign f_arrdiv32_fs205_xor0 = f_arrdiv32_mux2to1167_xor0 ^ b[13];
  assign f_arrdiv32_fs205_not0 = ~f_arrdiv32_mux2to1167_xor0;
  assign f_arrdiv32_fs205_and0 = f_arrdiv32_fs205_not0 & b[13];
  assign f_arrdiv32_fs205_xor1 = f_arrdiv32_fs204_or0 ^ f_arrdiv32_fs205_xor0;
  assign f_arrdiv32_fs205_not1 = ~f_arrdiv32_fs205_xor0;
  assign f_arrdiv32_fs205_and1 = f_arrdiv32_fs205_not1 & f_arrdiv32_fs204_or0;
  assign f_arrdiv32_fs205_or0 = f_arrdiv32_fs205_and1 | f_arrdiv32_fs205_and0;
  assign f_arrdiv32_fs206_xor0 = f_arrdiv32_mux2to1168_xor0 ^ b[14];
  assign f_arrdiv32_fs206_not0 = ~f_arrdiv32_mux2to1168_xor0;
  assign f_arrdiv32_fs206_and0 = f_arrdiv32_fs206_not0 & b[14];
  assign f_arrdiv32_fs206_xor1 = f_arrdiv32_fs205_or0 ^ f_arrdiv32_fs206_xor0;
  assign f_arrdiv32_fs206_not1 = ~f_arrdiv32_fs206_xor0;
  assign f_arrdiv32_fs206_and1 = f_arrdiv32_fs206_not1 & f_arrdiv32_fs205_or0;
  assign f_arrdiv32_fs206_or0 = f_arrdiv32_fs206_and1 | f_arrdiv32_fs206_and0;
  assign f_arrdiv32_fs207_xor0 = f_arrdiv32_mux2to1169_xor0 ^ b[15];
  assign f_arrdiv32_fs207_not0 = ~f_arrdiv32_mux2to1169_xor0;
  assign f_arrdiv32_fs207_and0 = f_arrdiv32_fs207_not0 & b[15];
  assign f_arrdiv32_fs207_xor1 = f_arrdiv32_fs206_or0 ^ f_arrdiv32_fs207_xor0;
  assign f_arrdiv32_fs207_not1 = ~f_arrdiv32_fs207_xor0;
  assign f_arrdiv32_fs207_and1 = f_arrdiv32_fs207_not1 & f_arrdiv32_fs206_or0;
  assign f_arrdiv32_fs207_or0 = f_arrdiv32_fs207_and1 | f_arrdiv32_fs207_and0;
  assign f_arrdiv32_fs208_xor0 = f_arrdiv32_mux2to1170_xor0 ^ b[16];
  assign f_arrdiv32_fs208_not0 = ~f_arrdiv32_mux2to1170_xor0;
  assign f_arrdiv32_fs208_and0 = f_arrdiv32_fs208_not0 & b[16];
  assign f_arrdiv32_fs208_xor1 = f_arrdiv32_fs207_or0 ^ f_arrdiv32_fs208_xor0;
  assign f_arrdiv32_fs208_not1 = ~f_arrdiv32_fs208_xor0;
  assign f_arrdiv32_fs208_and1 = f_arrdiv32_fs208_not1 & f_arrdiv32_fs207_or0;
  assign f_arrdiv32_fs208_or0 = f_arrdiv32_fs208_and1 | f_arrdiv32_fs208_and0;
  assign f_arrdiv32_fs209_xor0 = f_arrdiv32_mux2to1171_xor0 ^ b[17];
  assign f_arrdiv32_fs209_not0 = ~f_arrdiv32_mux2to1171_xor0;
  assign f_arrdiv32_fs209_and0 = f_arrdiv32_fs209_not0 & b[17];
  assign f_arrdiv32_fs209_xor1 = f_arrdiv32_fs208_or0 ^ f_arrdiv32_fs209_xor0;
  assign f_arrdiv32_fs209_not1 = ~f_arrdiv32_fs209_xor0;
  assign f_arrdiv32_fs209_and1 = f_arrdiv32_fs209_not1 & f_arrdiv32_fs208_or0;
  assign f_arrdiv32_fs209_or0 = f_arrdiv32_fs209_and1 | f_arrdiv32_fs209_and0;
  assign f_arrdiv32_fs210_xor0 = f_arrdiv32_mux2to1172_xor0 ^ b[18];
  assign f_arrdiv32_fs210_not0 = ~f_arrdiv32_mux2to1172_xor0;
  assign f_arrdiv32_fs210_and0 = f_arrdiv32_fs210_not0 & b[18];
  assign f_arrdiv32_fs210_xor1 = f_arrdiv32_fs209_or0 ^ f_arrdiv32_fs210_xor0;
  assign f_arrdiv32_fs210_not1 = ~f_arrdiv32_fs210_xor0;
  assign f_arrdiv32_fs210_and1 = f_arrdiv32_fs210_not1 & f_arrdiv32_fs209_or0;
  assign f_arrdiv32_fs210_or0 = f_arrdiv32_fs210_and1 | f_arrdiv32_fs210_and0;
  assign f_arrdiv32_fs211_xor0 = f_arrdiv32_mux2to1173_xor0 ^ b[19];
  assign f_arrdiv32_fs211_not0 = ~f_arrdiv32_mux2to1173_xor0;
  assign f_arrdiv32_fs211_and0 = f_arrdiv32_fs211_not0 & b[19];
  assign f_arrdiv32_fs211_xor1 = f_arrdiv32_fs210_or0 ^ f_arrdiv32_fs211_xor0;
  assign f_arrdiv32_fs211_not1 = ~f_arrdiv32_fs211_xor0;
  assign f_arrdiv32_fs211_and1 = f_arrdiv32_fs211_not1 & f_arrdiv32_fs210_or0;
  assign f_arrdiv32_fs211_or0 = f_arrdiv32_fs211_and1 | f_arrdiv32_fs211_and0;
  assign f_arrdiv32_fs212_xor0 = f_arrdiv32_mux2to1174_xor0 ^ b[20];
  assign f_arrdiv32_fs212_not0 = ~f_arrdiv32_mux2to1174_xor0;
  assign f_arrdiv32_fs212_and0 = f_arrdiv32_fs212_not0 & b[20];
  assign f_arrdiv32_fs212_xor1 = f_arrdiv32_fs211_or0 ^ f_arrdiv32_fs212_xor0;
  assign f_arrdiv32_fs212_not1 = ~f_arrdiv32_fs212_xor0;
  assign f_arrdiv32_fs212_and1 = f_arrdiv32_fs212_not1 & f_arrdiv32_fs211_or0;
  assign f_arrdiv32_fs212_or0 = f_arrdiv32_fs212_and1 | f_arrdiv32_fs212_and0;
  assign f_arrdiv32_fs213_xor0 = f_arrdiv32_mux2to1175_xor0 ^ b[21];
  assign f_arrdiv32_fs213_not0 = ~f_arrdiv32_mux2to1175_xor0;
  assign f_arrdiv32_fs213_and0 = f_arrdiv32_fs213_not0 & b[21];
  assign f_arrdiv32_fs213_xor1 = f_arrdiv32_fs212_or0 ^ f_arrdiv32_fs213_xor0;
  assign f_arrdiv32_fs213_not1 = ~f_arrdiv32_fs213_xor0;
  assign f_arrdiv32_fs213_and1 = f_arrdiv32_fs213_not1 & f_arrdiv32_fs212_or0;
  assign f_arrdiv32_fs213_or0 = f_arrdiv32_fs213_and1 | f_arrdiv32_fs213_and0;
  assign f_arrdiv32_fs214_xor0 = f_arrdiv32_mux2to1176_xor0 ^ b[22];
  assign f_arrdiv32_fs214_not0 = ~f_arrdiv32_mux2to1176_xor0;
  assign f_arrdiv32_fs214_and0 = f_arrdiv32_fs214_not0 & b[22];
  assign f_arrdiv32_fs214_xor1 = f_arrdiv32_fs213_or0 ^ f_arrdiv32_fs214_xor0;
  assign f_arrdiv32_fs214_not1 = ~f_arrdiv32_fs214_xor0;
  assign f_arrdiv32_fs214_and1 = f_arrdiv32_fs214_not1 & f_arrdiv32_fs213_or0;
  assign f_arrdiv32_fs214_or0 = f_arrdiv32_fs214_and1 | f_arrdiv32_fs214_and0;
  assign f_arrdiv32_fs215_xor0 = f_arrdiv32_mux2to1177_xor0 ^ b[23];
  assign f_arrdiv32_fs215_not0 = ~f_arrdiv32_mux2to1177_xor0;
  assign f_arrdiv32_fs215_and0 = f_arrdiv32_fs215_not0 & b[23];
  assign f_arrdiv32_fs215_xor1 = f_arrdiv32_fs214_or0 ^ f_arrdiv32_fs215_xor0;
  assign f_arrdiv32_fs215_not1 = ~f_arrdiv32_fs215_xor0;
  assign f_arrdiv32_fs215_and1 = f_arrdiv32_fs215_not1 & f_arrdiv32_fs214_or0;
  assign f_arrdiv32_fs215_or0 = f_arrdiv32_fs215_and1 | f_arrdiv32_fs215_and0;
  assign f_arrdiv32_fs216_xor0 = f_arrdiv32_mux2to1178_xor0 ^ b[24];
  assign f_arrdiv32_fs216_not0 = ~f_arrdiv32_mux2to1178_xor0;
  assign f_arrdiv32_fs216_and0 = f_arrdiv32_fs216_not0 & b[24];
  assign f_arrdiv32_fs216_xor1 = f_arrdiv32_fs215_or0 ^ f_arrdiv32_fs216_xor0;
  assign f_arrdiv32_fs216_not1 = ~f_arrdiv32_fs216_xor0;
  assign f_arrdiv32_fs216_and1 = f_arrdiv32_fs216_not1 & f_arrdiv32_fs215_or0;
  assign f_arrdiv32_fs216_or0 = f_arrdiv32_fs216_and1 | f_arrdiv32_fs216_and0;
  assign f_arrdiv32_fs217_xor0 = f_arrdiv32_mux2to1179_xor0 ^ b[25];
  assign f_arrdiv32_fs217_not0 = ~f_arrdiv32_mux2to1179_xor0;
  assign f_arrdiv32_fs217_and0 = f_arrdiv32_fs217_not0 & b[25];
  assign f_arrdiv32_fs217_xor1 = f_arrdiv32_fs216_or0 ^ f_arrdiv32_fs217_xor0;
  assign f_arrdiv32_fs217_not1 = ~f_arrdiv32_fs217_xor0;
  assign f_arrdiv32_fs217_and1 = f_arrdiv32_fs217_not1 & f_arrdiv32_fs216_or0;
  assign f_arrdiv32_fs217_or0 = f_arrdiv32_fs217_and1 | f_arrdiv32_fs217_and0;
  assign f_arrdiv32_fs218_xor0 = f_arrdiv32_mux2to1180_xor0 ^ b[26];
  assign f_arrdiv32_fs218_not0 = ~f_arrdiv32_mux2to1180_xor0;
  assign f_arrdiv32_fs218_and0 = f_arrdiv32_fs218_not0 & b[26];
  assign f_arrdiv32_fs218_xor1 = f_arrdiv32_fs217_or0 ^ f_arrdiv32_fs218_xor0;
  assign f_arrdiv32_fs218_not1 = ~f_arrdiv32_fs218_xor0;
  assign f_arrdiv32_fs218_and1 = f_arrdiv32_fs218_not1 & f_arrdiv32_fs217_or0;
  assign f_arrdiv32_fs218_or0 = f_arrdiv32_fs218_and1 | f_arrdiv32_fs218_and0;
  assign f_arrdiv32_fs219_xor0 = f_arrdiv32_mux2to1181_xor0 ^ b[27];
  assign f_arrdiv32_fs219_not0 = ~f_arrdiv32_mux2to1181_xor0;
  assign f_arrdiv32_fs219_and0 = f_arrdiv32_fs219_not0 & b[27];
  assign f_arrdiv32_fs219_xor1 = f_arrdiv32_fs218_or0 ^ f_arrdiv32_fs219_xor0;
  assign f_arrdiv32_fs219_not1 = ~f_arrdiv32_fs219_xor0;
  assign f_arrdiv32_fs219_and1 = f_arrdiv32_fs219_not1 & f_arrdiv32_fs218_or0;
  assign f_arrdiv32_fs219_or0 = f_arrdiv32_fs219_and1 | f_arrdiv32_fs219_and0;
  assign f_arrdiv32_fs220_xor0 = f_arrdiv32_mux2to1182_xor0 ^ b[28];
  assign f_arrdiv32_fs220_not0 = ~f_arrdiv32_mux2to1182_xor0;
  assign f_arrdiv32_fs220_and0 = f_arrdiv32_fs220_not0 & b[28];
  assign f_arrdiv32_fs220_xor1 = f_arrdiv32_fs219_or0 ^ f_arrdiv32_fs220_xor0;
  assign f_arrdiv32_fs220_not1 = ~f_arrdiv32_fs220_xor0;
  assign f_arrdiv32_fs220_and1 = f_arrdiv32_fs220_not1 & f_arrdiv32_fs219_or0;
  assign f_arrdiv32_fs220_or0 = f_arrdiv32_fs220_and1 | f_arrdiv32_fs220_and0;
  assign f_arrdiv32_fs221_xor0 = f_arrdiv32_mux2to1183_xor0 ^ b[29];
  assign f_arrdiv32_fs221_not0 = ~f_arrdiv32_mux2to1183_xor0;
  assign f_arrdiv32_fs221_and0 = f_arrdiv32_fs221_not0 & b[29];
  assign f_arrdiv32_fs221_xor1 = f_arrdiv32_fs220_or0 ^ f_arrdiv32_fs221_xor0;
  assign f_arrdiv32_fs221_not1 = ~f_arrdiv32_fs221_xor0;
  assign f_arrdiv32_fs221_and1 = f_arrdiv32_fs221_not1 & f_arrdiv32_fs220_or0;
  assign f_arrdiv32_fs221_or0 = f_arrdiv32_fs221_and1 | f_arrdiv32_fs221_and0;
  assign f_arrdiv32_fs222_xor0 = f_arrdiv32_mux2to1184_xor0 ^ b[30];
  assign f_arrdiv32_fs222_not0 = ~f_arrdiv32_mux2to1184_xor0;
  assign f_arrdiv32_fs222_and0 = f_arrdiv32_fs222_not0 & b[30];
  assign f_arrdiv32_fs222_xor1 = f_arrdiv32_fs221_or0 ^ f_arrdiv32_fs222_xor0;
  assign f_arrdiv32_fs222_not1 = ~f_arrdiv32_fs222_xor0;
  assign f_arrdiv32_fs222_and1 = f_arrdiv32_fs222_not1 & f_arrdiv32_fs221_or0;
  assign f_arrdiv32_fs222_or0 = f_arrdiv32_fs222_and1 | f_arrdiv32_fs222_and0;
  assign f_arrdiv32_fs223_xor0 = f_arrdiv32_mux2to1185_xor0 ^ b[31];
  assign f_arrdiv32_fs223_not0 = ~f_arrdiv32_mux2to1185_xor0;
  assign f_arrdiv32_fs223_and0 = f_arrdiv32_fs223_not0 & b[31];
  assign f_arrdiv32_fs223_xor1 = f_arrdiv32_fs222_or0 ^ f_arrdiv32_fs223_xor0;
  assign f_arrdiv32_fs223_not1 = ~f_arrdiv32_fs223_xor0;
  assign f_arrdiv32_fs223_and1 = f_arrdiv32_fs223_not1 & f_arrdiv32_fs222_or0;
  assign f_arrdiv32_fs223_or0 = f_arrdiv32_fs223_and1 | f_arrdiv32_fs223_and0;
  assign f_arrdiv32_mux2to1186_and0 = a[25] & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1186_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1186_and1 = f_arrdiv32_fs192_xor0 & f_arrdiv32_mux2to1186_not0;
  assign f_arrdiv32_mux2to1186_xor0 = f_arrdiv32_mux2to1186_and0 ^ f_arrdiv32_mux2to1186_and1;
  assign f_arrdiv32_mux2to1187_and0 = f_arrdiv32_mux2to1155_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1187_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1187_and1 = f_arrdiv32_fs193_xor1 & f_arrdiv32_mux2to1187_not0;
  assign f_arrdiv32_mux2to1187_xor0 = f_arrdiv32_mux2to1187_and0 ^ f_arrdiv32_mux2to1187_and1;
  assign f_arrdiv32_mux2to1188_and0 = f_arrdiv32_mux2to1156_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1188_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1188_and1 = f_arrdiv32_fs194_xor1 & f_arrdiv32_mux2to1188_not0;
  assign f_arrdiv32_mux2to1188_xor0 = f_arrdiv32_mux2to1188_and0 ^ f_arrdiv32_mux2to1188_and1;
  assign f_arrdiv32_mux2to1189_and0 = f_arrdiv32_mux2to1157_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1189_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1189_and1 = f_arrdiv32_fs195_xor1 & f_arrdiv32_mux2to1189_not0;
  assign f_arrdiv32_mux2to1189_xor0 = f_arrdiv32_mux2to1189_and0 ^ f_arrdiv32_mux2to1189_and1;
  assign f_arrdiv32_mux2to1190_and0 = f_arrdiv32_mux2to1158_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1190_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1190_and1 = f_arrdiv32_fs196_xor1 & f_arrdiv32_mux2to1190_not0;
  assign f_arrdiv32_mux2to1190_xor0 = f_arrdiv32_mux2to1190_and0 ^ f_arrdiv32_mux2to1190_and1;
  assign f_arrdiv32_mux2to1191_and0 = f_arrdiv32_mux2to1159_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1191_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1191_and1 = f_arrdiv32_fs197_xor1 & f_arrdiv32_mux2to1191_not0;
  assign f_arrdiv32_mux2to1191_xor0 = f_arrdiv32_mux2to1191_and0 ^ f_arrdiv32_mux2to1191_and1;
  assign f_arrdiv32_mux2to1192_and0 = f_arrdiv32_mux2to1160_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1192_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1192_and1 = f_arrdiv32_fs198_xor1 & f_arrdiv32_mux2to1192_not0;
  assign f_arrdiv32_mux2to1192_xor0 = f_arrdiv32_mux2to1192_and0 ^ f_arrdiv32_mux2to1192_and1;
  assign f_arrdiv32_mux2to1193_and0 = f_arrdiv32_mux2to1161_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1193_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1193_and1 = f_arrdiv32_fs199_xor1 & f_arrdiv32_mux2to1193_not0;
  assign f_arrdiv32_mux2to1193_xor0 = f_arrdiv32_mux2to1193_and0 ^ f_arrdiv32_mux2to1193_and1;
  assign f_arrdiv32_mux2to1194_and0 = f_arrdiv32_mux2to1162_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1194_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1194_and1 = f_arrdiv32_fs200_xor1 & f_arrdiv32_mux2to1194_not0;
  assign f_arrdiv32_mux2to1194_xor0 = f_arrdiv32_mux2to1194_and0 ^ f_arrdiv32_mux2to1194_and1;
  assign f_arrdiv32_mux2to1195_and0 = f_arrdiv32_mux2to1163_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1195_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1195_and1 = f_arrdiv32_fs201_xor1 & f_arrdiv32_mux2to1195_not0;
  assign f_arrdiv32_mux2to1195_xor0 = f_arrdiv32_mux2to1195_and0 ^ f_arrdiv32_mux2to1195_and1;
  assign f_arrdiv32_mux2to1196_and0 = f_arrdiv32_mux2to1164_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1196_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1196_and1 = f_arrdiv32_fs202_xor1 & f_arrdiv32_mux2to1196_not0;
  assign f_arrdiv32_mux2to1196_xor0 = f_arrdiv32_mux2to1196_and0 ^ f_arrdiv32_mux2to1196_and1;
  assign f_arrdiv32_mux2to1197_and0 = f_arrdiv32_mux2to1165_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1197_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1197_and1 = f_arrdiv32_fs203_xor1 & f_arrdiv32_mux2to1197_not0;
  assign f_arrdiv32_mux2to1197_xor0 = f_arrdiv32_mux2to1197_and0 ^ f_arrdiv32_mux2to1197_and1;
  assign f_arrdiv32_mux2to1198_and0 = f_arrdiv32_mux2to1166_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1198_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1198_and1 = f_arrdiv32_fs204_xor1 & f_arrdiv32_mux2to1198_not0;
  assign f_arrdiv32_mux2to1198_xor0 = f_arrdiv32_mux2to1198_and0 ^ f_arrdiv32_mux2to1198_and1;
  assign f_arrdiv32_mux2to1199_and0 = f_arrdiv32_mux2to1167_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1199_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1199_and1 = f_arrdiv32_fs205_xor1 & f_arrdiv32_mux2to1199_not0;
  assign f_arrdiv32_mux2to1199_xor0 = f_arrdiv32_mux2to1199_and0 ^ f_arrdiv32_mux2to1199_and1;
  assign f_arrdiv32_mux2to1200_and0 = f_arrdiv32_mux2to1168_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1200_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1200_and1 = f_arrdiv32_fs206_xor1 & f_arrdiv32_mux2to1200_not0;
  assign f_arrdiv32_mux2to1200_xor0 = f_arrdiv32_mux2to1200_and0 ^ f_arrdiv32_mux2to1200_and1;
  assign f_arrdiv32_mux2to1201_and0 = f_arrdiv32_mux2to1169_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1201_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1201_and1 = f_arrdiv32_fs207_xor1 & f_arrdiv32_mux2to1201_not0;
  assign f_arrdiv32_mux2to1201_xor0 = f_arrdiv32_mux2to1201_and0 ^ f_arrdiv32_mux2to1201_and1;
  assign f_arrdiv32_mux2to1202_and0 = f_arrdiv32_mux2to1170_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1202_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1202_and1 = f_arrdiv32_fs208_xor1 & f_arrdiv32_mux2to1202_not0;
  assign f_arrdiv32_mux2to1202_xor0 = f_arrdiv32_mux2to1202_and0 ^ f_arrdiv32_mux2to1202_and1;
  assign f_arrdiv32_mux2to1203_and0 = f_arrdiv32_mux2to1171_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1203_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1203_and1 = f_arrdiv32_fs209_xor1 & f_arrdiv32_mux2to1203_not0;
  assign f_arrdiv32_mux2to1203_xor0 = f_arrdiv32_mux2to1203_and0 ^ f_arrdiv32_mux2to1203_and1;
  assign f_arrdiv32_mux2to1204_and0 = f_arrdiv32_mux2to1172_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1204_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1204_and1 = f_arrdiv32_fs210_xor1 & f_arrdiv32_mux2to1204_not0;
  assign f_arrdiv32_mux2to1204_xor0 = f_arrdiv32_mux2to1204_and0 ^ f_arrdiv32_mux2to1204_and1;
  assign f_arrdiv32_mux2to1205_and0 = f_arrdiv32_mux2to1173_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1205_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1205_and1 = f_arrdiv32_fs211_xor1 & f_arrdiv32_mux2to1205_not0;
  assign f_arrdiv32_mux2to1205_xor0 = f_arrdiv32_mux2to1205_and0 ^ f_arrdiv32_mux2to1205_and1;
  assign f_arrdiv32_mux2to1206_and0 = f_arrdiv32_mux2to1174_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1206_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1206_and1 = f_arrdiv32_fs212_xor1 & f_arrdiv32_mux2to1206_not0;
  assign f_arrdiv32_mux2to1206_xor0 = f_arrdiv32_mux2to1206_and0 ^ f_arrdiv32_mux2to1206_and1;
  assign f_arrdiv32_mux2to1207_and0 = f_arrdiv32_mux2to1175_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1207_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1207_and1 = f_arrdiv32_fs213_xor1 & f_arrdiv32_mux2to1207_not0;
  assign f_arrdiv32_mux2to1207_xor0 = f_arrdiv32_mux2to1207_and0 ^ f_arrdiv32_mux2to1207_and1;
  assign f_arrdiv32_mux2to1208_and0 = f_arrdiv32_mux2to1176_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1208_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1208_and1 = f_arrdiv32_fs214_xor1 & f_arrdiv32_mux2to1208_not0;
  assign f_arrdiv32_mux2to1208_xor0 = f_arrdiv32_mux2to1208_and0 ^ f_arrdiv32_mux2to1208_and1;
  assign f_arrdiv32_mux2to1209_and0 = f_arrdiv32_mux2to1177_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1209_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1209_and1 = f_arrdiv32_fs215_xor1 & f_arrdiv32_mux2to1209_not0;
  assign f_arrdiv32_mux2to1209_xor0 = f_arrdiv32_mux2to1209_and0 ^ f_arrdiv32_mux2to1209_and1;
  assign f_arrdiv32_mux2to1210_and0 = f_arrdiv32_mux2to1178_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1210_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1210_and1 = f_arrdiv32_fs216_xor1 & f_arrdiv32_mux2to1210_not0;
  assign f_arrdiv32_mux2to1210_xor0 = f_arrdiv32_mux2to1210_and0 ^ f_arrdiv32_mux2to1210_and1;
  assign f_arrdiv32_mux2to1211_and0 = f_arrdiv32_mux2to1179_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1211_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1211_and1 = f_arrdiv32_fs217_xor1 & f_arrdiv32_mux2to1211_not0;
  assign f_arrdiv32_mux2to1211_xor0 = f_arrdiv32_mux2to1211_and0 ^ f_arrdiv32_mux2to1211_and1;
  assign f_arrdiv32_mux2to1212_and0 = f_arrdiv32_mux2to1180_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1212_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1212_and1 = f_arrdiv32_fs218_xor1 & f_arrdiv32_mux2to1212_not0;
  assign f_arrdiv32_mux2to1212_xor0 = f_arrdiv32_mux2to1212_and0 ^ f_arrdiv32_mux2to1212_and1;
  assign f_arrdiv32_mux2to1213_and0 = f_arrdiv32_mux2to1181_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1213_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1213_and1 = f_arrdiv32_fs219_xor1 & f_arrdiv32_mux2to1213_not0;
  assign f_arrdiv32_mux2to1213_xor0 = f_arrdiv32_mux2to1213_and0 ^ f_arrdiv32_mux2to1213_and1;
  assign f_arrdiv32_mux2to1214_and0 = f_arrdiv32_mux2to1182_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1214_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1214_and1 = f_arrdiv32_fs220_xor1 & f_arrdiv32_mux2to1214_not0;
  assign f_arrdiv32_mux2to1214_xor0 = f_arrdiv32_mux2to1214_and0 ^ f_arrdiv32_mux2to1214_and1;
  assign f_arrdiv32_mux2to1215_and0 = f_arrdiv32_mux2to1183_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1215_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1215_and1 = f_arrdiv32_fs221_xor1 & f_arrdiv32_mux2to1215_not0;
  assign f_arrdiv32_mux2to1215_xor0 = f_arrdiv32_mux2to1215_and0 ^ f_arrdiv32_mux2to1215_and1;
  assign f_arrdiv32_mux2to1216_and0 = f_arrdiv32_mux2to1184_xor0 & f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1216_not0 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_mux2to1216_and1 = f_arrdiv32_fs222_xor1 & f_arrdiv32_mux2to1216_not0;
  assign f_arrdiv32_mux2to1216_xor0 = f_arrdiv32_mux2to1216_and0 ^ f_arrdiv32_mux2to1216_and1;
  assign f_arrdiv32_not6 = ~f_arrdiv32_fs223_or0;
  assign f_arrdiv32_fs224_xor0 = a[24] ^ b[0];
  assign f_arrdiv32_fs224_not0 = ~a[24];
  assign f_arrdiv32_fs224_and0 = f_arrdiv32_fs224_not0 & b[0];
  assign f_arrdiv32_fs224_not1 = ~f_arrdiv32_fs224_xor0;
  assign f_arrdiv32_fs225_xor0 = f_arrdiv32_mux2to1186_xor0 ^ b[1];
  assign f_arrdiv32_fs225_not0 = ~f_arrdiv32_mux2to1186_xor0;
  assign f_arrdiv32_fs225_and0 = f_arrdiv32_fs225_not0 & b[1];
  assign f_arrdiv32_fs225_xor1 = f_arrdiv32_fs224_and0 ^ f_arrdiv32_fs225_xor0;
  assign f_arrdiv32_fs225_not1 = ~f_arrdiv32_fs225_xor0;
  assign f_arrdiv32_fs225_and1 = f_arrdiv32_fs225_not1 & f_arrdiv32_fs224_and0;
  assign f_arrdiv32_fs225_or0 = f_arrdiv32_fs225_and1 | f_arrdiv32_fs225_and0;
  assign f_arrdiv32_fs226_xor0 = f_arrdiv32_mux2to1187_xor0 ^ b[2];
  assign f_arrdiv32_fs226_not0 = ~f_arrdiv32_mux2to1187_xor0;
  assign f_arrdiv32_fs226_and0 = f_arrdiv32_fs226_not0 & b[2];
  assign f_arrdiv32_fs226_xor1 = f_arrdiv32_fs225_or0 ^ f_arrdiv32_fs226_xor0;
  assign f_arrdiv32_fs226_not1 = ~f_arrdiv32_fs226_xor0;
  assign f_arrdiv32_fs226_and1 = f_arrdiv32_fs226_not1 & f_arrdiv32_fs225_or0;
  assign f_arrdiv32_fs226_or0 = f_arrdiv32_fs226_and1 | f_arrdiv32_fs226_and0;
  assign f_arrdiv32_fs227_xor0 = f_arrdiv32_mux2to1188_xor0 ^ b[3];
  assign f_arrdiv32_fs227_not0 = ~f_arrdiv32_mux2to1188_xor0;
  assign f_arrdiv32_fs227_and0 = f_arrdiv32_fs227_not0 & b[3];
  assign f_arrdiv32_fs227_xor1 = f_arrdiv32_fs226_or0 ^ f_arrdiv32_fs227_xor0;
  assign f_arrdiv32_fs227_not1 = ~f_arrdiv32_fs227_xor0;
  assign f_arrdiv32_fs227_and1 = f_arrdiv32_fs227_not1 & f_arrdiv32_fs226_or0;
  assign f_arrdiv32_fs227_or0 = f_arrdiv32_fs227_and1 | f_arrdiv32_fs227_and0;
  assign f_arrdiv32_fs228_xor0 = f_arrdiv32_mux2to1189_xor0 ^ b[4];
  assign f_arrdiv32_fs228_not0 = ~f_arrdiv32_mux2to1189_xor0;
  assign f_arrdiv32_fs228_and0 = f_arrdiv32_fs228_not0 & b[4];
  assign f_arrdiv32_fs228_xor1 = f_arrdiv32_fs227_or0 ^ f_arrdiv32_fs228_xor0;
  assign f_arrdiv32_fs228_not1 = ~f_arrdiv32_fs228_xor0;
  assign f_arrdiv32_fs228_and1 = f_arrdiv32_fs228_not1 & f_arrdiv32_fs227_or0;
  assign f_arrdiv32_fs228_or0 = f_arrdiv32_fs228_and1 | f_arrdiv32_fs228_and0;
  assign f_arrdiv32_fs229_xor0 = f_arrdiv32_mux2to1190_xor0 ^ b[5];
  assign f_arrdiv32_fs229_not0 = ~f_arrdiv32_mux2to1190_xor0;
  assign f_arrdiv32_fs229_and0 = f_arrdiv32_fs229_not0 & b[5];
  assign f_arrdiv32_fs229_xor1 = f_arrdiv32_fs228_or0 ^ f_arrdiv32_fs229_xor0;
  assign f_arrdiv32_fs229_not1 = ~f_arrdiv32_fs229_xor0;
  assign f_arrdiv32_fs229_and1 = f_arrdiv32_fs229_not1 & f_arrdiv32_fs228_or0;
  assign f_arrdiv32_fs229_or0 = f_arrdiv32_fs229_and1 | f_arrdiv32_fs229_and0;
  assign f_arrdiv32_fs230_xor0 = f_arrdiv32_mux2to1191_xor0 ^ b[6];
  assign f_arrdiv32_fs230_not0 = ~f_arrdiv32_mux2to1191_xor0;
  assign f_arrdiv32_fs230_and0 = f_arrdiv32_fs230_not0 & b[6];
  assign f_arrdiv32_fs230_xor1 = f_arrdiv32_fs229_or0 ^ f_arrdiv32_fs230_xor0;
  assign f_arrdiv32_fs230_not1 = ~f_arrdiv32_fs230_xor0;
  assign f_arrdiv32_fs230_and1 = f_arrdiv32_fs230_not1 & f_arrdiv32_fs229_or0;
  assign f_arrdiv32_fs230_or0 = f_arrdiv32_fs230_and1 | f_arrdiv32_fs230_and0;
  assign f_arrdiv32_fs231_xor0 = f_arrdiv32_mux2to1192_xor0 ^ b[7];
  assign f_arrdiv32_fs231_not0 = ~f_arrdiv32_mux2to1192_xor0;
  assign f_arrdiv32_fs231_and0 = f_arrdiv32_fs231_not0 & b[7];
  assign f_arrdiv32_fs231_xor1 = f_arrdiv32_fs230_or0 ^ f_arrdiv32_fs231_xor0;
  assign f_arrdiv32_fs231_not1 = ~f_arrdiv32_fs231_xor0;
  assign f_arrdiv32_fs231_and1 = f_arrdiv32_fs231_not1 & f_arrdiv32_fs230_or0;
  assign f_arrdiv32_fs231_or0 = f_arrdiv32_fs231_and1 | f_arrdiv32_fs231_and0;
  assign f_arrdiv32_fs232_xor0 = f_arrdiv32_mux2to1193_xor0 ^ b[8];
  assign f_arrdiv32_fs232_not0 = ~f_arrdiv32_mux2to1193_xor0;
  assign f_arrdiv32_fs232_and0 = f_arrdiv32_fs232_not0 & b[8];
  assign f_arrdiv32_fs232_xor1 = f_arrdiv32_fs231_or0 ^ f_arrdiv32_fs232_xor0;
  assign f_arrdiv32_fs232_not1 = ~f_arrdiv32_fs232_xor0;
  assign f_arrdiv32_fs232_and1 = f_arrdiv32_fs232_not1 & f_arrdiv32_fs231_or0;
  assign f_arrdiv32_fs232_or0 = f_arrdiv32_fs232_and1 | f_arrdiv32_fs232_and0;
  assign f_arrdiv32_fs233_xor0 = f_arrdiv32_mux2to1194_xor0 ^ b[9];
  assign f_arrdiv32_fs233_not0 = ~f_arrdiv32_mux2to1194_xor0;
  assign f_arrdiv32_fs233_and0 = f_arrdiv32_fs233_not0 & b[9];
  assign f_arrdiv32_fs233_xor1 = f_arrdiv32_fs232_or0 ^ f_arrdiv32_fs233_xor0;
  assign f_arrdiv32_fs233_not1 = ~f_arrdiv32_fs233_xor0;
  assign f_arrdiv32_fs233_and1 = f_arrdiv32_fs233_not1 & f_arrdiv32_fs232_or0;
  assign f_arrdiv32_fs233_or0 = f_arrdiv32_fs233_and1 | f_arrdiv32_fs233_and0;
  assign f_arrdiv32_fs234_xor0 = f_arrdiv32_mux2to1195_xor0 ^ b[10];
  assign f_arrdiv32_fs234_not0 = ~f_arrdiv32_mux2to1195_xor0;
  assign f_arrdiv32_fs234_and0 = f_arrdiv32_fs234_not0 & b[10];
  assign f_arrdiv32_fs234_xor1 = f_arrdiv32_fs233_or0 ^ f_arrdiv32_fs234_xor0;
  assign f_arrdiv32_fs234_not1 = ~f_arrdiv32_fs234_xor0;
  assign f_arrdiv32_fs234_and1 = f_arrdiv32_fs234_not1 & f_arrdiv32_fs233_or0;
  assign f_arrdiv32_fs234_or0 = f_arrdiv32_fs234_and1 | f_arrdiv32_fs234_and0;
  assign f_arrdiv32_fs235_xor0 = f_arrdiv32_mux2to1196_xor0 ^ b[11];
  assign f_arrdiv32_fs235_not0 = ~f_arrdiv32_mux2to1196_xor0;
  assign f_arrdiv32_fs235_and0 = f_arrdiv32_fs235_not0 & b[11];
  assign f_arrdiv32_fs235_xor1 = f_arrdiv32_fs234_or0 ^ f_arrdiv32_fs235_xor0;
  assign f_arrdiv32_fs235_not1 = ~f_arrdiv32_fs235_xor0;
  assign f_arrdiv32_fs235_and1 = f_arrdiv32_fs235_not1 & f_arrdiv32_fs234_or0;
  assign f_arrdiv32_fs235_or0 = f_arrdiv32_fs235_and1 | f_arrdiv32_fs235_and0;
  assign f_arrdiv32_fs236_xor0 = f_arrdiv32_mux2to1197_xor0 ^ b[12];
  assign f_arrdiv32_fs236_not0 = ~f_arrdiv32_mux2to1197_xor0;
  assign f_arrdiv32_fs236_and0 = f_arrdiv32_fs236_not0 & b[12];
  assign f_arrdiv32_fs236_xor1 = f_arrdiv32_fs235_or0 ^ f_arrdiv32_fs236_xor0;
  assign f_arrdiv32_fs236_not1 = ~f_arrdiv32_fs236_xor0;
  assign f_arrdiv32_fs236_and1 = f_arrdiv32_fs236_not1 & f_arrdiv32_fs235_or0;
  assign f_arrdiv32_fs236_or0 = f_arrdiv32_fs236_and1 | f_arrdiv32_fs236_and0;
  assign f_arrdiv32_fs237_xor0 = f_arrdiv32_mux2to1198_xor0 ^ b[13];
  assign f_arrdiv32_fs237_not0 = ~f_arrdiv32_mux2to1198_xor0;
  assign f_arrdiv32_fs237_and0 = f_arrdiv32_fs237_not0 & b[13];
  assign f_arrdiv32_fs237_xor1 = f_arrdiv32_fs236_or0 ^ f_arrdiv32_fs237_xor0;
  assign f_arrdiv32_fs237_not1 = ~f_arrdiv32_fs237_xor0;
  assign f_arrdiv32_fs237_and1 = f_arrdiv32_fs237_not1 & f_arrdiv32_fs236_or0;
  assign f_arrdiv32_fs237_or0 = f_arrdiv32_fs237_and1 | f_arrdiv32_fs237_and0;
  assign f_arrdiv32_fs238_xor0 = f_arrdiv32_mux2to1199_xor0 ^ b[14];
  assign f_arrdiv32_fs238_not0 = ~f_arrdiv32_mux2to1199_xor0;
  assign f_arrdiv32_fs238_and0 = f_arrdiv32_fs238_not0 & b[14];
  assign f_arrdiv32_fs238_xor1 = f_arrdiv32_fs237_or0 ^ f_arrdiv32_fs238_xor0;
  assign f_arrdiv32_fs238_not1 = ~f_arrdiv32_fs238_xor0;
  assign f_arrdiv32_fs238_and1 = f_arrdiv32_fs238_not1 & f_arrdiv32_fs237_or0;
  assign f_arrdiv32_fs238_or0 = f_arrdiv32_fs238_and1 | f_arrdiv32_fs238_and0;
  assign f_arrdiv32_fs239_xor0 = f_arrdiv32_mux2to1200_xor0 ^ b[15];
  assign f_arrdiv32_fs239_not0 = ~f_arrdiv32_mux2to1200_xor0;
  assign f_arrdiv32_fs239_and0 = f_arrdiv32_fs239_not0 & b[15];
  assign f_arrdiv32_fs239_xor1 = f_arrdiv32_fs238_or0 ^ f_arrdiv32_fs239_xor0;
  assign f_arrdiv32_fs239_not1 = ~f_arrdiv32_fs239_xor0;
  assign f_arrdiv32_fs239_and1 = f_arrdiv32_fs239_not1 & f_arrdiv32_fs238_or0;
  assign f_arrdiv32_fs239_or0 = f_arrdiv32_fs239_and1 | f_arrdiv32_fs239_and0;
  assign f_arrdiv32_fs240_xor0 = f_arrdiv32_mux2to1201_xor0 ^ b[16];
  assign f_arrdiv32_fs240_not0 = ~f_arrdiv32_mux2to1201_xor0;
  assign f_arrdiv32_fs240_and0 = f_arrdiv32_fs240_not0 & b[16];
  assign f_arrdiv32_fs240_xor1 = f_arrdiv32_fs239_or0 ^ f_arrdiv32_fs240_xor0;
  assign f_arrdiv32_fs240_not1 = ~f_arrdiv32_fs240_xor0;
  assign f_arrdiv32_fs240_and1 = f_arrdiv32_fs240_not1 & f_arrdiv32_fs239_or0;
  assign f_arrdiv32_fs240_or0 = f_arrdiv32_fs240_and1 | f_arrdiv32_fs240_and0;
  assign f_arrdiv32_fs241_xor0 = f_arrdiv32_mux2to1202_xor0 ^ b[17];
  assign f_arrdiv32_fs241_not0 = ~f_arrdiv32_mux2to1202_xor0;
  assign f_arrdiv32_fs241_and0 = f_arrdiv32_fs241_not0 & b[17];
  assign f_arrdiv32_fs241_xor1 = f_arrdiv32_fs240_or0 ^ f_arrdiv32_fs241_xor0;
  assign f_arrdiv32_fs241_not1 = ~f_arrdiv32_fs241_xor0;
  assign f_arrdiv32_fs241_and1 = f_arrdiv32_fs241_not1 & f_arrdiv32_fs240_or0;
  assign f_arrdiv32_fs241_or0 = f_arrdiv32_fs241_and1 | f_arrdiv32_fs241_and0;
  assign f_arrdiv32_fs242_xor0 = f_arrdiv32_mux2to1203_xor0 ^ b[18];
  assign f_arrdiv32_fs242_not0 = ~f_arrdiv32_mux2to1203_xor0;
  assign f_arrdiv32_fs242_and0 = f_arrdiv32_fs242_not0 & b[18];
  assign f_arrdiv32_fs242_xor1 = f_arrdiv32_fs241_or0 ^ f_arrdiv32_fs242_xor0;
  assign f_arrdiv32_fs242_not1 = ~f_arrdiv32_fs242_xor0;
  assign f_arrdiv32_fs242_and1 = f_arrdiv32_fs242_not1 & f_arrdiv32_fs241_or0;
  assign f_arrdiv32_fs242_or0 = f_arrdiv32_fs242_and1 | f_arrdiv32_fs242_and0;
  assign f_arrdiv32_fs243_xor0 = f_arrdiv32_mux2to1204_xor0 ^ b[19];
  assign f_arrdiv32_fs243_not0 = ~f_arrdiv32_mux2to1204_xor0;
  assign f_arrdiv32_fs243_and0 = f_arrdiv32_fs243_not0 & b[19];
  assign f_arrdiv32_fs243_xor1 = f_arrdiv32_fs242_or0 ^ f_arrdiv32_fs243_xor0;
  assign f_arrdiv32_fs243_not1 = ~f_arrdiv32_fs243_xor0;
  assign f_arrdiv32_fs243_and1 = f_arrdiv32_fs243_not1 & f_arrdiv32_fs242_or0;
  assign f_arrdiv32_fs243_or0 = f_arrdiv32_fs243_and1 | f_arrdiv32_fs243_and0;
  assign f_arrdiv32_fs244_xor0 = f_arrdiv32_mux2to1205_xor0 ^ b[20];
  assign f_arrdiv32_fs244_not0 = ~f_arrdiv32_mux2to1205_xor0;
  assign f_arrdiv32_fs244_and0 = f_arrdiv32_fs244_not0 & b[20];
  assign f_arrdiv32_fs244_xor1 = f_arrdiv32_fs243_or0 ^ f_arrdiv32_fs244_xor0;
  assign f_arrdiv32_fs244_not1 = ~f_arrdiv32_fs244_xor0;
  assign f_arrdiv32_fs244_and1 = f_arrdiv32_fs244_not1 & f_arrdiv32_fs243_or0;
  assign f_arrdiv32_fs244_or0 = f_arrdiv32_fs244_and1 | f_arrdiv32_fs244_and0;
  assign f_arrdiv32_fs245_xor0 = f_arrdiv32_mux2to1206_xor0 ^ b[21];
  assign f_arrdiv32_fs245_not0 = ~f_arrdiv32_mux2to1206_xor0;
  assign f_arrdiv32_fs245_and0 = f_arrdiv32_fs245_not0 & b[21];
  assign f_arrdiv32_fs245_xor1 = f_arrdiv32_fs244_or0 ^ f_arrdiv32_fs245_xor0;
  assign f_arrdiv32_fs245_not1 = ~f_arrdiv32_fs245_xor0;
  assign f_arrdiv32_fs245_and1 = f_arrdiv32_fs245_not1 & f_arrdiv32_fs244_or0;
  assign f_arrdiv32_fs245_or0 = f_arrdiv32_fs245_and1 | f_arrdiv32_fs245_and0;
  assign f_arrdiv32_fs246_xor0 = f_arrdiv32_mux2to1207_xor0 ^ b[22];
  assign f_arrdiv32_fs246_not0 = ~f_arrdiv32_mux2to1207_xor0;
  assign f_arrdiv32_fs246_and0 = f_arrdiv32_fs246_not0 & b[22];
  assign f_arrdiv32_fs246_xor1 = f_arrdiv32_fs245_or0 ^ f_arrdiv32_fs246_xor0;
  assign f_arrdiv32_fs246_not1 = ~f_arrdiv32_fs246_xor0;
  assign f_arrdiv32_fs246_and1 = f_arrdiv32_fs246_not1 & f_arrdiv32_fs245_or0;
  assign f_arrdiv32_fs246_or0 = f_arrdiv32_fs246_and1 | f_arrdiv32_fs246_and0;
  assign f_arrdiv32_fs247_xor0 = f_arrdiv32_mux2to1208_xor0 ^ b[23];
  assign f_arrdiv32_fs247_not0 = ~f_arrdiv32_mux2to1208_xor0;
  assign f_arrdiv32_fs247_and0 = f_arrdiv32_fs247_not0 & b[23];
  assign f_arrdiv32_fs247_xor1 = f_arrdiv32_fs246_or0 ^ f_arrdiv32_fs247_xor0;
  assign f_arrdiv32_fs247_not1 = ~f_arrdiv32_fs247_xor0;
  assign f_arrdiv32_fs247_and1 = f_arrdiv32_fs247_not1 & f_arrdiv32_fs246_or0;
  assign f_arrdiv32_fs247_or0 = f_arrdiv32_fs247_and1 | f_arrdiv32_fs247_and0;
  assign f_arrdiv32_fs248_xor0 = f_arrdiv32_mux2to1209_xor0 ^ b[24];
  assign f_arrdiv32_fs248_not0 = ~f_arrdiv32_mux2to1209_xor0;
  assign f_arrdiv32_fs248_and0 = f_arrdiv32_fs248_not0 & b[24];
  assign f_arrdiv32_fs248_xor1 = f_arrdiv32_fs247_or0 ^ f_arrdiv32_fs248_xor0;
  assign f_arrdiv32_fs248_not1 = ~f_arrdiv32_fs248_xor0;
  assign f_arrdiv32_fs248_and1 = f_arrdiv32_fs248_not1 & f_arrdiv32_fs247_or0;
  assign f_arrdiv32_fs248_or0 = f_arrdiv32_fs248_and1 | f_arrdiv32_fs248_and0;
  assign f_arrdiv32_fs249_xor0 = f_arrdiv32_mux2to1210_xor0 ^ b[25];
  assign f_arrdiv32_fs249_not0 = ~f_arrdiv32_mux2to1210_xor0;
  assign f_arrdiv32_fs249_and0 = f_arrdiv32_fs249_not0 & b[25];
  assign f_arrdiv32_fs249_xor1 = f_arrdiv32_fs248_or0 ^ f_arrdiv32_fs249_xor0;
  assign f_arrdiv32_fs249_not1 = ~f_arrdiv32_fs249_xor0;
  assign f_arrdiv32_fs249_and1 = f_arrdiv32_fs249_not1 & f_arrdiv32_fs248_or0;
  assign f_arrdiv32_fs249_or0 = f_arrdiv32_fs249_and1 | f_arrdiv32_fs249_and0;
  assign f_arrdiv32_fs250_xor0 = f_arrdiv32_mux2to1211_xor0 ^ b[26];
  assign f_arrdiv32_fs250_not0 = ~f_arrdiv32_mux2to1211_xor0;
  assign f_arrdiv32_fs250_and0 = f_arrdiv32_fs250_not0 & b[26];
  assign f_arrdiv32_fs250_xor1 = f_arrdiv32_fs249_or0 ^ f_arrdiv32_fs250_xor0;
  assign f_arrdiv32_fs250_not1 = ~f_arrdiv32_fs250_xor0;
  assign f_arrdiv32_fs250_and1 = f_arrdiv32_fs250_not1 & f_arrdiv32_fs249_or0;
  assign f_arrdiv32_fs250_or0 = f_arrdiv32_fs250_and1 | f_arrdiv32_fs250_and0;
  assign f_arrdiv32_fs251_xor0 = f_arrdiv32_mux2to1212_xor0 ^ b[27];
  assign f_arrdiv32_fs251_not0 = ~f_arrdiv32_mux2to1212_xor0;
  assign f_arrdiv32_fs251_and0 = f_arrdiv32_fs251_not0 & b[27];
  assign f_arrdiv32_fs251_xor1 = f_arrdiv32_fs250_or0 ^ f_arrdiv32_fs251_xor0;
  assign f_arrdiv32_fs251_not1 = ~f_arrdiv32_fs251_xor0;
  assign f_arrdiv32_fs251_and1 = f_arrdiv32_fs251_not1 & f_arrdiv32_fs250_or0;
  assign f_arrdiv32_fs251_or0 = f_arrdiv32_fs251_and1 | f_arrdiv32_fs251_and0;
  assign f_arrdiv32_fs252_xor0 = f_arrdiv32_mux2to1213_xor0 ^ b[28];
  assign f_arrdiv32_fs252_not0 = ~f_arrdiv32_mux2to1213_xor0;
  assign f_arrdiv32_fs252_and0 = f_arrdiv32_fs252_not0 & b[28];
  assign f_arrdiv32_fs252_xor1 = f_arrdiv32_fs251_or0 ^ f_arrdiv32_fs252_xor0;
  assign f_arrdiv32_fs252_not1 = ~f_arrdiv32_fs252_xor0;
  assign f_arrdiv32_fs252_and1 = f_arrdiv32_fs252_not1 & f_arrdiv32_fs251_or0;
  assign f_arrdiv32_fs252_or0 = f_arrdiv32_fs252_and1 | f_arrdiv32_fs252_and0;
  assign f_arrdiv32_fs253_xor0 = f_arrdiv32_mux2to1214_xor0 ^ b[29];
  assign f_arrdiv32_fs253_not0 = ~f_arrdiv32_mux2to1214_xor0;
  assign f_arrdiv32_fs253_and0 = f_arrdiv32_fs253_not0 & b[29];
  assign f_arrdiv32_fs253_xor1 = f_arrdiv32_fs252_or0 ^ f_arrdiv32_fs253_xor0;
  assign f_arrdiv32_fs253_not1 = ~f_arrdiv32_fs253_xor0;
  assign f_arrdiv32_fs253_and1 = f_arrdiv32_fs253_not1 & f_arrdiv32_fs252_or0;
  assign f_arrdiv32_fs253_or0 = f_arrdiv32_fs253_and1 | f_arrdiv32_fs253_and0;
  assign f_arrdiv32_fs254_xor0 = f_arrdiv32_mux2to1215_xor0 ^ b[30];
  assign f_arrdiv32_fs254_not0 = ~f_arrdiv32_mux2to1215_xor0;
  assign f_arrdiv32_fs254_and0 = f_arrdiv32_fs254_not0 & b[30];
  assign f_arrdiv32_fs254_xor1 = f_arrdiv32_fs253_or0 ^ f_arrdiv32_fs254_xor0;
  assign f_arrdiv32_fs254_not1 = ~f_arrdiv32_fs254_xor0;
  assign f_arrdiv32_fs254_and1 = f_arrdiv32_fs254_not1 & f_arrdiv32_fs253_or0;
  assign f_arrdiv32_fs254_or0 = f_arrdiv32_fs254_and1 | f_arrdiv32_fs254_and0;
  assign f_arrdiv32_fs255_xor0 = f_arrdiv32_mux2to1216_xor0 ^ b[31];
  assign f_arrdiv32_fs255_not0 = ~f_arrdiv32_mux2to1216_xor0;
  assign f_arrdiv32_fs255_and0 = f_arrdiv32_fs255_not0 & b[31];
  assign f_arrdiv32_fs255_xor1 = f_arrdiv32_fs254_or0 ^ f_arrdiv32_fs255_xor0;
  assign f_arrdiv32_fs255_not1 = ~f_arrdiv32_fs255_xor0;
  assign f_arrdiv32_fs255_and1 = f_arrdiv32_fs255_not1 & f_arrdiv32_fs254_or0;
  assign f_arrdiv32_fs255_or0 = f_arrdiv32_fs255_and1 | f_arrdiv32_fs255_and0;
  assign f_arrdiv32_mux2to1217_and0 = a[24] & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1217_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1217_and1 = f_arrdiv32_fs224_xor0 & f_arrdiv32_mux2to1217_not0;
  assign f_arrdiv32_mux2to1217_xor0 = f_arrdiv32_mux2to1217_and0 ^ f_arrdiv32_mux2to1217_and1;
  assign f_arrdiv32_mux2to1218_and0 = f_arrdiv32_mux2to1186_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1218_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1218_and1 = f_arrdiv32_fs225_xor1 & f_arrdiv32_mux2to1218_not0;
  assign f_arrdiv32_mux2to1218_xor0 = f_arrdiv32_mux2to1218_and0 ^ f_arrdiv32_mux2to1218_and1;
  assign f_arrdiv32_mux2to1219_and0 = f_arrdiv32_mux2to1187_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1219_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1219_and1 = f_arrdiv32_fs226_xor1 & f_arrdiv32_mux2to1219_not0;
  assign f_arrdiv32_mux2to1219_xor0 = f_arrdiv32_mux2to1219_and0 ^ f_arrdiv32_mux2to1219_and1;
  assign f_arrdiv32_mux2to1220_and0 = f_arrdiv32_mux2to1188_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1220_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1220_and1 = f_arrdiv32_fs227_xor1 & f_arrdiv32_mux2to1220_not0;
  assign f_arrdiv32_mux2to1220_xor0 = f_arrdiv32_mux2to1220_and0 ^ f_arrdiv32_mux2to1220_and1;
  assign f_arrdiv32_mux2to1221_and0 = f_arrdiv32_mux2to1189_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1221_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1221_and1 = f_arrdiv32_fs228_xor1 & f_arrdiv32_mux2to1221_not0;
  assign f_arrdiv32_mux2to1221_xor0 = f_arrdiv32_mux2to1221_and0 ^ f_arrdiv32_mux2to1221_and1;
  assign f_arrdiv32_mux2to1222_and0 = f_arrdiv32_mux2to1190_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1222_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1222_and1 = f_arrdiv32_fs229_xor1 & f_arrdiv32_mux2to1222_not0;
  assign f_arrdiv32_mux2to1222_xor0 = f_arrdiv32_mux2to1222_and0 ^ f_arrdiv32_mux2to1222_and1;
  assign f_arrdiv32_mux2to1223_and0 = f_arrdiv32_mux2to1191_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1223_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1223_and1 = f_arrdiv32_fs230_xor1 & f_arrdiv32_mux2to1223_not0;
  assign f_arrdiv32_mux2to1223_xor0 = f_arrdiv32_mux2to1223_and0 ^ f_arrdiv32_mux2to1223_and1;
  assign f_arrdiv32_mux2to1224_and0 = f_arrdiv32_mux2to1192_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1224_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1224_and1 = f_arrdiv32_fs231_xor1 & f_arrdiv32_mux2to1224_not0;
  assign f_arrdiv32_mux2to1224_xor0 = f_arrdiv32_mux2to1224_and0 ^ f_arrdiv32_mux2to1224_and1;
  assign f_arrdiv32_mux2to1225_and0 = f_arrdiv32_mux2to1193_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1225_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1225_and1 = f_arrdiv32_fs232_xor1 & f_arrdiv32_mux2to1225_not0;
  assign f_arrdiv32_mux2to1225_xor0 = f_arrdiv32_mux2to1225_and0 ^ f_arrdiv32_mux2to1225_and1;
  assign f_arrdiv32_mux2to1226_and0 = f_arrdiv32_mux2to1194_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1226_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1226_and1 = f_arrdiv32_fs233_xor1 & f_arrdiv32_mux2to1226_not0;
  assign f_arrdiv32_mux2to1226_xor0 = f_arrdiv32_mux2to1226_and0 ^ f_arrdiv32_mux2to1226_and1;
  assign f_arrdiv32_mux2to1227_and0 = f_arrdiv32_mux2to1195_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1227_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1227_and1 = f_arrdiv32_fs234_xor1 & f_arrdiv32_mux2to1227_not0;
  assign f_arrdiv32_mux2to1227_xor0 = f_arrdiv32_mux2to1227_and0 ^ f_arrdiv32_mux2to1227_and1;
  assign f_arrdiv32_mux2to1228_and0 = f_arrdiv32_mux2to1196_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1228_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1228_and1 = f_arrdiv32_fs235_xor1 & f_arrdiv32_mux2to1228_not0;
  assign f_arrdiv32_mux2to1228_xor0 = f_arrdiv32_mux2to1228_and0 ^ f_arrdiv32_mux2to1228_and1;
  assign f_arrdiv32_mux2to1229_and0 = f_arrdiv32_mux2to1197_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1229_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1229_and1 = f_arrdiv32_fs236_xor1 & f_arrdiv32_mux2to1229_not0;
  assign f_arrdiv32_mux2to1229_xor0 = f_arrdiv32_mux2to1229_and0 ^ f_arrdiv32_mux2to1229_and1;
  assign f_arrdiv32_mux2to1230_and0 = f_arrdiv32_mux2to1198_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1230_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1230_and1 = f_arrdiv32_fs237_xor1 & f_arrdiv32_mux2to1230_not0;
  assign f_arrdiv32_mux2to1230_xor0 = f_arrdiv32_mux2to1230_and0 ^ f_arrdiv32_mux2to1230_and1;
  assign f_arrdiv32_mux2to1231_and0 = f_arrdiv32_mux2to1199_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1231_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1231_and1 = f_arrdiv32_fs238_xor1 & f_arrdiv32_mux2to1231_not0;
  assign f_arrdiv32_mux2to1231_xor0 = f_arrdiv32_mux2to1231_and0 ^ f_arrdiv32_mux2to1231_and1;
  assign f_arrdiv32_mux2to1232_and0 = f_arrdiv32_mux2to1200_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1232_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1232_and1 = f_arrdiv32_fs239_xor1 & f_arrdiv32_mux2to1232_not0;
  assign f_arrdiv32_mux2to1232_xor0 = f_arrdiv32_mux2to1232_and0 ^ f_arrdiv32_mux2to1232_and1;
  assign f_arrdiv32_mux2to1233_and0 = f_arrdiv32_mux2to1201_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1233_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1233_and1 = f_arrdiv32_fs240_xor1 & f_arrdiv32_mux2to1233_not0;
  assign f_arrdiv32_mux2to1233_xor0 = f_arrdiv32_mux2to1233_and0 ^ f_arrdiv32_mux2to1233_and1;
  assign f_arrdiv32_mux2to1234_and0 = f_arrdiv32_mux2to1202_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1234_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1234_and1 = f_arrdiv32_fs241_xor1 & f_arrdiv32_mux2to1234_not0;
  assign f_arrdiv32_mux2to1234_xor0 = f_arrdiv32_mux2to1234_and0 ^ f_arrdiv32_mux2to1234_and1;
  assign f_arrdiv32_mux2to1235_and0 = f_arrdiv32_mux2to1203_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1235_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1235_and1 = f_arrdiv32_fs242_xor1 & f_arrdiv32_mux2to1235_not0;
  assign f_arrdiv32_mux2to1235_xor0 = f_arrdiv32_mux2to1235_and0 ^ f_arrdiv32_mux2to1235_and1;
  assign f_arrdiv32_mux2to1236_and0 = f_arrdiv32_mux2to1204_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1236_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1236_and1 = f_arrdiv32_fs243_xor1 & f_arrdiv32_mux2to1236_not0;
  assign f_arrdiv32_mux2to1236_xor0 = f_arrdiv32_mux2to1236_and0 ^ f_arrdiv32_mux2to1236_and1;
  assign f_arrdiv32_mux2to1237_and0 = f_arrdiv32_mux2to1205_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1237_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1237_and1 = f_arrdiv32_fs244_xor1 & f_arrdiv32_mux2to1237_not0;
  assign f_arrdiv32_mux2to1237_xor0 = f_arrdiv32_mux2to1237_and0 ^ f_arrdiv32_mux2to1237_and1;
  assign f_arrdiv32_mux2to1238_and0 = f_arrdiv32_mux2to1206_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1238_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1238_and1 = f_arrdiv32_fs245_xor1 & f_arrdiv32_mux2to1238_not0;
  assign f_arrdiv32_mux2to1238_xor0 = f_arrdiv32_mux2to1238_and0 ^ f_arrdiv32_mux2to1238_and1;
  assign f_arrdiv32_mux2to1239_and0 = f_arrdiv32_mux2to1207_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1239_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1239_and1 = f_arrdiv32_fs246_xor1 & f_arrdiv32_mux2to1239_not0;
  assign f_arrdiv32_mux2to1239_xor0 = f_arrdiv32_mux2to1239_and0 ^ f_arrdiv32_mux2to1239_and1;
  assign f_arrdiv32_mux2to1240_and0 = f_arrdiv32_mux2to1208_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1240_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1240_and1 = f_arrdiv32_fs247_xor1 & f_arrdiv32_mux2to1240_not0;
  assign f_arrdiv32_mux2to1240_xor0 = f_arrdiv32_mux2to1240_and0 ^ f_arrdiv32_mux2to1240_and1;
  assign f_arrdiv32_mux2to1241_and0 = f_arrdiv32_mux2to1209_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1241_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1241_and1 = f_arrdiv32_fs248_xor1 & f_arrdiv32_mux2to1241_not0;
  assign f_arrdiv32_mux2to1241_xor0 = f_arrdiv32_mux2to1241_and0 ^ f_arrdiv32_mux2to1241_and1;
  assign f_arrdiv32_mux2to1242_and0 = f_arrdiv32_mux2to1210_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1242_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1242_and1 = f_arrdiv32_fs249_xor1 & f_arrdiv32_mux2to1242_not0;
  assign f_arrdiv32_mux2to1242_xor0 = f_arrdiv32_mux2to1242_and0 ^ f_arrdiv32_mux2to1242_and1;
  assign f_arrdiv32_mux2to1243_and0 = f_arrdiv32_mux2to1211_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1243_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1243_and1 = f_arrdiv32_fs250_xor1 & f_arrdiv32_mux2to1243_not0;
  assign f_arrdiv32_mux2to1243_xor0 = f_arrdiv32_mux2to1243_and0 ^ f_arrdiv32_mux2to1243_and1;
  assign f_arrdiv32_mux2to1244_and0 = f_arrdiv32_mux2to1212_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1244_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1244_and1 = f_arrdiv32_fs251_xor1 & f_arrdiv32_mux2to1244_not0;
  assign f_arrdiv32_mux2to1244_xor0 = f_arrdiv32_mux2to1244_and0 ^ f_arrdiv32_mux2to1244_and1;
  assign f_arrdiv32_mux2to1245_and0 = f_arrdiv32_mux2to1213_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1245_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1245_and1 = f_arrdiv32_fs252_xor1 & f_arrdiv32_mux2to1245_not0;
  assign f_arrdiv32_mux2to1245_xor0 = f_arrdiv32_mux2to1245_and0 ^ f_arrdiv32_mux2to1245_and1;
  assign f_arrdiv32_mux2to1246_and0 = f_arrdiv32_mux2to1214_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1246_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1246_and1 = f_arrdiv32_fs253_xor1 & f_arrdiv32_mux2to1246_not0;
  assign f_arrdiv32_mux2to1246_xor0 = f_arrdiv32_mux2to1246_and0 ^ f_arrdiv32_mux2to1246_and1;
  assign f_arrdiv32_mux2to1247_and0 = f_arrdiv32_mux2to1215_xor0 & f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1247_not0 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_mux2to1247_and1 = f_arrdiv32_fs254_xor1 & f_arrdiv32_mux2to1247_not0;
  assign f_arrdiv32_mux2to1247_xor0 = f_arrdiv32_mux2to1247_and0 ^ f_arrdiv32_mux2to1247_and1;
  assign f_arrdiv32_not7 = ~f_arrdiv32_fs255_or0;
  assign f_arrdiv32_fs256_xor0 = a[23] ^ b[0];
  assign f_arrdiv32_fs256_not0 = ~a[23];
  assign f_arrdiv32_fs256_and0 = f_arrdiv32_fs256_not0 & b[0];
  assign f_arrdiv32_fs256_not1 = ~f_arrdiv32_fs256_xor0;
  assign f_arrdiv32_fs257_xor0 = f_arrdiv32_mux2to1217_xor0 ^ b[1];
  assign f_arrdiv32_fs257_not0 = ~f_arrdiv32_mux2to1217_xor0;
  assign f_arrdiv32_fs257_and0 = f_arrdiv32_fs257_not0 & b[1];
  assign f_arrdiv32_fs257_xor1 = f_arrdiv32_fs256_and0 ^ f_arrdiv32_fs257_xor0;
  assign f_arrdiv32_fs257_not1 = ~f_arrdiv32_fs257_xor0;
  assign f_arrdiv32_fs257_and1 = f_arrdiv32_fs257_not1 & f_arrdiv32_fs256_and0;
  assign f_arrdiv32_fs257_or0 = f_arrdiv32_fs257_and1 | f_arrdiv32_fs257_and0;
  assign f_arrdiv32_fs258_xor0 = f_arrdiv32_mux2to1218_xor0 ^ b[2];
  assign f_arrdiv32_fs258_not0 = ~f_arrdiv32_mux2to1218_xor0;
  assign f_arrdiv32_fs258_and0 = f_arrdiv32_fs258_not0 & b[2];
  assign f_arrdiv32_fs258_xor1 = f_arrdiv32_fs257_or0 ^ f_arrdiv32_fs258_xor0;
  assign f_arrdiv32_fs258_not1 = ~f_arrdiv32_fs258_xor0;
  assign f_arrdiv32_fs258_and1 = f_arrdiv32_fs258_not1 & f_arrdiv32_fs257_or0;
  assign f_arrdiv32_fs258_or0 = f_arrdiv32_fs258_and1 | f_arrdiv32_fs258_and0;
  assign f_arrdiv32_fs259_xor0 = f_arrdiv32_mux2to1219_xor0 ^ b[3];
  assign f_arrdiv32_fs259_not0 = ~f_arrdiv32_mux2to1219_xor0;
  assign f_arrdiv32_fs259_and0 = f_arrdiv32_fs259_not0 & b[3];
  assign f_arrdiv32_fs259_xor1 = f_arrdiv32_fs258_or0 ^ f_arrdiv32_fs259_xor0;
  assign f_arrdiv32_fs259_not1 = ~f_arrdiv32_fs259_xor0;
  assign f_arrdiv32_fs259_and1 = f_arrdiv32_fs259_not1 & f_arrdiv32_fs258_or0;
  assign f_arrdiv32_fs259_or0 = f_arrdiv32_fs259_and1 | f_arrdiv32_fs259_and0;
  assign f_arrdiv32_fs260_xor0 = f_arrdiv32_mux2to1220_xor0 ^ b[4];
  assign f_arrdiv32_fs260_not0 = ~f_arrdiv32_mux2to1220_xor0;
  assign f_arrdiv32_fs260_and0 = f_arrdiv32_fs260_not0 & b[4];
  assign f_arrdiv32_fs260_xor1 = f_arrdiv32_fs259_or0 ^ f_arrdiv32_fs260_xor0;
  assign f_arrdiv32_fs260_not1 = ~f_arrdiv32_fs260_xor0;
  assign f_arrdiv32_fs260_and1 = f_arrdiv32_fs260_not1 & f_arrdiv32_fs259_or0;
  assign f_arrdiv32_fs260_or0 = f_arrdiv32_fs260_and1 | f_arrdiv32_fs260_and0;
  assign f_arrdiv32_fs261_xor0 = f_arrdiv32_mux2to1221_xor0 ^ b[5];
  assign f_arrdiv32_fs261_not0 = ~f_arrdiv32_mux2to1221_xor0;
  assign f_arrdiv32_fs261_and0 = f_arrdiv32_fs261_not0 & b[5];
  assign f_arrdiv32_fs261_xor1 = f_arrdiv32_fs260_or0 ^ f_arrdiv32_fs261_xor0;
  assign f_arrdiv32_fs261_not1 = ~f_arrdiv32_fs261_xor0;
  assign f_arrdiv32_fs261_and1 = f_arrdiv32_fs261_not1 & f_arrdiv32_fs260_or0;
  assign f_arrdiv32_fs261_or0 = f_arrdiv32_fs261_and1 | f_arrdiv32_fs261_and0;
  assign f_arrdiv32_fs262_xor0 = f_arrdiv32_mux2to1222_xor0 ^ b[6];
  assign f_arrdiv32_fs262_not0 = ~f_arrdiv32_mux2to1222_xor0;
  assign f_arrdiv32_fs262_and0 = f_arrdiv32_fs262_not0 & b[6];
  assign f_arrdiv32_fs262_xor1 = f_arrdiv32_fs261_or0 ^ f_arrdiv32_fs262_xor0;
  assign f_arrdiv32_fs262_not1 = ~f_arrdiv32_fs262_xor0;
  assign f_arrdiv32_fs262_and1 = f_arrdiv32_fs262_not1 & f_arrdiv32_fs261_or0;
  assign f_arrdiv32_fs262_or0 = f_arrdiv32_fs262_and1 | f_arrdiv32_fs262_and0;
  assign f_arrdiv32_fs263_xor0 = f_arrdiv32_mux2to1223_xor0 ^ b[7];
  assign f_arrdiv32_fs263_not0 = ~f_arrdiv32_mux2to1223_xor0;
  assign f_arrdiv32_fs263_and0 = f_arrdiv32_fs263_not0 & b[7];
  assign f_arrdiv32_fs263_xor1 = f_arrdiv32_fs262_or0 ^ f_arrdiv32_fs263_xor0;
  assign f_arrdiv32_fs263_not1 = ~f_arrdiv32_fs263_xor0;
  assign f_arrdiv32_fs263_and1 = f_arrdiv32_fs263_not1 & f_arrdiv32_fs262_or0;
  assign f_arrdiv32_fs263_or0 = f_arrdiv32_fs263_and1 | f_arrdiv32_fs263_and0;
  assign f_arrdiv32_fs264_xor0 = f_arrdiv32_mux2to1224_xor0 ^ b[8];
  assign f_arrdiv32_fs264_not0 = ~f_arrdiv32_mux2to1224_xor0;
  assign f_arrdiv32_fs264_and0 = f_arrdiv32_fs264_not0 & b[8];
  assign f_arrdiv32_fs264_xor1 = f_arrdiv32_fs263_or0 ^ f_arrdiv32_fs264_xor0;
  assign f_arrdiv32_fs264_not1 = ~f_arrdiv32_fs264_xor0;
  assign f_arrdiv32_fs264_and1 = f_arrdiv32_fs264_not1 & f_arrdiv32_fs263_or0;
  assign f_arrdiv32_fs264_or0 = f_arrdiv32_fs264_and1 | f_arrdiv32_fs264_and0;
  assign f_arrdiv32_fs265_xor0 = f_arrdiv32_mux2to1225_xor0 ^ b[9];
  assign f_arrdiv32_fs265_not0 = ~f_arrdiv32_mux2to1225_xor0;
  assign f_arrdiv32_fs265_and0 = f_arrdiv32_fs265_not0 & b[9];
  assign f_arrdiv32_fs265_xor1 = f_arrdiv32_fs264_or0 ^ f_arrdiv32_fs265_xor0;
  assign f_arrdiv32_fs265_not1 = ~f_arrdiv32_fs265_xor0;
  assign f_arrdiv32_fs265_and1 = f_arrdiv32_fs265_not1 & f_arrdiv32_fs264_or0;
  assign f_arrdiv32_fs265_or0 = f_arrdiv32_fs265_and1 | f_arrdiv32_fs265_and0;
  assign f_arrdiv32_fs266_xor0 = f_arrdiv32_mux2to1226_xor0 ^ b[10];
  assign f_arrdiv32_fs266_not0 = ~f_arrdiv32_mux2to1226_xor0;
  assign f_arrdiv32_fs266_and0 = f_arrdiv32_fs266_not0 & b[10];
  assign f_arrdiv32_fs266_xor1 = f_arrdiv32_fs265_or0 ^ f_arrdiv32_fs266_xor0;
  assign f_arrdiv32_fs266_not1 = ~f_arrdiv32_fs266_xor0;
  assign f_arrdiv32_fs266_and1 = f_arrdiv32_fs266_not1 & f_arrdiv32_fs265_or0;
  assign f_arrdiv32_fs266_or0 = f_arrdiv32_fs266_and1 | f_arrdiv32_fs266_and0;
  assign f_arrdiv32_fs267_xor0 = f_arrdiv32_mux2to1227_xor0 ^ b[11];
  assign f_arrdiv32_fs267_not0 = ~f_arrdiv32_mux2to1227_xor0;
  assign f_arrdiv32_fs267_and0 = f_arrdiv32_fs267_not0 & b[11];
  assign f_arrdiv32_fs267_xor1 = f_arrdiv32_fs266_or0 ^ f_arrdiv32_fs267_xor0;
  assign f_arrdiv32_fs267_not1 = ~f_arrdiv32_fs267_xor0;
  assign f_arrdiv32_fs267_and1 = f_arrdiv32_fs267_not1 & f_arrdiv32_fs266_or0;
  assign f_arrdiv32_fs267_or0 = f_arrdiv32_fs267_and1 | f_arrdiv32_fs267_and0;
  assign f_arrdiv32_fs268_xor0 = f_arrdiv32_mux2to1228_xor0 ^ b[12];
  assign f_arrdiv32_fs268_not0 = ~f_arrdiv32_mux2to1228_xor0;
  assign f_arrdiv32_fs268_and0 = f_arrdiv32_fs268_not0 & b[12];
  assign f_arrdiv32_fs268_xor1 = f_arrdiv32_fs267_or0 ^ f_arrdiv32_fs268_xor0;
  assign f_arrdiv32_fs268_not1 = ~f_arrdiv32_fs268_xor0;
  assign f_arrdiv32_fs268_and1 = f_arrdiv32_fs268_not1 & f_arrdiv32_fs267_or0;
  assign f_arrdiv32_fs268_or0 = f_arrdiv32_fs268_and1 | f_arrdiv32_fs268_and0;
  assign f_arrdiv32_fs269_xor0 = f_arrdiv32_mux2to1229_xor0 ^ b[13];
  assign f_arrdiv32_fs269_not0 = ~f_arrdiv32_mux2to1229_xor0;
  assign f_arrdiv32_fs269_and0 = f_arrdiv32_fs269_not0 & b[13];
  assign f_arrdiv32_fs269_xor1 = f_arrdiv32_fs268_or0 ^ f_arrdiv32_fs269_xor0;
  assign f_arrdiv32_fs269_not1 = ~f_arrdiv32_fs269_xor0;
  assign f_arrdiv32_fs269_and1 = f_arrdiv32_fs269_not1 & f_arrdiv32_fs268_or0;
  assign f_arrdiv32_fs269_or0 = f_arrdiv32_fs269_and1 | f_arrdiv32_fs269_and0;
  assign f_arrdiv32_fs270_xor0 = f_arrdiv32_mux2to1230_xor0 ^ b[14];
  assign f_arrdiv32_fs270_not0 = ~f_arrdiv32_mux2to1230_xor0;
  assign f_arrdiv32_fs270_and0 = f_arrdiv32_fs270_not0 & b[14];
  assign f_arrdiv32_fs270_xor1 = f_arrdiv32_fs269_or0 ^ f_arrdiv32_fs270_xor0;
  assign f_arrdiv32_fs270_not1 = ~f_arrdiv32_fs270_xor0;
  assign f_arrdiv32_fs270_and1 = f_arrdiv32_fs270_not1 & f_arrdiv32_fs269_or0;
  assign f_arrdiv32_fs270_or0 = f_arrdiv32_fs270_and1 | f_arrdiv32_fs270_and0;
  assign f_arrdiv32_fs271_xor0 = f_arrdiv32_mux2to1231_xor0 ^ b[15];
  assign f_arrdiv32_fs271_not0 = ~f_arrdiv32_mux2to1231_xor0;
  assign f_arrdiv32_fs271_and0 = f_arrdiv32_fs271_not0 & b[15];
  assign f_arrdiv32_fs271_xor1 = f_arrdiv32_fs270_or0 ^ f_arrdiv32_fs271_xor0;
  assign f_arrdiv32_fs271_not1 = ~f_arrdiv32_fs271_xor0;
  assign f_arrdiv32_fs271_and1 = f_arrdiv32_fs271_not1 & f_arrdiv32_fs270_or0;
  assign f_arrdiv32_fs271_or0 = f_arrdiv32_fs271_and1 | f_arrdiv32_fs271_and0;
  assign f_arrdiv32_fs272_xor0 = f_arrdiv32_mux2to1232_xor0 ^ b[16];
  assign f_arrdiv32_fs272_not0 = ~f_arrdiv32_mux2to1232_xor0;
  assign f_arrdiv32_fs272_and0 = f_arrdiv32_fs272_not0 & b[16];
  assign f_arrdiv32_fs272_xor1 = f_arrdiv32_fs271_or0 ^ f_arrdiv32_fs272_xor0;
  assign f_arrdiv32_fs272_not1 = ~f_arrdiv32_fs272_xor0;
  assign f_arrdiv32_fs272_and1 = f_arrdiv32_fs272_not1 & f_arrdiv32_fs271_or0;
  assign f_arrdiv32_fs272_or0 = f_arrdiv32_fs272_and1 | f_arrdiv32_fs272_and0;
  assign f_arrdiv32_fs273_xor0 = f_arrdiv32_mux2to1233_xor0 ^ b[17];
  assign f_arrdiv32_fs273_not0 = ~f_arrdiv32_mux2to1233_xor0;
  assign f_arrdiv32_fs273_and0 = f_arrdiv32_fs273_not0 & b[17];
  assign f_arrdiv32_fs273_xor1 = f_arrdiv32_fs272_or0 ^ f_arrdiv32_fs273_xor0;
  assign f_arrdiv32_fs273_not1 = ~f_arrdiv32_fs273_xor0;
  assign f_arrdiv32_fs273_and1 = f_arrdiv32_fs273_not1 & f_arrdiv32_fs272_or0;
  assign f_arrdiv32_fs273_or0 = f_arrdiv32_fs273_and1 | f_arrdiv32_fs273_and0;
  assign f_arrdiv32_fs274_xor0 = f_arrdiv32_mux2to1234_xor0 ^ b[18];
  assign f_arrdiv32_fs274_not0 = ~f_arrdiv32_mux2to1234_xor0;
  assign f_arrdiv32_fs274_and0 = f_arrdiv32_fs274_not0 & b[18];
  assign f_arrdiv32_fs274_xor1 = f_arrdiv32_fs273_or0 ^ f_arrdiv32_fs274_xor0;
  assign f_arrdiv32_fs274_not1 = ~f_arrdiv32_fs274_xor0;
  assign f_arrdiv32_fs274_and1 = f_arrdiv32_fs274_not1 & f_arrdiv32_fs273_or0;
  assign f_arrdiv32_fs274_or0 = f_arrdiv32_fs274_and1 | f_arrdiv32_fs274_and0;
  assign f_arrdiv32_fs275_xor0 = f_arrdiv32_mux2to1235_xor0 ^ b[19];
  assign f_arrdiv32_fs275_not0 = ~f_arrdiv32_mux2to1235_xor0;
  assign f_arrdiv32_fs275_and0 = f_arrdiv32_fs275_not0 & b[19];
  assign f_arrdiv32_fs275_xor1 = f_arrdiv32_fs274_or0 ^ f_arrdiv32_fs275_xor0;
  assign f_arrdiv32_fs275_not1 = ~f_arrdiv32_fs275_xor0;
  assign f_arrdiv32_fs275_and1 = f_arrdiv32_fs275_not1 & f_arrdiv32_fs274_or0;
  assign f_arrdiv32_fs275_or0 = f_arrdiv32_fs275_and1 | f_arrdiv32_fs275_and0;
  assign f_arrdiv32_fs276_xor0 = f_arrdiv32_mux2to1236_xor0 ^ b[20];
  assign f_arrdiv32_fs276_not0 = ~f_arrdiv32_mux2to1236_xor0;
  assign f_arrdiv32_fs276_and0 = f_arrdiv32_fs276_not0 & b[20];
  assign f_arrdiv32_fs276_xor1 = f_arrdiv32_fs275_or0 ^ f_arrdiv32_fs276_xor0;
  assign f_arrdiv32_fs276_not1 = ~f_arrdiv32_fs276_xor0;
  assign f_arrdiv32_fs276_and1 = f_arrdiv32_fs276_not1 & f_arrdiv32_fs275_or0;
  assign f_arrdiv32_fs276_or0 = f_arrdiv32_fs276_and1 | f_arrdiv32_fs276_and0;
  assign f_arrdiv32_fs277_xor0 = f_arrdiv32_mux2to1237_xor0 ^ b[21];
  assign f_arrdiv32_fs277_not0 = ~f_arrdiv32_mux2to1237_xor0;
  assign f_arrdiv32_fs277_and0 = f_arrdiv32_fs277_not0 & b[21];
  assign f_arrdiv32_fs277_xor1 = f_arrdiv32_fs276_or0 ^ f_arrdiv32_fs277_xor0;
  assign f_arrdiv32_fs277_not1 = ~f_arrdiv32_fs277_xor0;
  assign f_arrdiv32_fs277_and1 = f_arrdiv32_fs277_not1 & f_arrdiv32_fs276_or0;
  assign f_arrdiv32_fs277_or0 = f_arrdiv32_fs277_and1 | f_arrdiv32_fs277_and0;
  assign f_arrdiv32_fs278_xor0 = f_arrdiv32_mux2to1238_xor0 ^ b[22];
  assign f_arrdiv32_fs278_not0 = ~f_arrdiv32_mux2to1238_xor0;
  assign f_arrdiv32_fs278_and0 = f_arrdiv32_fs278_not0 & b[22];
  assign f_arrdiv32_fs278_xor1 = f_arrdiv32_fs277_or0 ^ f_arrdiv32_fs278_xor0;
  assign f_arrdiv32_fs278_not1 = ~f_arrdiv32_fs278_xor0;
  assign f_arrdiv32_fs278_and1 = f_arrdiv32_fs278_not1 & f_arrdiv32_fs277_or0;
  assign f_arrdiv32_fs278_or0 = f_arrdiv32_fs278_and1 | f_arrdiv32_fs278_and0;
  assign f_arrdiv32_fs279_xor0 = f_arrdiv32_mux2to1239_xor0 ^ b[23];
  assign f_arrdiv32_fs279_not0 = ~f_arrdiv32_mux2to1239_xor0;
  assign f_arrdiv32_fs279_and0 = f_arrdiv32_fs279_not0 & b[23];
  assign f_arrdiv32_fs279_xor1 = f_arrdiv32_fs278_or0 ^ f_arrdiv32_fs279_xor0;
  assign f_arrdiv32_fs279_not1 = ~f_arrdiv32_fs279_xor0;
  assign f_arrdiv32_fs279_and1 = f_arrdiv32_fs279_not1 & f_arrdiv32_fs278_or0;
  assign f_arrdiv32_fs279_or0 = f_arrdiv32_fs279_and1 | f_arrdiv32_fs279_and0;
  assign f_arrdiv32_fs280_xor0 = f_arrdiv32_mux2to1240_xor0 ^ b[24];
  assign f_arrdiv32_fs280_not0 = ~f_arrdiv32_mux2to1240_xor0;
  assign f_arrdiv32_fs280_and0 = f_arrdiv32_fs280_not0 & b[24];
  assign f_arrdiv32_fs280_xor1 = f_arrdiv32_fs279_or0 ^ f_arrdiv32_fs280_xor0;
  assign f_arrdiv32_fs280_not1 = ~f_arrdiv32_fs280_xor0;
  assign f_arrdiv32_fs280_and1 = f_arrdiv32_fs280_not1 & f_arrdiv32_fs279_or0;
  assign f_arrdiv32_fs280_or0 = f_arrdiv32_fs280_and1 | f_arrdiv32_fs280_and0;
  assign f_arrdiv32_fs281_xor0 = f_arrdiv32_mux2to1241_xor0 ^ b[25];
  assign f_arrdiv32_fs281_not0 = ~f_arrdiv32_mux2to1241_xor0;
  assign f_arrdiv32_fs281_and0 = f_arrdiv32_fs281_not0 & b[25];
  assign f_arrdiv32_fs281_xor1 = f_arrdiv32_fs280_or0 ^ f_arrdiv32_fs281_xor0;
  assign f_arrdiv32_fs281_not1 = ~f_arrdiv32_fs281_xor0;
  assign f_arrdiv32_fs281_and1 = f_arrdiv32_fs281_not1 & f_arrdiv32_fs280_or0;
  assign f_arrdiv32_fs281_or0 = f_arrdiv32_fs281_and1 | f_arrdiv32_fs281_and0;
  assign f_arrdiv32_fs282_xor0 = f_arrdiv32_mux2to1242_xor0 ^ b[26];
  assign f_arrdiv32_fs282_not0 = ~f_arrdiv32_mux2to1242_xor0;
  assign f_arrdiv32_fs282_and0 = f_arrdiv32_fs282_not0 & b[26];
  assign f_arrdiv32_fs282_xor1 = f_arrdiv32_fs281_or0 ^ f_arrdiv32_fs282_xor0;
  assign f_arrdiv32_fs282_not1 = ~f_arrdiv32_fs282_xor0;
  assign f_arrdiv32_fs282_and1 = f_arrdiv32_fs282_not1 & f_arrdiv32_fs281_or0;
  assign f_arrdiv32_fs282_or0 = f_arrdiv32_fs282_and1 | f_arrdiv32_fs282_and0;
  assign f_arrdiv32_fs283_xor0 = f_arrdiv32_mux2to1243_xor0 ^ b[27];
  assign f_arrdiv32_fs283_not0 = ~f_arrdiv32_mux2to1243_xor0;
  assign f_arrdiv32_fs283_and0 = f_arrdiv32_fs283_not0 & b[27];
  assign f_arrdiv32_fs283_xor1 = f_arrdiv32_fs282_or0 ^ f_arrdiv32_fs283_xor0;
  assign f_arrdiv32_fs283_not1 = ~f_arrdiv32_fs283_xor0;
  assign f_arrdiv32_fs283_and1 = f_arrdiv32_fs283_not1 & f_arrdiv32_fs282_or0;
  assign f_arrdiv32_fs283_or0 = f_arrdiv32_fs283_and1 | f_arrdiv32_fs283_and0;
  assign f_arrdiv32_fs284_xor0 = f_arrdiv32_mux2to1244_xor0 ^ b[28];
  assign f_arrdiv32_fs284_not0 = ~f_arrdiv32_mux2to1244_xor0;
  assign f_arrdiv32_fs284_and0 = f_arrdiv32_fs284_not0 & b[28];
  assign f_arrdiv32_fs284_xor1 = f_arrdiv32_fs283_or0 ^ f_arrdiv32_fs284_xor0;
  assign f_arrdiv32_fs284_not1 = ~f_arrdiv32_fs284_xor0;
  assign f_arrdiv32_fs284_and1 = f_arrdiv32_fs284_not1 & f_arrdiv32_fs283_or0;
  assign f_arrdiv32_fs284_or0 = f_arrdiv32_fs284_and1 | f_arrdiv32_fs284_and0;
  assign f_arrdiv32_fs285_xor0 = f_arrdiv32_mux2to1245_xor0 ^ b[29];
  assign f_arrdiv32_fs285_not0 = ~f_arrdiv32_mux2to1245_xor0;
  assign f_arrdiv32_fs285_and0 = f_arrdiv32_fs285_not0 & b[29];
  assign f_arrdiv32_fs285_xor1 = f_arrdiv32_fs284_or0 ^ f_arrdiv32_fs285_xor0;
  assign f_arrdiv32_fs285_not1 = ~f_arrdiv32_fs285_xor0;
  assign f_arrdiv32_fs285_and1 = f_arrdiv32_fs285_not1 & f_arrdiv32_fs284_or0;
  assign f_arrdiv32_fs285_or0 = f_arrdiv32_fs285_and1 | f_arrdiv32_fs285_and0;
  assign f_arrdiv32_fs286_xor0 = f_arrdiv32_mux2to1246_xor0 ^ b[30];
  assign f_arrdiv32_fs286_not0 = ~f_arrdiv32_mux2to1246_xor0;
  assign f_arrdiv32_fs286_and0 = f_arrdiv32_fs286_not0 & b[30];
  assign f_arrdiv32_fs286_xor1 = f_arrdiv32_fs285_or0 ^ f_arrdiv32_fs286_xor0;
  assign f_arrdiv32_fs286_not1 = ~f_arrdiv32_fs286_xor0;
  assign f_arrdiv32_fs286_and1 = f_arrdiv32_fs286_not1 & f_arrdiv32_fs285_or0;
  assign f_arrdiv32_fs286_or0 = f_arrdiv32_fs286_and1 | f_arrdiv32_fs286_and0;
  assign f_arrdiv32_fs287_xor0 = f_arrdiv32_mux2to1247_xor0 ^ b[31];
  assign f_arrdiv32_fs287_not0 = ~f_arrdiv32_mux2to1247_xor0;
  assign f_arrdiv32_fs287_and0 = f_arrdiv32_fs287_not0 & b[31];
  assign f_arrdiv32_fs287_xor1 = f_arrdiv32_fs286_or0 ^ f_arrdiv32_fs287_xor0;
  assign f_arrdiv32_fs287_not1 = ~f_arrdiv32_fs287_xor0;
  assign f_arrdiv32_fs287_and1 = f_arrdiv32_fs287_not1 & f_arrdiv32_fs286_or0;
  assign f_arrdiv32_fs287_or0 = f_arrdiv32_fs287_and1 | f_arrdiv32_fs287_and0;
  assign f_arrdiv32_mux2to1248_and0 = a[23] & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1248_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1248_and1 = f_arrdiv32_fs256_xor0 & f_arrdiv32_mux2to1248_not0;
  assign f_arrdiv32_mux2to1248_xor0 = f_arrdiv32_mux2to1248_and0 ^ f_arrdiv32_mux2to1248_and1;
  assign f_arrdiv32_mux2to1249_and0 = f_arrdiv32_mux2to1217_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1249_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1249_and1 = f_arrdiv32_fs257_xor1 & f_arrdiv32_mux2to1249_not0;
  assign f_arrdiv32_mux2to1249_xor0 = f_arrdiv32_mux2to1249_and0 ^ f_arrdiv32_mux2to1249_and1;
  assign f_arrdiv32_mux2to1250_and0 = f_arrdiv32_mux2to1218_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1250_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1250_and1 = f_arrdiv32_fs258_xor1 & f_arrdiv32_mux2to1250_not0;
  assign f_arrdiv32_mux2to1250_xor0 = f_arrdiv32_mux2to1250_and0 ^ f_arrdiv32_mux2to1250_and1;
  assign f_arrdiv32_mux2to1251_and0 = f_arrdiv32_mux2to1219_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1251_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1251_and1 = f_arrdiv32_fs259_xor1 & f_arrdiv32_mux2to1251_not0;
  assign f_arrdiv32_mux2to1251_xor0 = f_arrdiv32_mux2to1251_and0 ^ f_arrdiv32_mux2to1251_and1;
  assign f_arrdiv32_mux2to1252_and0 = f_arrdiv32_mux2to1220_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1252_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1252_and1 = f_arrdiv32_fs260_xor1 & f_arrdiv32_mux2to1252_not0;
  assign f_arrdiv32_mux2to1252_xor0 = f_arrdiv32_mux2to1252_and0 ^ f_arrdiv32_mux2to1252_and1;
  assign f_arrdiv32_mux2to1253_and0 = f_arrdiv32_mux2to1221_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1253_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1253_and1 = f_arrdiv32_fs261_xor1 & f_arrdiv32_mux2to1253_not0;
  assign f_arrdiv32_mux2to1253_xor0 = f_arrdiv32_mux2to1253_and0 ^ f_arrdiv32_mux2to1253_and1;
  assign f_arrdiv32_mux2to1254_and0 = f_arrdiv32_mux2to1222_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1254_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1254_and1 = f_arrdiv32_fs262_xor1 & f_arrdiv32_mux2to1254_not0;
  assign f_arrdiv32_mux2to1254_xor0 = f_arrdiv32_mux2to1254_and0 ^ f_arrdiv32_mux2to1254_and1;
  assign f_arrdiv32_mux2to1255_and0 = f_arrdiv32_mux2to1223_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1255_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1255_and1 = f_arrdiv32_fs263_xor1 & f_arrdiv32_mux2to1255_not0;
  assign f_arrdiv32_mux2to1255_xor0 = f_arrdiv32_mux2to1255_and0 ^ f_arrdiv32_mux2to1255_and1;
  assign f_arrdiv32_mux2to1256_and0 = f_arrdiv32_mux2to1224_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1256_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1256_and1 = f_arrdiv32_fs264_xor1 & f_arrdiv32_mux2to1256_not0;
  assign f_arrdiv32_mux2to1256_xor0 = f_arrdiv32_mux2to1256_and0 ^ f_arrdiv32_mux2to1256_and1;
  assign f_arrdiv32_mux2to1257_and0 = f_arrdiv32_mux2to1225_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1257_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1257_and1 = f_arrdiv32_fs265_xor1 & f_arrdiv32_mux2to1257_not0;
  assign f_arrdiv32_mux2to1257_xor0 = f_arrdiv32_mux2to1257_and0 ^ f_arrdiv32_mux2to1257_and1;
  assign f_arrdiv32_mux2to1258_and0 = f_arrdiv32_mux2to1226_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1258_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1258_and1 = f_arrdiv32_fs266_xor1 & f_arrdiv32_mux2to1258_not0;
  assign f_arrdiv32_mux2to1258_xor0 = f_arrdiv32_mux2to1258_and0 ^ f_arrdiv32_mux2to1258_and1;
  assign f_arrdiv32_mux2to1259_and0 = f_arrdiv32_mux2to1227_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1259_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1259_and1 = f_arrdiv32_fs267_xor1 & f_arrdiv32_mux2to1259_not0;
  assign f_arrdiv32_mux2to1259_xor0 = f_arrdiv32_mux2to1259_and0 ^ f_arrdiv32_mux2to1259_and1;
  assign f_arrdiv32_mux2to1260_and0 = f_arrdiv32_mux2to1228_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1260_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1260_and1 = f_arrdiv32_fs268_xor1 & f_arrdiv32_mux2to1260_not0;
  assign f_arrdiv32_mux2to1260_xor0 = f_arrdiv32_mux2to1260_and0 ^ f_arrdiv32_mux2to1260_and1;
  assign f_arrdiv32_mux2to1261_and0 = f_arrdiv32_mux2to1229_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1261_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1261_and1 = f_arrdiv32_fs269_xor1 & f_arrdiv32_mux2to1261_not0;
  assign f_arrdiv32_mux2to1261_xor0 = f_arrdiv32_mux2to1261_and0 ^ f_arrdiv32_mux2to1261_and1;
  assign f_arrdiv32_mux2to1262_and0 = f_arrdiv32_mux2to1230_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1262_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1262_and1 = f_arrdiv32_fs270_xor1 & f_arrdiv32_mux2to1262_not0;
  assign f_arrdiv32_mux2to1262_xor0 = f_arrdiv32_mux2to1262_and0 ^ f_arrdiv32_mux2to1262_and1;
  assign f_arrdiv32_mux2to1263_and0 = f_arrdiv32_mux2to1231_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1263_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1263_and1 = f_arrdiv32_fs271_xor1 & f_arrdiv32_mux2to1263_not0;
  assign f_arrdiv32_mux2to1263_xor0 = f_arrdiv32_mux2to1263_and0 ^ f_arrdiv32_mux2to1263_and1;
  assign f_arrdiv32_mux2to1264_and0 = f_arrdiv32_mux2to1232_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1264_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1264_and1 = f_arrdiv32_fs272_xor1 & f_arrdiv32_mux2to1264_not0;
  assign f_arrdiv32_mux2to1264_xor0 = f_arrdiv32_mux2to1264_and0 ^ f_arrdiv32_mux2to1264_and1;
  assign f_arrdiv32_mux2to1265_and0 = f_arrdiv32_mux2to1233_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1265_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1265_and1 = f_arrdiv32_fs273_xor1 & f_arrdiv32_mux2to1265_not0;
  assign f_arrdiv32_mux2to1265_xor0 = f_arrdiv32_mux2to1265_and0 ^ f_arrdiv32_mux2to1265_and1;
  assign f_arrdiv32_mux2to1266_and0 = f_arrdiv32_mux2to1234_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1266_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1266_and1 = f_arrdiv32_fs274_xor1 & f_arrdiv32_mux2to1266_not0;
  assign f_arrdiv32_mux2to1266_xor0 = f_arrdiv32_mux2to1266_and0 ^ f_arrdiv32_mux2to1266_and1;
  assign f_arrdiv32_mux2to1267_and0 = f_arrdiv32_mux2to1235_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1267_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1267_and1 = f_arrdiv32_fs275_xor1 & f_arrdiv32_mux2to1267_not0;
  assign f_arrdiv32_mux2to1267_xor0 = f_arrdiv32_mux2to1267_and0 ^ f_arrdiv32_mux2to1267_and1;
  assign f_arrdiv32_mux2to1268_and0 = f_arrdiv32_mux2to1236_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1268_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1268_and1 = f_arrdiv32_fs276_xor1 & f_arrdiv32_mux2to1268_not0;
  assign f_arrdiv32_mux2to1268_xor0 = f_arrdiv32_mux2to1268_and0 ^ f_arrdiv32_mux2to1268_and1;
  assign f_arrdiv32_mux2to1269_and0 = f_arrdiv32_mux2to1237_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1269_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1269_and1 = f_arrdiv32_fs277_xor1 & f_arrdiv32_mux2to1269_not0;
  assign f_arrdiv32_mux2to1269_xor0 = f_arrdiv32_mux2to1269_and0 ^ f_arrdiv32_mux2to1269_and1;
  assign f_arrdiv32_mux2to1270_and0 = f_arrdiv32_mux2to1238_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1270_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1270_and1 = f_arrdiv32_fs278_xor1 & f_arrdiv32_mux2to1270_not0;
  assign f_arrdiv32_mux2to1270_xor0 = f_arrdiv32_mux2to1270_and0 ^ f_arrdiv32_mux2to1270_and1;
  assign f_arrdiv32_mux2to1271_and0 = f_arrdiv32_mux2to1239_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1271_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1271_and1 = f_arrdiv32_fs279_xor1 & f_arrdiv32_mux2to1271_not0;
  assign f_arrdiv32_mux2to1271_xor0 = f_arrdiv32_mux2to1271_and0 ^ f_arrdiv32_mux2to1271_and1;
  assign f_arrdiv32_mux2to1272_and0 = f_arrdiv32_mux2to1240_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1272_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1272_and1 = f_arrdiv32_fs280_xor1 & f_arrdiv32_mux2to1272_not0;
  assign f_arrdiv32_mux2to1272_xor0 = f_arrdiv32_mux2to1272_and0 ^ f_arrdiv32_mux2to1272_and1;
  assign f_arrdiv32_mux2to1273_and0 = f_arrdiv32_mux2to1241_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1273_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1273_and1 = f_arrdiv32_fs281_xor1 & f_arrdiv32_mux2to1273_not0;
  assign f_arrdiv32_mux2to1273_xor0 = f_arrdiv32_mux2to1273_and0 ^ f_arrdiv32_mux2to1273_and1;
  assign f_arrdiv32_mux2to1274_and0 = f_arrdiv32_mux2to1242_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1274_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1274_and1 = f_arrdiv32_fs282_xor1 & f_arrdiv32_mux2to1274_not0;
  assign f_arrdiv32_mux2to1274_xor0 = f_arrdiv32_mux2to1274_and0 ^ f_arrdiv32_mux2to1274_and1;
  assign f_arrdiv32_mux2to1275_and0 = f_arrdiv32_mux2to1243_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1275_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1275_and1 = f_arrdiv32_fs283_xor1 & f_arrdiv32_mux2to1275_not0;
  assign f_arrdiv32_mux2to1275_xor0 = f_arrdiv32_mux2to1275_and0 ^ f_arrdiv32_mux2to1275_and1;
  assign f_arrdiv32_mux2to1276_and0 = f_arrdiv32_mux2to1244_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1276_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1276_and1 = f_arrdiv32_fs284_xor1 & f_arrdiv32_mux2to1276_not0;
  assign f_arrdiv32_mux2to1276_xor0 = f_arrdiv32_mux2to1276_and0 ^ f_arrdiv32_mux2to1276_and1;
  assign f_arrdiv32_mux2to1277_and0 = f_arrdiv32_mux2to1245_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1277_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1277_and1 = f_arrdiv32_fs285_xor1 & f_arrdiv32_mux2to1277_not0;
  assign f_arrdiv32_mux2to1277_xor0 = f_arrdiv32_mux2to1277_and0 ^ f_arrdiv32_mux2to1277_and1;
  assign f_arrdiv32_mux2to1278_and0 = f_arrdiv32_mux2to1246_xor0 & f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1278_not0 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_mux2to1278_and1 = f_arrdiv32_fs286_xor1 & f_arrdiv32_mux2to1278_not0;
  assign f_arrdiv32_mux2to1278_xor0 = f_arrdiv32_mux2to1278_and0 ^ f_arrdiv32_mux2to1278_and1;
  assign f_arrdiv32_not8 = ~f_arrdiv32_fs287_or0;
  assign f_arrdiv32_fs288_xor0 = a[22] ^ b[0];
  assign f_arrdiv32_fs288_not0 = ~a[22];
  assign f_arrdiv32_fs288_and0 = f_arrdiv32_fs288_not0 & b[0];
  assign f_arrdiv32_fs288_not1 = ~f_arrdiv32_fs288_xor0;
  assign f_arrdiv32_fs289_xor0 = f_arrdiv32_mux2to1248_xor0 ^ b[1];
  assign f_arrdiv32_fs289_not0 = ~f_arrdiv32_mux2to1248_xor0;
  assign f_arrdiv32_fs289_and0 = f_arrdiv32_fs289_not0 & b[1];
  assign f_arrdiv32_fs289_xor1 = f_arrdiv32_fs288_and0 ^ f_arrdiv32_fs289_xor0;
  assign f_arrdiv32_fs289_not1 = ~f_arrdiv32_fs289_xor0;
  assign f_arrdiv32_fs289_and1 = f_arrdiv32_fs289_not1 & f_arrdiv32_fs288_and0;
  assign f_arrdiv32_fs289_or0 = f_arrdiv32_fs289_and1 | f_arrdiv32_fs289_and0;
  assign f_arrdiv32_fs290_xor0 = f_arrdiv32_mux2to1249_xor0 ^ b[2];
  assign f_arrdiv32_fs290_not0 = ~f_arrdiv32_mux2to1249_xor0;
  assign f_arrdiv32_fs290_and0 = f_arrdiv32_fs290_not0 & b[2];
  assign f_arrdiv32_fs290_xor1 = f_arrdiv32_fs289_or0 ^ f_arrdiv32_fs290_xor0;
  assign f_arrdiv32_fs290_not1 = ~f_arrdiv32_fs290_xor0;
  assign f_arrdiv32_fs290_and1 = f_arrdiv32_fs290_not1 & f_arrdiv32_fs289_or0;
  assign f_arrdiv32_fs290_or0 = f_arrdiv32_fs290_and1 | f_arrdiv32_fs290_and0;
  assign f_arrdiv32_fs291_xor0 = f_arrdiv32_mux2to1250_xor0 ^ b[3];
  assign f_arrdiv32_fs291_not0 = ~f_arrdiv32_mux2to1250_xor0;
  assign f_arrdiv32_fs291_and0 = f_arrdiv32_fs291_not0 & b[3];
  assign f_arrdiv32_fs291_xor1 = f_arrdiv32_fs290_or0 ^ f_arrdiv32_fs291_xor0;
  assign f_arrdiv32_fs291_not1 = ~f_arrdiv32_fs291_xor0;
  assign f_arrdiv32_fs291_and1 = f_arrdiv32_fs291_not1 & f_arrdiv32_fs290_or0;
  assign f_arrdiv32_fs291_or0 = f_arrdiv32_fs291_and1 | f_arrdiv32_fs291_and0;
  assign f_arrdiv32_fs292_xor0 = f_arrdiv32_mux2to1251_xor0 ^ b[4];
  assign f_arrdiv32_fs292_not0 = ~f_arrdiv32_mux2to1251_xor0;
  assign f_arrdiv32_fs292_and0 = f_arrdiv32_fs292_not0 & b[4];
  assign f_arrdiv32_fs292_xor1 = f_arrdiv32_fs291_or0 ^ f_arrdiv32_fs292_xor0;
  assign f_arrdiv32_fs292_not1 = ~f_arrdiv32_fs292_xor0;
  assign f_arrdiv32_fs292_and1 = f_arrdiv32_fs292_not1 & f_arrdiv32_fs291_or0;
  assign f_arrdiv32_fs292_or0 = f_arrdiv32_fs292_and1 | f_arrdiv32_fs292_and0;
  assign f_arrdiv32_fs293_xor0 = f_arrdiv32_mux2to1252_xor0 ^ b[5];
  assign f_arrdiv32_fs293_not0 = ~f_arrdiv32_mux2to1252_xor0;
  assign f_arrdiv32_fs293_and0 = f_arrdiv32_fs293_not0 & b[5];
  assign f_arrdiv32_fs293_xor1 = f_arrdiv32_fs292_or0 ^ f_arrdiv32_fs293_xor0;
  assign f_arrdiv32_fs293_not1 = ~f_arrdiv32_fs293_xor0;
  assign f_arrdiv32_fs293_and1 = f_arrdiv32_fs293_not1 & f_arrdiv32_fs292_or0;
  assign f_arrdiv32_fs293_or0 = f_arrdiv32_fs293_and1 | f_arrdiv32_fs293_and0;
  assign f_arrdiv32_fs294_xor0 = f_arrdiv32_mux2to1253_xor0 ^ b[6];
  assign f_arrdiv32_fs294_not0 = ~f_arrdiv32_mux2to1253_xor0;
  assign f_arrdiv32_fs294_and0 = f_arrdiv32_fs294_not0 & b[6];
  assign f_arrdiv32_fs294_xor1 = f_arrdiv32_fs293_or0 ^ f_arrdiv32_fs294_xor0;
  assign f_arrdiv32_fs294_not1 = ~f_arrdiv32_fs294_xor0;
  assign f_arrdiv32_fs294_and1 = f_arrdiv32_fs294_not1 & f_arrdiv32_fs293_or0;
  assign f_arrdiv32_fs294_or0 = f_arrdiv32_fs294_and1 | f_arrdiv32_fs294_and0;
  assign f_arrdiv32_fs295_xor0 = f_arrdiv32_mux2to1254_xor0 ^ b[7];
  assign f_arrdiv32_fs295_not0 = ~f_arrdiv32_mux2to1254_xor0;
  assign f_arrdiv32_fs295_and0 = f_arrdiv32_fs295_not0 & b[7];
  assign f_arrdiv32_fs295_xor1 = f_arrdiv32_fs294_or0 ^ f_arrdiv32_fs295_xor0;
  assign f_arrdiv32_fs295_not1 = ~f_arrdiv32_fs295_xor0;
  assign f_arrdiv32_fs295_and1 = f_arrdiv32_fs295_not1 & f_arrdiv32_fs294_or0;
  assign f_arrdiv32_fs295_or0 = f_arrdiv32_fs295_and1 | f_arrdiv32_fs295_and0;
  assign f_arrdiv32_fs296_xor0 = f_arrdiv32_mux2to1255_xor0 ^ b[8];
  assign f_arrdiv32_fs296_not0 = ~f_arrdiv32_mux2to1255_xor0;
  assign f_arrdiv32_fs296_and0 = f_arrdiv32_fs296_not0 & b[8];
  assign f_arrdiv32_fs296_xor1 = f_arrdiv32_fs295_or0 ^ f_arrdiv32_fs296_xor0;
  assign f_arrdiv32_fs296_not1 = ~f_arrdiv32_fs296_xor0;
  assign f_arrdiv32_fs296_and1 = f_arrdiv32_fs296_not1 & f_arrdiv32_fs295_or0;
  assign f_arrdiv32_fs296_or0 = f_arrdiv32_fs296_and1 | f_arrdiv32_fs296_and0;
  assign f_arrdiv32_fs297_xor0 = f_arrdiv32_mux2to1256_xor0 ^ b[9];
  assign f_arrdiv32_fs297_not0 = ~f_arrdiv32_mux2to1256_xor0;
  assign f_arrdiv32_fs297_and0 = f_arrdiv32_fs297_not0 & b[9];
  assign f_arrdiv32_fs297_xor1 = f_arrdiv32_fs296_or0 ^ f_arrdiv32_fs297_xor0;
  assign f_arrdiv32_fs297_not1 = ~f_arrdiv32_fs297_xor0;
  assign f_arrdiv32_fs297_and1 = f_arrdiv32_fs297_not1 & f_arrdiv32_fs296_or0;
  assign f_arrdiv32_fs297_or0 = f_arrdiv32_fs297_and1 | f_arrdiv32_fs297_and0;
  assign f_arrdiv32_fs298_xor0 = f_arrdiv32_mux2to1257_xor0 ^ b[10];
  assign f_arrdiv32_fs298_not0 = ~f_arrdiv32_mux2to1257_xor0;
  assign f_arrdiv32_fs298_and0 = f_arrdiv32_fs298_not0 & b[10];
  assign f_arrdiv32_fs298_xor1 = f_arrdiv32_fs297_or0 ^ f_arrdiv32_fs298_xor0;
  assign f_arrdiv32_fs298_not1 = ~f_arrdiv32_fs298_xor0;
  assign f_arrdiv32_fs298_and1 = f_arrdiv32_fs298_not1 & f_arrdiv32_fs297_or0;
  assign f_arrdiv32_fs298_or0 = f_arrdiv32_fs298_and1 | f_arrdiv32_fs298_and0;
  assign f_arrdiv32_fs299_xor0 = f_arrdiv32_mux2to1258_xor0 ^ b[11];
  assign f_arrdiv32_fs299_not0 = ~f_arrdiv32_mux2to1258_xor0;
  assign f_arrdiv32_fs299_and0 = f_arrdiv32_fs299_not0 & b[11];
  assign f_arrdiv32_fs299_xor1 = f_arrdiv32_fs298_or0 ^ f_arrdiv32_fs299_xor0;
  assign f_arrdiv32_fs299_not1 = ~f_arrdiv32_fs299_xor0;
  assign f_arrdiv32_fs299_and1 = f_arrdiv32_fs299_not1 & f_arrdiv32_fs298_or0;
  assign f_arrdiv32_fs299_or0 = f_arrdiv32_fs299_and1 | f_arrdiv32_fs299_and0;
  assign f_arrdiv32_fs300_xor0 = f_arrdiv32_mux2to1259_xor0 ^ b[12];
  assign f_arrdiv32_fs300_not0 = ~f_arrdiv32_mux2to1259_xor0;
  assign f_arrdiv32_fs300_and0 = f_arrdiv32_fs300_not0 & b[12];
  assign f_arrdiv32_fs300_xor1 = f_arrdiv32_fs299_or0 ^ f_arrdiv32_fs300_xor0;
  assign f_arrdiv32_fs300_not1 = ~f_arrdiv32_fs300_xor0;
  assign f_arrdiv32_fs300_and1 = f_arrdiv32_fs300_not1 & f_arrdiv32_fs299_or0;
  assign f_arrdiv32_fs300_or0 = f_arrdiv32_fs300_and1 | f_arrdiv32_fs300_and0;
  assign f_arrdiv32_fs301_xor0 = f_arrdiv32_mux2to1260_xor0 ^ b[13];
  assign f_arrdiv32_fs301_not0 = ~f_arrdiv32_mux2to1260_xor0;
  assign f_arrdiv32_fs301_and0 = f_arrdiv32_fs301_not0 & b[13];
  assign f_arrdiv32_fs301_xor1 = f_arrdiv32_fs300_or0 ^ f_arrdiv32_fs301_xor0;
  assign f_arrdiv32_fs301_not1 = ~f_arrdiv32_fs301_xor0;
  assign f_arrdiv32_fs301_and1 = f_arrdiv32_fs301_not1 & f_arrdiv32_fs300_or0;
  assign f_arrdiv32_fs301_or0 = f_arrdiv32_fs301_and1 | f_arrdiv32_fs301_and0;
  assign f_arrdiv32_fs302_xor0 = f_arrdiv32_mux2to1261_xor0 ^ b[14];
  assign f_arrdiv32_fs302_not0 = ~f_arrdiv32_mux2to1261_xor0;
  assign f_arrdiv32_fs302_and0 = f_arrdiv32_fs302_not0 & b[14];
  assign f_arrdiv32_fs302_xor1 = f_arrdiv32_fs301_or0 ^ f_arrdiv32_fs302_xor0;
  assign f_arrdiv32_fs302_not1 = ~f_arrdiv32_fs302_xor0;
  assign f_arrdiv32_fs302_and1 = f_arrdiv32_fs302_not1 & f_arrdiv32_fs301_or0;
  assign f_arrdiv32_fs302_or0 = f_arrdiv32_fs302_and1 | f_arrdiv32_fs302_and0;
  assign f_arrdiv32_fs303_xor0 = f_arrdiv32_mux2to1262_xor0 ^ b[15];
  assign f_arrdiv32_fs303_not0 = ~f_arrdiv32_mux2to1262_xor0;
  assign f_arrdiv32_fs303_and0 = f_arrdiv32_fs303_not0 & b[15];
  assign f_arrdiv32_fs303_xor1 = f_arrdiv32_fs302_or0 ^ f_arrdiv32_fs303_xor0;
  assign f_arrdiv32_fs303_not1 = ~f_arrdiv32_fs303_xor0;
  assign f_arrdiv32_fs303_and1 = f_arrdiv32_fs303_not1 & f_arrdiv32_fs302_or0;
  assign f_arrdiv32_fs303_or0 = f_arrdiv32_fs303_and1 | f_arrdiv32_fs303_and0;
  assign f_arrdiv32_fs304_xor0 = f_arrdiv32_mux2to1263_xor0 ^ b[16];
  assign f_arrdiv32_fs304_not0 = ~f_arrdiv32_mux2to1263_xor0;
  assign f_arrdiv32_fs304_and0 = f_arrdiv32_fs304_not0 & b[16];
  assign f_arrdiv32_fs304_xor1 = f_arrdiv32_fs303_or0 ^ f_arrdiv32_fs304_xor0;
  assign f_arrdiv32_fs304_not1 = ~f_arrdiv32_fs304_xor0;
  assign f_arrdiv32_fs304_and1 = f_arrdiv32_fs304_not1 & f_arrdiv32_fs303_or0;
  assign f_arrdiv32_fs304_or0 = f_arrdiv32_fs304_and1 | f_arrdiv32_fs304_and0;
  assign f_arrdiv32_fs305_xor0 = f_arrdiv32_mux2to1264_xor0 ^ b[17];
  assign f_arrdiv32_fs305_not0 = ~f_arrdiv32_mux2to1264_xor0;
  assign f_arrdiv32_fs305_and0 = f_arrdiv32_fs305_not0 & b[17];
  assign f_arrdiv32_fs305_xor1 = f_arrdiv32_fs304_or0 ^ f_arrdiv32_fs305_xor0;
  assign f_arrdiv32_fs305_not1 = ~f_arrdiv32_fs305_xor0;
  assign f_arrdiv32_fs305_and1 = f_arrdiv32_fs305_not1 & f_arrdiv32_fs304_or0;
  assign f_arrdiv32_fs305_or0 = f_arrdiv32_fs305_and1 | f_arrdiv32_fs305_and0;
  assign f_arrdiv32_fs306_xor0 = f_arrdiv32_mux2to1265_xor0 ^ b[18];
  assign f_arrdiv32_fs306_not0 = ~f_arrdiv32_mux2to1265_xor0;
  assign f_arrdiv32_fs306_and0 = f_arrdiv32_fs306_not0 & b[18];
  assign f_arrdiv32_fs306_xor1 = f_arrdiv32_fs305_or0 ^ f_arrdiv32_fs306_xor0;
  assign f_arrdiv32_fs306_not1 = ~f_arrdiv32_fs306_xor0;
  assign f_arrdiv32_fs306_and1 = f_arrdiv32_fs306_not1 & f_arrdiv32_fs305_or0;
  assign f_arrdiv32_fs306_or0 = f_arrdiv32_fs306_and1 | f_arrdiv32_fs306_and0;
  assign f_arrdiv32_fs307_xor0 = f_arrdiv32_mux2to1266_xor0 ^ b[19];
  assign f_arrdiv32_fs307_not0 = ~f_arrdiv32_mux2to1266_xor0;
  assign f_arrdiv32_fs307_and0 = f_arrdiv32_fs307_not0 & b[19];
  assign f_arrdiv32_fs307_xor1 = f_arrdiv32_fs306_or0 ^ f_arrdiv32_fs307_xor0;
  assign f_arrdiv32_fs307_not1 = ~f_arrdiv32_fs307_xor0;
  assign f_arrdiv32_fs307_and1 = f_arrdiv32_fs307_not1 & f_arrdiv32_fs306_or0;
  assign f_arrdiv32_fs307_or0 = f_arrdiv32_fs307_and1 | f_arrdiv32_fs307_and0;
  assign f_arrdiv32_fs308_xor0 = f_arrdiv32_mux2to1267_xor0 ^ b[20];
  assign f_arrdiv32_fs308_not0 = ~f_arrdiv32_mux2to1267_xor0;
  assign f_arrdiv32_fs308_and0 = f_arrdiv32_fs308_not0 & b[20];
  assign f_arrdiv32_fs308_xor1 = f_arrdiv32_fs307_or0 ^ f_arrdiv32_fs308_xor0;
  assign f_arrdiv32_fs308_not1 = ~f_arrdiv32_fs308_xor0;
  assign f_arrdiv32_fs308_and1 = f_arrdiv32_fs308_not1 & f_arrdiv32_fs307_or0;
  assign f_arrdiv32_fs308_or0 = f_arrdiv32_fs308_and1 | f_arrdiv32_fs308_and0;
  assign f_arrdiv32_fs309_xor0 = f_arrdiv32_mux2to1268_xor0 ^ b[21];
  assign f_arrdiv32_fs309_not0 = ~f_arrdiv32_mux2to1268_xor0;
  assign f_arrdiv32_fs309_and0 = f_arrdiv32_fs309_not0 & b[21];
  assign f_arrdiv32_fs309_xor1 = f_arrdiv32_fs308_or0 ^ f_arrdiv32_fs309_xor0;
  assign f_arrdiv32_fs309_not1 = ~f_arrdiv32_fs309_xor0;
  assign f_arrdiv32_fs309_and1 = f_arrdiv32_fs309_not1 & f_arrdiv32_fs308_or0;
  assign f_arrdiv32_fs309_or0 = f_arrdiv32_fs309_and1 | f_arrdiv32_fs309_and0;
  assign f_arrdiv32_fs310_xor0 = f_arrdiv32_mux2to1269_xor0 ^ b[22];
  assign f_arrdiv32_fs310_not0 = ~f_arrdiv32_mux2to1269_xor0;
  assign f_arrdiv32_fs310_and0 = f_arrdiv32_fs310_not0 & b[22];
  assign f_arrdiv32_fs310_xor1 = f_arrdiv32_fs309_or0 ^ f_arrdiv32_fs310_xor0;
  assign f_arrdiv32_fs310_not1 = ~f_arrdiv32_fs310_xor0;
  assign f_arrdiv32_fs310_and1 = f_arrdiv32_fs310_not1 & f_arrdiv32_fs309_or0;
  assign f_arrdiv32_fs310_or0 = f_arrdiv32_fs310_and1 | f_arrdiv32_fs310_and0;
  assign f_arrdiv32_fs311_xor0 = f_arrdiv32_mux2to1270_xor0 ^ b[23];
  assign f_arrdiv32_fs311_not0 = ~f_arrdiv32_mux2to1270_xor0;
  assign f_arrdiv32_fs311_and0 = f_arrdiv32_fs311_not0 & b[23];
  assign f_arrdiv32_fs311_xor1 = f_arrdiv32_fs310_or0 ^ f_arrdiv32_fs311_xor0;
  assign f_arrdiv32_fs311_not1 = ~f_arrdiv32_fs311_xor0;
  assign f_arrdiv32_fs311_and1 = f_arrdiv32_fs311_not1 & f_arrdiv32_fs310_or0;
  assign f_arrdiv32_fs311_or0 = f_arrdiv32_fs311_and1 | f_arrdiv32_fs311_and0;
  assign f_arrdiv32_fs312_xor0 = f_arrdiv32_mux2to1271_xor0 ^ b[24];
  assign f_arrdiv32_fs312_not0 = ~f_arrdiv32_mux2to1271_xor0;
  assign f_arrdiv32_fs312_and0 = f_arrdiv32_fs312_not0 & b[24];
  assign f_arrdiv32_fs312_xor1 = f_arrdiv32_fs311_or0 ^ f_arrdiv32_fs312_xor0;
  assign f_arrdiv32_fs312_not1 = ~f_arrdiv32_fs312_xor0;
  assign f_arrdiv32_fs312_and1 = f_arrdiv32_fs312_not1 & f_arrdiv32_fs311_or0;
  assign f_arrdiv32_fs312_or0 = f_arrdiv32_fs312_and1 | f_arrdiv32_fs312_and0;
  assign f_arrdiv32_fs313_xor0 = f_arrdiv32_mux2to1272_xor0 ^ b[25];
  assign f_arrdiv32_fs313_not0 = ~f_arrdiv32_mux2to1272_xor0;
  assign f_arrdiv32_fs313_and0 = f_arrdiv32_fs313_not0 & b[25];
  assign f_arrdiv32_fs313_xor1 = f_arrdiv32_fs312_or0 ^ f_arrdiv32_fs313_xor0;
  assign f_arrdiv32_fs313_not1 = ~f_arrdiv32_fs313_xor0;
  assign f_arrdiv32_fs313_and1 = f_arrdiv32_fs313_not1 & f_arrdiv32_fs312_or0;
  assign f_arrdiv32_fs313_or0 = f_arrdiv32_fs313_and1 | f_arrdiv32_fs313_and0;
  assign f_arrdiv32_fs314_xor0 = f_arrdiv32_mux2to1273_xor0 ^ b[26];
  assign f_arrdiv32_fs314_not0 = ~f_arrdiv32_mux2to1273_xor0;
  assign f_arrdiv32_fs314_and0 = f_arrdiv32_fs314_not0 & b[26];
  assign f_arrdiv32_fs314_xor1 = f_arrdiv32_fs313_or0 ^ f_arrdiv32_fs314_xor0;
  assign f_arrdiv32_fs314_not1 = ~f_arrdiv32_fs314_xor0;
  assign f_arrdiv32_fs314_and1 = f_arrdiv32_fs314_not1 & f_arrdiv32_fs313_or0;
  assign f_arrdiv32_fs314_or0 = f_arrdiv32_fs314_and1 | f_arrdiv32_fs314_and0;
  assign f_arrdiv32_fs315_xor0 = f_arrdiv32_mux2to1274_xor0 ^ b[27];
  assign f_arrdiv32_fs315_not0 = ~f_arrdiv32_mux2to1274_xor0;
  assign f_arrdiv32_fs315_and0 = f_arrdiv32_fs315_not0 & b[27];
  assign f_arrdiv32_fs315_xor1 = f_arrdiv32_fs314_or0 ^ f_arrdiv32_fs315_xor0;
  assign f_arrdiv32_fs315_not1 = ~f_arrdiv32_fs315_xor0;
  assign f_arrdiv32_fs315_and1 = f_arrdiv32_fs315_not1 & f_arrdiv32_fs314_or0;
  assign f_arrdiv32_fs315_or0 = f_arrdiv32_fs315_and1 | f_arrdiv32_fs315_and0;
  assign f_arrdiv32_fs316_xor0 = f_arrdiv32_mux2to1275_xor0 ^ b[28];
  assign f_arrdiv32_fs316_not0 = ~f_arrdiv32_mux2to1275_xor0;
  assign f_arrdiv32_fs316_and0 = f_arrdiv32_fs316_not0 & b[28];
  assign f_arrdiv32_fs316_xor1 = f_arrdiv32_fs315_or0 ^ f_arrdiv32_fs316_xor0;
  assign f_arrdiv32_fs316_not1 = ~f_arrdiv32_fs316_xor0;
  assign f_arrdiv32_fs316_and1 = f_arrdiv32_fs316_not1 & f_arrdiv32_fs315_or0;
  assign f_arrdiv32_fs316_or0 = f_arrdiv32_fs316_and1 | f_arrdiv32_fs316_and0;
  assign f_arrdiv32_fs317_xor0 = f_arrdiv32_mux2to1276_xor0 ^ b[29];
  assign f_arrdiv32_fs317_not0 = ~f_arrdiv32_mux2to1276_xor0;
  assign f_arrdiv32_fs317_and0 = f_arrdiv32_fs317_not0 & b[29];
  assign f_arrdiv32_fs317_xor1 = f_arrdiv32_fs316_or0 ^ f_arrdiv32_fs317_xor0;
  assign f_arrdiv32_fs317_not1 = ~f_arrdiv32_fs317_xor0;
  assign f_arrdiv32_fs317_and1 = f_arrdiv32_fs317_not1 & f_arrdiv32_fs316_or0;
  assign f_arrdiv32_fs317_or0 = f_arrdiv32_fs317_and1 | f_arrdiv32_fs317_and0;
  assign f_arrdiv32_fs318_xor0 = f_arrdiv32_mux2to1277_xor0 ^ b[30];
  assign f_arrdiv32_fs318_not0 = ~f_arrdiv32_mux2to1277_xor0;
  assign f_arrdiv32_fs318_and0 = f_arrdiv32_fs318_not0 & b[30];
  assign f_arrdiv32_fs318_xor1 = f_arrdiv32_fs317_or0 ^ f_arrdiv32_fs318_xor0;
  assign f_arrdiv32_fs318_not1 = ~f_arrdiv32_fs318_xor0;
  assign f_arrdiv32_fs318_and1 = f_arrdiv32_fs318_not1 & f_arrdiv32_fs317_or0;
  assign f_arrdiv32_fs318_or0 = f_arrdiv32_fs318_and1 | f_arrdiv32_fs318_and0;
  assign f_arrdiv32_fs319_xor0 = f_arrdiv32_mux2to1278_xor0 ^ b[31];
  assign f_arrdiv32_fs319_not0 = ~f_arrdiv32_mux2to1278_xor0;
  assign f_arrdiv32_fs319_and0 = f_arrdiv32_fs319_not0 & b[31];
  assign f_arrdiv32_fs319_xor1 = f_arrdiv32_fs318_or0 ^ f_arrdiv32_fs319_xor0;
  assign f_arrdiv32_fs319_not1 = ~f_arrdiv32_fs319_xor0;
  assign f_arrdiv32_fs319_and1 = f_arrdiv32_fs319_not1 & f_arrdiv32_fs318_or0;
  assign f_arrdiv32_fs319_or0 = f_arrdiv32_fs319_and1 | f_arrdiv32_fs319_and0;
  assign f_arrdiv32_mux2to1279_and0 = a[22] & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1279_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1279_and1 = f_arrdiv32_fs288_xor0 & f_arrdiv32_mux2to1279_not0;
  assign f_arrdiv32_mux2to1279_xor0 = f_arrdiv32_mux2to1279_and0 ^ f_arrdiv32_mux2to1279_and1;
  assign f_arrdiv32_mux2to1280_and0 = f_arrdiv32_mux2to1248_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1280_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1280_and1 = f_arrdiv32_fs289_xor1 & f_arrdiv32_mux2to1280_not0;
  assign f_arrdiv32_mux2to1280_xor0 = f_arrdiv32_mux2to1280_and0 ^ f_arrdiv32_mux2to1280_and1;
  assign f_arrdiv32_mux2to1281_and0 = f_arrdiv32_mux2to1249_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1281_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1281_and1 = f_arrdiv32_fs290_xor1 & f_arrdiv32_mux2to1281_not0;
  assign f_arrdiv32_mux2to1281_xor0 = f_arrdiv32_mux2to1281_and0 ^ f_arrdiv32_mux2to1281_and1;
  assign f_arrdiv32_mux2to1282_and0 = f_arrdiv32_mux2to1250_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1282_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1282_and1 = f_arrdiv32_fs291_xor1 & f_arrdiv32_mux2to1282_not0;
  assign f_arrdiv32_mux2to1282_xor0 = f_arrdiv32_mux2to1282_and0 ^ f_arrdiv32_mux2to1282_and1;
  assign f_arrdiv32_mux2to1283_and0 = f_arrdiv32_mux2to1251_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1283_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1283_and1 = f_arrdiv32_fs292_xor1 & f_arrdiv32_mux2to1283_not0;
  assign f_arrdiv32_mux2to1283_xor0 = f_arrdiv32_mux2to1283_and0 ^ f_arrdiv32_mux2to1283_and1;
  assign f_arrdiv32_mux2to1284_and0 = f_arrdiv32_mux2to1252_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1284_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1284_and1 = f_arrdiv32_fs293_xor1 & f_arrdiv32_mux2to1284_not0;
  assign f_arrdiv32_mux2to1284_xor0 = f_arrdiv32_mux2to1284_and0 ^ f_arrdiv32_mux2to1284_and1;
  assign f_arrdiv32_mux2to1285_and0 = f_arrdiv32_mux2to1253_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1285_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1285_and1 = f_arrdiv32_fs294_xor1 & f_arrdiv32_mux2to1285_not0;
  assign f_arrdiv32_mux2to1285_xor0 = f_arrdiv32_mux2to1285_and0 ^ f_arrdiv32_mux2to1285_and1;
  assign f_arrdiv32_mux2to1286_and0 = f_arrdiv32_mux2to1254_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1286_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1286_and1 = f_arrdiv32_fs295_xor1 & f_arrdiv32_mux2to1286_not0;
  assign f_arrdiv32_mux2to1286_xor0 = f_arrdiv32_mux2to1286_and0 ^ f_arrdiv32_mux2to1286_and1;
  assign f_arrdiv32_mux2to1287_and0 = f_arrdiv32_mux2to1255_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1287_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1287_and1 = f_arrdiv32_fs296_xor1 & f_arrdiv32_mux2to1287_not0;
  assign f_arrdiv32_mux2to1287_xor0 = f_arrdiv32_mux2to1287_and0 ^ f_arrdiv32_mux2to1287_and1;
  assign f_arrdiv32_mux2to1288_and0 = f_arrdiv32_mux2to1256_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1288_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1288_and1 = f_arrdiv32_fs297_xor1 & f_arrdiv32_mux2to1288_not0;
  assign f_arrdiv32_mux2to1288_xor0 = f_arrdiv32_mux2to1288_and0 ^ f_arrdiv32_mux2to1288_and1;
  assign f_arrdiv32_mux2to1289_and0 = f_arrdiv32_mux2to1257_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1289_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1289_and1 = f_arrdiv32_fs298_xor1 & f_arrdiv32_mux2to1289_not0;
  assign f_arrdiv32_mux2to1289_xor0 = f_arrdiv32_mux2to1289_and0 ^ f_arrdiv32_mux2to1289_and1;
  assign f_arrdiv32_mux2to1290_and0 = f_arrdiv32_mux2to1258_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1290_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1290_and1 = f_arrdiv32_fs299_xor1 & f_arrdiv32_mux2to1290_not0;
  assign f_arrdiv32_mux2to1290_xor0 = f_arrdiv32_mux2to1290_and0 ^ f_arrdiv32_mux2to1290_and1;
  assign f_arrdiv32_mux2to1291_and0 = f_arrdiv32_mux2to1259_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1291_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1291_and1 = f_arrdiv32_fs300_xor1 & f_arrdiv32_mux2to1291_not0;
  assign f_arrdiv32_mux2to1291_xor0 = f_arrdiv32_mux2to1291_and0 ^ f_arrdiv32_mux2to1291_and1;
  assign f_arrdiv32_mux2to1292_and0 = f_arrdiv32_mux2to1260_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1292_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1292_and1 = f_arrdiv32_fs301_xor1 & f_arrdiv32_mux2to1292_not0;
  assign f_arrdiv32_mux2to1292_xor0 = f_arrdiv32_mux2to1292_and0 ^ f_arrdiv32_mux2to1292_and1;
  assign f_arrdiv32_mux2to1293_and0 = f_arrdiv32_mux2to1261_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1293_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1293_and1 = f_arrdiv32_fs302_xor1 & f_arrdiv32_mux2to1293_not0;
  assign f_arrdiv32_mux2to1293_xor0 = f_arrdiv32_mux2to1293_and0 ^ f_arrdiv32_mux2to1293_and1;
  assign f_arrdiv32_mux2to1294_and0 = f_arrdiv32_mux2to1262_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1294_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1294_and1 = f_arrdiv32_fs303_xor1 & f_arrdiv32_mux2to1294_not0;
  assign f_arrdiv32_mux2to1294_xor0 = f_arrdiv32_mux2to1294_and0 ^ f_arrdiv32_mux2to1294_and1;
  assign f_arrdiv32_mux2to1295_and0 = f_arrdiv32_mux2to1263_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1295_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1295_and1 = f_arrdiv32_fs304_xor1 & f_arrdiv32_mux2to1295_not0;
  assign f_arrdiv32_mux2to1295_xor0 = f_arrdiv32_mux2to1295_and0 ^ f_arrdiv32_mux2to1295_and1;
  assign f_arrdiv32_mux2to1296_and0 = f_arrdiv32_mux2to1264_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1296_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1296_and1 = f_arrdiv32_fs305_xor1 & f_arrdiv32_mux2to1296_not0;
  assign f_arrdiv32_mux2to1296_xor0 = f_arrdiv32_mux2to1296_and0 ^ f_arrdiv32_mux2to1296_and1;
  assign f_arrdiv32_mux2to1297_and0 = f_arrdiv32_mux2to1265_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1297_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1297_and1 = f_arrdiv32_fs306_xor1 & f_arrdiv32_mux2to1297_not0;
  assign f_arrdiv32_mux2to1297_xor0 = f_arrdiv32_mux2to1297_and0 ^ f_arrdiv32_mux2to1297_and1;
  assign f_arrdiv32_mux2to1298_and0 = f_arrdiv32_mux2to1266_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1298_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1298_and1 = f_arrdiv32_fs307_xor1 & f_arrdiv32_mux2to1298_not0;
  assign f_arrdiv32_mux2to1298_xor0 = f_arrdiv32_mux2to1298_and0 ^ f_arrdiv32_mux2to1298_and1;
  assign f_arrdiv32_mux2to1299_and0 = f_arrdiv32_mux2to1267_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1299_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1299_and1 = f_arrdiv32_fs308_xor1 & f_arrdiv32_mux2to1299_not0;
  assign f_arrdiv32_mux2to1299_xor0 = f_arrdiv32_mux2to1299_and0 ^ f_arrdiv32_mux2to1299_and1;
  assign f_arrdiv32_mux2to1300_and0 = f_arrdiv32_mux2to1268_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1300_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1300_and1 = f_arrdiv32_fs309_xor1 & f_arrdiv32_mux2to1300_not0;
  assign f_arrdiv32_mux2to1300_xor0 = f_arrdiv32_mux2to1300_and0 ^ f_arrdiv32_mux2to1300_and1;
  assign f_arrdiv32_mux2to1301_and0 = f_arrdiv32_mux2to1269_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1301_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1301_and1 = f_arrdiv32_fs310_xor1 & f_arrdiv32_mux2to1301_not0;
  assign f_arrdiv32_mux2to1301_xor0 = f_arrdiv32_mux2to1301_and0 ^ f_arrdiv32_mux2to1301_and1;
  assign f_arrdiv32_mux2to1302_and0 = f_arrdiv32_mux2to1270_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1302_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1302_and1 = f_arrdiv32_fs311_xor1 & f_arrdiv32_mux2to1302_not0;
  assign f_arrdiv32_mux2to1302_xor0 = f_arrdiv32_mux2to1302_and0 ^ f_arrdiv32_mux2to1302_and1;
  assign f_arrdiv32_mux2to1303_and0 = f_arrdiv32_mux2to1271_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1303_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1303_and1 = f_arrdiv32_fs312_xor1 & f_arrdiv32_mux2to1303_not0;
  assign f_arrdiv32_mux2to1303_xor0 = f_arrdiv32_mux2to1303_and0 ^ f_arrdiv32_mux2to1303_and1;
  assign f_arrdiv32_mux2to1304_and0 = f_arrdiv32_mux2to1272_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1304_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1304_and1 = f_arrdiv32_fs313_xor1 & f_arrdiv32_mux2to1304_not0;
  assign f_arrdiv32_mux2to1304_xor0 = f_arrdiv32_mux2to1304_and0 ^ f_arrdiv32_mux2to1304_and1;
  assign f_arrdiv32_mux2to1305_and0 = f_arrdiv32_mux2to1273_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1305_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1305_and1 = f_arrdiv32_fs314_xor1 & f_arrdiv32_mux2to1305_not0;
  assign f_arrdiv32_mux2to1305_xor0 = f_arrdiv32_mux2to1305_and0 ^ f_arrdiv32_mux2to1305_and1;
  assign f_arrdiv32_mux2to1306_and0 = f_arrdiv32_mux2to1274_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1306_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1306_and1 = f_arrdiv32_fs315_xor1 & f_arrdiv32_mux2to1306_not0;
  assign f_arrdiv32_mux2to1306_xor0 = f_arrdiv32_mux2to1306_and0 ^ f_arrdiv32_mux2to1306_and1;
  assign f_arrdiv32_mux2to1307_and0 = f_arrdiv32_mux2to1275_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1307_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1307_and1 = f_arrdiv32_fs316_xor1 & f_arrdiv32_mux2to1307_not0;
  assign f_arrdiv32_mux2to1307_xor0 = f_arrdiv32_mux2to1307_and0 ^ f_arrdiv32_mux2to1307_and1;
  assign f_arrdiv32_mux2to1308_and0 = f_arrdiv32_mux2to1276_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1308_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1308_and1 = f_arrdiv32_fs317_xor1 & f_arrdiv32_mux2to1308_not0;
  assign f_arrdiv32_mux2to1308_xor0 = f_arrdiv32_mux2to1308_and0 ^ f_arrdiv32_mux2to1308_and1;
  assign f_arrdiv32_mux2to1309_and0 = f_arrdiv32_mux2to1277_xor0 & f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1309_not0 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_mux2to1309_and1 = f_arrdiv32_fs318_xor1 & f_arrdiv32_mux2to1309_not0;
  assign f_arrdiv32_mux2to1309_xor0 = f_arrdiv32_mux2to1309_and0 ^ f_arrdiv32_mux2to1309_and1;
  assign f_arrdiv32_not9 = ~f_arrdiv32_fs319_or0;
  assign f_arrdiv32_fs320_xor0 = a[21] ^ b[0];
  assign f_arrdiv32_fs320_not0 = ~a[21];
  assign f_arrdiv32_fs320_and0 = f_arrdiv32_fs320_not0 & b[0];
  assign f_arrdiv32_fs320_not1 = ~f_arrdiv32_fs320_xor0;
  assign f_arrdiv32_fs321_xor0 = f_arrdiv32_mux2to1279_xor0 ^ b[1];
  assign f_arrdiv32_fs321_not0 = ~f_arrdiv32_mux2to1279_xor0;
  assign f_arrdiv32_fs321_and0 = f_arrdiv32_fs321_not0 & b[1];
  assign f_arrdiv32_fs321_xor1 = f_arrdiv32_fs320_and0 ^ f_arrdiv32_fs321_xor0;
  assign f_arrdiv32_fs321_not1 = ~f_arrdiv32_fs321_xor0;
  assign f_arrdiv32_fs321_and1 = f_arrdiv32_fs321_not1 & f_arrdiv32_fs320_and0;
  assign f_arrdiv32_fs321_or0 = f_arrdiv32_fs321_and1 | f_arrdiv32_fs321_and0;
  assign f_arrdiv32_fs322_xor0 = f_arrdiv32_mux2to1280_xor0 ^ b[2];
  assign f_arrdiv32_fs322_not0 = ~f_arrdiv32_mux2to1280_xor0;
  assign f_arrdiv32_fs322_and0 = f_arrdiv32_fs322_not0 & b[2];
  assign f_arrdiv32_fs322_xor1 = f_arrdiv32_fs321_or0 ^ f_arrdiv32_fs322_xor0;
  assign f_arrdiv32_fs322_not1 = ~f_arrdiv32_fs322_xor0;
  assign f_arrdiv32_fs322_and1 = f_arrdiv32_fs322_not1 & f_arrdiv32_fs321_or0;
  assign f_arrdiv32_fs322_or0 = f_arrdiv32_fs322_and1 | f_arrdiv32_fs322_and0;
  assign f_arrdiv32_fs323_xor0 = f_arrdiv32_mux2to1281_xor0 ^ b[3];
  assign f_arrdiv32_fs323_not0 = ~f_arrdiv32_mux2to1281_xor0;
  assign f_arrdiv32_fs323_and0 = f_arrdiv32_fs323_not0 & b[3];
  assign f_arrdiv32_fs323_xor1 = f_arrdiv32_fs322_or0 ^ f_arrdiv32_fs323_xor0;
  assign f_arrdiv32_fs323_not1 = ~f_arrdiv32_fs323_xor0;
  assign f_arrdiv32_fs323_and1 = f_arrdiv32_fs323_not1 & f_arrdiv32_fs322_or0;
  assign f_arrdiv32_fs323_or0 = f_arrdiv32_fs323_and1 | f_arrdiv32_fs323_and0;
  assign f_arrdiv32_fs324_xor0 = f_arrdiv32_mux2to1282_xor0 ^ b[4];
  assign f_arrdiv32_fs324_not0 = ~f_arrdiv32_mux2to1282_xor0;
  assign f_arrdiv32_fs324_and0 = f_arrdiv32_fs324_not0 & b[4];
  assign f_arrdiv32_fs324_xor1 = f_arrdiv32_fs323_or0 ^ f_arrdiv32_fs324_xor0;
  assign f_arrdiv32_fs324_not1 = ~f_arrdiv32_fs324_xor0;
  assign f_arrdiv32_fs324_and1 = f_arrdiv32_fs324_not1 & f_arrdiv32_fs323_or0;
  assign f_arrdiv32_fs324_or0 = f_arrdiv32_fs324_and1 | f_arrdiv32_fs324_and0;
  assign f_arrdiv32_fs325_xor0 = f_arrdiv32_mux2to1283_xor0 ^ b[5];
  assign f_arrdiv32_fs325_not0 = ~f_arrdiv32_mux2to1283_xor0;
  assign f_arrdiv32_fs325_and0 = f_arrdiv32_fs325_not0 & b[5];
  assign f_arrdiv32_fs325_xor1 = f_arrdiv32_fs324_or0 ^ f_arrdiv32_fs325_xor0;
  assign f_arrdiv32_fs325_not1 = ~f_arrdiv32_fs325_xor0;
  assign f_arrdiv32_fs325_and1 = f_arrdiv32_fs325_not1 & f_arrdiv32_fs324_or0;
  assign f_arrdiv32_fs325_or0 = f_arrdiv32_fs325_and1 | f_arrdiv32_fs325_and0;
  assign f_arrdiv32_fs326_xor0 = f_arrdiv32_mux2to1284_xor0 ^ b[6];
  assign f_arrdiv32_fs326_not0 = ~f_arrdiv32_mux2to1284_xor0;
  assign f_arrdiv32_fs326_and0 = f_arrdiv32_fs326_not0 & b[6];
  assign f_arrdiv32_fs326_xor1 = f_arrdiv32_fs325_or0 ^ f_arrdiv32_fs326_xor0;
  assign f_arrdiv32_fs326_not1 = ~f_arrdiv32_fs326_xor0;
  assign f_arrdiv32_fs326_and1 = f_arrdiv32_fs326_not1 & f_arrdiv32_fs325_or0;
  assign f_arrdiv32_fs326_or0 = f_arrdiv32_fs326_and1 | f_arrdiv32_fs326_and0;
  assign f_arrdiv32_fs327_xor0 = f_arrdiv32_mux2to1285_xor0 ^ b[7];
  assign f_arrdiv32_fs327_not0 = ~f_arrdiv32_mux2to1285_xor0;
  assign f_arrdiv32_fs327_and0 = f_arrdiv32_fs327_not0 & b[7];
  assign f_arrdiv32_fs327_xor1 = f_arrdiv32_fs326_or0 ^ f_arrdiv32_fs327_xor0;
  assign f_arrdiv32_fs327_not1 = ~f_arrdiv32_fs327_xor0;
  assign f_arrdiv32_fs327_and1 = f_arrdiv32_fs327_not1 & f_arrdiv32_fs326_or0;
  assign f_arrdiv32_fs327_or0 = f_arrdiv32_fs327_and1 | f_arrdiv32_fs327_and0;
  assign f_arrdiv32_fs328_xor0 = f_arrdiv32_mux2to1286_xor0 ^ b[8];
  assign f_arrdiv32_fs328_not0 = ~f_arrdiv32_mux2to1286_xor0;
  assign f_arrdiv32_fs328_and0 = f_arrdiv32_fs328_not0 & b[8];
  assign f_arrdiv32_fs328_xor1 = f_arrdiv32_fs327_or0 ^ f_arrdiv32_fs328_xor0;
  assign f_arrdiv32_fs328_not1 = ~f_arrdiv32_fs328_xor0;
  assign f_arrdiv32_fs328_and1 = f_arrdiv32_fs328_not1 & f_arrdiv32_fs327_or0;
  assign f_arrdiv32_fs328_or0 = f_arrdiv32_fs328_and1 | f_arrdiv32_fs328_and0;
  assign f_arrdiv32_fs329_xor0 = f_arrdiv32_mux2to1287_xor0 ^ b[9];
  assign f_arrdiv32_fs329_not0 = ~f_arrdiv32_mux2to1287_xor0;
  assign f_arrdiv32_fs329_and0 = f_arrdiv32_fs329_not0 & b[9];
  assign f_arrdiv32_fs329_xor1 = f_arrdiv32_fs328_or0 ^ f_arrdiv32_fs329_xor0;
  assign f_arrdiv32_fs329_not1 = ~f_arrdiv32_fs329_xor0;
  assign f_arrdiv32_fs329_and1 = f_arrdiv32_fs329_not1 & f_arrdiv32_fs328_or0;
  assign f_arrdiv32_fs329_or0 = f_arrdiv32_fs329_and1 | f_arrdiv32_fs329_and0;
  assign f_arrdiv32_fs330_xor0 = f_arrdiv32_mux2to1288_xor0 ^ b[10];
  assign f_arrdiv32_fs330_not0 = ~f_arrdiv32_mux2to1288_xor0;
  assign f_arrdiv32_fs330_and0 = f_arrdiv32_fs330_not0 & b[10];
  assign f_arrdiv32_fs330_xor1 = f_arrdiv32_fs329_or0 ^ f_arrdiv32_fs330_xor0;
  assign f_arrdiv32_fs330_not1 = ~f_arrdiv32_fs330_xor0;
  assign f_arrdiv32_fs330_and1 = f_arrdiv32_fs330_not1 & f_arrdiv32_fs329_or0;
  assign f_arrdiv32_fs330_or0 = f_arrdiv32_fs330_and1 | f_arrdiv32_fs330_and0;
  assign f_arrdiv32_fs331_xor0 = f_arrdiv32_mux2to1289_xor0 ^ b[11];
  assign f_arrdiv32_fs331_not0 = ~f_arrdiv32_mux2to1289_xor0;
  assign f_arrdiv32_fs331_and0 = f_arrdiv32_fs331_not0 & b[11];
  assign f_arrdiv32_fs331_xor1 = f_arrdiv32_fs330_or0 ^ f_arrdiv32_fs331_xor0;
  assign f_arrdiv32_fs331_not1 = ~f_arrdiv32_fs331_xor0;
  assign f_arrdiv32_fs331_and1 = f_arrdiv32_fs331_not1 & f_arrdiv32_fs330_or0;
  assign f_arrdiv32_fs331_or0 = f_arrdiv32_fs331_and1 | f_arrdiv32_fs331_and0;
  assign f_arrdiv32_fs332_xor0 = f_arrdiv32_mux2to1290_xor0 ^ b[12];
  assign f_arrdiv32_fs332_not0 = ~f_arrdiv32_mux2to1290_xor0;
  assign f_arrdiv32_fs332_and0 = f_arrdiv32_fs332_not0 & b[12];
  assign f_arrdiv32_fs332_xor1 = f_arrdiv32_fs331_or0 ^ f_arrdiv32_fs332_xor0;
  assign f_arrdiv32_fs332_not1 = ~f_arrdiv32_fs332_xor0;
  assign f_arrdiv32_fs332_and1 = f_arrdiv32_fs332_not1 & f_arrdiv32_fs331_or0;
  assign f_arrdiv32_fs332_or0 = f_arrdiv32_fs332_and1 | f_arrdiv32_fs332_and0;
  assign f_arrdiv32_fs333_xor0 = f_arrdiv32_mux2to1291_xor0 ^ b[13];
  assign f_arrdiv32_fs333_not0 = ~f_arrdiv32_mux2to1291_xor0;
  assign f_arrdiv32_fs333_and0 = f_arrdiv32_fs333_not0 & b[13];
  assign f_arrdiv32_fs333_xor1 = f_arrdiv32_fs332_or0 ^ f_arrdiv32_fs333_xor0;
  assign f_arrdiv32_fs333_not1 = ~f_arrdiv32_fs333_xor0;
  assign f_arrdiv32_fs333_and1 = f_arrdiv32_fs333_not1 & f_arrdiv32_fs332_or0;
  assign f_arrdiv32_fs333_or0 = f_arrdiv32_fs333_and1 | f_arrdiv32_fs333_and0;
  assign f_arrdiv32_fs334_xor0 = f_arrdiv32_mux2to1292_xor0 ^ b[14];
  assign f_arrdiv32_fs334_not0 = ~f_arrdiv32_mux2to1292_xor0;
  assign f_arrdiv32_fs334_and0 = f_arrdiv32_fs334_not0 & b[14];
  assign f_arrdiv32_fs334_xor1 = f_arrdiv32_fs333_or0 ^ f_arrdiv32_fs334_xor0;
  assign f_arrdiv32_fs334_not1 = ~f_arrdiv32_fs334_xor0;
  assign f_arrdiv32_fs334_and1 = f_arrdiv32_fs334_not1 & f_arrdiv32_fs333_or0;
  assign f_arrdiv32_fs334_or0 = f_arrdiv32_fs334_and1 | f_arrdiv32_fs334_and0;
  assign f_arrdiv32_fs335_xor0 = f_arrdiv32_mux2to1293_xor0 ^ b[15];
  assign f_arrdiv32_fs335_not0 = ~f_arrdiv32_mux2to1293_xor0;
  assign f_arrdiv32_fs335_and0 = f_arrdiv32_fs335_not0 & b[15];
  assign f_arrdiv32_fs335_xor1 = f_arrdiv32_fs334_or0 ^ f_arrdiv32_fs335_xor0;
  assign f_arrdiv32_fs335_not1 = ~f_arrdiv32_fs335_xor0;
  assign f_arrdiv32_fs335_and1 = f_arrdiv32_fs335_not1 & f_arrdiv32_fs334_or0;
  assign f_arrdiv32_fs335_or0 = f_arrdiv32_fs335_and1 | f_arrdiv32_fs335_and0;
  assign f_arrdiv32_fs336_xor0 = f_arrdiv32_mux2to1294_xor0 ^ b[16];
  assign f_arrdiv32_fs336_not0 = ~f_arrdiv32_mux2to1294_xor0;
  assign f_arrdiv32_fs336_and0 = f_arrdiv32_fs336_not0 & b[16];
  assign f_arrdiv32_fs336_xor1 = f_arrdiv32_fs335_or0 ^ f_arrdiv32_fs336_xor0;
  assign f_arrdiv32_fs336_not1 = ~f_arrdiv32_fs336_xor0;
  assign f_arrdiv32_fs336_and1 = f_arrdiv32_fs336_not1 & f_arrdiv32_fs335_or0;
  assign f_arrdiv32_fs336_or0 = f_arrdiv32_fs336_and1 | f_arrdiv32_fs336_and0;
  assign f_arrdiv32_fs337_xor0 = f_arrdiv32_mux2to1295_xor0 ^ b[17];
  assign f_arrdiv32_fs337_not0 = ~f_arrdiv32_mux2to1295_xor0;
  assign f_arrdiv32_fs337_and0 = f_arrdiv32_fs337_not0 & b[17];
  assign f_arrdiv32_fs337_xor1 = f_arrdiv32_fs336_or0 ^ f_arrdiv32_fs337_xor0;
  assign f_arrdiv32_fs337_not1 = ~f_arrdiv32_fs337_xor0;
  assign f_arrdiv32_fs337_and1 = f_arrdiv32_fs337_not1 & f_arrdiv32_fs336_or0;
  assign f_arrdiv32_fs337_or0 = f_arrdiv32_fs337_and1 | f_arrdiv32_fs337_and0;
  assign f_arrdiv32_fs338_xor0 = f_arrdiv32_mux2to1296_xor0 ^ b[18];
  assign f_arrdiv32_fs338_not0 = ~f_arrdiv32_mux2to1296_xor0;
  assign f_arrdiv32_fs338_and0 = f_arrdiv32_fs338_not0 & b[18];
  assign f_arrdiv32_fs338_xor1 = f_arrdiv32_fs337_or0 ^ f_arrdiv32_fs338_xor0;
  assign f_arrdiv32_fs338_not1 = ~f_arrdiv32_fs338_xor0;
  assign f_arrdiv32_fs338_and1 = f_arrdiv32_fs338_not1 & f_arrdiv32_fs337_or0;
  assign f_arrdiv32_fs338_or0 = f_arrdiv32_fs338_and1 | f_arrdiv32_fs338_and0;
  assign f_arrdiv32_fs339_xor0 = f_arrdiv32_mux2to1297_xor0 ^ b[19];
  assign f_arrdiv32_fs339_not0 = ~f_arrdiv32_mux2to1297_xor0;
  assign f_arrdiv32_fs339_and0 = f_arrdiv32_fs339_not0 & b[19];
  assign f_arrdiv32_fs339_xor1 = f_arrdiv32_fs338_or0 ^ f_arrdiv32_fs339_xor0;
  assign f_arrdiv32_fs339_not1 = ~f_arrdiv32_fs339_xor0;
  assign f_arrdiv32_fs339_and1 = f_arrdiv32_fs339_not1 & f_arrdiv32_fs338_or0;
  assign f_arrdiv32_fs339_or0 = f_arrdiv32_fs339_and1 | f_arrdiv32_fs339_and0;
  assign f_arrdiv32_fs340_xor0 = f_arrdiv32_mux2to1298_xor0 ^ b[20];
  assign f_arrdiv32_fs340_not0 = ~f_arrdiv32_mux2to1298_xor0;
  assign f_arrdiv32_fs340_and0 = f_arrdiv32_fs340_not0 & b[20];
  assign f_arrdiv32_fs340_xor1 = f_arrdiv32_fs339_or0 ^ f_arrdiv32_fs340_xor0;
  assign f_arrdiv32_fs340_not1 = ~f_arrdiv32_fs340_xor0;
  assign f_arrdiv32_fs340_and1 = f_arrdiv32_fs340_not1 & f_arrdiv32_fs339_or0;
  assign f_arrdiv32_fs340_or0 = f_arrdiv32_fs340_and1 | f_arrdiv32_fs340_and0;
  assign f_arrdiv32_fs341_xor0 = f_arrdiv32_mux2to1299_xor0 ^ b[21];
  assign f_arrdiv32_fs341_not0 = ~f_arrdiv32_mux2to1299_xor0;
  assign f_arrdiv32_fs341_and0 = f_arrdiv32_fs341_not0 & b[21];
  assign f_arrdiv32_fs341_xor1 = f_arrdiv32_fs340_or0 ^ f_arrdiv32_fs341_xor0;
  assign f_arrdiv32_fs341_not1 = ~f_arrdiv32_fs341_xor0;
  assign f_arrdiv32_fs341_and1 = f_arrdiv32_fs341_not1 & f_arrdiv32_fs340_or0;
  assign f_arrdiv32_fs341_or0 = f_arrdiv32_fs341_and1 | f_arrdiv32_fs341_and0;
  assign f_arrdiv32_fs342_xor0 = f_arrdiv32_mux2to1300_xor0 ^ b[22];
  assign f_arrdiv32_fs342_not0 = ~f_arrdiv32_mux2to1300_xor0;
  assign f_arrdiv32_fs342_and0 = f_arrdiv32_fs342_not0 & b[22];
  assign f_arrdiv32_fs342_xor1 = f_arrdiv32_fs341_or0 ^ f_arrdiv32_fs342_xor0;
  assign f_arrdiv32_fs342_not1 = ~f_arrdiv32_fs342_xor0;
  assign f_arrdiv32_fs342_and1 = f_arrdiv32_fs342_not1 & f_arrdiv32_fs341_or0;
  assign f_arrdiv32_fs342_or0 = f_arrdiv32_fs342_and1 | f_arrdiv32_fs342_and0;
  assign f_arrdiv32_fs343_xor0 = f_arrdiv32_mux2to1301_xor0 ^ b[23];
  assign f_arrdiv32_fs343_not0 = ~f_arrdiv32_mux2to1301_xor0;
  assign f_arrdiv32_fs343_and0 = f_arrdiv32_fs343_not0 & b[23];
  assign f_arrdiv32_fs343_xor1 = f_arrdiv32_fs342_or0 ^ f_arrdiv32_fs343_xor0;
  assign f_arrdiv32_fs343_not1 = ~f_arrdiv32_fs343_xor0;
  assign f_arrdiv32_fs343_and1 = f_arrdiv32_fs343_not1 & f_arrdiv32_fs342_or0;
  assign f_arrdiv32_fs343_or0 = f_arrdiv32_fs343_and1 | f_arrdiv32_fs343_and0;
  assign f_arrdiv32_fs344_xor0 = f_arrdiv32_mux2to1302_xor0 ^ b[24];
  assign f_arrdiv32_fs344_not0 = ~f_arrdiv32_mux2to1302_xor0;
  assign f_arrdiv32_fs344_and0 = f_arrdiv32_fs344_not0 & b[24];
  assign f_arrdiv32_fs344_xor1 = f_arrdiv32_fs343_or0 ^ f_arrdiv32_fs344_xor0;
  assign f_arrdiv32_fs344_not1 = ~f_arrdiv32_fs344_xor0;
  assign f_arrdiv32_fs344_and1 = f_arrdiv32_fs344_not1 & f_arrdiv32_fs343_or0;
  assign f_arrdiv32_fs344_or0 = f_arrdiv32_fs344_and1 | f_arrdiv32_fs344_and0;
  assign f_arrdiv32_fs345_xor0 = f_arrdiv32_mux2to1303_xor0 ^ b[25];
  assign f_arrdiv32_fs345_not0 = ~f_arrdiv32_mux2to1303_xor0;
  assign f_arrdiv32_fs345_and0 = f_arrdiv32_fs345_not0 & b[25];
  assign f_arrdiv32_fs345_xor1 = f_arrdiv32_fs344_or0 ^ f_arrdiv32_fs345_xor0;
  assign f_arrdiv32_fs345_not1 = ~f_arrdiv32_fs345_xor0;
  assign f_arrdiv32_fs345_and1 = f_arrdiv32_fs345_not1 & f_arrdiv32_fs344_or0;
  assign f_arrdiv32_fs345_or0 = f_arrdiv32_fs345_and1 | f_arrdiv32_fs345_and0;
  assign f_arrdiv32_fs346_xor0 = f_arrdiv32_mux2to1304_xor0 ^ b[26];
  assign f_arrdiv32_fs346_not0 = ~f_arrdiv32_mux2to1304_xor0;
  assign f_arrdiv32_fs346_and0 = f_arrdiv32_fs346_not0 & b[26];
  assign f_arrdiv32_fs346_xor1 = f_arrdiv32_fs345_or0 ^ f_arrdiv32_fs346_xor0;
  assign f_arrdiv32_fs346_not1 = ~f_arrdiv32_fs346_xor0;
  assign f_arrdiv32_fs346_and1 = f_arrdiv32_fs346_not1 & f_arrdiv32_fs345_or0;
  assign f_arrdiv32_fs346_or0 = f_arrdiv32_fs346_and1 | f_arrdiv32_fs346_and0;
  assign f_arrdiv32_fs347_xor0 = f_arrdiv32_mux2to1305_xor0 ^ b[27];
  assign f_arrdiv32_fs347_not0 = ~f_arrdiv32_mux2to1305_xor0;
  assign f_arrdiv32_fs347_and0 = f_arrdiv32_fs347_not0 & b[27];
  assign f_arrdiv32_fs347_xor1 = f_arrdiv32_fs346_or0 ^ f_arrdiv32_fs347_xor0;
  assign f_arrdiv32_fs347_not1 = ~f_arrdiv32_fs347_xor0;
  assign f_arrdiv32_fs347_and1 = f_arrdiv32_fs347_not1 & f_arrdiv32_fs346_or0;
  assign f_arrdiv32_fs347_or0 = f_arrdiv32_fs347_and1 | f_arrdiv32_fs347_and0;
  assign f_arrdiv32_fs348_xor0 = f_arrdiv32_mux2to1306_xor0 ^ b[28];
  assign f_arrdiv32_fs348_not0 = ~f_arrdiv32_mux2to1306_xor0;
  assign f_arrdiv32_fs348_and0 = f_arrdiv32_fs348_not0 & b[28];
  assign f_arrdiv32_fs348_xor1 = f_arrdiv32_fs347_or0 ^ f_arrdiv32_fs348_xor0;
  assign f_arrdiv32_fs348_not1 = ~f_arrdiv32_fs348_xor0;
  assign f_arrdiv32_fs348_and1 = f_arrdiv32_fs348_not1 & f_arrdiv32_fs347_or0;
  assign f_arrdiv32_fs348_or0 = f_arrdiv32_fs348_and1 | f_arrdiv32_fs348_and0;
  assign f_arrdiv32_fs349_xor0 = f_arrdiv32_mux2to1307_xor0 ^ b[29];
  assign f_arrdiv32_fs349_not0 = ~f_arrdiv32_mux2to1307_xor0;
  assign f_arrdiv32_fs349_and0 = f_arrdiv32_fs349_not0 & b[29];
  assign f_arrdiv32_fs349_xor1 = f_arrdiv32_fs348_or0 ^ f_arrdiv32_fs349_xor0;
  assign f_arrdiv32_fs349_not1 = ~f_arrdiv32_fs349_xor0;
  assign f_arrdiv32_fs349_and1 = f_arrdiv32_fs349_not1 & f_arrdiv32_fs348_or0;
  assign f_arrdiv32_fs349_or0 = f_arrdiv32_fs349_and1 | f_arrdiv32_fs349_and0;
  assign f_arrdiv32_fs350_xor0 = f_arrdiv32_mux2to1308_xor0 ^ b[30];
  assign f_arrdiv32_fs350_not0 = ~f_arrdiv32_mux2to1308_xor0;
  assign f_arrdiv32_fs350_and0 = f_arrdiv32_fs350_not0 & b[30];
  assign f_arrdiv32_fs350_xor1 = f_arrdiv32_fs349_or0 ^ f_arrdiv32_fs350_xor0;
  assign f_arrdiv32_fs350_not1 = ~f_arrdiv32_fs350_xor0;
  assign f_arrdiv32_fs350_and1 = f_arrdiv32_fs350_not1 & f_arrdiv32_fs349_or0;
  assign f_arrdiv32_fs350_or0 = f_arrdiv32_fs350_and1 | f_arrdiv32_fs350_and0;
  assign f_arrdiv32_fs351_xor0 = f_arrdiv32_mux2to1309_xor0 ^ b[31];
  assign f_arrdiv32_fs351_not0 = ~f_arrdiv32_mux2to1309_xor0;
  assign f_arrdiv32_fs351_and0 = f_arrdiv32_fs351_not0 & b[31];
  assign f_arrdiv32_fs351_xor1 = f_arrdiv32_fs350_or0 ^ f_arrdiv32_fs351_xor0;
  assign f_arrdiv32_fs351_not1 = ~f_arrdiv32_fs351_xor0;
  assign f_arrdiv32_fs351_and1 = f_arrdiv32_fs351_not1 & f_arrdiv32_fs350_or0;
  assign f_arrdiv32_fs351_or0 = f_arrdiv32_fs351_and1 | f_arrdiv32_fs351_and0;
  assign f_arrdiv32_mux2to1310_and0 = a[21] & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1310_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1310_and1 = f_arrdiv32_fs320_xor0 & f_arrdiv32_mux2to1310_not0;
  assign f_arrdiv32_mux2to1310_xor0 = f_arrdiv32_mux2to1310_and0 ^ f_arrdiv32_mux2to1310_and1;
  assign f_arrdiv32_mux2to1311_and0 = f_arrdiv32_mux2to1279_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1311_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1311_and1 = f_arrdiv32_fs321_xor1 & f_arrdiv32_mux2to1311_not0;
  assign f_arrdiv32_mux2to1311_xor0 = f_arrdiv32_mux2to1311_and0 ^ f_arrdiv32_mux2to1311_and1;
  assign f_arrdiv32_mux2to1312_and0 = f_arrdiv32_mux2to1280_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1312_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1312_and1 = f_arrdiv32_fs322_xor1 & f_arrdiv32_mux2to1312_not0;
  assign f_arrdiv32_mux2to1312_xor0 = f_arrdiv32_mux2to1312_and0 ^ f_arrdiv32_mux2to1312_and1;
  assign f_arrdiv32_mux2to1313_and0 = f_arrdiv32_mux2to1281_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1313_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1313_and1 = f_arrdiv32_fs323_xor1 & f_arrdiv32_mux2to1313_not0;
  assign f_arrdiv32_mux2to1313_xor0 = f_arrdiv32_mux2to1313_and0 ^ f_arrdiv32_mux2to1313_and1;
  assign f_arrdiv32_mux2to1314_and0 = f_arrdiv32_mux2to1282_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1314_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1314_and1 = f_arrdiv32_fs324_xor1 & f_arrdiv32_mux2to1314_not0;
  assign f_arrdiv32_mux2to1314_xor0 = f_arrdiv32_mux2to1314_and0 ^ f_arrdiv32_mux2to1314_and1;
  assign f_arrdiv32_mux2to1315_and0 = f_arrdiv32_mux2to1283_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1315_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1315_and1 = f_arrdiv32_fs325_xor1 & f_arrdiv32_mux2to1315_not0;
  assign f_arrdiv32_mux2to1315_xor0 = f_arrdiv32_mux2to1315_and0 ^ f_arrdiv32_mux2to1315_and1;
  assign f_arrdiv32_mux2to1316_and0 = f_arrdiv32_mux2to1284_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1316_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1316_and1 = f_arrdiv32_fs326_xor1 & f_arrdiv32_mux2to1316_not0;
  assign f_arrdiv32_mux2to1316_xor0 = f_arrdiv32_mux2to1316_and0 ^ f_arrdiv32_mux2to1316_and1;
  assign f_arrdiv32_mux2to1317_and0 = f_arrdiv32_mux2to1285_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1317_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1317_and1 = f_arrdiv32_fs327_xor1 & f_arrdiv32_mux2to1317_not0;
  assign f_arrdiv32_mux2to1317_xor0 = f_arrdiv32_mux2to1317_and0 ^ f_arrdiv32_mux2to1317_and1;
  assign f_arrdiv32_mux2to1318_and0 = f_arrdiv32_mux2to1286_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1318_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1318_and1 = f_arrdiv32_fs328_xor1 & f_arrdiv32_mux2to1318_not0;
  assign f_arrdiv32_mux2to1318_xor0 = f_arrdiv32_mux2to1318_and0 ^ f_arrdiv32_mux2to1318_and1;
  assign f_arrdiv32_mux2to1319_and0 = f_arrdiv32_mux2to1287_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1319_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1319_and1 = f_arrdiv32_fs329_xor1 & f_arrdiv32_mux2to1319_not0;
  assign f_arrdiv32_mux2to1319_xor0 = f_arrdiv32_mux2to1319_and0 ^ f_arrdiv32_mux2to1319_and1;
  assign f_arrdiv32_mux2to1320_and0 = f_arrdiv32_mux2to1288_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1320_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1320_and1 = f_arrdiv32_fs330_xor1 & f_arrdiv32_mux2to1320_not0;
  assign f_arrdiv32_mux2to1320_xor0 = f_arrdiv32_mux2to1320_and0 ^ f_arrdiv32_mux2to1320_and1;
  assign f_arrdiv32_mux2to1321_and0 = f_arrdiv32_mux2to1289_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1321_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1321_and1 = f_arrdiv32_fs331_xor1 & f_arrdiv32_mux2to1321_not0;
  assign f_arrdiv32_mux2to1321_xor0 = f_arrdiv32_mux2to1321_and0 ^ f_arrdiv32_mux2to1321_and1;
  assign f_arrdiv32_mux2to1322_and0 = f_arrdiv32_mux2to1290_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1322_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1322_and1 = f_arrdiv32_fs332_xor1 & f_arrdiv32_mux2to1322_not0;
  assign f_arrdiv32_mux2to1322_xor0 = f_arrdiv32_mux2to1322_and0 ^ f_arrdiv32_mux2to1322_and1;
  assign f_arrdiv32_mux2to1323_and0 = f_arrdiv32_mux2to1291_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1323_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1323_and1 = f_arrdiv32_fs333_xor1 & f_arrdiv32_mux2to1323_not0;
  assign f_arrdiv32_mux2to1323_xor0 = f_arrdiv32_mux2to1323_and0 ^ f_arrdiv32_mux2to1323_and1;
  assign f_arrdiv32_mux2to1324_and0 = f_arrdiv32_mux2to1292_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1324_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1324_and1 = f_arrdiv32_fs334_xor1 & f_arrdiv32_mux2to1324_not0;
  assign f_arrdiv32_mux2to1324_xor0 = f_arrdiv32_mux2to1324_and0 ^ f_arrdiv32_mux2to1324_and1;
  assign f_arrdiv32_mux2to1325_and0 = f_arrdiv32_mux2to1293_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1325_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1325_and1 = f_arrdiv32_fs335_xor1 & f_arrdiv32_mux2to1325_not0;
  assign f_arrdiv32_mux2to1325_xor0 = f_arrdiv32_mux2to1325_and0 ^ f_arrdiv32_mux2to1325_and1;
  assign f_arrdiv32_mux2to1326_and0 = f_arrdiv32_mux2to1294_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1326_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1326_and1 = f_arrdiv32_fs336_xor1 & f_arrdiv32_mux2to1326_not0;
  assign f_arrdiv32_mux2to1326_xor0 = f_arrdiv32_mux2to1326_and0 ^ f_arrdiv32_mux2to1326_and1;
  assign f_arrdiv32_mux2to1327_and0 = f_arrdiv32_mux2to1295_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1327_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1327_and1 = f_arrdiv32_fs337_xor1 & f_arrdiv32_mux2to1327_not0;
  assign f_arrdiv32_mux2to1327_xor0 = f_arrdiv32_mux2to1327_and0 ^ f_arrdiv32_mux2to1327_and1;
  assign f_arrdiv32_mux2to1328_and0 = f_arrdiv32_mux2to1296_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1328_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1328_and1 = f_arrdiv32_fs338_xor1 & f_arrdiv32_mux2to1328_not0;
  assign f_arrdiv32_mux2to1328_xor0 = f_arrdiv32_mux2to1328_and0 ^ f_arrdiv32_mux2to1328_and1;
  assign f_arrdiv32_mux2to1329_and0 = f_arrdiv32_mux2to1297_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1329_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1329_and1 = f_arrdiv32_fs339_xor1 & f_arrdiv32_mux2to1329_not0;
  assign f_arrdiv32_mux2to1329_xor0 = f_arrdiv32_mux2to1329_and0 ^ f_arrdiv32_mux2to1329_and1;
  assign f_arrdiv32_mux2to1330_and0 = f_arrdiv32_mux2to1298_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1330_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1330_and1 = f_arrdiv32_fs340_xor1 & f_arrdiv32_mux2to1330_not0;
  assign f_arrdiv32_mux2to1330_xor0 = f_arrdiv32_mux2to1330_and0 ^ f_arrdiv32_mux2to1330_and1;
  assign f_arrdiv32_mux2to1331_and0 = f_arrdiv32_mux2to1299_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1331_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1331_and1 = f_arrdiv32_fs341_xor1 & f_arrdiv32_mux2to1331_not0;
  assign f_arrdiv32_mux2to1331_xor0 = f_arrdiv32_mux2to1331_and0 ^ f_arrdiv32_mux2to1331_and1;
  assign f_arrdiv32_mux2to1332_and0 = f_arrdiv32_mux2to1300_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1332_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1332_and1 = f_arrdiv32_fs342_xor1 & f_arrdiv32_mux2to1332_not0;
  assign f_arrdiv32_mux2to1332_xor0 = f_arrdiv32_mux2to1332_and0 ^ f_arrdiv32_mux2to1332_and1;
  assign f_arrdiv32_mux2to1333_and0 = f_arrdiv32_mux2to1301_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1333_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1333_and1 = f_arrdiv32_fs343_xor1 & f_arrdiv32_mux2to1333_not0;
  assign f_arrdiv32_mux2to1333_xor0 = f_arrdiv32_mux2to1333_and0 ^ f_arrdiv32_mux2to1333_and1;
  assign f_arrdiv32_mux2to1334_and0 = f_arrdiv32_mux2to1302_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1334_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1334_and1 = f_arrdiv32_fs344_xor1 & f_arrdiv32_mux2to1334_not0;
  assign f_arrdiv32_mux2to1334_xor0 = f_arrdiv32_mux2to1334_and0 ^ f_arrdiv32_mux2to1334_and1;
  assign f_arrdiv32_mux2to1335_and0 = f_arrdiv32_mux2to1303_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1335_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1335_and1 = f_arrdiv32_fs345_xor1 & f_arrdiv32_mux2to1335_not0;
  assign f_arrdiv32_mux2to1335_xor0 = f_arrdiv32_mux2to1335_and0 ^ f_arrdiv32_mux2to1335_and1;
  assign f_arrdiv32_mux2to1336_and0 = f_arrdiv32_mux2to1304_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1336_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1336_and1 = f_arrdiv32_fs346_xor1 & f_arrdiv32_mux2to1336_not0;
  assign f_arrdiv32_mux2to1336_xor0 = f_arrdiv32_mux2to1336_and0 ^ f_arrdiv32_mux2to1336_and1;
  assign f_arrdiv32_mux2to1337_and0 = f_arrdiv32_mux2to1305_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1337_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1337_and1 = f_arrdiv32_fs347_xor1 & f_arrdiv32_mux2to1337_not0;
  assign f_arrdiv32_mux2to1337_xor0 = f_arrdiv32_mux2to1337_and0 ^ f_arrdiv32_mux2to1337_and1;
  assign f_arrdiv32_mux2to1338_and0 = f_arrdiv32_mux2to1306_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1338_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1338_and1 = f_arrdiv32_fs348_xor1 & f_arrdiv32_mux2to1338_not0;
  assign f_arrdiv32_mux2to1338_xor0 = f_arrdiv32_mux2to1338_and0 ^ f_arrdiv32_mux2to1338_and1;
  assign f_arrdiv32_mux2to1339_and0 = f_arrdiv32_mux2to1307_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1339_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1339_and1 = f_arrdiv32_fs349_xor1 & f_arrdiv32_mux2to1339_not0;
  assign f_arrdiv32_mux2to1339_xor0 = f_arrdiv32_mux2to1339_and0 ^ f_arrdiv32_mux2to1339_and1;
  assign f_arrdiv32_mux2to1340_and0 = f_arrdiv32_mux2to1308_xor0 & f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1340_not0 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_mux2to1340_and1 = f_arrdiv32_fs350_xor1 & f_arrdiv32_mux2to1340_not0;
  assign f_arrdiv32_mux2to1340_xor0 = f_arrdiv32_mux2to1340_and0 ^ f_arrdiv32_mux2to1340_and1;
  assign f_arrdiv32_not10 = ~f_arrdiv32_fs351_or0;
  assign f_arrdiv32_fs352_xor0 = a[20] ^ b[0];
  assign f_arrdiv32_fs352_not0 = ~a[20];
  assign f_arrdiv32_fs352_and0 = f_arrdiv32_fs352_not0 & b[0];
  assign f_arrdiv32_fs352_not1 = ~f_arrdiv32_fs352_xor0;
  assign f_arrdiv32_fs353_xor0 = f_arrdiv32_mux2to1310_xor0 ^ b[1];
  assign f_arrdiv32_fs353_not0 = ~f_arrdiv32_mux2to1310_xor0;
  assign f_arrdiv32_fs353_and0 = f_arrdiv32_fs353_not0 & b[1];
  assign f_arrdiv32_fs353_xor1 = f_arrdiv32_fs352_and0 ^ f_arrdiv32_fs353_xor0;
  assign f_arrdiv32_fs353_not1 = ~f_arrdiv32_fs353_xor0;
  assign f_arrdiv32_fs353_and1 = f_arrdiv32_fs353_not1 & f_arrdiv32_fs352_and0;
  assign f_arrdiv32_fs353_or0 = f_arrdiv32_fs353_and1 | f_arrdiv32_fs353_and0;
  assign f_arrdiv32_fs354_xor0 = f_arrdiv32_mux2to1311_xor0 ^ b[2];
  assign f_arrdiv32_fs354_not0 = ~f_arrdiv32_mux2to1311_xor0;
  assign f_arrdiv32_fs354_and0 = f_arrdiv32_fs354_not0 & b[2];
  assign f_arrdiv32_fs354_xor1 = f_arrdiv32_fs353_or0 ^ f_arrdiv32_fs354_xor0;
  assign f_arrdiv32_fs354_not1 = ~f_arrdiv32_fs354_xor0;
  assign f_arrdiv32_fs354_and1 = f_arrdiv32_fs354_not1 & f_arrdiv32_fs353_or0;
  assign f_arrdiv32_fs354_or0 = f_arrdiv32_fs354_and1 | f_arrdiv32_fs354_and0;
  assign f_arrdiv32_fs355_xor0 = f_arrdiv32_mux2to1312_xor0 ^ b[3];
  assign f_arrdiv32_fs355_not0 = ~f_arrdiv32_mux2to1312_xor0;
  assign f_arrdiv32_fs355_and0 = f_arrdiv32_fs355_not0 & b[3];
  assign f_arrdiv32_fs355_xor1 = f_arrdiv32_fs354_or0 ^ f_arrdiv32_fs355_xor0;
  assign f_arrdiv32_fs355_not1 = ~f_arrdiv32_fs355_xor0;
  assign f_arrdiv32_fs355_and1 = f_arrdiv32_fs355_not1 & f_arrdiv32_fs354_or0;
  assign f_arrdiv32_fs355_or0 = f_arrdiv32_fs355_and1 | f_arrdiv32_fs355_and0;
  assign f_arrdiv32_fs356_xor0 = f_arrdiv32_mux2to1313_xor0 ^ b[4];
  assign f_arrdiv32_fs356_not0 = ~f_arrdiv32_mux2to1313_xor0;
  assign f_arrdiv32_fs356_and0 = f_arrdiv32_fs356_not0 & b[4];
  assign f_arrdiv32_fs356_xor1 = f_arrdiv32_fs355_or0 ^ f_arrdiv32_fs356_xor0;
  assign f_arrdiv32_fs356_not1 = ~f_arrdiv32_fs356_xor0;
  assign f_arrdiv32_fs356_and1 = f_arrdiv32_fs356_not1 & f_arrdiv32_fs355_or0;
  assign f_arrdiv32_fs356_or0 = f_arrdiv32_fs356_and1 | f_arrdiv32_fs356_and0;
  assign f_arrdiv32_fs357_xor0 = f_arrdiv32_mux2to1314_xor0 ^ b[5];
  assign f_arrdiv32_fs357_not0 = ~f_arrdiv32_mux2to1314_xor0;
  assign f_arrdiv32_fs357_and0 = f_arrdiv32_fs357_not0 & b[5];
  assign f_arrdiv32_fs357_xor1 = f_arrdiv32_fs356_or0 ^ f_arrdiv32_fs357_xor0;
  assign f_arrdiv32_fs357_not1 = ~f_arrdiv32_fs357_xor0;
  assign f_arrdiv32_fs357_and1 = f_arrdiv32_fs357_not1 & f_arrdiv32_fs356_or0;
  assign f_arrdiv32_fs357_or0 = f_arrdiv32_fs357_and1 | f_arrdiv32_fs357_and0;
  assign f_arrdiv32_fs358_xor0 = f_arrdiv32_mux2to1315_xor0 ^ b[6];
  assign f_arrdiv32_fs358_not0 = ~f_arrdiv32_mux2to1315_xor0;
  assign f_arrdiv32_fs358_and0 = f_arrdiv32_fs358_not0 & b[6];
  assign f_arrdiv32_fs358_xor1 = f_arrdiv32_fs357_or0 ^ f_arrdiv32_fs358_xor0;
  assign f_arrdiv32_fs358_not1 = ~f_arrdiv32_fs358_xor0;
  assign f_arrdiv32_fs358_and1 = f_arrdiv32_fs358_not1 & f_arrdiv32_fs357_or0;
  assign f_arrdiv32_fs358_or0 = f_arrdiv32_fs358_and1 | f_arrdiv32_fs358_and0;
  assign f_arrdiv32_fs359_xor0 = f_arrdiv32_mux2to1316_xor0 ^ b[7];
  assign f_arrdiv32_fs359_not0 = ~f_arrdiv32_mux2to1316_xor0;
  assign f_arrdiv32_fs359_and0 = f_arrdiv32_fs359_not0 & b[7];
  assign f_arrdiv32_fs359_xor1 = f_arrdiv32_fs358_or0 ^ f_arrdiv32_fs359_xor0;
  assign f_arrdiv32_fs359_not1 = ~f_arrdiv32_fs359_xor0;
  assign f_arrdiv32_fs359_and1 = f_arrdiv32_fs359_not1 & f_arrdiv32_fs358_or0;
  assign f_arrdiv32_fs359_or0 = f_arrdiv32_fs359_and1 | f_arrdiv32_fs359_and0;
  assign f_arrdiv32_fs360_xor0 = f_arrdiv32_mux2to1317_xor0 ^ b[8];
  assign f_arrdiv32_fs360_not0 = ~f_arrdiv32_mux2to1317_xor0;
  assign f_arrdiv32_fs360_and0 = f_arrdiv32_fs360_not0 & b[8];
  assign f_arrdiv32_fs360_xor1 = f_arrdiv32_fs359_or0 ^ f_arrdiv32_fs360_xor0;
  assign f_arrdiv32_fs360_not1 = ~f_arrdiv32_fs360_xor0;
  assign f_arrdiv32_fs360_and1 = f_arrdiv32_fs360_not1 & f_arrdiv32_fs359_or0;
  assign f_arrdiv32_fs360_or0 = f_arrdiv32_fs360_and1 | f_arrdiv32_fs360_and0;
  assign f_arrdiv32_fs361_xor0 = f_arrdiv32_mux2to1318_xor0 ^ b[9];
  assign f_arrdiv32_fs361_not0 = ~f_arrdiv32_mux2to1318_xor0;
  assign f_arrdiv32_fs361_and0 = f_arrdiv32_fs361_not0 & b[9];
  assign f_arrdiv32_fs361_xor1 = f_arrdiv32_fs360_or0 ^ f_arrdiv32_fs361_xor0;
  assign f_arrdiv32_fs361_not1 = ~f_arrdiv32_fs361_xor0;
  assign f_arrdiv32_fs361_and1 = f_arrdiv32_fs361_not1 & f_arrdiv32_fs360_or0;
  assign f_arrdiv32_fs361_or0 = f_arrdiv32_fs361_and1 | f_arrdiv32_fs361_and0;
  assign f_arrdiv32_fs362_xor0 = f_arrdiv32_mux2to1319_xor0 ^ b[10];
  assign f_arrdiv32_fs362_not0 = ~f_arrdiv32_mux2to1319_xor0;
  assign f_arrdiv32_fs362_and0 = f_arrdiv32_fs362_not0 & b[10];
  assign f_arrdiv32_fs362_xor1 = f_arrdiv32_fs361_or0 ^ f_arrdiv32_fs362_xor0;
  assign f_arrdiv32_fs362_not1 = ~f_arrdiv32_fs362_xor0;
  assign f_arrdiv32_fs362_and1 = f_arrdiv32_fs362_not1 & f_arrdiv32_fs361_or0;
  assign f_arrdiv32_fs362_or0 = f_arrdiv32_fs362_and1 | f_arrdiv32_fs362_and0;
  assign f_arrdiv32_fs363_xor0 = f_arrdiv32_mux2to1320_xor0 ^ b[11];
  assign f_arrdiv32_fs363_not0 = ~f_arrdiv32_mux2to1320_xor0;
  assign f_arrdiv32_fs363_and0 = f_arrdiv32_fs363_not0 & b[11];
  assign f_arrdiv32_fs363_xor1 = f_arrdiv32_fs362_or0 ^ f_arrdiv32_fs363_xor0;
  assign f_arrdiv32_fs363_not1 = ~f_arrdiv32_fs363_xor0;
  assign f_arrdiv32_fs363_and1 = f_arrdiv32_fs363_not1 & f_arrdiv32_fs362_or0;
  assign f_arrdiv32_fs363_or0 = f_arrdiv32_fs363_and1 | f_arrdiv32_fs363_and0;
  assign f_arrdiv32_fs364_xor0 = f_arrdiv32_mux2to1321_xor0 ^ b[12];
  assign f_arrdiv32_fs364_not0 = ~f_arrdiv32_mux2to1321_xor0;
  assign f_arrdiv32_fs364_and0 = f_arrdiv32_fs364_not0 & b[12];
  assign f_arrdiv32_fs364_xor1 = f_arrdiv32_fs363_or0 ^ f_arrdiv32_fs364_xor0;
  assign f_arrdiv32_fs364_not1 = ~f_arrdiv32_fs364_xor0;
  assign f_arrdiv32_fs364_and1 = f_arrdiv32_fs364_not1 & f_arrdiv32_fs363_or0;
  assign f_arrdiv32_fs364_or0 = f_arrdiv32_fs364_and1 | f_arrdiv32_fs364_and0;
  assign f_arrdiv32_fs365_xor0 = f_arrdiv32_mux2to1322_xor0 ^ b[13];
  assign f_arrdiv32_fs365_not0 = ~f_arrdiv32_mux2to1322_xor0;
  assign f_arrdiv32_fs365_and0 = f_arrdiv32_fs365_not0 & b[13];
  assign f_arrdiv32_fs365_xor1 = f_arrdiv32_fs364_or0 ^ f_arrdiv32_fs365_xor0;
  assign f_arrdiv32_fs365_not1 = ~f_arrdiv32_fs365_xor0;
  assign f_arrdiv32_fs365_and1 = f_arrdiv32_fs365_not1 & f_arrdiv32_fs364_or0;
  assign f_arrdiv32_fs365_or0 = f_arrdiv32_fs365_and1 | f_arrdiv32_fs365_and0;
  assign f_arrdiv32_fs366_xor0 = f_arrdiv32_mux2to1323_xor0 ^ b[14];
  assign f_arrdiv32_fs366_not0 = ~f_arrdiv32_mux2to1323_xor0;
  assign f_arrdiv32_fs366_and0 = f_arrdiv32_fs366_not0 & b[14];
  assign f_arrdiv32_fs366_xor1 = f_arrdiv32_fs365_or0 ^ f_arrdiv32_fs366_xor0;
  assign f_arrdiv32_fs366_not1 = ~f_arrdiv32_fs366_xor0;
  assign f_arrdiv32_fs366_and1 = f_arrdiv32_fs366_not1 & f_arrdiv32_fs365_or0;
  assign f_arrdiv32_fs366_or0 = f_arrdiv32_fs366_and1 | f_arrdiv32_fs366_and0;
  assign f_arrdiv32_fs367_xor0 = f_arrdiv32_mux2to1324_xor0 ^ b[15];
  assign f_arrdiv32_fs367_not0 = ~f_arrdiv32_mux2to1324_xor0;
  assign f_arrdiv32_fs367_and0 = f_arrdiv32_fs367_not0 & b[15];
  assign f_arrdiv32_fs367_xor1 = f_arrdiv32_fs366_or0 ^ f_arrdiv32_fs367_xor0;
  assign f_arrdiv32_fs367_not1 = ~f_arrdiv32_fs367_xor0;
  assign f_arrdiv32_fs367_and1 = f_arrdiv32_fs367_not1 & f_arrdiv32_fs366_or0;
  assign f_arrdiv32_fs367_or0 = f_arrdiv32_fs367_and1 | f_arrdiv32_fs367_and0;
  assign f_arrdiv32_fs368_xor0 = f_arrdiv32_mux2to1325_xor0 ^ b[16];
  assign f_arrdiv32_fs368_not0 = ~f_arrdiv32_mux2to1325_xor0;
  assign f_arrdiv32_fs368_and0 = f_arrdiv32_fs368_not0 & b[16];
  assign f_arrdiv32_fs368_xor1 = f_arrdiv32_fs367_or0 ^ f_arrdiv32_fs368_xor0;
  assign f_arrdiv32_fs368_not1 = ~f_arrdiv32_fs368_xor0;
  assign f_arrdiv32_fs368_and1 = f_arrdiv32_fs368_not1 & f_arrdiv32_fs367_or0;
  assign f_arrdiv32_fs368_or0 = f_arrdiv32_fs368_and1 | f_arrdiv32_fs368_and0;
  assign f_arrdiv32_fs369_xor0 = f_arrdiv32_mux2to1326_xor0 ^ b[17];
  assign f_arrdiv32_fs369_not0 = ~f_arrdiv32_mux2to1326_xor0;
  assign f_arrdiv32_fs369_and0 = f_arrdiv32_fs369_not0 & b[17];
  assign f_arrdiv32_fs369_xor1 = f_arrdiv32_fs368_or0 ^ f_arrdiv32_fs369_xor0;
  assign f_arrdiv32_fs369_not1 = ~f_arrdiv32_fs369_xor0;
  assign f_arrdiv32_fs369_and1 = f_arrdiv32_fs369_not1 & f_arrdiv32_fs368_or0;
  assign f_arrdiv32_fs369_or0 = f_arrdiv32_fs369_and1 | f_arrdiv32_fs369_and0;
  assign f_arrdiv32_fs370_xor0 = f_arrdiv32_mux2to1327_xor0 ^ b[18];
  assign f_arrdiv32_fs370_not0 = ~f_arrdiv32_mux2to1327_xor0;
  assign f_arrdiv32_fs370_and0 = f_arrdiv32_fs370_not0 & b[18];
  assign f_arrdiv32_fs370_xor1 = f_arrdiv32_fs369_or0 ^ f_arrdiv32_fs370_xor0;
  assign f_arrdiv32_fs370_not1 = ~f_arrdiv32_fs370_xor0;
  assign f_arrdiv32_fs370_and1 = f_arrdiv32_fs370_not1 & f_arrdiv32_fs369_or0;
  assign f_arrdiv32_fs370_or0 = f_arrdiv32_fs370_and1 | f_arrdiv32_fs370_and0;
  assign f_arrdiv32_fs371_xor0 = f_arrdiv32_mux2to1328_xor0 ^ b[19];
  assign f_arrdiv32_fs371_not0 = ~f_arrdiv32_mux2to1328_xor0;
  assign f_arrdiv32_fs371_and0 = f_arrdiv32_fs371_not0 & b[19];
  assign f_arrdiv32_fs371_xor1 = f_arrdiv32_fs370_or0 ^ f_arrdiv32_fs371_xor0;
  assign f_arrdiv32_fs371_not1 = ~f_arrdiv32_fs371_xor0;
  assign f_arrdiv32_fs371_and1 = f_arrdiv32_fs371_not1 & f_arrdiv32_fs370_or0;
  assign f_arrdiv32_fs371_or0 = f_arrdiv32_fs371_and1 | f_arrdiv32_fs371_and0;
  assign f_arrdiv32_fs372_xor0 = f_arrdiv32_mux2to1329_xor0 ^ b[20];
  assign f_arrdiv32_fs372_not0 = ~f_arrdiv32_mux2to1329_xor0;
  assign f_arrdiv32_fs372_and0 = f_arrdiv32_fs372_not0 & b[20];
  assign f_arrdiv32_fs372_xor1 = f_arrdiv32_fs371_or0 ^ f_arrdiv32_fs372_xor0;
  assign f_arrdiv32_fs372_not1 = ~f_arrdiv32_fs372_xor0;
  assign f_arrdiv32_fs372_and1 = f_arrdiv32_fs372_not1 & f_arrdiv32_fs371_or0;
  assign f_arrdiv32_fs372_or0 = f_arrdiv32_fs372_and1 | f_arrdiv32_fs372_and0;
  assign f_arrdiv32_fs373_xor0 = f_arrdiv32_mux2to1330_xor0 ^ b[21];
  assign f_arrdiv32_fs373_not0 = ~f_arrdiv32_mux2to1330_xor0;
  assign f_arrdiv32_fs373_and0 = f_arrdiv32_fs373_not0 & b[21];
  assign f_arrdiv32_fs373_xor1 = f_arrdiv32_fs372_or0 ^ f_arrdiv32_fs373_xor0;
  assign f_arrdiv32_fs373_not1 = ~f_arrdiv32_fs373_xor0;
  assign f_arrdiv32_fs373_and1 = f_arrdiv32_fs373_not1 & f_arrdiv32_fs372_or0;
  assign f_arrdiv32_fs373_or0 = f_arrdiv32_fs373_and1 | f_arrdiv32_fs373_and0;
  assign f_arrdiv32_fs374_xor0 = f_arrdiv32_mux2to1331_xor0 ^ b[22];
  assign f_arrdiv32_fs374_not0 = ~f_arrdiv32_mux2to1331_xor0;
  assign f_arrdiv32_fs374_and0 = f_arrdiv32_fs374_not0 & b[22];
  assign f_arrdiv32_fs374_xor1 = f_arrdiv32_fs373_or0 ^ f_arrdiv32_fs374_xor0;
  assign f_arrdiv32_fs374_not1 = ~f_arrdiv32_fs374_xor0;
  assign f_arrdiv32_fs374_and1 = f_arrdiv32_fs374_not1 & f_arrdiv32_fs373_or0;
  assign f_arrdiv32_fs374_or0 = f_arrdiv32_fs374_and1 | f_arrdiv32_fs374_and0;
  assign f_arrdiv32_fs375_xor0 = f_arrdiv32_mux2to1332_xor0 ^ b[23];
  assign f_arrdiv32_fs375_not0 = ~f_arrdiv32_mux2to1332_xor0;
  assign f_arrdiv32_fs375_and0 = f_arrdiv32_fs375_not0 & b[23];
  assign f_arrdiv32_fs375_xor1 = f_arrdiv32_fs374_or0 ^ f_arrdiv32_fs375_xor0;
  assign f_arrdiv32_fs375_not1 = ~f_arrdiv32_fs375_xor0;
  assign f_arrdiv32_fs375_and1 = f_arrdiv32_fs375_not1 & f_arrdiv32_fs374_or0;
  assign f_arrdiv32_fs375_or0 = f_arrdiv32_fs375_and1 | f_arrdiv32_fs375_and0;
  assign f_arrdiv32_fs376_xor0 = f_arrdiv32_mux2to1333_xor0 ^ b[24];
  assign f_arrdiv32_fs376_not0 = ~f_arrdiv32_mux2to1333_xor0;
  assign f_arrdiv32_fs376_and0 = f_arrdiv32_fs376_not0 & b[24];
  assign f_arrdiv32_fs376_xor1 = f_arrdiv32_fs375_or0 ^ f_arrdiv32_fs376_xor0;
  assign f_arrdiv32_fs376_not1 = ~f_arrdiv32_fs376_xor0;
  assign f_arrdiv32_fs376_and1 = f_arrdiv32_fs376_not1 & f_arrdiv32_fs375_or0;
  assign f_arrdiv32_fs376_or0 = f_arrdiv32_fs376_and1 | f_arrdiv32_fs376_and0;
  assign f_arrdiv32_fs377_xor0 = f_arrdiv32_mux2to1334_xor0 ^ b[25];
  assign f_arrdiv32_fs377_not0 = ~f_arrdiv32_mux2to1334_xor0;
  assign f_arrdiv32_fs377_and0 = f_arrdiv32_fs377_not0 & b[25];
  assign f_arrdiv32_fs377_xor1 = f_arrdiv32_fs376_or0 ^ f_arrdiv32_fs377_xor0;
  assign f_arrdiv32_fs377_not1 = ~f_arrdiv32_fs377_xor0;
  assign f_arrdiv32_fs377_and1 = f_arrdiv32_fs377_not1 & f_arrdiv32_fs376_or0;
  assign f_arrdiv32_fs377_or0 = f_arrdiv32_fs377_and1 | f_arrdiv32_fs377_and0;
  assign f_arrdiv32_fs378_xor0 = f_arrdiv32_mux2to1335_xor0 ^ b[26];
  assign f_arrdiv32_fs378_not0 = ~f_arrdiv32_mux2to1335_xor0;
  assign f_arrdiv32_fs378_and0 = f_arrdiv32_fs378_not0 & b[26];
  assign f_arrdiv32_fs378_xor1 = f_arrdiv32_fs377_or0 ^ f_arrdiv32_fs378_xor0;
  assign f_arrdiv32_fs378_not1 = ~f_arrdiv32_fs378_xor0;
  assign f_arrdiv32_fs378_and1 = f_arrdiv32_fs378_not1 & f_arrdiv32_fs377_or0;
  assign f_arrdiv32_fs378_or0 = f_arrdiv32_fs378_and1 | f_arrdiv32_fs378_and0;
  assign f_arrdiv32_fs379_xor0 = f_arrdiv32_mux2to1336_xor0 ^ b[27];
  assign f_arrdiv32_fs379_not0 = ~f_arrdiv32_mux2to1336_xor0;
  assign f_arrdiv32_fs379_and0 = f_arrdiv32_fs379_not0 & b[27];
  assign f_arrdiv32_fs379_xor1 = f_arrdiv32_fs378_or0 ^ f_arrdiv32_fs379_xor0;
  assign f_arrdiv32_fs379_not1 = ~f_arrdiv32_fs379_xor0;
  assign f_arrdiv32_fs379_and1 = f_arrdiv32_fs379_not1 & f_arrdiv32_fs378_or0;
  assign f_arrdiv32_fs379_or0 = f_arrdiv32_fs379_and1 | f_arrdiv32_fs379_and0;
  assign f_arrdiv32_fs380_xor0 = f_arrdiv32_mux2to1337_xor0 ^ b[28];
  assign f_arrdiv32_fs380_not0 = ~f_arrdiv32_mux2to1337_xor0;
  assign f_arrdiv32_fs380_and0 = f_arrdiv32_fs380_not0 & b[28];
  assign f_arrdiv32_fs380_xor1 = f_arrdiv32_fs379_or0 ^ f_arrdiv32_fs380_xor0;
  assign f_arrdiv32_fs380_not1 = ~f_arrdiv32_fs380_xor0;
  assign f_arrdiv32_fs380_and1 = f_arrdiv32_fs380_not1 & f_arrdiv32_fs379_or0;
  assign f_arrdiv32_fs380_or0 = f_arrdiv32_fs380_and1 | f_arrdiv32_fs380_and0;
  assign f_arrdiv32_fs381_xor0 = f_arrdiv32_mux2to1338_xor0 ^ b[29];
  assign f_arrdiv32_fs381_not0 = ~f_arrdiv32_mux2to1338_xor0;
  assign f_arrdiv32_fs381_and0 = f_arrdiv32_fs381_not0 & b[29];
  assign f_arrdiv32_fs381_xor1 = f_arrdiv32_fs380_or0 ^ f_arrdiv32_fs381_xor0;
  assign f_arrdiv32_fs381_not1 = ~f_arrdiv32_fs381_xor0;
  assign f_arrdiv32_fs381_and1 = f_arrdiv32_fs381_not1 & f_arrdiv32_fs380_or0;
  assign f_arrdiv32_fs381_or0 = f_arrdiv32_fs381_and1 | f_arrdiv32_fs381_and0;
  assign f_arrdiv32_fs382_xor0 = f_arrdiv32_mux2to1339_xor0 ^ b[30];
  assign f_arrdiv32_fs382_not0 = ~f_arrdiv32_mux2to1339_xor0;
  assign f_arrdiv32_fs382_and0 = f_arrdiv32_fs382_not0 & b[30];
  assign f_arrdiv32_fs382_xor1 = f_arrdiv32_fs381_or0 ^ f_arrdiv32_fs382_xor0;
  assign f_arrdiv32_fs382_not1 = ~f_arrdiv32_fs382_xor0;
  assign f_arrdiv32_fs382_and1 = f_arrdiv32_fs382_not1 & f_arrdiv32_fs381_or0;
  assign f_arrdiv32_fs382_or0 = f_arrdiv32_fs382_and1 | f_arrdiv32_fs382_and0;
  assign f_arrdiv32_fs383_xor0 = f_arrdiv32_mux2to1340_xor0 ^ b[31];
  assign f_arrdiv32_fs383_not0 = ~f_arrdiv32_mux2to1340_xor0;
  assign f_arrdiv32_fs383_and0 = f_arrdiv32_fs383_not0 & b[31];
  assign f_arrdiv32_fs383_xor1 = f_arrdiv32_fs382_or0 ^ f_arrdiv32_fs383_xor0;
  assign f_arrdiv32_fs383_not1 = ~f_arrdiv32_fs383_xor0;
  assign f_arrdiv32_fs383_and1 = f_arrdiv32_fs383_not1 & f_arrdiv32_fs382_or0;
  assign f_arrdiv32_fs383_or0 = f_arrdiv32_fs383_and1 | f_arrdiv32_fs383_and0;
  assign f_arrdiv32_mux2to1341_and0 = a[20] & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1341_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1341_and1 = f_arrdiv32_fs352_xor0 & f_arrdiv32_mux2to1341_not0;
  assign f_arrdiv32_mux2to1341_xor0 = f_arrdiv32_mux2to1341_and0 ^ f_arrdiv32_mux2to1341_and1;
  assign f_arrdiv32_mux2to1342_and0 = f_arrdiv32_mux2to1310_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1342_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1342_and1 = f_arrdiv32_fs353_xor1 & f_arrdiv32_mux2to1342_not0;
  assign f_arrdiv32_mux2to1342_xor0 = f_arrdiv32_mux2to1342_and0 ^ f_arrdiv32_mux2to1342_and1;
  assign f_arrdiv32_mux2to1343_and0 = f_arrdiv32_mux2to1311_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1343_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1343_and1 = f_arrdiv32_fs354_xor1 & f_arrdiv32_mux2to1343_not0;
  assign f_arrdiv32_mux2to1343_xor0 = f_arrdiv32_mux2to1343_and0 ^ f_arrdiv32_mux2to1343_and1;
  assign f_arrdiv32_mux2to1344_and0 = f_arrdiv32_mux2to1312_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1344_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1344_and1 = f_arrdiv32_fs355_xor1 & f_arrdiv32_mux2to1344_not0;
  assign f_arrdiv32_mux2to1344_xor0 = f_arrdiv32_mux2to1344_and0 ^ f_arrdiv32_mux2to1344_and1;
  assign f_arrdiv32_mux2to1345_and0 = f_arrdiv32_mux2to1313_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1345_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1345_and1 = f_arrdiv32_fs356_xor1 & f_arrdiv32_mux2to1345_not0;
  assign f_arrdiv32_mux2to1345_xor0 = f_arrdiv32_mux2to1345_and0 ^ f_arrdiv32_mux2to1345_and1;
  assign f_arrdiv32_mux2to1346_and0 = f_arrdiv32_mux2to1314_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1346_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1346_and1 = f_arrdiv32_fs357_xor1 & f_arrdiv32_mux2to1346_not0;
  assign f_arrdiv32_mux2to1346_xor0 = f_arrdiv32_mux2to1346_and0 ^ f_arrdiv32_mux2to1346_and1;
  assign f_arrdiv32_mux2to1347_and0 = f_arrdiv32_mux2to1315_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1347_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1347_and1 = f_arrdiv32_fs358_xor1 & f_arrdiv32_mux2to1347_not0;
  assign f_arrdiv32_mux2to1347_xor0 = f_arrdiv32_mux2to1347_and0 ^ f_arrdiv32_mux2to1347_and1;
  assign f_arrdiv32_mux2to1348_and0 = f_arrdiv32_mux2to1316_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1348_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1348_and1 = f_arrdiv32_fs359_xor1 & f_arrdiv32_mux2to1348_not0;
  assign f_arrdiv32_mux2to1348_xor0 = f_arrdiv32_mux2to1348_and0 ^ f_arrdiv32_mux2to1348_and1;
  assign f_arrdiv32_mux2to1349_and0 = f_arrdiv32_mux2to1317_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1349_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1349_and1 = f_arrdiv32_fs360_xor1 & f_arrdiv32_mux2to1349_not0;
  assign f_arrdiv32_mux2to1349_xor0 = f_arrdiv32_mux2to1349_and0 ^ f_arrdiv32_mux2to1349_and1;
  assign f_arrdiv32_mux2to1350_and0 = f_arrdiv32_mux2to1318_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1350_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1350_and1 = f_arrdiv32_fs361_xor1 & f_arrdiv32_mux2to1350_not0;
  assign f_arrdiv32_mux2to1350_xor0 = f_arrdiv32_mux2to1350_and0 ^ f_arrdiv32_mux2to1350_and1;
  assign f_arrdiv32_mux2to1351_and0 = f_arrdiv32_mux2to1319_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1351_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1351_and1 = f_arrdiv32_fs362_xor1 & f_arrdiv32_mux2to1351_not0;
  assign f_arrdiv32_mux2to1351_xor0 = f_arrdiv32_mux2to1351_and0 ^ f_arrdiv32_mux2to1351_and1;
  assign f_arrdiv32_mux2to1352_and0 = f_arrdiv32_mux2to1320_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1352_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1352_and1 = f_arrdiv32_fs363_xor1 & f_arrdiv32_mux2to1352_not0;
  assign f_arrdiv32_mux2to1352_xor0 = f_arrdiv32_mux2to1352_and0 ^ f_arrdiv32_mux2to1352_and1;
  assign f_arrdiv32_mux2to1353_and0 = f_arrdiv32_mux2to1321_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1353_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1353_and1 = f_arrdiv32_fs364_xor1 & f_arrdiv32_mux2to1353_not0;
  assign f_arrdiv32_mux2to1353_xor0 = f_arrdiv32_mux2to1353_and0 ^ f_arrdiv32_mux2to1353_and1;
  assign f_arrdiv32_mux2to1354_and0 = f_arrdiv32_mux2to1322_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1354_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1354_and1 = f_arrdiv32_fs365_xor1 & f_arrdiv32_mux2to1354_not0;
  assign f_arrdiv32_mux2to1354_xor0 = f_arrdiv32_mux2to1354_and0 ^ f_arrdiv32_mux2to1354_and1;
  assign f_arrdiv32_mux2to1355_and0 = f_arrdiv32_mux2to1323_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1355_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1355_and1 = f_arrdiv32_fs366_xor1 & f_arrdiv32_mux2to1355_not0;
  assign f_arrdiv32_mux2to1355_xor0 = f_arrdiv32_mux2to1355_and0 ^ f_arrdiv32_mux2to1355_and1;
  assign f_arrdiv32_mux2to1356_and0 = f_arrdiv32_mux2to1324_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1356_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1356_and1 = f_arrdiv32_fs367_xor1 & f_arrdiv32_mux2to1356_not0;
  assign f_arrdiv32_mux2to1356_xor0 = f_arrdiv32_mux2to1356_and0 ^ f_arrdiv32_mux2to1356_and1;
  assign f_arrdiv32_mux2to1357_and0 = f_arrdiv32_mux2to1325_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1357_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1357_and1 = f_arrdiv32_fs368_xor1 & f_arrdiv32_mux2to1357_not0;
  assign f_arrdiv32_mux2to1357_xor0 = f_arrdiv32_mux2to1357_and0 ^ f_arrdiv32_mux2to1357_and1;
  assign f_arrdiv32_mux2to1358_and0 = f_arrdiv32_mux2to1326_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1358_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1358_and1 = f_arrdiv32_fs369_xor1 & f_arrdiv32_mux2to1358_not0;
  assign f_arrdiv32_mux2to1358_xor0 = f_arrdiv32_mux2to1358_and0 ^ f_arrdiv32_mux2to1358_and1;
  assign f_arrdiv32_mux2to1359_and0 = f_arrdiv32_mux2to1327_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1359_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1359_and1 = f_arrdiv32_fs370_xor1 & f_arrdiv32_mux2to1359_not0;
  assign f_arrdiv32_mux2to1359_xor0 = f_arrdiv32_mux2to1359_and0 ^ f_arrdiv32_mux2to1359_and1;
  assign f_arrdiv32_mux2to1360_and0 = f_arrdiv32_mux2to1328_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1360_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1360_and1 = f_arrdiv32_fs371_xor1 & f_arrdiv32_mux2to1360_not0;
  assign f_arrdiv32_mux2to1360_xor0 = f_arrdiv32_mux2to1360_and0 ^ f_arrdiv32_mux2to1360_and1;
  assign f_arrdiv32_mux2to1361_and0 = f_arrdiv32_mux2to1329_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1361_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1361_and1 = f_arrdiv32_fs372_xor1 & f_arrdiv32_mux2to1361_not0;
  assign f_arrdiv32_mux2to1361_xor0 = f_arrdiv32_mux2to1361_and0 ^ f_arrdiv32_mux2to1361_and1;
  assign f_arrdiv32_mux2to1362_and0 = f_arrdiv32_mux2to1330_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1362_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1362_and1 = f_arrdiv32_fs373_xor1 & f_arrdiv32_mux2to1362_not0;
  assign f_arrdiv32_mux2to1362_xor0 = f_arrdiv32_mux2to1362_and0 ^ f_arrdiv32_mux2to1362_and1;
  assign f_arrdiv32_mux2to1363_and0 = f_arrdiv32_mux2to1331_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1363_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1363_and1 = f_arrdiv32_fs374_xor1 & f_arrdiv32_mux2to1363_not0;
  assign f_arrdiv32_mux2to1363_xor0 = f_arrdiv32_mux2to1363_and0 ^ f_arrdiv32_mux2to1363_and1;
  assign f_arrdiv32_mux2to1364_and0 = f_arrdiv32_mux2to1332_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1364_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1364_and1 = f_arrdiv32_fs375_xor1 & f_arrdiv32_mux2to1364_not0;
  assign f_arrdiv32_mux2to1364_xor0 = f_arrdiv32_mux2to1364_and0 ^ f_arrdiv32_mux2to1364_and1;
  assign f_arrdiv32_mux2to1365_and0 = f_arrdiv32_mux2to1333_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1365_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1365_and1 = f_arrdiv32_fs376_xor1 & f_arrdiv32_mux2to1365_not0;
  assign f_arrdiv32_mux2to1365_xor0 = f_arrdiv32_mux2to1365_and0 ^ f_arrdiv32_mux2to1365_and1;
  assign f_arrdiv32_mux2to1366_and0 = f_arrdiv32_mux2to1334_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1366_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1366_and1 = f_arrdiv32_fs377_xor1 & f_arrdiv32_mux2to1366_not0;
  assign f_arrdiv32_mux2to1366_xor0 = f_arrdiv32_mux2to1366_and0 ^ f_arrdiv32_mux2to1366_and1;
  assign f_arrdiv32_mux2to1367_and0 = f_arrdiv32_mux2to1335_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1367_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1367_and1 = f_arrdiv32_fs378_xor1 & f_arrdiv32_mux2to1367_not0;
  assign f_arrdiv32_mux2to1367_xor0 = f_arrdiv32_mux2to1367_and0 ^ f_arrdiv32_mux2to1367_and1;
  assign f_arrdiv32_mux2to1368_and0 = f_arrdiv32_mux2to1336_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1368_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1368_and1 = f_arrdiv32_fs379_xor1 & f_arrdiv32_mux2to1368_not0;
  assign f_arrdiv32_mux2to1368_xor0 = f_arrdiv32_mux2to1368_and0 ^ f_arrdiv32_mux2to1368_and1;
  assign f_arrdiv32_mux2to1369_and0 = f_arrdiv32_mux2to1337_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1369_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1369_and1 = f_arrdiv32_fs380_xor1 & f_arrdiv32_mux2to1369_not0;
  assign f_arrdiv32_mux2to1369_xor0 = f_arrdiv32_mux2to1369_and0 ^ f_arrdiv32_mux2to1369_and1;
  assign f_arrdiv32_mux2to1370_and0 = f_arrdiv32_mux2to1338_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1370_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1370_and1 = f_arrdiv32_fs381_xor1 & f_arrdiv32_mux2to1370_not0;
  assign f_arrdiv32_mux2to1370_xor0 = f_arrdiv32_mux2to1370_and0 ^ f_arrdiv32_mux2to1370_and1;
  assign f_arrdiv32_mux2to1371_and0 = f_arrdiv32_mux2to1339_xor0 & f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1371_not0 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_mux2to1371_and1 = f_arrdiv32_fs382_xor1 & f_arrdiv32_mux2to1371_not0;
  assign f_arrdiv32_mux2to1371_xor0 = f_arrdiv32_mux2to1371_and0 ^ f_arrdiv32_mux2to1371_and1;
  assign f_arrdiv32_not11 = ~f_arrdiv32_fs383_or0;
  assign f_arrdiv32_fs384_xor0 = a[19] ^ b[0];
  assign f_arrdiv32_fs384_not0 = ~a[19];
  assign f_arrdiv32_fs384_and0 = f_arrdiv32_fs384_not0 & b[0];
  assign f_arrdiv32_fs384_not1 = ~f_arrdiv32_fs384_xor0;
  assign f_arrdiv32_fs385_xor0 = f_arrdiv32_mux2to1341_xor0 ^ b[1];
  assign f_arrdiv32_fs385_not0 = ~f_arrdiv32_mux2to1341_xor0;
  assign f_arrdiv32_fs385_and0 = f_arrdiv32_fs385_not0 & b[1];
  assign f_arrdiv32_fs385_xor1 = f_arrdiv32_fs384_and0 ^ f_arrdiv32_fs385_xor0;
  assign f_arrdiv32_fs385_not1 = ~f_arrdiv32_fs385_xor0;
  assign f_arrdiv32_fs385_and1 = f_arrdiv32_fs385_not1 & f_arrdiv32_fs384_and0;
  assign f_arrdiv32_fs385_or0 = f_arrdiv32_fs385_and1 | f_arrdiv32_fs385_and0;
  assign f_arrdiv32_fs386_xor0 = f_arrdiv32_mux2to1342_xor0 ^ b[2];
  assign f_arrdiv32_fs386_not0 = ~f_arrdiv32_mux2to1342_xor0;
  assign f_arrdiv32_fs386_and0 = f_arrdiv32_fs386_not0 & b[2];
  assign f_arrdiv32_fs386_xor1 = f_arrdiv32_fs385_or0 ^ f_arrdiv32_fs386_xor0;
  assign f_arrdiv32_fs386_not1 = ~f_arrdiv32_fs386_xor0;
  assign f_arrdiv32_fs386_and1 = f_arrdiv32_fs386_not1 & f_arrdiv32_fs385_or0;
  assign f_arrdiv32_fs386_or0 = f_arrdiv32_fs386_and1 | f_arrdiv32_fs386_and0;
  assign f_arrdiv32_fs387_xor0 = f_arrdiv32_mux2to1343_xor0 ^ b[3];
  assign f_arrdiv32_fs387_not0 = ~f_arrdiv32_mux2to1343_xor0;
  assign f_arrdiv32_fs387_and0 = f_arrdiv32_fs387_not0 & b[3];
  assign f_arrdiv32_fs387_xor1 = f_arrdiv32_fs386_or0 ^ f_arrdiv32_fs387_xor0;
  assign f_arrdiv32_fs387_not1 = ~f_arrdiv32_fs387_xor0;
  assign f_arrdiv32_fs387_and1 = f_arrdiv32_fs387_not1 & f_arrdiv32_fs386_or0;
  assign f_arrdiv32_fs387_or0 = f_arrdiv32_fs387_and1 | f_arrdiv32_fs387_and0;
  assign f_arrdiv32_fs388_xor0 = f_arrdiv32_mux2to1344_xor0 ^ b[4];
  assign f_arrdiv32_fs388_not0 = ~f_arrdiv32_mux2to1344_xor0;
  assign f_arrdiv32_fs388_and0 = f_arrdiv32_fs388_not0 & b[4];
  assign f_arrdiv32_fs388_xor1 = f_arrdiv32_fs387_or0 ^ f_arrdiv32_fs388_xor0;
  assign f_arrdiv32_fs388_not1 = ~f_arrdiv32_fs388_xor0;
  assign f_arrdiv32_fs388_and1 = f_arrdiv32_fs388_not1 & f_arrdiv32_fs387_or0;
  assign f_arrdiv32_fs388_or0 = f_arrdiv32_fs388_and1 | f_arrdiv32_fs388_and0;
  assign f_arrdiv32_fs389_xor0 = f_arrdiv32_mux2to1345_xor0 ^ b[5];
  assign f_arrdiv32_fs389_not0 = ~f_arrdiv32_mux2to1345_xor0;
  assign f_arrdiv32_fs389_and0 = f_arrdiv32_fs389_not0 & b[5];
  assign f_arrdiv32_fs389_xor1 = f_arrdiv32_fs388_or0 ^ f_arrdiv32_fs389_xor0;
  assign f_arrdiv32_fs389_not1 = ~f_arrdiv32_fs389_xor0;
  assign f_arrdiv32_fs389_and1 = f_arrdiv32_fs389_not1 & f_arrdiv32_fs388_or0;
  assign f_arrdiv32_fs389_or0 = f_arrdiv32_fs389_and1 | f_arrdiv32_fs389_and0;
  assign f_arrdiv32_fs390_xor0 = f_arrdiv32_mux2to1346_xor0 ^ b[6];
  assign f_arrdiv32_fs390_not0 = ~f_arrdiv32_mux2to1346_xor0;
  assign f_arrdiv32_fs390_and0 = f_arrdiv32_fs390_not0 & b[6];
  assign f_arrdiv32_fs390_xor1 = f_arrdiv32_fs389_or0 ^ f_arrdiv32_fs390_xor0;
  assign f_arrdiv32_fs390_not1 = ~f_arrdiv32_fs390_xor0;
  assign f_arrdiv32_fs390_and1 = f_arrdiv32_fs390_not1 & f_arrdiv32_fs389_or0;
  assign f_arrdiv32_fs390_or0 = f_arrdiv32_fs390_and1 | f_arrdiv32_fs390_and0;
  assign f_arrdiv32_fs391_xor0 = f_arrdiv32_mux2to1347_xor0 ^ b[7];
  assign f_arrdiv32_fs391_not0 = ~f_arrdiv32_mux2to1347_xor0;
  assign f_arrdiv32_fs391_and0 = f_arrdiv32_fs391_not0 & b[7];
  assign f_arrdiv32_fs391_xor1 = f_arrdiv32_fs390_or0 ^ f_arrdiv32_fs391_xor0;
  assign f_arrdiv32_fs391_not1 = ~f_arrdiv32_fs391_xor0;
  assign f_arrdiv32_fs391_and1 = f_arrdiv32_fs391_not1 & f_arrdiv32_fs390_or0;
  assign f_arrdiv32_fs391_or0 = f_arrdiv32_fs391_and1 | f_arrdiv32_fs391_and0;
  assign f_arrdiv32_fs392_xor0 = f_arrdiv32_mux2to1348_xor0 ^ b[8];
  assign f_arrdiv32_fs392_not0 = ~f_arrdiv32_mux2to1348_xor0;
  assign f_arrdiv32_fs392_and0 = f_arrdiv32_fs392_not0 & b[8];
  assign f_arrdiv32_fs392_xor1 = f_arrdiv32_fs391_or0 ^ f_arrdiv32_fs392_xor0;
  assign f_arrdiv32_fs392_not1 = ~f_arrdiv32_fs392_xor0;
  assign f_arrdiv32_fs392_and1 = f_arrdiv32_fs392_not1 & f_arrdiv32_fs391_or0;
  assign f_arrdiv32_fs392_or0 = f_arrdiv32_fs392_and1 | f_arrdiv32_fs392_and0;
  assign f_arrdiv32_fs393_xor0 = f_arrdiv32_mux2to1349_xor0 ^ b[9];
  assign f_arrdiv32_fs393_not0 = ~f_arrdiv32_mux2to1349_xor0;
  assign f_arrdiv32_fs393_and0 = f_arrdiv32_fs393_not0 & b[9];
  assign f_arrdiv32_fs393_xor1 = f_arrdiv32_fs392_or0 ^ f_arrdiv32_fs393_xor0;
  assign f_arrdiv32_fs393_not1 = ~f_arrdiv32_fs393_xor0;
  assign f_arrdiv32_fs393_and1 = f_arrdiv32_fs393_not1 & f_arrdiv32_fs392_or0;
  assign f_arrdiv32_fs393_or0 = f_arrdiv32_fs393_and1 | f_arrdiv32_fs393_and0;
  assign f_arrdiv32_fs394_xor0 = f_arrdiv32_mux2to1350_xor0 ^ b[10];
  assign f_arrdiv32_fs394_not0 = ~f_arrdiv32_mux2to1350_xor0;
  assign f_arrdiv32_fs394_and0 = f_arrdiv32_fs394_not0 & b[10];
  assign f_arrdiv32_fs394_xor1 = f_arrdiv32_fs393_or0 ^ f_arrdiv32_fs394_xor0;
  assign f_arrdiv32_fs394_not1 = ~f_arrdiv32_fs394_xor0;
  assign f_arrdiv32_fs394_and1 = f_arrdiv32_fs394_not1 & f_arrdiv32_fs393_or0;
  assign f_arrdiv32_fs394_or0 = f_arrdiv32_fs394_and1 | f_arrdiv32_fs394_and0;
  assign f_arrdiv32_fs395_xor0 = f_arrdiv32_mux2to1351_xor0 ^ b[11];
  assign f_arrdiv32_fs395_not0 = ~f_arrdiv32_mux2to1351_xor0;
  assign f_arrdiv32_fs395_and0 = f_arrdiv32_fs395_not0 & b[11];
  assign f_arrdiv32_fs395_xor1 = f_arrdiv32_fs394_or0 ^ f_arrdiv32_fs395_xor0;
  assign f_arrdiv32_fs395_not1 = ~f_arrdiv32_fs395_xor0;
  assign f_arrdiv32_fs395_and1 = f_arrdiv32_fs395_not1 & f_arrdiv32_fs394_or0;
  assign f_arrdiv32_fs395_or0 = f_arrdiv32_fs395_and1 | f_arrdiv32_fs395_and0;
  assign f_arrdiv32_fs396_xor0 = f_arrdiv32_mux2to1352_xor0 ^ b[12];
  assign f_arrdiv32_fs396_not0 = ~f_arrdiv32_mux2to1352_xor0;
  assign f_arrdiv32_fs396_and0 = f_arrdiv32_fs396_not0 & b[12];
  assign f_arrdiv32_fs396_xor1 = f_arrdiv32_fs395_or0 ^ f_arrdiv32_fs396_xor0;
  assign f_arrdiv32_fs396_not1 = ~f_arrdiv32_fs396_xor0;
  assign f_arrdiv32_fs396_and1 = f_arrdiv32_fs396_not1 & f_arrdiv32_fs395_or0;
  assign f_arrdiv32_fs396_or0 = f_arrdiv32_fs396_and1 | f_arrdiv32_fs396_and0;
  assign f_arrdiv32_fs397_xor0 = f_arrdiv32_mux2to1353_xor0 ^ b[13];
  assign f_arrdiv32_fs397_not0 = ~f_arrdiv32_mux2to1353_xor0;
  assign f_arrdiv32_fs397_and0 = f_arrdiv32_fs397_not0 & b[13];
  assign f_arrdiv32_fs397_xor1 = f_arrdiv32_fs396_or0 ^ f_arrdiv32_fs397_xor0;
  assign f_arrdiv32_fs397_not1 = ~f_arrdiv32_fs397_xor0;
  assign f_arrdiv32_fs397_and1 = f_arrdiv32_fs397_not1 & f_arrdiv32_fs396_or0;
  assign f_arrdiv32_fs397_or0 = f_arrdiv32_fs397_and1 | f_arrdiv32_fs397_and0;
  assign f_arrdiv32_fs398_xor0 = f_arrdiv32_mux2to1354_xor0 ^ b[14];
  assign f_arrdiv32_fs398_not0 = ~f_arrdiv32_mux2to1354_xor0;
  assign f_arrdiv32_fs398_and0 = f_arrdiv32_fs398_not0 & b[14];
  assign f_arrdiv32_fs398_xor1 = f_arrdiv32_fs397_or0 ^ f_arrdiv32_fs398_xor0;
  assign f_arrdiv32_fs398_not1 = ~f_arrdiv32_fs398_xor0;
  assign f_arrdiv32_fs398_and1 = f_arrdiv32_fs398_not1 & f_arrdiv32_fs397_or0;
  assign f_arrdiv32_fs398_or0 = f_arrdiv32_fs398_and1 | f_arrdiv32_fs398_and0;
  assign f_arrdiv32_fs399_xor0 = f_arrdiv32_mux2to1355_xor0 ^ b[15];
  assign f_arrdiv32_fs399_not0 = ~f_arrdiv32_mux2to1355_xor0;
  assign f_arrdiv32_fs399_and0 = f_arrdiv32_fs399_not0 & b[15];
  assign f_arrdiv32_fs399_xor1 = f_arrdiv32_fs398_or0 ^ f_arrdiv32_fs399_xor0;
  assign f_arrdiv32_fs399_not1 = ~f_arrdiv32_fs399_xor0;
  assign f_arrdiv32_fs399_and1 = f_arrdiv32_fs399_not1 & f_arrdiv32_fs398_or0;
  assign f_arrdiv32_fs399_or0 = f_arrdiv32_fs399_and1 | f_arrdiv32_fs399_and0;
  assign f_arrdiv32_fs400_xor0 = f_arrdiv32_mux2to1356_xor0 ^ b[16];
  assign f_arrdiv32_fs400_not0 = ~f_arrdiv32_mux2to1356_xor0;
  assign f_arrdiv32_fs400_and0 = f_arrdiv32_fs400_not0 & b[16];
  assign f_arrdiv32_fs400_xor1 = f_arrdiv32_fs399_or0 ^ f_arrdiv32_fs400_xor0;
  assign f_arrdiv32_fs400_not1 = ~f_arrdiv32_fs400_xor0;
  assign f_arrdiv32_fs400_and1 = f_arrdiv32_fs400_not1 & f_arrdiv32_fs399_or0;
  assign f_arrdiv32_fs400_or0 = f_arrdiv32_fs400_and1 | f_arrdiv32_fs400_and0;
  assign f_arrdiv32_fs401_xor0 = f_arrdiv32_mux2to1357_xor0 ^ b[17];
  assign f_arrdiv32_fs401_not0 = ~f_arrdiv32_mux2to1357_xor0;
  assign f_arrdiv32_fs401_and0 = f_arrdiv32_fs401_not0 & b[17];
  assign f_arrdiv32_fs401_xor1 = f_arrdiv32_fs400_or0 ^ f_arrdiv32_fs401_xor0;
  assign f_arrdiv32_fs401_not1 = ~f_arrdiv32_fs401_xor0;
  assign f_arrdiv32_fs401_and1 = f_arrdiv32_fs401_not1 & f_arrdiv32_fs400_or0;
  assign f_arrdiv32_fs401_or0 = f_arrdiv32_fs401_and1 | f_arrdiv32_fs401_and0;
  assign f_arrdiv32_fs402_xor0 = f_arrdiv32_mux2to1358_xor0 ^ b[18];
  assign f_arrdiv32_fs402_not0 = ~f_arrdiv32_mux2to1358_xor0;
  assign f_arrdiv32_fs402_and0 = f_arrdiv32_fs402_not0 & b[18];
  assign f_arrdiv32_fs402_xor1 = f_arrdiv32_fs401_or0 ^ f_arrdiv32_fs402_xor0;
  assign f_arrdiv32_fs402_not1 = ~f_arrdiv32_fs402_xor0;
  assign f_arrdiv32_fs402_and1 = f_arrdiv32_fs402_not1 & f_arrdiv32_fs401_or0;
  assign f_arrdiv32_fs402_or0 = f_arrdiv32_fs402_and1 | f_arrdiv32_fs402_and0;
  assign f_arrdiv32_fs403_xor0 = f_arrdiv32_mux2to1359_xor0 ^ b[19];
  assign f_arrdiv32_fs403_not0 = ~f_arrdiv32_mux2to1359_xor0;
  assign f_arrdiv32_fs403_and0 = f_arrdiv32_fs403_not0 & b[19];
  assign f_arrdiv32_fs403_xor1 = f_arrdiv32_fs402_or0 ^ f_arrdiv32_fs403_xor0;
  assign f_arrdiv32_fs403_not1 = ~f_arrdiv32_fs403_xor0;
  assign f_arrdiv32_fs403_and1 = f_arrdiv32_fs403_not1 & f_arrdiv32_fs402_or0;
  assign f_arrdiv32_fs403_or0 = f_arrdiv32_fs403_and1 | f_arrdiv32_fs403_and0;
  assign f_arrdiv32_fs404_xor0 = f_arrdiv32_mux2to1360_xor0 ^ b[20];
  assign f_arrdiv32_fs404_not0 = ~f_arrdiv32_mux2to1360_xor0;
  assign f_arrdiv32_fs404_and0 = f_arrdiv32_fs404_not0 & b[20];
  assign f_arrdiv32_fs404_xor1 = f_arrdiv32_fs403_or0 ^ f_arrdiv32_fs404_xor0;
  assign f_arrdiv32_fs404_not1 = ~f_arrdiv32_fs404_xor0;
  assign f_arrdiv32_fs404_and1 = f_arrdiv32_fs404_not1 & f_arrdiv32_fs403_or0;
  assign f_arrdiv32_fs404_or0 = f_arrdiv32_fs404_and1 | f_arrdiv32_fs404_and0;
  assign f_arrdiv32_fs405_xor0 = f_arrdiv32_mux2to1361_xor0 ^ b[21];
  assign f_arrdiv32_fs405_not0 = ~f_arrdiv32_mux2to1361_xor0;
  assign f_arrdiv32_fs405_and0 = f_arrdiv32_fs405_not0 & b[21];
  assign f_arrdiv32_fs405_xor1 = f_arrdiv32_fs404_or0 ^ f_arrdiv32_fs405_xor0;
  assign f_arrdiv32_fs405_not1 = ~f_arrdiv32_fs405_xor0;
  assign f_arrdiv32_fs405_and1 = f_arrdiv32_fs405_not1 & f_arrdiv32_fs404_or0;
  assign f_arrdiv32_fs405_or0 = f_arrdiv32_fs405_and1 | f_arrdiv32_fs405_and0;
  assign f_arrdiv32_fs406_xor0 = f_arrdiv32_mux2to1362_xor0 ^ b[22];
  assign f_arrdiv32_fs406_not0 = ~f_arrdiv32_mux2to1362_xor0;
  assign f_arrdiv32_fs406_and0 = f_arrdiv32_fs406_not0 & b[22];
  assign f_arrdiv32_fs406_xor1 = f_arrdiv32_fs405_or0 ^ f_arrdiv32_fs406_xor0;
  assign f_arrdiv32_fs406_not1 = ~f_arrdiv32_fs406_xor0;
  assign f_arrdiv32_fs406_and1 = f_arrdiv32_fs406_not1 & f_arrdiv32_fs405_or0;
  assign f_arrdiv32_fs406_or0 = f_arrdiv32_fs406_and1 | f_arrdiv32_fs406_and0;
  assign f_arrdiv32_fs407_xor0 = f_arrdiv32_mux2to1363_xor0 ^ b[23];
  assign f_arrdiv32_fs407_not0 = ~f_arrdiv32_mux2to1363_xor0;
  assign f_arrdiv32_fs407_and0 = f_arrdiv32_fs407_not0 & b[23];
  assign f_arrdiv32_fs407_xor1 = f_arrdiv32_fs406_or0 ^ f_arrdiv32_fs407_xor0;
  assign f_arrdiv32_fs407_not1 = ~f_arrdiv32_fs407_xor0;
  assign f_arrdiv32_fs407_and1 = f_arrdiv32_fs407_not1 & f_arrdiv32_fs406_or0;
  assign f_arrdiv32_fs407_or0 = f_arrdiv32_fs407_and1 | f_arrdiv32_fs407_and0;
  assign f_arrdiv32_fs408_xor0 = f_arrdiv32_mux2to1364_xor0 ^ b[24];
  assign f_arrdiv32_fs408_not0 = ~f_arrdiv32_mux2to1364_xor0;
  assign f_arrdiv32_fs408_and0 = f_arrdiv32_fs408_not0 & b[24];
  assign f_arrdiv32_fs408_xor1 = f_arrdiv32_fs407_or0 ^ f_arrdiv32_fs408_xor0;
  assign f_arrdiv32_fs408_not1 = ~f_arrdiv32_fs408_xor0;
  assign f_arrdiv32_fs408_and1 = f_arrdiv32_fs408_not1 & f_arrdiv32_fs407_or0;
  assign f_arrdiv32_fs408_or0 = f_arrdiv32_fs408_and1 | f_arrdiv32_fs408_and0;
  assign f_arrdiv32_fs409_xor0 = f_arrdiv32_mux2to1365_xor0 ^ b[25];
  assign f_arrdiv32_fs409_not0 = ~f_arrdiv32_mux2to1365_xor0;
  assign f_arrdiv32_fs409_and0 = f_arrdiv32_fs409_not0 & b[25];
  assign f_arrdiv32_fs409_xor1 = f_arrdiv32_fs408_or0 ^ f_arrdiv32_fs409_xor0;
  assign f_arrdiv32_fs409_not1 = ~f_arrdiv32_fs409_xor0;
  assign f_arrdiv32_fs409_and1 = f_arrdiv32_fs409_not1 & f_arrdiv32_fs408_or0;
  assign f_arrdiv32_fs409_or0 = f_arrdiv32_fs409_and1 | f_arrdiv32_fs409_and0;
  assign f_arrdiv32_fs410_xor0 = f_arrdiv32_mux2to1366_xor0 ^ b[26];
  assign f_arrdiv32_fs410_not0 = ~f_arrdiv32_mux2to1366_xor0;
  assign f_arrdiv32_fs410_and0 = f_arrdiv32_fs410_not0 & b[26];
  assign f_arrdiv32_fs410_xor1 = f_arrdiv32_fs409_or0 ^ f_arrdiv32_fs410_xor0;
  assign f_arrdiv32_fs410_not1 = ~f_arrdiv32_fs410_xor0;
  assign f_arrdiv32_fs410_and1 = f_arrdiv32_fs410_not1 & f_arrdiv32_fs409_or0;
  assign f_arrdiv32_fs410_or0 = f_arrdiv32_fs410_and1 | f_arrdiv32_fs410_and0;
  assign f_arrdiv32_fs411_xor0 = f_arrdiv32_mux2to1367_xor0 ^ b[27];
  assign f_arrdiv32_fs411_not0 = ~f_arrdiv32_mux2to1367_xor0;
  assign f_arrdiv32_fs411_and0 = f_arrdiv32_fs411_not0 & b[27];
  assign f_arrdiv32_fs411_xor1 = f_arrdiv32_fs410_or0 ^ f_arrdiv32_fs411_xor0;
  assign f_arrdiv32_fs411_not1 = ~f_arrdiv32_fs411_xor0;
  assign f_arrdiv32_fs411_and1 = f_arrdiv32_fs411_not1 & f_arrdiv32_fs410_or0;
  assign f_arrdiv32_fs411_or0 = f_arrdiv32_fs411_and1 | f_arrdiv32_fs411_and0;
  assign f_arrdiv32_fs412_xor0 = f_arrdiv32_mux2to1368_xor0 ^ b[28];
  assign f_arrdiv32_fs412_not0 = ~f_arrdiv32_mux2to1368_xor0;
  assign f_arrdiv32_fs412_and0 = f_arrdiv32_fs412_not0 & b[28];
  assign f_arrdiv32_fs412_xor1 = f_arrdiv32_fs411_or0 ^ f_arrdiv32_fs412_xor0;
  assign f_arrdiv32_fs412_not1 = ~f_arrdiv32_fs412_xor0;
  assign f_arrdiv32_fs412_and1 = f_arrdiv32_fs412_not1 & f_arrdiv32_fs411_or0;
  assign f_arrdiv32_fs412_or0 = f_arrdiv32_fs412_and1 | f_arrdiv32_fs412_and0;
  assign f_arrdiv32_fs413_xor0 = f_arrdiv32_mux2to1369_xor0 ^ b[29];
  assign f_arrdiv32_fs413_not0 = ~f_arrdiv32_mux2to1369_xor0;
  assign f_arrdiv32_fs413_and0 = f_arrdiv32_fs413_not0 & b[29];
  assign f_arrdiv32_fs413_xor1 = f_arrdiv32_fs412_or0 ^ f_arrdiv32_fs413_xor0;
  assign f_arrdiv32_fs413_not1 = ~f_arrdiv32_fs413_xor0;
  assign f_arrdiv32_fs413_and1 = f_arrdiv32_fs413_not1 & f_arrdiv32_fs412_or0;
  assign f_arrdiv32_fs413_or0 = f_arrdiv32_fs413_and1 | f_arrdiv32_fs413_and0;
  assign f_arrdiv32_fs414_xor0 = f_arrdiv32_mux2to1370_xor0 ^ b[30];
  assign f_arrdiv32_fs414_not0 = ~f_arrdiv32_mux2to1370_xor0;
  assign f_arrdiv32_fs414_and0 = f_arrdiv32_fs414_not0 & b[30];
  assign f_arrdiv32_fs414_xor1 = f_arrdiv32_fs413_or0 ^ f_arrdiv32_fs414_xor0;
  assign f_arrdiv32_fs414_not1 = ~f_arrdiv32_fs414_xor0;
  assign f_arrdiv32_fs414_and1 = f_arrdiv32_fs414_not1 & f_arrdiv32_fs413_or0;
  assign f_arrdiv32_fs414_or0 = f_arrdiv32_fs414_and1 | f_arrdiv32_fs414_and0;
  assign f_arrdiv32_fs415_xor0 = f_arrdiv32_mux2to1371_xor0 ^ b[31];
  assign f_arrdiv32_fs415_not0 = ~f_arrdiv32_mux2to1371_xor0;
  assign f_arrdiv32_fs415_and0 = f_arrdiv32_fs415_not0 & b[31];
  assign f_arrdiv32_fs415_xor1 = f_arrdiv32_fs414_or0 ^ f_arrdiv32_fs415_xor0;
  assign f_arrdiv32_fs415_not1 = ~f_arrdiv32_fs415_xor0;
  assign f_arrdiv32_fs415_and1 = f_arrdiv32_fs415_not1 & f_arrdiv32_fs414_or0;
  assign f_arrdiv32_fs415_or0 = f_arrdiv32_fs415_and1 | f_arrdiv32_fs415_and0;
  assign f_arrdiv32_mux2to1372_and0 = a[19] & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1372_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1372_and1 = f_arrdiv32_fs384_xor0 & f_arrdiv32_mux2to1372_not0;
  assign f_arrdiv32_mux2to1372_xor0 = f_arrdiv32_mux2to1372_and0 ^ f_arrdiv32_mux2to1372_and1;
  assign f_arrdiv32_mux2to1373_and0 = f_arrdiv32_mux2to1341_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1373_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1373_and1 = f_arrdiv32_fs385_xor1 & f_arrdiv32_mux2to1373_not0;
  assign f_arrdiv32_mux2to1373_xor0 = f_arrdiv32_mux2to1373_and0 ^ f_arrdiv32_mux2to1373_and1;
  assign f_arrdiv32_mux2to1374_and0 = f_arrdiv32_mux2to1342_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1374_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1374_and1 = f_arrdiv32_fs386_xor1 & f_arrdiv32_mux2to1374_not0;
  assign f_arrdiv32_mux2to1374_xor0 = f_arrdiv32_mux2to1374_and0 ^ f_arrdiv32_mux2to1374_and1;
  assign f_arrdiv32_mux2to1375_and0 = f_arrdiv32_mux2to1343_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1375_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1375_and1 = f_arrdiv32_fs387_xor1 & f_arrdiv32_mux2to1375_not0;
  assign f_arrdiv32_mux2to1375_xor0 = f_arrdiv32_mux2to1375_and0 ^ f_arrdiv32_mux2to1375_and1;
  assign f_arrdiv32_mux2to1376_and0 = f_arrdiv32_mux2to1344_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1376_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1376_and1 = f_arrdiv32_fs388_xor1 & f_arrdiv32_mux2to1376_not0;
  assign f_arrdiv32_mux2to1376_xor0 = f_arrdiv32_mux2to1376_and0 ^ f_arrdiv32_mux2to1376_and1;
  assign f_arrdiv32_mux2to1377_and0 = f_arrdiv32_mux2to1345_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1377_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1377_and1 = f_arrdiv32_fs389_xor1 & f_arrdiv32_mux2to1377_not0;
  assign f_arrdiv32_mux2to1377_xor0 = f_arrdiv32_mux2to1377_and0 ^ f_arrdiv32_mux2to1377_and1;
  assign f_arrdiv32_mux2to1378_and0 = f_arrdiv32_mux2to1346_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1378_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1378_and1 = f_arrdiv32_fs390_xor1 & f_arrdiv32_mux2to1378_not0;
  assign f_arrdiv32_mux2to1378_xor0 = f_arrdiv32_mux2to1378_and0 ^ f_arrdiv32_mux2to1378_and1;
  assign f_arrdiv32_mux2to1379_and0 = f_arrdiv32_mux2to1347_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1379_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1379_and1 = f_arrdiv32_fs391_xor1 & f_arrdiv32_mux2to1379_not0;
  assign f_arrdiv32_mux2to1379_xor0 = f_arrdiv32_mux2to1379_and0 ^ f_arrdiv32_mux2to1379_and1;
  assign f_arrdiv32_mux2to1380_and0 = f_arrdiv32_mux2to1348_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1380_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1380_and1 = f_arrdiv32_fs392_xor1 & f_arrdiv32_mux2to1380_not0;
  assign f_arrdiv32_mux2to1380_xor0 = f_arrdiv32_mux2to1380_and0 ^ f_arrdiv32_mux2to1380_and1;
  assign f_arrdiv32_mux2to1381_and0 = f_arrdiv32_mux2to1349_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1381_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1381_and1 = f_arrdiv32_fs393_xor1 & f_arrdiv32_mux2to1381_not0;
  assign f_arrdiv32_mux2to1381_xor0 = f_arrdiv32_mux2to1381_and0 ^ f_arrdiv32_mux2to1381_and1;
  assign f_arrdiv32_mux2to1382_and0 = f_arrdiv32_mux2to1350_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1382_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1382_and1 = f_arrdiv32_fs394_xor1 & f_arrdiv32_mux2to1382_not0;
  assign f_arrdiv32_mux2to1382_xor0 = f_arrdiv32_mux2to1382_and0 ^ f_arrdiv32_mux2to1382_and1;
  assign f_arrdiv32_mux2to1383_and0 = f_arrdiv32_mux2to1351_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1383_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1383_and1 = f_arrdiv32_fs395_xor1 & f_arrdiv32_mux2to1383_not0;
  assign f_arrdiv32_mux2to1383_xor0 = f_arrdiv32_mux2to1383_and0 ^ f_arrdiv32_mux2to1383_and1;
  assign f_arrdiv32_mux2to1384_and0 = f_arrdiv32_mux2to1352_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1384_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1384_and1 = f_arrdiv32_fs396_xor1 & f_arrdiv32_mux2to1384_not0;
  assign f_arrdiv32_mux2to1384_xor0 = f_arrdiv32_mux2to1384_and0 ^ f_arrdiv32_mux2to1384_and1;
  assign f_arrdiv32_mux2to1385_and0 = f_arrdiv32_mux2to1353_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1385_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1385_and1 = f_arrdiv32_fs397_xor1 & f_arrdiv32_mux2to1385_not0;
  assign f_arrdiv32_mux2to1385_xor0 = f_arrdiv32_mux2to1385_and0 ^ f_arrdiv32_mux2to1385_and1;
  assign f_arrdiv32_mux2to1386_and0 = f_arrdiv32_mux2to1354_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1386_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1386_and1 = f_arrdiv32_fs398_xor1 & f_arrdiv32_mux2to1386_not0;
  assign f_arrdiv32_mux2to1386_xor0 = f_arrdiv32_mux2to1386_and0 ^ f_arrdiv32_mux2to1386_and1;
  assign f_arrdiv32_mux2to1387_and0 = f_arrdiv32_mux2to1355_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1387_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1387_and1 = f_arrdiv32_fs399_xor1 & f_arrdiv32_mux2to1387_not0;
  assign f_arrdiv32_mux2to1387_xor0 = f_arrdiv32_mux2to1387_and0 ^ f_arrdiv32_mux2to1387_and1;
  assign f_arrdiv32_mux2to1388_and0 = f_arrdiv32_mux2to1356_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1388_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1388_and1 = f_arrdiv32_fs400_xor1 & f_arrdiv32_mux2to1388_not0;
  assign f_arrdiv32_mux2to1388_xor0 = f_arrdiv32_mux2to1388_and0 ^ f_arrdiv32_mux2to1388_and1;
  assign f_arrdiv32_mux2to1389_and0 = f_arrdiv32_mux2to1357_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1389_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1389_and1 = f_arrdiv32_fs401_xor1 & f_arrdiv32_mux2to1389_not0;
  assign f_arrdiv32_mux2to1389_xor0 = f_arrdiv32_mux2to1389_and0 ^ f_arrdiv32_mux2to1389_and1;
  assign f_arrdiv32_mux2to1390_and0 = f_arrdiv32_mux2to1358_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1390_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1390_and1 = f_arrdiv32_fs402_xor1 & f_arrdiv32_mux2to1390_not0;
  assign f_arrdiv32_mux2to1390_xor0 = f_arrdiv32_mux2to1390_and0 ^ f_arrdiv32_mux2to1390_and1;
  assign f_arrdiv32_mux2to1391_and0 = f_arrdiv32_mux2to1359_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1391_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1391_and1 = f_arrdiv32_fs403_xor1 & f_arrdiv32_mux2to1391_not0;
  assign f_arrdiv32_mux2to1391_xor0 = f_arrdiv32_mux2to1391_and0 ^ f_arrdiv32_mux2to1391_and1;
  assign f_arrdiv32_mux2to1392_and0 = f_arrdiv32_mux2to1360_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1392_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1392_and1 = f_arrdiv32_fs404_xor1 & f_arrdiv32_mux2to1392_not0;
  assign f_arrdiv32_mux2to1392_xor0 = f_arrdiv32_mux2to1392_and0 ^ f_arrdiv32_mux2to1392_and1;
  assign f_arrdiv32_mux2to1393_and0 = f_arrdiv32_mux2to1361_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1393_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1393_and1 = f_arrdiv32_fs405_xor1 & f_arrdiv32_mux2to1393_not0;
  assign f_arrdiv32_mux2to1393_xor0 = f_arrdiv32_mux2to1393_and0 ^ f_arrdiv32_mux2to1393_and1;
  assign f_arrdiv32_mux2to1394_and0 = f_arrdiv32_mux2to1362_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1394_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1394_and1 = f_arrdiv32_fs406_xor1 & f_arrdiv32_mux2to1394_not0;
  assign f_arrdiv32_mux2to1394_xor0 = f_arrdiv32_mux2to1394_and0 ^ f_arrdiv32_mux2to1394_and1;
  assign f_arrdiv32_mux2to1395_and0 = f_arrdiv32_mux2to1363_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1395_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1395_and1 = f_arrdiv32_fs407_xor1 & f_arrdiv32_mux2to1395_not0;
  assign f_arrdiv32_mux2to1395_xor0 = f_arrdiv32_mux2to1395_and0 ^ f_arrdiv32_mux2to1395_and1;
  assign f_arrdiv32_mux2to1396_and0 = f_arrdiv32_mux2to1364_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1396_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1396_and1 = f_arrdiv32_fs408_xor1 & f_arrdiv32_mux2to1396_not0;
  assign f_arrdiv32_mux2to1396_xor0 = f_arrdiv32_mux2to1396_and0 ^ f_arrdiv32_mux2to1396_and1;
  assign f_arrdiv32_mux2to1397_and0 = f_arrdiv32_mux2to1365_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1397_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1397_and1 = f_arrdiv32_fs409_xor1 & f_arrdiv32_mux2to1397_not0;
  assign f_arrdiv32_mux2to1397_xor0 = f_arrdiv32_mux2to1397_and0 ^ f_arrdiv32_mux2to1397_and1;
  assign f_arrdiv32_mux2to1398_and0 = f_arrdiv32_mux2to1366_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1398_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1398_and1 = f_arrdiv32_fs410_xor1 & f_arrdiv32_mux2to1398_not0;
  assign f_arrdiv32_mux2to1398_xor0 = f_arrdiv32_mux2to1398_and0 ^ f_arrdiv32_mux2to1398_and1;
  assign f_arrdiv32_mux2to1399_and0 = f_arrdiv32_mux2to1367_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1399_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1399_and1 = f_arrdiv32_fs411_xor1 & f_arrdiv32_mux2to1399_not0;
  assign f_arrdiv32_mux2to1399_xor0 = f_arrdiv32_mux2to1399_and0 ^ f_arrdiv32_mux2to1399_and1;
  assign f_arrdiv32_mux2to1400_and0 = f_arrdiv32_mux2to1368_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1400_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1400_and1 = f_arrdiv32_fs412_xor1 & f_arrdiv32_mux2to1400_not0;
  assign f_arrdiv32_mux2to1400_xor0 = f_arrdiv32_mux2to1400_and0 ^ f_arrdiv32_mux2to1400_and1;
  assign f_arrdiv32_mux2to1401_and0 = f_arrdiv32_mux2to1369_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1401_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1401_and1 = f_arrdiv32_fs413_xor1 & f_arrdiv32_mux2to1401_not0;
  assign f_arrdiv32_mux2to1401_xor0 = f_arrdiv32_mux2to1401_and0 ^ f_arrdiv32_mux2to1401_and1;
  assign f_arrdiv32_mux2to1402_and0 = f_arrdiv32_mux2to1370_xor0 & f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1402_not0 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_mux2to1402_and1 = f_arrdiv32_fs414_xor1 & f_arrdiv32_mux2to1402_not0;
  assign f_arrdiv32_mux2to1402_xor0 = f_arrdiv32_mux2to1402_and0 ^ f_arrdiv32_mux2to1402_and1;
  assign f_arrdiv32_not12 = ~f_arrdiv32_fs415_or0;
  assign f_arrdiv32_fs416_xor0 = a[18] ^ b[0];
  assign f_arrdiv32_fs416_not0 = ~a[18];
  assign f_arrdiv32_fs416_and0 = f_arrdiv32_fs416_not0 & b[0];
  assign f_arrdiv32_fs416_not1 = ~f_arrdiv32_fs416_xor0;
  assign f_arrdiv32_fs417_xor0 = f_arrdiv32_mux2to1372_xor0 ^ b[1];
  assign f_arrdiv32_fs417_not0 = ~f_arrdiv32_mux2to1372_xor0;
  assign f_arrdiv32_fs417_and0 = f_arrdiv32_fs417_not0 & b[1];
  assign f_arrdiv32_fs417_xor1 = f_arrdiv32_fs416_and0 ^ f_arrdiv32_fs417_xor0;
  assign f_arrdiv32_fs417_not1 = ~f_arrdiv32_fs417_xor0;
  assign f_arrdiv32_fs417_and1 = f_arrdiv32_fs417_not1 & f_arrdiv32_fs416_and0;
  assign f_arrdiv32_fs417_or0 = f_arrdiv32_fs417_and1 | f_arrdiv32_fs417_and0;
  assign f_arrdiv32_fs418_xor0 = f_arrdiv32_mux2to1373_xor0 ^ b[2];
  assign f_arrdiv32_fs418_not0 = ~f_arrdiv32_mux2to1373_xor0;
  assign f_arrdiv32_fs418_and0 = f_arrdiv32_fs418_not0 & b[2];
  assign f_arrdiv32_fs418_xor1 = f_arrdiv32_fs417_or0 ^ f_arrdiv32_fs418_xor0;
  assign f_arrdiv32_fs418_not1 = ~f_arrdiv32_fs418_xor0;
  assign f_arrdiv32_fs418_and1 = f_arrdiv32_fs418_not1 & f_arrdiv32_fs417_or0;
  assign f_arrdiv32_fs418_or0 = f_arrdiv32_fs418_and1 | f_arrdiv32_fs418_and0;
  assign f_arrdiv32_fs419_xor0 = f_arrdiv32_mux2to1374_xor0 ^ b[3];
  assign f_arrdiv32_fs419_not0 = ~f_arrdiv32_mux2to1374_xor0;
  assign f_arrdiv32_fs419_and0 = f_arrdiv32_fs419_not0 & b[3];
  assign f_arrdiv32_fs419_xor1 = f_arrdiv32_fs418_or0 ^ f_arrdiv32_fs419_xor0;
  assign f_arrdiv32_fs419_not1 = ~f_arrdiv32_fs419_xor0;
  assign f_arrdiv32_fs419_and1 = f_arrdiv32_fs419_not1 & f_arrdiv32_fs418_or0;
  assign f_arrdiv32_fs419_or0 = f_arrdiv32_fs419_and1 | f_arrdiv32_fs419_and0;
  assign f_arrdiv32_fs420_xor0 = f_arrdiv32_mux2to1375_xor0 ^ b[4];
  assign f_arrdiv32_fs420_not0 = ~f_arrdiv32_mux2to1375_xor0;
  assign f_arrdiv32_fs420_and0 = f_arrdiv32_fs420_not0 & b[4];
  assign f_arrdiv32_fs420_xor1 = f_arrdiv32_fs419_or0 ^ f_arrdiv32_fs420_xor0;
  assign f_arrdiv32_fs420_not1 = ~f_arrdiv32_fs420_xor0;
  assign f_arrdiv32_fs420_and1 = f_arrdiv32_fs420_not1 & f_arrdiv32_fs419_or0;
  assign f_arrdiv32_fs420_or0 = f_arrdiv32_fs420_and1 | f_arrdiv32_fs420_and0;
  assign f_arrdiv32_fs421_xor0 = f_arrdiv32_mux2to1376_xor0 ^ b[5];
  assign f_arrdiv32_fs421_not0 = ~f_arrdiv32_mux2to1376_xor0;
  assign f_arrdiv32_fs421_and0 = f_arrdiv32_fs421_not0 & b[5];
  assign f_arrdiv32_fs421_xor1 = f_arrdiv32_fs420_or0 ^ f_arrdiv32_fs421_xor0;
  assign f_arrdiv32_fs421_not1 = ~f_arrdiv32_fs421_xor0;
  assign f_arrdiv32_fs421_and1 = f_arrdiv32_fs421_not1 & f_arrdiv32_fs420_or0;
  assign f_arrdiv32_fs421_or0 = f_arrdiv32_fs421_and1 | f_arrdiv32_fs421_and0;
  assign f_arrdiv32_fs422_xor0 = f_arrdiv32_mux2to1377_xor0 ^ b[6];
  assign f_arrdiv32_fs422_not0 = ~f_arrdiv32_mux2to1377_xor0;
  assign f_arrdiv32_fs422_and0 = f_arrdiv32_fs422_not0 & b[6];
  assign f_arrdiv32_fs422_xor1 = f_arrdiv32_fs421_or0 ^ f_arrdiv32_fs422_xor0;
  assign f_arrdiv32_fs422_not1 = ~f_arrdiv32_fs422_xor0;
  assign f_arrdiv32_fs422_and1 = f_arrdiv32_fs422_not1 & f_arrdiv32_fs421_or0;
  assign f_arrdiv32_fs422_or0 = f_arrdiv32_fs422_and1 | f_arrdiv32_fs422_and0;
  assign f_arrdiv32_fs423_xor0 = f_arrdiv32_mux2to1378_xor0 ^ b[7];
  assign f_arrdiv32_fs423_not0 = ~f_arrdiv32_mux2to1378_xor0;
  assign f_arrdiv32_fs423_and0 = f_arrdiv32_fs423_not0 & b[7];
  assign f_arrdiv32_fs423_xor1 = f_arrdiv32_fs422_or0 ^ f_arrdiv32_fs423_xor0;
  assign f_arrdiv32_fs423_not1 = ~f_arrdiv32_fs423_xor0;
  assign f_arrdiv32_fs423_and1 = f_arrdiv32_fs423_not1 & f_arrdiv32_fs422_or0;
  assign f_arrdiv32_fs423_or0 = f_arrdiv32_fs423_and1 | f_arrdiv32_fs423_and0;
  assign f_arrdiv32_fs424_xor0 = f_arrdiv32_mux2to1379_xor0 ^ b[8];
  assign f_arrdiv32_fs424_not0 = ~f_arrdiv32_mux2to1379_xor0;
  assign f_arrdiv32_fs424_and0 = f_arrdiv32_fs424_not0 & b[8];
  assign f_arrdiv32_fs424_xor1 = f_arrdiv32_fs423_or0 ^ f_arrdiv32_fs424_xor0;
  assign f_arrdiv32_fs424_not1 = ~f_arrdiv32_fs424_xor0;
  assign f_arrdiv32_fs424_and1 = f_arrdiv32_fs424_not1 & f_arrdiv32_fs423_or0;
  assign f_arrdiv32_fs424_or0 = f_arrdiv32_fs424_and1 | f_arrdiv32_fs424_and0;
  assign f_arrdiv32_fs425_xor0 = f_arrdiv32_mux2to1380_xor0 ^ b[9];
  assign f_arrdiv32_fs425_not0 = ~f_arrdiv32_mux2to1380_xor0;
  assign f_arrdiv32_fs425_and0 = f_arrdiv32_fs425_not0 & b[9];
  assign f_arrdiv32_fs425_xor1 = f_arrdiv32_fs424_or0 ^ f_arrdiv32_fs425_xor0;
  assign f_arrdiv32_fs425_not1 = ~f_arrdiv32_fs425_xor0;
  assign f_arrdiv32_fs425_and1 = f_arrdiv32_fs425_not1 & f_arrdiv32_fs424_or0;
  assign f_arrdiv32_fs425_or0 = f_arrdiv32_fs425_and1 | f_arrdiv32_fs425_and0;
  assign f_arrdiv32_fs426_xor0 = f_arrdiv32_mux2to1381_xor0 ^ b[10];
  assign f_arrdiv32_fs426_not0 = ~f_arrdiv32_mux2to1381_xor0;
  assign f_arrdiv32_fs426_and0 = f_arrdiv32_fs426_not0 & b[10];
  assign f_arrdiv32_fs426_xor1 = f_arrdiv32_fs425_or0 ^ f_arrdiv32_fs426_xor0;
  assign f_arrdiv32_fs426_not1 = ~f_arrdiv32_fs426_xor0;
  assign f_arrdiv32_fs426_and1 = f_arrdiv32_fs426_not1 & f_arrdiv32_fs425_or0;
  assign f_arrdiv32_fs426_or0 = f_arrdiv32_fs426_and1 | f_arrdiv32_fs426_and0;
  assign f_arrdiv32_fs427_xor0 = f_arrdiv32_mux2to1382_xor0 ^ b[11];
  assign f_arrdiv32_fs427_not0 = ~f_arrdiv32_mux2to1382_xor0;
  assign f_arrdiv32_fs427_and0 = f_arrdiv32_fs427_not0 & b[11];
  assign f_arrdiv32_fs427_xor1 = f_arrdiv32_fs426_or0 ^ f_arrdiv32_fs427_xor0;
  assign f_arrdiv32_fs427_not1 = ~f_arrdiv32_fs427_xor0;
  assign f_arrdiv32_fs427_and1 = f_arrdiv32_fs427_not1 & f_arrdiv32_fs426_or0;
  assign f_arrdiv32_fs427_or0 = f_arrdiv32_fs427_and1 | f_arrdiv32_fs427_and0;
  assign f_arrdiv32_fs428_xor0 = f_arrdiv32_mux2to1383_xor0 ^ b[12];
  assign f_arrdiv32_fs428_not0 = ~f_arrdiv32_mux2to1383_xor0;
  assign f_arrdiv32_fs428_and0 = f_arrdiv32_fs428_not0 & b[12];
  assign f_arrdiv32_fs428_xor1 = f_arrdiv32_fs427_or0 ^ f_arrdiv32_fs428_xor0;
  assign f_arrdiv32_fs428_not1 = ~f_arrdiv32_fs428_xor0;
  assign f_arrdiv32_fs428_and1 = f_arrdiv32_fs428_not1 & f_arrdiv32_fs427_or0;
  assign f_arrdiv32_fs428_or0 = f_arrdiv32_fs428_and1 | f_arrdiv32_fs428_and0;
  assign f_arrdiv32_fs429_xor0 = f_arrdiv32_mux2to1384_xor0 ^ b[13];
  assign f_arrdiv32_fs429_not0 = ~f_arrdiv32_mux2to1384_xor0;
  assign f_arrdiv32_fs429_and0 = f_arrdiv32_fs429_not0 & b[13];
  assign f_arrdiv32_fs429_xor1 = f_arrdiv32_fs428_or0 ^ f_arrdiv32_fs429_xor0;
  assign f_arrdiv32_fs429_not1 = ~f_arrdiv32_fs429_xor0;
  assign f_arrdiv32_fs429_and1 = f_arrdiv32_fs429_not1 & f_arrdiv32_fs428_or0;
  assign f_arrdiv32_fs429_or0 = f_arrdiv32_fs429_and1 | f_arrdiv32_fs429_and0;
  assign f_arrdiv32_fs430_xor0 = f_arrdiv32_mux2to1385_xor0 ^ b[14];
  assign f_arrdiv32_fs430_not0 = ~f_arrdiv32_mux2to1385_xor0;
  assign f_arrdiv32_fs430_and0 = f_arrdiv32_fs430_not0 & b[14];
  assign f_arrdiv32_fs430_xor1 = f_arrdiv32_fs429_or0 ^ f_arrdiv32_fs430_xor0;
  assign f_arrdiv32_fs430_not1 = ~f_arrdiv32_fs430_xor0;
  assign f_arrdiv32_fs430_and1 = f_arrdiv32_fs430_not1 & f_arrdiv32_fs429_or0;
  assign f_arrdiv32_fs430_or0 = f_arrdiv32_fs430_and1 | f_arrdiv32_fs430_and0;
  assign f_arrdiv32_fs431_xor0 = f_arrdiv32_mux2to1386_xor0 ^ b[15];
  assign f_arrdiv32_fs431_not0 = ~f_arrdiv32_mux2to1386_xor0;
  assign f_arrdiv32_fs431_and0 = f_arrdiv32_fs431_not0 & b[15];
  assign f_arrdiv32_fs431_xor1 = f_arrdiv32_fs430_or0 ^ f_arrdiv32_fs431_xor0;
  assign f_arrdiv32_fs431_not1 = ~f_arrdiv32_fs431_xor0;
  assign f_arrdiv32_fs431_and1 = f_arrdiv32_fs431_not1 & f_arrdiv32_fs430_or0;
  assign f_arrdiv32_fs431_or0 = f_arrdiv32_fs431_and1 | f_arrdiv32_fs431_and0;
  assign f_arrdiv32_fs432_xor0 = f_arrdiv32_mux2to1387_xor0 ^ b[16];
  assign f_arrdiv32_fs432_not0 = ~f_arrdiv32_mux2to1387_xor0;
  assign f_arrdiv32_fs432_and0 = f_arrdiv32_fs432_not0 & b[16];
  assign f_arrdiv32_fs432_xor1 = f_arrdiv32_fs431_or0 ^ f_arrdiv32_fs432_xor0;
  assign f_arrdiv32_fs432_not1 = ~f_arrdiv32_fs432_xor0;
  assign f_arrdiv32_fs432_and1 = f_arrdiv32_fs432_not1 & f_arrdiv32_fs431_or0;
  assign f_arrdiv32_fs432_or0 = f_arrdiv32_fs432_and1 | f_arrdiv32_fs432_and0;
  assign f_arrdiv32_fs433_xor0 = f_arrdiv32_mux2to1388_xor0 ^ b[17];
  assign f_arrdiv32_fs433_not0 = ~f_arrdiv32_mux2to1388_xor0;
  assign f_arrdiv32_fs433_and0 = f_arrdiv32_fs433_not0 & b[17];
  assign f_arrdiv32_fs433_xor1 = f_arrdiv32_fs432_or0 ^ f_arrdiv32_fs433_xor0;
  assign f_arrdiv32_fs433_not1 = ~f_arrdiv32_fs433_xor0;
  assign f_arrdiv32_fs433_and1 = f_arrdiv32_fs433_not1 & f_arrdiv32_fs432_or0;
  assign f_arrdiv32_fs433_or0 = f_arrdiv32_fs433_and1 | f_arrdiv32_fs433_and0;
  assign f_arrdiv32_fs434_xor0 = f_arrdiv32_mux2to1389_xor0 ^ b[18];
  assign f_arrdiv32_fs434_not0 = ~f_arrdiv32_mux2to1389_xor0;
  assign f_arrdiv32_fs434_and0 = f_arrdiv32_fs434_not0 & b[18];
  assign f_arrdiv32_fs434_xor1 = f_arrdiv32_fs433_or0 ^ f_arrdiv32_fs434_xor0;
  assign f_arrdiv32_fs434_not1 = ~f_arrdiv32_fs434_xor0;
  assign f_arrdiv32_fs434_and1 = f_arrdiv32_fs434_not1 & f_arrdiv32_fs433_or0;
  assign f_arrdiv32_fs434_or0 = f_arrdiv32_fs434_and1 | f_arrdiv32_fs434_and0;
  assign f_arrdiv32_fs435_xor0 = f_arrdiv32_mux2to1390_xor0 ^ b[19];
  assign f_arrdiv32_fs435_not0 = ~f_arrdiv32_mux2to1390_xor0;
  assign f_arrdiv32_fs435_and0 = f_arrdiv32_fs435_not0 & b[19];
  assign f_arrdiv32_fs435_xor1 = f_arrdiv32_fs434_or0 ^ f_arrdiv32_fs435_xor0;
  assign f_arrdiv32_fs435_not1 = ~f_arrdiv32_fs435_xor0;
  assign f_arrdiv32_fs435_and1 = f_arrdiv32_fs435_not1 & f_arrdiv32_fs434_or0;
  assign f_arrdiv32_fs435_or0 = f_arrdiv32_fs435_and1 | f_arrdiv32_fs435_and0;
  assign f_arrdiv32_fs436_xor0 = f_arrdiv32_mux2to1391_xor0 ^ b[20];
  assign f_arrdiv32_fs436_not0 = ~f_arrdiv32_mux2to1391_xor0;
  assign f_arrdiv32_fs436_and0 = f_arrdiv32_fs436_not0 & b[20];
  assign f_arrdiv32_fs436_xor1 = f_arrdiv32_fs435_or0 ^ f_arrdiv32_fs436_xor0;
  assign f_arrdiv32_fs436_not1 = ~f_arrdiv32_fs436_xor0;
  assign f_arrdiv32_fs436_and1 = f_arrdiv32_fs436_not1 & f_arrdiv32_fs435_or0;
  assign f_arrdiv32_fs436_or0 = f_arrdiv32_fs436_and1 | f_arrdiv32_fs436_and0;
  assign f_arrdiv32_fs437_xor0 = f_arrdiv32_mux2to1392_xor0 ^ b[21];
  assign f_arrdiv32_fs437_not0 = ~f_arrdiv32_mux2to1392_xor0;
  assign f_arrdiv32_fs437_and0 = f_arrdiv32_fs437_not0 & b[21];
  assign f_arrdiv32_fs437_xor1 = f_arrdiv32_fs436_or0 ^ f_arrdiv32_fs437_xor0;
  assign f_arrdiv32_fs437_not1 = ~f_arrdiv32_fs437_xor0;
  assign f_arrdiv32_fs437_and1 = f_arrdiv32_fs437_not1 & f_arrdiv32_fs436_or0;
  assign f_arrdiv32_fs437_or0 = f_arrdiv32_fs437_and1 | f_arrdiv32_fs437_and0;
  assign f_arrdiv32_fs438_xor0 = f_arrdiv32_mux2to1393_xor0 ^ b[22];
  assign f_arrdiv32_fs438_not0 = ~f_arrdiv32_mux2to1393_xor0;
  assign f_arrdiv32_fs438_and0 = f_arrdiv32_fs438_not0 & b[22];
  assign f_arrdiv32_fs438_xor1 = f_arrdiv32_fs437_or0 ^ f_arrdiv32_fs438_xor0;
  assign f_arrdiv32_fs438_not1 = ~f_arrdiv32_fs438_xor0;
  assign f_arrdiv32_fs438_and1 = f_arrdiv32_fs438_not1 & f_arrdiv32_fs437_or0;
  assign f_arrdiv32_fs438_or0 = f_arrdiv32_fs438_and1 | f_arrdiv32_fs438_and0;
  assign f_arrdiv32_fs439_xor0 = f_arrdiv32_mux2to1394_xor0 ^ b[23];
  assign f_arrdiv32_fs439_not0 = ~f_arrdiv32_mux2to1394_xor0;
  assign f_arrdiv32_fs439_and0 = f_arrdiv32_fs439_not0 & b[23];
  assign f_arrdiv32_fs439_xor1 = f_arrdiv32_fs438_or0 ^ f_arrdiv32_fs439_xor0;
  assign f_arrdiv32_fs439_not1 = ~f_arrdiv32_fs439_xor0;
  assign f_arrdiv32_fs439_and1 = f_arrdiv32_fs439_not1 & f_arrdiv32_fs438_or0;
  assign f_arrdiv32_fs439_or0 = f_arrdiv32_fs439_and1 | f_arrdiv32_fs439_and0;
  assign f_arrdiv32_fs440_xor0 = f_arrdiv32_mux2to1395_xor0 ^ b[24];
  assign f_arrdiv32_fs440_not0 = ~f_arrdiv32_mux2to1395_xor0;
  assign f_arrdiv32_fs440_and0 = f_arrdiv32_fs440_not0 & b[24];
  assign f_arrdiv32_fs440_xor1 = f_arrdiv32_fs439_or0 ^ f_arrdiv32_fs440_xor0;
  assign f_arrdiv32_fs440_not1 = ~f_arrdiv32_fs440_xor0;
  assign f_arrdiv32_fs440_and1 = f_arrdiv32_fs440_not1 & f_arrdiv32_fs439_or0;
  assign f_arrdiv32_fs440_or0 = f_arrdiv32_fs440_and1 | f_arrdiv32_fs440_and0;
  assign f_arrdiv32_fs441_xor0 = f_arrdiv32_mux2to1396_xor0 ^ b[25];
  assign f_arrdiv32_fs441_not0 = ~f_arrdiv32_mux2to1396_xor0;
  assign f_arrdiv32_fs441_and0 = f_arrdiv32_fs441_not0 & b[25];
  assign f_arrdiv32_fs441_xor1 = f_arrdiv32_fs440_or0 ^ f_arrdiv32_fs441_xor0;
  assign f_arrdiv32_fs441_not1 = ~f_arrdiv32_fs441_xor0;
  assign f_arrdiv32_fs441_and1 = f_arrdiv32_fs441_not1 & f_arrdiv32_fs440_or0;
  assign f_arrdiv32_fs441_or0 = f_arrdiv32_fs441_and1 | f_arrdiv32_fs441_and0;
  assign f_arrdiv32_fs442_xor0 = f_arrdiv32_mux2to1397_xor0 ^ b[26];
  assign f_arrdiv32_fs442_not0 = ~f_arrdiv32_mux2to1397_xor0;
  assign f_arrdiv32_fs442_and0 = f_arrdiv32_fs442_not0 & b[26];
  assign f_arrdiv32_fs442_xor1 = f_arrdiv32_fs441_or0 ^ f_arrdiv32_fs442_xor0;
  assign f_arrdiv32_fs442_not1 = ~f_arrdiv32_fs442_xor0;
  assign f_arrdiv32_fs442_and1 = f_arrdiv32_fs442_not1 & f_arrdiv32_fs441_or0;
  assign f_arrdiv32_fs442_or0 = f_arrdiv32_fs442_and1 | f_arrdiv32_fs442_and0;
  assign f_arrdiv32_fs443_xor0 = f_arrdiv32_mux2to1398_xor0 ^ b[27];
  assign f_arrdiv32_fs443_not0 = ~f_arrdiv32_mux2to1398_xor0;
  assign f_arrdiv32_fs443_and0 = f_arrdiv32_fs443_not0 & b[27];
  assign f_arrdiv32_fs443_xor1 = f_arrdiv32_fs442_or0 ^ f_arrdiv32_fs443_xor0;
  assign f_arrdiv32_fs443_not1 = ~f_arrdiv32_fs443_xor0;
  assign f_arrdiv32_fs443_and1 = f_arrdiv32_fs443_not1 & f_arrdiv32_fs442_or0;
  assign f_arrdiv32_fs443_or0 = f_arrdiv32_fs443_and1 | f_arrdiv32_fs443_and0;
  assign f_arrdiv32_fs444_xor0 = f_arrdiv32_mux2to1399_xor0 ^ b[28];
  assign f_arrdiv32_fs444_not0 = ~f_arrdiv32_mux2to1399_xor0;
  assign f_arrdiv32_fs444_and0 = f_arrdiv32_fs444_not0 & b[28];
  assign f_arrdiv32_fs444_xor1 = f_arrdiv32_fs443_or0 ^ f_arrdiv32_fs444_xor0;
  assign f_arrdiv32_fs444_not1 = ~f_arrdiv32_fs444_xor0;
  assign f_arrdiv32_fs444_and1 = f_arrdiv32_fs444_not1 & f_arrdiv32_fs443_or0;
  assign f_arrdiv32_fs444_or0 = f_arrdiv32_fs444_and1 | f_arrdiv32_fs444_and0;
  assign f_arrdiv32_fs445_xor0 = f_arrdiv32_mux2to1400_xor0 ^ b[29];
  assign f_arrdiv32_fs445_not0 = ~f_arrdiv32_mux2to1400_xor0;
  assign f_arrdiv32_fs445_and0 = f_arrdiv32_fs445_not0 & b[29];
  assign f_arrdiv32_fs445_xor1 = f_arrdiv32_fs444_or0 ^ f_arrdiv32_fs445_xor0;
  assign f_arrdiv32_fs445_not1 = ~f_arrdiv32_fs445_xor0;
  assign f_arrdiv32_fs445_and1 = f_arrdiv32_fs445_not1 & f_arrdiv32_fs444_or0;
  assign f_arrdiv32_fs445_or0 = f_arrdiv32_fs445_and1 | f_arrdiv32_fs445_and0;
  assign f_arrdiv32_fs446_xor0 = f_arrdiv32_mux2to1401_xor0 ^ b[30];
  assign f_arrdiv32_fs446_not0 = ~f_arrdiv32_mux2to1401_xor0;
  assign f_arrdiv32_fs446_and0 = f_arrdiv32_fs446_not0 & b[30];
  assign f_arrdiv32_fs446_xor1 = f_arrdiv32_fs445_or0 ^ f_arrdiv32_fs446_xor0;
  assign f_arrdiv32_fs446_not1 = ~f_arrdiv32_fs446_xor0;
  assign f_arrdiv32_fs446_and1 = f_arrdiv32_fs446_not1 & f_arrdiv32_fs445_or0;
  assign f_arrdiv32_fs446_or0 = f_arrdiv32_fs446_and1 | f_arrdiv32_fs446_and0;
  assign f_arrdiv32_fs447_xor0 = f_arrdiv32_mux2to1402_xor0 ^ b[31];
  assign f_arrdiv32_fs447_not0 = ~f_arrdiv32_mux2to1402_xor0;
  assign f_arrdiv32_fs447_and0 = f_arrdiv32_fs447_not0 & b[31];
  assign f_arrdiv32_fs447_xor1 = f_arrdiv32_fs446_or0 ^ f_arrdiv32_fs447_xor0;
  assign f_arrdiv32_fs447_not1 = ~f_arrdiv32_fs447_xor0;
  assign f_arrdiv32_fs447_and1 = f_arrdiv32_fs447_not1 & f_arrdiv32_fs446_or0;
  assign f_arrdiv32_fs447_or0 = f_arrdiv32_fs447_and1 | f_arrdiv32_fs447_and0;
  assign f_arrdiv32_mux2to1403_and0 = a[18] & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1403_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1403_and1 = f_arrdiv32_fs416_xor0 & f_arrdiv32_mux2to1403_not0;
  assign f_arrdiv32_mux2to1403_xor0 = f_arrdiv32_mux2to1403_and0 ^ f_arrdiv32_mux2to1403_and1;
  assign f_arrdiv32_mux2to1404_and0 = f_arrdiv32_mux2to1372_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1404_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1404_and1 = f_arrdiv32_fs417_xor1 & f_arrdiv32_mux2to1404_not0;
  assign f_arrdiv32_mux2to1404_xor0 = f_arrdiv32_mux2to1404_and0 ^ f_arrdiv32_mux2to1404_and1;
  assign f_arrdiv32_mux2to1405_and0 = f_arrdiv32_mux2to1373_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1405_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1405_and1 = f_arrdiv32_fs418_xor1 & f_arrdiv32_mux2to1405_not0;
  assign f_arrdiv32_mux2to1405_xor0 = f_arrdiv32_mux2to1405_and0 ^ f_arrdiv32_mux2to1405_and1;
  assign f_arrdiv32_mux2to1406_and0 = f_arrdiv32_mux2to1374_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1406_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1406_and1 = f_arrdiv32_fs419_xor1 & f_arrdiv32_mux2to1406_not0;
  assign f_arrdiv32_mux2to1406_xor0 = f_arrdiv32_mux2to1406_and0 ^ f_arrdiv32_mux2to1406_and1;
  assign f_arrdiv32_mux2to1407_and0 = f_arrdiv32_mux2to1375_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1407_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1407_and1 = f_arrdiv32_fs420_xor1 & f_arrdiv32_mux2to1407_not0;
  assign f_arrdiv32_mux2to1407_xor0 = f_arrdiv32_mux2to1407_and0 ^ f_arrdiv32_mux2to1407_and1;
  assign f_arrdiv32_mux2to1408_and0 = f_arrdiv32_mux2to1376_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1408_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1408_and1 = f_arrdiv32_fs421_xor1 & f_arrdiv32_mux2to1408_not0;
  assign f_arrdiv32_mux2to1408_xor0 = f_arrdiv32_mux2to1408_and0 ^ f_arrdiv32_mux2to1408_and1;
  assign f_arrdiv32_mux2to1409_and0 = f_arrdiv32_mux2to1377_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1409_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1409_and1 = f_arrdiv32_fs422_xor1 & f_arrdiv32_mux2to1409_not0;
  assign f_arrdiv32_mux2to1409_xor0 = f_arrdiv32_mux2to1409_and0 ^ f_arrdiv32_mux2to1409_and1;
  assign f_arrdiv32_mux2to1410_and0 = f_arrdiv32_mux2to1378_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1410_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1410_and1 = f_arrdiv32_fs423_xor1 & f_arrdiv32_mux2to1410_not0;
  assign f_arrdiv32_mux2to1410_xor0 = f_arrdiv32_mux2to1410_and0 ^ f_arrdiv32_mux2to1410_and1;
  assign f_arrdiv32_mux2to1411_and0 = f_arrdiv32_mux2to1379_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1411_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1411_and1 = f_arrdiv32_fs424_xor1 & f_arrdiv32_mux2to1411_not0;
  assign f_arrdiv32_mux2to1411_xor0 = f_arrdiv32_mux2to1411_and0 ^ f_arrdiv32_mux2to1411_and1;
  assign f_arrdiv32_mux2to1412_and0 = f_arrdiv32_mux2to1380_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1412_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1412_and1 = f_arrdiv32_fs425_xor1 & f_arrdiv32_mux2to1412_not0;
  assign f_arrdiv32_mux2to1412_xor0 = f_arrdiv32_mux2to1412_and0 ^ f_arrdiv32_mux2to1412_and1;
  assign f_arrdiv32_mux2to1413_and0 = f_arrdiv32_mux2to1381_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1413_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1413_and1 = f_arrdiv32_fs426_xor1 & f_arrdiv32_mux2to1413_not0;
  assign f_arrdiv32_mux2to1413_xor0 = f_arrdiv32_mux2to1413_and0 ^ f_arrdiv32_mux2to1413_and1;
  assign f_arrdiv32_mux2to1414_and0 = f_arrdiv32_mux2to1382_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1414_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1414_and1 = f_arrdiv32_fs427_xor1 & f_arrdiv32_mux2to1414_not0;
  assign f_arrdiv32_mux2to1414_xor0 = f_arrdiv32_mux2to1414_and0 ^ f_arrdiv32_mux2to1414_and1;
  assign f_arrdiv32_mux2to1415_and0 = f_arrdiv32_mux2to1383_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1415_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1415_and1 = f_arrdiv32_fs428_xor1 & f_arrdiv32_mux2to1415_not0;
  assign f_arrdiv32_mux2to1415_xor0 = f_arrdiv32_mux2to1415_and0 ^ f_arrdiv32_mux2to1415_and1;
  assign f_arrdiv32_mux2to1416_and0 = f_arrdiv32_mux2to1384_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1416_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1416_and1 = f_arrdiv32_fs429_xor1 & f_arrdiv32_mux2to1416_not0;
  assign f_arrdiv32_mux2to1416_xor0 = f_arrdiv32_mux2to1416_and0 ^ f_arrdiv32_mux2to1416_and1;
  assign f_arrdiv32_mux2to1417_and0 = f_arrdiv32_mux2to1385_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1417_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1417_and1 = f_arrdiv32_fs430_xor1 & f_arrdiv32_mux2to1417_not0;
  assign f_arrdiv32_mux2to1417_xor0 = f_arrdiv32_mux2to1417_and0 ^ f_arrdiv32_mux2to1417_and1;
  assign f_arrdiv32_mux2to1418_and0 = f_arrdiv32_mux2to1386_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1418_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1418_and1 = f_arrdiv32_fs431_xor1 & f_arrdiv32_mux2to1418_not0;
  assign f_arrdiv32_mux2to1418_xor0 = f_arrdiv32_mux2to1418_and0 ^ f_arrdiv32_mux2to1418_and1;
  assign f_arrdiv32_mux2to1419_and0 = f_arrdiv32_mux2to1387_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1419_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1419_and1 = f_arrdiv32_fs432_xor1 & f_arrdiv32_mux2to1419_not0;
  assign f_arrdiv32_mux2to1419_xor0 = f_arrdiv32_mux2to1419_and0 ^ f_arrdiv32_mux2to1419_and1;
  assign f_arrdiv32_mux2to1420_and0 = f_arrdiv32_mux2to1388_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1420_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1420_and1 = f_arrdiv32_fs433_xor1 & f_arrdiv32_mux2to1420_not0;
  assign f_arrdiv32_mux2to1420_xor0 = f_arrdiv32_mux2to1420_and0 ^ f_arrdiv32_mux2to1420_and1;
  assign f_arrdiv32_mux2to1421_and0 = f_arrdiv32_mux2to1389_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1421_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1421_and1 = f_arrdiv32_fs434_xor1 & f_arrdiv32_mux2to1421_not0;
  assign f_arrdiv32_mux2to1421_xor0 = f_arrdiv32_mux2to1421_and0 ^ f_arrdiv32_mux2to1421_and1;
  assign f_arrdiv32_mux2to1422_and0 = f_arrdiv32_mux2to1390_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1422_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1422_and1 = f_arrdiv32_fs435_xor1 & f_arrdiv32_mux2to1422_not0;
  assign f_arrdiv32_mux2to1422_xor0 = f_arrdiv32_mux2to1422_and0 ^ f_arrdiv32_mux2to1422_and1;
  assign f_arrdiv32_mux2to1423_and0 = f_arrdiv32_mux2to1391_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1423_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1423_and1 = f_arrdiv32_fs436_xor1 & f_arrdiv32_mux2to1423_not0;
  assign f_arrdiv32_mux2to1423_xor0 = f_arrdiv32_mux2to1423_and0 ^ f_arrdiv32_mux2to1423_and1;
  assign f_arrdiv32_mux2to1424_and0 = f_arrdiv32_mux2to1392_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1424_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1424_and1 = f_arrdiv32_fs437_xor1 & f_arrdiv32_mux2to1424_not0;
  assign f_arrdiv32_mux2to1424_xor0 = f_arrdiv32_mux2to1424_and0 ^ f_arrdiv32_mux2to1424_and1;
  assign f_arrdiv32_mux2to1425_and0 = f_arrdiv32_mux2to1393_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1425_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1425_and1 = f_arrdiv32_fs438_xor1 & f_arrdiv32_mux2to1425_not0;
  assign f_arrdiv32_mux2to1425_xor0 = f_arrdiv32_mux2to1425_and0 ^ f_arrdiv32_mux2to1425_and1;
  assign f_arrdiv32_mux2to1426_and0 = f_arrdiv32_mux2to1394_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1426_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1426_and1 = f_arrdiv32_fs439_xor1 & f_arrdiv32_mux2to1426_not0;
  assign f_arrdiv32_mux2to1426_xor0 = f_arrdiv32_mux2to1426_and0 ^ f_arrdiv32_mux2to1426_and1;
  assign f_arrdiv32_mux2to1427_and0 = f_arrdiv32_mux2to1395_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1427_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1427_and1 = f_arrdiv32_fs440_xor1 & f_arrdiv32_mux2to1427_not0;
  assign f_arrdiv32_mux2to1427_xor0 = f_arrdiv32_mux2to1427_and0 ^ f_arrdiv32_mux2to1427_and1;
  assign f_arrdiv32_mux2to1428_and0 = f_arrdiv32_mux2to1396_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1428_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1428_and1 = f_arrdiv32_fs441_xor1 & f_arrdiv32_mux2to1428_not0;
  assign f_arrdiv32_mux2to1428_xor0 = f_arrdiv32_mux2to1428_and0 ^ f_arrdiv32_mux2to1428_and1;
  assign f_arrdiv32_mux2to1429_and0 = f_arrdiv32_mux2to1397_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1429_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1429_and1 = f_arrdiv32_fs442_xor1 & f_arrdiv32_mux2to1429_not0;
  assign f_arrdiv32_mux2to1429_xor0 = f_arrdiv32_mux2to1429_and0 ^ f_arrdiv32_mux2to1429_and1;
  assign f_arrdiv32_mux2to1430_and0 = f_arrdiv32_mux2to1398_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1430_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1430_and1 = f_arrdiv32_fs443_xor1 & f_arrdiv32_mux2to1430_not0;
  assign f_arrdiv32_mux2to1430_xor0 = f_arrdiv32_mux2to1430_and0 ^ f_arrdiv32_mux2to1430_and1;
  assign f_arrdiv32_mux2to1431_and0 = f_arrdiv32_mux2to1399_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1431_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1431_and1 = f_arrdiv32_fs444_xor1 & f_arrdiv32_mux2to1431_not0;
  assign f_arrdiv32_mux2to1431_xor0 = f_arrdiv32_mux2to1431_and0 ^ f_arrdiv32_mux2to1431_and1;
  assign f_arrdiv32_mux2to1432_and0 = f_arrdiv32_mux2to1400_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1432_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1432_and1 = f_arrdiv32_fs445_xor1 & f_arrdiv32_mux2to1432_not0;
  assign f_arrdiv32_mux2to1432_xor0 = f_arrdiv32_mux2to1432_and0 ^ f_arrdiv32_mux2to1432_and1;
  assign f_arrdiv32_mux2to1433_and0 = f_arrdiv32_mux2to1401_xor0 & f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1433_not0 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_mux2to1433_and1 = f_arrdiv32_fs446_xor1 & f_arrdiv32_mux2to1433_not0;
  assign f_arrdiv32_mux2to1433_xor0 = f_arrdiv32_mux2to1433_and0 ^ f_arrdiv32_mux2to1433_and1;
  assign f_arrdiv32_not13 = ~f_arrdiv32_fs447_or0;
  assign f_arrdiv32_fs448_xor0 = a[17] ^ b[0];
  assign f_arrdiv32_fs448_not0 = ~a[17];
  assign f_arrdiv32_fs448_and0 = f_arrdiv32_fs448_not0 & b[0];
  assign f_arrdiv32_fs448_not1 = ~f_arrdiv32_fs448_xor0;
  assign f_arrdiv32_fs449_xor0 = f_arrdiv32_mux2to1403_xor0 ^ b[1];
  assign f_arrdiv32_fs449_not0 = ~f_arrdiv32_mux2to1403_xor0;
  assign f_arrdiv32_fs449_and0 = f_arrdiv32_fs449_not0 & b[1];
  assign f_arrdiv32_fs449_xor1 = f_arrdiv32_fs448_and0 ^ f_arrdiv32_fs449_xor0;
  assign f_arrdiv32_fs449_not1 = ~f_arrdiv32_fs449_xor0;
  assign f_arrdiv32_fs449_and1 = f_arrdiv32_fs449_not1 & f_arrdiv32_fs448_and0;
  assign f_arrdiv32_fs449_or0 = f_arrdiv32_fs449_and1 | f_arrdiv32_fs449_and0;
  assign f_arrdiv32_fs450_xor0 = f_arrdiv32_mux2to1404_xor0 ^ b[2];
  assign f_arrdiv32_fs450_not0 = ~f_arrdiv32_mux2to1404_xor0;
  assign f_arrdiv32_fs450_and0 = f_arrdiv32_fs450_not0 & b[2];
  assign f_arrdiv32_fs450_xor1 = f_arrdiv32_fs449_or0 ^ f_arrdiv32_fs450_xor0;
  assign f_arrdiv32_fs450_not1 = ~f_arrdiv32_fs450_xor0;
  assign f_arrdiv32_fs450_and1 = f_arrdiv32_fs450_not1 & f_arrdiv32_fs449_or0;
  assign f_arrdiv32_fs450_or0 = f_arrdiv32_fs450_and1 | f_arrdiv32_fs450_and0;
  assign f_arrdiv32_fs451_xor0 = f_arrdiv32_mux2to1405_xor0 ^ b[3];
  assign f_arrdiv32_fs451_not0 = ~f_arrdiv32_mux2to1405_xor0;
  assign f_arrdiv32_fs451_and0 = f_arrdiv32_fs451_not0 & b[3];
  assign f_arrdiv32_fs451_xor1 = f_arrdiv32_fs450_or0 ^ f_arrdiv32_fs451_xor0;
  assign f_arrdiv32_fs451_not1 = ~f_arrdiv32_fs451_xor0;
  assign f_arrdiv32_fs451_and1 = f_arrdiv32_fs451_not1 & f_arrdiv32_fs450_or0;
  assign f_arrdiv32_fs451_or0 = f_arrdiv32_fs451_and1 | f_arrdiv32_fs451_and0;
  assign f_arrdiv32_fs452_xor0 = f_arrdiv32_mux2to1406_xor0 ^ b[4];
  assign f_arrdiv32_fs452_not0 = ~f_arrdiv32_mux2to1406_xor0;
  assign f_arrdiv32_fs452_and0 = f_arrdiv32_fs452_not0 & b[4];
  assign f_arrdiv32_fs452_xor1 = f_arrdiv32_fs451_or0 ^ f_arrdiv32_fs452_xor0;
  assign f_arrdiv32_fs452_not1 = ~f_arrdiv32_fs452_xor0;
  assign f_arrdiv32_fs452_and1 = f_arrdiv32_fs452_not1 & f_arrdiv32_fs451_or0;
  assign f_arrdiv32_fs452_or0 = f_arrdiv32_fs452_and1 | f_arrdiv32_fs452_and0;
  assign f_arrdiv32_fs453_xor0 = f_arrdiv32_mux2to1407_xor0 ^ b[5];
  assign f_arrdiv32_fs453_not0 = ~f_arrdiv32_mux2to1407_xor0;
  assign f_arrdiv32_fs453_and0 = f_arrdiv32_fs453_not0 & b[5];
  assign f_arrdiv32_fs453_xor1 = f_arrdiv32_fs452_or0 ^ f_arrdiv32_fs453_xor0;
  assign f_arrdiv32_fs453_not1 = ~f_arrdiv32_fs453_xor0;
  assign f_arrdiv32_fs453_and1 = f_arrdiv32_fs453_not1 & f_arrdiv32_fs452_or0;
  assign f_arrdiv32_fs453_or0 = f_arrdiv32_fs453_and1 | f_arrdiv32_fs453_and0;
  assign f_arrdiv32_fs454_xor0 = f_arrdiv32_mux2to1408_xor0 ^ b[6];
  assign f_arrdiv32_fs454_not0 = ~f_arrdiv32_mux2to1408_xor0;
  assign f_arrdiv32_fs454_and0 = f_arrdiv32_fs454_not0 & b[6];
  assign f_arrdiv32_fs454_xor1 = f_arrdiv32_fs453_or0 ^ f_arrdiv32_fs454_xor0;
  assign f_arrdiv32_fs454_not1 = ~f_arrdiv32_fs454_xor0;
  assign f_arrdiv32_fs454_and1 = f_arrdiv32_fs454_not1 & f_arrdiv32_fs453_or0;
  assign f_arrdiv32_fs454_or0 = f_arrdiv32_fs454_and1 | f_arrdiv32_fs454_and0;
  assign f_arrdiv32_fs455_xor0 = f_arrdiv32_mux2to1409_xor0 ^ b[7];
  assign f_arrdiv32_fs455_not0 = ~f_arrdiv32_mux2to1409_xor0;
  assign f_arrdiv32_fs455_and0 = f_arrdiv32_fs455_not0 & b[7];
  assign f_arrdiv32_fs455_xor1 = f_arrdiv32_fs454_or0 ^ f_arrdiv32_fs455_xor0;
  assign f_arrdiv32_fs455_not1 = ~f_arrdiv32_fs455_xor0;
  assign f_arrdiv32_fs455_and1 = f_arrdiv32_fs455_not1 & f_arrdiv32_fs454_or0;
  assign f_arrdiv32_fs455_or0 = f_arrdiv32_fs455_and1 | f_arrdiv32_fs455_and0;
  assign f_arrdiv32_fs456_xor0 = f_arrdiv32_mux2to1410_xor0 ^ b[8];
  assign f_arrdiv32_fs456_not0 = ~f_arrdiv32_mux2to1410_xor0;
  assign f_arrdiv32_fs456_and0 = f_arrdiv32_fs456_not0 & b[8];
  assign f_arrdiv32_fs456_xor1 = f_arrdiv32_fs455_or0 ^ f_arrdiv32_fs456_xor0;
  assign f_arrdiv32_fs456_not1 = ~f_arrdiv32_fs456_xor0;
  assign f_arrdiv32_fs456_and1 = f_arrdiv32_fs456_not1 & f_arrdiv32_fs455_or0;
  assign f_arrdiv32_fs456_or0 = f_arrdiv32_fs456_and1 | f_arrdiv32_fs456_and0;
  assign f_arrdiv32_fs457_xor0 = f_arrdiv32_mux2to1411_xor0 ^ b[9];
  assign f_arrdiv32_fs457_not0 = ~f_arrdiv32_mux2to1411_xor0;
  assign f_arrdiv32_fs457_and0 = f_arrdiv32_fs457_not0 & b[9];
  assign f_arrdiv32_fs457_xor1 = f_arrdiv32_fs456_or0 ^ f_arrdiv32_fs457_xor0;
  assign f_arrdiv32_fs457_not1 = ~f_arrdiv32_fs457_xor0;
  assign f_arrdiv32_fs457_and1 = f_arrdiv32_fs457_not1 & f_arrdiv32_fs456_or0;
  assign f_arrdiv32_fs457_or0 = f_arrdiv32_fs457_and1 | f_arrdiv32_fs457_and0;
  assign f_arrdiv32_fs458_xor0 = f_arrdiv32_mux2to1412_xor0 ^ b[10];
  assign f_arrdiv32_fs458_not0 = ~f_arrdiv32_mux2to1412_xor0;
  assign f_arrdiv32_fs458_and0 = f_arrdiv32_fs458_not0 & b[10];
  assign f_arrdiv32_fs458_xor1 = f_arrdiv32_fs457_or0 ^ f_arrdiv32_fs458_xor0;
  assign f_arrdiv32_fs458_not1 = ~f_arrdiv32_fs458_xor0;
  assign f_arrdiv32_fs458_and1 = f_arrdiv32_fs458_not1 & f_arrdiv32_fs457_or0;
  assign f_arrdiv32_fs458_or0 = f_arrdiv32_fs458_and1 | f_arrdiv32_fs458_and0;
  assign f_arrdiv32_fs459_xor0 = f_arrdiv32_mux2to1413_xor0 ^ b[11];
  assign f_arrdiv32_fs459_not0 = ~f_arrdiv32_mux2to1413_xor0;
  assign f_arrdiv32_fs459_and0 = f_arrdiv32_fs459_not0 & b[11];
  assign f_arrdiv32_fs459_xor1 = f_arrdiv32_fs458_or0 ^ f_arrdiv32_fs459_xor0;
  assign f_arrdiv32_fs459_not1 = ~f_arrdiv32_fs459_xor0;
  assign f_arrdiv32_fs459_and1 = f_arrdiv32_fs459_not1 & f_arrdiv32_fs458_or0;
  assign f_arrdiv32_fs459_or0 = f_arrdiv32_fs459_and1 | f_arrdiv32_fs459_and0;
  assign f_arrdiv32_fs460_xor0 = f_arrdiv32_mux2to1414_xor0 ^ b[12];
  assign f_arrdiv32_fs460_not0 = ~f_arrdiv32_mux2to1414_xor0;
  assign f_arrdiv32_fs460_and0 = f_arrdiv32_fs460_not0 & b[12];
  assign f_arrdiv32_fs460_xor1 = f_arrdiv32_fs459_or0 ^ f_arrdiv32_fs460_xor0;
  assign f_arrdiv32_fs460_not1 = ~f_arrdiv32_fs460_xor0;
  assign f_arrdiv32_fs460_and1 = f_arrdiv32_fs460_not1 & f_arrdiv32_fs459_or0;
  assign f_arrdiv32_fs460_or0 = f_arrdiv32_fs460_and1 | f_arrdiv32_fs460_and0;
  assign f_arrdiv32_fs461_xor0 = f_arrdiv32_mux2to1415_xor0 ^ b[13];
  assign f_arrdiv32_fs461_not0 = ~f_arrdiv32_mux2to1415_xor0;
  assign f_arrdiv32_fs461_and0 = f_arrdiv32_fs461_not0 & b[13];
  assign f_arrdiv32_fs461_xor1 = f_arrdiv32_fs460_or0 ^ f_arrdiv32_fs461_xor0;
  assign f_arrdiv32_fs461_not1 = ~f_arrdiv32_fs461_xor0;
  assign f_arrdiv32_fs461_and1 = f_arrdiv32_fs461_not1 & f_arrdiv32_fs460_or0;
  assign f_arrdiv32_fs461_or0 = f_arrdiv32_fs461_and1 | f_arrdiv32_fs461_and0;
  assign f_arrdiv32_fs462_xor0 = f_arrdiv32_mux2to1416_xor0 ^ b[14];
  assign f_arrdiv32_fs462_not0 = ~f_arrdiv32_mux2to1416_xor0;
  assign f_arrdiv32_fs462_and0 = f_arrdiv32_fs462_not0 & b[14];
  assign f_arrdiv32_fs462_xor1 = f_arrdiv32_fs461_or0 ^ f_arrdiv32_fs462_xor0;
  assign f_arrdiv32_fs462_not1 = ~f_arrdiv32_fs462_xor0;
  assign f_arrdiv32_fs462_and1 = f_arrdiv32_fs462_not1 & f_arrdiv32_fs461_or0;
  assign f_arrdiv32_fs462_or0 = f_arrdiv32_fs462_and1 | f_arrdiv32_fs462_and0;
  assign f_arrdiv32_fs463_xor0 = f_arrdiv32_mux2to1417_xor0 ^ b[15];
  assign f_arrdiv32_fs463_not0 = ~f_arrdiv32_mux2to1417_xor0;
  assign f_arrdiv32_fs463_and0 = f_arrdiv32_fs463_not0 & b[15];
  assign f_arrdiv32_fs463_xor1 = f_arrdiv32_fs462_or0 ^ f_arrdiv32_fs463_xor0;
  assign f_arrdiv32_fs463_not1 = ~f_arrdiv32_fs463_xor0;
  assign f_arrdiv32_fs463_and1 = f_arrdiv32_fs463_not1 & f_arrdiv32_fs462_or0;
  assign f_arrdiv32_fs463_or0 = f_arrdiv32_fs463_and1 | f_arrdiv32_fs463_and0;
  assign f_arrdiv32_fs464_xor0 = f_arrdiv32_mux2to1418_xor0 ^ b[16];
  assign f_arrdiv32_fs464_not0 = ~f_arrdiv32_mux2to1418_xor0;
  assign f_arrdiv32_fs464_and0 = f_arrdiv32_fs464_not0 & b[16];
  assign f_arrdiv32_fs464_xor1 = f_arrdiv32_fs463_or0 ^ f_arrdiv32_fs464_xor0;
  assign f_arrdiv32_fs464_not1 = ~f_arrdiv32_fs464_xor0;
  assign f_arrdiv32_fs464_and1 = f_arrdiv32_fs464_not1 & f_arrdiv32_fs463_or0;
  assign f_arrdiv32_fs464_or0 = f_arrdiv32_fs464_and1 | f_arrdiv32_fs464_and0;
  assign f_arrdiv32_fs465_xor0 = f_arrdiv32_mux2to1419_xor0 ^ b[17];
  assign f_arrdiv32_fs465_not0 = ~f_arrdiv32_mux2to1419_xor0;
  assign f_arrdiv32_fs465_and0 = f_arrdiv32_fs465_not0 & b[17];
  assign f_arrdiv32_fs465_xor1 = f_arrdiv32_fs464_or0 ^ f_arrdiv32_fs465_xor0;
  assign f_arrdiv32_fs465_not1 = ~f_arrdiv32_fs465_xor0;
  assign f_arrdiv32_fs465_and1 = f_arrdiv32_fs465_not1 & f_arrdiv32_fs464_or0;
  assign f_arrdiv32_fs465_or0 = f_arrdiv32_fs465_and1 | f_arrdiv32_fs465_and0;
  assign f_arrdiv32_fs466_xor0 = f_arrdiv32_mux2to1420_xor0 ^ b[18];
  assign f_arrdiv32_fs466_not0 = ~f_arrdiv32_mux2to1420_xor0;
  assign f_arrdiv32_fs466_and0 = f_arrdiv32_fs466_not0 & b[18];
  assign f_arrdiv32_fs466_xor1 = f_arrdiv32_fs465_or0 ^ f_arrdiv32_fs466_xor0;
  assign f_arrdiv32_fs466_not1 = ~f_arrdiv32_fs466_xor0;
  assign f_arrdiv32_fs466_and1 = f_arrdiv32_fs466_not1 & f_arrdiv32_fs465_or0;
  assign f_arrdiv32_fs466_or0 = f_arrdiv32_fs466_and1 | f_arrdiv32_fs466_and0;
  assign f_arrdiv32_fs467_xor0 = f_arrdiv32_mux2to1421_xor0 ^ b[19];
  assign f_arrdiv32_fs467_not0 = ~f_arrdiv32_mux2to1421_xor0;
  assign f_arrdiv32_fs467_and0 = f_arrdiv32_fs467_not0 & b[19];
  assign f_arrdiv32_fs467_xor1 = f_arrdiv32_fs466_or0 ^ f_arrdiv32_fs467_xor0;
  assign f_arrdiv32_fs467_not1 = ~f_arrdiv32_fs467_xor0;
  assign f_arrdiv32_fs467_and1 = f_arrdiv32_fs467_not1 & f_arrdiv32_fs466_or0;
  assign f_arrdiv32_fs467_or0 = f_arrdiv32_fs467_and1 | f_arrdiv32_fs467_and0;
  assign f_arrdiv32_fs468_xor0 = f_arrdiv32_mux2to1422_xor0 ^ b[20];
  assign f_arrdiv32_fs468_not0 = ~f_arrdiv32_mux2to1422_xor0;
  assign f_arrdiv32_fs468_and0 = f_arrdiv32_fs468_not0 & b[20];
  assign f_arrdiv32_fs468_xor1 = f_arrdiv32_fs467_or0 ^ f_arrdiv32_fs468_xor0;
  assign f_arrdiv32_fs468_not1 = ~f_arrdiv32_fs468_xor0;
  assign f_arrdiv32_fs468_and1 = f_arrdiv32_fs468_not1 & f_arrdiv32_fs467_or0;
  assign f_arrdiv32_fs468_or0 = f_arrdiv32_fs468_and1 | f_arrdiv32_fs468_and0;
  assign f_arrdiv32_fs469_xor0 = f_arrdiv32_mux2to1423_xor0 ^ b[21];
  assign f_arrdiv32_fs469_not0 = ~f_arrdiv32_mux2to1423_xor0;
  assign f_arrdiv32_fs469_and0 = f_arrdiv32_fs469_not0 & b[21];
  assign f_arrdiv32_fs469_xor1 = f_arrdiv32_fs468_or0 ^ f_arrdiv32_fs469_xor0;
  assign f_arrdiv32_fs469_not1 = ~f_arrdiv32_fs469_xor0;
  assign f_arrdiv32_fs469_and1 = f_arrdiv32_fs469_not1 & f_arrdiv32_fs468_or0;
  assign f_arrdiv32_fs469_or0 = f_arrdiv32_fs469_and1 | f_arrdiv32_fs469_and0;
  assign f_arrdiv32_fs470_xor0 = f_arrdiv32_mux2to1424_xor0 ^ b[22];
  assign f_arrdiv32_fs470_not0 = ~f_arrdiv32_mux2to1424_xor0;
  assign f_arrdiv32_fs470_and0 = f_arrdiv32_fs470_not0 & b[22];
  assign f_arrdiv32_fs470_xor1 = f_arrdiv32_fs469_or0 ^ f_arrdiv32_fs470_xor0;
  assign f_arrdiv32_fs470_not1 = ~f_arrdiv32_fs470_xor0;
  assign f_arrdiv32_fs470_and1 = f_arrdiv32_fs470_not1 & f_arrdiv32_fs469_or0;
  assign f_arrdiv32_fs470_or0 = f_arrdiv32_fs470_and1 | f_arrdiv32_fs470_and0;
  assign f_arrdiv32_fs471_xor0 = f_arrdiv32_mux2to1425_xor0 ^ b[23];
  assign f_arrdiv32_fs471_not0 = ~f_arrdiv32_mux2to1425_xor0;
  assign f_arrdiv32_fs471_and0 = f_arrdiv32_fs471_not0 & b[23];
  assign f_arrdiv32_fs471_xor1 = f_arrdiv32_fs470_or0 ^ f_arrdiv32_fs471_xor0;
  assign f_arrdiv32_fs471_not1 = ~f_arrdiv32_fs471_xor0;
  assign f_arrdiv32_fs471_and1 = f_arrdiv32_fs471_not1 & f_arrdiv32_fs470_or0;
  assign f_arrdiv32_fs471_or0 = f_arrdiv32_fs471_and1 | f_arrdiv32_fs471_and0;
  assign f_arrdiv32_fs472_xor0 = f_arrdiv32_mux2to1426_xor0 ^ b[24];
  assign f_arrdiv32_fs472_not0 = ~f_arrdiv32_mux2to1426_xor0;
  assign f_arrdiv32_fs472_and0 = f_arrdiv32_fs472_not0 & b[24];
  assign f_arrdiv32_fs472_xor1 = f_arrdiv32_fs471_or0 ^ f_arrdiv32_fs472_xor0;
  assign f_arrdiv32_fs472_not1 = ~f_arrdiv32_fs472_xor0;
  assign f_arrdiv32_fs472_and1 = f_arrdiv32_fs472_not1 & f_arrdiv32_fs471_or0;
  assign f_arrdiv32_fs472_or0 = f_arrdiv32_fs472_and1 | f_arrdiv32_fs472_and0;
  assign f_arrdiv32_fs473_xor0 = f_arrdiv32_mux2to1427_xor0 ^ b[25];
  assign f_arrdiv32_fs473_not0 = ~f_arrdiv32_mux2to1427_xor0;
  assign f_arrdiv32_fs473_and0 = f_arrdiv32_fs473_not0 & b[25];
  assign f_arrdiv32_fs473_xor1 = f_arrdiv32_fs472_or0 ^ f_arrdiv32_fs473_xor0;
  assign f_arrdiv32_fs473_not1 = ~f_arrdiv32_fs473_xor0;
  assign f_arrdiv32_fs473_and1 = f_arrdiv32_fs473_not1 & f_arrdiv32_fs472_or0;
  assign f_arrdiv32_fs473_or0 = f_arrdiv32_fs473_and1 | f_arrdiv32_fs473_and0;
  assign f_arrdiv32_fs474_xor0 = f_arrdiv32_mux2to1428_xor0 ^ b[26];
  assign f_arrdiv32_fs474_not0 = ~f_arrdiv32_mux2to1428_xor0;
  assign f_arrdiv32_fs474_and0 = f_arrdiv32_fs474_not0 & b[26];
  assign f_arrdiv32_fs474_xor1 = f_arrdiv32_fs473_or0 ^ f_arrdiv32_fs474_xor0;
  assign f_arrdiv32_fs474_not1 = ~f_arrdiv32_fs474_xor0;
  assign f_arrdiv32_fs474_and1 = f_arrdiv32_fs474_not1 & f_arrdiv32_fs473_or0;
  assign f_arrdiv32_fs474_or0 = f_arrdiv32_fs474_and1 | f_arrdiv32_fs474_and0;
  assign f_arrdiv32_fs475_xor0 = f_arrdiv32_mux2to1429_xor0 ^ b[27];
  assign f_arrdiv32_fs475_not0 = ~f_arrdiv32_mux2to1429_xor0;
  assign f_arrdiv32_fs475_and0 = f_arrdiv32_fs475_not0 & b[27];
  assign f_arrdiv32_fs475_xor1 = f_arrdiv32_fs474_or0 ^ f_arrdiv32_fs475_xor0;
  assign f_arrdiv32_fs475_not1 = ~f_arrdiv32_fs475_xor0;
  assign f_arrdiv32_fs475_and1 = f_arrdiv32_fs475_not1 & f_arrdiv32_fs474_or0;
  assign f_arrdiv32_fs475_or0 = f_arrdiv32_fs475_and1 | f_arrdiv32_fs475_and0;
  assign f_arrdiv32_fs476_xor0 = f_arrdiv32_mux2to1430_xor0 ^ b[28];
  assign f_arrdiv32_fs476_not0 = ~f_arrdiv32_mux2to1430_xor0;
  assign f_arrdiv32_fs476_and0 = f_arrdiv32_fs476_not0 & b[28];
  assign f_arrdiv32_fs476_xor1 = f_arrdiv32_fs475_or0 ^ f_arrdiv32_fs476_xor0;
  assign f_arrdiv32_fs476_not1 = ~f_arrdiv32_fs476_xor0;
  assign f_arrdiv32_fs476_and1 = f_arrdiv32_fs476_not1 & f_arrdiv32_fs475_or0;
  assign f_arrdiv32_fs476_or0 = f_arrdiv32_fs476_and1 | f_arrdiv32_fs476_and0;
  assign f_arrdiv32_fs477_xor0 = f_arrdiv32_mux2to1431_xor0 ^ b[29];
  assign f_arrdiv32_fs477_not0 = ~f_arrdiv32_mux2to1431_xor0;
  assign f_arrdiv32_fs477_and0 = f_arrdiv32_fs477_not0 & b[29];
  assign f_arrdiv32_fs477_xor1 = f_arrdiv32_fs476_or0 ^ f_arrdiv32_fs477_xor0;
  assign f_arrdiv32_fs477_not1 = ~f_arrdiv32_fs477_xor0;
  assign f_arrdiv32_fs477_and1 = f_arrdiv32_fs477_not1 & f_arrdiv32_fs476_or0;
  assign f_arrdiv32_fs477_or0 = f_arrdiv32_fs477_and1 | f_arrdiv32_fs477_and0;
  assign f_arrdiv32_fs478_xor0 = f_arrdiv32_mux2to1432_xor0 ^ b[30];
  assign f_arrdiv32_fs478_not0 = ~f_arrdiv32_mux2to1432_xor0;
  assign f_arrdiv32_fs478_and0 = f_arrdiv32_fs478_not0 & b[30];
  assign f_arrdiv32_fs478_xor1 = f_arrdiv32_fs477_or0 ^ f_arrdiv32_fs478_xor0;
  assign f_arrdiv32_fs478_not1 = ~f_arrdiv32_fs478_xor0;
  assign f_arrdiv32_fs478_and1 = f_arrdiv32_fs478_not1 & f_arrdiv32_fs477_or0;
  assign f_arrdiv32_fs478_or0 = f_arrdiv32_fs478_and1 | f_arrdiv32_fs478_and0;
  assign f_arrdiv32_fs479_xor0 = f_arrdiv32_mux2to1433_xor0 ^ b[31];
  assign f_arrdiv32_fs479_not0 = ~f_arrdiv32_mux2to1433_xor0;
  assign f_arrdiv32_fs479_and0 = f_arrdiv32_fs479_not0 & b[31];
  assign f_arrdiv32_fs479_xor1 = f_arrdiv32_fs478_or0 ^ f_arrdiv32_fs479_xor0;
  assign f_arrdiv32_fs479_not1 = ~f_arrdiv32_fs479_xor0;
  assign f_arrdiv32_fs479_and1 = f_arrdiv32_fs479_not1 & f_arrdiv32_fs478_or0;
  assign f_arrdiv32_fs479_or0 = f_arrdiv32_fs479_and1 | f_arrdiv32_fs479_and0;
  assign f_arrdiv32_mux2to1434_and0 = a[17] & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1434_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1434_and1 = f_arrdiv32_fs448_xor0 & f_arrdiv32_mux2to1434_not0;
  assign f_arrdiv32_mux2to1434_xor0 = f_arrdiv32_mux2to1434_and0 ^ f_arrdiv32_mux2to1434_and1;
  assign f_arrdiv32_mux2to1435_and0 = f_arrdiv32_mux2to1403_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1435_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1435_and1 = f_arrdiv32_fs449_xor1 & f_arrdiv32_mux2to1435_not0;
  assign f_arrdiv32_mux2to1435_xor0 = f_arrdiv32_mux2to1435_and0 ^ f_arrdiv32_mux2to1435_and1;
  assign f_arrdiv32_mux2to1436_and0 = f_arrdiv32_mux2to1404_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1436_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1436_and1 = f_arrdiv32_fs450_xor1 & f_arrdiv32_mux2to1436_not0;
  assign f_arrdiv32_mux2to1436_xor0 = f_arrdiv32_mux2to1436_and0 ^ f_arrdiv32_mux2to1436_and1;
  assign f_arrdiv32_mux2to1437_and0 = f_arrdiv32_mux2to1405_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1437_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1437_and1 = f_arrdiv32_fs451_xor1 & f_arrdiv32_mux2to1437_not0;
  assign f_arrdiv32_mux2to1437_xor0 = f_arrdiv32_mux2to1437_and0 ^ f_arrdiv32_mux2to1437_and1;
  assign f_arrdiv32_mux2to1438_and0 = f_arrdiv32_mux2to1406_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1438_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1438_and1 = f_arrdiv32_fs452_xor1 & f_arrdiv32_mux2to1438_not0;
  assign f_arrdiv32_mux2to1438_xor0 = f_arrdiv32_mux2to1438_and0 ^ f_arrdiv32_mux2to1438_and1;
  assign f_arrdiv32_mux2to1439_and0 = f_arrdiv32_mux2to1407_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1439_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1439_and1 = f_arrdiv32_fs453_xor1 & f_arrdiv32_mux2to1439_not0;
  assign f_arrdiv32_mux2to1439_xor0 = f_arrdiv32_mux2to1439_and0 ^ f_arrdiv32_mux2to1439_and1;
  assign f_arrdiv32_mux2to1440_and0 = f_arrdiv32_mux2to1408_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1440_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1440_and1 = f_arrdiv32_fs454_xor1 & f_arrdiv32_mux2to1440_not0;
  assign f_arrdiv32_mux2to1440_xor0 = f_arrdiv32_mux2to1440_and0 ^ f_arrdiv32_mux2to1440_and1;
  assign f_arrdiv32_mux2to1441_and0 = f_arrdiv32_mux2to1409_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1441_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1441_and1 = f_arrdiv32_fs455_xor1 & f_arrdiv32_mux2to1441_not0;
  assign f_arrdiv32_mux2to1441_xor0 = f_arrdiv32_mux2to1441_and0 ^ f_arrdiv32_mux2to1441_and1;
  assign f_arrdiv32_mux2to1442_and0 = f_arrdiv32_mux2to1410_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1442_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1442_and1 = f_arrdiv32_fs456_xor1 & f_arrdiv32_mux2to1442_not0;
  assign f_arrdiv32_mux2to1442_xor0 = f_arrdiv32_mux2to1442_and0 ^ f_arrdiv32_mux2to1442_and1;
  assign f_arrdiv32_mux2to1443_and0 = f_arrdiv32_mux2to1411_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1443_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1443_and1 = f_arrdiv32_fs457_xor1 & f_arrdiv32_mux2to1443_not0;
  assign f_arrdiv32_mux2to1443_xor0 = f_arrdiv32_mux2to1443_and0 ^ f_arrdiv32_mux2to1443_and1;
  assign f_arrdiv32_mux2to1444_and0 = f_arrdiv32_mux2to1412_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1444_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1444_and1 = f_arrdiv32_fs458_xor1 & f_arrdiv32_mux2to1444_not0;
  assign f_arrdiv32_mux2to1444_xor0 = f_arrdiv32_mux2to1444_and0 ^ f_arrdiv32_mux2to1444_and1;
  assign f_arrdiv32_mux2to1445_and0 = f_arrdiv32_mux2to1413_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1445_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1445_and1 = f_arrdiv32_fs459_xor1 & f_arrdiv32_mux2to1445_not0;
  assign f_arrdiv32_mux2to1445_xor0 = f_arrdiv32_mux2to1445_and0 ^ f_arrdiv32_mux2to1445_and1;
  assign f_arrdiv32_mux2to1446_and0 = f_arrdiv32_mux2to1414_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1446_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1446_and1 = f_arrdiv32_fs460_xor1 & f_arrdiv32_mux2to1446_not0;
  assign f_arrdiv32_mux2to1446_xor0 = f_arrdiv32_mux2to1446_and0 ^ f_arrdiv32_mux2to1446_and1;
  assign f_arrdiv32_mux2to1447_and0 = f_arrdiv32_mux2to1415_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1447_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1447_and1 = f_arrdiv32_fs461_xor1 & f_arrdiv32_mux2to1447_not0;
  assign f_arrdiv32_mux2to1447_xor0 = f_arrdiv32_mux2to1447_and0 ^ f_arrdiv32_mux2to1447_and1;
  assign f_arrdiv32_mux2to1448_and0 = f_arrdiv32_mux2to1416_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1448_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1448_and1 = f_arrdiv32_fs462_xor1 & f_arrdiv32_mux2to1448_not0;
  assign f_arrdiv32_mux2to1448_xor0 = f_arrdiv32_mux2to1448_and0 ^ f_arrdiv32_mux2to1448_and1;
  assign f_arrdiv32_mux2to1449_and0 = f_arrdiv32_mux2to1417_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1449_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1449_and1 = f_arrdiv32_fs463_xor1 & f_arrdiv32_mux2to1449_not0;
  assign f_arrdiv32_mux2to1449_xor0 = f_arrdiv32_mux2to1449_and0 ^ f_arrdiv32_mux2to1449_and1;
  assign f_arrdiv32_mux2to1450_and0 = f_arrdiv32_mux2to1418_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1450_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1450_and1 = f_arrdiv32_fs464_xor1 & f_arrdiv32_mux2to1450_not0;
  assign f_arrdiv32_mux2to1450_xor0 = f_arrdiv32_mux2to1450_and0 ^ f_arrdiv32_mux2to1450_and1;
  assign f_arrdiv32_mux2to1451_and0 = f_arrdiv32_mux2to1419_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1451_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1451_and1 = f_arrdiv32_fs465_xor1 & f_arrdiv32_mux2to1451_not0;
  assign f_arrdiv32_mux2to1451_xor0 = f_arrdiv32_mux2to1451_and0 ^ f_arrdiv32_mux2to1451_and1;
  assign f_arrdiv32_mux2to1452_and0 = f_arrdiv32_mux2to1420_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1452_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1452_and1 = f_arrdiv32_fs466_xor1 & f_arrdiv32_mux2to1452_not0;
  assign f_arrdiv32_mux2to1452_xor0 = f_arrdiv32_mux2to1452_and0 ^ f_arrdiv32_mux2to1452_and1;
  assign f_arrdiv32_mux2to1453_and0 = f_arrdiv32_mux2to1421_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1453_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1453_and1 = f_arrdiv32_fs467_xor1 & f_arrdiv32_mux2to1453_not0;
  assign f_arrdiv32_mux2to1453_xor0 = f_arrdiv32_mux2to1453_and0 ^ f_arrdiv32_mux2to1453_and1;
  assign f_arrdiv32_mux2to1454_and0 = f_arrdiv32_mux2to1422_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1454_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1454_and1 = f_arrdiv32_fs468_xor1 & f_arrdiv32_mux2to1454_not0;
  assign f_arrdiv32_mux2to1454_xor0 = f_arrdiv32_mux2to1454_and0 ^ f_arrdiv32_mux2to1454_and1;
  assign f_arrdiv32_mux2to1455_and0 = f_arrdiv32_mux2to1423_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1455_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1455_and1 = f_arrdiv32_fs469_xor1 & f_arrdiv32_mux2to1455_not0;
  assign f_arrdiv32_mux2to1455_xor0 = f_arrdiv32_mux2to1455_and0 ^ f_arrdiv32_mux2to1455_and1;
  assign f_arrdiv32_mux2to1456_and0 = f_arrdiv32_mux2to1424_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1456_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1456_and1 = f_arrdiv32_fs470_xor1 & f_arrdiv32_mux2to1456_not0;
  assign f_arrdiv32_mux2to1456_xor0 = f_arrdiv32_mux2to1456_and0 ^ f_arrdiv32_mux2to1456_and1;
  assign f_arrdiv32_mux2to1457_and0 = f_arrdiv32_mux2to1425_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1457_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1457_and1 = f_arrdiv32_fs471_xor1 & f_arrdiv32_mux2to1457_not0;
  assign f_arrdiv32_mux2to1457_xor0 = f_arrdiv32_mux2to1457_and0 ^ f_arrdiv32_mux2to1457_and1;
  assign f_arrdiv32_mux2to1458_and0 = f_arrdiv32_mux2to1426_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1458_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1458_and1 = f_arrdiv32_fs472_xor1 & f_arrdiv32_mux2to1458_not0;
  assign f_arrdiv32_mux2to1458_xor0 = f_arrdiv32_mux2to1458_and0 ^ f_arrdiv32_mux2to1458_and1;
  assign f_arrdiv32_mux2to1459_and0 = f_arrdiv32_mux2to1427_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1459_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1459_and1 = f_arrdiv32_fs473_xor1 & f_arrdiv32_mux2to1459_not0;
  assign f_arrdiv32_mux2to1459_xor0 = f_arrdiv32_mux2to1459_and0 ^ f_arrdiv32_mux2to1459_and1;
  assign f_arrdiv32_mux2to1460_and0 = f_arrdiv32_mux2to1428_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1460_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1460_and1 = f_arrdiv32_fs474_xor1 & f_arrdiv32_mux2to1460_not0;
  assign f_arrdiv32_mux2to1460_xor0 = f_arrdiv32_mux2to1460_and0 ^ f_arrdiv32_mux2to1460_and1;
  assign f_arrdiv32_mux2to1461_and0 = f_arrdiv32_mux2to1429_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1461_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1461_and1 = f_arrdiv32_fs475_xor1 & f_arrdiv32_mux2to1461_not0;
  assign f_arrdiv32_mux2to1461_xor0 = f_arrdiv32_mux2to1461_and0 ^ f_arrdiv32_mux2to1461_and1;
  assign f_arrdiv32_mux2to1462_and0 = f_arrdiv32_mux2to1430_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1462_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1462_and1 = f_arrdiv32_fs476_xor1 & f_arrdiv32_mux2to1462_not0;
  assign f_arrdiv32_mux2to1462_xor0 = f_arrdiv32_mux2to1462_and0 ^ f_arrdiv32_mux2to1462_and1;
  assign f_arrdiv32_mux2to1463_and0 = f_arrdiv32_mux2to1431_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1463_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1463_and1 = f_arrdiv32_fs477_xor1 & f_arrdiv32_mux2to1463_not0;
  assign f_arrdiv32_mux2to1463_xor0 = f_arrdiv32_mux2to1463_and0 ^ f_arrdiv32_mux2to1463_and1;
  assign f_arrdiv32_mux2to1464_and0 = f_arrdiv32_mux2to1432_xor0 & f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1464_not0 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_mux2to1464_and1 = f_arrdiv32_fs478_xor1 & f_arrdiv32_mux2to1464_not0;
  assign f_arrdiv32_mux2to1464_xor0 = f_arrdiv32_mux2to1464_and0 ^ f_arrdiv32_mux2to1464_and1;
  assign f_arrdiv32_not14 = ~f_arrdiv32_fs479_or0;
  assign f_arrdiv32_fs480_xor0 = a[16] ^ b[0];
  assign f_arrdiv32_fs480_not0 = ~a[16];
  assign f_arrdiv32_fs480_and0 = f_arrdiv32_fs480_not0 & b[0];
  assign f_arrdiv32_fs480_not1 = ~f_arrdiv32_fs480_xor0;
  assign f_arrdiv32_fs481_xor0 = f_arrdiv32_mux2to1434_xor0 ^ b[1];
  assign f_arrdiv32_fs481_not0 = ~f_arrdiv32_mux2to1434_xor0;
  assign f_arrdiv32_fs481_and0 = f_arrdiv32_fs481_not0 & b[1];
  assign f_arrdiv32_fs481_xor1 = f_arrdiv32_fs480_and0 ^ f_arrdiv32_fs481_xor0;
  assign f_arrdiv32_fs481_not1 = ~f_arrdiv32_fs481_xor0;
  assign f_arrdiv32_fs481_and1 = f_arrdiv32_fs481_not1 & f_arrdiv32_fs480_and0;
  assign f_arrdiv32_fs481_or0 = f_arrdiv32_fs481_and1 | f_arrdiv32_fs481_and0;
  assign f_arrdiv32_fs482_xor0 = f_arrdiv32_mux2to1435_xor0 ^ b[2];
  assign f_arrdiv32_fs482_not0 = ~f_arrdiv32_mux2to1435_xor0;
  assign f_arrdiv32_fs482_and0 = f_arrdiv32_fs482_not0 & b[2];
  assign f_arrdiv32_fs482_xor1 = f_arrdiv32_fs481_or0 ^ f_arrdiv32_fs482_xor0;
  assign f_arrdiv32_fs482_not1 = ~f_arrdiv32_fs482_xor0;
  assign f_arrdiv32_fs482_and1 = f_arrdiv32_fs482_not1 & f_arrdiv32_fs481_or0;
  assign f_arrdiv32_fs482_or0 = f_arrdiv32_fs482_and1 | f_arrdiv32_fs482_and0;
  assign f_arrdiv32_fs483_xor0 = f_arrdiv32_mux2to1436_xor0 ^ b[3];
  assign f_arrdiv32_fs483_not0 = ~f_arrdiv32_mux2to1436_xor0;
  assign f_arrdiv32_fs483_and0 = f_arrdiv32_fs483_not0 & b[3];
  assign f_arrdiv32_fs483_xor1 = f_arrdiv32_fs482_or0 ^ f_arrdiv32_fs483_xor0;
  assign f_arrdiv32_fs483_not1 = ~f_arrdiv32_fs483_xor0;
  assign f_arrdiv32_fs483_and1 = f_arrdiv32_fs483_not1 & f_arrdiv32_fs482_or0;
  assign f_arrdiv32_fs483_or0 = f_arrdiv32_fs483_and1 | f_arrdiv32_fs483_and0;
  assign f_arrdiv32_fs484_xor0 = f_arrdiv32_mux2to1437_xor0 ^ b[4];
  assign f_arrdiv32_fs484_not0 = ~f_arrdiv32_mux2to1437_xor0;
  assign f_arrdiv32_fs484_and0 = f_arrdiv32_fs484_not0 & b[4];
  assign f_arrdiv32_fs484_xor1 = f_arrdiv32_fs483_or0 ^ f_arrdiv32_fs484_xor0;
  assign f_arrdiv32_fs484_not1 = ~f_arrdiv32_fs484_xor0;
  assign f_arrdiv32_fs484_and1 = f_arrdiv32_fs484_not1 & f_arrdiv32_fs483_or0;
  assign f_arrdiv32_fs484_or0 = f_arrdiv32_fs484_and1 | f_arrdiv32_fs484_and0;
  assign f_arrdiv32_fs485_xor0 = f_arrdiv32_mux2to1438_xor0 ^ b[5];
  assign f_arrdiv32_fs485_not0 = ~f_arrdiv32_mux2to1438_xor0;
  assign f_arrdiv32_fs485_and0 = f_arrdiv32_fs485_not0 & b[5];
  assign f_arrdiv32_fs485_xor1 = f_arrdiv32_fs484_or0 ^ f_arrdiv32_fs485_xor0;
  assign f_arrdiv32_fs485_not1 = ~f_arrdiv32_fs485_xor0;
  assign f_arrdiv32_fs485_and1 = f_arrdiv32_fs485_not1 & f_arrdiv32_fs484_or0;
  assign f_arrdiv32_fs485_or0 = f_arrdiv32_fs485_and1 | f_arrdiv32_fs485_and0;
  assign f_arrdiv32_fs486_xor0 = f_arrdiv32_mux2to1439_xor0 ^ b[6];
  assign f_arrdiv32_fs486_not0 = ~f_arrdiv32_mux2to1439_xor0;
  assign f_arrdiv32_fs486_and0 = f_arrdiv32_fs486_not0 & b[6];
  assign f_arrdiv32_fs486_xor1 = f_arrdiv32_fs485_or0 ^ f_arrdiv32_fs486_xor0;
  assign f_arrdiv32_fs486_not1 = ~f_arrdiv32_fs486_xor0;
  assign f_arrdiv32_fs486_and1 = f_arrdiv32_fs486_not1 & f_arrdiv32_fs485_or0;
  assign f_arrdiv32_fs486_or0 = f_arrdiv32_fs486_and1 | f_arrdiv32_fs486_and0;
  assign f_arrdiv32_fs487_xor0 = f_arrdiv32_mux2to1440_xor0 ^ b[7];
  assign f_arrdiv32_fs487_not0 = ~f_arrdiv32_mux2to1440_xor0;
  assign f_arrdiv32_fs487_and0 = f_arrdiv32_fs487_not0 & b[7];
  assign f_arrdiv32_fs487_xor1 = f_arrdiv32_fs486_or0 ^ f_arrdiv32_fs487_xor0;
  assign f_arrdiv32_fs487_not1 = ~f_arrdiv32_fs487_xor0;
  assign f_arrdiv32_fs487_and1 = f_arrdiv32_fs487_not1 & f_arrdiv32_fs486_or0;
  assign f_arrdiv32_fs487_or0 = f_arrdiv32_fs487_and1 | f_arrdiv32_fs487_and0;
  assign f_arrdiv32_fs488_xor0 = f_arrdiv32_mux2to1441_xor0 ^ b[8];
  assign f_arrdiv32_fs488_not0 = ~f_arrdiv32_mux2to1441_xor0;
  assign f_arrdiv32_fs488_and0 = f_arrdiv32_fs488_not0 & b[8];
  assign f_arrdiv32_fs488_xor1 = f_arrdiv32_fs487_or0 ^ f_arrdiv32_fs488_xor0;
  assign f_arrdiv32_fs488_not1 = ~f_arrdiv32_fs488_xor0;
  assign f_arrdiv32_fs488_and1 = f_arrdiv32_fs488_not1 & f_arrdiv32_fs487_or0;
  assign f_arrdiv32_fs488_or0 = f_arrdiv32_fs488_and1 | f_arrdiv32_fs488_and0;
  assign f_arrdiv32_fs489_xor0 = f_arrdiv32_mux2to1442_xor0 ^ b[9];
  assign f_arrdiv32_fs489_not0 = ~f_arrdiv32_mux2to1442_xor0;
  assign f_arrdiv32_fs489_and0 = f_arrdiv32_fs489_not0 & b[9];
  assign f_arrdiv32_fs489_xor1 = f_arrdiv32_fs488_or0 ^ f_arrdiv32_fs489_xor0;
  assign f_arrdiv32_fs489_not1 = ~f_arrdiv32_fs489_xor0;
  assign f_arrdiv32_fs489_and1 = f_arrdiv32_fs489_not1 & f_arrdiv32_fs488_or0;
  assign f_arrdiv32_fs489_or0 = f_arrdiv32_fs489_and1 | f_arrdiv32_fs489_and0;
  assign f_arrdiv32_fs490_xor0 = f_arrdiv32_mux2to1443_xor0 ^ b[10];
  assign f_arrdiv32_fs490_not0 = ~f_arrdiv32_mux2to1443_xor0;
  assign f_arrdiv32_fs490_and0 = f_arrdiv32_fs490_not0 & b[10];
  assign f_arrdiv32_fs490_xor1 = f_arrdiv32_fs489_or0 ^ f_arrdiv32_fs490_xor0;
  assign f_arrdiv32_fs490_not1 = ~f_arrdiv32_fs490_xor0;
  assign f_arrdiv32_fs490_and1 = f_arrdiv32_fs490_not1 & f_arrdiv32_fs489_or0;
  assign f_arrdiv32_fs490_or0 = f_arrdiv32_fs490_and1 | f_arrdiv32_fs490_and0;
  assign f_arrdiv32_fs491_xor0 = f_arrdiv32_mux2to1444_xor0 ^ b[11];
  assign f_arrdiv32_fs491_not0 = ~f_arrdiv32_mux2to1444_xor0;
  assign f_arrdiv32_fs491_and0 = f_arrdiv32_fs491_not0 & b[11];
  assign f_arrdiv32_fs491_xor1 = f_arrdiv32_fs490_or0 ^ f_arrdiv32_fs491_xor0;
  assign f_arrdiv32_fs491_not1 = ~f_arrdiv32_fs491_xor0;
  assign f_arrdiv32_fs491_and1 = f_arrdiv32_fs491_not1 & f_arrdiv32_fs490_or0;
  assign f_arrdiv32_fs491_or0 = f_arrdiv32_fs491_and1 | f_arrdiv32_fs491_and0;
  assign f_arrdiv32_fs492_xor0 = f_arrdiv32_mux2to1445_xor0 ^ b[12];
  assign f_arrdiv32_fs492_not0 = ~f_arrdiv32_mux2to1445_xor0;
  assign f_arrdiv32_fs492_and0 = f_arrdiv32_fs492_not0 & b[12];
  assign f_arrdiv32_fs492_xor1 = f_arrdiv32_fs491_or0 ^ f_arrdiv32_fs492_xor0;
  assign f_arrdiv32_fs492_not1 = ~f_arrdiv32_fs492_xor0;
  assign f_arrdiv32_fs492_and1 = f_arrdiv32_fs492_not1 & f_arrdiv32_fs491_or0;
  assign f_arrdiv32_fs492_or0 = f_arrdiv32_fs492_and1 | f_arrdiv32_fs492_and0;
  assign f_arrdiv32_fs493_xor0 = f_arrdiv32_mux2to1446_xor0 ^ b[13];
  assign f_arrdiv32_fs493_not0 = ~f_arrdiv32_mux2to1446_xor0;
  assign f_arrdiv32_fs493_and0 = f_arrdiv32_fs493_not0 & b[13];
  assign f_arrdiv32_fs493_xor1 = f_arrdiv32_fs492_or0 ^ f_arrdiv32_fs493_xor0;
  assign f_arrdiv32_fs493_not1 = ~f_arrdiv32_fs493_xor0;
  assign f_arrdiv32_fs493_and1 = f_arrdiv32_fs493_not1 & f_arrdiv32_fs492_or0;
  assign f_arrdiv32_fs493_or0 = f_arrdiv32_fs493_and1 | f_arrdiv32_fs493_and0;
  assign f_arrdiv32_fs494_xor0 = f_arrdiv32_mux2to1447_xor0 ^ b[14];
  assign f_arrdiv32_fs494_not0 = ~f_arrdiv32_mux2to1447_xor0;
  assign f_arrdiv32_fs494_and0 = f_arrdiv32_fs494_not0 & b[14];
  assign f_arrdiv32_fs494_xor1 = f_arrdiv32_fs493_or0 ^ f_arrdiv32_fs494_xor0;
  assign f_arrdiv32_fs494_not1 = ~f_arrdiv32_fs494_xor0;
  assign f_arrdiv32_fs494_and1 = f_arrdiv32_fs494_not1 & f_arrdiv32_fs493_or0;
  assign f_arrdiv32_fs494_or0 = f_arrdiv32_fs494_and1 | f_arrdiv32_fs494_and0;
  assign f_arrdiv32_fs495_xor0 = f_arrdiv32_mux2to1448_xor0 ^ b[15];
  assign f_arrdiv32_fs495_not0 = ~f_arrdiv32_mux2to1448_xor0;
  assign f_arrdiv32_fs495_and0 = f_arrdiv32_fs495_not0 & b[15];
  assign f_arrdiv32_fs495_xor1 = f_arrdiv32_fs494_or0 ^ f_arrdiv32_fs495_xor0;
  assign f_arrdiv32_fs495_not1 = ~f_arrdiv32_fs495_xor0;
  assign f_arrdiv32_fs495_and1 = f_arrdiv32_fs495_not1 & f_arrdiv32_fs494_or0;
  assign f_arrdiv32_fs495_or0 = f_arrdiv32_fs495_and1 | f_arrdiv32_fs495_and0;
  assign f_arrdiv32_fs496_xor0 = f_arrdiv32_mux2to1449_xor0 ^ b[16];
  assign f_arrdiv32_fs496_not0 = ~f_arrdiv32_mux2to1449_xor0;
  assign f_arrdiv32_fs496_and0 = f_arrdiv32_fs496_not0 & b[16];
  assign f_arrdiv32_fs496_xor1 = f_arrdiv32_fs495_or0 ^ f_arrdiv32_fs496_xor0;
  assign f_arrdiv32_fs496_not1 = ~f_arrdiv32_fs496_xor0;
  assign f_arrdiv32_fs496_and1 = f_arrdiv32_fs496_not1 & f_arrdiv32_fs495_or0;
  assign f_arrdiv32_fs496_or0 = f_arrdiv32_fs496_and1 | f_arrdiv32_fs496_and0;
  assign f_arrdiv32_fs497_xor0 = f_arrdiv32_mux2to1450_xor0 ^ b[17];
  assign f_arrdiv32_fs497_not0 = ~f_arrdiv32_mux2to1450_xor0;
  assign f_arrdiv32_fs497_and0 = f_arrdiv32_fs497_not0 & b[17];
  assign f_arrdiv32_fs497_xor1 = f_arrdiv32_fs496_or0 ^ f_arrdiv32_fs497_xor0;
  assign f_arrdiv32_fs497_not1 = ~f_arrdiv32_fs497_xor0;
  assign f_arrdiv32_fs497_and1 = f_arrdiv32_fs497_not1 & f_arrdiv32_fs496_or0;
  assign f_arrdiv32_fs497_or0 = f_arrdiv32_fs497_and1 | f_arrdiv32_fs497_and0;
  assign f_arrdiv32_fs498_xor0 = f_arrdiv32_mux2to1451_xor0 ^ b[18];
  assign f_arrdiv32_fs498_not0 = ~f_arrdiv32_mux2to1451_xor0;
  assign f_arrdiv32_fs498_and0 = f_arrdiv32_fs498_not0 & b[18];
  assign f_arrdiv32_fs498_xor1 = f_arrdiv32_fs497_or0 ^ f_arrdiv32_fs498_xor0;
  assign f_arrdiv32_fs498_not1 = ~f_arrdiv32_fs498_xor0;
  assign f_arrdiv32_fs498_and1 = f_arrdiv32_fs498_not1 & f_arrdiv32_fs497_or0;
  assign f_arrdiv32_fs498_or0 = f_arrdiv32_fs498_and1 | f_arrdiv32_fs498_and0;
  assign f_arrdiv32_fs499_xor0 = f_arrdiv32_mux2to1452_xor0 ^ b[19];
  assign f_arrdiv32_fs499_not0 = ~f_arrdiv32_mux2to1452_xor0;
  assign f_arrdiv32_fs499_and0 = f_arrdiv32_fs499_not0 & b[19];
  assign f_arrdiv32_fs499_xor1 = f_arrdiv32_fs498_or0 ^ f_arrdiv32_fs499_xor0;
  assign f_arrdiv32_fs499_not1 = ~f_arrdiv32_fs499_xor0;
  assign f_arrdiv32_fs499_and1 = f_arrdiv32_fs499_not1 & f_arrdiv32_fs498_or0;
  assign f_arrdiv32_fs499_or0 = f_arrdiv32_fs499_and1 | f_arrdiv32_fs499_and0;
  assign f_arrdiv32_fs500_xor0 = f_arrdiv32_mux2to1453_xor0 ^ b[20];
  assign f_arrdiv32_fs500_not0 = ~f_arrdiv32_mux2to1453_xor0;
  assign f_arrdiv32_fs500_and0 = f_arrdiv32_fs500_not0 & b[20];
  assign f_arrdiv32_fs500_xor1 = f_arrdiv32_fs499_or0 ^ f_arrdiv32_fs500_xor0;
  assign f_arrdiv32_fs500_not1 = ~f_arrdiv32_fs500_xor0;
  assign f_arrdiv32_fs500_and1 = f_arrdiv32_fs500_not1 & f_arrdiv32_fs499_or0;
  assign f_arrdiv32_fs500_or0 = f_arrdiv32_fs500_and1 | f_arrdiv32_fs500_and0;
  assign f_arrdiv32_fs501_xor0 = f_arrdiv32_mux2to1454_xor0 ^ b[21];
  assign f_arrdiv32_fs501_not0 = ~f_arrdiv32_mux2to1454_xor0;
  assign f_arrdiv32_fs501_and0 = f_arrdiv32_fs501_not0 & b[21];
  assign f_arrdiv32_fs501_xor1 = f_arrdiv32_fs500_or0 ^ f_arrdiv32_fs501_xor0;
  assign f_arrdiv32_fs501_not1 = ~f_arrdiv32_fs501_xor0;
  assign f_arrdiv32_fs501_and1 = f_arrdiv32_fs501_not1 & f_arrdiv32_fs500_or0;
  assign f_arrdiv32_fs501_or0 = f_arrdiv32_fs501_and1 | f_arrdiv32_fs501_and0;
  assign f_arrdiv32_fs502_xor0 = f_arrdiv32_mux2to1455_xor0 ^ b[22];
  assign f_arrdiv32_fs502_not0 = ~f_arrdiv32_mux2to1455_xor0;
  assign f_arrdiv32_fs502_and0 = f_arrdiv32_fs502_not0 & b[22];
  assign f_arrdiv32_fs502_xor1 = f_arrdiv32_fs501_or0 ^ f_arrdiv32_fs502_xor0;
  assign f_arrdiv32_fs502_not1 = ~f_arrdiv32_fs502_xor0;
  assign f_arrdiv32_fs502_and1 = f_arrdiv32_fs502_not1 & f_arrdiv32_fs501_or0;
  assign f_arrdiv32_fs502_or0 = f_arrdiv32_fs502_and1 | f_arrdiv32_fs502_and0;
  assign f_arrdiv32_fs503_xor0 = f_arrdiv32_mux2to1456_xor0 ^ b[23];
  assign f_arrdiv32_fs503_not0 = ~f_arrdiv32_mux2to1456_xor0;
  assign f_arrdiv32_fs503_and0 = f_arrdiv32_fs503_not0 & b[23];
  assign f_arrdiv32_fs503_xor1 = f_arrdiv32_fs502_or0 ^ f_arrdiv32_fs503_xor0;
  assign f_arrdiv32_fs503_not1 = ~f_arrdiv32_fs503_xor0;
  assign f_arrdiv32_fs503_and1 = f_arrdiv32_fs503_not1 & f_arrdiv32_fs502_or0;
  assign f_arrdiv32_fs503_or0 = f_arrdiv32_fs503_and1 | f_arrdiv32_fs503_and0;
  assign f_arrdiv32_fs504_xor0 = f_arrdiv32_mux2to1457_xor0 ^ b[24];
  assign f_arrdiv32_fs504_not0 = ~f_arrdiv32_mux2to1457_xor0;
  assign f_arrdiv32_fs504_and0 = f_arrdiv32_fs504_not0 & b[24];
  assign f_arrdiv32_fs504_xor1 = f_arrdiv32_fs503_or0 ^ f_arrdiv32_fs504_xor0;
  assign f_arrdiv32_fs504_not1 = ~f_arrdiv32_fs504_xor0;
  assign f_arrdiv32_fs504_and1 = f_arrdiv32_fs504_not1 & f_arrdiv32_fs503_or0;
  assign f_arrdiv32_fs504_or0 = f_arrdiv32_fs504_and1 | f_arrdiv32_fs504_and0;
  assign f_arrdiv32_fs505_xor0 = f_arrdiv32_mux2to1458_xor0 ^ b[25];
  assign f_arrdiv32_fs505_not0 = ~f_arrdiv32_mux2to1458_xor0;
  assign f_arrdiv32_fs505_and0 = f_arrdiv32_fs505_not0 & b[25];
  assign f_arrdiv32_fs505_xor1 = f_arrdiv32_fs504_or0 ^ f_arrdiv32_fs505_xor0;
  assign f_arrdiv32_fs505_not1 = ~f_arrdiv32_fs505_xor0;
  assign f_arrdiv32_fs505_and1 = f_arrdiv32_fs505_not1 & f_arrdiv32_fs504_or0;
  assign f_arrdiv32_fs505_or0 = f_arrdiv32_fs505_and1 | f_arrdiv32_fs505_and0;
  assign f_arrdiv32_fs506_xor0 = f_arrdiv32_mux2to1459_xor0 ^ b[26];
  assign f_arrdiv32_fs506_not0 = ~f_arrdiv32_mux2to1459_xor0;
  assign f_arrdiv32_fs506_and0 = f_arrdiv32_fs506_not0 & b[26];
  assign f_arrdiv32_fs506_xor1 = f_arrdiv32_fs505_or0 ^ f_arrdiv32_fs506_xor0;
  assign f_arrdiv32_fs506_not1 = ~f_arrdiv32_fs506_xor0;
  assign f_arrdiv32_fs506_and1 = f_arrdiv32_fs506_not1 & f_arrdiv32_fs505_or0;
  assign f_arrdiv32_fs506_or0 = f_arrdiv32_fs506_and1 | f_arrdiv32_fs506_and0;
  assign f_arrdiv32_fs507_xor0 = f_arrdiv32_mux2to1460_xor0 ^ b[27];
  assign f_arrdiv32_fs507_not0 = ~f_arrdiv32_mux2to1460_xor0;
  assign f_arrdiv32_fs507_and0 = f_arrdiv32_fs507_not0 & b[27];
  assign f_arrdiv32_fs507_xor1 = f_arrdiv32_fs506_or0 ^ f_arrdiv32_fs507_xor0;
  assign f_arrdiv32_fs507_not1 = ~f_arrdiv32_fs507_xor0;
  assign f_arrdiv32_fs507_and1 = f_arrdiv32_fs507_not1 & f_arrdiv32_fs506_or0;
  assign f_arrdiv32_fs507_or0 = f_arrdiv32_fs507_and1 | f_arrdiv32_fs507_and0;
  assign f_arrdiv32_fs508_xor0 = f_arrdiv32_mux2to1461_xor0 ^ b[28];
  assign f_arrdiv32_fs508_not0 = ~f_arrdiv32_mux2to1461_xor0;
  assign f_arrdiv32_fs508_and0 = f_arrdiv32_fs508_not0 & b[28];
  assign f_arrdiv32_fs508_xor1 = f_arrdiv32_fs507_or0 ^ f_arrdiv32_fs508_xor0;
  assign f_arrdiv32_fs508_not1 = ~f_arrdiv32_fs508_xor0;
  assign f_arrdiv32_fs508_and1 = f_arrdiv32_fs508_not1 & f_arrdiv32_fs507_or0;
  assign f_arrdiv32_fs508_or0 = f_arrdiv32_fs508_and1 | f_arrdiv32_fs508_and0;
  assign f_arrdiv32_fs509_xor0 = f_arrdiv32_mux2to1462_xor0 ^ b[29];
  assign f_arrdiv32_fs509_not0 = ~f_arrdiv32_mux2to1462_xor0;
  assign f_arrdiv32_fs509_and0 = f_arrdiv32_fs509_not0 & b[29];
  assign f_arrdiv32_fs509_xor1 = f_arrdiv32_fs508_or0 ^ f_arrdiv32_fs509_xor0;
  assign f_arrdiv32_fs509_not1 = ~f_arrdiv32_fs509_xor0;
  assign f_arrdiv32_fs509_and1 = f_arrdiv32_fs509_not1 & f_arrdiv32_fs508_or0;
  assign f_arrdiv32_fs509_or0 = f_arrdiv32_fs509_and1 | f_arrdiv32_fs509_and0;
  assign f_arrdiv32_fs510_xor0 = f_arrdiv32_mux2to1463_xor0 ^ b[30];
  assign f_arrdiv32_fs510_not0 = ~f_arrdiv32_mux2to1463_xor0;
  assign f_arrdiv32_fs510_and0 = f_arrdiv32_fs510_not0 & b[30];
  assign f_arrdiv32_fs510_xor1 = f_arrdiv32_fs509_or0 ^ f_arrdiv32_fs510_xor0;
  assign f_arrdiv32_fs510_not1 = ~f_arrdiv32_fs510_xor0;
  assign f_arrdiv32_fs510_and1 = f_arrdiv32_fs510_not1 & f_arrdiv32_fs509_or0;
  assign f_arrdiv32_fs510_or0 = f_arrdiv32_fs510_and1 | f_arrdiv32_fs510_and0;
  assign f_arrdiv32_fs511_xor0 = f_arrdiv32_mux2to1464_xor0 ^ b[31];
  assign f_arrdiv32_fs511_not0 = ~f_arrdiv32_mux2to1464_xor0;
  assign f_arrdiv32_fs511_and0 = f_arrdiv32_fs511_not0 & b[31];
  assign f_arrdiv32_fs511_xor1 = f_arrdiv32_fs510_or0 ^ f_arrdiv32_fs511_xor0;
  assign f_arrdiv32_fs511_not1 = ~f_arrdiv32_fs511_xor0;
  assign f_arrdiv32_fs511_and1 = f_arrdiv32_fs511_not1 & f_arrdiv32_fs510_or0;
  assign f_arrdiv32_fs511_or0 = f_arrdiv32_fs511_and1 | f_arrdiv32_fs511_and0;
  assign f_arrdiv32_mux2to1465_and0 = a[16] & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1465_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1465_and1 = f_arrdiv32_fs480_xor0 & f_arrdiv32_mux2to1465_not0;
  assign f_arrdiv32_mux2to1465_xor0 = f_arrdiv32_mux2to1465_and0 ^ f_arrdiv32_mux2to1465_and1;
  assign f_arrdiv32_mux2to1466_and0 = f_arrdiv32_mux2to1434_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1466_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1466_and1 = f_arrdiv32_fs481_xor1 & f_arrdiv32_mux2to1466_not0;
  assign f_arrdiv32_mux2to1466_xor0 = f_arrdiv32_mux2to1466_and0 ^ f_arrdiv32_mux2to1466_and1;
  assign f_arrdiv32_mux2to1467_and0 = f_arrdiv32_mux2to1435_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1467_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1467_and1 = f_arrdiv32_fs482_xor1 & f_arrdiv32_mux2to1467_not0;
  assign f_arrdiv32_mux2to1467_xor0 = f_arrdiv32_mux2to1467_and0 ^ f_arrdiv32_mux2to1467_and1;
  assign f_arrdiv32_mux2to1468_and0 = f_arrdiv32_mux2to1436_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1468_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1468_and1 = f_arrdiv32_fs483_xor1 & f_arrdiv32_mux2to1468_not0;
  assign f_arrdiv32_mux2to1468_xor0 = f_arrdiv32_mux2to1468_and0 ^ f_arrdiv32_mux2to1468_and1;
  assign f_arrdiv32_mux2to1469_and0 = f_arrdiv32_mux2to1437_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1469_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1469_and1 = f_arrdiv32_fs484_xor1 & f_arrdiv32_mux2to1469_not0;
  assign f_arrdiv32_mux2to1469_xor0 = f_arrdiv32_mux2to1469_and0 ^ f_arrdiv32_mux2to1469_and1;
  assign f_arrdiv32_mux2to1470_and0 = f_arrdiv32_mux2to1438_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1470_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1470_and1 = f_arrdiv32_fs485_xor1 & f_arrdiv32_mux2to1470_not0;
  assign f_arrdiv32_mux2to1470_xor0 = f_arrdiv32_mux2to1470_and0 ^ f_arrdiv32_mux2to1470_and1;
  assign f_arrdiv32_mux2to1471_and0 = f_arrdiv32_mux2to1439_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1471_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1471_and1 = f_arrdiv32_fs486_xor1 & f_arrdiv32_mux2to1471_not0;
  assign f_arrdiv32_mux2to1471_xor0 = f_arrdiv32_mux2to1471_and0 ^ f_arrdiv32_mux2to1471_and1;
  assign f_arrdiv32_mux2to1472_and0 = f_arrdiv32_mux2to1440_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1472_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1472_and1 = f_arrdiv32_fs487_xor1 & f_arrdiv32_mux2to1472_not0;
  assign f_arrdiv32_mux2to1472_xor0 = f_arrdiv32_mux2to1472_and0 ^ f_arrdiv32_mux2to1472_and1;
  assign f_arrdiv32_mux2to1473_and0 = f_arrdiv32_mux2to1441_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1473_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1473_and1 = f_arrdiv32_fs488_xor1 & f_arrdiv32_mux2to1473_not0;
  assign f_arrdiv32_mux2to1473_xor0 = f_arrdiv32_mux2to1473_and0 ^ f_arrdiv32_mux2to1473_and1;
  assign f_arrdiv32_mux2to1474_and0 = f_arrdiv32_mux2to1442_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1474_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1474_and1 = f_arrdiv32_fs489_xor1 & f_arrdiv32_mux2to1474_not0;
  assign f_arrdiv32_mux2to1474_xor0 = f_arrdiv32_mux2to1474_and0 ^ f_arrdiv32_mux2to1474_and1;
  assign f_arrdiv32_mux2to1475_and0 = f_arrdiv32_mux2to1443_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1475_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1475_and1 = f_arrdiv32_fs490_xor1 & f_arrdiv32_mux2to1475_not0;
  assign f_arrdiv32_mux2to1475_xor0 = f_arrdiv32_mux2to1475_and0 ^ f_arrdiv32_mux2to1475_and1;
  assign f_arrdiv32_mux2to1476_and0 = f_arrdiv32_mux2to1444_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1476_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1476_and1 = f_arrdiv32_fs491_xor1 & f_arrdiv32_mux2to1476_not0;
  assign f_arrdiv32_mux2to1476_xor0 = f_arrdiv32_mux2to1476_and0 ^ f_arrdiv32_mux2to1476_and1;
  assign f_arrdiv32_mux2to1477_and0 = f_arrdiv32_mux2to1445_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1477_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1477_and1 = f_arrdiv32_fs492_xor1 & f_arrdiv32_mux2to1477_not0;
  assign f_arrdiv32_mux2to1477_xor0 = f_arrdiv32_mux2to1477_and0 ^ f_arrdiv32_mux2to1477_and1;
  assign f_arrdiv32_mux2to1478_and0 = f_arrdiv32_mux2to1446_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1478_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1478_and1 = f_arrdiv32_fs493_xor1 & f_arrdiv32_mux2to1478_not0;
  assign f_arrdiv32_mux2to1478_xor0 = f_arrdiv32_mux2to1478_and0 ^ f_arrdiv32_mux2to1478_and1;
  assign f_arrdiv32_mux2to1479_and0 = f_arrdiv32_mux2to1447_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1479_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1479_and1 = f_arrdiv32_fs494_xor1 & f_arrdiv32_mux2to1479_not0;
  assign f_arrdiv32_mux2to1479_xor0 = f_arrdiv32_mux2to1479_and0 ^ f_arrdiv32_mux2to1479_and1;
  assign f_arrdiv32_mux2to1480_and0 = f_arrdiv32_mux2to1448_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1480_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1480_and1 = f_arrdiv32_fs495_xor1 & f_arrdiv32_mux2to1480_not0;
  assign f_arrdiv32_mux2to1480_xor0 = f_arrdiv32_mux2to1480_and0 ^ f_arrdiv32_mux2to1480_and1;
  assign f_arrdiv32_mux2to1481_and0 = f_arrdiv32_mux2to1449_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1481_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1481_and1 = f_arrdiv32_fs496_xor1 & f_arrdiv32_mux2to1481_not0;
  assign f_arrdiv32_mux2to1481_xor0 = f_arrdiv32_mux2to1481_and0 ^ f_arrdiv32_mux2to1481_and1;
  assign f_arrdiv32_mux2to1482_and0 = f_arrdiv32_mux2to1450_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1482_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1482_and1 = f_arrdiv32_fs497_xor1 & f_arrdiv32_mux2to1482_not0;
  assign f_arrdiv32_mux2to1482_xor0 = f_arrdiv32_mux2to1482_and0 ^ f_arrdiv32_mux2to1482_and1;
  assign f_arrdiv32_mux2to1483_and0 = f_arrdiv32_mux2to1451_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1483_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1483_and1 = f_arrdiv32_fs498_xor1 & f_arrdiv32_mux2to1483_not0;
  assign f_arrdiv32_mux2to1483_xor0 = f_arrdiv32_mux2to1483_and0 ^ f_arrdiv32_mux2to1483_and1;
  assign f_arrdiv32_mux2to1484_and0 = f_arrdiv32_mux2to1452_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1484_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1484_and1 = f_arrdiv32_fs499_xor1 & f_arrdiv32_mux2to1484_not0;
  assign f_arrdiv32_mux2to1484_xor0 = f_arrdiv32_mux2to1484_and0 ^ f_arrdiv32_mux2to1484_and1;
  assign f_arrdiv32_mux2to1485_and0 = f_arrdiv32_mux2to1453_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1485_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1485_and1 = f_arrdiv32_fs500_xor1 & f_arrdiv32_mux2to1485_not0;
  assign f_arrdiv32_mux2to1485_xor0 = f_arrdiv32_mux2to1485_and0 ^ f_arrdiv32_mux2to1485_and1;
  assign f_arrdiv32_mux2to1486_and0 = f_arrdiv32_mux2to1454_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1486_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1486_and1 = f_arrdiv32_fs501_xor1 & f_arrdiv32_mux2to1486_not0;
  assign f_arrdiv32_mux2to1486_xor0 = f_arrdiv32_mux2to1486_and0 ^ f_arrdiv32_mux2to1486_and1;
  assign f_arrdiv32_mux2to1487_and0 = f_arrdiv32_mux2to1455_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1487_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1487_and1 = f_arrdiv32_fs502_xor1 & f_arrdiv32_mux2to1487_not0;
  assign f_arrdiv32_mux2to1487_xor0 = f_arrdiv32_mux2to1487_and0 ^ f_arrdiv32_mux2to1487_and1;
  assign f_arrdiv32_mux2to1488_and0 = f_arrdiv32_mux2to1456_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1488_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1488_and1 = f_arrdiv32_fs503_xor1 & f_arrdiv32_mux2to1488_not0;
  assign f_arrdiv32_mux2to1488_xor0 = f_arrdiv32_mux2to1488_and0 ^ f_arrdiv32_mux2to1488_and1;
  assign f_arrdiv32_mux2to1489_and0 = f_arrdiv32_mux2to1457_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1489_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1489_and1 = f_arrdiv32_fs504_xor1 & f_arrdiv32_mux2to1489_not0;
  assign f_arrdiv32_mux2to1489_xor0 = f_arrdiv32_mux2to1489_and0 ^ f_arrdiv32_mux2to1489_and1;
  assign f_arrdiv32_mux2to1490_and0 = f_arrdiv32_mux2to1458_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1490_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1490_and1 = f_arrdiv32_fs505_xor1 & f_arrdiv32_mux2to1490_not0;
  assign f_arrdiv32_mux2to1490_xor0 = f_arrdiv32_mux2to1490_and0 ^ f_arrdiv32_mux2to1490_and1;
  assign f_arrdiv32_mux2to1491_and0 = f_arrdiv32_mux2to1459_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1491_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1491_and1 = f_arrdiv32_fs506_xor1 & f_arrdiv32_mux2to1491_not0;
  assign f_arrdiv32_mux2to1491_xor0 = f_arrdiv32_mux2to1491_and0 ^ f_arrdiv32_mux2to1491_and1;
  assign f_arrdiv32_mux2to1492_and0 = f_arrdiv32_mux2to1460_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1492_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1492_and1 = f_arrdiv32_fs507_xor1 & f_arrdiv32_mux2to1492_not0;
  assign f_arrdiv32_mux2to1492_xor0 = f_arrdiv32_mux2to1492_and0 ^ f_arrdiv32_mux2to1492_and1;
  assign f_arrdiv32_mux2to1493_and0 = f_arrdiv32_mux2to1461_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1493_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1493_and1 = f_arrdiv32_fs508_xor1 & f_arrdiv32_mux2to1493_not0;
  assign f_arrdiv32_mux2to1493_xor0 = f_arrdiv32_mux2to1493_and0 ^ f_arrdiv32_mux2to1493_and1;
  assign f_arrdiv32_mux2to1494_and0 = f_arrdiv32_mux2to1462_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1494_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1494_and1 = f_arrdiv32_fs509_xor1 & f_arrdiv32_mux2to1494_not0;
  assign f_arrdiv32_mux2to1494_xor0 = f_arrdiv32_mux2to1494_and0 ^ f_arrdiv32_mux2to1494_and1;
  assign f_arrdiv32_mux2to1495_and0 = f_arrdiv32_mux2to1463_xor0 & f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1495_not0 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_mux2to1495_and1 = f_arrdiv32_fs510_xor1 & f_arrdiv32_mux2to1495_not0;
  assign f_arrdiv32_mux2to1495_xor0 = f_arrdiv32_mux2to1495_and0 ^ f_arrdiv32_mux2to1495_and1;
  assign f_arrdiv32_not15 = ~f_arrdiv32_fs511_or0;
  assign f_arrdiv32_fs512_xor0 = a[15] ^ b[0];
  assign f_arrdiv32_fs512_not0 = ~a[15];
  assign f_arrdiv32_fs512_and0 = f_arrdiv32_fs512_not0 & b[0];
  assign f_arrdiv32_fs512_not1 = ~f_arrdiv32_fs512_xor0;
  assign f_arrdiv32_fs513_xor0 = f_arrdiv32_mux2to1465_xor0 ^ b[1];
  assign f_arrdiv32_fs513_not0 = ~f_arrdiv32_mux2to1465_xor0;
  assign f_arrdiv32_fs513_and0 = f_arrdiv32_fs513_not0 & b[1];
  assign f_arrdiv32_fs513_xor1 = f_arrdiv32_fs512_and0 ^ f_arrdiv32_fs513_xor0;
  assign f_arrdiv32_fs513_not1 = ~f_arrdiv32_fs513_xor0;
  assign f_arrdiv32_fs513_and1 = f_arrdiv32_fs513_not1 & f_arrdiv32_fs512_and0;
  assign f_arrdiv32_fs513_or0 = f_arrdiv32_fs513_and1 | f_arrdiv32_fs513_and0;
  assign f_arrdiv32_fs514_xor0 = f_arrdiv32_mux2to1466_xor0 ^ b[2];
  assign f_arrdiv32_fs514_not0 = ~f_arrdiv32_mux2to1466_xor0;
  assign f_arrdiv32_fs514_and0 = f_arrdiv32_fs514_not0 & b[2];
  assign f_arrdiv32_fs514_xor1 = f_arrdiv32_fs513_or0 ^ f_arrdiv32_fs514_xor0;
  assign f_arrdiv32_fs514_not1 = ~f_arrdiv32_fs514_xor0;
  assign f_arrdiv32_fs514_and1 = f_arrdiv32_fs514_not1 & f_arrdiv32_fs513_or0;
  assign f_arrdiv32_fs514_or0 = f_arrdiv32_fs514_and1 | f_arrdiv32_fs514_and0;
  assign f_arrdiv32_fs515_xor0 = f_arrdiv32_mux2to1467_xor0 ^ b[3];
  assign f_arrdiv32_fs515_not0 = ~f_arrdiv32_mux2to1467_xor0;
  assign f_arrdiv32_fs515_and0 = f_arrdiv32_fs515_not0 & b[3];
  assign f_arrdiv32_fs515_xor1 = f_arrdiv32_fs514_or0 ^ f_arrdiv32_fs515_xor0;
  assign f_arrdiv32_fs515_not1 = ~f_arrdiv32_fs515_xor0;
  assign f_arrdiv32_fs515_and1 = f_arrdiv32_fs515_not1 & f_arrdiv32_fs514_or0;
  assign f_arrdiv32_fs515_or0 = f_arrdiv32_fs515_and1 | f_arrdiv32_fs515_and0;
  assign f_arrdiv32_fs516_xor0 = f_arrdiv32_mux2to1468_xor0 ^ b[4];
  assign f_arrdiv32_fs516_not0 = ~f_arrdiv32_mux2to1468_xor0;
  assign f_arrdiv32_fs516_and0 = f_arrdiv32_fs516_not0 & b[4];
  assign f_arrdiv32_fs516_xor1 = f_arrdiv32_fs515_or0 ^ f_arrdiv32_fs516_xor0;
  assign f_arrdiv32_fs516_not1 = ~f_arrdiv32_fs516_xor0;
  assign f_arrdiv32_fs516_and1 = f_arrdiv32_fs516_not1 & f_arrdiv32_fs515_or0;
  assign f_arrdiv32_fs516_or0 = f_arrdiv32_fs516_and1 | f_arrdiv32_fs516_and0;
  assign f_arrdiv32_fs517_xor0 = f_arrdiv32_mux2to1469_xor0 ^ b[5];
  assign f_arrdiv32_fs517_not0 = ~f_arrdiv32_mux2to1469_xor0;
  assign f_arrdiv32_fs517_and0 = f_arrdiv32_fs517_not0 & b[5];
  assign f_arrdiv32_fs517_xor1 = f_arrdiv32_fs516_or0 ^ f_arrdiv32_fs517_xor0;
  assign f_arrdiv32_fs517_not1 = ~f_arrdiv32_fs517_xor0;
  assign f_arrdiv32_fs517_and1 = f_arrdiv32_fs517_not1 & f_arrdiv32_fs516_or0;
  assign f_arrdiv32_fs517_or0 = f_arrdiv32_fs517_and1 | f_arrdiv32_fs517_and0;
  assign f_arrdiv32_fs518_xor0 = f_arrdiv32_mux2to1470_xor0 ^ b[6];
  assign f_arrdiv32_fs518_not0 = ~f_arrdiv32_mux2to1470_xor0;
  assign f_arrdiv32_fs518_and0 = f_arrdiv32_fs518_not0 & b[6];
  assign f_arrdiv32_fs518_xor1 = f_arrdiv32_fs517_or0 ^ f_arrdiv32_fs518_xor0;
  assign f_arrdiv32_fs518_not1 = ~f_arrdiv32_fs518_xor0;
  assign f_arrdiv32_fs518_and1 = f_arrdiv32_fs518_not1 & f_arrdiv32_fs517_or0;
  assign f_arrdiv32_fs518_or0 = f_arrdiv32_fs518_and1 | f_arrdiv32_fs518_and0;
  assign f_arrdiv32_fs519_xor0 = f_arrdiv32_mux2to1471_xor0 ^ b[7];
  assign f_arrdiv32_fs519_not0 = ~f_arrdiv32_mux2to1471_xor0;
  assign f_arrdiv32_fs519_and0 = f_arrdiv32_fs519_not0 & b[7];
  assign f_arrdiv32_fs519_xor1 = f_arrdiv32_fs518_or0 ^ f_arrdiv32_fs519_xor0;
  assign f_arrdiv32_fs519_not1 = ~f_arrdiv32_fs519_xor0;
  assign f_arrdiv32_fs519_and1 = f_arrdiv32_fs519_not1 & f_arrdiv32_fs518_or0;
  assign f_arrdiv32_fs519_or0 = f_arrdiv32_fs519_and1 | f_arrdiv32_fs519_and0;
  assign f_arrdiv32_fs520_xor0 = f_arrdiv32_mux2to1472_xor0 ^ b[8];
  assign f_arrdiv32_fs520_not0 = ~f_arrdiv32_mux2to1472_xor0;
  assign f_arrdiv32_fs520_and0 = f_arrdiv32_fs520_not0 & b[8];
  assign f_arrdiv32_fs520_xor1 = f_arrdiv32_fs519_or0 ^ f_arrdiv32_fs520_xor0;
  assign f_arrdiv32_fs520_not1 = ~f_arrdiv32_fs520_xor0;
  assign f_arrdiv32_fs520_and1 = f_arrdiv32_fs520_not1 & f_arrdiv32_fs519_or0;
  assign f_arrdiv32_fs520_or0 = f_arrdiv32_fs520_and1 | f_arrdiv32_fs520_and0;
  assign f_arrdiv32_fs521_xor0 = f_arrdiv32_mux2to1473_xor0 ^ b[9];
  assign f_arrdiv32_fs521_not0 = ~f_arrdiv32_mux2to1473_xor0;
  assign f_arrdiv32_fs521_and0 = f_arrdiv32_fs521_not0 & b[9];
  assign f_arrdiv32_fs521_xor1 = f_arrdiv32_fs520_or0 ^ f_arrdiv32_fs521_xor0;
  assign f_arrdiv32_fs521_not1 = ~f_arrdiv32_fs521_xor0;
  assign f_arrdiv32_fs521_and1 = f_arrdiv32_fs521_not1 & f_arrdiv32_fs520_or0;
  assign f_arrdiv32_fs521_or0 = f_arrdiv32_fs521_and1 | f_arrdiv32_fs521_and0;
  assign f_arrdiv32_fs522_xor0 = f_arrdiv32_mux2to1474_xor0 ^ b[10];
  assign f_arrdiv32_fs522_not0 = ~f_arrdiv32_mux2to1474_xor0;
  assign f_arrdiv32_fs522_and0 = f_arrdiv32_fs522_not0 & b[10];
  assign f_arrdiv32_fs522_xor1 = f_arrdiv32_fs521_or0 ^ f_arrdiv32_fs522_xor0;
  assign f_arrdiv32_fs522_not1 = ~f_arrdiv32_fs522_xor0;
  assign f_arrdiv32_fs522_and1 = f_arrdiv32_fs522_not1 & f_arrdiv32_fs521_or0;
  assign f_arrdiv32_fs522_or0 = f_arrdiv32_fs522_and1 | f_arrdiv32_fs522_and0;
  assign f_arrdiv32_fs523_xor0 = f_arrdiv32_mux2to1475_xor0 ^ b[11];
  assign f_arrdiv32_fs523_not0 = ~f_arrdiv32_mux2to1475_xor0;
  assign f_arrdiv32_fs523_and0 = f_arrdiv32_fs523_not0 & b[11];
  assign f_arrdiv32_fs523_xor1 = f_arrdiv32_fs522_or0 ^ f_arrdiv32_fs523_xor0;
  assign f_arrdiv32_fs523_not1 = ~f_arrdiv32_fs523_xor0;
  assign f_arrdiv32_fs523_and1 = f_arrdiv32_fs523_not1 & f_arrdiv32_fs522_or0;
  assign f_arrdiv32_fs523_or0 = f_arrdiv32_fs523_and1 | f_arrdiv32_fs523_and0;
  assign f_arrdiv32_fs524_xor0 = f_arrdiv32_mux2to1476_xor0 ^ b[12];
  assign f_arrdiv32_fs524_not0 = ~f_arrdiv32_mux2to1476_xor0;
  assign f_arrdiv32_fs524_and0 = f_arrdiv32_fs524_not0 & b[12];
  assign f_arrdiv32_fs524_xor1 = f_arrdiv32_fs523_or0 ^ f_arrdiv32_fs524_xor0;
  assign f_arrdiv32_fs524_not1 = ~f_arrdiv32_fs524_xor0;
  assign f_arrdiv32_fs524_and1 = f_arrdiv32_fs524_not1 & f_arrdiv32_fs523_or0;
  assign f_arrdiv32_fs524_or0 = f_arrdiv32_fs524_and1 | f_arrdiv32_fs524_and0;
  assign f_arrdiv32_fs525_xor0 = f_arrdiv32_mux2to1477_xor0 ^ b[13];
  assign f_arrdiv32_fs525_not0 = ~f_arrdiv32_mux2to1477_xor0;
  assign f_arrdiv32_fs525_and0 = f_arrdiv32_fs525_not0 & b[13];
  assign f_arrdiv32_fs525_xor1 = f_arrdiv32_fs524_or0 ^ f_arrdiv32_fs525_xor0;
  assign f_arrdiv32_fs525_not1 = ~f_arrdiv32_fs525_xor0;
  assign f_arrdiv32_fs525_and1 = f_arrdiv32_fs525_not1 & f_arrdiv32_fs524_or0;
  assign f_arrdiv32_fs525_or0 = f_arrdiv32_fs525_and1 | f_arrdiv32_fs525_and0;
  assign f_arrdiv32_fs526_xor0 = f_arrdiv32_mux2to1478_xor0 ^ b[14];
  assign f_arrdiv32_fs526_not0 = ~f_arrdiv32_mux2to1478_xor0;
  assign f_arrdiv32_fs526_and0 = f_arrdiv32_fs526_not0 & b[14];
  assign f_arrdiv32_fs526_xor1 = f_arrdiv32_fs525_or0 ^ f_arrdiv32_fs526_xor0;
  assign f_arrdiv32_fs526_not1 = ~f_arrdiv32_fs526_xor0;
  assign f_arrdiv32_fs526_and1 = f_arrdiv32_fs526_not1 & f_arrdiv32_fs525_or0;
  assign f_arrdiv32_fs526_or0 = f_arrdiv32_fs526_and1 | f_arrdiv32_fs526_and0;
  assign f_arrdiv32_fs527_xor0 = f_arrdiv32_mux2to1479_xor0 ^ b[15];
  assign f_arrdiv32_fs527_not0 = ~f_arrdiv32_mux2to1479_xor0;
  assign f_arrdiv32_fs527_and0 = f_arrdiv32_fs527_not0 & b[15];
  assign f_arrdiv32_fs527_xor1 = f_arrdiv32_fs526_or0 ^ f_arrdiv32_fs527_xor0;
  assign f_arrdiv32_fs527_not1 = ~f_arrdiv32_fs527_xor0;
  assign f_arrdiv32_fs527_and1 = f_arrdiv32_fs527_not1 & f_arrdiv32_fs526_or0;
  assign f_arrdiv32_fs527_or0 = f_arrdiv32_fs527_and1 | f_arrdiv32_fs527_and0;
  assign f_arrdiv32_fs528_xor0 = f_arrdiv32_mux2to1480_xor0 ^ b[16];
  assign f_arrdiv32_fs528_not0 = ~f_arrdiv32_mux2to1480_xor0;
  assign f_arrdiv32_fs528_and0 = f_arrdiv32_fs528_not0 & b[16];
  assign f_arrdiv32_fs528_xor1 = f_arrdiv32_fs527_or0 ^ f_arrdiv32_fs528_xor0;
  assign f_arrdiv32_fs528_not1 = ~f_arrdiv32_fs528_xor0;
  assign f_arrdiv32_fs528_and1 = f_arrdiv32_fs528_not1 & f_arrdiv32_fs527_or0;
  assign f_arrdiv32_fs528_or0 = f_arrdiv32_fs528_and1 | f_arrdiv32_fs528_and0;
  assign f_arrdiv32_fs529_xor0 = f_arrdiv32_mux2to1481_xor0 ^ b[17];
  assign f_arrdiv32_fs529_not0 = ~f_arrdiv32_mux2to1481_xor0;
  assign f_arrdiv32_fs529_and0 = f_arrdiv32_fs529_not0 & b[17];
  assign f_arrdiv32_fs529_xor1 = f_arrdiv32_fs528_or0 ^ f_arrdiv32_fs529_xor0;
  assign f_arrdiv32_fs529_not1 = ~f_arrdiv32_fs529_xor0;
  assign f_arrdiv32_fs529_and1 = f_arrdiv32_fs529_not1 & f_arrdiv32_fs528_or0;
  assign f_arrdiv32_fs529_or0 = f_arrdiv32_fs529_and1 | f_arrdiv32_fs529_and0;
  assign f_arrdiv32_fs530_xor0 = f_arrdiv32_mux2to1482_xor0 ^ b[18];
  assign f_arrdiv32_fs530_not0 = ~f_arrdiv32_mux2to1482_xor0;
  assign f_arrdiv32_fs530_and0 = f_arrdiv32_fs530_not0 & b[18];
  assign f_arrdiv32_fs530_xor1 = f_arrdiv32_fs529_or0 ^ f_arrdiv32_fs530_xor0;
  assign f_arrdiv32_fs530_not1 = ~f_arrdiv32_fs530_xor0;
  assign f_arrdiv32_fs530_and1 = f_arrdiv32_fs530_not1 & f_arrdiv32_fs529_or0;
  assign f_arrdiv32_fs530_or0 = f_arrdiv32_fs530_and1 | f_arrdiv32_fs530_and0;
  assign f_arrdiv32_fs531_xor0 = f_arrdiv32_mux2to1483_xor0 ^ b[19];
  assign f_arrdiv32_fs531_not0 = ~f_arrdiv32_mux2to1483_xor0;
  assign f_arrdiv32_fs531_and0 = f_arrdiv32_fs531_not0 & b[19];
  assign f_arrdiv32_fs531_xor1 = f_arrdiv32_fs530_or0 ^ f_arrdiv32_fs531_xor0;
  assign f_arrdiv32_fs531_not1 = ~f_arrdiv32_fs531_xor0;
  assign f_arrdiv32_fs531_and1 = f_arrdiv32_fs531_not1 & f_arrdiv32_fs530_or0;
  assign f_arrdiv32_fs531_or0 = f_arrdiv32_fs531_and1 | f_arrdiv32_fs531_and0;
  assign f_arrdiv32_fs532_xor0 = f_arrdiv32_mux2to1484_xor0 ^ b[20];
  assign f_arrdiv32_fs532_not0 = ~f_arrdiv32_mux2to1484_xor0;
  assign f_arrdiv32_fs532_and0 = f_arrdiv32_fs532_not0 & b[20];
  assign f_arrdiv32_fs532_xor1 = f_arrdiv32_fs531_or0 ^ f_arrdiv32_fs532_xor0;
  assign f_arrdiv32_fs532_not1 = ~f_arrdiv32_fs532_xor0;
  assign f_arrdiv32_fs532_and1 = f_arrdiv32_fs532_not1 & f_arrdiv32_fs531_or0;
  assign f_arrdiv32_fs532_or0 = f_arrdiv32_fs532_and1 | f_arrdiv32_fs532_and0;
  assign f_arrdiv32_fs533_xor0 = f_arrdiv32_mux2to1485_xor0 ^ b[21];
  assign f_arrdiv32_fs533_not0 = ~f_arrdiv32_mux2to1485_xor0;
  assign f_arrdiv32_fs533_and0 = f_arrdiv32_fs533_not0 & b[21];
  assign f_arrdiv32_fs533_xor1 = f_arrdiv32_fs532_or0 ^ f_arrdiv32_fs533_xor0;
  assign f_arrdiv32_fs533_not1 = ~f_arrdiv32_fs533_xor0;
  assign f_arrdiv32_fs533_and1 = f_arrdiv32_fs533_not1 & f_arrdiv32_fs532_or0;
  assign f_arrdiv32_fs533_or0 = f_arrdiv32_fs533_and1 | f_arrdiv32_fs533_and0;
  assign f_arrdiv32_fs534_xor0 = f_arrdiv32_mux2to1486_xor0 ^ b[22];
  assign f_arrdiv32_fs534_not0 = ~f_arrdiv32_mux2to1486_xor0;
  assign f_arrdiv32_fs534_and0 = f_arrdiv32_fs534_not0 & b[22];
  assign f_arrdiv32_fs534_xor1 = f_arrdiv32_fs533_or0 ^ f_arrdiv32_fs534_xor0;
  assign f_arrdiv32_fs534_not1 = ~f_arrdiv32_fs534_xor0;
  assign f_arrdiv32_fs534_and1 = f_arrdiv32_fs534_not1 & f_arrdiv32_fs533_or0;
  assign f_arrdiv32_fs534_or0 = f_arrdiv32_fs534_and1 | f_arrdiv32_fs534_and0;
  assign f_arrdiv32_fs535_xor0 = f_arrdiv32_mux2to1487_xor0 ^ b[23];
  assign f_arrdiv32_fs535_not0 = ~f_arrdiv32_mux2to1487_xor0;
  assign f_arrdiv32_fs535_and0 = f_arrdiv32_fs535_not0 & b[23];
  assign f_arrdiv32_fs535_xor1 = f_arrdiv32_fs534_or0 ^ f_arrdiv32_fs535_xor0;
  assign f_arrdiv32_fs535_not1 = ~f_arrdiv32_fs535_xor0;
  assign f_arrdiv32_fs535_and1 = f_arrdiv32_fs535_not1 & f_arrdiv32_fs534_or0;
  assign f_arrdiv32_fs535_or0 = f_arrdiv32_fs535_and1 | f_arrdiv32_fs535_and0;
  assign f_arrdiv32_fs536_xor0 = f_arrdiv32_mux2to1488_xor0 ^ b[24];
  assign f_arrdiv32_fs536_not0 = ~f_arrdiv32_mux2to1488_xor0;
  assign f_arrdiv32_fs536_and0 = f_arrdiv32_fs536_not0 & b[24];
  assign f_arrdiv32_fs536_xor1 = f_arrdiv32_fs535_or0 ^ f_arrdiv32_fs536_xor0;
  assign f_arrdiv32_fs536_not1 = ~f_arrdiv32_fs536_xor0;
  assign f_arrdiv32_fs536_and1 = f_arrdiv32_fs536_not1 & f_arrdiv32_fs535_or0;
  assign f_arrdiv32_fs536_or0 = f_arrdiv32_fs536_and1 | f_arrdiv32_fs536_and0;
  assign f_arrdiv32_fs537_xor0 = f_arrdiv32_mux2to1489_xor0 ^ b[25];
  assign f_arrdiv32_fs537_not0 = ~f_arrdiv32_mux2to1489_xor0;
  assign f_arrdiv32_fs537_and0 = f_arrdiv32_fs537_not0 & b[25];
  assign f_arrdiv32_fs537_xor1 = f_arrdiv32_fs536_or0 ^ f_arrdiv32_fs537_xor0;
  assign f_arrdiv32_fs537_not1 = ~f_arrdiv32_fs537_xor0;
  assign f_arrdiv32_fs537_and1 = f_arrdiv32_fs537_not1 & f_arrdiv32_fs536_or0;
  assign f_arrdiv32_fs537_or0 = f_arrdiv32_fs537_and1 | f_arrdiv32_fs537_and0;
  assign f_arrdiv32_fs538_xor0 = f_arrdiv32_mux2to1490_xor0 ^ b[26];
  assign f_arrdiv32_fs538_not0 = ~f_arrdiv32_mux2to1490_xor0;
  assign f_arrdiv32_fs538_and0 = f_arrdiv32_fs538_not0 & b[26];
  assign f_arrdiv32_fs538_xor1 = f_arrdiv32_fs537_or0 ^ f_arrdiv32_fs538_xor0;
  assign f_arrdiv32_fs538_not1 = ~f_arrdiv32_fs538_xor0;
  assign f_arrdiv32_fs538_and1 = f_arrdiv32_fs538_not1 & f_arrdiv32_fs537_or0;
  assign f_arrdiv32_fs538_or0 = f_arrdiv32_fs538_and1 | f_arrdiv32_fs538_and0;
  assign f_arrdiv32_fs539_xor0 = f_arrdiv32_mux2to1491_xor0 ^ b[27];
  assign f_arrdiv32_fs539_not0 = ~f_arrdiv32_mux2to1491_xor0;
  assign f_arrdiv32_fs539_and0 = f_arrdiv32_fs539_not0 & b[27];
  assign f_arrdiv32_fs539_xor1 = f_arrdiv32_fs538_or0 ^ f_arrdiv32_fs539_xor0;
  assign f_arrdiv32_fs539_not1 = ~f_arrdiv32_fs539_xor0;
  assign f_arrdiv32_fs539_and1 = f_arrdiv32_fs539_not1 & f_arrdiv32_fs538_or0;
  assign f_arrdiv32_fs539_or0 = f_arrdiv32_fs539_and1 | f_arrdiv32_fs539_and0;
  assign f_arrdiv32_fs540_xor0 = f_arrdiv32_mux2to1492_xor0 ^ b[28];
  assign f_arrdiv32_fs540_not0 = ~f_arrdiv32_mux2to1492_xor0;
  assign f_arrdiv32_fs540_and0 = f_arrdiv32_fs540_not0 & b[28];
  assign f_arrdiv32_fs540_xor1 = f_arrdiv32_fs539_or0 ^ f_arrdiv32_fs540_xor0;
  assign f_arrdiv32_fs540_not1 = ~f_arrdiv32_fs540_xor0;
  assign f_arrdiv32_fs540_and1 = f_arrdiv32_fs540_not1 & f_arrdiv32_fs539_or0;
  assign f_arrdiv32_fs540_or0 = f_arrdiv32_fs540_and1 | f_arrdiv32_fs540_and0;
  assign f_arrdiv32_fs541_xor0 = f_arrdiv32_mux2to1493_xor0 ^ b[29];
  assign f_arrdiv32_fs541_not0 = ~f_arrdiv32_mux2to1493_xor0;
  assign f_arrdiv32_fs541_and0 = f_arrdiv32_fs541_not0 & b[29];
  assign f_arrdiv32_fs541_xor1 = f_arrdiv32_fs540_or0 ^ f_arrdiv32_fs541_xor0;
  assign f_arrdiv32_fs541_not1 = ~f_arrdiv32_fs541_xor0;
  assign f_arrdiv32_fs541_and1 = f_arrdiv32_fs541_not1 & f_arrdiv32_fs540_or0;
  assign f_arrdiv32_fs541_or0 = f_arrdiv32_fs541_and1 | f_arrdiv32_fs541_and0;
  assign f_arrdiv32_fs542_xor0 = f_arrdiv32_mux2to1494_xor0 ^ b[30];
  assign f_arrdiv32_fs542_not0 = ~f_arrdiv32_mux2to1494_xor0;
  assign f_arrdiv32_fs542_and0 = f_arrdiv32_fs542_not0 & b[30];
  assign f_arrdiv32_fs542_xor1 = f_arrdiv32_fs541_or0 ^ f_arrdiv32_fs542_xor0;
  assign f_arrdiv32_fs542_not1 = ~f_arrdiv32_fs542_xor0;
  assign f_arrdiv32_fs542_and1 = f_arrdiv32_fs542_not1 & f_arrdiv32_fs541_or0;
  assign f_arrdiv32_fs542_or0 = f_arrdiv32_fs542_and1 | f_arrdiv32_fs542_and0;
  assign f_arrdiv32_fs543_xor0 = f_arrdiv32_mux2to1495_xor0 ^ b[31];
  assign f_arrdiv32_fs543_not0 = ~f_arrdiv32_mux2to1495_xor0;
  assign f_arrdiv32_fs543_and0 = f_arrdiv32_fs543_not0 & b[31];
  assign f_arrdiv32_fs543_xor1 = f_arrdiv32_fs542_or0 ^ f_arrdiv32_fs543_xor0;
  assign f_arrdiv32_fs543_not1 = ~f_arrdiv32_fs543_xor0;
  assign f_arrdiv32_fs543_and1 = f_arrdiv32_fs543_not1 & f_arrdiv32_fs542_or0;
  assign f_arrdiv32_fs543_or0 = f_arrdiv32_fs543_and1 | f_arrdiv32_fs543_and0;
  assign f_arrdiv32_mux2to1496_and0 = a[15] & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1496_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1496_and1 = f_arrdiv32_fs512_xor0 & f_arrdiv32_mux2to1496_not0;
  assign f_arrdiv32_mux2to1496_xor0 = f_arrdiv32_mux2to1496_and0 ^ f_arrdiv32_mux2to1496_and1;
  assign f_arrdiv32_mux2to1497_and0 = f_arrdiv32_mux2to1465_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1497_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1497_and1 = f_arrdiv32_fs513_xor1 & f_arrdiv32_mux2to1497_not0;
  assign f_arrdiv32_mux2to1497_xor0 = f_arrdiv32_mux2to1497_and0 ^ f_arrdiv32_mux2to1497_and1;
  assign f_arrdiv32_mux2to1498_and0 = f_arrdiv32_mux2to1466_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1498_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1498_and1 = f_arrdiv32_fs514_xor1 & f_arrdiv32_mux2to1498_not0;
  assign f_arrdiv32_mux2to1498_xor0 = f_arrdiv32_mux2to1498_and0 ^ f_arrdiv32_mux2to1498_and1;
  assign f_arrdiv32_mux2to1499_and0 = f_arrdiv32_mux2to1467_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1499_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1499_and1 = f_arrdiv32_fs515_xor1 & f_arrdiv32_mux2to1499_not0;
  assign f_arrdiv32_mux2to1499_xor0 = f_arrdiv32_mux2to1499_and0 ^ f_arrdiv32_mux2to1499_and1;
  assign f_arrdiv32_mux2to1500_and0 = f_arrdiv32_mux2to1468_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1500_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1500_and1 = f_arrdiv32_fs516_xor1 & f_arrdiv32_mux2to1500_not0;
  assign f_arrdiv32_mux2to1500_xor0 = f_arrdiv32_mux2to1500_and0 ^ f_arrdiv32_mux2to1500_and1;
  assign f_arrdiv32_mux2to1501_and0 = f_arrdiv32_mux2to1469_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1501_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1501_and1 = f_arrdiv32_fs517_xor1 & f_arrdiv32_mux2to1501_not0;
  assign f_arrdiv32_mux2to1501_xor0 = f_arrdiv32_mux2to1501_and0 ^ f_arrdiv32_mux2to1501_and1;
  assign f_arrdiv32_mux2to1502_and0 = f_arrdiv32_mux2to1470_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1502_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1502_and1 = f_arrdiv32_fs518_xor1 & f_arrdiv32_mux2to1502_not0;
  assign f_arrdiv32_mux2to1502_xor0 = f_arrdiv32_mux2to1502_and0 ^ f_arrdiv32_mux2to1502_and1;
  assign f_arrdiv32_mux2to1503_and0 = f_arrdiv32_mux2to1471_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1503_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1503_and1 = f_arrdiv32_fs519_xor1 & f_arrdiv32_mux2to1503_not0;
  assign f_arrdiv32_mux2to1503_xor0 = f_arrdiv32_mux2to1503_and0 ^ f_arrdiv32_mux2to1503_and1;
  assign f_arrdiv32_mux2to1504_and0 = f_arrdiv32_mux2to1472_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1504_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1504_and1 = f_arrdiv32_fs520_xor1 & f_arrdiv32_mux2to1504_not0;
  assign f_arrdiv32_mux2to1504_xor0 = f_arrdiv32_mux2to1504_and0 ^ f_arrdiv32_mux2to1504_and1;
  assign f_arrdiv32_mux2to1505_and0 = f_arrdiv32_mux2to1473_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1505_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1505_and1 = f_arrdiv32_fs521_xor1 & f_arrdiv32_mux2to1505_not0;
  assign f_arrdiv32_mux2to1505_xor0 = f_arrdiv32_mux2to1505_and0 ^ f_arrdiv32_mux2to1505_and1;
  assign f_arrdiv32_mux2to1506_and0 = f_arrdiv32_mux2to1474_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1506_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1506_and1 = f_arrdiv32_fs522_xor1 & f_arrdiv32_mux2to1506_not0;
  assign f_arrdiv32_mux2to1506_xor0 = f_arrdiv32_mux2to1506_and0 ^ f_arrdiv32_mux2to1506_and1;
  assign f_arrdiv32_mux2to1507_and0 = f_arrdiv32_mux2to1475_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1507_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1507_and1 = f_arrdiv32_fs523_xor1 & f_arrdiv32_mux2to1507_not0;
  assign f_arrdiv32_mux2to1507_xor0 = f_arrdiv32_mux2to1507_and0 ^ f_arrdiv32_mux2to1507_and1;
  assign f_arrdiv32_mux2to1508_and0 = f_arrdiv32_mux2to1476_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1508_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1508_and1 = f_arrdiv32_fs524_xor1 & f_arrdiv32_mux2to1508_not0;
  assign f_arrdiv32_mux2to1508_xor0 = f_arrdiv32_mux2to1508_and0 ^ f_arrdiv32_mux2to1508_and1;
  assign f_arrdiv32_mux2to1509_and0 = f_arrdiv32_mux2to1477_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1509_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1509_and1 = f_arrdiv32_fs525_xor1 & f_arrdiv32_mux2to1509_not0;
  assign f_arrdiv32_mux2to1509_xor0 = f_arrdiv32_mux2to1509_and0 ^ f_arrdiv32_mux2to1509_and1;
  assign f_arrdiv32_mux2to1510_and0 = f_arrdiv32_mux2to1478_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1510_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1510_and1 = f_arrdiv32_fs526_xor1 & f_arrdiv32_mux2to1510_not0;
  assign f_arrdiv32_mux2to1510_xor0 = f_arrdiv32_mux2to1510_and0 ^ f_arrdiv32_mux2to1510_and1;
  assign f_arrdiv32_mux2to1511_and0 = f_arrdiv32_mux2to1479_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1511_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1511_and1 = f_arrdiv32_fs527_xor1 & f_arrdiv32_mux2to1511_not0;
  assign f_arrdiv32_mux2to1511_xor0 = f_arrdiv32_mux2to1511_and0 ^ f_arrdiv32_mux2to1511_and1;
  assign f_arrdiv32_mux2to1512_and0 = f_arrdiv32_mux2to1480_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1512_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1512_and1 = f_arrdiv32_fs528_xor1 & f_arrdiv32_mux2to1512_not0;
  assign f_arrdiv32_mux2to1512_xor0 = f_arrdiv32_mux2to1512_and0 ^ f_arrdiv32_mux2to1512_and1;
  assign f_arrdiv32_mux2to1513_and0 = f_arrdiv32_mux2to1481_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1513_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1513_and1 = f_arrdiv32_fs529_xor1 & f_arrdiv32_mux2to1513_not0;
  assign f_arrdiv32_mux2to1513_xor0 = f_arrdiv32_mux2to1513_and0 ^ f_arrdiv32_mux2to1513_and1;
  assign f_arrdiv32_mux2to1514_and0 = f_arrdiv32_mux2to1482_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1514_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1514_and1 = f_arrdiv32_fs530_xor1 & f_arrdiv32_mux2to1514_not0;
  assign f_arrdiv32_mux2to1514_xor0 = f_arrdiv32_mux2to1514_and0 ^ f_arrdiv32_mux2to1514_and1;
  assign f_arrdiv32_mux2to1515_and0 = f_arrdiv32_mux2to1483_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1515_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1515_and1 = f_arrdiv32_fs531_xor1 & f_arrdiv32_mux2to1515_not0;
  assign f_arrdiv32_mux2to1515_xor0 = f_arrdiv32_mux2to1515_and0 ^ f_arrdiv32_mux2to1515_and1;
  assign f_arrdiv32_mux2to1516_and0 = f_arrdiv32_mux2to1484_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1516_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1516_and1 = f_arrdiv32_fs532_xor1 & f_arrdiv32_mux2to1516_not0;
  assign f_arrdiv32_mux2to1516_xor0 = f_arrdiv32_mux2to1516_and0 ^ f_arrdiv32_mux2to1516_and1;
  assign f_arrdiv32_mux2to1517_and0 = f_arrdiv32_mux2to1485_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1517_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1517_and1 = f_arrdiv32_fs533_xor1 & f_arrdiv32_mux2to1517_not0;
  assign f_arrdiv32_mux2to1517_xor0 = f_arrdiv32_mux2to1517_and0 ^ f_arrdiv32_mux2to1517_and1;
  assign f_arrdiv32_mux2to1518_and0 = f_arrdiv32_mux2to1486_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1518_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1518_and1 = f_arrdiv32_fs534_xor1 & f_arrdiv32_mux2to1518_not0;
  assign f_arrdiv32_mux2to1518_xor0 = f_arrdiv32_mux2to1518_and0 ^ f_arrdiv32_mux2to1518_and1;
  assign f_arrdiv32_mux2to1519_and0 = f_arrdiv32_mux2to1487_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1519_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1519_and1 = f_arrdiv32_fs535_xor1 & f_arrdiv32_mux2to1519_not0;
  assign f_arrdiv32_mux2to1519_xor0 = f_arrdiv32_mux2to1519_and0 ^ f_arrdiv32_mux2to1519_and1;
  assign f_arrdiv32_mux2to1520_and0 = f_arrdiv32_mux2to1488_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1520_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1520_and1 = f_arrdiv32_fs536_xor1 & f_arrdiv32_mux2to1520_not0;
  assign f_arrdiv32_mux2to1520_xor0 = f_arrdiv32_mux2to1520_and0 ^ f_arrdiv32_mux2to1520_and1;
  assign f_arrdiv32_mux2to1521_and0 = f_arrdiv32_mux2to1489_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1521_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1521_and1 = f_arrdiv32_fs537_xor1 & f_arrdiv32_mux2to1521_not0;
  assign f_arrdiv32_mux2to1521_xor0 = f_arrdiv32_mux2to1521_and0 ^ f_arrdiv32_mux2to1521_and1;
  assign f_arrdiv32_mux2to1522_and0 = f_arrdiv32_mux2to1490_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1522_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1522_and1 = f_arrdiv32_fs538_xor1 & f_arrdiv32_mux2to1522_not0;
  assign f_arrdiv32_mux2to1522_xor0 = f_arrdiv32_mux2to1522_and0 ^ f_arrdiv32_mux2to1522_and1;
  assign f_arrdiv32_mux2to1523_and0 = f_arrdiv32_mux2to1491_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1523_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1523_and1 = f_arrdiv32_fs539_xor1 & f_arrdiv32_mux2to1523_not0;
  assign f_arrdiv32_mux2to1523_xor0 = f_arrdiv32_mux2to1523_and0 ^ f_arrdiv32_mux2to1523_and1;
  assign f_arrdiv32_mux2to1524_and0 = f_arrdiv32_mux2to1492_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1524_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1524_and1 = f_arrdiv32_fs540_xor1 & f_arrdiv32_mux2to1524_not0;
  assign f_arrdiv32_mux2to1524_xor0 = f_arrdiv32_mux2to1524_and0 ^ f_arrdiv32_mux2to1524_and1;
  assign f_arrdiv32_mux2to1525_and0 = f_arrdiv32_mux2to1493_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1525_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1525_and1 = f_arrdiv32_fs541_xor1 & f_arrdiv32_mux2to1525_not0;
  assign f_arrdiv32_mux2to1525_xor0 = f_arrdiv32_mux2to1525_and0 ^ f_arrdiv32_mux2to1525_and1;
  assign f_arrdiv32_mux2to1526_and0 = f_arrdiv32_mux2to1494_xor0 & f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1526_not0 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_mux2to1526_and1 = f_arrdiv32_fs542_xor1 & f_arrdiv32_mux2to1526_not0;
  assign f_arrdiv32_mux2to1526_xor0 = f_arrdiv32_mux2to1526_and0 ^ f_arrdiv32_mux2to1526_and1;
  assign f_arrdiv32_not16 = ~f_arrdiv32_fs543_or0;
  assign f_arrdiv32_fs544_xor0 = a[14] ^ b[0];
  assign f_arrdiv32_fs544_not0 = ~a[14];
  assign f_arrdiv32_fs544_and0 = f_arrdiv32_fs544_not0 & b[0];
  assign f_arrdiv32_fs544_not1 = ~f_arrdiv32_fs544_xor0;
  assign f_arrdiv32_fs545_xor0 = f_arrdiv32_mux2to1496_xor0 ^ b[1];
  assign f_arrdiv32_fs545_not0 = ~f_arrdiv32_mux2to1496_xor0;
  assign f_arrdiv32_fs545_and0 = f_arrdiv32_fs545_not0 & b[1];
  assign f_arrdiv32_fs545_xor1 = f_arrdiv32_fs544_and0 ^ f_arrdiv32_fs545_xor0;
  assign f_arrdiv32_fs545_not1 = ~f_arrdiv32_fs545_xor0;
  assign f_arrdiv32_fs545_and1 = f_arrdiv32_fs545_not1 & f_arrdiv32_fs544_and0;
  assign f_arrdiv32_fs545_or0 = f_arrdiv32_fs545_and1 | f_arrdiv32_fs545_and0;
  assign f_arrdiv32_fs546_xor0 = f_arrdiv32_mux2to1497_xor0 ^ b[2];
  assign f_arrdiv32_fs546_not0 = ~f_arrdiv32_mux2to1497_xor0;
  assign f_arrdiv32_fs546_and0 = f_arrdiv32_fs546_not0 & b[2];
  assign f_arrdiv32_fs546_xor1 = f_arrdiv32_fs545_or0 ^ f_arrdiv32_fs546_xor0;
  assign f_arrdiv32_fs546_not1 = ~f_arrdiv32_fs546_xor0;
  assign f_arrdiv32_fs546_and1 = f_arrdiv32_fs546_not1 & f_arrdiv32_fs545_or0;
  assign f_arrdiv32_fs546_or0 = f_arrdiv32_fs546_and1 | f_arrdiv32_fs546_and0;
  assign f_arrdiv32_fs547_xor0 = f_arrdiv32_mux2to1498_xor0 ^ b[3];
  assign f_arrdiv32_fs547_not0 = ~f_arrdiv32_mux2to1498_xor0;
  assign f_arrdiv32_fs547_and0 = f_arrdiv32_fs547_not0 & b[3];
  assign f_arrdiv32_fs547_xor1 = f_arrdiv32_fs546_or0 ^ f_arrdiv32_fs547_xor0;
  assign f_arrdiv32_fs547_not1 = ~f_arrdiv32_fs547_xor0;
  assign f_arrdiv32_fs547_and1 = f_arrdiv32_fs547_not1 & f_arrdiv32_fs546_or0;
  assign f_arrdiv32_fs547_or0 = f_arrdiv32_fs547_and1 | f_arrdiv32_fs547_and0;
  assign f_arrdiv32_fs548_xor0 = f_arrdiv32_mux2to1499_xor0 ^ b[4];
  assign f_arrdiv32_fs548_not0 = ~f_arrdiv32_mux2to1499_xor0;
  assign f_arrdiv32_fs548_and0 = f_arrdiv32_fs548_not0 & b[4];
  assign f_arrdiv32_fs548_xor1 = f_arrdiv32_fs547_or0 ^ f_arrdiv32_fs548_xor0;
  assign f_arrdiv32_fs548_not1 = ~f_arrdiv32_fs548_xor0;
  assign f_arrdiv32_fs548_and1 = f_arrdiv32_fs548_not1 & f_arrdiv32_fs547_or0;
  assign f_arrdiv32_fs548_or0 = f_arrdiv32_fs548_and1 | f_arrdiv32_fs548_and0;
  assign f_arrdiv32_fs549_xor0 = f_arrdiv32_mux2to1500_xor0 ^ b[5];
  assign f_arrdiv32_fs549_not0 = ~f_arrdiv32_mux2to1500_xor0;
  assign f_arrdiv32_fs549_and0 = f_arrdiv32_fs549_not0 & b[5];
  assign f_arrdiv32_fs549_xor1 = f_arrdiv32_fs548_or0 ^ f_arrdiv32_fs549_xor0;
  assign f_arrdiv32_fs549_not1 = ~f_arrdiv32_fs549_xor0;
  assign f_arrdiv32_fs549_and1 = f_arrdiv32_fs549_not1 & f_arrdiv32_fs548_or0;
  assign f_arrdiv32_fs549_or0 = f_arrdiv32_fs549_and1 | f_arrdiv32_fs549_and0;
  assign f_arrdiv32_fs550_xor0 = f_arrdiv32_mux2to1501_xor0 ^ b[6];
  assign f_arrdiv32_fs550_not0 = ~f_arrdiv32_mux2to1501_xor0;
  assign f_arrdiv32_fs550_and0 = f_arrdiv32_fs550_not0 & b[6];
  assign f_arrdiv32_fs550_xor1 = f_arrdiv32_fs549_or0 ^ f_arrdiv32_fs550_xor0;
  assign f_arrdiv32_fs550_not1 = ~f_arrdiv32_fs550_xor0;
  assign f_arrdiv32_fs550_and1 = f_arrdiv32_fs550_not1 & f_arrdiv32_fs549_or0;
  assign f_arrdiv32_fs550_or0 = f_arrdiv32_fs550_and1 | f_arrdiv32_fs550_and0;
  assign f_arrdiv32_fs551_xor0 = f_arrdiv32_mux2to1502_xor0 ^ b[7];
  assign f_arrdiv32_fs551_not0 = ~f_arrdiv32_mux2to1502_xor0;
  assign f_arrdiv32_fs551_and0 = f_arrdiv32_fs551_not0 & b[7];
  assign f_arrdiv32_fs551_xor1 = f_arrdiv32_fs550_or0 ^ f_arrdiv32_fs551_xor0;
  assign f_arrdiv32_fs551_not1 = ~f_arrdiv32_fs551_xor0;
  assign f_arrdiv32_fs551_and1 = f_arrdiv32_fs551_not1 & f_arrdiv32_fs550_or0;
  assign f_arrdiv32_fs551_or0 = f_arrdiv32_fs551_and1 | f_arrdiv32_fs551_and0;
  assign f_arrdiv32_fs552_xor0 = f_arrdiv32_mux2to1503_xor0 ^ b[8];
  assign f_arrdiv32_fs552_not0 = ~f_arrdiv32_mux2to1503_xor0;
  assign f_arrdiv32_fs552_and0 = f_arrdiv32_fs552_not0 & b[8];
  assign f_arrdiv32_fs552_xor1 = f_arrdiv32_fs551_or0 ^ f_arrdiv32_fs552_xor0;
  assign f_arrdiv32_fs552_not1 = ~f_arrdiv32_fs552_xor0;
  assign f_arrdiv32_fs552_and1 = f_arrdiv32_fs552_not1 & f_arrdiv32_fs551_or0;
  assign f_arrdiv32_fs552_or0 = f_arrdiv32_fs552_and1 | f_arrdiv32_fs552_and0;
  assign f_arrdiv32_fs553_xor0 = f_arrdiv32_mux2to1504_xor0 ^ b[9];
  assign f_arrdiv32_fs553_not0 = ~f_arrdiv32_mux2to1504_xor0;
  assign f_arrdiv32_fs553_and0 = f_arrdiv32_fs553_not0 & b[9];
  assign f_arrdiv32_fs553_xor1 = f_arrdiv32_fs552_or0 ^ f_arrdiv32_fs553_xor0;
  assign f_arrdiv32_fs553_not1 = ~f_arrdiv32_fs553_xor0;
  assign f_arrdiv32_fs553_and1 = f_arrdiv32_fs553_not1 & f_arrdiv32_fs552_or0;
  assign f_arrdiv32_fs553_or0 = f_arrdiv32_fs553_and1 | f_arrdiv32_fs553_and0;
  assign f_arrdiv32_fs554_xor0 = f_arrdiv32_mux2to1505_xor0 ^ b[10];
  assign f_arrdiv32_fs554_not0 = ~f_arrdiv32_mux2to1505_xor0;
  assign f_arrdiv32_fs554_and0 = f_arrdiv32_fs554_not0 & b[10];
  assign f_arrdiv32_fs554_xor1 = f_arrdiv32_fs553_or0 ^ f_arrdiv32_fs554_xor0;
  assign f_arrdiv32_fs554_not1 = ~f_arrdiv32_fs554_xor0;
  assign f_arrdiv32_fs554_and1 = f_arrdiv32_fs554_not1 & f_arrdiv32_fs553_or0;
  assign f_arrdiv32_fs554_or0 = f_arrdiv32_fs554_and1 | f_arrdiv32_fs554_and0;
  assign f_arrdiv32_fs555_xor0 = f_arrdiv32_mux2to1506_xor0 ^ b[11];
  assign f_arrdiv32_fs555_not0 = ~f_arrdiv32_mux2to1506_xor0;
  assign f_arrdiv32_fs555_and0 = f_arrdiv32_fs555_not0 & b[11];
  assign f_arrdiv32_fs555_xor1 = f_arrdiv32_fs554_or0 ^ f_arrdiv32_fs555_xor0;
  assign f_arrdiv32_fs555_not1 = ~f_arrdiv32_fs555_xor0;
  assign f_arrdiv32_fs555_and1 = f_arrdiv32_fs555_not1 & f_arrdiv32_fs554_or0;
  assign f_arrdiv32_fs555_or0 = f_arrdiv32_fs555_and1 | f_arrdiv32_fs555_and0;
  assign f_arrdiv32_fs556_xor0 = f_arrdiv32_mux2to1507_xor0 ^ b[12];
  assign f_arrdiv32_fs556_not0 = ~f_arrdiv32_mux2to1507_xor0;
  assign f_arrdiv32_fs556_and0 = f_arrdiv32_fs556_not0 & b[12];
  assign f_arrdiv32_fs556_xor1 = f_arrdiv32_fs555_or0 ^ f_arrdiv32_fs556_xor0;
  assign f_arrdiv32_fs556_not1 = ~f_arrdiv32_fs556_xor0;
  assign f_arrdiv32_fs556_and1 = f_arrdiv32_fs556_not1 & f_arrdiv32_fs555_or0;
  assign f_arrdiv32_fs556_or0 = f_arrdiv32_fs556_and1 | f_arrdiv32_fs556_and0;
  assign f_arrdiv32_fs557_xor0 = f_arrdiv32_mux2to1508_xor0 ^ b[13];
  assign f_arrdiv32_fs557_not0 = ~f_arrdiv32_mux2to1508_xor0;
  assign f_arrdiv32_fs557_and0 = f_arrdiv32_fs557_not0 & b[13];
  assign f_arrdiv32_fs557_xor1 = f_arrdiv32_fs556_or0 ^ f_arrdiv32_fs557_xor0;
  assign f_arrdiv32_fs557_not1 = ~f_arrdiv32_fs557_xor0;
  assign f_arrdiv32_fs557_and1 = f_arrdiv32_fs557_not1 & f_arrdiv32_fs556_or0;
  assign f_arrdiv32_fs557_or0 = f_arrdiv32_fs557_and1 | f_arrdiv32_fs557_and0;
  assign f_arrdiv32_fs558_xor0 = f_arrdiv32_mux2to1509_xor0 ^ b[14];
  assign f_arrdiv32_fs558_not0 = ~f_arrdiv32_mux2to1509_xor0;
  assign f_arrdiv32_fs558_and0 = f_arrdiv32_fs558_not0 & b[14];
  assign f_arrdiv32_fs558_xor1 = f_arrdiv32_fs557_or0 ^ f_arrdiv32_fs558_xor0;
  assign f_arrdiv32_fs558_not1 = ~f_arrdiv32_fs558_xor0;
  assign f_arrdiv32_fs558_and1 = f_arrdiv32_fs558_not1 & f_arrdiv32_fs557_or0;
  assign f_arrdiv32_fs558_or0 = f_arrdiv32_fs558_and1 | f_arrdiv32_fs558_and0;
  assign f_arrdiv32_fs559_xor0 = f_arrdiv32_mux2to1510_xor0 ^ b[15];
  assign f_arrdiv32_fs559_not0 = ~f_arrdiv32_mux2to1510_xor0;
  assign f_arrdiv32_fs559_and0 = f_arrdiv32_fs559_not0 & b[15];
  assign f_arrdiv32_fs559_xor1 = f_arrdiv32_fs558_or0 ^ f_arrdiv32_fs559_xor0;
  assign f_arrdiv32_fs559_not1 = ~f_arrdiv32_fs559_xor0;
  assign f_arrdiv32_fs559_and1 = f_arrdiv32_fs559_not1 & f_arrdiv32_fs558_or0;
  assign f_arrdiv32_fs559_or0 = f_arrdiv32_fs559_and1 | f_arrdiv32_fs559_and0;
  assign f_arrdiv32_fs560_xor0 = f_arrdiv32_mux2to1511_xor0 ^ b[16];
  assign f_arrdiv32_fs560_not0 = ~f_arrdiv32_mux2to1511_xor0;
  assign f_arrdiv32_fs560_and0 = f_arrdiv32_fs560_not0 & b[16];
  assign f_arrdiv32_fs560_xor1 = f_arrdiv32_fs559_or0 ^ f_arrdiv32_fs560_xor0;
  assign f_arrdiv32_fs560_not1 = ~f_arrdiv32_fs560_xor0;
  assign f_arrdiv32_fs560_and1 = f_arrdiv32_fs560_not1 & f_arrdiv32_fs559_or0;
  assign f_arrdiv32_fs560_or0 = f_arrdiv32_fs560_and1 | f_arrdiv32_fs560_and0;
  assign f_arrdiv32_fs561_xor0 = f_arrdiv32_mux2to1512_xor0 ^ b[17];
  assign f_arrdiv32_fs561_not0 = ~f_arrdiv32_mux2to1512_xor0;
  assign f_arrdiv32_fs561_and0 = f_arrdiv32_fs561_not0 & b[17];
  assign f_arrdiv32_fs561_xor1 = f_arrdiv32_fs560_or0 ^ f_arrdiv32_fs561_xor0;
  assign f_arrdiv32_fs561_not1 = ~f_arrdiv32_fs561_xor0;
  assign f_arrdiv32_fs561_and1 = f_arrdiv32_fs561_not1 & f_arrdiv32_fs560_or0;
  assign f_arrdiv32_fs561_or0 = f_arrdiv32_fs561_and1 | f_arrdiv32_fs561_and0;
  assign f_arrdiv32_fs562_xor0 = f_arrdiv32_mux2to1513_xor0 ^ b[18];
  assign f_arrdiv32_fs562_not0 = ~f_arrdiv32_mux2to1513_xor0;
  assign f_arrdiv32_fs562_and0 = f_arrdiv32_fs562_not0 & b[18];
  assign f_arrdiv32_fs562_xor1 = f_arrdiv32_fs561_or0 ^ f_arrdiv32_fs562_xor0;
  assign f_arrdiv32_fs562_not1 = ~f_arrdiv32_fs562_xor0;
  assign f_arrdiv32_fs562_and1 = f_arrdiv32_fs562_not1 & f_arrdiv32_fs561_or0;
  assign f_arrdiv32_fs562_or0 = f_arrdiv32_fs562_and1 | f_arrdiv32_fs562_and0;
  assign f_arrdiv32_fs563_xor0 = f_arrdiv32_mux2to1514_xor0 ^ b[19];
  assign f_arrdiv32_fs563_not0 = ~f_arrdiv32_mux2to1514_xor0;
  assign f_arrdiv32_fs563_and0 = f_arrdiv32_fs563_not0 & b[19];
  assign f_arrdiv32_fs563_xor1 = f_arrdiv32_fs562_or0 ^ f_arrdiv32_fs563_xor0;
  assign f_arrdiv32_fs563_not1 = ~f_arrdiv32_fs563_xor0;
  assign f_arrdiv32_fs563_and1 = f_arrdiv32_fs563_not1 & f_arrdiv32_fs562_or0;
  assign f_arrdiv32_fs563_or0 = f_arrdiv32_fs563_and1 | f_arrdiv32_fs563_and0;
  assign f_arrdiv32_fs564_xor0 = f_arrdiv32_mux2to1515_xor0 ^ b[20];
  assign f_arrdiv32_fs564_not0 = ~f_arrdiv32_mux2to1515_xor0;
  assign f_arrdiv32_fs564_and0 = f_arrdiv32_fs564_not0 & b[20];
  assign f_arrdiv32_fs564_xor1 = f_arrdiv32_fs563_or0 ^ f_arrdiv32_fs564_xor0;
  assign f_arrdiv32_fs564_not1 = ~f_arrdiv32_fs564_xor0;
  assign f_arrdiv32_fs564_and1 = f_arrdiv32_fs564_not1 & f_arrdiv32_fs563_or0;
  assign f_arrdiv32_fs564_or0 = f_arrdiv32_fs564_and1 | f_arrdiv32_fs564_and0;
  assign f_arrdiv32_fs565_xor0 = f_arrdiv32_mux2to1516_xor0 ^ b[21];
  assign f_arrdiv32_fs565_not0 = ~f_arrdiv32_mux2to1516_xor0;
  assign f_arrdiv32_fs565_and0 = f_arrdiv32_fs565_not0 & b[21];
  assign f_arrdiv32_fs565_xor1 = f_arrdiv32_fs564_or0 ^ f_arrdiv32_fs565_xor0;
  assign f_arrdiv32_fs565_not1 = ~f_arrdiv32_fs565_xor0;
  assign f_arrdiv32_fs565_and1 = f_arrdiv32_fs565_not1 & f_arrdiv32_fs564_or0;
  assign f_arrdiv32_fs565_or0 = f_arrdiv32_fs565_and1 | f_arrdiv32_fs565_and0;
  assign f_arrdiv32_fs566_xor0 = f_arrdiv32_mux2to1517_xor0 ^ b[22];
  assign f_arrdiv32_fs566_not0 = ~f_arrdiv32_mux2to1517_xor0;
  assign f_arrdiv32_fs566_and0 = f_arrdiv32_fs566_not0 & b[22];
  assign f_arrdiv32_fs566_xor1 = f_arrdiv32_fs565_or0 ^ f_arrdiv32_fs566_xor0;
  assign f_arrdiv32_fs566_not1 = ~f_arrdiv32_fs566_xor0;
  assign f_arrdiv32_fs566_and1 = f_arrdiv32_fs566_not1 & f_arrdiv32_fs565_or0;
  assign f_arrdiv32_fs566_or0 = f_arrdiv32_fs566_and1 | f_arrdiv32_fs566_and0;
  assign f_arrdiv32_fs567_xor0 = f_arrdiv32_mux2to1518_xor0 ^ b[23];
  assign f_arrdiv32_fs567_not0 = ~f_arrdiv32_mux2to1518_xor0;
  assign f_arrdiv32_fs567_and0 = f_arrdiv32_fs567_not0 & b[23];
  assign f_arrdiv32_fs567_xor1 = f_arrdiv32_fs566_or0 ^ f_arrdiv32_fs567_xor0;
  assign f_arrdiv32_fs567_not1 = ~f_arrdiv32_fs567_xor0;
  assign f_arrdiv32_fs567_and1 = f_arrdiv32_fs567_not1 & f_arrdiv32_fs566_or0;
  assign f_arrdiv32_fs567_or0 = f_arrdiv32_fs567_and1 | f_arrdiv32_fs567_and0;
  assign f_arrdiv32_fs568_xor0 = f_arrdiv32_mux2to1519_xor0 ^ b[24];
  assign f_arrdiv32_fs568_not0 = ~f_arrdiv32_mux2to1519_xor0;
  assign f_arrdiv32_fs568_and0 = f_arrdiv32_fs568_not0 & b[24];
  assign f_arrdiv32_fs568_xor1 = f_arrdiv32_fs567_or0 ^ f_arrdiv32_fs568_xor0;
  assign f_arrdiv32_fs568_not1 = ~f_arrdiv32_fs568_xor0;
  assign f_arrdiv32_fs568_and1 = f_arrdiv32_fs568_not1 & f_arrdiv32_fs567_or0;
  assign f_arrdiv32_fs568_or0 = f_arrdiv32_fs568_and1 | f_arrdiv32_fs568_and0;
  assign f_arrdiv32_fs569_xor0 = f_arrdiv32_mux2to1520_xor0 ^ b[25];
  assign f_arrdiv32_fs569_not0 = ~f_arrdiv32_mux2to1520_xor0;
  assign f_arrdiv32_fs569_and0 = f_arrdiv32_fs569_not0 & b[25];
  assign f_arrdiv32_fs569_xor1 = f_arrdiv32_fs568_or0 ^ f_arrdiv32_fs569_xor0;
  assign f_arrdiv32_fs569_not1 = ~f_arrdiv32_fs569_xor0;
  assign f_arrdiv32_fs569_and1 = f_arrdiv32_fs569_not1 & f_arrdiv32_fs568_or0;
  assign f_arrdiv32_fs569_or0 = f_arrdiv32_fs569_and1 | f_arrdiv32_fs569_and0;
  assign f_arrdiv32_fs570_xor0 = f_arrdiv32_mux2to1521_xor0 ^ b[26];
  assign f_arrdiv32_fs570_not0 = ~f_arrdiv32_mux2to1521_xor0;
  assign f_arrdiv32_fs570_and0 = f_arrdiv32_fs570_not0 & b[26];
  assign f_arrdiv32_fs570_xor1 = f_arrdiv32_fs569_or0 ^ f_arrdiv32_fs570_xor0;
  assign f_arrdiv32_fs570_not1 = ~f_arrdiv32_fs570_xor0;
  assign f_arrdiv32_fs570_and1 = f_arrdiv32_fs570_not1 & f_arrdiv32_fs569_or0;
  assign f_arrdiv32_fs570_or0 = f_arrdiv32_fs570_and1 | f_arrdiv32_fs570_and0;
  assign f_arrdiv32_fs571_xor0 = f_arrdiv32_mux2to1522_xor0 ^ b[27];
  assign f_arrdiv32_fs571_not0 = ~f_arrdiv32_mux2to1522_xor0;
  assign f_arrdiv32_fs571_and0 = f_arrdiv32_fs571_not0 & b[27];
  assign f_arrdiv32_fs571_xor1 = f_arrdiv32_fs570_or0 ^ f_arrdiv32_fs571_xor0;
  assign f_arrdiv32_fs571_not1 = ~f_arrdiv32_fs571_xor0;
  assign f_arrdiv32_fs571_and1 = f_arrdiv32_fs571_not1 & f_arrdiv32_fs570_or0;
  assign f_arrdiv32_fs571_or0 = f_arrdiv32_fs571_and1 | f_arrdiv32_fs571_and0;
  assign f_arrdiv32_fs572_xor0 = f_arrdiv32_mux2to1523_xor0 ^ b[28];
  assign f_arrdiv32_fs572_not0 = ~f_arrdiv32_mux2to1523_xor0;
  assign f_arrdiv32_fs572_and0 = f_arrdiv32_fs572_not0 & b[28];
  assign f_arrdiv32_fs572_xor1 = f_arrdiv32_fs571_or0 ^ f_arrdiv32_fs572_xor0;
  assign f_arrdiv32_fs572_not1 = ~f_arrdiv32_fs572_xor0;
  assign f_arrdiv32_fs572_and1 = f_arrdiv32_fs572_not1 & f_arrdiv32_fs571_or0;
  assign f_arrdiv32_fs572_or0 = f_arrdiv32_fs572_and1 | f_arrdiv32_fs572_and0;
  assign f_arrdiv32_fs573_xor0 = f_arrdiv32_mux2to1524_xor0 ^ b[29];
  assign f_arrdiv32_fs573_not0 = ~f_arrdiv32_mux2to1524_xor0;
  assign f_arrdiv32_fs573_and0 = f_arrdiv32_fs573_not0 & b[29];
  assign f_arrdiv32_fs573_xor1 = f_arrdiv32_fs572_or0 ^ f_arrdiv32_fs573_xor0;
  assign f_arrdiv32_fs573_not1 = ~f_arrdiv32_fs573_xor0;
  assign f_arrdiv32_fs573_and1 = f_arrdiv32_fs573_not1 & f_arrdiv32_fs572_or0;
  assign f_arrdiv32_fs573_or0 = f_arrdiv32_fs573_and1 | f_arrdiv32_fs573_and0;
  assign f_arrdiv32_fs574_xor0 = f_arrdiv32_mux2to1525_xor0 ^ b[30];
  assign f_arrdiv32_fs574_not0 = ~f_arrdiv32_mux2to1525_xor0;
  assign f_arrdiv32_fs574_and0 = f_arrdiv32_fs574_not0 & b[30];
  assign f_arrdiv32_fs574_xor1 = f_arrdiv32_fs573_or0 ^ f_arrdiv32_fs574_xor0;
  assign f_arrdiv32_fs574_not1 = ~f_arrdiv32_fs574_xor0;
  assign f_arrdiv32_fs574_and1 = f_arrdiv32_fs574_not1 & f_arrdiv32_fs573_or0;
  assign f_arrdiv32_fs574_or0 = f_arrdiv32_fs574_and1 | f_arrdiv32_fs574_and0;
  assign f_arrdiv32_fs575_xor0 = f_arrdiv32_mux2to1526_xor0 ^ b[31];
  assign f_arrdiv32_fs575_not0 = ~f_arrdiv32_mux2to1526_xor0;
  assign f_arrdiv32_fs575_and0 = f_arrdiv32_fs575_not0 & b[31];
  assign f_arrdiv32_fs575_xor1 = f_arrdiv32_fs574_or0 ^ f_arrdiv32_fs575_xor0;
  assign f_arrdiv32_fs575_not1 = ~f_arrdiv32_fs575_xor0;
  assign f_arrdiv32_fs575_and1 = f_arrdiv32_fs575_not1 & f_arrdiv32_fs574_or0;
  assign f_arrdiv32_fs575_or0 = f_arrdiv32_fs575_and1 | f_arrdiv32_fs575_and0;
  assign f_arrdiv32_mux2to1527_and0 = a[14] & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1527_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1527_and1 = f_arrdiv32_fs544_xor0 & f_arrdiv32_mux2to1527_not0;
  assign f_arrdiv32_mux2to1527_xor0 = f_arrdiv32_mux2to1527_and0 ^ f_arrdiv32_mux2to1527_and1;
  assign f_arrdiv32_mux2to1528_and0 = f_arrdiv32_mux2to1496_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1528_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1528_and1 = f_arrdiv32_fs545_xor1 & f_arrdiv32_mux2to1528_not0;
  assign f_arrdiv32_mux2to1528_xor0 = f_arrdiv32_mux2to1528_and0 ^ f_arrdiv32_mux2to1528_and1;
  assign f_arrdiv32_mux2to1529_and0 = f_arrdiv32_mux2to1497_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1529_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1529_and1 = f_arrdiv32_fs546_xor1 & f_arrdiv32_mux2to1529_not0;
  assign f_arrdiv32_mux2to1529_xor0 = f_arrdiv32_mux2to1529_and0 ^ f_arrdiv32_mux2to1529_and1;
  assign f_arrdiv32_mux2to1530_and0 = f_arrdiv32_mux2to1498_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1530_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1530_and1 = f_arrdiv32_fs547_xor1 & f_arrdiv32_mux2to1530_not0;
  assign f_arrdiv32_mux2to1530_xor0 = f_arrdiv32_mux2to1530_and0 ^ f_arrdiv32_mux2to1530_and1;
  assign f_arrdiv32_mux2to1531_and0 = f_arrdiv32_mux2to1499_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1531_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1531_and1 = f_arrdiv32_fs548_xor1 & f_arrdiv32_mux2to1531_not0;
  assign f_arrdiv32_mux2to1531_xor0 = f_arrdiv32_mux2to1531_and0 ^ f_arrdiv32_mux2to1531_and1;
  assign f_arrdiv32_mux2to1532_and0 = f_arrdiv32_mux2to1500_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1532_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1532_and1 = f_arrdiv32_fs549_xor1 & f_arrdiv32_mux2to1532_not0;
  assign f_arrdiv32_mux2to1532_xor0 = f_arrdiv32_mux2to1532_and0 ^ f_arrdiv32_mux2to1532_and1;
  assign f_arrdiv32_mux2to1533_and0 = f_arrdiv32_mux2to1501_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1533_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1533_and1 = f_arrdiv32_fs550_xor1 & f_arrdiv32_mux2to1533_not0;
  assign f_arrdiv32_mux2to1533_xor0 = f_arrdiv32_mux2to1533_and0 ^ f_arrdiv32_mux2to1533_and1;
  assign f_arrdiv32_mux2to1534_and0 = f_arrdiv32_mux2to1502_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1534_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1534_and1 = f_arrdiv32_fs551_xor1 & f_arrdiv32_mux2to1534_not0;
  assign f_arrdiv32_mux2to1534_xor0 = f_arrdiv32_mux2to1534_and0 ^ f_arrdiv32_mux2to1534_and1;
  assign f_arrdiv32_mux2to1535_and0 = f_arrdiv32_mux2to1503_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1535_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1535_and1 = f_arrdiv32_fs552_xor1 & f_arrdiv32_mux2to1535_not0;
  assign f_arrdiv32_mux2to1535_xor0 = f_arrdiv32_mux2to1535_and0 ^ f_arrdiv32_mux2to1535_and1;
  assign f_arrdiv32_mux2to1536_and0 = f_arrdiv32_mux2to1504_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1536_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1536_and1 = f_arrdiv32_fs553_xor1 & f_arrdiv32_mux2to1536_not0;
  assign f_arrdiv32_mux2to1536_xor0 = f_arrdiv32_mux2to1536_and0 ^ f_arrdiv32_mux2to1536_and1;
  assign f_arrdiv32_mux2to1537_and0 = f_arrdiv32_mux2to1505_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1537_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1537_and1 = f_arrdiv32_fs554_xor1 & f_arrdiv32_mux2to1537_not0;
  assign f_arrdiv32_mux2to1537_xor0 = f_arrdiv32_mux2to1537_and0 ^ f_arrdiv32_mux2to1537_and1;
  assign f_arrdiv32_mux2to1538_and0 = f_arrdiv32_mux2to1506_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1538_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1538_and1 = f_arrdiv32_fs555_xor1 & f_arrdiv32_mux2to1538_not0;
  assign f_arrdiv32_mux2to1538_xor0 = f_arrdiv32_mux2to1538_and0 ^ f_arrdiv32_mux2to1538_and1;
  assign f_arrdiv32_mux2to1539_and0 = f_arrdiv32_mux2to1507_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1539_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1539_and1 = f_arrdiv32_fs556_xor1 & f_arrdiv32_mux2to1539_not0;
  assign f_arrdiv32_mux2to1539_xor0 = f_arrdiv32_mux2to1539_and0 ^ f_arrdiv32_mux2to1539_and1;
  assign f_arrdiv32_mux2to1540_and0 = f_arrdiv32_mux2to1508_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1540_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1540_and1 = f_arrdiv32_fs557_xor1 & f_arrdiv32_mux2to1540_not0;
  assign f_arrdiv32_mux2to1540_xor0 = f_arrdiv32_mux2to1540_and0 ^ f_arrdiv32_mux2to1540_and1;
  assign f_arrdiv32_mux2to1541_and0 = f_arrdiv32_mux2to1509_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1541_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1541_and1 = f_arrdiv32_fs558_xor1 & f_arrdiv32_mux2to1541_not0;
  assign f_arrdiv32_mux2to1541_xor0 = f_arrdiv32_mux2to1541_and0 ^ f_arrdiv32_mux2to1541_and1;
  assign f_arrdiv32_mux2to1542_and0 = f_arrdiv32_mux2to1510_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1542_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1542_and1 = f_arrdiv32_fs559_xor1 & f_arrdiv32_mux2to1542_not0;
  assign f_arrdiv32_mux2to1542_xor0 = f_arrdiv32_mux2to1542_and0 ^ f_arrdiv32_mux2to1542_and1;
  assign f_arrdiv32_mux2to1543_and0 = f_arrdiv32_mux2to1511_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1543_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1543_and1 = f_arrdiv32_fs560_xor1 & f_arrdiv32_mux2to1543_not0;
  assign f_arrdiv32_mux2to1543_xor0 = f_arrdiv32_mux2to1543_and0 ^ f_arrdiv32_mux2to1543_and1;
  assign f_arrdiv32_mux2to1544_and0 = f_arrdiv32_mux2to1512_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1544_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1544_and1 = f_arrdiv32_fs561_xor1 & f_arrdiv32_mux2to1544_not0;
  assign f_arrdiv32_mux2to1544_xor0 = f_arrdiv32_mux2to1544_and0 ^ f_arrdiv32_mux2to1544_and1;
  assign f_arrdiv32_mux2to1545_and0 = f_arrdiv32_mux2to1513_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1545_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1545_and1 = f_arrdiv32_fs562_xor1 & f_arrdiv32_mux2to1545_not0;
  assign f_arrdiv32_mux2to1545_xor0 = f_arrdiv32_mux2to1545_and0 ^ f_arrdiv32_mux2to1545_and1;
  assign f_arrdiv32_mux2to1546_and0 = f_arrdiv32_mux2to1514_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1546_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1546_and1 = f_arrdiv32_fs563_xor1 & f_arrdiv32_mux2to1546_not0;
  assign f_arrdiv32_mux2to1546_xor0 = f_arrdiv32_mux2to1546_and0 ^ f_arrdiv32_mux2to1546_and1;
  assign f_arrdiv32_mux2to1547_and0 = f_arrdiv32_mux2to1515_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1547_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1547_and1 = f_arrdiv32_fs564_xor1 & f_arrdiv32_mux2to1547_not0;
  assign f_arrdiv32_mux2to1547_xor0 = f_arrdiv32_mux2to1547_and0 ^ f_arrdiv32_mux2to1547_and1;
  assign f_arrdiv32_mux2to1548_and0 = f_arrdiv32_mux2to1516_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1548_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1548_and1 = f_arrdiv32_fs565_xor1 & f_arrdiv32_mux2to1548_not0;
  assign f_arrdiv32_mux2to1548_xor0 = f_arrdiv32_mux2to1548_and0 ^ f_arrdiv32_mux2to1548_and1;
  assign f_arrdiv32_mux2to1549_and0 = f_arrdiv32_mux2to1517_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1549_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1549_and1 = f_arrdiv32_fs566_xor1 & f_arrdiv32_mux2to1549_not0;
  assign f_arrdiv32_mux2to1549_xor0 = f_arrdiv32_mux2to1549_and0 ^ f_arrdiv32_mux2to1549_and1;
  assign f_arrdiv32_mux2to1550_and0 = f_arrdiv32_mux2to1518_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1550_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1550_and1 = f_arrdiv32_fs567_xor1 & f_arrdiv32_mux2to1550_not0;
  assign f_arrdiv32_mux2to1550_xor0 = f_arrdiv32_mux2to1550_and0 ^ f_arrdiv32_mux2to1550_and1;
  assign f_arrdiv32_mux2to1551_and0 = f_arrdiv32_mux2to1519_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1551_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1551_and1 = f_arrdiv32_fs568_xor1 & f_arrdiv32_mux2to1551_not0;
  assign f_arrdiv32_mux2to1551_xor0 = f_arrdiv32_mux2to1551_and0 ^ f_arrdiv32_mux2to1551_and1;
  assign f_arrdiv32_mux2to1552_and0 = f_arrdiv32_mux2to1520_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1552_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1552_and1 = f_arrdiv32_fs569_xor1 & f_arrdiv32_mux2to1552_not0;
  assign f_arrdiv32_mux2to1552_xor0 = f_arrdiv32_mux2to1552_and0 ^ f_arrdiv32_mux2to1552_and1;
  assign f_arrdiv32_mux2to1553_and0 = f_arrdiv32_mux2to1521_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1553_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1553_and1 = f_arrdiv32_fs570_xor1 & f_arrdiv32_mux2to1553_not0;
  assign f_arrdiv32_mux2to1553_xor0 = f_arrdiv32_mux2to1553_and0 ^ f_arrdiv32_mux2to1553_and1;
  assign f_arrdiv32_mux2to1554_and0 = f_arrdiv32_mux2to1522_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1554_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1554_and1 = f_arrdiv32_fs571_xor1 & f_arrdiv32_mux2to1554_not0;
  assign f_arrdiv32_mux2to1554_xor0 = f_arrdiv32_mux2to1554_and0 ^ f_arrdiv32_mux2to1554_and1;
  assign f_arrdiv32_mux2to1555_and0 = f_arrdiv32_mux2to1523_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1555_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1555_and1 = f_arrdiv32_fs572_xor1 & f_arrdiv32_mux2to1555_not0;
  assign f_arrdiv32_mux2to1555_xor0 = f_arrdiv32_mux2to1555_and0 ^ f_arrdiv32_mux2to1555_and1;
  assign f_arrdiv32_mux2to1556_and0 = f_arrdiv32_mux2to1524_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1556_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1556_and1 = f_arrdiv32_fs573_xor1 & f_arrdiv32_mux2to1556_not0;
  assign f_arrdiv32_mux2to1556_xor0 = f_arrdiv32_mux2to1556_and0 ^ f_arrdiv32_mux2to1556_and1;
  assign f_arrdiv32_mux2to1557_and0 = f_arrdiv32_mux2to1525_xor0 & f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1557_not0 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_mux2to1557_and1 = f_arrdiv32_fs574_xor1 & f_arrdiv32_mux2to1557_not0;
  assign f_arrdiv32_mux2to1557_xor0 = f_arrdiv32_mux2to1557_and0 ^ f_arrdiv32_mux2to1557_and1;
  assign f_arrdiv32_not17 = ~f_arrdiv32_fs575_or0;
  assign f_arrdiv32_fs576_xor0 = a[13] ^ b[0];
  assign f_arrdiv32_fs576_not0 = ~a[13];
  assign f_arrdiv32_fs576_and0 = f_arrdiv32_fs576_not0 & b[0];
  assign f_arrdiv32_fs576_not1 = ~f_arrdiv32_fs576_xor0;
  assign f_arrdiv32_fs577_xor0 = f_arrdiv32_mux2to1527_xor0 ^ b[1];
  assign f_arrdiv32_fs577_not0 = ~f_arrdiv32_mux2to1527_xor0;
  assign f_arrdiv32_fs577_and0 = f_arrdiv32_fs577_not0 & b[1];
  assign f_arrdiv32_fs577_xor1 = f_arrdiv32_fs576_and0 ^ f_arrdiv32_fs577_xor0;
  assign f_arrdiv32_fs577_not1 = ~f_arrdiv32_fs577_xor0;
  assign f_arrdiv32_fs577_and1 = f_arrdiv32_fs577_not1 & f_arrdiv32_fs576_and0;
  assign f_arrdiv32_fs577_or0 = f_arrdiv32_fs577_and1 | f_arrdiv32_fs577_and0;
  assign f_arrdiv32_fs578_xor0 = f_arrdiv32_mux2to1528_xor0 ^ b[2];
  assign f_arrdiv32_fs578_not0 = ~f_arrdiv32_mux2to1528_xor0;
  assign f_arrdiv32_fs578_and0 = f_arrdiv32_fs578_not0 & b[2];
  assign f_arrdiv32_fs578_xor1 = f_arrdiv32_fs577_or0 ^ f_arrdiv32_fs578_xor0;
  assign f_arrdiv32_fs578_not1 = ~f_arrdiv32_fs578_xor0;
  assign f_arrdiv32_fs578_and1 = f_arrdiv32_fs578_not1 & f_arrdiv32_fs577_or0;
  assign f_arrdiv32_fs578_or0 = f_arrdiv32_fs578_and1 | f_arrdiv32_fs578_and0;
  assign f_arrdiv32_fs579_xor0 = f_arrdiv32_mux2to1529_xor0 ^ b[3];
  assign f_arrdiv32_fs579_not0 = ~f_arrdiv32_mux2to1529_xor0;
  assign f_arrdiv32_fs579_and0 = f_arrdiv32_fs579_not0 & b[3];
  assign f_arrdiv32_fs579_xor1 = f_arrdiv32_fs578_or0 ^ f_arrdiv32_fs579_xor0;
  assign f_arrdiv32_fs579_not1 = ~f_arrdiv32_fs579_xor0;
  assign f_arrdiv32_fs579_and1 = f_arrdiv32_fs579_not1 & f_arrdiv32_fs578_or0;
  assign f_arrdiv32_fs579_or0 = f_arrdiv32_fs579_and1 | f_arrdiv32_fs579_and0;
  assign f_arrdiv32_fs580_xor0 = f_arrdiv32_mux2to1530_xor0 ^ b[4];
  assign f_arrdiv32_fs580_not0 = ~f_arrdiv32_mux2to1530_xor0;
  assign f_arrdiv32_fs580_and0 = f_arrdiv32_fs580_not0 & b[4];
  assign f_arrdiv32_fs580_xor1 = f_arrdiv32_fs579_or0 ^ f_arrdiv32_fs580_xor0;
  assign f_arrdiv32_fs580_not1 = ~f_arrdiv32_fs580_xor0;
  assign f_arrdiv32_fs580_and1 = f_arrdiv32_fs580_not1 & f_arrdiv32_fs579_or0;
  assign f_arrdiv32_fs580_or0 = f_arrdiv32_fs580_and1 | f_arrdiv32_fs580_and0;
  assign f_arrdiv32_fs581_xor0 = f_arrdiv32_mux2to1531_xor0 ^ b[5];
  assign f_arrdiv32_fs581_not0 = ~f_arrdiv32_mux2to1531_xor0;
  assign f_arrdiv32_fs581_and0 = f_arrdiv32_fs581_not0 & b[5];
  assign f_arrdiv32_fs581_xor1 = f_arrdiv32_fs580_or0 ^ f_arrdiv32_fs581_xor0;
  assign f_arrdiv32_fs581_not1 = ~f_arrdiv32_fs581_xor0;
  assign f_arrdiv32_fs581_and1 = f_arrdiv32_fs581_not1 & f_arrdiv32_fs580_or0;
  assign f_arrdiv32_fs581_or0 = f_arrdiv32_fs581_and1 | f_arrdiv32_fs581_and0;
  assign f_arrdiv32_fs582_xor0 = f_arrdiv32_mux2to1532_xor0 ^ b[6];
  assign f_arrdiv32_fs582_not0 = ~f_arrdiv32_mux2to1532_xor0;
  assign f_arrdiv32_fs582_and0 = f_arrdiv32_fs582_not0 & b[6];
  assign f_arrdiv32_fs582_xor1 = f_arrdiv32_fs581_or0 ^ f_arrdiv32_fs582_xor0;
  assign f_arrdiv32_fs582_not1 = ~f_arrdiv32_fs582_xor0;
  assign f_arrdiv32_fs582_and1 = f_arrdiv32_fs582_not1 & f_arrdiv32_fs581_or0;
  assign f_arrdiv32_fs582_or0 = f_arrdiv32_fs582_and1 | f_arrdiv32_fs582_and0;
  assign f_arrdiv32_fs583_xor0 = f_arrdiv32_mux2to1533_xor0 ^ b[7];
  assign f_arrdiv32_fs583_not0 = ~f_arrdiv32_mux2to1533_xor0;
  assign f_arrdiv32_fs583_and0 = f_arrdiv32_fs583_not0 & b[7];
  assign f_arrdiv32_fs583_xor1 = f_arrdiv32_fs582_or0 ^ f_arrdiv32_fs583_xor0;
  assign f_arrdiv32_fs583_not1 = ~f_arrdiv32_fs583_xor0;
  assign f_arrdiv32_fs583_and1 = f_arrdiv32_fs583_not1 & f_arrdiv32_fs582_or0;
  assign f_arrdiv32_fs583_or0 = f_arrdiv32_fs583_and1 | f_arrdiv32_fs583_and0;
  assign f_arrdiv32_fs584_xor0 = f_arrdiv32_mux2to1534_xor0 ^ b[8];
  assign f_arrdiv32_fs584_not0 = ~f_arrdiv32_mux2to1534_xor0;
  assign f_arrdiv32_fs584_and0 = f_arrdiv32_fs584_not0 & b[8];
  assign f_arrdiv32_fs584_xor1 = f_arrdiv32_fs583_or0 ^ f_arrdiv32_fs584_xor0;
  assign f_arrdiv32_fs584_not1 = ~f_arrdiv32_fs584_xor0;
  assign f_arrdiv32_fs584_and1 = f_arrdiv32_fs584_not1 & f_arrdiv32_fs583_or0;
  assign f_arrdiv32_fs584_or0 = f_arrdiv32_fs584_and1 | f_arrdiv32_fs584_and0;
  assign f_arrdiv32_fs585_xor0 = f_arrdiv32_mux2to1535_xor0 ^ b[9];
  assign f_arrdiv32_fs585_not0 = ~f_arrdiv32_mux2to1535_xor0;
  assign f_arrdiv32_fs585_and0 = f_arrdiv32_fs585_not0 & b[9];
  assign f_arrdiv32_fs585_xor1 = f_arrdiv32_fs584_or0 ^ f_arrdiv32_fs585_xor0;
  assign f_arrdiv32_fs585_not1 = ~f_arrdiv32_fs585_xor0;
  assign f_arrdiv32_fs585_and1 = f_arrdiv32_fs585_not1 & f_arrdiv32_fs584_or0;
  assign f_arrdiv32_fs585_or0 = f_arrdiv32_fs585_and1 | f_arrdiv32_fs585_and0;
  assign f_arrdiv32_fs586_xor0 = f_arrdiv32_mux2to1536_xor0 ^ b[10];
  assign f_arrdiv32_fs586_not0 = ~f_arrdiv32_mux2to1536_xor0;
  assign f_arrdiv32_fs586_and0 = f_arrdiv32_fs586_not0 & b[10];
  assign f_arrdiv32_fs586_xor1 = f_arrdiv32_fs585_or0 ^ f_arrdiv32_fs586_xor0;
  assign f_arrdiv32_fs586_not1 = ~f_arrdiv32_fs586_xor0;
  assign f_arrdiv32_fs586_and1 = f_arrdiv32_fs586_not1 & f_arrdiv32_fs585_or0;
  assign f_arrdiv32_fs586_or0 = f_arrdiv32_fs586_and1 | f_arrdiv32_fs586_and0;
  assign f_arrdiv32_fs587_xor0 = f_arrdiv32_mux2to1537_xor0 ^ b[11];
  assign f_arrdiv32_fs587_not0 = ~f_arrdiv32_mux2to1537_xor0;
  assign f_arrdiv32_fs587_and0 = f_arrdiv32_fs587_not0 & b[11];
  assign f_arrdiv32_fs587_xor1 = f_arrdiv32_fs586_or0 ^ f_arrdiv32_fs587_xor0;
  assign f_arrdiv32_fs587_not1 = ~f_arrdiv32_fs587_xor0;
  assign f_arrdiv32_fs587_and1 = f_arrdiv32_fs587_not1 & f_arrdiv32_fs586_or0;
  assign f_arrdiv32_fs587_or0 = f_arrdiv32_fs587_and1 | f_arrdiv32_fs587_and0;
  assign f_arrdiv32_fs588_xor0 = f_arrdiv32_mux2to1538_xor0 ^ b[12];
  assign f_arrdiv32_fs588_not0 = ~f_arrdiv32_mux2to1538_xor0;
  assign f_arrdiv32_fs588_and0 = f_arrdiv32_fs588_not0 & b[12];
  assign f_arrdiv32_fs588_xor1 = f_arrdiv32_fs587_or0 ^ f_arrdiv32_fs588_xor0;
  assign f_arrdiv32_fs588_not1 = ~f_arrdiv32_fs588_xor0;
  assign f_arrdiv32_fs588_and1 = f_arrdiv32_fs588_not1 & f_arrdiv32_fs587_or0;
  assign f_arrdiv32_fs588_or0 = f_arrdiv32_fs588_and1 | f_arrdiv32_fs588_and0;
  assign f_arrdiv32_fs589_xor0 = f_arrdiv32_mux2to1539_xor0 ^ b[13];
  assign f_arrdiv32_fs589_not0 = ~f_arrdiv32_mux2to1539_xor0;
  assign f_arrdiv32_fs589_and0 = f_arrdiv32_fs589_not0 & b[13];
  assign f_arrdiv32_fs589_xor1 = f_arrdiv32_fs588_or0 ^ f_arrdiv32_fs589_xor0;
  assign f_arrdiv32_fs589_not1 = ~f_arrdiv32_fs589_xor0;
  assign f_arrdiv32_fs589_and1 = f_arrdiv32_fs589_not1 & f_arrdiv32_fs588_or0;
  assign f_arrdiv32_fs589_or0 = f_arrdiv32_fs589_and1 | f_arrdiv32_fs589_and0;
  assign f_arrdiv32_fs590_xor0 = f_arrdiv32_mux2to1540_xor0 ^ b[14];
  assign f_arrdiv32_fs590_not0 = ~f_arrdiv32_mux2to1540_xor0;
  assign f_arrdiv32_fs590_and0 = f_arrdiv32_fs590_not0 & b[14];
  assign f_arrdiv32_fs590_xor1 = f_arrdiv32_fs589_or0 ^ f_arrdiv32_fs590_xor0;
  assign f_arrdiv32_fs590_not1 = ~f_arrdiv32_fs590_xor0;
  assign f_arrdiv32_fs590_and1 = f_arrdiv32_fs590_not1 & f_arrdiv32_fs589_or0;
  assign f_arrdiv32_fs590_or0 = f_arrdiv32_fs590_and1 | f_arrdiv32_fs590_and0;
  assign f_arrdiv32_fs591_xor0 = f_arrdiv32_mux2to1541_xor0 ^ b[15];
  assign f_arrdiv32_fs591_not0 = ~f_arrdiv32_mux2to1541_xor0;
  assign f_arrdiv32_fs591_and0 = f_arrdiv32_fs591_not0 & b[15];
  assign f_arrdiv32_fs591_xor1 = f_arrdiv32_fs590_or0 ^ f_arrdiv32_fs591_xor0;
  assign f_arrdiv32_fs591_not1 = ~f_arrdiv32_fs591_xor0;
  assign f_arrdiv32_fs591_and1 = f_arrdiv32_fs591_not1 & f_arrdiv32_fs590_or0;
  assign f_arrdiv32_fs591_or0 = f_arrdiv32_fs591_and1 | f_arrdiv32_fs591_and0;
  assign f_arrdiv32_fs592_xor0 = f_arrdiv32_mux2to1542_xor0 ^ b[16];
  assign f_arrdiv32_fs592_not0 = ~f_arrdiv32_mux2to1542_xor0;
  assign f_arrdiv32_fs592_and0 = f_arrdiv32_fs592_not0 & b[16];
  assign f_arrdiv32_fs592_xor1 = f_arrdiv32_fs591_or0 ^ f_arrdiv32_fs592_xor0;
  assign f_arrdiv32_fs592_not1 = ~f_arrdiv32_fs592_xor0;
  assign f_arrdiv32_fs592_and1 = f_arrdiv32_fs592_not1 & f_arrdiv32_fs591_or0;
  assign f_arrdiv32_fs592_or0 = f_arrdiv32_fs592_and1 | f_arrdiv32_fs592_and0;
  assign f_arrdiv32_fs593_xor0 = f_arrdiv32_mux2to1543_xor0 ^ b[17];
  assign f_arrdiv32_fs593_not0 = ~f_arrdiv32_mux2to1543_xor0;
  assign f_arrdiv32_fs593_and0 = f_arrdiv32_fs593_not0 & b[17];
  assign f_arrdiv32_fs593_xor1 = f_arrdiv32_fs592_or0 ^ f_arrdiv32_fs593_xor0;
  assign f_arrdiv32_fs593_not1 = ~f_arrdiv32_fs593_xor0;
  assign f_arrdiv32_fs593_and1 = f_arrdiv32_fs593_not1 & f_arrdiv32_fs592_or0;
  assign f_arrdiv32_fs593_or0 = f_arrdiv32_fs593_and1 | f_arrdiv32_fs593_and0;
  assign f_arrdiv32_fs594_xor0 = f_arrdiv32_mux2to1544_xor0 ^ b[18];
  assign f_arrdiv32_fs594_not0 = ~f_arrdiv32_mux2to1544_xor0;
  assign f_arrdiv32_fs594_and0 = f_arrdiv32_fs594_not0 & b[18];
  assign f_arrdiv32_fs594_xor1 = f_arrdiv32_fs593_or0 ^ f_arrdiv32_fs594_xor0;
  assign f_arrdiv32_fs594_not1 = ~f_arrdiv32_fs594_xor0;
  assign f_arrdiv32_fs594_and1 = f_arrdiv32_fs594_not1 & f_arrdiv32_fs593_or0;
  assign f_arrdiv32_fs594_or0 = f_arrdiv32_fs594_and1 | f_arrdiv32_fs594_and0;
  assign f_arrdiv32_fs595_xor0 = f_arrdiv32_mux2to1545_xor0 ^ b[19];
  assign f_arrdiv32_fs595_not0 = ~f_arrdiv32_mux2to1545_xor0;
  assign f_arrdiv32_fs595_and0 = f_arrdiv32_fs595_not0 & b[19];
  assign f_arrdiv32_fs595_xor1 = f_arrdiv32_fs594_or0 ^ f_arrdiv32_fs595_xor0;
  assign f_arrdiv32_fs595_not1 = ~f_arrdiv32_fs595_xor0;
  assign f_arrdiv32_fs595_and1 = f_arrdiv32_fs595_not1 & f_arrdiv32_fs594_or0;
  assign f_arrdiv32_fs595_or0 = f_arrdiv32_fs595_and1 | f_arrdiv32_fs595_and0;
  assign f_arrdiv32_fs596_xor0 = f_arrdiv32_mux2to1546_xor0 ^ b[20];
  assign f_arrdiv32_fs596_not0 = ~f_arrdiv32_mux2to1546_xor0;
  assign f_arrdiv32_fs596_and0 = f_arrdiv32_fs596_not0 & b[20];
  assign f_arrdiv32_fs596_xor1 = f_arrdiv32_fs595_or0 ^ f_arrdiv32_fs596_xor0;
  assign f_arrdiv32_fs596_not1 = ~f_arrdiv32_fs596_xor0;
  assign f_arrdiv32_fs596_and1 = f_arrdiv32_fs596_not1 & f_arrdiv32_fs595_or0;
  assign f_arrdiv32_fs596_or0 = f_arrdiv32_fs596_and1 | f_arrdiv32_fs596_and0;
  assign f_arrdiv32_fs597_xor0 = f_arrdiv32_mux2to1547_xor0 ^ b[21];
  assign f_arrdiv32_fs597_not0 = ~f_arrdiv32_mux2to1547_xor0;
  assign f_arrdiv32_fs597_and0 = f_arrdiv32_fs597_not0 & b[21];
  assign f_arrdiv32_fs597_xor1 = f_arrdiv32_fs596_or0 ^ f_arrdiv32_fs597_xor0;
  assign f_arrdiv32_fs597_not1 = ~f_arrdiv32_fs597_xor0;
  assign f_arrdiv32_fs597_and1 = f_arrdiv32_fs597_not1 & f_arrdiv32_fs596_or0;
  assign f_arrdiv32_fs597_or0 = f_arrdiv32_fs597_and1 | f_arrdiv32_fs597_and0;
  assign f_arrdiv32_fs598_xor0 = f_arrdiv32_mux2to1548_xor0 ^ b[22];
  assign f_arrdiv32_fs598_not0 = ~f_arrdiv32_mux2to1548_xor0;
  assign f_arrdiv32_fs598_and0 = f_arrdiv32_fs598_not0 & b[22];
  assign f_arrdiv32_fs598_xor1 = f_arrdiv32_fs597_or0 ^ f_arrdiv32_fs598_xor0;
  assign f_arrdiv32_fs598_not1 = ~f_arrdiv32_fs598_xor0;
  assign f_arrdiv32_fs598_and1 = f_arrdiv32_fs598_not1 & f_arrdiv32_fs597_or0;
  assign f_arrdiv32_fs598_or0 = f_arrdiv32_fs598_and1 | f_arrdiv32_fs598_and0;
  assign f_arrdiv32_fs599_xor0 = f_arrdiv32_mux2to1549_xor0 ^ b[23];
  assign f_arrdiv32_fs599_not0 = ~f_arrdiv32_mux2to1549_xor0;
  assign f_arrdiv32_fs599_and0 = f_arrdiv32_fs599_not0 & b[23];
  assign f_arrdiv32_fs599_xor1 = f_arrdiv32_fs598_or0 ^ f_arrdiv32_fs599_xor0;
  assign f_arrdiv32_fs599_not1 = ~f_arrdiv32_fs599_xor0;
  assign f_arrdiv32_fs599_and1 = f_arrdiv32_fs599_not1 & f_arrdiv32_fs598_or0;
  assign f_arrdiv32_fs599_or0 = f_arrdiv32_fs599_and1 | f_arrdiv32_fs599_and0;
  assign f_arrdiv32_fs600_xor0 = f_arrdiv32_mux2to1550_xor0 ^ b[24];
  assign f_arrdiv32_fs600_not0 = ~f_arrdiv32_mux2to1550_xor0;
  assign f_arrdiv32_fs600_and0 = f_arrdiv32_fs600_not0 & b[24];
  assign f_arrdiv32_fs600_xor1 = f_arrdiv32_fs599_or0 ^ f_arrdiv32_fs600_xor0;
  assign f_arrdiv32_fs600_not1 = ~f_arrdiv32_fs600_xor0;
  assign f_arrdiv32_fs600_and1 = f_arrdiv32_fs600_not1 & f_arrdiv32_fs599_or0;
  assign f_arrdiv32_fs600_or0 = f_arrdiv32_fs600_and1 | f_arrdiv32_fs600_and0;
  assign f_arrdiv32_fs601_xor0 = f_arrdiv32_mux2to1551_xor0 ^ b[25];
  assign f_arrdiv32_fs601_not0 = ~f_arrdiv32_mux2to1551_xor0;
  assign f_arrdiv32_fs601_and0 = f_arrdiv32_fs601_not0 & b[25];
  assign f_arrdiv32_fs601_xor1 = f_arrdiv32_fs600_or0 ^ f_arrdiv32_fs601_xor0;
  assign f_arrdiv32_fs601_not1 = ~f_arrdiv32_fs601_xor0;
  assign f_arrdiv32_fs601_and1 = f_arrdiv32_fs601_not1 & f_arrdiv32_fs600_or0;
  assign f_arrdiv32_fs601_or0 = f_arrdiv32_fs601_and1 | f_arrdiv32_fs601_and0;
  assign f_arrdiv32_fs602_xor0 = f_arrdiv32_mux2to1552_xor0 ^ b[26];
  assign f_arrdiv32_fs602_not0 = ~f_arrdiv32_mux2to1552_xor0;
  assign f_arrdiv32_fs602_and0 = f_arrdiv32_fs602_not0 & b[26];
  assign f_arrdiv32_fs602_xor1 = f_arrdiv32_fs601_or0 ^ f_arrdiv32_fs602_xor0;
  assign f_arrdiv32_fs602_not1 = ~f_arrdiv32_fs602_xor0;
  assign f_arrdiv32_fs602_and1 = f_arrdiv32_fs602_not1 & f_arrdiv32_fs601_or0;
  assign f_arrdiv32_fs602_or0 = f_arrdiv32_fs602_and1 | f_arrdiv32_fs602_and0;
  assign f_arrdiv32_fs603_xor0 = f_arrdiv32_mux2to1553_xor0 ^ b[27];
  assign f_arrdiv32_fs603_not0 = ~f_arrdiv32_mux2to1553_xor0;
  assign f_arrdiv32_fs603_and0 = f_arrdiv32_fs603_not0 & b[27];
  assign f_arrdiv32_fs603_xor1 = f_arrdiv32_fs602_or0 ^ f_arrdiv32_fs603_xor0;
  assign f_arrdiv32_fs603_not1 = ~f_arrdiv32_fs603_xor0;
  assign f_arrdiv32_fs603_and1 = f_arrdiv32_fs603_not1 & f_arrdiv32_fs602_or0;
  assign f_arrdiv32_fs603_or0 = f_arrdiv32_fs603_and1 | f_arrdiv32_fs603_and0;
  assign f_arrdiv32_fs604_xor0 = f_arrdiv32_mux2to1554_xor0 ^ b[28];
  assign f_arrdiv32_fs604_not0 = ~f_arrdiv32_mux2to1554_xor0;
  assign f_arrdiv32_fs604_and0 = f_arrdiv32_fs604_not0 & b[28];
  assign f_arrdiv32_fs604_xor1 = f_arrdiv32_fs603_or0 ^ f_arrdiv32_fs604_xor0;
  assign f_arrdiv32_fs604_not1 = ~f_arrdiv32_fs604_xor0;
  assign f_arrdiv32_fs604_and1 = f_arrdiv32_fs604_not1 & f_arrdiv32_fs603_or0;
  assign f_arrdiv32_fs604_or0 = f_arrdiv32_fs604_and1 | f_arrdiv32_fs604_and0;
  assign f_arrdiv32_fs605_xor0 = f_arrdiv32_mux2to1555_xor0 ^ b[29];
  assign f_arrdiv32_fs605_not0 = ~f_arrdiv32_mux2to1555_xor0;
  assign f_arrdiv32_fs605_and0 = f_arrdiv32_fs605_not0 & b[29];
  assign f_arrdiv32_fs605_xor1 = f_arrdiv32_fs604_or0 ^ f_arrdiv32_fs605_xor0;
  assign f_arrdiv32_fs605_not1 = ~f_arrdiv32_fs605_xor0;
  assign f_arrdiv32_fs605_and1 = f_arrdiv32_fs605_not1 & f_arrdiv32_fs604_or0;
  assign f_arrdiv32_fs605_or0 = f_arrdiv32_fs605_and1 | f_arrdiv32_fs605_and0;
  assign f_arrdiv32_fs606_xor0 = f_arrdiv32_mux2to1556_xor0 ^ b[30];
  assign f_arrdiv32_fs606_not0 = ~f_arrdiv32_mux2to1556_xor0;
  assign f_arrdiv32_fs606_and0 = f_arrdiv32_fs606_not0 & b[30];
  assign f_arrdiv32_fs606_xor1 = f_arrdiv32_fs605_or0 ^ f_arrdiv32_fs606_xor0;
  assign f_arrdiv32_fs606_not1 = ~f_arrdiv32_fs606_xor0;
  assign f_arrdiv32_fs606_and1 = f_arrdiv32_fs606_not1 & f_arrdiv32_fs605_or0;
  assign f_arrdiv32_fs606_or0 = f_arrdiv32_fs606_and1 | f_arrdiv32_fs606_and0;
  assign f_arrdiv32_fs607_xor0 = f_arrdiv32_mux2to1557_xor0 ^ b[31];
  assign f_arrdiv32_fs607_not0 = ~f_arrdiv32_mux2to1557_xor0;
  assign f_arrdiv32_fs607_and0 = f_arrdiv32_fs607_not0 & b[31];
  assign f_arrdiv32_fs607_xor1 = f_arrdiv32_fs606_or0 ^ f_arrdiv32_fs607_xor0;
  assign f_arrdiv32_fs607_not1 = ~f_arrdiv32_fs607_xor0;
  assign f_arrdiv32_fs607_and1 = f_arrdiv32_fs607_not1 & f_arrdiv32_fs606_or0;
  assign f_arrdiv32_fs607_or0 = f_arrdiv32_fs607_and1 | f_arrdiv32_fs607_and0;
  assign f_arrdiv32_mux2to1558_and0 = a[13] & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1558_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1558_and1 = f_arrdiv32_fs576_xor0 & f_arrdiv32_mux2to1558_not0;
  assign f_arrdiv32_mux2to1558_xor0 = f_arrdiv32_mux2to1558_and0 ^ f_arrdiv32_mux2to1558_and1;
  assign f_arrdiv32_mux2to1559_and0 = f_arrdiv32_mux2to1527_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1559_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1559_and1 = f_arrdiv32_fs577_xor1 & f_arrdiv32_mux2to1559_not0;
  assign f_arrdiv32_mux2to1559_xor0 = f_arrdiv32_mux2to1559_and0 ^ f_arrdiv32_mux2to1559_and1;
  assign f_arrdiv32_mux2to1560_and0 = f_arrdiv32_mux2to1528_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1560_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1560_and1 = f_arrdiv32_fs578_xor1 & f_arrdiv32_mux2to1560_not0;
  assign f_arrdiv32_mux2to1560_xor0 = f_arrdiv32_mux2to1560_and0 ^ f_arrdiv32_mux2to1560_and1;
  assign f_arrdiv32_mux2to1561_and0 = f_arrdiv32_mux2to1529_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1561_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1561_and1 = f_arrdiv32_fs579_xor1 & f_arrdiv32_mux2to1561_not0;
  assign f_arrdiv32_mux2to1561_xor0 = f_arrdiv32_mux2to1561_and0 ^ f_arrdiv32_mux2to1561_and1;
  assign f_arrdiv32_mux2to1562_and0 = f_arrdiv32_mux2to1530_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1562_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1562_and1 = f_arrdiv32_fs580_xor1 & f_arrdiv32_mux2to1562_not0;
  assign f_arrdiv32_mux2to1562_xor0 = f_arrdiv32_mux2to1562_and0 ^ f_arrdiv32_mux2to1562_and1;
  assign f_arrdiv32_mux2to1563_and0 = f_arrdiv32_mux2to1531_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1563_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1563_and1 = f_arrdiv32_fs581_xor1 & f_arrdiv32_mux2to1563_not0;
  assign f_arrdiv32_mux2to1563_xor0 = f_arrdiv32_mux2to1563_and0 ^ f_arrdiv32_mux2to1563_and1;
  assign f_arrdiv32_mux2to1564_and0 = f_arrdiv32_mux2to1532_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1564_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1564_and1 = f_arrdiv32_fs582_xor1 & f_arrdiv32_mux2to1564_not0;
  assign f_arrdiv32_mux2to1564_xor0 = f_arrdiv32_mux2to1564_and0 ^ f_arrdiv32_mux2to1564_and1;
  assign f_arrdiv32_mux2to1565_and0 = f_arrdiv32_mux2to1533_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1565_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1565_and1 = f_arrdiv32_fs583_xor1 & f_arrdiv32_mux2to1565_not0;
  assign f_arrdiv32_mux2to1565_xor0 = f_arrdiv32_mux2to1565_and0 ^ f_arrdiv32_mux2to1565_and1;
  assign f_arrdiv32_mux2to1566_and0 = f_arrdiv32_mux2to1534_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1566_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1566_and1 = f_arrdiv32_fs584_xor1 & f_arrdiv32_mux2to1566_not0;
  assign f_arrdiv32_mux2to1566_xor0 = f_arrdiv32_mux2to1566_and0 ^ f_arrdiv32_mux2to1566_and1;
  assign f_arrdiv32_mux2to1567_and0 = f_arrdiv32_mux2to1535_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1567_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1567_and1 = f_arrdiv32_fs585_xor1 & f_arrdiv32_mux2to1567_not0;
  assign f_arrdiv32_mux2to1567_xor0 = f_arrdiv32_mux2to1567_and0 ^ f_arrdiv32_mux2to1567_and1;
  assign f_arrdiv32_mux2to1568_and0 = f_arrdiv32_mux2to1536_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1568_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1568_and1 = f_arrdiv32_fs586_xor1 & f_arrdiv32_mux2to1568_not0;
  assign f_arrdiv32_mux2to1568_xor0 = f_arrdiv32_mux2to1568_and0 ^ f_arrdiv32_mux2to1568_and1;
  assign f_arrdiv32_mux2to1569_and0 = f_arrdiv32_mux2to1537_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1569_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1569_and1 = f_arrdiv32_fs587_xor1 & f_arrdiv32_mux2to1569_not0;
  assign f_arrdiv32_mux2to1569_xor0 = f_arrdiv32_mux2to1569_and0 ^ f_arrdiv32_mux2to1569_and1;
  assign f_arrdiv32_mux2to1570_and0 = f_arrdiv32_mux2to1538_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1570_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1570_and1 = f_arrdiv32_fs588_xor1 & f_arrdiv32_mux2to1570_not0;
  assign f_arrdiv32_mux2to1570_xor0 = f_arrdiv32_mux2to1570_and0 ^ f_arrdiv32_mux2to1570_and1;
  assign f_arrdiv32_mux2to1571_and0 = f_arrdiv32_mux2to1539_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1571_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1571_and1 = f_arrdiv32_fs589_xor1 & f_arrdiv32_mux2to1571_not0;
  assign f_arrdiv32_mux2to1571_xor0 = f_arrdiv32_mux2to1571_and0 ^ f_arrdiv32_mux2to1571_and1;
  assign f_arrdiv32_mux2to1572_and0 = f_arrdiv32_mux2to1540_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1572_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1572_and1 = f_arrdiv32_fs590_xor1 & f_arrdiv32_mux2to1572_not0;
  assign f_arrdiv32_mux2to1572_xor0 = f_arrdiv32_mux2to1572_and0 ^ f_arrdiv32_mux2to1572_and1;
  assign f_arrdiv32_mux2to1573_and0 = f_arrdiv32_mux2to1541_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1573_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1573_and1 = f_arrdiv32_fs591_xor1 & f_arrdiv32_mux2to1573_not0;
  assign f_arrdiv32_mux2to1573_xor0 = f_arrdiv32_mux2to1573_and0 ^ f_arrdiv32_mux2to1573_and1;
  assign f_arrdiv32_mux2to1574_and0 = f_arrdiv32_mux2to1542_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1574_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1574_and1 = f_arrdiv32_fs592_xor1 & f_arrdiv32_mux2to1574_not0;
  assign f_arrdiv32_mux2to1574_xor0 = f_arrdiv32_mux2to1574_and0 ^ f_arrdiv32_mux2to1574_and1;
  assign f_arrdiv32_mux2to1575_and0 = f_arrdiv32_mux2to1543_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1575_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1575_and1 = f_arrdiv32_fs593_xor1 & f_arrdiv32_mux2to1575_not0;
  assign f_arrdiv32_mux2to1575_xor0 = f_arrdiv32_mux2to1575_and0 ^ f_arrdiv32_mux2to1575_and1;
  assign f_arrdiv32_mux2to1576_and0 = f_arrdiv32_mux2to1544_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1576_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1576_and1 = f_arrdiv32_fs594_xor1 & f_arrdiv32_mux2to1576_not0;
  assign f_arrdiv32_mux2to1576_xor0 = f_arrdiv32_mux2to1576_and0 ^ f_arrdiv32_mux2to1576_and1;
  assign f_arrdiv32_mux2to1577_and0 = f_arrdiv32_mux2to1545_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1577_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1577_and1 = f_arrdiv32_fs595_xor1 & f_arrdiv32_mux2to1577_not0;
  assign f_arrdiv32_mux2to1577_xor0 = f_arrdiv32_mux2to1577_and0 ^ f_arrdiv32_mux2to1577_and1;
  assign f_arrdiv32_mux2to1578_and0 = f_arrdiv32_mux2to1546_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1578_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1578_and1 = f_arrdiv32_fs596_xor1 & f_arrdiv32_mux2to1578_not0;
  assign f_arrdiv32_mux2to1578_xor0 = f_arrdiv32_mux2to1578_and0 ^ f_arrdiv32_mux2to1578_and1;
  assign f_arrdiv32_mux2to1579_and0 = f_arrdiv32_mux2to1547_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1579_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1579_and1 = f_arrdiv32_fs597_xor1 & f_arrdiv32_mux2to1579_not0;
  assign f_arrdiv32_mux2to1579_xor0 = f_arrdiv32_mux2to1579_and0 ^ f_arrdiv32_mux2to1579_and1;
  assign f_arrdiv32_mux2to1580_and0 = f_arrdiv32_mux2to1548_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1580_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1580_and1 = f_arrdiv32_fs598_xor1 & f_arrdiv32_mux2to1580_not0;
  assign f_arrdiv32_mux2to1580_xor0 = f_arrdiv32_mux2to1580_and0 ^ f_arrdiv32_mux2to1580_and1;
  assign f_arrdiv32_mux2to1581_and0 = f_arrdiv32_mux2to1549_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1581_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1581_and1 = f_arrdiv32_fs599_xor1 & f_arrdiv32_mux2to1581_not0;
  assign f_arrdiv32_mux2to1581_xor0 = f_arrdiv32_mux2to1581_and0 ^ f_arrdiv32_mux2to1581_and1;
  assign f_arrdiv32_mux2to1582_and0 = f_arrdiv32_mux2to1550_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1582_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1582_and1 = f_arrdiv32_fs600_xor1 & f_arrdiv32_mux2to1582_not0;
  assign f_arrdiv32_mux2to1582_xor0 = f_arrdiv32_mux2to1582_and0 ^ f_arrdiv32_mux2to1582_and1;
  assign f_arrdiv32_mux2to1583_and0 = f_arrdiv32_mux2to1551_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1583_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1583_and1 = f_arrdiv32_fs601_xor1 & f_arrdiv32_mux2to1583_not0;
  assign f_arrdiv32_mux2to1583_xor0 = f_arrdiv32_mux2to1583_and0 ^ f_arrdiv32_mux2to1583_and1;
  assign f_arrdiv32_mux2to1584_and0 = f_arrdiv32_mux2to1552_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1584_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1584_and1 = f_arrdiv32_fs602_xor1 & f_arrdiv32_mux2to1584_not0;
  assign f_arrdiv32_mux2to1584_xor0 = f_arrdiv32_mux2to1584_and0 ^ f_arrdiv32_mux2to1584_and1;
  assign f_arrdiv32_mux2to1585_and0 = f_arrdiv32_mux2to1553_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1585_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1585_and1 = f_arrdiv32_fs603_xor1 & f_arrdiv32_mux2to1585_not0;
  assign f_arrdiv32_mux2to1585_xor0 = f_arrdiv32_mux2to1585_and0 ^ f_arrdiv32_mux2to1585_and1;
  assign f_arrdiv32_mux2to1586_and0 = f_arrdiv32_mux2to1554_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1586_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1586_and1 = f_arrdiv32_fs604_xor1 & f_arrdiv32_mux2to1586_not0;
  assign f_arrdiv32_mux2to1586_xor0 = f_arrdiv32_mux2to1586_and0 ^ f_arrdiv32_mux2to1586_and1;
  assign f_arrdiv32_mux2to1587_and0 = f_arrdiv32_mux2to1555_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1587_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1587_and1 = f_arrdiv32_fs605_xor1 & f_arrdiv32_mux2to1587_not0;
  assign f_arrdiv32_mux2to1587_xor0 = f_arrdiv32_mux2to1587_and0 ^ f_arrdiv32_mux2to1587_and1;
  assign f_arrdiv32_mux2to1588_and0 = f_arrdiv32_mux2to1556_xor0 & f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1588_not0 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_mux2to1588_and1 = f_arrdiv32_fs606_xor1 & f_arrdiv32_mux2to1588_not0;
  assign f_arrdiv32_mux2to1588_xor0 = f_arrdiv32_mux2to1588_and0 ^ f_arrdiv32_mux2to1588_and1;
  assign f_arrdiv32_not18 = ~f_arrdiv32_fs607_or0;
  assign f_arrdiv32_fs608_xor0 = a[12] ^ b[0];
  assign f_arrdiv32_fs608_not0 = ~a[12];
  assign f_arrdiv32_fs608_and0 = f_arrdiv32_fs608_not0 & b[0];
  assign f_arrdiv32_fs608_not1 = ~f_arrdiv32_fs608_xor0;
  assign f_arrdiv32_fs609_xor0 = f_arrdiv32_mux2to1558_xor0 ^ b[1];
  assign f_arrdiv32_fs609_not0 = ~f_arrdiv32_mux2to1558_xor0;
  assign f_arrdiv32_fs609_and0 = f_arrdiv32_fs609_not0 & b[1];
  assign f_arrdiv32_fs609_xor1 = f_arrdiv32_fs608_and0 ^ f_arrdiv32_fs609_xor0;
  assign f_arrdiv32_fs609_not1 = ~f_arrdiv32_fs609_xor0;
  assign f_arrdiv32_fs609_and1 = f_arrdiv32_fs609_not1 & f_arrdiv32_fs608_and0;
  assign f_arrdiv32_fs609_or0 = f_arrdiv32_fs609_and1 | f_arrdiv32_fs609_and0;
  assign f_arrdiv32_fs610_xor0 = f_arrdiv32_mux2to1559_xor0 ^ b[2];
  assign f_arrdiv32_fs610_not0 = ~f_arrdiv32_mux2to1559_xor0;
  assign f_arrdiv32_fs610_and0 = f_arrdiv32_fs610_not0 & b[2];
  assign f_arrdiv32_fs610_xor1 = f_arrdiv32_fs609_or0 ^ f_arrdiv32_fs610_xor0;
  assign f_arrdiv32_fs610_not1 = ~f_arrdiv32_fs610_xor0;
  assign f_arrdiv32_fs610_and1 = f_arrdiv32_fs610_not1 & f_arrdiv32_fs609_or0;
  assign f_arrdiv32_fs610_or0 = f_arrdiv32_fs610_and1 | f_arrdiv32_fs610_and0;
  assign f_arrdiv32_fs611_xor0 = f_arrdiv32_mux2to1560_xor0 ^ b[3];
  assign f_arrdiv32_fs611_not0 = ~f_arrdiv32_mux2to1560_xor0;
  assign f_arrdiv32_fs611_and0 = f_arrdiv32_fs611_not0 & b[3];
  assign f_arrdiv32_fs611_xor1 = f_arrdiv32_fs610_or0 ^ f_arrdiv32_fs611_xor0;
  assign f_arrdiv32_fs611_not1 = ~f_arrdiv32_fs611_xor0;
  assign f_arrdiv32_fs611_and1 = f_arrdiv32_fs611_not1 & f_arrdiv32_fs610_or0;
  assign f_arrdiv32_fs611_or0 = f_arrdiv32_fs611_and1 | f_arrdiv32_fs611_and0;
  assign f_arrdiv32_fs612_xor0 = f_arrdiv32_mux2to1561_xor0 ^ b[4];
  assign f_arrdiv32_fs612_not0 = ~f_arrdiv32_mux2to1561_xor0;
  assign f_arrdiv32_fs612_and0 = f_arrdiv32_fs612_not0 & b[4];
  assign f_arrdiv32_fs612_xor1 = f_arrdiv32_fs611_or0 ^ f_arrdiv32_fs612_xor0;
  assign f_arrdiv32_fs612_not1 = ~f_arrdiv32_fs612_xor0;
  assign f_arrdiv32_fs612_and1 = f_arrdiv32_fs612_not1 & f_arrdiv32_fs611_or0;
  assign f_arrdiv32_fs612_or0 = f_arrdiv32_fs612_and1 | f_arrdiv32_fs612_and0;
  assign f_arrdiv32_fs613_xor0 = f_arrdiv32_mux2to1562_xor0 ^ b[5];
  assign f_arrdiv32_fs613_not0 = ~f_arrdiv32_mux2to1562_xor0;
  assign f_arrdiv32_fs613_and0 = f_arrdiv32_fs613_not0 & b[5];
  assign f_arrdiv32_fs613_xor1 = f_arrdiv32_fs612_or0 ^ f_arrdiv32_fs613_xor0;
  assign f_arrdiv32_fs613_not1 = ~f_arrdiv32_fs613_xor0;
  assign f_arrdiv32_fs613_and1 = f_arrdiv32_fs613_not1 & f_arrdiv32_fs612_or0;
  assign f_arrdiv32_fs613_or0 = f_arrdiv32_fs613_and1 | f_arrdiv32_fs613_and0;
  assign f_arrdiv32_fs614_xor0 = f_arrdiv32_mux2to1563_xor0 ^ b[6];
  assign f_arrdiv32_fs614_not0 = ~f_arrdiv32_mux2to1563_xor0;
  assign f_arrdiv32_fs614_and0 = f_arrdiv32_fs614_not0 & b[6];
  assign f_arrdiv32_fs614_xor1 = f_arrdiv32_fs613_or0 ^ f_arrdiv32_fs614_xor0;
  assign f_arrdiv32_fs614_not1 = ~f_arrdiv32_fs614_xor0;
  assign f_arrdiv32_fs614_and1 = f_arrdiv32_fs614_not1 & f_arrdiv32_fs613_or0;
  assign f_arrdiv32_fs614_or0 = f_arrdiv32_fs614_and1 | f_arrdiv32_fs614_and0;
  assign f_arrdiv32_fs615_xor0 = f_arrdiv32_mux2to1564_xor0 ^ b[7];
  assign f_arrdiv32_fs615_not0 = ~f_arrdiv32_mux2to1564_xor0;
  assign f_arrdiv32_fs615_and0 = f_arrdiv32_fs615_not0 & b[7];
  assign f_arrdiv32_fs615_xor1 = f_arrdiv32_fs614_or0 ^ f_arrdiv32_fs615_xor0;
  assign f_arrdiv32_fs615_not1 = ~f_arrdiv32_fs615_xor0;
  assign f_arrdiv32_fs615_and1 = f_arrdiv32_fs615_not1 & f_arrdiv32_fs614_or0;
  assign f_arrdiv32_fs615_or0 = f_arrdiv32_fs615_and1 | f_arrdiv32_fs615_and0;
  assign f_arrdiv32_fs616_xor0 = f_arrdiv32_mux2to1565_xor0 ^ b[8];
  assign f_arrdiv32_fs616_not0 = ~f_arrdiv32_mux2to1565_xor0;
  assign f_arrdiv32_fs616_and0 = f_arrdiv32_fs616_not0 & b[8];
  assign f_arrdiv32_fs616_xor1 = f_arrdiv32_fs615_or0 ^ f_arrdiv32_fs616_xor0;
  assign f_arrdiv32_fs616_not1 = ~f_arrdiv32_fs616_xor0;
  assign f_arrdiv32_fs616_and1 = f_arrdiv32_fs616_not1 & f_arrdiv32_fs615_or0;
  assign f_arrdiv32_fs616_or0 = f_arrdiv32_fs616_and1 | f_arrdiv32_fs616_and0;
  assign f_arrdiv32_fs617_xor0 = f_arrdiv32_mux2to1566_xor0 ^ b[9];
  assign f_arrdiv32_fs617_not0 = ~f_arrdiv32_mux2to1566_xor0;
  assign f_arrdiv32_fs617_and0 = f_arrdiv32_fs617_not0 & b[9];
  assign f_arrdiv32_fs617_xor1 = f_arrdiv32_fs616_or0 ^ f_arrdiv32_fs617_xor0;
  assign f_arrdiv32_fs617_not1 = ~f_arrdiv32_fs617_xor0;
  assign f_arrdiv32_fs617_and1 = f_arrdiv32_fs617_not1 & f_arrdiv32_fs616_or0;
  assign f_arrdiv32_fs617_or0 = f_arrdiv32_fs617_and1 | f_arrdiv32_fs617_and0;
  assign f_arrdiv32_fs618_xor0 = f_arrdiv32_mux2to1567_xor0 ^ b[10];
  assign f_arrdiv32_fs618_not0 = ~f_arrdiv32_mux2to1567_xor0;
  assign f_arrdiv32_fs618_and0 = f_arrdiv32_fs618_not0 & b[10];
  assign f_arrdiv32_fs618_xor1 = f_arrdiv32_fs617_or0 ^ f_arrdiv32_fs618_xor0;
  assign f_arrdiv32_fs618_not1 = ~f_arrdiv32_fs618_xor0;
  assign f_arrdiv32_fs618_and1 = f_arrdiv32_fs618_not1 & f_arrdiv32_fs617_or0;
  assign f_arrdiv32_fs618_or0 = f_arrdiv32_fs618_and1 | f_arrdiv32_fs618_and0;
  assign f_arrdiv32_fs619_xor0 = f_arrdiv32_mux2to1568_xor0 ^ b[11];
  assign f_arrdiv32_fs619_not0 = ~f_arrdiv32_mux2to1568_xor0;
  assign f_arrdiv32_fs619_and0 = f_arrdiv32_fs619_not0 & b[11];
  assign f_arrdiv32_fs619_xor1 = f_arrdiv32_fs618_or0 ^ f_arrdiv32_fs619_xor0;
  assign f_arrdiv32_fs619_not1 = ~f_arrdiv32_fs619_xor0;
  assign f_arrdiv32_fs619_and1 = f_arrdiv32_fs619_not1 & f_arrdiv32_fs618_or0;
  assign f_arrdiv32_fs619_or0 = f_arrdiv32_fs619_and1 | f_arrdiv32_fs619_and0;
  assign f_arrdiv32_fs620_xor0 = f_arrdiv32_mux2to1569_xor0 ^ b[12];
  assign f_arrdiv32_fs620_not0 = ~f_arrdiv32_mux2to1569_xor0;
  assign f_arrdiv32_fs620_and0 = f_arrdiv32_fs620_not0 & b[12];
  assign f_arrdiv32_fs620_xor1 = f_arrdiv32_fs619_or0 ^ f_arrdiv32_fs620_xor0;
  assign f_arrdiv32_fs620_not1 = ~f_arrdiv32_fs620_xor0;
  assign f_arrdiv32_fs620_and1 = f_arrdiv32_fs620_not1 & f_arrdiv32_fs619_or0;
  assign f_arrdiv32_fs620_or0 = f_arrdiv32_fs620_and1 | f_arrdiv32_fs620_and0;
  assign f_arrdiv32_fs621_xor0 = f_arrdiv32_mux2to1570_xor0 ^ b[13];
  assign f_arrdiv32_fs621_not0 = ~f_arrdiv32_mux2to1570_xor0;
  assign f_arrdiv32_fs621_and0 = f_arrdiv32_fs621_not0 & b[13];
  assign f_arrdiv32_fs621_xor1 = f_arrdiv32_fs620_or0 ^ f_arrdiv32_fs621_xor0;
  assign f_arrdiv32_fs621_not1 = ~f_arrdiv32_fs621_xor0;
  assign f_arrdiv32_fs621_and1 = f_arrdiv32_fs621_not1 & f_arrdiv32_fs620_or0;
  assign f_arrdiv32_fs621_or0 = f_arrdiv32_fs621_and1 | f_arrdiv32_fs621_and0;
  assign f_arrdiv32_fs622_xor0 = f_arrdiv32_mux2to1571_xor0 ^ b[14];
  assign f_arrdiv32_fs622_not0 = ~f_arrdiv32_mux2to1571_xor0;
  assign f_arrdiv32_fs622_and0 = f_arrdiv32_fs622_not0 & b[14];
  assign f_arrdiv32_fs622_xor1 = f_arrdiv32_fs621_or0 ^ f_arrdiv32_fs622_xor0;
  assign f_arrdiv32_fs622_not1 = ~f_arrdiv32_fs622_xor0;
  assign f_arrdiv32_fs622_and1 = f_arrdiv32_fs622_not1 & f_arrdiv32_fs621_or0;
  assign f_arrdiv32_fs622_or0 = f_arrdiv32_fs622_and1 | f_arrdiv32_fs622_and0;
  assign f_arrdiv32_fs623_xor0 = f_arrdiv32_mux2to1572_xor0 ^ b[15];
  assign f_arrdiv32_fs623_not0 = ~f_arrdiv32_mux2to1572_xor0;
  assign f_arrdiv32_fs623_and0 = f_arrdiv32_fs623_not0 & b[15];
  assign f_arrdiv32_fs623_xor1 = f_arrdiv32_fs622_or0 ^ f_arrdiv32_fs623_xor0;
  assign f_arrdiv32_fs623_not1 = ~f_arrdiv32_fs623_xor0;
  assign f_arrdiv32_fs623_and1 = f_arrdiv32_fs623_not1 & f_arrdiv32_fs622_or0;
  assign f_arrdiv32_fs623_or0 = f_arrdiv32_fs623_and1 | f_arrdiv32_fs623_and0;
  assign f_arrdiv32_fs624_xor0 = f_arrdiv32_mux2to1573_xor0 ^ b[16];
  assign f_arrdiv32_fs624_not0 = ~f_arrdiv32_mux2to1573_xor0;
  assign f_arrdiv32_fs624_and0 = f_arrdiv32_fs624_not0 & b[16];
  assign f_arrdiv32_fs624_xor1 = f_arrdiv32_fs623_or0 ^ f_arrdiv32_fs624_xor0;
  assign f_arrdiv32_fs624_not1 = ~f_arrdiv32_fs624_xor0;
  assign f_arrdiv32_fs624_and1 = f_arrdiv32_fs624_not1 & f_arrdiv32_fs623_or0;
  assign f_arrdiv32_fs624_or0 = f_arrdiv32_fs624_and1 | f_arrdiv32_fs624_and0;
  assign f_arrdiv32_fs625_xor0 = f_arrdiv32_mux2to1574_xor0 ^ b[17];
  assign f_arrdiv32_fs625_not0 = ~f_arrdiv32_mux2to1574_xor0;
  assign f_arrdiv32_fs625_and0 = f_arrdiv32_fs625_not0 & b[17];
  assign f_arrdiv32_fs625_xor1 = f_arrdiv32_fs624_or0 ^ f_arrdiv32_fs625_xor0;
  assign f_arrdiv32_fs625_not1 = ~f_arrdiv32_fs625_xor0;
  assign f_arrdiv32_fs625_and1 = f_arrdiv32_fs625_not1 & f_arrdiv32_fs624_or0;
  assign f_arrdiv32_fs625_or0 = f_arrdiv32_fs625_and1 | f_arrdiv32_fs625_and0;
  assign f_arrdiv32_fs626_xor0 = f_arrdiv32_mux2to1575_xor0 ^ b[18];
  assign f_arrdiv32_fs626_not0 = ~f_arrdiv32_mux2to1575_xor0;
  assign f_arrdiv32_fs626_and0 = f_arrdiv32_fs626_not0 & b[18];
  assign f_arrdiv32_fs626_xor1 = f_arrdiv32_fs625_or0 ^ f_arrdiv32_fs626_xor0;
  assign f_arrdiv32_fs626_not1 = ~f_arrdiv32_fs626_xor0;
  assign f_arrdiv32_fs626_and1 = f_arrdiv32_fs626_not1 & f_arrdiv32_fs625_or0;
  assign f_arrdiv32_fs626_or0 = f_arrdiv32_fs626_and1 | f_arrdiv32_fs626_and0;
  assign f_arrdiv32_fs627_xor0 = f_arrdiv32_mux2to1576_xor0 ^ b[19];
  assign f_arrdiv32_fs627_not0 = ~f_arrdiv32_mux2to1576_xor0;
  assign f_arrdiv32_fs627_and0 = f_arrdiv32_fs627_not0 & b[19];
  assign f_arrdiv32_fs627_xor1 = f_arrdiv32_fs626_or0 ^ f_arrdiv32_fs627_xor0;
  assign f_arrdiv32_fs627_not1 = ~f_arrdiv32_fs627_xor0;
  assign f_arrdiv32_fs627_and1 = f_arrdiv32_fs627_not1 & f_arrdiv32_fs626_or0;
  assign f_arrdiv32_fs627_or0 = f_arrdiv32_fs627_and1 | f_arrdiv32_fs627_and0;
  assign f_arrdiv32_fs628_xor0 = f_arrdiv32_mux2to1577_xor0 ^ b[20];
  assign f_arrdiv32_fs628_not0 = ~f_arrdiv32_mux2to1577_xor0;
  assign f_arrdiv32_fs628_and0 = f_arrdiv32_fs628_not0 & b[20];
  assign f_arrdiv32_fs628_xor1 = f_arrdiv32_fs627_or0 ^ f_arrdiv32_fs628_xor0;
  assign f_arrdiv32_fs628_not1 = ~f_arrdiv32_fs628_xor0;
  assign f_arrdiv32_fs628_and1 = f_arrdiv32_fs628_not1 & f_arrdiv32_fs627_or0;
  assign f_arrdiv32_fs628_or0 = f_arrdiv32_fs628_and1 | f_arrdiv32_fs628_and0;
  assign f_arrdiv32_fs629_xor0 = f_arrdiv32_mux2to1578_xor0 ^ b[21];
  assign f_arrdiv32_fs629_not0 = ~f_arrdiv32_mux2to1578_xor0;
  assign f_arrdiv32_fs629_and0 = f_arrdiv32_fs629_not0 & b[21];
  assign f_arrdiv32_fs629_xor1 = f_arrdiv32_fs628_or0 ^ f_arrdiv32_fs629_xor0;
  assign f_arrdiv32_fs629_not1 = ~f_arrdiv32_fs629_xor0;
  assign f_arrdiv32_fs629_and1 = f_arrdiv32_fs629_not1 & f_arrdiv32_fs628_or0;
  assign f_arrdiv32_fs629_or0 = f_arrdiv32_fs629_and1 | f_arrdiv32_fs629_and0;
  assign f_arrdiv32_fs630_xor0 = f_arrdiv32_mux2to1579_xor0 ^ b[22];
  assign f_arrdiv32_fs630_not0 = ~f_arrdiv32_mux2to1579_xor0;
  assign f_arrdiv32_fs630_and0 = f_arrdiv32_fs630_not0 & b[22];
  assign f_arrdiv32_fs630_xor1 = f_arrdiv32_fs629_or0 ^ f_arrdiv32_fs630_xor0;
  assign f_arrdiv32_fs630_not1 = ~f_arrdiv32_fs630_xor0;
  assign f_arrdiv32_fs630_and1 = f_arrdiv32_fs630_not1 & f_arrdiv32_fs629_or0;
  assign f_arrdiv32_fs630_or0 = f_arrdiv32_fs630_and1 | f_arrdiv32_fs630_and0;
  assign f_arrdiv32_fs631_xor0 = f_arrdiv32_mux2to1580_xor0 ^ b[23];
  assign f_arrdiv32_fs631_not0 = ~f_arrdiv32_mux2to1580_xor0;
  assign f_arrdiv32_fs631_and0 = f_arrdiv32_fs631_not0 & b[23];
  assign f_arrdiv32_fs631_xor1 = f_arrdiv32_fs630_or0 ^ f_arrdiv32_fs631_xor0;
  assign f_arrdiv32_fs631_not1 = ~f_arrdiv32_fs631_xor0;
  assign f_arrdiv32_fs631_and1 = f_arrdiv32_fs631_not1 & f_arrdiv32_fs630_or0;
  assign f_arrdiv32_fs631_or0 = f_arrdiv32_fs631_and1 | f_arrdiv32_fs631_and0;
  assign f_arrdiv32_fs632_xor0 = f_arrdiv32_mux2to1581_xor0 ^ b[24];
  assign f_arrdiv32_fs632_not0 = ~f_arrdiv32_mux2to1581_xor0;
  assign f_arrdiv32_fs632_and0 = f_arrdiv32_fs632_not0 & b[24];
  assign f_arrdiv32_fs632_xor1 = f_arrdiv32_fs631_or0 ^ f_arrdiv32_fs632_xor0;
  assign f_arrdiv32_fs632_not1 = ~f_arrdiv32_fs632_xor0;
  assign f_arrdiv32_fs632_and1 = f_arrdiv32_fs632_not1 & f_arrdiv32_fs631_or0;
  assign f_arrdiv32_fs632_or0 = f_arrdiv32_fs632_and1 | f_arrdiv32_fs632_and0;
  assign f_arrdiv32_fs633_xor0 = f_arrdiv32_mux2to1582_xor0 ^ b[25];
  assign f_arrdiv32_fs633_not0 = ~f_arrdiv32_mux2to1582_xor0;
  assign f_arrdiv32_fs633_and0 = f_arrdiv32_fs633_not0 & b[25];
  assign f_arrdiv32_fs633_xor1 = f_arrdiv32_fs632_or0 ^ f_arrdiv32_fs633_xor0;
  assign f_arrdiv32_fs633_not1 = ~f_arrdiv32_fs633_xor0;
  assign f_arrdiv32_fs633_and1 = f_arrdiv32_fs633_not1 & f_arrdiv32_fs632_or0;
  assign f_arrdiv32_fs633_or0 = f_arrdiv32_fs633_and1 | f_arrdiv32_fs633_and0;
  assign f_arrdiv32_fs634_xor0 = f_arrdiv32_mux2to1583_xor0 ^ b[26];
  assign f_arrdiv32_fs634_not0 = ~f_arrdiv32_mux2to1583_xor0;
  assign f_arrdiv32_fs634_and0 = f_arrdiv32_fs634_not0 & b[26];
  assign f_arrdiv32_fs634_xor1 = f_arrdiv32_fs633_or0 ^ f_arrdiv32_fs634_xor0;
  assign f_arrdiv32_fs634_not1 = ~f_arrdiv32_fs634_xor0;
  assign f_arrdiv32_fs634_and1 = f_arrdiv32_fs634_not1 & f_arrdiv32_fs633_or0;
  assign f_arrdiv32_fs634_or0 = f_arrdiv32_fs634_and1 | f_arrdiv32_fs634_and0;
  assign f_arrdiv32_fs635_xor0 = f_arrdiv32_mux2to1584_xor0 ^ b[27];
  assign f_arrdiv32_fs635_not0 = ~f_arrdiv32_mux2to1584_xor0;
  assign f_arrdiv32_fs635_and0 = f_arrdiv32_fs635_not0 & b[27];
  assign f_arrdiv32_fs635_xor1 = f_arrdiv32_fs634_or0 ^ f_arrdiv32_fs635_xor0;
  assign f_arrdiv32_fs635_not1 = ~f_arrdiv32_fs635_xor0;
  assign f_arrdiv32_fs635_and1 = f_arrdiv32_fs635_not1 & f_arrdiv32_fs634_or0;
  assign f_arrdiv32_fs635_or0 = f_arrdiv32_fs635_and1 | f_arrdiv32_fs635_and0;
  assign f_arrdiv32_fs636_xor0 = f_arrdiv32_mux2to1585_xor0 ^ b[28];
  assign f_arrdiv32_fs636_not0 = ~f_arrdiv32_mux2to1585_xor0;
  assign f_arrdiv32_fs636_and0 = f_arrdiv32_fs636_not0 & b[28];
  assign f_arrdiv32_fs636_xor1 = f_arrdiv32_fs635_or0 ^ f_arrdiv32_fs636_xor0;
  assign f_arrdiv32_fs636_not1 = ~f_arrdiv32_fs636_xor0;
  assign f_arrdiv32_fs636_and1 = f_arrdiv32_fs636_not1 & f_arrdiv32_fs635_or0;
  assign f_arrdiv32_fs636_or0 = f_arrdiv32_fs636_and1 | f_arrdiv32_fs636_and0;
  assign f_arrdiv32_fs637_xor0 = f_arrdiv32_mux2to1586_xor0 ^ b[29];
  assign f_arrdiv32_fs637_not0 = ~f_arrdiv32_mux2to1586_xor0;
  assign f_arrdiv32_fs637_and0 = f_arrdiv32_fs637_not0 & b[29];
  assign f_arrdiv32_fs637_xor1 = f_arrdiv32_fs636_or0 ^ f_arrdiv32_fs637_xor0;
  assign f_arrdiv32_fs637_not1 = ~f_arrdiv32_fs637_xor0;
  assign f_arrdiv32_fs637_and1 = f_arrdiv32_fs637_not1 & f_arrdiv32_fs636_or0;
  assign f_arrdiv32_fs637_or0 = f_arrdiv32_fs637_and1 | f_arrdiv32_fs637_and0;
  assign f_arrdiv32_fs638_xor0 = f_arrdiv32_mux2to1587_xor0 ^ b[30];
  assign f_arrdiv32_fs638_not0 = ~f_arrdiv32_mux2to1587_xor0;
  assign f_arrdiv32_fs638_and0 = f_arrdiv32_fs638_not0 & b[30];
  assign f_arrdiv32_fs638_xor1 = f_arrdiv32_fs637_or0 ^ f_arrdiv32_fs638_xor0;
  assign f_arrdiv32_fs638_not1 = ~f_arrdiv32_fs638_xor0;
  assign f_arrdiv32_fs638_and1 = f_arrdiv32_fs638_not1 & f_arrdiv32_fs637_or0;
  assign f_arrdiv32_fs638_or0 = f_arrdiv32_fs638_and1 | f_arrdiv32_fs638_and0;
  assign f_arrdiv32_fs639_xor0 = f_arrdiv32_mux2to1588_xor0 ^ b[31];
  assign f_arrdiv32_fs639_not0 = ~f_arrdiv32_mux2to1588_xor0;
  assign f_arrdiv32_fs639_and0 = f_arrdiv32_fs639_not0 & b[31];
  assign f_arrdiv32_fs639_xor1 = f_arrdiv32_fs638_or0 ^ f_arrdiv32_fs639_xor0;
  assign f_arrdiv32_fs639_not1 = ~f_arrdiv32_fs639_xor0;
  assign f_arrdiv32_fs639_and1 = f_arrdiv32_fs639_not1 & f_arrdiv32_fs638_or0;
  assign f_arrdiv32_fs639_or0 = f_arrdiv32_fs639_and1 | f_arrdiv32_fs639_and0;
  assign f_arrdiv32_mux2to1589_and0 = a[12] & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1589_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1589_and1 = f_arrdiv32_fs608_xor0 & f_arrdiv32_mux2to1589_not0;
  assign f_arrdiv32_mux2to1589_xor0 = f_arrdiv32_mux2to1589_and0 ^ f_arrdiv32_mux2to1589_and1;
  assign f_arrdiv32_mux2to1590_and0 = f_arrdiv32_mux2to1558_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1590_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1590_and1 = f_arrdiv32_fs609_xor1 & f_arrdiv32_mux2to1590_not0;
  assign f_arrdiv32_mux2to1590_xor0 = f_arrdiv32_mux2to1590_and0 ^ f_arrdiv32_mux2to1590_and1;
  assign f_arrdiv32_mux2to1591_and0 = f_arrdiv32_mux2to1559_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1591_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1591_and1 = f_arrdiv32_fs610_xor1 & f_arrdiv32_mux2to1591_not0;
  assign f_arrdiv32_mux2to1591_xor0 = f_arrdiv32_mux2to1591_and0 ^ f_arrdiv32_mux2to1591_and1;
  assign f_arrdiv32_mux2to1592_and0 = f_arrdiv32_mux2to1560_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1592_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1592_and1 = f_arrdiv32_fs611_xor1 & f_arrdiv32_mux2to1592_not0;
  assign f_arrdiv32_mux2to1592_xor0 = f_arrdiv32_mux2to1592_and0 ^ f_arrdiv32_mux2to1592_and1;
  assign f_arrdiv32_mux2to1593_and0 = f_arrdiv32_mux2to1561_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1593_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1593_and1 = f_arrdiv32_fs612_xor1 & f_arrdiv32_mux2to1593_not0;
  assign f_arrdiv32_mux2to1593_xor0 = f_arrdiv32_mux2to1593_and0 ^ f_arrdiv32_mux2to1593_and1;
  assign f_arrdiv32_mux2to1594_and0 = f_arrdiv32_mux2to1562_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1594_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1594_and1 = f_arrdiv32_fs613_xor1 & f_arrdiv32_mux2to1594_not0;
  assign f_arrdiv32_mux2to1594_xor0 = f_arrdiv32_mux2to1594_and0 ^ f_arrdiv32_mux2to1594_and1;
  assign f_arrdiv32_mux2to1595_and0 = f_arrdiv32_mux2to1563_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1595_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1595_and1 = f_arrdiv32_fs614_xor1 & f_arrdiv32_mux2to1595_not0;
  assign f_arrdiv32_mux2to1595_xor0 = f_arrdiv32_mux2to1595_and0 ^ f_arrdiv32_mux2to1595_and1;
  assign f_arrdiv32_mux2to1596_and0 = f_arrdiv32_mux2to1564_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1596_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1596_and1 = f_arrdiv32_fs615_xor1 & f_arrdiv32_mux2to1596_not0;
  assign f_arrdiv32_mux2to1596_xor0 = f_arrdiv32_mux2to1596_and0 ^ f_arrdiv32_mux2to1596_and1;
  assign f_arrdiv32_mux2to1597_and0 = f_arrdiv32_mux2to1565_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1597_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1597_and1 = f_arrdiv32_fs616_xor1 & f_arrdiv32_mux2to1597_not0;
  assign f_arrdiv32_mux2to1597_xor0 = f_arrdiv32_mux2to1597_and0 ^ f_arrdiv32_mux2to1597_and1;
  assign f_arrdiv32_mux2to1598_and0 = f_arrdiv32_mux2to1566_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1598_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1598_and1 = f_arrdiv32_fs617_xor1 & f_arrdiv32_mux2to1598_not0;
  assign f_arrdiv32_mux2to1598_xor0 = f_arrdiv32_mux2to1598_and0 ^ f_arrdiv32_mux2to1598_and1;
  assign f_arrdiv32_mux2to1599_and0 = f_arrdiv32_mux2to1567_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1599_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1599_and1 = f_arrdiv32_fs618_xor1 & f_arrdiv32_mux2to1599_not0;
  assign f_arrdiv32_mux2to1599_xor0 = f_arrdiv32_mux2to1599_and0 ^ f_arrdiv32_mux2to1599_and1;
  assign f_arrdiv32_mux2to1600_and0 = f_arrdiv32_mux2to1568_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1600_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1600_and1 = f_arrdiv32_fs619_xor1 & f_arrdiv32_mux2to1600_not0;
  assign f_arrdiv32_mux2to1600_xor0 = f_arrdiv32_mux2to1600_and0 ^ f_arrdiv32_mux2to1600_and1;
  assign f_arrdiv32_mux2to1601_and0 = f_arrdiv32_mux2to1569_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1601_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1601_and1 = f_arrdiv32_fs620_xor1 & f_arrdiv32_mux2to1601_not0;
  assign f_arrdiv32_mux2to1601_xor0 = f_arrdiv32_mux2to1601_and0 ^ f_arrdiv32_mux2to1601_and1;
  assign f_arrdiv32_mux2to1602_and0 = f_arrdiv32_mux2to1570_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1602_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1602_and1 = f_arrdiv32_fs621_xor1 & f_arrdiv32_mux2to1602_not0;
  assign f_arrdiv32_mux2to1602_xor0 = f_arrdiv32_mux2to1602_and0 ^ f_arrdiv32_mux2to1602_and1;
  assign f_arrdiv32_mux2to1603_and0 = f_arrdiv32_mux2to1571_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1603_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1603_and1 = f_arrdiv32_fs622_xor1 & f_arrdiv32_mux2to1603_not0;
  assign f_arrdiv32_mux2to1603_xor0 = f_arrdiv32_mux2to1603_and0 ^ f_arrdiv32_mux2to1603_and1;
  assign f_arrdiv32_mux2to1604_and0 = f_arrdiv32_mux2to1572_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1604_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1604_and1 = f_arrdiv32_fs623_xor1 & f_arrdiv32_mux2to1604_not0;
  assign f_arrdiv32_mux2to1604_xor0 = f_arrdiv32_mux2to1604_and0 ^ f_arrdiv32_mux2to1604_and1;
  assign f_arrdiv32_mux2to1605_and0 = f_arrdiv32_mux2to1573_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1605_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1605_and1 = f_arrdiv32_fs624_xor1 & f_arrdiv32_mux2to1605_not0;
  assign f_arrdiv32_mux2to1605_xor0 = f_arrdiv32_mux2to1605_and0 ^ f_arrdiv32_mux2to1605_and1;
  assign f_arrdiv32_mux2to1606_and0 = f_arrdiv32_mux2to1574_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1606_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1606_and1 = f_arrdiv32_fs625_xor1 & f_arrdiv32_mux2to1606_not0;
  assign f_arrdiv32_mux2to1606_xor0 = f_arrdiv32_mux2to1606_and0 ^ f_arrdiv32_mux2to1606_and1;
  assign f_arrdiv32_mux2to1607_and0 = f_arrdiv32_mux2to1575_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1607_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1607_and1 = f_arrdiv32_fs626_xor1 & f_arrdiv32_mux2to1607_not0;
  assign f_arrdiv32_mux2to1607_xor0 = f_arrdiv32_mux2to1607_and0 ^ f_arrdiv32_mux2to1607_and1;
  assign f_arrdiv32_mux2to1608_and0 = f_arrdiv32_mux2to1576_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1608_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1608_and1 = f_arrdiv32_fs627_xor1 & f_arrdiv32_mux2to1608_not0;
  assign f_arrdiv32_mux2to1608_xor0 = f_arrdiv32_mux2to1608_and0 ^ f_arrdiv32_mux2to1608_and1;
  assign f_arrdiv32_mux2to1609_and0 = f_arrdiv32_mux2to1577_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1609_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1609_and1 = f_arrdiv32_fs628_xor1 & f_arrdiv32_mux2to1609_not0;
  assign f_arrdiv32_mux2to1609_xor0 = f_arrdiv32_mux2to1609_and0 ^ f_arrdiv32_mux2to1609_and1;
  assign f_arrdiv32_mux2to1610_and0 = f_arrdiv32_mux2to1578_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1610_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1610_and1 = f_arrdiv32_fs629_xor1 & f_arrdiv32_mux2to1610_not0;
  assign f_arrdiv32_mux2to1610_xor0 = f_arrdiv32_mux2to1610_and0 ^ f_arrdiv32_mux2to1610_and1;
  assign f_arrdiv32_mux2to1611_and0 = f_arrdiv32_mux2to1579_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1611_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1611_and1 = f_arrdiv32_fs630_xor1 & f_arrdiv32_mux2to1611_not0;
  assign f_arrdiv32_mux2to1611_xor0 = f_arrdiv32_mux2to1611_and0 ^ f_arrdiv32_mux2to1611_and1;
  assign f_arrdiv32_mux2to1612_and0 = f_arrdiv32_mux2to1580_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1612_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1612_and1 = f_arrdiv32_fs631_xor1 & f_arrdiv32_mux2to1612_not0;
  assign f_arrdiv32_mux2to1612_xor0 = f_arrdiv32_mux2to1612_and0 ^ f_arrdiv32_mux2to1612_and1;
  assign f_arrdiv32_mux2to1613_and0 = f_arrdiv32_mux2to1581_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1613_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1613_and1 = f_arrdiv32_fs632_xor1 & f_arrdiv32_mux2to1613_not0;
  assign f_arrdiv32_mux2to1613_xor0 = f_arrdiv32_mux2to1613_and0 ^ f_arrdiv32_mux2to1613_and1;
  assign f_arrdiv32_mux2to1614_and0 = f_arrdiv32_mux2to1582_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1614_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1614_and1 = f_arrdiv32_fs633_xor1 & f_arrdiv32_mux2to1614_not0;
  assign f_arrdiv32_mux2to1614_xor0 = f_arrdiv32_mux2to1614_and0 ^ f_arrdiv32_mux2to1614_and1;
  assign f_arrdiv32_mux2to1615_and0 = f_arrdiv32_mux2to1583_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1615_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1615_and1 = f_arrdiv32_fs634_xor1 & f_arrdiv32_mux2to1615_not0;
  assign f_arrdiv32_mux2to1615_xor0 = f_arrdiv32_mux2to1615_and0 ^ f_arrdiv32_mux2to1615_and1;
  assign f_arrdiv32_mux2to1616_and0 = f_arrdiv32_mux2to1584_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1616_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1616_and1 = f_arrdiv32_fs635_xor1 & f_arrdiv32_mux2to1616_not0;
  assign f_arrdiv32_mux2to1616_xor0 = f_arrdiv32_mux2to1616_and0 ^ f_arrdiv32_mux2to1616_and1;
  assign f_arrdiv32_mux2to1617_and0 = f_arrdiv32_mux2to1585_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1617_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1617_and1 = f_arrdiv32_fs636_xor1 & f_arrdiv32_mux2to1617_not0;
  assign f_arrdiv32_mux2to1617_xor0 = f_arrdiv32_mux2to1617_and0 ^ f_arrdiv32_mux2to1617_and1;
  assign f_arrdiv32_mux2to1618_and0 = f_arrdiv32_mux2to1586_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1618_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1618_and1 = f_arrdiv32_fs637_xor1 & f_arrdiv32_mux2to1618_not0;
  assign f_arrdiv32_mux2to1618_xor0 = f_arrdiv32_mux2to1618_and0 ^ f_arrdiv32_mux2to1618_and1;
  assign f_arrdiv32_mux2to1619_and0 = f_arrdiv32_mux2to1587_xor0 & f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1619_not0 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_mux2to1619_and1 = f_arrdiv32_fs638_xor1 & f_arrdiv32_mux2to1619_not0;
  assign f_arrdiv32_mux2to1619_xor0 = f_arrdiv32_mux2to1619_and0 ^ f_arrdiv32_mux2to1619_and1;
  assign f_arrdiv32_not19 = ~f_arrdiv32_fs639_or0;
  assign f_arrdiv32_fs640_xor0 = a[11] ^ b[0];
  assign f_arrdiv32_fs640_not0 = ~a[11];
  assign f_arrdiv32_fs640_and0 = f_arrdiv32_fs640_not0 & b[0];
  assign f_arrdiv32_fs640_not1 = ~f_arrdiv32_fs640_xor0;
  assign f_arrdiv32_fs641_xor0 = f_arrdiv32_mux2to1589_xor0 ^ b[1];
  assign f_arrdiv32_fs641_not0 = ~f_arrdiv32_mux2to1589_xor0;
  assign f_arrdiv32_fs641_and0 = f_arrdiv32_fs641_not0 & b[1];
  assign f_arrdiv32_fs641_xor1 = f_arrdiv32_fs640_and0 ^ f_arrdiv32_fs641_xor0;
  assign f_arrdiv32_fs641_not1 = ~f_arrdiv32_fs641_xor0;
  assign f_arrdiv32_fs641_and1 = f_arrdiv32_fs641_not1 & f_arrdiv32_fs640_and0;
  assign f_arrdiv32_fs641_or0 = f_arrdiv32_fs641_and1 | f_arrdiv32_fs641_and0;
  assign f_arrdiv32_fs642_xor0 = f_arrdiv32_mux2to1590_xor0 ^ b[2];
  assign f_arrdiv32_fs642_not0 = ~f_arrdiv32_mux2to1590_xor0;
  assign f_arrdiv32_fs642_and0 = f_arrdiv32_fs642_not0 & b[2];
  assign f_arrdiv32_fs642_xor1 = f_arrdiv32_fs641_or0 ^ f_arrdiv32_fs642_xor0;
  assign f_arrdiv32_fs642_not1 = ~f_arrdiv32_fs642_xor0;
  assign f_arrdiv32_fs642_and1 = f_arrdiv32_fs642_not1 & f_arrdiv32_fs641_or0;
  assign f_arrdiv32_fs642_or0 = f_arrdiv32_fs642_and1 | f_arrdiv32_fs642_and0;
  assign f_arrdiv32_fs643_xor0 = f_arrdiv32_mux2to1591_xor0 ^ b[3];
  assign f_arrdiv32_fs643_not0 = ~f_arrdiv32_mux2to1591_xor0;
  assign f_arrdiv32_fs643_and0 = f_arrdiv32_fs643_not0 & b[3];
  assign f_arrdiv32_fs643_xor1 = f_arrdiv32_fs642_or0 ^ f_arrdiv32_fs643_xor0;
  assign f_arrdiv32_fs643_not1 = ~f_arrdiv32_fs643_xor0;
  assign f_arrdiv32_fs643_and1 = f_arrdiv32_fs643_not1 & f_arrdiv32_fs642_or0;
  assign f_arrdiv32_fs643_or0 = f_arrdiv32_fs643_and1 | f_arrdiv32_fs643_and0;
  assign f_arrdiv32_fs644_xor0 = f_arrdiv32_mux2to1592_xor0 ^ b[4];
  assign f_arrdiv32_fs644_not0 = ~f_arrdiv32_mux2to1592_xor0;
  assign f_arrdiv32_fs644_and0 = f_arrdiv32_fs644_not0 & b[4];
  assign f_arrdiv32_fs644_xor1 = f_arrdiv32_fs643_or0 ^ f_arrdiv32_fs644_xor0;
  assign f_arrdiv32_fs644_not1 = ~f_arrdiv32_fs644_xor0;
  assign f_arrdiv32_fs644_and1 = f_arrdiv32_fs644_not1 & f_arrdiv32_fs643_or0;
  assign f_arrdiv32_fs644_or0 = f_arrdiv32_fs644_and1 | f_arrdiv32_fs644_and0;
  assign f_arrdiv32_fs645_xor0 = f_arrdiv32_mux2to1593_xor0 ^ b[5];
  assign f_arrdiv32_fs645_not0 = ~f_arrdiv32_mux2to1593_xor0;
  assign f_arrdiv32_fs645_and0 = f_arrdiv32_fs645_not0 & b[5];
  assign f_arrdiv32_fs645_xor1 = f_arrdiv32_fs644_or0 ^ f_arrdiv32_fs645_xor0;
  assign f_arrdiv32_fs645_not1 = ~f_arrdiv32_fs645_xor0;
  assign f_arrdiv32_fs645_and1 = f_arrdiv32_fs645_not1 & f_arrdiv32_fs644_or0;
  assign f_arrdiv32_fs645_or0 = f_arrdiv32_fs645_and1 | f_arrdiv32_fs645_and0;
  assign f_arrdiv32_fs646_xor0 = f_arrdiv32_mux2to1594_xor0 ^ b[6];
  assign f_arrdiv32_fs646_not0 = ~f_arrdiv32_mux2to1594_xor0;
  assign f_arrdiv32_fs646_and0 = f_arrdiv32_fs646_not0 & b[6];
  assign f_arrdiv32_fs646_xor1 = f_arrdiv32_fs645_or0 ^ f_arrdiv32_fs646_xor0;
  assign f_arrdiv32_fs646_not1 = ~f_arrdiv32_fs646_xor0;
  assign f_arrdiv32_fs646_and1 = f_arrdiv32_fs646_not1 & f_arrdiv32_fs645_or0;
  assign f_arrdiv32_fs646_or0 = f_arrdiv32_fs646_and1 | f_arrdiv32_fs646_and0;
  assign f_arrdiv32_fs647_xor0 = f_arrdiv32_mux2to1595_xor0 ^ b[7];
  assign f_arrdiv32_fs647_not0 = ~f_arrdiv32_mux2to1595_xor0;
  assign f_arrdiv32_fs647_and0 = f_arrdiv32_fs647_not0 & b[7];
  assign f_arrdiv32_fs647_xor1 = f_arrdiv32_fs646_or0 ^ f_arrdiv32_fs647_xor0;
  assign f_arrdiv32_fs647_not1 = ~f_arrdiv32_fs647_xor0;
  assign f_arrdiv32_fs647_and1 = f_arrdiv32_fs647_not1 & f_arrdiv32_fs646_or0;
  assign f_arrdiv32_fs647_or0 = f_arrdiv32_fs647_and1 | f_arrdiv32_fs647_and0;
  assign f_arrdiv32_fs648_xor0 = f_arrdiv32_mux2to1596_xor0 ^ b[8];
  assign f_arrdiv32_fs648_not0 = ~f_arrdiv32_mux2to1596_xor0;
  assign f_arrdiv32_fs648_and0 = f_arrdiv32_fs648_not0 & b[8];
  assign f_arrdiv32_fs648_xor1 = f_arrdiv32_fs647_or0 ^ f_arrdiv32_fs648_xor0;
  assign f_arrdiv32_fs648_not1 = ~f_arrdiv32_fs648_xor0;
  assign f_arrdiv32_fs648_and1 = f_arrdiv32_fs648_not1 & f_arrdiv32_fs647_or0;
  assign f_arrdiv32_fs648_or0 = f_arrdiv32_fs648_and1 | f_arrdiv32_fs648_and0;
  assign f_arrdiv32_fs649_xor0 = f_arrdiv32_mux2to1597_xor0 ^ b[9];
  assign f_arrdiv32_fs649_not0 = ~f_arrdiv32_mux2to1597_xor0;
  assign f_arrdiv32_fs649_and0 = f_arrdiv32_fs649_not0 & b[9];
  assign f_arrdiv32_fs649_xor1 = f_arrdiv32_fs648_or0 ^ f_arrdiv32_fs649_xor0;
  assign f_arrdiv32_fs649_not1 = ~f_arrdiv32_fs649_xor0;
  assign f_arrdiv32_fs649_and1 = f_arrdiv32_fs649_not1 & f_arrdiv32_fs648_or0;
  assign f_arrdiv32_fs649_or0 = f_arrdiv32_fs649_and1 | f_arrdiv32_fs649_and0;
  assign f_arrdiv32_fs650_xor0 = f_arrdiv32_mux2to1598_xor0 ^ b[10];
  assign f_arrdiv32_fs650_not0 = ~f_arrdiv32_mux2to1598_xor0;
  assign f_arrdiv32_fs650_and0 = f_arrdiv32_fs650_not0 & b[10];
  assign f_arrdiv32_fs650_xor1 = f_arrdiv32_fs649_or0 ^ f_arrdiv32_fs650_xor0;
  assign f_arrdiv32_fs650_not1 = ~f_arrdiv32_fs650_xor0;
  assign f_arrdiv32_fs650_and1 = f_arrdiv32_fs650_not1 & f_arrdiv32_fs649_or0;
  assign f_arrdiv32_fs650_or0 = f_arrdiv32_fs650_and1 | f_arrdiv32_fs650_and0;
  assign f_arrdiv32_fs651_xor0 = f_arrdiv32_mux2to1599_xor0 ^ b[11];
  assign f_arrdiv32_fs651_not0 = ~f_arrdiv32_mux2to1599_xor0;
  assign f_arrdiv32_fs651_and0 = f_arrdiv32_fs651_not0 & b[11];
  assign f_arrdiv32_fs651_xor1 = f_arrdiv32_fs650_or0 ^ f_arrdiv32_fs651_xor0;
  assign f_arrdiv32_fs651_not1 = ~f_arrdiv32_fs651_xor0;
  assign f_arrdiv32_fs651_and1 = f_arrdiv32_fs651_not1 & f_arrdiv32_fs650_or0;
  assign f_arrdiv32_fs651_or0 = f_arrdiv32_fs651_and1 | f_arrdiv32_fs651_and0;
  assign f_arrdiv32_fs652_xor0 = f_arrdiv32_mux2to1600_xor0 ^ b[12];
  assign f_arrdiv32_fs652_not0 = ~f_arrdiv32_mux2to1600_xor0;
  assign f_arrdiv32_fs652_and0 = f_arrdiv32_fs652_not0 & b[12];
  assign f_arrdiv32_fs652_xor1 = f_arrdiv32_fs651_or0 ^ f_arrdiv32_fs652_xor0;
  assign f_arrdiv32_fs652_not1 = ~f_arrdiv32_fs652_xor0;
  assign f_arrdiv32_fs652_and1 = f_arrdiv32_fs652_not1 & f_arrdiv32_fs651_or0;
  assign f_arrdiv32_fs652_or0 = f_arrdiv32_fs652_and1 | f_arrdiv32_fs652_and0;
  assign f_arrdiv32_fs653_xor0 = f_arrdiv32_mux2to1601_xor0 ^ b[13];
  assign f_arrdiv32_fs653_not0 = ~f_arrdiv32_mux2to1601_xor0;
  assign f_arrdiv32_fs653_and0 = f_arrdiv32_fs653_not0 & b[13];
  assign f_arrdiv32_fs653_xor1 = f_arrdiv32_fs652_or0 ^ f_arrdiv32_fs653_xor0;
  assign f_arrdiv32_fs653_not1 = ~f_arrdiv32_fs653_xor0;
  assign f_arrdiv32_fs653_and1 = f_arrdiv32_fs653_not1 & f_arrdiv32_fs652_or0;
  assign f_arrdiv32_fs653_or0 = f_arrdiv32_fs653_and1 | f_arrdiv32_fs653_and0;
  assign f_arrdiv32_fs654_xor0 = f_arrdiv32_mux2to1602_xor0 ^ b[14];
  assign f_arrdiv32_fs654_not0 = ~f_arrdiv32_mux2to1602_xor0;
  assign f_arrdiv32_fs654_and0 = f_arrdiv32_fs654_not0 & b[14];
  assign f_arrdiv32_fs654_xor1 = f_arrdiv32_fs653_or0 ^ f_arrdiv32_fs654_xor0;
  assign f_arrdiv32_fs654_not1 = ~f_arrdiv32_fs654_xor0;
  assign f_arrdiv32_fs654_and1 = f_arrdiv32_fs654_not1 & f_arrdiv32_fs653_or0;
  assign f_arrdiv32_fs654_or0 = f_arrdiv32_fs654_and1 | f_arrdiv32_fs654_and0;
  assign f_arrdiv32_fs655_xor0 = f_arrdiv32_mux2to1603_xor0 ^ b[15];
  assign f_arrdiv32_fs655_not0 = ~f_arrdiv32_mux2to1603_xor0;
  assign f_arrdiv32_fs655_and0 = f_arrdiv32_fs655_not0 & b[15];
  assign f_arrdiv32_fs655_xor1 = f_arrdiv32_fs654_or0 ^ f_arrdiv32_fs655_xor0;
  assign f_arrdiv32_fs655_not1 = ~f_arrdiv32_fs655_xor0;
  assign f_arrdiv32_fs655_and1 = f_arrdiv32_fs655_not1 & f_arrdiv32_fs654_or0;
  assign f_arrdiv32_fs655_or0 = f_arrdiv32_fs655_and1 | f_arrdiv32_fs655_and0;
  assign f_arrdiv32_fs656_xor0 = f_arrdiv32_mux2to1604_xor0 ^ b[16];
  assign f_arrdiv32_fs656_not0 = ~f_arrdiv32_mux2to1604_xor0;
  assign f_arrdiv32_fs656_and0 = f_arrdiv32_fs656_not0 & b[16];
  assign f_arrdiv32_fs656_xor1 = f_arrdiv32_fs655_or0 ^ f_arrdiv32_fs656_xor0;
  assign f_arrdiv32_fs656_not1 = ~f_arrdiv32_fs656_xor0;
  assign f_arrdiv32_fs656_and1 = f_arrdiv32_fs656_not1 & f_arrdiv32_fs655_or0;
  assign f_arrdiv32_fs656_or0 = f_arrdiv32_fs656_and1 | f_arrdiv32_fs656_and0;
  assign f_arrdiv32_fs657_xor0 = f_arrdiv32_mux2to1605_xor0 ^ b[17];
  assign f_arrdiv32_fs657_not0 = ~f_arrdiv32_mux2to1605_xor0;
  assign f_arrdiv32_fs657_and0 = f_arrdiv32_fs657_not0 & b[17];
  assign f_arrdiv32_fs657_xor1 = f_arrdiv32_fs656_or0 ^ f_arrdiv32_fs657_xor0;
  assign f_arrdiv32_fs657_not1 = ~f_arrdiv32_fs657_xor0;
  assign f_arrdiv32_fs657_and1 = f_arrdiv32_fs657_not1 & f_arrdiv32_fs656_or0;
  assign f_arrdiv32_fs657_or0 = f_arrdiv32_fs657_and1 | f_arrdiv32_fs657_and0;
  assign f_arrdiv32_fs658_xor0 = f_arrdiv32_mux2to1606_xor0 ^ b[18];
  assign f_arrdiv32_fs658_not0 = ~f_arrdiv32_mux2to1606_xor0;
  assign f_arrdiv32_fs658_and0 = f_arrdiv32_fs658_not0 & b[18];
  assign f_arrdiv32_fs658_xor1 = f_arrdiv32_fs657_or0 ^ f_arrdiv32_fs658_xor0;
  assign f_arrdiv32_fs658_not1 = ~f_arrdiv32_fs658_xor0;
  assign f_arrdiv32_fs658_and1 = f_arrdiv32_fs658_not1 & f_arrdiv32_fs657_or0;
  assign f_arrdiv32_fs658_or0 = f_arrdiv32_fs658_and1 | f_arrdiv32_fs658_and0;
  assign f_arrdiv32_fs659_xor0 = f_arrdiv32_mux2to1607_xor0 ^ b[19];
  assign f_arrdiv32_fs659_not0 = ~f_arrdiv32_mux2to1607_xor0;
  assign f_arrdiv32_fs659_and0 = f_arrdiv32_fs659_not0 & b[19];
  assign f_arrdiv32_fs659_xor1 = f_arrdiv32_fs658_or0 ^ f_arrdiv32_fs659_xor0;
  assign f_arrdiv32_fs659_not1 = ~f_arrdiv32_fs659_xor0;
  assign f_arrdiv32_fs659_and1 = f_arrdiv32_fs659_not1 & f_arrdiv32_fs658_or0;
  assign f_arrdiv32_fs659_or0 = f_arrdiv32_fs659_and1 | f_arrdiv32_fs659_and0;
  assign f_arrdiv32_fs660_xor0 = f_arrdiv32_mux2to1608_xor0 ^ b[20];
  assign f_arrdiv32_fs660_not0 = ~f_arrdiv32_mux2to1608_xor0;
  assign f_arrdiv32_fs660_and0 = f_arrdiv32_fs660_not0 & b[20];
  assign f_arrdiv32_fs660_xor1 = f_arrdiv32_fs659_or0 ^ f_arrdiv32_fs660_xor0;
  assign f_arrdiv32_fs660_not1 = ~f_arrdiv32_fs660_xor0;
  assign f_arrdiv32_fs660_and1 = f_arrdiv32_fs660_not1 & f_arrdiv32_fs659_or0;
  assign f_arrdiv32_fs660_or0 = f_arrdiv32_fs660_and1 | f_arrdiv32_fs660_and0;
  assign f_arrdiv32_fs661_xor0 = f_arrdiv32_mux2to1609_xor0 ^ b[21];
  assign f_arrdiv32_fs661_not0 = ~f_arrdiv32_mux2to1609_xor0;
  assign f_arrdiv32_fs661_and0 = f_arrdiv32_fs661_not0 & b[21];
  assign f_arrdiv32_fs661_xor1 = f_arrdiv32_fs660_or0 ^ f_arrdiv32_fs661_xor0;
  assign f_arrdiv32_fs661_not1 = ~f_arrdiv32_fs661_xor0;
  assign f_arrdiv32_fs661_and1 = f_arrdiv32_fs661_not1 & f_arrdiv32_fs660_or0;
  assign f_arrdiv32_fs661_or0 = f_arrdiv32_fs661_and1 | f_arrdiv32_fs661_and0;
  assign f_arrdiv32_fs662_xor0 = f_arrdiv32_mux2to1610_xor0 ^ b[22];
  assign f_arrdiv32_fs662_not0 = ~f_arrdiv32_mux2to1610_xor0;
  assign f_arrdiv32_fs662_and0 = f_arrdiv32_fs662_not0 & b[22];
  assign f_arrdiv32_fs662_xor1 = f_arrdiv32_fs661_or0 ^ f_arrdiv32_fs662_xor0;
  assign f_arrdiv32_fs662_not1 = ~f_arrdiv32_fs662_xor0;
  assign f_arrdiv32_fs662_and1 = f_arrdiv32_fs662_not1 & f_arrdiv32_fs661_or0;
  assign f_arrdiv32_fs662_or0 = f_arrdiv32_fs662_and1 | f_arrdiv32_fs662_and0;
  assign f_arrdiv32_fs663_xor0 = f_arrdiv32_mux2to1611_xor0 ^ b[23];
  assign f_arrdiv32_fs663_not0 = ~f_arrdiv32_mux2to1611_xor0;
  assign f_arrdiv32_fs663_and0 = f_arrdiv32_fs663_not0 & b[23];
  assign f_arrdiv32_fs663_xor1 = f_arrdiv32_fs662_or0 ^ f_arrdiv32_fs663_xor0;
  assign f_arrdiv32_fs663_not1 = ~f_arrdiv32_fs663_xor0;
  assign f_arrdiv32_fs663_and1 = f_arrdiv32_fs663_not1 & f_arrdiv32_fs662_or0;
  assign f_arrdiv32_fs663_or0 = f_arrdiv32_fs663_and1 | f_arrdiv32_fs663_and0;
  assign f_arrdiv32_fs664_xor0 = f_arrdiv32_mux2to1612_xor0 ^ b[24];
  assign f_arrdiv32_fs664_not0 = ~f_arrdiv32_mux2to1612_xor0;
  assign f_arrdiv32_fs664_and0 = f_arrdiv32_fs664_not0 & b[24];
  assign f_arrdiv32_fs664_xor1 = f_arrdiv32_fs663_or0 ^ f_arrdiv32_fs664_xor0;
  assign f_arrdiv32_fs664_not1 = ~f_arrdiv32_fs664_xor0;
  assign f_arrdiv32_fs664_and1 = f_arrdiv32_fs664_not1 & f_arrdiv32_fs663_or0;
  assign f_arrdiv32_fs664_or0 = f_arrdiv32_fs664_and1 | f_arrdiv32_fs664_and0;
  assign f_arrdiv32_fs665_xor0 = f_arrdiv32_mux2to1613_xor0 ^ b[25];
  assign f_arrdiv32_fs665_not0 = ~f_arrdiv32_mux2to1613_xor0;
  assign f_arrdiv32_fs665_and0 = f_arrdiv32_fs665_not0 & b[25];
  assign f_arrdiv32_fs665_xor1 = f_arrdiv32_fs664_or0 ^ f_arrdiv32_fs665_xor0;
  assign f_arrdiv32_fs665_not1 = ~f_arrdiv32_fs665_xor0;
  assign f_arrdiv32_fs665_and1 = f_arrdiv32_fs665_not1 & f_arrdiv32_fs664_or0;
  assign f_arrdiv32_fs665_or0 = f_arrdiv32_fs665_and1 | f_arrdiv32_fs665_and0;
  assign f_arrdiv32_fs666_xor0 = f_arrdiv32_mux2to1614_xor0 ^ b[26];
  assign f_arrdiv32_fs666_not0 = ~f_arrdiv32_mux2to1614_xor0;
  assign f_arrdiv32_fs666_and0 = f_arrdiv32_fs666_not0 & b[26];
  assign f_arrdiv32_fs666_xor1 = f_arrdiv32_fs665_or0 ^ f_arrdiv32_fs666_xor0;
  assign f_arrdiv32_fs666_not1 = ~f_arrdiv32_fs666_xor0;
  assign f_arrdiv32_fs666_and1 = f_arrdiv32_fs666_not1 & f_arrdiv32_fs665_or0;
  assign f_arrdiv32_fs666_or0 = f_arrdiv32_fs666_and1 | f_arrdiv32_fs666_and0;
  assign f_arrdiv32_fs667_xor0 = f_arrdiv32_mux2to1615_xor0 ^ b[27];
  assign f_arrdiv32_fs667_not0 = ~f_arrdiv32_mux2to1615_xor0;
  assign f_arrdiv32_fs667_and0 = f_arrdiv32_fs667_not0 & b[27];
  assign f_arrdiv32_fs667_xor1 = f_arrdiv32_fs666_or0 ^ f_arrdiv32_fs667_xor0;
  assign f_arrdiv32_fs667_not1 = ~f_arrdiv32_fs667_xor0;
  assign f_arrdiv32_fs667_and1 = f_arrdiv32_fs667_not1 & f_arrdiv32_fs666_or0;
  assign f_arrdiv32_fs667_or0 = f_arrdiv32_fs667_and1 | f_arrdiv32_fs667_and0;
  assign f_arrdiv32_fs668_xor0 = f_arrdiv32_mux2to1616_xor0 ^ b[28];
  assign f_arrdiv32_fs668_not0 = ~f_arrdiv32_mux2to1616_xor0;
  assign f_arrdiv32_fs668_and0 = f_arrdiv32_fs668_not0 & b[28];
  assign f_arrdiv32_fs668_xor1 = f_arrdiv32_fs667_or0 ^ f_arrdiv32_fs668_xor0;
  assign f_arrdiv32_fs668_not1 = ~f_arrdiv32_fs668_xor0;
  assign f_arrdiv32_fs668_and1 = f_arrdiv32_fs668_not1 & f_arrdiv32_fs667_or0;
  assign f_arrdiv32_fs668_or0 = f_arrdiv32_fs668_and1 | f_arrdiv32_fs668_and0;
  assign f_arrdiv32_fs669_xor0 = f_arrdiv32_mux2to1617_xor0 ^ b[29];
  assign f_arrdiv32_fs669_not0 = ~f_arrdiv32_mux2to1617_xor0;
  assign f_arrdiv32_fs669_and0 = f_arrdiv32_fs669_not0 & b[29];
  assign f_arrdiv32_fs669_xor1 = f_arrdiv32_fs668_or0 ^ f_arrdiv32_fs669_xor0;
  assign f_arrdiv32_fs669_not1 = ~f_arrdiv32_fs669_xor0;
  assign f_arrdiv32_fs669_and1 = f_arrdiv32_fs669_not1 & f_arrdiv32_fs668_or0;
  assign f_arrdiv32_fs669_or0 = f_arrdiv32_fs669_and1 | f_arrdiv32_fs669_and0;
  assign f_arrdiv32_fs670_xor0 = f_arrdiv32_mux2to1618_xor0 ^ b[30];
  assign f_arrdiv32_fs670_not0 = ~f_arrdiv32_mux2to1618_xor0;
  assign f_arrdiv32_fs670_and0 = f_arrdiv32_fs670_not0 & b[30];
  assign f_arrdiv32_fs670_xor1 = f_arrdiv32_fs669_or0 ^ f_arrdiv32_fs670_xor0;
  assign f_arrdiv32_fs670_not1 = ~f_arrdiv32_fs670_xor0;
  assign f_arrdiv32_fs670_and1 = f_arrdiv32_fs670_not1 & f_arrdiv32_fs669_or0;
  assign f_arrdiv32_fs670_or0 = f_arrdiv32_fs670_and1 | f_arrdiv32_fs670_and0;
  assign f_arrdiv32_fs671_xor0 = f_arrdiv32_mux2to1619_xor0 ^ b[31];
  assign f_arrdiv32_fs671_not0 = ~f_arrdiv32_mux2to1619_xor0;
  assign f_arrdiv32_fs671_and0 = f_arrdiv32_fs671_not0 & b[31];
  assign f_arrdiv32_fs671_xor1 = f_arrdiv32_fs670_or0 ^ f_arrdiv32_fs671_xor0;
  assign f_arrdiv32_fs671_not1 = ~f_arrdiv32_fs671_xor0;
  assign f_arrdiv32_fs671_and1 = f_arrdiv32_fs671_not1 & f_arrdiv32_fs670_or0;
  assign f_arrdiv32_fs671_or0 = f_arrdiv32_fs671_and1 | f_arrdiv32_fs671_and0;
  assign f_arrdiv32_mux2to1620_and0 = a[11] & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1620_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1620_and1 = f_arrdiv32_fs640_xor0 & f_arrdiv32_mux2to1620_not0;
  assign f_arrdiv32_mux2to1620_xor0 = f_arrdiv32_mux2to1620_and0 ^ f_arrdiv32_mux2to1620_and1;
  assign f_arrdiv32_mux2to1621_and0 = f_arrdiv32_mux2to1589_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1621_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1621_and1 = f_arrdiv32_fs641_xor1 & f_arrdiv32_mux2to1621_not0;
  assign f_arrdiv32_mux2to1621_xor0 = f_arrdiv32_mux2to1621_and0 ^ f_arrdiv32_mux2to1621_and1;
  assign f_arrdiv32_mux2to1622_and0 = f_arrdiv32_mux2to1590_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1622_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1622_and1 = f_arrdiv32_fs642_xor1 & f_arrdiv32_mux2to1622_not0;
  assign f_arrdiv32_mux2to1622_xor0 = f_arrdiv32_mux2to1622_and0 ^ f_arrdiv32_mux2to1622_and1;
  assign f_arrdiv32_mux2to1623_and0 = f_arrdiv32_mux2to1591_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1623_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1623_and1 = f_arrdiv32_fs643_xor1 & f_arrdiv32_mux2to1623_not0;
  assign f_arrdiv32_mux2to1623_xor0 = f_arrdiv32_mux2to1623_and0 ^ f_arrdiv32_mux2to1623_and1;
  assign f_arrdiv32_mux2to1624_and0 = f_arrdiv32_mux2to1592_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1624_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1624_and1 = f_arrdiv32_fs644_xor1 & f_arrdiv32_mux2to1624_not0;
  assign f_arrdiv32_mux2to1624_xor0 = f_arrdiv32_mux2to1624_and0 ^ f_arrdiv32_mux2to1624_and1;
  assign f_arrdiv32_mux2to1625_and0 = f_arrdiv32_mux2to1593_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1625_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1625_and1 = f_arrdiv32_fs645_xor1 & f_arrdiv32_mux2to1625_not0;
  assign f_arrdiv32_mux2to1625_xor0 = f_arrdiv32_mux2to1625_and0 ^ f_arrdiv32_mux2to1625_and1;
  assign f_arrdiv32_mux2to1626_and0 = f_arrdiv32_mux2to1594_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1626_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1626_and1 = f_arrdiv32_fs646_xor1 & f_arrdiv32_mux2to1626_not0;
  assign f_arrdiv32_mux2to1626_xor0 = f_arrdiv32_mux2to1626_and0 ^ f_arrdiv32_mux2to1626_and1;
  assign f_arrdiv32_mux2to1627_and0 = f_arrdiv32_mux2to1595_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1627_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1627_and1 = f_arrdiv32_fs647_xor1 & f_arrdiv32_mux2to1627_not0;
  assign f_arrdiv32_mux2to1627_xor0 = f_arrdiv32_mux2to1627_and0 ^ f_arrdiv32_mux2to1627_and1;
  assign f_arrdiv32_mux2to1628_and0 = f_arrdiv32_mux2to1596_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1628_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1628_and1 = f_arrdiv32_fs648_xor1 & f_arrdiv32_mux2to1628_not0;
  assign f_arrdiv32_mux2to1628_xor0 = f_arrdiv32_mux2to1628_and0 ^ f_arrdiv32_mux2to1628_and1;
  assign f_arrdiv32_mux2to1629_and0 = f_arrdiv32_mux2to1597_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1629_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1629_and1 = f_arrdiv32_fs649_xor1 & f_arrdiv32_mux2to1629_not0;
  assign f_arrdiv32_mux2to1629_xor0 = f_arrdiv32_mux2to1629_and0 ^ f_arrdiv32_mux2to1629_and1;
  assign f_arrdiv32_mux2to1630_and0 = f_arrdiv32_mux2to1598_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1630_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1630_and1 = f_arrdiv32_fs650_xor1 & f_arrdiv32_mux2to1630_not0;
  assign f_arrdiv32_mux2to1630_xor0 = f_arrdiv32_mux2to1630_and0 ^ f_arrdiv32_mux2to1630_and1;
  assign f_arrdiv32_mux2to1631_and0 = f_arrdiv32_mux2to1599_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1631_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1631_and1 = f_arrdiv32_fs651_xor1 & f_arrdiv32_mux2to1631_not0;
  assign f_arrdiv32_mux2to1631_xor0 = f_arrdiv32_mux2to1631_and0 ^ f_arrdiv32_mux2to1631_and1;
  assign f_arrdiv32_mux2to1632_and0 = f_arrdiv32_mux2to1600_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1632_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1632_and1 = f_arrdiv32_fs652_xor1 & f_arrdiv32_mux2to1632_not0;
  assign f_arrdiv32_mux2to1632_xor0 = f_arrdiv32_mux2to1632_and0 ^ f_arrdiv32_mux2to1632_and1;
  assign f_arrdiv32_mux2to1633_and0 = f_arrdiv32_mux2to1601_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1633_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1633_and1 = f_arrdiv32_fs653_xor1 & f_arrdiv32_mux2to1633_not0;
  assign f_arrdiv32_mux2to1633_xor0 = f_arrdiv32_mux2to1633_and0 ^ f_arrdiv32_mux2to1633_and1;
  assign f_arrdiv32_mux2to1634_and0 = f_arrdiv32_mux2to1602_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1634_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1634_and1 = f_arrdiv32_fs654_xor1 & f_arrdiv32_mux2to1634_not0;
  assign f_arrdiv32_mux2to1634_xor0 = f_arrdiv32_mux2to1634_and0 ^ f_arrdiv32_mux2to1634_and1;
  assign f_arrdiv32_mux2to1635_and0 = f_arrdiv32_mux2to1603_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1635_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1635_and1 = f_arrdiv32_fs655_xor1 & f_arrdiv32_mux2to1635_not0;
  assign f_arrdiv32_mux2to1635_xor0 = f_arrdiv32_mux2to1635_and0 ^ f_arrdiv32_mux2to1635_and1;
  assign f_arrdiv32_mux2to1636_and0 = f_arrdiv32_mux2to1604_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1636_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1636_and1 = f_arrdiv32_fs656_xor1 & f_arrdiv32_mux2to1636_not0;
  assign f_arrdiv32_mux2to1636_xor0 = f_arrdiv32_mux2to1636_and0 ^ f_arrdiv32_mux2to1636_and1;
  assign f_arrdiv32_mux2to1637_and0 = f_arrdiv32_mux2to1605_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1637_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1637_and1 = f_arrdiv32_fs657_xor1 & f_arrdiv32_mux2to1637_not0;
  assign f_arrdiv32_mux2to1637_xor0 = f_arrdiv32_mux2to1637_and0 ^ f_arrdiv32_mux2to1637_and1;
  assign f_arrdiv32_mux2to1638_and0 = f_arrdiv32_mux2to1606_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1638_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1638_and1 = f_arrdiv32_fs658_xor1 & f_arrdiv32_mux2to1638_not0;
  assign f_arrdiv32_mux2to1638_xor0 = f_arrdiv32_mux2to1638_and0 ^ f_arrdiv32_mux2to1638_and1;
  assign f_arrdiv32_mux2to1639_and0 = f_arrdiv32_mux2to1607_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1639_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1639_and1 = f_arrdiv32_fs659_xor1 & f_arrdiv32_mux2to1639_not0;
  assign f_arrdiv32_mux2to1639_xor0 = f_arrdiv32_mux2to1639_and0 ^ f_arrdiv32_mux2to1639_and1;
  assign f_arrdiv32_mux2to1640_and0 = f_arrdiv32_mux2to1608_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1640_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1640_and1 = f_arrdiv32_fs660_xor1 & f_arrdiv32_mux2to1640_not0;
  assign f_arrdiv32_mux2to1640_xor0 = f_arrdiv32_mux2to1640_and0 ^ f_arrdiv32_mux2to1640_and1;
  assign f_arrdiv32_mux2to1641_and0 = f_arrdiv32_mux2to1609_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1641_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1641_and1 = f_arrdiv32_fs661_xor1 & f_arrdiv32_mux2to1641_not0;
  assign f_arrdiv32_mux2to1641_xor0 = f_arrdiv32_mux2to1641_and0 ^ f_arrdiv32_mux2to1641_and1;
  assign f_arrdiv32_mux2to1642_and0 = f_arrdiv32_mux2to1610_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1642_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1642_and1 = f_arrdiv32_fs662_xor1 & f_arrdiv32_mux2to1642_not0;
  assign f_arrdiv32_mux2to1642_xor0 = f_arrdiv32_mux2to1642_and0 ^ f_arrdiv32_mux2to1642_and1;
  assign f_arrdiv32_mux2to1643_and0 = f_arrdiv32_mux2to1611_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1643_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1643_and1 = f_arrdiv32_fs663_xor1 & f_arrdiv32_mux2to1643_not0;
  assign f_arrdiv32_mux2to1643_xor0 = f_arrdiv32_mux2to1643_and0 ^ f_arrdiv32_mux2to1643_and1;
  assign f_arrdiv32_mux2to1644_and0 = f_arrdiv32_mux2to1612_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1644_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1644_and1 = f_arrdiv32_fs664_xor1 & f_arrdiv32_mux2to1644_not0;
  assign f_arrdiv32_mux2to1644_xor0 = f_arrdiv32_mux2to1644_and0 ^ f_arrdiv32_mux2to1644_and1;
  assign f_arrdiv32_mux2to1645_and0 = f_arrdiv32_mux2to1613_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1645_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1645_and1 = f_arrdiv32_fs665_xor1 & f_arrdiv32_mux2to1645_not0;
  assign f_arrdiv32_mux2to1645_xor0 = f_arrdiv32_mux2to1645_and0 ^ f_arrdiv32_mux2to1645_and1;
  assign f_arrdiv32_mux2to1646_and0 = f_arrdiv32_mux2to1614_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1646_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1646_and1 = f_arrdiv32_fs666_xor1 & f_arrdiv32_mux2to1646_not0;
  assign f_arrdiv32_mux2to1646_xor0 = f_arrdiv32_mux2to1646_and0 ^ f_arrdiv32_mux2to1646_and1;
  assign f_arrdiv32_mux2to1647_and0 = f_arrdiv32_mux2to1615_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1647_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1647_and1 = f_arrdiv32_fs667_xor1 & f_arrdiv32_mux2to1647_not0;
  assign f_arrdiv32_mux2to1647_xor0 = f_arrdiv32_mux2to1647_and0 ^ f_arrdiv32_mux2to1647_and1;
  assign f_arrdiv32_mux2to1648_and0 = f_arrdiv32_mux2to1616_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1648_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1648_and1 = f_arrdiv32_fs668_xor1 & f_arrdiv32_mux2to1648_not0;
  assign f_arrdiv32_mux2to1648_xor0 = f_arrdiv32_mux2to1648_and0 ^ f_arrdiv32_mux2to1648_and1;
  assign f_arrdiv32_mux2to1649_and0 = f_arrdiv32_mux2to1617_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1649_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1649_and1 = f_arrdiv32_fs669_xor1 & f_arrdiv32_mux2to1649_not0;
  assign f_arrdiv32_mux2to1649_xor0 = f_arrdiv32_mux2to1649_and0 ^ f_arrdiv32_mux2to1649_and1;
  assign f_arrdiv32_mux2to1650_and0 = f_arrdiv32_mux2to1618_xor0 & f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1650_not0 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_mux2to1650_and1 = f_arrdiv32_fs670_xor1 & f_arrdiv32_mux2to1650_not0;
  assign f_arrdiv32_mux2to1650_xor0 = f_arrdiv32_mux2to1650_and0 ^ f_arrdiv32_mux2to1650_and1;
  assign f_arrdiv32_not20 = ~f_arrdiv32_fs671_or0;
  assign f_arrdiv32_fs672_xor0 = a[10] ^ b[0];
  assign f_arrdiv32_fs672_not0 = ~a[10];
  assign f_arrdiv32_fs672_and0 = f_arrdiv32_fs672_not0 & b[0];
  assign f_arrdiv32_fs672_not1 = ~f_arrdiv32_fs672_xor0;
  assign f_arrdiv32_fs673_xor0 = f_arrdiv32_mux2to1620_xor0 ^ b[1];
  assign f_arrdiv32_fs673_not0 = ~f_arrdiv32_mux2to1620_xor0;
  assign f_arrdiv32_fs673_and0 = f_arrdiv32_fs673_not0 & b[1];
  assign f_arrdiv32_fs673_xor1 = f_arrdiv32_fs672_and0 ^ f_arrdiv32_fs673_xor0;
  assign f_arrdiv32_fs673_not1 = ~f_arrdiv32_fs673_xor0;
  assign f_arrdiv32_fs673_and1 = f_arrdiv32_fs673_not1 & f_arrdiv32_fs672_and0;
  assign f_arrdiv32_fs673_or0 = f_arrdiv32_fs673_and1 | f_arrdiv32_fs673_and0;
  assign f_arrdiv32_fs674_xor0 = f_arrdiv32_mux2to1621_xor0 ^ b[2];
  assign f_arrdiv32_fs674_not0 = ~f_arrdiv32_mux2to1621_xor0;
  assign f_arrdiv32_fs674_and0 = f_arrdiv32_fs674_not0 & b[2];
  assign f_arrdiv32_fs674_xor1 = f_arrdiv32_fs673_or0 ^ f_arrdiv32_fs674_xor0;
  assign f_arrdiv32_fs674_not1 = ~f_arrdiv32_fs674_xor0;
  assign f_arrdiv32_fs674_and1 = f_arrdiv32_fs674_not1 & f_arrdiv32_fs673_or0;
  assign f_arrdiv32_fs674_or0 = f_arrdiv32_fs674_and1 | f_arrdiv32_fs674_and0;
  assign f_arrdiv32_fs675_xor0 = f_arrdiv32_mux2to1622_xor0 ^ b[3];
  assign f_arrdiv32_fs675_not0 = ~f_arrdiv32_mux2to1622_xor0;
  assign f_arrdiv32_fs675_and0 = f_arrdiv32_fs675_not0 & b[3];
  assign f_arrdiv32_fs675_xor1 = f_arrdiv32_fs674_or0 ^ f_arrdiv32_fs675_xor0;
  assign f_arrdiv32_fs675_not1 = ~f_arrdiv32_fs675_xor0;
  assign f_arrdiv32_fs675_and1 = f_arrdiv32_fs675_not1 & f_arrdiv32_fs674_or0;
  assign f_arrdiv32_fs675_or0 = f_arrdiv32_fs675_and1 | f_arrdiv32_fs675_and0;
  assign f_arrdiv32_fs676_xor0 = f_arrdiv32_mux2to1623_xor0 ^ b[4];
  assign f_arrdiv32_fs676_not0 = ~f_arrdiv32_mux2to1623_xor0;
  assign f_arrdiv32_fs676_and0 = f_arrdiv32_fs676_not0 & b[4];
  assign f_arrdiv32_fs676_xor1 = f_arrdiv32_fs675_or0 ^ f_arrdiv32_fs676_xor0;
  assign f_arrdiv32_fs676_not1 = ~f_arrdiv32_fs676_xor0;
  assign f_arrdiv32_fs676_and1 = f_arrdiv32_fs676_not1 & f_arrdiv32_fs675_or0;
  assign f_arrdiv32_fs676_or0 = f_arrdiv32_fs676_and1 | f_arrdiv32_fs676_and0;
  assign f_arrdiv32_fs677_xor0 = f_arrdiv32_mux2to1624_xor0 ^ b[5];
  assign f_arrdiv32_fs677_not0 = ~f_arrdiv32_mux2to1624_xor0;
  assign f_arrdiv32_fs677_and0 = f_arrdiv32_fs677_not0 & b[5];
  assign f_arrdiv32_fs677_xor1 = f_arrdiv32_fs676_or0 ^ f_arrdiv32_fs677_xor0;
  assign f_arrdiv32_fs677_not1 = ~f_arrdiv32_fs677_xor0;
  assign f_arrdiv32_fs677_and1 = f_arrdiv32_fs677_not1 & f_arrdiv32_fs676_or0;
  assign f_arrdiv32_fs677_or0 = f_arrdiv32_fs677_and1 | f_arrdiv32_fs677_and0;
  assign f_arrdiv32_fs678_xor0 = f_arrdiv32_mux2to1625_xor0 ^ b[6];
  assign f_arrdiv32_fs678_not0 = ~f_arrdiv32_mux2to1625_xor0;
  assign f_arrdiv32_fs678_and0 = f_arrdiv32_fs678_not0 & b[6];
  assign f_arrdiv32_fs678_xor1 = f_arrdiv32_fs677_or0 ^ f_arrdiv32_fs678_xor0;
  assign f_arrdiv32_fs678_not1 = ~f_arrdiv32_fs678_xor0;
  assign f_arrdiv32_fs678_and1 = f_arrdiv32_fs678_not1 & f_arrdiv32_fs677_or0;
  assign f_arrdiv32_fs678_or0 = f_arrdiv32_fs678_and1 | f_arrdiv32_fs678_and0;
  assign f_arrdiv32_fs679_xor0 = f_arrdiv32_mux2to1626_xor0 ^ b[7];
  assign f_arrdiv32_fs679_not0 = ~f_arrdiv32_mux2to1626_xor0;
  assign f_arrdiv32_fs679_and0 = f_arrdiv32_fs679_not0 & b[7];
  assign f_arrdiv32_fs679_xor1 = f_arrdiv32_fs678_or0 ^ f_arrdiv32_fs679_xor0;
  assign f_arrdiv32_fs679_not1 = ~f_arrdiv32_fs679_xor0;
  assign f_arrdiv32_fs679_and1 = f_arrdiv32_fs679_not1 & f_arrdiv32_fs678_or0;
  assign f_arrdiv32_fs679_or0 = f_arrdiv32_fs679_and1 | f_arrdiv32_fs679_and0;
  assign f_arrdiv32_fs680_xor0 = f_arrdiv32_mux2to1627_xor0 ^ b[8];
  assign f_arrdiv32_fs680_not0 = ~f_arrdiv32_mux2to1627_xor0;
  assign f_arrdiv32_fs680_and0 = f_arrdiv32_fs680_not0 & b[8];
  assign f_arrdiv32_fs680_xor1 = f_arrdiv32_fs679_or0 ^ f_arrdiv32_fs680_xor0;
  assign f_arrdiv32_fs680_not1 = ~f_arrdiv32_fs680_xor0;
  assign f_arrdiv32_fs680_and1 = f_arrdiv32_fs680_not1 & f_arrdiv32_fs679_or0;
  assign f_arrdiv32_fs680_or0 = f_arrdiv32_fs680_and1 | f_arrdiv32_fs680_and0;
  assign f_arrdiv32_fs681_xor0 = f_arrdiv32_mux2to1628_xor0 ^ b[9];
  assign f_arrdiv32_fs681_not0 = ~f_arrdiv32_mux2to1628_xor0;
  assign f_arrdiv32_fs681_and0 = f_arrdiv32_fs681_not0 & b[9];
  assign f_arrdiv32_fs681_xor1 = f_arrdiv32_fs680_or0 ^ f_arrdiv32_fs681_xor0;
  assign f_arrdiv32_fs681_not1 = ~f_arrdiv32_fs681_xor0;
  assign f_arrdiv32_fs681_and1 = f_arrdiv32_fs681_not1 & f_arrdiv32_fs680_or0;
  assign f_arrdiv32_fs681_or0 = f_arrdiv32_fs681_and1 | f_arrdiv32_fs681_and0;
  assign f_arrdiv32_fs682_xor0 = f_arrdiv32_mux2to1629_xor0 ^ b[10];
  assign f_arrdiv32_fs682_not0 = ~f_arrdiv32_mux2to1629_xor0;
  assign f_arrdiv32_fs682_and0 = f_arrdiv32_fs682_not0 & b[10];
  assign f_arrdiv32_fs682_xor1 = f_arrdiv32_fs681_or0 ^ f_arrdiv32_fs682_xor0;
  assign f_arrdiv32_fs682_not1 = ~f_arrdiv32_fs682_xor0;
  assign f_arrdiv32_fs682_and1 = f_arrdiv32_fs682_not1 & f_arrdiv32_fs681_or0;
  assign f_arrdiv32_fs682_or0 = f_arrdiv32_fs682_and1 | f_arrdiv32_fs682_and0;
  assign f_arrdiv32_fs683_xor0 = f_arrdiv32_mux2to1630_xor0 ^ b[11];
  assign f_arrdiv32_fs683_not0 = ~f_arrdiv32_mux2to1630_xor0;
  assign f_arrdiv32_fs683_and0 = f_arrdiv32_fs683_not0 & b[11];
  assign f_arrdiv32_fs683_xor1 = f_arrdiv32_fs682_or0 ^ f_arrdiv32_fs683_xor0;
  assign f_arrdiv32_fs683_not1 = ~f_arrdiv32_fs683_xor0;
  assign f_arrdiv32_fs683_and1 = f_arrdiv32_fs683_not1 & f_arrdiv32_fs682_or0;
  assign f_arrdiv32_fs683_or0 = f_arrdiv32_fs683_and1 | f_arrdiv32_fs683_and0;
  assign f_arrdiv32_fs684_xor0 = f_arrdiv32_mux2to1631_xor0 ^ b[12];
  assign f_arrdiv32_fs684_not0 = ~f_arrdiv32_mux2to1631_xor0;
  assign f_arrdiv32_fs684_and0 = f_arrdiv32_fs684_not0 & b[12];
  assign f_arrdiv32_fs684_xor1 = f_arrdiv32_fs683_or0 ^ f_arrdiv32_fs684_xor0;
  assign f_arrdiv32_fs684_not1 = ~f_arrdiv32_fs684_xor0;
  assign f_arrdiv32_fs684_and1 = f_arrdiv32_fs684_not1 & f_arrdiv32_fs683_or0;
  assign f_arrdiv32_fs684_or0 = f_arrdiv32_fs684_and1 | f_arrdiv32_fs684_and0;
  assign f_arrdiv32_fs685_xor0 = f_arrdiv32_mux2to1632_xor0 ^ b[13];
  assign f_arrdiv32_fs685_not0 = ~f_arrdiv32_mux2to1632_xor0;
  assign f_arrdiv32_fs685_and0 = f_arrdiv32_fs685_not0 & b[13];
  assign f_arrdiv32_fs685_xor1 = f_arrdiv32_fs684_or0 ^ f_arrdiv32_fs685_xor0;
  assign f_arrdiv32_fs685_not1 = ~f_arrdiv32_fs685_xor0;
  assign f_arrdiv32_fs685_and1 = f_arrdiv32_fs685_not1 & f_arrdiv32_fs684_or0;
  assign f_arrdiv32_fs685_or0 = f_arrdiv32_fs685_and1 | f_arrdiv32_fs685_and0;
  assign f_arrdiv32_fs686_xor0 = f_arrdiv32_mux2to1633_xor0 ^ b[14];
  assign f_arrdiv32_fs686_not0 = ~f_arrdiv32_mux2to1633_xor0;
  assign f_arrdiv32_fs686_and0 = f_arrdiv32_fs686_not0 & b[14];
  assign f_arrdiv32_fs686_xor1 = f_arrdiv32_fs685_or0 ^ f_arrdiv32_fs686_xor0;
  assign f_arrdiv32_fs686_not1 = ~f_arrdiv32_fs686_xor0;
  assign f_arrdiv32_fs686_and1 = f_arrdiv32_fs686_not1 & f_arrdiv32_fs685_or0;
  assign f_arrdiv32_fs686_or0 = f_arrdiv32_fs686_and1 | f_arrdiv32_fs686_and0;
  assign f_arrdiv32_fs687_xor0 = f_arrdiv32_mux2to1634_xor0 ^ b[15];
  assign f_arrdiv32_fs687_not0 = ~f_arrdiv32_mux2to1634_xor0;
  assign f_arrdiv32_fs687_and0 = f_arrdiv32_fs687_not0 & b[15];
  assign f_arrdiv32_fs687_xor1 = f_arrdiv32_fs686_or0 ^ f_arrdiv32_fs687_xor0;
  assign f_arrdiv32_fs687_not1 = ~f_arrdiv32_fs687_xor0;
  assign f_arrdiv32_fs687_and1 = f_arrdiv32_fs687_not1 & f_arrdiv32_fs686_or0;
  assign f_arrdiv32_fs687_or0 = f_arrdiv32_fs687_and1 | f_arrdiv32_fs687_and0;
  assign f_arrdiv32_fs688_xor0 = f_arrdiv32_mux2to1635_xor0 ^ b[16];
  assign f_arrdiv32_fs688_not0 = ~f_arrdiv32_mux2to1635_xor0;
  assign f_arrdiv32_fs688_and0 = f_arrdiv32_fs688_not0 & b[16];
  assign f_arrdiv32_fs688_xor1 = f_arrdiv32_fs687_or0 ^ f_arrdiv32_fs688_xor0;
  assign f_arrdiv32_fs688_not1 = ~f_arrdiv32_fs688_xor0;
  assign f_arrdiv32_fs688_and1 = f_arrdiv32_fs688_not1 & f_arrdiv32_fs687_or0;
  assign f_arrdiv32_fs688_or0 = f_arrdiv32_fs688_and1 | f_arrdiv32_fs688_and0;
  assign f_arrdiv32_fs689_xor0 = f_arrdiv32_mux2to1636_xor0 ^ b[17];
  assign f_arrdiv32_fs689_not0 = ~f_arrdiv32_mux2to1636_xor0;
  assign f_arrdiv32_fs689_and0 = f_arrdiv32_fs689_not0 & b[17];
  assign f_arrdiv32_fs689_xor1 = f_arrdiv32_fs688_or0 ^ f_arrdiv32_fs689_xor0;
  assign f_arrdiv32_fs689_not1 = ~f_arrdiv32_fs689_xor0;
  assign f_arrdiv32_fs689_and1 = f_arrdiv32_fs689_not1 & f_arrdiv32_fs688_or0;
  assign f_arrdiv32_fs689_or0 = f_arrdiv32_fs689_and1 | f_arrdiv32_fs689_and0;
  assign f_arrdiv32_fs690_xor0 = f_arrdiv32_mux2to1637_xor0 ^ b[18];
  assign f_arrdiv32_fs690_not0 = ~f_arrdiv32_mux2to1637_xor0;
  assign f_arrdiv32_fs690_and0 = f_arrdiv32_fs690_not0 & b[18];
  assign f_arrdiv32_fs690_xor1 = f_arrdiv32_fs689_or0 ^ f_arrdiv32_fs690_xor0;
  assign f_arrdiv32_fs690_not1 = ~f_arrdiv32_fs690_xor0;
  assign f_arrdiv32_fs690_and1 = f_arrdiv32_fs690_not1 & f_arrdiv32_fs689_or0;
  assign f_arrdiv32_fs690_or0 = f_arrdiv32_fs690_and1 | f_arrdiv32_fs690_and0;
  assign f_arrdiv32_fs691_xor0 = f_arrdiv32_mux2to1638_xor0 ^ b[19];
  assign f_arrdiv32_fs691_not0 = ~f_arrdiv32_mux2to1638_xor0;
  assign f_arrdiv32_fs691_and0 = f_arrdiv32_fs691_not0 & b[19];
  assign f_arrdiv32_fs691_xor1 = f_arrdiv32_fs690_or0 ^ f_arrdiv32_fs691_xor0;
  assign f_arrdiv32_fs691_not1 = ~f_arrdiv32_fs691_xor0;
  assign f_arrdiv32_fs691_and1 = f_arrdiv32_fs691_not1 & f_arrdiv32_fs690_or0;
  assign f_arrdiv32_fs691_or0 = f_arrdiv32_fs691_and1 | f_arrdiv32_fs691_and0;
  assign f_arrdiv32_fs692_xor0 = f_arrdiv32_mux2to1639_xor0 ^ b[20];
  assign f_arrdiv32_fs692_not0 = ~f_arrdiv32_mux2to1639_xor0;
  assign f_arrdiv32_fs692_and0 = f_arrdiv32_fs692_not0 & b[20];
  assign f_arrdiv32_fs692_xor1 = f_arrdiv32_fs691_or0 ^ f_arrdiv32_fs692_xor0;
  assign f_arrdiv32_fs692_not1 = ~f_arrdiv32_fs692_xor0;
  assign f_arrdiv32_fs692_and1 = f_arrdiv32_fs692_not1 & f_arrdiv32_fs691_or0;
  assign f_arrdiv32_fs692_or0 = f_arrdiv32_fs692_and1 | f_arrdiv32_fs692_and0;
  assign f_arrdiv32_fs693_xor0 = f_arrdiv32_mux2to1640_xor0 ^ b[21];
  assign f_arrdiv32_fs693_not0 = ~f_arrdiv32_mux2to1640_xor0;
  assign f_arrdiv32_fs693_and0 = f_arrdiv32_fs693_not0 & b[21];
  assign f_arrdiv32_fs693_xor1 = f_arrdiv32_fs692_or0 ^ f_arrdiv32_fs693_xor0;
  assign f_arrdiv32_fs693_not1 = ~f_arrdiv32_fs693_xor0;
  assign f_arrdiv32_fs693_and1 = f_arrdiv32_fs693_not1 & f_arrdiv32_fs692_or0;
  assign f_arrdiv32_fs693_or0 = f_arrdiv32_fs693_and1 | f_arrdiv32_fs693_and0;
  assign f_arrdiv32_fs694_xor0 = f_arrdiv32_mux2to1641_xor0 ^ b[22];
  assign f_arrdiv32_fs694_not0 = ~f_arrdiv32_mux2to1641_xor0;
  assign f_arrdiv32_fs694_and0 = f_arrdiv32_fs694_not0 & b[22];
  assign f_arrdiv32_fs694_xor1 = f_arrdiv32_fs693_or0 ^ f_arrdiv32_fs694_xor0;
  assign f_arrdiv32_fs694_not1 = ~f_arrdiv32_fs694_xor0;
  assign f_arrdiv32_fs694_and1 = f_arrdiv32_fs694_not1 & f_arrdiv32_fs693_or0;
  assign f_arrdiv32_fs694_or0 = f_arrdiv32_fs694_and1 | f_arrdiv32_fs694_and0;
  assign f_arrdiv32_fs695_xor0 = f_arrdiv32_mux2to1642_xor0 ^ b[23];
  assign f_arrdiv32_fs695_not0 = ~f_arrdiv32_mux2to1642_xor0;
  assign f_arrdiv32_fs695_and0 = f_arrdiv32_fs695_not0 & b[23];
  assign f_arrdiv32_fs695_xor1 = f_arrdiv32_fs694_or0 ^ f_arrdiv32_fs695_xor0;
  assign f_arrdiv32_fs695_not1 = ~f_arrdiv32_fs695_xor0;
  assign f_arrdiv32_fs695_and1 = f_arrdiv32_fs695_not1 & f_arrdiv32_fs694_or0;
  assign f_arrdiv32_fs695_or0 = f_arrdiv32_fs695_and1 | f_arrdiv32_fs695_and0;
  assign f_arrdiv32_fs696_xor0 = f_arrdiv32_mux2to1643_xor0 ^ b[24];
  assign f_arrdiv32_fs696_not0 = ~f_arrdiv32_mux2to1643_xor0;
  assign f_arrdiv32_fs696_and0 = f_arrdiv32_fs696_not0 & b[24];
  assign f_arrdiv32_fs696_xor1 = f_arrdiv32_fs695_or0 ^ f_arrdiv32_fs696_xor0;
  assign f_arrdiv32_fs696_not1 = ~f_arrdiv32_fs696_xor0;
  assign f_arrdiv32_fs696_and1 = f_arrdiv32_fs696_not1 & f_arrdiv32_fs695_or0;
  assign f_arrdiv32_fs696_or0 = f_arrdiv32_fs696_and1 | f_arrdiv32_fs696_and0;
  assign f_arrdiv32_fs697_xor0 = f_arrdiv32_mux2to1644_xor0 ^ b[25];
  assign f_arrdiv32_fs697_not0 = ~f_arrdiv32_mux2to1644_xor0;
  assign f_arrdiv32_fs697_and0 = f_arrdiv32_fs697_not0 & b[25];
  assign f_arrdiv32_fs697_xor1 = f_arrdiv32_fs696_or0 ^ f_arrdiv32_fs697_xor0;
  assign f_arrdiv32_fs697_not1 = ~f_arrdiv32_fs697_xor0;
  assign f_arrdiv32_fs697_and1 = f_arrdiv32_fs697_not1 & f_arrdiv32_fs696_or0;
  assign f_arrdiv32_fs697_or0 = f_arrdiv32_fs697_and1 | f_arrdiv32_fs697_and0;
  assign f_arrdiv32_fs698_xor0 = f_arrdiv32_mux2to1645_xor0 ^ b[26];
  assign f_arrdiv32_fs698_not0 = ~f_arrdiv32_mux2to1645_xor0;
  assign f_arrdiv32_fs698_and0 = f_arrdiv32_fs698_not0 & b[26];
  assign f_arrdiv32_fs698_xor1 = f_arrdiv32_fs697_or0 ^ f_arrdiv32_fs698_xor0;
  assign f_arrdiv32_fs698_not1 = ~f_arrdiv32_fs698_xor0;
  assign f_arrdiv32_fs698_and1 = f_arrdiv32_fs698_not1 & f_arrdiv32_fs697_or0;
  assign f_arrdiv32_fs698_or0 = f_arrdiv32_fs698_and1 | f_arrdiv32_fs698_and0;
  assign f_arrdiv32_fs699_xor0 = f_arrdiv32_mux2to1646_xor0 ^ b[27];
  assign f_arrdiv32_fs699_not0 = ~f_arrdiv32_mux2to1646_xor0;
  assign f_arrdiv32_fs699_and0 = f_arrdiv32_fs699_not0 & b[27];
  assign f_arrdiv32_fs699_xor1 = f_arrdiv32_fs698_or0 ^ f_arrdiv32_fs699_xor0;
  assign f_arrdiv32_fs699_not1 = ~f_arrdiv32_fs699_xor0;
  assign f_arrdiv32_fs699_and1 = f_arrdiv32_fs699_not1 & f_arrdiv32_fs698_or0;
  assign f_arrdiv32_fs699_or0 = f_arrdiv32_fs699_and1 | f_arrdiv32_fs699_and0;
  assign f_arrdiv32_fs700_xor0 = f_arrdiv32_mux2to1647_xor0 ^ b[28];
  assign f_arrdiv32_fs700_not0 = ~f_arrdiv32_mux2to1647_xor0;
  assign f_arrdiv32_fs700_and0 = f_arrdiv32_fs700_not0 & b[28];
  assign f_arrdiv32_fs700_xor1 = f_arrdiv32_fs699_or0 ^ f_arrdiv32_fs700_xor0;
  assign f_arrdiv32_fs700_not1 = ~f_arrdiv32_fs700_xor0;
  assign f_arrdiv32_fs700_and1 = f_arrdiv32_fs700_not1 & f_arrdiv32_fs699_or0;
  assign f_arrdiv32_fs700_or0 = f_arrdiv32_fs700_and1 | f_arrdiv32_fs700_and0;
  assign f_arrdiv32_fs701_xor0 = f_arrdiv32_mux2to1648_xor0 ^ b[29];
  assign f_arrdiv32_fs701_not0 = ~f_arrdiv32_mux2to1648_xor0;
  assign f_arrdiv32_fs701_and0 = f_arrdiv32_fs701_not0 & b[29];
  assign f_arrdiv32_fs701_xor1 = f_arrdiv32_fs700_or0 ^ f_arrdiv32_fs701_xor0;
  assign f_arrdiv32_fs701_not1 = ~f_arrdiv32_fs701_xor0;
  assign f_arrdiv32_fs701_and1 = f_arrdiv32_fs701_not1 & f_arrdiv32_fs700_or0;
  assign f_arrdiv32_fs701_or0 = f_arrdiv32_fs701_and1 | f_arrdiv32_fs701_and0;
  assign f_arrdiv32_fs702_xor0 = f_arrdiv32_mux2to1649_xor0 ^ b[30];
  assign f_arrdiv32_fs702_not0 = ~f_arrdiv32_mux2to1649_xor0;
  assign f_arrdiv32_fs702_and0 = f_arrdiv32_fs702_not0 & b[30];
  assign f_arrdiv32_fs702_xor1 = f_arrdiv32_fs701_or0 ^ f_arrdiv32_fs702_xor0;
  assign f_arrdiv32_fs702_not1 = ~f_arrdiv32_fs702_xor0;
  assign f_arrdiv32_fs702_and1 = f_arrdiv32_fs702_not1 & f_arrdiv32_fs701_or0;
  assign f_arrdiv32_fs702_or0 = f_arrdiv32_fs702_and1 | f_arrdiv32_fs702_and0;
  assign f_arrdiv32_fs703_xor0 = f_arrdiv32_mux2to1650_xor0 ^ b[31];
  assign f_arrdiv32_fs703_not0 = ~f_arrdiv32_mux2to1650_xor0;
  assign f_arrdiv32_fs703_and0 = f_arrdiv32_fs703_not0 & b[31];
  assign f_arrdiv32_fs703_xor1 = f_arrdiv32_fs702_or0 ^ f_arrdiv32_fs703_xor0;
  assign f_arrdiv32_fs703_not1 = ~f_arrdiv32_fs703_xor0;
  assign f_arrdiv32_fs703_and1 = f_arrdiv32_fs703_not1 & f_arrdiv32_fs702_or0;
  assign f_arrdiv32_fs703_or0 = f_arrdiv32_fs703_and1 | f_arrdiv32_fs703_and0;
  assign f_arrdiv32_mux2to1651_and0 = a[10] & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1651_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1651_and1 = f_arrdiv32_fs672_xor0 & f_arrdiv32_mux2to1651_not0;
  assign f_arrdiv32_mux2to1651_xor0 = f_arrdiv32_mux2to1651_and0 ^ f_arrdiv32_mux2to1651_and1;
  assign f_arrdiv32_mux2to1652_and0 = f_arrdiv32_mux2to1620_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1652_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1652_and1 = f_arrdiv32_fs673_xor1 & f_arrdiv32_mux2to1652_not0;
  assign f_arrdiv32_mux2to1652_xor0 = f_arrdiv32_mux2to1652_and0 ^ f_arrdiv32_mux2to1652_and1;
  assign f_arrdiv32_mux2to1653_and0 = f_arrdiv32_mux2to1621_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1653_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1653_and1 = f_arrdiv32_fs674_xor1 & f_arrdiv32_mux2to1653_not0;
  assign f_arrdiv32_mux2to1653_xor0 = f_arrdiv32_mux2to1653_and0 ^ f_arrdiv32_mux2to1653_and1;
  assign f_arrdiv32_mux2to1654_and0 = f_arrdiv32_mux2to1622_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1654_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1654_and1 = f_arrdiv32_fs675_xor1 & f_arrdiv32_mux2to1654_not0;
  assign f_arrdiv32_mux2to1654_xor0 = f_arrdiv32_mux2to1654_and0 ^ f_arrdiv32_mux2to1654_and1;
  assign f_arrdiv32_mux2to1655_and0 = f_arrdiv32_mux2to1623_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1655_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1655_and1 = f_arrdiv32_fs676_xor1 & f_arrdiv32_mux2to1655_not0;
  assign f_arrdiv32_mux2to1655_xor0 = f_arrdiv32_mux2to1655_and0 ^ f_arrdiv32_mux2to1655_and1;
  assign f_arrdiv32_mux2to1656_and0 = f_arrdiv32_mux2to1624_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1656_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1656_and1 = f_arrdiv32_fs677_xor1 & f_arrdiv32_mux2to1656_not0;
  assign f_arrdiv32_mux2to1656_xor0 = f_arrdiv32_mux2to1656_and0 ^ f_arrdiv32_mux2to1656_and1;
  assign f_arrdiv32_mux2to1657_and0 = f_arrdiv32_mux2to1625_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1657_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1657_and1 = f_arrdiv32_fs678_xor1 & f_arrdiv32_mux2to1657_not0;
  assign f_arrdiv32_mux2to1657_xor0 = f_arrdiv32_mux2to1657_and0 ^ f_arrdiv32_mux2to1657_and1;
  assign f_arrdiv32_mux2to1658_and0 = f_arrdiv32_mux2to1626_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1658_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1658_and1 = f_arrdiv32_fs679_xor1 & f_arrdiv32_mux2to1658_not0;
  assign f_arrdiv32_mux2to1658_xor0 = f_arrdiv32_mux2to1658_and0 ^ f_arrdiv32_mux2to1658_and1;
  assign f_arrdiv32_mux2to1659_and0 = f_arrdiv32_mux2to1627_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1659_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1659_and1 = f_arrdiv32_fs680_xor1 & f_arrdiv32_mux2to1659_not0;
  assign f_arrdiv32_mux2to1659_xor0 = f_arrdiv32_mux2to1659_and0 ^ f_arrdiv32_mux2to1659_and1;
  assign f_arrdiv32_mux2to1660_and0 = f_arrdiv32_mux2to1628_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1660_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1660_and1 = f_arrdiv32_fs681_xor1 & f_arrdiv32_mux2to1660_not0;
  assign f_arrdiv32_mux2to1660_xor0 = f_arrdiv32_mux2to1660_and0 ^ f_arrdiv32_mux2to1660_and1;
  assign f_arrdiv32_mux2to1661_and0 = f_arrdiv32_mux2to1629_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1661_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1661_and1 = f_arrdiv32_fs682_xor1 & f_arrdiv32_mux2to1661_not0;
  assign f_arrdiv32_mux2to1661_xor0 = f_arrdiv32_mux2to1661_and0 ^ f_arrdiv32_mux2to1661_and1;
  assign f_arrdiv32_mux2to1662_and0 = f_arrdiv32_mux2to1630_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1662_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1662_and1 = f_arrdiv32_fs683_xor1 & f_arrdiv32_mux2to1662_not0;
  assign f_arrdiv32_mux2to1662_xor0 = f_arrdiv32_mux2to1662_and0 ^ f_arrdiv32_mux2to1662_and1;
  assign f_arrdiv32_mux2to1663_and0 = f_arrdiv32_mux2to1631_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1663_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1663_and1 = f_arrdiv32_fs684_xor1 & f_arrdiv32_mux2to1663_not0;
  assign f_arrdiv32_mux2to1663_xor0 = f_arrdiv32_mux2to1663_and0 ^ f_arrdiv32_mux2to1663_and1;
  assign f_arrdiv32_mux2to1664_and0 = f_arrdiv32_mux2to1632_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1664_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1664_and1 = f_arrdiv32_fs685_xor1 & f_arrdiv32_mux2to1664_not0;
  assign f_arrdiv32_mux2to1664_xor0 = f_arrdiv32_mux2to1664_and0 ^ f_arrdiv32_mux2to1664_and1;
  assign f_arrdiv32_mux2to1665_and0 = f_arrdiv32_mux2to1633_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1665_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1665_and1 = f_arrdiv32_fs686_xor1 & f_arrdiv32_mux2to1665_not0;
  assign f_arrdiv32_mux2to1665_xor0 = f_arrdiv32_mux2to1665_and0 ^ f_arrdiv32_mux2to1665_and1;
  assign f_arrdiv32_mux2to1666_and0 = f_arrdiv32_mux2to1634_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1666_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1666_and1 = f_arrdiv32_fs687_xor1 & f_arrdiv32_mux2to1666_not0;
  assign f_arrdiv32_mux2to1666_xor0 = f_arrdiv32_mux2to1666_and0 ^ f_arrdiv32_mux2to1666_and1;
  assign f_arrdiv32_mux2to1667_and0 = f_arrdiv32_mux2to1635_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1667_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1667_and1 = f_arrdiv32_fs688_xor1 & f_arrdiv32_mux2to1667_not0;
  assign f_arrdiv32_mux2to1667_xor0 = f_arrdiv32_mux2to1667_and0 ^ f_arrdiv32_mux2to1667_and1;
  assign f_arrdiv32_mux2to1668_and0 = f_arrdiv32_mux2to1636_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1668_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1668_and1 = f_arrdiv32_fs689_xor1 & f_arrdiv32_mux2to1668_not0;
  assign f_arrdiv32_mux2to1668_xor0 = f_arrdiv32_mux2to1668_and0 ^ f_arrdiv32_mux2to1668_and1;
  assign f_arrdiv32_mux2to1669_and0 = f_arrdiv32_mux2to1637_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1669_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1669_and1 = f_arrdiv32_fs690_xor1 & f_arrdiv32_mux2to1669_not0;
  assign f_arrdiv32_mux2to1669_xor0 = f_arrdiv32_mux2to1669_and0 ^ f_arrdiv32_mux2to1669_and1;
  assign f_arrdiv32_mux2to1670_and0 = f_arrdiv32_mux2to1638_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1670_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1670_and1 = f_arrdiv32_fs691_xor1 & f_arrdiv32_mux2to1670_not0;
  assign f_arrdiv32_mux2to1670_xor0 = f_arrdiv32_mux2to1670_and0 ^ f_arrdiv32_mux2to1670_and1;
  assign f_arrdiv32_mux2to1671_and0 = f_arrdiv32_mux2to1639_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1671_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1671_and1 = f_arrdiv32_fs692_xor1 & f_arrdiv32_mux2to1671_not0;
  assign f_arrdiv32_mux2to1671_xor0 = f_arrdiv32_mux2to1671_and0 ^ f_arrdiv32_mux2to1671_and1;
  assign f_arrdiv32_mux2to1672_and0 = f_arrdiv32_mux2to1640_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1672_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1672_and1 = f_arrdiv32_fs693_xor1 & f_arrdiv32_mux2to1672_not0;
  assign f_arrdiv32_mux2to1672_xor0 = f_arrdiv32_mux2to1672_and0 ^ f_arrdiv32_mux2to1672_and1;
  assign f_arrdiv32_mux2to1673_and0 = f_arrdiv32_mux2to1641_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1673_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1673_and1 = f_arrdiv32_fs694_xor1 & f_arrdiv32_mux2to1673_not0;
  assign f_arrdiv32_mux2to1673_xor0 = f_arrdiv32_mux2to1673_and0 ^ f_arrdiv32_mux2to1673_and1;
  assign f_arrdiv32_mux2to1674_and0 = f_arrdiv32_mux2to1642_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1674_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1674_and1 = f_arrdiv32_fs695_xor1 & f_arrdiv32_mux2to1674_not0;
  assign f_arrdiv32_mux2to1674_xor0 = f_arrdiv32_mux2to1674_and0 ^ f_arrdiv32_mux2to1674_and1;
  assign f_arrdiv32_mux2to1675_and0 = f_arrdiv32_mux2to1643_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1675_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1675_and1 = f_arrdiv32_fs696_xor1 & f_arrdiv32_mux2to1675_not0;
  assign f_arrdiv32_mux2to1675_xor0 = f_arrdiv32_mux2to1675_and0 ^ f_arrdiv32_mux2to1675_and1;
  assign f_arrdiv32_mux2to1676_and0 = f_arrdiv32_mux2to1644_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1676_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1676_and1 = f_arrdiv32_fs697_xor1 & f_arrdiv32_mux2to1676_not0;
  assign f_arrdiv32_mux2to1676_xor0 = f_arrdiv32_mux2to1676_and0 ^ f_arrdiv32_mux2to1676_and1;
  assign f_arrdiv32_mux2to1677_and0 = f_arrdiv32_mux2to1645_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1677_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1677_and1 = f_arrdiv32_fs698_xor1 & f_arrdiv32_mux2to1677_not0;
  assign f_arrdiv32_mux2to1677_xor0 = f_arrdiv32_mux2to1677_and0 ^ f_arrdiv32_mux2to1677_and1;
  assign f_arrdiv32_mux2to1678_and0 = f_arrdiv32_mux2to1646_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1678_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1678_and1 = f_arrdiv32_fs699_xor1 & f_arrdiv32_mux2to1678_not0;
  assign f_arrdiv32_mux2to1678_xor0 = f_arrdiv32_mux2to1678_and0 ^ f_arrdiv32_mux2to1678_and1;
  assign f_arrdiv32_mux2to1679_and0 = f_arrdiv32_mux2to1647_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1679_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1679_and1 = f_arrdiv32_fs700_xor1 & f_arrdiv32_mux2to1679_not0;
  assign f_arrdiv32_mux2to1679_xor0 = f_arrdiv32_mux2to1679_and0 ^ f_arrdiv32_mux2to1679_and1;
  assign f_arrdiv32_mux2to1680_and0 = f_arrdiv32_mux2to1648_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1680_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1680_and1 = f_arrdiv32_fs701_xor1 & f_arrdiv32_mux2to1680_not0;
  assign f_arrdiv32_mux2to1680_xor0 = f_arrdiv32_mux2to1680_and0 ^ f_arrdiv32_mux2to1680_and1;
  assign f_arrdiv32_mux2to1681_and0 = f_arrdiv32_mux2to1649_xor0 & f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1681_not0 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_mux2to1681_and1 = f_arrdiv32_fs702_xor1 & f_arrdiv32_mux2to1681_not0;
  assign f_arrdiv32_mux2to1681_xor0 = f_arrdiv32_mux2to1681_and0 ^ f_arrdiv32_mux2to1681_and1;
  assign f_arrdiv32_not21 = ~f_arrdiv32_fs703_or0;
  assign f_arrdiv32_fs704_xor0 = a[9] ^ b[0];
  assign f_arrdiv32_fs704_not0 = ~a[9];
  assign f_arrdiv32_fs704_and0 = f_arrdiv32_fs704_not0 & b[0];
  assign f_arrdiv32_fs704_not1 = ~f_arrdiv32_fs704_xor0;
  assign f_arrdiv32_fs705_xor0 = f_arrdiv32_mux2to1651_xor0 ^ b[1];
  assign f_arrdiv32_fs705_not0 = ~f_arrdiv32_mux2to1651_xor0;
  assign f_arrdiv32_fs705_and0 = f_arrdiv32_fs705_not0 & b[1];
  assign f_arrdiv32_fs705_xor1 = f_arrdiv32_fs704_and0 ^ f_arrdiv32_fs705_xor0;
  assign f_arrdiv32_fs705_not1 = ~f_arrdiv32_fs705_xor0;
  assign f_arrdiv32_fs705_and1 = f_arrdiv32_fs705_not1 & f_arrdiv32_fs704_and0;
  assign f_arrdiv32_fs705_or0 = f_arrdiv32_fs705_and1 | f_arrdiv32_fs705_and0;
  assign f_arrdiv32_fs706_xor0 = f_arrdiv32_mux2to1652_xor0 ^ b[2];
  assign f_arrdiv32_fs706_not0 = ~f_arrdiv32_mux2to1652_xor0;
  assign f_arrdiv32_fs706_and0 = f_arrdiv32_fs706_not0 & b[2];
  assign f_arrdiv32_fs706_xor1 = f_arrdiv32_fs705_or0 ^ f_arrdiv32_fs706_xor0;
  assign f_arrdiv32_fs706_not1 = ~f_arrdiv32_fs706_xor0;
  assign f_arrdiv32_fs706_and1 = f_arrdiv32_fs706_not1 & f_arrdiv32_fs705_or0;
  assign f_arrdiv32_fs706_or0 = f_arrdiv32_fs706_and1 | f_arrdiv32_fs706_and0;
  assign f_arrdiv32_fs707_xor0 = f_arrdiv32_mux2to1653_xor0 ^ b[3];
  assign f_arrdiv32_fs707_not0 = ~f_arrdiv32_mux2to1653_xor0;
  assign f_arrdiv32_fs707_and0 = f_arrdiv32_fs707_not0 & b[3];
  assign f_arrdiv32_fs707_xor1 = f_arrdiv32_fs706_or0 ^ f_arrdiv32_fs707_xor0;
  assign f_arrdiv32_fs707_not1 = ~f_arrdiv32_fs707_xor0;
  assign f_arrdiv32_fs707_and1 = f_arrdiv32_fs707_not1 & f_arrdiv32_fs706_or0;
  assign f_arrdiv32_fs707_or0 = f_arrdiv32_fs707_and1 | f_arrdiv32_fs707_and0;
  assign f_arrdiv32_fs708_xor0 = f_arrdiv32_mux2to1654_xor0 ^ b[4];
  assign f_arrdiv32_fs708_not0 = ~f_arrdiv32_mux2to1654_xor0;
  assign f_arrdiv32_fs708_and0 = f_arrdiv32_fs708_not0 & b[4];
  assign f_arrdiv32_fs708_xor1 = f_arrdiv32_fs707_or0 ^ f_arrdiv32_fs708_xor0;
  assign f_arrdiv32_fs708_not1 = ~f_arrdiv32_fs708_xor0;
  assign f_arrdiv32_fs708_and1 = f_arrdiv32_fs708_not1 & f_arrdiv32_fs707_or0;
  assign f_arrdiv32_fs708_or0 = f_arrdiv32_fs708_and1 | f_arrdiv32_fs708_and0;
  assign f_arrdiv32_fs709_xor0 = f_arrdiv32_mux2to1655_xor0 ^ b[5];
  assign f_arrdiv32_fs709_not0 = ~f_arrdiv32_mux2to1655_xor0;
  assign f_arrdiv32_fs709_and0 = f_arrdiv32_fs709_not0 & b[5];
  assign f_arrdiv32_fs709_xor1 = f_arrdiv32_fs708_or0 ^ f_arrdiv32_fs709_xor0;
  assign f_arrdiv32_fs709_not1 = ~f_arrdiv32_fs709_xor0;
  assign f_arrdiv32_fs709_and1 = f_arrdiv32_fs709_not1 & f_arrdiv32_fs708_or0;
  assign f_arrdiv32_fs709_or0 = f_arrdiv32_fs709_and1 | f_arrdiv32_fs709_and0;
  assign f_arrdiv32_fs710_xor0 = f_arrdiv32_mux2to1656_xor0 ^ b[6];
  assign f_arrdiv32_fs710_not0 = ~f_arrdiv32_mux2to1656_xor0;
  assign f_arrdiv32_fs710_and0 = f_arrdiv32_fs710_not0 & b[6];
  assign f_arrdiv32_fs710_xor1 = f_arrdiv32_fs709_or0 ^ f_arrdiv32_fs710_xor0;
  assign f_arrdiv32_fs710_not1 = ~f_arrdiv32_fs710_xor0;
  assign f_arrdiv32_fs710_and1 = f_arrdiv32_fs710_not1 & f_arrdiv32_fs709_or0;
  assign f_arrdiv32_fs710_or0 = f_arrdiv32_fs710_and1 | f_arrdiv32_fs710_and0;
  assign f_arrdiv32_fs711_xor0 = f_arrdiv32_mux2to1657_xor0 ^ b[7];
  assign f_arrdiv32_fs711_not0 = ~f_arrdiv32_mux2to1657_xor0;
  assign f_arrdiv32_fs711_and0 = f_arrdiv32_fs711_not0 & b[7];
  assign f_arrdiv32_fs711_xor1 = f_arrdiv32_fs710_or0 ^ f_arrdiv32_fs711_xor0;
  assign f_arrdiv32_fs711_not1 = ~f_arrdiv32_fs711_xor0;
  assign f_arrdiv32_fs711_and1 = f_arrdiv32_fs711_not1 & f_arrdiv32_fs710_or0;
  assign f_arrdiv32_fs711_or0 = f_arrdiv32_fs711_and1 | f_arrdiv32_fs711_and0;
  assign f_arrdiv32_fs712_xor0 = f_arrdiv32_mux2to1658_xor0 ^ b[8];
  assign f_arrdiv32_fs712_not0 = ~f_arrdiv32_mux2to1658_xor0;
  assign f_arrdiv32_fs712_and0 = f_arrdiv32_fs712_not0 & b[8];
  assign f_arrdiv32_fs712_xor1 = f_arrdiv32_fs711_or0 ^ f_arrdiv32_fs712_xor0;
  assign f_arrdiv32_fs712_not1 = ~f_arrdiv32_fs712_xor0;
  assign f_arrdiv32_fs712_and1 = f_arrdiv32_fs712_not1 & f_arrdiv32_fs711_or0;
  assign f_arrdiv32_fs712_or0 = f_arrdiv32_fs712_and1 | f_arrdiv32_fs712_and0;
  assign f_arrdiv32_fs713_xor0 = f_arrdiv32_mux2to1659_xor0 ^ b[9];
  assign f_arrdiv32_fs713_not0 = ~f_arrdiv32_mux2to1659_xor0;
  assign f_arrdiv32_fs713_and0 = f_arrdiv32_fs713_not0 & b[9];
  assign f_arrdiv32_fs713_xor1 = f_arrdiv32_fs712_or0 ^ f_arrdiv32_fs713_xor0;
  assign f_arrdiv32_fs713_not1 = ~f_arrdiv32_fs713_xor0;
  assign f_arrdiv32_fs713_and1 = f_arrdiv32_fs713_not1 & f_arrdiv32_fs712_or0;
  assign f_arrdiv32_fs713_or0 = f_arrdiv32_fs713_and1 | f_arrdiv32_fs713_and0;
  assign f_arrdiv32_fs714_xor0 = f_arrdiv32_mux2to1660_xor0 ^ b[10];
  assign f_arrdiv32_fs714_not0 = ~f_arrdiv32_mux2to1660_xor0;
  assign f_arrdiv32_fs714_and0 = f_arrdiv32_fs714_not0 & b[10];
  assign f_arrdiv32_fs714_xor1 = f_arrdiv32_fs713_or0 ^ f_arrdiv32_fs714_xor0;
  assign f_arrdiv32_fs714_not1 = ~f_arrdiv32_fs714_xor0;
  assign f_arrdiv32_fs714_and1 = f_arrdiv32_fs714_not1 & f_arrdiv32_fs713_or0;
  assign f_arrdiv32_fs714_or0 = f_arrdiv32_fs714_and1 | f_arrdiv32_fs714_and0;
  assign f_arrdiv32_fs715_xor0 = f_arrdiv32_mux2to1661_xor0 ^ b[11];
  assign f_arrdiv32_fs715_not0 = ~f_arrdiv32_mux2to1661_xor0;
  assign f_arrdiv32_fs715_and0 = f_arrdiv32_fs715_not0 & b[11];
  assign f_arrdiv32_fs715_xor1 = f_arrdiv32_fs714_or0 ^ f_arrdiv32_fs715_xor0;
  assign f_arrdiv32_fs715_not1 = ~f_arrdiv32_fs715_xor0;
  assign f_arrdiv32_fs715_and1 = f_arrdiv32_fs715_not1 & f_arrdiv32_fs714_or0;
  assign f_arrdiv32_fs715_or0 = f_arrdiv32_fs715_and1 | f_arrdiv32_fs715_and0;
  assign f_arrdiv32_fs716_xor0 = f_arrdiv32_mux2to1662_xor0 ^ b[12];
  assign f_arrdiv32_fs716_not0 = ~f_arrdiv32_mux2to1662_xor0;
  assign f_arrdiv32_fs716_and0 = f_arrdiv32_fs716_not0 & b[12];
  assign f_arrdiv32_fs716_xor1 = f_arrdiv32_fs715_or0 ^ f_arrdiv32_fs716_xor0;
  assign f_arrdiv32_fs716_not1 = ~f_arrdiv32_fs716_xor0;
  assign f_arrdiv32_fs716_and1 = f_arrdiv32_fs716_not1 & f_arrdiv32_fs715_or0;
  assign f_arrdiv32_fs716_or0 = f_arrdiv32_fs716_and1 | f_arrdiv32_fs716_and0;
  assign f_arrdiv32_fs717_xor0 = f_arrdiv32_mux2to1663_xor0 ^ b[13];
  assign f_arrdiv32_fs717_not0 = ~f_arrdiv32_mux2to1663_xor0;
  assign f_arrdiv32_fs717_and0 = f_arrdiv32_fs717_not0 & b[13];
  assign f_arrdiv32_fs717_xor1 = f_arrdiv32_fs716_or0 ^ f_arrdiv32_fs717_xor0;
  assign f_arrdiv32_fs717_not1 = ~f_arrdiv32_fs717_xor0;
  assign f_arrdiv32_fs717_and1 = f_arrdiv32_fs717_not1 & f_arrdiv32_fs716_or0;
  assign f_arrdiv32_fs717_or0 = f_arrdiv32_fs717_and1 | f_arrdiv32_fs717_and0;
  assign f_arrdiv32_fs718_xor0 = f_arrdiv32_mux2to1664_xor0 ^ b[14];
  assign f_arrdiv32_fs718_not0 = ~f_arrdiv32_mux2to1664_xor0;
  assign f_arrdiv32_fs718_and0 = f_arrdiv32_fs718_not0 & b[14];
  assign f_arrdiv32_fs718_xor1 = f_arrdiv32_fs717_or0 ^ f_arrdiv32_fs718_xor0;
  assign f_arrdiv32_fs718_not1 = ~f_arrdiv32_fs718_xor0;
  assign f_arrdiv32_fs718_and1 = f_arrdiv32_fs718_not1 & f_arrdiv32_fs717_or0;
  assign f_arrdiv32_fs718_or0 = f_arrdiv32_fs718_and1 | f_arrdiv32_fs718_and0;
  assign f_arrdiv32_fs719_xor0 = f_arrdiv32_mux2to1665_xor0 ^ b[15];
  assign f_arrdiv32_fs719_not0 = ~f_arrdiv32_mux2to1665_xor0;
  assign f_arrdiv32_fs719_and0 = f_arrdiv32_fs719_not0 & b[15];
  assign f_arrdiv32_fs719_xor1 = f_arrdiv32_fs718_or0 ^ f_arrdiv32_fs719_xor0;
  assign f_arrdiv32_fs719_not1 = ~f_arrdiv32_fs719_xor0;
  assign f_arrdiv32_fs719_and1 = f_arrdiv32_fs719_not1 & f_arrdiv32_fs718_or0;
  assign f_arrdiv32_fs719_or0 = f_arrdiv32_fs719_and1 | f_arrdiv32_fs719_and0;
  assign f_arrdiv32_fs720_xor0 = f_arrdiv32_mux2to1666_xor0 ^ b[16];
  assign f_arrdiv32_fs720_not0 = ~f_arrdiv32_mux2to1666_xor0;
  assign f_arrdiv32_fs720_and0 = f_arrdiv32_fs720_not0 & b[16];
  assign f_arrdiv32_fs720_xor1 = f_arrdiv32_fs719_or0 ^ f_arrdiv32_fs720_xor0;
  assign f_arrdiv32_fs720_not1 = ~f_arrdiv32_fs720_xor0;
  assign f_arrdiv32_fs720_and1 = f_arrdiv32_fs720_not1 & f_arrdiv32_fs719_or0;
  assign f_arrdiv32_fs720_or0 = f_arrdiv32_fs720_and1 | f_arrdiv32_fs720_and0;
  assign f_arrdiv32_fs721_xor0 = f_arrdiv32_mux2to1667_xor0 ^ b[17];
  assign f_arrdiv32_fs721_not0 = ~f_arrdiv32_mux2to1667_xor0;
  assign f_arrdiv32_fs721_and0 = f_arrdiv32_fs721_not0 & b[17];
  assign f_arrdiv32_fs721_xor1 = f_arrdiv32_fs720_or0 ^ f_arrdiv32_fs721_xor0;
  assign f_arrdiv32_fs721_not1 = ~f_arrdiv32_fs721_xor0;
  assign f_arrdiv32_fs721_and1 = f_arrdiv32_fs721_not1 & f_arrdiv32_fs720_or0;
  assign f_arrdiv32_fs721_or0 = f_arrdiv32_fs721_and1 | f_arrdiv32_fs721_and0;
  assign f_arrdiv32_fs722_xor0 = f_arrdiv32_mux2to1668_xor0 ^ b[18];
  assign f_arrdiv32_fs722_not0 = ~f_arrdiv32_mux2to1668_xor0;
  assign f_arrdiv32_fs722_and0 = f_arrdiv32_fs722_not0 & b[18];
  assign f_arrdiv32_fs722_xor1 = f_arrdiv32_fs721_or0 ^ f_arrdiv32_fs722_xor0;
  assign f_arrdiv32_fs722_not1 = ~f_arrdiv32_fs722_xor0;
  assign f_arrdiv32_fs722_and1 = f_arrdiv32_fs722_not1 & f_arrdiv32_fs721_or0;
  assign f_arrdiv32_fs722_or0 = f_arrdiv32_fs722_and1 | f_arrdiv32_fs722_and0;
  assign f_arrdiv32_fs723_xor0 = f_arrdiv32_mux2to1669_xor0 ^ b[19];
  assign f_arrdiv32_fs723_not0 = ~f_arrdiv32_mux2to1669_xor0;
  assign f_arrdiv32_fs723_and0 = f_arrdiv32_fs723_not0 & b[19];
  assign f_arrdiv32_fs723_xor1 = f_arrdiv32_fs722_or0 ^ f_arrdiv32_fs723_xor0;
  assign f_arrdiv32_fs723_not1 = ~f_arrdiv32_fs723_xor0;
  assign f_arrdiv32_fs723_and1 = f_arrdiv32_fs723_not1 & f_arrdiv32_fs722_or0;
  assign f_arrdiv32_fs723_or0 = f_arrdiv32_fs723_and1 | f_arrdiv32_fs723_and0;
  assign f_arrdiv32_fs724_xor0 = f_arrdiv32_mux2to1670_xor0 ^ b[20];
  assign f_arrdiv32_fs724_not0 = ~f_arrdiv32_mux2to1670_xor0;
  assign f_arrdiv32_fs724_and0 = f_arrdiv32_fs724_not0 & b[20];
  assign f_arrdiv32_fs724_xor1 = f_arrdiv32_fs723_or0 ^ f_arrdiv32_fs724_xor0;
  assign f_arrdiv32_fs724_not1 = ~f_arrdiv32_fs724_xor0;
  assign f_arrdiv32_fs724_and1 = f_arrdiv32_fs724_not1 & f_arrdiv32_fs723_or0;
  assign f_arrdiv32_fs724_or0 = f_arrdiv32_fs724_and1 | f_arrdiv32_fs724_and0;
  assign f_arrdiv32_fs725_xor0 = f_arrdiv32_mux2to1671_xor0 ^ b[21];
  assign f_arrdiv32_fs725_not0 = ~f_arrdiv32_mux2to1671_xor0;
  assign f_arrdiv32_fs725_and0 = f_arrdiv32_fs725_not0 & b[21];
  assign f_arrdiv32_fs725_xor1 = f_arrdiv32_fs724_or0 ^ f_arrdiv32_fs725_xor0;
  assign f_arrdiv32_fs725_not1 = ~f_arrdiv32_fs725_xor0;
  assign f_arrdiv32_fs725_and1 = f_arrdiv32_fs725_not1 & f_arrdiv32_fs724_or0;
  assign f_arrdiv32_fs725_or0 = f_arrdiv32_fs725_and1 | f_arrdiv32_fs725_and0;
  assign f_arrdiv32_fs726_xor0 = f_arrdiv32_mux2to1672_xor0 ^ b[22];
  assign f_arrdiv32_fs726_not0 = ~f_arrdiv32_mux2to1672_xor0;
  assign f_arrdiv32_fs726_and0 = f_arrdiv32_fs726_not0 & b[22];
  assign f_arrdiv32_fs726_xor1 = f_arrdiv32_fs725_or0 ^ f_arrdiv32_fs726_xor0;
  assign f_arrdiv32_fs726_not1 = ~f_arrdiv32_fs726_xor0;
  assign f_arrdiv32_fs726_and1 = f_arrdiv32_fs726_not1 & f_arrdiv32_fs725_or0;
  assign f_arrdiv32_fs726_or0 = f_arrdiv32_fs726_and1 | f_arrdiv32_fs726_and0;
  assign f_arrdiv32_fs727_xor0 = f_arrdiv32_mux2to1673_xor0 ^ b[23];
  assign f_arrdiv32_fs727_not0 = ~f_arrdiv32_mux2to1673_xor0;
  assign f_arrdiv32_fs727_and0 = f_arrdiv32_fs727_not0 & b[23];
  assign f_arrdiv32_fs727_xor1 = f_arrdiv32_fs726_or0 ^ f_arrdiv32_fs727_xor0;
  assign f_arrdiv32_fs727_not1 = ~f_arrdiv32_fs727_xor0;
  assign f_arrdiv32_fs727_and1 = f_arrdiv32_fs727_not1 & f_arrdiv32_fs726_or0;
  assign f_arrdiv32_fs727_or0 = f_arrdiv32_fs727_and1 | f_arrdiv32_fs727_and0;
  assign f_arrdiv32_fs728_xor0 = f_arrdiv32_mux2to1674_xor0 ^ b[24];
  assign f_arrdiv32_fs728_not0 = ~f_arrdiv32_mux2to1674_xor0;
  assign f_arrdiv32_fs728_and0 = f_arrdiv32_fs728_not0 & b[24];
  assign f_arrdiv32_fs728_xor1 = f_arrdiv32_fs727_or0 ^ f_arrdiv32_fs728_xor0;
  assign f_arrdiv32_fs728_not1 = ~f_arrdiv32_fs728_xor0;
  assign f_arrdiv32_fs728_and1 = f_arrdiv32_fs728_not1 & f_arrdiv32_fs727_or0;
  assign f_arrdiv32_fs728_or0 = f_arrdiv32_fs728_and1 | f_arrdiv32_fs728_and0;
  assign f_arrdiv32_fs729_xor0 = f_arrdiv32_mux2to1675_xor0 ^ b[25];
  assign f_arrdiv32_fs729_not0 = ~f_arrdiv32_mux2to1675_xor0;
  assign f_arrdiv32_fs729_and0 = f_arrdiv32_fs729_not0 & b[25];
  assign f_arrdiv32_fs729_xor1 = f_arrdiv32_fs728_or0 ^ f_arrdiv32_fs729_xor0;
  assign f_arrdiv32_fs729_not1 = ~f_arrdiv32_fs729_xor0;
  assign f_arrdiv32_fs729_and1 = f_arrdiv32_fs729_not1 & f_arrdiv32_fs728_or0;
  assign f_arrdiv32_fs729_or0 = f_arrdiv32_fs729_and1 | f_arrdiv32_fs729_and0;
  assign f_arrdiv32_fs730_xor0 = f_arrdiv32_mux2to1676_xor0 ^ b[26];
  assign f_arrdiv32_fs730_not0 = ~f_arrdiv32_mux2to1676_xor0;
  assign f_arrdiv32_fs730_and0 = f_arrdiv32_fs730_not0 & b[26];
  assign f_arrdiv32_fs730_xor1 = f_arrdiv32_fs729_or0 ^ f_arrdiv32_fs730_xor0;
  assign f_arrdiv32_fs730_not1 = ~f_arrdiv32_fs730_xor0;
  assign f_arrdiv32_fs730_and1 = f_arrdiv32_fs730_not1 & f_arrdiv32_fs729_or0;
  assign f_arrdiv32_fs730_or0 = f_arrdiv32_fs730_and1 | f_arrdiv32_fs730_and0;
  assign f_arrdiv32_fs731_xor0 = f_arrdiv32_mux2to1677_xor0 ^ b[27];
  assign f_arrdiv32_fs731_not0 = ~f_arrdiv32_mux2to1677_xor0;
  assign f_arrdiv32_fs731_and0 = f_arrdiv32_fs731_not0 & b[27];
  assign f_arrdiv32_fs731_xor1 = f_arrdiv32_fs730_or0 ^ f_arrdiv32_fs731_xor0;
  assign f_arrdiv32_fs731_not1 = ~f_arrdiv32_fs731_xor0;
  assign f_arrdiv32_fs731_and1 = f_arrdiv32_fs731_not1 & f_arrdiv32_fs730_or0;
  assign f_arrdiv32_fs731_or0 = f_arrdiv32_fs731_and1 | f_arrdiv32_fs731_and0;
  assign f_arrdiv32_fs732_xor0 = f_arrdiv32_mux2to1678_xor0 ^ b[28];
  assign f_arrdiv32_fs732_not0 = ~f_arrdiv32_mux2to1678_xor0;
  assign f_arrdiv32_fs732_and0 = f_arrdiv32_fs732_not0 & b[28];
  assign f_arrdiv32_fs732_xor1 = f_arrdiv32_fs731_or0 ^ f_arrdiv32_fs732_xor0;
  assign f_arrdiv32_fs732_not1 = ~f_arrdiv32_fs732_xor0;
  assign f_arrdiv32_fs732_and1 = f_arrdiv32_fs732_not1 & f_arrdiv32_fs731_or0;
  assign f_arrdiv32_fs732_or0 = f_arrdiv32_fs732_and1 | f_arrdiv32_fs732_and0;
  assign f_arrdiv32_fs733_xor0 = f_arrdiv32_mux2to1679_xor0 ^ b[29];
  assign f_arrdiv32_fs733_not0 = ~f_arrdiv32_mux2to1679_xor0;
  assign f_arrdiv32_fs733_and0 = f_arrdiv32_fs733_not0 & b[29];
  assign f_arrdiv32_fs733_xor1 = f_arrdiv32_fs732_or0 ^ f_arrdiv32_fs733_xor0;
  assign f_arrdiv32_fs733_not1 = ~f_arrdiv32_fs733_xor0;
  assign f_arrdiv32_fs733_and1 = f_arrdiv32_fs733_not1 & f_arrdiv32_fs732_or0;
  assign f_arrdiv32_fs733_or0 = f_arrdiv32_fs733_and1 | f_arrdiv32_fs733_and0;
  assign f_arrdiv32_fs734_xor0 = f_arrdiv32_mux2to1680_xor0 ^ b[30];
  assign f_arrdiv32_fs734_not0 = ~f_arrdiv32_mux2to1680_xor0;
  assign f_arrdiv32_fs734_and0 = f_arrdiv32_fs734_not0 & b[30];
  assign f_arrdiv32_fs734_xor1 = f_arrdiv32_fs733_or0 ^ f_arrdiv32_fs734_xor0;
  assign f_arrdiv32_fs734_not1 = ~f_arrdiv32_fs734_xor0;
  assign f_arrdiv32_fs734_and1 = f_arrdiv32_fs734_not1 & f_arrdiv32_fs733_or0;
  assign f_arrdiv32_fs734_or0 = f_arrdiv32_fs734_and1 | f_arrdiv32_fs734_and0;
  assign f_arrdiv32_fs735_xor0 = f_arrdiv32_mux2to1681_xor0 ^ b[31];
  assign f_arrdiv32_fs735_not0 = ~f_arrdiv32_mux2to1681_xor0;
  assign f_arrdiv32_fs735_and0 = f_arrdiv32_fs735_not0 & b[31];
  assign f_arrdiv32_fs735_xor1 = f_arrdiv32_fs734_or0 ^ f_arrdiv32_fs735_xor0;
  assign f_arrdiv32_fs735_not1 = ~f_arrdiv32_fs735_xor0;
  assign f_arrdiv32_fs735_and1 = f_arrdiv32_fs735_not1 & f_arrdiv32_fs734_or0;
  assign f_arrdiv32_fs735_or0 = f_arrdiv32_fs735_and1 | f_arrdiv32_fs735_and0;
  assign f_arrdiv32_mux2to1682_and0 = a[9] & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1682_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1682_and1 = f_arrdiv32_fs704_xor0 & f_arrdiv32_mux2to1682_not0;
  assign f_arrdiv32_mux2to1682_xor0 = f_arrdiv32_mux2to1682_and0 ^ f_arrdiv32_mux2to1682_and1;
  assign f_arrdiv32_mux2to1683_and0 = f_arrdiv32_mux2to1651_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1683_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1683_and1 = f_arrdiv32_fs705_xor1 & f_arrdiv32_mux2to1683_not0;
  assign f_arrdiv32_mux2to1683_xor0 = f_arrdiv32_mux2to1683_and0 ^ f_arrdiv32_mux2to1683_and1;
  assign f_arrdiv32_mux2to1684_and0 = f_arrdiv32_mux2to1652_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1684_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1684_and1 = f_arrdiv32_fs706_xor1 & f_arrdiv32_mux2to1684_not0;
  assign f_arrdiv32_mux2to1684_xor0 = f_arrdiv32_mux2to1684_and0 ^ f_arrdiv32_mux2to1684_and1;
  assign f_arrdiv32_mux2to1685_and0 = f_arrdiv32_mux2to1653_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1685_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1685_and1 = f_arrdiv32_fs707_xor1 & f_arrdiv32_mux2to1685_not0;
  assign f_arrdiv32_mux2to1685_xor0 = f_arrdiv32_mux2to1685_and0 ^ f_arrdiv32_mux2to1685_and1;
  assign f_arrdiv32_mux2to1686_and0 = f_arrdiv32_mux2to1654_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1686_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1686_and1 = f_arrdiv32_fs708_xor1 & f_arrdiv32_mux2to1686_not0;
  assign f_arrdiv32_mux2to1686_xor0 = f_arrdiv32_mux2to1686_and0 ^ f_arrdiv32_mux2to1686_and1;
  assign f_arrdiv32_mux2to1687_and0 = f_arrdiv32_mux2to1655_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1687_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1687_and1 = f_arrdiv32_fs709_xor1 & f_arrdiv32_mux2to1687_not0;
  assign f_arrdiv32_mux2to1687_xor0 = f_arrdiv32_mux2to1687_and0 ^ f_arrdiv32_mux2to1687_and1;
  assign f_arrdiv32_mux2to1688_and0 = f_arrdiv32_mux2to1656_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1688_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1688_and1 = f_arrdiv32_fs710_xor1 & f_arrdiv32_mux2to1688_not0;
  assign f_arrdiv32_mux2to1688_xor0 = f_arrdiv32_mux2to1688_and0 ^ f_arrdiv32_mux2to1688_and1;
  assign f_arrdiv32_mux2to1689_and0 = f_arrdiv32_mux2to1657_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1689_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1689_and1 = f_arrdiv32_fs711_xor1 & f_arrdiv32_mux2to1689_not0;
  assign f_arrdiv32_mux2to1689_xor0 = f_arrdiv32_mux2to1689_and0 ^ f_arrdiv32_mux2to1689_and1;
  assign f_arrdiv32_mux2to1690_and0 = f_arrdiv32_mux2to1658_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1690_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1690_and1 = f_arrdiv32_fs712_xor1 & f_arrdiv32_mux2to1690_not0;
  assign f_arrdiv32_mux2to1690_xor0 = f_arrdiv32_mux2to1690_and0 ^ f_arrdiv32_mux2to1690_and1;
  assign f_arrdiv32_mux2to1691_and0 = f_arrdiv32_mux2to1659_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1691_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1691_and1 = f_arrdiv32_fs713_xor1 & f_arrdiv32_mux2to1691_not0;
  assign f_arrdiv32_mux2to1691_xor0 = f_arrdiv32_mux2to1691_and0 ^ f_arrdiv32_mux2to1691_and1;
  assign f_arrdiv32_mux2to1692_and0 = f_arrdiv32_mux2to1660_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1692_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1692_and1 = f_arrdiv32_fs714_xor1 & f_arrdiv32_mux2to1692_not0;
  assign f_arrdiv32_mux2to1692_xor0 = f_arrdiv32_mux2to1692_and0 ^ f_arrdiv32_mux2to1692_and1;
  assign f_arrdiv32_mux2to1693_and0 = f_arrdiv32_mux2to1661_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1693_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1693_and1 = f_arrdiv32_fs715_xor1 & f_arrdiv32_mux2to1693_not0;
  assign f_arrdiv32_mux2to1693_xor0 = f_arrdiv32_mux2to1693_and0 ^ f_arrdiv32_mux2to1693_and1;
  assign f_arrdiv32_mux2to1694_and0 = f_arrdiv32_mux2to1662_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1694_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1694_and1 = f_arrdiv32_fs716_xor1 & f_arrdiv32_mux2to1694_not0;
  assign f_arrdiv32_mux2to1694_xor0 = f_arrdiv32_mux2to1694_and0 ^ f_arrdiv32_mux2to1694_and1;
  assign f_arrdiv32_mux2to1695_and0 = f_arrdiv32_mux2to1663_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1695_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1695_and1 = f_arrdiv32_fs717_xor1 & f_arrdiv32_mux2to1695_not0;
  assign f_arrdiv32_mux2to1695_xor0 = f_arrdiv32_mux2to1695_and0 ^ f_arrdiv32_mux2to1695_and1;
  assign f_arrdiv32_mux2to1696_and0 = f_arrdiv32_mux2to1664_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1696_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1696_and1 = f_arrdiv32_fs718_xor1 & f_arrdiv32_mux2to1696_not0;
  assign f_arrdiv32_mux2to1696_xor0 = f_arrdiv32_mux2to1696_and0 ^ f_arrdiv32_mux2to1696_and1;
  assign f_arrdiv32_mux2to1697_and0 = f_arrdiv32_mux2to1665_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1697_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1697_and1 = f_arrdiv32_fs719_xor1 & f_arrdiv32_mux2to1697_not0;
  assign f_arrdiv32_mux2to1697_xor0 = f_arrdiv32_mux2to1697_and0 ^ f_arrdiv32_mux2to1697_and1;
  assign f_arrdiv32_mux2to1698_and0 = f_arrdiv32_mux2to1666_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1698_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1698_and1 = f_arrdiv32_fs720_xor1 & f_arrdiv32_mux2to1698_not0;
  assign f_arrdiv32_mux2to1698_xor0 = f_arrdiv32_mux2to1698_and0 ^ f_arrdiv32_mux2to1698_and1;
  assign f_arrdiv32_mux2to1699_and0 = f_arrdiv32_mux2to1667_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1699_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1699_and1 = f_arrdiv32_fs721_xor1 & f_arrdiv32_mux2to1699_not0;
  assign f_arrdiv32_mux2to1699_xor0 = f_arrdiv32_mux2to1699_and0 ^ f_arrdiv32_mux2to1699_and1;
  assign f_arrdiv32_mux2to1700_and0 = f_arrdiv32_mux2to1668_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1700_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1700_and1 = f_arrdiv32_fs722_xor1 & f_arrdiv32_mux2to1700_not0;
  assign f_arrdiv32_mux2to1700_xor0 = f_arrdiv32_mux2to1700_and0 ^ f_arrdiv32_mux2to1700_and1;
  assign f_arrdiv32_mux2to1701_and0 = f_arrdiv32_mux2to1669_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1701_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1701_and1 = f_arrdiv32_fs723_xor1 & f_arrdiv32_mux2to1701_not0;
  assign f_arrdiv32_mux2to1701_xor0 = f_arrdiv32_mux2to1701_and0 ^ f_arrdiv32_mux2to1701_and1;
  assign f_arrdiv32_mux2to1702_and0 = f_arrdiv32_mux2to1670_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1702_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1702_and1 = f_arrdiv32_fs724_xor1 & f_arrdiv32_mux2to1702_not0;
  assign f_arrdiv32_mux2to1702_xor0 = f_arrdiv32_mux2to1702_and0 ^ f_arrdiv32_mux2to1702_and1;
  assign f_arrdiv32_mux2to1703_and0 = f_arrdiv32_mux2to1671_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1703_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1703_and1 = f_arrdiv32_fs725_xor1 & f_arrdiv32_mux2to1703_not0;
  assign f_arrdiv32_mux2to1703_xor0 = f_arrdiv32_mux2to1703_and0 ^ f_arrdiv32_mux2to1703_and1;
  assign f_arrdiv32_mux2to1704_and0 = f_arrdiv32_mux2to1672_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1704_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1704_and1 = f_arrdiv32_fs726_xor1 & f_arrdiv32_mux2to1704_not0;
  assign f_arrdiv32_mux2to1704_xor0 = f_arrdiv32_mux2to1704_and0 ^ f_arrdiv32_mux2to1704_and1;
  assign f_arrdiv32_mux2to1705_and0 = f_arrdiv32_mux2to1673_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1705_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1705_and1 = f_arrdiv32_fs727_xor1 & f_arrdiv32_mux2to1705_not0;
  assign f_arrdiv32_mux2to1705_xor0 = f_arrdiv32_mux2to1705_and0 ^ f_arrdiv32_mux2to1705_and1;
  assign f_arrdiv32_mux2to1706_and0 = f_arrdiv32_mux2to1674_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1706_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1706_and1 = f_arrdiv32_fs728_xor1 & f_arrdiv32_mux2to1706_not0;
  assign f_arrdiv32_mux2to1706_xor0 = f_arrdiv32_mux2to1706_and0 ^ f_arrdiv32_mux2to1706_and1;
  assign f_arrdiv32_mux2to1707_and0 = f_arrdiv32_mux2to1675_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1707_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1707_and1 = f_arrdiv32_fs729_xor1 & f_arrdiv32_mux2to1707_not0;
  assign f_arrdiv32_mux2to1707_xor0 = f_arrdiv32_mux2to1707_and0 ^ f_arrdiv32_mux2to1707_and1;
  assign f_arrdiv32_mux2to1708_and0 = f_arrdiv32_mux2to1676_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1708_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1708_and1 = f_arrdiv32_fs730_xor1 & f_arrdiv32_mux2to1708_not0;
  assign f_arrdiv32_mux2to1708_xor0 = f_arrdiv32_mux2to1708_and0 ^ f_arrdiv32_mux2to1708_and1;
  assign f_arrdiv32_mux2to1709_and0 = f_arrdiv32_mux2to1677_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1709_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1709_and1 = f_arrdiv32_fs731_xor1 & f_arrdiv32_mux2to1709_not0;
  assign f_arrdiv32_mux2to1709_xor0 = f_arrdiv32_mux2to1709_and0 ^ f_arrdiv32_mux2to1709_and1;
  assign f_arrdiv32_mux2to1710_and0 = f_arrdiv32_mux2to1678_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1710_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1710_and1 = f_arrdiv32_fs732_xor1 & f_arrdiv32_mux2to1710_not0;
  assign f_arrdiv32_mux2to1710_xor0 = f_arrdiv32_mux2to1710_and0 ^ f_arrdiv32_mux2to1710_and1;
  assign f_arrdiv32_mux2to1711_and0 = f_arrdiv32_mux2to1679_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1711_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1711_and1 = f_arrdiv32_fs733_xor1 & f_arrdiv32_mux2to1711_not0;
  assign f_arrdiv32_mux2to1711_xor0 = f_arrdiv32_mux2to1711_and0 ^ f_arrdiv32_mux2to1711_and1;
  assign f_arrdiv32_mux2to1712_and0 = f_arrdiv32_mux2to1680_xor0 & f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1712_not0 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_mux2to1712_and1 = f_arrdiv32_fs734_xor1 & f_arrdiv32_mux2to1712_not0;
  assign f_arrdiv32_mux2to1712_xor0 = f_arrdiv32_mux2to1712_and0 ^ f_arrdiv32_mux2to1712_and1;
  assign f_arrdiv32_not22 = ~f_arrdiv32_fs735_or0;
  assign f_arrdiv32_fs736_xor0 = a[8] ^ b[0];
  assign f_arrdiv32_fs736_not0 = ~a[8];
  assign f_arrdiv32_fs736_and0 = f_arrdiv32_fs736_not0 & b[0];
  assign f_arrdiv32_fs736_not1 = ~f_arrdiv32_fs736_xor0;
  assign f_arrdiv32_fs737_xor0 = f_arrdiv32_mux2to1682_xor0 ^ b[1];
  assign f_arrdiv32_fs737_not0 = ~f_arrdiv32_mux2to1682_xor0;
  assign f_arrdiv32_fs737_and0 = f_arrdiv32_fs737_not0 & b[1];
  assign f_arrdiv32_fs737_xor1 = f_arrdiv32_fs736_and0 ^ f_arrdiv32_fs737_xor0;
  assign f_arrdiv32_fs737_not1 = ~f_arrdiv32_fs737_xor0;
  assign f_arrdiv32_fs737_and1 = f_arrdiv32_fs737_not1 & f_arrdiv32_fs736_and0;
  assign f_arrdiv32_fs737_or0 = f_arrdiv32_fs737_and1 | f_arrdiv32_fs737_and0;
  assign f_arrdiv32_fs738_xor0 = f_arrdiv32_mux2to1683_xor0 ^ b[2];
  assign f_arrdiv32_fs738_not0 = ~f_arrdiv32_mux2to1683_xor0;
  assign f_arrdiv32_fs738_and0 = f_arrdiv32_fs738_not0 & b[2];
  assign f_arrdiv32_fs738_xor1 = f_arrdiv32_fs737_or0 ^ f_arrdiv32_fs738_xor0;
  assign f_arrdiv32_fs738_not1 = ~f_arrdiv32_fs738_xor0;
  assign f_arrdiv32_fs738_and1 = f_arrdiv32_fs738_not1 & f_arrdiv32_fs737_or0;
  assign f_arrdiv32_fs738_or0 = f_arrdiv32_fs738_and1 | f_arrdiv32_fs738_and0;
  assign f_arrdiv32_fs739_xor0 = f_arrdiv32_mux2to1684_xor0 ^ b[3];
  assign f_arrdiv32_fs739_not0 = ~f_arrdiv32_mux2to1684_xor0;
  assign f_arrdiv32_fs739_and0 = f_arrdiv32_fs739_not0 & b[3];
  assign f_arrdiv32_fs739_xor1 = f_arrdiv32_fs738_or0 ^ f_arrdiv32_fs739_xor0;
  assign f_arrdiv32_fs739_not1 = ~f_arrdiv32_fs739_xor0;
  assign f_arrdiv32_fs739_and1 = f_arrdiv32_fs739_not1 & f_arrdiv32_fs738_or0;
  assign f_arrdiv32_fs739_or0 = f_arrdiv32_fs739_and1 | f_arrdiv32_fs739_and0;
  assign f_arrdiv32_fs740_xor0 = f_arrdiv32_mux2to1685_xor0 ^ b[4];
  assign f_arrdiv32_fs740_not0 = ~f_arrdiv32_mux2to1685_xor0;
  assign f_arrdiv32_fs740_and0 = f_arrdiv32_fs740_not0 & b[4];
  assign f_arrdiv32_fs740_xor1 = f_arrdiv32_fs739_or0 ^ f_arrdiv32_fs740_xor0;
  assign f_arrdiv32_fs740_not1 = ~f_arrdiv32_fs740_xor0;
  assign f_arrdiv32_fs740_and1 = f_arrdiv32_fs740_not1 & f_arrdiv32_fs739_or0;
  assign f_arrdiv32_fs740_or0 = f_arrdiv32_fs740_and1 | f_arrdiv32_fs740_and0;
  assign f_arrdiv32_fs741_xor0 = f_arrdiv32_mux2to1686_xor0 ^ b[5];
  assign f_arrdiv32_fs741_not0 = ~f_arrdiv32_mux2to1686_xor0;
  assign f_arrdiv32_fs741_and0 = f_arrdiv32_fs741_not0 & b[5];
  assign f_arrdiv32_fs741_xor1 = f_arrdiv32_fs740_or0 ^ f_arrdiv32_fs741_xor0;
  assign f_arrdiv32_fs741_not1 = ~f_arrdiv32_fs741_xor0;
  assign f_arrdiv32_fs741_and1 = f_arrdiv32_fs741_not1 & f_arrdiv32_fs740_or0;
  assign f_arrdiv32_fs741_or0 = f_arrdiv32_fs741_and1 | f_arrdiv32_fs741_and0;
  assign f_arrdiv32_fs742_xor0 = f_arrdiv32_mux2to1687_xor0 ^ b[6];
  assign f_arrdiv32_fs742_not0 = ~f_arrdiv32_mux2to1687_xor0;
  assign f_arrdiv32_fs742_and0 = f_arrdiv32_fs742_not0 & b[6];
  assign f_arrdiv32_fs742_xor1 = f_arrdiv32_fs741_or0 ^ f_arrdiv32_fs742_xor0;
  assign f_arrdiv32_fs742_not1 = ~f_arrdiv32_fs742_xor0;
  assign f_arrdiv32_fs742_and1 = f_arrdiv32_fs742_not1 & f_arrdiv32_fs741_or0;
  assign f_arrdiv32_fs742_or0 = f_arrdiv32_fs742_and1 | f_arrdiv32_fs742_and0;
  assign f_arrdiv32_fs743_xor0 = f_arrdiv32_mux2to1688_xor0 ^ b[7];
  assign f_arrdiv32_fs743_not0 = ~f_arrdiv32_mux2to1688_xor0;
  assign f_arrdiv32_fs743_and0 = f_arrdiv32_fs743_not0 & b[7];
  assign f_arrdiv32_fs743_xor1 = f_arrdiv32_fs742_or0 ^ f_arrdiv32_fs743_xor0;
  assign f_arrdiv32_fs743_not1 = ~f_arrdiv32_fs743_xor0;
  assign f_arrdiv32_fs743_and1 = f_arrdiv32_fs743_not1 & f_arrdiv32_fs742_or0;
  assign f_arrdiv32_fs743_or0 = f_arrdiv32_fs743_and1 | f_arrdiv32_fs743_and0;
  assign f_arrdiv32_fs744_xor0 = f_arrdiv32_mux2to1689_xor0 ^ b[8];
  assign f_arrdiv32_fs744_not0 = ~f_arrdiv32_mux2to1689_xor0;
  assign f_arrdiv32_fs744_and0 = f_arrdiv32_fs744_not0 & b[8];
  assign f_arrdiv32_fs744_xor1 = f_arrdiv32_fs743_or0 ^ f_arrdiv32_fs744_xor0;
  assign f_arrdiv32_fs744_not1 = ~f_arrdiv32_fs744_xor0;
  assign f_arrdiv32_fs744_and1 = f_arrdiv32_fs744_not1 & f_arrdiv32_fs743_or0;
  assign f_arrdiv32_fs744_or0 = f_arrdiv32_fs744_and1 | f_arrdiv32_fs744_and0;
  assign f_arrdiv32_fs745_xor0 = f_arrdiv32_mux2to1690_xor0 ^ b[9];
  assign f_arrdiv32_fs745_not0 = ~f_arrdiv32_mux2to1690_xor0;
  assign f_arrdiv32_fs745_and0 = f_arrdiv32_fs745_not0 & b[9];
  assign f_arrdiv32_fs745_xor1 = f_arrdiv32_fs744_or0 ^ f_arrdiv32_fs745_xor0;
  assign f_arrdiv32_fs745_not1 = ~f_arrdiv32_fs745_xor0;
  assign f_arrdiv32_fs745_and1 = f_arrdiv32_fs745_not1 & f_arrdiv32_fs744_or0;
  assign f_arrdiv32_fs745_or0 = f_arrdiv32_fs745_and1 | f_arrdiv32_fs745_and0;
  assign f_arrdiv32_fs746_xor0 = f_arrdiv32_mux2to1691_xor0 ^ b[10];
  assign f_arrdiv32_fs746_not0 = ~f_arrdiv32_mux2to1691_xor0;
  assign f_arrdiv32_fs746_and0 = f_arrdiv32_fs746_not0 & b[10];
  assign f_arrdiv32_fs746_xor1 = f_arrdiv32_fs745_or0 ^ f_arrdiv32_fs746_xor0;
  assign f_arrdiv32_fs746_not1 = ~f_arrdiv32_fs746_xor0;
  assign f_arrdiv32_fs746_and1 = f_arrdiv32_fs746_not1 & f_arrdiv32_fs745_or0;
  assign f_arrdiv32_fs746_or0 = f_arrdiv32_fs746_and1 | f_arrdiv32_fs746_and0;
  assign f_arrdiv32_fs747_xor0 = f_arrdiv32_mux2to1692_xor0 ^ b[11];
  assign f_arrdiv32_fs747_not0 = ~f_arrdiv32_mux2to1692_xor0;
  assign f_arrdiv32_fs747_and0 = f_arrdiv32_fs747_not0 & b[11];
  assign f_arrdiv32_fs747_xor1 = f_arrdiv32_fs746_or0 ^ f_arrdiv32_fs747_xor0;
  assign f_arrdiv32_fs747_not1 = ~f_arrdiv32_fs747_xor0;
  assign f_arrdiv32_fs747_and1 = f_arrdiv32_fs747_not1 & f_arrdiv32_fs746_or0;
  assign f_arrdiv32_fs747_or0 = f_arrdiv32_fs747_and1 | f_arrdiv32_fs747_and0;
  assign f_arrdiv32_fs748_xor0 = f_arrdiv32_mux2to1693_xor0 ^ b[12];
  assign f_arrdiv32_fs748_not0 = ~f_arrdiv32_mux2to1693_xor0;
  assign f_arrdiv32_fs748_and0 = f_arrdiv32_fs748_not0 & b[12];
  assign f_arrdiv32_fs748_xor1 = f_arrdiv32_fs747_or0 ^ f_arrdiv32_fs748_xor0;
  assign f_arrdiv32_fs748_not1 = ~f_arrdiv32_fs748_xor0;
  assign f_arrdiv32_fs748_and1 = f_arrdiv32_fs748_not1 & f_arrdiv32_fs747_or0;
  assign f_arrdiv32_fs748_or0 = f_arrdiv32_fs748_and1 | f_arrdiv32_fs748_and0;
  assign f_arrdiv32_fs749_xor0 = f_arrdiv32_mux2to1694_xor0 ^ b[13];
  assign f_arrdiv32_fs749_not0 = ~f_arrdiv32_mux2to1694_xor0;
  assign f_arrdiv32_fs749_and0 = f_arrdiv32_fs749_not0 & b[13];
  assign f_arrdiv32_fs749_xor1 = f_arrdiv32_fs748_or0 ^ f_arrdiv32_fs749_xor0;
  assign f_arrdiv32_fs749_not1 = ~f_arrdiv32_fs749_xor0;
  assign f_arrdiv32_fs749_and1 = f_arrdiv32_fs749_not1 & f_arrdiv32_fs748_or0;
  assign f_arrdiv32_fs749_or0 = f_arrdiv32_fs749_and1 | f_arrdiv32_fs749_and0;
  assign f_arrdiv32_fs750_xor0 = f_arrdiv32_mux2to1695_xor0 ^ b[14];
  assign f_arrdiv32_fs750_not0 = ~f_arrdiv32_mux2to1695_xor0;
  assign f_arrdiv32_fs750_and0 = f_arrdiv32_fs750_not0 & b[14];
  assign f_arrdiv32_fs750_xor1 = f_arrdiv32_fs749_or0 ^ f_arrdiv32_fs750_xor0;
  assign f_arrdiv32_fs750_not1 = ~f_arrdiv32_fs750_xor0;
  assign f_arrdiv32_fs750_and1 = f_arrdiv32_fs750_not1 & f_arrdiv32_fs749_or0;
  assign f_arrdiv32_fs750_or0 = f_arrdiv32_fs750_and1 | f_arrdiv32_fs750_and0;
  assign f_arrdiv32_fs751_xor0 = f_arrdiv32_mux2to1696_xor0 ^ b[15];
  assign f_arrdiv32_fs751_not0 = ~f_arrdiv32_mux2to1696_xor0;
  assign f_arrdiv32_fs751_and0 = f_arrdiv32_fs751_not0 & b[15];
  assign f_arrdiv32_fs751_xor1 = f_arrdiv32_fs750_or0 ^ f_arrdiv32_fs751_xor0;
  assign f_arrdiv32_fs751_not1 = ~f_arrdiv32_fs751_xor0;
  assign f_arrdiv32_fs751_and1 = f_arrdiv32_fs751_not1 & f_arrdiv32_fs750_or0;
  assign f_arrdiv32_fs751_or0 = f_arrdiv32_fs751_and1 | f_arrdiv32_fs751_and0;
  assign f_arrdiv32_fs752_xor0 = f_arrdiv32_mux2to1697_xor0 ^ b[16];
  assign f_arrdiv32_fs752_not0 = ~f_arrdiv32_mux2to1697_xor0;
  assign f_arrdiv32_fs752_and0 = f_arrdiv32_fs752_not0 & b[16];
  assign f_arrdiv32_fs752_xor1 = f_arrdiv32_fs751_or0 ^ f_arrdiv32_fs752_xor0;
  assign f_arrdiv32_fs752_not1 = ~f_arrdiv32_fs752_xor0;
  assign f_arrdiv32_fs752_and1 = f_arrdiv32_fs752_not1 & f_arrdiv32_fs751_or0;
  assign f_arrdiv32_fs752_or0 = f_arrdiv32_fs752_and1 | f_arrdiv32_fs752_and0;
  assign f_arrdiv32_fs753_xor0 = f_arrdiv32_mux2to1698_xor0 ^ b[17];
  assign f_arrdiv32_fs753_not0 = ~f_arrdiv32_mux2to1698_xor0;
  assign f_arrdiv32_fs753_and0 = f_arrdiv32_fs753_not0 & b[17];
  assign f_arrdiv32_fs753_xor1 = f_arrdiv32_fs752_or0 ^ f_arrdiv32_fs753_xor0;
  assign f_arrdiv32_fs753_not1 = ~f_arrdiv32_fs753_xor0;
  assign f_arrdiv32_fs753_and1 = f_arrdiv32_fs753_not1 & f_arrdiv32_fs752_or0;
  assign f_arrdiv32_fs753_or0 = f_arrdiv32_fs753_and1 | f_arrdiv32_fs753_and0;
  assign f_arrdiv32_fs754_xor0 = f_arrdiv32_mux2to1699_xor0 ^ b[18];
  assign f_arrdiv32_fs754_not0 = ~f_arrdiv32_mux2to1699_xor0;
  assign f_arrdiv32_fs754_and0 = f_arrdiv32_fs754_not0 & b[18];
  assign f_arrdiv32_fs754_xor1 = f_arrdiv32_fs753_or0 ^ f_arrdiv32_fs754_xor0;
  assign f_arrdiv32_fs754_not1 = ~f_arrdiv32_fs754_xor0;
  assign f_arrdiv32_fs754_and1 = f_arrdiv32_fs754_not1 & f_arrdiv32_fs753_or0;
  assign f_arrdiv32_fs754_or0 = f_arrdiv32_fs754_and1 | f_arrdiv32_fs754_and0;
  assign f_arrdiv32_fs755_xor0 = f_arrdiv32_mux2to1700_xor0 ^ b[19];
  assign f_arrdiv32_fs755_not0 = ~f_arrdiv32_mux2to1700_xor0;
  assign f_arrdiv32_fs755_and0 = f_arrdiv32_fs755_not0 & b[19];
  assign f_arrdiv32_fs755_xor1 = f_arrdiv32_fs754_or0 ^ f_arrdiv32_fs755_xor0;
  assign f_arrdiv32_fs755_not1 = ~f_arrdiv32_fs755_xor0;
  assign f_arrdiv32_fs755_and1 = f_arrdiv32_fs755_not1 & f_arrdiv32_fs754_or0;
  assign f_arrdiv32_fs755_or0 = f_arrdiv32_fs755_and1 | f_arrdiv32_fs755_and0;
  assign f_arrdiv32_fs756_xor0 = f_arrdiv32_mux2to1701_xor0 ^ b[20];
  assign f_arrdiv32_fs756_not0 = ~f_arrdiv32_mux2to1701_xor0;
  assign f_arrdiv32_fs756_and0 = f_arrdiv32_fs756_not0 & b[20];
  assign f_arrdiv32_fs756_xor1 = f_arrdiv32_fs755_or0 ^ f_arrdiv32_fs756_xor0;
  assign f_arrdiv32_fs756_not1 = ~f_arrdiv32_fs756_xor0;
  assign f_arrdiv32_fs756_and1 = f_arrdiv32_fs756_not1 & f_arrdiv32_fs755_or0;
  assign f_arrdiv32_fs756_or0 = f_arrdiv32_fs756_and1 | f_arrdiv32_fs756_and0;
  assign f_arrdiv32_fs757_xor0 = f_arrdiv32_mux2to1702_xor0 ^ b[21];
  assign f_arrdiv32_fs757_not0 = ~f_arrdiv32_mux2to1702_xor0;
  assign f_arrdiv32_fs757_and0 = f_arrdiv32_fs757_not0 & b[21];
  assign f_arrdiv32_fs757_xor1 = f_arrdiv32_fs756_or0 ^ f_arrdiv32_fs757_xor0;
  assign f_arrdiv32_fs757_not1 = ~f_arrdiv32_fs757_xor0;
  assign f_arrdiv32_fs757_and1 = f_arrdiv32_fs757_not1 & f_arrdiv32_fs756_or0;
  assign f_arrdiv32_fs757_or0 = f_arrdiv32_fs757_and1 | f_arrdiv32_fs757_and0;
  assign f_arrdiv32_fs758_xor0 = f_arrdiv32_mux2to1703_xor0 ^ b[22];
  assign f_arrdiv32_fs758_not0 = ~f_arrdiv32_mux2to1703_xor0;
  assign f_arrdiv32_fs758_and0 = f_arrdiv32_fs758_not0 & b[22];
  assign f_arrdiv32_fs758_xor1 = f_arrdiv32_fs757_or0 ^ f_arrdiv32_fs758_xor0;
  assign f_arrdiv32_fs758_not1 = ~f_arrdiv32_fs758_xor0;
  assign f_arrdiv32_fs758_and1 = f_arrdiv32_fs758_not1 & f_arrdiv32_fs757_or0;
  assign f_arrdiv32_fs758_or0 = f_arrdiv32_fs758_and1 | f_arrdiv32_fs758_and0;
  assign f_arrdiv32_fs759_xor0 = f_arrdiv32_mux2to1704_xor0 ^ b[23];
  assign f_arrdiv32_fs759_not0 = ~f_arrdiv32_mux2to1704_xor0;
  assign f_arrdiv32_fs759_and0 = f_arrdiv32_fs759_not0 & b[23];
  assign f_arrdiv32_fs759_xor1 = f_arrdiv32_fs758_or0 ^ f_arrdiv32_fs759_xor0;
  assign f_arrdiv32_fs759_not1 = ~f_arrdiv32_fs759_xor0;
  assign f_arrdiv32_fs759_and1 = f_arrdiv32_fs759_not1 & f_arrdiv32_fs758_or0;
  assign f_arrdiv32_fs759_or0 = f_arrdiv32_fs759_and1 | f_arrdiv32_fs759_and0;
  assign f_arrdiv32_fs760_xor0 = f_arrdiv32_mux2to1705_xor0 ^ b[24];
  assign f_arrdiv32_fs760_not0 = ~f_arrdiv32_mux2to1705_xor0;
  assign f_arrdiv32_fs760_and0 = f_arrdiv32_fs760_not0 & b[24];
  assign f_arrdiv32_fs760_xor1 = f_arrdiv32_fs759_or0 ^ f_arrdiv32_fs760_xor0;
  assign f_arrdiv32_fs760_not1 = ~f_arrdiv32_fs760_xor0;
  assign f_arrdiv32_fs760_and1 = f_arrdiv32_fs760_not1 & f_arrdiv32_fs759_or0;
  assign f_arrdiv32_fs760_or0 = f_arrdiv32_fs760_and1 | f_arrdiv32_fs760_and0;
  assign f_arrdiv32_fs761_xor0 = f_arrdiv32_mux2to1706_xor0 ^ b[25];
  assign f_arrdiv32_fs761_not0 = ~f_arrdiv32_mux2to1706_xor0;
  assign f_arrdiv32_fs761_and0 = f_arrdiv32_fs761_not0 & b[25];
  assign f_arrdiv32_fs761_xor1 = f_arrdiv32_fs760_or0 ^ f_arrdiv32_fs761_xor0;
  assign f_arrdiv32_fs761_not1 = ~f_arrdiv32_fs761_xor0;
  assign f_arrdiv32_fs761_and1 = f_arrdiv32_fs761_not1 & f_arrdiv32_fs760_or0;
  assign f_arrdiv32_fs761_or0 = f_arrdiv32_fs761_and1 | f_arrdiv32_fs761_and0;
  assign f_arrdiv32_fs762_xor0 = f_arrdiv32_mux2to1707_xor0 ^ b[26];
  assign f_arrdiv32_fs762_not0 = ~f_arrdiv32_mux2to1707_xor0;
  assign f_arrdiv32_fs762_and0 = f_arrdiv32_fs762_not0 & b[26];
  assign f_arrdiv32_fs762_xor1 = f_arrdiv32_fs761_or0 ^ f_arrdiv32_fs762_xor0;
  assign f_arrdiv32_fs762_not1 = ~f_arrdiv32_fs762_xor0;
  assign f_arrdiv32_fs762_and1 = f_arrdiv32_fs762_not1 & f_arrdiv32_fs761_or0;
  assign f_arrdiv32_fs762_or0 = f_arrdiv32_fs762_and1 | f_arrdiv32_fs762_and0;
  assign f_arrdiv32_fs763_xor0 = f_arrdiv32_mux2to1708_xor0 ^ b[27];
  assign f_arrdiv32_fs763_not0 = ~f_arrdiv32_mux2to1708_xor0;
  assign f_arrdiv32_fs763_and0 = f_arrdiv32_fs763_not0 & b[27];
  assign f_arrdiv32_fs763_xor1 = f_arrdiv32_fs762_or0 ^ f_arrdiv32_fs763_xor0;
  assign f_arrdiv32_fs763_not1 = ~f_arrdiv32_fs763_xor0;
  assign f_arrdiv32_fs763_and1 = f_arrdiv32_fs763_not1 & f_arrdiv32_fs762_or0;
  assign f_arrdiv32_fs763_or0 = f_arrdiv32_fs763_and1 | f_arrdiv32_fs763_and0;
  assign f_arrdiv32_fs764_xor0 = f_arrdiv32_mux2to1709_xor0 ^ b[28];
  assign f_arrdiv32_fs764_not0 = ~f_arrdiv32_mux2to1709_xor0;
  assign f_arrdiv32_fs764_and0 = f_arrdiv32_fs764_not0 & b[28];
  assign f_arrdiv32_fs764_xor1 = f_arrdiv32_fs763_or0 ^ f_arrdiv32_fs764_xor0;
  assign f_arrdiv32_fs764_not1 = ~f_arrdiv32_fs764_xor0;
  assign f_arrdiv32_fs764_and1 = f_arrdiv32_fs764_not1 & f_arrdiv32_fs763_or0;
  assign f_arrdiv32_fs764_or0 = f_arrdiv32_fs764_and1 | f_arrdiv32_fs764_and0;
  assign f_arrdiv32_fs765_xor0 = f_arrdiv32_mux2to1710_xor0 ^ b[29];
  assign f_arrdiv32_fs765_not0 = ~f_arrdiv32_mux2to1710_xor0;
  assign f_arrdiv32_fs765_and0 = f_arrdiv32_fs765_not0 & b[29];
  assign f_arrdiv32_fs765_xor1 = f_arrdiv32_fs764_or0 ^ f_arrdiv32_fs765_xor0;
  assign f_arrdiv32_fs765_not1 = ~f_arrdiv32_fs765_xor0;
  assign f_arrdiv32_fs765_and1 = f_arrdiv32_fs765_not1 & f_arrdiv32_fs764_or0;
  assign f_arrdiv32_fs765_or0 = f_arrdiv32_fs765_and1 | f_arrdiv32_fs765_and0;
  assign f_arrdiv32_fs766_xor0 = f_arrdiv32_mux2to1711_xor0 ^ b[30];
  assign f_arrdiv32_fs766_not0 = ~f_arrdiv32_mux2to1711_xor0;
  assign f_arrdiv32_fs766_and0 = f_arrdiv32_fs766_not0 & b[30];
  assign f_arrdiv32_fs766_xor1 = f_arrdiv32_fs765_or0 ^ f_arrdiv32_fs766_xor0;
  assign f_arrdiv32_fs766_not1 = ~f_arrdiv32_fs766_xor0;
  assign f_arrdiv32_fs766_and1 = f_arrdiv32_fs766_not1 & f_arrdiv32_fs765_or0;
  assign f_arrdiv32_fs766_or0 = f_arrdiv32_fs766_and1 | f_arrdiv32_fs766_and0;
  assign f_arrdiv32_fs767_xor0 = f_arrdiv32_mux2to1712_xor0 ^ b[31];
  assign f_arrdiv32_fs767_not0 = ~f_arrdiv32_mux2to1712_xor0;
  assign f_arrdiv32_fs767_and0 = f_arrdiv32_fs767_not0 & b[31];
  assign f_arrdiv32_fs767_xor1 = f_arrdiv32_fs766_or0 ^ f_arrdiv32_fs767_xor0;
  assign f_arrdiv32_fs767_not1 = ~f_arrdiv32_fs767_xor0;
  assign f_arrdiv32_fs767_and1 = f_arrdiv32_fs767_not1 & f_arrdiv32_fs766_or0;
  assign f_arrdiv32_fs767_or0 = f_arrdiv32_fs767_and1 | f_arrdiv32_fs767_and0;
  assign f_arrdiv32_mux2to1713_and0 = a[8] & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1713_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1713_and1 = f_arrdiv32_fs736_xor0 & f_arrdiv32_mux2to1713_not0;
  assign f_arrdiv32_mux2to1713_xor0 = f_arrdiv32_mux2to1713_and0 ^ f_arrdiv32_mux2to1713_and1;
  assign f_arrdiv32_mux2to1714_and0 = f_arrdiv32_mux2to1682_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1714_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1714_and1 = f_arrdiv32_fs737_xor1 & f_arrdiv32_mux2to1714_not0;
  assign f_arrdiv32_mux2to1714_xor0 = f_arrdiv32_mux2to1714_and0 ^ f_arrdiv32_mux2to1714_and1;
  assign f_arrdiv32_mux2to1715_and0 = f_arrdiv32_mux2to1683_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1715_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1715_and1 = f_arrdiv32_fs738_xor1 & f_arrdiv32_mux2to1715_not0;
  assign f_arrdiv32_mux2to1715_xor0 = f_arrdiv32_mux2to1715_and0 ^ f_arrdiv32_mux2to1715_and1;
  assign f_arrdiv32_mux2to1716_and0 = f_arrdiv32_mux2to1684_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1716_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1716_and1 = f_arrdiv32_fs739_xor1 & f_arrdiv32_mux2to1716_not0;
  assign f_arrdiv32_mux2to1716_xor0 = f_arrdiv32_mux2to1716_and0 ^ f_arrdiv32_mux2to1716_and1;
  assign f_arrdiv32_mux2to1717_and0 = f_arrdiv32_mux2to1685_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1717_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1717_and1 = f_arrdiv32_fs740_xor1 & f_arrdiv32_mux2to1717_not0;
  assign f_arrdiv32_mux2to1717_xor0 = f_arrdiv32_mux2to1717_and0 ^ f_arrdiv32_mux2to1717_and1;
  assign f_arrdiv32_mux2to1718_and0 = f_arrdiv32_mux2to1686_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1718_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1718_and1 = f_arrdiv32_fs741_xor1 & f_arrdiv32_mux2to1718_not0;
  assign f_arrdiv32_mux2to1718_xor0 = f_arrdiv32_mux2to1718_and0 ^ f_arrdiv32_mux2to1718_and1;
  assign f_arrdiv32_mux2to1719_and0 = f_arrdiv32_mux2to1687_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1719_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1719_and1 = f_arrdiv32_fs742_xor1 & f_arrdiv32_mux2to1719_not0;
  assign f_arrdiv32_mux2to1719_xor0 = f_arrdiv32_mux2to1719_and0 ^ f_arrdiv32_mux2to1719_and1;
  assign f_arrdiv32_mux2to1720_and0 = f_arrdiv32_mux2to1688_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1720_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1720_and1 = f_arrdiv32_fs743_xor1 & f_arrdiv32_mux2to1720_not0;
  assign f_arrdiv32_mux2to1720_xor0 = f_arrdiv32_mux2to1720_and0 ^ f_arrdiv32_mux2to1720_and1;
  assign f_arrdiv32_mux2to1721_and0 = f_arrdiv32_mux2to1689_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1721_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1721_and1 = f_arrdiv32_fs744_xor1 & f_arrdiv32_mux2to1721_not0;
  assign f_arrdiv32_mux2to1721_xor0 = f_arrdiv32_mux2to1721_and0 ^ f_arrdiv32_mux2to1721_and1;
  assign f_arrdiv32_mux2to1722_and0 = f_arrdiv32_mux2to1690_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1722_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1722_and1 = f_arrdiv32_fs745_xor1 & f_arrdiv32_mux2to1722_not0;
  assign f_arrdiv32_mux2to1722_xor0 = f_arrdiv32_mux2to1722_and0 ^ f_arrdiv32_mux2to1722_and1;
  assign f_arrdiv32_mux2to1723_and0 = f_arrdiv32_mux2to1691_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1723_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1723_and1 = f_arrdiv32_fs746_xor1 & f_arrdiv32_mux2to1723_not0;
  assign f_arrdiv32_mux2to1723_xor0 = f_arrdiv32_mux2to1723_and0 ^ f_arrdiv32_mux2to1723_and1;
  assign f_arrdiv32_mux2to1724_and0 = f_arrdiv32_mux2to1692_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1724_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1724_and1 = f_arrdiv32_fs747_xor1 & f_arrdiv32_mux2to1724_not0;
  assign f_arrdiv32_mux2to1724_xor0 = f_arrdiv32_mux2to1724_and0 ^ f_arrdiv32_mux2to1724_and1;
  assign f_arrdiv32_mux2to1725_and0 = f_arrdiv32_mux2to1693_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1725_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1725_and1 = f_arrdiv32_fs748_xor1 & f_arrdiv32_mux2to1725_not0;
  assign f_arrdiv32_mux2to1725_xor0 = f_arrdiv32_mux2to1725_and0 ^ f_arrdiv32_mux2to1725_and1;
  assign f_arrdiv32_mux2to1726_and0 = f_arrdiv32_mux2to1694_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1726_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1726_and1 = f_arrdiv32_fs749_xor1 & f_arrdiv32_mux2to1726_not0;
  assign f_arrdiv32_mux2to1726_xor0 = f_arrdiv32_mux2to1726_and0 ^ f_arrdiv32_mux2to1726_and1;
  assign f_arrdiv32_mux2to1727_and0 = f_arrdiv32_mux2to1695_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1727_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1727_and1 = f_arrdiv32_fs750_xor1 & f_arrdiv32_mux2to1727_not0;
  assign f_arrdiv32_mux2to1727_xor0 = f_arrdiv32_mux2to1727_and0 ^ f_arrdiv32_mux2to1727_and1;
  assign f_arrdiv32_mux2to1728_and0 = f_arrdiv32_mux2to1696_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1728_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1728_and1 = f_arrdiv32_fs751_xor1 & f_arrdiv32_mux2to1728_not0;
  assign f_arrdiv32_mux2to1728_xor0 = f_arrdiv32_mux2to1728_and0 ^ f_arrdiv32_mux2to1728_and1;
  assign f_arrdiv32_mux2to1729_and0 = f_arrdiv32_mux2to1697_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1729_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1729_and1 = f_arrdiv32_fs752_xor1 & f_arrdiv32_mux2to1729_not0;
  assign f_arrdiv32_mux2to1729_xor0 = f_arrdiv32_mux2to1729_and0 ^ f_arrdiv32_mux2to1729_and1;
  assign f_arrdiv32_mux2to1730_and0 = f_arrdiv32_mux2to1698_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1730_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1730_and1 = f_arrdiv32_fs753_xor1 & f_arrdiv32_mux2to1730_not0;
  assign f_arrdiv32_mux2to1730_xor0 = f_arrdiv32_mux2to1730_and0 ^ f_arrdiv32_mux2to1730_and1;
  assign f_arrdiv32_mux2to1731_and0 = f_arrdiv32_mux2to1699_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1731_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1731_and1 = f_arrdiv32_fs754_xor1 & f_arrdiv32_mux2to1731_not0;
  assign f_arrdiv32_mux2to1731_xor0 = f_arrdiv32_mux2to1731_and0 ^ f_arrdiv32_mux2to1731_and1;
  assign f_arrdiv32_mux2to1732_and0 = f_arrdiv32_mux2to1700_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1732_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1732_and1 = f_arrdiv32_fs755_xor1 & f_arrdiv32_mux2to1732_not0;
  assign f_arrdiv32_mux2to1732_xor0 = f_arrdiv32_mux2to1732_and0 ^ f_arrdiv32_mux2to1732_and1;
  assign f_arrdiv32_mux2to1733_and0 = f_arrdiv32_mux2to1701_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1733_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1733_and1 = f_arrdiv32_fs756_xor1 & f_arrdiv32_mux2to1733_not0;
  assign f_arrdiv32_mux2to1733_xor0 = f_arrdiv32_mux2to1733_and0 ^ f_arrdiv32_mux2to1733_and1;
  assign f_arrdiv32_mux2to1734_and0 = f_arrdiv32_mux2to1702_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1734_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1734_and1 = f_arrdiv32_fs757_xor1 & f_arrdiv32_mux2to1734_not0;
  assign f_arrdiv32_mux2to1734_xor0 = f_arrdiv32_mux2to1734_and0 ^ f_arrdiv32_mux2to1734_and1;
  assign f_arrdiv32_mux2to1735_and0 = f_arrdiv32_mux2to1703_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1735_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1735_and1 = f_arrdiv32_fs758_xor1 & f_arrdiv32_mux2to1735_not0;
  assign f_arrdiv32_mux2to1735_xor0 = f_arrdiv32_mux2to1735_and0 ^ f_arrdiv32_mux2to1735_and1;
  assign f_arrdiv32_mux2to1736_and0 = f_arrdiv32_mux2to1704_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1736_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1736_and1 = f_arrdiv32_fs759_xor1 & f_arrdiv32_mux2to1736_not0;
  assign f_arrdiv32_mux2to1736_xor0 = f_arrdiv32_mux2to1736_and0 ^ f_arrdiv32_mux2to1736_and1;
  assign f_arrdiv32_mux2to1737_and0 = f_arrdiv32_mux2to1705_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1737_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1737_and1 = f_arrdiv32_fs760_xor1 & f_arrdiv32_mux2to1737_not0;
  assign f_arrdiv32_mux2to1737_xor0 = f_arrdiv32_mux2to1737_and0 ^ f_arrdiv32_mux2to1737_and1;
  assign f_arrdiv32_mux2to1738_and0 = f_arrdiv32_mux2to1706_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1738_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1738_and1 = f_arrdiv32_fs761_xor1 & f_arrdiv32_mux2to1738_not0;
  assign f_arrdiv32_mux2to1738_xor0 = f_arrdiv32_mux2to1738_and0 ^ f_arrdiv32_mux2to1738_and1;
  assign f_arrdiv32_mux2to1739_and0 = f_arrdiv32_mux2to1707_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1739_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1739_and1 = f_arrdiv32_fs762_xor1 & f_arrdiv32_mux2to1739_not0;
  assign f_arrdiv32_mux2to1739_xor0 = f_arrdiv32_mux2to1739_and0 ^ f_arrdiv32_mux2to1739_and1;
  assign f_arrdiv32_mux2to1740_and0 = f_arrdiv32_mux2to1708_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1740_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1740_and1 = f_arrdiv32_fs763_xor1 & f_arrdiv32_mux2to1740_not0;
  assign f_arrdiv32_mux2to1740_xor0 = f_arrdiv32_mux2to1740_and0 ^ f_arrdiv32_mux2to1740_and1;
  assign f_arrdiv32_mux2to1741_and0 = f_arrdiv32_mux2to1709_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1741_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1741_and1 = f_arrdiv32_fs764_xor1 & f_arrdiv32_mux2to1741_not0;
  assign f_arrdiv32_mux2to1741_xor0 = f_arrdiv32_mux2to1741_and0 ^ f_arrdiv32_mux2to1741_and1;
  assign f_arrdiv32_mux2to1742_and0 = f_arrdiv32_mux2to1710_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1742_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1742_and1 = f_arrdiv32_fs765_xor1 & f_arrdiv32_mux2to1742_not0;
  assign f_arrdiv32_mux2to1742_xor0 = f_arrdiv32_mux2to1742_and0 ^ f_arrdiv32_mux2to1742_and1;
  assign f_arrdiv32_mux2to1743_and0 = f_arrdiv32_mux2to1711_xor0 & f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1743_not0 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_mux2to1743_and1 = f_arrdiv32_fs766_xor1 & f_arrdiv32_mux2to1743_not0;
  assign f_arrdiv32_mux2to1743_xor0 = f_arrdiv32_mux2to1743_and0 ^ f_arrdiv32_mux2to1743_and1;
  assign f_arrdiv32_not23 = ~f_arrdiv32_fs767_or0;
  assign f_arrdiv32_fs768_xor0 = a[7] ^ b[0];
  assign f_arrdiv32_fs768_not0 = ~a[7];
  assign f_arrdiv32_fs768_and0 = f_arrdiv32_fs768_not0 & b[0];
  assign f_arrdiv32_fs768_not1 = ~f_arrdiv32_fs768_xor0;
  assign f_arrdiv32_fs769_xor0 = f_arrdiv32_mux2to1713_xor0 ^ b[1];
  assign f_arrdiv32_fs769_not0 = ~f_arrdiv32_mux2to1713_xor0;
  assign f_arrdiv32_fs769_and0 = f_arrdiv32_fs769_not0 & b[1];
  assign f_arrdiv32_fs769_xor1 = f_arrdiv32_fs768_and0 ^ f_arrdiv32_fs769_xor0;
  assign f_arrdiv32_fs769_not1 = ~f_arrdiv32_fs769_xor0;
  assign f_arrdiv32_fs769_and1 = f_arrdiv32_fs769_not1 & f_arrdiv32_fs768_and0;
  assign f_arrdiv32_fs769_or0 = f_arrdiv32_fs769_and1 | f_arrdiv32_fs769_and0;
  assign f_arrdiv32_fs770_xor0 = f_arrdiv32_mux2to1714_xor0 ^ b[2];
  assign f_arrdiv32_fs770_not0 = ~f_arrdiv32_mux2to1714_xor0;
  assign f_arrdiv32_fs770_and0 = f_arrdiv32_fs770_not0 & b[2];
  assign f_arrdiv32_fs770_xor1 = f_arrdiv32_fs769_or0 ^ f_arrdiv32_fs770_xor0;
  assign f_arrdiv32_fs770_not1 = ~f_arrdiv32_fs770_xor0;
  assign f_arrdiv32_fs770_and1 = f_arrdiv32_fs770_not1 & f_arrdiv32_fs769_or0;
  assign f_arrdiv32_fs770_or0 = f_arrdiv32_fs770_and1 | f_arrdiv32_fs770_and0;
  assign f_arrdiv32_fs771_xor0 = f_arrdiv32_mux2to1715_xor0 ^ b[3];
  assign f_arrdiv32_fs771_not0 = ~f_arrdiv32_mux2to1715_xor0;
  assign f_arrdiv32_fs771_and0 = f_arrdiv32_fs771_not0 & b[3];
  assign f_arrdiv32_fs771_xor1 = f_arrdiv32_fs770_or0 ^ f_arrdiv32_fs771_xor0;
  assign f_arrdiv32_fs771_not1 = ~f_arrdiv32_fs771_xor0;
  assign f_arrdiv32_fs771_and1 = f_arrdiv32_fs771_not1 & f_arrdiv32_fs770_or0;
  assign f_arrdiv32_fs771_or0 = f_arrdiv32_fs771_and1 | f_arrdiv32_fs771_and0;
  assign f_arrdiv32_fs772_xor0 = f_arrdiv32_mux2to1716_xor0 ^ b[4];
  assign f_arrdiv32_fs772_not0 = ~f_arrdiv32_mux2to1716_xor0;
  assign f_arrdiv32_fs772_and0 = f_arrdiv32_fs772_not0 & b[4];
  assign f_arrdiv32_fs772_xor1 = f_arrdiv32_fs771_or0 ^ f_arrdiv32_fs772_xor0;
  assign f_arrdiv32_fs772_not1 = ~f_arrdiv32_fs772_xor0;
  assign f_arrdiv32_fs772_and1 = f_arrdiv32_fs772_not1 & f_arrdiv32_fs771_or0;
  assign f_arrdiv32_fs772_or0 = f_arrdiv32_fs772_and1 | f_arrdiv32_fs772_and0;
  assign f_arrdiv32_fs773_xor0 = f_arrdiv32_mux2to1717_xor0 ^ b[5];
  assign f_arrdiv32_fs773_not0 = ~f_arrdiv32_mux2to1717_xor0;
  assign f_arrdiv32_fs773_and0 = f_arrdiv32_fs773_not0 & b[5];
  assign f_arrdiv32_fs773_xor1 = f_arrdiv32_fs772_or0 ^ f_arrdiv32_fs773_xor0;
  assign f_arrdiv32_fs773_not1 = ~f_arrdiv32_fs773_xor0;
  assign f_arrdiv32_fs773_and1 = f_arrdiv32_fs773_not1 & f_arrdiv32_fs772_or0;
  assign f_arrdiv32_fs773_or0 = f_arrdiv32_fs773_and1 | f_arrdiv32_fs773_and0;
  assign f_arrdiv32_fs774_xor0 = f_arrdiv32_mux2to1718_xor0 ^ b[6];
  assign f_arrdiv32_fs774_not0 = ~f_arrdiv32_mux2to1718_xor0;
  assign f_arrdiv32_fs774_and0 = f_arrdiv32_fs774_not0 & b[6];
  assign f_arrdiv32_fs774_xor1 = f_arrdiv32_fs773_or0 ^ f_arrdiv32_fs774_xor0;
  assign f_arrdiv32_fs774_not1 = ~f_arrdiv32_fs774_xor0;
  assign f_arrdiv32_fs774_and1 = f_arrdiv32_fs774_not1 & f_arrdiv32_fs773_or0;
  assign f_arrdiv32_fs774_or0 = f_arrdiv32_fs774_and1 | f_arrdiv32_fs774_and0;
  assign f_arrdiv32_fs775_xor0 = f_arrdiv32_mux2to1719_xor0 ^ b[7];
  assign f_arrdiv32_fs775_not0 = ~f_arrdiv32_mux2to1719_xor0;
  assign f_arrdiv32_fs775_and0 = f_arrdiv32_fs775_not0 & b[7];
  assign f_arrdiv32_fs775_xor1 = f_arrdiv32_fs774_or0 ^ f_arrdiv32_fs775_xor0;
  assign f_arrdiv32_fs775_not1 = ~f_arrdiv32_fs775_xor0;
  assign f_arrdiv32_fs775_and1 = f_arrdiv32_fs775_not1 & f_arrdiv32_fs774_or0;
  assign f_arrdiv32_fs775_or0 = f_arrdiv32_fs775_and1 | f_arrdiv32_fs775_and0;
  assign f_arrdiv32_fs776_xor0 = f_arrdiv32_mux2to1720_xor0 ^ b[8];
  assign f_arrdiv32_fs776_not0 = ~f_arrdiv32_mux2to1720_xor0;
  assign f_arrdiv32_fs776_and0 = f_arrdiv32_fs776_not0 & b[8];
  assign f_arrdiv32_fs776_xor1 = f_arrdiv32_fs775_or0 ^ f_arrdiv32_fs776_xor0;
  assign f_arrdiv32_fs776_not1 = ~f_arrdiv32_fs776_xor0;
  assign f_arrdiv32_fs776_and1 = f_arrdiv32_fs776_not1 & f_arrdiv32_fs775_or0;
  assign f_arrdiv32_fs776_or0 = f_arrdiv32_fs776_and1 | f_arrdiv32_fs776_and0;
  assign f_arrdiv32_fs777_xor0 = f_arrdiv32_mux2to1721_xor0 ^ b[9];
  assign f_arrdiv32_fs777_not0 = ~f_arrdiv32_mux2to1721_xor0;
  assign f_arrdiv32_fs777_and0 = f_arrdiv32_fs777_not0 & b[9];
  assign f_arrdiv32_fs777_xor1 = f_arrdiv32_fs776_or0 ^ f_arrdiv32_fs777_xor0;
  assign f_arrdiv32_fs777_not1 = ~f_arrdiv32_fs777_xor0;
  assign f_arrdiv32_fs777_and1 = f_arrdiv32_fs777_not1 & f_arrdiv32_fs776_or0;
  assign f_arrdiv32_fs777_or0 = f_arrdiv32_fs777_and1 | f_arrdiv32_fs777_and0;
  assign f_arrdiv32_fs778_xor0 = f_arrdiv32_mux2to1722_xor0 ^ b[10];
  assign f_arrdiv32_fs778_not0 = ~f_arrdiv32_mux2to1722_xor0;
  assign f_arrdiv32_fs778_and0 = f_arrdiv32_fs778_not0 & b[10];
  assign f_arrdiv32_fs778_xor1 = f_arrdiv32_fs777_or0 ^ f_arrdiv32_fs778_xor0;
  assign f_arrdiv32_fs778_not1 = ~f_arrdiv32_fs778_xor0;
  assign f_arrdiv32_fs778_and1 = f_arrdiv32_fs778_not1 & f_arrdiv32_fs777_or0;
  assign f_arrdiv32_fs778_or0 = f_arrdiv32_fs778_and1 | f_arrdiv32_fs778_and0;
  assign f_arrdiv32_fs779_xor0 = f_arrdiv32_mux2to1723_xor0 ^ b[11];
  assign f_arrdiv32_fs779_not0 = ~f_arrdiv32_mux2to1723_xor0;
  assign f_arrdiv32_fs779_and0 = f_arrdiv32_fs779_not0 & b[11];
  assign f_arrdiv32_fs779_xor1 = f_arrdiv32_fs778_or0 ^ f_arrdiv32_fs779_xor0;
  assign f_arrdiv32_fs779_not1 = ~f_arrdiv32_fs779_xor0;
  assign f_arrdiv32_fs779_and1 = f_arrdiv32_fs779_not1 & f_arrdiv32_fs778_or0;
  assign f_arrdiv32_fs779_or0 = f_arrdiv32_fs779_and1 | f_arrdiv32_fs779_and0;
  assign f_arrdiv32_fs780_xor0 = f_arrdiv32_mux2to1724_xor0 ^ b[12];
  assign f_arrdiv32_fs780_not0 = ~f_arrdiv32_mux2to1724_xor0;
  assign f_arrdiv32_fs780_and0 = f_arrdiv32_fs780_not0 & b[12];
  assign f_arrdiv32_fs780_xor1 = f_arrdiv32_fs779_or0 ^ f_arrdiv32_fs780_xor0;
  assign f_arrdiv32_fs780_not1 = ~f_arrdiv32_fs780_xor0;
  assign f_arrdiv32_fs780_and1 = f_arrdiv32_fs780_not1 & f_arrdiv32_fs779_or0;
  assign f_arrdiv32_fs780_or0 = f_arrdiv32_fs780_and1 | f_arrdiv32_fs780_and0;
  assign f_arrdiv32_fs781_xor0 = f_arrdiv32_mux2to1725_xor0 ^ b[13];
  assign f_arrdiv32_fs781_not0 = ~f_arrdiv32_mux2to1725_xor0;
  assign f_arrdiv32_fs781_and0 = f_arrdiv32_fs781_not0 & b[13];
  assign f_arrdiv32_fs781_xor1 = f_arrdiv32_fs780_or0 ^ f_arrdiv32_fs781_xor0;
  assign f_arrdiv32_fs781_not1 = ~f_arrdiv32_fs781_xor0;
  assign f_arrdiv32_fs781_and1 = f_arrdiv32_fs781_not1 & f_arrdiv32_fs780_or0;
  assign f_arrdiv32_fs781_or0 = f_arrdiv32_fs781_and1 | f_arrdiv32_fs781_and0;
  assign f_arrdiv32_fs782_xor0 = f_arrdiv32_mux2to1726_xor0 ^ b[14];
  assign f_arrdiv32_fs782_not0 = ~f_arrdiv32_mux2to1726_xor0;
  assign f_arrdiv32_fs782_and0 = f_arrdiv32_fs782_not0 & b[14];
  assign f_arrdiv32_fs782_xor1 = f_arrdiv32_fs781_or0 ^ f_arrdiv32_fs782_xor0;
  assign f_arrdiv32_fs782_not1 = ~f_arrdiv32_fs782_xor0;
  assign f_arrdiv32_fs782_and1 = f_arrdiv32_fs782_not1 & f_arrdiv32_fs781_or0;
  assign f_arrdiv32_fs782_or0 = f_arrdiv32_fs782_and1 | f_arrdiv32_fs782_and0;
  assign f_arrdiv32_fs783_xor0 = f_arrdiv32_mux2to1727_xor0 ^ b[15];
  assign f_arrdiv32_fs783_not0 = ~f_arrdiv32_mux2to1727_xor0;
  assign f_arrdiv32_fs783_and0 = f_arrdiv32_fs783_not0 & b[15];
  assign f_arrdiv32_fs783_xor1 = f_arrdiv32_fs782_or0 ^ f_arrdiv32_fs783_xor0;
  assign f_arrdiv32_fs783_not1 = ~f_arrdiv32_fs783_xor0;
  assign f_arrdiv32_fs783_and1 = f_arrdiv32_fs783_not1 & f_arrdiv32_fs782_or0;
  assign f_arrdiv32_fs783_or0 = f_arrdiv32_fs783_and1 | f_arrdiv32_fs783_and0;
  assign f_arrdiv32_fs784_xor0 = f_arrdiv32_mux2to1728_xor0 ^ b[16];
  assign f_arrdiv32_fs784_not0 = ~f_arrdiv32_mux2to1728_xor0;
  assign f_arrdiv32_fs784_and0 = f_arrdiv32_fs784_not0 & b[16];
  assign f_arrdiv32_fs784_xor1 = f_arrdiv32_fs783_or0 ^ f_arrdiv32_fs784_xor0;
  assign f_arrdiv32_fs784_not1 = ~f_arrdiv32_fs784_xor0;
  assign f_arrdiv32_fs784_and1 = f_arrdiv32_fs784_not1 & f_arrdiv32_fs783_or0;
  assign f_arrdiv32_fs784_or0 = f_arrdiv32_fs784_and1 | f_arrdiv32_fs784_and0;
  assign f_arrdiv32_fs785_xor0 = f_arrdiv32_mux2to1729_xor0 ^ b[17];
  assign f_arrdiv32_fs785_not0 = ~f_arrdiv32_mux2to1729_xor0;
  assign f_arrdiv32_fs785_and0 = f_arrdiv32_fs785_not0 & b[17];
  assign f_arrdiv32_fs785_xor1 = f_arrdiv32_fs784_or0 ^ f_arrdiv32_fs785_xor0;
  assign f_arrdiv32_fs785_not1 = ~f_arrdiv32_fs785_xor0;
  assign f_arrdiv32_fs785_and1 = f_arrdiv32_fs785_not1 & f_arrdiv32_fs784_or0;
  assign f_arrdiv32_fs785_or0 = f_arrdiv32_fs785_and1 | f_arrdiv32_fs785_and0;
  assign f_arrdiv32_fs786_xor0 = f_arrdiv32_mux2to1730_xor0 ^ b[18];
  assign f_arrdiv32_fs786_not0 = ~f_arrdiv32_mux2to1730_xor0;
  assign f_arrdiv32_fs786_and0 = f_arrdiv32_fs786_not0 & b[18];
  assign f_arrdiv32_fs786_xor1 = f_arrdiv32_fs785_or0 ^ f_arrdiv32_fs786_xor0;
  assign f_arrdiv32_fs786_not1 = ~f_arrdiv32_fs786_xor0;
  assign f_arrdiv32_fs786_and1 = f_arrdiv32_fs786_not1 & f_arrdiv32_fs785_or0;
  assign f_arrdiv32_fs786_or0 = f_arrdiv32_fs786_and1 | f_arrdiv32_fs786_and0;
  assign f_arrdiv32_fs787_xor0 = f_arrdiv32_mux2to1731_xor0 ^ b[19];
  assign f_arrdiv32_fs787_not0 = ~f_arrdiv32_mux2to1731_xor0;
  assign f_arrdiv32_fs787_and0 = f_arrdiv32_fs787_not0 & b[19];
  assign f_arrdiv32_fs787_xor1 = f_arrdiv32_fs786_or0 ^ f_arrdiv32_fs787_xor0;
  assign f_arrdiv32_fs787_not1 = ~f_arrdiv32_fs787_xor0;
  assign f_arrdiv32_fs787_and1 = f_arrdiv32_fs787_not1 & f_arrdiv32_fs786_or0;
  assign f_arrdiv32_fs787_or0 = f_arrdiv32_fs787_and1 | f_arrdiv32_fs787_and0;
  assign f_arrdiv32_fs788_xor0 = f_arrdiv32_mux2to1732_xor0 ^ b[20];
  assign f_arrdiv32_fs788_not0 = ~f_arrdiv32_mux2to1732_xor0;
  assign f_arrdiv32_fs788_and0 = f_arrdiv32_fs788_not0 & b[20];
  assign f_arrdiv32_fs788_xor1 = f_arrdiv32_fs787_or0 ^ f_arrdiv32_fs788_xor0;
  assign f_arrdiv32_fs788_not1 = ~f_arrdiv32_fs788_xor0;
  assign f_arrdiv32_fs788_and1 = f_arrdiv32_fs788_not1 & f_arrdiv32_fs787_or0;
  assign f_arrdiv32_fs788_or0 = f_arrdiv32_fs788_and1 | f_arrdiv32_fs788_and0;
  assign f_arrdiv32_fs789_xor0 = f_arrdiv32_mux2to1733_xor0 ^ b[21];
  assign f_arrdiv32_fs789_not0 = ~f_arrdiv32_mux2to1733_xor0;
  assign f_arrdiv32_fs789_and0 = f_arrdiv32_fs789_not0 & b[21];
  assign f_arrdiv32_fs789_xor1 = f_arrdiv32_fs788_or0 ^ f_arrdiv32_fs789_xor0;
  assign f_arrdiv32_fs789_not1 = ~f_arrdiv32_fs789_xor0;
  assign f_arrdiv32_fs789_and1 = f_arrdiv32_fs789_not1 & f_arrdiv32_fs788_or0;
  assign f_arrdiv32_fs789_or0 = f_arrdiv32_fs789_and1 | f_arrdiv32_fs789_and0;
  assign f_arrdiv32_fs790_xor0 = f_arrdiv32_mux2to1734_xor0 ^ b[22];
  assign f_arrdiv32_fs790_not0 = ~f_arrdiv32_mux2to1734_xor0;
  assign f_arrdiv32_fs790_and0 = f_arrdiv32_fs790_not0 & b[22];
  assign f_arrdiv32_fs790_xor1 = f_arrdiv32_fs789_or0 ^ f_arrdiv32_fs790_xor0;
  assign f_arrdiv32_fs790_not1 = ~f_arrdiv32_fs790_xor0;
  assign f_arrdiv32_fs790_and1 = f_arrdiv32_fs790_not1 & f_arrdiv32_fs789_or0;
  assign f_arrdiv32_fs790_or0 = f_arrdiv32_fs790_and1 | f_arrdiv32_fs790_and0;
  assign f_arrdiv32_fs791_xor0 = f_arrdiv32_mux2to1735_xor0 ^ b[23];
  assign f_arrdiv32_fs791_not0 = ~f_arrdiv32_mux2to1735_xor0;
  assign f_arrdiv32_fs791_and0 = f_arrdiv32_fs791_not0 & b[23];
  assign f_arrdiv32_fs791_xor1 = f_arrdiv32_fs790_or0 ^ f_arrdiv32_fs791_xor0;
  assign f_arrdiv32_fs791_not1 = ~f_arrdiv32_fs791_xor0;
  assign f_arrdiv32_fs791_and1 = f_arrdiv32_fs791_not1 & f_arrdiv32_fs790_or0;
  assign f_arrdiv32_fs791_or0 = f_arrdiv32_fs791_and1 | f_arrdiv32_fs791_and0;
  assign f_arrdiv32_fs792_xor0 = f_arrdiv32_mux2to1736_xor0 ^ b[24];
  assign f_arrdiv32_fs792_not0 = ~f_arrdiv32_mux2to1736_xor0;
  assign f_arrdiv32_fs792_and0 = f_arrdiv32_fs792_not0 & b[24];
  assign f_arrdiv32_fs792_xor1 = f_arrdiv32_fs791_or0 ^ f_arrdiv32_fs792_xor0;
  assign f_arrdiv32_fs792_not1 = ~f_arrdiv32_fs792_xor0;
  assign f_arrdiv32_fs792_and1 = f_arrdiv32_fs792_not1 & f_arrdiv32_fs791_or0;
  assign f_arrdiv32_fs792_or0 = f_arrdiv32_fs792_and1 | f_arrdiv32_fs792_and0;
  assign f_arrdiv32_fs793_xor0 = f_arrdiv32_mux2to1737_xor0 ^ b[25];
  assign f_arrdiv32_fs793_not0 = ~f_arrdiv32_mux2to1737_xor0;
  assign f_arrdiv32_fs793_and0 = f_arrdiv32_fs793_not0 & b[25];
  assign f_arrdiv32_fs793_xor1 = f_arrdiv32_fs792_or0 ^ f_arrdiv32_fs793_xor0;
  assign f_arrdiv32_fs793_not1 = ~f_arrdiv32_fs793_xor0;
  assign f_arrdiv32_fs793_and1 = f_arrdiv32_fs793_not1 & f_arrdiv32_fs792_or0;
  assign f_arrdiv32_fs793_or0 = f_arrdiv32_fs793_and1 | f_arrdiv32_fs793_and0;
  assign f_arrdiv32_fs794_xor0 = f_arrdiv32_mux2to1738_xor0 ^ b[26];
  assign f_arrdiv32_fs794_not0 = ~f_arrdiv32_mux2to1738_xor0;
  assign f_arrdiv32_fs794_and0 = f_arrdiv32_fs794_not0 & b[26];
  assign f_arrdiv32_fs794_xor1 = f_arrdiv32_fs793_or0 ^ f_arrdiv32_fs794_xor0;
  assign f_arrdiv32_fs794_not1 = ~f_arrdiv32_fs794_xor0;
  assign f_arrdiv32_fs794_and1 = f_arrdiv32_fs794_not1 & f_arrdiv32_fs793_or0;
  assign f_arrdiv32_fs794_or0 = f_arrdiv32_fs794_and1 | f_arrdiv32_fs794_and0;
  assign f_arrdiv32_fs795_xor0 = f_arrdiv32_mux2to1739_xor0 ^ b[27];
  assign f_arrdiv32_fs795_not0 = ~f_arrdiv32_mux2to1739_xor0;
  assign f_arrdiv32_fs795_and0 = f_arrdiv32_fs795_not0 & b[27];
  assign f_arrdiv32_fs795_xor1 = f_arrdiv32_fs794_or0 ^ f_arrdiv32_fs795_xor0;
  assign f_arrdiv32_fs795_not1 = ~f_arrdiv32_fs795_xor0;
  assign f_arrdiv32_fs795_and1 = f_arrdiv32_fs795_not1 & f_arrdiv32_fs794_or0;
  assign f_arrdiv32_fs795_or0 = f_arrdiv32_fs795_and1 | f_arrdiv32_fs795_and0;
  assign f_arrdiv32_fs796_xor0 = f_arrdiv32_mux2to1740_xor0 ^ b[28];
  assign f_arrdiv32_fs796_not0 = ~f_arrdiv32_mux2to1740_xor0;
  assign f_arrdiv32_fs796_and0 = f_arrdiv32_fs796_not0 & b[28];
  assign f_arrdiv32_fs796_xor1 = f_arrdiv32_fs795_or0 ^ f_arrdiv32_fs796_xor0;
  assign f_arrdiv32_fs796_not1 = ~f_arrdiv32_fs796_xor0;
  assign f_arrdiv32_fs796_and1 = f_arrdiv32_fs796_not1 & f_arrdiv32_fs795_or0;
  assign f_arrdiv32_fs796_or0 = f_arrdiv32_fs796_and1 | f_arrdiv32_fs796_and0;
  assign f_arrdiv32_fs797_xor0 = f_arrdiv32_mux2to1741_xor0 ^ b[29];
  assign f_arrdiv32_fs797_not0 = ~f_arrdiv32_mux2to1741_xor0;
  assign f_arrdiv32_fs797_and0 = f_arrdiv32_fs797_not0 & b[29];
  assign f_arrdiv32_fs797_xor1 = f_arrdiv32_fs796_or0 ^ f_arrdiv32_fs797_xor0;
  assign f_arrdiv32_fs797_not1 = ~f_arrdiv32_fs797_xor0;
  assign f_arrdiv32_fs797_and1 = f_arrdiv32_fs797_not1 & f_arrdiv32_fs796_or0;
  assign f_arrdiv32_fs797_or0 = f_arrdiv32_fs797_and1 | f_arrdiv32_fs797_and0;
  assign f_arrdiv32_fs798_xor0 = f_arrdiv32_mux2to1742_xor0 ^ b[30];
  assign f_arrdiv32_fs798_not0 = ~f_arrdiv32_mux2to1742_xor0;
  assign f_arrdiv32_fs798_and0 = f_arrdiv32_fs798_not0 & b[30];
  assign f_arrdiv32_fs798_xor1 = f_arrdiv32_fs797_or0 ^ f_arrdiv32_fs798_xor0;
  assign f_arrdiv32_fs798_not1 = ~f_arrdiv32_fs798_xor0;
  assign f_arrdiv32_fs798_and1 = f_arrdiv32_fs798_not1 & f_arrdiv32_fs797_or0;
  assign f_arrdiv32_fs798_or0 = f_arrdiv32_fs798_and1 | f_arrdiv32_fs798_and0;
  assign f_arrdiv32_fs799_xor0 = f_arrdiv32_mux2to1743_xor0 ^ b[31];
  assign f_arrdiv32_fs799_not0 = ~f_arrdiv32_mux2to1743_xor0;
  assign f_arrdiv32_fs799_and0 = f_arrdiv32_fs799_not0 & b[31];
  assign f_arrdiv32_fs799_xor1 = f_arrdiv32_fs798_or0 ^ f_arrdiv32_fs799_xor0;
  assign f_arrdiv32_fs799_not1 = ~f_arrdiv32_fs799_xor0;
  assign f_arrdiv32_fs799_and1 = f_arrdiv32_fs799_not1 & f_arrdiv32_fs798_or0;
  assign f_arrdiv32_fs799_or0 = f_arrdiv32_fs799_and1 | f_arrdiv32_fs799_and0;
  assign f_arrdiv32_mux2to1744_and0 = a[7] & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1744_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1744_and1 = f_arrdiv32_fs768_xor0 & f_arrdiv32_mux2to1744_not0;
  assign f_arrdiv32_mux2to1744_xor0 = f_arrdiv32_mux2to1744_and0 ^ f_arrdiv32_mux2to1744_and1;
  assign f_arrdiv32_mux2to1745_and0 = f_arrdiv32_mux2to1713_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1745_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1745_and1 = f_arrdiv32_fs769_xor1 & f_arrdiv32_mux2to1745_not0;
  assign f_arrdiv32_mux2to1745_xor0 = f_arrdiv32_mux2to1745_and0 ^ f_arrdiv32_mux2to1745_and1;
  assign f_arrdiv32_mux2to1746_and0 = f_arrdiv32_mux2to1714_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1746_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1746_and1 = f_arrdiv32_fs770_xor1 & f_arrdiv32_mux2to1746_not0;
  assign f_arrdiv32_mux2to1746_xor0 = f_arrdiv32_mux2to1746_and0 ^ f_arrdiv32_mux2to1746_and1;
  assign f_arrdiv32_mux2to1747_and0 = f_arrdiv32_mux2to1715_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1747_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1747_and1 = f_arrdiv32_fs771_xor1 & f_arrdiv32_mux2to1747_not0;
  assign f_arrdiv32_mux2to1747_xor0 = f_arrdiv32_mux2to1747_and0 ^ f_arrdiv32_mux2to1747_and1;
  assign f_arrdiv32_mux2to1748_and0 = f_arrdiv32_mux2to1716_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1748_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1748_and1 = f_arrdiv32_fs772_xor1 & f_arrdiv32_mux2to1748_not0;
  assign f_arrdiv32_mux2to1748_xor0 = f_arrdiv32_mux2to1748_and0 ^ f_arrdiv32_mux2to1748_and1;
  assign f_arrdiv32_mux2to1749_and0 = f_arrdiv32_mux2to1717_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1749_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1749_and1 = f_arrdiv32_fs773_xor1 & f_arrdiv32_mux2to1749_not0;
  assign f_arrdiv32_mux2to1749_xor0 = f_arrdiv32_mux2to1749_and0 ^ f_arrdiv32_mux2to1749_and1;
  assign f_arrdiv32_mux2to1750_and0 = f_arrdiv32_mux2to1718_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1750_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1750_and1 = f_arrdiv32_fs774_xor1 & f_arrdiv32_mux2to1750_not0;
  assign f_arrdiv32_mux2to1750_xor0 = f_arrdiv32_mux2to1750_and0 ^ f_arrdiv32_mux2to1750_and1;
  assign f_arrdiv32_mux2to1751_and0 = f_arrdiv32_mux2to1719_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1751_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1751_and1 = f_arrdiv32_fs775_xor1 & f_arrdiv32_mux2to1751_not0;
  assign f_arrdiv32_mux2to1751_xor0 = f_arrdiv32_mux2to1751_and0 ^ f_arrdiv32_mux2to1751_and1;
  assign f_arrdiv32_mux2to1752_and0 = f_arrdiv32_mux2to1720_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1752_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1752_and1 = f_arrdiv32_fs776_xor1 & f_arrdiv32_mux2to1752_not0;
  assign f_arrdiv32_mux2to1752_xor0 = f_arrdiv32_mux2to1752_and0 ^ f_arrdiv32_mux2to1752_and1;
  assign f_arrdiv32_mux2to1753_and0 = f_arrdiv32_mux2to1721_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1753_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1753_and1 = f_arrdiv32_fs777_xor1 & f_arrdiv32_mux2to1753_not0;
  assign f_arrdiv32_mux2to1753_xor0 = f_arrdiv32_mux2to1753_and0 ^ f_arrdiv32_mux2to1753_and1;
  assign f_arrdiv32_mux2to1754_and0 = f_arrdiv32_mux2to1722_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1754_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1754_and1 = f_arrdiv32_fs778_xor1 & f_arrdiv32_mux2to1754_not0;
  assign f_arrdiv32_mux2to1754_xor0 = f_arrdiv32_mux2to1754_and0 ^ f_arrdiv32_mux2to1754_and1;
  assign f_arrdiv32_mux2to1755_and0 = f_arrdiv32_mux2to1723_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1755_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1755_and1 = f_arrdiv32_fs779_xor1 & f_arrdiv32_mux2to1755_not0;
  assign f_arrdiv32_mux2to1755_xor0 = f_arrdiv32_mux2to1755_and0 ^ f_arrdiv32_mux2to1755_and1;
  assign f_arrdiv32_mux2to1756_and0 = f_arrdiv32_mux2to1724_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1756_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1756_and1 = f_arrdiv32_fs780_xor1 & f_arrdiv32_mux2to1756_not0;
  assign f_arrdiv32_mux2to1756_xor0 = f_arrdiv32_mux2to1756_and0 ^ f_arrdiv32_mux2to1756_and1;
  assign f_arrdiv32_mux2to1757_and0 = f_arrdiv32_mux2to1725_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1757_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1757_and1 = f_arrdiv32_fs781_xor1 & f_arrdiv32_mux2to1757_not0;
  assign f_arrdiv32_mux2to1757_xor0 = f_arrdiv32_mux2to1757_and0 ^ f_arrdiv32_mux2to1757_and1;
  assign f_arrdiv32_mux2to1758_and0 = f_arrdiv32_mux2to1726_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1758_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1758_and1 = f_arrdiv32_fs782_xor1 & f_arrdiv32_mux2to1758_not0;
  assign f_arrdiv32_mux2to1758_xor0 = f_arrdiv32_mux2to1758_and0 ^ f_arrdiv32_mux2to1758_and1;
  assign f_arrdiv32_mux2to1759_and0 = f_arrdiv32_mux2to1727_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1759_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1759_and1 = f_arrdiv32_fs783_xor1 & f_arrdiv32_mux2to1759_not0;
  assign f_arrdiv32_mux2to1759_xor0 = f_arrdiv32_mux2to1759_and0 ^ f_arrdiv32_mux2to1759_and1;
  assign f_arrdiv32_mux2to1760_and0 = f_arrdiv32_mux2to1728_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1760_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1760_and1 = f_arrdiv32_fs784_xor1 & f_arrdiv32_mux2to1760_not0;
  assign f_arrdiv32_mux2to1760_xor0 = f_arrdiv32_mux2to1760_and0 ^ f_arrdiv32_mux2to1760_and1;
  assign f_arrdiv32_mux2to1761_and0 = f_arrdiv32_mux2to1729_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1761_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1761_and1 = f_arrdiv32_fs785_xor1 & f_arrdiv32_mux2to1761_not0;
  assign f_arrdiv32_mux2to1761_xor0 = f_arrdiv32_mux2to1761_and0 ^ f_arrdiv32_mux2to1761_and1;
  assign f_arrdiv32_mux2to1762_and0 = f_arrdiv32_mux2to1730_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1762_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1762_and1 = f_arrdiv32_fs786_xor1 & f_arrdiv32_mux2to1762_not0;
  assign f_arrdiv32_mux2to1762_xor0 = f_arrdiv32_mux2to1762_and0 ^ f_arrdiv32_mux2to1762_and1;
  assign f_arrdiv32_mux2to1763_and0 = f_arrdiv32_mux2to1731_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1763_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1763_and1 = f_arrdiv32_fs787_xor1 & f_arrdiv32_mux2to1763_not0;
  assign f_arrdiv32_mux2to1763_xor0 = f_arrdiv32_mux2to1763_and0 ^ f_arrdiv32_mux2to1763_and1;
  assign f_arrdiv32_mux2to1764_and0 = f_arrdiv32_mux2to1732_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1764_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1764_and1 = f_arrdiv32_fs788_xor1 & f_arrdiv32_mux2to1764_not0;
  assign f_arrdiv32_mux2to1764_xor0 = f_arrdiv32_mux2to1764_and0 ^ f_arrdiv32_mux2to1764_and1;
  assign f_arrdiv32_mux2to1765_and0 = f_arrdiv32_mux2to1733_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1765_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1765_and1 = f_arrdiv32_fs789_xor1 & f_arrdiv32_mux2to1765_not0;
  assign f_arrdiv32_mux2to1765_xor0 = f_arrdiv32_mux2to1765_and0 ^ f_arrdiv32_mux2to1765_and1;
  assign f_arrdiv32_mux2to1766_and0 = f_arrdiv32_mux2to1734_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1766_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1766_and1 = f_arrdiv32_fs790_xor1 & f_arrdiv32_mux2to1766_not0;
  assign f_arrdiv32_mux2to1766_xor0 = f_arrdiv32_mux2to1766_and0 ^ f_arrdiv32_mux2to1766_and1;
  assign f_arrdiv32_mux2to1767_and0 = f_arrdiv32_mux2to1735_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1767_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1767_and1 = f_arrdiv32_fs791_xor1 & f_arrdiv32_mux2to1767_not0;
  assign f_arrdiv32_mux2to1767_xor0 = f_arrdiv32_mux2to1767_and0 ^ f_arrdiv32_mux2to1767_and1;
  assign f_arrdiv32_mux2to1768_and0 = f_arrdiv32_mux2to1736_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1768_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1768_and1 = f_arrdiv32_fs792_xor1 & f_arrdiv32_mux2to1768_not0;
  assign f_arrdiv32_mux2to1768_xor0 = f_arrdiv32_mux2to1768_and0 ^ f_arrdiv32_mux2to1768_and1;
  assign f_arrdiv32_mux2to1769_and0 = f_arrdiv32_mux2to1737_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1769_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1769_and1 = f_arrdiv32_fs793_xor1 & f_arrdiv32_mux2to1769_not0;
  assign f_arrdiv32_mux2to1769_xor0 = f_arrdiv32_mux2to1769_and0 ^ f_arrdiv32_mux2to1769_and1;
  assign f_arrdiv32_mux2to1770_and0 = f_arrdiv32_mux2to1738_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1770_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1770_and1 = f_arrdiv32_fs794_xor1 & f_arrdiv32_mux2to1770_not0;
  assign f_arrdiv32_mux2to1770_xor0 = f_arrdiv32_mux2to1770_and0 ^ f_arrdiv32_mux2to1770_and1;
  assign f_arrdiv32_mux2to1771_and0 = f_arrdiv32_mux2to1739_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1771_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1771_and1 = f_arrdiv32_fs795_xor1 & f_arrdiv32_mux2to1771_not0;
  assign f_arrdiv32_mux2to1771_xor0 = f_arrdiv32_mux2to1771_and0 ^ f_arrdiv32_mux2to1771_and1;
  assign f_arrdiv32_mux2to1772_and0 = f_arrdiv32_mux2to1740_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1772_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1772_and1 = f_arrdiv32_fs796_xor1 & f_arrdiv32_mux2to1772_not0;
  assign f_arrdiv32_mux2to1772_xor0 = f_arrdiv32_mux2to1772_and0 ^ f_arrdiv32_mux2to1772_and1;
  assign f_arrdiv32_mux2to1773_and0 = f_arrdiv32_mux2to1741_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1773_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1773_and1 = f_arrdiv32_fs797_xor1 & f_arrdiv32_mux2to1773_not0;
  assign f_arrdiv32_mux2to1773_xor0 = f_arrdiv32_mux2to1773_and0 ^ f_arrdiv32_mux2to1773_and1;
  assign f_arrdiv32_mux2to1774_and0 = f_arrdiv32_mux2to1742_xor0 & f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1774_not0 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_mux2to1774_and1 = f_arrdiv32_fs798_xor1 & f_arrdiv32_mux2to1774_not0;
  assign f_arrdiv32_mux2to1774_xor0 = f_arrdiv32_mux2to1774_and0 ^ f_arrdiv32_mux2to1774_and1;
  assign f_arrdiv32_not24 = ~f_arrdiv32_fs799_or0;
  assign f_arrdiv32_fs800_xor0 = a[6] ^ b[0];
  assign f_arrdiv32_fs800_not0 = ~a[6];
  assign f_arrdiv32_fs800_and0 = f_arrdiv32_fs800_not0 & b[0];
  assign f_arrdiv32_fs800_not1 = ~f_arrdiv32_fs800_xor0;
  assign f_arrdiv32_fs801_xor0 = f_arrdiv32_mux2to1744_xor0 ^ b[1];
  assign f_arrdiv32_fs801_not0 = ~f_arrdiv32_mux2to1744_xor0;
  assign f_arrdiv32_fs801_and0 = f_arrdiv32_fs801_not0 & b[1];
  assign f_arrdiv32_fs801_xor1 = f_arrdiv32_fs800_and0 ^ f_arrdiv32_fs801_xor0;
  assign f_arrdiv32_fs801_not1 = ~f_arrdiv32_fs801_xor0;
  assign f_arrdiv32_fs801_and1 = f_arrdiv32_fs801_not1 & f_arrdiv32_fs800_and0;
  assign f_arrdiv32_fs801_or0 = f_arrdiv32_fs801_and1 | f_arrdiv32_fs801_and0;
  assign f_arrdiv32_fs802_xor0 = f_arrdiv32_mux2to1745_xor0 ^ b[2];
  assign f_arrdiv32_fs802_not0 = ~f_arrdiv32_mux2to1745_xor0;
  assign f_arrdiv32_fs802_and0 = f_arrdiv32_fs802_not0 & b[2];
  assign f_arrdiv32_fs802_xor1 = f_arrdiv32_fs801_or0 ^ f_arrdiv32_fs802_xor0;
  assign f_arrdiv32_fs802_not1 = ~f_arrdiv32_fs802_xor0;
  assign f_arrdiv32_fs802_and1 = f_arrdiv32_fs802_not1 & f_arrdiv32_fs801_or0;
  assign f_arrdiv32_fs802_or0 = f_arrdiv32_fs802_and1 | f_arrdiv32_fs802_and0;
  assign f_arrdiv32_fs803_xor0 = f_arrdiv32_mux2to1746_xor0 ^ b[3];
  assign f_arrdiv32_fs803_not0 = ~f_arrdiv32_mux2to1746_xor0;
  assign f_arrdiv32_fs803_and0 = f_arrdiv32_fs803_not0 & b[3];
  assign f_arrdiv32_fs803_xor1 = f_arrdiv32_fs802_or0 ^ f_arrdiv32_fs803_xor0;
  assign f_arrdiv32_fs803_not1 = ~f_arrdiv32_fs803_xor0;
  assign f_arrdiv32_fs803_and1 = f_arrdiv32_fs803_not1 & f_arrdiv32_fs802_or0;
  assign f_arrdiv32_fs803_or0 = f_arrdiv32_fs803_and1 | f_arrdiv32_fs803_and0;
  assign f_arrdiv32_fs804_xor0 = f_arrdiv32_mux2to1747_xor0 ^ b[4];
  assign f_arrdiv32_fs804_not0 = ~f_arrdiv32_mux2to1747_xor0;
  assign f_arrdiv32_fs804_and0 = f_arrdiv32_fs804_not0 & b[4];
  assign f_arrdiv32_fs804_xor1 = f_arrdiv32_fs803_or0 ^ f_arrdiv32_fs804_xor0;
  assign f_arrdiv32_fs804_not1 = ~f_arrdiv32_fs804_xor0;
  assign f_arrdiv32_fs804_and1 = f_arrdiv32_fs804_not1 & f_arrdiv32_fs803_or0;
  assign f_arrdiv32_fs804_or0 = f_arrdiv32_fs804_and1 | f_arrdiv32_fs804_and0;
  assign f_arrdiv32_fs805_xor0 = f_arrdiv32_mux2to1748_xor0 ^ b[5];
  assign f_arrdiv32_fs805_not0 = ~f_arrdiv32_mux2to1748_xor0;
  assign f_arrdiv32_fs805_and0 = f_arrdiv32_fs805_not0 & b[5];
  assign f_arrdiv32_fs805_xor1 = f_arrdiv32_fs804_or0 ^ f_arrdiv32_fs805_xor0;
  assign f_arrdiv32_fs805_not1 = ~f_arrdiv32_fs805_xor0;
  assign f_arrdiv32_fs805_and1 = f_arrdiv32_fs805_not1 & f_arrdiv32_fs804_or0;
  assign f_arrdiv32_fs805_or0 = f_arrdiv32_fs805_and1 | f_arrdiv32_fs805_and0;
  assign f_arrdiv32_fs806_xor0 = f_arrdiv32_mux2to1749_xor0 ^ b[6];
  assign f_arrdiv32_fs806_not0 = ~f_arrdiv32_mux2to1749_xor0;
  assign f_arrdiv32_fs806_and0 = f_arrdiv32_fs806_not0 & b[6];
  assign f_arrdiv32_fs806_xor1 = f_arrdiv32_fs805_or0 ^ f_arrdiv32_fs806_xor0;
  assign f_arrdiv32_fs806_not1 = ~f_arrdiv32_fs806_xor0;
  assign f_arrdiv32_fs806_and1 = f_arrdiv32_fs806_not1 & f_arrdiv32_fs805_or0;
  assign f_arrdiv32_fs806_or0 = f_arrdiv32_fs806_and1 | f_arrdiv32_fs806_and0;
  assign f_arrdiv32_fs807_xor0 = f_arrdiv32_mux2to1750_xor0 ^ b[7];
  assign f_arrdiv32_fs807_not0 = ~f_arrdiv32_mux2to1750_xor0;
  assign f_arrdiv32_fs807_and0 = f_arrdiv32_fs807_not0 & b[7];
  assign f_arrdiv32_fs807_xor1 = f_arrdiv32_fs806_or0 ^ f_arrdiv32_fs807_xor0;
  assign f_arrdiv32_fs807_not1 = ~f_arrdiv32_fs807_xor0;
  assign f_arrdiv32_fs807_and1 = f_arrdiv32_fs807_not1 & f_arrdiv32_fs806_or0;
  assign f_arrdiv32_fs807_or0 = f_arrdiv32_fs807_and1 | f_arrdiv32_fs807_and0;
  assign f_arrdiv32_fs808_xor0 = f_arrdiv32_mux2to1751_xor0 ^ b[8];
  assign f_arrdiv32_fs808_not0 = ~f_arrdiv32_mux2to1751_xor0;
  assign f_arrdiv32_fs808_and0 = f_arrdiv32_fs808_not0 & b[8];
  assign f_arrdiv32_fs808_xor1 = f_arrdiv32_fs807_or0 ^ f_arrdiv32_fs808_xor0;
  assign f_arrdiv32_fs808_not1 = ~f_arrdiv32_fs808_xor0;
  assign f_arrdiv32_fs808_and1 = f_arrdiv32_fs808_not1 & f_arrdiv32_fs807_or0;
  assign f_arrdiv32_fs808_or0 = f_arrdiv32_fs808_and1 | f_arrdiv32_fs808_and0;
  assign f_arrdiv32_fs809_xor0 = f_arrdiv32_mux2to1752_xor0 ^ b[9];
  assign f_arrdiv32_fs809_not0 = ~f_arrdiv32_mux2to1752_xor0;
  assign f_arrdiv32_fs809_and0 = f_arrdiv32_fs809_not0 & b[9];
  assign f_arrdiv32_fs809_xor1 = f_arrdiv32_fs808_or0 ^ f_arrdiv32_fs809_xor0;
  assign f_arrdiv32_fs809_not1 = ~f_arrdiv32_fs809_xor0;
  assign f_arrdiv32_fs809_and1 = f_arrdiv32_fs809_not1 & f_arrdiv32_fs808_or0;
  assign f_arrdiv32_fs809_or0 = f_arrdiv32_fs809_and1 | f_arrdiv32_fs809_and0;
  assign f_arrdiv32_fs810_xor0 = f_arrdiv32_mux2to1753_xor0 ^ b[10];
  assign f_arrdiv32_fs810_not0 = ~f_arrdiv32_mux2to1753_xor0;
  assign f_arrdiv32_fs810_and0 = f_arrdiv32_fs810_not0 & b[10];
  assign f_arrdiv32_fs810_xor1 = f_arrdiv32_fs809_or0 ^ f_arrdiv32_fs810_xor0;
  assign f_arrdiv32_fs810_not1 = ~f_arrdiv32_fs810_xor0;
  assign f_arrdiv32_fs810_and1 = f_arrdiv32_fs810_not1 & f_arrdiv32_fs809_or0;
  assign f_arrdiv32_fs810_or0 = f_arrdiv32_fs810_and1 | f_arrdiv32_fs810_and0;
  assign f_arrdiv32_fs811_xor0 = f_arrdiv32_mux2to1754_xor0 ^ b[11];
  assign f_arrdiv32_fs811_not0 = ~f_arrdiv32_mux2to1754_xor0;
  assign f_arrdiv32_fs811_and0 = f_arrdiv32_fs811_not0 & b[11];
  assign f_arrdiv32_fs811_xor1 = f_arrdiv32_fs810_or0 ^ f_arrdiv32_fs811_xor0;
  assign f_arrdiv32_fs811_not1 = ~f_arrdiv32_fs811_xor0;
  assign f_arrdiv32_fs811_and1 = f_arrdiv32_fs811_not1 & f_arrdiv32_fs810_or0;
  assign f_arrdiv32_fs811_or0 = f_arrdiv32_fs811_and1 | f_arrdiv32_fs811_and0;
  assign f_arrdiv32_fs812_xor0 = f_arrdiv32_mux2to1755_xor0 ^ b[12];
  assign f_arrdiv32_fs812_not0 = ~f_arrdiv32_mux2to1755_xor0;
  assign f_arrdiv32_fs812_and0 = f_arrdiv32_fs812_not0 & b[12];
  assign f_arrdiv32_fs812_xor1 = f_arrdiv32_fs811_or0 ^ f_arrdiv32_fs812_xor0;
  assign f_arrdiv32_fs812_not1 = ~f_arrdiv32_fs812_xor0;
  assign f_arrdiv32_fs812_and1 = f_arrdiv32_fs812_not1 & f_arrdiv32_fs811_or0;
  assign f_arrdiv32_fs812_or0 = f_arrdiv32_fs812_and1 | f_arrdiv32_fs812_and0;
  assign f_arrdiv32_fs813_xor0 = f_arrdiv32_mux2to1756_xor0 ^ b[13];
  assign f_arrdiv32_fs813_not0 = ~f_arrdiv32_mux2to1756_xor0;
  assign f_arrdiv32_fs813_and0 = f_arrdiv32_fs813_not0 & b[13];
  assign f_arrdiv32_fs813_xor1 = f_arrdiv32_fs812_or0 ^ f_arrdiv32_fs813_xor0;
  assign f_arrdiv32_fs813_not1 = ~f_arrdiv32_fs813_xor0;
  assign f_arrdiv32_fs813_and1 = f_arrdiv32_fs813_not1 & f_arrdiv32_fs812_or0;
  assign f_arrdiv32_fs813_or0 = f_arrdiv32_fs813_and1 | f_arrdiv32_fs813_and0;
  assign f_arrdiv32_fs814_xor0 = f_arrdiv32_mux2to1757_xor0 ^ b[14];
  assign f_arrdiv32_fs814_not0 = ~f_arrdiv32_mux2to1757_xor0;
  assign f_arrdiv32_fs814_and0 = f_arrdiv32_fs814_not0 & b[14];
  assign f_arrdiv32_fs814_xor1 = f_arrdiv32_fs813_or0 ^ f_arrdiv32_fs814_xor0;
  assign f_arrdiv32_fs814_not1 = ~f_arrdiv32_fs814_xor0;
  assign f_arrdiv32_fs814_and1 = f_arrdiv32_fs814_not1 & f_arrdiv32_fs813_or0;
  assign f_arrdiv32_fs814_or0 = f_arrdiv32_fs814_and1 | f_arrdiv32_fs814_and0;
  assign f_arrdiv32_fs815_xor0 = f_arrdiv32_mux2to1758_xor0 ^ b[15];
  assign f_arrdiv32_fs815_not0 = ~f_arrdiv32_mux2to1758_xor0;
  assign f_arrdiv32_fs815_and0 = f_arrdiv32_fs815_not0 & b[15];
  assign f_arrdiv32_fs815_xor1 = f_arrdiv32_fs814_or0 ^ f_arrdiv32_fs815_xor0;
  assign f_arrdiv32_fs815_not1 = ~f_arrdiv32_fs815_xor0;
  assign f_arrdiv32_fs815_and1 = f_arrdiv32_fs815_not1 & f_arrdiv32_fs814_or0;
  assign f_arrdiv32_fs815_or0 = f_arrdiv32_fs815_and1 | f_arrdiv32_fs815_and0;
  assign f_arrdiv32_fs816_xor0 = f_arrdiv32_mux2to1759_xor0 ^ b[16];
  assign f_arrdiv32_fs816_not0 = ~f_arrdiv32_mux2to1759_xor0;
  assign f_arrdiv32_fs816_and0 = f_arrdiv32_fs816_not0 & b[16];
  assign f_arrdiv32_fs816_xor1 = f_arrdiv32_fs815_or0 ^ f_arrdiv32_fs816_xor0;
  assign f_arrdiv32_fs816_not1 = ~f_arrdiv32_fs816_xor0;
  assign f_arrdiv32_fs816_and1 = f_arrdiv32_fs816_not1 & f_arrdiv32_fs815_or0;
  assign f_arrdiv32_fs816_or0 = f_arrdiv32_fs816_and1 | f_arrdiv32_fs816_and0;
  assign f_arrdiv32_fs817_xor0 = f_arrdiv32_mux2to1760_xor0 ^ b[17];
  assign f_arrdiv32_fs817_not0 = ~f_arrdiv32_mux2to1760_xor0;
  assign f_arrdiv32_fs817_and0 = f_arrdiv32_fs817_not0 & b[17];
  assign f_arrdiv32_fs817_xor1 = f_arrdiv32_fs816_or0 ^ f_arrdiv32_fs817_xor0;
  assign f_arrdiv32_fs817_not1 = ~f_arrdiv32_fs817_xor0;
  assign f_arrdiv32_fs817_and1 = f_arrdiv32_fs817_not1 & f_arrdiv32_fs816_or0;
  assign f_arrdiv32_fs817_or0 = f_arrdiv32_fs817_and1 | f_arrdiv32_fs817_and0;
  assign f_arrdiv32_fs818_xor0 = f_arrdiv32_mux2to1761_xor0 ^ b[18];
  assign f_arrdiv32_fs818_not0 = ~f_arrdiv32_mux2to1761_xor0;
  assign f_arrdiv32_fs818_and0 = f_arrdiv32_fs818_not0 & b[18];
  assign f_arrdiv32_fs818_xor1 = f_arrdiv32_fs817_or0 ^ f_arrdiv32_fs818_xor0;
  assign f_arrdiv32_fs818_not1 = ~f_arrdiv32_fs818_xor0;
  assign f_arrdiv32_fs818_and1 = f_arrdiv32_fs818_not1 & f_arrdiv32_fs817_or0;
  assign f_arrdiv32_fs818_or0 = f_arrdiv32_fs818_and1 | f_arrdiv32_fs818_and0;
  assign f_arrdiv32_fs819_xor0 = f_arrdiv32_mux2to1762_xor0 ^ b[19];
  assign f_arrdiv32_fs819_not0 = ~f_arrdiv32_mux2to1762_xor0;
  assign f_arrdiv32_fs819_and0 = f_arrdiv32_fs819_not0 & b[19];
  assign f_arrdiv32_fs819_xor1 = f_arrdiv32_fs818_or0 ^ f_arrdiv32_fs819_xor0;
  assign f_arrdiv32_fs819_not1 = ~f_arrdiv32_fs819_xor0;
  assign f_arrdiv32_fs819_and1 = f_arrdiv32_fs819_not1 & f_arrdiv32_fs818_or0;
  assign f_arrdiv32_fs819_or0 = f_arrdiv32_fs819_and1 | f_arrdiv32_fs819_and0;
  assign f_arrdiv32_fs820_xor0 = f_arrdiv32_mux2to1763_xor0 ^ b[20];
  assign f_arrdiv32_fs820_not0 = ~f_arrdiv32_mux2to1763_xor0;
  assign f_arrdiv32_fs820_and0 = f_arrdiv32_fs820_not0 & b[20];
  assign f_arrdiv32_fs820_xor1 = f_arrdiv32_fs819_or0 ^ f_arrdiv32_fs820_xor0;
  assign f_arrdiv32_fs820_not1 = ~f_arrdiv32_fs820_xor0;
  assign f_arrdiv32_fs820_and1 = f_arrdiv32_fs820_not1 & f_arrdiv32_fs819_or0;
  assign f_arrdiv32_fs820_or0 = f_arrdiv32_fs820_and1 | f_arrdiv32_fs820_and0;
  assign f_arrdiv32_fs821_xor0 = f_arrdiv32_mux2to1764_xor0 ^ b[21];
  assign f_arrdiv32_fs821_not0 = ~f_arrdiv32_mux2to1764_xor0;
  assign f_arrdiv32_fs821_and0 = f_arrdiv32_fs821_not0 & b[21];
  assign f_arrdiv32_fs821_xor1 = f_arrdiv32_fs820_or0 ^ f_arrdiv32_fs821_xor0;
  assign f_arrdiv32_fs821_not1 = ~f_arrdiv32_fs821_xor0;
  assign f_arrdiv32_fs821_and1 = f_arrdiv32_fs821_not1 & f_arrdiv32_fs820_or0;
  assign f_arrdiv32_fs821_or0 = f_arrdiv32_fs821_and1 | f_arrdiv32_fs821_and0;
  assign f_arrdiv32_fs822_xor0 = f_arrdiv32_mux2to1765_xor0 ^ b[22];
  assign f_arrdiv32_fs822_not0 = ~f_arrdiv32_mux2to1765_xor0;
  assign f_arrdiv32_fs822_and0 = f_arrdiv32_fs822_not0 & b[22];
  assign f_arrdiv32_fs822_xor1 = f_arrdiv32_fs821_or0 ^ f_arrdiv32_fs822_xor0;
  assign f_arrdiv32_fs822_not1 = ~f_arrdiv32_fs822_xor0;
  assign f_arrdiv32_fs822_and1 = f_arrdiv32_fs822_not1 & f_arrdiv32_fs821_or0;
  assign f_arrdiv32_fs822_or0 = f_arrdiv32_fs822_and1 | f_arrdiv32_fs822_and0;
  assign f_arrdiv32_fs823_xor0 = f_arrdiv32_mux2to1766_xor0 ^ b[23];
  assign f_arrdiv32_fs823_not0 = ~f_arrdiv32_mux2to1766_xor0;
  assign f_arrdiv32_fs823_and0 = f_arrdiv32_fs823_not0 & b[23];
  assign f_arrdiv32_fs823_xor1 = f_arrdiv32_fs822_or0 ^ f_arrdiv32_fs823_xor0;
  assign f_arrdiv32_fs823_not1 = ~f_arrdiv32_fs823_xor0;
  assign f_arrdiv32_fs823_and1 = f_arrdiv32_fs823_not1 & f_arrdiv32_fs822_or0;
  assign f_arrdiv32_fs823_or0 = f_arrdiv32_fs823_and1 | f_arrdiv32_fs823_and0;
  assign f_arrdiv32_fs824_xor0 = f_arrdiv32_mux2to1767_xor0 ^ b[24];
  assign f_arrdiv32_fs824_not0 = ~f_arrdiv32_mux2to1767_xor0;
  assign f_arrdiv32_fs824_and0 = f_arrdiv32_fs824_not0 & b[24];
  assign f_arrdiv32_fs824_xor1 = f_arrdiv32_fs823_or0 ^ f_arrdiv32_fs824_xor0;
  assign f_arrdiv32_fs824_not1 = ~f_arrdiv32_fs824_xor0;
  assign f_arrdiv32_fs824_and1 = f_arrdiv32_fs824_not1 & f_arrdiv32_fs823_or0;
  assign f_arrdiv32_fs824_or0 = f_arrdiv32_fs824_and1 | f_arrdiv32_fs824_and0;
  assign f_arrdiv32_fs825_xor0 = f_arrdiv32_mux2to1768_xor0 ^ b[25];
  assign f_arrdiv32_fs825_not0 = ~f_arrdiv32_mux2to1768_xor0;
  assign f_arrdiv32_fs825_and0 = f_arrdiv32_fs825_not0 & b[25];
  assign f_arrdiv32_fs825_xor1 = f_arrdiv32_fs824_or0 ^ f_arrdiv32_fs825_xor0;
  assign f_arrdiv32_fs825_not1 = ~f_arrdiv32_fs825_xor0;
  assign f_arrdiv32_fs825_and1 = f_arrdiv32_fs825_not1 & f_arrdiv32_fs824_or0;
  assign f_arrdiv32_fs825_or0 = f_arrdiv32_fs825_and1 | f_arrdiv32_fs825_and0;
  assign f_arrdiv32_fs826_xor0 = f_arrdiv32_mux2to1769_xor0 ^ b[26];
  assign f_arrdiv32_fs826_not0 = ~f_arrdiv32_mux2to1769_xor0;
  assign f_arrdiv32_fs826_and0 = f_arrdiv32_fs826_not0 & b[26];
  assign f_arrdiv32_fs826_xor1 = f_arrdiv32_fs825_or0 ^ f_arrdiv32_fs826_xor0;
  assign f_arrdiv32_fs826_not1 = ~f_arrdiv32_fs826_xor0;
  assign f_arrdiv32_fs826_and1 = f_arrdiv32_fs826_not1 & f_arrdiv32_fs825_or0;
  assign f_arrdiv32_fs826_or0 = f_arrdiv32_fs826_and1 | f_arrdiv32_fs826_and0;
  assign f_arrdiv32_fs827_xor0 = f_arrdiv32_mux2to1770_xor0 ^ b[27];
  assign f_arrdiv32_fs827_not0 = ~f_arrdiv32_mux2to1770_xor0;
  assign f_arrdiv32_fs827_and0 = f_arrdiv32_fs827_not0 & b[27];
  assign f_arrdiv32_fs827_xor1 = f_arrdiv32_fs826_or0 ^ f_arrdiv32_fs827_xor0;
  assign f_arrdiv32_fs827_not1 = ~f_arrdiv32_fs827_xor0;
  assign f_arrdiv32_fs827_and1 = f_arrdiv32_fs827_not1 & f_arrdiv32_fs826_or0;
  assign f_arrdiv32_fs827_or0 = f_arrdiv32_fs827_and1 | f_arrdiv32_fs827_and0;
  assign f_arrdiv32_fs828_xor0 = f_arrdiv32_mux2to1771_xor0 ^ b[28];
  assign f_arrdiv32_fs828_not0 = ~f_arrdiv32_mux2to1771_xor0;
  assign f_arrdiv32_fs828_and0 = f_arrdiv32_fs828_not0 & b[28];
  assign f_arrdiv32_fs828_xor1 = f_arrdiv32_fs827_or0 ^ f_arrdiv32_fs828_xor0;
  assign f_arrdiv32_fs828_not1 = ~f_arrdiv32_fs828_xor0;
  assign f_arrdiv32_fs828_and1 = f_arrdiv32_fs828_not1 & f_arrdiv32_fs827_or0;
  assign f_arrdiv32_fs828_or0 = f_arrdiv32_fs828_and1 | f_arrdiv32_fs828_and0;
  assign f_arrdiv32_fs829_xor0 = f_arrdiv32_mux2to1772_xor0 ^ b[29];
  assign f_arrdiv32_fs829_not0 = ~f_arrdiv32_mux2to1772_xor0;
  assign f_arrdiv32_fs829_and0 = f_arrdiv32_fs829_not0 & b[29];
  assign f_arrdiv32_fs829_xor1 = f_arrdiv32_fs828_or0 ^ f_arrdiv32_fs829_xor0;
  assign f_arrdiv32_fs829_not1 = ~f_arrdiv32_fs829_xor0;
  assign f_arrdiv32_fs829_and1 = f_arrdiv32_fs829_not1 & f_arrdiv32_fs828_or0;
  assign f_arrdiv32_fs829_or0 = f_arrdiv32_fs829_and1 | f_arrdiv32_fs829_and0;
  assign f_arrdiv32_fs830_xor0 = f_arrdiv32_mux2to1773_xor0 ^ b[30];
  assign f_arrdiv32_fs830_not0 = ~f_arrdiv32_mux2to1773_xor0;
  assign f_arrdiv32_fs830_and0 = f_arrdiv32_fs830_not0 & b[30];
  assign f_arrdiv32_fs830_xor1 = f_arrdiv32_fs829_or0 ^ f_arrdiv32_fs830_xor0;
  assign f_arrdiv32_fs830_not1 = ~f_arrdiv32_fs830_xor0;
  assign f_arrdiv32_fs830_and1 = f_arrdiv32_fs830_not1 & f_arrdiv32_fs829_or0;
  assign f_arrdiv32_fs830_or0 = f_arrdiv32_fs830_and1 | f_arrdiv32_fs830_and0;
  assign f_arrdiv32_fs831_xor0 = f_arrdiv32_mux2to1774_xor0 ^ b[31];
  assign f_arrdiv32_fs831_not0 = ~f_arrdiv32_mux2to1774_xor0;
  assign f_arrdiv32_fs831_and0 = f_arrdiv32_fs831_not0 & b[31];
  assign f_arrdiv32_fs831_xor1 = f_arrdiv32_fs830_or0 ^ f_arrdiv32_fs831_xor0;
  assign f_arrdiv32_fs831_not1 = ~f_arrdiv32_fs831_xor0;
  assign f_arrdiv32_fs831_and1 = f_arrdiv32_fs831_not1 & f_arrdiv32_fs830_or0;
  assign f_arrdiv32_fs831_or0 = f_arrdiv32_fs831_and1 | f_arrdiv32_fs831_and0;
  assign f_arrdiv32_mux2to1775_and0 = a[6] & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1775_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1775_and1 = f_arrdiv32_fs800_xor0 & f_arrdiv32_mux2to1775_not0;
  assign f_arrdiv32_mux2to1775_xor0 = f_arrdiv32_mux2to1775_and0 ^ f_arrdiv32_mux2to1775_and1;
  assign f_arrdiv32_mux2to1776_and0 = f_arrdiv32_mux2to1744_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1776_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1776_and1 = f_arrdiv32_fs801_xor1 & f_arrdiv32_mux2to1776_not0;
  assign f_arrdiv32_mux2to1776_xor0 = f_arrdiv32_mux2to1776_and0 ^ f_arrdiv32_mux2to1776_and1;
  assign f_arrdiv32_mux2to1777_and0 = f_arrdiv32_mux2to1745_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1777_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1777_and1 = f_arrdiv32_fs802_xor1 & f_arrdiv32_mux2to1777_not0;
  assign f_arrdiv32_mux2to1777_xor0 = f_arrdiv32_mux2to1777_and0 ^ f_arrdiv32_mux2to1777_and1;
  assign f_arrdiv32_mux2to1778_and0 = f_arrdiv32_mux2to1746_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1778_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1778_and1 = f_arrdiv32_fs803_xor1 & f_arrdiv32_mux2to1778_not0;
  assign f_arrdiv32_mux2to1778_xor0 = f_arrdiv32_mux2to1778_and0 ^ f_arrdiv32_mux2to1778_and1;
  assign f_arrdiv32_mux2to1779_and0 = f_arrdiv32_mux2to1747_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1779_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1779_and1 = f_arrdiv32_fs804_xor1 & f_arrdiv32_mux2to1779_not0;
  assign f_arrdiv32_mux2to1779_xor0 = f_arrdiv32_mux2to1779_and0 ^ f_arrdiv32_mux2to1779_and1;
  assign f_arrdiv32_mux2to1780_and0 = f_arrdiv32_mux2to1748_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1780_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1780_and1 = f_arrdiv32_fs805_xor1 & f_arrdiv32_mux2to1780_not0;
  assign f_arrdiv32_mux2to1780_xor0 = f_arrdiv32_mux2to1780_and0 ^ f_arrdiv32_mux2to1780_and1;
  assign f_arrdiv32_mux2to1781_and0 = f_arrdiv32_mux2to1749_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1781_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1781_and1 = f_arrdiv32_fs806_xor1 & f_arrdiv32_mux2to1781_not0;
  assign f_arrdiv32_mux2to1781_xor0 = f_arrdiv32_mux2to1781_and0 ^ f_arrdiv32_mux2to1781_and1;
  assign f_arrdiv32_mux2to1782_and0 = f_arrdiv32_mux2to1750_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1782_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1782_and1 = f_arrdiv32_fs807_xor1 & f_arrdiv32_mux2to1782_not0;
  assign f_arrdiv32_mux2to1782_xor0 = f_arrdiv32_mux2to1782_and0 ^ f_arrdiv32_mux2to1782_and1;
  assign f_arrdiv32_mux2to1783_and0 = f_arrdiv32_mux2to1751_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1783_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1783_and1 = f_arrdiv32_fs808_xor1 & f_arrdiv32_mux2to1783_not0;
  assign f_arrdiv32_mux2to1783_xor0 = f_arrdiv32_mux2to1783_and0 ^ f_arrdiv32_mux2to1783_and1;
  assign f_arrdiv32_mux2to1784_and0 = f_arrdiv32_mux2to1752_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1784_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1784_and1 = f_arrdiv32_fs809_xor1 & f_arrdiv32_mux2to1784_not0;
  assign f_arrdiv32_mux2to1784_xor0 = f_arrdiv32_mux2to1784_and0 ^ f_arrdiv32_mux2to1784_and1;
  assign f_arrdiv32_mux2to1785_and0 = f_arrdiv32_mux2to1753_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1785_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1785_and1 = f_arrdiv32_fs810_xor1 & f_arrdiv32_mux2to1785_not0;
  assign f_arrdiv32_mux2to1785_xor0 = f_arrdiv32_mux2to1785_and0 ^ f_arrdiv32_mux2to1785_and1;
  assign f_arrdiv32_mux2to1786_and0 = f_arrdiv32_mux2to1754_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1786_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1786_and1 = f_arrdiv32_fs811_xor1 & f_arrdiv32_mux2to1786_not0;
  assign f_arrdiv32_mux2to1786_xor0 = f_arrdiv32_mux2to1786_and0 ^ f_arrdiv32_mux2to1786_and1;
  assign f_arrdiv32_mux2to1787_and0 = f_arrdiv32_mux2to1755_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1787_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1787_and1 = f_arrdiv32_fs812_xor1 & f_arrdiv32_mux2to1787_not0;
  assign f_arrdiv32_mux2to1787_xor0 = f_arrdiv32_mux2to1787_and0 ^ f_arrdiv32_mux2to1787_and1;
  assign f_arrdiv32_mux2to1788_and0 = f_arrdiv32_mux2to1756_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1788_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1788_and1 = f_arrdiv32_fs813_xor1 & f_arrdiv32_mux2to1788_not0;
  assign f_arrdiv32_mux2to1788_xor0 = f_arrdiv32_mux2to1788_and0 ^ f_arrdiv32_mux2to1788_and1;
  assign f_arrdiv32_mux2to1789_and0 = f_arrdiv32_mux2to1757_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1789_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1789_and1 = f_arrdiv32_fs814_xor1 & f_arrdiv32_mux2to1789_not0;
  assign f_arrdiv32_mux2to1789_xor0 = f_arrdiv32_mux2to1789_and0 ^ f_arrdiv32_mux2to1789_and1;
  assign f_arrdiv32_mux2to1790_and0 = f_arrdiv32_mux2to1758_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1790_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1790_and1 = f_arrdiv32_fs815_xor1 & f_arrdiv32_mux2to1790_not0;
  assign f_arrdiv32_mux2to1790_xor0 = f_arrdiv32_mux2to1790_and0 ^ f_arrdiv32_mux2to1790_and1;
  assign f_arrdiv32_mux2to1791_and0 = f_arrdiv32_mux2to1759_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1791_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1791_and1 = f_arrdiv32_fs816_xor1 & f_arrdiv32_mux2to1791_not0;
  assign f_arrdiv32_mux2to1791_xor0 = f_arrdiv32_mux2to1791_and0 ^ f_arrdiv32_mux2to1791_and1;
  assign f_arrdiv32_mux2to1792_and0 = f_arrdiv32_mux2to1760_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1792_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1792_and1 = f_arrdiv32_fs817_xor1 & f_arrdiv32_mux2to1792_not0;
  assign f_arrdiv32_mux2to1792_xor0 = f_arrdiv32_mux2to1792_and0 ^ f_arrdiv32_mux2to1792_and1;
  assign f_arrdiv32_mux2to1793_and0 = f_arrdiv32_mux2to1761_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1793_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1793_and1 = f_arrdiv32_fs818_xor1 & f_arrdiv32_mux2to1793_not0;
  assign f_arrdiv32_mux2to1793_xor0 = f_arrdiv32_mux2to1793_and0 ^ f_arrdiv32_mux2to1793_and1;
  assign f_arrdiv32_mux2to1794_and0 = f_arrdiv32_mux2to1762_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1794_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1794_and1 = f_arrdiv32_fs819_xor1 & f_arrdiv32_mux2to1794_not0;
  assign f_arrdiv32_mux2to1794_xor0 = f_arrdiv32_mux2to1794_and0 ^ f_arrdiv32_mux2to1794_and1;
  assign f_arrdiv32_mux2to1795_and0 = f_arrdiv32_mux2to1763_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1795_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1795_and1 = f_arrdiv32_fs820_xor1 & f_arrdiv32_mux2to1795_not0;
  assign f_arrdiv32_mux2to1795_xor0 = f_arrdiv32_mux2to1795_and0 ^ f_arrdiv32_mux2to1795_and1;
  assign f_arrdiv32_mux2to1796_and0 = f_arrdiv32_mux2to1764_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1796_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1796_and1 = f_arrdiv32_fs821_xor1 & f_arrdiv32_mux2to1796_not0;
  assign f_arrdiv32_mux2to1796_xor0 = f_arrdiv32_mux2to1796_and0 ^ f_arrdiv32_mux2to1796_and1;
  assign f_arrdiv32_mux2to1797_and0 = f_arrdiv32_mux2to1765_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1797_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1797_and1 = f_arrdiv32_fs822_xor1 & f_arrdiv32_mux2to1797_not0;
  assign f_arrdiv32_mux2to1797_xor0 = f_arrdiv32_mux2to1797_and0 ^ f_arrdiv32_mux2to1797_and1;
  assign f_arrdiv32_mux2to1798_and0 = f_arrdiv32_mux2to1766_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1798_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1798_and1 = f_arrdiv32_fs823_xor1 & f_arrdiv32_mux2to1798_not0;
  assign f_arrdiv32_mux2to1798_xor0 = f_arrdiv32_mux2to1798_and0 ^ f_arrdiv32_mux2to1798_and1;
  assign f_arrdiv32_mux2to1799_and0 = f_arrdiv32_mux2to1767_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1799_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1799_and1 = f_arrdiv32_fs824_xor1 & f_arrdiv32_mux2to1799_not0;
  assign f_arrdiv32_mux2to1799_xor0 = f_arrdiv32_mux2to1799_and0 ^ f_arrdiv32_mux2to1799_and1;
  assign f_arrdiv32_mux2to1800_and0 = f_arrdiv32_mux2to1768_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1800_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1800_and1 = f_arrdiv32_fs825_xor1 & f_arrdiv32_mux2to1800_not0;
  assign f_arrdiv32_mux2to1800_xor0 = f_arrdiv32_mux2to1800_and0 ^ f_arrdiv32_mux2to1800_and1;
  assign f_arrdiv32_mux2to1801_and0 = f_arrdiv32_mux2to1769_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1801_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1801_and1 = f_arrdiv32_fs826_xor1 & f_arrdiv32_mux2to1801_not0;
  assign f_arrdiv32_mux2to1801_xor0 = f_arrdiv32_mux2to1801_and0 ^ f_arrdiv32_mux2to1801_and1;
  assign f_arrdiv32_mux2to1802_and0 = f_arrdiv32_mux2to1770_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1802_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1802_and1 = f_arrdiv32_fs827_xor1 & f_arrdiv32_mux2to1802_not0;
  assign f_arrdiv32_mux2to1802_xor0 = f_arrdiv32_mux2to1802_and0 ^ f_arrdiv32_mux2to1802_and1;
  assign f_arrdiv32_mux2to1803_and0 = f_arrdiv32_mux2to1771_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1803_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1803_and1 = f_arrdiv32_fs828_xor1 & f_arrdiv32_mux2to1803_not0;
  assign f_arrdiv32_mux2to1803_xor0 = f_arrdiv32_mux2to1803_and0 ^ f_arrdiv32_mux2to1803_and1;
  assign f_arrdiv32_mux2to1804_and0 = f_arrdiv32_mux2to1772_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1804_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1804_and1 = f_arrdiv32_fs829_xor1 & f_arrdiv32_mux2to1804_not0;
  assign f_arrdiv32_mux2to1804_xor0 = f_arrdiv32_mux2to1804_and0 ^ f_arrdiv32_mux2to1804_and1;
  assign f_arrdiv32_mux2to1805_and0 = f_arrdiv32_mux2to1773_xor0 & f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1805_not0 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_mux2to1805_and1 = f_arrdiv32_fs830_xor1 & f_arrdiv32_mux2to1805_not0;
  assign f_arrdiv32_mux2to1805_xor0 = f_arrdiv32_mux2to1805_and0 ^ f_arrdiv32_mux2to1805_and1;
  assign f_arrdiv32_not25 = ~f_arrdiv32_fs831_or0;
  assign f_arrdiv32_fs832_xor0 = a[5] ^ b[0];
  assign f_arrdiv32_fs832_not0 = ~a[5];
  assign f_arrdiv32_fs832_and0 = f_arrdiv32_fs832_not0 & b[0];
  assign f_arrdiv32_fs832_not1 = ~f_arrdiv32_fs832_xor0;
  assign f_arrdiv32_fs833_xor0 = f_arrdiv32_mux2to1775_xor0 ^ b[1];
  assign f_arrdiv32_fs833_not0 = ~f_arrdiv32_mux2to1775_xor0;
  assign f_arrdiv32_fs833_and0 = f_arrdiv32_fs833_not0 & b[1];
  assign f_arrdiv32_fs833_xor1 = f_arrdiv32_fs832_and0 ^ f_arrdiv32_fs833_xor0;
  assign f_arrdiv32_fs833_not1 = ~f_arrdiv32_fs833_xor0;
  assign f_arrdiv32_fs833_and1 = f_arrdiv32_fs833_not1 & f_arrdiv32_fs832_and0;
  assign f_arrdiv32_fs833_or0 = f_arrdiv32_fs833_and1 | f_arrdiv32_fs833_and0;
  assign f_arrdiv32_fs834_xor0 = f_arrdiv32_mux2to1776_xor0 ^ b[2];
  assign f_arrdiv32_fs834_not0 = ~f_arrdiv32_mux2to1776_xor0;
  assign f_arrdiv32_fs834_and0 = f_arrdiv32_fs834_not0 & b[2];
  assign f_arrdiv32_fs834_xor1 = f_arrdiv32_fs833_or0 ^ f_arrdiv32_fs834_xor0;
  assign f_arrdiv32_fs834_not1 = ~f_arrdiv32_fs834_xor0;
  assign f_arrdiv32_fs834_and1 = f_arrdiv32_fs834_not1 & f_arrdiv32_fs833_or0;
  assign f_arrdiv32_fs834_or0 = f_arrdiv32_fs834_and1 | f_arrdiv32_fs834_and0;
  assign f_arrdiv32_fs835_xor0 = f_arrdiv32_mux2to1777_xor0 ^ b[3];
  assign f_arrdiv32_fs835_not0 = ~f_arrdiv32_mux2to1777_xor0;
  assign f_arrdiv32_fs835_and0 = f_arrdiv32_fs835_not0 & b[3];
  assign f_arrdiv32_fs835_xor1 = f_arrdiv32_fs834_or0 ^ f_arrdiv32_fs835_xor0;
  assign f_arrdiv32_fs835_not1 = ~f_arrdiv32_fs835_xor0;
  assign f_arrdiv32_fs835_and1 = f_arrdiv32_fs835_not1 & f_arrdiv32_fs834_or0;
  assign f_arrdiv32_fs835_or0 = f_arrdiv32_fs835_and1 | f_arrdiv32_fs835_and0;
  assign f_arrdiv32_fs836_xor0 = f_arrdiv32_mux2to1778_xor0 ^ b[4];
  assign f_arrdiv32_fs836_not0 = ~f_arrdiv32_mux2to1778_xor0;
  assign f_arrdiv32_fs836_and0 = f_arrdiv32_fs836_not0 & b[4];
  assign f_arrdiv32_fs836_xor1 = f_arrdiv32_fs835_or0 ^ f_arrdiv32_fs836_xor0;
  assign f_arrdiv32_fs836_not1 = ~f_arrdiv32_fs836_xor0;
  assign f_arrdiv32_fs836_and1 = f_arrdiv32_fs836_not1 & f_arrdiv32_fs835_or0;
  assign f_arrdiv32_fs836_or0 = f_arrdiv32_fs836_and1 | f_arrdiv32_fs836_and0;
  assign f_arrdiv32_fs837_xor0 = f_arrdiv32_mux2to1779_xor0 ^ b[5];
  assign f_arrdiv32_fs837_not0 = ~f_arrdiv32_mux2to1779_xor0;
  assign f_arrdiv32_fs837_and0 = f_arrdiv32_fs837_not0 & b[5];
  assign f_arrdiv32_fs837_xor1 = f_arrdiv32_fs836_or0 ^ f_arrdiv32_fs837_xor0;
  assign f_arrdiv32_fs837_not1 = ~f_arrdiv32_fs837_xor0;
  assign f_arrdiv32_fs837_and1 = f_arrdiv32_fs837_not1 & f_arrdiv32_fs836_or0;
  assign f_arrdiv32_fs837_or0 = f_arrdiv32_fs837_and1 | f_arrdiv32_fs837_and0;
  assign f_arrdiv32_fs838_xor0 = f_arrdiv32_mux2to1780_xor0 ^ b[6];
  assign f_arrdiv32_fs838_not0 = ~f_arrdiv32_mux2to1780_xor0;
  assign f_arrdiv32_fs838_and0 = f_arrdiv32_fs838_not0 & b[6];
  assign f_arrdiv32_fs838_xor1 = f_arrdiv32_fs837_or0 ^ f_arrdiv32_fs838_xor0;
  assign f_arrdiv32_fs838_not1 = ~f_arrdiv32_fs838_xor0;
  assign f_arrdiv32_fs838_and1 = f_arrdiv32_fs838_not1 & f_arrdiv32_fs837_or0;
  assign f_arrdiv32_fs838_or0 = f_arrdiv32_fs838_and1 | f_arrdiv32_fs838_and0;
  assign f_arrdiv32_fs839_xor0 = f_arrdiv32_mux2to1781_xor0 ^ b[7];
  assign f_arrdiv32_fs839_not0 = ~f_arrdiv32_mux2to1781_xor0;
  assign f_arrdiv32_fs839_and0 = f_arrdiv32_fs839_not0 & b[7];
  assign f_arrdiv32_fs839_xor1 = f_arrdiv32_fs838_or0 ^ f_arrdiv32_fs839_xor0;
  assign f_arrdiv32_fs839_not1 = ~f_arrdiv32_fs839_xor0;
  assign f_arrdiv32_fs839_and1 = f_arrdiv32_fs839_not1 & f_arrdiv32_fs838_or0;
  assign f_arrdiv32_fs839_or0 = f_arrdiv32_fs839_and1 | f_arrdiv32_fs839_and0;
  assign f_arrdiv32_fs840_xor0 = f_arrdiv32_mux2to1782_xor0 ^ b[8];
  assign f_arrdiv32_fs840_not0 = ~f_arrdiv32_mux2to1782_xor0;
  assign f_arrdiv32_fs840_and0 = f_arrdiv32_fs840_not0 & b[8];
  assign f_arrdiv32_fs840_xor1 = f_arrdiv32_fs839_or0 ^ f_arrdiv32_fs840_xor0;
  assign f_arrdiv32_fs840_not1 = ~f_arrdiv32_fs840_xor0;
  assign f_arrdiv32_fs840_and1 = f_arrdiv32_fs840_not1 & f_arrdiv32_fs839_or0;
  assign f_arrdiv32_fs840_or0 = f_arrdiv32_fs840_and1 | f_arrdiv32_fs840_and0;
  assign f_arrdiv32_fs841_xor0 = f_arrdiv32_mux2to1783_xor0 ^ b[9];
  assign f_arrdiv32_fs841_not0 = ~f_arrdiv32_mux2to1783_xor0;
  assign f_arrdiv32_fs841_and0 = f_arrdiv32_fs841_not0 & b[9];
  assign f_arrdiv32_fs841_xor1 = f_arrdiv32_fs840_or0 ^ f_arrdiv32_fs841_xor0;
  assign f_arrdiv32_fs841_not1 = ~f_arrdiv32_fs841_xor0;
  assign f_arrdiv32_fs841_and1 = f_arrdiv32_fs841_not1 & f_arrdiv32_fs840_or0;
  assign f_arrdiv32_fs841_or0 = f_arrdiv32_fs841_and1 | f_arrdiv32_fs841_and0;
  assign f_arrdiv32_fs842_xor0 = f_arrdiv32_mux2to1784_xor0 ^ b[10];
  assign f_arrdiv32_fs842_not0 = ~f_arrdiv32_mux2to1784_xor0;
  assign f_arrdiv32_fs842_and0 = f_arrdiv32_fs842_not0 & b[10];
  assign f_arrdiv32_fs842_xor1 = f_arrdiv32_fs841_or0 ^ f_arrdiv32_fs842_xor0;
  assign f_arrdiv32_fs842_not1 = ~f_arrdiv32_fs842_xor0;
  assign f_arrdiv32_fs842_and1 = f_arrdiv32_fs842_not1 & f_arrdiv32_fs841_or0;
  assign f_arrdiv32_fs842_or0 = f_arrdiv32_fs842_and1 | f_arrdiv32_fs842_and0;
  assign f_arrdiv32_fs843_xor0 = f_arrdiv32_mux2to1785_xor0 ^ b[11];
  assign f_arrdiv32_fs843_not0 = ~f_arrdiv32_mux2to1785_xor0;
  assign f_arrdiv32_fs843_and0 = f_arrdiv32_fs843_not0 & b[11];
  assign f_arrdiv32_fs843_xor1 = f_arrdiv32_fs842_or0 ^ f_arrdiv32_fs843_xor0;
  assign f_arrdiv32_fs843_not1 = ~f_arrdiv32_fs843_xor0;
  assign f_arrdiv32_fs843_and1 = f_arrdiv32_fs843_not1 & f_arrdiv32_fs842_or0;
  assign f_arrdiv32_fs843_or0 = f_arrdiv32_fs843_and1 | f_arrdiv32_fs843_and0;
  assign f_arrdiv32_fs844_xor0 = f_arrdiv32_mux2to1786_xor0 ^ b[12];
  assign f_arrdiv32_fs844_not0 = ~f_arrdiv32_mux2to1786_xor0;
  assign f_arrdiv32_fs844_and0 = f_arrdiv32_fs844_not0 & b[12];
  assign f_arrdiv32_fs844_xor1 = f_arrdiv32_fs843_or0 ^ f_arrdiv32_fs844_xor0;
  assign f_arrdiv32_fs844_not1 = ~f_arrdiv32_fs844_xor0;
  assign f_arrdiv32_fs844_and1 = f_arrdiv32_fs844_not1 & f_arrdiv32_fs843_or0;
  assign f_arrdiv32_fs844_or0 = f_arrdiv32_fs844_and1 | f_arrdiv32_fs844_and0;
  assign f_arrdiv32_fs845_xor0 = f_arrdiv32_mux2to1787_xor0 ^ b[13];
  assign f_arrdiv32_fs845_not0 = ~f_arrdiv32_mux2to1787_xor0;
  assign f_arrdiv32_fs845_and0 = f_arrdiv32_fs845_not0 & b[13];
  assign f_arrdiv32_fs845_xor1 = f_arrdiv32_fs844_or0 ^ f_arrdiv32_fs845_xor0;
  assign f_arrdiv32_fs845_not1 = ~f_arrdiv32_fs845_xor0;
  assign f_arrdiv32_fs845_and1 = f_arrdiv32_fs845_not1 & f_arrdiv32_fs844_or0;
  assign f_arrdiv32_fs845_or0 = f_arrdiv32_fs845_and1 | f_arrdiv32_fs845_and0;
  assign f_arrdiv32_fs846_xor0 = f_arrdiv32_mux2to1788_xor0 ^ b[14];
  assign f_arrdiv32_fs846_not0 = ~f_arrdiv32_mux2to1788_xor0;
  assign f_arrdiv32_fs846_and0 = f_arrdiv32_fs846_not0 & b[14];
  assign f_arrdiv32_fs846_xor1 = f_arrdiv32_fs845_or0 ^ f_arrdiv32_fs846_xor0;
  assign f_arrdiv32_fs846_not1 = ~f_arrdiv32_fs846_xor0;
  assign f_arrdiv32_fs846_and1 = f_arrdiv32_fs846_not1 & f_arrdiv32_fs845_or0;
  assign f_arrdiv32_fs846_or0 = f_arrdiv32_fs846_and1 | f_arrdiv32_fs846_and0;
  assign f_arrdiv32_fs847_xor0 = f_arrdiv32_mux2to1789_xor0 ^ b[15];
  assign f_arrdiv32_fs847_not0 = ~f_arrdiv32_mux2to1789_xor0;
  assign f_arrdiv32_fs847_and0 = f_arrdiv32_fs847_not0 & b[15];
  assign f_arrdiv32_fs847_xor1 = f_arrdiv32_fs846_or0 ^ f_arrdiv32_fs847_xor0;
  assign f_arrdiv32_fs847_not1 = ~f_arrdiv32_fs847_xor0;
  assign f_arrdiv32_fs847_and1 = f_arrdiv32_fs847_not1 & f_arrdiv32_fs846_or0;
  assign f_arrdiv32_fs847_or0 = f_arrdiv32_fs847_and1 | f_arrdiv32_fs847_and0;
  assign f_arrdiv32_fs848_xor0 = f_arrdiv32_mux2to1790_xor0 ^ b[16];
  assign f_arrdiv32_fs848_not0 = ~f_arrdiv32_mux2to1790_xor0;
  assign f_arrdiv32_fs848_and0 = f_arrdiv32_fs848_not0 & b[16];
  assign f_arrdiv32_fs848_xor1 = f_arrdiv32_fs847_or0 ^ f_arrdiv32_fs848_xor0;
  assign f_arrdiv32_fs848_not1 = ~f_arrdiv32_fs848_xor0;
  assign f_arrdiv32_fs848_and1 = f_arrdiv32_fs848_not1 & f_arrdiv32_fs847_or0;
  assign f_arrdiv32_fs848_or0 = f_arrdiv32_fs848_and1 | f_arrdiv32_fs848_and0;
  assign f_arrdiv32_fs849_xor0 = f_arrdiv32_mux2to1791_xor0 ^ b[17];
  assign f_arrdiv32_fs849_not0 = ~f_arrdiv32_mux2to1791_xor0;
  assign f_arrdiv32_fs849_and0 = f_arrdiv32_fs849_not0 & b[17];
  assign f_arrdiv32_fs849_xor1 = f_arrdiv32_fs848_or0 ^ f_arrdiv32_fs849_xor0;
  assign f_arrdiv32_fs849_not1 = ~f_arrdiv32_fs849_xor0;
  assign f_arrdiv32_fs849_and1 = f_arrdiv32_fs849_not1 & f_arrdiv32_fs848_or0;
  assign f_arrdiv32_fs849_or0 = f_arrdiv32_fs849_and1 | f_arrdiv32_fs849_and0;
  assign f_arrdiv32_fs850_xor0 = f_arrdiv32_mux2to1792_xor0 ^ b[18];
  assign f_arrdiv32_fs850_not0 = ~f_arrdiv32_mux2to1792_xor0;
  assign f_arrdiv32_fs850_and0 = f_arrdiv32_fs850_not0 & b[18];
  assign f_arrdiv32_fs850_xor1 = f_arrdiv32_fs849_or0 ^ f_arrdiv32_fs850_xor0;
  assign f_arrdiv32_fs850_not1 = ~f_arrdiv32_fs850_xor0;
  assign f_arrdiv32_fs850_and1 = f_arrdiv32_fs850_not1 & f_arrdiv32_fs849_or0;
  assign f_arrdiv32_fs850_or0 = f_arrdiv32_fs850_and1 | f_arrdiv32_fs850_and0;
  assign f_arrdiv32_fs851_xor0 = f_arrdiv32_mux2to1793_xor0 ^ b[19];
  assign f_arrdiv32_fs851_not0 = ~f_arrdiv32_mux2to1793_xor0;
  assign f_arrdiv32_fs851_and0 = f_arrdiv32_fs851_not0 & b[19];
  assign f_arrdiv32_fs851_xor1 = f_arrdiv32_fs850_or0 ^ f_arrdiv32_fs851_xor0;
  assign f_arrdiv32_fs851_not1 = ~f_arrdiv32_fs851_xor0;
  assign f_arrdiv32_fs851_and1 = f_arrdiv32_fs851_not1 & f_arrdiv32_fs850_or0;
  assign f_arrdiv32_fs851_or0 = f_arrdiv32_fs851_and1 | f_arrdiv32_fs851_and0;
  assign f_arrdiv32_fs852_xor0 = f_arrdiv32_mux2to1794_xor0 ^ b[20];
  assign f_arrdiv32_fs852_not0 = ~f_arrdiv32_mux2to1794_xor0;
  assign f_arrdiv32_fs852_and0 = f_arrdiv32_fs852_not0 & b[20];
  assign f_arrdiv32_fs852_xor1 = f_arrdiv32_fs851_or0 ^ f_arrdiv32_fs852_xor0;
  assign f_arrdiv32_fs852_not1 = ~f_arrdiv32_fs852_xor0;
  assign f_arrdiv32_fs852_and1 = f_arrdiv32_fs852_not1 & f_arrdiv32_fs851_or0;
  assign f_arrdiv32_fs852_or0 = f_arrdiv32_fs852_and1 | f_arrdiv32_fs852_and0;
  assign f_arrdiv32_fs853_xor0 = f_arrdiv32_mux2to1795_xor0 ^ b[21];
  assign f_arrdiv32_fs853_not0 = ~f_arrdiv32_mux2to1795_xor0;
  assign f_arrdiv32_fs853_and0 = f_arrdiv32_fs853_not0 & b[21];
  assign f_arrdiv32_fs853_xor1 = f_arrdiv32_fs852_or0 ^ f_arrdiv32_fs853_xor0;
  assign f_arrdiv32_fs853_not1 = ~f_arrdiv32_fs853_xor0;
  assign f_arrdiv32_fs853_and1 = f_arrdiv32_fs853_not1 & f_arrdiv32_fs852_or0;
  assign f_arrdiv32_fs853_or0 = f_arrdiv32_fs853_and1 | f_arrdiv32_fs853_and0;
  assign f_arrdiv32_fs854_xor0 = f_arrdiv32_mux2to1796_xor0 ^ b[22];
  assign f_arrdiv32_fs854_not0 = ~f_arrdiv32_mux2to1796_xor0;
  assign f_arrdiv32_fs854_and0 = f_arrdiv32_fs854_not0 & b[22];
  assign f_arrdiv32_fs854_xor1 = f_arrdiv32_fs853_or0 ^ f_arrdiv32_fs854_xor0;
  assign f_arrdiv32_fs854_not1 = ~f_arrdiv32_fs854_xor0;
  assign f_arrdiv32_fs854_and1 = f_arrdiv32_fs854_not1 & f_arrdiv32_fs853_or0;
  assign f_arrdiv32_fs854_or0 = f_arrdiv32_fs854_and1 | f_arrdiv32_fs854_and0;
  assign f_arrdiv32_fs855_xor0 = f_arrdiv32_mux2to1797_xor0 ^ b[23];
  assign f_arrdiv32_fs855_not0 = ~f_arrdiv32_mux2to1797_xor0;
  assign f_arrdiv32_fs855_and0 = f_arrdiv32_fs855_not0 & b[23];
  assign f_arrdiv32_fs855_xor1 = f_arrdiv32_fs854_or0 ^ f_arrdiv32_fs855_xor0;
  assign f_arrdiv32_fs855_not1 = ~f_arrdiv32_fs855_xor0;
  assign f_arrdiv32_fs855_and1 = f_arrdiv32_fs855_not1 & f_arrdiv32_fs854_or0;
  assign f_arrdiv32_fs855_or0 = f_arrdiv32_fs855_and1 | f_arrdiv32_fs855_and0;
  assign f_arrdiv32_fs856_xor0 = f_arrdiv32_mux2to1798_xor0 ^ b[24];
  assign f_arrdiv32_fs856_not0 = ~f_arrdiv32_mux2to1798_xor0;
  assign f_arrdiv32_fs856_and0 = f_arrdiv32_fs856_not0 & b[24];
  assign f_arrdiv32_fs856_xor1 = f_arrdiv32_fs855_or0 ^ f_arrdiv32_fs856_xor0;
  assign f_arrdiv32_fs856_not1 = ~f_arrdiv32_fs856_xor0;
  assign f_arrdiv32_fs856_and1 = f_arrdiv32_fs856_not1 & f_arrdiv32_fs855_or0;
  assign f_arrdiv32_fs856_or0 = f_arrdiv32_fs856_and1 | f_arrdiv32_fs856_and0;
  assign f_arrdiv32_fs857_xor0 = f_arrdiv32_mux2to1799_xor0 ^ b[25];
  assign f_arrdiv32_fs857_not0 = ~f_arrdiv32_mux2to1799_xor0;
  assign f_arrdiv32_fs857_and0 = f_arrdiv32_fs857_not0 & b[25];
  assign f_arrdiv32_fs857_xor1 = f_arrdiv32_fs856_or0 ^ f_arrdiv32_fs857_xor0;
  assign f_arrdiv32_fs857_not1 = ~f_arrdiv32_fs857_xor0;
  assign f_arrdiv32_fs857_and1 = f_arrdiv32_fs857_not1 & f_arrdiv32_fs856_or0;
  assign f_arrdiv32_fs857_or0 = f_arrdiv32_fs857_and1 | f_arrdiv32_fs857_and0;
  assign f_arrdiv32_fs858_xor0 = f_arrdiv32_mux2to1800_xor0 ^ b[26];
  assign f_arrdiv32_fs858_not0 = ~f_arrdiv32_mux2to1800_xor0;
  assign f_arrdiv32_fs858_and0 = f_arrdiv32_fs858_not0 & b[26];
  assign f_arrdiv32_fs858_xor1 = f_arrdiv32_fs857_or0 ^ f_arrdiv32_fs858_xor0;
  assign f_arrdiv32_fs858_not1 = ~f_arrdiv32_fs858_xor0;
  assign f_arrdiv32_fs858_and1 = f_arrdiv32_fs858_not1 & f_arrdiv32_fs857_or0;
  assign f_arrdiv32_fs858_or0 = f_arrdiv32_fs858_and1 | f_arrdiv32_fs858_and0;
  assign f_arrdiv32_fs859_xor0 = f_arrdiv32_mux2to1801_xor0 ^ b[27];
  assign f_arrdiv32_fs859_not0 = ~f_arrdiv32_mux2to1801_xor0;
  assign f_arrdiv32_fs859_and0 = f_arrdiv32_fs859_not0 & b[27];
  assign f_arrdiv32_fs859_xor1 = f_arrdiv32_fs858_or0 ^ f_arrdiv32_fs859_xor0;
  assign f_arrdiv32_fs859_not1 = ~f_arrdiv32_fs859_xor0;
  assign f_arrdiv32_fs859_and1 = f_arrdiv32_fs859_not1 & f_arrdiv32_fs858_or0;
  assign f_arrdiv32_fs859_or0 = f_arrdiv32_fs859_and1 | f_arrdiv32_fs859_and0;
  assign f_arrdiv32_fs860_xor0 = f_arrdiv32_mux2to1802_xor0 ^ b[28];
  assign f_arrdiv32_fs860_not0 = ~f_arrdiv32_mux2to1802_xor0;
  assign f_arrdiv32_fs860_and0 = f_arrdiv32_fs860_not0 & b[28];
  assign f_arrdiv32_fs860_xor1 = f_arrdiv32_fs859_or0 ^ f_arrdiv32_fs860_xor0;
  assign f_arrdiv32_fs860_not1 = ~f_arrdiv32_fs860_xor0;
  assign f_arrdiv32_fs860_and1 = f_arrdiv32_fs860_not1 & f_arrdiv32_fs859_or0;
  assign f_arrdiv32_fs860_or0 = f_arrdiv32_fs860_and1 | f_arrdiv32_fs860_and0;
  assign f_arrdiv32_fs861_xor0 = f_arrdiv32_mux2to1803_xor0 ^ b[29];
  assign f_arrdiv32_fs861_not0 = ~f_arrdiv32_mux2to1803_xor0;
  assign f_arrdiv32_fs861_and0 = f_arrdiv32_fs861_not0 & b[29];
  assign f_arrdiv32_fs861_xor1 = f_arrdiv32_fs860_or0 ^ f_arrdiv32_fs861_xor0;
  assign f_arrdiv32_fs861_not1 = ~f_arrdiv32_fs861_xor0;
  assign f_arrdiv32_fs861_and1 = f_arrdiv32_fs861_not1 & f_arrdiv32_fs860_or0;
  assign f_arrdiv32_fs861_or0 = f_arrdiv32_fs861_and1 | f_arrdiv32_fs861_and0;
  assign f_arrdiv32_fs862_xor0 = f_arrdiv32_mux2to1804_xor0 ^ b[30];
  assign f_arrdiv32_fs862_not0 = ~f_arrdiv32_mux2to1804_xor0;
  assign f_arrdiv32_fs862_and0 = f_arrdiv32_fs862_not0 & b[30];
  assign f_arrdiv32_fs862_xor1 = f_arrdiv32_fs861_or0 ^ f_arrdiv32_fs862_xor0;
  assign f_arrdiv32_fs862_not1 = ~f_arrdiv32_fs862_xor0;
  assign f_arrdiv32_fs862_and1 = f_arrdiv32_fs862_not1 & f_arrdiv32_fs861_or0;
  assign f_arrdiv32_fs862_or0 = f_arrdiv32_fs862_and1 | f_arrdiv32_fs862_and0;
  assign f_arrdiv32_fs863_xor0 = f_arrdiv32_mux2to1805_xor0 ^ b[31];
  assign f_arrdiv32_fs863_not0 = ~f_arrdiv32_mux2to1805_xor0;
  assign f_arrdiv32_fs863_and0 = f_arrdiv32_fs863_not0 & b[31];
  assign f_arrdiv32_fs863_xor1 = f_arrdiv32_fs862_or0 ^ f_arrdiv32_fs863_xor0;
  assign f_arrdiv32_fs863_not1 = ~f_arrdiv32_fs863_xor0;
  assign f_arrdiv32_fs863_and1 = f_arrdiv32_fs863_not1 & f_arrdiv32_fs862_or0;
  assign f_arrdiv32_fs863_or0 = f_arrdiv32_fs863_and1 | f_arrdiv32_fs863_and0;
  assign f_arrdiv32_mux2to1806_and0 = a[5] & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1806_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1806_and1 = f_arrdiv32_fs832_xor0 & f_arrdiv32_mux2to1806_not0;
  assign f_arrdiv32_mux2to1806_xor0 = f_arrdiv32_mux2to1806_and0 ^ f_arrdiv32_mux2to1806_and1;
  assign f_arrdiv32_mux2to1807_and0 = f_arrdiv32_mux2to1775_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1807_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1807_and1 = f_arrdiv32_fs833_xor1 & f_arrdiv32_mux2to1807_not0;
  assign f_arrdiv32_mux2to1807_xor0 = f_arrdiv32_mux2to1807_and0 ^ f_arrdiv32_mux2to1807_and1;
  assign f_arrdiv32_mux2to1808_and0 = f_arrdiv32_mux2to1776_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1808_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1808_and1 = f_arrdiv32_fs834_xor1 & f_arrdiv32_mux2to1808_not0;
  assign f_arrdiv32_mux2to1808_xor0 = f_arrdiv32_mux2to1808_and0 ^ f_arrdiv32_mux2to1808_and1;
  assign f_arrdiv32_mux2to1809_and0 = f_arrdiv32_mux2to1777_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1809_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1809_and1 = f_arrdiv32_fs835_xor1 & f_arrdiv32_mux2to1809_not0;
  assign f_arrdiv32_mux2to1809_xor0 = f_arrdiv32_mux2to1809_and0 ^ f_arrdiv32_mux2to1809_and1;
  assign f_arrdiv32_mux2to1810_and0 = f_arrdiv32_mux2to1778_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1810_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1810_and1 = f_arrdiv32_fs836_xor1 & f_arrdiv32_mux2to1810_not0;
  assign f_arrdiv32_mux2to1810_xor0 = f_arrdiv32_mux2to1810_and0 ^ f_arrdiv32_mux2to1810_and1;
  assign f_arrdiv32_mux2to1811_and0 = f_arrdiv32_mux2to1779_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1811_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1811_and1 = f_arrdiv32_fs837_xor1 & f_arrdiv32_mux2to1811_not0;
  assign f_arrdiv32_mux2to1811_xor0 = f_arrdiv32_mux2to1811_and0 ^ f_arrdiv32_mux2to1811_and1;
  assign f_arrdiv32_mux2to1812_and0 = f_arrdiv32_mux2to1780_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1812_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1812_and1 = f_arrdiv32_fs838_xor1 & f_arrdiv32_mux2to1812_not0;
  assign f_arrdiv32_mux2to1812_xor0 = f_arrdiv32_mux2to1812_and0 ^ f_arrdiv32_mux2to1812_and1;
  assign f_arrdiv32_mux2to1813_and0 = f_arrdiv32_mux2to1781_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1813_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1813_and1 = f_arrdiv32_fs839_xor1 & f_arrdiv32_mux2to1813_not0;
  assign f_arrdiv32_mux2to1813_xor0 = f_arrdiv32_mux2to1813_and0 ^ f_arrdiv32_mux2to1813_and1;
  assign f_arrdiv32_mux2to1814_and0 = f_arrdiv32_mux2to1782_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1814_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1814_and1 = f_arrdiv32_fs840_xor1 & f_arrdiv32_mux2to1814_not0;
  assign f_arrdiv32_mux2to1814_xor0 = f_arrdiv32_mux2to1814_and0 ^ f_arrdiv32_mux2to1814_and1;
  assign f_arrdiv32_mux2to1815_and0 = f_arrdiv32_mux2to1783_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1815_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1815_and1 = f_arrdiv32_fs841_xor1 & f_arrdiv32_mux2to1815_not0;
  assign f_arrdiv32_mux2to1815_xor0 = f_arrdiv32_mux2to1815_and0 ^ f_arrdiv32_mux2to1815_and1;
  assign f_arrdiv32_mux2to1816_and0 = f_arrdiv32_mux2to1784_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1816_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1816_and1 = f_arrdiv32_fs842_xor1 & f_arrdiv32_mux2to1816_not0;
  assign f_arrdiv32_mux2to1816_xor0 = f_arrdiv32_mux2to1816_and0 ^ f_arrdiv32_mux2to1816_and1;
  assign f_arrdiv32_mux2to1817_and0 = f_arrdiv32_mux2to1785_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1817_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1817_and1 = f_arrdiv32_fs843_xor1 & f_arrdiv32_mux2to1817_not0;
  assign f_arrdiv32_mux2to1817_xor0 = f_arrdiv32_mux2to1817_and0 ^ f_arrdiv32_mux2to1817_and1;
  assign f_arrdiv32_mux2to1818_and0 = f_arrdiv32_mux2to1786_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1818_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1818_and1 = f_arrdiv32_fs844_xor1 & f_arrdiv32_mux2to1818_not0;
  assign f_arrdiv32_mux2to1818_xor0 = f_arrdiv32_mux2to1818_and0 ^ f_arrdiv32_mux2to1818_and1;
  assign f_arrdiv32_mux2to1819_and0 = f_arrdiv32_mux2to1787_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1819_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1819_and1 = f_arrdiv32_fs845_xor1 & f_arrdiv32_mux2to1819_not0;
  assign f_arrdiv32_mux2to1819_xor0 = f_arrdiv32_mux2to1819_and0 ^ f_arrdiv32_mux2to1819_and1;
  assign f_arrdiv32_mux2to1820_and0 = f_arrdiv32_mux2to1788_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1820_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1820_and1 = f_arrdiv32_fs846_xor1 & f_arrdiv32_mux2to1820_not0;
  assign f_arrdiv32_mux2to1820_xor0 = f_arrdiv32_mux2to1820_and0 ^ f_arrdiv32_mux2to1820_and1;
  assign f_arrdiv32_mux2to1821_and0 = f_arrdiv32_mux2to1789_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1821_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1821_and1 = f_arrdiv32_fs847_xor1 & f_arrdiv32_mux2to1821_not0;
  assign f_arrdiv32_mux2to1821_xor0 = f_arrdiv32_mux2to1821_and0 ^ f_arrdiv32_mux2to1821_and1;
  assign f_arrdiv32_mux2to1822_and0 = f_arrdiv32_mux2to1790_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1822_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1822_and1 = f_arrdiv32_fs848_xor1 & f_arrdiv32_mux2to1822_not0;
  assign f_arrdiv32_mux2to1822_xor0 = f_arrdiv32_mux2to1822_and0 ^ f_arrdiv32_mux2to1822_and1;
  assign f_arrdiv32_mux2to1823_and0 = f_arrdiv32_mux2to1791_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1823_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1823_and1 = f_arrdiv32_fs849_xor1 & f_arrdiv32_mux2to1823_not0;
  assign f_arrdiv32_mux2to1823_xor0 = f_arrdiv32_mux2to1823_and0 ^ f_arrdiv32_mux2to1823_and1;
  assign f_arrdiv32_mux2to1824_and0 = f_arrdiv32_mux2to1792_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1824_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1824_and1 = f_arrdiv32_fs850_xor1 & f_arrdiv32_mux2to1824_not0;
  assign f_arrdiv32_mux2to1824_xor0 = f_arrdiv32_mux2to1824_and0 ^ f_arrdiv32_mux2to1824_and1;
  assign f_arrdiv32_mux2to1825_and0 = f_arrdiv32_mux2to1793_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1825_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1825_and1 = f_arrdiv32_fs851_xor1 & f_arrdiv32_mux2to1825_not0;
  assign f_arrdiv32_mux2to1825_xor0 = f_arrdiv32_mux2to1825_and0 ^ f_arrdiv32_mux2to1825_and1;
  assign f_arrdiv32_mux2to1826_and0 = f_arrdiv32_mux2to1794_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1826_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1826_and1 = f_arrdiv32_fs852_xor1 & f_arrdiv32_mux2to1826_not0;
  assign f_arrdiv32_mux2to1826_xor0 = f_arrdiv32_mux2to1826_and0 ^ f_arrdiv32_mux2to1826_and1;
  assign f_arrdiv32_mux2to1827_and0 = f_arrdiv32_mux2to1795_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1827_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1827_and1 = f_arrdiv32_fs853_xor1 & f_arrdiv32_mux2to1827_not0;
  assign f_arrdiv32_mux2to1827_xor0 = f_arrdiv32_mux2to1827_and0 ^ f_arrdiv32_mux2to1827_and1;
  assign f_arrdiv32_mux2to1828_and0 = f_arrdiv32_mux2to1796_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1828_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1828_and1 = f_arrdiv32_fs854_xor1 & f_arrdiv32_mux2to1828_not0;
  assign f_arrdiv32_mux2to1828_xor0 = f_arrdiv32_mux2to1828_and0 ^ f_arrdiv32_mux2to1828_and1;
  assign f_arrdiv32_mux2to1829_and0 = f_arrdiv32_mux2to1797_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1829_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1829_and1 = f_arrdiv32_fs855_xor1 & f_arrdiv32_mux2to1829_not0;
  assign f_arrdiv32_mux2to1829_xor0 = f_arrdiv32_mux2to1829_and0 ^ f_arrdiv32_mux2to1829_and1;
  assign f_arrdiv32_mux2to1830_and0 = f_arrdiv32_mux2to1798_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1830_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1830_and1 = f_arrdiv32_fs856_xor1 & f_arrdiv32_mux2to1830_not0;
  assign f_arrdiv32_mux2to1830_xor0 = f_arrdiv32_mux2to1830_and0 ^ f_arrdiv32_mux2to1830_and1;
  assign f_arrdiv32_mux2to1831_and0 = f_arrdiv32_mux2to1799_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1831_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1831_and1 = f_arrdiv32_fs857_xor1 & f_arrdiv32_mux2to1831_not0;
  assign f_arrdiv32_mux2to1831_xor0 = f_arrdiv32_mux2to1831_and0 ^ f_arrdiv32_mux2to1831_and1;
  assign f_arrdiv32_mux2to1832_and0 = f_arrdiv32_mux2to1800_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1832_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1832_and1 = f_arrdiv32_fs858_xor1 & f_arrdiv32_mux2to1832_not0;
  assign f_arrdiv32_mux2to1832_xor0 = f_arrdiv32_mux2to1832_and0 ^ f_arrdiv32_mux2to1832_and1;
  assign f_arrdiv32_mux2to1833_and0 = f_arrdiv32_mux2to1801_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1833_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1833_and1 = f_arrdiv32_fs859_xor1 & f_arrdiv32_mux2to1833_not0;
  assign f_arrdiv32_mux2to1833_xor0 = f_arrdiv32_mux2to1833_and0 ^ f_arrdiv32_mux2to1833_and1;
  assign f_arrdiv32_mux2to1834_and0 = f_arrdiv32_mux2to1802_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1834_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1834_and1 = f_arrdiv32_fs860_xor1 & f_arrdiv32_mux2to1834_not0;
  assign f_arrdiv32_mux2to1834_xor0 = f_arrdiv32_mux2to1834_and0 ^ f_arrdiv32_mux2to1834_and1;
  assign f_arrdiv32_mux2to1835_and0 = f_arrdiv32_mux2to1803_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1835_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1835_and1 = f_arrdiv32_fs861_xor1 & f_arrdiv32_mux2to1835_not0;
  assign f_arrdiv32_mux2to1835_xor0 = f_arrdiv32_mux2to1835_and0 ^ f_arrdiv32_mux2to1835_and1;
  assign f_arrdiv32_mux2to1836_and0 = f_arrdiv32_mux2to1804_xor0 & f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1836_not0 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_mux2to1836_and1 = f_arrdiv32_fs862_xor1 & f_arrdiv32_mux2to1836_not0;
  assign f_arrdiv32_mux2to1836_xor0 = f_arrdiv32_mux2to1836_and0 ^ f_arrdiv32_mux2to1836_and1;
  assign f_arrdiv32_not26 = ~f_arrdiv32_fs863_or0;
  assign f_arrdiv32_fs864_xor0 = a[4] ^ b[0];
  assign f_arrdiv32_fs864_not0 = ~a[4];
  assign f_arrdiv32_fs864_and0 = f_arrdiv32_fs864_not0 & b[0];
  assign f_arrdiv32_fs864_not1 = ~f_arrdiv32_fs864_xor0;
  assign f_arrdiv32_fs865_xor0 = f_arrdiv32_mux2to1806_xor0 ^ b[1];
  assign f_arrdiv32_fs865_not0 = ~f_arrdiv32_mux2to1806_xor0;
  assign f_arrdiv32_fs865_and0 = f_arrdiv32_fs865_not0 & b[1];
  assign f_arrdiv32_fs865_xor1 = f_arrdiv32_fs864_and0 ^ f_arrdiv32_fs865_xor0;
  assign f_arrdiv32_fs865_not1 = ~f_arrdiv32_fs865_xor0;
  assign f_arrdiv32_fs865_and1 = f_arrdiv32_fs865_not1 & f_arrdiv32_fs864_and0;
  assign f_arrdiv32_fs865_or0 = f_arrdiv32_fs865_and1 | f_arrdiv32_fs865_and0;
  assign f_arrdiv32_fs866_xor0 = f_arrdiv32_mux2to1807_xor0 ^ b[2];
  assign f_arrdiv32_fs866_not0 = ~f_arrdiv32_mux2to1807_xor0;
  assign f_arrdiv32_fs866_and0 = f_arrdiv32_fs866_not0 & b[2];
  assign f_arrdiv32_fs866_xor1 = f_arrdiv32_fs865_or0 ^ f_arrdiv32_fs866_xor0;
  assign f_arrdiv32_fs866_not1 = ~f_arrdiv32_fs866_xor0;
  assign f_arrdiv32_fs866_and1 = f_arrdiv32_fs866_not1 & f_arrdiv32_fs865_or0;
  assign f_arrdiv32_fs866_or0 = f_arrdiv32_fs866_and1 | f_arrdiv32_fs866_and0;
  assign f_arrdiv32_fs867_xor0 = f_arrdiv32_mux2to1808_xor0 ^ b[3];
  assign f_arrdiv32_fs867_not0 = ~f_arrdiv32_mux2to1808_xor0;
  assign f_arrdiv32_fs867_and0 = f_arrdiv32_fs867_not0 & b[3];
  assign f_arrdiv32_fs867_xor1 = f_arrdiv32_fs866_or0 ^ f_arrdiv32_fs867_xor0;
  assign f_arrdiv32_fs867_not1 = ~f_arrdiv32_fs867_xor0;
  assign f_arrdiv32_fs867_and1 = f_arrdiv32_fs867_not1 & f_arrdiv32_fs866_or0;
  assign f_arrdiv32_fs867_or0 = f_arrdiv32_fs867_and1 | f_arrdiv32_fs867_and0;
  assign f_arrdiv32_fs868_xor0 = f_arrdiv32_mux2to1809_xor0 ^ b[4];
  assign f_arrdiv32_fs868_not0 = ~f_arrdiv32_mux2to1809_xor0;
  assign f_arrdiv32_fs868_and0 = f_arrdiv32_fs868_not0 & b[4];
  assign f_arrdiv32_fs868_xor1 = f_arrdiv32_fs867_or0 ^ f_arrdiv32_fs868_xor0;
  assign f_arrdiv32_fs868_not1 = ~f_arrdiv32_fs868_xor0;
  assign f_arrdiv32_fs868_and1 = f_arrdiv32_fs868_not1 & f_arrdiv32_fs867_or0;
  assign f_arrdiv32_fs868_or0 = f_arrdiv32_fs868_and1 | f_arrdiv32_fs868_and0;
  assign f_arrdiv32_fs869_xor0 = f_arrdiv32_mux2to1810_xor0 ^ b[5];
  assign f_arrdiv32_fs869_not0 = ~f_arrdiv32_mux2to1810_xor0;
  assign f_arrdiv32_fs869_and0 = f_arrdiv32_fs869_not0 & b[5];
  assign f_arrdiv32_fs869_xor1 = f_arrdiv32_fs868_or0 ^ f_arrdiv32_fs869_xor0;
  assign f_arrdiv32_fs869_not1 = ~f_arrdiv32_fs869_xor0;
  assign f_arrdiv32_fs869_and1 = f_arrdiv32_fs869_not1 & f_arrdiv32_fs868_or0;
  assign f_arrdiv32_fs869_or0 = f_arrdiv32_fs869_and1 | f_arrdiv32_fs869_and0;
  assign f_arrdiv32_fs870_xor0 = f_arrdiv32_mux2to1811_xor0 ^ b[6];
  assign f_arrdiv32_fs870_not0 = ~f_arrdiv32_mux2to1811_xor0;
  assign f_arrdiv32_fs870_and0 = f_arrdiv32_fs870_not0 & b[6];
  assign f_arrdiv32_fs870_xor1 = f_arrdiv32_fs869_or0 ^ f_arrdiv32_fs870_xor0;
  assign f_arrdiv32_fs870_not1 = ~f_arrdiv32_fs870_xor0;
  assign f_arrdiv32_fs870_and1 = f_arrdiv32_fs870_not1 & f_arrdiv32_fs869_or0;
  assign f_arrdiv32_fs870_or0 = f_arrdiv32_fs870_and1 | f_arrdiv32_fs870_and0;
  assign f_arrdiv32_fs871_xor0 = f_arrdiv32_mux2to1812_xor0 ^ b[7];
  assign f_arrdiv32_fs871_not0 = ~f_arrdiv32_mux2to1812_xor0;
  assign f_arrdiv32_fs871_and0 = f_arrdiv32_fs871_not0 & b[7];
  assign f_arrdiv32_fs871_xor1 = f_arrdiv32_fs870_or0 ^ f_arrdiv32_fs871_xor0;
  assign f_arrdiv32_fs871_not1 = ~f_arrdiv32_fs871_xor0;
  assign f_arrdiv32_fs871_and1 = f_arrdiv32_fs871_not1 & f_arrdiv32_fs870_or0;
  assign f_arrdiv32_fs871_or0 = f_arrdiv32_fs871_and1 | f_arrdiv32_fs871_and0;
  assign f_arrdiv32_fs872_xor0 = f_arrdiv32_mux2to1813_xor0 ^ b[8];
  assign f_arrdiv32_fs872_not0 = ~f_arrdiv32_mux2to1813_xor0;
  assign f_arrdiv32_fs872_and0 = f_arrdiv32_fs872_not0 & b[8];
  assign f_arrdiv32_fs872_xor1 = f_arrdiv32_fs871_or0 ^ f_arrdiv32_fs872_xor0;
  assign f_arrdiv32_fs872_not1 = ~f_arrdiv32_fs872_xor0;
  assign f_arrdiv32_fs872_and1 = f_arrdiv32_fs872_not1 & f_arrdiv32_fs871_or0;
  assign f_arrdiv32_fs872_or0 = f_arrdiv32_fs872_and1 | f_arrdiv32_fs872_and0;
  assign f_arrdiv32_fs873_xor0 = f_arrdiv32_mux2to1814_xor0 ^ b[9];
  assign f_arrdiv32_fs873_not0 = ~f_arrdiv32_mux2to1814_xor0;
  assign f_arrdiv32_fs873_and0 = f_arrdiv32_fs873_not0 & b[9];
  assign f_arrdiv32_fs873_xor1 = f_arrdiv32_fs872_or0 ^ f_arrdiv32_fs873_xor0;
  assign f_arrdiv32_fs873_not1 = ~f_arrdiv32_fs873_xor0;
  assign f_arrdiv32_fs873_and1 = f_arrdiv32_fs873_not1 & f_arrdiv32_fs872_or0;
  assign f_arrdiv32_fs873_or0 = f_arrdiv32_fs873_and1 | f_arrdiv32_fs873_and0;
  assign f_arrdiv32_fs874_xor0 = f_arrdiv32_mux2to1815_xor0 ^ b[10];
  assign f_arrdiv32_fs874_not0 = ~f_arrdiv32_mux2to1815_xor0;
  assign f_arrdiv32_fs874_and0 = f_arrdiv32_fs874_not0 & b[10];
  assign f_arrdiv32_fs874_xor1 = f_arrdiv32_fs873_or0 ^ f_arrdiv32_fs874_xor0;
  assign f_arrdiv32_fs874_not1 = ~f_arrdiv32_fs874_xor0;
  assign f_arrdiv32_fs874_and1 = f_arrdiv32_fs874_not1 & f_arrdiv32_fs873_or0;
  assign f_arrdiv32_fs874_or0 = f_arrdiv32_fs874_and1 | f_arrdiv32_fs874_and0;
  assign f_arrdiv32_fs875_xor0 = f_arrdiv32_mux2to1816_xor0 ^ b[11];
  assign f_arrdiv32_fs875_not0 = ~f_arrdiv32_mux2to1816_xor0;
  assign f_arrdiv32_fs875_and0 = f_arrdiv32_fs875_not0 & b[11];
  assign f_arrdiv32_fs875_xor1 = f_arrdiv32_fs874_or0 ^ f_arrdiv32_fs875_xor0;
  assign f_arrdiv32_fs875_not1 = ~f_arrdiv32_fs875_xor0;
  assign f_arrdiv32_fs875_and1 = f_arrdiv32_fs875_not1 & f_arrdiv32_fs874_or0;
  assign f_arrdiv32_fs875_or0 = f_arrdiv32_fs875_and1 | f_arrdiv32_fs875_and0;
  assign f_arrdiv32_fs876_xor0 = f_arrdiv32_mux2to1817_xor0 ^ b[12];
  assign f_arrdiv32_fs876_not0 = ~f_arrdiv32_mux2to1817_xor0;
  assign f_arrdiv32_fs876_and0 = f_arrdiv32_fs876_not0 & b[12];
  assign f_arrdiv32_fs876_xor1 = f_arrdiv32_fs875_or0 ^ f_arrdiv32_fs876_xor0;
  assign f_arrdiv32_fs876_not1 = ~f_arrdiv32_fs876_xor0;
  assign f_arrdiv32_fs876_and1 = f_arrdiv32_fs876_not1 & f_arrdiv32_fs875_or0;
  assign f_arrdiv32_fs876_or0 = f_arrdiv32_fs876_and1 | f_arrdiv32_fs876_and0;
  assign f_arrdiv32_fs877_xor0 = f_arrdiv32_mux2to1818_xor0 ^ b[13];
  assign f_arrdiv32_fs877_not0 = ~f_arrdiv32_mux2to1818_xor0;
  assign f_arrdiv32_fs877_and0 = f_arrdiv32_fs877_not0 & b[13];
  assign f_arrdiv32_fs877_xor1 = f_arrdiv32_fs876_or0 ^ f_arrdiv32_fs877_xor0;
  assign f_arrdiv32_fs877_not1 = ~f_arrdiv32_fs877_xor0;
  assign f_arrdiv32_fs877_and1 = f_arrdiv32_fs877_not1 & f_arrdiv32_fs876_or0;
  assign f_arrdiv32_fs877_or0 = f_arrdiv32_fs877_and1 | f_arrdiv32_fs877_and0;
  assign f_arrdiv32_fs878_xor0 = f_arrdiv32_mux2to1819_xor0 ^ b[14];
  assign f_arrdiv32_fs878_not0 = ~f_arrdiv32_mux2to1819_xor0;
  assign f_arrdiv32_fs878_and0 = f_arrdiv32_fs878_not0 & b[14];
  assign f_arrdiv32_fs878_xor1 = f_arrdiv32_fs877_or0 ^ f_arrdiv32_fs878_xor0;
  assign f_arrdiv32_fs878_not1 = ~f_arrdiv32_fs878_xor0;
  assign f_arrdiv32_fs878_and1 = f_arrdiv32_fs878_not1 & f_arrdiv32_fs877_or0;
  assign f_arrdiv32_fs878_or0 = f_arrdiv32_fs878_and1 | f_arrdiv32_fs878_and0;
  assign f_arrdiv32_fs879_xor0 = f_arrdiv32_mux2to1820_xor0 ^ b[15];
  assign f_arrdiv32_fs879_not0 = ~f_arrdiv32_mux2to1820_xor0;
  assign f_arrdiv32_fs879_and0 = f_arrdiv32_fs879_not0 & b[15];
  assign f_arrdiv32_fs879_xor1 = f_arrdiv32_fs878_or0 ^ f_arrdiv32_fs879_xor0;
  assign f_arrdiv32_fs879_not1 = ~f_arrdiv32_fs879_xor0;
  assign f_arrdiv32_fs879_and1 = f_arrdiv32_fs879_not1 & f_arrdiv32_fs878_or0;
  assign f_arrdiv32_fs879_or0 = f_arrdiv32_fs879_and1 | f_arrdiv32_fs879_and0;
  assign f_arrdiv32_fs880_xor0 = f_arrdiv32_mux2to1821_xor0 ^ b[16];
  assign f_arrdiv32_fs880_not0 = ~f_arrdiv32_mux2to1821_xor0;
  assign f_arrdiv32_fs880_and0 = f_arrdiv32_fs880_not0 & b[16];
  assign f_arrdiv32_fs880_xor1 = f_arrdiv32_fs879_or0 ^ f_arrdiv32_fs880_xor0;
  assign f_arrdiv32_fs880_not1 = ~f_arrdiv32_fs880_xor0;
  assign f_arrdiv32_fs880_and1 = f_arrdiv32_fs880_not1 & f_arrdiv32_fs879_or0;
  assign f_arrdiv32_fs880_or0 = f_arrdiv32_fs880_and1 | f_arrdiv32_fs880_and0;
  assign f_arrdiv32_fs881_xor0 = f_arrdiv32_mux2to1822_xor0 ^ b[17];
  assign f_arrdiv32_fs881_not0 = ~f_arrdiv32_mux2to1822_xor0;
  assign f_arrdiv32_fs881_and0 = f_arrdiv32_fs881_not0 & b[17];
  assign f_arrdiv32_fs881_xor1 = f_arrdiv32_fs880_or0 ^ f_arrdiv32_fs881_xor0;
  assign f_arrdiv32_fs881_not1 = ~f_arrdiv32_fs881_xor0;
  assign f_arrdiv32_fs881_and1 = f_arrdiv32_fs881_not1 & f_arrdiv32_fs880_or0;
  assign f_arrdiv32_fs881_or0 = f_arrdiv32_fs881_and1 | f_arrdiv32_fs881_and0;
  assign f_arrdiv32_fs882_xor0 = f_arrdiv32_mux2to1823_xor0 ^ b[18];
  assign f_arrdiv32_fs882_not0 = ~f_arrdiv32_mux2to1823_xor0;
  assign f_arrdiv32_fs882_and0 = f_arrdiv32_fs882_not0 & b[18];
  assign f_arrdiv32_fs882_xor1 = f_arrdiv32_fs881_or0 ^ f_arrdiv32_fs882_xor0;
  assign f_arrdiv32_fs882_not1 = ~f_arrdiv32_fs882_xor0;
  assign f_arrdiv32_fs882_and1 = f_arrdiv32_fs882_not1 & f_arrdiv32_fs881_or0;
  assign f_arrdiv32_fs882_or0 = f_arrdiv32_fs882_and1 | f_arrdiv32_fs882_and0;
  assign f_arrdiv32_fs883_xor0 = f_arrdiv32_mux2to1824_xor0 ^ b[19];
  assign f_arrdiv32_fs883_not0 = ~f_arrdiv32_mux2to1824_xor0;
  assign f_arrdiv32_fs883_and0 = f_arrdiv32_fs883_not0 & b[19];
  assign f_arrdiv32_fs883_xor1 = f_arrdiv32_fs882_or0 ^ f_arrdiv32_fs883_xor0;
  assign f_arrdiv32_fs883_not1 = ~f_arrdiv32_fs883_xor0;
  assign f_arrdiv32_fs883_and1 = f_arrdiv32_fs883_not1 & f_arrdiv32_fs882_or0;
  assign f_arrdiv32_fs883_or0 = f_arrdiv32_fs883_and1 | f_arrdiv32_fs883_and0;
  assign f_arrdiv32_fs884_xor0 = f_arrdiv32_mux2to1825_xor0 ^ b[20];
  assign f_arrdiv32_fs884_not0 = ~f_arrdiv32_mux2to1825_xor0;
  assign f_arrdiv32_fs884_and0 = f_arrdiv32_fs884_not0 & b[20];
  assign f_arrdiv32_fs884_xor1 = f_arrdiv32_fs883_or0 ^ f_arrdiv32_fs884_xor0;
  assign f_arrdiv32_fs884_not1 = ~f_arrdiv32_fs884_xor0;
  assign f_arrdiv32_fs884_and1 = f_arrdiv32_fs884_not1 & f_arrdiv32_fs883_or0;
  assign f_arrdiv32_fs884_or0 = f_arrdiv32_fs884_and1 | f_arrdiv32_fs884_and0;
  assign f_arrdiv32_fs885_xor0 = f_arrdiv32_mux2to1826_xor0 ^ b[21];
  assign f_arrdiv32_fs885_not0 = ~f_arrdiv32_mux2to1826_xor0;
  assign f_arrdiv32_fs885_and0 = f_arrdiv32_fs885_not0 & b[21];
  assign f_arrdiv32_fs885_xor1 = f_arrdiv32_fs884_or0 ^ f_arrdiv32_fs885_xor0;
  assign f_arrdiv32_fs885_not1 = ~f_arrdiv32_fs885_xor0;
  assign f_arrdiv32_fs885_and1 = f_arrdiv32_fs885_not1 & f_arrdiv32_fs884_or0;
  assign f_arrdiv32_fs885_or0 = f_arrdiv32_fs885_and1 | f_arrdiv32_fs885_and0;
  assign f_arrdiv32_fs886_xor0 = f_arrdiv32_mux2to1827_xor0 ^ b[22];
  assign f_arrdiv32_fs886_not0 = ~f_arrdiv32_mux2to1827_xor0;
  assign f_arrdiv32_fs886_and0 = f_arrdiv32_fs886_not0 & b[22];
  assign f_arrdiv32_fs886_xor1 = f_arrdiv32_fs885_or0 ^ f_arrdiv32_fs886_xor0;
  assign f_arrdiv32_fs886_not1 = ~f_arrdiv32_fs886_xor0;
  assign f_arrdiv32_fs886_and1 = f_arrdiv32_fs886_not1 & f_arrdiv32_fs885_or0;
  assign f_arrdiv32_fs886_or0 = f_arrdiv32_fs886_and1 | f_arrdiv32_fs886_and0;
  assign f_arrdiv32_fs887_xor0 = f_arrdiv32_mux2to1828_xor0 ^ b[23];
  assign f_arrdiv32_fs887_not0 = ~f_arrdiv32_mux2to1828_xor0;
  assign f_arrdiv32_fs887_and0 = f_arrdiv32_fs887_not0 & b[23];
  assign f_arrdiv32_fs887_xor1 = f_arrdiv32_fs886_or0 ^ f_arrdiv32_fs887_xor0;
  assign f_arrdiv32_fs887_not1 = ~f_arrdiv32_fs887_xor0;
  assign f_arrdiv32_fs887_and1 = f_arrdiv32_fs887_not1 & f_arrdiv32_fs886_or0;
  assign f_arrdiv32_fs887_or0 = f_arrdiv32_fs887_and1 | f_arrdiv32_fs887_and0;
  assign f_arrdiv32_fs888_xor0 = f_arrdiv32_mux2to1829_xor0 ^ b[24];
  assign f_arrdiv32_fs888_not0 = ~f_arrdiv32_mux2to1829_xor0;
  assign f_arrdiv32_fs888_and0 = f_arrdiv32_fs888_not0 & b[24];
  assign f_arrdiv32_fs888_xor1 = f_arrdiv32_fs887_or0 ^ f_arrdiv32_fs888_xor0;
  assign f_arrdiv32_fs888_not1 = ~f_arrdiv32_fs888_xor0;
  assign f_arrdiv32_fs888_and1 = f_arrdiv32_fs888_not1 & f_arrdiv32_fs887_or0;
  assign f_arrdiv32_fs888_or0 = f_arrdiv32_fs888_and1 | f_arrdiv32_fs888_and0;
  assign f_arrdiv32_fs889_xor0 = f_arrdiv32_mux2to1830_xor0 ^ b[25];
  assign f_arrdiv32_fs889_not0 = ~f_arrdiv32_mux2to1830_xor0;
  assign f_arrdiv32_fs889_and0 = f_arrdiv32_fs889_not0 & b[25];
  assign f_arrdiv32_fs889_xor1 = f_arrdiv32_fs888_or0 ^ f_arrdiv32_fs889_xor0;
  assign f_arrdiv32_fs889_not1 = ~f_arrdiv32_fs889_xor0;
  assign f_arrdiv32_fs889_and1 = f_arrdiv32_fs889_not1 & f_arrdiv32_fs888_or0;
  assign f_arrdiv32_fs889_or0 = f_arrdiv32_fs889_and1 | f_arrdiv32_fs889_and0;
  assign f_arrdiv32_fs890_xor0 = f_arrdiv32_mux2to1831_xor0 ^ b[26];
  assign f_arrdiv32_fs890_not0 = ~f_arrdiv32_mux2to1831_xor0;
  assign f_arrdiv32_fs890_and0 = f_arrdiv32_fs890_not0 & b[26];
  assign f_arrdiv32_fs890_xor1 = f_arrdiv32_fs889_or0 ^ f_arrdiv32_fs890_xor0;
  assign f_arrdiv32_fs890_not1 = ~f_arrdiv32_fs890_xor0;
  assign f_arrdiv32_fs890_and1 = f_arrdiv32_fs890_not1 & f_arrdiv32_fs889_or0;
  assign f_arrdiv32_fs890_or0 = f_arrdiv32_fs890_and1 | f_arrdiv32_fs890_and0;
  assign f_arrdiv32_fs891_xor0 = f_arrdiv32_mux2to1832_xor0 ^ b[27];
  assign f_arrdiv32_fs891_not0 = ~f_arrdiv32_mux2to1832_xor0;
  assign f_arrdiv32_fs891_and0 = f_arrdiv32_fs891_not0 & b[27];
  assign f_arrdiv32_fs891_xor1 = f_arrdiv32_fs890_or0 ^ f_arrdiv32_fs891_xor0;
  assign f_arrdiv32_fs891_not1 = ~f_arrdiv32_fs891_xor0;
  assign f_arrdiv32_fs891_and1 = f_arrdiv32_fs891_not1 & f_arrdiv32_fs890_or0;
  assign f_arrdiv32_fs891_or0 = f_arrdiv32_fs891_and1 | f_arrdiv32_fs891_and0;
  assign f_arrdiv32_fs892_xor0 = f_arrdiv32_mux2to1833_xor0 ^ b[28];
  assign f_arrdiv32_fs892_not0 = ~f_arrdiv32_mux2to1833_xor0;
  assign f_arrdiv32_fs892_and0 = f_arrdiv32_fs892_not0 & b[28];
  assign f_arrdiv32_fs892_xor1 = f_arrdiv32_fs891_or0 ^ f_arrdiv32_fs892_xor0;
  assign f_arrdiv32_fs892_not1 = ~f_arrdiv32_fs892_xor0;
  assign f_arrdiv32_fs892_and1 = f_arrdiv32_fs892_not1 & f_arrdiv32_fs891_or0;
  assign f_arrdiv32_fs892_or0 = f_arrdiv32_fs892_and1 | f_arrdiv32_fs892_and0;
  assign f_arrdiv32_fs893_xor0 = f_arrdiv32_mux2to1834_xor0 ^ b[29];
  assign f_arrdiv32_fs893_not0 = ~f_arrdiv32_mux2to1834_xor0;
  assign f_arrdiv32_fs893_and0 = f_arrdiv32_fs893_not0 & b[29];
  assign f_arrdiv32_fs893_xor1 = f_arrdiv32_fs892_or0 ^ f_arrdiv32_fs893_xor0;
  assign f_arrdiv32_fs893_not1 = ~f_arrdiv32_fs893_xor0;
  assign f_arrdiv32_fs893_and1 = f_arrdiv32_fs893_not1 & f_arrdiv32_fs892_or0;
  assign f_arrdiv32_fs893_or0 = f_arrdiv32_fs893_and1 | f_arrdiv32_fs893_and0;
  assign f_arrdiv32_fs894_xor0 = f_arrdiv32_mux2to1835_xor0 ^ b[30];
  assign f_arrdiv32_fs894_not0 = ~f_arrdiv32_mux2to1835_xor0;
  assign f_arrdiv32_fs894_and0 = f_arrdiv32_fs894_not0 & b[30];
  assign f_arrdiv32_fs894_xor1 = f_arrdiv32_fs893_or0 ^ f_arrdiv32_fs894_xor0;
  assign f_arrdiv32_fs894_not1 = ~f_arrdiv32_fs894_xor0;
  assign f_arrdiv32_fs894_and1 = f_arrdiv32_fs894_not1 & f_arrdiv32_fs893_or0;
  assign f_arrdiv32_fs894_or0 = f_arrdiv32_fs894_and1 | f_arrdiv32_fs894_and0;
  assign f_arrdiv32_fs895_xor0 = f_arrdiv32_mux2to1836_xor0 ^ b[31];
  assign f_arrdiv32_fs895_not0 = ~f_arrdiv32_mux2to1836_xor0;
  assign f_arrdiv32_fs895_and0 = f_arrdiv32_fs895_not0 & b[31];
  assign f_arrdiv32_fs895_xor1 = f_arrdiv32_fs894_or0 ^ f_arrdiv32_fs895_xor0;
  assign f_arrdiv32_fs895_not1 = ~f_arrdiv32_fs895_xor0;
  assign f_arrdiv32_fs895_and1 = f_arrdiv32_fs895_not1 & f_arrdiv32_fs894_or0;
  assign f_arrdiv32_fs895_or0 = f_arrdiv32_fs895_and1 | f_arrdiv32_fs895_and0;
  assign f_arrdiv32_mux2to1837_and0 = a[4] & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1837_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1837_and1 = f_arrdiv32_fs864_xor0 & f_arrdiv32_mux2to1837_not0;
  assign f_arrdiv32_mux2to1837_xor0 = f_arrdiv32_mux2to1837_and0 ^ f_arrdiv32_mux2to1837_and1;
  assign f_arrdiv32_mux2to1838_and0 = f_arrdiv32_mux2to1806_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1838_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1838_and1 = f_arrdiv32_fs865_xor1 & f_arrdiv32_mux2to1838_not0;
  assign f_arrdiv32_mux2to1838_xor0 = f_arrdiv32_mux2to1838_and0 ^ f_arrdiv32_mux2to1838_and1;
  assign f_arrdiv32_mux2to1839_and0 = f_arrdiv32_mux2to1807_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1839_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1839_and1 = f_arrdiv32_fs866_xor1 & f_arrdiv32_mux2to1839_not0;
  assign f_arrdiv32_mux2to1839_xor0 = f_arrdiv32_mux2to1839_and0 ^ f_arrdiv32_mux2to1839_and1;
  assign f_arrdiv32_mux2to1840_and0 = f_arrdiv32_mux2to1808_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1840_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1840_and1 = f_arrdiv32_fs867_xor1 & f_arrdiv32_mux2to1840_not0;
  assign f_arrdiv32_mux2to1840_xor0 = f_arrdiv32_mux2to1840_and0 ^ f_arrdiv32_mux2to1840_and1;
  assign f_arrdiv32_mux2to1841_and0 = f_arrdiv32_mux2to1809_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1841_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1841_and1 = f_arrdiv32_fs868_xor1 & f_arrdiv32_mux2to1841_not0;
  assign f_arrdiv32_mux2to1841_xor0 = f_arrdiv32_mux2to1841_and0 ^ f_arrdiv32_mux2to1841_and1;
  assign f_arrdiv32_mux2to1842_and0 = f_arrdiv32_mux2to1810_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1842_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1842_and1 = f_arrdiv32_fs869_xor1 & f_arrdiv32_mux2to1842_not0;
  assign f_arrdiv32_mux2to1842_xor0 = f_arrdiv32_mux2to1842_and0 ^ f_arrdiv32_mux2to1842_and1;
  assign f_arrdiv32_mux2to1843_and0 = f_arrdiv32_mux2to1811_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1843_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1843_and1 = f_arrdiv32_fs870_xor1 & f_arrdiv32_mux2to1843_not0;
  assign f_arrdiv32_mux2to1843_xor0 = f_arrdiv32_mux2to1843_and0 ^ f_arrdiv32_mux2to1843_and1;
  assign f_arrdiv32_mux2to1844_and0 = f_arrdiv32_mux2to1812_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1844_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1844_and1 = f_arrdiv32_fs871_xor1 & f_arrdiv32_mux2to1844_not0;
  assign f_arrdiv32_mux2to1844_xor0 = f_arrdiv32_mux2to1844_and0 ^ f_arrdiv32_mux2to1844_and1;
  assign f_arrdiv32_mux2to1845_and0 = f_arrdiv32_mux2to1813_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1845_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1845_and1 = f_arrdiv32_fs872_xor1 & f_arrdiv32_mux2to1845_not0;
  assign f_arrdiv32_mux2to1845_xor0 = f_arrdiv32_mux2to1845_and0 ^ f_arrdiv32_mux2to1845_and1;
  assign f_arrdiv32_mux2to1846_and0 = f_arrdiv32_mux2to1814_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1846_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1846_and1 = f_arrdiv32_fs873_xor1 & f_arrdiv32_mux2to1846_not0;
  assign f_arrdiv32_mux2to1846_xor0 = f_arrdiv32_mux2to1846_and0 ^ f_arrdiv32_mux2to1846_and1;
  assign f_arrdiv32_mux2to1847_and0 = f_arrdiv32_mux2to1815_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1847_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1847_and1 = f_arrdiv32_fs874_xor1 & f_arrdiv32_mux2to1847_not0;
  assign f_arrdiv32_mux2to1847_xor0 = f_arrdiv32_mux2to1847_and0 ^ f_arrdiv32_mux2to1847_and1;
  assign f_arrdiv32_mux2to1848_and0 = f_arrdiv32_mux2to1816_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1848_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1848_and1 = f_arrdiv32_fs875_xor1 & f_arrdiv32_mux2to1848_not0;
  assign f_arrdiv32_mux2to1848_xor0 = f_arrdiv32_mux2to1848_and0 ^ f_arrdiv32_mux2to1848_and1;
  assign f_arrdiv32_mux2to1849_and0 = f_arrdiv32_mux2to1817_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1849_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1849_and1 = f_arrdiv32_fs876_xor1 & f_arrdiv32_mux2to1849_not0;
  assign f_arrdiv32_mux2to1849_xor0 = f_arrdiv32_mux2to1849_and0 ^ f_arrdiv32_mux2to1849_and1;
  assign f_arrdiv32_mux2to1850_and0 = f_arrdiv32_mux2to1818_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1850_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1850_and1 = f_arrdiv32_fs877_xor1 & f_arrdiv32_mux2to1850_not0;
  assign f_arrdiv32_mux2to1850_xor0 = f_arrdiv32_mux2to1850_and0 ^ f_arrdiv32_mux2to1850_and1;
  assign f_arrdiv32_mux2to1851_and0 = f_arrdiv32_mux2to1819_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1851_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1851_and1 = f_arrdiv32_fs878_xor1 & f_arrdiv32_mux2to1851_not0;
  assign f_arrdiv32_mux2to1851_xor0 = f_arrdiv32_mux2to1851_and0 ^ f_arrdiv32_mux2to1851_and1;
  assign f_arrdiv32_mux2to1852_and0 = f_arrdiv32_mux2to1820_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1852_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1852_and1 = f_arrdiv32_fs879_xor1 & f_arrdiv32_mux2to1852_not0;
  assign f_arrdiv32_mux2to1852_xor0 = f_arrdiv32_mux2to1852_and0 ^ f_arrdiv32_mux2to1852_and1;
  assign f_arrdiv32_mux2to1853_and0 = f_arrdiv32_mux2to1821_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1853_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1853_and1 = f_arrdiv32_fs880_xor1 & f_arrdiv32_mux2to1853_not0;
  assign f_arrdiv32_mux2to1853_xor0 = f_arrdiv32_mux2to1853_and0 ^ f_arrdiv32_mux2to1853_and1;
  assign f_arrdiv32_mux2to1854_and0 = f_arrdiv32_mux2to1822_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1854_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1854_and1 = f_arrdiv32_fs881_xor1 & f_arrdiv32_mux2to1854_not0;
  assign f_arrdiv32_mux2to1854_xor0 = f_arrdiv32_mux2to1854_and0 ^ f_arrdiv32_mux2to1854_and1;
  assign f_arrdiv32_mux2to1855_and0 = f_arrdiv32_mux2to1823_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1855_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1855_and1 = f_arrdiv32_fs882_xor1 & f_arrdiv32_mux2to1855_not0;
  assign f_arrdiv32_mux2to1855_xor0 = f_arrdiv32_mux2to1855_and0 ^ f_arrdiv32_mux2to1855_and1;
  assign f_arrdiv32_mux2to1856_and0 = f_arrdiv32_mux2to1824_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1856_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1856_and1 = f_arrdiv32_fs883_xor1 & f_arrdiv32_mux2to1856_not0;
  assign f_arrdiv32_mux2to1856_xor0 = f_arrdiv32_mux2to1856_and0 ^ f_arrdiv32_mux2to1856_and1;
  assign f_arrdiv32_mux2to1857_and0 = f_arrdiv32_mux2to1825_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1857_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1857_and1 = f_arrdiv32_fs884_xor1 & f_arrdiv32_mux2to1857_not0;
  assign f_arrdiv32_mux2to1857_xor0 = f_arrdiv32_mux2to1857_and0 ^ f_arrdiv32_mux2to1857_and1;
  assign f_arrdiv32_mux2to1858_and0 = f_arrdiv32_mux2to1826_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1858_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1858_and1 = f_arrdiv32_fs885_xor1 & f_arrdiv32_mux2to1858_not0;
  assign f_arrdiv32_mux2to1858_xor0 = f_arrdiv32_mux2to1858_and0 ^ f_arrdiv32_mux2to1858_and1;
  assign f_arrdiv32_mux2to1859_and0 = f_arrdiv32_mux2to1827_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1859_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1859_and1 = f_arrdiv32_fs886_xor1 & f_arrdiv32_mux2to1859_not0;
  assign f_arrdiv32_mux2to1859_xor0 = f_arrdiv32_mux2to1859_and0 ^ f_arrdiv32_mux2to1859_and1;
  assign f_arrdiv32_mux2to1860_and0 = f_arrdiv32_mux2to1828_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1860_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1860_and1 = f_arrdiv32_fs887_xor1 & f_arrdiv32_mux2to1860_not0;
  assign f_arrdiv32_mux2to1860_xor0 = f_arrdiv32_mux2to1860_and0 ^ f_arrdiv32_mux2to1860_and1;
  assign f_arrdiv32_mux2to1861_and0 = f_arrdiv32_mux2to1829_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1861_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1861_and1 = f_arrdiv32_fs888_xor1 & f_arrdiv32_mux2to1861_not0;
  assign f_arrdiv32_mux2to1861_xor0 = f_arrdiv32_mux2to1861_and0 ^ f_arrdiv32_mux2to1861_and1;
  assign f_arrdiv32_mux2to1862_and0 = f_arrdiv32_mux2to1830_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1862_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1862_and1 = f_arrdiv32_fs889_xor1 & f_arrdiv32_mux2to1862_not0;
  assign f_arrdiv32_mux2to1862_xor0 = f_arrdiv32_mux2to1862_and0 ^ f_arrdiv32_mux2to1862_and1;
  assign f_arrdiv32_mux2to1863_and0 = f_arrdiv32_mux2to1831_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1863_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1863_and1 = f_arrdiv32_fs890_xor1 & f_arrdiv32_mux2to1863_not0;
  assign f_arrdiv32_mux2to1863_xor0 = f_arrdiv32_mux2to1863_and0 ^ f_arrdiv32_mux2to1863_and1;
  assign f_arrdiv32_mux2to1864_and0 = f_arrdiv32_mux2to1832_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1864_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1864_and1 = f_arrdiv32_fs891_xor1 & f_arrdiv32_mux2to1864_not0;
  assign f_arrdiv32_mux2to1864_xor0 = f_arrdiv32_mux2to1864_and0 ^ f_arrdiv32_mux2to1864_and1;
  assign f_arrdiv32_mux2to1865_and0 = f_arrdiv32_mux2to1833_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1865_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1865_and1 = f_arrdiv32_fs892_xor1 & f_arrdiv32_mux2to1865_not0;
  assign f_arrdiv32_mux2to1865_xor0 = f_arrdiv32_mux2to1865_and0 ^ f_arrdiv32_mux2to1865_and1;
  assign f_arrdiv32_mux2to1866_and0 = f_arrdiv32_mux2to1834_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1866_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1866_and1 = f_arrdiv32_fs893_xor1 & f_arrdiv32_mux2to1866_not0;
  assign f_arrdiv32_mux2to1866_xor0 = f_arrdiv32_mux2to1866_and0 ^ f_arrdiv32_mux2to1866_and1;
  assign f_arrdiv32_mux2to1867_and0 = f_arrdiv32_mux2to1835_xor0 & f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1867_not0 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_mux2to1867_and1 = f_arrdiv32_fs894_xor1 & f_arrdiv32_mux2to1867_not0;
  assign f_arrdiv32_mux2to1867_xor0 = f_arrdiv32_mux2to1867_and0 ^ f_arrdiv32_mux2to1867_and1;
  assign f_arrdiv32_not27 = ~f_arrdiv32_fs895_or0;
  assign f_arrdiv32_fs896_xor0 = a[3] ^ b[0];
  assign f_arrdiv32_fs896_not0 = ~a[3];
  assign f_arrdiv32_fs896_and0 = f_arrdiv32_fs896_not0 & b[0];
  assign f_arrdiv32_fs896_not1 = ~f_arrdiv32_fs896_xor0;
  assign f_arrdiv32_fs897_xor0 = f_arrdiv32_mux2to1837_xor0 ^ b[1];
  assign f_arrdiv32_fs897_not0 = ~f_arrdiv32_mux2to1837_xor0;
  assign f_arrdiv32_fs897_and0 = f_arrdiv32_fs897_not0 & b[1];
  assign f_arrdiv32_fs897_xor1 = f_arrdiv32_fs896_and0 ^ f_arrdiv32_fs897_xor0;
  assign f_arrdiv32_fs897_not1 = ~f_arrdiv32_fs897_xor0;
  assign f_arrdiv32_fs897_and1 = f_arrdiv32_fs897_not1 & f_arrdiv32_fs896_and0;
  assign f_arrdiv32_fs897_or0 = f_arrdiv32_fs897_and1 | f_arrdiv32_fs897_and0;
  assign f_arrdiv32_fs898_xor0 = f_arrdiv32_mux2to1838_xor0 ^ b[2];
  assign f_arrdiv32_fs898_not0 = ~f_arrdiv32_mux2to1838_xor0;
  assign f_arrdiv32_fs898_and0 = f_arrdiv32_fs898_not0 & b[2];
  assign f_arrdiv32_fs898_xor1 = f_arrdiv32_fs897_or0 ^ f_arrdiv32_fs898_xor0;
  assign f_arrdiv32_fs898_not1 = ~f_arrdiv32_fs898_xor0;
  assign f_arrdiv32_fs898_and1 = f_arrdiv32_fs898_not1 & f_arrdiv32_fs897_or0;
  assign f_arrdiv32_fs898_or0 = f_arrdiv32_fs898_and1 | f_arrdiv32_fs898_and0;
  assign f_arrdiv32_fs899_xor0 = f_arrdiv32_mux2to1839_xor0 ^ b[3];
  assign f_arrdiv32_fs899_not0 = ~f_arrdiv32_mux2to1839_xor0;
  assign f_arrdiv32_fs899_and0 = f_arrdiv32_fs899_not0 & b[3];
  assign f_arrdiv32_fs899_xor1 = f_arrdiv32_fs898_or0 ^ f_arrdiv32_fs899_xor0;
  assign f_arrdiv32_fs899_not1 = ~f_arrdiv32_fs899_xor0;
  assign f_arrdiv32_fs899_and1 = f_arrdiv32_fs899_not1 & f_arrdiv32_fs898_or0;
  assign f_arrdiv32_fs899_or0 = f_arrdiv32_fs899_and1 | f_arrdiv32_fs899_and0;
  assign f_arrdiv32_fs900_xor0 = f_arrdiv32_mux2to1840_xor0 ^ b[4];
  assign f_arrdiv32_fs900_not0 = ~f_arrdiv32_mux2to1840_xor0;
  assign f_arrdiv32_fs900_and0 = f_arrdiv32_fs900_not0 & b[4];
  assign f_arrdiv32_fs900_xor1 = f_arrdiv32_fs899_or0 ^ f_arrdiv32_fs900_xor0;
  assign f_arrdiv32_fs900_not1 = ~f_arrdiv32_fs900_xor0;
  assign f_arrdiv32_fs900_and1 = f_arrdiv32_fs900_not1 & f_arrdiv32_fs899_or0;
  assign f_arrdiv32_fs900_or0 = f_arrdiv32_fs900_and1 | f_arrdiv32_fs900_and0;
  assign f_arrdiv32_fs901_xor0 = f_arrdiv32_mux2to1841_xor0 ^ b[5];
  assign f_arrdiv32_fs901_not0 = ~f_arrdiv32_mux2to1841_xor0;
  assign f_arrdiv32_fs901_and0 = f_arrdiv32_fs901_not0 & b[5];
  assign f_arrdiv32_fs901_xor1 = f_arrdiv32_fs900_or0 ^ f_arrdiv32_fs901_xor0;
  assign f_arrdiv32_fs901_not1 = ~f_arrdiv32_fs901_xor0;
  assign f_arrdiv32_fs901_and1 = f_arrdiv32_fs901_not1 & f_arrdiv32_fs900_or0;
  assign f_arrdiv32_fs901_or0 = f_arrdiv32_fs901_and1 | f_arrdiv32_fs901_and0;
  assign f_arrdiv32_fs902_xor0 = f_arrdiv32_mux2to1842_xor0 ^ b[6];
  assign f_arrdiv32_fs902_not0 = ~f_arrdiv32_mux2to1842_xor0;
  assign f_arrdiv32_fs902_and0 = f_arrdiv32_fs902_not0 & b[6];
  assign f_arrdiv32_fs902_xor1 = f_arrdiv32_fs901_or0 ^ f_arrdiv32_fs902_xor0;
  assign f_arrdiv32_fs902_not1 = ~f_arrdiv32_fs902_xor0;
  assign f_arrdiv32_fs902_and1 = f_arrdiv32_fs902_not1 & f_arrdiv32_fs901_or0;
  assign f_arrdiv32_fs902_or0 = f_arrdiv32_fs902_and1 | f_arrdiv32_fs902_and0;
  assign f_arrdiv32_fs903_xor0 = f_arrdiv32_mux2to1843_xor0 ^ b[7];
  assign f_arrdiv32_fs903_not0 = ~f_arrdiv32_mux2to1843_xor0;
  assign f_arrdiv32_fs903_and0 = f_arrdiv32_fs903_not0 & b[7];
  assign f_arrdiv32_fs903_xor1 = f_arrdiv32_fs902_or0 ^ f_arrdiv32_fs903_xor0;
  assign f_arrdiv32_fs903_not1 = ~f_arrdiv32_fs903_xor0;
  assign f_arrdiv32_fs903_and1 = f_arrdiv32_fs903_not1 & f_arrdiv32_fs902_or0;
  assign f_arrdiv32_fs903_or0 = f_arrdiv32_fs903_and1 | f_arrdiv32_fs903_and0;
  assign f_arrdiv32_fs904_xor0 = f_arrdiv32_mux2to1844_xor0 ^ b[8];
  assign f_arrdiv32_fs904_not0 = ~f_arrdiv32_mux2to1844_xor0;
  assign f_arrdiv32_fs904_and0 = f_arrdiv32_fs904_not0 & b[8];
  assign f_arrdiv32_fs904_xor1 = f_arrdiv32_fs903_or0 ^ f_arrdiv32_fs904_xor0;
  assign f_arrdiv32_fs904_not1 = ~f_arrdiv32_fs904_xor0;
  assign f_arrdiv32_fs904_and1 = f_arrdiv32_fs904_not1 & f_arrdiv32_fs903_or0;
  assign f_arrdiv32_fs904_or0 = f_arrdiv32_fs904_and1 | f_arrdiv32_fs904_and0;
  assign f_arrdiv32_fs905_xor0 = f_arrdiv32_mux2to1845_xor0 ^ b[9];
  assign f_arrdiv32_fs905_not0 = ~f_arrdiv32_mux2to1845_xor0;
  assign f_arrdiv32_fs905_and0 = f_arrdiv32_fs905_not0 & b[9];
  assign f_arrdiv32_fs905_xor1 = f_arrdiv32_fs904_or0 ^ f_arrdiv32_fs905_xor0;
  assign f_arrdiv32_fs905_not1 = ~f_arrdiv32_fs905_xor0;
  assign f_arrdiv32_fs905_and1 = f_arrdiv32_fs905_not1 & f_arrdiv32_fs904_or0;
  assign f_arrdiv32_fs905_or0 = f_arrdiv32_fs905_and1 | f_arrdiv32_fs905_and0;
  assign f_arrdiv32_fs906_xor0 = f_arrdiv32_mux2to1846_xor0 ^ b[10];
  assign f_arrdiv32_fs906_not0 = ~f_arrdiv32_mux2to1846_xor0;
  assign f_arrdiv32_fs906_and0 = f_arrdiv32_fs906_not0 & b[10];
  assign f_arrdiv32_fs906_xor1 = f_arrdiv32_fs905_or0 ^ f_arrdiv32_fs906_xor0;
  assign f_arrdiv32_fs906_not1 = ~f_arrdiv32_fs906_xor0;
  assign f_arrdiv32_fs906_and1 = f_arrdiv32_fs906_not1 & f_arrdiv32_fs905_or0;
  assign f_arrdiv32_fs906_or0 = f_arrdiv32_fs906_and1 | f_arrdiv32_fs906_and0;
  assign f_arrdiv32_fs907_xor0 = f_arrdiv32_mux2to1847_xor0 ^ b[11];
  assign f_arrdiv32_fs907_not0 = ~f_arrdiv32_mux2to1847_xor0;
  assign f_arrdiv32_fs907_and0 = f_arrdiv32_fs907_not0 & b[11];
  assign f_arrdiv32_fs907_xor1 = f_arrdiv32_fs906_or0 ^ f_arrdiv32_fs907_xor0;
  assign f_arrdiv32_fs907_not1 = ~f_arrdiv32_fs907_xor0;
  assign f_arrdiv32_fs907_and1 = f_arrdiv32_fs907_not1 & f_arrdiv32_fs906_or0;
  assign f_arrdiv32_fs907_or0 = f_arrdiv32_fs907_and1 | f_arrdiv32_fs907_and0;
  assign f_arrdiv32_fs908_xor0 = f_arrdiv32_mux2to1848_xor0 ^ b[12];
  assign f_arrdiv32_fs908_not0 = ~f_arrdiv32_mux2to1848_xor0;
  assign f_arrdiv32_fs908_and0 = f_arrdiv32_fs908_not0 & b[12];
  assign f_arrdiv32_fs908_xor1 = f_arrdiv32_fs907_or0 ^ f_arrdiv32_fs908_xor0;
  assign f_arrdiv32_fs908_not1 = ~f_arrdiv32_fs908_xor0;
  assign f_arrdiv32_fs908_and1 = f_arrdiv32_fs908_not1 & f_arrdiv32_fs907_or0;
  assign f_arrdiv32_fs908_or0 = f_arrdiv32_fs908_and1 | f_arrdiv32_fs908_and0;
  assign f_arrdiv32_fs909_xor0 = f_arrdiv32_mux2to1849_xor0 ^ b[13];
  assign f_arrdiv32_fs909_not0 = ~f_arrdiv32_mux2to1849_xor0;
  assign f_arrdiv32_fs909_and0 = f_arrdiv32_fs909_not0 & b[13];
  assign f_arrdiv32_fs909_xor1 = f_arrdiv32_fs908_or0 ^ f_arrdiv32_fs909_xor0;
  assign f_arrdiv32_fs909_not1 = ~f_arrdiv32_fs909_xor0;
  assign f_arrdiv32_fs909_and1 = f_arrdiv32_fs909_not1 & f_arrdiv32_fs908_or0;
  assign f_arrdiv32_fs909_or0 = f_arrdiv32_fs909_and1 | f_arrdiv32_fs909_and0;
  assign f_arrdiv32_fs910_xor0 = f_arrdiv32_mux2to1850_xor0 ^ b[14];
  assign f_arrdiv32_fs910_not0 = ~f_arrdiv32_mux2to1850_xor0;
  assign f_arrdiv32_fs910_and0 = f_arrdiv32_fs910_not0 & b[14];
  assign f_arrdiv32_fs910_xor1 = f_arrdiv32_fs909_or0 ^ f_arrdiv32_fs910_xor0;
  assign f_arrdiv32_fs910_not1 = ~f_arrdiv32_fs910_xor0;
  assign f_arrdiv32_fs910_and1 = f_arrdiv32_fs910_not1 & f_arrdiv32_fs909_or0;
  assign f_arrdiv32_fs910_or0 = f_arrdiv32_fs910_and1 | f_arrdiv32_fs910_and0;
  assign f_arrdiv32_fs911_xor0 = f_arrdiv32_mux2to1851_xor0 ^ b[15];
  assign f_arrdiv32_fs911_not0 = ~f_arrdiv32_mux2to1851_xor0;
  assign f_arrdiv32_fs911_and0 = f_arrdiv32_fs911_not0 & b[15];
  assign f_arrdiv32_fs911_xor1 = f_arrdiv32_fs910_or0 ^ f_arrdiv32_fs911_xor0;
  assign f_arrdiv32_fs911_not1 = ~f_arrdiv32_fs911_xor0;
  assign f_arrdiv32_fs911_and1 = f_arrdiv32_fs911_not1 & f_arrdiv32_fs910_or0;
  assign f_arrdiv32_fs911_or0 = f_arrdiv32_fs911_and1 | f_arrdiv32_fs911_and0;
  assign f_arrdiv32_fs912_xor0 = f_arrdiv32_mux2to1852_xor0 ^ b[16];
  assign f_arrdiv32_fs912_not0 = ~f_arrdiv32_mux2to1852_xor0;
  assign f_arrdiv32_fs912_and0 = f_arrdiv32_fs912_not0 & b[16];
  assign f_arrdiv32_fs912_xor1 = f_arrdiv32_fs911_or0 ^ f_arrdiv32_fs912_xor0;
  assign f_arrdiv32_fs912_not1 = ~f_arrdiv32_fs912_xor0;
  assign f_arrdiv32_fs912_and1 = f_arrdiv32_fs912_not1 & f_arrdiv32_fs911_or0;
  assign f_arrdiv32_fs912_or0 = f_arrdiv32_fs912_and1 | f_arrdiv32_fs912_and0;
  assign f_arrdiv32_fs913_xor0 = f_arrdiv32_mux2to1853_xor0 ^ b[17];
  assign f_arrdiv32_fs913_not0 = ~f_arrdiv32_mux2to1853_xor0;
  assign f_arrdiv32_fs913_and0 = f_arrdiv32_fs913_not0 & b[17];
  assign f_arrdiv32_fs913_xor1 = f_arrdiv32_fs912_or0 ^ f_arrdiv32_fs913_xor0;
  assign f_arrdiv32_fs913_not1 = ~f_arrdiv32_fs913_xor0;
  assign f_arrdiv32_fs913_and1 = f_arrdiv32_fs913_not1 & f_arrdiv32_fs912_or0;
  assign f_arrdiv32_fs913_or0 = f_arrdiv32_fs913_and1 | f_arrdiv32_fs913_and0;
  assign f_arrdiv32_fs914_xor0 = f_arrdiv32_mux2to1854_xor0 ^ b[18];
  assign f_arrdiv32_fs914_not0 = ~f_arrdiv32_mux2to1854_xor0;
  assign f_arrdiv32_fs914_and0 = f_arrdiv32_fs914_not0 & b[18];
  assign f_arrdiv32_fs914_xor1 = f_arrdiv32_fs913_or0 ^ f_arrdiv32_fs914_xor0;
  assign f_arrdiv32_fs914_not1 = ~f_arrdiv32_fs914_xor0;
  assign f_arrdiv32_fs914_and1 = f_arrdiv32_fs914_not1 & f_arrdiv32_fs913_or0;
  assign f_arrdiv32_fs914_or0 = f_arrdiv32_fs914_and1 | f_arrdiv32_fs914_and0;
  assign f_arrdiv32_fs915_xor0 = f_arrdiv32_mux2to1855_xor0 ^ b[19];
  assign f_arrdiv32_fs915_not0 = ~f_arrdiv32_mux2to1855_xor0;
  assign f_arrdiv32_fs915_and0 = f_arrdiv32_fs915_not0 & b[19];
  assign f_arrdiv32_fs915_xor1 = f_arrdiv32_fs914_or0 ^ f_arrdiv32_fs915_xor0;
  assign f_arrdiv32_fs915_not1 = ~f_arrdiv32_fs915_xor0;
  assign f_arrdiv32_fs915_and1 = f_arrdiv32_fs915_not1 & f_arrdiv32_fs914_or0;
  assign f_arrdiv32_fs915_or0 = f_arrdiv32_fs915_and1 | f_arrdiv32_fs915_and0;
  assign f_arrdiv32_fs916_xor0 = f_arrdiv32_mux2to1856_xor0 ^ b[20];
  assign f_arrdiv32_fs916_not0 = ~f_arrdiv32_mux2to1856_xor0;
  assign f_arrdiv32_fs916_and0 = f_arrdiv32_fs916_not0 & b[20];
  assign f_arrdiv32_fs916_xor1 = f_arrdiv32_fs915_or0 ^ f_arrdiv32_fs916_xor0;
  assign f_arrdiv32_fs916_not1 = ~f_arrdiv32_fs916_xor0;
  assign f_arrdiv32_fs916_and1 = f_arrdiv32_fs916_not1 & f_arrdiv32_fs915_or0;
  assign f_arrdiv32_fs916_or0 = f_arrdiv32_fs916_and1 | f_arrdiv32_fs916_and0;
  assign f_arrdiv32_fs917_xor0 = f_arrdiv32_mux2to1857_xor0 ^ b[21];
  assign f_arrdiv32_fs917_not0 = ~f_arrdiv32_mux2to1857_xor0;
  assign f_arrdiv32_fs917_and0 = f_arrdiv32_fs917_not0 & b[21];
  assign f_arrdiv32_fs917_xor1 = f_arrdiv32_fs916_or0 ^ f_arrdiv32_fs917_xor0;
  assign f_arrdiv32_fs917_not1 = ~f_arrdiv32_fs917_xor0;
  assign f_arrdiv32_fs917_and1 = f_arrdiv32_fs917_not1 & f_arrdiv32_fs916_or0;
  assign f_arrdiv32_fs917_or0 = f_arrdiv32_fs917_and1 | f_arrdiv32_fs917_and0;
  assign f_arrdiv32_fs918_xor0 = f_arrdiv32_mux2to1858_xor0 ^ b[22];
  assign f_arrdiv32_fs918_not0 = ~f_arrdiv32_mux2to1858_xor0;
  assign f_arrdiv32_fs918_and0 = f_arrdiv32_fs918_not0 & b[22];
  assign f_arrdiv32_fs918_xor1 = f_arrdiv32_fs917_or0 ^ f_arrdiv32_fs918_xor0;
  assign f_arrdiv32_fs918_not1 = ~f_arrdiv32_fs918_xor0;
  assign f_arrdiv32_fs918_and1 = f_arrdiv32_fs918_not1 & f_arrdiv32_fs917_or0;
  assign f_arrdiv32_fs918_or0 = f_arrdiv32_fs918_and1 | f_arrdiv32_fs918_and0;
  assign f_arrdiv32_fs919_xor0 = f_arrdiv32_mux2to1859_xor0 ^ b[23];
  assign f_arrdiv32_fs919_not0 = ~f_arrdiv32_mux2to1859_xor0;
  assign f_arrdiv32_fs919_and0 = f_arrdiv32_fs919_not0 & b[23];
  assign f_arrdiv32_fs919_xor1 = f_arrdiv32_fs918_or0 ^ f_arrdiv32_fs919_xor0;
  assign f_arrdiv32_fs919_not1 = ~f_arrdiv32_fs919_xor0;
  assign f_arrdiv32_fs919_and1 = f_arrdiv32_fs919_not1 & f_arrdiv32_fs918_or0;
  assign f_arrdiv32_fs919_or0 = f_arrdiv32_fs919_and1 | f_arrdiv32_fs919_and0;
  assign f_arrdiv32_fs920_xor0 = f_arrdiv32_mux2to1860_xor0 ^ b[24];
  assign f_arrdiv32_fs920_not0 = ~f_arrdiv32_mux2to1860_xor0;
  assign f_arrdiv32_fs920_and0 = f_arrdiv32_fs920_not0 & b[24];
  assign f_arrdiv32_fs920_xor1 = f_arrdiv32_fs919_or0 ^ f_arrdiv32_fs920_xor0;
  assign f_arrdiv32_fs920_not1 = ~f_arrdiv32_fs920_xor0;
  assign f_arrdiv32_fs920_and1 = f_arrdiv32_fs920_not1 & f_arrdiv32_fs919_or0;
  assign f_arrdiv32_fs920_or0 = f_arrdiv32_fs920_and1 | f_arrdiv32_fs920_and0;
  assign f_arrdiv32_fs921_xor0 = f_arrdiv32_mux2to1861_xor0 ^ b[25];
  assign f_arrdiv32_fs921_not0 = ~f_arrdiv32_mux2to1861_xor0;
  assign f_arrdiv32_fs921_and0 = f_arrdiv32_fs921_not0 & b[25];
  assign f_arrdiv32_fs921_xor1 = f_arrdiv32_fs920_or0 ^ f_arrdiv32_fs921_xor0;
  assign f_arrdiv32_fs921_not1 = ~f_arrdiv32_fs921_xor0;
  assign f_arrdiv32_fs921_and1 = f_arrdiv32_fs921_not1 & f_arrdiv32_fs920_or0;
  assign f_arrdiv32_fs921_or0 = f_arrdiv32_fs921_and1 | f_arrdiv32_fs921_and0;
  assign f_arrdiv32_fs922_xor0 = f_arrdiv32_mux2to1862_xor0 ^ b[26];
  assign f_arrdiv32_fs922_not0 = ~f_arrdiv32_mux2to1862_xor0;
  assign f_arrdiv32_fs922_and0 = f_arrdiv32_fs922_not0 & b[26];
  assign f_arrdiv32_fs922_xor1 = f_arrdiv32_fs921_or0 ^ f_arrdiv32_fs922_xor0;
  assign f_arrdiv32_fs922_not1 = ~f_arrdiv32_fs922_xor0;
  assign f_arrdiv32_fs922_and1 = f_arrdiv32_fs922_not1 & f_arrdiv32_fs921_or0;
  assign f_arrdiv32_fs922_or0 = f_arrdiv32_fs922_and1 | f_arrdiv32_fs922_and0;
  assign f_arrdiv32_fs923_xor0 = f_arrdiv32_mux2to1863_xor0 ^ b[27];
  assign f_arrdiv32_fs923_not0 = ~f_arrdiv32_mux2to1863_xor0;
  assign f_arrdiv32_fs923_and0 = f_arrdiv32_fs923_not0 & b[27];
  assign f_arrdiv32_fs923_xor1 = f_arrdiv32_fs922_or0 ^ f_arrdiv32_fs923_xor0;
  assign f_arrdiv32_fs923_not1 = ~f_arrdiv32_fs923_xor0;
  assign f_arrdiv32_fs923_and1 = f_arrdiv32_fs923_not1 & f_arrdiv32_fs922_or0;
  assign f_arrdiv32_fs923_or0 = f_arrdiv32_fs923_and1 | f_arrdiv32_fs923_and0;
  assign f_arrdiv32_fs924_xor0 = f_arrdiv32_mux2to1864_xor0 ^ b[28];
  assign f_arrdiv32_fs924_not0 = ~f_arrdiv32_mux2to1864_xor0;
  assign f_arrdiv32_fs924_and0 = f_arrdiv32_fs924_not0 & b[28];
  assign f_arrdiv32_fs924_xor1 = f_arrdiv32_fs923_or0 ^ f_arrdiv32_fs924_xor0;
  assign f_arrdiv32_fs924_not1 = ~f_arrdiv32_fs924_xor0;
  assign f_arrdiv32_fs924_and1 = f_arrdiv32_fs924_not1 & f_arrdiv32_fs923_or0;
  assign f_arrdiv32_fs924_or0 = f_arrdiv32_fs924_and1 | f_arrdiv32_fs924_and0;
  assign f_arrdiv32_fs925_xor0 = f_arrdiv32_mux2to1865_xor0 ^ b[29];
  assign f_arrdiv32_fs925_not0 = ~f_arrdiv32_mux2to1865_xor0;
  assign f_arrdiv32_fs925_and0 = f_arrdiv32_fs925_not0 & b[29];
  assign f_arrdiv32_fs925_xor1 = f_arrdiv32_fs924_or0 ^ f_arrdiv32_fs925_xor0;
  assign f_arrdiv32_fs925_not1 = ~f_arrdiv32_fs925_xor0;
  assign f_arrdiv32_fs925_and1 = f_arrdiv32_fs925_not1 & f_arrdiv32_fs924_or0;
  assign f_arrdiv32_fs925_or0 = f_arrdiv32_fs925_and1 | f_arrdiv32_fs925_and0;
  assign f_arrdiv32_fs926_xor0 = f_arrdiv32_mux2to1866_xor0 ^ b[30];
  assign f_arrdiv32_fs926_not0 = ~f_arrdiv32_mux2to1866_xor0;
  assign f_arrdiv32_fs926_and0 = f_arrdiv32_fs926_not0 & b[30];
  assign f_arrdiv32_fs926_xor1 = f_arrdiv32_fs925_or0 ^ f_arrdiv32_fs926_xor0;
  assign f_arrdiv32_fs926_not1 = ~f_arrdiv32_fs926_xor0;
  assign f_arrdiv32_fs926_and1 = f_arrdiv32_fs926_not1 & f_arrdiv32_fs925_or0;
  assign f_arrdiv32_fs926_or0 = f_arrdiv32_fs926_and1 | f_arrdiv32_fs926_and0;
  assign f_arrdiv32_fs927_xor0 = f_arrdiv32_mux2to1867_xor0 ^ b[31];
  assign f_arrdiv32_fs927_not0 = ~f_arrdiv32_mux2to1867_xor0;
  assign f_arrdiv32_fs927_and0 = f_arrdiv32_fs927_not0 & b[31];
  assign f_arrdiv32_fs927_xor1 = f_arrdiv32_fs926_or0 ^ f_arrdiv32_fs927_xor0;
  assign f_arrdiv32_fs927_not1 = ~f_arrdiv32_fs927_xor0;
  assign f_arrdiv32_fs927_and1 = f_arrdiv32_fs927_not1 & f_arrdiv32_fs926_or0;
  assign f_arrdiv32_fs927_or0 = f_arrdiv32_fs927_and1 | f_arrdiv32_fs927_and0;
  assign f_arrdiv32_mux2to1868_and0 = a[3] & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1868_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1868_and1 = f_arrdiv32_fs896_xor0 & f_arrdiv32_mux2to1868_not0;
  assign f_arrdiv32_mux2to1868_xor0 = f_arrdiv32_mux2to1868_and0 ^ f_arrdiv32_mux2to1868_and1;
  assign f_arrdiv32_mux2to1869_and0 = f_arrdiv32_mux2to1837_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1869_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1869_and1 = f_arrdiv32_fs897_xor1 & f_arrdiv32_mux2to1869_not0;
  assign f_arrdiv32_mux2to1869_xor0 = f_arrdiv32_mux2to1869_and0 ^ f_arrdiv32_mux2to1869_and1;
  assign f_arrdiv32_mux2to1870_and0 = f_arrdiv32_mux2to1838_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1870_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1870_and1 = f_arrdiv32_fs898_xor1 & f_arrdiv32_mux2to1870_not0;
  assign f_arrdiv32_mux2to1870_xor0 = f_arrdiv32_mux2to1870_and0 ^ f_arrdiv32_mux2to1870_and1;
  assign f_arrdiv32_mux2to1871_and0 = f_arrdiv32_mux2to1839_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1871_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1871_and1 = f_arrdiv32_fs899_xor1 & f_arrdiv32_mux2to1871_not0;
  assign f_arrdiv32_mux2to1871_xor0 = f_arrdiv32_mux2to1871_and0 ^ f_arrdiv32_mux2to1871_and1;
  assign f_arrdiv32_mux2to1872_and0 = f_arrdiv32_mux2to1840_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1872_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1872_and1 = f_arrdiv32_fs900_xor1 & f_arrdiv32_mux2to1872_not0;
  assign f_arrdiv32_mux2to1872_xor0 = f_arrdiv32_mux2to1872_and0 ^ f_arrdiv32_mux2to1872_and1;
  assign f_arrdiv32_mux2to1873_and0 = f_arrdiv32_mux2to1841_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1873_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1873_and1 = f_arrdiv32_fs901_xor1 & f_arrdiv32_mux2to1873_not0;
  assign f_arrdiv32_mux2to1873_xor0 = f_arrdiv32_mux2to1873_and0 ^ f_arrdiv32_mux2to1873_and1;
  assign f_arrdiv32_mux2to1874_and0 = f_arrdiv32_mux2to1842_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1874_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1874_and1 = f_arrdiv32_fs902_xor1 & f_arrdiv32_mux2to1874_not0;
  assign f_arrdiv32_mux2to1874_xor0 = f_arrdiv32_mux2to1874_and0 ^ f_arrdiv32_mux2to1874_and1;
  assign f_arrdiv32_mux2to1875_and0 = f_arrdiv32_mux2to1843_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1875_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1875_and1 = f_arrdiv32_fs903_xor1 & f_arrdiv32_mux2to1875_not0;
  assign f_arrdiv32_mux2to1875_xor0 = f_arrdiv32_mux2to1875_and0 ^ f_arrdiv32_mux2to1875_and1;
  assign f_arrdiv32_mux2to1876_and0 = f_arrdiv32_mux2to1844_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1876_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1876_and1 = f_arrdiv32_fs904_xor1 & f_arrdiv32_mux2to1876_not0;
  assign f_arrdiv32_mux2to1876_xor0 = f_arrdiv32_mux2to1876_and0 ^ f_arrdiv32_mux2to1876_and1;
  assign f_arrdiv32_mux2to1877_and0 = f_arrdiv32_mux2to1845_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1877_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1877_and1 = f_arrdiv32_fs905_xor1 & f_arrdiv32_mux2to1877_not0;
  assign f_arrdiv32_mux2to1877_xor0 = f_arrdiv32_mux2to1877_and0 ^ f_arrdiv32_mux2to1877_and1;
  assign f_arrdiv32_mux2to1878_and0 = f_arrdiv32_mux2to1846_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1878_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1878_and1 = f_arrdiv32_fs906_xor1 & f_arrdiv32_mux2to1878_not0;
  assign f_arrdiv32_mux2to1878_xor0 = f_arrdiv32_mux2to1878_and0 ^ f_arrdiv32_mux2to1878_and1;
  assign f_arrdiv32_mux2to1879_and0 = f_arrdiv32_mux2to1847_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1879_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1879_and1 = f_arrdiv32_fs907_xor1 & f_arrdiv32_mux2to1879_not0;
  assign f_arrdiv32_mux2to1879_xor0 = f_arrdiv32_mux2to1879_and0 ^ f_arrdiv32_mux2to1879_and1;
  assign f_arrdiv32_mux2to1880_and0 = f_arrdiv32_mux2to1848_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1880_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1880_and1 = f_arrdiv32_fs908_xor1 & f_arrdiv32_mux2to1880_not0;
  assign f_arrdiv32_mux2to1880_xor0 = f_arrdiv32_mux2to1880_and0 ^ f_arrdiv32_mux2to1880_and1;
  assign f_arrdiv32_mux2to1881_and0 = f_arrdiv32_mux2to1849_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1881_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1881_and1 = f_arrdiv32_fs909_xor1 & f_arrdiv32_mux2to1881_not0;
  assign f_arrdiv32_mux2to1881_xor0 = f_arrdiv32_mux2to1881_and0 ^ f_arrdiv32_mux2to1881_and1;
  assign f_arrdiv32_mux2to1882_and0 = f_arrdiv32_mux2to1850_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1882_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1882_and1 = f_arrdiv32_fs910_xor1 & f_arrdiv32_mux2to1882_not0;
  assign f_arrdiv32_mux2to1882_xor0 = f_arrdiv32_mux2to1882_and0 ^ f_arrdiv32_mux2to1882_and1;
  assign f_arrdiv32_mux2to1883_and0 = f_arrdiv32_mux2to1851_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1883_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1883_and1 = f_arrdiv32_fs911_xor1 & f_arrdiv32_mux2to1883_not0;
  assign f_arrdiv32_mux2to1883_xor0 = f_arrdiv32_mux2to1883_and0 ^ f_arrdiv32_mux2to1883_and1;
  assign f_arrdiv32_mux2to1884_and0 = f_arrdiv32_mux2to1852_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1884_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1884_and1 = f_arrdiv32_fs912_xor1 & f_arrdiv32_mux2to1884_not0;
  assign f_arrdiv32_mux2to1884_xor0 = f_arrdiv32_mux2to1884_and0 ^ f_arrdiv32_mux2to1884_and1;
  assign f_arrdiv32_mux2to1885_and0 = f_arrdiv32_mux2to1853_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1885_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1885_and1 = f_arrdiv32_fs913_xor1 & f_arrdiv32_mux2to1885_not0;
  assign f_arrdiv32_mux2to1885_xor0 = f_arrdiv32_mux2to1885_and0 ^ f_arrdiv32_mux2to1885_and1;
  assign f_arrdiv32_mux2to1886_and0 = f_arrdiv32_mux2to1854_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1886_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1886_and1 = f_arrdiv32_fs914_xor1 & f_arrdiv32_mux2to1886_not0;
  assign f_arrdiv32_mux2to1886_xor0 = f_arrdiv32_mux2to1886_and0 ^ f_arrdiv32_mux2to1886_and1;
  assign f_arrdiv32_mux2to1887_and0 = f_arrdiv32_mux2to1855_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1887_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1887_and1 = f_arrdiv32_fs915_xor1 & f_arrdiv32_mux2to1887_not0;
  assign f_arrdiv32_mux2to1887_xor0 = f_arrdiv32_mux2to1887_and0 ^ f_arrdiv32_mux2to1887_and1;
  assign f_arrdiv32_mux2to1888_and0 = f_arrdiv32_mux2to1856_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1888_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1888_and1 = f_arrdiv32_fs916_xor1 & f_arrdiv32_mux2to1888_not0;
  assign f_arrdiv32_mux2to1888_xor0 = f_arrdiv32_mux2to1888_and0 ^ f_arrdiv32_mux2to1888_and1;
  assign f_arrdiv32_mux2to1889_and0 = f_arrdiv32_mux2to1857_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1889_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1889_and1 = f_arrdiv32_fs917_xor1 & f_arrdiv32_mux2to1889_not0;
  assign f_arrdiv32_mux2to1889_xor0 = f_arrdiv32_mux2to1889_and0 ^ f_arrdiv32_mux2to1889_and1;
  assign f_arrdiv32_mux2to1890_and0 = f_arrdiv32_mux2to1858_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1890_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1890_and1 = f_arrdiv32_fs918_xor1 & f_arrdiv32_mux2to1890_not0;
  assign f_arrdiv32_mux2to1890_xor0 = f_arrdiv32_mux2to1890_and0 ^ f_arrdiv32_mux2to1890_and1;
  assign f_arrdiv32_mux2to1891_and0 = f_arrdiv32_mux2to1859_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1891_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1891_and1 = f_arrdiv32_fs919_xor1 & f_arrdiv32_mux2to1891_not0;
  assign f_arrdiv32_mux2to1891_xor0 = f_arrdiv32_mux2to1891_and0 ^ f_arrdiv32_mux2to1891_and1;
  assign f_arrdiv32_mux2to1892_and0 = f_arrdiv32_mux2to1860_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1892_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1892_and1 = f_arrdiv32_fs920_xor1 & f_arrdiv32_mux2to1892_not0;
  assign f_arrdiv32_mux2to1892_xor0 = f_arrdiv32_mux2to1892_and0 ^ f_arrdiv32_mux2to1892_and1;
  assign f_arrdiv32_mux2to1893_and0 = f_arrdiv32_mux2to1861_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1893_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1893_and1 = f_arrdiv32_fs921_xor1 & f_arrdiv32_mux2to1893_not0;
  assign f_arrdiv32_mux2to1893_xor0 = f_arrdiv32_mux2to1893_and0 ^ f_arrdiv32_mux2to1893_and1;
  assign f_arrdiv32_mux2to1894_and0 = f_arrdiv32_mux2to1862_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1894_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1894_and1 = f_arrdiv32_fs922_xor1 & f_arrdiv32_mux2to1894_not0;
  assign f_arrdiv32_mux2to1894_xor0 = f_arrdiv32_mux2to1894_and0 ^ f_arrdiv32_mux2to1894_and1;
  assign f_arrdiv32_mux2to1895_and0 = f_arrdiv32_mux2to1863_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1895_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1895_and1 = f_arrdiv32_fs923_xor1 & f_arrdiv32_mux2to1895_not0;
  assign f_arrdiv32_mux2to1895_xor0 = f_arrdiv32_mux2to1895_and0 ^ f_arrdiv32_mux2to1895_and1;
  assign f_arrdiv32_mux2to1896_and0 = f_arrdiv32_mux2to1864_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1896_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1896_and1 = f_arrdiv32_fs924_xor1 & f_arrdiv32_mux2to1896_not0;
  assign f_arrdiv32_mux2to1896_xor0 = f_arrdiv32_mux2to1896_and0 ^ f_arrdiv32_mux2to1896_and1;
  assign f_arrdiv32_mux2to1897_and0 = f_arrdiv32_mux2to1865_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1897_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1897_and1 = f_arrdiv32_fs925_xor1 & f_arrdiv32_mux2to1897_not0;
  assign f_arrdiv32_mux2to1897_xor0 = f_arrdiv32_mux2to1897_and0 ^ f_arrdiv32_mux2to1897_and1;
  assign f_arrdiv32_mux2to1898_and0 = f_arrdiv32_mux2to1866_xor0 & f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1898_not0 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_mux2to1898_and1 = f_arrdiv32_fs926_xor1 & f_arrdiv32_mux2to1898_not0;
  assign f_arrdiv32_mux2to1898_xor0 = f_arrdiv32_mux2to1898_and0 ^ f_arrdiv32_mux2to1898_and1;
  assign f_arrdiv32_not28 = ~f_arrdiv32_fs927_or0;
  assign f_arrdiv32_fs928_xor0 = a[2] ^ b[0];
  assign f_arrdiv32_fs928_not0 = ~a[2];
  assign f_arrdiv32_fs928_and0 = f_arrdiv32_fs928_not0 & b[0];
  assign f_arrdiv32_fs928_not1 = ~f_arrdiv32_fs928_xor0;
  assign f_arrdiv32_fs929_xor0 = f_arrdiv32_mux2to1868_xor0 ^ b[1];
  assign f_arrdiv32_fs929_not0 = ~f_arrdiv32_mux2to1868_xor0;
  assign f_arrdiv32_fs929_and0 = f_arrdiv32_fs929_not0 & b[1];
  assign f_arrdiv32_fs929_xor1 = f_arrdiv32_fs928_and0 ^ f_arrdiv32_fs929_xor0;
  assign f_arrdiv32_fs929_not1 = ~f_arrdiv32_fs929_xor0;
  assign f_arrdiv32_fs929_and1 = f_arrdiv32_fs929_not1 & f_arrdiv32_fs928_and0;
  assign f_arrdiv32_fs929_or0 = f_arrdiv32_fs929_and1 | f_arrdiv32_fs929_and0;
  assign f_arrdiv32_fs930_xor0 = f_arrdiv32_mux2to1869_xor0 ^ b[2];
  assign f_arrdiv32_fs930_not0 = ~f_arrdiv32_mux2to1869_xor0;
  assign f_arrdiv32_fs930_and0 = f_arrdiv32_fs930_not0 & b[2];
  assign f_arrdiv32_fs930_xor1 = f_arrdiv32_fs929_or0 ^ f_arrdiv32_fs930_xor0;
  assign f_arrdiv32_fs930_not1 = ~f_arrdiv32_fs930_xor0;
  assign f_arrdiv32_fs930_and1 = f_arrdiv32_fs930_not1 & f_arrdiv32_fs929_or0;
  assign f_arrdiv32_fs930_or0 = f_arrdiv32_fs930_and1 | f_arrdiv32_fs930_and0;
  assign f_arrdiv32_fs931_xor0 = f_arrdiv32_mux2to1870_xor0 ^ b[3];
  assign f_arrdiv32_fs931_not0 = ~f_arrdiv32_mux2to1870_xor0;
  assign f_arrdiv32_fs931_and0 = f_arrdiv32_fs931_not0 & b[3];
  assign f_arrdiv32_fs931_xor1 = f_arrdiv32_fs930_or0 ^ f_arrdiv32_fs931_xor0;
  assign f_arrdiv32_fs931_not1 = ~f_arrdiv32_fs931_xor0;
  assign f_arrdiv32_fs931_and1 = f_arrdiv32_fs931_not1 & f_arrdiv32_fs930_or0;
  assign f_arrdiv32_fs931_or0 = f_arrdiv32_fs931_and1 | f_arrdiv32_fs931_and0;
  assign f_arrdiv32_fs932_xor0 = f_arrdiv32_mux2to1871_xor0 ^ b[4];
  assign f_arrdiv32_fs932_not0 = ~f_arrdiv32_mux2to1871_xor0;
  assign f_arrdiv32_fs932_and0 = f_arrdiv32_fs932_not0 & b[4];
  assign f_arrdiv32_fs932_xor1 = f_arrdiv32_fs931_or0 ^ f_arrdiv32_fs932_xor0;
  assign f_arrdiv32_fs932_not1 = ~f_arrdiv32_fs932_xor0;
  assign f_arrdiv32_fs932_and1 = f_arrdiv32_fs932_not1 & f_arrdiv32_fs931_or0;
  assign f_arrdiv32_fs932_or0 = f_arrdiv32_fs932_and1 | f_arrdiv32_fs932_and0;
  assign f_arrdiv32_fs933_xor0 = f_arrdiv32_mux2to1872_xor0 ^ b[5];
  assign f_arrdiv32_fs933_not0 = ~f_arrdiv32_mux2to1872_xor0;
  assign f_arrdiv32_fs933_and0 = f_arrdiv32_fs933_not0 & b[5];
  assign f_arrdiv32_fs933_xor1 = f_arrdiv32_fs932_or0 ^ f_arrdiv32_fs933_xor0;
  assign f_arrdiv32_fs933_not1 = ~f_arrdiv32_fs933_xor0;
  assign f_arrdiv32_fs933_and1 = f_arrdiv32_fs933_not1 & f_arrdiv32_fs932_or0;
  assign f_arrdiv32_fs933_or0 = f_arrdiv32_fs933_and1 | f_arrdiv32_fs933_and0;
  assign f_arrdiv32_fs934_xor0 = f_arrdiv32_mux2to1873_xor0 ^ b[6];
  assign f_arrdiv32_fs934_not0 = ~f_arrdiv32_mux2to1873_xor0;
  assign f_arrdiv32_fs934_and0 = f_arrdiv32_fs934_not0 & b[6];
  assign f_arrdiv32_fs934_xor1 = f_arrdiv32_fs933_or0 ^ f_arrdiv32_fs934_xor0;
  assign f_arrdiv32_fs934_not1 = ~f_arrdiv32_fs934_xor0;
  assign f_arrdiv32_fs934_and1 = f_arrdiv32_fs934_not1 & f_arrdiv32_fs933_or0;
  assign f_arrdiv32_fs934_or0 = f_arrdiv32_fs934_and1 | f_arrdiv32_fs934_and0;
  assign f_arrdiv32_fs935_xor0 = f_arrdiv32_mux2to1874_xor0 ^ b[7];
  assign f_arrdiv32_fs935_not0 = ~f_arrdiv32_mux2to1874_xor0;
  assign f_arrdiv32_fs935_and0 = f_arrdiv32_fs935_not0 & b[7];
  assign f_arrdiv32_fs935_xor1 = f_arrdiv32_fs934_or0 ^ f_arrdiv32_fs935_xor0;
  assign f_arrdiv32_fs935_not1 = ~f_arrdiv32_fs935_xor0;
  assign f_arrdiv32_fs935_and1 = f_arrdiv32_fs935_not1 & f_arrdiv32_fs934_or0;
  assign f_arrdiv32_fs935_or0 = f_arrdiv32_fs935_and1 | f_arrdiv32_fs935_and0;
  assign f_arrdiv32_fs936_xor0 = f_arrdiv32_mux2to1875_xor0 ^ b[8];
  assign f_arrdiv32_fs936_not0 = ~f_arrdiv32_mux2to1875_xor0;
  assign f_arrdiv32_fs936_and0 = f_arrdiv32_fs936_not0 & b[8];
  assign f_arrdiv32_fs936_xor1 = f_arrdiv32_fs935_or0 ^ f_arrdiv32_fs936_xor0;
  assign f_arrdiv32_fs936_not1 = ~f_arrdiv32_fs936_xor0;
  assign f_arrdiv32_fs936_and1 = f_arrdiv32_fs936_not1 & f_arrdiv32_fs935_or0;
  assign f_arrdiv32_fs936_or0 = f_arrdiv32_fs936_and1 | f_arrdiv32_fs936_and0;
  assign f_arrdiv32_fs937_xor0 = f_arrdiv32_mux2to1876_xor0 ^ b[9];
  assign f_arrdiv32_fs937_not0 = ~f_arrdiv32_mux2to1876_xor0;
  assign f_arrdiv32_fs937_and0 = f_arrdiv32_fs937_not0 & b[9];
  assign f_arrdiv32_fs937_xor1 = f_arrdiv32_fs936_or0 ^ f_arrdiv32_fs937_xor0;
  assign f_arrdiv32_fs937_not1 = ~f_arrdiv32_fs937_xor0;
  assign f_arrdiv32_fs937_and1 = f_arrdiv32_fs937_not1 & f_arrdiv32_fs936_or0;
  assign f_arrdiv32_fs937_or0 = f_arrdiv32_fs937_and1 | f_arrdiv32_fs937_and0;
  assign f_arrdiv32_fs938_xor0 = f_arrdiv32_mux2to1877_xor0 ^ b[10];
  assign f_arrdiv32_fs938_not0 = ~f_arrdiv32_mux2to1877_xor0;
  assign f_arrdiv32_fs938_and0 = f_arrdiv32_fs938_not0 & b[10];
  assign f_arrdiv32_fs938_xor1 = f_arrdiv32_fs937_or0 ^ f_arrdiv32_fs938_xor0;
  assign f_arrdiv32_fs938_not1 = ~f_arrdiv32_fs938_xor0;
  assign f_arrdiv32_fs938_and1 = f_arrdiv32_fs938_not1 & f_arrdiv32_fs937_or0;
  assign f_arrdiv32_fs938_or0 = f_arrdiv32_fs938_and1 | f_arrdiv32_fs938_and0;
  assign f_arrdiv32_fs939_xor0 = f_arrdiv32_mux2to1878_xor0 ^ b[11];
  assign f_arrdiv32_fs939_not0 = ~f_arrdiv32_mux2to1878_xor0;
  assign f_arrdiv32_fs939_and0 = f_arrdiv32_fs939_not0 & b[11];
  assign f_arrdiv32_fs939_xor1 = f_arrdiv32_fs938_or0 ^ f_arrdiv32_fs939_xor0;
  assign f_arrdiv32_fs939_not1 = ~f_arrdiv32_fs939_xor0;
  assign f_arrdiv32_fs939_and1 = f_arrdiv32_fs939_not1 & f_arrdiv32_fs938_or0;
  assign f_arrdiv32_fs939_or0 = f_arrdiv32_fs939_and1 | f_arrdiv32_fs939_and0;
  assign f_arrdiv32_fs940_xor0 = f_arrdiv32_mux2to1879_xor0 ^ b[12];
  assign f_arrdiv32_fs940_not0 = ~f_arrdiv32_mux2to1879_xor0;
  assign f_arrdiv32_fs940_and0 = f_arrdiv32_fs940_not0 & b[12];
  assign f_arrdiv32_fs940_xor1 = f_arrdiv32_fs939_or0 ^ f_arrdiv32_fs940_xor0;
  assign f_arrdiv32_fs940_not1 = ~f_arrdiv32_fs940_xor0;
  assign f_arrdiv32_fs940_and1 = f_arrdiv32_fs940_not1 & f_arrdiv32_fs939_or0;
  assign f_arrdiv32_fs940_or0 = f_arrdiv32_fs940_and1 | f_arrdiv32_fs940_and0;
  assign f_arrdiv32_fs941_xor0 = f_arrdiv32_mux2to1880_xor0 ^ b[13];
  assign f_arrdiv32_fs941_not0 = ~f_arrdiv32_mux2to1880_xor0;
  assign f_arrdiv32_fs941_and0 = f_arrdiv32_fs941_not0 & b[13];
  assign f_arrdiv32_fs941_xor1 = f_arrdiv32_fs940_or0 ^ f_arrdiv32_fs941_xor0;
  assign f_arrdiv32_fs941_not1 = ~f_arrdiv32_fs941_xor0;
  assign f_arrdiv32_fs941_and1 = f_arrdiv32_fs941_not1 & f_arrdiv32_fs940_or0;
  assign f_arrdiv32_fs941_or0 = f_arrdiv32_fs941_and1 | f_arrdiv32_fs941_and0;
  assign f_arrdiv32_fs942_xor0 = f_arrdiv32_mux2to1881_xor0 ^ b[14];
  assign f_arrdiv32_fs942_not0 = ~f_arrdiv32_mux2to1881_xor0;
  assign f_arrdiv32_fs942_and0 = f_arrdiv32_fs942_not0 & b[14];
  assign f_arrdiv32_fs942_xor1 = f_arrdiv32_fs941_or0 ^ f_arrdiv32_fs942_xor0;
  assign f_arrdiv32_fs942_not1 = ~f_arrdiv32_fs942_xor0;
  assign f_arrdiv32_fs942_and1 = f_arrdiv32_fs942_not1 & f_arrdiv32_fs941_or0;
  assign f_arrdiv32_fs942_or0 = f_arrdiv32_fs942_and1 | f_arrdiv32_fs942_and0;
  assign f_arrdiv32_fs943_xor0 = f_arrdiv32_mux2to1882_xor0 ^ b[15];
  assign f_arrdiv32_fs943_not0 = ~f_arrdiv32_mux2to1882_xor0;
  assign f_arrdiv32_fs943_and0 = f_arrdiv32_fs943_not0 & b[15];
  assign f_arrdiv32_fs943_xor1 = f_arrdiv32_fs942_or0 ^ f_arrdiv32_fs943_xor0;
  assign f_arrdiv32_fs943_not1 = ~f_arrdiv32_fs943_xor0;
  assign f_arrdiv32_fs943_and1 = f_arrdiv32_fs943_not1 & f_arrdiv32_fs942_or0;
  assign f_arrdiv32_fs943_or0 = f_arrdiv32_fs943_and1 | f_arrdiv32_fs943_and0;
  assign f_arrdiv32_fs944_xor0 = f_arrdiv32_mux2to1883_xor0 ^ b[16];
  assign f_arrdiv32_fs944_not0 = ~f_arrdiv32_mux2to1883_xor0;
  assign f_arrdiv32_fs944_and0 = f_arrdiv32_fs944_not0 & b[16];
  assign f_arrdiv32_fs944_xor1 = f_arrdiv32_fs943_or0 ^ f_arrdiv32_fs944_xor0;
  assign f_arrdiv32_fs944_not1 = ~f_arrdiv32_fs944_xor0;
  assign f_arrdiv32_fs944_and1 = f_arrdiv32_fs944_not1 & f_arrdiv32_fs943_or0;
  assign f_arrdiv32_fs944_or0 = f_arrdiv32_fs944_and1 | f_arrdiv32_fs944_and0;
  assign f_arrdiv32_fs945_xor0 = f_arrdiv32_mux2to1884_xor0 ^ b[17];
  assign f_arrdiv32_fs945_not0 = ~f_arrdiv32_mux2to1884_xor0;
  assign f_arrdiv32_fs945_and0 = f_arrdiv32_fs945_not0 & b[17];
  assign f_arrdiv32_fs945_xor1 = f_arrdiv32_fs944_or0 ^ f_arrdiv32_fs945_xor0;
  assign f_arrdiv32_fs945_not1 = ~f_arrdiv32_fs945_xor0;
  assign f_arrdiv32_fs945_and1 = f_arrdiv32_fs945_not1 & f_arrdiv32_fs944_or0;
  assign f_arrdiv32_fs945_or0 = f_arrdiv32_fs945_and1 | f_arrdiv32_fs945_and0;
  assign f_arrdiv32_fs946_xor0 = f_arrdiv32_mux2to1885_xor0 ^ b[18];
  assign f_arrdiv32_fs946_not0 = ~f_arrdiv32_mux2to1885_xor0;
  assign f_arrdiv32_fs946_and0 = f_arrdiv32_fs946_not0 & b[18];
  assign f_arrdiv32_fs946_xor1 = f_arrdiv32_fs945_or0 ^ f_arrdiv32_fs946_xor0;
  assign f_arrdiv32_fs946_not1 = ~f_arrdiv32_fs946_xor0;
  assign f_arrdiv32_fs946_and1 = f_arrdiv32_fs946_not1 & f_arrdiv32_fs945_or0;
  assign f_arrdiv32_fs946_or0 = f_arrdiv32_fs946_and1 | f_arrdiv32_fs946_and0;
  assign f_arrdiv32_fs947_xor0 = f_arrdiv32_mux2to1886_xor0 ^ b[19];
  assign f_arrdiv32_fs947_not0 = ~f_arrdiv32_mux2to1886_xor0;
  assign f_arrdiv32_fs947_and0 = f_arrdiv32_fs947_not0 & b[19];
  assign f_arrdiv32_fs947_xor1 = f_arrdiv32_fs946_or0 ^ f_arrdiv32_fs947_xor0;
  assign f_arrdiv32_fs947_not1 = ~f_arrdiv32_fs947_xor0;
  assign f_arrdiv32_fs947_and1 = f_arrdiv32_fs947_not1 & f_arrdiv32_fs946_or0;
  assign f_arrdiv32_fs947_or0 = f_arrdiv32_fs947_and1 | f_arrdiv32_fs947_and0;
  assign f_arrdiv32_fs948_xor0 = f_arrdiv32_mux2to1887_xor0 ^ b[20];
  assign f_arrdiv32_fs948_not0 = ~f_arrdiv32_mux2to1887_xor0;
  assign f_arrdiv32_fs948_and0 = f_arrdiv32_fs948_not0 & b[20];
  assign f_arrdiv32_fs948_xor1 = f_arrdiv32_fs947_or0 ^ f_arrdiv32_fs948_xor0;
  assign f_arrdiv32_fs948_not1 = ~f_arrdiv32_fs948_xor0;
  assign f_arrdiv32_fs948_and1 = f_arrdiv32_fs948_not1 & f_arrdiv32_fs947_or0;
  assign f_arrdiv32_fs948_or0 = f_arrdiv32_fs948_and1 | f_arrdiv32_fs948_and0;
  assign f_arrdiv32_fs949_xor0 = f_arrdiv32_mux2to1888_xor0 ^ b[21];
  assign f_arrdiv32_fs949_not0 = ~f_arrdiv32_mux2to1888_xor0;
  assign f_arrdiv32_fs949_and0 = f_arrdiv32_fs949_not0 & b[21];
  assign f_arrdiv32_fs949_xor1 = f_arrdiv32_fs948_or0 ^ f_arrdiv32_fs949_xor0;
  assign f_arrdiv32_fs949_not1 = ~f_arrdiv32_fs949_xor0;
  assign f_arrdiv32_fs949_and1 = f_arrdiv32_fs949_not1 & f_arrdiv32_fs948_or0;
  assign f_arrdiv32_fs949_or0 = f_arrdiv32_fs949_and1 | f_arrdiv32_fs949_and0;
  assign f_arrdiv32_fs950_xor0 = f_arrdiv32_mux2to1889_xor0 ^ b[22];
  assign f_arrdiv32_fs950_not0 = ~f_arrdiv32_mux2to1889_xor0;
  assign f_arrdiv32_fs950_and0 = f_arrdiv32_fs950_not0 & b[22];
  assign f_arrdiv32_fs950_xor1 = f_arrdiv32_fs949_or0 ^ f_arrdiv32_fs950_xor0;
  assign f_arrdiv32_fs950_not1 = ~f_arrdiv32_fs950_xor0;
  assign f_arrdiv32_fs950_and1 = f_arrdiv32_fs950_not1 & f_arrdiv32_fs949_or0;
  assign f_arrdiv32_fs950_or0 = f_arrdiv32_fs950_and1 | f_arrdiv32_fs950_and0;
  assign f_arrdiv32_fs951_xor0 = f_arrdiv32_mux2to1890_xor0 ^ b[23];
  assign f_arrdiv32_fs951_not0 = ~f_arrdiv32_mux2to1890_xor0;
  assign f_arrdiv32_fs951_and0 = f_arrdiv32_fs951_not0 & b[23];
  assign f_arrdiv32_fs951_xor1 = f_arrdiv32_fs950_or0 ^ f_arrdiv32_fs951_xor0;
  assign f_arrdiv32_fs951_not1 = ~f_arrdiv32_fs951_xor0;
  assign f_arrdiv32_fs951_and1 = f_arrdiv32_fs951_not1 & f_arrdiv32_fs950_or0;
  assign f_arrdiv32_fs951_or0 = f_arrdiv32_fs951_and1 | f_arrdiv32_fs951_and0;
  assign f_arrdiv32_fs952_xor0 = f_arrdiv32_mux2to1891_xor0 ^ b[24];
  assign f_arrdiv32_fs952_not0 = ~f_arrdiv32_mux2to1891_xor0;
  assign f_arrdiv32_fs952_and0 = f_arrdiv32_fs952_not0 & b[24];
  assign f_arrdiv32_fs952_xor1 = f_arrdiv32_fs951_or0 ^ f_arrdiv32_fs952_xor0;
  assign f_arrdiv32_fs952_not1 = ~f_arrdiv32_fs952_xor0;
  assign f_arrdiv32_fs952_and1 = f_arrdiv32_fs952_not1 & f_arrdiv32_fs951_or0;
  assign f_arrdiv32_fs952_or0 = f_arrdiv32_fs952_and1 | f_arrdiv32_fs952_and0;
  assign f_arrdiv32_fs953_xor0 = f_arrdiv32_mux2to1892_xor0 ^ b[25];
  assign f_arrdiv32_fs953_not0 = ~f_arrdiv32_mux2to1892_xor0;
  assign f_arrdiv32_fs953_and0 = f_arrdiv32_fs953_not0 & b[25];
  assign f_arrdiv32_fs953_xor1 = f_arrdiv32_fs952_or0 ^ f_arrdiv32_fs953_xor0;
  assign f_arrdiv32_fs953_not1 = ~f_arrdiv32_fs953_xor0;
  assign f_arrdiv32_fs953_and1 = f_arrdiv32_fs953_not1 & f_arrdiv32_fs952_or0;
  assign f_arrdiv32_fs953_or0 = f_arrdiv32_fs953_and1 | f_arrdiv32_fs953_and0;
  assign f_arrdiv32_fs954_xor0 = f_arrdiv32_mux2to1893_xor0 ^ b[26];
  assign f_arrdiv32_fs954_not0 = ~f_arrdiv32_mux2to1893_xor0;
  assign f_arrdiv32_fs954_and0 = f_arrdiv32_fs954_not0 & b[26];
  assign f_arrdiv32_fs954_xor1 = f_arrdiv32_fs953_or0 ^ f_arrdiv32_fs954_xor0;
  assign f_arrdiv32_fs954_not1 = ~f_arrdiv32_fs954_xor0;
  assign f_arrdiv32_fs954_and1 = f_arrdiv32_fs954_not1 & f_arrdiv32_fs953_or0;
  assign f_arrdiv32_fs954_or0 = f_arrdiv32_fs954_and1 | f_arrdiv32_fs954_and0;
  assign f_arrdiv32_fs955_xor0 = f_arrdiv32_mux2to1894_xor0 ^ b[27];
  assign f_arrdiv32_fs955_not0 = ~f_arrdiv32_mux2to1894_xor0;
  assign f_arrdiv32_fs955_and0 = f_arrdiv32_fs955_not0 & b[27];
  assign f_arrdiv32_fs955_xor1 = f_arrdiv32_fs954_or0 ^ f_arrdiv32_fs955_xor0;
  assign f_arrdiv32_fs955_not1 = ~f_arrdiv32_fs955_xor0;
  assign f_arrdiv32_fs955_and1 = f_arrdiv32_fs955_not1 & f_arrdiv32_fs954_or0;
  assign f_arrdiv32_fs955_or0 = f_arrdiv32_fs955_and1 | f_arrdiv32_fs955_and0;
  assign f_arrdiv32_fs956_xor0 = f_arrdiv32_mux2to1895_xor0 ^ b[28];
  assign f_arrdiv32_fs956_not0 = ~f_arrdiv32_mux2to1895_xor0;
  assign f_arrdiv32_fs956_and0 = f_arrdiv32_fs956_not0 & b[28];
  assign f_arrdiv32_fs956_xor1 = f_arrdiv32_fs955_or0 ^ f_arrdiv32_fs956_xor0;
  assign f_arrdiv32_fs956_not1 = ~f_arrdiv32_fs956_xor0;
  assign f_arrdiv32_fs956_and1 = f_arrdiv32_fs956_not1 & f_arrdiv32_fs955_or0;
  assign f_arrdiv32_fs956_or0 = f_arrdiv32_fs956_and1 | f_arrdiv32_fs956_and0;
  assign f_arrdiv32_fs957_xor0 = f_arrdiv32_mux2to1896_xor0 ^ b[29];
  assign f_arrdiv32_fs957_not0 = ~f_arrdiv32_mux2to1896_xor0;
  assign f_arrdiv32_fs957_and0 = f_arrdiv32_fs957_not0 & b[29];
  assign f_arrdiv32_fs957_xor1 = f_arrdiv32_fs956_or0 ^ f_arrdiv32_fs957_xor0;
  assign f_arrdiv32_fs957_not1 = ~f_arrdiv32_fs957_xor0;
  assign f_arrdiv32_fs957_and1 = f_arrdiv32_fs957_not1 & f_arrdiv32_fs956_or0;
  assign f_arrdiv32_fs957_or0 = f_arrdiv32_fs957_and1 | f_arrdiv32_fs957_and0;
  assign f_arrdiv32_fs958_xor0 = f_arrdiv32_mux2to1897_xor0 ^ b[30];
  assign f_arrdiv32_fs958_not0 = ~f_arrdiv32_mux2to1897_xor0;
  assign f_arrdiv32_fs958_and0 = f_arrdiv32_fs958_not0 & b[30];
  assign f_arrdiv32_fs958_xor1 = f_arrdiv32_fs957_or0 ^ f_arrdiv32_fs958_xor0;
  assign f_arrdiv32_fs958_not1 = ~f_arrdiv32_fs958_xor0;
  assign f_arrdiv32_fs958_and1 = f_arrdiv32_fs958_not1 & f_arrdiv32_fs957_or0;
  assign f_arrdiv32_fs958_or0 = f_arrdiv32_fs958_and1 | f_arrdiv32_fs958_and0;
  assign f_arrdiv32_fs959_xor0 = f_arrdiv32_mux2to1898_xor0 ^ b[31];
  assign f_arrdiv32_fs959_not0 = ~f_arrdiv32_mux2to1898_xor0;
  assign f_arrdiv32_fs959_and0 = f_arrdiv32_fs959_not0 & b[31];
  assign f_arrdiv32_fs959_xor1 = f_arrdiv32_fs958_or0 ^ f_arrdiv32_fs959_xor0;
  assign f_arrdiv32_fs959_not1 = ~f_arrdiv32_fs959_xor0;
  assign f_arrdiv32_fs959_and1 = f_arrdiv32_fs959_not1 & f_arrdiv32_fs958_or0;
  assign f_arrdiv32_fs959_or0 = f_arrdiv32_fs959_and1 | f_arrdiv32_fs959_and0;
  assign f_arrdiv32_mux2to1899_and0 = a[2] & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1899_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1899_and1 = f_arrdiv32_fs928_xor0 & f_arrdiv32_mux2to1899_not0;
  assign f_arrdiv32_mux2to1899_xor0 = f_arrdiv32_mux2to1899_and0 ^ f_arrdiv32_mux2to1899_and1;
  assign f_arrdiv32_mux2to1900_and0 = f_arrdiv32_mux2to1868_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1900_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1900_and1 = f_arrdiv32_fs929_xor1 & f_arrdiv32_mux2to1900_not0;
  assign f_arrdiv32_mux2to1900_xor0 = f_arrdiv32_mux2to1900_and0 ^ f_arrdiv32_mux2to1900_and1;
  assign f_arrdiv32_mux2to1901_and0 = f_arrdiv32_mux2to1869_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1901_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1901_and1 = f_arrdiv32_fs930_xor1 & f_arrdiv32_mux2to1901_not0;
  assign f_arrdiv32_mux2to1901_xor0 = f_arrdiv32_mux2to1901_and0 ^ f_arrdiv32_mux2to1901_and1;
  assign f_arrdiv32_mux2to1902_and0 = f_arrdiv32_mux2to1870_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1902_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1902_and1 = f_arrdiv32_fs931_xor1 & f_arrdiv32_mux2to1902_not0;
  assign f_arrdiv32_mux2to1902_xor0 = f_arrdiv32_mux2to1902_and0 ^ f_arrdiv32_mux2to1902_and1;
  assign f_arrdiv32_mux2to1903_and0 = f_arrdiv32_mux2to1871_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1903_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1903_and1 = f_arrdiv32_fs932_xor1 & f_arrdiv32_mux2to1903_not0;
  assign f_arrdiv32_mux2to1903_xor0 = f_arrdiv32_mux2to1903_and0 ^ f_arrdiv32_mux2to1903_and1;
  assign f_arrdiv32_mux2to1904_and0 = f_arrdiv32_mux2to1872_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1904_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1904_and1 = f_arrdiv32_fs933_xor1 & f_arrdiv32_mux2to1904_not0;
  assign f_arrdiv32_mux2to1904_xor0 = f_arrdiv32_mux2to1904_and0 ^ f_arrdiv32_mux2to1904_and1;
  assign f_arrdiv32_mux2to1905_and0 = f_arrdiv32_mux2to1873_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1905_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1905_and1 = f_arrdiv32_fs934_xor1 & f_arrdiv32_mux2to1905_not0;
  assign f_arrdiv32_mux2to1905_xor0 = f_arrdiv32_mux2to1905_and0 ^ f_arrdiv32_mux2to1905_and1;
  assign f_arrdiv32_mux2to1906_and0 = f_arrdiv32_mux2to1874_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1906_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1906_and1 = f_arrdiv32_fs935_xor1 & f_arrdiv32_mux2to1906_not0;
  assign f_arrdiv32_mux2to1906_xor0 = f_arrdiv32_mux2to1906_and0 ^ f_arrdiv32_mux2to1906_and1;
  assign f_arrdiv32_mux2to1907_and0 = f_arrdiv32_mux2to1875_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1907_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1907_and1 = f_arrdiv32_fs936_xor1 & f_arrdiv32_mux2to1907_not0;
  assign f_arrdiv32_mux2to1907_xor0 = f_arrdiv32_mux2to1907_and0 ^ f_arrdiv32_mux2to1907_and1;
  assign f_arrdiv32_mux2to1908_and0 = f_arrdiv32_mux2to1876_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1908_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1908_and1 = f_arrdiv32_fs937_xor1 & f_arrdiv32_mux2to1908_not0;
  assign f_arrdiv32_mux2to1908_xor0 = f_arrdiv32_mux2to1908_and0 ^ f_arrdiv32_mux2to1908_and1;
  assign f_arrdiv32_mux2to1909_and0 = f_arrdiv32_mux2to1877_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1909_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1909_and1 = f_arrdiv32_fs938_xor1 & f_arrdiv32_mux2to1909_not0;
  assign f_arrdiv32_mux2to1909_xor0 = f_arrdiv32_mux2to1909_and0 ^ f_arrdiv32_mux2to1909_and1;
  assign f_arrdiv32_mux2to1910_and0 = f_arrdiv32_mux2to1878_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1910_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1910_and1 = f_arrdiv32_fs939_xor1 & f_arrdiv32_mux2to1910_not0;
  assign f_arrdiv32_mux2to1910_xor0 = f_arrdiv32_mux2to1910_and0 ^ f_arrdiv32_mux2to1910_and1;
  assign f_arrdiv32_mux2to1911_and0 = f_arrdiv32_mux2to1879_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1911_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1911_and1 = f_arrdiv32_fs940_xor1 & f_arrdiv32_mux2to1911_not0;
  assign f_arrdiv32_mux2to1911_xor0 = f_arrdiv32_mux2to1911_and0 ^ f_arrdiv32_mux2to1911_and1;
  assign f_arrdiv32_mux2to1912_and0 = f_arrdiv32_mux2to1880_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1912_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1912_and1 = f_arrdiv32_fs941_xor1 & f_arrdiv32_mux2to1912_not0;
  assign f_arrdiv32_mux2to1912_xor0 = f_arrdiv32_mux2to1912_and0 ^ f_arrdiv32_mux2to1912_and1;
  assign f_arrdiv32_mux2to1913_and0 = f_arrdiv32_mux2to1881_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1913_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1913_and1 = f_arrdiv32_fs942_xor1 & f_arrdiv32_mux2to1913_not0;
  assign f_arrdiv32_mux2to1913_xor0 = f_arrdiv32_mux2to1913_and0 ^ f_arrdiv32_mux2to1913_and1;
  assign f_arrdiv32_mux2to1914_and0 = f_arrdiv32_mux2to1882_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1914_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1914_and1 = f_arrdiv32_fs943_xor1 & f_arrdiv32_mux2to1914_not0;
  assign f_arrdiv32_mux2to1914_xor0 = f_arrdiv32_mux2to1914_and0 ^ f_arrdiv32_mux2to1914_and1;
  assign f_arrdiv32_mux2to1915_and0 = f_arrdiv32_mux2to1883_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1915_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1915_and1 = f_arrdiv32_fs944_xor1 & f_arrdiv32_mux2to1915_not0;
  assign f_arrdiv32_mux2to1915_xor0 = f_arrdiv32_mux2to1915_and0 ^ f_arrdiv32_mux2to1915_and1;
  assign f_arrdiv32_mux2to1916_and0 = f_arrdiv32_mux2to1884_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1916_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1916_and1 = f_arrdiv32_fs945_xor1 & f_arrdiv32_mux2to1916_not0;
  assign f_arrdiv32_mux2to1916_xor0 = f_arrdiv32_mux2to1916_and0 ^ f_arrdiv32_mux2to1916_and1;
  assign f_arrdiv32_mux2to1917_and0 = f_arrdiv32_mux2to1885_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1917_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1917_and1 = f_arrdiv32_fs946_xor1 & f_arrdiv32_mux2to1917_not0;
  assign f_arrdiv32_mux2to1917_xor0 = f_arrdiv32_mux2to1917_and0 ^ f_arrdiv32_mux2to1917_and1;
  assign f_arrdiv32_mux2to1918_and0 = f_arrdiv32_mux2to1886_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1918_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1918_and1 = f_arrdiv32_fs947_xor1 & f_arrdiv32_mux2to1918_not0;
  assign f_arrdiv32_mux2to1918_xor0 = f_arrdiv32_mux2to1918_and0 ^ f_arrdiv32_mux2to1918_and1;
  assign f_arrdiv32_mux2to1919_and0 = f_arrdiv32_mux2to1887_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1919_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1919_and1 = f_arrdiv32_fs948_xor1 & f_arrdiv32_mux2to1919_not0;
  assign f_arrdiv32_mux2to1919_xor0 = f_arrdiv32_mux2to1919_and0 ^ f_arrdiv32_mux2to1919_and1;
  assign f_arrdiv32_mux2to1920_and0 = f_arrdiv32_mux2to1888_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1920_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1920_and1 = f_arrdiv32_fs949_xor1 & f_arrdiv32_mux2to1920_not0;
  assign f_arrdiv32_mux2to1920_xor0 = f_arrdiv32_mux2to1920_and0 ^ f_arrdiv32_mux2to1920_and1;
  assign f_arrdiv32_mux2to1921_and0 = f_arrdiv32_mux2to1889_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1921_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1921_and1 = f_arrdiv32_fs950_xor1 & f_arrdiv32_mux2to1921_not0;
  assign f_arrdiv32_mux2to1921_xor0 = f_arrdiv32_mux2to1921_and0 ^ f_arrdiv32_mux2to1921_and1;
  assign f_arrdiv32_mux2to1922_and0 = f_arrdiv32_mux2to1890_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1922_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1922_and1 = f_arrdiv32_fs951_xor1 & f_arrdiv32_mux2to1922_not0;
  assign f_arrdiv32_mux2to1922_xor0 = f_arrdiv32_mux2to1922_and0 ^ f_arrdiv32_mux2to1922_and1;
  assign f_arrdiv32_mux2to1923_and0 = f_arrdiv32_mux2to1891_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1923_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1923_and1 = f_arrdiv32_fs952_xor1 & f_arrdiv32_mux2to1923_not0;
  assign f_arrdiv32_mux2to1923_xor0 = f_arrdiv32_mux2to1923_and0 ^ f_arrdiv32_mux2to1923_and1;
  assign f_arrdiv32_mux2to1924_and0 = f_arrdiv32_mux2to1892_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1924_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1924_and1 = f_arrdiv32_fs953_xor1 & f_arrdiv32_mux2to1924_not0;
  assign f_arrdiv32_mux2to1924_xor0 = f_arrdiv32_mux2to1924_and0 ^ f_arrdiv32_mux2to1924_and1;
  assign f_arrdiv32_mux2to1925_and0 = f_arrdiv32_mux2to1893_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1925_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1925_and1 = f_arrdiv32_fs954_xor1 & f_arrdiv32_mux2to1925_not0;
  assign f_arrdiv32_mux2to1925_xor0 = f_arrdiv32_mux2to1925_and0 ^ f_arrdiv32_mux2to1925_and1;
  assign f_arrdiv32_mux2to1926_and0 = f_arrdiv32_mux2to1894_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1926_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1926_and1 = f_arrdiv32_fs955_xor1 & f_arrdiv32_mux2to1926_not0;
  assign f_arrdiv32_mux2to1926_xor0 = f_arrdiv32_mux2to1926_and0 ^ f_arrdiv32_mux2to1926_and1;
  assign f_arrdiv32_mux2to1927_and0 = f_arrdiv32_mux2to1895_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1927_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1927_and1 = f_arrdiv32_fs956_xor1 & f_arrdiv32_mux2to1927_not0;
  assign f_arrdiv32_mux2to1927_xor0 = f_arrdiv32_mux2to1927_and0 ^ f_arrdiv32_mux2to1927_and1;
  assign f_arrdiv32_mux2to1928_and0 = f_arrdiv32_mux2to1896_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1928_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1928_and1 = f_arrdiv32_fs957_xor1 & f_arrdiv32_mux2to1928_not0;
  assign f_arrdiv32_mux2to1928_xor0 = f_arrdiv32_mux2to1928_and0 ^ f_arrdiv32_mux2to1928_and1;
  assign f_arrdiv32_mux2to1929_and0 = f_arrdiv32_mux2to1897_xor0 & f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1929_not0 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_mux2to1929_and1 = f_arrdiv32_fs958_xor1 & f_arrdiv32_mux2to1929_not0;
  assign f_arrdiv32_mux2to1929_xor0 = f_arrdiv32_mux2to1929_and0 ^ f_arrdiv32_mux2to1929_and1;
  assign f_arrdiv32_not29 = ~f_arrdiv32_fs959_or0;
  assign f_arrdiv32_fs960_xor0 = a[1] ^ b[0];
  assign f_arrdiv32_fs960_not0 = ~a[1];
  assign f_arrdiv32_fs960_and0 = f_arrdiv32_fs960_not0 & b[0];
  assign f_arrdiv32_fs960_not1 = ~f_arrdiv32_fs960_xor0;
  assign f_arrdiv32_fs961_xor0 = f_arrdiv32_mux2to1899_xor0 ^ b[1];
  assign f_arrdiv32_fs961_not0 = ~f_arrdiv32_mux2to1899_xor0;
  assign f_arrdiv32_fs961_and0 = f_arrdiv32_fs961_not0 & b[1];
  assign f_arrdiv32_fs961_xor1 = f_arrdiv32_fs960_and0 ^ f_arrdiv32_fs961_xor0;
  assign f_arrdiv32_fs961_not1 = ~f_arrdiv32_fs961_xor0;
  assign f_arrdiv32_fs961_and1 = f_arrdiv32_fs961_not1 & f_arrdiv32_fs960_and0;
  assign f_arrdiv32_fs961_or0 = f_arrdiv32_fs961_and1 | f_arrdiv32_fs961_and0;
  assign f_arrdiv32_fs962_xor0 = f_arrdiv32_mux2to1900_xor0 ^ b[2];
  assign f_arrdiv32_fs962_not0 = ~f_arrdiv32_mux2to1900_xor0;
  assign f_arrdiv32_fs962_and0 = f_arrdiv32_fs962_not0 & b[2];
  assign f_arrdiv32_fs962_xor1 = f_arrdiv32_fs961_or0 ^ f_arrdiv32_fs962_xor0;
  assign f_arrdiv32_fs962_not1 = ~f_arrdiv32_fs962_xor0;
  assign f_arrdiv32_fs962_and1 = f_arrdiv32_fs962_not1 & f_arrdiv32_fs961_or0;
  assign f_arrdiv32_fs962_or0 = f_arrdiv32_fs962_and1 | f_arrdiv32_fs962_and0;
  assign f_arrdiv32_fs963_xor0 = f_arrdiv32_mux2to1901_xor0 ^ b[3];
  assign f_arrdiv32_fs963_not0 = ~f_arrdiv32_mux2to1901_xor0;
  assign f_arrdiv32_fs963_and0 = f_arrdiv32_fs963_not0 & b[3];
  assign f_arrdiv32_fs963_xor1 = f_arrdiv32_fs962_or0 ^ f_arrdiv32_fs963_xor0;
  assign f_arrdiv32_fs963_not1 = ~f_arrdiv32_fs963_xor0;
  assign f_arrdiv32_fs963_and1 = f_arrdiv32_fs963_not1 & f_arrdiv32_fs962_or0;
  assign f_arrdiv32_fs963_or0 = f_arrdiv32_fs963_and1 | f_arrdiv32_fs963_and0;
  assign f_arrdiv32_fs964_xor0 = f_arrdiv32_mux2to1902_xor0 ^ b[4];
  assign f_arrdiv32_fs964_not0 = ~f_arrdiv32_mux2to1902_xor0;
  assign f_arrdiv32_fs964_and0 = f_arrdiv32_fs964_not0 & b[4];
  assign f_arrdiv32_fs964_xor1 = f_arrdiv32_fs963_or0 ^ f_arrdiv32_fs964_xor0;
  assign f_arrdiv32_fs964_not1 = ~f_arrdiv32_fs964_xor0;
  assign f_arrdiv32_fs964_and1 = f_arrdiv32_fs964_not1 & f_arrdiv32_fs963_or0;
  assign f_arrdiv32_fs964_or0 = f_arrdiv32_fs964_and1 | f_arrdiv32_fs964_and0;
  assign f_arrdiv32_fs965_xor0 = f_arrdiv32_mux2to1903_xor0 ^ b[5];
  assign f_arrdiv32_fs965_not0 = ~f_arrdiv32_mux2to1903_xor0;
  assign f_arrdiv32_fs965_and0 = f_arrdiv32_fs965_not0 & b[5];
  assign f_arrdiv32_fs965_xor1 = f_arrdiv32_fs964_or0 ^ f_arrdiv32_fs965_xor0;
  assign f_arrdiv32_fs965_not1 = ~f_arrdiv32_fs965_xor0;
  assign f_arrdiv32_fs965_and1 = f_arrdiv32_fs965_not1 & f_arrdiv32_fs964_or0;
  assign f_arrdiv32_fs965_or0 = f_arrdiv32_fs965_and1 | f_arrdiv32_fs965_and0;
  assign f_arrdiv32_fs966_xor0 = f_arrdiv32_mux2to1904_xor0 ^ b[6];
  assign f_arrdiv32_fs966_not0 = ~f_arrdiv32_mux2to1904_xor0;
  assign f_arrdiv32_fs966_and0 = f_arrdiv32_fs966_not0 & b[6];
  assign f_arrdiv32_fs966_xor1 = f_arrdiv32_fs965_or0 ^ f_arrdiv32_fs966_xor0;
  assign f_arrdiv32_fs966_not1 = ~f_arrdiv32_fs966_xor0;
  assign f_arrdiv32_fs966_and1 = f_arrdiv32_fs966_not1 & f_arrdiv32_fs965_or0;
  assign f_arrdiv32_fs966_or0 = f_arrdiv32_fs966_and1 | f_arrdiv32_fs966_and0;
  assign f_arrdiv32_fs967_xor0 = f_arrdiv32_mux2to1905_xor0 ^ b[7];
  assign f_arrdiv32_fs967_not0 = ~f_arrdiv32_mux2to1905_xor0;
  assign f_arrdiv32_fs967_and0 = f_arrdiv32_fs967_not0 & b[7];
  assign f_arrdiv32_fs967_xor1 = f_arrdiv32_fs966_or0 ^ f_arrdiv32_fs967_xor0;
  assign f_arrdiv32_fs967_not1 = ~f_arrdiv32_fs967_xor0;
  assign f_arrdiv32_fs967_and1 = f_arrdiv32_fs967_not1 & f_arrdiv32_fs966_or0;
  assign f_arrdiv32_fs967_or0 = f_arrdiv32_fs967_and1 | f_arrdiv32_fs967_and0;
  assign f_arrdiv32_fs968_xor0 = f_arrdiv32_mux2to1906_xor0 ^ b[8];
  assign f_arrdiv32_fs968_not0 = ~f_arrdiv32_mux2to1906_xor0;
  assign f_arrdiv32_fs968_and0 = f_arrdiv32_fs968_not0 & b[8];
  assign f_arrdiv32_fs968_xor1 = f_arrdiv32_fs967_or0 ^ f_arrdiv32_fs968_xor0;
  assign f_arrdiv32_fs968_not1 = ~f_arrdiv32_fs968_xor0;
  assign f_arrdiv32_fs968_and1 = f_arrdiv32_fs968_not1 & f_arrdiv32_fs967_or0;
  assign f_arrdiv32_fs968_or0 = f_arrdiv32_fs968_and1 | f_arrdiv32_fs968_and0;
  assign f_arrdiv32_fs969_xor0 = f_arrdiv32_mux2to1907_xor0 ^ b[9];
  assign f_arrdiv32_fs969_not0 = ~f_arrdiv32_mux2to1907_xor0;
  assign f_arrdiv32_fs969_and0 = f_arrdiv32_fs969_not0 & b[9];
  assign f_arrdiv32_fs969_xor1 = f_arrdiv32_fs968_or0 ^ f_arrdiv32_fs969_xor0;
  assign f_arrdiv32_fs969_not1 = ~f_arrdiv32_fs969_xor0;
  assign f_arrdiv32_fs969_and1 = f_arrdiv32_fs969_not1 & f_arrdiv32_fs968_or0;
  assign f_arrdiv32_fs969_or0 = f_arrdiv32_fs969_and1 | f_arrdiv32_fs969_and0;
  assign f_arrdiv32_fs970_xor0 = f_arrdiv32_mux2to1908_xor0 ^ b[10];
  assign f_arrdiv32_fs970_not0 = ~f_arrdiv32_mux2to1908_xor0;
  assign f_arrdiv32_fs970_and0 = f_arrdiv32_fs970_not0 & b[10];
  assign f_arrdiv32_fs970_xor1 = f_arrdiv32_fs969_or0 ^ f_arrdiv32_fs970_xor0;
  assign f_arrdiv32_fs970_not1 = ~f_arrdiv32_fs970_xor0;
  assign f_arrdiv32_fs970_and1 = f_arrdiv32_fs970_not1 & f_arrdiv32_fs969_or0;
  assign f_arrdiv32_fs970_or0 = f_arrdiv32_fs970_and1 | f_arrdiv32_fs970_and0;
  assign f_arrdiv32_fs971_xor0 = f_arrdiv32_mux2to1909_xor0 ^ b[11];
  assign f_arrdiv32_fs971_not0 = ~f_arrdiv32_mux2to1909_xor0;
  assign f_arrdiv32_fs971_and0 = f_arrdiv32_fs971_not0 & b[11];
  assign f_arrdiv32_fs971_xor1 = f_arrdiv32_fs970_or0 ^ f_arrdiv32_fs971_xor0;
  assign f_arrdiv32_fs971_not1 = ~f_arrdiv32_fs971_xor0;
  assign f_arrdiv32_fs971_and1 = f_arrdiv32_fs971_not1 & f_arrdiv32_fs970_or0;
  assign f_arrdiv32_fs971_or0 = f_arrdiv32_fs971_and1 | f_arrdiv32_fs971_and0;
  assign f_arrdiv32_fs972_xor0 = f_arrdiv32_mux2to1910_xor0 ^ b[12];
  assign f_arrdiv32_fs972_not0 = ~f_arrdiv32_mux2to1910_xor0;
  assign f_arrdiv32_fs972_and0 = f_arrdiv32_fs972_not0 & b[12];
  assign f_arrdiv32_fs972_xor1 = f_arrdiv32_fs971_or0 ^ f_arrdiv32_fs972_xor0;
  assign f_arrdiv32_fs972_not1 = ~f_arrdiv32_fs972_xor0;
  assign f_arrdiv32_fs972_and1 = f_arrdiv32_fs972_not1 & f_arrdiv32_fs971_or0;
  assign f_arrdiv32_fs972_or0 = f_arrdiv32_fs972_and1 | f_arrdiv32_fs972_and0;
  assign f_arrdiv32_fs973_xor0 = f_arrdiv32_mux2to1911_xor0 ^ b[13];
  assign f_arrdiv32_fs973_not0 = ~f_arrdiv32_mux2to1911_xor0;
  assign f_arrdiv32_fs973_and0 = f_arrdiv32_fs973_not0 & b[13];
  assign f_arrdiv32_fs973_xor1 = f_arrdiv32_fs972_or0 ^ f_arrdiv32_fs973_xor0;
  assign f_arrdiv32_fs973_not1 = ~f_arrdiv32_fs973_xor0;
  assign f_arrdiv32_fs973_and1 = f_arrdiv32_fs973_not1 & f_arrdiv32_fs972_or0;
  assign f_arrdiv32_fs973_or0 = f_arrdiv32_fs973_and1 | f_arrdiv32_fs973_and0;
  assign f_arrdiv32_fs974_xor0 = f_arrdiv32_mux2to1912_xor0 ^ b[14];
  assign f_arrdiv32_fs974_not0 = ~f_arrdiv32_mux2to1912_xor0;
  assign f_arrdiv32_fs974_and0 = f_arrdiv32_fs974_not0 & b[14];
  assign f_arrdiv32_fs974_xor1 = f_arrdiv32_fs973_or0 ^ f_arrdiv32_fs974_xor0;
  assign f_arrdiv32_fs974_not1 = ~f_arrdiv32_fs974_xor0;
  assign f_arrdiv32_fs974_and1 = f_arrdiv32_fs974_not1 & f_arrdiv32_fs973_or0;
  assign f_arrdiv32_fs974_or0 = f_arrdiv32_fs974_and1 | f_arrdiv32_fs974_and0;
  assign f_arrdiv32_fs975_xor0 = f_arrdiv32_mux2to1913_xor0 ^ b[15];
  assign f_arrdiv32_fs975_not0 = ~f_arrdiv32_mux2to1913_xor0;
  assign f_arrdiv32_fs975_and0 = f_arrdiv32_fs975_not0 & b[15];
  assign f_arrdiv32_fs975_xor1 = f_arrdiv32_fs974_or0 ^ f_arrdiv32_fs975_xor0;
  assign f_arrdiv32_fs975_not1 = ~f_arrdiv32_fs975_xor0;
  assign f_arrdiv32_fs975_and1 = f_arrdiv32_fs975_not1 & f_arrdiv32_fs974_or0;
  assign f_arrdiv32_fs975_or0 = f_arrdiv32_fs975_and1 | f_arrdiv32_fs975_and0;
  assign f_arrdiv32_fs976_xor0 = f_arrdiv32_mux2to1914_xor0 ^ b[16];
  assign f_arrdiv32_fs976_not0 = ~f_arrdiv32_mux2to1914_xor0;
  assign f_arrdiv32_fs976_and0 = f_arrdiv32_fs976_not0 & b[16];
  assign f_arrdiv32_fs976_xor1 = f_arrdiv32_fs975_or0 ^ f_arrdiv32_fs976_xor0;
  assign f_arrdiv32_fs976_not1 = ~f_arrdiv32_fs976_xor0;
  assign f_arrdiv32_fs976_and1 = f_arrdiv32_fs976_not1 & f_arrdiv32_fs975_or0;
  assign f_arrdiv32_fs976_or0 = f_arrdiv32_fs976_and1 | f_arrdiv32_fs976_and0;
  assign f_arrdiv32_fs977_xor0 = f_arrdiv32_mux2to1915_xor0 ^ b[17];
  assign f_arrdiv32_fs977_not0 = ~f_arrdiv32_mux2to1915_xor0;
  assign f_arrdiv32_fs977_and0 = f_arrdiv32_fs977_not0 & b[17];
  assign f_arrdiv32_fs977_xor1 = f_arrdiv32_fs976_or0 ^ f_arrdiv32_fs977_xor0;
  assign f_arrdiv32_fs977_not1 = ~f_arrdiv32_fs977_xor0;
  assign f_arrdiv32_fs977_and1 = f_arrdiv32_fs977_not1 & f_arrdiv32_fs976_or0;
  assign f_arrdiv32_fs977_or0 = f_arrdiv32_fs977_and1 | f_arrdiv32_fs977_and0;
  assign f_arrdiv32_fs978_xor0 = f_arrdiv32_mux2to1916_xor0 ^ b[18];
  assign f_arrdiv32_fs978_not0 = ~f_arrdiv32_mux2to1916_xor0;
  assign f_arrdiv32_fs978_and0 = f_arrdiv32_fs978_not0 & b[18];
  assign f_arrdiv32_fs978_xor1 = f_arrdiv32_fs977_or0 ^ f_arrdiv32_fs978_xor0;
  assign f_arrdiv32_fs978_not1 = ~f_arrdiv32_fs978_xor0;
  assign f_arrdiv32_fs978_and1 = f_arrdiv32_fs978_not1 & f_arrdiv32_fs977_or0;
  assign f_arrdiv32_fs978_or0 = f_arrdiv32_fs978_and1 | f_arrdiv32_fs978_and0;
  assign f_arrdiv32_fs979_xor0 = f_arrdiv32_mux2to1917_xor0 ^ b[19];
  assign f_arrdiv32_fs979_not0 = ~f_arrdiv32_mux2to1917_xor0;
  assign f_arrdiv32_fs979_and0 = f_arrdiv32_fs979_not0 & b[19];
  assign f_arrdiv32_fs979_xor1 = f_arrdiv32_fs978_or0 ^ f_arrdiv32_fs979_xor0;
  assign f_arrdiv32_fs979_not1 = ~f_arrdiv32_fs979_xor0;
  assign f_arrdiv32_fs979_and1 = f_arrdiv32_fs979_not1 & f_arrdiv32_fs978_or0;
  assign f_arrdiv32_fs979_or0 = f_arrdiv32_fs979_and1 | f_arrdiv32_fs979_and0;
  assign f_arrdiv32_fs980_xor0 = f_arrdiv32_mux2to1918_xor0 ^ b[20];
  assign f_arrdiv32_fs980_not0 = ~f_arrdiv32_mux2to1918_xor0;
  assign f_arrdiv32_fs980_and0 = f_arrdiv32_fs980_not0 & b[20];
  assign f_arrdiv32_fs980_xor1 = f_arrdiv32_fs979_or0 ^ f_arrdiv32_fs980_xor0;
  assign f_arrdiv32_fs980_not1 = ~f_arrdiv32_fs980_xor0;
  assign f_arrdiv32_fs980_and1 = f_arrdiv32_fs980_not1 & f_arrdiv32_fs979_or0;
  assign f_arrdiv32_fs980_or0 = f_arrdiv32_fs980_and1 | f_arrdiv32_fs980_and0;
  assign f_arrdiv32_fs981_xor0 = f_arrdiv32_mux2to1919_xor0 ^ b[21];
  assign f_arrdiv32_fs981_not0 = ~f_arrdiv32_mux2to1919_xor0;
  assign f_arrdiv32_fs981_and0 = f_arrdiv32_fs981_not0 & b[21];
  assign f_arrdiv32_fs981_xor1 = f_arrdiv32_fs980_or0 ^ f_arrdiv32_fs981_xor0;
  assign f_arrdiv32_fs981_not1 = ~f_arrdiv32_fs981_xor0;
  assign f_arrdiv32_fs981_and1 = f_arrdiv32_fs981_not1 & f_arrdiv32_fs980_or0;
  assign f_arrdiv32_fs981_or0 = f_arrdiv32_fs981_and1 | f_arrdiv32_fs981_and0;
  assign f_arrdiv32_fs982_xor0 = f_arrdiv32_mux2to1920_xor0 ^ b[22];
  assign f_arrdiv32_fs982_not0 = ~f_arrdiv32_mux2to1920_xor0;
  assign f_arrdiv32_fs982_and0 = f_arrdiv32_fs982_not0 & b[22];
  assign f_arrdiv32_fs982_xor1 = f_arrdiv32_fs981_or0 ^ f_arrdiv32_fs982_xor0;
  assign f_arrdiv32_fs982_not1 = ~f_arrdiv32_fs982_xor0;
  assign f_arrdiv32_fs982_and1 = f_arrdiv32_fs982_not1 & f_arrdiv32_fs981_or0;
  assign f_arrdiv32_fs982_or0 = f_arrdiv32_fs982_and1 | f_arrdiv32_fs982_and0;
  assign f_arrdiv32_fs983_xor0 = f_arrdiv32_mux2to1921_xor0 ^ b[23];
  assign f_arrdiv32_fs983_not0 = ~f_arrdiv32_mux2to1921_xor0;
  assign f_arrdiv32_fs983_and0 = f_arrdiv32_fs983_not0 & b[23];
  assign f_arrdiv32_fs983_xor1 = f_arrdiv32_fs982_or0 ^ f_arrdiv32_fs983_xor0;
  assign f_arrdiv32_fs983_not1 = ~f_arrdiv32_fs983_xor0;
  assign f_arrdiv32_fs983_and1 = f_arrdiv32_fs983_not1 & f_arrdiv32_fs982_or0;
  assign f_arrdiv32_fs983_or0 = f_arrdiv32_fs983_and1 | f_arrdiv32_fs983_and0;
  assign f_arrdiv32_fs984_xor0 = f_arrdiv32_mux2to1922_xor0 ^ b[24];
  assign f_arrdiv32_fs984_not0 = ~f_arrdiv32_mux2to1922_xor0;
  assign f_arrdiv32_fs984_and0 = f_arrdiv32_fs984_not0 & b[24];
  assign f_arrdiv32_fs984_xor1 = f_arrdiv32_fs983_or0 ^ f_arrdiv32_fs984_xor0;
  assign f_arrdiv32_fs984_not1 = ~f_arrdiv32_fs984_xor0;
  assign f_arrdiv32_fs984_and1 = f_arrdiv32_fs984_not1 & f_arrdiv32_fs983_or0;
  assign f_arrdiv32_fs984_or0 = f_arrdiv32_fs984_and1 | f_arrdiv32_fs984_and0;
  assign f_arrdiv32_fs985_xor0 = f_arrdiv32_mux2to1923_xor0 ^ b[25];
  assign f_arrdiv32_fs985_not0 = ~f_arrdiv32_mux2to1923_xor0;
  assign f_arrdiv32_fs985_and0 = f_arrdiv32_fs985_not0 & b[25];
  assign f_arrdiv32_fs985_xor1 = f_arrdiv32_fs984_or0 ^ f_arrdiv32_fs985_xor0;
  assign f_arrdiv32_fs985_not1 = ~f_arrdiv32_fs985_xor0;
  assign f_arrdiv32_fs985_and1 = f_arrdiv32_fs985_not1 & f_arrdiv32_fs984_or0;
  assign f_arrdiv32_fs985_or0 = f_arrdiv32_fs985_and1 | f_arrdiv32_fs985_and0;
  assign f_arrdiv32_fs986_xor0 = f_arrdiv32_mux2to1924_xor0 ^ b[26];
  assign f_arrdiv32_fs986_not0 = ~f_arrdiv32_mux2to1924_xor0;
  assign f_arrdiv32_fs986_and0 = f_arrdiv32_fs986_not0 & b[26];
  assign f_arrdiv32_fs986_xor1 = f_arrdiv32_fs985_or0 ^ f_arrdiv32_fs986_xor0;
  assign f_arrdiv32_fs986_not1 = ~f_arrdiv32_fs986_xor0;
  assign f_arrdiv32_fs986_and1 = f_arrdiv32_fs986_not1 & f_arrdiv32_fs985_or0;
  assign f_arrdiv32_fs986_or0 = f_arrdiv32_fs986_and1 | f_arrdiv32_fs986_and0;
  assign f_arrdiv32_fs987_xor0 = f_arrdiv32_mux2to1925_xor0 ^ b[27];
  assign f_arrdiv32_fs987_not0 = ~f_arrdiv32_mux2to1925_xor0;
  assign f_arrdiv32_fs987_and0 = f_arrdiv32_fs987_not0 & b[27];
  assign f_arrdiv32_fs987_xor1 = f_arrdiv32_fs986_or0 ^ f_arrdiv32_fs987_xor0;
  assign f_arrdiv32_fs987_not1 = ~f_arrdiv32_fs987_xor0;
  assign f_arrdiv32_fs987_and1 = f_arrdiv32_fs987_not1 & f_arrdiv32_fs986_or0;
  assign f_arrdiv32_fs987_or0 = f_arrdiv32_fs987_and1 | f_arrdiv32_fs987_and0;
  assign f_arrdiv32_fs988_xor0 = f_arrdiv32_mux2to1926_xor0 ^ b[28];
  assign f_arrdiv32_fs988_not0 = ~f_arrdiv32_mux2to1926_xor0;
  assign f_arrdiv32_fs988_and0 = f_arrdiv32_fs988_not0 & b[28];
  assign f_arrdiv32_fs988_xor1 = f_arrdiv32_fs987_or0 ^ f_arrdiv32_fs988_xor0;
  assign f_arrdiv32_fs988_not1 = ~f_arrdiv32_fs988_xor0;
  assign f_arrdiv32_fs988_and1 = f_arrdiv32_fs988_not1 & f_arrdiv32_fs987_or0;
  assign f_arrdiv32_fs988_or0 = f_arrdiv32_fs988_and1 | f_arrdiv32_fs988_and0;
  assign f_arrdiv32_fs989_xor0 = f_arrdiv32_mux2to1927_xor0 ^ b[29];
  assign f_arrdiv32_fs989_not0 = ~f_arrdiv32_mux2to1927_xor0;
  assign f_arrdiv32_fs989_and0 = f_arrdiv32_fs989_not0 & b[29];
  assign f_arrdiv32_fs989_xor1 = f_arrdiv32_fs988_or0 ^ f_arrdiv32_fs989_xor0;
  assign f_arrdiv32_fs989_not1 = ~f_arrdiv32_fs989_xor0;
  assign f_arrdiv32_fs989_and1 = f_arrdiv32_fs989_not1 & f_arrdiv32_fs988_or0;
  assign f_arrdiv32_fs989_or0 = f_arrdiv32_fs989_and1 | f_arrdiv32_fs989_and0;
  assign f_arrdiv32_fs990_xor0 = f_arrdiv32_mux2to1928_xor0 ^ b[30];
  assign f_arrdiv32_fs990_not0 = ~f_arrdiv32_mux2to1928_xor0;
  assign f_arrdiv32_fs990_and0 = f_arrdiv32_fs990_not0 & b[30];
  assign f_arrdiv32_fs990_xor1 = f_arrdiv32_fs989_or0 ^ f_arrdiv32_fs990_xor0;
  assign f_arrdiv32_fs990_not1 = ~f_arrdiv32_fs990_xor0;
  assign f_arrdiv32_fs990_and1 = f_arrdiv32_fs990_not1 & f_arrdiv32_fs989_or0;
  assign f_arrdiv32_fs990_or0 = f_arrdiv32_fs990_and1 | f_arrdiv32_fs990_and0;
  assign f_arrdiv32_fs991_xor0 = f_arrdiv32_mux2to1929_xor0 ^ b[31];
  assign f_arrdiv32_fs991_not0 = ~f_arrdiv32_mux2to1929_xor0;
  assign f_arrdiv32_fs991_and0 = f_arrdiv32_fs991_not0 & b[31];
  assign f_arrdiv32_fs991_xor1 = f_arrdiv32_fs990_or0 ^ f_arrdiv32_fs991_xor0;
  assign f_arrdiv32_fs991_not1 = ~f_arrdiv32_fs991_xor0;
  assign f_arrdiv32_fs991_and1 = f_arrdiv32_fs991_not1 & f_arrdiv32_fs990_or0;
  assign f_arrdiv32_fs991_or0 = f_arrdiv32_fs991_and1 | f_arrdiv32_fs991_and0;
  assign f_arrdiv32_mux2to1930_and0 = a[1] & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1930_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1930_and1 = f_arrdiv32_fs960_xor0 & f_arrdiv32_mux2to1930_not0;
  assign f_arrdiv32_mux2to1930_xor0 = f_arrdiv32_mux2to1930_and0 ^ f_arrdiv32_mux2to1930_and1;
  assign f_arrdiv32_mux2to1931_and0 = f_arrdiv32_mux2to1899_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1931_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1931_and1 = f_arrdiv32_fs961_xor1 & f_arrdiv32_mux2to1931_not0;
  assign f_arrdiv32_mux2to1931_xor0 = f_arrdiv32_mux2to1931_and0 ^ f_arrdiv32_mux2to1931_and1;
  assign f_arrdiv32_mux2to1932_and0 = f_arrdiv32_mux2to1900_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1932_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1932_and1 = f_arrdiv32_fs962_xor1 & f_arrdiv32_mux2to1932_not0;
  assign f_arrdiv32_mux2to1932_xor0 = f_arrdiv32_mux2to1932_and0 ^ f_arrdiv32_mux2to1932_and1;
  assign f_arrdiv32_mux2to1933_and0 = f_arrdiv32_mux2to1901_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1933_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1933_and1 = f_arrdiv32_fs963_xor1 & f_arrdiv32_mux2to1933_not0;
  assign f_arrdiv32_mux2to1933_xor0 = f_arrdiv32_mux2to1933_and0 ^ f_arrdiv32_mux2to1933_and1;
  assign f_arrdiv32_mux2to1934_and0 = f_arrdiv32_mux2to1902_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1934_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1934_and1 = f_arrdiv32_fs964_xor1 & f_arrdiv32_mux2to1934_not0;
  assign f_arrdiv32_mux2to1934_xor0 = f_arrdiv32_mux2to1934_and0 ^ f_arrdiv32_mux2to1934_and1;
  assign f_arrdiv32_mux2to1935_and0 = f_arrdiv32_mux2to1903_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1935_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1935_and1 = f_arrdiv32_fs965_xor1 & f_arrdiv32_mux2to1935_not0;
  assign f_arrdiv32_mux2to1935_xor0 = f_arrdiv32_mux2to1935_and0 ^ f_arrdiv32_mux2to1935_and1;
  assign f_arrdiv32_mux2to1936_and0 = f_arrdiv32_mux2to1904_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1936_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1936_and1 = f_arrdiv32_fs966_xor1 & f_arrdiv32_mux2to1936_not0;
  assign f_arrdiv32_mux2to1936_xor0 = f_arrdiv32_mux2to1936_and0 ^ f_arrdiv32_mux2to1936_and1;
  assign f_arrdiv32_mux2to1937_and0 = f_arrdiv32_mux2to1905_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1937_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1937_and1 = f_arrdiv32_fs967_xor1 & f_arrdiv32_mux2to1937_not0;
  assign f_arrdiv32_mux2to1937_xor0 = f_arrdiv32_mux2to1937_and0 ^ f_arrdiv32_mux2to1937_and1;
  assign f_arrdiv32_mux2to1938_and0 = f_arrdiv32_mux2to1906_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1938_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1938_and1 = f_arrdiv32_fs968_xor1 & f_arrdiv32_mux2to1938_not0;
  assign f_arrdiv32_mux2to1938_xor0 = f_arrdiv32_mux2to1938_and0 ^ f_arrdiv32_mux2to1938_and1;
  assign f_arrdiv32_mux2to1939_and0 = f_arrdiv32_mux2to1907_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1939_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1939_and1 = f_arrdiv32_fs969_xor1 & f_arrdiv32_mux2to1939_not0;
  assign f_arrdiv32_mux2to1939_xor0 = f_arrdiv32_mux2to1939_and0 ^ f_arrdiv32_mux2to1939_and1;
  assign f_arrdiv32_mux2to1940_and0 = f_arrdiv32_mux2to1908_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1940_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1940_and1 = f_arrdiv32_fs970_xor1 & f_arrdiv32_mux2to1940_not0;
  assign f_arrdiv32_mux2to1940_xor0 = f_arrdiv32_mux2to1940_and0 ^ f_arrdiv32_mux2to1940_and1;
  assign f_arrdiv32_mux2to1941_and0 = f_arrdiv32_mux2to1909_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1941_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1941_and1 = f_arrdiv32_fs971_xor1 & f_arrdiv32_mux2to1941_not0;
  assign f_arrdiv32_mux2to1941_xor0 = f_arrdiv32_mux2to1941_and0 ^ f_arrdiv32_mux2to1941_and1;
  assign f_arrdiv32_mux2to1942_and0 = f_arrdiv32_mux2to1910_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1942_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1942_and1 = f_arrdiv32_fs972_xor1 & f_arrdiv32_mux2to1942_not0;
  assign f_arrdiv32_mux2to1942_xor0 = f_arrdiv32_mux2to1942_and0 ^ f_arrdiv32_mux2to1942_and1;
  assign f_arrdiv32_mux2to1943_and0 = f_arrdiv32_mux2to1911_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1943_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1943_and1 = f_arrdiv32_fs973_xor1 & f_arrdiv32_mux2to1943_not0;
  assign f_arrdiv32_mux2to1943_xor0 = f_arrdiv32_mux2to1943_and0 ^ f_arrdiv32_mux2to1943_and1;
  assign f_arrdiv32_mux2to1944_and0 = f_arrdiv32_mux2to1912_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1944_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1944_and1 = f_arrdiv32_fs974_xor1 & f_arrdiv32_mux2to1944_not0;
  assign f_arrdiv32_mux2to1944_xor0 = f_arrdiv32_mux2to1944_and0 ^ f_arrdiv32_mux2to1944_and1;
  assign f_arrdiv32_mux2to1945_and0 = f_arrdiv32_mux2to1913_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1945_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1945_and1 = f_arrdiv32_fs975_xor1 & f_arrdiv32_mux2to1945_not0;
  assign f_arrdiv32_mux2to1945_xor0 = f_arrdiv32_mux2to1945_and0 ^ f_arrdiv32_mux2to1945_and1;
  assign f_arrdiv32_mux2to1946_and0 = f_arrdiv32_mux2to1914_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1946_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1946_and1 = f_arrdiv32_fs976_xor1 & f_arrdiv32_mux2to1946_not0;
  assign f_arrdiv32_mux2to1946_xor0 = f_arrdiv32_mux2to1946_and0 ^ f_arrdiv32_mux2to1946_and1;
  assign f_arrdiv32_mux2to1947_and0 = f_arrdiv32_mux2to1915_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1947_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1947_and1 = f_arrdiv32_fs977_xor1 & f_arrdiv32_mux2to1947_not0;
  assign f_arrdiv32_mux2to1947_xor0 = f_arrdiv32_mux2to1947_and0 ^ f_arrdiv32_mux2to1947_and1;
  assign f_arrdiv32_mux2to1948_and0 = f_arrdiv32_mux2to1916_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1948_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1948_and1 = f_arrdiv32_fs978_xor1 & f_arrdiv32_mux2to1948_not0;
  assign f_arrdiv32_mux2to1948_xor0 = f_arrdiv32_mux2to1948_and0 ^ f_arrdiv32_mux2to1948_and1;
  assign f_arrdiv32_mux2to1949_and0 = f_arrdiv32_mux2to1917_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1949_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1949_and1 = f_arrdiv32_fs979_xor1 & f_arrdiv32_mux2to1949_not0;
  assign f_arrdiv32_mux2to1949_xor0 = f_arrdiv32_mux2to1949_and0 ^ f_arrdiv32_mux2to1949_and1;
  assign f_arrdiv32_mux2to1950_and0 = f_arrdiv32_mux2to1918_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1950_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1950_and1 = f_arrdiv32_fs980_xor1 & f_arrdiv32_mux2to1950_not0;
  assign f_arrdiv32_mux2to1950_xor0 = f_arrdiv32_mux2to1950_and0 ^ f_arrdiv32_mux2to1950_and1;
  assign f_arrdiv32_mux2to1951_and0 = f_arrdiv32_mux2to1919_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1951_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1951_and1 = f_arrdiv32_fs981_xor1 & f_arrdiv32_mux2to1951_not0;
  assign f_arrdiv32_mux2to1951_xor0 = f_arrdiv32_mux2to1951_and0 ^ f_arrdiv32_mux2to1951_and1;
  assign f_arrdiv32_mux2to1952_and0 = f_arrdiv32_mux2to1920_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1952_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1952_and1 = f_arrdiv32_fs982_xor1 & f_arrdiv32_mux2to1952_not0;
  assign f_arrdiv32_mux2to1952_xor0 = f_arrdiv32_mux2to1952_and0 ^ f_arrdiv32_mux2to1952_and1;
  assign f_arrdiv32_mux2to1953_and0 = f_arrdiv32_mux2to1921_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1953_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1953_and1 = f_arrdiv32_fs983_xor1 & f_arrdiv32_mux2to1953_not0;
  assign f_arrdiv32_mux2to1953_xor0 = f_arrdiv32_mux2to1953_and0 ^ f_arrdiv32_mux2to1953_and1;
  assign f_arrdiv32_mux2to1954_and0 = f_arrdiv32_mux2to1922_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1954_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1954_and1 = f_arrdiv32_fs984_xor1 & f_arrdiv32_mux2to1954_not0;
  assign f_arrdiv32_mux2to1954_xor0 = f_arrdiv32_mux2to1954_and0 ^ f_arrdiv32_mux2to1954_and1;
  assign f_arrdiv32_mux2to1955_and0 = f_arrdiv32_mux2to1923_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1955_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1955_and1 = f_arrdiv32_fs985_xor1 & f_arrdiv32_mux2to1955_not0;
  assign f_arrdiv32_mux2to1955_xor0 = f_arrdiv32_mux2to1955_and0 ^ f_arrdiv32_mux2to1955_and1;
  assign f_arrdiv32_mux2to1956_and0 = f_arrdiv32_mux2to1924_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1956_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1956_and1 = f_arrdiv32_fs986_xor1 & f_arrdiv32_mux2to1956_not0;
  assign f_arrdiv32_mux2to1956_xor0 = f_arrdiv32_mux2to1956_and0 ^ f_arrdiv32_mux2to1956_and1;
  assign f_arrdiv32_mux2to1957_and0 = f_arrdiv32_mux2to1925_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1957_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1957_and1 = f_arrdiv32_fs987_xor1 & f_arrdiv32_mux2to1957_not0;
  assign f_arrdiv32_mux2to1957_xor0 = f_arrdiv32_mux2to1957_and0 ^ f_arrdiv32_mux2to1957_and1;
  assign f_arrdiv32_mux2to1958_and0 = f_arrdiv32_mux2to1926_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1958_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1958_and1 = f_arrdiv32_fs988_xor1 & f_arrdiv32_mux2to1958_not0;
  assign f_arrdiv32_mux2to1958_xor0 = f_arrdiv32_mux2to1958_and0 ^ f_arrdiv32_mux2to1958_and1;
  assign f_arrdiv32_mux2to1959_and0 = f_arrdiv32_mux2to1927_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1959_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1959_and1 = f_arrdiv32_fs989_xor1 & f_arrdiv32_mux2to1959_not0;
  assign f_arrdiv32_mux2to1959_xor0 = f_arrdiv32_mux2to1959_and0 ^ f_arrdiv32_mux2to1959_and1;
  assign f_arrdiv32_mux2to1960_and0 = f_arrdiv32_mux2to1928_xor0 & f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1960_not0 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_mux2to1960_and1 = f_arrdiv32_fs990_xor1 & f_arrdiv32_mux2to1960_not0;
  assign f_arrdiv32_mux2to1960_xor0 = f_arrdiv32_mux2to1960_and0 ^ f_arrdiv32_mux2to1960_and1;
  assign f_arrdiv32_not30 = ~f_arrdiv32_fs991_or0;
  assign f_arrdiv32_fs992_xor0 = a[0] ^ b[0];
  assign f_arrdiv32_fs992_not0 = ~a[0];
  assign f_arrdiv32_fs992_and0 = f_arrdiv32_fs992_not0 & b[0];
  assign f_arrdiv32_fs992_not1 = ~f_arrdiv32_fs992_xor0;
  assign f_arrdiv32_fs993_xor0 = f_arrdiv32_mux2to1930_xor0 ^ b[1];
  assign f_arrdiv32_fs993_not0 = ~f_arrdiv32_mux2to1930_xor0;
  assign f_arrdiv32_fs993_and0 = f_arrdiv32_fs993_not0 & b[1];
  assign f_arrdiv32_fs993_xor1 = f_arrdiv32_fs992_and0 ^ f_arrdiv32_fs993_xor0;
  assign f_arrdiv32_fs993_not1 = ~f_arrdiv32_fs993_xor0;
  assign f_arrdiv32_fs993_and1 = f_arrdiv32_fs993_not1 & f_arrdiv32_fs992_and0;
  assign f_arrdiv32_fs993_or0 = f_arrdiv32_fs993_and1 | f_arrdiv32_fs993_and0;
  assign f_arrdiv32_fs994_xor0 = f_arrdiv32_mux2to1931_xor0 ^ b[2];
  assign f_arrdiv32_fs994_not0 = ~f_arrdiv32_mux2to1931_xor0;
  assign f_arrdiv32_fs994_and0 = f_arrdiv32_fs994_not0 & b[2];
  assign f_arrdiv32_fs994_xor1 = f_arrdiv32_fs993_or0 ^ f_arrdiv32_fs994_xor0;
  assign f_arrdiv32_fs994_not1 = ~f_arrdiv32_fs994_xor0;
  assign f_arrdiv32_fs994_and1 = f_arrdiv32_fs994_not1 & f_arrdiv32_fs993_or0;
  assign f_arrdiv32_fs994_or0 = f_arrdiv32_fs994_and1 | f_arrdiv32_fs994_and0;
  assign f_arrdiv32_fs995_xor0 = f_arrdiv32_mux2to1932_xor0 ^ b[3];
  assign f_arrdiv32_fs995_not0 = ~f_arrdiv32_mux2to1932_xor0;
  assign f_arrdiv32_fs995_and0 = f_arrdiv32_fs995_not0 & b[3];
  assign f_arrdiv32_fs995_xor1 = f_arrdiv32_fs994_or0 ^ f_arrdiv32_fs995_xor0;
  assign f_arrdiv32_fs995_not1 = ~f_arrdiv32_fs995_xor0;
  assign f_arrdiv32_fs995_and1 = f_arrdiv32_fs995_not1 & f_arrdiv32_fs994_or0;
  assign f_arrdiv32_fs995_or0 = f_arrdiv32_fs995_and1 | f_arrdiv32_fs995_and0;
  assign f_arrdiv32_fs996_xor0 = f_arrdiv32_mux2to1933_xor0 ^ b[4];
  assign f_arrdiv32_fs996_not0 = ~f_arrdiv32_mux2to1933_xor0;
  assign f_arrdiv32_fs996_and0 = f_arrdiv32_fs996_not0 & b[4];
  assign f_arrdiv32_fs996_xor1 = f_arrdiv32_fs995_or0 ^ f_arrdiv32_fs996_xor0;
  assign f_arrdiv32_fs996_not1 = ~f_arrdiv32_fs996_xor0;
  assign f_arrdiv32_fs996_and1 = f_arrdiv32_fs996_not1 & f_arrdiv32_fs995_or0;
  assign f_arrdiv32_fs996_or0 = f_arrdiv32_fs996_and1 | f_arrdiv32_fs996_and0;
  assign f_arrdiv32_fs997_xor0 = f_arrdiv32_mux2to1934_xor0 ^ b[5];
  assign f_arrdiv32_fs997_not0 = ~f_arrdiv32_mux2to1934_xor0;
  assign f_arrdiv32_fs997_and0 = f_arrdiv32_fs997_not0 & b[5];
  assign f_arrdiv32_fs997_xor1 = f_arrdiv32_fs996_or0 ^ f_arrdiv32_fs997_xor0;
  assign f_arrdiv32_fs997_not1 = ~f_arrdiv32_fs997_xor0;
  assign f_arrdiv32_fs997_and1 = f_arrdiv32_fs997_not1 & f_arrdiv32_fs996_or0;
  assign f_arrdiv32_fs997_or0 = f_arrdiv32_fs997_and1 | f_arrdiv32_fs997_and0;
  assign f_arrdiv32_fs998_xor0 = f_arrdiv32_mux2to1935_xor0 ^ b[6];
  assign f_arrdiv32_fs998_not0 = ~f_arrdiv32_mux2to1935_xor0;
  assign f_arrdiv32_fs998_and0 = f_arrdiv32_fs998_not0 & b[6];
  assign f_arrdiv32_fs998_xor1 = f_arrdiv32_fs997_or0 ^ f_arrdiv32_fs998_xor0;
  assign f_arrdiv32_fs998_not1 = ~f_arrdiv32_fs998_xor0;
  assign f_arrdiv32_fs998_and1 = f_arrdiv32_fs998_not1 & f_arrdiv32_fs997_or0;
  assign f_arrdiv32_fs998_or0 = f_arrdiv32_fs998_and1 | f_arrdiv32_fs998_and0;
  assign f_arrdiv32_fs999_xor0 = f_arrdiv32_mux2to1936_xor0 ^ b[7];
  assign f_arrdiv32_fs999_not0 = ~f_arrdiv32_mux2to1936_xor0;
  assign f_arrdiv32_fs999_and0 = f_arrdiv32_fs999_not0 & b[7];
  assign f_arrdiv32_fs999_xor1 = f_arrdiv32_fs998_or0 ^ f_arrdiv32_fs999_xor0;
  assign f_arrdiv32_fs999_not1 = ~f_arrdiv32_fs999_xor0;
  assign f_arrdiv32_fs999_and1 = f_arrdiv32_fs999_not1 & f_arrdiv32_fs998_or0;
  assign f_arrdiv32_fs999_or0 = f_arrdiv32_fs999_and1 | f_arrdiv32_fs999_and0;
  assign f_arrdiv32_fs1000_xor0 = f_arrdiv32_mux2to1937_xor0 ^ b[8];
  assign f_arrdiv32_fs1000_not0 = ~f_arrdiv32_mux2to1937_xor0;
  assign f_arrdiv32_fs1000_and0 = f_arrdiv32_fs1000_not0 & b[8];
  assign f_arrdiv32_fs1000_xor1 = f_arrdiv32_fs999_or0 ^ f_arrdiv32_fs1000_xor0;
  assign f_arrdiv32_fs1000_not1 = ~f_arrdiv32_fs1000_xor0;
  assign f_arrdiv32_fs1000_and1 = f_arrdiv32_fs1000_not1 & f_arrdiv32_fs999_or0;
  assign f_arrdiv32_fs1000_or0 = f_arrdiv32_fs1000_and1 | f_arrdiv32_fs1000_and0;
  assign f_arrdiv32_fs1001_xor0 = f_arrdiv32_mux2to1938_xor0 ^ b[9];
  assign f_arrdiv32_fs1001_not0 = ~f_arrdiv32_mux2to1938_xor0;
  assign f_arrdiv32_fs1001_and0 = f_arrdiv32_fs1001_not0 & b[9];
  assign f_arrdiv32_fs1001_xor1 = f_arrdiv32_fs1000_or0 ^ f_arrdiv32_fs1001_xor0;
  assign f_arrdiv32_fs1001_not1 = ~f_arrdiv32_fs1001_xor0;
  assign f_arrdiv32_fs1001_and1 = f_arrdiv32_fs1001_not1 & f_arrdiv32_fs1000_or0;
  assign f_arrdiv32_fs1001_or0 = f_arrdiv32_fs1001_and1 | f_arrdiv32_fs1001_and0;
  assign f_arrdiv32_fs1002_xor0 = f_arrdiv32_mux2to1939_xor0 ^ b[10];
  assign f_arrdiv32_fs1002_not0 = ~f_arrdiv32_mux2to1939_xor0;
  assign f_arrdiv32_fs1002_and0 = f_arrdiv32_fs1002_not0 & b[10];
  assign f_arrdiv32_fs1002_xor1 = f_arrdiv32_fs1001_or0 ^ f_arrdiv32_fs1002_xor0;
  assign f_arrdiv32_fs1002_not1 = ~f_arrdiv32_fs1002_xor0;
  assign f_arrdiv32_fs1002_and1 = f_arrdiv32_fs1002_not1 & f_arrdiv32_fs1001_or0;
  assign f_arrdiv32_fs1002_or0 = f_arrdiv32_fs1002_and1 | f_arrdiv32_fs1002_and0;
  assign f_arrdiv32_fs1003_xor0 = f_arrdiv32_mux2to1940_xor0 ^ b[11];
  assign f_arrdiv32_fs1003_not0 = ~f_arrdiv32_mux2to1940_xor0;
  assign f_arrdiv32_fs1003_and0 = f_arrdiv32_fs1003_not0 & b[11];
  assign f_arrdiv32_fs1003_xor1 = f_arrdiv32_fs1002_or0 ^ f_arrdiv32_fs1003_xor0;
  assign f_arrdiv32_fs1003_not1 = ~f_arrdiv32_fs1003_xor0;
  assign f_arrdiv32_fs1003_and1 = f_arrdiv32_fs1003_not1 & f_arrdiv32_fs1002_or0;
  assign f_arrdiv32_fs1003_or0 = f_arrdiv32_fs1003_and1 | f_arrdiv32_fs1003_and0;
  assign f_arrdiv32_fs1004_xor0 = f_arrdiv32_mux2to1941_xor0 ^ b[12];
  assign f_arrdiv32_fs1004_not0 = ~f_arrdiv32_mux2to1941_xor0;
  assign f_arrdiv32_fs1004_and0 = f_arrdiv32_fs1004_not0 & b[12];
  assign f_arrdiv32_fs1004_xor1 = f_arrdiv32_fs1003_or0 ^ f_arrdiv32_fs1004_xor0;
  assign f_arrdiv32_fs1004_not1 = ~f_arrdiv32_fs1004_xor0;
  assign f_arrdiv32_fs1004_and1 = f_arrdiv32_fs1004_not1 & f_arrdiv32_fs1003_or0;
  assign f_arrdiv32_fs1004_or0 = f_arrdiv32_fs1004_and1 | f_arrdiv32_fs1004_and0;
  assign f_arrdiv32_fs1005_xor0 = f_arrdiv32_mux2to1942_xor0 ^ b[13];
  assign f_arrdiv32_fs1005_not0 = ~f_arrdiv32_mux2to1942_xor0;
  assign f_arrdiv32_fs1005_and0 = f_arrdiv32_fs1005_not0 & b[13];
  assign f_arrdiv32_fs1005_xor1 = f_arrdiv32_fs1004_or0 ^ f_arrdiv32_fs1005_xor0;
  assign f_arrdiv32_fs1005_not1 = ~f_arrdiv32_fs1005_xor0;
  assign f_arrdiv32_fs1005_and1 = f_arrdiv32_fs1005_not1 & f_arrdiv32_fs1004_or0;
  assign f_arrdiv32_fs1005_or0 = f_arrdiv32_fs1005_and1 | f_arrdiv32_fs1005_and0;
  assign f_arrdiv32_fs1006_xor0 = f_arrdiv32_mux2to1943_xor0 ^ b[14];
  assign f_arrdiv32_fs1006_not0 = ~f_arrdiv32_mux2to1943_xor0;
  assign f_arrdiv32_fs1006_and0 = f_arrdiv32_fs1006_not0 & b[14];
  assign f_arrdiv32_fs1006_xor1 = f_arrdiv32_fs1005_or0 ^ f_arrdiv32_fs1006_xor0;
  assign f_arrdiv32_fs1006_not1 = ~f_arrdiv32_fs1006_xor0;
  assign f_arrdiv32_fs1006_and1 = f_arrdiv32_fs1006_not1 & f_arrdiv32_fs1005_or0;
  assign f_arrdiv32_fs1006_or0 = f_arrdiv32_fs1006_and1 | f_arrdiv32_fs1006_and0;
  assign f_arrdiv32_fs1007_xor0 = f_arrdiv32_mux2to1944_xor0 ^ b[15];
  assign f_arrdiv32_fs1007_not0 = ~f_arrdiv32_mux2to1944_xor0;
  assign f_arrdiv32_fs1007_and0 = f_arrdiv32_fs1007_not0 & b[15];
  assign f_arrdiv32_fs1007_xor1 = f_arrdiv32_fs1006_or0 ^ f_arrdiv32_fs1007_xor0;
  assign f_arrdiv32_fs1007_not1 = ~f_arrdiv32_fs1007_xor0;
  assign f_arrdiv32_fs1007_and1 = f_arrdiv32_fs1007_not1 & f_arrdiv32_fs1006_or0;
  assign f_arrdiv32_fs1007_or0 = f_arrdiv32_fs1007_and1 | f_arrdiv32_fs1007_and0;
  assign f_arrdiv32_fs1008_xor0 = f_arrdiv32_mux2to1945_xor0 ^ b[16];
  assign f_arrdiv32_fs1008_not0 = ~f_arrdiv32_mux2to1945_xor0;
  assign f_arrdiv32_fs1008_and0 = f_arrdiv32_fs1008_not0 & b[16];
  assign f_arrdiv32_fs1008_xor1 = f_arrdiv32_fs1007_or0 ^ f_arrdiv32_fs1008_xor0;
  assign f_arrdiv32_fs1008_not1 = ~f_arrdiv32_fs1008_xor0;
  assign f_arrdiv32_fs1008_and1 = f_arrdiv32_fs1008_not1 & f_arrdiv32_fs1007_or0;
  assign f_arrdiv32_fs1008_or0 = f_arrdiv32_fs1008_and1 | f_arrdiv32_fs1008_and0;
  assign f_arrdiv32_fs1009_xor0 = f_arrdiv32_mux2to1946_xor0 ^ b[17];
  assign f_arrdiv32_fs1009_not0 = ~f_arrdiv32_mux2to1946_xor0;
  assign f_arrdiv32_fs1009_and0 = f_arrdiv32_fs1009_not0 & b[17];
  assign f_arrdiv32_fs1009_xor1 = f_arrdiv32_fs1008_or0 ^ f_arrdiv32_fs1009_xor0;
  assign f_arrdiv32_fs1009_not1 = ~f_arrdiv32_fs1009_xor0;
  assign f_arrdiv32_fs1009_and1 = f_arrdiv32_fs1009_not1 & f_arrdiv32_fs1008_or0;
  assign f_arrdiv32_fs1009_or0 = f_arrdiv32_fs1009_and1 | f_arrdiv32_fs1009_and0;
  assign f_arrdiv32_fs1010_xor0 = f_arrdiv32_mux2to1947_xor0 ^ b[18];
  assign f_arrdiv32_fs1010_not0 = ~f_arrdiv32_mux2to1947_xor0;
  assign f_arrdiv32_fs1010_and0 = f_arrdiv32_fs1010_not0 & b[18];
  assign f_arrdiv32_fs1010_xor1 = f_arrdiv32_fs1009_or0 ^ f_arrdiv32_fs1010_xor0;
  assign f_arrdiv32_fs1010_not1 = ~f_arrdiv32_fs1010_xor0;
  assign f_arrdiv32_fs1010_and1 = f_arrdiv32_fs1010_not1 & f_arrdiv32_fs1009_or0;
  assign f_arrdiv32_fs1010_or0 = f_arrdiv32_fs1010_and1 | f_arrdiv32_fs1010_and0;
  assign f_arrdiv32_fs1011_xor0 = f_arrdiv32_mux2to1948_xor0 ^ b[19];
  assign f_arrdiv32_fs1011_not0 = ~f_arrdiv32_mux2to1948_xor0;
  assign f_arrdiv32_fs1011_and0 = f_arrdiv32_fs1011_not0 & b[19];
  assign f_arrdiv32_fs1011_xor1 = f_arrdiv32_fs1010_or0 ^ f_arrdiv32_fs1011_xor0;
  assign f_arrdiv32_fs1011_not1 = ~f_arrdiv32_fs1011_xor0;
  assign f_arrdiv32_fs1011_and1 = f_arrdiv32_fs1011_not1 & f_arrdiv32_fs1010_or0;
  assign f_arrdiv32_fs1011_or0 = f_arrdiv32_fs1011_and1 | f_arrdiv32_fs1011_and0;
  assign f_arrdiv32_fs1012_xor0 = f_arrdiv32_mux2to1949_xor0 ^ b[20];
  assign f_arrdiv32_fs1012_not0 = ~f_arrdiv32_mux2to1949_xor0;
  assign f_arrdiv32_fs1012_and0 = f_arrdiv32_fs1012_not0 & b[20];
  assign f_arrdiv32_fs1012_xor1 = f_arrdiv32_fs1011_or0 ^ f_arrdiv32_fs1012_xor0;
  assign f_arrdiv32_fs1012_not1 = ~f_arrdiv32_fs1012_xor0;
  assign f_arrdiv32_fs1012_and1 = f_arrdiv32_fs1012_not1 & f_arrdiv32_fs1011_or0;
  assign f_arrdiv32_fs1012_or0 = f_arrdiv32_fs1012_and1 | f_arrdiv32_fs1012_and0;
  assign f_arrdiv32_fs1013_xor0 = f_arrdiv32_mux2to1950_xor0 ^ b[21];
  assign f_arrdiv32_fs1013_not0 = ~f_arrdiv32_mux2to1950_xor0;
  assign f_arrdiv32_fs1013_and0 = f_arrdiv32_fs1013_not0 & b[21];
  assign f_arrdiv32_fs1013_xor1 = f_arrdiv32_fs1012_or0 ^ f_arrdiv32_fs1013_xor0;
  assign f_arrdiv32_fs1013_not1 = ~f_arrdiv32_fs1013_xor0;
  assign f_arrdiv32_fs1013_and1 = f_arrdiv32_fs1013_not1 & f_arrdiv32_fs1012_or0;
  assign f_arrdiv32_fs1013_or0 = f_arrdiv32_fs1013_and1 | f_arrdiv32_fs1013_and0;
  assign f_arrdiv32_fs1014_xor0 = f_arrdiv32_mux2to1951_xor0 ^ b[22];
  assign f_arrdiv32_fs1014_not0 = ~f_arrdiv32_mux2to1951_xor0;
  assign f_arrdiv32_fs1014_and0 = f_arrdiv32_fs1014_not0 & b[22];
  assign f_arrdiv32_fs1014_xor1 = f_arrdiv32_fs1013_or0 ^ f_arrdiv32_fs1014_xor0;
  assign f_arrdiv32_fs1014_not1 = ~f_arrdiv32_fs1014_xor0;
  assign f_arrdiv32_fs1014_and1 = f_arrdiv32_fs1014_not1 & f_arrdiv32_fs1013_or0;
  assign f_arrdiv32_fs1014_or0 = f_arrdiv32_fs1014_and1 | f_arrdiv32_fs1014_and0;
  assign f_arrdiv32_fs1015_xor0 = f_arrdiv32_mux2to1952_xor0 ^ b[23];
  assign f_arrdiv32_fs1015_not0 = ~f_arrdiv32_mux2to1952_xor0;
  assign f_arrdiv32_fs1015_and0 = f_arrdiv32_fs1015_not0 & b[23];
  assign f_arrdiv32_fs1015_xor1 = f_arrdiv32_fs1014_or0 ^ f_arrdiv32_fs1015_xor0;
  assign f_arrdiv32_fs1015_not1 = ~f_arrdiv32_fs1015_xor0;
  assign f_arrdiv32_fs1015_and1 = f_arrdiv32_fs1015_not1 & f_arrdiv32_fs1014_or0;
  assign f_arrdiv32_fs1015_or0 = f_arrdiv32_fs1015_and1 | f_arrdiv32_fs1015_and0;
  assign f_arrdiv32_fs1016_xor0 = f_arrdiv32_mux2to1953_xor0 ^ b[24];
  assign f_arrdiv32_fs1016_not0 = ~f_arrdiv32_mux2to1953_xor0;
  assign f_arrdiv32_fs1016_and0 = f_arrdiv32_fs1016_not0 & b[24];
  assign f_arrdiv32_fs1016_xor1 = f_arrdiv32_fs1015_or0 ^ f_arrdiv32_fs1016_xor0;
  assign f_arrdiv32_fs1016_not1 = ~f_arrdiv32_fs1016_xor0;
  assign f_arrdiv32_fs1016_and1 = f_arrdiv32_fs1016_not1 & f_arrdiv32_fs1015_or0;
  assign f_arrdiv32_fs1016_or0 = f_arrdiv32_fs1016_and1 | f_arrdiv32_fs1016_and0;
  assign f_arrdiv32_fs1017_xor0 = f_arrdiv32_mux2to1954_xor0 ^ b[25];
  assign f_arrdiv32_fs1017_not0 = ~f_arrdiv32_mux2to1954_xor0;
  assign f_arrdiv32_fs1017_and0 = f_arrdiv32_fs1017_not0 & b[25];
  assign f_arrdiv32_fs1017_xor1 = f_arrdiv32_fs1016_or0 ^ f_arrdiv32_fs1017_xor0;
  assign f_arrdiv32_fs1017_not1 = ~f_arrdiv32_fs1017_xor0;
  assign f_arrdiv32_fs1017_and1 = f_arrdiv32_fs1017_not1 & f_arrdiv32_fs1016_or0;
  assign f_arrdiv32_fs1017_or0 = f_arrdiv32_fs1017_and1 | f_arrdiv32_fs1017_and0;
  assign f_arrdiv32_fs1018_xor0 = f_arrdiv32_mux2to1955_xor0 ^ b[26];
  assign f_arrdiv32_fs1018_not0 = ~f_arrdiv32_mux2to1955_xor0;
  assign f_arrdiv32_fs1018_and0 = f_arrdiv32_fs1018_not0 & b[26];
  assign f_arrdiv32_fs1018_xor1 = f_arrdiv32_fs1017_or0 ^ f_arrdiv32_fs1018_xor0;
  assign f_arrdiv32_fs1018_not1 = ~f_arrdiv32_fs1018_xor0;
  assign f_arrdiv32_fs1018_and1 = f_arrdiv32_fs1018_not1 & f_arrdiv32_fs1017_or0;
  assign f_arrdiv32_fs1018_or0 = f_arrdiv32_fs1018_and1 | f_arrdiv32_fs1018_and0;
  assign f_arrdiv32_fs1019_xor0 = f_arrdiv32_mux2to1956_xor0 ^ b[27];
  assign f_arrdiv32_fs1019_not0 = ~f_arrdiv32_mux2to1956_xor0;
  assign f_arrdiv32_fs1019_and0 = f_arrdiv32_fs1019_not0 & b[27];
  assign f_arrdiv32_fs1019_xor1 = f_arrdiv32_fs1018_or0 ^ f_arrdiv32_fs1019_xor0;
  assign f_arrdiv32_fs1019_not1 = ~f_arrdiv32_fs1019_xor0;
  assign f_arrdiv32_fs1019_and1 = f_arrdiv32_fs1019_not1 & f_arrdiv32_fs1018_or0;
  assign f_arrdiv32_fs1019_or0 = f_arrdiv32_fs1019_and1 | f_arrdiv32_fs1019_and0;
  assign f_arrdiv32_fs1020_xor0 = f_arrdiv32_mux2to1957_xor0 ^ b[28];
  assign f_arrdiv32_fs1020_not0 = ~f_arrdiv32_mux2to1957_xor0;
  assign f_arrdiv32_fs1020_and0 = f_arrdiv32_fs1020_not0 & b[28];
  assign f_arrdiv32_fs1020_xor1 = f_arrdiv32_fs1019_or0 ^ f_arrdiv32_fs1020_xor0;
  assign f_arrdiv32_fs1020_not1 = ~f_arrdiv32_fs1020_xor0;
  assign f_arrdiv32_fs1020_and1 = f_arrdiv32_fs1020_not1 & f_arrdiv32_fs1019_or0;
  assign f_arrdiv32_fs1020_or0 = f_arrdiv32_fs1020_and1 | f_arrdiv32_fs1020_and0;
  assign f_arrdiv32_fs1021_xor0 = f_arrdiv32_mux2to1958_xor0 ^ b[29];
  assign f_arrdiv32_fs1021_not0 = ~f_arrdiv32_mux2to1958_xor0;
  assign f_arrdiv32_fs1021_and0 = f_arrdiv32_fs1021_not0 & b[29];
  assign f_arrdiv32_fs1021_xor1 = f_arrdiv32_fs1020_or0 ^ f_arrdiv32_fs1021_xor0;
  assign f_arrdiv32_fs1021_not1 = ~f_arrdiv32_fs1021_xor0;
  assign f_arrdiv32_fs1021_and1 = f_arrdiv32_fs1021_not1 & f_arrdiv32_fs1020_or0;
  assign f_arrdiv32_fs1021_or0 = f_arrdiv32_fs1021_and1 | f_arrdiv32_fs1021_and0;
  assign f_arrdiv32_fs1022_xor0 = f_arrdiv32_mux2to1959_xor0 ^ b[30];
  assign f_arrdiv32_fs1022_not0 = ~f_arrdiv32_mux2to1959_xor0;
  assign f_arrdiv32_fs1022_and0 = f_arrdiv32_fs1022_not0 & b[30];
  assign f_arrdiv32_fs1022_xor1 = f_arrdiv32_fs1021_or0 ^ f_arrdiv32_fs1022_xor0;
  assign f_arrdiv32_fs1022_not1 = ~f_arrdiv32_fs1022_xor0;
  assign f_arrdiv32_fs1022_and1 = f_arrdiv32_fs1022_not1 & f_arrdiv32_fs1021_or0;
  assign f_arrdiv32_fs1022_or0 = f_arrdiv32_fs1022_and1 | f_arrdiv32_fs1022_and0;
  assign f_arrdiv32_fs1023_xor0 = f_arrdiv32_mux2to1960_xor0 ^ b[31];
  assign f_arrdiv32_fs1023_not0 = ~f_arrdiv32_mux2to1960_xor0;
  assign f_arrdiv32_fs1023_and0 = f_arrdiv32_fs1023_not0 & b[31];
  assign f_arrdiv32_fs1023_xor1 = f_arrdiv32_fs1022_or0 ^ f_arrdiv32_fs1023_xor0;
  assign f_arrdiv32_fs1023_not1 = ~f_arrdiv32_fs1023_xor0;
  assign f_arrdiv32_fs1023_and1 = f_arrdiv32_fs1023_not1 & f_arrdiv32_fs1022_or0;
  assign f_arrdiv32_fs1023_or0 = f_arrdiv32_fs1023_and1 | f_arrdiv32_fs1023_and0;
  assign f_arrdiv32_not31 = ~f_arrdiv32_fs1023_or0;

  assign f_arrdiv32_out[0] = f_arrdiv32_not31;
  assign f_arrdiv32_out[1] = f_arrdiv32_not30;
  assign f_arrdiv32_out[2] = f_arrdiv32_not29;
  assign f_arrdiv32_out[3] = f_arrdiv32_not28;
  assign f_arrdiv32_out[4] = f_arrdiv32_not27;
  assign f_arrdiv32_out[5] = f_arrdiv32_not26;
  assign f_arrdiv32_out[6] = f_arrdiv32_not25;
  assign f_arrdiv32_out[7] = f_arrdiv32_not24;
  assign f_arrdiv32_out[8] = f_arrdiv32_not23;
  assign f_arrdiv32_out[9] = f_arrdiv32_not22;
  assign f_arrdiv32_out[10] = f_arrdiv32_not21;
  assign f_arrdiv32_out[11] = f_arrdiv32_not20;
  assign f_arrdiv32_out[12] = f_arrdiv32_not19;
  assign f_arrdiv32_out[13] = f_arrdiv32_not18;
  assign f_arrdiv32_out[14] = f_arrdiv32_not17;
  assign f_arrdiv32_out[15] = f_arrdiv32_not16;
  assign f_arrdiv32_out[16] = f_arrdiv32_not15;
  assign f_arrdiv32_out[17] = f_arrdiv32_not14;
  assign f_arrdiv32_out[18] = f_arrdiv32_not13;
  assign f_arrdiv32_out[19] = f_arrdiv32_not12;
  assign f_arrdiv32_out[20] = f_arrdiv32_not11;
  assign f_arrdiv32_out[21] = f_arrdiv32_not10;
  assign f_arrdiv32_out[22] = f_arrdiv32_not9;
  assign f_arrdiv32_out[23] = f_arrdiv32_not8;
  assign f_arrdiv32_out[24] = f_arrdiv32_not7;
  assign f_arrdiv32_out[25] = f_arrdiv32_not6;
  assign f_arrdiv32_out[26] = f_arrdiv32_not5;
  assign f_arrdiv32_out[27] = f_arrdiv32_not4;
  assign f_arrdiv32_out[28] = f_arrdiv32_not3;
  assign f_arrdiv32_out[29] = f_arrdiv32_not2;
  assign f_arrdiv32_out[30] = f_arrdiv32_not1;
  assign f_arrdiv32_out[31] = f_arrdiv32_not0;
endmodule