module f_u_dadda_mul6(input [5:0] a, input [5:0] b, output [11:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire f_u_dadda_mul6_and_4_0_a_4;
  wire f_u_dadda_mul6_and_4_0_b_0;
  wire f_u_dadda_mul6_and_4_0_y0;
  wire f_u_dadda_mul6_and_3_1_a_3;
  wire f_u_dadda_mul6_and_3_1_b_1;
  wire f_u_dadda_mul6_and_3_1_y0;
  wire f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_4_0_y0;
  wire f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_3_1_y0;
  wire f_u_dadda_mul6_ha0_y0;
  wire f_u_dadda_mul6_ha0_y1;
  wire f_u_dadda_mul6_and_5_0_a_5;
  wire f_u_dadda_mul6_and_5_0_b_0;
  wire f_u_dadda_mul6_and_5_0_y0;
  wire f_u_dadda_mul6_and_4_1_a_4;
  wire f_u_dadda_mul6_and_4_1_b_1;
  wire f_u_dadda_mul6_and_4_1_y0;
  wire f_u_dadda_mul6_fa0_f_u_dadda_mul6_ha0_y1;
  wire f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_5_0_y0;
  wire f_u_dadda_mul6_fa0_y0;
  wire f_u_dadda_mul6_fa0_y1;
  wire f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_4_1_y0;
  wire f_u_dadda_mul6_fa0_y2;
  wire f_u_dadda_mul6_fa0_y3;
  wire f_u_dadda_mul6_fa0_y4;
  wire f_u_dadda_mul6_and_3_2_a_3;
  wire f_u_dadda_mul6_and_3_2_b_2;
  wire f_u_dadda_mul6_and_3_2_y0;
  wire f_u_dadda_mul6_and_2_3_a_2;
  wire f_u_dadda_mul6_and_2_3_b_3;
  wire f_u_dadda_mul6_and_2_3_y0;
  wire f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_3_2_y0;
  wire f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_2_3_y0;
  wire f_u_dadda_mul6_ha1_y0;
  wire f_u_dadda_mul6_ha1_y1;
  wire f_u_dadda_mul6_and_5_1_a_5;
  wire f_u_dadda_mul6_and_5_1_b_1;
  wire f_u_dadda_mul6_and_5_1_y0;
  wire f_u_dadda_mul6_fa1_f_u_dadda_mul6_ha1_y1;
  wire f_u_dadda_mul6_fa1_f_u_dadda_mul6_fa0_y4;
  wire f_u_dadda_mul6_fa1_y0;
  wire f_u_dadda_mul6_fa1_y1;
  wire f_u_dadda_mul6_fa1_f_u_dadda_mul6_and_5_1_y0;
  wire f_u_dadda_mul6_fa1_y2;
  wire f_u_dadda_mul6_fa1_y3;
  wire f_u_dadda_mul6_fa1_y4;
  wire f_u_dadda_mul6_and_4_2_a_4;
  wire f_u_dadda_mul6_and_4_2_b_2;
  wire f_u_dadda_mul6_and_4_2_y0;
  wire f_u_dadda_mul6_and_3_3_a_3;
  wire f_u_dadda_mul6_and_3_3_b_3;
  wire f_u_dadda_mul6_and_3_3_y0;
  wire f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_4_2_y0;
  wire f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_3_3_y0;
  wire f_u_dadda_mul6_ha2_y0;
  wire f_u_dadda_mul6_ha2_y1;
  wire f_u_dadda_mul6_and_5_2_a_5;
  wire f_u_dadda_mul6_and_5_2_b_2;
  wire f_u_dadda_mul6_and_5_2_y0;
  wire f_u_dadda_mul6_fa2_f_u_dadda_mul6_ha2_y1;
  wire f_u_dadda_mul6_fa2_f_u_dadda_mul6_fa1_y4;
  wire f_u_dadda_mul6_fa2_y0;
  wire f_u_dadda_mul6_fa2_y1;
  wire f_u_dadda_mul6_fa2_f_u_dadda_mul6_and_5_2_y0;
  wire f_u_dadda_mul6_fa2_y2;
  wire f_u_dadda_mul6_fa2_y3;
  wire f_u_dadda_mul6_fa2_y4;
  wire f_u_dadda_mul6_and_2_0_a_2;
  wire f_u_dadda_mul6_and_2_0_b_0;
  wire f_u_dadda_mul6_and_2_0_y0;
  wire f_u_dadda_mul6_and_1_1_a_1;
  wire f_u_dadda_mul6_and_1_1_b_1;
  wire f_u_dadda_mul6_and_1_1_y0;
  wire f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_2_0_y0;
  wire f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_1_1_y0;
  wire f_u_dadda_mul6_ha3_y0;
  wire f_u_dadda_mul6_ha3_y1;
  wire f_u_dadda_mul6_and_3_0_a_3;
  wire f_u_dadda_mul6_and_3_0_b_0;
  wire f_u_dadda_mul6_and_3_0_y0;
  wire f_u_dadda_mul6_and_2_1_a_2;
  wire f_u_dadda_mul6_and_2_1_b_1;
  wire f_u_dadda_mul6_and_2_1_y0;
  wire f_u_dadda_mul6_fa3_f_u_dadda_mul6_ha3_y1;
  wire f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_3_0_y0;
  wire f_u_dadda_mul6_fa3_y0;
  wire f_u_dadda_mul6_fa3_y1;
  wire f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_2_1_y0;
  wire f_u_dadda_mul6_fa3_y2;
  wire f_u_dadda_mul6_fa3_y3;
  wire f_u_dadda_mul6_fa3_y4;
  wire f_u_dadda_mul6_and_1_2_a_1;
  wire f_u_dadda_mul6_and_1_2_b_2;
  wire f_u_dadda_mul6_and_1_2_y0;
  wire f_u_dadda_mul6_and_0_3_a_0;
  wire f_u_dadda_mul6_and_0_3_b_3;
  wire f_u_dadda_mul6_and_0_3_y0;
  wire f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_1_2_y0;
  wire f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_0_3_y0;
  wire f_u_dadda_mul6_ha4_y0;
  wire f_u_dadda_mul6_ha4_y1;
  wire f_u_dadda_mul6_and_2_2_a_2;
  wire f_u_dadda_mul6_and_2_2_b_2;
  wire f_u_dadda_mul6_and_2_2_y0;
  wire f_u_dadda_mul6_fa4_f_u_dadda_mul6_ha4_y1;
  wire f_u_dadda_mul6_fa4_f_u_dadda_mul6_fa3_y4;
  wire f_u_dadda_mul6_fa4_y0;
  wire f_u_dadda_mul6_fa4_y1;
  wire f_u_dadda_mul6_fa4_f_u_dadda_mul6_and_2_2_y0;
  wire f_u_dadda_mul6_fa4_y2;
  wire f_u_dadda_mul6_fa4_y3;
  wire f_u_dadda_mul6_fa4_y4;
  wire f_u_dadda_mul6_and_1_3_a_1;
  wire f_u_dadda_mul6_and_1_3_b_3;
  wire f_u_dadda_mul6_and_1_3_y0;
  wire f_u_dadda_mul6_and_0_4_a_0;
  wire f_u_dadda_mul6_and_0_4_b_4;
  wire f_u_dadda_mul6_and_0_4_y0;
  wire f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_1_3_y0;
  wire f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_0_4_y0;
  wire f_u_dadda_mul6_fa5_y0;
  wire f_u_dadda_mul6_fa5_y1;
  wire f_u_dadda_mul6_fa5_f_u_dadda_mul6_ha0_y0;
  wire f_u_dadda_mul6_fa5_y2;
  wire f_u_dadda_mul6_fa5_y3;
  wire f_u_dadda_mul6_fa5_y4;
  wire f_u_dadda_mul6_and_1_4_a_1;
  wire f_u_dadda_mul6_and_1_4_b_4;
  wire f_u_dadda_mul6_and_1_4_y0;
  wire f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa5_y4;
  wire f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa4_y4;
  wire f_u_dadda_mul6_fa6_y0;
  wire f_u_dadda_mul6_fa6_y1;
  wire f_u_dadda_mul6_fa6_f_u_dadda_mul6_and_1_4_y0;
  wire f_u_dadda_mul6_fa6_y2;
  wire f_u_dadda_mul6_fa6_y3;
  wire f_u_dadda_mul6_fa6_y4;
  wire f_u_dadda_mul6_and_0_5_a_0;
  wire f_u_dadda_mul6_and_0_5_b_5;
  wire f_u_dadda_mul6_and_0_5_y0;
  wire f_u_dadda_mul6_fa7_f_u_dadda_mul6_and_0_5_y0;
  wire f_u_dadda_mul6_fa7_f_u_dadda_mul6_fa0_y2;
  wire f_u_dadda_mul6_fa7_y0;
  wire f_u_dadda_mul6_fa7_y1;
  wire f_u_dadda_mul6_fa7_f_u_dadda_mul6_ha1_y0;
  wire f_u_dadda_mul6_fa7_y2;
  wire f_u_dadda_mul6_fa7_y3;
  wire f_u_dadda_mul6_fa7_y4;
  wire f_u_dadda_mul6_and_2_4_a_2;
  wire f_u_dadda_mul6_and_2_4_b_4;
  wire f_u_dadda_mul6_and_2_4_y0;
  wire f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa7_y4;
  wire f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa6_y4;
  wire f_u_dadda_mul6_fa8_y0;
  wire f_u_dadda_mul6_fa8_y1;
  wire f_u_dadda_mul6_fa8_f_u_dadda_mul6_and_2_4_y0;
  wire f_u_dadda_mul6_fa8_y2;
  wire f_u_dadda_mul6_fa8_y3;
  wire f_u_dadda_mul6_fa8_y4;
  wire f_u_dadda_mul6_and_1_5_a_1;
  wire f_u_dadda_mul6_and_1_5_b_5;
  wire f_u_dadda_mul6_and_1_5_y0;
  wire f_u_dadda_mul6_fa9_f_u_dadda_mul6_and_1_5_y0;
  wire f_u_dadda_mul6_fa9_f_u_dadda_mul6_fa1_y2;
  wire f_u_dadda_mul6_fa9_y0;
  wire f_u_dadda_mul6_fa9_y1;
  wire f_u_dadda_mul6_fa9_f_u_dadda_mul6_ha2_y0;
  wire f_u_dadda_mul6_fa9_y2;
  wire f_u_dadda_mul6_fa9_y3;
  wire f_u_dadda_mul6_fa9_y4;
  wire f_u_dadda_mul6_and_4_3_a_4;
  wire f_u_dadda_mul6_and_4_3_b_3;
  wire f_u_dadda_mul6_and_4_3_y0;
  wire f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa9_y4;
  wire f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa8_y4;
  wire f_u_dadda_mul6_fa10_y0;
  wire f_u_dadda_mul6_fa10_y1;
  wire f_u_dadda_mul6_fa10_f_u_dadda_mul6_and_4_3_y0;
  wire f_u_dadda_mul6_fa10_y2;
  wire f_u_dadda_mul6_fa10_y3;
  wire f_u_dadda_mul6_fa10_y4;
  wire f_u_dadda_mul6_and_3_4_a_3;
  wire f_u_dadda_mul6_and_3_4_b_4;
  wire f_u_dadda_mul6_and_3_4_y0;
  wire f_u_dadda_mul6_and_2_5_a_2;
  wire f_u_dadda_mul6_and_2_5_b_5;
  wire f_u_dadda_mul6_and_2_5_y0;
  wire f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_3_4_y0;
  wire f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_2_5_y0;
  wire f_u_dadda_mul6_fa11_y0;
  wire f_u_dadda_mul6_fa11_y1;
  wire f_u_dadda_mul6_fa11_f_u_dadda_mul6_fa2_y2;
  wire f_u_dadda_mul6_fa11_y2;
  wire f_u_dadda_mul6_fa11_y3;
  wire f_u_dadda_mul6_fa11_y4;
  wire f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa11_y4;
  wire f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa10_y4;
  wire f_u_dadda_mul6_fa12_y0;
  wire f_u_dadda_mul6_fa12_y1;
  wire f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa2_y4;
  wire f_u_dadda_mul6_fa12_y2;
  wire f_u_dadda_mul6_fa12_y3;
  wire f_u_dadda_mul6_fa12_y4;
  wire f_u_dadda_mul6_and_5_3_a_5;
  wire f_u_dadda_mul6_and_5_3_b_3;
  wire f_u_dadda_mul6_and_5_3_y0;
  wire f_u_dadda_mul6_and_4_4_a_4;
  wire f_u_dadda_mul6_and_4_4_b_4;
  wire f_u_dadda_mul6_and_4_4_y0;
  wire f_u_dadda_mul6_and_3_5_a_3;
  wire f_u_dadda_mul6_and_3_5_b_5;
  wire f_u_dadda_mul6_and_3_5_y0;
  wire f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_5_3_y0;
  wire f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_4_4_y0;
  wire f_u_dadda_mul6_fa13_y0;
  wire f_u_dadda_mul6_fa13_y1;
  wire f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_3_5_y0;
  wire f_u_dadda_mul6_fa13_y2;
  wire f_u_dadda_mul6_fa13_y3;
  wire f_u_dadda_mul6_fa13_y4;
  wire f_u_dadda_mul6_and_5_4_a_5;
  wire f_u_dadda_mul6_and_5_4_b_4;
  wire f_u_dadda_mul6_and_5_4_y0;
  wire f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa13_y4;
  wire f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa12_y4;
  wire f_u_dadda_mul6_fa14_y0;
  wire f_u_dadda_mul6_fa14_y1;
  wire f_u_dadda_mul6_fa14_f_u_dadda_mul6_and_5_4_y0;
  wire f_u_dadda_mul6_fa14_y2;
  wire f_u_dadda_mul6_fa14_y3;
  wire f_u_dadda_mul6_fa14_y4;
  wire f_u_dadda_mul6_and_0_0_a_0;
  wire f_u_dadda_mul6_and_0_0_b_0;
  wire f_u_dadda_mul6_and_0_0_y0;
  wire f_u_dadda_mul6_and_1_0_a_1;
  wire f_u_dadda_mul6_and_1_0_b_0;
  wire f_u_dadda_mul6_and_1_0_y0;
  wire f_u_dadda_mul6_and_0_2_a_0;
  wire f_u_dadda_mul6_and_0_2_b_2;
  wire f_u_dadda_mul6_and_0_2_y0;
  wire f_u_dadda_mul6_and_4_5_a_4;
  wire f_u_dadda_mul6_and_4_5_b_5;
  wire f_u_dadda_mul6_and_4_5_y0;
  wire f_u_dadda_mul6_and_0_1_a_0;
  wire f_u_dadda_mul6_and_0_1_b_1;
  wire f_u_dadda_mul6_and_0_1_y0;
  wire f_u_dadda_mul6_and_5_5_a_5;
  wire f_u_dadda_mul6_and_5_5_b_5;
  wire f_u_dadda_mul6_and_5_5_y0;
  wire f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_1_0_y0;
  wire f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_0_1_y0;
  wire f_u_dadda_mul6_u_rca10_ha_y0;
  wire f_u_dadda_mul6_u_rca10_ha_y1;
  wire f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_and_0_2_y0;
  wire f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_ha3_y0;
  wire f_u_dadda_mul6_u_rca10_fa1_y0;
  wire f_u_dadda_mul6_u_rca10_fa1_y1;
  wire f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_u_rca10_ha_y1;
  wire f_u_dadda_mul6_u_rca10_fa1_y2;
  wire f_u_dadda_mul6_u_rca10_fa1_y3;
  wire f_u_dadda_mul6_u_rca10_fa1_y4;
  wire f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_fa3_y2;
  wire f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_ha4_y0;
  wire f_u_dadda_mul6_u_rca10_fa2_y0;
  wire f_u_dadda_mul6_u_rca10_fa2_y1;
  wire f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_u_rca10_fa1_y4;
  wire f_u_dadda_mul6_u_rca10_fa2_y2;
  wire f_u_dadda_mul6_u_rca10_fa2_y3;
  wire f_u_dadda_mul6_u_rca10_fa2_y4;
  wire f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa4_y2;
  wire f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa5_y2;
  wire f_u_dadda_mul6_u_rca10_fa3_y0;
  wire f_u_dadda_mul6_u_rca10_fa3_y1;
  wire f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_u_rca10_fa2_y4;
  wire f_u_dadda_mul6_u_rca10_fa3_y2;
  wire f_u_dadda_mul6_u_rca10_fa3_y3;
  wire f_u_dadda_mul6_u_rca10_fa3_y4;
  wire f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa6_y2;
  wire f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa7_y2;
  wire f_u_dadda_mul6_u_rca10_fa4_y0;
  wire f_u_dadda_mul6_u_rca10_fa4_y1;
  wire f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_u_rca10_fa3_y4;
  wire f_u_dadda_mul6_u_rca10_fa4_y2;
  wire f_u_dadda_mul6_u_rca10_fa4_y3;
  wire f_u_dadda_mul6_u_rca10_fa4_y4;
  wire f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa8_y2;
  wire f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa9_y2;
  wire f_u_dadda_mul6_u_rca10_fa5_y0;
  wire f_u_dadda_mul6_u_rca10_fa5_y1;
  wire f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_u_rca10_fa4_y4;
  wire f_u_dadda_mul6_u_rca10_fa5_y2;
  wire f_u_dadda_mul6_u_rca10_fa5_y3;
  wire f_u_dadda_mul6_u_rca10_fa5_y4;
  wire f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa10_y2;
  wire f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa11_y2;
  wire f_u_dadda_mul6_u_rca10_fa6_y0;
  wire f_u_dadda_mul6_u_rca10_fa6_y1;
  wire f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_u_rca10_fa5_y4;
  wire f_u_dadda_mul6_u_rca10_fa6_y2;
  wire f_u_dadda_mul6_u_rca10_fa6_y3;
  wire f_u_dadda_mul6_u_rca10_fa6_y4;
  wire f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa12_y2;
  wire f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa13_y2;
  wire f_u_dadda_mul6_u_rca10_fa7_y0;
  wire f_u_dadda_mul6_u_rca10_fa7_y1;
  wire f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_u_rca10_fa6_y4;
  wire f_u_dadda_mul6_u_rca10_fa7_y2;
  wire f_u_dadda_mul6_u_rca10_fa7_y3;
  wire f_u_dadda_mul6_u_rca10_fa7_y4;
  wire f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_and_4_5_y0;
  wire f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_fa14_y2;
  wire f_u_dadda_mul6_u_rca10_fa8_y0;
  wire f_u_dadda_mul6_u_rca10_fa8_y1;
  wire f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_u_rca10_fa7_y4;
  wire f_u_dadda_mul6_u_rca10_fa8_y2;
  wire f_u_dadda_mul6_u_rca10_fa8_y3;
  wire f_u_dadda_mul6_u_rca10_fa8_y4;
  wire f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_fa14_y4;
  wire f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_and_5_5_y0;
  wire f_u_dadda_mul6_u_rca10_fa9_y0;
  wire f_u_dadda_mul6_u_rca10_fa9_y1;
  wire f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_u_rca10_fa8_y4;
  wire f_u_dadda_mul6_u_rca10_fa9_y2;
  wire f_u_dadda_mul6_u_rca10_fa9_y3;
  wire f_u_dadda_mul6_u_rca10_fa9_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign f_u_dadda_mul6_and_4_0_a_4 = a_4;
  assign f_u_dadda_mul6_and_4_0_b_0 = b_0;
  assign f_u_dadda_mul6_and_4_0_y0 = f_u_dadda_mul6_and_4_0_a_4 & f_u_dadda_mul6_and_4_0_b_0;
  assign f_u_dadda_mul6_and_3_1_a_3 = a_3;
  assign f_u_dadda_mul6_and_3_1_b_1 = b_1;
  assign f_u_dadda_mul6_and_3_1_y0 = f_u_dadda_mul6_and_3_1_a_3 & f_u_dadda_mul6_and_3_1_b_1;
  assign f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_4_0_y0 = f_u_dadda_mul6_and_4_0_y0;
  assign f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_3_1_y0 = f_u_dadda_mul6_and_3_1_y0;
  assign f_u_dadda_mul6_ha0_y0 = f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_4_0_y0 ^ f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_3_1_y0;
  assign f_u_dadda_mul6_ha0_y1 = f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_4_0_y0 & f_u_dadda_mul6_ha0_f_u_dadda_mul6_and_3_1_y0;
  assign f_u_dadda_mul6_and_5_0_a_5 = a_5;
  assign f_u_dadda_mul6_and_5_0_b_0 = b_0;
  assign f_u_dadda_mul6_and_5_0_y0 = f_u_dadda_mul6_and_5_0_a_5 & f_u_dadda_mul6_and_5_0_b_0;
  assign f_u_dadda_mul6_and_4_1_a_4 = a_4;
  assign f_u_dadda_mul6_and_4_1_b_1 = b_1;
  assign f_u_dadda_mul6_and_4_1_y0 = f_u_dadda_mul6_and_4_1_a_4 & f_u_dadda_mul6_and_4_1_b_1;
  assign f_u_dadda_mul6_fa0_f_u_dadda_mul6_ha0_y1 = f_u_dadda_mul6_ha0_y1;
  assign f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_5_0_y0 = f_u_dadda_mul6_and_5_0_y0;
  assign f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_4_1_y0 = f_u_dadda_mul6_and_4_1_y0;
  assign f_u_dadda_mul6_fa0_y0 = f_u_dadda_mul6_fa0_f_u_dadda_mul6_ha0_y1 ^ f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_5_0_y0;
  assign f_u_dadda_mul6_fa0_y1 = f_u_dadda_mul6_fa0_f_u_dadda_mul6_ha0_y1 & f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_5_0_y0;
  assign f_u_dadda_mul6_fa0_y2 = f_u_dadda_mul6_fa0_y0 ^ f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_4_1_y0;
  assign f_u_dadda_mul6_fa0_y3 = f_u_dadda_mul6_fa0_y0 & f_u_dadda_mul6_fa0_f_u_dadda_mul6_and_4_1_y0;
  assign f_u_dadda_mul6_fa0_y4 = f_u_dadda_mul6_fa0_y1 | f_u_dadda_mul6_fa0_y3;
  assign f_u_dadda_mul6_and_3_2_a_3 = a_3;
  assign f_u_dadda_mul6_and_3_2_b_2 = b_2;
  assign f_u_dadda_mul6_and_3_2_y0 = f_u_dadda_mul6_and_3_2_a_3 & f_u_dadda_mul6_and_3_2_b_2;
  assign f_u_dadda_mul6_and_2_3_a_2 = a_2;
  assign f_u_dadda_mul6_and_2_3_b_3 = b_3;
  assign f_u_dadda_mul6_and_2_3_y0 = f_u_dadda_mul6_and_2_3_a_2 & f_u_dadda_mul6_and_2_3_b_3;
  assign f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_3_2_y0 = f_u_dadda_mul6_and_3_2_y0;
  assign f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_2_3_y0 = f_u_dadda_mul6_and_2_3_y0;
  assign f_u_dadda_mul6_ha1_y0 = f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_3_2_y0 ^ f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_2_3_y0;
  assign f_u_dadda_mul6_ha1_y1 = f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_3_2_y0 & f_u_dadda_mul6_ha1_f_u_dadda_mul6_and_2_3_y0;
  assign f_u_dadda_mul6_and_5_1_a_5 = a_5;
  assign f_u_dadda_mul6_and_5_1_b_1 = b_1;
  assign f_u_dadda_mul6_and_5_1_y0 = f_u_dadda_mul6_and_5_1_a_5 & f_u_dadda_mul6_and_5_1_b_1;
  assign f_u_dadda_mul6_fa1_f_u_dadda_mul6_ha1_y1 = f_u_dadda_mul6_ha1_y1;
  assign f_u_dadda_mul6_fa1_f_u_dadda_mul6_fa0_y4 = f_u_dadda_mul6_fa0_y4;
  assign f_u_dadda_mul6_fa1_f_u_dadda_mul6_and_5_1_y0 = f_u_dadda_mul6_and_5_1_y0;
  assign f_u_dadda_mul6_fa1_y0 = f_u_dadda_mul6_fa1_f_u_dadda_mul6_ha1_y1 ^ f_u_dadda_mul6_fa1_f_u_dadda_mul6_fa0_y4;
  assign f_u_dadda_mul6_fa1_y1 = f_u_dadda_mul6_fa1_f_u_dadda_mul6_ha1_y1 & f_u_dadda_mul6_fa1_f_u_dadda_mul6_fa0_y4;
  assign f_u_dadda_mul6_fa1_y2 = f_u_dadda_mul6_fa1_y0 ^ f_u_dadda_mul6_fa1_f_u_dadda_mul6_and_5_1_y0;
  assign f_u_dadda_mul6_fa1_y3 = f_u_dadda_mul6_fa1_y0 & f_u_dadda_mul6_fa1_f_u_dadda_mul6_and_5_1_y0;
  assign f_u_dadda_mul6_fa1_y4 = f_u_dadda_mul6_fa1_y1 | f_u_dadda_mul6_fa1_y3;
  assign f_u_dadda_mul6_and_4_2_a_4 = a_4;
  assign f_u_dadda_mul6_and_4_2_b_2 = b_2;
  assign f_u_dadda_mul6_and_4_2_y0 = f_u_dadda_mul6_and_4_2_a_4 & f_u_dadda_mul6_and_4_2_b_2;
  assign f_u_dadda_mul6_and_3_3_a_3 = a_3;
  assign f_u_dadda_mul6_and_3_3_b_3 = b_3;
  assign f_u_dadda_mul6_and_3_3_y0 = f_u_dadda_mul6_and_3_3_a_3 & f_u_dadda_mul6_and_3_3_b_3;
  assign f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_4_2_y0 = f_u_dadda_mul6_and_4_2_y0;
  assign f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_3_3_y0 = f_u_dadda_mul6_and_3_3_y0;
  assign f_u_dadda_mul6_ha2_y0 = f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_4_2_y0 ^ f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_3_3_y0;
  assign f_u_dadda_mul6_ha2_y1 = f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_4_2_y0 & f_u_dadda_mul6_ha2_f_u_dadda_mul6_and_3_3_y0;
  assign f_u_dadda_mul6_and_5_2_a_5 = a_5;
  assign f_u_dadda_mul6_and_5_2_b_2 = b_2;
  assign f_u_dadda_mul6_and_5_2_y0 = f_u_dadda_mul6_and_5_2_a_5 & f_u_dadda_mul6_and_5_2_b_2;
  assign f_u_dadda_mul6_fa2_f_u_dadda_mul6_ha2_y1 = f_u_dadda_mul6_ha2_y1;
  assign f_u_dadda_mul6_fa2_f_u_dadda_mul6_fa1_y4 = f_u_dadda_mul6_fa1_y4;
  assign f_u_dadda_mul6_fa2_f_u_dadda_mul6_and_5_2_y0 = f_u_dadda_mul6_and_5_2_y0;
  assign f_u_dadda_mul6_fa2_y0 = f_u_dadda_mul6_fa2_f_u_dadda_mul6_ha2_y1 ^ f_u_dadda_mul6_fa2_f_u_dadda_mul6_fa1_y4;
  assign f_u_dadda_mul6_fa2_y1 = f_u_dadda_mul6_fa2_f_u_dadda_mul6_ha2_y1 & f_u_dadda_mul6_fa2_f_u_dadda_mul6_fa1_y4;
  assign f_u_dadda_mul6_fa2_y2 = f_u_dadda_mul6_fa2_y0 ^ f_u_dadda_mul6_fa2_f_u_dadda_mul6_and_5_2_y0;
  assign f_u_dadda_mul6_fa2_y3 = f_u_dadda_mul6_fa2_y0 & f_u_dadda_mul6_fa2_f_u_dadda_mul6_and_5_2_y0;
  assign f_u_dadda_mul6_fa2_y4 = f_u_dadda_mul6_fa2_y1 | f_u_dadda_mul6_fa2_y3;
  assign f_u_dadda_mul6_and_2_0_a_2 = a_2;
  assign f_u_dadda_mul6_and_2_0_b_0 = b_0;
  assign f_u_dadda_mul6_and_2_0_y0 = f_u_dadda_mul6_and_2_0_a_2 & f_u_dadda_mul6_and_2_0_b_0;
  assign f_u_dadda_mul6_and_1_1_a_1 = a_1;
  assign f_u_dadda_mul6_and_1_1_b_1 = b_1;
  assign f_u_dadda_mul6_and_1_1_y0 = f_u_dadda_mul6_and_1_1_a_1 & f_u_dadda_mul6_and_1_1_b_1;
  assign f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_2_0_y0 = f_u_dadda_mul6_and_2_0_y0;
  assign f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_1_1_y0 = f_u_dadda_mul6_and_1_1_y0;
  assign f_u_dadda_mul6_ha3_y0 = f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_2_0_y0 ^ f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_1_1_y0;
  assign f_u_dadda_mul6_ha3_y1 = f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_2_0_y0 & f_u_dadda_mul6_ha3_f_u_dadda_mul6_and_1_1_y0;
  assign f_u_dadda_mul6_and_3_0_a_3 = a_3;
  assign f_u_dadda_mul6_and_3_0_b_0 = b_0;
  assign f_u_dadda_mul6_and_3_0_y0 = f_u_dadda_mul6_and_3_0_a_3 & f_u_dadda_mul6_and_3_0_b_0;
  assign f_u_dadda_mul6_and_2_1_a_2 = a_2;
  assign f_u_dadda_mul6_and_2_1_b_1 = b_1;
  assign f_u_dadda_mul6_and_2_1_y0 = f_u_dadda_mul6_and_2_1_a_2 & f_u_dadda_mul6_and_2_1_b_1;
  assign f_u_dadda_mul6_fa3_f_u_dadda_mul6_ha3_y1 = f_u_dadda_mul6_ha3_y1;
  assign f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_3_0_y0 = f_u_dadda_mul6_and_3_0_y0;
  assign f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_2_1_y0 = f_u_dadda_mul6_and_2_1_y0;
  assign f_u_dadda_mul6_fa3_y0 = f_u_dadda_mul6_fa3_f_u_dadda_mul6_ha3_y1 ^ f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_3_0_y0;
  assign f_u_dadda_mul6_fa3_y1 = f_u_dadda_mul6_fa3_f_u_dadda_mul6_ha3_y1 & f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_3_0_y0;
  assign f_u_dadda_mul6_fa3_y2 = f_u_dadda_mul6_fa3_y0 ^ f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_2_1_y0;
  assign f_u_dadda_mul6_fa3_y3 = f_u_dadda_mul6_fa3_y0 & f_u_dadda_mul6_fa3_f_u_dadda_mul6_and_2_1_y0;
  assign f_u_dadda_mul6_fa3_y4 = f_u_dadda_mul6_fa3_y1 | f_u_dadda_mul6_fa3_y3;
  assign f_u_dadda_mul6_and_1_2_a_1 = a_1;
  assign f_u_dadda_mul6_and_1_2_b_2 = b_2;
  assign f_u_dadda_mul6_and_1_2_y0 = f_u_dadda_mul6_and_1_2_a_1 & f_u_dadda_mul6_and_1_2_b_2;
  assign f_u_dadda_mul6_and_0_3_a_0 = a_0;
  assign f_u_dadda_mul6_and_0_3_b_3 = b_3;
  assign f_u_dadda_mul6_and_0_3_y0 = f_u_dadda_mul6_and_0_3_a_0 & f_u_dadda_mul6_and_0_3_b_3;
  assign f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_1_2_y0 = f_u_dadda_mul6_and_1_2_y0;
  assign f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_0_3_y0 = f_u_dadda_mul6_and_0_3_y0;
  assign f_u_dadda_mul6_ha4_y0 = f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_1_2_y0 ^ f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_0_3_y0;
  assign f_u_dadda_mul6_ha4_y1 = f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_1_2_y0 & f_u_dadda_mul6_ha4_f_u_dadda_mul6_and_0_3_y0;
  assign f_u_dadda_mul6_and_2_2_a_2 = a_2;
  assign f_u_dadda_mul6_and_2_2_b_2 = b_2;
  assign f_u_dadda_mul6_and_2_2_y0 = f_u_dadda_mul6_and_2_2_a_2 & f_u_dadda_mul6_and_2_2_b_2;
  assign f_u_dadda_mul6_fa4_f_u_dadda_mul6_ha4_y1 = f_u_dadda_mul6_ha4_y1;
  assign f_u_dadda_mul6_fa4_f_u_dadda_mul6_fa3_y4 = f_u_dadda_mul6_fa3_y4;
  assign f_u_dadda_mul6_fa4_f_u_dadda_mul6_and_2_2_y0 = f_u_dadda_mul6_and_2_2_y0;
  assign f_u_dadda_mul6_fa4_y0 = f_u_dadda_mul6_fa4_f_u_dadda_mul6_ha4_y1 ^ f_u_dadda_mul6_fa4_f_u_dadda_mul6_fa3_y4;
  assign f_u_dadda_mul6_fa4_y1 = f_u_dadda_mul6_fa4_f_u_dadda_mul6_ha4_y1 & f_u_dadda_mul6_fa4_f_u_dadda_mul6_fa3_y4;
  assign f_u_dadda_mul6_fa4_y2 = f_u_dadda_mul6_fa4_y0 ^ f_u_dadda_mul6_fa4_f_u_dadda_mul6_and_2_2_y0;
  assign f_u_dadda_mul6_fa4_y3 = f_u_dadda_mul6_fa4_y0 & f_u_dadda_mul6_fa4_f_u_dadda_mul6_and_2_2_y0;
  assign f_u_dadda_mul6_fa4_y4 = f_u_dadda_mul6_fa4_y1 | f_u_dadda_mul6_fa4_y3;
  assign f_u_dadda_mul6_and_1_3_a_1 = a_1;
  assign f_u_dadda_mul6_and_1_3_b_3 = b_3;
  assign f_u_dadda_mul6_and_1_3_y0 = f_u_dadda_mul6_and_1_3_a_1 & f_u_dadda_mul6_and_1_3_b_3;
  assign f_u_dadda_mul6_and_0_4_a_0 = a_0;
  assign f_u_dadda_mul6_and_0_4_b_4 = b_4;
  assign f_u_dadda_mul6_and_0_4_y0 = f_u_dadda_mul6_and_0_4_a_0 & f_u_dadda_mul6_and_0_4_b_4;
  assign f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_1_3_y0 = f_u_dadda_mul6_and_1_3_y0;
  assign f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_0_4_y0 = f_u_dadda_mul6_and_0_4_y0;
  assign f_u_dadda_mul6_fa5_f_u_dadda_mul6_ha0_y0 = f_u_dadda_mul6_ha0_y0;
  assign f_u_dadda_mul6_fa5_y0 = f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_1_3_y0 ^ f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_0_4_y0;
  assign f_u_dadda_mul6_fa5_y1 = f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_1_3_y0 & f_u_dadda_mul6_fa5_f_u_dadda_mul6_and_0_4_y0;
  assign f_u_dadda_mul6_fa5_y2 = f_u_dadda_mul6_fa5_y0 ^ f_u_dadda_mul6_fa5_f_u_dadda_mul6_ha0_y0;
  assign f_u_dadda_mul6_fa5_y3 = f_u_dadda_mul6_fa5_y0 & f_u_dadda_mul6_fa5_f_u_dadda_mul6_ha0_y0;
  assign f_u_dadda_mul6_fa5_y4 = f_u_dadda_mul6_fa5_y1 | f_u_dadda_mul6_fa5_y3;
  assign f_u_dadda_mul6_and_1_4_a_1 = a_1;
  assign f_u_dadda_mul6_and_1_4_b_4 = b_4;
  assign f_u_dadda_mul6_and_1_4_y0 = f_u_dadda_mul6_and_1_4_a_1 & f_u_dadda_mul6_and_1_4_b_4;
  assign f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa5_y4 = f_u_dadda_mul6_fa5_y4;
  assign f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa4_y4 = f_u_dadda_mul6_fa4_y4;
  assign f_u_dadda_mul6_fa6_f_u_dadda_mul6_and_1_4_y0 = f_u_dadda_mul6_and_1_4_y0;
  assign f_u_dadda_mul6_fa6_y0 = f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa5_y4 ^ f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa4_y4;
  assign f_u_dadda_mul6_fa6_y1 = f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa5_y4 & f_u_dadda_mul6_fa6_f_u_dadda_mul6_fa4_y4;
  assign f_u_dadda_mul6_fa6_y2 = f_u_dadda_mul6_fa6_y0 ^ f_u_dadda_mul6_fa6_f_u_dadda_mul6_and_1_4_y0;
  assign f_u_dadda_mul6_fa6_y3 = f_u_dadda_mul6_fa6_y0 & f_u_dadda_mul6_fa6_f_u_dadda_mul6_and_1_4_y0;
  assign f_u_dadda_mul6_fa6_y4 = f_u_dadda_mul6_fa6_y1 | f_u_dadda_mul6_fa6_y3;
  assign f_u_dadda_mul6_and_0_5_a_0 = a_0;
  assign f_u_dadda_mul6_and_0_5_b_5 = b_5;
  assign f_u_dadda_mul6_and_0_5_y0 = f_u_dadda_mul6_and_0_5_a_0 & f_u_dadda_mul6_and_0_5_b_5;
  assign f_u_dadda_mul6_fa7_f_u_dadda_mul6_and_0_5_y0 = f_u_dadda_mul6_and_0_5_y0;
  assign f_u_dadda_mul6_fa7_f_u_dadda_mul6_fa0_y2 = f_u_dadda_mul6_fa0_y2;
  assign f_u_dadda_mul6_fa7_f_u_dadda_mul6_ha1_y0 = f_u_dadda_mul6_ha1_y0;
  assign f_u_dadda_mul6_fa7_y0 = f_u_dadda_mul6_fa7_f_u_dadda_mul6_and_0_5_y0 ^ f_u_dadda_mul6_fa7_f_u_dadda_mul6_fa0_y2;
  assign f_u_dadda_mul6_fa7_y1 = f_u_dadda_mul6_fa7_f_u_dadda_mul6_and_0_5_y0 & f_u_dadda_mul6_fa7_f_u_dadda_mul6_fa0_y2;
  assign f_u_dadda_mul6_fa7_y2 = f_u_dadda_mul6_fa7_y0 ^ f_u_dadda_mul6_fa7_f_u_dadda_mul6_ha1_y0;
  assign f_u_dadda_mul6_fa7_y3 = f_u_dadda_mul6_fa7_y0 & f_u_dadda_mul6_fa7_f_u_dadda_mul6_ha1_y0;
  assign f_u_dadda_mul6_fa7_y4 = f_u_dadda_mul6_fa7_y1 | f_u_dadda_mul6_fa7_y3;
  assign f_u_dadda_mul6_and_2_4_a_2 = a_2;
  assign f_u_dadda_mul6_and_2_4_b_4 = b_4;
  assign f_u_dadda_mul6_and_2_4_y0 = f_u_dadda_mul6_and_2_4_a_2 & f_u_dadda_mul6_and_2_4_b_4;
  assign f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa7_y4 = f_u_dadda_mul6_fa7_y4;
  assign f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa6_y4 = f_u_dadda_mul6_fa6_y4;
  assign f_u_dadda_mul6_fa8_f_u_dadda_mul6_and_2_4_y0 = f_u_dadda_mul6_and_2_4_y0;
  assign f_u_dadda_mul6_fa8_y0 = f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa7_y4 ^ f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa6_y4;
  assign f_u_dadda_mul6_fa8_y1 = f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa7_y4 & f_u_dadda_mul6_fa8_f_u_dadda_mul6_fa6_y4;
  assign f_u_dadda_mul6_fa8_y2 = f_u_dadda_mul6_fa8_y0 ^ f_u_dadda_mul6_fa8_f_u_dadda_mul6_and_2_4_y0;
  assign f_u_dadda_mul6_fa8_y3 = f_u_dadda_mul6_fa8_y0 & f_u_dadda_mul6_fa8_f_u_dadda_mul6_and_2_4_y0;
  assign f_u_dadda_mul6_fa8_y4 = f_u_dadda_mul6_fa8_y1 | f_u_dadda_mul6_fa8_y3;
  assign f_u_dadda_mul6_and_1_5_a_1 = a_1;
  assign f_u_dadda_mul6_and_1_5_b_5 = b_5;
  assign f_u_dadda_mul6_and_1_5_y0 = f_u_dadda_mul6_and_1_5_a_1 & f_u_dadda_mul6_and_1_5_b_5;
  assign f_u_dadda_mul6_fa9_f_u_dadda_mul6_and_1_5_y0 = f_u_dadda_mul6_and_1_5_y0;
  assign f_u_dadda_mul6_fa9_f_u_dadda_mul6_fa1_y2 = f_u_dadda_mul6_fa1_y2;
  assign f_u_dadda_mul6_fa9_f_u_dadda_mul6_ha2_y0 = f_u_dadda_mul6_ha2_y0;
  assign f_u_dadda_mul6_fa9_y0 = f_u_dadda_mul6_fa9_f_u_dadda_mul6_and_1_5_y0 ^ f_u_dadda_mul6_fa9_f_u_dadda_mul6_fa1_y2;
  assign f_u_dadda_mul6_fa9_y1 = f_u_dadda_mul6_fa9_f_u_dadda_mul6_and_1_5_y0 & f_u_dadda_mul6_fa9_f_u_dadda_mul6_fa1_y2;
  assign f_u_dadda_mul6_fa9_y2 = f_u_dadda_mul6_fa9_y0 ^ f_u_dadda_mul6_fa9_f_u_dadda_mul6_ha2_y0;
  assign f_u_dadda_mul6_fa9_y3 = f_u_dadda_mul6_fa9_y0 & f_u_dadda_mul6_fa9_f_u_dadda_mul6_ha2_y0;
  assign f_u_dadda_mul6_fa9_y4 = f_u_dadda_mul6_fa9_y1 | f_u_dadda_mul6_fa9_y3;
  assign f_u_dadda_mul6_and_4_3_a_4 = a_4;
  assign f_u_dadda_mul6_and_4_3_b_3 = b_3;
  assign f_u_dadda_mul6_and_4_3_y0 = f_u_dadda_mul6_and_4_3_a_4 & f_u_dadda_mul6_and_4_3_b_3;
  assign f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa9_y4 = f_u_dadda_mul6_fa9_y4;
  assign f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa8_y4 = f_u_dadda_mul6_fa8_y4;
  assign f_u_dadda_mul6_fa10_f_u_dadda_mul6_and_4_3_y0 = f_u_dadda_mul6_and_4_3_y0;
  assign f_u_dadda_mul6_fa10_y0 = f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa9_y4 ^ f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa8_y4;
  assign f_u_dadda_mul6_fa10_y1 = f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa9_y4 & f_u_dadda_mul6_fa10_f_u_dadda_mul6_fa8_y4;
  assign f_u_dadda_mul6_fa10_y2 = f_u_dadda_mul6_fa10_y0 ^ f_u_dadda_mul6_fa10_f_u_dadda_mul6_and_4_3_y0;
  assign f_u_dadda_mul6_fa10_y3 = f_u_dadda_mul6_fa10_y0 & f_u_dadda_mul6_fa10_f_u_dadda_mul6_and_4_3_y0;
  assign f_u_dadda_mul6_fa10_y4 = f_u_dadda_mul6_fa10_y1 | f_u_dadda_mul6_fa10_y3;
  assign f_u_dadda_mul6_and_3_4_a_3 = a_3;
  assign f_u_dadda_mul6_and_3_4_b_4 = b_4;
  assign f_u_dadda_mul6_and_3_4_y0 = f_u_dadda_mul6_and_3_4_a_3 & f_u_dadda_mul6_and_3_4_b_4;
  assign f_u_dadda_mul6_and_2_5_a_2 = a_2;
  assign f_u_dadda_mul6_and_2_5_b_5 = b_5;
  assign f_u_dadda_mul6_and_2_5_y0 = f_u_dadda_mul6_and_2_5_a_2 & f_u_dadda_mul6_and_2_5_b_5;
  assign f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_3_4_y0 = f_u_dadda_mul6_and_3_4_y0;
  assign f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_2_5_y0 = f_u_dadda_mul6_and_2_5_y0;
  assign f_u_dadda_mul6_fa11_f_u_dadda_mul6_fa2_y2 = f_u_dadda_mul6_fa2_y2;
  assign f_u_dadda_mul6_fa11_y0 = f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_3_4_y0 ^ f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_2_5_y0;
  assign f_u_dadda_mul6_fa11_y1 = f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_3_4_y0 & f_u_dadda_mul6_fa11_f_u_dadda_mul6_and_2_5_y0;
  assign f_u_dadda_mul6_fa11_y2 = f_u_dadda_mul6_fa11_y0 ^ f_u_dadda_mul6_fa11_f_u_dadda_mul6_fa2_y2;
  assign f_u_dadda_mul6_fa11_y3 = f_u_dadda_mul6_fa11_y0 & f_u_dadda_mul6_fa11_f_u_dadda_mul6_fa2_y2;
  assign f_u_dadda_mul6_fa11_y4 = f_u_dadda_mul6_fa11_y1 | f_u_dadda_mul6_fa11_y3;
  assign f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa11_y4 = f_u_dadda_mul6_fa11_y4;
  assign f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa10_y4 = f_u_dadda_mul6_fa10_y4;
  assign f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa2_y4 = f_u_dadda_mul6_fa2_y4;
  assign f_u_dadda_mul6_fa12_y0 = f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa11_y4 ^ f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa10_y4;
  assign f_u_dadda_mul6_fa12_y1 = f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa11_y4 & f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa10_y4;
  assign f_u_dadda_mul6_fa12_y2 = f_u_dadda_mul6_fa12_y0 ^ f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa2_y4;
  assign f_u_dadda_mul6_fa12_y3 = f_u_dadda_mul6_fa12_y0 & f_u_dadda_mul6_fa12_f_u_dadda_mul6_fa2_y4;
  assign f_u_dadda_mul6_fa12_y4 = f_u_dadda_mul6_fa12_y1 | f_u_dadda_mul6_fa12_y3;
  assign f_u_dadda_mul6_and_5_3_a_5 = a_5;
  assign f_u_dadda_mul6_and_5_3_b_3 = b_3;
  assign f_u_dadda_mul6_and_5_3_y0 = f_u_dadda_mul6_and_5_3_a_5 & f_u_dadda_mul6_and_5_3_b_3;
  assign f_u_dadda_mul6_and_4_4_a_4 = a_4;
  assign f_u_dadda_mul6_and_4_4_b_4 = b_4;
  assign f_u_dadda_mul6_and_4_4_y0 = f_u_dadda_mul6_and_4_4_a_4 & f_u_dadda_mul6_and_4_4_b_4;
  assign f_u_dadda_mul6_and_3_5_a_3 = a_3;
  assign f_u_dadda_mul6_and_3_5_b_5 = b_5;
  assign f_u_dadda_mul6_and_3_5_y0 = f_u_dadda_mul6_and_3_5_a_3 & f_u_dadda_mul6_and_3_5_b_5;
  assign f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_5_3_y0 = f_u_dadda_mul6_and_5_3_y0;
  assign f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_4_4_y0 = f_u_dadda_mul6_and_4_4_y0;
  assign f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_3_5_y0 = f_u_dadda_mul6_and_3_5_y0;
  assign f_u_dadda_mul6_fa13_y0 = f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_5_3_y0 ^ f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_4_4_y0;
  assign f_u_dadda_mul6_fa13_y1 = f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_5_3_y0 & f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_4_4_y0;
  assign f_u_dadda_mul6_fa13_y2 = f_u_dadda_mul6_fa13_y0 ^ f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_3_5_y0;
  assign f_u_dadda_mul6_fa13_y3 = f_u_dadda_mul6_fa13_y0 & f_u_dadda_mul6_fa13_f_u_dadda_mul6_and_3_5_y0;
  assign f_u_dadda_mul6_fa13_y4 = f_u_dadda_mul6_fa13_y1 | f_u_dadda_mul6_fa13_y3;
  assign f_u_dadda_mul6_and_5_4_a_5 = a_5;
  assign f_u_dadda_mul6_and_5_4_b_4 = b_4;
  assign f_u_dadda_mul6_and_5_4_y0 = f_u_dadda_mul6_and_5_4_a_5 & f_u_dadda_mul6_and_5_4_b_4;
  assign f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa13_y4 = f_u_dadda_mul6_fa13_y4;
  assign f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa12_y4 = f_u_dadda_mul6_fa12_y4;
  assign f_u_dadda_mul6_fa14_f_u_dadda_mul6_and_5_4_y0 = f_u_dadda_mul6_and_5_4_y0;
  assign f_u_dadda_mul6_fa14_y0 = f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa13_y4 ^ f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa12_y4;
  assign f_u_dadda_mul6_fa14_y1 = f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa13_y4 & f_u_dadda_mul6_fa14_f_u_dadda_mul6_fa12_y4;
  assign f_u_dadda_mul6_fa14_y2 = f_u_dadda_mul6_fa14_y0 ^ f_u_dadda_mul6_fa14_f_u_dadda_mul6_and_5_4_y0;
  assign f_u_dadda_mul6_fa14_y3 = f_u_dadda_mul6_fa14_y0 & f_u_dadda_mul6_fa14_f_u_dadda_mul6_and_5_4_y0;
  assign f_u_dadda_mul6_fa14_y4 = f_u_dadda_mul6_fa14_y1 | f_u_dadda_mul6_fa14_y3;
  assign f_u_dadda_mul6_and_0_0_a_0 = a_0;
  assign f_u_dadda_mul6_and_0_0_b_0 = b_0;
  assign f_u_dadda_mul6_and_0_0_y0 = f_u_dadda_mul6_and_0_0_a_0 & f_u_dadda_mul6_and_0_0_b_0;
  assign f_u_dadda_mul6_and_1_0_a_1 = a_1;
  assign f_u_dadda_mul6_and_1_0_b_0 = b_0;
  assign f_u_dadda_mul6_and_1_0_y0 = f_u_dadda_mul6_and_1_0_a_1 & f_u_dadda_mul6_and_1_0_b_0;
  assign f_u_dadda_mul6_and_0_2_a_0 = a_0;
  assign f_u_dadda_mul6_and_0_2_b_2 = b_2;
  assign f_u_dadda_mul6_and_0_2_y0 = f_u_dadda_mul6_and_0_2_a_0 & f_u_dadda_mul6_and_0_2_b_2;
  assign f_u_dadda_mul6_and_4_5_a_4 = a_4;
  assign f_u_dadda_mul6_and_4_5_b_5 = b_5;
  assign f_u_dadda_mul6_and_4_5_y0 = f_u_dadda_mul6_and_4_5_a_4 & f_u_dadda_mul6_and_4_5_b_5;
  assign f_u_dadda_mul6_and_0_1_a_0 = a_0;
  assign f_u_dadda_mul6_and_0_1_b_1 = b_1;
  assign f_u_dadda_mul6_and_0_1_y0 = f_u_dadda_mul6_and_0_1_a_0 & f_u_dadda_mul6_and_0_1_b_1;
  assign f_u_dadda_mul6_and_5_5_a_5 = a_5;
  assign f_u_dadda_mul6_and_5_5_b_5 = b_5;
  assign f_u_dadda_mul6_and_5_5_y0 = f_u_dadda_mul6_and_5_5_a_5 & f_u_dadda_mul6_and_5_5_b_5;
  assign f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_1_0_y0 = f_u_dadda_mul6_and_1_0_y0;
  assign f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_0_1_y0 = f_u_dadda_mul6_and_0_1_y0;
  assign f_u_dadda_mul6_u_rca10_ha_y0 = f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_1_0_y0 ^ f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_0_1_y0;
  assign f_u_dadda_mul6_u_rca10_ha_y1 = f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_1_0_y0 & f_u_dadda_mul6_u_rca10_ha_f_u_dadda_mul6_and_0_1_y0;
  assign f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_and_0_2_y0 = f_u_dadda_mul6_and_0_2_y0;
  assign f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_ha3_y0 = f_u_dadda_mul6_ha3_y0;
  assign f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_u_rca10_ha_y1 = f_u_dadda_mul6_u_rca10_ha_y1;
  assign f_u_dadda_mul6_u_rca10_fa1_y0 = f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_and_0_2_y0 ^ f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_ha3_y0;
  assign f_u_dadda_mul6_u_rca10_fa1_y1 = f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_and_0_2_y0 & f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_ha3_y0;
  assign f_u_dadda_mul6_u_rca10_fa1_y2 = f_u_dadda_mul6_u_rca10_fa1_y0 ^ f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_u_rca10_ha_y1;
  assign f_u_dadda_mul6_u_rca10_fa1_y3 = f_u_dadda_mul6_u_rca10_fa1_y0 & f_u_dadda_mul6_u_rca10_fa1_f_u_dadda_mul6_u_rca10_ha_y1;
  assign f_u_dadda_mul6_u_rca10_fa1_y4 = f_u_dadda_mul6_u_rca10_fa1_y1 | f_u_dadda_mul6_u_rca10_fa1_y3;
  assign f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_fa3_y2 = f_u_dadda_mul6_fa3_y2;
  assign f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_ha4_y0 = f_u_dadda_mul6_ha4_y0;
  assign f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_u_rca10_fa1_y4 = f_u_dadda_mul6_u_rca10_fa1_y4;
  assign f_u_dadda_mul6_u_rca10_fa2_y0 = f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_fa3_y2 ^ f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_ha4_y0;
  assign f_u_dadda_mul6_u_rca10_fa2_y1 = f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_fa3_y2 & f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_ha4_y0;
  assign f_u_dadda_mul6_u_rca10_fa2_y2 = f_u_dadda_mul6_u_rca10_fa2_y0 ^ f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_u_rca10_fa1_y4;
  assign f_u_dadda_mul6_u_rca10_fa2_y3 = f_u_dadda_mul6_u_rca10_fa2_y0 & f_u_dadda_mul6_u_rca10_fa2_f_u_dadda_mul6_u_rca10_fa1_y4;
  assign f_u_dadda_mul6_u_rca10_fa2_y4 = f_u_dadda_mul6_u_rca10_fa2_y1 | f_u_dadda_mul6_u_rca10_fa2_y3;
  assign f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa4_y2 = f_u_dadda_mul6_fa4_y2;
  assign f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa5_y2 = f_u_dadda_mul6_fa5_y2;
  assign f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_u_rca10_fa2_y4 = f_u_dadda_mul6_u_rca10_fa2_y4;
  assign f_u_dadda_mul6_u_rca10_fa3_y0 = f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa4_y2 ^ f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa5_y2;
  assign f_u_dadda_mul6_u_rca10_fa3_y1 = f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa4_y2 & f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_fa5_y2;
  assign f_u_dadda_mul6_u_rca10_fa3_y2 = f_u_dadda_mul6_u_rca10_fa3_y0 ^ f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_u_rca10_fa2_y4;
  assign f_u_dadda_mul6_u_rca10_fa3_y3 = f_u_dadda_mul6_u_rca10_fa3_y0 & f_u_dadda_mul6_u_rca10_fa3_f_u_dadda_mul6_u_rca10_fa2_y4;
  assign f_u_dadda_mul6_u_rca10_fa3_y4 = f_u_dadda_mul6_u_rca10_fa3_y1 | f_u_dadda_mul6_u_rca10_fa3_y3;
  assign f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa6_y2 = f_u_dadda_mul6_fa6_y2;
  assign f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa7_y2 = f_u_dadda_mul6_fa7_y2;
  assign f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_u_rca10_fa3_y4 = f_u_dadda_mul6_u_rca10_fa3_y4;
  assign f_u_dadda_mul6_u_rca10_fa4_y0 = f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa6_y2 ^ f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa7_y2;
  assign f_u_dadda_mul6_u_rca10_fa4_y1 = f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa6_y2 & f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_fa7_y2;
  assign f_u_dadda_mul6_u_rca10_fa4_y2 = f_u_dadda_mul6_u_rca10_fa4_y0 ^ f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_u_rca10_fa3_y4;
  assign f_u_dadda_mul6_u_rca10_fa4_y3 = f_u_dadda_mul6_u_rca10_fa4_y0 & f_u_dadda_mul6_u_rca10_fa4_f_u_dadda_mul6_u_rca10_fa3_y4;
  assign f_u_dadda_mul6_u_rca10_fa4_y4 = f_u_dadda_mul6_u_rca10_fa4_y1 | f_u_dadda_mul6_u_rca10_fa4_y3;
  assign f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa8_y2 = f_u_dadda_mul6_fa8_y2;
  assign f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa9_y2 = f_u_dadda_mul6_fa9_y2;
  assign f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_u_rca10_fa4_y4 = f_u_dadda_mul6_u_rca10_fa4_y4;
  assign f_u_dadda_mul6_u_rca10_fa5_y0 = f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa8_y2 ^ f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa9_y2;
  assign f_u_dadda_mul6_u_rca10_fa5_y1 = f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa8_y2 & f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_fa9_y2;
  assign f_u_dadda_mul6_u_rca10_fa5_y2 = f_u_dadda_mul6_u_rca10_fa5_y0 ^ f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_u_rca10_fa4_y4;
  assign f_u_dadda_mul6_u_rca10_fa5_y3 = f_u_dadda_mul6_u_rca10_fa5_y0 & f_u_dadda_mul6_u_rca10_fa5_f_u_dadda_mul6_u_rca10_fa4_y4;
  assign f_u_dadda_mul6_u_rca10_fa5_y4 = f_u_dadda_mul6_u_rca10_fa5_y1 | f_u_dadda_mul6_u_rca10_fa5_y3;
  assign f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa10_y2 = f_u_dadda_mul6_fa10_y2;
  assign f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa11_y2 = f_u_dadda_mul6_fa11_y2;
  assign f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_u_rca10_fa5_y4 = f_u_dadda_mul6_u_rca10_fa5_y4;
  assign f_u_dadda_mul6_u_rca10_fa6_y0 = f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa10_y2 ^ f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa11_y2;
  assign f_u_dadda_mul6_u_rca10_fa6_y1 = f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa10_y2 & f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_fa11_y2;
  assign f_u_dadda_mul6_u_rca10_fa6_y2 = f_u_dadda_mul6_u_rca10_fa6_y0 ^ f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_u_rca10_fa5_y4;
  assign f_u_dadda_mul6_u_rca10_fa6_y3 = f_u_dadda_mul6_u_rca10_fa6_y0 & f_u_dadda_mul6_u_rca10_fa6_f_u_dadda_mul6_u_rca10_fa5_y4;
  assign f_u_dadda_mul6_u_rca10_fa6_y4 = f_u_dadda_mul6_u_rca10_fa6_y1 | f_u_dadda_mul6_u_rca10_fa6_y3;
  assign f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa12_y2 = f_u_dadda_mul6_fa12_y2;
  assign f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa13_y2 = f_u_dadda_mul6_fa13_y2;
  assign f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_u_rca10_fa6_y4 = f_u_dadda_mul6_u_rca10_fa6_y4;
  assign f_u_dadda_mul6_u_rca10_fa7_y0 = f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa12_y2 ^ f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa13_y2;
  assign f_u_dadda_mul6_u_rca10_fa7_y1 = f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa12_y2 & f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_fa13_y2;
  assign f_u_dadda_mul6_u_rca10_fa7_y2 = f_u_dadda_mul6_u_rca10_fa7_y0 ^ f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_u_rca10_fa6_y4;
  assign f_u_dadda_mul6_u_rca10_fa7_y3 = f_u_dadda_mul6_u_rca10_fa7_y0 & f_u_dadda_mul6_u_rca10_fa7_f_u_dadda_mul6_u_rca10_fa6_y4;
  assign f_u_dadda_mul6_u_rca10_fa7_y4 = f_u_dadda_mul6_u_rca10_fa7_y1 | f_u_dadda_mul6_u_rca10_fa7_y3;
  assign f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_and_4_5_y0 = f_u_dadda_mul6_and_4_5_y0;
  assign f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_fa14_y2 = f_u_dadda_mul6_fa14_y2;
  assign f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_u_rca10_fa7_y4 = f_u_dadda_mul6_u_rca10_fa7_y4;
  assign f_u_dadda_mul6_u_rca10_fa8_y0 = f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_and_4_5_y0 ^ f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_fa14_y2;
  assign f_u_dadda_mul6_u_rca10_fa8_y1 = f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_and_4_5_y0 & f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_fa14_y2;
  assign f_u_dadda_mul6_u_rca10_fa8_y2 = f_u_dadda_mul6_u_rca10_fa8_y0 ^ f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_u_rca10_fa7_y4;
  assign f_u_dadda_mul6_u_rca10_fa8_y3 = f_u_dadda_mul6_u_rca10_fa8_y0 & f_u_dadda_mul6_u_rca10_fa8_f_u_dadda_mul6_u_rca10_fa7_y4;
  assign f_u_dadda_mul6_u_rca10_fa8_y4 = f_u_dadda_mul6_u_rca10_fa8_y1 | f_u_dadda_mul6_u_rca10_fa8_y3;
  assign f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_fa14_y4 = f_u_dadda_mul6_fa14_y4;
  assign f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_and_5_5_y0 = f_u_dadda_mul6_and_5_5_y0;
  assign f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_u_rca10_fa8_y4 = f_u_dadda_mul6_u_rca10_fa8_y4;
  assign f_u_dadda_mul6_u_rca10_fa9_y0 = f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_fa14_y4 ^ f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_and_5_5_y0;
  assign f_u_dadda_mul6_u_rca10_fa9_y1 = f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_fa14_y4 & f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_and_5_5_y0;
  assign f_u_dadda_mul6_u_rca10_fa9_y2 = f_u_dadda_mul6_u_rca10_fa9_y0 ^ f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_u_rca10_fa8_y4;
  assign f_u_dadda_mul6_u_rca10_fa9_y3 = f_u_dadda_mul6_u_rca10_fa9_y0 & f_u_dadda_mul6_u_rca10_fa9_f_u_dadda_mul6_u_rca10_fa8_y4;
  assign f_u_dadda_mul6_u_rca10_fa9_y4 = f_u_dadda_mul6_u_rca10_fa9_y1 | f_u_dadda_mul6_u_rca10_fa9_y3;


  assign out[0] = f_u_dadda_mul6_and_0_0_y0;
  assign out[1] = f_u_dadda_mul6_u_rca10_ha_y0;
  assign out[2] = f_u_dadda_mul6_u_rca10_fa1_y2;
  assign out[3] = f_u_dadda_mul6_u_rca10_fa2_y2;
  assign out[4] = f_u_dadda_mul6_u_rca10_fa3_y2;
  assign out[5] = f_u_dadda_mul6_u_rca10_fa4_y2;
  assign out[6] = f_u_dadda_mul6_u_rca10_fa5_y2;
  assign out[7] = f_u_dadda_mul6_u_rca10_fa6_y2;
  assign out[8] = f_u_dadda_mul6_u_rca10_fa7_y2;
  assign out[9] = f_u_dadda_mul6_u_rca10_fa8_y2;
  assign out[10] = f_u_dadda_mul6_u_rca10_fa9_y2;
  assign out[11] = f_u_dadda_mul6_u_rca10_fa9_y4;
endmodule