module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fs(input [0:0] a, input [0:0] b, input [0:0] bin, output [0:0] fs_xor1, output [0:0] fs_or0);
  wire [0:0] fs_xor0;
  wire [0:0] fs_not0;
  wire [0:0] fs_and0;
  wire [0:0] fs_not1;
  wire [0:0] fs_and1;
  xor_gate xor_gate_fs_xor0(.a(a[0]), .b(b[0]), .out(fs_xor0));
  not_gate not_gate_fs_not0(.a(a[0]), .out(fs_not0));
  and_gate and_gate_fs_and0(.a(fs_not0[0]), .b(b[0]), .out(fs_and0));
  xor_gate xor_gate_fs_xor1(.a(bin[0]), .b(fs_xor0[0]), .out(fs_xor1));
  not_gate not_gate_fs_not1(.a(fs_xor0[0]), .out(fs_not1));
  and_gate and_gate_fs_and1(.a(fs_not1[0]), .b(bin[0]), .out(fs_and1));
  or_gate or_gate_fs_or0(.a(fs_and1[0]), .b(fs_and0[0]), .out(fs_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module h_arrdiv24(input [23:0] a, input [23:0] b, output [23:0] h_arrdiv24_out);
  wire [0:0] h_arrdiv24_fs0_xor0;
  wire [0:0] h_arrdiv24_fs0_and0;
  wire [0:0] h_arrdiv24_fs1_xor1;
  wire [0:0] h_arrdiv24_fs1_or0;
  wire [0:0] h_arrdiv24_fs2_xor1;
  wire [0:0] h_arrdiv24_fs2_or0;
  wire [0:0] h_arrdiv24_fs3_xor1;
  wire [0:0] h_arrdiv24_fs3_or0;
  wire [0:0] h_arrdiv24_fs4_xor1;
  wire [0:0] h_arrdiv24_fs4_or0;
  wire [0:0] h_arrdiv24_fs5_xor1;
  wire [0:0] h_arrdiv24_fs5_or0;
  wire [0:0] h_arrdiv24_fs6_xor1;
  wire [0:0] h_arrdiv24_fs6_or0;
  wire [0:0] h_arrdiv24_fs7_xor1;
  wire [0:0] h_arrdiv24_fs7_or0;
  wire [0:0] h_arrdiv24_fs8_xor1;
  wire [0:0] h_arrdiv24_fs8_or0;
  wire [0:0] h_arrdiv24_fs9_xor1;
  wire [0:0] h_arrdiv24_fs9_or0;
  wire [0:0] h_arrdiv24_fs10_xor1;
  wire [0:0] h_arrdiv24_fs10_or0;
  wire [0:0] h_arrdiv24_fs11_xor1;
  wire [0:0] h_arrdiv24_fs11_or0;
  wire [0:0] h_arrdiv24_fs12_xor1;
  wire [0:0] h_arrdiv24_fs12_or0;
  wire [0:0] h_arrdiv24_fs13_xor1;
  wire [0:0] h_arrdiv24_fs13_or0;
  wire [0:0] h_arrdiv24_fs14_xor1;
  wire [0:0] h_arrdiv24_fs14_or0;
  wire [0:0] h_arrdiv24_fs15_xor1;
  wire [0:0] h_arrdiv24_fs15_or0;
  wire [0:0] h_arrdiv24_fs16_xor1;
  wire [0:0] h_arrdiv24_fs16_or0;
  wire [0:0] h_arrdiv24_fs17_xor1;
  wire [0:0] h_arrdiv24_fs17_or0;
  wire [0:0] h_arrdiv24_fs18_xor1;
  wire [0:0] h_arrdiv24_fs18_or0;
  wire [0:0] h_arrdiv24_fs19_xor1;
  wire [0:0] h_arrdiv24_fs19_or0;
  wire [0:0] h_arrdiv24_fs20_xor1;
  wire [0:0] h_arrdiv24_fs20_or0;
  wire [0:0] h_arrdiv24_fs21_xor1;
  wire [0:0] h_arrdiv24_fs21_or0;
  wire [0:0] h_arrdiv24_fs22_xor1;
  wire [0:0] h_arrdiv24_fs22_or0;
  wire [0:0] h_arrdiv24_fs23_xor1;
  wire [0:0] h_arrdiv24_fs23_or0;
  wire [0:0] h_arrdiv24_mux2to10_xor0;
  wire [0:0] h_arrdiv24_mux2to11_and1;
  wire [0:0] h_arrdiv24_mux2to12_and1;
  wire [0:0] h_arrdiv24_mux2to13_and1;
  wire [0:0] h_arrdiv24_mux2to14_and1;
  wire [0:0] h_arrdiv24_mux2to15_and1;
  wire [0:0] h_arrdiv24_mux2to16_and1;
  wire [0:0] h_arrdiv24_mux2to17_and1;
  wire [0:0] h_arrdiv24_mux2to18_and1;
  wire [0:0] h_arrdiv24_mux2to19_and1;
  wire [0:0] h_arrdiv24_mux2to110_and1;
  wire [0:0] h_arrdiv24_mux2to111_and1;
  wire [0:0] h_arrdiv24_mux2to112_and1;
  wire [0:0] h_arrdiv24_mux2to113_and1;
  wire [0:0] h_arrdiv24_mux2to114_and1;
  wire [0:0] h_arrdiv24_mux2to115_and1;
  wire [0:0] h_arrdiv24_mux2to116_and1;
  wire [0:0] h_arrdiv24_mux2to117_and1;
  wire [0:0] h_arrdiv24_mux2to118_and1;
  wire [0:0] h_arrdiv24_mux2to119_and1;
  wire [0:0] h_arrdiv24_mux2to120_and1;
  wire [0:0] h_arrdiv24_mux2to121_and1;
  wire [0:0] h_arrdiv24_mux2to122_and1;
  wire [0:0] h_arrdiv24_not0;
  wire [0:0] h_arrdiv24_fs24_xor0;
  wire [0:0] h_arrdiv24_fs24_and0;
  wire [0:0] h_arrdiv24_fs25_xor1;
  wire [0:0] h_arrdiv24_fs25_or0;
  wire [0:0] h_arrdiv24_fs26_xor1;
  wire [0:0] h_arrdiv24_fs26_or0;
  wire [0:0] h_arrdiv24_fs27_xor1;
  wire [0:0] h_arrdiv24_fs27_or0;
  wire [0:0] h_arrdiv24_fs28_xor1;
  wire [0:0] h_arrdiv24_fs28_or0;
  wire [0:0] h_arrdiv24_fs29_xor1;
  wire [0:0] h_arrdiv24_fs29_or0;
  wire [0:0] h_arrdiv24_fs30_xor1;
  wire [0:0] h_arrdiv24_fs30_or0;
  wire [0:0] h_arrdiv24_fs31_xor1;
  wire [0:0] h_arrdiv24_fs31_or0;
  wire [0:0] h_arrdiv24_fs32_xor1;
  wire [0:0] h_arrdiv24_fs32_or0;
  wire [0:0] h_arrdiv24_fs33_xor1;
  wire [0:0] h_arrdiv24_fs33_or0;
  wire [0:0] h_arrdiv24_fs34_xor1;
  wire [0:0] h_arrdiv24_fs34_or0;
  wire [0:0] h_arrdiv24_fs35_xor1;
  wire [0:0] h_arrdiv24_fs35_or0;
  wire [0:0] h_arrdiv24_fs36_xor1;
  wire [0:0] h_arrdiv24_fs36_or0;
  wire [0:0] h_arrdiv24_fs37_xor1;
  wire [0:0] h_arrdiv24_fs37_or0;
  wire [0:0] h_arrdiv24_fs38_xor1;
  wire [0:0] h_arrdiv24_fs38_or0;
  wire [0:0] h_arrdiv24_fs39_xor1;
  wire [0:0] h_arrdiv24_fs39_or0;
  wire [0:0] h_arrdiv24_fs40_xor1;
  wire [0:0] h_arrdiv24_fs40_or0;
  wire [0:0] h_arrdiv24_fs41_xor1;
  wire [0:0] h_arrdiv24_fs41_or0;
  wire [0:0] h_arrdiv24_fs42_xor1;
  wire [0:0] h_arrdiv24_fs42_or0;
  wire [0:0] h_arrdiv24_fs43_xor1;
  wire [0:0] h_arrdiv24_fs43_or0;
  wire [0:0] h_arrdiv24_fs44_xor1;
  wire [0:0] h_arrdiv24_fs44_or0;
  wire [0:0] h_arrdiv24_fs45_xor1;
  wire [0:0] h_arrdiv24_fs45_or0;
  wire [0:0] h_arrdiv24_fs46_xor1;
  wire [0:0] h_arrdiv24_fs46_or0;
  wire [0:0] h_arrdiv24_fs47_xor1;
  wire [0:0] h_arrdiv24_fs47_or0;
  wire [0:0] h_arrdiv24_mux2to123_xor0;
  wire [0:0] h_arrdiv24_mux2to124_xor0;
  wire [0:0] h_arrdiv24_mux2to125_xor0;
  wire [0:0] h_arrdiv24_mux2to126_xor0;
  wire [0:0] h_arrdiv24_mux2to127_xor0;
  wire [0:0] h_arrdiv24_mux2to128_xor0;
  wire [0:0] h_arrdiv24_mux2to129_xor0;
  wire [0:0] h_arrdiv24_mux2to130_xor0;
  wire [0:0] h_arrdiv24_mux2to131_xor0;
  wire [0:0] h_arrdiv24_mux2to132_xor0;
  wire [0:0] h_arrdiv24_mux2to133_xor0;
  wire [0:0] h_arrdiv24_mux2to134_xor0;
  wire [0:0] h_arrdiv24_mux2to135_xor0;
  wire [0:0] h_arrdiv24_mux2to136_xor0;
  wire [0:0] h_arrdiv24_mux2to137_xor0;
  wire [0:0] h_arrdiv24_mux2to138_xor0;
  wire [0:0] h_arrdiv24_mux2to139_xor0;
  wire [0:0] h_arrdiv24_mux2to140_xor0;
  wire [0:0] h_arrdiv24_mux2to141_xor0;
  wire [0:0] h_arrdiv24_mux2to142_xor0;
  wire [0:0] h_arrdiv24_mux2to143_xor0;
  wire [0:0] h_arrdiv24_mux2to144_xor0;
  wire [0:0] h_arrdiv24_mux2to145_xor0;
  wire [0:0] h_arrdiv24_not1;
  wire [0:0] h_arrdiv24_fs48_xor0;
  wire [0:0] h_arrdiv24_fs48_and0;
  wire [0:0] h_arrdiv24_fs49_xor1;
  wire [0:0] h_arrdiv24_fs49_or0;
  wire [0:0] h_arrdiv24_fs50_xor1;
  wire [0:0] h_arrdiv24_fs50_or0;
  wire [0:0] h_arrdiv24_fs51_xor1;
  wire [0:0] h_arrdiv24_fs51_or0;
  wire [0:0] h_arrdiv24_fs52_xor1;
  wire [0:0] h_arrdiv24_fs52_or0;
  wire [0:0] h_arrdiv24_fs53_xor1;
  wire [0:0] h_arrdiv24_fs53_or0;
  wire [0:0] h_arrdiv24_fs54_xor1;
  wire [0:0] h_arrdiv24_fs54_or0;
  wire [0:0] h_arrdiv24_fs55_xor1;
  wire [0:0] h_arrdiv24_fs55_or0;
  wire [0:0] h_arrdiv24_fs56_xor1;
  wire [0:0] h_arrdiv24_fs56_or0;
  wire [0:0] h_arrdiv24_fs57_xor1;
  wire [0:0] h_arrdiv24_fs57_or0;
  wire [0:0] h_arrdiv24_fs58_xor1;
  wire [0:0] h_arrdiv24_fs58_or0;
  wire [0:0] h_arrdiv24_fs59_xor1;
  wire [0:0] h_arrdiv24_fs59_or0;
  wire [0:0] h_arrdiv24_fs60_xor1;
  wire [0:0] h_arrdiv24_fs60_or0;
  wire [0:0] h_arrdiv24_fs61_xor1;
  wire [0:0] h_arrdiv24_fs61_or0;
  wire [0:0] h_arrdiv24_fs62_xor1;
  wire [0:0] h_arrdiv24_fs62_or0;
  wire [0:0] h_arrdiv24_fs63_xor1;
  wire [0:0] h_arrdiv24_fs63_or0;
  wire [0:0] h_arrdiv24_fs64_xor1;
  wire [0:0] h_arrdiv24_fs64_or0;
  wire [0:0] h_arrdiv24_fs65_xor1;
  wire [0:0] h_arrdiv24_fs65_or0;
  wire [0:0] h_arrdiv24_fs66_xor1;
  wire [0:0] h_arrdiv24_fs66_or0;
  wire [0:0] h_arrdiv24_fs67_xor1;
  wire [0:0] h_arrdiv24_fs67_or0;
  wire [0:0] h_arrdiv24_fs68_xor1;
  wire [0:0] h_arrdiv24_fs68_or0;
  wire [0:0] h_arrdiv24_fs69_xor1;
  wire [0:0] h_arrdiv24_fs69_or0;
  wire [0:0] h_arrdiv24_fs70_xor1;
  wire [0:0] h_arrdiv24_fs70_or0;
  wire [0:0] h_arrdiv24_fs71_xor1;
  wire [0:0] h_arrdiv24_fs71_or0;
  wire [0:0] h_arrdiv24_mux2to146_xor0;
  wire [0:0] h_arrdiv24_mux2to147_xor0;
  wire [0:0] h_arrdiv24_mux2to148_xor0;
  wire [0:0] h_arrdiv24_mux2to149_xor0;
  wire [0:0] h_arrdiv24_mux2to150_xor0;
  wire [0:0] h_arrdiv24_mux2to151_xor0;
  wire [0:0] h_arrdiv24_mux2to152_xor0;
  wire [0:0] h_arrdiv24_mux2to153_xor0;
  wire [0:0] h_arrdiv24_mux2to154_xor0;
  wire [0:0] h_arrdiv24_mux2to155_xor0;
  wire [0:0] h_arrdiv24_mux2to156_xor0;
  wire [0:0] h_arrdiv24_mux2to157_xor0;
  wire [0:0] h_arrdiv24_mux2to158_xor0;
  wire [0:0] h_arrdiv24_mux2to159_xor0;
  wire [0:0] h_arrdiv24_mux2to160_xor0;
  wire [0:0] h_arrdiv24_mux2to161_xor0;
  wire [0:0] h_arrdiv24_mux2to162_xor0;
  wire [0:0] h_arrdiv24_mux2to163_xor0;
  wire [0:0] h_arrdiv24_mux2to164_xor0;
  wire [0:0] h_arrdiv24_mux2to165_xor0;
  wire [0:0] h_arrdiv24_mux2to166_xor0;
  wire [0:0] h_arrdiv24_mux2to167_xor0;
  wire [0:0] h_arrdiv24_mux2to168_xor0;
  wire [0:0] h_arrdiv24_not2;
  wire [0:0] h_arrdiv24_fs72_xor0;
  wire [0:0] h_arrdiv24_fs72_and0;
  wire [0:0] h_arrdiv24_fs73_xor1;
  wire [0:0] h_arrdiv24_fs73_or0;
  wire [0:0] h_arrdiv24_fs74_xor1;
  wire [0:0] h_arrdiv24_fs74_or0;
  wire [0:0] h_arrdiv24_fs75_xor1;
  wire [0:0] h_arrdiv24_fs75_or0;
  wire [0:0] h_arrdiv24_fs76_xor1;
  wire [0:0] h_arrdiv24_fs76_or0;
  wire [0:0] h_arrdiv24_fs77_xor1;
  wire [0:0] h_arrdiv24_fs77_or0;
  wire [0:0] h_arrdiv24_fs78_xor1;
  wire [0:0] h_arrdiv24_fs78_or0;
  wire [0:0] h_arrdiv24_fs79_xor1;
  wire [0:0] h_arrdiv24_fs79_or0;
  wire [0:0] h_arrdiv24_fs80_xor1;
  wire [0:0] h_arrdiv24_fs80_or0;
  wire [0:0] h_arrdiv24_fs81_xor1;
  wire [0:0] h_arrdiv24_fs81_or0;
  wire [0:0] h_arrdiv24_fs82_xor1;
  wire [0:0] h_arrdiv24_fs82_or0;
  wire [0:0] h_arrdiv24_fs83_xor1;
  wire [0:0] h_arrdiv24_fs83_or0;
  wire [0:0] h_arrdiv24_fs84_xor1;
  wire [0:0] h_arrdiv24_fs84_or0;
  wire [0:0] h_arrdiv24_fs85_xor1;
  wire [0:0] h_arrdiv24_fs85_or0;
  wire [0:0] h_arrdiv24_fs86_xor1;
  wire [0:0] h_arrdiv24_fs86_or0;
  wire [0:0] h_arrdiv24_fs87_xor1;
  wire [0:0] h_arrdiv24_fs87_or0;
  wire [0:0] h_arrdiv24_fs88_xor1;
  wire [0:0] h_arrdiv24_fs88_or0;
  wire [0:0] h_arrdiv24_fs89_xor1;
  wire [0:0] h_arrdiv24_fs89_or0;
  wire [0:0] h_arrdiv24_fs90_xor1;
  wire [0:0] h_arrdiv24_fs90_or0;
  wire [0:0] h_arrdiv24_fs91_xor1;
  wire [0:0] h_arrdiv24_fs91_or0;
  wire [0:0] h_arrdiv24_fs92_xor1;
  wire [0:0] h_arrdiv24_fs92_or0;
  wire [0:0] h_arrdiv24_fs93_xor1;
  wire [0:0] h_arrdiv24_fs93_or0;
  wire [0:0] h_arrdiv24_fs94_xor1;
  wire [0:0] h_arrdiv24_fs94_or0;
  wire [0:0] h_arrdiv24_fs95_xor1;
  wire [0:0] h_arrdiv24_fs95_or0;
  wire [0:0] h_arrdiv24_mux2to169_xor0;
  wire [0:0] h_arrdiv24_mux2to170_xor0;
  wire [0:0] h_arrdiv24_mux2to171_xor0;
  wire [0:0] h_arrdiv24_mux2to172_xor0;
  wire [0:0] h_arrdiv24_mux2to173_xor0;
  wire [0:0] h_arrdiv24_mux2to174_xor0;
  wire [0:0] h_arrdiv24_mux2to175_xor0;
  wire [0:0] h_arrdiv24_mux2to176_xor0;
  wire [0:0] h_arrdiv24_mux2to177_xor0;
  wire [0:0] h_arrdiv24_mux2to178_xor0;
  wire [0:0] h_arrdiv24_mux2to179_xor0;
  wire [0:0] h_arrdiv24_mux2to180_xor0;
  wire [0:0] h_arrdiv24_mux2to181_xor0;
  wire [0:0] h_arrdiv24_mux2to182_xor0;
  wire [0:0] h_arrdiv24_mux2to183_xor0;
  wire [0:0] h_arrdiv24_mux2to184_xor0;
  wire [0:0] h_arrdiv24_mux2to185_xor0;
  wire [0:0] h_arrdiv24_mux2to186_xor0;
  wire [0:0] h_arrdiv24_mux2to187_xor0;
  wire [0:0] h_arrdiv24_mux2to188_xor0;
  wire [0:0] h_arrdiv24_mux2to189_xor0;
  wire [0:0] h_arrdiv24_mux2to190_xor0;
  wire [0:0] h_arrdiv24_mux2to191_xor0;
  wire [0:0] h_arrdiv24_not3;
  wire [0:0] h_arrdiv24_fs96_xor0;
  wire [0:0] h_arrdiv24_fs96_and0;
  wire [0:0] h_arrdiv24_fs97_xor1;
  wire [0:0] h_arrdiv24_fs97_or0;
  wire [0:0] h_arrdiv24_fs98_xor1;
  wire [0:0] h_arrdiv24_fs98_or0;
  wire [0:0] h_arrdiv24_fs99_xor1;
  wire [0:0] h_arrdiv24_fs99_or0;
  wire [0:0] h_arrdiv24_fs100_xor1;
  wire [0:0] h_arrdiv24_fs100_or0;
  wire [0:0] h_arrdiv24_fs101_xor1;
  wire [0:0] h_arrdiv24_fs101_or0;
  wire [0:0] h_arrdiv24_fs102_xor1;
  wire [0:0] h_arrdiv24_fs102_or0;
  wire [0:0] h_arrdiv24_fs103_xor1;
  wire [0:0] h_arrdiv24_fs103_or0;
  wire [0:0] h_arrdiv24_fs104_xor1;
  wire [0:0] h_arrdiv24_fs104_or0;
  wire [0:0] h_arrdiv24_fs105_xor1;
  wire [0:0] h_arrdiv24_fs105_or0;
  wire [0:0] h_arrdiv24_fs106_xor1;
  wire [0:0] h_arrdiv24_fs106_or0;
  wire [0:0] h_arrdiv24_fs107_xor1;
  wire [0:0] h_arrdiv24_fs107_or0;
  wire [0:0] h_arrdiv24_fs108_xor1;
  wire [0:0] h_arrdiv24_fs108_or0;
  wire [0:0] h_arrdiv24_fs109_xor1;
  wire [0:0] h_arrdiv24_fs109_or0;
  wire [0:0] h_arrdiv24_fs110_xor1;
  wire [0:0] h_arrdiv24_fs110_or0;
  wire [0:0] h_arrdiv24_fs111_xor1;
  wire [0:0] h_arrdiv24_fs111_or0;
  wire [0:0] h_arrdiv24_fs112_xor1;
  wire [0:0] h_arrdiv24_fs112_or0;
  wire [0:0] h_arrdiv24_fs113_xor1;
  wire [0:0] h_arrdiv24_fs113_or0;
  wire [0:0] h_arrdiv24_fs114_xor1;
  wire [0:0] h_arrdiv24_fs114_or0;
  wire [0:0] h_arrdiv24_fs115_xor1;
  wire [0:0] h_arrdiv24_fs115_or0;
  wire [0:0] h_arrdiv24_fs116_xor1;
  wire [0:0] h_arrdiv24_fs116_or0;
  wire [0:0] h_arrdiv24_fs117_xor1;
  wire [0:0] h_arrdiv24_fs117_or0;
  wire [0:0] h_arrdiv24_fs118_xor1;
  wire [0:0] h_arrdiv24_fs118_or0;
  wire [0:0] h_arrdiv24_fs119_xor1;
  wire [0:0] h_arrdiv24_fs119_or0;
  wire [0:0] h_arrdiv24_mux2to192_xor0;
  wire [0:0] h_arrdiv24_mux2to193_xor0;
  wire [0:0] h_arrdiv24_mux2to194_xor0;
  wire [0:0] h_arrdiv24_mux2to195_xor0;
  wire [0:0] h_arrdiv24_mux2to196_xor0;
  wire [0:0] h_arrdiv24_mux2to197_xor0;
  wire [0:0] h_arrdiv24_mux2to198_xor0;
  wire [0:0] h_arrdiv24_mux2to199_xor0;
  wire [0:0] h_arrdiv24_mux2to1100_xor0;
  wire [0:0] h_arrdiv24_mux2to1101_xor0;
  wire [0:0] h_arrdiv24_mux2to1102_xor0;
  wire [0:0] h_arrdiv24_mux2to1103_xor0;
  wire [0:0] h_arrdiv24_mux2to1104_xor0;
  wire [0:0] h_arrdiv24_mux2to1105_xor0;
  wire [0:0] h_arrdiv24_mux2to1106_xor0;
  wire [0:0] h_arrdiv24_mux2to1107_xor0;
  wire [0:0] h_arrdiv24_mux2to1108_xor0;
  wire [0:0] h_arrdiv24_mux2to1109_xor0;
  wire [0:0] h_arrdiv24_mux2to1110_xor0;
  wire [0:0] h_arrdiv24_mux2to1111_xor0;
  wire [0:0] h_arrdiv24_mux2to1112_xor0;
  wire [0:0] h_arrdiv24_mux2to1113_xor0;
  wire [0:0] h_arrdiv24_mux2to1114_xor0;
  wire [0:0] h_arrdiv24_not4;
  wire [0:0] h_arrdiv24_fs120_xor0;
  wire [0:0] h_arrdiv24_fs120_and0;
  wire [0:0] h_arrdiv24_fs121_xor1;
  wire [0:0] h_arrdiv24_fs121_or0;
  wire [0:0] h_arrdiv24_fs122_xor1;
  wire [0:0] h_arrdiv24_fs122_or0;
  wire [0:0] h_arrdiv24_fs123_xor1;
  wire [0:0] h_arrdiv24_fs123_or0;
  wire [0:0] h_arrdiv24_fs124_xor1;
  wire [0:0] h_arrdiv24_fs124_or0;
  wire [0:0] h_arrdiv24_fs125_xor1;
  wire [0:0] h_arrdiv24_fs125_or0;
  wire [0:0] h_arrdiv24_fs126_xor1;
  wire [0:0] h_arrdiv24_fs126_or0;
  wire [0:0] h_arrdiv24_fs127_xor1;
  wire [0:0] h_arrdiv24_fs127_or0;
  wire [0:0] h_arrdiv24_fs128_xor1;
  wire [0:0] h_arrdiv24_fs128_or0;
  wire [0:0] h_arrdiv24_fs129_xor1;
  wire [0:0] h_arrdiv24_fs129_or0;
  wire [0:0] h_arrdiv24_fs130_xor1;
  wire [0:0] h_arrdiv24_fs130_or0;
  wire [0:0] h_arrdiv24_fs131_xor1;
  wire [0:0] h_arrdiv24_fs131_or0;
  wire [0:0] h_arrdiv24_fs132_xor1;
  wire [0:0] h_arrdiv24_fs132_or0;
  wire [0:0] h_arrdiv24_fs133_xor1;
  wire [0:0] h_arrdiv24_fs133_or0;
  wire [0:0] h_arrdiv24_fs134_xor1;
  wire [0:0] h_arrdiv24_fs134_or0;
  wire [0:0] h_arrdiv24_fs135_xor1;
  wire [0:0] h_arrdiv24_fs135_or0;
  wire [0:0] h_arrdiv24_fs136_xor1;
  wire [0:0] h_arrdiv24_fs136_or0;
  wire [0:0] h_arrdiv24_fs137_xor1;
  wire [0:0] h_arrdiv24_fs137_or0;
  wire [0:0] h_arrdiv24_fs138_xor1;
  wire [0:0] h_arrdiv24_fs138_or0;
  wire [0:0] h_arrdiv24_fs139_xor1;
  wire [0:0] h_arrdiv24_fs139_or0;
  wire [0:0] h_arrdiv24_fs140_xor1;
  wire [0:0] h_arrdiv24_fs140_or0;
  wire [0:0] h_arrdiv24_fs141_xor1;
  wire [0:0] h_arrdiv24_fs141_or0;
  wire [0:0] h_arrdiv24_fs142_xor1;
  wire [0:0] h_arrdiv24_fs142_or0;
  wire [0:0] h_arrdiv24_fs143_xor1;
  wire [0:0] h_arrdiv24_fs143_or0;
  wire [0:0] h_arrdiv24_mux2to1115_xor0;
  wire [0:0] h_arrdiv24_mux2to1116_xor0;
  wire [0:0] h_arrdiv24_mux2to1117_xor0;
  wire [0:0] h_arrdiv24_mux2to1118_xor0;
  wire [0:0] h_arrdiv24_mux2to1119_xor0;
  wire [0:0] h_arrdiv24_mux2to1120_xor0;
  wire [0:0] h_arrdiv24_mux2to1121_xor0;
  wire [0:0] h_arrdiv24_mux2to1122_xor0;
  wire [0:0] h_arrdiv24_mux2to1123_xor0;
  wire [0:0] h_arrdiv24_mux2to1124_xor0;
  wire [0:0] h_arrdiv24_mux2to1125_xor0;
  wire [0:0] h_arrdiv24_mux2to1126_xor0;
  wire [0:0] h_arrdiv24_mux2to1127_xor0;
  wire [0:0] h_arrdiv24_mux2to1128_xor0;
  wire [0:0] h_arrdiv24_mux2to1129_xor0;
  wire [0:0] h_arrdiv24_mux2to1130_xor0;
  wire [0:0] h_arrdiv24_mux2to1131_xor0;
  wire [0:0] h_arrdiv24_mux2to1132_xor0;
  wire [0:0] h_arrdiv24_mux2to1133_xor0;
  wire [0:0] h_arrdiv24_mux2to1134_xor0;
  wire [0:0] h_arrdiv24_mux2to1135_xor0;
  wire [0:0] h_arrdiv24_mux2to1136_xor0;
  wire [0:0] h_arrdiv24_mux2to1137_xor0;
  wire [0:0] h_arrdiv24_not5;
  wire [0:0] h_arrdiv24_fs144_xor0;
  wire [0:0] h_arrdiv24_fs144_and0;
  wire [0:0] h_arrdiv24_fs145_xor1;
  wire [0:0] h_arrdiv24_fs145_or0;
  wire [0:0] h_arrdiv24_fs146_xor1;
  wire [0:0] h_arrdiv24_fs146_or0;
  wire [0:0] h_arrdiv24_fs147_xor1;
  wire [0:0] h_arrdiv24_fs147_or0;
  wire [0:0] h_arrdiv24_fs148_xor1;
  wire [0:0] h_arrdiv24_fs148_or0;
  wire [0:0] h_arrdiv24_fs149_xor1;
  wire [0:0] h_arrdiv24_fs149_or0;
  wire [0:0] h_arrdiv24_fs150_xor1;
  wire [0:0] h_arrdiv24_fs150_or0;
  wire [0:0] h_arrdiv24_fs151_xor1;
  wire [0:0] h_arrdiv24_fs151_or0;
  wire [0:0] h_arrdiv24_fs152_xor1;
  wire [0:0] h_arrdiv24_fs152_or0;
  wire [0:0] h_arrdiv24_fs153_xor1;
  wire [0:0] h_arrdiv24_fs153_or0;
  wire [0:0] h_arrdiv24_fs154_xor1;
  wire [0:0] h_arrdiv24_fs154_or0;
  wire [0:0] h_arrdiv24_fs155_xor1;
  wire [0:0] h_arrdiv24_fs155_or0;
  wire [0:0] h_arrdiv24_fs156_xor1;
  wire [0:0] h_arrdiv24_fs156_or0;
  wire [0:0] h_arrdiv24_fs157_xor1;
  wire [0:0] h_arrdiv24_fs157_or0;
  wire [0:0] h_arrdiv24_fs158_xor1;
  wire [0:0] h_arrdiv24_fs158_or0;
  wire [0:0] h_arrdiv24_fs159_xor1;
  wire [0:0] h_arrdiv24_fs159_or0;
  wire [0:0] h_arrdiv24_fs160_xor1;
  wire [0:0] h_arrdiv24_fs160_or0;
  wire [0:0] h_arrdiv24_fs161_xor1;
  wire [0:0] h_arrdiv24_fs161_or0;
  wire [0:0] h_arrdiv24_fs162_xor1;
  wire [0:0] h_arrdiv24_fs162_or0;
  wire [0:0] h_arrdiv24_fs163_xor1;
  wire [0:0] h_arrdiv24_fs163_or0;
  wire [0:0] h_arrdiv24_fs164_xor1;
  wire [0:0] h_arrdiv24_fs164_or0;
  wire [0:0] h_arrdiv24_fs165_xor1;
  wire [0:0] h_arrdiv24_fs165_or0;
  wire [0:0] h_arrdiv24_fs166_xor1;
  wire [0:0] h_arrdiv24_fs166_or0;
  wire [0:0] h_arrdiv24_fs167_xor1;
  wire [0:0] h_arrdiv24_fs167_or0;
  wire [0:0] h_arrdiv24_mux2to1138_xor0;
  wire [0:0] h_arrdiv24_mux2to1139_xor0;
  wire [0:0] h_arrdiv24_mux2to1140_xor0;
  wire [0:0] h_arrdiv24_mux2to1141_xor0;
  wire [0:0] h_arrdiv24_mux2to1142_xor0;
  wire [0:0] h_arrdiv24_mux2to1143_xor0;
  wire [0:0] h_arrdiv24_mux2to1144_xor0;
  wire [0:0] h_arrdiv24_mux2to1145_xor0;
  wire [0:0] h_arrdiv24_mux2to1146_xor0;
  wire [0:0] h_arrdiv24_mux2to1147_xor0;
  wire [0:0] h_arrdiv24_mux2to1148_xor0;
  wire [0:0] h_arrdiv24_mux2to1149_xor0;
  wire [0:0] h_arrdiv24_mux2to1150_xor0;
  wire [0:0] h_arrdiv24_mux2to1151_xor0;
  wire [0:0] h_arrdiv24_mux2to1152_xor0;
  wire [0:0] h_arrdiv24_mux2to1153_xor0;
  wire [0:0] h_arrdiv24_mux2to1154_xor0;
  wire [0:0] h_arrdiv24_mux2to1155_xor0;
  wire [0:0] h_arrdiv24_mux2to1156_xor0;
  wire [0:0] h_arrdiv24_mux2to1157_xor0;
  wire [0:0] h_arrdiv24_mux2to1158_xor0;
  wire [0:0] h_arrdiv24_mux2to1159_xor0;
  wire [0:0] h_arrdiv24_mux2to1160_xor0;
  wire [0:0] h_arrdiv24_not6;
  wire [0:0] h_arrdiv24_fs168_xor0;
  wire [0:0] h_arrdiv24_fs168_and0;
  wire [0:0] h_arrdiv24_fs169_xor1;
  wire [0:0] h_arrdiv24_fs169_or0;
  wire [0:0] h_arrdiv24_fs170_xor1;
  wire [0:0] h_arrdiv24_fs170_or0;
  wire [0:0] h_arrdiv24_fs171_xor1;
  wire [0:0] h_arrdiv24_fs171_or0;
  wire [0:0] h_arrdiv24_fs172_xor1;
  wire [0:0] h_arrdiv24_fs172_or0;
  wire [0:0] h_arrdiv24_fs173_xor1;
  wire [0:0] h_arrdiv24_fs173_or0;
  wire [0:0] h_arrdiv24_fs174_xor1;
  wire [0:0] h_arrdiv24_fs174_or0;
  wire [0:0] h_arrdiv24_fs175_xor1;
  wire [0:0] h_arrdiv24_fs175_or0;
  wire [0:0] h_arrdiv24_fs176_xor1;
  wire [0:0] h_arrdiv24_fs176_or0;
  wire [0:0] h_arrdiv24_fs177_xor1;
  wire [0:0] h_arrdiv24_fs177_or0;
  wire [0:0] h_arrdiv24_fs178_xor1;
  wire [0:0] h_arrdiv24_fs178_or0;
  wire [0:0] h_arrdiv24_fs179_xor1;
  wire [0:0] h_arrdiv24_fs179_or0;
  wire [0:0] h_arrdiv24_fs180_xor1;
  wire [0:0] h_arrdiv24_fs180_or0;
  wire [0:0] h_arrdiv24_fs181_xor1;
  wire [0:0] h_arrdiv24_fs181_or0;
  wire [0:0] h_arrdiv24_fs182_xor1;
  wire [0:0] h_arrdiv24_fs182_or0;
  wire [0:0] h_arrdiv24_fs183_xor1;
  wire [0:0] h_arrdiv24_fs183_or0;
  wire [0:0] h_arrdiv24_fs184_xor1;
  wire [0:0] h_arrdiv24_fs184_or0;
  wire [0:0] h_arrdiv24_fs185_xor1;
  wire [0:0] h_arrdiv24_fs185_or0;
  wire [0:0] h_arrdiv24_fs186_xor1;
  wire [0:0] h_arrdiv24_fs186_or0;
  wire [0:0] h_arrdiv24_fs187_xor1;
  wire [0:0] h_arrdiv24_fs187_or0;
  wire [0:0] h_arrdiv24_fs188_xor1;
  wire [0:0] h_arrdiv24_fs188_or0;
  wire [0:0] h_arrdiv24_fs189_xor1;
  wire [0:0] h_arrdiv24_fs189_or0;
  wire [0:0] h_arrdiv24_fs190_xor1;
  wire [0:0] h_arrdiv24_fs190_or0;
  wire [0:0] h_arrdiv24_fs191_xor1;
  wire [0:0] h_arrdiv24_fs191_or0;
  wire [0:0] h_arrdiv24_mux2to1161_xor0;
  wire [0:0] h_arrdiv24_mux2to1162_xor0;
  wire [0:0] h_arrdiv24_mux2to1163_xor0;
  wire [0:0] h_arrdiv24_mux2to1164_xor0;
  wire [0:0] h_arrdiv24_mux2to1165_xor0;
  wire [0:0] h_arrdiv24_mux2to1166_xor0;
  wire [0:0] h_arrdiv24_mux2to1167_xor0;
  wire [0:0] h_arrdiv24_mux2to1168_xor0;
  wire [0:0] h_arrdiv24_mux2to1169_xor0;
  wire [0:0] h_arrdiv24_mux2to1170_xor0;
  wire [0:0] h_arrdiv24_mux2to1171_xor0;
  wire [0:0] h_arrdiv24_mux2to1172_xor0;
  wire [0:0] h_arrdiv24_mux2to1173_xor0;
  wire [0:0] h_arrdiv24_mux2to1174_xor0;
  wire [0:0] h_arrdiv24_mux2to1175_xor0;
  wire [0:0] h_arrdiv24_mux2to1176_xor0;
  wire [0:0] h_arrdiv24_mux2to1177_xor0;
  wire [0:0] h_arrdiv24_mux2to1178_xor0;
  wire [0:0] h_arrdiv24_mux2to1179_xor0;
  wire [0:0] h_arrdiv24_mux2to1180_xor0;
  wire [0:0] h_arrdiv24_mux2to1181_xor0;
  wire [0:0] h_arrdiv24_mux2to1182_xor0;
  wire [0:0] h_arrdiv24_mux2to1183_xor0;
  wire [0:0] h_arrdiv24_not7;
  wire [0:0] h_arrdiv24_fs192_xor0;
  wire [0:0] h_arrdiv24_fs192_and0;
  wire [0:0] h_arrdiv24_fs193_xor1;
  wire [0:0] h_arrdiv24_fs193_or0;
  wire [0:0] h_arrdiv24_fs194_xor1;
  wire [0:0] h_arrdiv24_fs194_or0;
  wire [0:0] h_arrdiv24_fs195_xor1;
  wire [0:0] h_arrdiv24_fs195_or0;
  wire [0:0] h_arrdiv24_fs196_xor1;
  wire [0:0] h_arrdiv24_fs196_or0;
  wire [0:0] h_arrdiv24_fs197_xor1;
  wire [0:0] h_arrdiv24_fs197_or0;
  wire [0:0] h_arrdiv24_fs198_xor1;
  wire [0:0] h_arrdiv24_fs198_or0;
  wire [0:0] h_arrdiv24_fs199_xor1;
  wire [0:0] h_arrdiv24_fs199_or0;
  wire [0:0] h_arrdiv24_fs200_xor1;
  wire [0:0] h_arrdiv24_fs200_or0;
  wire [0:0] h_arrdiv24_fs201_xor1;
  wire [0:0] h_arrdiv24_fs201_or0;
  wire [0:0] h_arrdiv24_fs202_xor1;
  wire [0:0] h_arrdiv24_fs202_or0;
  wire [0:0] h_arrdiv24_fs203_xor1;
  wire [0:0] h_arrdiv24_fs203_or0;
  wire [0:0] h_arrdiv24_fs204_xor1;
  wire [0:0] h_arrdiv24_fs204_or0;
  wire [0:0] h_arrdiv24_fs205_xor1;
  wire [0:0] h_arrdiv24_fs205_or0;
  wire [0:0] h_arrdiv24_fs206_xor1;
  wire [0:0] h_arrdiv24_fs206_or0;
  wire [0:0] h_arrdiv24_fs207_xor1;
  wire [0:0] h_arrdiv24_fs207_or0;
  wire [0:0] h_arrdiv24_fs208_xor1;
  wire [0:0] h_arrdiv24_fs208_or0;
  wire [0:0] h_arrdiv24_fs209_xor1;
  wire [0:0] h_arrdiv24_fs209_or0;
  wire [0:0] h_arrdiv24_fs210_xor1;
  wire [0:0] h_arrdiv24_fs210_or0;
  wire [0:0] h_arrdiv24_fs211_xor1;
  wire [0:0] h_arrdiv24_fs211_or0;
  wire [0:0] h_arrdiv24_fs212_xor1;
  wire [0:0] h_arrdiv24_fs212_or0;
  wire [0:0] h_arrdiv24_fs213_xor1;
  wire [0:0] h_arrdiv24_fs213_or0;
  wire [0:0] h_arrdiv24_fs214_xor1;
  wire [0:0] h_arrdiv24_fs214_or0;
  wire [0:0] h_arrdiv24_fs215_xor1;
  wire [0:0] h_arrdiv24_fs215_or0;
  wire [0:0] h_arrdiv24_mux2to1184_xor0;
  wire [0:0] h_arrdiv24_mux2to1185_xor0;
  wire [0:0] h_arrdiv24_mux2to1186_xor0;
  wire [0:0] h_arrdiv24_mux2to1187_xor0;
  wire [0:0] h_arrdiv24_mux2to1188_xor0;
  wire [0:0] h_arrdiv24_mux2to1189_xor0;
  wire [0:0] h_arrdiv24_mux2to1190_xor0;
  wire [0:0] h_arrdiv24_mux2to1191_xor0;
  wire [0:0] h_arrdiv24_mux2to1192_xor0;
  wire [0:0] h_arrdiv24_mux2to1193_xor0;
  wire [0:0] h_arrdiv24_mux2to1194_xor0;
  wire [0:0] h_arrdiv24_mux2to1195_xor0;
  wire [0:0] h_arrdiv24_mux2to1196_xor0;
  wire [0:0] h_arrdiv24_mux2to1197_xor0;
  wire [0:0] h_arrdiv24_mux2to1198_xor0;
  wire [0:0] h_arrdiv24_mux2to1199_xor0;
  wire [0:0] h_arrdiv24_mux2to1200_xor0;
  wire [0:0] h_arrdiv24_mux2to1201_xor0;
  wire [0:0] h_arrdiv24_mux2to1202_xor0;
  wire [0:0] h_arrdiv24_mux2to1203_xor0;
  wire [0:0] h_arrdiv24_mux2to1204_xor0;
  wire [0:0] h_arrdiv24_mux2to1205_xor0;
  wire [0:0] h_arrdiv24_mux2to1206_xor0;
  wire [0:0] h_arrdiv24_not8;
  wire [0:0] h_arrdiv24_fs216_xor0;
  wire [0:0] h_arrdiv24_fs216_and0;
  wire [0:0] h_arrdiv24_fs217_xor1;
  wire [0:0] h_arrdiv24_fs217_or0;
  wire [0:0] h_arrdiv24_fs218_xor1;
  wire [0:0] h_arrdiv24_fs218_or0;
  wire [0:0] h_arrdiv24_fs219_xor1;
  wire [0:0] h_arrdiv24_fs219_or0;
  wire [0:0] h_arrdiv24_fs220_xor1;
  wire [0:0] h_arrdiv24_fs220_or0;
  wire [0:0] h_arrdiv24_fs221_xor1;
  wire [0:0] h_arrdiv24_fs221_or0;
  wire [0:0] h_arrdiv24_fs222_xor1;
  wire [0:0] h_arrdiv24_fs222_or0;
  wire [0:0] h_arrdiv24_fs223_xor1;
  wire [0:0] h_arrdiv24_fs223_or0;
  wire [0:0] h_arrdiv24_fs224_xor1;
  wire [0:0] h_arrdiv24_fs224_or0;
  wire [0:0] h_arrdiv24_fs225_xor1;
  wire [0:0] h_arrdiv24_fs225_or0;
  wire [0:0] h_arrdiv24_fs226_xor1;
  wire [0:0] h_arrdiv24_fs226_or0;
  wire [0:0] h_arrdiv24_fs227_xor1;
  wire [0:0] h_arrdiv24_fs227_or0;
  wire [0:0] h_arrdiv24_fs228_xor1;
  wire [0:0] h_arrdiv24_fs228_or0;
  wire [0:0] h_arrdiv24_fs229_xor1;
  wire [0:0] h_arrdiv24_fs229_or0;
  wire [0:0] h_arrdiv24_fs230_xor1;
  wire [0:0] h_arrdiv24_fs230_or0;
  wire [0:0] h_arrdiv24_fs231_xor1;
  wire [0:0] h_arrdiv24_fs231_or0;
  wire [0:0] h_arrdiv24_fs232_xor1;
  wire [0:0] h_arrdiv24_fs232_or0;
  wire [0:0] h_arrdiv24_fs233_xor1;
  wire [0:0] h_arrdiv24_fs233_or0;
  wire [0:0] h_arrdiv24_fs234_xor1;
  wire [0:0] h_arrdiv24_fs234_or0;
  wire [0:0] h_arrdiv24_fs235_xor1;
  wire [0:0] h_arrdiv24_fs235_or0;
  wire [0:0] h_arrdiv24_fs236_xor1;
  wire [0:0] h_arrdiv24_fs236_or0;
  wire [0:0] h_arrdiv24_fs237_xor1;
  wire [0:0] h_arrdiv24_fs237_or0;
  wire [0:0] h_arrdiv24_fs238_xor1;
  wire [0:0] h_arrdiv24_fs238_or0;
  wire [0:0] h_arrdiv24_fs239_xor1;
  wire [0:0] h_arrdiv24_fs239_or0;
  wire [0:0] h_arrdiv24_mux2to1207_xor0;
  wire [0:0] h_arrdiv24_mux2to1208_xor0;
  wire [0:0] h_arrdiv24_mux2to1209_xor0;
  wire [0:0] h_arrdiv24_mux2to1210_xor0;
  wire [0:0] h_arrdiv24_mux2to1211_xor0;
  wire [0:0] h_arrdiv24_mux2to1212_xor0;
  wire [0:0] h_arrdiv24_mux2to1213_xor0;
  wire [0:0] h_arrdiv24_mux2to1214_xor0;
  wire [0:0] h_arrdiv24_mux2to1215_xor0;
  wire [0:0] h_arrdiv24_mux2to1216_xor0;
  wire [0:0] h_arrdiv24_mux2to1217_xor0;
  wire [0:0] h_arrdiv24_mux2to1218_xor0;
  wire [0:0] h_arrdiv24_mux2to1219_xor0;
  wire [0:0] h_arrdiv24_mux2to1220_xor0;
  wire [0:0] h_arrdiv24_mux2to1221_xor0;
  wire [0:0] h_arrdiv24_mux2to1222_xor0;
  wire [0:0] h_arrdiv24_mux2to1223_xor0;
  wire [0:0] h_arrdiv24_mux2to1224_xor0;
  wire [0:0] h_arrdiv24_mux2to1225_xor0;
  wire [0:0] h_arrdiv24_mux2to1226_xor0;
  wire [0:0] h_arrdiv24_mux2to1227_xor0;
  wire [0:0] h_arrdiv24_mux2to1228_xor0;
  wire [0:0] h_arrdiv24_mux2to1229_xor0;
  wire [0:0] h_arrdiv24_not9;
  wire [0:0] h_arrdiv24_fs240_xor0;
  wire [0:0] h_arrdiv24_fs240_and0;
  wire [0:0] h_arrdiv24_fs241_xor1;
  wire [0:0] h_arrdiv24_fs241_or0;
  wire [0:0] h_arrdiv24_fs242_xor1;
  wire [0:0] h_arrdiv24_fs242_or0;
  wire [0:0] h_arrdiv24_fs243_xor1;
  wire [0:0] h_arrdiv24_fs243_or0;
  wire [0:0] h_arrdiv24_fs244_xor1;
  wire [0:0] h_arrdiv24_fs244_or0;
  wire [0:0] h_arrdiv24_fs245_xor1;
  wire [0:0] h_arrdiv24_fs245_or0;
  wire [0:0] h_arrdiv24_fs246_xor1;
  wire [0:0] h_arrdiv24_fs246_or0;
  wire [0:0] h_arrdiv24_fs247_xor1;
  wire [0:0] h_arrdiv24_fs247_or0;
  wire [0:0] h_arrdiv24_fs248_xor1;
  wire [0:0] h_arrdiv24_fs248_or0;
  wire [0:0] h_arrdiv24_fs249_xor1;
  wire [0:0] h_arrdiv24_fs249_or0;
  wire [0:0] h_arrdiv24_fs250_xor1;
  wire [0:0] h_arrdiv24_fs250_or0;
  wire [0:0] h_arrdiv24_fs251_xor1;
  wire [0:0] h_arrdiv24_fs251_or0;
  wire [0:0] h_arrdiv24_fs252_xor1;
  wire [0:0] h_arrdiv24_fs252_or0;
  wire [0:0] h_arrdiv24_fs253_xor1;
  wire [0:0] h_arrdiv24_fs253_or0;
  wire [0:0] h_arrdiv24_fs254_xor1;
  wire [0:0] h_arrdiv24_fs254_or0;
  wire [0:0] h_arrdiv24_fs255_xor1;
  wire [0:0] h_arrdiv24_fs255_or0;
  wire [0:0] h_arrdiv24_fs256_xor1;
  wire [0:0] h_arrdiv24_fs256_or0;
  wire [0:0] h_arrdiv24_fs257_xor1;
  wire [0:0] h_arrdiv24_fs257_or0;
  wire [0:0] h_arrdiv24_fs258_xor1;
  wire [0:0] h_arrdiv24_fs258_or0;
  wire [0:0] h_arrdiv24_fs259_xor1;
  wire [0:0] h_arrdiv24_fs259_or0;
  wire [0:0] h_arrdiv24_fs260_xor1;
  wire [0:0] h_arrdiv24_fs260_or0;
  wire [0:0] h_arrdiv24_fs261_xor1;
  wire [0:0] h_arrdiv24_fs261_or0;
  wire [0:0] h_arrdiv24_fs262_xor1;
  wire [0:0] h_arrdiv24_fs262_or0;
  wire [0:0] h_arrdiv24_fs263_xor1;
  wire [0:0] h_arrdiv24_fs263_or0;
  wire [0:0] h_arrdiv24_mux2to1230_xor0;
  wire [0:0] h_arrdiv24_mux2to1231_xor0;
  wire [0:0] h_arrdiv24_mux2to1232_xor0;
  wire [0:0] h_arrdiv24_mux2to1233_xor0;
  wire [0:0] h_arrdiv24_mux2to1234_xor0;
  wire [0:0] h_arrdiv24_mux2to1235_xor0;
  wire [0:0] h_arrdiv24_mux2to1236_xor0;
  wire [0:0] h_arrdiv24_mux2to1237_xor0;
  wire [0:0] h_arrdiv24_mux2to1238_xor0;
  wire [0:0] h_arrdiv24_mux2to1239_xor0;
  wire [0:0] h_arrdiv24_mux2to1240_xor0;
  wire [0:0] h_arrdiv24_mux2to1241_xor0;
  wire [0:0] h_arrdiv24_mux2to1242_xor0;
  wire [0:0] h_arrdiv24_mux2to1243_xor0;
  wire [0:0] h_arrdiv24_mux2to1244_xor0;
  wire [0:0] h_arrdiv24_mux2to1245_xor0;
  wire [0:0] h_arrdiv24_mux2to1246_xor0;
  wire [0:0] h_arrdiv24_mux2to1247_xor0;
  wire [0:0] h_arrdiv24_mux2to1248_xor0;
  wire [0:0] h_arrdiv24_mux2to1249_xor0;
  wire [0:0] h_arrdiv24_mux2to1250_xor0;
  wire [0:0] h_arrdiv24_mux2to1251_xor0;
  wire [0:0] h_arrdiv24_mux2to1252_xor0;
  wire [0:0] h_arrdiv24_not10;
  wire [0:0] h_arrdiv24_fs264_xor0;
  wire [0:0] h_arrdiv24_fs264_and0;
  wire [0:0] h_arrdiv24_fs265_xor1;
  wire [0:0] h_arrdiv24_fs265_or0;
  wire [0:0] h_arrdiv24_fs266_xor1;
  wire [0:0] h_arrdiv24_fs266_or0;
  wire [0:0] h_arrdiv24_fs267_xor1;
  wire [0:0] h_arrdiv24_fs267_or0;
  wire [0:0] h_arrdiv24_fs268_xor1;
  wire [0:0] h_arrdiv24_fs268_or0;
  wire [0:0] h_arrdiv24_fs269_xor1;
  wire [0:0] h_arrdiv24_fs269_or0;
  wire [0:0] h_arrdiv24_fs270_xor1;
  wire [0:0] h_arrdiv24_fs270_or0;
  wire [0:0] h_arrdiv24_fs271_xor1;
  wire [0:0] h_arrdiv24_fs271_or0;
  wire [0:0] h_arrdiv24_fs272_xor1;
  wire [0:0] h_arrdiv24_fs272_or0;
  wire [0:0] h_arrdiv24_fs273_xor1;
  wire [0:0] h_arrdiv24_fs273_or0;
  wire [0:0] h_arrdiv24_fs274_xor1;
  wire [0:0] h_arrdiv24_fs274_or0;
  wire [0:0] h_arrdiv24_fs275_xor1;
  wire [0:0] h_arrdiv24_fs275_or0;
  wire [0:0] h_arrdiv24_fs276_xor1;
  wire [0:0] h_arrdiv24_fs276_or0;
  wire [0:0] h_arrdiv24_fs277_xor1;
  wire [0:0] h_arrdiv24_fs277_or0;
  wire [0:0] h_arrdiv24_fs278_xor1;
  wire [0:0] h_arrdiv24_fs278_or0;
  wire [0:0] h_arrdiv24_fs279_xor1;
  wire [0:0] h_arrdiv24_fs279_or0;
  wire [0:0] h_arrdiv24_fs280_xor1;
  wire [0:0] h_arrdiv24_fs280_or0;
  wire [0:0] h_arrdiv24_fs281_xor1;
  wire [0:0] h_arrdiv24_fs281_or0;
  wire [0:0] h_arrdiv24_fs282_xor1;
  wire [0:0] h_arrdiv24_fs282_or0;
  wire [0:0] h_arrdiv24_fs283_xor1;
  wire [0:0] h_arrdiv24_fs283_or0;
  wire [0:0] h_arrdiv24_fs284_xor1;
  wire [0:0] h_arrdiv24_fs284_or0;
  wire [0:0] h_arrdiv24_fs285_xor1;
  wire [0:0] h_arrdiv24_fs285_or0;
  wire [0:0] h_arrdiv24_fs286_xor1;
  wire [0:0] h_arrdiv24_fs286_or0;
  wire [0:0] h_arrdiv24_fs287_xor1;
  wire [0:0] h_arrdiv24_fs287_or0;
  wire [0:0] h_arrdiv24_mux2to1253_xor0;
  wire [0:0] h_arrdiv24_mux2to1254_xor0;
  wire [0:0] h_arrdiv24_mux2to1255_xor0;
  wire [0:0] h_arrdiv24_mux2to1256_xor0;
  wire [0:0] h_arrdiv24_mux2to1257_xor0;
  wire [0:0] h_arrdiv24_mux2to1258_xor0;
  wire [0:0] h_arrdiv24_mux2to1259_xor0;
  wire [0:0] h_arrdiv24_mux2to1260_xor0;
  wire [0:0] h_arrdiv24_mux2to1261_xor0;
  wire [0:0] h_arrdiv24_mux2to1262_xor0;
  wire [0:0] h_arrdiv24_mux2to1263_xor0;
  wire [0:0] h_arrdiv24_mux2to1264_xor0;
  wire [0:0] h_arrdiv24_mux2to1265_xor0;
  wire [0:0] h_arrdiv24_mux2to1266_xor0;
  wire [0:0] h_arrdiv24_mux2to1267_xor0;
  wire [0:0] h_arrdiv24_mux2to1268_xor0;
  wire [0:0] h_arrdiv24_mux2to1269_xor0;
  wire [0:0] h_arrdiv24_mux2to1270_xor0;
  wire [0:0] h_arrdiv24_mux2to1271_xor0;
  wire [0:0] h_arrdiv24_mux2to1272_xor0;
  wire [0:0] h_arrdiv24_mux2to1273_xor0;
  wire [0:0] h_arrdiv24_mux2to1274_xor0;
  wire [0:0] h_arrdiv24_mux2to1275_xor0;
  wire [0:0] h_arrdiv24_not11;
  wire [0:0] h_arrdiv24_fs288_xor0;
  wire [0:0] h_arrdiv24_fs288_and0;
  wire [0:0] h_arrdiv24_fs289_xor1;
  wire [0:0] h_arrdiv24_fs289_or0;
  wire [0:0] h_arrdiv24_fs290_xor1;
  wire [0:0] h_arrdiv24_fs290_or0;
  wire [0:0] h_arrdiv24_fs291_xor1;
  wire [0:0] h_arrdiv24_fs291_or0;
  wire [0:0] h_arrdiv24_fs292_xor1;
  wire [0:0] h_arrdiv24_fs292_or0;
  wire [0:0] h_arrdiv24_fs293_xor1;
  wire [0:0] h_arrdiv24_fs293_or0;
  wire [0:0] h_arrdiv24_fs294_xor1;
  wire [0:0] h_arrdiv24_fs294_or0;
  wire [0:0] h_arrdiv24_fs295_xor1;
  wire [0:0] h_arrdiv24_fs295_or0;
  wire [0:0] h_arrdiv24_fs296_xor1;
  wire [0:0] h_arrdiv24_fs296_or0;
  wire [0:0] h_arrdiv24_fs297_xor1;
  wire [0:0] h_arrdiv24_fs297_or0;
  wire [0:0] h_arrdiv24_fs298_xor1;
  wire [0:0] h_arrdiv24_fs298_or0;
  wire [0:0] h_arrdiv24_fs299_xor1;
  wire [0:0] h_arrdiv24_fs299_or0;
  wire [0:0] h_arrdiv24_fs300_xor1;
  wire [0:0] h_arrdiv24_fs300_or0;
  wire [0:0] h_arrdiv24_fs301_xor1;
  wire [0:0] h_arrdiv24_fs301_or0;
  wire [0:0] h_arrdiv24_fs302_xor1;
  wire [0:0] h_arrdiv24_fs302_or0;
  wire [0:0] h_arrdiv24_fs303_xor1;
  wire [0:0] h_arrdiv24_fs303_or0;
  wire [0:0] h_arrdiv24_fs304_xor1;
  wire [0:0] h_arrdiv24_fs304_or0;
  wire [0:0] h_arrdiv24_fs305_xor1;
  wire [0:0] h_arrdiv24_fs305_or0;
  wire [0:0] h_arrdiv24_fs306_xor1;
  wire [0:0] h_arrdiv24_fs306_or0;
  wire [0:0] h_arrdiv24_fs307_xor1;
  wire [0:0] h_arrdiv24_fs307_or0;
  wire [0:0] h_arrdiv24_fs308_xor1;
  wire [0:0] h_arrdiv24_fs308_or0;
  wire [0:0] h_arrdiv24_fs309_xor1;
  wire [0:0] h_arrdiv24_fs309_or0;
  wire [0:0] h_arrdiv24_fs310_xor1;
  wire [0:0] h_arrdiv24_fs310_or0;
  wire [0:0] h_arrdiv24_fs311_xor1;
  wire [0:0] h_arrdiv24_fs311_or0;
  wire [0:0] h_arrdiv24_mux2to1276_xor0;
  wire [0:0] h_arrdiv24_mux2to1277_xor0;
  wire [0:0] h_arrdiv24_mux2to1278_xor0;
  wire [0:0] h_arrdiv24_mux2to1279_xor0;
  wire [0:0] h_arrdiv24_mux2to1280_xor0;
  wire [0:0] h_arrdiv24_mux2to1281_xor0;
  wire [0:0] h_arrdiv24_mux2to1282_xor0;
  wire [0:0] h_arrdiv24_mux2to1283_xor0;
  wire [0:0] h_arrdiv24_mux2to1284_xor0;
  wire [0:0] h_arrdiv24_mux2to1285_xor0;
  wire [0:0] h_arrdiv24_mux2to1286_xor0;
  wire [0:0] h_arrdiv24_mux2to1287_xor0;
  wire [0:0] h_arrdiv24_mux2to1288_xor0;
  wire [0:0] h_arrdiv24_mux2to1289_xor0;
  wire [0:0] h_arrdiv24_mux2to1290_xor0;
  wire [0:0] h_arrdiv24_mux2to1291_xor0;
  wire [0:0] h_arrdiv24_mux2to1292_xor0;
  wire [0:0] h_arrdiv24_mux2to1293_xor0;
  wire [0:0] h_arrdiv24_mux2to1294_xor0;
  wire [0:0] h_arrdiv24_mux2to1295_xor0;
  wire [0:0] h_arrdiv24_mux2to1296_xor0;
  wire [0:0] h_arrdiv24_mux2to1297_xor0;
  wire [0:0] h_arrdiv24_mux2to1298_xor0;
  wire [0:0] h_arrdiv24_not12;
  wire [0:0] h_arrdiv24_fs312_xor0;
  wire [0:0] h_arrdiv24_fs312_and0;
  wire [0:0] h_arrdiv24_fs313_xor1;
  wire [0:0] h_arrdiv24_fs313_or0;
  wire [0:0] h_arrdiv24_fs314_xor1;
  wire [0:0] h_arrdiv24_fs314_or0;
  wire [0:0] h_arrdiv24_fs315_xor1;
  wire [0:0] h_arrdiv24_fs315_or0;
  wire [0:0] h_arrdiv24_fs316_xor1;
  wire [0:0] h_arrdiv24_fs316_or0;
  wire [0:0] h_arrdiv24_fs317_xor1;
  wire [0:0] h_arrdiv24_fs317_or0;
  wire [0:0] h_arrdiv24_fs318_xor1;
  wire [0:0] h_arrdiv24_fs318_or0;
  wire [0:0] h_arrdiv24_fs319_xor1;
  wire [0:0] h_arrdiv24_fs319_or0;
  wire [0:0] h_arrdiv24_fs320_xor1;
  wire [0:0] h_arrdiv24_fs320_or0;
  wire [0:0] h_arrdiv24_fs321_xor1;
  wire [0:0] h_arrdiv24_fs321_or0;
  wire [0:0] h_arrdiv24_fs322_xor1;
  wire [0:0] h_arrdiv24_fs322_or0;
  wire [0:0] h_arrdiv24_fs323_xor1;
  wire [0:0] h_arrdiv24_fs323_or0;
  wire [0:0] h_arrdiv24_fs324_xor1;
  wire [0:0] h_arrdiv24_fs324_or0;
  wire [0:0] h_arrdiv24_fs325_xor1;
  wire [0:0] h_arrdiv24_fs325_or0;
  wire [0:0] h_arrdiv24_fs326_xor1;
  wire [0:0] h_arrdiv24_fs326_or0;
  wire [0:0] h_arrdiv24_fs327_xor1;
  wire [0:0] h_arrdiv24_fs327_or0;
  wire [0:0] h_arrdiv24_fs328_xor1;
  wire [0:0] h_arrdiv24_fs328_or0;
  wire [0:0] h_arrdiv24_fs329_xor1;
  wire [0:0] h_arrdiv24_fs329_or0;
  wire [0:0] h_arrdiv24_fs330_xor1;
  wire [0:0] h_arrdiv24_fs330_or0;
  wire [0:0] h_arrdiv24_fs331_xor1;
  wire [0:0] h_arrdiv24_fs331_or0;
  wire [0:0] h_arrdiv24_fs332_xor1;
  wire [0:0] h_arrdiv24_fs332_or0;
  wire [0:0] h_arrdiv24_fs333_xor1;
  wire [0:0] h_arrdiv24_fs333_or0;
  wire [0:0] h_arrdiv24_fs334_xor1;
  wire [0:0] h_arrdiv24_fs334_or0;
  wire [0:0] h_arrdiv24_fs335_xor1;
  wire [0:0] h_arrdiv24_fs335_or0;
  wire [0:0] h_arrdiv24_mux2to1299_xor0;
  wire [0:0] h_arrdiv24_mux2to1300_xor0;
  wire [0:0] h_arrdiv24_mux2to1301_xor0;
  wire [0:0] h_arrdiv24_mux2to1302_xor0;
  wire [0:0] h_arrdiv24_mux2to1303_xor0;
  wire [0:0] h_arrdiv24_mux2to1304_xor0;
  wire [0:0] h_arrdiv24_mux2to1305_xor0;
  wire [0:0] h_arrdiv24_mux2to1306_xor0;
  wire [0:0] h_arrdiv24_mux2to1307_xor0;
  wire [0:0] h_arrdiv24_mux2to1308_xor0;
  wire [0:0] h_arrdiv24_mux2to1309_xor0;
  wire [0:0] h_arrdiv24_mux2to1310_xor0;
  wire [0:0] h_arrdiv24_mux2to1311_xor0;
  wire [0:0] h_arrdiv24_mux2to1312_xor0;
  wire [0:0] h_arrdiv24_mux2to1313_xor0;
  wire [0:0] h_arrdiv24_mux2to1314_xor0;
  wire [0:0] h_arrdiv24_mux2to1315_xor0;
  wire [0:0] h_arrdiv24_mux2to1316_xor0;
  wire [0:0] h_arrdiv24_mux2to1317_xor0;
  wire [0:0] h_arrdiv24_mux2to1318_xor0;
  wire [0:0] h_arrdiv24_mux2to1319_xor0;
  wire [0:0] h_arrdiv24_mux2to1320_xor0;
  wire [0:0] h_arrdiv24_mux2to1321_xor0;
  wire [0:0] h_arrdiv24_not13;
  wire [0:0] h_arrdiv24_fs336_xor0;
  wire [0:0] h_arrdiv24_fs336_and0;
  wire [0:0] h_arrdiv24_fs337_xor1;
  wire [0:0] h_arrdiv24_fs337_or0;
  wire [0:0] h_arrdiv24_fs338_xor1;
  wire [0:0] h_arrdiv24_fs338_or0;
  wire [0:0] h_arrdiv24_fs339_xor1;
  wire [0:0] h_arrdiv24_fs339_or0;
  wire [0:0] h_arrdiv24_fs340_xor1;
  wire [0:0] h_arrdiv24_fs340_or0;
  wire [0:0] h_arrdiv24_fs341_xor1;
  wire [0:0] h_arrdiv24_fs341_or0;
  wire [0:0] h_arrdiv24_fs342_xor1;
  wire [0:0] h_arrdiv24_fs342_or0;
  wire [0:0] h_arrdiv24_fs343_xor1;
  wire [0:0] h_arrdiv24_fs343_or0;
  wire [0:0] h_arrdiv24_fs344_xor1;
  wire [0:0] h_arrdiv24_fs344_or0;
  wire [0:0] h_arrdiv24_fs345_xor1;
  wire [0:0] h_arrdiv24_fs345_or0;
  wire [0:0] h_arrdiv24_fs346_xor1;
  wire [0:0] h_arrdiv24_fs346_or0;
  wire [0:0] h_arrdiv24_fs347_xor1;
  wire [0:0] h_arrdiv24_fs347_or0;
  wire [0:0] h_arrdiv24_fs348_xor1;
  wire [0:0] h_arrdiv24_fs348_or0;
  wire [0:0] h_arrdiv24_fs349_xor1;
  wire [0:0] h_arrdiv24_fs349_or0;
  wire [0:0] h_arrdiv24_fs350_xor1;
  wire [0:0] h_arrdiv24_fs350_or0;
  wire [0:0] h_arrdiv24_fs351_xor1;
  wire [0:0] h_arrdiv24_fs351_or0;
  wire [0:0] h_arrdiv24_fs352_xor1;
  wire [0:0] h_arrdiv24_fs352_or0;
  wire [0:0] h_arrdiv24_fs353_xor1;
  wire [0:0] h_arrdiv24_fs353_or0;
  wire [0:0] h_arrdiv24_fs354_xor1;
  wire [0:0] h_arrdiv24_fs354_or0;
  wire [0:0] h_arrdiv24_fs355_xor1;
  wire [0:0] h_arrdiv24_fs355_or0;
  wire [0:0] h_arrdiv24_fs356_xor1;
  wire [0:0] h_arrdiv24_fs356_or0;
  wire [0:0] h_arrdiv24_fs357_xor1;
  wire [0:0] h_arrdiv24_fs357_or0;
  wire [0:0] h_arrdiv24_fs358_xor1;
  wire [0:0] h_arrdiv24_fs358_or0;
  wire [0:0] h_arrdiv24_fs359_xor1;
  wire [0:0] h_arrdiv24_fs359_or0;
  wire [0:0] h_arrdiv24_mux2to1322_xor0;
  wire [0:0] h_arrdiv24_mux2to1323_xor0;
  wire [0:0] h_arrdiv24_mux2to1324_xor0;
  wire [0:0] h_arrdiv24_mux2to1325_xor0;
  wire [0:0] h_arrdiv24_mux2to1326_xor0;
  wire [0:0] h_arrdiv24_mux2to1327_xor0;
  wire [0:0] h_arrdiv24_mux2to1328_xor0;
  wire [0:0] h_arrdiv24_mux2to1329_xor0;
  wire [0:0] h_arrdiv24_mux2to1330_xor0;
  wire [0:0] h_arrdiv24_mux2to1331_xor0;
  wire [0:0] h_arrdiv24_mux2to1332_xor0;
  wire [0:0] h_arrdiv24_mux2to1333_xor0;
  wire [0:0] h_arrdiv24_mux2to1334_xor0;
  wire [0:0] h_arrdiv24_mux2to1335_xor0;
  wire [0:0] h_arrdiv24_mux2to1336_xor0;
  wire [0:0] h_arrdiv24_mux2to1337_xor0;
  wire [0:0] h_arrdiv24_mux2to1338_xor0;
  wire [0:0] h_arrdiv24_mux2to1339_xor0;
  wire [0:0] h_arrdiv24_mux2to1340_xor0;
  wire [0:0] h_arrdiv24_mux2to1341_xor0;
  wire [0:0] h_arrdiv24_mux2to1342_xor0;
  wire [0:0] h_arrdiv24_mux2to1343_xor0;
  wire [0:0] h_arrdiv24_mux2to1344_xor0;
  wire [0:0] h_arrdiv24_not14;
  wire [0:0] h_arrdiv24_fs360_xor0;
  wire [0:0] h_arrdiv24_fs360_and0;
  wire [0:0] h_arrdiv24_fs361_xor1;
  wire [0:0] h_arrdiv24_fs361_or0;
  wire [0:0] h_arrdiv24_fs362_xor1;
  wire [0:0] h_arrdiv24_fs362_or0;
  wire [0:0] h_arrdiv24_fs363_xor1;
  wire [0:0] h_arrdiv24_fs363_or0;
  wire [0:0] h_arrdiv24_fs364_xor1;
  wire [0:0] h_arrdiv24_fs364_or0;
  wire [0:0] h_arrdiv24_fs365_xor1;
  wire [0:0] h_arrdiv24_fs365_or0;
  wire [0:0] h_arrdiv24_fs366_xor1;
  wire [0:0] h_arrdiv24_fs366_or0;
  wire [0:0] h_arrdiv24_fs367_xor1;
  wire [0:0] h_arrdiv24_fs367_or0;
  wire [0:0] h_arrdiv24_fs368_xor1;
  wire [0:0] h_arrdiv24_fs368_or0;
  wire [0:0] h_arrdiv24_fs369_xor1;
  wire [0:0] h_arrdiv24_fs369_or0;
  wire [0:0] h_arrdiv24_fs370_xor1;
  wire [0:0] h_arrdiv24_fs370_or0;
  wire [0:0] h_arrdiv24_fs371_xor1;
  wire [0:0] h_arrdiv24_fs371_or0;
  wire [0:0] h_arrdiv24_fs372_xor1;
  wire [0:0] h_arrdiv24_fs372_or0;
  wire [0:0] h_arrdiv24_fs373_xor1;
  wire [0:0] h_arrdiv24_fs373_or0;
  wire [0:0] h_arrdiv24_fs374_xor1;
  wire [0:0] h_arrdiv24_fs374_or0;
  wire [0:0] h_arrdiv24_fs375_xor1;
  wire [0:0] h_arrdiv24_fs375_or0;
  wire [0:0] h_arrdiv24_fs376_xor1;
  wire [0:0] h_arrdiv24_fs376_or0;
  wire [0:0] h_arrdiv24_fs377_xor1;
  wire [0:0] h_arrdiv24_fs377_or0;
  wire [0:0] h_arrdiv24_fs378_xor1;
  wire [0:0] h_arrdiv24_fs378_or0;
  wire [0:0] h_arrdiv24_fs379_xor1;
  wire [0:0] h_arrdiv24_fs379_or0;
  wire [0:0] h_arrdiv24_fs380_xor1;
  wire [0:0] h_arrdiv24_fs380_or0;
  wire [0:0] h_arrdiv24_fs381_xor1;
  wire [0:0] h_arrdiv24_fs381_or0;
  wire [0:0] h_arrdiv24_fs382_xor1;
  wire [0:0] h_arrdiv24_fs382_or0;
  wire [0:0] h_arrdiv24_fs383_xor1;
  wire [0:0] h_arrdiv24_fs383_or0;
  wire [0:0] h_arrdiv24_mux2to1345_xor0;
  wire [0:0] h_arrdiv24_mux2to1346_xor0;
  wire [0:0] h_arrdiv24_mux2to1347_xor0;
  wire [0:0] h_arrdiv24_mux2to1348_xor0;
  wire [0:0] h_arrdiv24_mux2to1349_xor0;
  wire [0:0] h_arrdiv24_mux2to1350_xor0;
  wire [0:0] h_arrdiv24_mux2to1351_xor0;
  wire [0:0] h_arrdiv24_mux2to1352_xor0;
  wire [0:0] h_arrdiv24_mux2to1353_xor0;
  wire [0:0] h_arrdiv24_mux2to1354_xor0;
  wire [0:0] h_arrdiv24_mux2to1355_xor0;
  wire [0:0] h_arrdiv24_mux2to1356_xor0;
  wire [0:0] h_arrdiv24_mux2to1357_xor0;
  wire [0:0] h_arrdiv24_mux2to1358_xor0;
  wire [0:0] h_arrdiv24_mux2to1359_xor0;
  wire [0:0] h_arrdiv24_mux2to1360_xor0;
  wire [0:0] h_arrdiv24_mux2to1361_xor0;
  wire [0:0] h_arrdiv24_mux2to1362_xor0;
  wire [0:0] h_arrdiv24_mux2to1363_xor0;
  wire [0:0] h_arrdiv24_mux2to1364_xor0;
  wire [0:0] h_arrdiv24_mux2to1365_xor0;
  wire [0:0] h_arrdiv24_mux2to1366_xor0;
  wire [0:0] h_arrdiv24_mux2to1367_xor0;
  wire [0:0] h_arrdiv24_not15;
  wire [0:0] h_arrdiv24_fs384_xor0;
  wire [0:0] h_arrdiv24_fs384_and0;
  wire [0:0] h_arrdiv24_fs385_xor1;
  wire [0:0] h_arrdiv24_fs385_or0;
  wire [0:0] h_arrdiv24_fs386_xor1;
  wire [0:0] h_arrdiv24_fs386_or0;
  wire [0:0] h_arrdiv24_fs387_xor1;
  wire [0:0] h_arrdiv24_fs387_or0;
  wire [0:0] h_arrdiv24_fs388_xor1;
  wire [0:0] h_arrdiv24_fs388_or0;
  wire [0:0] h_arrdiv24_fs389_xor1;
  wire [0:0] h_arrdiv24_fs389_or0;
  wire [0:0] h_arrdiv24_fs390_xor1;
  wire [0:0] h_arrdiv24_fs390_or0;
  wire [0:0] h_arrdiv24_fs391_xor1;
  wire [0:0] h_arrdiv24_fs391_or0;
  wire [0:0] h_arrdiv24_fs392_xor1;
  wire [0:0] h_arrdiv24_fs392_or0;
  wire [0:0] h_arrdiv24_fs393_xor1;
  wire [0:0] h_arrdiv24_fs393_or0;
  wire [0:0] h_arrdiv24_fs394_xor1;
  wire [0:0] h_arrdiv24_fs394_or0;
  wire [0:0] h_arrdiv24_fs395_xor1;
  wire [0:0] h_arrdiv24_fs395_or0;
  wire [0:0] h_arrdiv24_fs396_xor1;
  wire [0:0] h_arrdiv24_fs396_or0;
  wire [0:0] h_arrdiv24_fs397_xor1;
  wire [0:0] h_arrdiv24_fs397_or0;
  wire [0:0] h_arrdiv24_fs398_xor1;
  wire [0:0] h_arrdiv24_fs398_or0;
  wire [0:0] h_arrdiv24_fs399_xor1;
  wire [0:0] h_arrdiv24_fs399_or0;
  wire [0:0] h_arrdiv24_fs400_xor1;
  wire [0:0] h_arrdiv24_fs400_or0;
  wire [0:0] h_arrdiv24_fs401_xor1;
  wire [0:0] h_arrdiv24_fs401_or0;
  wire [0:0] h_arrdiv24_fs402_xor1;
  wire [0:0] h_arrdiv24_fs402_or0;
  wire [0:0] h_arrdiv24_fs403_xor1;
  wire [0:0] h_arrdiv24_fs403_or0;
  wire [0:0] h_arrdiv24_fs404_xor1;
  wire [0:0] h_arrdiv24_fs404_or0;
  wire [0:0] h_arrdiv24_fs405_xor1;
  wire [0:0] h_arrdiv24_fs405_or0;
  wire [0:0] h_arrdiv24_fs406_xor1;
  wire [0:0] h_arrdiv24_fs406_or0;
  wire [0:0] h_arrdiv24_fs407_xor1;
  wire [0:0] h_arrdiv24_fs407_or0;
  wire [0:0] h_arrdiv24_mux2to1368_xor0;
  wire [0:0] h_arrdiv24_mux2to1369_xor0;
  wire [0:0] h_arrdiv24_mux2to1370_xor0;
  wire [0:0] h_arrdiv24_mux2to1371_xor0;
  wire [0:0] h_arrdiv24_mux2to1372_xor0;
  wire [0:0] h_arrdiv24_mux2to1373_xor0;
  wire [0:0] h_arrdiv24_mux2to1374_xor0;
  wire [0:0] h_arrdiv24_mux2to1375_xor0;
  wire [0:0] h_arrdiv24_mux2to1376_xor0;
  wire [0:0] h_arrdiv24_mux2to1377_xor0;
  wire [0:0] h_arrdiv24_mux2to1378_xor0;
  wire [0:0] h_arrdiv24_mux2to1379_xor0;
  wire [0:0] h_arrdiv24_mux2to1380_xor0;
  wire [0:0] h_arrdiv24_mux2to1381_xor0;
  wire [0:0] h_arrdiv24_mux2to1382_xor0;
  wire [0:0] h_arrdiv24_mux2to1383_xor0;
  wire [0:0] h_arrdiv24_mux2to1384_xor0;
  wire [0:0] h_arrdiv24_mux2to1385_xor0;
  wire [0:0] h_arrdiv24_mux2to1386_xor0;
  wire [0:0] h_arrdiv24_mux2to1387_xor0;
  wire [0:0] h_arrdiv24_mux2to1388_xor0;
  wire [0:0] h_arrdiv24_mux2to1389_xor0;
  wire [0:0] h_arrdiv24_mux2to1390_xor0;
  wire [0:0] h_arrdiv24_not16;
  wire [0:0] h_arrdiv24_fs408_xor0;
  wire [0:0] h_arrdiv24_fs408_and0;
  wire [0:0] h_arrdiv24_fs409_xor1;
  wire [0:0] h_arrdiv24_fs409_or0;
  wire [0:0] h_arrdiv24_fs410_xor1;
  wire [0:0] h_arrdiv24_fs410_or0;
  wire [0:0] h_arrdiv24_fs411_xor1;
  wire [0:0] h_arrdiv24_fs411_or0;
  wire [0:0] h_arrdiv24_fs412_xor1;
  wire [0:0] h_arrdiv24_fs412_or0;
  wire [0:0] h_arrdiv24_fs413_xor1;
  wire [0:0] h_arrdiv24_fs413_or0;
  wire [0:0] h_arrdiv24_fs414_xor1;
  wire [0:0] h_arrdiv24_fs414_or0;
  wire [0:0] h_arrdiv24_fs415_xor1;
  wire [0:0] h_arrdiv24_fs415_or0;
  wire [0:0] h_arrdiv24_fs416_xor1;
  wire [0:0] h_arrdiv24_fs416_or0;
  wire [0:0] h_arrdiv24_fs417_xor1;
  wire [0:0] h_arrdiv24_fs417_or0;
  wire [0:0] h_arrdiv24_fs418_xor1;
  wire [0:0] h_arrdiv24_fs418_or0;
  wire [0:0] h_arrdiv24_fs419_xor1;
  wire [0:0] h_arrdiv24_fs419_or0;
  wire [0:0] h_arrdiv24_fs420_xor1;
  wire [0:0] h_arrdiv24_fs420_or0;
  wire [0:0] h_arrdiv24_fs421_xor1;
  wire [0:0] h_arrdiv24_fs421_or0;
  wire [0:0] h_arrdiv24_fs422_xor1;
  wire [0:0] h_arrdiv24_fs422_or0;
  wire [0:0] h_arrdiv24_fs423_xor1;
  wire [0:0] h_arrdiv24_fs423_or0;
  wire [0:0] h_arrdiv24_fs424_xor1;
  wire [0:0] h_arrdiv24_fs424_or0;
  wire [0:0] h_arrdiv24_fs425_xor1;
  wire [0:0] h_arrdiv24_fs425_or0;
  wire [0:0] h_arrdiv24_fs426_xor1;
  wire [0:0] h_arrdiv24_fs426_or0;
  wire [0:0] h_arrdiv24_fs427_xor1;
  wire [0:0] h_arrdiv24_fs427_or0;
  wire [0:0] h_arrdiv24_fs428_xor1;
  wire [0:0] h_arrdiv24_fs428_or0;
  wire [0:0] h_arrdiv24_fs429_xor1;
  wire [0:0] h_arrdiv24_fs429_or0;
  wire [0:0] h_arrdiv24_fs430_xor1;
  wire [0:0] h_arrdiv24_fs430_or0;
  wire [0:0] h_arrdiv24_fs431_xor1;
  wire [0:0] h_arrdiv24_fs431_or0;
  wire [0:0] h_arrdiv24_mux2to1391_xor0;
  wire [0:0] h_arrdiv24_mux2to1392_xor0;
  wire [0:0] h_arrdiv24_mux2to1393_xor0;
  wire [0:0] h_arrdiv24_mux2to1394_xor0;
  wire [0:0] h_arrdiv24_mux2to1395_xor0;
  wire [0:0] h_arrdiv24_mux2to1396_xor0;
  wire [0:0] h_arrdiv24_mux2to1397_xor0;
  wire [0:0] h_arrdiv24_mux2to1398_xor0;
  wire [0:0] h_arrdiv24_mux2to1399_xor0;
  wire [0:0] h_arrdiv24_mux2to1400_xor0;
  wire [0:0] h_arrdiv24_mux2to1401_xor0;
  wire [0:0] h_arrdiv24_mux2to1402_xor0;
  wire [0:0] h_arrdiv24_mux2to1403_xor0;
  wire [0:0] h_arrdiv24_mux2to1404_xor0;
  wire [0:0] h_arrdiv24_mux2to1405_xor0;
  wire [0:0] h_arrdiv24_mux2to1406_xor0;
  wire [0:0] h_arrdiv24_mux2to1407_xor0;
  wire [0:0] h_arrdiv24_mux2to1408_xor0;
  wire [0:0] h_arrdiv24_mux2to1409_xor0;
  wire [0:0] h_arrdiv24_mux2to1410_xor0;
  wire [0:0] h_arrdiv24_mux2to1411_xor0;
  wire [0:0] h_arrdiv24_mux2to1412_xor0;
  wire [0:0] h_arrdiv24_mux2to1413_xor0;
  wire [0:0] h_arrdiv24_not17;
  wire [0:0] h_arrdiv24_fs432_xor0;
  wire [0:0] h_arrdiv24_fs432_and0;
  wire [0:0] h_arrdiv24_fs433_xor1;
  wire [0:0] h_arrdiv24_fs433_or0;
  wire [0:0] h_arrdiv24_fs434_xor1;
  wire [0:0] h_arrdiv24_fs434_or0;
  wire [0:0] h_arrdiv24_fs435_xor1;
  wire [0:0] h_arrdiv24_fs435_or0;
  wire [0:0] h_arrdiv24_fs436_xor1;
  wire [0:0] h_arrdiv24_fs436_or0;
  wire [0:0] h_arrdiv24_fs437_xor1;
  wire [0:0] h_arrdiv24_fs437_or0;
  wire [0:0] h_arrdiv24_fs438_xor1;
  wire [0:0] h_arrdiv24_fs438_or0;
  wire [0:0] h_arrdiv24_fs439_xor1;
  wire [0:0] h_arrdiv24_fs439_or0;
  wire [0:0] h_arrdiv24_fs440_xor1;
  wire [0:0] h_arrdiv24_fs440_or0;
  wire [0:0] h_arrdiv24_fs441_xor1;
  wire [0:0] h_arrdiv24_fs441_or0;
  wire [0:0] h_arrdiv24_fs442_xor1;
  wire [0:0] h_arrdiv24_fs442_or0;
  wire [0:0] h_arrdiv24_fs443_xor1;
  wire [0:0] h_arrdiv24_fs443_or0;
  wire [0:0] h_arrdiv24_fs444_xor1;
  wire [0:0] h_arrdiv24_fs444_or0;
  wire [0:0] h_arrdiv24_fs445_xor1;
  wire [0:0] h_arrdiv24_fs445_or0;
  wire [0:0] h_arrdiv24_fs446_xor1;
  wire [0:0] h_arrdiv24_fs446_or0;
  wire [0:0] h_arrdiv24_fs447_xor1;
  wire [0:0] h_arrdiv24_fs447_or0;
  wire [0:0] h_arrdiv24_fs448_xor1;
  wire [0:0] h_arrdiv24_fs448_or0;
  wire [0:0] h_arrdiv24_fs449_xor1;
  wire [0:0] h_arrdiv24_fs449_or0;
  wire [0:0] h_arrdiv24_fs450_xor1;
  wire [0:0] h_arrdiv24_fs450_or0;
  wire [0:0] h_arrdiv24_fs451_xor1;
  wire [0:0] h_arrdiv24_fs451_or0;
  wire [0:0] h_arrdiv24_fs452_xor1;
  wire [0:0] h_arrdiv24_fs452_or0;
  wire [0:0] h_arrdiv24_fs453_xor1;
  wire [0:0] h_arrdiv24_fs453_or0;
  wire [0:0] h_arrdiv24_fs454_xor1;
  wire [0:0] h_arrdiv24_fs454_or0;
  wire [0:0] h_arrdiv24_fs455_xor1;
  wire [0:0] h_arrdiv24_fs455_or0;
  wire [0:0] h_arrdiv24_mux2to1414_xor0;
  wire [0:0] h_arrdiv24_mux2to1415_xor0;
  wire [0:0] h_arrdiv24_mux2to1416_xor0;
  wire [0:0] h_arrdiv24_mux2to1417_xor0;
  wire [0:0] h_arrdiv24_mux2to1418_xor0;
  wire [0:0] h_arrdiv24_mux2to1419_xor0;
  wire [0:0] h_arrdiv24_mux2to1420_xor0;
  wire [0:0] h_arrdiv24_mux2to1421_xor0;
  wire [0:0] h_arrdiv24_mux2to1422_xor0;
  wire [0:0] h_arrdiv24_mux2to1423_xor0;
  wire [0:0] h_arrdiv24_mux2to1424_xor0;
  wire [0:0] h_arrdiv24_mux2to1425_xor0;
  wire [0:0] h_arrdiv24_mux2to1426_xor0;
  wire [0:0] h_arrdiv24_mux2to1427_xor0;
  wire [0:0] h_arrdiv24_mux2to1428_xor0;
  wire [0:0] h_arrdiv24_mux2to1429_xor0;
  wire [0:0] h_arrdiv24_mux2to1430_xor0;
  wire [0:0] h_arrdiv24_mux2to1431_xor0;
  wire [0:0] h_arrdiv24_mux2to1432_xor0;
  wire [0:0] h_arrdiv24_mux2to1433_xor0;
  wire [0:0] h_arrdiv24_mux2to1434_xor0;
  wire [0:0] h_arrdiv24_mux2to1435_xor0;
  wire [0:0] h_arrdiv24_mux2to1436_xor0;
  wire [0:0] h_arrdiv24_not18;
  wire [0:0] h_arrdiv24_fs456_xor0;
  wire [0:0] h_arrdiv24_fs456_and0;
  wire [0:0] h_arrdiv24_fs457_xor1;
  wire [0:0] h_arrdiv24_fs457_or0;
  wire [0:0] h_arrdiv24_fs458_xor1;
  wire [0:0] h_arrdiv24_fs458_or0;
  wire [0:0] h_arrdiv24_fs459_xor1;
  wire [0:0] h_arrdiv24_fs459_or0;
  wire [0:0] h_arrdiv24_fs460_xor1;
  wire [0:0] h_arrdiv24_fs460_or0;
  wire [0:0] h_arrdiv24_fs461_xor1;
  wire [0:0] h_arrdiv24_fs461_or0;
  wire [0:0] h_arrdiv24_fs462_xor1;
  wire [0:0] h_arrdiv24_fs462_or0;
  wire [0:0] h_arrdiv24_fs463_xor1;
  wire [0:0] h_arrdiv24_fs463_or0;
  wire [0:0] h_arrdiv24_fs464_xor1;
  wire [0:0] h_arrdiv24_fs464_or0;
  wire [0:0] h_arrdiv24_fs465_xor1;
  wire [0:0] h_arrdiv24_fs465_or0;
  wire [0:0] h_arrdiv24_fs466_xor1;
  wire [0:0] h_arrdiv24_fs466_or0;
  wire [0:0] h_arrdiv24_fs467_xor1;
  wire [0:0] h_arrdiv24_fs467_or0;
  wire [0:0] h_arrdiv24_fs468_xor1;
  wire [0:0] h_arrdiv24_fs468_or0;
  wire [0:0] h_arrdiv24_fs469_xor1;
  wire [0:0] h_arrdiv24_fs469_or0;
  wire [0:0] h_arrdiv24_fs470_xor1;
  wire [0:0] h_arrdiv24_fs470_or0;
  wire [0:0] h_arrdiv24_fs471_xor1;
  wire [0:0] h_arrdiv24_fs471_or0;
  wire [0:0] h_arrdiv24_fs472_xor1;
  wire [0:0] h_arrdiv24_fs472_or0;
  wire [0:0] h_arrdiv24_fs473_xor1;
  wire [0:0] h_arrdiv24_fs473_or0;
  wire [0:0] h_arrdiv24_fs474_xor1;
  wire [0:0] h_arrdiv24_fs474_or0;
  wire [0:0] h_arrdiv24_fs475_xor1;
  wire [0:0] h_arrdiv24_fs475_or0;
  wire [0:0] h_arrdiv24_fs476_xor1;
  wire [0:0] h_arrdiv24_fs476_or0;
  wire [0:0] h_arrdiv24_fs477_xor1;
  wire [0:0] h_arrdiv24_fs477_or0;
  wire [0:0] h_arrdiv24_fs478_xor1;
  wire [0:0] h_arrdiv24_fs478_or0;
  wire [0:0] h_arrdiv24_fs479_xor1;
  wire [0:0] h_arrdiv24_fs479_or0;
  wire [0:0] h_arrdiv24_mux2to1437_xor0;
  wire [0:0] h_arrdiv24_mux2to1438_xor0;
  wire [0:0] h_arrdiv24_mux2to1439_xor0;
  wire [0:0] h_arrdiv24_mux2to1440_xor0;
  wire [0:0] h_arrdiv24_mux2to1441_xor0;
  wire [0:0] h_arrdiv24_mux2to1442_xor0;
  wire [0:0] h_arrdiv24_mux2to1443_xor0;
  wire [0:0] h_arrdiv24_mux2to1444_xor0;
  wire [0:0] h_arrdiv24_mux2to1445_xor0;
  wire [0:0] h_arrdiv24_mux2to1446_xor0;
  wire [0:0] h_arrdiv24_mux2to1447_xor0;
  wire [0:0] h_arrdiv24_mux2to1448_xor0;
  wire [0:0] h_arrdiv24_mux2to1449_xor0;
  wire [0:0] h_arrdiv24_mux2to1450_xor0;
  wire [0:0] h_arrdiv24_mux2to1451_xor0;
  wire [0:0] h_arrdiv24_mux2to1452_xor0;
  wire [0:0] h_arrdiv24_mux2to1453_xor0;
  wire [0:0] h_arrdiv24_mux2to1454_xor0;
  wire [0:0] h_arrdiv24_mux2to1455_xor0;
  wire [0:0] h_arrdiv24_mux2to1456_xor0;
  wire [0:0] h_arrdiv24_mux2to1457_xor0;
  wire [0:0] h_arrdiv24_mux2to1458_xor0;
  wire [0:0] h_arrdiv24_mux2to1459_xor0;
  wire [0:0] h_arrdiv24_not19;
  wire [0:0] h_arrdiv24_fs480_xor0;
  wire [0:0] h_arrdiv24_fs480_and0;
  wire [0:0] h_arrdiv24_fs481_xor1;
  wire [0:0] h_arrdiv24_fs481_or0;
  wire [0:0] h_arrdiv24_fs482_xor1;
  wire [0:0] h_arrdiv24_fs482_or0;
  wire [0:0] h_arrdiv24_fs483_xor1;
  wire [0:0] h_arrdiv24_fs483_or0;
  wire [0:0] h_arrdiv24_fs484_xor1;
  wire [0:0] h_arrdiv24_fs484_or0;
  wire [0:0] h_arrdiv24_fs485_xor1;
  wire [0:0] h_arrdiv24_fs485_or0;
  wire [0:0] h_arrdiv24_fs486_xor1;
  wire [0:0] h_arrdiv24_fs486_or0;
  wire [0:0] h_arrdiv24_fs487_xor1;
  wire [0:0] h_arrdiv24_fs487_or0;
  wire [0:0] h_arrdiv24_fs488_xor1;
  wire [0:0] h_arrdiv24_fs488_or0;
  wire [0:0] h_arrdiv24_fs489_xor1;
  wire [0:0] h_arrdiv24_fs489_or0;
  wire [0:0] h_arrdiv24_fs490_xor1;
  wire [0:0] h_arrdiv24_fs490_or0;
  wire [0:0] h_arrdiv24_fs491_xor1;
  wire [0:0] h_arrdiv24_fs491_or0;
  wire [0:0] h_arrdiv24_fs492_xor1;
  wire [0:0] h_arrdiv24_fs492_or0;
  wire [0:0] h_arrdiv24_fs493_xor1;
  wire [0:0] h_arrdiv24_fs493_or0;
  wire [0:0] h_arrdiv24_fs494_xor1;
  wire [0:0] h_arrdiv24_fs494_or0;
  wire [0:0] h_arrdiv24_fs495_xor1;
  wire [0:0] h_arrdiv24_fs495_or0;
  wire [0:0] h_arrdiv24_fs496_xor1;
  wire [0:0] h_arrdiv24_fs496_or0;
  wire [0:0] h_arrdiv24_fs497_xor1;
  wire [0:0] h_arrdiv24_fs497_or0;
  wire [0:0] h_arrdiv24_fs498_xor1;
  wire [0:0] h_arrdiv24_fs498_or0;
  wire [0:0] h_arrdiv24_fs499_xor1;
  wire [0:0] h_arrdiv24_fs499_or0;
  wire [0:0] h_arrdiv24_fs500_xor1;
  wire [0:0] h_arrdiv24_fs500_or0;
  wire [0:0] h_arrdiv24_fs501_xor1;
  wire [0:0] h_arrdiv24_fs501_or0;
  wire [0:0] h_arrdiv24_fs502_xor1;
  wire [0:0] h_arrdiv24_fs502_or0;
  wire [0:0] h_arrdiv24_fs503_xor1;
  wire [0:0] h_arrdiv24_fs503_or0;
  wire [0:0] h_arrdiv24_mux2to1460_xor0;
  wire [0:0] h_arrdiv24_mux2to1461_xor0;
  wire [0:0] h_arrdiv24_mux2to1462_xor0;
  wire [0:0] h_arrdiv24_mux2to1463_xor0;
  wire [0:0] h_arrdiv24_mux2to1464_xor0;
  wire [0:0] h_arrdiv24_mux2to1465_xor0;
  wire [0:0] h_arrdiv24_mux2to1466_xor0;
  wire [0:0] h_arrdiv24_mux2to1467_xor0;
  wire [0:0] h_arrdiv24_mux2to1468_xor0;
  wire [0:0] h_arrdiv24_mux2to1469_xor0;
  wire [0:0] h_arrdiv24_mux2to1470_xor0;
  wire [0:0] h_arrdiv24_mux2to1471_xor0;
  wire [0:0] h_arrdiv24_mux2to1472_xor0;
  wire [0:0] h_arrdiv24_mux2to1473_xor0;
  wire [0:0] h_arrdiv24_mux2to1474_xor0;
  wire [0:0] h_arrdiv24_mux2to1475_xor0;
  wire [0:0] h_arrdiv24_mux2to1476_xor0;
  wire [0:0] h_arrdiv24_mux2to1477_xor0;
  wire [0:0] h_arrdiv24_mux2to1478_xor0;
  wire [0:0] h_arrdiv24_mux2to1479_xor0;
  wire [0:0] h_arrdiv24_mux2to1480_xor0;
  wire [0:0] h_arrdiv24_mux2to1481_xor0;
  wire [0:0] h_arrdiv24_mux2to1482_xor0;
  wire [0:0] h_arrdiv24_not20;
  wire [0:0] h_arrdiv24_fs504_xor0;
  wire [0:0] h_arrdiv24_fs504_and0;
  wire [0:0] h_arrdiv24_fs505_xor1;
  wire [0:0] h_arrdiv24_fs505_or0;
  wire [0:0] h_arrdiv24_fs506_xor1;
  wire [0:0] h_arrdiv24_fs506_or0;
  wire [0:0] h_arrdiv24_fs507_xor1;
  wire [0:0] h_arrdiv24_fs507_or0;
  wire [0:0] h_arrdiv24_fs508_xor1;
  wire [0:0] h_arrdiv24_fs508_or0;
  wire [0:0] h_arrdiv24_fs509_xor1;
  wire [0:0] h_arrdiv24_fs509_or0;
  wire [0:0] h_arrdiv24_fs510_xor1;
  wire [0:0] h_arrdiv24_fs510_or0;
  wire [0:0] h_arrdiv24_fs511_xor1;
  wire [0:0] h_arrdiv24_fs511_or0;
  wire [0:0] h_arrdiv24_fs512_xor1;
  wire [0:0] h_arrdiv24_fs512_or0;
  wire [0:0] h_arrdiv24_fs513_xor1;
  wire [0:0] h_arrdiv24_fs513_or0;
  wire [0:0] h_arrdiv24_fs514_xor1;
  wire [0:0] h_arrdiv24_fs514_or0;
  wire [0:0] h_arrdiv24_fs515_xor1;
  wire [0:0] h_arrdiv24_fs515_or0;
  wire [0:0] h_arrdiv24_fs516_xor1;
  wire [0:0] h_arrdiv24_fs516_or0;
  wire [0:0] h_arrdiv24_fs517_xor1;
  wire [0:0] h_arrdiv24_fs517_or0;
  wire [0:0] h_arrdiv24_fs518_xor1;
  wire [0:0] h_arrdiv24_fs518_or0;
  wire [0:0] h_arrdiv24_fs519_xor1;
  wire [0:0] h_arrdiv24_fs519_or0;
  wire [0:0] h_arrdiv24_fs520_xor1;
  wire [0:0] h_arrdiv24_fs520_or0;
  wire [0:0] h_arrdiv24_fs521_xor1;
  wire [0:0] h_arrdiv24_fs521_or0;
  wire [0:0] h_arrdiv24_fs522_xor1;
  wire [0:0] h_arrdiv24_fs522_or0;
  wire [0:0] h_arrdiv24_fs523_xor1;
  wire [0:0] h_arrdiv24_fs523_or0;
  wire [0:0] h_arrdiv24_fs524_xor1;
  wire [0:0] h_arrdiv24_fs524_or0;
  wire [0:0] h_arrdiv24_fs525_xor1;
  wire [0:0] h_arrdiv24_fs525_or0;
  wire [0:0] h_arrdiv24_fs526_xor1;
  wire [0:0] h_arrdiv24_fs526_or0;
  wire [0:0] h_arrdiv24_fs527_xor1;
  wire [0:0] h_arrdiv24_fs527_or0;
  wire [0:0] h_arrdiv24_mux2to1483_xor0;
  wire [0:0] h_arrdiv24_mux2to1484_xor0;
  wire [0:0] h_arrdiv24_mux2to1485_xor0;
  wire [0:0] h_arrdiv24_mux2to1486_xor0;
  wire [0:0] h_arrdiv24_mux2to1487_xor0;
  wire [0:0] h_arrdiv24_mux2to1488_xor0;
  wire [0:0] h_arrdiv24_mux2to1489_xor0;
  wire [0:0] h_arrdiv24_mux2to1490_xor0;
  wire [0:0] h_arrdiv24_mux2to1491_xor0;
  wire [0:0] h_arrdiv24_mux2to1492_xor0;
  wire [0:0] h_arrdiv24_mux2to1493_xor0;
  wire [0:0] h_arrdiv24_mux2to1494_xor0;
  wire [0:0] h_arrdiv24_mux2to1495_xor0;
  wire [0:0] h_arrdiv24_mux2to1496_xor0;
  wire [0:0] h_arrdiv24_mux2to1497_xor0;
  wire [0:0] h_arrdiv24_mux2to1498_xor0;
  wire [0:0] h_arrdiv24_mux2to1499_xor0;
  wire [0:0] h_arrdiv24_mux2to1500_xor0;
  wire [0:0] h_arrdiv24_mux2to1501_xor0;
  wire [0:0] h_arrdiv24_mux2to1502_xor0;
  wire [0:0] h_arrdiv24_mux2to1503_xor0;
  wire [0:0] h_arrdiv24_mux2to1504_xor0;
  wire [0:0] h_arrdiv24_mux2to1505_xor0;
  wire [0:0] h_arrdiv24_not21;
  wire [0:0] h_arrdiv24_fs528_xor0;
  wire [0:0] h_arrdiv24_fs528_and0;
  wire [0:0] h_arrdiv24_fs529_xor1;
  wire [0:0] h_arrdiv24_fs529_or0;
  wire [0:0] h_arrdiv24_fs530_xor1;
  wire [0:0] h_arrdiv24_fs530_or0;
  wire [0:0] h_arrdiv24_fs531_xor1;
  wire [0:0] h_arrdiv24_fs531_or0;
  wire [0:0] h_arrdiv24_fs532_xor1;
  wire [0:0] h_arrdiv24_fs532_or0;
  wire [0:0] h_arrdiv24_fs533_xor1;
  wire [0:0] h_arrdiv24_fs533_or0;
  wire [0:0] h_arrdiv24_fs534_xor1;
  wire [0:0] h_arrdiv24_fs534_or0;
  wire [0:0] h_arrdiv24_fs535_xor1;
  wire [0:0] h_arrdiv24_fs535_or0;
  wire [0:0] h_arrdiv24_fs536_xor1;
  wire [0:0] h_arrdiv24_fs536_or0;
  wire [0:0] h_arrdiv24_fs537_xor1;
  wire [0:0] h_arrdiv24_fs537_or0;
  wire [0:0] h_arrdiv24_fs538_xor1;
  wire [0:0] h_arrdiv24_fs538_or0;
  wire [0:0] h_arrdiv24_fs539_xor1;
  wire [0:0] h_arrdiv24_fs539_or0;
  wire [0:0] h_arrdiv24_fs540_xor1;
  wire [0:0] h_arrdiv24_fs540_or0;
  wire [0:0] h_arrdiv24_fs541_xor1;
  wire [0:0] h_arrdiv24_fs541_or0;
  wire [0:0] h_arrdiv24_fs542_xor1;
  wire [0:0] h_arrdiv24_fs542_or0;
  wire [0:0] h_arrdiv24_fs543_xor1;
  wire [0:0] h_arrdiv24_fs543_or0;
  wire [0:0] h_arrdiv24_fs544_xor1;
  wire [0:0] h_arrdiv24_fs544_or0;
  wire [0:0] h_arrdiv24_fs545_xor1;
  wire [0:0] h_arrdiv24_fs545_or0;
  wire [0:0] h_arrdiv24_fs546_xor1;
  wire [0:0] h_arrdiv24_fs546_or0;
  wire [0:0] h_arrdiv24_fs547_xor1;
  wire [0:0] h_arrdiv24_fs547_or0;
  wire [0:0] h_arrdiv24_fs548_xor1;
  wire [0:0] h_arrdiv24_fs548_or0;
  wire [0:0] h_arrdiv24_fs549_xor1;
  wire [0:0] h_arrdiv24_fs549_or0;
  wire [0:0] h_arrdiv24_fs550_xor1;
  wire [0:0] h_arrdiv24_fs550_or0;
  wire [0:0] h_arrdiv24_fs551_xor1;
  wire [0:0] h_arrdiv24_fs551_or0;
  wire [0:0] h_arrdiv24_mux2to1506_xor0;
  wire [0:0] h_arrdiv24_mux2to1507_xor0;
  wire [0:0] h_arrdiv24_mux2to1508_xor0;
  wire [0:0] h_arrdiv24_mux2to1509_xor0;
  wire [0:0] h_arrdiv24_mux2to1510_xor0;
  wire [0:0] h_arrdiv24_mux2to1511_xor0;
  wire [0:0] h_arrdiv24_mux2to1512_xor0;
  wire [0:0] h_arrdiv24_mux2to1513_xor0;
  wire [0:0] h_arrdiv24_mux2to1514_xor0;
  wire [0:0] h_arrdiv24_mux2to1515_xor0;
  wire [0:0] h_arrdiv24_mux2to1516_xor0;
  wire [0:0] h_arrdiv24_mux2to1517_xor0;
  wire [0:0] h_arrdiv24_mux2to1518_xor0;
  wire [0:0] h_arrdiv24_mux2to1519_xor0;
  wire [0:0] h_arrdiv24_mux2to1520_xor0;
  wire [0:0] h_arrdiv24_mux2to1521_xor0;
  wire [0:0] h_arrdiv24_mux2to1522_xor0;
  wire [0:0] h_arrdiv24_mux2to1523_xor0;
  wire [0:0] h_arrdiv24_mux2to1524_xor0;
  wire [0:0] h_arrdiv24_mux2to1525_xor0;
  wire [0:0] h_arrdiv24_mux2to1526_xor0;
  wire [0:0] h_arrdiv24_mux2to1527_xor0;
  wire [0:0] h_arrdiv24_mux2to1528_xor0;
  wire [0:0] h_arrdiv24_not22;
  wire [0:0] h_arrdiv24_fs552_xor0;
  wire [0:0] h_arrdiv24_fs552_and0;
  wire [0:0] h_arrdiv24_fs553_xor1;
  wire [0:0] h_arrdiv24_fs553_or0;
  wire [0:0] h_arrdiv24_fs554_xor1;
  wire [0:0] h_arrdiv24_fs554_or0;
  wire [0:0] h_arrdiv24_fs555_xor1;
  wire [0:0] h_arrdiv24_fs555_or0;
  wire [0:0] h_arrdiv24_fs556_xor1;
  wire [0:0] h_arrdiv24_fs556_or0;
  wire [0:0] h_arrdiv24_fs557_xor1;
  wire [0:0] h_arrdiv24_fs557_or0;
  wire [0:0] h_arrdiv24_fs558_xor1;
  wire [0:0] h_arrdiv24_fs558_or0;
  wire [0:0] h_arrdiv24_fs559_xor1;
  wire [0:0] h_arrdiv24_fs559_or0;
  wire [0:0] h_arrdiv24_fs560_xor1;
  wire [0:0] h_arrdiv24_fs560_or0;
  wire [0:0] h_arrdiv24_fs561_xor1;
  wire [0:0] h_arrdiv24_fs561_or0;
  wire [0:0] h_arrdiv24_fs562_xor1;
  wire [0:0] h_arrdiv24_fs562_or0;
  wire [0:0] h_arrdiv24_fs563_xor1;
  wire [0:0] h_arrdiv24_fs563_or0;
  wire [0:0] h_arrdiv24_fs564_xor1;
  wire [0:0] h_arrdiv24_fs564_or0;
  wire [0:0] h_arrdiv24_fs565_xor1;
  wire [0:0] h_arrdiv24_fs565_or0;
  wire [0:0] h_arrdiv24_fs566_xor1;
  wire [0:0] h_arrdiv24_fs566_or0;
  wire [0:0] h_arrdiv24_fs567_xor1;
  wire [0:0] h_arrdiv24_fs567_or0;
  wire [0:0] h_arrdiv24_fs568_xor1;
  wire [0:0] h_arrdiv24_fs568_or0;
  wire [0:0] h_arrdiv24_fs569_xor1;
  wire [0:0] h_arrdiv24_fs569_or0;
  wire [0:0] h_arrdiv24_fs570_xor1;
  wire [0:0] h_arrdiv24_fs570_or0;
  wire [0:0] h_arrdiv24_fs571_xor1;
  wire [0:0] h_arrdiv24_fs571_or0;
  wire [0:0] h_arrdiv24_fs572_xor1;
  wire [0:0] h_arrdiv24_fs572_or0;
  wire [0:0] h_arrdiv24_fs573_xor1;
  wire [0:0] h_arrdiv24_fs573_or0;
  wire [0:0] h_arrdiv24_fs574_xor1;
  wire [0:0] h_arrdiv24_fs574_or0;
  wire [0:0] h_arrdiv24_fs575_xor1;
  wire [0:0] h_arrdiv24_fs575_or0;
  wire [0:0] h_arrdiv24_not23;

  fs fs_h_arrdiv24_fs0_out(.a(a[23]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs0_xor0), .fs_or0(h_arrdiv24_fs0_and0));
  fs fs_h_arrdiv24_fs1_out(.a(1'b0), .b(b[1]), .bin(h_arrdiv24_fs0_and0[0]), .fs_xor1(h_arrdiv24_fs1_xor1), .fs_or0(h_arrdiv24_fs1_or0));
  fs fs_h_arrdiv24_fs2_out(.a(1'b0), .b(b[2]), .bin(h_arrdiv24_fs1_or0[0]), .fs_xor1(h_arrdiv24_fs2_xor1), .fs_or0(h_arrdiv24_fs2_or0));
  fs fs_h_arrdiv24_fs3_out(.a(1'b0), .b(b[3]), .bin(h_arrdiv24_fs2_or0[0]), .fs_xor1(h_arrdiv24_fs3_xor1), .fs_or0(h_arrdiv24_fs3_or0));
  fs fs_h_arrdiv24_fs4_out(.a(1'b0), .b(b[4]), .bin(h_arrdiv24_fs3_or0[0]), .fs_xor1(h_arrdiv24_fs4_xor1), .fs_or0(h_arrdiv24_fs4_or0));
  fs fs_h_arrdiv24_fs5_out(.a(1'b0), .b(b[5]), .bin(h_arrdiv24_fs4_or0[0]), .fs_xor1(h_arrdiv24_fs5_xor1), .fs_or0(h_arrdiv24_fs5_or0));
  fs fs_h_arrdiv24_fs6_out(.a(1'b0), .b(b[6]), .bin(h_arrdiv24_fs5_or0[0]), .fs_xor1(h_arrdiv24_fs6_xor1), .fs_or0(h_arrdiv24_fs6_or0));
  fs fs_h_arrdiv24_fs7_out(.a(1'b0), .b(b[7]), .bin(h_arrdiv24_fs6_or0[0]), .fs_xor1(h_arrdiv24_fs7_xor1), .fs_or0(h_arrdiv24_fs7_or0));
  fs fs_h_arrdiv24_fs8_out(.a(1'b0), .b(b[8]), .bin(h_arrdiv24_fs7_or0[0]), .fs_xor1(h_arrdiv24_fs8_xor1), .fs_or0(h_arrdiv24_fs8_or0));
  fs fs_h_arrdiv24_fs9_out(.a(1'b0), .b(b[9]), .bin(h_arrdiv24_fs8_or0[0]), .fs_xor1(h_arrdiv24_fs9_xor1), .fs_or0(h_arrdiv24_fs9_or0));
  fs fs_h_arrdiv24_fs10_out(.a(1'b0), .b(b[10]), .bin(h_arrdiv24_fs9_or0[0]), .fs_xor1(h_arrdiv24_fs10_xor1), .fs_or0(h_arrdiv24_fs10_or0));
  fs fs_h_arrdiv24_fs11_out(.a(1'b0), .b(b[11]), .bin(h_arrdiv24_fs10_or0[0]), .fs_xor1(h_arrdiv24_fs11_xor1), .fs_or0(h_arrdiv24_fs11_or0));
  fs fs_h_arrdiv24_fs12_out(.a(1'b0), .b(b[12]), .bin(h_arrdiv24_fs11_or0[0]), .fs_xor1(h_arrdiv24_fs12_xor1), .fs_or0(h_arrdiv24_fs12_or0));
  fs fs_h_arrdiv24_fs13_out(.a(1'b0), .b(b[13]), .bin(h_arrdiv24_fs12_or0[0]), .fs_xor1(h_arrdiv24_fs13_xor1), .fs_or0(h_arrdiv24_fs13_or0));
  fs fs_h_arrdiv24_fs14_out(.a(1'b0), .b(b[14]), .bin(h_arrdiv24_fs13_or0[0]), .fs_xor1(h_arrdiv24_fs14_xor1), .fs_or0(h_arrdiv24_fs14_or0));
  fs fs_h_arrdiv24_fs15_out(.a(1'b0), .b(b[15]), .bin(h_arrdiv24_fs14_or0[0]), .fs_xor1(h_arrdiv24_fs15_xor1), .fs_or0(h_arrdiv24_fs15_or0));
  fs fs_h_arrdiv24_fs16_out(.a(1'b0), .b(b[16]), .bin(h_arrdiv24_fs15_or0[0]), .fs_xor1(h_arrdiv24_fs16_xor1), .fs_or0(h_arrdiv24_fs16_or0));
  fs fs_h_arrdiv24_fs17_out(.a(1'b0), .b(b[17]), .bin(h_arrdiv24_fs16_or0[0]), .fs_xor1(h_arrdiv24_fs17_xor1), .fs_or0(h_arrdiv24_fs17_or0));
  fs fs_h_arrdiv24_fs18_out(.a(1'b0), .b(b[18]), .bin(h_arrdiv24_fs17_or0[0]), .fs_xor1(h_arrdiv24_fs18_xor1), .fs_or0(h_arrdiv24_fs18_or0));
  fs fs_h_arrdiv24_fs19_out(.a(1'b0), .b(b[19]), .bin(h_arrdiv24_fs18_or0[0]), .fs_xor1(h_arrdiv24_fs19_xor1), .fs_or0(h_arrdiv24_fs19_or0));
  fs fs_h_arrdiv24_fs20_out(.a(1'b0), .b(b[20]), .bin(h_arrdiv24_fs19_or0[0]), .fs_xor1(h_arrdiv24_fs20_xor1), .fs_or0(h_arrdiv24_fs20_or0));
  fs fs_h_arrdiv24_fs21_out(.a(1'b0), .b(b[21]), .bin(h_arrdiv24_fs20_or0[0]), .fs_xor1(h_arrdiv24_fs21_xor1), .fs_or0(h_arrdiv24_fs21_or0));
  fs fs_h_arrdiv24_fs22_out(.a(1'b0), .b(b[22]), .bin(h_arrdiv24_fs21_or0[0]), .fs_xor1(h_arrdiv24_fs22_xor1), .fs_or0(h_arrdiv24_fs22_or0));
  fs fs_h_arrdiv24_fs23_out(.a(1'b0), .b(b[23]), .bin(h_arrdiv24_fs22_or0[0]), .fs_xor1(h_arrdiv24_fs23_xor1), .fs_or0(h_arrdiv24_fs23_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to10_out(.d0(h_arrdiv24_fs0_xor0[0]), .d1(a[23]), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to10_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to11_out(.d0(h_arrdiv24_fs1_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to11_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to12_out(.d0(h_arrdiv24_fs2_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to12_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to13_out(.d0(h_arrdiv24_fs3_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to13_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to14_out(.d0(h_arrdiv24_fs4_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to14_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to15_out(.d0(h_arrdiv24_fs5_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to15_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to16_out(.d0(h_arrdiv24_fs6_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to16_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to17_out(.d0(h_arrdiv24_fs7_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to17_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to18_out(.d0(h_arrdiv24_fs8_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to18_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to19_out(.d0(h_arrdiv24_fs9_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to19_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to110_out(.d0(h_arrdiv24_fs10_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to110_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to111_out(.d0(h_arrdiv24_fs11_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to111_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to112_out(.d0(h_arrdiv24_fs12_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to112_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to113_out(.d0(h_arrdiv24_fs13_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to113_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to114_out(.d0(h_arrdiv24_fs14_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to114_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to115_out(.d0(h_arrdiv24_fs15_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to115_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to116_out(.d0(h_arrdiv24_fs16_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to116_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to117_out(.d0(h_arrdiv24_fs17_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to117_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to118_out(.d0(h_arrdiv24_fs18_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to118_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to119_out(.d0(h_arrdiv24_fs19_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to119_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to120_out(.d0(h_arrdiv24_fs20_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to120_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to121_out(.d0(h_arrdiv24_fs21_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to121_and1));
  mux2to1 mux2to1_h_arrdiv24_mux2to122_out(.d0(h_arrdiv24_fs22_xor1[0]), .d1(1'b0), .sel(h_arrdiv24_fs23_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to122_and1));
  not_gate not_gate_h_arrdiv24_not0(.a(h_arrdiv24_fs23_or0[0]), .out(h_arrdiv24_not0));
  fs fs_h_arrdiv24_fs24_out(.a(a[22]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs24_xor0), .fs_or0(h_arrdiv24_fs24_and0));
  fs fs_h_arrdiv24_fs25_out(.a(h_arrdiv24_mux2to10_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs24_and0[0]), .fs_xor1(h_arrdiv24_fs25_xor1), .fs_or0(h_arrdiv24_fs25_or0));
  fs fs_h_arrdiv24_fs26_out(.a(h_arrdiv24_mux2to11_and1[0]), .b(b[2]), .bin(h_arrdiv24_fs25_or0[0]), .fs_xor1(h_arrdiv24_fs26_xor1), .fs_or0(h_arrdiv24_fs26_or0));
  fs fs_h_arrdiv24_fs27_out(.a(h_arrdiv24_mux2to12_and1[0]), .b(b[3]), .bin(h_arrdiv24_fs26_or0[0]), .fs_xor1(h_arrdiv24_fs27_xor1), .fs_or0(h_arrdiv24_fs27_or0));
  fs fs_h_arrdiv24_fs28_out(.a(h_arrdiv24_mux2to13_and1[0]), .b(b[4]), .bin(h_arrdiv24_fs27_or0[0]), .fs_xor1(h_arrdiv24_fs28_xor1), .fs_or0(h_arrdiv24_fs28_or0));
  fs fs_h_arrdiv24_fs29_out(.a(h_arrdiv24_mux2to14_and1[0]), .b(b[5]), .bin(h_arrdiv24_fs28_or0[0]), .fs_xor1(h_arrdiv24_fs29_xor1), .fs_or0(h_arrdiv24_fs29_or0));
  fs fs_h_arrdiv24_fs30_out(.a(h_arrdiv24_mux2to15_and1[0]), .b(b[6]), .bin(h_arrdiv24_fs29_or0[0]), .fs_xor1(h_arrdiv24_fs30_xor1), .fs_or0(h_arrdiv24_fs30_or0));
  fs fs_h_arrdiv24_fs31_out(.a(h_arrdiv24_mux2to16_and1[0]), .b(b[7]), .bin(h_arrdiv24_fs30_or0[0]), .fs_xor1(h_arrdiv24_fs31_xor1), .fs_or0(h_arrdiv24_fs31_or0));
  fs fs_h_arrdiv24_fs32_out(.a(h_arrdiv24_mux2to17_and1[0]), .b(b[8]), .bin(h_arrdiv24_fs31_or0[0]), .fs_xor1(h_arrdiv24_fs32_xor1), .fs_or0(h_arrdiv24_fs32_or0));
  fs fs_h_arrdiv24_fs33_out(.a(h_arrdiv24_mux2to18_and1[0]), .b(b[9]), .bin(h_arrdiv24_fs32_or0[0]), .fs_xor1(h_arrdiv24_fs33_xor1), .fs_or0(h_arrdiv24_fs33_or0));
  fs fs_h_arrdiv24_fs34_out(.a(h_arrdiv24_mux2to19_and1[0]), .b(b[10]), .bin(h_arrdiv24_fs33_or0[0]), .fs_xor1(h_arrdiv24_fs34_xor1), .fs_or0(h_arrdiv24_fs34_or0));
  fs fs_h_arrdiv24_fs35_out(.a(h_arrdiv24_mux2to110_and1[0]), .b(b[11]), .bin(h_arrdiv24_fs34_or0[0]), .fs_xor1(h_arrdiv24_fs35_xor1), .fs_or0(h_arrdiv24_fs35_or0));
  fs fs_h_arrdiv24_fs36_out(.a(h_arrdiv24_mux2to111_and1[0]), .b(b[12]), .bin(h_arrdiv24_fs35_or0[0]), .fs_xor1(h_arrdiv24_fs36_xor1), .fs_or0(h_arrdiv24_fs36_or0));
  fs fs_h_arrdiv24_fs37_out(.a(h_arrdiv24_mux2to112_and1[0]), .b(b[13]), .bin(h_arrdiv24_fs36_or0[0]), .fs_xor1(h_arrdiv24_fs37_xor1), .fs_or0(h_arrdiv24_fs37_or0));
  fs fs_h_arrdiv24_fs38_out(.a(h_arrdiv24_mux2to113_and1[0]), .b(b[14]), .bin(h_arrdiv24_fs37_or0[0]), .fs_xor1(h_arrdiv24_fs38_xor1), .fs_or0(h_arrdiv24_fs38_or0));
  fs fs_h_arrdiv24_fs39_out(.a(h_arrdiv24_mux2to114_and1[0]), .b(b[15]), .bin(h_arrdiv24_fs38_or0[0]), .fs_xor1(h_arrdiv24_fs39_xor1), .fs_or0(h_arrdiv24_fs39_or0));
  fs fs_h_arrdiv24_fs40_out(.a(h_arrdiv24_mux2to115_and1[0]), .b(b[16]), .bin(h_arrdiv24_fs39_or0[0]), .fs_xor1(h_arrdiv24_fs40_xor1), .fs_or0(h_arrdiv24_fs40_or0));
  fs fs_h_arrdiv24_fs41_out(.a(h_arrdiv24_mux2to116_and1[0]), .b(b[17]), .bin(h_arrdiv24_fs40_or0[0]), .fs_xor1(h_arrdiv24_fs41_xor1), .fs_or0(h_arrdiv24_fs41_or0));
  fs fs_h_arrdiv24_fs42_out(.a(h_arrdiv24_mux2to117_and1[0]), .b(b[18]), .bin(h_arrdiv24_fs41_or0[0]), .fs_xor1(h_arrdiv24_fs42_xor1), .fs_or0(h_arrdiv24_fs42_or0));
  fs fs_h_arrdiv24_fs43_out(.a(h_arrdiv24_mux2to118_and1[0]), .b(b[19]), .bin(h_arrdiv24_fs42_or0[0]), .fs_xor1(h_arrdiv24_fs43_xor1), .fs_or0(h_arrdiv24_fs43_or0));
  fs fs_h_arrdiv24_fs44_out(.a(h_arrdiv24_mux2to119_and1[0]), .b(b[20]), .bin(h_arrdiv24_fs43_or0[0]), .fs_xor1(h_arrdiv24_fs44_xor1), .fs_or0(h_arrdiv24_fs44_or0));
  fs fs_h_arrdiv24_fs45_out(.a(h_arrdiv24_mux2to120_and1[0]), .b(b[21]), .bin(h_arrdiv24_fs44_or0[0]), .fs_xor1(h_arrdiv24_fs45_xor1), .fs_or0(h_arrdiv24_fs45_or0));
  fs fs_h_arrdiv24_fs46_out(.a(h_arrdiv24_mux2to121_and1[0]), .b(b[22]), .bin(h_arrdiv24_fs45_or0[0]), .fs_xor1(h_arrdiv24_fs46_xor1), .fs_or0(h_arrdiv24_fs46_or0));
  fs fs_h_arrdiv24_fs47_out(.a(h_arrdiv24_mux2to122_and1[0]), .b(b[23]), .bin(h_arrdiv24_fs46_or0[0]), .fs_xor1(h_arrdiv24_fs47_xor1), .fs_or0(h_arrdiv24_fs47_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to123_out(.d0(h_arrdiv24_fs24_xor0[0]), .d1(a[22]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to123_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to124_out(.d0(h_arrdiv24_fs25_xor1[0]), .d1(h_arrdiv24_mux2to10_xor0[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to124_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to125_out(.d0(h_arrdiv24_fs26_xor1[0]), .d1(h_arrdiv24_mux2to11_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to125_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to126_out(.d0(h_arrdiv24_fs27_xor1[0]), .d1(h_arrdiv24_mux2to12_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to126_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to127_out(.d0(h_arrdiv24_fs28_xor1[0]), .d1(h_arrdiv24_mux2to13_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to127_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to128_out(.d0(h_arrdiv24_fs29_xor1[0]), .d1(h_arrdiv24_mux2to14_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to128_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to129_out(.d0(h_arrdiv24_fs30_xor1[0]), .d1(h_arrdiv24_mux2to15_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to129_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to130_out(.d0(h_arrdiv24_fs31_xor1[0]), .d1(h_arrdiv24_mux2to16_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to130_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to131_out(.d0(h_arrdiv24_fs32_xor1[0]), .d1(h_arrdiv24_mux2to17_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to131_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to132_out(.d0(h_arrdiv24_fs33_xor1[0]), .d1(h_arrdiv24_mux2to18_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to132_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to133_out(.d0(h_arrdiv24_fs34_xor1[0]), .d1(h_arrdiv24_mux2to19_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to133_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to134_out(.d0(h_arrdiv24_fs35_xor1[0]), .d1(h_arrdiv24_mux2to110_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to134_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to135_out(.d0(h_arrdiv24_fs36_xor1[0]), .d1(h_arrdiv24_mux2to111_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to135_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to136_out(.d0(h_arrdiv24_fs37_xor1[0]), .d1(h_arrdiv24_mux2to112_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to136_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to137_out(.d0(h_arrdiv24_fs38_xor1[0]), .d1(h_arrdiv24_mux2to113_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to137_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to138_out(.d0(h_arrdiv24_fs39_xor1[0]), .d1(h_arrdiv24_mux2to114_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to138_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to139_out(.d0(h_arrdiv24_fs40_xor1[0]), .d1(h_arrdiv24_mux2to115_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to139_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to140_out(.d0(h_arrdiv24_fs41_xor1[0]), .d1(h_arrdiv24_mux2to116_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to140_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to141_out(.d0(h_arrdiv24_fs42_xor1[0]), .d1(h_arrdiv24_mux2to117_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to141_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to142_out(.d0(h_arrdiv24_fs43_xor1[0]), .d1(h_arrdiv24_mux2to118_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to142_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to143_out(.d0(h_arrdiv24_fs44_xor1[0]), .d1(h_arrdiv24_mux2to119_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to143_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to144_out(.d0(h_arrdiv24_fs45_xor1[0]), .d1(h_arrdiv24_mux2to120_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to144_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to145_out(.d0(h_arrdiv24_fs46_xor1[0]), .d1(h_arrdiv24_mux2to121_and1[0]), .sel(h_arrdiv24_fs47_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to145_xor0));
  not_gate not_gate_h_arrdiv24_not1(.a(h_arrdiv24_fs47_or0[0]), .out(h_arrdiv24_not1));
  fs fs_h_arrdiv24_fs48_out(.a(a[21]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs48_xor0), .fs_or0(h_arrdiv24_fs48_and0));
  fs fs_h_arrdiv24_fs49_out(.a(h_arrdiv24_mux2to123_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs48_and0[0]), .fs_xor1(h_arrdiv24_fs49_xor1), .fs_or0(h_arrdiv24_fs49_or0));
  fs fs_h_arrdiv24_fs50_out(.a(h_arrdiv24_mux2to124_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs49_or0[0]), .fs_xor1(h_arrdiv24_fs50_xor1), .fs_or0(h_arrdiv24_fs50_or0));
  fs fs_h_arrdiv24_fs51_out(.a(h_arrdiv24_mux2to125_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs50_or0[0]), .fs_xor1(h_arrdiv24_fs51_xor1), .fs_or0(h_arrdiv24_fs51_or0));
  fs fs_h_arrdiv24_fs52_out(.a(h_arrdiv24_mux2to126_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs51_or0[0]), .fs_xor1(h_arrdiv24_fs52_xor1), .fs_or0(h_arrdiv24_fs52_or0));
  fs fs_h_arrdiv24_fs53_out(.a(h_arrdiv24_mux2to127_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs52_or0[0]), .fs_xor1(h_arrdiv24_fs53_xor1), .fs_or0(h_arrdiv24_fs53_or0));
  fs fs_h_arrdiv24_fs54_out(.a(h_arrdiv24_mux2to128_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs53_or0[0]), .fs_xor1(h_arrdiv24_fs54_xor1), .fs_or0(h_arrdiv24_fs54_or0));
  fs fs_h_arrdiv24_fs55_out(.a(h_arrdiv24_mux2to129_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs54_or0[0]), .fs_xor1(h_arrdiv24_fs55_xor1), .fs_or0(h_arrdiv24_fs55_or0));
  fs fs_h_arrdiv24_fs56_out(.a(h_arrdiv24_mux2to130_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs55_or0[0]), .fs_xor1(h_arrdiv24_fs56_xor1), .fs_or0(h_arrdiv24_fs56_or0));
  fs fs_h_arrdiv24_fs57_out(.a(h_arrdiv24_mux2to131_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs56_or0[0]), .fs_xor1(h_arrdiv24_fs57_xor1), .fs_or0(h_arrdiv24_fs57_or0));
  fs fs_h_arrdiv24_fs58_out(.a(h_arrdiv24_mux2to132_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs57_or0[0]), .fs_xor1(h_arrdiv24_fs58_xor1), .fs_or0(h_arrdiv24_fs58_or0));
  fs fs_h_arrdiv24_fs59_out(.a(h_arrdiv24_mux2to133_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs58_or0[0]), .fs_xor1(h_arrdiv24_fs59_xor1), .fs_or0(h_arrdiv24_fs59_or0));
  fs fs_h_arrdiv24_fs60_out(.a(h_arrdiv24_mux2to134_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs59_or0[0]), .fs_xor1(h_arrdiv24_fs60_xor1), .fs_or0(h_arrdiv24_fs60_or0));
  fs fs_h_arrdiv24_fs61_out(.a(h_arrdiv24_mux2to135_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs60_or0[0]), .fs_xor1(h_arrdiv24_fs61_xor1), .fs_or0(h_arrdiv24_fs61_or0));
  fs fs_h_arrdiv24_fs62_out(.a(h_arrdiv24_mux2to136_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs61_or0[0]), .fs_xor1(h_arrdiv24_fs62_xor1), .fs_or0(h_arrdiv24_fs62_or0));
  fs fs_h_arrdiv24_fs63_out(.a(h_arrdiv24_mux2to137_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs62_or0[0]), .fs_xor1(h_arrdiv24_fs63_xor1), .fs_or0(h_arrdiv24_fs63_or0));
  fs fs_h_arrdiv24_fs64_out(.a(h_arrdiv24_mux2to138_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs63_or0[0]), .fs_xor1(h_arrdiv24_fs64_xor1), .fs_or0(h_arrdiv24_fs64_or0));
  fs fs_h_arrdiv24_fs65_out(.a(h_arrdiv24_mux2to139_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs64_or0[0]), .fs_xor1(h_arrdiv24_fs65_xor1), .fs_or0(h_arrdiv24_fs65_or0));
  fs fs_h_arrdiv24_fs66_out(.a(h_arrdiv24_mux2to140_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs65_or0[0]), .fs_xor1(h_arrdiv24_fs66_xor1), .fs_or0(h_arrdiv24_fs66_or0));
  fs fs_h_arrdiv24_fs67_out(.a(h_arrdiv24_mux2to141_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs66_or0[0]), .fs_xor1(h_arrdiv24_fs67_xor1), .fs_or0(h_arrdiv24_fs67_or0));
  fs fs_h_arrdiv24_fs68_out(.a(h_arrdiv24_mux2to142_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs67_or0[0]), .fs_xor1(h_arrdiv24_fs68_xor1), .fs_or0(h_arrdiv24_fs68_or0));
  fs fs_h_arrdiv24_fs69_out(.a(h_arrdiv24_mux2to143_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs68_or0[0]), .fs_xor1(h_arrdiv24_fs69_xor1), .fs_or0(h_arrdiv24_fs69_or0));
  fs fs_h_arrdiv24_fs70_out(.a(h_arrdiv24_mux2to144_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs69_or0[0]), .fs_xor1(h_arrdiv24_fs70_xor1), .fs_or0(h_arrdiv24_fs70_or0));
  fs fs_h_arrdiv24_fs71_out(.a(h_arrdiv24_mux2to145_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs70_or0[0]), .fs_xor1(h_arrdiv24_fs71_xor1), .fs_or0(h_arrdiv24_fs71_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to146_out(.d0(h_arrdiv24_fs48_xor0[0]), .d1(a[21]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to146_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to147_out(.d0(h_arrdiv24_fs49_xor1[0]), .d1(h_arrdiv24_mux2to123_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to147_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to148_out(.d0(h_arrdiv24_fs50_xor1[0]), .d1(h_arrdiv24_mux2to124_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to148_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to149_out(.d0(h_arrdiv24_fs51_xor1[0]), .d1(h_arrdiv24_mux2to125_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to149_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to150_out(.d0(h_arrdiv24_fs52_xor1[0]), .d1(h_arrdiv24_mux2to126_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to150_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to151_out(.d0(h_arrdiv24_fs53_xor1[0]), .d1(h_arrdiv24_mux2to127_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to151_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to152_out(.d0(h_arrdiv24_fs54_xor1[0]), .d1(h_arrdiv24_mux2to128_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to152_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to153_out(.d0(h_arrdiv24_fs55_xor1[0]), .d1(h_arrdiv24_mux2to129_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to153_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to154_out(.d0(h_arrdiv24_fs56_xor1[0]), .d1(h_arrdiv24_mux2to130_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to154_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to155_out(.d0(h_arrdiv24_fs57_xor1[0]), .d1(h_arrdiv24_mux2to131_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to155_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to156_out(.d0(h_arrdiv24_fs58_xor1[0]), .d1(h_arrdiv24_mux2to132_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to156_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to157_out(.d0(h_arrdiv24_fs59_xor1[0]), .d1(h_arrdiv24_mux2to133_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to157_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to158_out(.d0(h_arrdiv24_fs60_xor1[0]), .d1(h_arrdiv24_mux2to134_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to158_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to159_out(.d0(h_arrdiv24_fs61_xor1[0]), .d1(h_arrdiv24_mux2to135_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to159_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to160_out(.d0(h_arrdiv24_fs62_xor1[0]), .d1(h_arrdiv24_mux2to136_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to160_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to161_out(.d0(h_arrdiv24_fs63_xor1[0]), .d1(h_arrdiv24_mux2to137_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to161_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to162_out(.d0(h_arrdiv24_fs64_xor1[0]), .d1(h_arrdiv24_mux2to138_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to162_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to163_out(.d0(h_arrdiv24_fs65_xor1[0]), .d1(h_arrdiv24_mux2to139_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to163_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to164_out(.d0(h_arrdiv24_fs66_xor1[0]), .d1(h_arrdiv24_mux2to140_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to164_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to165_out(.d0(h_arrdiv24_fs67_xor1[0]), .d1(h_arrdiv24_mux2to141_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to165_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to166_out(.d0(h_arrdiv24_fs68_xor1[0]), .d1(h_arrdiv24_mux2to142_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to166_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to167_out(.d0(h_arrdiv24_fs69_xor1[0]), .d1(h_arrdiv24_mux2to143_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to167_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to168_out(.d0(h_arrdiv24_fs70_xor1[0]), .d1(h_arrdiv24_mux2to144_xor0[0]), .sel(h_arrdiv24_fs71_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to168_xor0));
  not_gate not_gate_h_arrdiv24_not2(.a(h_arrdiv24_fs71_or0[0]), .out(h_arrdiv24_not2));
  fs fs_h_arrdiv24_fs72_out(.a(a[20]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs72_xor0), .fs_or0(h_arrdiv24_fs72_and0));
  fs fs_h_arrdiv24_fs73_out(.a(h_arrdiv24_mux2to146_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs72_and0[0]), .fs_xor1(h_arrdiv24_fs73_xor1), .fs_or0(h_arrdiv24_fs73_or0));
  fs fs_h_arrdiv24_fs74_out(.a(h_arrdiv24_mux2to147_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs73_or0[0]), .fs_xor1(h_arrdiv24_fs74_xor1), .fs_or0(h_arrdiv24_fs74_or0));
  fs fs_h_arrdiv24_fs75_out(.a(h_arrdiv24_mux2to148_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs74_or0[0]), .fs_xor1(h_arrdiv24_fs75_xor1), .fs_or0(h_arrdiv24_fs75_or0));
  fs fs_h_arrdiv24_fs76_out(.a(h_arrdiv24_mux2to149_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs75_or0[0]), .fs_xor1(h_arrdiv24_fs76_xor1), .fs_or0(h_arrdiv24_fs76_or0));
  fs fs_h_arrdiv24_fs77_out(.a(h_arrdiv24_mux2to150_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs76_or0[0]), .fs_xor1(h_arrdiv24_fs77_xor1), .fs_or0(h_arrdiv24_fs77_or0));
  fs fs_h_arrdiv24_fs78_out(.a(h_arrdiv24_mux2to151_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs77_or0[0]), .fs_xor1(h_arrdiv24_fs78_xor1), .fs_or0(h_arrdiv24_fs78_or0));
  fs fs_h_arrdiv24_fs79_out(.a(h_arrdiv24_mux2to152_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs78_or0[0]), .fs_xor1(h_arrdiv24_fs79_xor1), .fs_or0(h_arrdiv24_fs79_or0));
  fs fs_h_arrdiv24_fs80_out(.a(h_arrdiv24_mux2to153_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs79_or0[0]), .fs_xor1(h_arrdiv24_fs80_xor1), .fs_or0(h_arrdiv24_fs80_or0));
  fs fs_h_arrdiv24_fs81_out(.a(h_arrdiv24_mux2to154_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs80_or0[0]), .fs_xor1(h_arrdiv24_fs81_xor1), .fs_or0(h_arrdiv24_fs81_or0));
  fs fs_h_arrdiv24_fs82_out(.a(h_arrdiv24_mux2to155_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs81_or0[0]), .fs_xor1(h_arrdiv24_fs82_xor1), .fs_or0(h_arrdiv24_fs82_or0));
  fs fs_h_arrdiv24_fs83_out(.a(h_arrdiv24_mux2to156_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs82_or0[0]), .fs_xor1(h_arrdiv24_fs83_xor1), .fs_or0(h_arrdiv24_fs83_or0));
  fs fs_h_arrdiv24_fs84_out(.a(h_arrdiv24_mux2to157_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs83_or0[0]), .fs_xor1(h_arrdiv24_fs84_xor1), .fs_or0(h_arrdiv24_fs84_or0));
  fs fs_h_arrdiv24_fs85_out(.a(h_arrdiv24_mux2to158_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs84_or0[0]), .fs_xor1(h_arrdiv24_fs85_xor1), .fs_or0(h_arrdiv24_fs85_or0));
  fs fs_h_arrdiv24_fs86_out(.a(h_arrdiv24_mux2to159_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs85_or0[0]), .fs_xor1(h_arrdiv24_fs86_xor1), .fs_or0(h_arrdiv24_fs86_or0));
  fs fs_h_arrdiv24_fs87_out(.a(h_arrdiv24_mux2to160_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs86_or0[0]), .fs_xor1(h_arrdiv24_fs87_xor1), .fs_or0(h_arrdiv24_fs87_or0));
  fs fs_h_arrdiv24_fs88_out(.a(h_arrdiv24_mux2to161_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs87_or0[0]), .fs_xor1(h_arrdiv24_fs88_xor1), .fs_or0(h_arrdiv24_fs88_or0));
  fs fs_h_arrdiv24_fs89_out(.a(h_arrdiv24_mux2to162_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs88_or0[0]), .fs_xor1(h_arrdiv24_fs89_xor1), .fs_or0(h_arrdiv24_fs89_or0));
  fs fs_h_arrdiv24_fs90_out(.a(h_arrdiv24_mux2to163_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs89_or0[0]), .fs_xor1(h_arrdiv24_fs90_xor1), .fs_or0(h_arrdiv24_fs90_or0));
  fs fs_h_arrdiv24_fs91_out(.a(h_arrdiv24_mux2to164_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs90_or0[0]), .fs_xor1(h_arrdiv24_fs91_xor1), .fs_or0(h_arrdiv24_fs91_or0));
  fs fs_h_arrdiv24_fs92_out(.a(h_arrdiv24_mux2to165_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs91_or0[0]), .fs_xor1(h_arrdiv24_fs92_xor1), .fs_or0(h_arrdiv24_fs92_or0));
  fs fs_h_arrdiv24_fs93_out(.a(h_arrdiv24_mux2to166_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs92_or0[0]), .fs_xor1(h_arrdiv24_fs93_xor1), .fs_or0(h_arrdiv24_fs93_or0));
  fs fs_h_arrdiv24_fs94_out(.a(h_arrdiv24_mux2to167_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs93_or0[0]), .fs_xor1(h_arrdiv24_fs94_xor1), .fs_or0(h_arrdiv24_fs94_or0));
  fs fs_h_arrdiv24_fs95_out(.a(h_arrdiv24_mux2to168_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs94_or0[0]), .fs_xor1(h_arrdiv24_fs95_xor1), .fs_or0(h_arrdiv24_fs95_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to169_out(.d0(h_arrdiv24_fs72_xor0[0]), .d1(a[20]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to169_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to170_out(.d0(h_arrdiv24_fs73_xor1[0]), .d1(h_arrdiv24_mux2to146_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to170_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to171_out(.d0(h_arrdiv24_fs74_xor1[0]), .d1(h_arrdiv24_mux2to147_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to171_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to172_out(.d0(h_arrdiv24_fs75_xor1[0]), .d1(h_arrdiv24_mux2to148_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to172_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to173_out(.d0(h_arrdiv24_fs76_xor1[0]), .d1(h_arrdiv24_mux2to149_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to173_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to174_out(.d0(h_arrdiv24_fs77_xor1[0]), .d1(h_arrdiv24_mux2to150_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to174_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to175_out(.d0(h_arrdiv24_fs78_xor1[0]), .d1(h_arrdiv24_mux2to151_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to175_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to176_out(.d0(h_arrdiv24_fs79_xor1[0]), .d1(h_arrdiv24_mux2to152_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to176_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to177_out(.d0(h_arrdiv24_fs80_xor1[0]), .d1(h_arrdiv24_mux2to153_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to177_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to178_out(.d0(h_arrdiv24_fs81_xor1[0]), .d1(h_arrdiv24_mux2to154_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to178_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to179_out(.d0(h_arrdiv24_fs82_xor1[0]), .d1(h_arrdiv24_mux2to155_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to179_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to180_out(.d0(h_arrdiv24_fs83_xor1[0]), .d1(h_arrdiv24_mux2to156_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to180_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to181_out(.d0(h_arrdiv24_fs84_xor1[0]), .d1(h_arrdiv24_mux2to157_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to181_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to182_out(.d0(h_arrdiv24_fs85_xor1[0]), .d1(h_arrdiv24_mux2to158_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to182_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to183_out(.d0(h_arrdiv24_fs86_xor1[0]), .d1(h_arrdiv24_mux2to159_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to183_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to184_out(.d0(h_arrdiv24_fs87_xor1[0]), .d1(h_arrdiv24_mux2to160_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to184_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to185_out(.d0(h_arrdiv24_fs88_xor1[0]), .d1(h_arrdiv24_mux2to161_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to185_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to186_out(.d0(h_arrdiv24_fs89_xor1[0]), .d1(h_arrdiv24_mux2to162_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to186_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to187_out(.d0(h_arrdiv24_fs90_xor1[0]), .d1(h_arrdiv24_mux2to163_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to187_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to188_out(.d0(h_arrdiv24_fs91_xor1[0]), .d1(h_arrdiv24_mux2to164_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to188_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to189_out(.d0(h_arrdiv24_fs92_xor1[0]), .d1(h_arrdiv24_mux2to165_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to189_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to190_out(.d0(h_arrdiv24_fs93_xor1[0]), .d1(h_arrdiv24_mux2to166_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to190_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to191_out(.d0(h_arrdiv24_fs94_xor1[0]), .d1(h_arrdiv24_mux2to167_xor0[0]), .sel(h_arrdiv24_fs95_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to191_xor0));
  not_gate not_gate_h_arrdiv24_not3(.a(h_arrdiv24_fs95_or0[0]), .out(h_arrdiv24_not3));
  fs fs_h_arrdiv24_fs96_out(.a(a[19]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs96_xor0), .fs_or0(h_arrdiv24_fs96_and0));
  fs fs_h_arrdiv24_fs97_out(.a(h_arrdiv24_mux2to169_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs96_and0[0]), .fs_xor1(h_arrdiv24_fs97_xor1), .fs_or0(h_arrdiv24_fs97_or0));
  fs fs_h_arrdiv24_fs98_out(.a(h_arrdiv24_mux2to170_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs97_or0[0]), .fs_xor1(h_arrdiv24_fs98_xor1), .fs_or0(h_arrdiv24_fs98_or0));
  fs fs_h_arrdiv24_fs99_out(.a(h_arrdiv24_mux2to171_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs98_or0[0]), .fs_xor1(h_arrdiv24_fs99_xor1), .fs_or0(h_arrdiv24_fs99_or0));
  fs fs_h_arrdiv24_fs100_out(.a(h_arrdiv24_mux2to172_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs99_or0[0]), .fs_xor1(h_arrdiv24_fs100_xor1), .fs_or0(h_arrdiv24_fs100_or0));
  fs fs_h_arrdiv24_fs101_out(.a(h_arrdiv24_mux2to173_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs100_or0[0]), .fs_xor1(h_arrdiv24_fs101_xor1), .fs_or0(h_arrdiv24_fs101_or0));
  fs fs_h_arrdiv24_fs102_out(.a(h_arrdiv24_mux2to174_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs101_or0[0]), .fs_xor1(h_arrdiv24_fs102_xor1), .fs_or0(h_arrdiv24_fs102_or0));
  fs fs_h_arrdiv24_fs103_out(.a(h_arrdiv24_mux2to175_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs102_or0[0]), .fs_xor1(h_arrdiv24_fs103_xor1), .fs_or0(h_arrdiv24_fs103_or0));
  fs fs_h_arrdiv24_fs104_out(.a(h_arrdiv24_mux2to176_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs103_or0[0]), .fs_xor1(h_arrdiv24_fs104_xor1), .fs_or0(h_arrdiv24_fs104_or0));
  fs fs_h_arrdiv24_fs105_out(.a(h_arrdiv24_mux2to177_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs104_or0[0]), .fs_xor1(h_arrdiv24_fs105_xor1), .fs_or0(h_arrdiv24_fs105_or0));
  fs fs_h_arrdiv24_fs106_out(.a(h_arrdiv24_mux2to178_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs105_or0[0]), .fs_xor1(h_arrdiv24_fs106_xor1), .fs_or0(h_arrdiv24_fs106_or0));
  fs fs_h_arrdiv24_fs107_out(.a(h_arrdiv24_mux2to179_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs106_or0[0]), .fs_xor1(h_arrdiv24_fs107_xor1), .fs_or0(h_arrdiv24_fs107_or0));
  fs fs_h_arrdiv24_fs108_out(.a(h_arrdiv24_mux2to180_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs107_or0[0]), .fs_xor1(h_arrdiv24_fs108_xor1), .fs_or0(h_arrdiv24_fs108_or0));
  fs fs_h_arrdiv24_fs109_out(.a(h_arrdiv24_mux2to181_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs108_or0[0]), .fs_xor1(h_arrdiv24_fs109_xor1), .fs_or0(h_arrdiv24_fs109_or0));
  fs fs_h_arrdiv24_fs110_out(.a(h_arrdiv24_mux2to182_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs109_or0[0]), .fs_xor1(h_arrdiv24_fs110_xor1), .fs_or0(h_arrdiv24_fs110_or0));
  fs fs_h_arrdiv24_fs111_out(.a(h_arrdiv24_mux2to183_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs110_or0[0]), .fs_xor1(h_arrdiv24_fs111_xor1), .fs_or0(h_arrdiv24_fs111_or0));
  fs fs_h_arrdiv24_fs112_out(.a(h_arrdiv24_mux2to184_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs111_or0[0]), .fs_xor1(h_arrdiv24_fs112_xor1), .fs_or0(h_arrdiv24_fs112_or0));
  fs fs_h_arrdiv24_fs113_out(.a(h_arrdiv24_mux2to185_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs112_or0[0]), .fs_xor1(h_arrdiv24_fs113_xor1), .fs_or0(h_arrdiv24_fs113_or0));
  fs fs_h_arrdiv24_fs114_out(.a(h_arrdiv24_mux2to186_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs113_or0[0]), .fs_xor1(h_arrdiv24_fs114_xor1), .fs_or0(h_arrdiv24_fs114_or0));
  fs fs_h_arrdiv24_fs115_out(.a(h_arrdiv24_mux2to187_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs114_or0[0]), .fs_xor1(h_arrdiv24_fs115_xor1), .fs_or0(h_arrdiv24_fs115_or0));
  fs fs_h_arrdiv24_fs116_out(.a(h_arrdiv24_mux2to188_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs115_or0[0]), .fs_xor1(h_arrdiv24_fs116_xor1), .fs_or0(h_arrdiv24_fs116_or0));
  fs fs_h_arrdiv24_fs117_out(.a(h_arrdiv24_mux2to189_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs116_or0[0]), .fs_xor1(h_arrdiv24_fs117_xor1), .fs_or0(h_arrdiv24_fs117_or0));
  fs fs_h_arrdiv24_fs118_out(.a(h_arrdiv24_mux2to190_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs117_or0[0]), .fs_xor1(h_arrdiv24_fs118_xor1), .fs_or0(h_arrdiv24_fs118_or0));
  fs fs_h_arrdiv24_fs119_out(.a(h_arrdiv24_mux2to191_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs118_or0[0]), .fs_xor1(h_arrdiv24_fs119_xor1), .fs_or0(h_arrdiv24_fs119_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to192_out(.d0(h_arrdiv24_fs96_xor0[0]), .d1(a[19]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to192_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to193_out(.d0(h_arrdiv24_fs97_xor1[0]), .d1(h_arrdiv24_mux2to169_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to193_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to194_out(.d0(h_arrdiv24_fs98_xor1[0]), .d1(h_arrdiv24_mux2to170_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to194_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to195_out(.d0(h_arrdiv24_fs99_xor1[0]), .d1(h_arrdiv24_mux2to171_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to195_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to196_out(.d0(h_arrdiv24_fs100_xor1[0]), .d1(h_arrdiv24_mux2to172_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to196_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to197_out(.d0(h_arrdiv24_fs101_xor1[0]), .d1(h_arrdiv24_mux2to173_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to197_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to198_out(.d0(h_arrdiv24_fs102_xor1[0]), .d1(h_arrdiv24_mux2to174_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to198_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to199_out(.d0(h_arrdiv24_fs103_xor1[0]), .d1(h_arrdiv24_mux2to175_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to199_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1100_out(.d0(h_arrdiv24_fs104_xor1[0]), .d1(h_arrdiv24_mux2to176_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1100_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1101_out(.d0(h_arrdiv24_fs105_xor1[0]), .d1(h_arrdiv24_mux2to177_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1101_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1102_out(.d0(h_arrdiv24_fs106_xor1[0]), .d1(h_arrdiv24_mux2to178_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1102_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1103_out(.d0(h_arrdiv24_fs107_xor1[0]), .d1(h_arrdiv24_mux2to179_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1103_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1104_out(.d0(h_arrdiv24_fs108_xor1[0]), .d1(h_arrdiv24_mux2to180_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1104_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1105_out(.d0(h_arrdiv24_fs109_xor1[0]), .d1(h_arrdiv24_mux2to181_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1105_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1106_out(.d0(h_arrdiv24_fs110_xor1[0]), .d1(h_arrdiv24_mux2to182_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1106_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1107_out(.d0(h_arrdiv24_fs111_xor1[0]), .d1(h_arrdiv24_mux2to183_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1107_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1108_out(.d0(h_arrdiv24_fs112_xor1[0]), .d1(h_arrdiv24_mux2to184_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1108_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1109_out(.d0(h_arrdiv24_fs113_xor1[0]), .d1(h_arrdiv24_mux2to185_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1109_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1110_out(.d0(h_arrdiv24_fs114_xor1[0]), .d1(h_arrdiv24_mux2to186_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1110_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1111_out(.d0(h_arrdiv24_fs115_xor1[0]), .d1(h_arrdiv24_mux2to187_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1111_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1112_out(.d0(h_arrdiv24_fs116_xor1[0]), .d1(h_arrdiv24_mux2to188_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1112_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1113_out(.d0(h_arrdiv24_fs117_xor1[0]), .d1(h_arrdiv24_mux2to189_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1113_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1114_out(.d0(h_arrdiv24_fs118_xor1[0]), .d1(h_arrdiv24_mux2to190_xor0[0]), .sel(h_arrdiv24_fs119_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1114_xor0));
  not_gate not_gate_h_arrdiv24_not4(.a(h_arrdiv24_fs119_or0[0]), .out(h_arrdiv24_not4));
  fs fs_h_arrdiv24_fs120_out(.a(a[18]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs120_xor0), .fs_or0(h_arrdiv24_fs120_and0));
  fs fs_h_arrdiv24_fs121_out(.a(h_arrdiv24_mux2to192_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs120_and0[0]), .fs_xor1(h_arrdiv24_fs121_xor1), .fs_or0(h_arrdiv24_fs121_or0));
  fs fs_h_arrdiv24_fs122_out(.a(h_arrdiv24_mux2to193_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs121_or0[0]), .fs_xor1(h_arrdiv24_fs122_xor1), .fs_or0(h_arrdiv24_fs122_or0));
  fs fs_h_arrdiv24_fs123_out(.a(h_arrdiv24_mux2to194_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs122_or0[0]), .fs_xor1(h_arrdiv24_fs123_xor1), .fs_or0(h_arrdiv24_fs123_or0));
  fs fs_h_arrdiv24_fs124_out(.a(h_arrdiv24_mux2to195_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs123_or0[0]), .fs_xor1(h_arrdiv24_fs124_xor1), .fs_or0(h_arrdiv24_fs124_or0));
  fs fs_h_arrdiv24_fs125_out(.a(h_arrdiv24_mux2to196_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs124_or0[0]), .fs_xor1(h_arrdiv24_fs125_xor1), .fs_or0(h_arrdiv24_fs125_or0));
  fs fs_h_arrdiv24_fs126_out(.a(h_arrdiv24_mux2to197_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs125_or0[0]), .fs_xor1(h_arrdiv24_fs126_xor1), .fs_or0(h_arrdiv24_fs126_or0));
  fs fs_h_arrdiv24_fs127_out(.a(h_arrdiv24_mux2to198_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs126_or0[0]), .fs_xor1(h_arrdiv24_fs127_xor1), .fs_or0(h_arrdiv24_fs127_or0));
  fs fs_h_arrdiv24_fs128_out(.a(h_arrdiv24_mux2to199_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs127_or0[0]), .fs_xor1(h_arrdiv24_fs128_xor1), .fs_or0(h_arrdiv24_fs128_or0));
  fs fs_h_arrdiv24_fs129_out(.a(h_arrdiv24_mux2to1100_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs128_or0[0]), .fs_xor1(h_arrdiv24_fs129_xor1), .fs_or0(h_arrdiv24_fs129_or0));
  fs fs_h_arrdiv24_fs130_out(.a(h_arrdiv24_mux2to1101_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs129_or0[0]), .fs_xor1(h_arrdiv24_fs130_xor1), .fs_or0(h_arrdiv24_fs130_or0));
  fs fs_h_arrdiv24_fs131_out(.a(h_arrdiv24_mux2to1102_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs130_or0[0]), .fs_xor1(h_arrdiv24_fs131_xor1), .fs_or0(h_arrdiv24_fs131_or0));
  fs fs_h_arrdiv24_fs132_out(.a(h_arrdiv24_mux2to1103_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs131_or0[0]), .fs_xor1(h_arrdiv24_fs132_xor1), .fs_or0(h_arrdiv24_fs132_or0));
  fs fs_h_arrdiv24_fs133_out(.a(h_arrdiv24_mux2to1104_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs132_or0[0]), .fs_xor1(h_arrdiv24_fs133_xor1), .fs_or0(h_arrdiv24_fs133_or0));
  fs fs_h_arrdiv24_fs134_out(.a(h_arrdiv24_mux2to1105_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs133_or0[0]), .fs_xor1(h_arrdiv24_fs134_xor1), .fs_or0(h_arrdiv24_fs134_or0));
  fs fs_h_arrdiv24_fs135_out(.a(h_arrdiv24_mux2to1106_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs134_or0[0]), .fs_xor1(h_arrdiv24_fs135_xor1), .fs_or0(h_arrdiv24_fs135_or0));
  fs fs_h_arrdiv24_fs136_out(.a(h_arrdiv24_mux2to1107_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs135_or0[0]), .fs_xor1(h_arrdiv24_fs136_xor1), .fs_or0(h_arrdiv24_fs136_or0));
  fs fs_h_arrdiv24_fs137_out(.a(h_arrdiv24_mux2to1108_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs136_or0[0]), .fs_xor1(h_arrdiv24_fs137_xor1), .fs_or0(h_arrdiv24_fs137_or0));
  fs fs_h_arrdiv24_fs138_out(.a(h_arrdiv24_mux2to1109_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs137_or0[0]), .fs_xor1(h_arrdiv24_fs138_xor1), .fs_or0(h_arrdiv24_fs138_or0));
  fs fs_h_arrdiv24_fs139_out(.a(h_arrdiv24_mux2to1110_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs138_or0[0]), .fs_xor1(h_arrdiv24_fs139_xor1), .fs_or0(h_arrdiv24_fs139_or0));
  fs fs_h_arrdiv24_fs140_out(.a(h_arrdiv24_mux2to1111_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs139_or0[0]), .fs_xor1(h_arrdiv24_fs140_xor1), .fs_or0(h_arrdiv24_fs140_or0));
  fs fs_h_arrdiv24_fs141_out(.a(h_arrdiv24_mux2to1112_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs140_or0[0]), .fs_xor1(h_arrdiv24_fs141_xor1), .fs_or0(h_arrdiv24_fs141_or0));
  fs fs_h_arrdiv24_fs142_out(.a(h_arrdiv24_mux2to1113_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs141_or0[0]), .fs_xor1(h_arrdiv24_fs142_xor1), .fs_or0(h_arrdiv24_fs142_or0));
  fs fs_h_arrdiv24_fs143_out(.a(h_arrdiv24_mux2to1114_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs142_or0[0]), .fs_xor1(h_arrdiv24_fs143_xor1), .fs_or0(h_arrdiv24_fs143_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1115_out(.d0(h_arrdiv24_fs120_xor0[0]), .d1(a[18]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1115_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1116_out(.d0(h_arrdiv24_fs121_xor1[0]), .d1(h_arrdiv24_mux2to192_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1116_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1117_out(.d0(h_arrdiv24_fs122_xor1[0]), .d1(h_arrdiv24_mux2to193_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1117_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1118_out(.d0(h_arrdiv24_fs123_xor1[0]), .d1(h_arrdiv24_mux2to194_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1118_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1119_out(.d0(h_arrdiv24_fs124_xor1[0]), .d1(h_arrdiv24_mux2to195_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1119_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1120_out(.d0(h_arrdiv24_fs125_xor1[0]), .d1(h_arrdiv24_mux2to196_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1120_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1121_out(.d0(h_arrdiv24_fs126_xor1[0]), .d1(h_arrdiv24_mux2to197_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1121_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1122_out(.d0(h_arrdiv24_fs127_xor1[0]), .d1(h_arrdiv24_mux2to198_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1122_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1123_out(.d0(h_arrdiv24_fs128_xor1[0]), .d1(h_arrdiv24_mux2to199_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1123_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1124_out(.d0(h_arrdiv24_fs129_xor1[0]), .d1(h_arrdiv24_mux2to1100_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1124_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1125_out(.d0(h_arrdiv24_fs130_xor1[0]), .d1(h_arrdiv24_mux2to1101_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1125_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1126_out(.d0(h_arrdiv24_fs131_xor1[0]), .d1(h_arrdiv24_mux2to1102_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1126_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1127_out(.d0(h_arrdiv24_fs132_xor1[0]), .d1(h_arrdiv24_mux2to1103_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1127_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1128_out(.d0(h_arrdiv24_fs133_xor1[0]), .d1(h_arrdiv24_mux2to1104_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1128_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1129_out(.d0(h_arrdiv24_fs134_xor1[0]), .d1(h_arrdiv24_mux2to1105_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1129_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1130_out(.d0(h_arrdiv24_fs135_xor1[0]), .d1(h_arrdiv24_mux2to1106_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1130_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1131_out(.d0(h_arrdiv24_fs136_xor1[0]), .d1(h_arrdiv24_mux2to1107_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1131_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1132_out(.d0(h_arrdiv24_fs137_xor1[0]), .d1(h_arrdiv24_mux2to1108_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1132_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1133_out(.d0(h_arrdiv24_fs138_xor1[0]), .d1(h_arrdiv24_mux2to1109_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1133_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1134_out(.d0(h_arrdiv24_fs139_xor1[0]), .d1(h_arrdiv24_mux2to1110_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1134_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1135_out(.d0(h_arrdiv24_fs140_xor1[0]), .d1(h_arrdiv24_mux2to1111_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1135_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1136_out(.d0(h_arrdiv24_fs141_xor1[0]), .d1(h_arrdiv24_mux2to1112_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1136_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1137_out(.d0(h_arrdiv24_fs142_xor1[0]), .d1(h_arrdiv24_mux2to1113_xor0[0]), .sel(h_arrdiv24_fs143_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1137_xor0));
  not_gate not_gate_h_arrdiv24_not5(.a(h_arrdiv24_fs143_or0[0]), .out(h_arrdiv24_not5));
  fs fs_h_arrdiv24_fs144_out(.a(a[17]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs144_xor0), .fs_or0(h_arrdiv24_fs144_and0));
  fs fs_h_arrdiv24_fs145_out(.a(h_arrdiv24_mux2to1115_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs144_and0[0]), .fs_xor1(h_arrdiv24_fs145_xor1), .fs_or0(h_arrdiv24_fs145_or0));
  fs fs_h_arrdiv24_fs146_out(.a(h_arrdiv24_mux2to1116_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs145_or0[0]), .fs_xor1(h_arrdiv24_fs146_xor1), .fs_or0(h_arrdiv24_fs146_or0));
  fs fs_h_arrdiv24_fs147_out(.a(h_arrdiv24_mux2to1117_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs146_or0[0]), .fs_xor1(h_arrdiv24_fs147_xor1), .fs_or0(h_arrdiv24_fs147_or0));
  fs fs_h_arrdiv24_fs148_out(.a(h_arrdiv24_mux2to1118_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs147_or0[0]), .fs_xor1(h_arrdiv24_fs148_xor1), .fs_or0(h_arrdiv24_fs148_or0));
  fs fs_h_arrdiv24_fs149_out(.a(h_arrdiv24_mux2to1119_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs148_or0[0]), .fs_xor1(h_arrdiv24_fs149_xor1), .fs_or0(h_arrdiv24_fs149_or0));
  fs fs_h_arrdiv24_fs150_out(.a(h_arrdiv24_mux2to1120_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs149_or0[0]), .fs_xor1(h_arrdiv24_fs150_xor1), .fs_or0(h_arrdiv24_fs150_or0));
  fs fs_h_arrdiv24_fs151_out(.a(h_arrdiv24_mux2to1121_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs150_or0[0]), .fs_xor1(h_arrdiv24_fs151_xor1), .fs_or0(h_arrdiv24_fs151_or0));
  fs fs_h_arrdiv24_fs152_out(.a(h_arrdiv24_mux2to1122_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs151_or0[0]), .fs_xor1(h_arrdiv24_fs152_xor1), .fs_or0(h_arrdiv24_fs152_or0));
  fs fs_h_arrdiv24_fs153_out(.a(h_arrdiv24_mux2to1123_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs152_or0[0]), .fs_xor1(h_arrdiv24_fs153_xor1), .fs_or0(h_arrdiv24_fs153_or0));
  fs fs_h_arrdiv24_fs154_out(.a(h_arrdiv24_mux2to1124_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs153_or0[0]), .fs_xor1(h_arrdiv24_fs154_xor1), .fs_or0(h_arrdiv24_fs154_or0));
  fs fs_h_arrdiv24_fs155_out(.a(h_arrdiv24_mux2to1125_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs154_or0[0]), .fs_xor1(h_arrdiv24_fs155_xor1), .fs_or0(h_arrdiv24_fs155_or0));
  fs fs_h_arrdiv24_fs156_out(.a(h_arrdiv24_mux2to1126_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs155_or0[0]), .fs_xor1(h_arrdiv24_fs156_xor1), .fs_or0(h_arrdiv24_fs156_or0));
  fs fs_h_arrdiv24_fs157_out(.a(h_arrdiv24_mux2to1127_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs156_or0[0]), .fs_xor1(h_arrdiv24_fs157_xor1), .fs_or0(h_arrdiv24_fs157_or0));
  fs fs_h_arrdiv24_fs158_out(.a(h_arrdiv24_mux2to1128_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs157_or0[0]), .fs_xor1(h_arrdiv24_fs158_xor1), .fs_or0(h_arrdiv24_fs158_or0));
  fs fs_h_arrdiv24_fs159_out(.a(h_arrdiv24_mux2to1129_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs158_or0[0]), .fs_xor1(h_arrdiv24_fs159_xor1), .fs_or0(h_arrdiv24_fs159_or0));
  fs fs_h_arrdiv24_fs160_out(.a(h_arrdiv24_mux2to1130_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs159_or0[0]), .fs_xor1(h_arrdiv24_fs160_xor1), .fs_or0(h_arrdiv24_fs160_or0));
  fs fs_h_arrdiv24_fs161_out(.a(h_arrdiv24_mux2to1131_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs160_or0[0]), .fs_xor1(h_arrdiv24_fs161_xor1), .fs_or0(h_arrdiv24_fs161_or0));
  fs fs_h_arrdiv24_fs162_out(.a(h_arrdiv24_mux2to1132_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs161_or0[0]), .fs_xor1(h_arrdiv24_fs162_xor1), .fs_or0(h_arrdiv24_fs162_or0));
  fs fs_h_arrdiv24_fs163_out(.a(h_arrdiv24_mux2to1133_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs162_or0[0]), .fs_xor1(h_arrdiv24_fs163_xor1), .fs_or0(h_arrdiv24_fs163_or0));
  fs fs_h_arrdiv24_fs164_out(.a(h_arrdiv24_mux2to1134_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs163_or0[0]), .fs_xor1(h_arrdiv24_fs164_xor1), .fs_or0(h_arrdiv24_fs164_or0));
  fs fs_h_arrdiv24_fs165_out(.a(h_arrdiv24_mux2to1135_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs164_or0[0]), .fs_xor1(h_arrdiv24_fs165_xor1), .fs_or0(h_arrdiv24_fs165_or0));
  fs fs_h_arrdiv24_fs166_out(.a(h_arrdiv24_mux2to1136_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs165_or0[0]), .fs_xor1(h_arrdiv24_fs166_xor1), .fs_or0(h_arrdiv24_fs166_or0));
  fs fs_h_arrdiv24_fs167_out(.a(h_arrdiv24_mux2to1137_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs166_or0[0]), .fs_xor1(h_arrdiv24_fs167_xor1), .fs_or0(h_arrdiv24_fs167_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1138_out(.d0(h_arrdiv24_fs144_xor0[0]), .d1(a[17]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1138_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1139_out(.d0(h_arrdiv24_fs145_xor1[0]), .d1(h_arrdiv24_mux2to1115_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1139_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1140_out(.d0(h_arrdiv24_fs146_xor1[0]), .d1(h_arrdiv24_mux2to1116_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1140_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1141_out(.d0(h_arrdiv24_fs147_xor1[0]), .d1(h_arrdiv24_mux2to1117_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1141_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1142_out(.d0(h_arrdiv24_fs148_xor1[0]), .d1(h_arrdiv24_mux2to1118_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1142_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1143_out(.d0(h_arrdiv24_fs149_xor1[0]), .d1(h_arrdiv24_mux2to1119_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1143_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1144_out(.d0(h_arrdiv24_fs150_xor1[0]), .d1(h_arrdiv24_mux2to1120_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1144_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1145_out(.d0(h_arrdiv24_fs151_xor1[0]), .d1(h_arrdiv24_mux2to1121_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1145_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1146_out(.d0(h_arrdiv24_fs152_xor1[0]), .d1(h_arrdiv24_mux2to1122_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1146_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1147_out(.d0(h_arrdiv24_fs153_xor1[0]), .d1(h_arrdiv24_mux2to1123_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1147_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1148_out(.d0(h_arrdiv24_fs154_xor1[0]), .d1(h_arrdiv24_mux2to1124_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1148_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1149_out(.d0(h_arrdiv24_fs155_xor1[0]), .d1(h_arrdiv24_mux2to1125_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1149_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1150_out(.d0(h_arrdiv24_fs156_xor1[0]), .d1(h_arrdiv24_mux2to1126_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1150_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1151_out(.d0(h_arrdiv24_fs157_xor1[0]), .d1(h_arrdiv24_mux2to1127_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1151_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1152_out(.d0(h_arrdiv24_fs158_xor1[0]), .d1(h_arrdiv24_mux2to1128_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1152_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1153_out(.d0(h_arrdiv24_fs159_xor1[0]), .d1(h_arrdiv24_mux2to1129_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1153_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1154_out(.d0(h_arrdiv24_fs160_xor1[0]), .d1(h_arrdiv24_mux2to1130_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1154_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1155_out(.d0(h_arrdiv24_fs161_xor1[0]), .d1(h_arrdiv24_mux2to1131_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1155_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1156_out(.d0(h_arrdiv24_fs162_xor1[0]), .d1(h_arrdiv24_mux2to1132_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1156_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1157_out(.d0(h_arrdiv24_fs163_xor1[0]), .d1(h_arrdiv24_mux2to1133_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1157_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1158_out(.d0(h_arrdiv24_fs164_xor1[0]), .d1(h_arrdiv24_mux2to1134_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1158_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1159_out(.d0(h_arrdiv24_fs165_xor1[0]), .d1(h_arrdiv24_mux2to1135_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1159_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1160_out(.d0(h_arrdiv24_fs166_xor1[0]), .d1(h_arrdiv24_mux2to1136_xor0[0]), .sel(h_arrdiv24_fs167_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1160_xor0));
  not_gate not_gate_h_arrdiv24_not6(.a(h_arrdiv24_fs167_or0[0]), .out(h_arrdiv24_not6));
  fs fs_h_arrdiv24_fs168_out(.a(a[16]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs168_xor0), .fs_or0(h_arrdiv24_fs168_and0));
  fs fs_h_arrdiv24_fs169_out(.a(h_arrdiv24_mux2to1138_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs168_and0[0]), .fs_xor1(h_arrdiv24_fs169_xor1), .fs_or0(h_arrdiv24_fs169_or0));
  fs fs_h_arrdiv24_fs170_out(.a(h_arrdiv24_mux2to1139_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs169_or0[0]), .fs_xor1(h_arrdiv24_fs170_xor1), .fs_or0(h_arrdiv24_fs170_or0));
  fs fs_h_arrdiv24_fs171_out(.a(h_arrdiv24_mux2to1140_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs170_or0[0]), .fs_xor1(h_arrdiv24_fs171_xor1), .fs_or0(h_arrdiv24_fs171_or0));
  fs fs_h_arrdiv24_fs172_out(.a(h_arrdiv24_mux2to1141_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs171_or0[0]), .fs_xor1(h_arrdiv24_fs172_xor1), .fs_or0(h_arrdiv24_fs172_or0));
  fs fs_h_arrdiv24_fs173_out(.a(h_arrdiv24_mux2to1142_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs172_or0[0]), .fs_xor1(h_arrdiv24_fs173_xor1), .fs_or0(h_arrdiv24_fs173_or0));
  fs fs_h_arrdiv24_fs174_out(.a(h_arrdiv24_mux2to1143_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs173_or0[0]), .fs_xor1(h_arrdiv24_fs174_xor1), .fs_or0(h_arrdiv24_fs174_or0));
  fs fs_h_arrdiv24_fs175_out(.a(h_arrdiv24_mux2to1144_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs174_or0[0]), .fs_xor1(h_arrdiv24_fs175_xor1), .fs_or0(h_arrdiv24_fs175_or0));
  fs fs_h_arrdiv24_fs176_out(.a(h_arrdiv24_mux2to1145_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs175_or0[0]), .fs_xor1(h_arrdiv24_fs176_xor1), .fs_or0(h_arrdiv24_fs176_or0));
  fs fs_h_arrdiv24_fs177_out(.a(h_arrdiv24_mux2to1146_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs176_or0[0]), .fs_xor1(h_arrdiv24_fs177_xor1), .fs_or0(h_arrdiv24_fs177_or0));
  fs fs_h_arrdiv24_fs178_out(.a(h_arrdiv24_mux2to1147_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs177_or0[0]), .fs_xor1(h_arrdiv24_fs178_xor1), .fs_or0(h_arrdiv24_fs178_or0));
  fs fs_h_arrdiv24_fs179_out(.a(h_arrdiv24_mux2to1148_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs178_or0[0]), .fs_xor1(h_arrdiv24_fs179_xor1), .fs_or0(h_arrdiv24_fs179_or0));
  fs fs_h_arrdiv24_fs180_out(.a(h_arrdiv24_mux2to1149_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs179_or0[0]), .fs_xor1(h_arrdiv24_fs180_xor1), .fs_or0(h_arrdiv24_fs180_or0));
  fs fs_h_arrdiv24_fs181_out(.a(h_arrdiv24_mux2to1150_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs180_or0[0]), .fs_xor1(h_arrdiv24_fs181_xor1), .fs_or0(h_arrdiv24_fs181_or0));
  fs fs_h_arrdiv24_fs182_out(.a(h_arrdiv24_mux2to1151_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs181_or0[0]), .fs_xor1(h_arrdiv24_fs182_xor1), .fs_or0(h_arrdiv24_fs182_or0));
  fs fs_h_arrdiv24_fs183_out(.a(h_arrdiv24_mux2to1152_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs182_or0[0]), .fs_xor1(h_arrdiv24_fs183_xor1), .fs_or0(h_arrdiv24_fs183_or0));
  fs fs_h_arrdiv24_fs184_out(.a(h_arrdiv24_mux2to1153_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs183_or0[0]), .fs_xor1(h_arrdiv24_fs184_xor1), .fs_or0(h_arrdiv24_fs184_or0));
  fs fs_h_arrdiv24_fs185_out(.a(h_arrdiv24_mux2to1154_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs184_or0[0]), .fs_xor1(h_arrdiv24_fs185_xor1), .fs_or0(h_arrdiv24_fs185_or0));
  fs fs_h_arrdiv24_fs186_out(.a(h_arrdiv24_mux2to1155_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs185_or0[0]), .fs_xor1(h_arrdiv24_fs186_xor1), .fs_or0(h_arrdiv24_fs186_or0));
  fs fs_h_arrdiv24_fs187_out(.a(h_arrdiv24_mux2to1156_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs186_or0[0]), .fs_xor1(h_arrdiv24_fs187_xor1), .fs_or0(h_arrdiv24_fs187_or0));
  fs fs_h_arrdiv24_fs188_out(.a(h_arrdiv24_mux2to1157_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs187_or0[0]), .fs_xor1(h_arrdiv24_fs188_xor1), .fs_or0(h_arrdiv24_fs188_or0));
  fs fs_h_arrdiv24_fs189_out(.a(h_arrdiv24_mux2to1158_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs188_or0[0]), .fs_xor1(h_arrdiv24_fs189_xor1), .fs_or0(h_arrdiv24_fs189_or0));
  fs fs_h_arrdiv24_fs190_out(.a(h_arrdiv24_mux2to1159_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs189_or0[0]), .fs_xor1(h_arrdiv24_fs190_xor1), .fs_or0(h_arrdiv24_fs190_or0));
  fs fs_h_arrdiv24_fs191_out(.a(h_arrdiv24_mux2to1160_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs190_or0[0]), .fs_xor1(h_arrdiv24_fs191_xor1), .fs_or0(h_arrdiv24_fs191_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1161_out(.d0(h_arrdiv24_fs168_xor0[0]), .d1(a[16]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1161_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1162_out(.d0(h_arrdiv24_fs169_xor1[0]), .d1(h_arrdiv24_mux2to1138_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1162_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1163_out(.d0(h_arrdiv24_fs170_xor1[0]), .d1(h_arrdiv24_mux2to1139_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1163_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1164_out(.d0(h_arrdiv24_fs171_xor1[0]), .d1(h_arrdiv24_mux2to1140_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1164_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1165_out(.d0(h_arrdiv24_fs172_xor1[0]), .d1(h_arrdiv24_mux2to1141_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1165_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1166_out(.d0(h_arrdiv24_fs173_xor1[0]), .d1(h_arrdiv24_mux2to1142_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1166_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1167_out(.d0(h_arrdiv24_fs174_xor1[0]), .d1(h_arrdiv24_mux2to1143_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1167_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1168_out(.d0(h_arrdiv24_fs175_xor1[0]), .d1(h_arrdiv24_mux2to1144_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1168_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1169_out(.d0(h_arrdiv24_fs176_xor1[0]), .d1(h_arrdiv24_mux2to1145_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1169_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1170_out(.d0(h_arrdiv24_fs177_xor1[0]), .d1(h_arrdiv24_mux2to1146_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1170_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1171_out(.d0(h_arrdiv24_fs178_xor1[0]), .d1(h_arrdiv24_mux2to1147_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1171_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1172_out(.d0(h_arrdiv24_fs179_xor1[0]), .d1(h_arrdiv24_mux2to1148_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1172_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1173_out(.d0(h_arrdiv24_fs180_xor1[0]), .d1(h_arrdiv24_mux2to1149_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1173_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1174_out(.d0(h_arrdiv24_fs181_xor1[0]), .d1(h_arrdiv24_mux2to1150_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1174_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1175_out(.d0(h_arrdiv24_fs182_xor1[0]), .d1(h_arrdiv24_mux2to1151_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1175_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1176_out(.d0(h_arrdiv24_fs183_xor1[0]), .d1(h_arrdiv24_mux2to1152_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1176_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1177_out(.d0(h_arrdiv24_fs184_xor1[0]), .d1(h_arrdiv24_mux2to1153_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1177_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1178_out(.d0(h_arrdiv24_fs185_xor1[0]), .d1(h_arrdiv24_mux2to1154_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1178_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1179_out(.d0(h_arrdiv24_fs186_xor1[0]), .d1(h_arrdiv24_mux2to1155_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1179_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1180_out(.d0(h_arrdiv24_fs187_xor1[0]), .d1(h_arrdiv24_mux2to1156_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1180_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1181_out(.d0(h_arrdiv24_fs188_xor1[0]), .d1(h_arrdiv24_mux2to1157_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1181_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1182_out(.d0(h_arrdiv24_fs189_xor1[0]), .d1(h_arrdiv24_mux2to1158_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1182_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1183_out(.d0(h_arrdiv24_fs190_xor1[0]), .d1(h_arrdiv24_mux2to1159_xor0[0]), .sel(h_arrdiv24_fs191_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1183_xor0));
  not_gate not_gate_h_arrdiv24_not7(.a(h_arrdiv24_fs191_or0[0]), .out(h_arrdiv24_not7));
  fs fs_h_arrdiv24_fs192_out(.a(a[15]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs192_xor0), .fs_or0(h_arrdiv24_fs192_and0));
  fs fs_h_arrdiv24_fs193_out(.a(h_arrdiv24_mux2to1161_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs192_and0[0]), .fs_xor1(h_arrdiv24_fs193_xor1), .fs_or0(h_arrdiv24_fs193_or0));
  fs fs_h_arrdiv24_fs194_out(.a(h_arrdiv24_mux2to1162_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs193_or0[0]), .fs_xor1(h_arrdiv24_fs194_xor1), .fs_or0(h_arrdiv24_fs194_or0));
  fs fs_h_arrdiv24_fs195_out(.a(h_arrdiv24_mux2to1163_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs194_or0[0]), .fs_xor1(h_arrdiv24_fs195_xor1), .fs_or0(h_arrdiv24_fs195_or0));
  fs fs_h_arrdiv24_fs196_out(.a(h_arrdiv24_mux2to1164_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs195_or0[0]), .fs_xor1(h_arrdiv24_fs196_xor1), .fs_or0(h_arrdiv24_fs196_or0));
  fs fs_h_arrdiv24_fs197_out(.a(h_arrdiv24_mux2to1165_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs196_or0[0]), .fs_xor1(h_arrdiv24_fs197_xor1), .fs_or0(h_arrdiv24_fs197_or0));
  fs fs_h_arrdiv24_fs198_out(.a(h_arrdiv24_mux2to1166_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs197_or0[0]), .fs_xor1(h_arrdiv24_fs198_xor1), .fs_or0(h_arrdiv24_fs198_or0));
  fs fs_h_arrdiv24_fs199_out(.a(h_arrdiv24_mux2to1167_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs198_or0[0]), .fs_xor1(h_arrdiv24_fs199_xor1), .fs_or0(h_arrdiv24_fs199_or0));
  fs fs_h_arrdiv24_fs200_out(.a(h_arrdiv24_mux2to1168_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs199_or0[0]), .fs_xor1(h_arrdiv24_fs200_xor1), .fs_or0(h_arrdiv24_fs200_or0));
  fs fs_h_arrdiv24_fs201_out(.a(h_arrdiv24_mux2to1169_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs200_or0[0]), .fs_xor1(h_arrdiv24_fs201_xor1), .fs_or0(h_arrdiv24_fs201_or0));
  fs fs_h_arrdiv24_fs202_out(.a(h_arrdiv24_mux2to1170_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs201_or0[0]), .fs_xor1(h_arrdiv24_fs202_xor1), .fs_or0(h_arrdiv24_fs202_or0));
  fs fs_h_arrdiv24_fs203_out(.a(h_arrdiv24_mux2to1171_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs202_or0[0]), .fs_xor1(h_arrdiv24_fs203_xor1), .fs_or0(h_arrdiv24_fs203_or0));
  fs fs_h_arrdiv24_fs204_out(.a(h_arrdiv24_mux2to1172_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs203_or0[0]), .fs_xor1(h_arrdiv24_fs204_xor1), .fs_or0(h_arrdiv24_fs204_or0));
  fs fs_h_arrdiv24_fs205_out(.a(h_arrdiv24_mux2to1173_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs204_or0[0]), .fs_xor1(h_arrdiv24_fs205_xor1), .fs_or0(h_arrdiv24_fs205_or0));
  fs fs_h_arrdiv24_fs206_out(.a(h_arrdiv24_mux2to1174_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs205_or0[0]), .fs_xor1(h_arrdiv24_fs206_xor1), .fs_or0(h_arrdiv24_fs206_or0));
  fs fs_h_arrdiv24_fs207_out(.a(h_arrdiv24_mux2to1175_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs206_or0[0]), .fs_xor1(h_arrdiv24_fs207_xor1), .fs_or0(h_arrdiv24_fs207_or0));
  fs fs_h_arrdiv24_fs208_out(.a(h_arrdiv24_mux2to1176_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs207_or0[0]), .fs_xor1(h_arrdiv24_fs208_xor1), .fs_or0(h_arrdiv24_fs208_or0));
  fs fs_h_arrdiv24_fs209_out(.a(h_arrdiv24_mux2to1177_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs208_or0[0]), .fs_xor1(h_arrdiv24_fs209_xor1), .fs_or0(h_arrdiv24_fs209_or0));
  fs fs_h_arrdiv24_fs210_out(.a(h_arrdiv24_mux2to1178_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs209_or0[0]), .fs_xor1(h_arrdiv24_fs210_xor1), .fs_or0(h_arrdiv24_fs210_or0));
  fs fs_h_arrdiv24_fs211_out(.a(h_arrdiv24_mux2to1179_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs210_or0[0]), .fs_xor1(h_arrdiv24_fs211_xor1), .fs_or0(h_arrdiv24_fs211_or0));
  fs fs_h_arrdiv24_fs212_out(.a(h_arrdiv24_mux2to1180_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs211_or0[0]), .fs_xor1(h_arrdiv24_fs212_xor1), .fs_or0(h_arrdiv24_fs212_or0));
  fs fs_h_arrdiv24_fs213_out(.a(h_arrdiv24_mux2to1181_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs212_or0[0]), .fs_xor1(h_arrdiv24_fs213_xor1), .fs_or0(h_arrdiv24_fs213_or0));
  fs fs_h_arrdiv24_fs214_out(.a(h_arrdiv24_mux2to1182_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs213_or0[0]), .fs_xor1(h_arrdiv24_fs214_xor1), .fs_or0(h_arrdiv24_fs214_or0));
  fs fs_h_arrdiv24_fs215_out(.a(h_arrdiv24_mux2to1183_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs214_or0[0]), .fs_xor1(h_arrdiv24_fs215_xor1), .fs_or0(h_arrdiv24_fs215_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1184_out(.d0(h_arrdiv24_fs192_xor0[0]), .d1(a[15]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1184_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1185_out(.d0(h_arrdiv24_fs193_xor1[0]), .d1(h_arrdiv24_mux2to1161_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1185_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1186_out(.d0(h_arrdiv24_fs194_xor1[0]), .d1(h_arrdiv24_mux2to1162_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1186_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1187_out(.d0(h_arrdiv24_fs195_xor1[0]), .d1(h_arrdiv24_mux2to1163_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1187_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1188_out(.d0(h_arrdiv24_fs196_xor1[0]), .d1(h_arrdiv24_mux2to1164_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1188_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1189_out(.d0(h_arrdiv24_fs197_xor1[0]), .d1(h_arrdiv24_mux2to1165_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1189_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1190_out(.d0(h_arrdiv24_fs198_xor1[0]), .d1(h_arrdiv24_mux2to1166_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1190_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1191_out(.d0(h_arrdiv24_fs199_xor1[0]), .d1(h_arrdiv24_mux2to1167_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1191_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1192_out(.d0(h_arrdiv24_fs200_xor1[0]), .d1(h_arrdiv24_mux2to1168_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1192_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1193_out(.d0(h_arrdiv24_fs201_xor1[0]), .d1(h_arrdiv24_mux2to1169_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1193_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1194_out(.d0(h_arrdiv24_fs202_xor1[0]), .d1(h_arrdiv24_mux2to1170_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1194_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1195_out(.d0(h_arrdiv24_fs203_xor1[0]), .d1(h_arrdiv24_mux2to1171_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1195_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1196_out(.d0(h_arrdiv24_fs204_xor1[0]), .d1(h_arrdiv24_mux2to1172_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1196_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1197_out(.d0(h_arrdiv24_fs205_xor1[0]), .d1(h_arrdiv24_mux2to1173_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1197_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1198_out(.d0(h_arrdiv24_fs206_xor1[0]), .d1(h_arrdiv24_mux2to1174_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1198_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1199_out(.d0(h_arrdiv24_fs207_xor1[0]), .d1(h_arrdiv24_mux2to1175_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1199_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1200_out(.d0(h_arrdiv24_fs208_xor1[0]), .d1(h_arrdiv24_mux2to1176_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1200_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1201_out(.d0(h_arrdiv24_fs209_xor1[0]), .d1(h_arrdiv24_mux2to1177_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1201_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1202_out(.d0(h_arrdiv24_fs210_xor1[0]), .d1(h_arrdiv24_mux2to1178_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1202_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1203_out(.d0(h_arrdiv24_fs211_xor1[0]), .d1(h_arrdiv24_mux2to1179_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1203_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1204_out(.d0(h_arrdiv24_fs212_xor1[0]), .d1(h_arrdiv24_mux2to1180_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1204_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1205_out(.d0(h_arrdiv24_fs213_xor1[0]), .d1(h_arrdiv24_mux2to1181_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1205_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1206_out(.d0(h_arrdiv24_fs214_xor1[0]), .d1(h_arrdiv24_mux2to1182_xor0[0]), .sel(h_arrdiv24_fs215_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1206_xor0));
  not_gate not_gate_h_arrdiv24_not8(.a(h_arrdiv24_fs215_or0[0]), .out(h_arrdiv24_not8));
  fs fs_h_arrdiv24_fs216_out(.a(a[14]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs216_xor0), .fs_or0(h_arrdiv24_fs216_and0));
  fs fs_h_arrdiv24_fs217_out(.a(h_arrdiv24_mux2to1184_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs216_and0[0]), .fs_xor1(h_arrdiv24_fs217_xor1), .fs_or0(h_arrdiv24_fs217_or0));
  fs fs_h_arrdiv24_fs218_out(.a(h_arrdiv24_mux2to1185_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs217_or0[0]), .fs_xor1(h_arrdiv24_fs218_xor1), .fs_or0(h_arrdiv24_fs218_or0));
  fs fs_h_arrdiv24_fs219_out(.a(h_arrdiv24_mux2to1186_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs218_or0[0]), .fs_xor1(h_arrdiv24_fs219_xor1), .fs_or0(h_arrdiv24_fs219_or0));
  fs fs_h_arrdiv24_fs220_out(.a(h_arrdiv24_mux2to1187_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs219_or0[0]), .fs_xor1(h_arrdiv24_fs220_xor1), .fs_or0(h_arrdiv24_fs220_or0));
  fs fs_h_arrdiv24_fs221_out(.a(h_arrdiv24_mux2to1188_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs220_or0[0]), .fs_xor1(h_arrdiv24_fs221_xor1), .fs_or0(h_arrdiv24_fs221_or0));
  fs fs_h_arrdiv24_fs222_out(.a(h_arrdiv24_mux2to1189_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs221_or0[0]), .fs_xor1(h_arrdiv24_fs222_xor1), .fs_or0(h_arrdiv24_fs222_or0));
  fs fs_h_arrdiv24_fs223_out(.a(h_arrdiv24_mux2to1190_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs222_or0[0]), .fs_xor1(h_arrdiv24_fs223_xor1), .fs_or0(h_arrdiv24_fs223_or0));
  fs fs_h_arrdiv24_fs224_out(.a(h_arrdiv24_mux2to1191_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs223_or0[0]), .fs_xor1(h_arrdiv24_fs224_xor1), .fs_or0(h_arrdiv24_fs224_or0));
  fs fs_h_arrdiv24_fs225_out(.a(h_arrdiv24_mux2to1192_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs224_or0[0]), .fs_xor1(h_arrdiv24_fs225_xor1), .fs_or0(h_arrdiv24_fs225_or0));
  fs fs_h_arrdiv24_fs226_out(.a(h_arrdiv24_mux2to1193_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs225_or0[0]), .fs_xor1(h_arrdiv24_fs226_xor1), .fs_or0(h_arrdiv24_fs226_or0));
  fs fs_h_arrdiv24_fs227_out(.a(h_arrdiv24_mux2to1194_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs226_or0[0]), .fs_xor1(h_arrdiv24_fs227_xor1), .fs_or0(h_arrdiv24_fs227_or0));
  fs fs_h_arrdiv24_fs228_out(.a(h_arrdiv24_mux2to1195_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs227_or0[0]), .fs_xor1(h_arrdiv24_fs228_xor1), .fs_or0(h_arrdiv24_fs228_or0));
  fs fs_h_arrdiv24_fs229_out(.a(h_arrdiv24_mux2to1196_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs228_or0[0]), .fs_xor1(h_arrdiv24_fs229_xor1), .fs_or0(h_arrdiv24_fs229_or0));
  fs fs_h_arrdiv24_fs230_out(.a(h_arrdiv24_mux2to1197_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs229_or0[0]), .fs_xor1(h_arrdiv24_fs230_xor1), .fs_or0(h_arrdiv24_fs230_or0));
  fs fs_h_arrdiv24_fs231_out(.a(h_arrdiv24_mux2to1198_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs230_or0[0]), .fs_xor1(h_arrdiv24_fs231_xor1), .fs_or0(h_arrdiv24_fs231_or0));
  fs fs_h_arrdiv24_fs232_out(.a(h_arrdiv24_mux2to1199_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs231_or0[0]), .fs_xor1(h_arrdiv24_fs232_xor1), .fs_or0(h_arrdiv24_fs232_or0));
  fs fs_h_arrdiv24_fs233_out(.a(h_arrdiv24_mux2to1200_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs232_or0[0]), .fs_xor1(h_arrdiv24_fs233_xor1), .fs_or0(h_arrdiv24_fs233_or0));
  fs fs_h_arrdiv24_fs234_out(.a(h_arrdiv24_mux2to1201_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs233_or0[0]), .fs_xor1(h_arrdiv24_fs234_xor1), .fs_or0(h_arrdiv24_fs234_or0));
  fs fs_h_arrdiv24_fs235_out(.a(h_arrdiv24_mux2to1202_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs234_or0[0]), .fs_xor1(h_arrdiv24_fs235_xor1), .fs_or0(h_arrdiv24_fs235_or0));
  fs fs_h_arrdiv24_fs236_out(.a(h_arrdiv24_mux2to1203_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs235_or0[0]), .fs_xor1(h_arrdiv24_fs236_xor1), .fs_or0(h_arrdiv24_fs236_or0));
  fs fs_h_arrdiv24_fs237_out(.a(h_arrdiv24_mux2to1204_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs236_or0[0]), .fs_xor1(h_arrdiv24_fs237_xor1), .fs_or0(h_arrdiv24_fs237_or0));
  fs fs_h_arrdiv24_fs238_out(.a(h_arrdiv24_mux2to1205_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs237_or0[0]), .fs_xor1(h_arrdiv24_fs238_xor1), .fs_or0(h_arrdiv24_fs238_or0));
  fs fs_h_arrdiv24_fs239_out(.a(h_arrdiv24_mux2to1206_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs238_or0[0]), .fs_xor1(h_arrdiv24_fs239_xor1), .fs_or0(h_arrdiv24_fs239_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1207_out(.d0(h_arrdiv24_fs216_xor0[0]), .d1(a[14]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1207_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1208_out(.d0(h_arrdiv24_fs217_xor1[0]), .d1(h_arrdiv24_mux2to1184_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1208_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1209_out(.d0(h_arrdiv24_fs218_xor1[0]), .d1(h_arrdiv24_mux2to1185_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1209_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1210_out(.d0(h_arrdiv24_fs219_xor1[0]), .d1(h_arrdiv24_mux2to1186_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1210_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1211_out(.d0(h_arrdiv24_fs220_xor1[0]), .d1(h_arrdiv24_mux2to1187_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1211_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1212_out(.d0(h_arrdiv24_fs221_xor1[0]), .d1(h_arrdiv24_mux2to1188_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1212_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1213_out(.d0(h_arrdiv24_fs222_xor1[0]), .d1(h_arrdiv24_mux2to1189_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1213_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1214_out(.d0(h_arrdiv24_fs223_xor1[0]), .d1(h_arrdiv24_mux2to1190_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1214_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1215_out(.d0(h_arrdiv24_fs224_xor1[0]), .d1(h_arrdiv24_mux2to1191_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1215_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1216_out(.d0(h_arrdiv24_fs225_xor1[0]), .d1(h_arrdiv24_mux2to1192_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1216_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1217_out(.d0(h_arrdiv24_fs226_xor1[0]), .d1(h_arrdiv24_mux2to1193_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1217_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1218_out(.d0(h_arrdiv24_fs227_xor1[0]), .d1(h_arrdiv24_mux2to1194_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1218_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1219_out(.d0(h_arrdiv24_fs228_xor1[0]), .d1(h_arrdiv24_mux2to1195_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1219_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1220_out(.d0(h_arrdiv24_fs229_xor1[0]), .d1(h_arrdiv24_mux2to1196_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1220_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1221_out(.d0(h_arrdiv24_fs230_xor1[0]), .d1(h_arrdiv24_mux2to1197_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1221_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1222_out(.d0(h_arrdiv24_fs231_xor1[0]), .d1(h_arrdiv24_mux2to1198_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1222_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1223_out(.d0(h_arrdiv24_fs232_xor1[0]), .d1(h_arrdiv24_mux2to1199_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1223_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1224_out(.d0(h_arrdiv24_fs233_xor1[0]), .d1(h_arrdiv24_mux2to1200_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1224_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1225_out(.d0(h_arrdiv24_fs234_xor1[0]), .d1(h_arrdiv24_mux2to1201_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1225_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1226_out(.d0(h_arrdiv24_fs235_xor1[0]), .d1(h_arrdiv24_mux2to1202_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1226_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1227_out(.d0(h_arrdiv24_fs236_xor1[0]), .d1(h_arrdiv24_mux2to1203_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1227_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1228_out(.d0(h_arrdiv24_fs237_xor1[0]), .d1(h_arrdiv24_mux2to1204_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1228_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1229_out(.d0(h_arrdiv24_fs238_xor1[0]), .d1(h_arrdiv24_mux2to1205_xor0[0]), .sel(h_arrdiv24_fs239_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1229_xor0));
  not_gate not_gate_h_arrdiv24_not9(.a(h_arrdiv24_fs239_or0[0]), .out(h_arrdiv24_not9));
  fs fs_h_arrdiv24_fs240_out(.a(a[13]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs240_xor0), .fs_or0(h_arrdiv24_fs240_and0));
  fs fs_h_arrdiv24_fs241_out(.a(h_arrdiv24_mux2to1207_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs240_and0[0]), .fs_xor1(h_arrdiv24_fs241_xor1), .fs_or0(h_arrdiv24_fs241_or0));
  fs fs_h_arrdiv24_fs242_out(.a(h_arrdiv24_mux2to1208_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs241_or0[0]), .fs_xor1(h_arrdiv24_fs242_xor1), .fs_or0(h_arrdiv24_fs242_or0));
  fs fs_h_arrdiv24_fs243_out(.a(h_arrdiv24_mux2to1209_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs242_or0[0]), .fs_xor1(h_arrdiv24_fs243_xor1), .fs_or0(h_arrdiv24_fs243_or0));
  fs fs_h_arrdiv24_fs244_out(.a(h_arrdiv24_mux2to1210_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs243_or0[0]), .fs_xor1(h_arrdiv24_fs244_xor1), .fs_or0(h_arrdiv24_fs244_or0));
  fs fs_h_arrdiv24_fs245_out(.a(h_arrdiv24_mux2to1211_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs244_or0[0]), .fs_xor1(h_arrdiv24_fs245_xor1), .fs_or0(h_arrdiv24_fs245_or0));
  fs fs_h_arrdiv24_fs246_out(.a(h_arrdiv24_mux2to1212_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs245_or0[0]), .fs_xor1(h_arrdiv24_fs246_xor1), .fs_or0(h_arrdiv24_fs246_or0));
  fs fs_h_arrdiv24_fs247_out(.a(h_arrdiv24_mux2to1213_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs246_or0[0]), .fs_xor1(h_arrdiv24_fs247_xor1), .fs_or0(h_arrdiv24_fs247_or0));
  fs fs_h_arrdiv24_fs248_out(.a(h_arrdiv24_mux2to1214_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs247_or0[0]), .fs_xor1(h_arrdiv24_fs248_xor1), .fs_or0(h_arrdiv24_fs248_or0));
  fs fs_h_arrdiv24_fs249_out(.a(h_arrdiv24_mux2to1215_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs248_or0[0]), .fs_xor1(h_arrdiv24_fs249_xor1), .fs_or0(h_arrdiv24_fs249_or0));
  fs fs_h_arrdiv24_fs250_out(.a(h_arrdiv24_mux2to1216_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs249_or0[0]), .fs_xor1(h_arrdiv24_fs250_xor1), .fs_or0(h_arrdiv24_fs250_or0));
  fs fs_h_arrdiv24_fs251_out(.a(h_arrdiv24_mux2to1217_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs250_or0[0]), .fs_xor1(h_arrdiv24_fs251_xor1), .fs_or0(h_arrdiv24_fs251_or0));
  fs fs_h_arrdiv24_fs252_out(.a(h_arrdiv24_mux2to1218_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs251_or0[0]), .fs_xor1(h_arrdiv24_fs252_xor1), .fs_or0(h_arrdiv24_fs252_or0));
  fs fs_h_arrdiv24_fs253_out(.a(h_arrdiv24_mux2to1219_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs252_or0[0]), .fs_xor1(h_arrdiv24_fs253_xor1), .fs_or0(h_arrdiv24_fs253_or0));
  fs fs_h_arrdiv24_fs254_out(.a(h_arrdiv24_mux2to1220_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs253_or0[0]), .fs_xor1(h_arrdiv24_fs254_xor1), .fs_or0(h_arrdiv24_fs254_or0));
  fs fs_h_arrdiv24_fs255_out(.a(h_arrdiv24_mux2to1221_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs254_or0[0]), .fs_xor1(h_arrdiv24_fs255_xor1), .fs_or0(h_arrdiv24_fs255_or0));
  fs fs_h_arrdiv24_fs256_out(.a(h_arrdiv24_mux2to1222_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs255_or0[0]), .fs_xor1(h_arrdiv24_fs256_xor1), .fs_or0(h_arrdiv24_fs256_or0));
  fs fs_h_arrdiv24_fs257_out(.a(h_arrdiv24_mux2to1223_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs256_or0[0]), .fs_xor1(h_arrdiv24_fs257_xor1), .fs_or0(h_arrdiv24_fs257_or0));
  fs fs_h_arrdiv24_fs258_out(.a(h_arrdiv24_mux2to1224_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs257_or0[0]), .fs_xor1(h_arrdiv24_fs258_xor1), .fs_or0(h_arrdiv24_fs258_or0));
  fs fs_h_arrdiv24_fs259_out(.a(h_arrdiv24_mux2to1225_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs258_or0[0]), .fs_xor1(h_arrdiv24_fs259_xor1), .fs_or0(h_arrdiv24_fs259_or0));
  fs fs_h_arrdiv24_fs260_out(.a(h_arrdiv24_mux2to1226_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs259_or0[0]), .fs_xor1(h_arrdiv24_fs260_xor1), .fs_or0(h_arrdiv24_fs260_or0));
  fs fs_h_arrdiv24_fs261_out(.a(h_arrdiv24_mux2to1227_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs260_or0[0]), .fs_xor1(h_arrdiv24_fs261_xor1), .fs_or0(h_arrdiv24_fs261_or0));
  fs fs_h_arrdiv24_fs262_out(.a(h_arrdiv24_mux2to1228_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs261_or0[0]), .fs_xor1(h_arrdiv24_fs262_xor1), .fs_or0(h_arrdiv24_fs262_or0));
  fs fs_h_arrdiv24_fs263_out(.a(h_arrdiv24_mux2to1229_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs262_or0[0]), .fs_xor1(h_arrdiv24_fs263_xor1), .fs_or0(h_arrdiv24_fs263_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1230_out(.d0(h_arrdiv24_fs240_xor0[0]), .d1(a[13]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1230_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1231_out(.d0(h_arrdiv24_fs241_xor1[0]), .d1(h_arrdiv24_mux2to1207_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1231_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1232_out(.d0(h_arrdiv24_fs242_xor1[0]), .d1(h_arrdiv24_mux2to1208_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1232_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1233_out(.d0(h_arrdiv24_fs243_xor1[0]), .d1(h_arrdiv24_mux2to1209_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1233_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1234_out(.d0(h_arrdiv24_fs244_xor1[0]), .d1(h_arrdiv24_mux2to1210_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1234_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1235_out(.d0(h_arrdiv24_fs245_xor1[0]), .d1(h_arrdiv24_mux2to1211_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1235_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1236_out(.d0(h_arrdiv24_fs246_xor1[0]), .d1(h_arrdiv24_mux2to1212_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1236_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1237_out(.d0(h_arrdiv24_fs247_xor1[0]), .d1(h_arrdiv24_mux2to1213_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1237_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1238_out(.d0(h_arrdiv24_fs248_xor1[0]), .d1(h_arrdiv24_mux2to1214_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1238_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1239_out(.d0(h_arrdiv24_fs249_xor1[0]), .d1(h_arrdiv24_mux2to1215_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1239_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1240_out(.d0(h_arrdiv24_fs250_xor1[0]), .d1(h_arrdiv24_mux2to1216_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1240_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1241_out(.d0(h_arrdiv24_fs251_xor1[0]), .d1(h_arrdiv24_mux2to1217_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1241_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1242_out(.d0(h_arrdiv24_fs252_xor1[0]), .d1(h_arrdiv24_mux2to1218_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1242_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1243_out(.d0(h_arrdiv24_fs253_xor1[0]), .d1(h_arrdiv24_mux2to1219_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1243_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1244_out(.d0(h_arrdiv24_fs254_xor1[0]), .d1(h_arrdiv24_mux2to1220_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1244_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1245_out(.d0(h_arrdiv24_fs255_xor1[0]), .d1(h_arrdiv24_mux2to1221_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1245_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1246_out(.d0(h_arrdiv24_fs256_xor1[0]), .d1(h_arrdiv24_mux2to1222_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1246_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1247_out(.d0(h_arrdiv24_fs257_xor1[0]), .d1(h_arrdiv24_mux2to1223_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1247_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1248_out(.d0(h_arrdiv24_fs258_xor1[0]), .d1(h_arrdiv24_mux2to1224_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1248_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1249_out(.d0(h_arrdiv24_fs259_xor1[0]), .d1(h_arrdiv24_mux2to1225_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1249_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1250_out(.d0(h_arrdiv24_fs260_xor1[0]), .d1(h_arrdiv24_mux2to1226_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1250_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1251_out(.d0(h_arrdiv24_fs261_xor1[0]), .d1(h_arrdiv24_mux2to1227_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1251_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1252_out(.d0(h_arrdiv24_fs262_xor1[0]), .d1(h_arrdiv24_mux2to1228_xor0[0]), .sel(h_arrdiv24_fs263_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1252_xor0));
  not_gate not_gate_h_arrdiv24_not10(.a(h_arrdiv24_fs263_or0[0]), .out(h_arrdiv24_not10));
  fs fs_h_arrdiv24_fs264_out(.a(a[12]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs264_xor0), .fs_or0(h_arrdiv24_fs264_and0));
  fs fs_h_arrdiv24_fs265_out(.a(h_arrdiv24_mux2to1230_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs264_and0[0]), .fs_xor1(h_arrdiv24_fs265_xor1), .fs_or0(h_arrdiv24_fs265_or0));
  fs fs_h_arrdiv24_fs266_out(.a(h_arrdiv24_mux2to1231_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs265_or0[0]), .fs_xor1(h_arrdiv24_fs266_xor1), .fs_or0(h_arrdiv24_fs266_or0));
  fs fs_h_arrdiv24_fs267_out(.a(h_arrdiv24_mux2to1232_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs266_or0[0]), .fs_xor1(h_arrdiv24_fs267_xor1), .fs_or0(h_arrdiv24_fs267_or0));
  fs fs_h_arrdiv24_fs268_out(.a(h_arrdiv24_mux2to1233_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs267_or0[0]), .fs_xor1(h_arrdiv24_fs268_xor1), .fs_or0(h_arrdiv24_fs268_or0));
  fs fs_h_arrdiv24_fs269_out(.a(h_arrdiv24_mux2to1234_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs268_or0[0]), .fs_xor1(h_arrdiv24_fs269_xor1), .fs_or0(h_arrdiv24_fs269_or0));
  fs fs_h_arrdiv24_fs270_out(.a(h_arrdiv24_mux2to1235_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs269_or0[0]), .fs_xor1(h_arrdiv24_fs270_xor1), .fs_or0(h_arrdiv24_fs270_or0));
  fs fs_h_arrdiv24_fs271_out(.a(h_arrdiv24_mux2to1236_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs270_or0[0]), .fs_xor1(h_arrdiv24_fs271_xor1), .fs_or0(h_arrdiv24_fs271_or0));
  fs fs_h_arrdiv24_fs272_out(.a(h_arrdiv24_mux2to1237_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs271_or0[0]), .fs_xor1(h_arrdiv24_fs272_xor1), .fs_or0(h_arrdiv24_fs272_or0));
  fs fs_h_arrdiv24_fs273_out(.a(h_arrdiv24_mux2to1238_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs272_or0[0]), .fs_xor1(h_arrdiv24_fs273_xor1), .fs_or0(h_arrdiv24_fs273_or0));
  fs fs_h_arrdiv24_fs274_out(.a(h_arrdiv24_mux2to1239_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs273_or0[0]), .fs_xor1(h_arrdiv24_fs274_xor1), .fs_or0(h_arrdiv24_fs274_or0));
  fs fs_h_arrdiv24_fs275_out(.a(h_arrdiv24_mux2to1240_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs274_or0[0]), .fs_xor1(h_arrdiv24_fs275_xor1), .fs_or0(h_arrdiv24_fs275_or0));
  fs fs_h_arrdiv24_fs276_out(.a(h_arrdiv24_mux2to1241_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs275_or0[0]), .fs_xor1(h_arrdiv24_fs276_xor1), .fs_or0(h_arrdiv24_fs276_or0));
  fs fs_h_arrdiv24_fs277_out(.a(h_arrdiv24_mux2to1242_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs276_or0[0]), .fs_xor1(h_arrdiv24_fs277_xor1), .fs_or0(h_arrdiv24_fs277_or0));
  fs fs_h_arrdiv24_fs278_out(.a(h_arrdiv24_mux2to1243_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs277_or0[0]), .fs_xor1(h_arrdiv24_fs278_xor1), .fs_or0(h_arrdiv24_fs278_or0));
  fs fs_h_arrdiv24_fs279_out(.a(h_arrdiv24_mux2to1244_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs278_or0[0]), .fs_xor1(h_arrdiv24_fs279_xor1), .fs_or0(h_arrdiv24_fs279_or0));
  fs fs_h_arrdiv24_fs280_out(.a(h_arrdiv24_mux2to1245_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs279_or0[0]), .fs_xor1(h_arrdiv24_fs280_xor1), .fs_or0(h_arrdiv24_fs280_or0));
  fs fs_h_arrdiv24_fs281_out(.a(h_arrdiv24_mux2to1246_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs280_or0[0]), .fs_xor1(h_arrdiv24_fs281_xor1), .fs_or0(h_arrdiv24_fs281_or0));
  fs fs_h_arrdiv24_fs282_out(.a(h_arrdiv24_mux2to1247_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs281_or0[0]), .fs_xor1(h_arrdiv24_fs282_xor1), .fs_or0(h_arrdiv24_fs282_or0));
  fs fs_h_arrdiv24_fs283_out(.a(h_arrdiv24_mux2to1248_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs282_or0[0]), .fs_xor1(h_arrdiv24_fs283_xor1), .fs_or0(h_arrdiv24_fs283_or0));
  fs fs_h_arrdiv24_fs284_out(.a(h_arrdiv24_mux2to1249_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs283_or0[0]), .fs_xor1(h_arrdiv24_fs284_xor1), .fs_or0(h_arrdiv24_fs284_or0));
  fs fs_h_arrdiv24_fs285_out(.a(h_arrdiv24_mux2to1250_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs284_or0[0]), .fs_xor1(h_arrdiv24_fs285_xor1), .fs_or0(h_arrdiv24_fs285_or0));
  fs fs_h_arrdiv24_fs286_out(.a(h_arrdiv24_mux2to1251_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs285_or0[0]), .fs_xor1(h_arrdiv24_fs286_xor1), .fs_or0(h_arrdiv24_fs286_or0));
  fs fs_h_arrdiv24_fs287_out(.a(h_arrdiv24_mux2to1252_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs286_or0[0]), .fs_xor1(h_arrdiv24_fs287_xor1), .fs_or0(h_arrdiv24_fs287_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1253_out(.d0(h_arrdiv24_fs264_xor0[0]), .d1(a[12]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1253_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1254_out(.d0(h_arrdiv24_fs265_xor1[0]), .d1(h_arrdiv24_mux2to1230_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1254_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1255_out(.d0(h_arrdiv24_fs266_xor1[0]), .d1(h_arrdiv24_mux2to1231_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1255_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1256_out(.d0(h_arrdiv24_fs267_xor1[0]), .d1(h_arrdiv24_mux2to1232_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1256_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1257_out(.d0(h_arrdiv24_fs268_xor1[0]), .d1(h_arrdiv24_mux2to1233_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1257_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1258_out(.d0(h_arrdiv24_fs269_xor1[0]), .d1(h_arrdiv24_mux2to1234_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1258_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1259_out(.d0(h_arrdiv24_fs270_xor1[0]), .d1(h_arrdiv24_mux2to1235_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1259_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1260_out(.d0(h_arrdiv24_fs271_xor1[0]), .d1(h_arrdiv24_mux2to1236_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1260_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1261_out(.d0(h_arrdiv24_fs272_xor1[0]), .d1(h_arrdiv24_mux2to1237_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1261_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1262_out(.d0(h_arrdiv24_fs273_xor1[0]), .d1(h_arrdiv24_mux2to1238_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1262_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1263_out(.d0(h_arrdiv24_fs274_xor1[0]), .d1(h_arrdiv24_mux2to1239_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1263_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1264_out(.d0(h_arrdiv24_fs275_xor1[0]), .d1(h_arrdiv24_mux2to1240_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1264_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1265_out(.d0(h_arrdiv24_fs276_xor1[0]), .d1(h_arrdiv24_mux2to1241_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1265_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1266_out(.d0(h_arrdiv24_fs277_xor1[0]), .d1(h_arrdiv24_mux2to1242_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1266_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1267_out(.d0(h_arrdiv24_fs278_xor1[0]), .d1(h_arrdiv24_mux2to1243_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1267_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1268_out(.d0(h_arrdiv24_fs279_xor1[0]), .d1(h_arrdiv24_mux2to1244_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1268_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1269_out(.d0(h_arrdiv24_fs280_xor1[0]), .d1(h_arrdiv24_mux2to1245_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1269_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1270_out(.d0(h_arrdiv24_fs281_xor1[0]), .d1(h_arrdiv24_mux2to1246_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1270_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1271_out(.d0(h_arrdiv24_fs282_xor1[0]), .d1(h_arrdiv24_mux2to1247_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1271_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1272_out(.d0(h_arrdiv24_fs283_xor1[0]), .d1(h_arrdiv24_mux2to1248_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1272_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1273_out(.d0(h_arrdiv24_fs284_xor1[0]), .d1(h_arrdiv24_mux2to1249_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1273_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1274_out(.d0(h_arrdiv24_fs285_xor1[0]), .d1(h_arrdiv24_mux2to1250_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1274_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1275_out(.d0(h_arrdiv24_fs286_xor1[0]), .d1(h_arrdiv24_mux2to1251_xor0[0]), .sel(h_arrdiv24_fs287_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1275_xor0));
  not_gate not_gate_h_arrdiv24_not11(.a(h_arrdiv24_fs287_or0[0]), .out(h_arrdiv24_not11));
  fs fs_h_arrdiv24_fs288_out(.a(a[11]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs288_xor0), .fs_or0(h_arrdiv24_fs288_and0));
  fs fs_h_arrdiv24_fs289_out(.a(h_arrdiv24_mux2to1253_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs288_and0[0]), .fs_xor1(h_arrdiv24_fs289_xor1), .fs_or0(h_arrdiv24_fs289_or0));
  fs fs_h_arrdiv24_fs290_out(.a(h_arrdiv24_mux2to1254_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs289_or0[0]), .fs_xor1(h_arrdiv24_fs290_xor1), .fs_or0(h_arrdiv24_fs290_or0));
  fs fs_h_arrdiv24_fs291_out(.a(h_arrdiv24_mux2to1255_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs290_or0[0]), .fs_xor1(h_arrdiv24_fs291_xor1), .fs_or0(h_arrdiv24_fs291_or0));
  fs fs_h_arrdiv24_fs292_out(.a(h_arrdiv24_mux2to1256_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs291_or0[0]), .fs_xor1(h_arrdiv24_fs292_xor1), .fs_or0(h_arrdiv24_fs292_or0));
  fs fs_h_arrdiv24_fs293_out(.a(h_arrdiv24_mux2to1257_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs292_or0[0]), .fs_xor1(h_arrdiv24_fs293_xor1), .fs_or0(h_arrdiv24_fs293_or0));
  fs fs_h_arrdiv24_fs294_out(.a(h_arrdiv24_mux2to1258_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs293_or0[0]), .fs_xor1(h_arrdiv24_fs294_xor1), .fs_or0(h_arrdiv24_fs294_or0));
  fs fs_h_arrdiv24_fs295_out(.a(h_arrdiv24_mux2to1259_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs294_or0[0]), .fs_xor1(h_arrdiv24_fs295_xor1), .fs_or0(h_arrdiv24_fs295_or0));
  fs fs_h_arrdiv24_fs296_out(.a(h_arrdiv24_mux2to1260_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs295_or0[0]), .fs_xor1(h_arrdiv24_fs296_xor1), .fs_or0(h_arrdiv24_fs296_or0));
  fs fs_h_arrdiv24_fs297_out(.a(h_arrdiv24_mux2to1261_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs296_or0[0]), .fs_xor1(h_arrdiv24_fs297_xor1), .fs_or0(h_arrdiv24_fs297_or0));
  fs fs_h_arrdiv24_fs298_out(.a(h_arrdiv24_mux2to1262_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs297_or0[0]), .fs_xor1(h_arrdiv24_fs298_xor1), .fs_or0(h_arrdiv24_fs298_or0));
  fs fs_h_arrdiv24_fs299_out(.a(h_arrdiv24_mux2to1263_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs298_or0[0]), .fs_xor1(h_arrdiv24_fs299_xor1), .fs_or0(h_arrdiv24_fs299_or0));
  fs fs_h_arrdiv24_fs300_out(.a(h_arrdiv24_mux2to1264_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs299_or0[0]), .fs_xor1(h_arrdiv24_fs300_xor1), .fs_or0(h_arrdiv24_fs300_or0));
  fs fs_h_arrdiv24_fs301_out(.a(h_arrdiv24_mux2to1265_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs300_or0[0]), .fs_xor1(h_arrdiv24_fs301_xor1), .fs_or0(h_arrdiv24_fs301_or0));
  fs fs_h_arrdiv24_fs302_out(.a(h_arrdiv24_mux2to1266_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs301_or0[0]), .fs_xor1(h_arrdiv24_fs302_xor1), .fs_or0(h_arrdiv24_fs302_or0));
  fs fs_h_arrdiv24_fs303_out(.a(h_arrdiv24_mux2to1267_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs302_or0[0]), .fs_xor1(h_arrdiv24_fs303_xor1), .fs_or0(h_arrdiv24_fs303_or0));
  fs fs_h_arrdiv24_fs304_out(.a(h_arrdiv24_mux2to1268_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs303_or0[0]), .fs_xor1(h_arrdiv24_fs304_xor1), .fs_or0(h_arrdiv24_fs304_or0));
  fs fs_h_arrdiv24_fs305_out(.a(h_arrdiv24_mux2to1269_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs304_or0[0]), .fs_xor1(h_arrdiv24_fs305_xor1), .fs_or0(h_arrdiv24_fs305_or0));
  fs fs_h_arrdiv24_fs306_out(.a(h_arrdiv24_mux2to1270_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs305_or0[0]), .fs_xor1(h_arrdiv24_fs306_xor1), .fs_or0(h_arrdiv24_fs306_or0));
  fs fs_h_arrdiv24_fs307_out(.a(h_arrdiv24_mux2to1271_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs306_or0[0]), .fs_xor1(h_arrdiv24_fs307_xor1), .fs_or0(h_arrdiv24_fs307_or0));
  fs fs_h_arrdiv24_fs308_out(.a(h_arrdiv24_mux2to1272_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs307_or0[0]), .fs_xor1(h_arrdiv24_fs308_xor1), .fs_or0(h_arrdiv24_fs308_or0));
  fs fs_h_arrdiv24_fs309_out(.a(h_arrdiv24_mux2to1273_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs308_or0[0]), .fs_xor1(h_arrdiv24_fs309_xor1), .fs_or0(h_arrdiv24_fs309_or0));
  fs fs_h_arrdiv24_fs310_out(.a(h_arrdiv24_mux2to1274_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs309_or0[0]), .fs_xor1(h_arrdiv24_fs310_xor1), .fs_or0(h_arrdiv24_fs310_or0));
  fs fs_h_arrdiv24_fs311_out(.a(h_arrdiv24_mux2to1275_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs310_or0[0]), .fs_xor1(h_arrdiv24_fs311_xor1), .fs_or0(h_arrdiv24_fs311_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1276_out(.d0(h_arrdiv24_fs288_xor0[0]), .d1(a[11]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1276_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1277_out(.d0(h_arrdiv24_fs289_xor1[0]), .d1(h_arrdiv24_mux2to1253_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1277_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1278_out(.d0(h_arrdiv24_fs290_xor1[0]), .d1(h_arrdiv24_mux2to1254_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1278_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1279_out(.d0(h_arrdiv24_fs291_xor1[0]), .d1(h_arrdiv24_mux2to1255_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1279_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1280_out(.d0(h_arrdiv24_fs292_xor1[0]), .d1(h_arrdiv24_mux2to1256_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1280_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1281_out(.d0(h_arrdiv24_fs293_xor1[0]), .d1(h_arrdiv24_mux2to1257_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1281_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1282_out(.d0(h_arrdiv24_fs294_xor1[0]), .d1(h_arrdiv24_mux2to1258_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1282_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1283_out(.d0(h_arrdiv24_fs295_xor1[0]), .d1(h_arrdiv24_mux2to1259_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1283_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1284_out(.d0(h_arrdiv24_fs296_xor1[0]), .d1(h_arrdiv24_mux2to1260_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1284_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1285_out(.d0(h_arrdiv24_fs297_xor1[0]), .d1(h_arrdiv24_mux2to1261_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1285_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1286_out(.d0(h_arrdiv24_fs298_xor1[0]), .d1(h_arrdiv24_mux2to1262_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1286_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1287_out(.d0(h_arrdiv24_fs299_xor1[0]), .d1(h_arrdiv24_mux2to1263_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1287_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1288_out(.d0(h_arrdiv24_fs300_xor1[0]), .d1(h_arrdiv24_mux2to1264_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1288_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1289_out(.d0(h_arrdiv24_fs301_xor1[0]), .d1(h_arrdiv24_mux2to1265_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1289_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1290_out(.d0(h_arrdiv24_fs302_xor1[0]), .d1(h_arrdiv24_mux2to1266_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1290_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1291_out(.d0(h_arrdiv24_fs303_xor1[0]), .d1(h_arrdiv24_mux2to1267_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1291_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1292_out(.d0(h_arrdiv24_fs304_xor1[0]), .d1(h_arrdiv24_mux2to1268_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1292_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1293_out(.d0(h_arrdiv24_fs305_xor1[0]), .d1(h_arrdiv24_mux2to1269_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1293_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1294_out(.d0(h_arrdiv24_fs306_xor1[0]), .d1(h_arrdiv24_mux2to1270_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1294_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1295_out(.d0(h_arrdiv24_fs307_xor1[0]), .d1(h_arrdiv24_mux2to1271_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1295_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1296_out(.d0(h_arrdiv24_fs308_xor1[0]), .d1(h_arrdiv24_mux2to1272_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1296_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1297_out(.d0(h_arrdiv24_fs309_xor1[0]), .d1(h_arrdiv24_mux2to1273_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1297_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1298_out(.d0(h_arrdiv24_fs310_xor1[0]), .d1(h_arrdiv24_mux2to1274_xor0[0]), .sel(h_arrdiv24_fs311_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1298_xor0));
  not_gate not_gate_h_arrdiv24_not12(.a(h_arrdiv24_fs311_or0[0]), .out(h_arrdiv24_not12));
  fs fs_h_arrdiv24_fs312_out(.a(a[10]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs312_xor0), .fs_or0(h_arrdiv24_fs312_and0));
  fs fs_h_arrdiv24_fs313_out(.a(h_arrdiv24_mux2to1276_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs312_and0[0]), .fs_xor1(h_arrdiv24_fs313_xor1), .fs_or0(h_arrdiv24_fs313_or0));
  fs fs_h_arrdiv24_fs314_out(.a(h_arrdiv24_mux2to1277_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs313_or0[0]), .fs_xor1(h_arrdiv24_fs314_xor1), .fs_or0(h_arrdiv24_fs314_or0));
  fs fs_h_arrdiv24_fs315_out(.a(h_arrdiv24_mux2to1278_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs314_or0[0]), .fs_xor1(h_arrdiv24_fs315_xor1), .fs_or0(h_arrdiv24_fs315_or0));
  fs fs_h_arrdiv24_fs316_out(.a(h_arrdiv24_mux2to1279_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs315_or0[0]), .fs_xor1(h_arrdiv24_fs316_xor1), .fs_or0(h_arrdiv24_fs316_or0));
  fs fs_h_arrdiv24_fs317_out(.a(h_arrdiv24_mux2to1280_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs316_or0[0]), .fs_xor1(h_arrdiv24_fs317_xor1), .fs_or0(h_arrdiv24_fs317_or0));
  fs fs_h_arrdiv24_fs318_out(.a(h_arrdiv24_mux2to1281_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs317_or0[0]), .fs_xor1(h_arrdiv24_fs318_xor1), .fs_or0(h_arrdiv24_fs318_or0));
  fs fs_h_arrdiv24_fs319_out(.a(h_arrdiv24_mux2to1282_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs318_or0[0]), .fs_xor1(h_arrdiv24_fs319_xor1), .fs_or0(h_arrdiv24_fs319_or0));
  fs fs_h_arrdiv24_fs320_out(.a(h_arrdiv24_mux2to1283_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs319_or0[0]), .fs_xor1(h_arrdiv24_fs320_xor1), .fs_or0(h_arrdiv24_fs320_or0));
  fs fs_h_arrdiv24_fs321_out(.a(h_arrdiv24_mux2to1284_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs320_or0[0]), .fs_xor1(h_arrdiv24_fs321_xor1), .fs_or0(h_arrdiv24_fs321_or0));
  fs fs_h_arrdiv24_fs322_out(.a(h_arrdiv24_mux2to1285_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs321_or0[0]), .fs_xor1(h_arrdiv24_fs322_xor1), .fs_or0(h_arrdiv24_fs322_or0));
  fs fs_h_arrdiv24_fs323_out(.a(h_arrdiv24_mux2to1286_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs322_or0[0]), .fs_xor1(h_arrdiv24_fs323_xor1), .fs_or0(h_arrdiv24_fs323_or0));
  fs fs_h_arrdiv24_fs324_out(.a(h_arrdiv24_mux2to1287_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs323_or0[0]), .fs_xor1(h_arrdiv24_fs324_xor1), .fs_or0(h_arrdiv24_fs324_or0));
  fs fs_h_arrdiv24_fs325_out(.a(h_arrdiv24_mux2to1288_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs324_or0[0]), .fs_xor1(h_arrdiv24_fs325_xor1), .fs_or0(h_arrdiv24_fs325_or0));
  fs fs_h_arrdiv24_fs326_out(.a(h_arrdiv24_mux2to1289_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs325_or0[0]), .fs_xor1(h_arrdiv24_fs326_xor1), .fs_or0(h_arrdiv24_fs326_or0));
  fs fs_h_arrdiv24_fs327_out(.a(h_arrdiv24_mux2to1290_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs326_or0[0]), .fs_xor1(h_arrdiv24_fs327_xor1), .fs_or0(h_arrdiv24_fs327_or0));
  fs fs_h_arrdiv24_fs328_out(.a(h_arrdiv24_mux2to1291_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs327_or0[0]), .fs_xor1(h_arrdiv24_fs328_xor1), .fs_or0(h_arrdiv24_fs328_or0));
  fs fs_h_arrdiv24_fs329_out(.a(h_arrdiv24_mux2to1292_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs328_or0[0]), .fs_xor1(h_arrdiv24_fs329_xor1), .fs_or0(h_arrdiv24_fs329_or0));
  fs fs_h_arrdiv24_fs330_out(.a(h_arrdiv24_mux2to1293_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs329_or0[0]), .fs_xor1(h_arrdiv24_fs330_xor1), .fs_or0(h_arrdiv24_fs330_or0));
  fs fs_h_arrdiv24_fs331_out(.a(h_arrdiv24_mux2to1294_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs330_or0[0]), .fs_xor1(h_arrdiv24_fs331_xor1), .fs_or0(h_arrdiv24_fs331_or0));
  fs fs_h_arrdiv24_fs332_out(.a(h_arrdiv24_mux2to1295_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs331_or0[0]), .fs_xor1(h_arrdiv24_fs332_xor1), .fs_or0(h_arrdiv24_fs332_or0));
  fs fs_h_arrdiv24_fs333_out(.a(h_arrdiv24_mux2to1296_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs332_or0[0]), .fs_xor1(h_arrdiv24_fs333_xor1), .fs_or0(h_arrdiv24_fs333_or0));
  fs fs_h_arrdiv24_fs334_out(.a(h_arrdiv24_mux2to1297_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs333_or0[0]), .fs_xor1(h_arrdiv24_fs334_xor1), .fs_or0(h_arrdiv24_fs334_or0));
  fs fs_h_arrdiv24_fs335_out(.a(h_arrdiv24_mux2to1298_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs334_or0[0]), .fs_xor1(h_arrdiv24_fs335_xor1), .fs_or0(h_arrdiv24_fs335_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1299_out(.d0(h_arrdiv24_fs312_xor0[0]), .d1(a[10]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1299_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1300_out(.d0(h_arrdiv24_fs313_xor1[0]), .d1(h_arrdiv24_mux2to1276_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1300_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1301_out(.d0(h_arrdiv24_fs314_xor1[0]), .d1(h_arrdiv24_mux2to1277_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1301_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1302_out(.d0(h_arrdiv24_fs315_xor1[0]), .d1(h_arrdiv24_mux2to1278_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1302_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1303_out(.d0(h_arrdiv24_fs316_xor1[0]), .d1(h_arrdiv24_mux2to1279_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1303_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1304_out(.d0(h_arrdiv24_fs317_xor1[0]), .d1(h_arrdiv24_mux2to1280_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1304_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1305_out(.d0(h_arrdiv24_fs318_xor1[0]), .d1(h_arrdiv24_mux2to1281_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1305_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1306_out(.d0(h_arrdiv24_fs319_xor1[0]), .d1(h_arrdiv24_mux2to1282_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1306_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1307_out(.d0(h_arrdiv24_fs320_xor1[0]), .d1(h_arrdiv24_mux2to1283_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1307_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1308_out(.d0(h_arrdiv24_fs321_xor1[0]), .d1(h_arrdiv24_mux2to1284_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1308_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1309_out(.d0(h_arrdiv24_fs322_xor1[0]), .d1(h_arrdiv24_mux2to1285_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1309_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1310_out(.d0(h_arrdiv24_fs323_xor1[0]), .d1(h_arrdiv24_mux2to1286_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1310_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1311_out(.d0(h_arrdiv24_fs324_xor1[0]), .d1(h_arrdiv24_mux2to1287_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1311_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1312_out(.d0(h_arrdiv24_fs325_xor1[0]), .d1(h_arrdiv24_mux2to1288_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1312_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1313_out(.d0(h_arrdiv24_fs326_xor1[0]), .d1(h_arrdiv24_mux2to1289_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1313_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1314_out(.d0(h_arrdiv24_fs327_xor1[0]), .d1(h_arrdiv24_mux2to1290_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1314_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1315_out(.d0(h_arrdiv24_fs328_xor1[0]), .d1(h_arrdiv24_mux2to1291_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1315_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1316_out(.d0(h_arrdiv24_fs329_xor1[0]), .d1(h_arrdiv24_mux2to1292_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1316_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1317_out(.d0(h_arrdiv24_fs330_xor1[0]), .d1(h_arrdiv24_mux2to1293_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1317_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1318_out(.d0(h_arrdiv24_fs331_xor1[0]), .d1(h_arrdiv24_mux2to1294_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1318_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1319_out(.d0(h_arrdiv24_fs332_xor1[0]), .d1(h_arrdiv24_mux2to1295_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1319_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1320_out(.d0(h_arrdiv24_fs333_xor1[0]), .d1(h_arrdiv24_mux2to1296_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1320_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1321_out(.d0(h_arrdiv24_fs334_xor1[0]), .d1(h_arrdiv24_mux2to1297_xor0[0]), .sel(h_arrdiv24_fs335_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1321_xor0));
  not_gate not_gate_h_arrdiv24_not13(.a(h_arrdiv24_fs335_or0[0]), .out(h_arrdiv24_not13));
  fs fs_h_arrdiv24_fs336_out(.a(a[9]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs336_xor0), .fs_or0(h_arrdiv24_fs336_and0));
  fs fs_h_arrdiv24_fs337_out(.a(h_arrdiv24_mux2to1299_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs336_and0[0]), .fs_xor1(h_arrdiv24_fs337_xor1), .fs_or0(h_arrdiv24_fs337_or0));
  fs fs_h_arrdiv24_fs338_out(.a(h_arrdiv24_mux2to1300_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs337_or0[0]), .fs_xor1(h_arrdiv24_fs338_xor1), .fs_or0(h_arrdiv24_fs338_or0));
  fs fs_h_arrdiv24_fs339_out(.a(h_arrdiv24_mux2to1301_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs338_or0[0]), .fs_xor1(h_arrdiv24_fs339_xor1), .fs_or0(h_arrdiv24_fs339_or0));
  fs fs_h_arrdiv24_fs340_out(.a(h_arrdiv24_mux2to1302_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs339_or0[0]), .fs_xor1(h_arrdiv24_fs340_xor1), .fs_or0(h_arrdiv24_fs340_or0));
  fs fs_h_arrdiv24_fs341_out(.a(h_arrdiv24_mux2to1303_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs340_or0[0]), .fs_xor1(h_arrdiv24_fs341_xor1), .fs_or0(h_arrdiv24_fs341_or0));
  fs fs_h_arrdiv24_fs342_out(.a(h_arrdiv24_mux2to1304_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs341_or0[0]), .fs_xor1(h_arrdiv24_fs342_xor1), .fs_or0(h_arrdiv24_fs342_or0));
  fs fs_h_arrdiv24_fs343_out(.a(h_arrdiv24_mux2to1305_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs342_or0[0]), .fs_xor1(h_arrdiv24_fs343_xor1), .fs_or0(h_arrdiv24_fs343_or0));
  fs fs_h_arrdiv24_fs344_out(.a(h_arrdiv24_mux2to1306_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs343_or0[0]), .fs_xor1(h_arrdiv24_fs344_xor1), .fs_or0(h_arrdiv24_fs344_or0));
  fs fs_h_arrdiv24_fs345_out(.a(h_arrdiv24_mux2to1307_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs344_or0[0]), .fs_xor1(h_arrdiv24_fs345_xor1), .fs_or0(h_arrdiv24_fs345_or0));
  fs fs_h_arrdiv24_fs346_out(.a(h_arrdiv24_mux2to1308_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs345_or0[0]), .fs_xor1(h_arrdiv24_fs346_xor1), .fs_or0(h_arrdiv24_fs346_or0));
  fs fs_h_arrdiv24_fs347_out(.a(h_arrdiv24_mux2to1309_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs346_or0[0]), .fs_xor1(h_arrdiv24_fs347_xor1), .fs_or0(h_arrdiv24_fs347_or0));
  fs fs_h_arrdiv24_fs348_out(.a(h_arrdiv24_mux2to1310_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs347_or0[0]), .fs_xor1(h_arrdiv24_fs348_xor1), .fs_or0(h_arrdiv24_fs348_or0));
  fs fs_h_arrdiv24_fs349_out(.a(h_arrdiv24_mux2to1311_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs348_or0[0]), .fs_xor1(h_arrdiv24_fs349_xor1), .fs_or0(h_arrdiv24_fs349_or0));
  fs fs_h_arrdiv24_fs350_out(.a(h_arrdiv24_mux2to1312_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs349_or0[0]), .fs_xor1(h_arrdiv24_fs350_xor1), .fs_or0(h_arrdiv24_fs350_or0));
  fs fs_h_arrdiv24_fs351_out(.a(h_arrdiv24_mux2to1313_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs350_or0[0]), .fs_xor1(h_arrdiv24_fs351_xor1), .fs_or0(h_arrdiv24_fs351_or0));
  fs fs_h_arrdiv24_fs352_out(.a(h_arrdiv24_mux2to1314_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs351_or0[0]), .fs_xor1(h_arrdiv24_fs352_xor1), .fs_or0(h_arrdiv24_fs352_or0));
  fs fs_h_arrdiv24_fs353_out(.a(h_arrdiv24_mux2to1315_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs352_or0[0]), .fs_xor1(h_arrdiv24_fs353_xor1), .fs_or0(h_arrdiv24_fs353_or0));
  fs fs_h_arrdiv24_fs354_out(.a(h_arrdiv24_mux2to1316_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs353_or0[0]), .fs_xor1(h_arrdiv24_fs354_xor1), .fs_or0(h_arrdiv24_fs354_or0));
  fs fs_h_arrdiv24_fs355_out(.a(h_arrdiv24_mux2to1317_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs354_or0[0]), .fs_xor1(h_arrdiv24_fs355_xor1), .fs_or0(h_arrdiv24_fs355_or0));
  fs fs_h_arrdiv24_fs356_out(.a(h_arrdiv24_mux2to1318_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs355_or0[0]), .fs_xor1(h_arrdiv24_fs356_xor1), .fs_or0(h_arrdiv24_fs356_or0));
  fs fs_h_arrdiv24_fs357_out(.a(h_arrdiv24_mux2to1319_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs356_or0[0]), .fs_xor1(h_arrdiv24_fs357_xor1), .fs_or0(h_arrdiv24_fs357_or0));
  fs fs_h_arrdiv24_fs358_out(.a(h_arrdiv24_mux2to1320_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs357_or0[0]), .fs_xor1(h_arrdiv24_fs358_xor1), .fs_or0(h_arrdiv24_fs358_or0));
  fs fs_h_arrdiv24_fs359_out(.a(h_arrdiv24_mux2to1321_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs358_or0[0]), .fs_xor1(h_arrdiv24_fs359_xor1), .fs_or0(h_arrdiv24_fs359_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1322_out(.d0(h_arrdiv24_fs336_xor0[0]), .d1(a[9]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1322_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1323_out(.d0(h_arrdiv24_fs337_xor1[0]), .d1(h_arrdiv24_mux2to1299_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1323_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1324_out(.d0(h_arrdiv24_fs338_xor1[0]), .d1(h_arrdiv24_mux2to1300_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1324_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1325_out(.d0(h_arrdiv24_fs339_xor1[0]), .d1(h_arrdiv24_mux2to1301_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1325_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1326_out(.d0(h_arrdiv24_fs340_xor1[0]), .d1(h_arrdiv24_mux2to1302_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1326_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1327_out(.d0(h_arrdiv24_fs341_xor1[0]), .d1(h_arrdiv24_mux2to1303_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1327_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1328_out(.d0(h_arrdiv24_fs342_xor1[0]), .d1(h_arrdiv24_mux2to1304_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1328_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1329_out(.d0(h_arrdiv24_fs343_xor1[0]), .d1(h_arrdiv24_mux2to1305_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1329_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1330_out(.d0(h_arrdiv24_fs344_xor1[0]), .d1(h_arrdiv24_mux2to1306_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1330_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1331_out(.d0(h_arrdiv24_fs345_xor1[0]), .d1(h_arrdiv24_mux2to1307_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1331_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1332_out(.d0(h_arrdiv24_fs346_xor1[0]), .d1(h_arrdiv24_mux2to1308_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1332_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1333_out(.d0(h_arrdiv24_fs347_xor1[0]), .d1(h_arrdiv24_mux2to1309_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1333_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1334_out(.d0(h_arrdiv24_fs348_xor1[0]), .d1(h_arrdiv24_mux2to1310_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1334_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1335_out(.d0(h_arrdiv24_fs349_xor1[0]), .d1(h_arrdiv24_mux2to1311_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1335_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1336_out(.d0(h_arrdiv24_fs350_xor1[0]), .d1(h_arrdiv24_mux2to1312_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1336_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1337_out(.d0(h_arrdiv24_fs351_xor1[0]), .d1(h_arrdiv24_mux2to1313_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1337_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1338_out(.d0(h_arrdiv24_fs352_xor1[0]), .d1(h_arrdiv24_mux2to1314_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1338_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1339_out(.d0(h_arrdiv24_fs353_xor1[0]), .d1(h_arrdiv24_mux2to1315_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1339_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1340_out(.d0(h_arrdiv24_fs354_xor1[0]), .d1(h_arrdiv24_mux2to1316_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1340_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1341_out(.d0(h_arrdiv24_fs355_xor1[0]), .d1(h_arrdiv24_mux2to1317_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1341_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1342_out(.d0(h_arrdiv24_fs356_xor1[0]), .d1(h_arrdiv24_mux2to1318_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1342_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1343_out(.d0(h_arrdiv24_fs357_xor1[0]), .d1(h_arrdiv24_mux2to1319_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1343_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1344_out(.d0(h_arrdiv24_fs358_xor1[0]), .d1(h_arrdiv24_mux2to1320_xor0[0]), .sel(h_arrdiv24_fs359_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1344_xor0));
  not_gate not_gate_h_arrdiv24_not14(.a(h_arrdiv24_fs359_or0[0]), .out(h_arrdiv24_not14));
  fs fs_h_arrdiv24_fs360_out(.a(a[8]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs360_xor0), .fs_or0(h_arrdiv24_fs360_and0));
  fs fs_h_arrdiv24_fs361_out(.a(h_arrdiv24_mux2to1322_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs360_and0[0]), .fs_xor1(h_arrdiv24_fs361_xor1), .fs_or0(h_arrdiv24_fs361_or0));
  fs fs_h_arrdiv24_fs362_out(.a(h_arrdiv24_mux2to1323_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs361_or0[0]), .fs_xor1(h_arrdiv24_fs362_xor1), .fs_or0(h_arrdiv24_fs362_or0));
  fs fs_h_arrdiv24_fs363_out(.a(h_arrdiv24_mux2to1324_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs362_or0[0]), .fs_xor1(h_arrdiv24_fs363_xor1), .fs_or0(h_arrdiv24_fs363_or0));
  fs fs_h_arrdiv24_fs364_out(.a(h_arrdiv24_mux2to1325_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs363_or0[0]), .fs_xor1(h_arrdiv24_fs364_xor1), .fs_or0(h_arrdiv24_fs364_or0));
  fs fs_h_arrdiv24_fs365_out(.a(h_arrdiv24_mux2to1326_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs364_or0[0]), .fs_xor1(h_arrdiv24_fs365_xor1), .fs_or0(h_arrdiv24_fs365_or0));
  fs fs_h_arrdiv24_fs366_out(.a(h_arrdiv24_mux2to1327_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs365_or0[0]), .fs_xor1(h_arrdiv24_fs366_xor1), .fs_or0(h_arrdiv24_fs366_or0));
  fs fs_h_arrdiv24_fs367_out(.a(h_arrdiv24_mux2to1328_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs366_or0[0]), .fs_xor1(h_arrdiv24_fs367_xor1), .fs_or0(h_arrdiv24_fs367_or0));
  fs fs_h_arrdiv24_fs368_out(.a(h_arrdiv24_mux2to1329_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs367_or0[0]), .fs_xor1(h_arrdiv24_fs368_xor1), .fs_or0(h_arrdiv24_fs368_or0));
  fs fs_h_arrdiv24_fs369_out(.a(h_arrdiv24_mux2to1330_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs368_or0[0]), .fs_xor1(h_arrdiv24_fs369_xor1), .fs_or0(h_arrdiv24_fs369_or0));
  fs fs_h_arrdiv24_fs370_out(.a(h_arrdiv24_mux2to1331_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs369_or0[0]), .fs_xor1(h_arrdiv24_fs370_xor1), .fs_or0(h_arrdiv24_fs370_or0));
  fs fs_h_arrdiv24_fs371_out(.a(h_arrdiv24_mux2to1332_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs370_or0[0]), .fs_xor1(h_arrdiv24_fs371_xor1), .fs_or0(h_arrdiv24_fs371_or0));
  fs fs_h_arrdiv24_fs372_out(.a(h_arrdiv24_mux2to1333_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs371_or0[0]), .fs_xor1(h_arrdiv24_fs372_xor1), .fs_or0(h_arrdiv24_fs372_or0));
  fs fs_h_arrdiv24_fs373_out(.a(h_arrdiv24_mux2to1334_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs372_or0[0]), .fs_xor1(h_arrdiv24_fs373_xor1), .fs_or0(h_arrdiv24_fs373_or0));
  fs fs_h_arrdiv24_fs374_out(.a(h_arrdiv24_mux2to1335_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs373_or0[0]), .fs_xor1(h_arrdiv24_fs374_xor1), .fs_or0(h_arrdiv24_fs374_or0));
  fs fs_h_arrdiv24_fs375_out(.a(h_arrdiv24_mux2to1336_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs374_or0[0]), .fs_xor1(h_arrdiv24_fs375_xor1), .fs_or0(h_arrdiv24_fs375_or0));
  fs fs_h_arrdiv24_fs376_out(.a(h_arrdiv24_mux2to1337_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs375_or0[0]), .fs_xor1(h_arrdiv24_fs376_xor1), .fs_or0(h_arrdiv24_fs376_or0));
  fs fs_h_arrdiv24_fs377_out(.a(h_arrdiv24_mux2to1338_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs376_or0[0]), .fs_xor1(h_arrdiv24_fs377_xor1), .fs_or0(h_arrdiv24_fs377_or0));
  fs fs_h_arrdiv24_fs378_out(.a(h_arrdiv24_mux2to1339_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs377_or0[0]), .fs_xor1(h_arrdiv24_fs378_xor1), .fs_or0(h_arrdiv24_fs378_or0));
  fs fs_h_arrdiv24_fs379_out(.a(h_arrdiv24_mux2to1340_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs378_or0[0]), .fs_xor1(h_arrdiv24_fs379_xor1), .fs_or0(h_arrdiv24_fs379_or0));
  fs fs_h_arrdiv24_fs380_out(.a(h_arrdiv24_mux2to1341_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs379_or0[0]), .fs_xor1(h_arrdiv24_fs380_xor1), .fs_or0(h_arrdiv24_fs380_or0));
  fs fs_h_arrdiv24_fs381_out(.a(h_arrdiv24_mux2to1342_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs380_or0[0]), .fs_xor1(h_arrdiv24_fs381_xor1), .fs_or0(h_arrdiv24_fs381_or0));
  fs fs_h_arrdiv24_fs382_out(.a(h_arrdiv24_mux2to1343_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs381_or0[0]), .fs_xor1(h_arrdiv24_fs382_xor1), .fs_or0(h_arrdiv24_fs382_or0));
  fs fs_h_arrdiv24_fs383_out(.a(h_arrdiv24_mux2to1344_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs382_or0[0]), .fs_xor1(h_arrdiv24_fs383_xor1), .fs_or0(h_arrdiv24_fs383_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1345_out(.d0(h_arrdiv24_fs360_xor0[0]), .d1(a[8]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1345_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1346_out(.d0(h_arrdiv24_fs361_xor1[0]), .d1(h_arrdiv24_mux2to1322_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1346_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1347_out(.d0(h_arrdiv24_fs362_xor1[0]), .d1(h_arrdiv24_mux2to1323_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1347_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1348_out(.d0(h_arrdiv24_fs363_xor1[0]), .d1(h_arrdiv24_mux2to1324_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1348_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1349_out(.d0(h_arrdiv24_fs364_xor1[0]), .d1(h_arrdiv24_mux2to1325_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1349_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1350_out(.d0(h_arrdiv24_fs365_xor1[0]), .d1(h_arrdiv24_mux2to1326_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1350_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1351_out(.d0(h_arrdiv24_fs366_xor1[0]), .d1(h_arrdiv24_mux2to1327_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1351_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1352_out(.d0(h_arrdiv24_fs367_xor1[0]), .d1(h_arrdiv24_mux2to1328_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1352_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1353_out(.d0(h_arrdiv24_fs368_xor1[0]), .d1(h_arrdiv24_mux2to1329_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1353_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1354_out(.d0(h_arrdiv24_fs369_xor1[0]), .d1(h_arrdiv24_mux2to1330_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1354_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1355_out(.d0(h_arrdiv24_fs370_xor1[0]), .d1(h_arrdiv24_mux2to1331_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1355_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1356_out(.d0(h_arrdiv24_fs371_xor1[0]), .d1(h_arrdiv24_mux2to1332_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1356_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1357_out(.d0(h_arrdiv24_fs372_xor1[0]), .d1(h_arrdiv24_mux2to1333_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1357_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1358_out(.d0(h_arrdiv24_fs373_xor1[0]), .d1(h_arrdiv24_mux2to1334_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1358_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1359_out(.d0(h_arrdiv24_fs374_xor1[0]), .d1(h_arrdiv24_mux2to1335_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1359_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1360_out(.d0(h_arrdiv24_fs375_xor1[0]), .d1(h_arrdiv24_mux2to1336_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1360_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1361_out(.d0(h_arrdiv24_fs376_xor1[0]), .d1(h_arrdiv24_mux2to1337_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1361_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1362_out(.d0(h_arrdiv24_fs377_xor1[0]), .d1(h_arrdiv24_mux2to1338_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1362_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1363_out(.d0(h_arrdiv24_fs378_xor1[0]), .d1(h_arrdiv24_mux2to1339_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1363_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1364_out(.d0(h_arrdiv24_fs379_xor1[0]), .d1(h_arrdiv24_mux2to1340_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1364_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1365_out(.d0(h_arrdiv24_fs380_xor1[0]), .d1(h_arrdiv24_mux2to1341_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1365_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1366_out(.d0(h_arrdiv24_fs381_xor1[0]), .d1(h_arrdiv24_mux2to1342_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1366_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1367_out(.d0(h_arrdiv24_fs382_xor1[0]), .d1(h_arrdiv24_mux2to1343_xor0[0]), .sel(h_arrdiv24_fs383_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1367_xor0));
  not_gate not_gate_h_arrdiv24_not15(.a(h_arrdiv24_fs383_or0[0]), .out(h_arrdiv24_not15));
  fs fs_h_arrdiv24_fs384_out(.a(a[7]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs384_xor0), .fs_or0(h_arrdiv24_fs384_and0));
  fs fs_h_arrdiv24_fs385_out(.a(h_arrdiv24_mux2to1345_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs384_and0[0]), .fs_xor1(h_arrdiv24_fs385_xor1), .fs_or0(h_arrdiv24_fs385_or0));
  fs fs_h_arrdiv24_fs386_out(.a(h_arrdiv24_mux2to1346_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs385_or0[0]), .fs_xor1(h_arrdiv24_fs386_xor1), .fs_or0(h_arrdiv24_fs386_or0));
  fs fs_h_arrdiv24_fs387_out(.a(h_arrdiv24_mux2to1347_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs386_or0[0]), .fs_xor1(h_arrdiv24_fs387_xor1), .fs_or0(h_arrdiv24_fs387_or0));
  fs fs_h_arrdiv24_fs388_out(.a(h_arrdiv24_mux2to1348_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs387_or0[0]), .fs_xor1(h_arrdiv24_fs388_xor1), .fs_or0(h_arrdiv24_fs388_or0));
  fs fs_h_arrdiv24_fs389_out(.a(h_arrdiv24_mux2to1349_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs388_or0[0]), .fs_xor1(h_arrdiv24_fs389_xor1), .fs_or0(h_arrdiv24_fs389_or0));
  fs fs_h_arrdiv24_fs390_out(.a(h_arrdiv24_mux2to1350_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs389_or0[0]), .fs_xor1(h_arrdiv24_fs390_xor1), .fs_or0(h_arrdiv24_fs390_or0));
  fs fs_h_arrdiv24_fs391_out(.a(h_arrdiv24_mux2to1351_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs390_or0[0]), .fs_xor1(h_arrdiv24_fs391_xor1), .fs_or0(h_arrdiv24_fs391_or0));
  fs fs_h_arrdiv24_fs392_out(.a(h_arrdiv24_mux2to1352_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs391_or0[0]), .fs_xor1(h_arrdiv24_fs392_xor1), .fs_or0(h_arrdiv24_fs392_or0));
  fs fs_h_arrdiv24_fs393_out(.a(h_arrdiv24_mux2to1353_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs392_or0[0]), .fs_xor1(h_arrdiv24_fs393_xor1), .fs_or0(h_arrdiv24_fs393_or0));
  fs fs_h_arrdiv24_fs394_out(.a(h_arrdiv24_mux2to1354_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs393_or0[0]), .fs_xor1(h_arrdiv24_fs394_xor1), .fs_or0(h_arrdiv24_fs394_or0));
  fs fs_h_arrdiv24_fs395_out(.a(h_arrdiv24_mux2to1355_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs394_or0[0]), .fs_xor1(h_arrdiv24_fs395_xor1), .fs_or0(h_arrdiv24_fs395_or0));
  fs fs_h_arrdiv24_fs396_out(.a(h_arrdiv24_mux2to1356_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs395_or0[0]), .fs_xor1(h_arrdiv24_fs396_xor1), .fs_or0(h_arrdiv24_fs396_or0));
  fs fs_h_arrdiv24_fs397_out(.a(h_arrdiv24_mux2to1357_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs396_or0[0]), .fs_xor1(h_arrdiv24_fs397_xor1), .fs_or0(h_arrdiv24_fs397_or0));
  fs fs_h_arrdiv24_fs398_out(.a(h_arrdiv24_mux2to1358_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs397_or0[0]), .fs_xor1(h_arrdiv24_fs398_xor1), .fs_or0(h_arrdiv24_fs398_or0));
  fs fs_h_arrdiv24_fs399_out(.a(h_arrdiv24_mux2to1359_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs398_or0[0]), .fs_xor1(h_arrdiv24_fs399_xor1), .fs_or0(h_arrdiv24_fs399_or0));
  fs fs_h_arrdiv24_fs400_out(.a(h_arrdiv24_mux2to1360_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs399_or0[0]), .fs_xor1(h_arrdiv24_fs400_xor1), .fs_or0(h_arrdiv24_fs400_or0));
  fs fs_h_arrdiv24_fs401_out(.a(h_arrdiv24_mux2to1361_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs400_or0[0]), .fs_xor1(h_arrdiv24_fs401_xor1), .fs_or0(h_arrdiv24_fs401_or0));
  fs fs_h_arrdiv24_fs402_out(.a(h_arrdiv24_mux2to1362_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs401_or0[0]), .fs_xor1(h_arrdiv24_fs402_xor1), .fs_or0(h_arrdiv24_fs402_or0));
  fs fs_h_arrdiv24_fs403_out(.a(h_arrdiv24_mux2to1363_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs402_or0[0]), .fs_xor1(h_arrdiv24_fs403_xor1), .fs_or0(h_arrdiv24_fs403_or0));
  fs fs_h_arrdiv24_fs404_out(.a(h_arrdiv24_mux2to1364_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs403_or0[0]), .fs_xor1(h_arrdiv24_fs404_xor1), .fs_or0(h_arrdiv24_fs404_or0));
  fs fs_h_arrdiv24_fs405_out(.a(h_arrdiv24_mux2to1365_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs404_or0[0]), .fs_xor1(h_arrdiv24_fs405_xor1), .fs_or0(h_arrdiv24_fs405_or0));
  fs fs_h_arrdiv24_fs406_out(.a(h_arrdiv24_mux2to1366_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs405_or0[0]), .fs_xor1(h_arrdiv24_fs406_xor1), .fs_or0(h_arrdiv24_fs406_or0));
  fs fs_h_arrdiv24_fs407_out(.a(h_arrdiv24_mux2to1367_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs406_or0[0]), .fs_xor1(h_arrdiv24_fs407_xor1), .fs_or0(h_arrdiv24_fs407_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1368_out(.d0(h_arrdiv24_fs384_xor0[0]), .d1(a[7]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1368_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1369_out(.d0(h_arrdiv24_fs385_xor1[0]), .d1(h_arrdiv24_mux2to1345_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1369_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1370_out(.d0(h_arrdiv24_fs386_xor1[0]), .d1(h_arrdiv24_mux2to1346_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1370_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1371_out(.d0(h_arrdiv24_fs387_xor1[0]), .d1(h_arrdiv24_mux2to1347_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1371_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1372_out(.d0(h_arrdiv24_fs388_xor1[0]), .d1(h_arrdiv24_mux2to1348_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1372_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1373_out(.d0(h_arrdiv24_fs389_xor1[0]), .d1(h_arrdiv24_mux2to1349_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1373_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1374_out(.d0(h_arrdiv24_fs390_xor1[0]), .d1(h_arrdiv24_mux2to1350_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1374_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1375_out(.d0(h_arrdiv24_fs391_xor1[0]), .d1(h_arrdiv24_mux2to1351_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1375_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1376_out(.d0(h_arrdiv24_fs392_xor1[0]), .d1(h_arrdiv24_mux2to1352_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1376_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1377_out(.d0(h_arrdiv24_fs393_xor1[0]), .d1(h_arrdiv24_mux2to1353_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1377_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1378_out(.d0(h_arrdiv24_fs394_xor1[0]), .d1(h_arrdiv24_mux2to1354_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1378_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1379_out(.d0(h_arrdiv24_fs395_xor1[0]), .d1(h_arrdiv24_mux2to1355_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1379_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1380_out(.d0(h_arrdiv24_fs396_xor1[0]), .d1(h_arrdiv24_mux2to1356_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1380_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1381_out(.d0(h_arrdiv24_fs397_xor1[0]), .d1(h_arrdiv24_mux2to1357_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1381_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1382_out(.d0(h_arrdiv24_fs398_xor1[0]), .d1(h_arrdiv24_mux2to1358_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1382_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1383_out(.d0(h_arrdiv24_fs399_xor1[0]), .d1(h_arrdiv24_mux2to1359_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1383_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1384_out(.d0(h_arrdiv24_fs400_xor1[0]), .d1(h_arrdiv24_mux2to1360_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1384_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1385_out(.d0(h_arrdiv24_fs401_xor1[0]), .d1(h_arrdiv24_mux2to1361_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1385_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1386_out(.d0(h_arrdiv24_fs402_xor1[0]), .d1(h_arrdiv24_mux2to1362_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1386_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1387_out(.d0(h_arrdiv24_fs403_xor1[0]), .d1(h_arrdiv24_mux2to1363_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1387_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1388_out(.d0(h_arrdiv24_fs404_xor1[0]), .d1(h_arrdiv24_mux2to1364_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1388_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1389_out(.d0(h_arrdiv24_fs405_xor1[0]), .d1(h_arrdiv24_mux2to1365_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1389_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1390_out(.d0(h_arrdiv24_fs406_xor1[0]), .d1(h_arrdiv24_mux2to1366_xor0[0]), .sel(h_arrdiv24_fs407_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1390_xor0));
  not_gate not_gate_h_arrdiv24_not16(.a(h_arrdiv24_fs407_or0[0]), .out(h_arrdiv24_not16));
  fs fs_h_arrdiv24_fs408_out(.a(a[6]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs408_xor0), .fs_or0(h_arrdiv24_fs408_and0));
  fs fs_h_arrdiv24_fs409_out(.a(h_arrdiv24_mux2to1368_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs408_and0[0]), .fs_xor1(h_arrdiv24_fs409_xor1), .fs_or0(h_arrdiv24_fs409_or0));
  fs fs_h_arrdiv24_fs410_out(.a(h_arrdiv24_mux2to1369_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs409_or0[0]), .fs_xor1(h_arrdiv24_fs410_xor1), .fs_or0(h_arrdiv24_fs410_or0));
  fs fs_h_arrdiv24_fs411_out(.a(h_arrdiv24_mux2to1370_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs410_or0[0]), .fs_xor1(h_arrdiv24_fs411_xor1), .fs_or0(h_arrdiv24_fs411_or0));
  fs fs_h_arrdiv24_fs412_out(.a(h_arrdiv24_mux2to1371_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs411_or0[0]), .fs_xor1(h_arrdiv24_fs412_xor1), .fs_or0(h_arrdiv24_fs412_or0));
  fs fs_h_arrdiv24_fs413_out(.a(h_arrdiv24_mux2to1372_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs412_or0[0]), .fs_xor1(h_arrdiv24_fs413_xor1), .fs_or0(h_arrdiv24_fs413_or0));
  fs fs_h_arrdiv24_fs414_out(.a(h_arrdiv24_mux2to1373_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs413_or0[0]), .fs_xor1(h_arrdiv24_fs414_xor1), .fs_or0(h_arrdiv24_fs414_or0));
  fs fs_h_arrdiv24_fs415_out(.a(h_arrdiv24_mux2to1374_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs414_or0[0]), .fs_xor1(h_arrdiv24_fs415_xor1), .fs_or0(h_arrdiv24_fs415_or0));
  fs fs_h_arrdiv24_fs416_out(.a(h_arrdiv24_mux2to1375_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs415_or0[0]), .fs_xor1(h_arrdiv24_fs416_xor1), .fs_or0(h_arrdiv24_fs416_or0));
  fs fs_h_arrdiv24_fs417_out(.a(h_arrdiv24_mux2to1376_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs416_or0[0]), .fs_xor1(h_arrdiv24_fs417_xor1), .fs_or0(h_arrdiv24_fs417_or0));
  fs fs_h_arrdiv24_fs418_out(.a(h_arrdiv24_mux2to1377_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs417_or0[0]), .fs_xor1(h_arrdiv24_fs418_xor1), .fs_or0(h_arrdiv24_fs418_or0));
  fs fs_h_arrdiv24_fs419_out(.a(h_arrdiv24_mux2to1378_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs418_or0[0]), .fs_xor1(h_arrdiv24_fs419_xor1), .fs_or0(h_arrdiv24_fs419_or0));
  fs fs_h_arrdiv24_fs420_out(.a(h_arrdiv24_mux2to1379_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs419_or0[0]), .fs_xor1(h_arrdiv24_fs420_xor1), .fs_or0(h_arrdiv24_fs420_or0));
  fs fs_h_arrdiv24_fs421_out(.a(h_arrdiv24_mux2to1380_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs420_or0[0]), .fs_xor1(h_arrdiv24_fs421_xor1), .fs_or0(h_arrdiv24_fs421_or0));
  fs fs_h_arrdiv24_fs422_out(.a(h_arrdiv24_mux2to1381_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs421_or0[0]), .fs_xor1(h_arrdiv24_fs422_xor1), .fs_or0(h_arrdiv24_fs422_or0));
  fs fs_h_arrdiv24_fs423_out(.a(h_arrdiv24_mux2to1382_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs422_or0[0]), .fs_xor1(h_arrdiv24_fs423_xor1), .fs_or0(h_arrdiv24_fs423_or0));
  fs fs_h_arrdiv24_fs424_out(.a(h_arrdiv24_mux2to1383_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs423_or0[0]), .fs_xor1(h_arrdiv24_fs424_xor1), .fs_or0(h_arrdiv24_fs424_or0));
  fs fs_h_arrdiv24_fs425_out(.a(h_arrdiv24_mux2to1384_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs424_or0[0]), .fs_xor1(h_arrdiv24_fs425_xor1), .fs_or0(h_arrdiv24_fs425_or0));
  fs fs_h_arrdiv24_fs426_out(.a(h_arrdiv24_mux2to1385_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs425_or0[0]), .fs_xor1(h_arrdiv24_fs426_xor1), .fs_or0(h_arrdiv24_fs426_or0));
  fs fs_h_arrdiv24_fs427_out(.a(h_arrdiv24_mux2to1386_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs426_or0[0]), .fs_xor1(h_arrdiv24_fs427_xor1), .fs_or0(h_arrdiv24_fs427_or0));
  fs fs_h_arrdiv24_fs428_out(.a(h_arrdiv24_mux2to1387_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs427_or0[0]), .fs_xor1(h_arrdiv24_fs428_xor1), .fs_or0(h_arrdiv24_fs428_or0));
  fs fs_h_arrdiv24_fs429_out(.a(h_arrdiv24_mux2to1388_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs428_or0[0]), .fs_xor1(h_arrdiv24_fs429_xor1), .fs_or0(h_arrdiv24_fs429_or0));
  fs fs_h_arrdiv24_fs430_out(.a(h_arrdiv24_mux2to1389_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs429_or0[0]), .fs_xor1(h_arrdiv24_fs430_xor1), .fs_or0(h_arrdiv24_fs430_or0));
  fs fs_h_arrdiv24_fs431_out(.a(h_arrdiv24_mux2to1390_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs430_or0[0]), .fs_xor1(h_arrdiv24_fs431_xor1), .fs_or0(h_arrdiv24_fs431_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1391_out(.d0(h_arrdiv24_fs408_xor0[0]), .d1(a[6]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1391_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1392_out(.d0(h_arrdiv24_fs409_xor1[0]), .d1(h_arrdiv24_mux2to1368_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1392_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1393_out(.d0(h_arrdiv24_fs410_xor1[0]), .d1(h_arrdiv24_mux2to1369_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1393_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1394_out(.d0(h_arrdiv24_fs411_xor1[0]), .d1(h_arrdiv24_mux2to1370_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1394_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1395_out(.d0(h_arrdiv24_fs412_xor1[0]), .d1(h_arrdiv24_mux2to1371_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1395_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1396_out(.d0(h_arrdiv24_fs413_xor1[0]), .d1(h_arrdiv24_mux2to1372_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1396_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1397_out(.d0(h_arrdiv24_fs414_xor1[0]), .d1(h_arrdiv24_mux2to1373_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1397_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1398_out(.d0(h_arrdiv24_fs415_xor1[0]), .d1(h_arrdiv24_mux2to1374_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1398_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1399_out(.d0(h_arrdiv24_fs416_xor1[0]), .d1(h_arrdiv24_mux2to1375_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1399_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1400_out(.d0(h_arrdiv24_fs417_xor1[0]), .d1(h_arrdiv24_mux2to1376_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1400_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1401_out(.d0(h_arrdiv24_fs418_xor1[0]), .d1(h_arrdiv24_mux2to1377_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1401_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1402_out(.d0(h_arrdiv24_fs419_xor1[0]), .d1(h_arrdiv24_mux2to1378_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1402_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1403_out(.d0(h_arrdiv24_fs420_xor1[0]), .d1(h_arrdiv24_mux2to1379_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1403_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1404_out(.d0(h_arrdiv24_fs421_xor1[0]), .d1(h_arrdiv24_mux2to1380_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1404_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1405_out(.d0(h_arrdiv24_fs422_xor1[0]), .d1(h_arrdiv24_mux2to1381_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1405_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1406_out(.d0(h_arrdiv24_fs423_xor1[0]), .d1(h_arrdiv24_mux2to1382_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1406_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1407_out(.d0(h_arrdiv24_fs424_xor1[0]), .d1(h_arrdiv24_mux2to1383_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1407_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1408_out(.d0(h_arrdiv24_fs425_xor1[0]), .d1(h_arrdiv24_mux2to1384_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1408_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1409_out(.d0(h_arrdiv24_fs426_xor1[0]), .d1(h_arrdiv24_mux2to1385_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1409_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1410_out(.d0(h_arrdiv24_fs427_xor1[0]), .d1(h_arrdiv24_mux2to1386_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1410_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1411_out(.d0(h_arrdiv24_fs428_xor1[0]), .d1(h_arrdiv24_mux2to1387_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1411_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1412_out(.d0(h_arrdiv24_fs429_xor1[0]), .d1(h_arrdiv24_mux2to1388_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1412_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1413_out(.d0(h_arrdiv24_fs430_xor1[0]), .d1(h_arrdiv24_mux2to1389_xor0[0]), .sel(h_arrdiv24_fs431_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1413_xor0));
  not_gate not_gate_h_arrdiv24_not17(.a(h_arrdiv24_fs431_or0[0]), .out(h_arrdiv24_not17));
  fs fs_h_arrdiv24_fs432_out(.a(a[5]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs432_xor0), .fs_or0(h_arrdiv24_fs432_and0));
  fs fs_h_arrdiv24_fs433_out(.a(h_arrdiv24_mux2to1391_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs432_and0[0]), .fs_xor1(h_arrdiv24_fs433_xor1), .fs_or0(h_arrdiv24_fs433_or0));
  fs fs_h_arrdiv24_fs434_out(.a(h_arrdiv24_mux2to1392_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs433_or0[0]), .fs_xor1(h_arrdiv24_fs434_xor1), .fs_or0(h_arrdiv24_fs434_or0));
  fs fs_h_arrdiv24_fs435_out(.a(h_arrdiv24_mux2to1393_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs434_or0[0]), .fs_xor1(h_arrdiv24_fs435_xor1), .fs_or0(h_arrdiv24_fs435_or0));
  fs fs_h_arrdiv24_fs436_out(.a(h_arrdiv24_mux2to1394_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs435_or0[0]), .fs_xor1(h_arrdiv24_fs436_xor1), .fs_or0(h_arrdiv24_fs436_or0));
  fs fs_h_arrdiv24_fs437_out(.a(h_arrdiv24_mux2to1395_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs436_or0[0]), .fs_xor1(h_arrdiv24_fs437_xor1), .fs_or0(h_arrdiv24_fs437_or0));
  fs fs_h_arrdiv24_fs438_out(.a(h_arrdiv24_mux2to1396_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs437_or0[0]), .fs_xor1(h_arrdiv24_fs438_xor1), .fs_or0(h_arrdiv24_fs438_or0));
  fs fs_h_arrdiv24_fs439_out(.a(h_arrdiv24_mux2to1397_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs438_or0[0]), .fs_xor1(h_arrdiv24_fs439_xor1), .fs_or0(h_arrdiv24_fs439_or0));
  fs fs_h_arrdiv24_fs440_out(.a(h_arrdiv24_mux2to1398_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs439_or0[0]), .fs_xor1(h_arrdiv24_fs440_xor1), .fs_or0(h_arrdiv24_fs440_or0));
  fs fs_h_arrdiv24_fs441_out(.a(h_arrdiv24_mux2to1399_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs440_or0[0]), .fs_xor1(h_arrdiv24_fs441_xor1), .fs_or0(h_arrdiv24_fs441_or0));
  fs fs_h_arrdiv24_fs442_out(.a(h_arrdiv24_mux2to1400_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs441_or0[0]), .fs_xor1(h_arrdiv24_fs442_xor1), .fs_or0(h_arrdiv24_fs442_or0));
  fs fs_h_arrdiv24_fs443_out(.a(h_arrdiv24_mux2to1401_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs442_or0[0]), .fs_xor1(h_arrdiv24_fs443_xor1), .fs_or0(h_arrdiv24_fs443_or0));
  fs fs_h_arrdiv24_fs444_out(.a(h_arrdiv24_mux2to1402_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs443_or0[0]), .fs_xor1(h_arrdiv24_fs444_xor1), .fs_or0(h_arrdiv24_fs444_or0));
  fs fs_h_arrdiv24_fs445_out(.a(h_arrdiv24_mux2to1403_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs444_or0[0]), .fs_xor1(h_arrdiv24_fs445_xor1), .fs_or0(h_arrdiv24_fs445_or0));
  fs fs_h_arrdiv24_fs446_out(.a(h_arrdiv24_mux2to1404_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs445_or0[0]), .fs_xor1(h_arrdiv24_fs446_xor1), .fs_or0(h_arrdiv24_fs446_or0));
  fs fs_h_arrdiv24_fs447_out(.a(h_arrdiv24_mux2to1405_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs446_or0[0]), .fs_xor1(h_arrdiv24_fs447_xor1), .fs_or0(h_arrdiv24_fs447_or0));
  fs fs_h_arrdiv24_fs448_out(.a(h_arrdiv24_mux2to1406_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs447_or0[0]), .fs_xor1(h_arrdiv24_fs448_xor1), .fs_or0(h_arrdiv24_fs448_or0));
  fs fs_h_arrdiv24_fs449_out(.a(h_arrdiv24_mux2to1407_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs448_or0[0]), .fs_xor1(h_arrdiv24_fs449_xor1), .fs_or0(h_arrdiv24_fs449_or0));
  fs fs_h_arrdiv24_fs450_out(.a(h_arrdiv24_mux2to1408_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs449_or0[0]), .fs_xor1(h_arrdiv24_fs450_xor1), .fs_or0(h_arrdiv24_fs450_or0));
  fs fs_h_arrdiv24_fs451_out(.a(h_arrdiv24_mux2to1409_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs450_or0[0]), .fs_xor1(h_arrdiv24_fs451_xor1), .fs_or0(h_arrdiv24_fs451_or0));
  fs fs_h_arrdiv24_fs452_out(.a(h_arrdiv24_mux2to1410_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs451_or0[0]), .fs_xor1(h_arrdiv24_fs452_xor1), .fs_or0(h_arrdiv24_fs452_or0));
  fs fs_h_arrdiv24_fs453_out(.a(h_arrdiv24_mux2to1411_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs452_or0[0]), .fs_xor1(h_arrdiv24_fs453_xor1), .fs_or0(h_arrdiv24_fs453_or0));
  fs fs_h_arrdiv24_fs454_out(.a(h_arrdiv24_mux2to1412_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs453_or0[0]), .fs_xor1(h_arrdiv24_fs454_xor1), .fs_or0(h_arrdiv24_fs454_or0));
  fs fs_h_arrdiv24_fs455_out(.a(h_arrdiv24_mux2to1413_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs454_or0[0]), .fs_xor1(h_arrdiv24_fs455_xor1), .fs_or0(h_arrdiv24_fs455_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1414_out(.d0(h_arrdiv24_fs432_xor0[0]), .d1(a[5]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1414_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1415_out(.d0(h_arrdiv24_fs433_xor1[0]), .d1(h_arrdiv24_mux2to1391_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1415_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1416_out(.d0(h_arrdiv24_fs434_xor1[0]), .d1(h_arrdiv24_mux2to1392_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1416_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1417_out(.d0(h_arrdiv24_fs435_xor1[0]), .d1(h_arrdiv24_mux2to1393_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1417_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1418_out(.d0(h_arrdiv24_fs436_xor1[0]), .d1(h_arrdiv24_mux2to1394_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1418_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1419_out(.d0(h_arrdiv24_fs437_xor1[0]), .d1(h_arrdiv24_mux2to1395_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1419_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1420_out(.d0(h_arrdiv24_fs438_xor1[0]), .d1(h_arrdiv24_mux2to1396_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1420_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1421_out(.d0(h_arrdiv24_fs439_xor1[0]), .d1(h_arrdiv24_mux2to1397_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1421_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1422_out(.d0(h_arrdiv24_fs440_xor1[0]), .d1(h_arrdiv24_mux2to1398_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1422_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1423_out(.d0(h_arrdiv24_fs441_xor1[0]), .d1(h_arrdiv24_mux2to1399_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1423_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1424_out(.d0(h_arrdiv24_fs442_xor1[0]), .d1(h_arrdiv24_mux2to1400_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1424_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1425_out(.d0(h_arrdiv24_fs443_xor1[0]), .d1(h_arrdiv24_mux2to1401_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1425_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1426_out(.d0(h_arrdiv24_fs444_xor1[0]), .d1(h_arrdiv24_mux2to1402_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1426_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1427_out(.d0(h_arrdiv24_fs445_xor1[0]), .d1(h_arrdiv24_mux2to1403_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1427_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1428_out(.d0(h_arrdiv24_fs446_xor1[0]), .d1(h_arrdiv24_mux2to1404_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1428_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1429_out(.d0(h_arrdiv24_fs447_xor1[0]), .d1(h_arrdiv24_mux2to1405_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1429_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1430_out(.d0(h_arrdiv24_fs448_xor1[0]), .d1(h_arrdiv24_mux2to1406_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1430_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1431_out(.d0(h_arrdiv24_fs449_xor1[0]), .d1(h_arrdiv24_mux2to1407_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1431_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1432_out(.d0(h_arrdiv24_fs450_xor1[0]), .d1(h_arrdiv24_mux2to1408_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1432_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1433_out(.d0(h_arrdiv24_fs451_xor1[0]), .d1(h_arrdiv24_mux2to1409_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1433_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1434_out(.d0(h_arrdiv24_fs452_xor1[0]), .d1(h_arrdiv24_mux2to1410_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1434_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1435_out(.d0(h_arrdiv24_fs453_xor1[0]), .d1(h_arrdiv24_mux2to1411_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1435_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1436_out(.d0(h_arrdiv24_fs454_xor1[0]), .d1(h_arrdiv24_mux2to1412_xor0[0]), .sel(h_arrdiv24_fs455_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1436_xor0));
  not_gate not_gate_h_arrdiv24_not18(.a(h_arrdiv24_fs455_or0[0]), .out(h_arrdiv24_not18));
  fs fs_h_arrdiv24_fs456_out(.a(a[4]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs456_xor0), .fs_or0(h_arrdiv24_fs456_and0));
  fs fs_h_arrdiv24_fs457_out(.a(h_arrdiv24_mux2to1414_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs456_and0[0]), .fs_xor1(h_arrdiv24_fs457_xor1), .fs_or0(h_arrdiv24_fs457_or0));
  fs fs_h_arrdiv24_fs458_out(.a(h_arrdiv24_mux2to1415_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs457_or0[0]), .fs_xor1(h_arrdiv24_fs458_xor1), .fs_or0(h_arrdiv24_fs458_or0));
  fs fs_h_arrdiv24_fs459_out(.a(h_arrdiv24_mux2to1416_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs458_or0[0]), .fs_xor1(h_arrdiv24_fs459_xor1), .fs_or0(h_arrdiv24_fs459_or0));
  fs fs_h_arrdiv24_fs460_out(.a(h_arrdiv24_mux2to1417_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs459_or0[0]), .fs_xor1(h_arrdiv24_fs460_xor1), .fs_or0(h_arrdiv24_fs460_or0));
  fs fs_h_arrdiv24_fs461_out(.a(h_arrdiv24_mux2to1418_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs460_or0[0]), .fs_xor1(h_arrdiv24_fs461_xor1), .fs_or0(h_arrdiv24_fs461_or0));
  fs fs_h_arrdiv24_fs462_out(.a(h_arrdiv24_mux2to1419_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs461_or0[0]), .fs_xor1(h_arrdiv24_fs462_xor1), .fs_or0(h_arrdiv24_fs462_or0));
  fs fs_h_arrdiv24_fs463_out(.a(h_arrdiv24_mux2to1420_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs462_or0[0]), .fs_xor1(h_arrdiv24_fs463_xor1), .fs_or0(h_arrdiv24_fs463_or0));
  fs fs_h_arrdiv24_fs464_out(.a(h_arrdiv24_mux2to1421_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs463_or0[0]), .fs_xor1(h_arrdiv24_fs464_xor1), .fs_or0(h_arrdiv24_fs464_or0));
  fs fs_h_arrdiv24_fs465_out(.a(h_arrdiv24_mux2to1422_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs464_or0[0]), .fs_xor1(h_arrdiv24_fs465_xor1), .fs_or0(h_arrdiv24_fs465_or0));
  fs fs_h_arrdiv24_fs466_out(.a(h_arrdiv24_mux2to1423_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs465_or0[0]), .fs_xor1(h_arrdiv24_fs466_xor1), .fs_or0(h_arrdiv24_fs466_or0));
  fs fs_h_arrdiv24_fs467_out(.a(h_arrdiv24_mux2to1424_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs466_or0[0]), .fs_xor1(h_arrdiv24_fs467_xor1), .fs_or0(h_arrdiv24_fs467_or0));
  fs fs_h_arrdiv24_fs468_out(.a(h_arrdiv24_mux2to1425_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs467_or0[0]), .fs_xor1(h_arrdiv24_fs468_xor1), .fs_or0(h_arrdiv24_fs468_or0));
  fs fs_h_arrdiv24_fs469_out(.a(h_arrdiv24_mux2to1426_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs468_or0[0]), .fs_xor1(h_arrdiv24_fs469_xor1), .fs_or0(h_arrdiv24_fs469_or0));
  fs fs_h_arrdiv24_fs470_out(.a(h_arrdiv24_mux2to1427_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs469_or0[0]), .fs_xor1(h_arrdiv24_fs470_xor1), .fs_or0(h_arrdiv24_fs470_or0));
  fs fs_h_arrdiv24_fs471_out(.a(h_arrdiv24_mux2to1428_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs470_or0[0]), .fs_xor1(h_arrdiv24_fs471_xor1), .fs_or0(h_arrdiv24_fs471_or0));
  fs fs_h_arrdiv24_fs472_out(.a(h_arrdiv24_mux2to1429_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs471_or0[0]), .fs_xor1(h_arrdiv24_fs472_xor1), .fs_or0(h_arrdiv24_fs472_or0));
  fs fs_h_arrdiv24_fs473_out(.a(h_arrdiv24_mux2to1430_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs472_or0[0]), .fs_xor1(h_arrdiv24_fs473_xor1), .fs_or0(h_arrdiv24_fs473_or0));
  fs fs_h_arrdiv24_fs474_out(.a(h_arrdiv24_mux2to1431_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs473_or0[0]), .fs_xor1(h_arrdiv24_fs474_xor1), .fs_or0(h_arrdiv24_fs474_or0));
  fs fs_h_arrdiv24_fs475_out(.a(h_arrdiv24_mux2to1432_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs474_or0[0]), .fs_xor1(h_arrdiv24_fs475_xor1), .fs_or0(h_arrdiv24_fs475_or0));
  fs fs_h_arrdiv24_fs476_out(.a(h_arrdiv24_mux2to1433_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs475_or0[0]), .fs_xor1(h_arrdiv24_fs476_xor1), .fs_or0(h_arrdiv24_fs476_or0));
  fs fs_h_arrdiv24_fs477_out(.a(h_arrdiv24_mux2to1434_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs476_or0[0]), .fs_xor1(h_arrdiv24_fs477_xor1), .fs_or0(h_arrdiv24_fs477_or0));
  fs fs_h_arrdiv24_fs478_out(.a(h_arrdiv24_mux2to1435_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs477_or0[0]), .fs_xor1(h_arrdiv24_fs478_xor1), .fs_or0(h_arrdiv24_fs478_or0));
  fs fs_h_arrdiv24_fs479_out(.a(h_arrdiv24_mux2to1436_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs478_or0[0]), .fs_xor1(h_arrdiv24_fs479_xor1), .fs_or0(h_arrdiv24_fs479_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1437_out(.d0(h_arrdiv24_fs456_xor0[0]), .d1(a[4]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1437_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1438_out(.d0(h_arrdiv24_fs457_xor1[0]), .d1(h_arrdiv24_mux2to1414_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1438_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1439_out(.d0(h_arrdiv24_fs458_xor1[0]), .d1(h_arrdiv24_mux2to1415_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1439_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1440_out(.d0(h_arrdiv24_fs459_xor1[0]), .d1(h_arrdiv24_mux2to1416_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1440_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1441_out(.d0(h_arrdiv24_fs460_xor1[0]), .d1(h_arrdiv24_mux2to1417_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1441_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1442_out(.d0(h_arrdiv24_fs461_xor1[0]), .d1(h_arrdiv24_mux2to1418_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1442_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1443_out(.d0(h_arrdiv24_fs462_xor1[0]), .d1(h_arrdiv24_mux2to1419_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1443_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1444_out(.d0(h_arrdiv24_fs463_xor1[0]), .d1(h_arrdiv24_mux2to1420_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1444_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1445_out(.d0(h_arrdiv24_fs464_xor1[0]), .d1(h_arrdiv24_mux2to1421_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1445_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1446_out(.d0(h_arrdiv24_fs465_xor1[0]), .d1(h_arrdiv24_mux2to1422_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1446_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1447_out(.d0(h_arrdiv24_fs466_xor1[0]), .d1(h_arrdiv24_mux2to1423_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1447_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1448_out(.d0(h_arrdiv24_fs467_xor1[0]), .d1(h_arrdiv24_mux2to1424_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1448_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1449_out(.d0(h_arrdiv24_fs468_xor1[0]), .d1(h_arrdiv24_mux2to1425_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1449_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1450_out(.d0(h_arrdiv24_fs469_xor1[0]), .d1(h_arrdiv24_mux2to1426_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1450_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1451_out(.d0(h_arrdiv24_fs470_xor1[0]), .d1(h_arrdiv24_mux2to1427_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1451_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1452_out(.d0(h_arrdiv24_fs471_xor1[0]), .d1(h_arrdiv24_mux2to1428_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1452_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1453_out(.d0(h_arrdiv24_fs472_xor1[0]), .d1(h_arrdiv24_mux2to1429_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1453_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1454_out(.d0(h_arrdiv24_fs473_xor1[0]), .d1(h_arrdiv24_mux2to1430_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1454_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1455_out(.d0(h_arrdiv24_fs474_xor1[0]), .d1(h_arrdiv24_mux2to1431_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1455_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1456_out(.d0(h_arrdiv24_fs475_xor1[0]), .d1(h_arrdiv24_mux2to1432_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1456_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1457_out(.d0(h_arrdiv24_fs476_xor1[0]), .d1(h_arrdiv24_mux2to1433_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1457_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1458_out(.d0(h_arrdiv24_fs477_xor1[0]), .d1(h_arrdiv24_mux2to1434_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1458_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1459_out(.d0(h_arrdiv24_fs478_xor1[0]), .d1(h_arrdiv24_mux2to1435_xor0[0]), .sel(h_arrdiv24_fs479_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1459_xor0));
  not_gate not_gate_h_arrdiv24_not19(.a(h_arrdiv24_fs479_or0[0]), .out(h_arrdiv24_not19));
  fs fs_h_arrdiv24_fs480_out(.a(a[3]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs480_xor0), .fs_or0(h_arrdiv24_fs480_and0));
  fs fs_h_arrdiv24_fs481_out(.a(h_arrdiv24_mux2to1437_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs480_and0[0]), .fs_xor1(h_arrdiv24_fs481_xor1), .fs_or0(h_arrdiv24_fs481_or0));
  fs fs_h_arrdiv24_fs482_out(.a(h_arrdiv24_mux2to1438_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs481_or0[0]), .fs_xor1(h_arrdiv24_fs482_xor1), .fs_or0(h_arrdiv24_fs482_or0));
  fs fs_h_arrdiv24_fs483_out(.a(h_arrdiv24_mux2to1439_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs482_or0[0]), .fs_xor1(h_arrdiv24_fs483_xor1), .fs_or0(h_arrdiv24_fs483_or0));
  fs fs_h_arrdiv24_fs484_out(.a(h_arrdiv24_mux2to1440_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs483_or0[0]), .fs_xor1(h_arrdiv24_fs484_xor1), .fs_or0(h_arrdiv24_fs484_or0));
  fs fs_h_arrdiv24_fs485_out(.a(h_arrdiv24_mux2to1441_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs484_or0[0]), .fs_xor1(h_arrdiv24_fs485_xor1), .fs_or0(h_arrdiv24_fs485_or0));
  fs fs_h_arrdiv24_fs486_out(.a(h_arrdiv24_mux2to1442_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs485_or0[0]), .fs_xor1(h_arrdiv24_fs486_xor1), .fs_or0(h_arrdiv24_fs486_or0));
  fs fs_h_arrdiv24_fs487_out(.a(h_arrdiv24_mux2to1443_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs486_or0[0]), .fs_xor1(h_arrdiv24_fs487_xor1), .fs_or0(h_arrdiv24_fs487_or0));
  fs fs_h_arrdiv24_fs488_out(.a(h_arrdiv24_mux2to1444_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs487_or0[0]), .fs_xor1(h_arrdiv24_fs488_xor1), .fs_or0(h_arrdiv24_fs488_or0));
  fs fs_h_arrdiv24_fs489_out(.a(h_arrdiv24_mux2to1445_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs488_or0[0]), .fs_xor1(h_arrdiv24_fs489_xor1), .fs_or0(h_arrdiv24_fs489_or0));
  fs fs_h_arrdiv24_fs490_out(.a(h_arrdiv24_mux2to1446_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs489_or0[0]), .fs_xor1(h_arrdiv24_fs490_xor1), .fs_or0(h_arrdiv24_fs490_or0));
  fs fs_h_arrdiv24_fs491_out(.a(h_arrdiv24_mux2to1447_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs490_or0[0]), .fs_xor1(h_arrdiv24_fs491_xor1), .fs_or0(h_arrdiv24_fs491_or0));
  fs fs_h_arrdiv24_fs492_out(.a(h_arrdiv24_mux2to1448_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs491_or0[0]), .fs_xor1(h_arrdiv24_fs492_xor1), .fs_or0(h_arrdiv24_fs492_or0));
  fs fs_h_arrdiv24_fs493_out(.a(h_arrdiv24_mux2to1449_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs492_or0[0]), .fs_xor1(h_arrdiv24_fs493_xor1), .fs_or0(h_arrdiv24_fs493_or0));
  fs fs_h_arrdiv24_fs494_out(.a(h_arrdiv24_mux2to1450_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs493_or0[0]), .fs_xor1(h_arrdiv24_fs494_xor1), .fs_or0(h_arrdiv24_fs494_or0));
  fs fs_h_arrdiv24_fs495_out(.a(h_arrdiv24_mux2to1451_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs494_or0[0]), .fs_xor1(h_arrdiv24_fs495_xor1), .fs_or0(h_arrdiv24_fs495_or0));
  fs fs_h_arrdiv24_fs496_out(.a(h_arrdiv24_mux2to1452_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs495_or0[0]), .fs_xor1(h_arrdiv24_fs496_xor1), .fs_or0(h_arrdiv24_fs496_or0));
  fs fs_h_arrdiv24_fs497_out(.a(h_arrdiv24_mux2to1453_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs496_or0[0]), .fs_xor1(h_arrdiv24_fs497_xor1), .fs_or0(h_arrdiv24_fs497_or0));
  fs fs_h_arrdiv24_fs498_out(.a(h_arrdiv24_mux2to1454_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs497_or0[0]), .fs_xor1(h_arrdiv24_fs498_xor1), .fs_or0(h_arrdiv24_fs498_or0));
  fs fs_h_arrdiv24_fs499_out(.a(h_arrdiv24_mux2to1455_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs498_or0[0]), .fs_xor1(h_arrdiv24_fs499_xor1), .fs_or0(h_arrdiv24_fs499_or0));
  fs fs_h_arrdiv24_fs500_out(.a(h_arrdiv24_mux2to1456_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs499_or0[0]), .fs_xor1(h_arrdiv24_fs500_xor1), .fs_or0(h_arrdiv24_fs500_or0));
  fs fs_h_arrdiv24_fs501_out(.a(h_arrdiv24_mux2to1457_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs500_or0[0]), .fs_xor1(h_arrdiv24_fs501_xor1), .fs_or0(h_arrdiv24_fs501_or0));
  fs fs_h_arrdiv24_fs502_out(.a(h_arrdiv24_mux2to1458_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs501_or0[0]), .fs_xor1(h_arrdiv24_fs502_xor1), .fs_or0(h_arrdiv24_fs502_or0));
  fs fs_h_arrdiv24_fs503_out(.a(h_arrdiv24_mux2to1459_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs502_or0[0]), .fs_xor1(h_arrdiv24_fs503_xor1), .fs_or0(h_arrdiv24_fs503_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1460_out(.d0(h_arrdiv24_fs480_xor0[0]), .d1(a[3]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1460_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1461_out(.d0(h_arrdiv24_fs481_xor1[0]), .d1(h_arrdiv24_mux2to1437_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1461_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1462_out(.d0(h_arrdiv24_fs482_xor1[0]), .d1(h_arrdiv24_mux2to1438_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1462_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1463_out(.d0(h_arrdiv24_fs483_xor1[0]), .d1(h_arrdiv24_mux2to1439_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1463_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1464_out(.d0(h_arrdiv24_fs484_xor1[0]), .d1(h_arrdiv24_mux2to1440_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1464_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1465_out(.d0(h_arrdiv24_fs485_xor1[0]), .d1(h_arrdiv24_mux2to1441_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1465_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1466_out(.d0(h_arrdiv24_fs486_xor1[0]), .d1(h_arrdiv24_mux2to1442_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1466_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1467_out(.d0(h_arrdiv24_fs487_xor1[0]), .d1(h_arrdiv24_mux2to1443_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1467_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1468_out(.d0(h_arrdiv24_fs488_xor1[0]), .d1(h_arrdiv24_mux2to1444_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1468_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1469_out(.d0(h_arrdiv24_fs489_xor1[0]), .d1(h_arrdiv24_mux2to1445_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1469_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1470_out(.d0(h_arrdiv24_fs490_xor1[0]), .d1(h_arrdiv24_mux2to1446_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1470_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1471_out(.d0(h_arrdiv24_fs491_xor1[0]), .d1(h_arrdiv24_mux2to1447_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1471_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1472_out(.d0(h_arrdiv24_fs492_xor1[0]), .d1(h_arrdiv24_mux2to1448_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1472_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1473_out(.d0(h_arrdiv24_fs493_xor1[0]), .d1(h_arrdiv24_mux2to1449_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1473_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1474_out(.d0(h_arrdiv24_fs494_xor1[0]), .d1(h_arrdiv24_mux2to1450_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1474_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1475_out(.d0(h_arrdiv24_fs495_xor1[0]), .d1(h_arrdiv24_mux2to1451_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1475_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1476_out(.d0(h_arrdiv24_fs496_xor1[0]), .d1(h_arrdiv24_mux2to1452_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1476_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1477_out(.d0(h_arrdiv24_fs497_xor1[0]), .d1(h_arrdiv24_mux2to1453_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1477_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1478_out(.d0(h_arrdiv24_fs498_xor1[0]), .d1(h_arrdiv24_mux2to1454_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1478_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1479_out(.d0(h_arrdiv24_fs499_xor1[0]), .d1(h_arrdiv24_mux2to1455_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1479_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1480_out(.d0(h_arrdiv24_fs500_xor1[0]), .d1(h_arrdiv24_mux2to1456_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1480_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1481_out(.d0(h_arrdiv24_fs501_xor1[0]), .d1(h_arrdiv24_mux2to1457_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1481_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1482_out(.d0(h_arrdiv24_fs502_xor1[0]), .d1(h_arrdiv24_mux2to1458_xor0[0]), .sel(h_arrdiv24_fs503_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1482_xor0));
  not_gate not_gate_h_arrdiv24_not20(.a(h_arrdiv24_fs503_or0[0]), .out(h_arrdiv24_not20));
  fs fs_h_arrdiv24_fs504_out(.a(a[2]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs504_xor0), .fs_or0(h_arrdiv24_fs504_and0));
  fs fs_h_arrdiv24_fs505_out(.a(h_arrdiv24_mux2to1460_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs504_and0[0]), .fs_xor1(h_arrdiv24_fs505_xor1), .fs_or0(h_arrdiv24_fs505_or0));
  fs fs_h_arrdiv24_fs506_out(.a(h_arrdiv24_mux2to1461_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs505_or0[0]), .fs_xor1(h_arrdiv24_fs506_xor1), .fs_or0(h_arrdiv24_fs506_or0));
  fs fs_h_arrdiv24_fs507_out(.a(h_arrdiv24_mux2to1462_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs506_or0[0]), .fs_xor1(h_arrdiv24_fs507_xor1), .fs_or0(h_arrdiv24_fs507_or0));
  fs fs_h_arrdiv24_fs508_out(.a(h_arrdiv24_mux2to1463_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs507_or0[0]), .fs_xor1(h_arrdiv24_fs508_xor1), .fs_or0(h_arrdiv24_fs508_or0));
  fs fs_h_arrdiv24_fs509_out(.a(h_arrdiv24_mux2to1464_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs508_or0[0]), .fs_xor1(h_arrdiv24_fs509_xor1), .fs_or0(h_arrdiv24_fs509_or0));
  fs fs_h_arrdiv24_fs510_out(.a(h_arrdiv24_mux2to1465_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs509_or0[0]), .fs_xor1(h_arrdiv24_fs510_xor1), .fs_or0(h_arrdiv24_fs510_or0));
  fs fs_h_arrdiv24_fs511_out(.a(h_arrdiv24_mux2to1466_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs510_or0[0]), .fs_xor1(h_arrdiv24_fs511_xor1), .fs_or0(h_arrdiv24_fs511_or0));
  fs fs_h_arrdiv24_fs512_out(.a(h_arrdiv24_mux2to1467_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs511_or0[0]), .fs_xor1(h_arrdiv24_fs512_xor1), .fs_or0(h_arrdiv24_fs512_or0));
  fs fs_h_arrdiv24_fs513_out(.a(h_arrdiv24_mux2to1468_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs512_or0[0]), .fs_xor1(h_arrdiv24_fs513_xor1), .fs_or0(h_arrdiv24_fs513_or0));
  fs fs_h_arrdiv24_fs514_out(.a(h_arrdiv24_mux2to1469_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs513_or0[0]), .fs_xor1(h_arrdiv24_fs514_xor1), .fs_or0(h_arrdiv24_fs514_or0));
  fs fs_h_arrdiv24_fs515_out(.a(h_arrdiv24_mux2to1470_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs514_or0[0]), .fs_xor1(h_arrdiv24_fs515_xor1), .fs_or0(h_arrdiv24_fs515_or0));
  fs fs_h_arrdiv24_fs516_out(.a(h_arrdiv24_mux2to1471_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs515_or0[0]), .fs_xor1(h_arrdiv24_fs516_xor1), .fs_or0(h_arrdiv24_fs516_or0));
  fs fs_h_arrdiv24_fs517_out(.a(h_arrdiv24_mux2to1472_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs516_or0[0]), .fs_xor1(h_arrdiv24_fs517_xor1), .fs_or0(h_arrdiv24_fs517_or0));
  fs fs_h_arrdiv24_fs518_out(.a(h_arrdiv24_mux2to1473_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs517_or0[0]), .fs_xor1(h_arrdiv24_fs518_xor1), .fs_or0(h_arrdiv24_fs518_or0));
  fs fs_h_arrdiv24_fs519_out(.a(h_arrdiv24_mux2to1474_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs518_or0[0]), .fs_xor1(h_arrdiv24_fs519_xor1), .fs_or0(h_arrdiv24_fs519_or0));
  fs fs_h_arrdiv24_fs520_out(.a(h_arrdiv24_mux2to1475_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs519_or0[0]), .fs_xor1(h_arrdiv24_fs520_xor1), .fs_or0(h_arrdiv24_fs520_or0));
  fs fs_h_arrdiv24_fs521_out(.a(h_arrdiv24_mux2to1476_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs520_or0[0]), .fs_xor1(h_arrdiv24_fs521_xor1), .fs_or0(h_arrdiv24_fs521_or0));
  fs fs_h_arrdiv24_fs522_out(.a(h_arrdiv24_mux2to1477_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs521_or0[0]), .fs_xor1(h_arrdiv24_fs522_xor1), .fs_or0(h_arrdiv24_fs522_or0));
  fs fs_h_arrdiv24_fs523_out(.a(h_arrdiv24_mux2to1478_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs522_or0[0]), .fs_xor1(h_arrdiv24_fs523_xor1), .fs_or0(h_arrdiv24_fs523_or0));
  fs fs_h_arrdiv24_fs524_out(.a(h_arrdiv24_mux2to1479_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs523_or0[0]), .fs_xor1(h_arrdiv24_fs524_xor1), .fs_or0(h_arrdiv24_fs524_or0));
  fs fs_h_arrdiv24_fs525_out(.a(h_arrdiv24_mux2to1480_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs524_or0[0]), .fs_xor1(h_arrdiv24_fs525_xor1), .fs_or0(h_arrdiv24_fs525_or0));
  fs fs_h_arrdiv24_fs526_out(.a(h_arrdiv24_mux2to1481_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs525_or0[0]), .fs_xor1(h_arrdiv24_fs526_xor1), .fs_or0(h_arrdiv24_fs526_or0));
  fs fs_h_arrdiv24_fs527_out(.a(h_arrdiv24_mux2to1482_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs526_or0[0]), .fs_xor1(h_arrdiv24_fs527_xor1), .fs_or0(h_arrdiv24_fs527_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1483_out(.d0(h_arrdiv24_fs504_xor0[0]), .d1(a[2]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1483_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1484_out(.d0(h_arrdiv24_fs505_xor1[0]), .d1(h_arrdiv24_mux2to1460_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1484_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1485_out(.d0(h_arrdiv24_fs506_xor1[0]), .d1(h_arrdiv24_mux2to1461_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1485_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1486_out(.d0(h_arrdiv24_fs507_xor1[0]), .d1(h_arrdiv24_mux2to1462_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1486_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1487_out(.d0(h_arrdiv24_fs508_xor1[0]), .d1(h_arrdiv24_mux2to1463_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1487_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1488_out(.d0(h_arrdiv24_fs509_xor1[0]), .d1(h_arrdiv24_mux2to1464_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1488_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1489_out(.d0(h_arrdiv24_fs510_xor1[0]), .d1(h_arrdiv24_mux2to1465_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1489_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1490_out(.d0(h_arrdiv24_fs511_xor1[0]), .d1(h_arrdiv24_mux2to1466_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1490_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1491_out(.d0(h_arrdiv24_fs512_xor1[0]), .d1(h_arrdiv24_mux2to1467_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1491_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1492_out(.d0(h_arrdiv24_fs513_xor1[0]), .d1(h_arrdiv24_mux2to1468_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1492_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1493_out(.d0(h_arrdiv24_fs514_xor1[0]), .d1(h_arrdiv24_mux2to1469_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1493_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1494_out(.d0(h_arrdiv24_fs515_xor1[0]), .d1(h_arrdiv24_mux2to1470_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1494_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1495_out(.d0(h_arrdiv24_fs516_xor1[0]), .d1(h_arrdiv24_mux2to1471_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1495_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1496_out(.d0(h_arrdiv24_fs517_xor1[0]), .d1(h_arrdiv24_mux2to1472_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1496_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1497_out(.d0(h_arrdiv24_fs518_xor1[0]), .d1(h_arrdiv24_mux2to1473_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1497_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1498_out(.d0(h_arrdiv24_fs519_xor1[0]), .d1(h_arrdiv24_mux2to1474_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1498_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1499_out(.d0(h_arrdiv24_fs520_xor1[0]), .d1(h_arrdiv24_mux2to1475_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1499_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1500_out(.d0(h_arrdiv24_fs521_xor1[0]), .d1(h_arrdiv24_mux2to1476_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1500_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1501_out(.d0(h_arrdiv24_fs522_xor1[0]), .d1(h_arrdiv24_mux2to1477_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1501_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1502_out(.d0(h_arrdiv24_fs523_xor1[0]), .d1(h_arrdiv24_mux2to1478_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1502_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1503_out(.d0(h_arrdiv24_fs524_xor1[0]), .d1(h_arrdiv24_mux2to1479_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1503_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1504_out(.d0(h_arrdiv24_fs525_xor1[0]), .d1(h_arrdiv24_mux2to1480_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1504_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1505_out(.d0(h_arrdiv24_fs526_xor1[0]), .d1(h_arrdiv24_mux2to1481_xor0[0]), .sel(h_arrdiv24_fs527_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1505_xor0));
  not_gate not_gate_h_arrdiv24_not21(.a(h_arrdiv24_fs527_or0[0]), .out(h_arrdiv24_not21));
  fs fs_h_arrdiv24_fs528_out(.a(a[1]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs528_xor0), .fs_or0(h_arrdiv24_fs528_and0));
  fs fs_h_arrdiv24_fs529_out(.a(h_arrdiv24_mux2to1483_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs528_and0[0]), .fs_xor1(h_arrdiv24_fs529_xor1), .fs_or0(h_arrdiv24_fs529_or0));
  fs fs_h_arrdiv24_fs530_out(.a(h_arrdiv24_mux2to1484_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs529_or0[0]), .fs_xor1(h_arrdiv24_fs530_xor1), .fs_or0(h_arrdiv24_fs530_or0));
  fs fs_h_arrdiv24_fs531_out(.a(h_arrdiv24_mux2to1485_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs530_or0[0]), .fs_xor1(h_arrdiv24_fs531_xor1), .fs_or0(h_arrdiv24_fs531_or0));
  fs fs_h_arrdiv24_fs532_out(.a(h_arrdiv24_mux2to1486_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs531_or0[0]), .fs_xor1(h_arrdiv24_fs532_xor1), .fs_or0(h_arrdiv24_fs532_or0));
  fs fs_h_arrdiv24_fs533_out(.a(h_arrdiv24_mux2to1487_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs532_or0[0]), .fs_xor1(h_arrdiv24_fs533_xor1), .fs_or0(h_arrdiv24_fs533_or0));
  fs fs_h_arrdiv24_fs534_out(.a(h_arrdiv24_mux2to1488_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs533_or0[0]), .fs_xor1(h_arrdiv24_fs534_xor1), .fs_or0(h_arrdiv24_fs534_or0));
  fs fs_h_arrdiv24_fs535_out(.a(h_arrdiv24_mux2to1489_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs534_or0[0]), .fs_xor1(h_arrdiv24_fs535_xor1), .fs_or0(h_arrdiv24_fs535_or0));
  fs fs_h_arrdiv24_fs536_out(.a(h_arrdiv24_mux2to1490_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs535_or0[0]), .fs_xor1(h_arrdiv24_fs536_xor1), .fs_or0(h_arrdiv24_fs536_or0));
  fs fs_h_arrdiv24_fs537_out(.a(h_arrdiv24_mux2to1491_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs536_or0[0]), .fs_xor1(h_arrdiv24_fs537_xor1), .fs_or0(h_arrdiv24_fs537_or0));
  fs fs_h_arrdiv24_fs538_out(.a(h_arrdiv24_mux2to1492_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs537_or0[0]), .fs_xor1(h_arrdiv24_fs538_xor1), .fs_or0(h_arrdiv24_fs538_or0));
  fs fs_h_arrdiv24_fs539_out(.a(h_arrdiv24_mux2to1493_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs538_or0[0]), .fs_xor1(h_arrdiv24_fs539_xor1), .fs_or0(h_arrdiv24_fs539_or0));
  fs fs_h_arrdiv24_fs540_out(.a(h_arrdiv24_mux2to1494_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs539_or0[0]), .fs_xor1(h_arrdiv24_fs540_xor1), .fs_or0(h_arrdiv24_fs540_or0));
  fs fs_h_arrdiv24_fs541_out(.a(h_arrdiv24_mux2to1495_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs540_or0[0]), .fs_xor1(h_arrdiv24_fs541_xor1), .fs_or0(h_arrdiv24_fs541_or0));
  fs fs_h_arrdiv24_fs542_out(.a(h_arrdiv24_mux2to1496_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs541_or0[0]), .fs_xor1(h_arrdiv24_fs542_xor1), .fs_or0(h_arrdiv24_fs542_or0));
  fs fs_h_arrdiv24_fs543_out(.a(h_arrdiv24_mux2to1497_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs542_or0[0]), .fs_xor1(h_arrdiv24_fs543_xor1), .fs_or0(h_arrdiv24_fs543_or0));
  fs fs_h_arrdiv24_fs544_out(.a(h_arrdiv24_mux2to1498_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs543_or0[0]), .fs_xor1(h_arrdiv24_fs544_xor1), .fs_or0(h_arrdiv24_fs544_or0));
  fs fs_h_arrdiv24_fs545_out(.a(h_arrdiv24_mux2to1499_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs544_or0[0]), .fs_xor1(h_arrdiv24_fs545_xor1), .fs_or0(h_arrdiv24_fs545_or0));
  fs fs_h_arrdiv24_fs546_out(.a(h_arrdiv24_mux2to1500_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs545_or0[0]), .fs_xor1(h_arrdiv24_fs546_xor1), .fs_or0(h_arrdiv24_fs546_or0));
  fs fs_h_arrdiv24_fs547_out(.a(h_arrdiv24_mux2to1501_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs546_or0[0]), .fs_xor1(h_arrdiv24_fs547_xor1), .fs_or0(h_arrdiv24_fs547_or0));
  fs fs_h_arrdiv24_fs548_out(.a(h_arrdiv24_mux2to1502_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs547_or0[0]), .fs_xor1(h_arrdiv24_fs548_xor1), .fs_or0(h_arrdiv24_fs548_or0));
  fs fs_h_arrdiv24_fs549_out(.a(h_arrdiv24_mux2to1503_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs548_or0[0]), .fs_xor1(h_arrdiv24_fs549_xor1), .fs_or0(h_arrdiv24_fs549_or0));
  fs fs_h_arrdiv24_fs550_out(.a(h_arrdiv24_mux2to1504_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs549_or0[0]), .fs_xor1(h_arrdiv24_fs550_xor1), .fs_or0(h_arrdiv24_fs550_or0));
  fs fs_h_arrdiv24_fs551_out(.a(h_arrdiv24_mux2to1505_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs550_or0[0]), .fs_xor1(h_arrdiv24_fs551_xor1), .fs_or0(h_arrdiv24_fs551_or0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1506_out(.d0(h_arrdiv24_fs528_xor0[0]), .d1(a[1]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1506_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1507_out(.d0(h_arrdiv24_fs529_xor1[0]), .d1(h_arrdiv24_mux2to1483_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1507_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1508_out(.d0(h_arrdiv24_fs530_xor1[0]), .d1(h_arrdiv24_mux2to1484_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1508_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1509_out(.d0(h_arrdiv24_fs531_xor1[0]), .d1(h_arrdiv24_mux2to1485_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1509_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1510_out(.d0(h_arrdiv24_fs532_xor1[0]), .d1(h_arrdiv24_mux2to1486_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1510_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1511_out(.d0(h_arrdiv24_fs533_xor1[0]), .d1(h_arrdiv24_mux2to1487_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1511_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1512_out(.d0(h_arrdiv24_fs534_xor1[0]), .d1(h_arrdiv24_mux2to1488_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1512_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1513_out(.d0(h_arrdiv24_fs535_xor1[0]), .d1(h_arrdiv24_mux2to1489_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1513_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1514_out(.d0(h_arrdiv24_fs536_xor1[0]), .d1(h_arrdiv24_mux2to1490_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1514_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1515_out(.d0(h_arrdiv24_fs537_xor1[0]), .d1(h_arrdiv24_mux2to1491_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1515_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1516_out(.d0(h_arrdiv24_fs538_xor1[0]), .d1(h_arrdiv24_mux2to1492_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1516_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1517_out(.d0(h_arrdiv24_fs539_xor1[0]), .d1(h_arrdiv24_mux2to1493_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1517_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1518_out(.d0(h_arrdiv24_fs540_xor1[0]), .d1(h_arrdiv24_mux2to1494_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1518_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1519_out(.d0(h_arrdiv24_fs541_xor1[0]), .d1(h_arrdiv24_mux2to1495_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1519_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1520_out(.d0(h_arrdiv24_fs542_xor1[0]), .d1(h_arrdiv24_mux2to1496_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1520_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1521_out(.d0(h_arrdiv24_fs543_xor1[0]), .d1(h_arrdiv24_mux2to1497_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1521_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1522_out(.d0(h_arrdiv24_fs544_xor1[0]), .d1(h_arrdiv24_mux2to1498_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1522_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1523_out(.d0(h_arrdiv24_fs545_xor1[0]), .d1(h_arrdiv24_mux2to1499_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1523_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1524_out(.d0(h_arrdiv24_fs546_xor1[0]), .d1(h_arrdiv24_mux2to1500_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1524_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1525_out(.d0(h_arrdiv24_fs547_xor1[0]), .d1(h_arrdiv24_mux2to1501_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1525_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1526_out(.d0(h_arrdiv24_fs548_xor1[0]), .d1(h_arrdiv24_mux2to1502_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1526_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1527_out(.d0(h_arrdiv24_fs549_xor1[0]), .d1(h_arrdiv24_mux2to1503_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1527_xor0));
  mux2to1 mux2to1_h_arrdiv24_mux2to1528_out(.d0(h_arrdiv24_fs550_xor1[0]), .d1(h_arrdiv24_mux2to1504_xor0[0]), .sel(h_arrdiv24_fs551_or0[0]), .mux2to1_xor0(h_arrdiv24_mux2to1528_xor0));
  not_gate not_gate_h_arrdiv24_not22(.a(h_arrdiv24_fs551_or0[0]), .out(h_arrdiv24_not22));
  fs fs_h_arrdiv24_fs552_out(.a(a[0]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv24_fs552_xor0), .fs_or0(h_arrdiv24_fs552_and0));
  fs fs_h_arrdiv24_fs553_out(.a(h_arrdiv24_mux2to1506_xor0[0]), .b(b[1]), .bin(h_arrdiv24_fs552_and0[0]), .fs_xor1(h_arrdiv24_fs553_xor1), .fs_or0(h_arrdiv24_fs553_or0));
  fs fs_h_arrdiv24_fs554_out(.a(h_arrdiv24_mux2to1507_xor0[0]), .b(b[2]), .bin(h_arrdiv24_fs553_or0[0]), .fs_xor1(h_arrdiv24_fs554_xor1), .fs_or0(h_arrdiv24_fs554_or0));
  fs fs_h_arrdiv24_fs555_out(.a(h_arrdiv24_mux2to1508_xor0[0]), .b(b[3]), .bin(h_arrdiv24_fs554_or0[0]), .fs_xor1(h_arrdiv24_fs555_xor1), .fs_or0(h_arrdiv24_fs555_or0));
  fs fs_h_arrdiv24_fs556_out(.a(h_arrdiv24_mux2to1509_xor0[0]), .b(b[4]), .bin(h_arrdiv24_fs555_or0[0]), .fs_xor1(h_arrdiv24_fs556_xor1), .fs_or0(h_arrdiv24_fs556_or0));
  fs fs_h_arrdiv24_fs557_out(.a(h_arrdiv24_mux2to1510_xor0[0]), .b(b[5]), .bin(h_arrdiv24_fs556_or0[0]), .fs_xor1(h_arrdiv24_fs557_xor1), .fs_or0(h_arrdiv24_fs557_or0));
  fs fs_h_arrdiv24_fs558_out(.a(h_arrdiv24_mux2to1511_xor0[0]), .b(b[6]), .bin(h_arrdiv24_fs557_or0[0]), .fs_xor1(h_arrdiv24_fs558_xor1), .fs_or0(h_arrdiv24_fs558_or0));
  fs fs_h_arrdiv24_fs559_out(.a(h_arrdiv24_mux2to1512_xor0[0]), .b(b[7]), .bin(h_arrdiv24_fs558_or0[0]), .fs_xor1(h_arrdiv24_fs559_xor1), .fs_or0(h_arrdiv24_fs559_or0));
  fs fs_h_arrdiv24_fs560_out(.a(h_arrdiv24_mux2to1513_xor0[0]), .b(b[8]), .bin(h_arrdiv24_fs559_or0[0]), .fs_xor1(h_arrdiv24_fs560_xor1), .fs_or0(h_arrdiv24_fs560_or0));
  fs fs_h_arrdiv24_fs561_out(.a(h_arrdiv24_mux2to1514_xor0[0]), .b(b[9]), .bin(h_arrdiv24_fs560_or0[0]), .fs_xor1(h_arrdiv24_fs561_xor1), .fs_or0(h_arrdiv24_fs561_or0));
  fs fs_h_arrdiv24_fs562_out(.a(h_arrdiv24_mux2to1515_xor0[0]), .b(b[10]), .bin(h_arrdiv24_fs561_or0[0]), .fs_xor1(h_arrdiv24_fs562_xor1), .fs_or0(h_arrdiv24_fs562_or0));
  fs fs_h_arrdiv24_fs563_out(.a(h_arrdiv24_mux2to1516_xor0[0]), .b(b[11]), .bin(h_arrdiv24_fs562_or0[0]), .fs_xor1(h_arrdiv24_fs563_xor1), .fs_or0(h_arrdiv24_fs563_or0));
  fs fs_h_arrdiv24_fs564_out(.a(h_arrdiv24_mux2to1517_xor0[0]), .b(b[12]), .bin(h_arrdiv24_fs563_or0[0]), .fs_xor1(h_arrdiv24_fs564_xor1), .fs_or0(h_arrdiv24_fs564_or0));
  fs fs_h_arrdiv24_fs565_out(.a(h_arrdiv24_mux2to1518_xor0[0]), .b(b[13]), .bin(h_arrdiv24_fs564_or0[0]), .fs_xor1(h_arrdiv24_fs565_xor1), .fs_or0(h_arrdiv24_fs565_or0));
  fs fs_h_arrdiv24_fs566_out(.a(h_arrdiv24_mux2to1519_xor0[0]), .b(b[14]), .bin(h_arrdiv24_fs565_or0[0]), .fs_xor1(h_arrdiv24_fs566_xor1), .fs_or0(h_arrdiv24_fs566_or0));
  fs fs_h_arrdiv24_fs567_out(.a(h_arrdiv24_mux2to1520_xor0[0]), .b(b[15]), .bin(h_arrdiv24_fs566_or0[0]), .fs_xor1(h_arrdiv24_fs567_xor1), .fs_or0(h_arrdiv24_fs567_or0));
  fs fs_h_arrdiv24_fs568_out(.a(h_arrdiv24_mux2to1521_xor0[0]), .b(b[16]), .bin(h_arrdiv24_fs567_or0[0]), .fs_xor1(h_arrdiv24_fs568_xor1), .fs_or0(h_arrdiv24_fs568_or0));
  fs fs_h_arrdiv24_fs569_out(.a(h_arrdiv24_mux2to1522_xor0[0]), .b(b[17]), .bin(h_arrdiv24_fs568_or0[0]), .fs_xor1(h_arrdiv24_fs569_xor1), .fs_or0(h_arrdiv24_fs569_or0));
  fs fs_h_arrdiv24_fs570_out(.a(h_arrdiv24_mux2to1523_xor0[0]), .b(b[18]), .bin(h_arrdiv24_fs569_or0[0]), .fs_xor1(h_arrdiv24_fs570_xor1), .fs_or0(h_arrdiv24_fs570_or0));
  fs fs_h_arrdiv24_fs571_out(.a(h_arrdiv24_mux2to1524_xor0[0]), .b(b[19]), .bin(h_arrdiv24_fs570_or0[0]), .fs_xor1(h_arrdiv24_fs571_xor1), .fs_or0(h_arrdiv24_fs571_or0));
  fs fs_h_arrdiv24_fs572_out(.a(h_arrdiv24_mux2to1525_xor0[0]), .b(b[20]), .bin(h_arrdiv24_fs571_or0[0]), .fs_xor1(h_arrdiv24_fs572_xor1), .fs_or0(h_arrdiv24_fs572_or0));
  fs fs_h_arrdiv24_fs573_out(.a(h_arrdiv24_mux2to1526_xor0[0]), .b(b[21]), .bin(h_arrdiv24_fs572_or0[0]), .fs_xor1(h_arrdiv24_fs573_xor1), .fs_or0(h_arrdiv24_fs573_or0));
  fs fs_h_arrdiv24_fs574_out(.a(h_arrdiv24_mux2to1527_xor0[0]), .b(b[22]), .bin(h_arrdiv24_fs573_or0[0]), .fs_xor1(h_arrdiv24_fs574_xor1), .fs_or0(h_arrdiv24_fs574_or0));
  fs fs_h_arrdiv24_fs575_out(.a(h_arrdiv24_mux2to1528_xor0[0]), .b(b[23]), .bin(h_arrdiv24_fs574_or0[0]), .fs_xor1(h_arrdiv24_fs575_xor1), .fs_or0(h_arrdiv24_fs575_or0));
  not_gate not_gate_h_arrdiv24_not23(.a(h_arrdiv24_fs575_or0[0]), .out(h_arrdiv24_not23));

  assign h_arrdiv24_out[0] = h_arrdiv24_not23[0];
  assign h_arrdiv24_out[1] = h_arrdiv24_not22[0];
  assign h_arrdiv24_out[2] = h_arrdiv24_not21[0];
  assign h_arrdiv24_out[3] = h_arrdiv24_not20[0];
  assign h_arrdiv24_out[4] = h_arrdiv24_not19[0];
  assign h_arrdiv24_out[5] = h_arrdiv24_not18[0];
  assign h_arrdiv24_out[6] = h_arrdiv24_not17[0];
  assign h_arrdiv24_out[7] = h_arrdiv24_not16[0];
  assign h_arrdiv24_out[8] = h_arrdiv24_not15[0];
  assign h_arrdiv24_out[9] = h_arrdiv24_not14[0];
  assign h_arrdiv24_out[10] = h_arrdiv24_not13[0];
  assign h_arrdiv24_out[11] = h_arrdiv24_not12[0];
  assign h_arrdiv24_out[12] = h_arrdiv24_not11[0];
  assign h_arrdiv24_out[13] = h_arrdiv24_not10[0];
  assign h_arrdiv24_out[14] = h_arrdiv24_not9[0];
  assign h_arrdiv24_out[15] = h_arrdiv24_not8[0];
  assign h_arrdiv24_out[16] = h_arrdiv24_not7[0];
  assign h_arrdiv24_out[17] = h_arrdiv24_not6[0];
  assign h_arrdiv24_out[18] = h_arrdiv24_not5[0];
  assign h_arrdiv24_out[19] = h_arrdiv24_not4[0];
  assign h_arrdiv24_out[20] = h_arrdiv24_not3[0];
  assign h_arrdiv24_out[21] = h_arrdiv24_not2[0];
  assign h_arrdiv24_out[22] = h_arrdiv24_not1[0];
  assign h_arrdiv24_out[23] = h_arrdiv24_not0[0];
endmodule