module f_u_arr_mul2(input [1:0] a, input [1:0] b, output [3:0] out);
  wire a_0;
  wire a_1;
  wire b_0;
  wire b_1;
  wire f_u_arr_mul2_and_0_0_a_0;
  wire f_u_arr_mul2_and_0_0_b_0;
  wire f_u_arr_mul2_and_0_0_y0;
  wire f_u_arr_mul2_and_1_0_a_1;
  wire f_u_arr_mul2_and_1_0_b_0;
  wire f_u_arr_mul2_and_1_0_y0;
  wire f_u_arr_mul2_and_0_1_a_0;
  wire f_u_arr_mul2_and_0_1_b_1;
  wire f_u_arr_mul2_and_0_1_y0;
  wire f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_0_1_y0;
  wire f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_1_0_y0;
  wire f_u_arr_mul2_ha_0_1_y0;
  wire f_u_arr_mul2_ha_0_1_y1;
  wire f_u_arr_mul2_and_1_1_a_1;
  wire f_u_arr_mul2_and_1_1_b_1;
  wire f_u_arr_mul2_and_1_1_y0;
  wire f_u_arr_mul2_ha_1_1_f_u_arr_mul2_and_1_1_y0;
  wire f_u_arr_mul2_ha_1_1_f_u_arr_mul2_ha_0_1_y1;
  wire f_u_arr_mul2_ha_1_1_y0;
  wire f_u_arr_mul2_ha_1_1_y1;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign f_u_arr_mul2_and_0_0_a_0 = a_0;
  assign f_u_arr_mul2_and_0_0_b_0 = b_0;
  assign f_u_arr_mul2_and_0_0_y0 = f_u_arr_mul2_and_0_0_a_0 & f_u_arr_mul2_and_0_0_b_0;
  assign f_u_arr_mul2_and_1_0_a_1 = a_1;
  assign f_u_arr_mul2_and_1_0_b_0 = b_0;
  assign f_u_arr_mul2_and_1_0_y0 = f_u_arr_mul2_and_1_0_a_1 & f_u_arr_mul2_and_1_0_b_0;
  assign f_u_arr_mul2_and_0_1_a_0 = a_0;
  assign f_u_arr_mul2_and_0_1_b_1 = b_1;
  assign f_u_arr_mul2_and_0_1_y0 = f_u_arr_mul2_and_0_1_a_0 & f_u_arr_mul2_and_0_1_b_1;
  assign f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_0_1_y0 = f_u_arr_mul2_and_0_1_y0;
  assign f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_1_0_y0 = f_u_arr_mul2_and_1_0_y0;
  assign f_u_arr_mul2_ha_0_1_y0 = f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_0_1_y0 ^ f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_1_0_y0;
  assign f_u_arr_mul2_ha_0_1_y1 = f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_0_1_y0 & f_u_arr_mul2_ha_0_1_f_u_arr_mul2_and_1_0_y0;
  assign f_u_arr_mul2_and_1_1_a_1 = a_1;
  assign f_u_arr_mul2_and_1_1_b_1 = b_1;
  assign f_u_arr_mul2_and_1_1_y0 = f_u_arr_mul2_and_1_1_a_1 & f_u_arr_mul2_and_1_1_b_1;
  assign f_u_arr_mul2_ha_1_1_f_u_arr_mul2_and_1_1_y0 = f_u_arr_mul2_and_1_1_y0;
  assign f_u_arr_mul2_ha_1_1_f_u_arr_mul2_ha_0_1_y1 = f_u_arr_mul2_ha_0_1_y1;
  assign f_u_arr_mul2_ha_1_1_y0 = f_u_arr_mul2_ha_1_1_f_u_arr_mul2_and_1_1_y0 ^ f_u_arr_mul2_ha_1_1_f_u_arr_mul2_ha_0_1_y1;
  assign f_u_arr_mul2_ha_1_1_y1 = f_u_arr_mul2_ha_1_1_f_u_arr_mul2_and_1_1_y0 & f_u_arr_mul2_ha_1_1_f_u_arr_mul2_ha_0_1_y1;

  assign out[0] = f_u_arr_mul2_and_0_0_y0;
  assign out[1] = f_u_arr_mul2_ha_0_1_y0;
  assign out[2] = f_u_arr_mul2_ha_1_1_y0;
  assign out[3] = f_u_arr_mul2_ha_1_1_y1;
endmodule