module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] pg_fa_xor0, output [0:0] pg_fa_and0, output [0:0] pg_fa_xor1);
  xor_gate xor_gate_pg_fa_xor0(.a(a[0]), .b(b[0]), .out(pg_fa_xor0));
  and_gate and_gate_pg_fa_and0(.a(a[0]), .b(b[0]), .out(pg_fa_and0));
  xor_gate xor_gate_pg_fa_xor1(.a(pg_fa_xor0[0]), .b(cin[0]), .out(pg_fa_xor1));
endmodule

module u_pg_rca24(input [23:0] a, input [23:0] b, output [24:0] u_pg_rca24_out);
  wire [0:0] u_pg_rca24_pg_fa0_xor0;
  wire [0:0] u_pg_rca24_pg_fa0_and0;
  wire [0:0] u_pg_rca24_pg_fa1_xor0;
  wire [0:0] u_pg_rca24_pg_fa1_and0;
  wire [0:0] u_pg_rca24_pg_fa1_xor1;
  wire [0:0] u_pg_rca24_and1;
  wire [0:0] u_pg_rca24_or1;
  wire [0:0] u_pg_rca24_pg_fa2_xor0;
  wire [0:0] u_pg_rca24_pg_fa2_and0;
  wire [0:0] u_pg_rca24_pg_fa2_xor1;
  wire [0:0] u_pg_rca24_and2;
  wire [0:0] u_pg_rca24_or2;
  wire [0:0] u_pg_rca24_pg_fa3_xor0;
  wire [0:0] u_pg_rca24_pg_fa3_and0;
  wire [0:0] u_pg_rca24_pg_fa3_xor1;
  wire [0:0] u_pg_rca24_and3;
  wire [0:0] u_pg_rca24_or3;
  wire [0:0] u_pg_rca24_pg_fa4_xor0;
  wire [0:0] u_pg_rca24_pg_fa4_and0;
  wire [0:0] u_pg_rca24_pg_fa4_xor1;
  wire [0:0] u_pg_rca24_and4;
  wire [0:0] u_pg_rca24_or4;
  wire [0:0] u_pg_rca24_pg_fa5_xor0;
  wire [0:0] u_pg_rca24_pg_fa5_and0;
  wire [0:0] u_pg_rca24_pg_fa5_xor1;
  wire [0:0] u_pg_rca24_and5;
  wire [0:0] u_pg_rca24_or5;
  wire [0:0] u_pg_rca24_pg_fa6_xor0;
  wire [0:0] u_pg_rca24_pg_fa6_and0;
  wire [0:0] u_pg_rca24_pg_fa6_xor1;
  wire [0:0] u_pg_rca24_and6;
  wire [0:0] u_pg_rca24_or6;
  wire [0:0] u_pg_rca24_pg_fa7_xor0;
  wire [0:0] u_pg_rca24_pg_fa7_and0;
  wire [0:0] u_pg_rca24_pg_fa7_xor1;
  wire [0:0] u_pg_rca24_and7;
  wire [0:0] u_pg_rca24_or7;
  wire [0:0] u_pg_rca24_pg_fa8_xor0;
  wire [0:0] u_pg_rca24_pg_fa8_and0;
  wire [0:0] u_pg_rca24_pg_fa8_xor1;
  wire [0:0] u_pg_rca24_and8;
  wire [0:0] u_pg_rca24_or8;
  wire [0:0] u_pg_rca24_pg_fa9_xor0;
  wire [0:0] u_pg_rca24_pg_fa9_and0;
  wire [0:0] u_pg_rca24_pg_fa9_xor1;
  wire [0:0] u_pg_rca24_and9;
  wire [0:0] u_pg_rca24_or9;
  wire [0:0] u_pg_rca24_pg_fa10_xor0;
  wire [0:0] u_pg_rca24_pg_fa10_and0;
  wire [0:0] u_pg_rca24_pg_fa10_xor1;
  wire [0:0] u_pg_rca24_and10;
  wire [0:0] u_pg_rca24_or10;
  wire [0:0] u_pg_rca24_pg_fa11_xor0;
  wire [0:0] u_pg_rca24_pg_fa11_and0;
  wire [0:0] u_pg_rca24_pg_fa11_xor1;
  wire [0:0] u_pg_rca24_and11;
  wire [0:0] u_pg_rca24_or11;
  wire [0:0] u_pg_rca24_pg_fa12_xor0;
  wire [0:0] u_pg_rca24_pg_fa12_and0;
  wire [0:0] u_pg_rca24_pg_fa12_xor1;
  wire [0:0] u_pg_rca24_and12;
  wire [0:0] u_pg_rca24_or12;
  wire [0:0] u_pg_rca24_pg_fa13_xor0;
  wire [0:0] u_pg_rca24_pg_fa13_and0;
  wire [0:0] u_pg_rca24_pg_fa13_xor1;
  wire [0:0] u_pg_rca24_and13;
  wire [0:0] u_pg_rca24_or13;
  wire [0:0] u_pg_rca24_pg_fa14_xor0;
  wire [0:0] u_pg_rca24_pg_fa14_and0;
  wire [0:0] u_pg_rca24_pg_fa14_xor1;
  wire [0:0] u_pg_rca24_and14;
  wire [0:0] u_pg_rca24_or14;
  wire [0:0] u_pg_rca24_pg_fa15_xor0;
  wire [0:0] u_pg_rca24_pg_fa15_and0;
  wire [0:0] u_pg_rca24_pg_fa15_xor1;
  wire [0:0] u_pg_rca24_and15;
  wire [0:0] u_pg_rca24_or15;
  wire [0:0] u_pg_rca24_pg_fa16_xor0;
  wire [0:0] u_pg_rca24_pg_fa16_and0;
  wire [0:0] u_pg_rca24_pg_fa16_xor1;
  wire [0:0] u_pg_rca24_and16;
  wire [0:0] u_pg_rca24_or16;
  wire [0:0] u_pg_rca24_pg_fa17_xor0;
  wire [0:0] u_pg_rca24_pg_fa17_and0;
  wire [0:0] u_pg_rca24_pg_fa17_xor1;
  wire [0:0] u_pg_rca24_and17;
  wire [0:0] u_pg_rca24_or17;
  wire [0:0] u_pg_rca24_pg_fa18_xor0;
  wire [0:0] u_pg_rca24_pg_fa18_and0;
  wire [0:0] u_pg_rca24_pg_fa18_xor1;
  wire [0:0] u_pg_rca24_and18;
  wire [0:0] u_pg_rca24_or18;
  wire [0:0] u_pg_rca24_pg_fa19_xor0;
  wire [0:0] u_pg_rca24_pg_fa19_and0;
  wire [0:0] u_pg_rca24_pg_fa19_xor1;
  wire [0:0] u_pg_rca24_and19;
  wire [0:0] u_pg_rca24_or19;
  wire [0:0] u_pg_rca24_pg_fa20_xor0;
  wire [0:0] u_pg_rca24_pg_fa20_and0;
  wire [0:0] u_pg_rca24_pg_fa20_xor1;
  wire [0:0] u_pg_rca24_and20;
  wire [0:0] u_pg_rca24_or20;
  wire [0:0] u_pg_rca24_pg_fa21_xor0;
  wire [0:0] u_pg_rca24_pg_fa21_and0;
  wire [0:0] u_pg_rca24_pg_fa21_xor1;
  wire [0:0] u_pg_rca24_and21;
  wire [0:0] u_pg_rca24_or21;
  wire [0:0] u_pg_rca24_pg_fa22_xor0;
  wire [0:0] u_pg_rca24_pg_fa22_and0;
  wire [0:0] u_pg_rca24_pg_fa22_xor1;
  wire [0:0] u_pg_rca24_and22;
  wire [0:0] u_pg_rca24_or22;
  wire [0:0] u_pg_rca24_pg_fa23_xor0;
  wire [0:0] u_pg_rca24_pg_fa23_and0;
  wire [0:0] u_pg_rca24_pg_fa23_xor1;
  wire [0:0] u_pg_rca24_and23;
  wire [0:0] u_pg_rca24_or23;

  pg_fa pg_fa_u_pg_rca24_pg_fa0_out(.a(a[0]), .b(b[0]), .cin(1'b0), .pg_fa_xor0(u_pg_rca24_pg_fa0_xor0), .pg_fa_and0(u_pg_rca24_pg_fa0_and0), .pg_fa_xor1());
  pg_fa pg_fa_u_pg_rca24_pg_fa1_out(.a(a[1]), .b(b[1]), .cin(u_pg_rca24_pg_fa0_and0[0]), .pg_fa_xor0(u_pg_rca24_pg_fa1_xor0), .pg_fa_and0(u_pg_rca24_pg_fa1_and0), .pg_fa_xor1(u_pg_rca24_pg_fa1_xor1));
  and_gate and_gate_u_pg_rca24_and1(.a(u_pg_rca24_pg_fa0_and0[0]), .b(u_pg_rca24_pg_fa1_xor0[0]), .out(u_pg_rca24_and1));
  or_gate or_gate_u_pg_rca24_or1(.a(u_pg_rca24_and1[0]), .b(u_pg_rca24_pg_fa1_and0[0]), .out(u_pg_rca24_or1));
  pg_fa pg_fa_u_pg_rca24_pg_fa2_out(.a(a[2]), .b(b[2]), .cin(u_pg_rca24_or1[0]), .pg_fa_xor0(u_pg_rca24_pg_fa2_xor0), .pg_fa_and0(u_pg_rca24_pg_fa2_and0), .pg_fa_xor1(u_pg_rca24_pg_fa2_xor1));
  and_gate and_gate_u_pg_rca24_and2(.a(u_pg_rca24_or1[0]), .b(u_pg_rca24_pg_fa2_xor0[0]), .out(u_pg_rca24_and2));
  or_gate or_gate_u_pg_rca24_or2(.a(u_pg_rca24_and2[0]), .b(u_pg_rca24_pg_fa2_and0[0]), .out(u_pg_rca24_or2));
  pg_fa pg_fa_u_pg_rca24_pg_fa3_out(.a(a[3]), .b(b[3]), .cin(u_pg_rca24_or2[0]), .pg_fa_xor0(u_pg_rca24_pg_fa3_xor0), .pg_fa_and0(u_pg_rca24_pg_fa3_and0), .pg_fa_xor1(u_pg_rca24_pg_fa3_xor1));
  and_gate and_gate_u_pg_rca24_and3(.a(u_pg_rca24_or2[0]), .b(u_pg_rca24_pg_fa3_xor0[0]), .out(u_pg_rca24_and3));
  or_gate or_gate_u_pg_rca24_or3(.a(u_pg_rca24_and3[0]), .b(u_pg_rca24_pg_fa3_and0[0]), .out(u_pg_rca24_or3));
  pg_fa pg_fa_u_pg_rca24_pg_fa4_out(.a(a[4]), .b(b[4]), .cin(u_pg_rca24_or3[0]), .pg_fa_xor0(u_pg_rca24_pg_fa4_xor0), .pg_fa_and0(u_pg_rca24_pg_fa4_and0), .pg_fa_xor1(u_pg_rca24_pg_fa4_xor1));
  and_gate and_gate_u_pg_rca24_and4(.a(u_pg_rca24_or3[0]), .b(u_pg_rca24_pg_fa4_xor0[0]), .out(u_pg_rca24_and4));
  or_gate or_gate_u_pg_rca24_or4(.a(u_pg_rca24_and4[0]), .b(u_pg_rca24_pg_fa4_and0[0]), .out(u_pg_rca24_or4));
  pg_fa pg_fa_u_pg_rca24_pg_fa5_out(.a(a[5]), .b(b[5]), .cin(u_pg_rca24_or4[0]), .pg_fa_xor0(u_pg_rca24_pg_fa5_xor0), .pg_fa_and0(u_pg_rca24_pg_fa5_and0), .pg_fa_xor1(u_pg_rca24_pg_fa5_xor1));
  and_gate and_gate_u_pg_rca24_and5(.a(u_pg_rca24_or4[0]), .b(u_pg_rca24_pg_fa5_xor0[0]), .out(u_pg_rca24_and5));
  or_gate or_gate_u_pg_rca24_or5(.a(u_pg_rca24_and5[0]), .b(u_pg_rca24_pg_fa5_and0[0]), .out(u_pg_rca24_or5));
  pg_fa pg_fa_u_pg_rca24_pg_fa6_out(.a(a[6]), .b(b[6]), .cin(u_pg_rca24_or5[0]), .pg_fa_xor0(u_pg_rca24_pg_fa6_xor0), .pg_fa_and0(u_pg_rca24_pg_fa6_and0), .pg_fa_xor1(u_pg_rca24_pg_fa6_xor1));
  and_gate and_gate_u_pg_rca24_and6(.a(u_pg_rca24_or5[0]), .b(u_pg_rca24_pg_fa6_xor0[0]), .out(u_pg_rca24_and6));
  or_gate or_gate_u_pg_rca24_or6(.a(u_pg_rca24_and6[0]), .b(u_pg_rca24_pg_fa6_and0[0]), .out(u_pg_rca24_or6));
  pg_fa pg_fa_u_pg_rca24_pg_fa7_out(.a(a[7]), .b(b[7]), .cin(u_pg_rca24_or6[0]), .pg_fa_xor0(u_pg_rca24_pg_fa7_xor0), .pg_fa_and0(u_pg_rca24_pg_fa7_and0), .pg_fa_xor1(u_pg_rca24_pg_fa7_xor1));
  and_gate and_gate_u_pg_rca24_and7(.a(u_pg_rca24_or6[0]), .b(u_pg_rca24_pg_fa7_xor0[0]), .out(u_pg_rca24_and7));
  or_gate or_gate_u_pg_rca24_or7(.a(u_pg_rca24_and7[0]), .b(u_pg_rca24_pg_fa7_and0[0]), .out(u_pg_rca24_or7));
  pg_fa pg_fa_u_pg_rca24_pg_fa8_out(.a(a[8]), .b(b[8]), .cin(u_pg_rca24_or7[0]), .pg_fa_xor0(u_pg_rca24_pg_fa8_xor0), .pg_fa_and0(u_pg_rca24_pg_fa8_and0), .pg_fa_xor1(u_pg_rca24_pg_fa8_xor1));
  and_gate and_gate_u_pg_rca24_and8(.a(u_pg_rca24_or7[0]), .b(u_pg_rca24_pg_fa8_xor0[0]), .out(u_pg_rca24_and8));
  or_gate or_gate_u_pg_rca24_or8(.a(u_pg_rca24_and8[0]), .b(u_pg_rca24_pg_fa8_and0[0]), .out(u_pg_rca24_or8));
  pg_fa pg_fa_u_pg_rca24_pg_fa9_out(.a(a[9]), .b(b[9]), .cin(u_pg_rca24_or8[0]), .pg_fa_xor0(u_pg_rca24_pg_fa9_xor0), .pg_fa_and0(u_pg_rca24_pg_fa9_and0), .pg_fa_xor1(u_pg_rca24_pg_fa9_xor1));
  and_gate and_gate_u_pg_rca24_and9(.a(u_pg_rca24_or8[0]), .b(u_pg_rca24_pg_fa9_xor0[0]), .out(u_pg_rca24_and9));
  or_gate or_gate_u_pg_rca24_or9(.a(u_pg_rca24_and9[0]), .b(u_pg_rca24_pg_fa9_and0[0]), .out(u_pg_rca24_or9));
  pg_fa pg_fa_u_pg_rca24_pg_fa10_out(.a(a[10]), .b(b[10]), .cin(u_pg_rca24_or9[0]), .pg_fa_xor0(u_pg_rca24_pg_fa10_xor0), .pg_fa_and0(u_pg_rca24_pg_fa10_and0), .pg_fa_xor1(u_pg_rca24_pg_fa10_xor1));
  and_gate and_gate_u_pg_rca24_and10(.a(u_pg_rca24_or9[0]), .b(u_pg_rca24_pg_fa10_xor0[0]), .out(u_pg_rca24_and10));
  or_gate or_gate_u_pg_rca24_or10(.a(u_pg_rca24_and10[0]), .b(u_pg_rca24_pg_fa10_and0[0]), .out(u_pg_rca24_or10));
  pg_fa pg_fa_u_pg_rca24_pg_fa11_out(.a(a[11]), .b(b[11]), .cin(u_pg_rca24_or10[0]), .pg_fa_xor0(u_pg_rca24_pg_fa11_xor0), .pg_fa_and0(u_pg_rca24_pg_fa11_and0), .pg_fa_xor1(u_pg_rca24_pg_fa11_xor1));
  and_gate and_gate_u_pg_rca24_and11(.a(u_pg_rca24_or10[0]), .b(u_pg_rca24_pg_fa11_xor0[0]), .out(u_pg_rca24_and11));
  or_gate or_gate_u_pg_rca24_or11(.a(u_pg_rca24_and11[0]), .b(u_pg_rca24_pg_fa11_and0[0]), .out(u_pg_rca24_or11));
  pg_fa pg_fa_u_pg_rca24_pg_fa12_out(.a(a[12]), .b(b[12]), .cin(u_pg_rca24_or11[0]), .pg_fa_xor0(u_pg_rca24_pg_fa12_xor0), .pg_fa_and0(u_pg_rca24_pg_fa12_and0), .pg_fa_xor1(u_pg_rca24_pg_fa12_xor1));
  and_gate and_gate_u_pg_rca24_and12(.a(u_pg_rca24_or11[0]), .b(u_pg_rca24_pg_fa12_xor0[0]), .out(u_pg_rca24_and12));
  or_gate or_gate_u_pg_rca24_or12(.a(u_pg_rca24_and12[0]), .b(u_pg_rca24_pg_fa12_and0[0]), .out(u_pg_rca24_or12));
  pg_fa pg_fa_u_pg_rca24_pg_fa13_out(.a(a[13]), .b(b[13]), .cin(u_pg_rca24_or12[0]), .pg_fa_xor0(u_pg_rca24_pg_fa13_xor0), .pg_fa_and0(u_pg_rca24_pg_fa13_and0), .pg_fa_xor1(u_pg_rca24_pg_fa13_xor1));
  and_gate and_gate_u_pg_rca24_and13(.a(u_pg_rca24_or12[0]), .b(u_pg_rca24_pg_fa13_xor0[0]), .out(u_pg_rca24_and13));
  or_gate or_gate_u_pg_rca24_or13(.a(u_pg_rca24_and13[0]), .b(u_pg_rca24_pg_fa13_and0[0]), .out(u_pg_rca24_or13));
  pg_fa pg_fa_u_pg_rca24_pg_fa14_out(.a(a[14]), .b(b[14]), .cin(u_pg_rca24_or13[0]), .pg_fa_xor0(u_pg_rca24_pg_fa14_xor0), .pg_fa_and0(u_pg_rca24_pg_fa14_and0), .pg_fa_xor1(u_pg_rca24_pg_fa14_xor1));
  and_gate and_gate_u_pg_rca24_and14(.a(u_pg_rca24_or13[0]), .b(u_pg_rca24_pg_fa14_xor0[0]), .out(u_pg_rca24_and14));
  or_gate or_gate_u_pg_rca24_or14(.a(u_pg_rca24_and14[0]), .b(u_pg_rca24_pg_fa14_and0[0]), .out(u_pg_rca24_or14));
  pg_fa pg_fa_u_pg_rca24_pg_fa15_out(.a(a[15]), .b(b[15]), .cin(u_pg_rca24_or14[0]), .pg_fa_xor0(u_pg_rca24_pg_fa15_xor0), .pg_fa_and0(u_pg_rca24_pg_fa15_and0), .pg_fa_xor1(u_pg_rca24_pg_fa15_xor1));
  and_gate and_gate_u_pg_rca24_and15(.a(u_pg_rca24_or14[0]), .b(u_pg_rca24_pg_fa15_xor0[0]), .out(u_pg_rca24_and15));
  or_gate or_gate_u_pg_rca24_or15(.a(u_pg_rca24_and15[0]), .b(u_pg_rca24_pg_fa15_and0[0]), .out(u_pg_rca24_or15));
  pg_fa pg_fa_u_pg_rca24_pg_fa16_out(.a(a[16]), .b(b[16]), .cin(u_pg_rca24_or15[0]), .pg_fa_xor0(u_pg_rca24_pg_fa16_xor0), .pg_fa_and0(u_pg_rca24_pg_fa16_and0), .pg_fa_xor1(u_pg_rca24_pg_fa16_xor1));
  and_gate and_gate_u_pg_rca24_and16(.a(u_pg_rca24_or15[0]), .b(u_pg_rca24_pg_fa16_xor0[0]), .out(u_pg_rca24_and16));
  or_gate or_gate_u_pg_rca24_or16(.a(u_pg_rca24_and16[0]), .b(u_pg_rca24_pg_fa16_and0[0]), .out(u_pg_rca24_or16));
  pg_fa pg_fa_u_pg_rca24_pg_fa17_out(.a(a[17]), .b(b[17]), .cin(u_pg_rca24_or16[0]), .pg_fa_xor0(u_pg_rca24_pg_fa17_xor0), .pg_fa_and0(u_pg_rca24_pg_fa17_and0), .pg_fa_xor1(u_pg_rca24_pg_fa17_xor1));
  and_gate and_gate_u_pg_rca24_and17(.a(u_pg_rca24_or16[0]), .b(u_pg_rca24_pg_fa17_xor0[0]), .out(u_pg_rca24_and17));
  or_gate or_gate_u_pg_rca24_or17(.a(u_pg_rca24_and17[0]), .b(u_pg_rca24_pg_fa17_and0[0]), .out(u_pg_rca24_or17));
  pg_fa pg_fa_u_pg_rca24_pg_fa18_out(.a(a[18]), .b(b[18]), .cin(u_pg_rca24_or17[0]), .pg_fa_xor0(u_pg_rca24_pg_fa18_xor0), .pg_fa_and0(u_pg_rca24_pg_fa18_and0), .pg_fa_xor1(u_pg_rca24_pg_fa18_xor1));
  and_gate and_gate_u_pg_rca24_and18(.a(u_pg_rca24_or17[0]), .b(u_pg_rca24_pg_fa18_xor0[0]), .out(u_pg_rca24_and18));
  or_gate or_gate_u_pg_rca24_or18(.a(u_pg_rca24_and18[0]), .b(u_pg_rca24_pg_fa18_and0[0]), .out(u_pg_rca24_or18));
  pg_fa pg_fa_u_pg_rca24_pg_fa19_out(.a(a[19]), .b(b[19]), .cin(u_pg_rca24_or18[0]), .pg_fa_xor0(u_pg_rca24_pg_fa19_xor0), .pg_fa_and0(u_pg_rca24_pg_fa19_and0), .pg_fa_xor1(u_pg_rca24_pg_fa19_xor1));
  and_gate and_gate_u_pg_rca24_and19(.a(u_pg_rca24_or18[0]), .b(u_pg_rca24_pg_fa19_xor0[0]), .out(u_pg_rca24_and19));
  or_gate or_gate_u_pg_rca24_or19(.a(u_pg_rca24_and19[0]), .b(u_pg_rca24_pg_fa19_and0[0]), .out(u_pg_rca24_or19));
  pg_fa pg_fa_u_pg_rca24_pg_fa20_out(.a(a[20]), .b(b[20]), .cin(u_pg_rca24_or19[0]), .pg_fa_xor0(u_pg_rca24_pg_fa20_xor0), .pg_fa_and0(u_pg_rca24_pg_fa20_and0), .pg_fa_xor1(u_pg_rca24_pg_fa20_xor1));
  and_gate and_gate_u_pg_rca24_and20(.a(u_pg_rca24_or19[0]), .b(u_pg_rca24_pg_fa20_xor0[0]), .out(u_pg_rca24_and20));
  or_gate or_gate_u_pg_rca24_or20(.a(u_pg_rca24_and20[0]), .b(u_pg_rca24_pg_fa20_and0[0]), .out(u_pg_rca24_or20));
  pg_fa pg_fa_u_pg_rca24_pg_fa21_out(.a(a[21]), .b(b[21]), .cin(u_pg_rca24_or20[0]), .pg_fa_xor0(u_pg_rca24_pg_fa21_xor0), .pg_fa_and0(u_pg_rca24_pg_fa21_and0), .pg_fa_xor1(u_pg_rca24_pg_fa21_xor1));
  and_gate and_gate_u_pg_rca24_and21(.a(u_pg_rca24_or20[0]), .b(u_pg_rca24_pg_fa21_xor0[0]), .out(u_pg_rca24_and21));
  or_gate or_gate_u_pg_rca24_or21(.a(u_pg_rca24_and21[0]), .b(u_pg_rca24_pg_fa21_and0[0]), .out(u_pg_rca24_or21));
  pg_fa pg_fa_u_pg_rca24_pg_fa22_out(.a(a[22]), .b(b[22]), .cin(u_pg_rca24_or21[0]), .pg_fa_xor0(u_pg_rca24_pg_fa22_xor0), .pg_fa_and0(u_pg_rca24_pg_fa22_and0), .pg_fa_xor1(u_pg_rca24_pg_fa22_xor1));
  and_gate and_gate_u_pg_rca24_and22(.a(u_pg_rca24_or21[0]), .b(u_pg_rca24_pg_fa22_xor0[0]), .out(u_pg_rca24_and22));
  or_gate or_gate_u_pg_rca24_or22(.a(u_pg_rca24_and22[0]), .b(u_pg_rca24_pg_fa22_and0[0]), .out(u_pg_rca24_or22));
  pg_fa pg_fa_u_pg_rca24_pg_fa23_out(.a(a[23]), .b(b[23]), .cin(u_pg_rca24_or22[0]), .pg_fa_xor0(u_pg_rca24_pg_fa23_xor0), .pg_fa_and0(u_pg_rca24_pg_fa23_and0), .pg_fa_xor1(u_pg_rca24_pg_fa23_xor1));
  and_gate and_gate_u_pg_rca24_and23(.a(u_pg_rca24_or22[0]), .b(u_pg_rca24_pg_fa23_xor0[0]), .out(u_pg_rca24_and23));
  or_gate or_gate_u_pg_rca24_or23(.a(u_pg_rca24_and23[0]), .b(u_pg_rca24_pg_fa23_and0[0]), .out(u_pg_rca24_or23));

  assign u_pg_rca24_out[0] = u_pg_rca24_pg_fa0_xor0[0];
  assign u_pg_rca24_out[1] = u_pg_rca24_pg_fa1_xor1[0];
  assign u_pg_rca24_out[2] = u_pg_rca24_pg_fa2_xor1[0];
  assign u_pg_rca24_out[3] = u_pg_rca24_pg_fa3_xor1[0];
  assign u_pg_rca24_out[4] = u_pg_rca24_pg_fa4_xor1[0];
  assign u_pg_rca24_out[5] = u_pg_rca24_pg_fa5_xor1[0];
  assign u_pg_rca24_out[6] = u_pg_rca24_pg_fa6_xor1[0];
  assign u_pg_rca24_out[7] = u_pg_rca24_pg_fa7_xor1[0];
  assign u_pg_rca24_out[8] = u_pg_rca24_pg_fa8_xor1[0];
  assign u_pg_rca24_out[9] = u_pg_rca24_pg_fa9_xor1[0];
  assign u_pg_rca24_out[10] = u_pg_rca24_pg_fa10_xor1[0];
  assign u_pg_rca24_out[11] = u_pg_rca24_pg_fa11_xor1[0];
  assign u_pg_rca24_out[12] = u_pg_rca24_pg_fa12_xor1[0];
  assign u_pg_rca24_out[13] = u_pg_rca24_pg_fa13_xor1[0];
  assign u_pg_rca24_out[14] = u_pg_rca24_pg_fa14_xor1[0];
  assign u_pg_rca24_out[15] = u_pg_rca24_pg_fa15_xor1[0];
  assign u_pg_rca24_out[16] = u_pg_rca24_pg_fa16_xor1[0];
  assign u_pg_rca24_out[17] = u_pg_rca24_pg_fa17_xor1[0];
  assign u_pg_rca24_out[18] = u_pg_rca24_pg_fa18_xor1[0];
  assign u_pg_rca24_out[19] = u_pg_rca24_pg_fa19_xor1[0];
  assign u_pg_rca24_out[20] = u_pg_rca24_pg_fa20_xor1[0];
  assign u_pg_rca24_out[21] = u_pg_rca24_pg_fa21_xor1[0];
  assign u_pg_rca24_out[22] = u_pg_rca24_pg_fa22_xor1[0];
  assign u_pg_rca24_out[23] = u_pg_rca24_pg_fa23_xor1[0];
  assign u_pg_rca24_out[24] = u_pg_rca24_or23[0];
endmodule

module u_csamul_pg_rca24(input [23:0] a, input [23:0] b, output [47:0] u_csamul_pg_rca24_out);
  wire [0:0] u_csamul_pg_rca24_and0_0;
  wire [0:0] u_csamul_pg_rca24_and1_0;
  wire [0:0] u_csamul_pg_rca24_and2_0;
  wire [0:0] u_csamul_pg_rca24_and3_0;
  wire [0:0] u_csamul_pg_rca24_and4_0;
  wire [0:0] u_csamul_pg_rca24_and5_0;
  wire [0:0] u_csamul_pg_rca24_and6_0;
  wire [0:0] u_csamul_pg_rca24_and7_0;
  wire [0:0] u_csamul_pg_rca24_and8_0;
  wire [0:0] u_csamul_pg_rca24_and9_0;
  wire [0:0] u_csamul_pg_rca24_and10_0;
  wire [0:0] u_csamul_pg_rca24_and11_0;
  wire [0:0] u_csamul_pg_rca24_and12_0;
  wire [0:0] u_csamul_pg_rca24_and13_0;
  wire [0:0] u_csamul_pg_rca24_and14_0;
  wire [0:0] u_csamul_pg_rca24_and15_0;
  wire [0:0] u_csamul_pg_rca24_and16_0;
  wire [0:0] u_csamul_pg_rca24_and17_0;
  wire [0:0] u_csamul_pg_rca24_and18_0;
  wire [0:0] u_csamul_pg_rca24_and19_0;
  wire [0:0] u_csamul_pg_rca24_and20_0;
  wire [0:0] u_csamul_pg_rca24_and21_0;
  wire [0:0] u_csamul_pg_rca24_and22_0;
  wire [0:0] u_csamul_pg_rca24_and23_0;
  wire [0:0] u_csamul_pg_rca24_and0_1;
  wire [0:0] u_csamul_pg_rca24_ha0_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha0_1_and0;
  wire [0:0] u_csamul_pg_rca24_and1_1;
  wire [0:0] u_csamul_pg_rca24_ha1_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha1_1_and0;
  wire [0:0] u_csamul_pg_rca24_and2_1;
  wire [0:0] u_csamul_pg_rca24_ha2_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha2_1_and0;
  wire [0:0] u_csamul_pg_rca24_and3_1;
  wire [0:0] u_csamul_pg_rca24_ha3_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha3_1_and0;
  wire [0:0] u_csamul_pg_rca24_and4_1;
  wire [0:0] u_csamul_pg_rca24_ha4_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha4_1_and0;
  wire [0:0] u_csamul_pg_rca24_and5_1;
  wire [0:0] u_csamul_pg_rca24_ha5_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha5_1_and0;
  wire [0:0] u_csamul_pg_rca24_and6_1;
  wire [0:0] u_csamul_pg_rca24_ha6_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha6_1_and0;
  wire [0:0] u_csamul_pg_rca24_and7_1;
  wire [0:0] u_csamul_pg_rca24_ha7_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha7_1_and0;
  wire [0:0] u_csamul_pg_rca24_and8_1;
  wire [0:0] u_csamul_pg_rca24_ha8_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha8_1_and0;
  wire [0:0] u_csamul_pg_rca24_and9_1;
  wire [0:0] u_csamul_pg_rca24_ha9_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha9_1_and0;
  wire [0:0] u_csamul_pg_rca24_and10_1;
  wire [0:0] u_csamul_pg_rca24_ha10_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha10_1_and0;
  wire [0:0] u_csamul_pg_rca24_and11_1;
  wire [0:0] u_csamul_pg_rca24_ha11_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha11_1_and0;
  wire [0:0] u_csamul_pg_rca24_and12_1;
  wire [0:0] u_csamul_pg_rca24_ha12_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha12_1_and0;
  wire [0:0] u_csamul_pg_rca24_and13_1;
  wire [0:0] u_csamul_pg_rca24_ha13_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha13_1_and0;
  wire [0:0] u_csamul_pg_rca24_and14_1;
  wire [0:0] u_csamul_pg_rca24_ha14_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha14_1_and0;
  wire [0:0] u_csamul_pg_rca24_and15_1;
  wire [0:0] u_csamul_pg_rca24_ha15_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha15_1_and0;
  wire [0:0] u_csamul_pg_rca24_and16_1;
  wire [0:0] u_csamul_pg_rca24_ha16_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha16_1_and0;
  wire [0:0] u_csamul_pg_rca24_and17_1;
  wire [0:0] u_csamul_pg_rca24_ha17_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha17_1_and0;
  wire [0:0] u_csamul_pg_rca24_and18_1;
  wire [0:0] u_csamul_pg_rca24_ha18_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha18_1_and0;
  wire [0:0] u_csamul_pg_rca24_and19_1;
  wire [0:0] u_csamul_pg_rca24_ha19_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha19_1_and0;
  wire [0:0] u_csamul_pg_rca24_and20_1;
  wire [0:0] u_csamul_pg_rca24_ha20_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha20_1_and0;
  wire [0:0] u_csamul_pg_rca24_and21_1;
  wire [0:0] u_csamul_pg_rca24_ha21_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha21_1_and0;
  wire [0:0] u_csamul_pg_rca24_and22_1;
  wire [0:0] u_csamul_pg_rca24_ha22_1_xor0;
  wire [0:0] u_csamul_pg_rca24_ha22_1_and0;
  wire [0:0] u_csamul_pg_rca24_and23_1;
  wire [0:0] u_csamul_pg_rca24_and0_2;
  wire [0:0] u_csamul_pg_rca24_fa0_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_2_or0;
  wire [0:0] u_csamul_pg_rca24_and1_2;
  wire [0:0] u_csamul_pg_rca24_fa1_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_2_or0;
  wire [0:0] u_csamul_pg_rca24_and2_2;
  wire [0:0] u_csamul_pg_rca24_fa2_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_2_or0;
  wire [0:0] u_csamul_pg_rca24_and3_2;
  wire [0:0] u_csamul_pg_rca24_fa3_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_2_or0;
  wire [0:0] u_csamul_pg_rca24_and4_2;
  wire [0:0] u_csamul_pg_rca24_fa4_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_2_or0;
  wire [0:0] u_csamul_pg_rca24_and5_2;
  wire [0:0] u_csamul_pg_rca24_fa5_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_2_or0;
  wire [0:0] u_csamul_pg_rca24_and6_2;
  wire [0:0] u_csamul_pg_rca24_fa6_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_2_or0;
  wire [0:0] u_csamul_pg_rca24_and7_2;
  wire [0:0] u_csamul_pg_rca24_fa7_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_2_or0;
  wire [0:0] u_csamul_pg_rca24_and8_2;
  wire [0:0] u_csamul_pg_rca24_fa8_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_2_or0;
  wire [0:0] u_csamul_pg_rca24_and9_2;
  wire [0:0] u_csamul_pg_rca24_fa9_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_2_or0;
  wire [0:0] u_csamul_pg_rca24_and10_2;
  wire [0:0] u_csamul_pg_rca24_fa10_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_2_or0;
  wire [0:0] u_csamul_pg_rca24_and11_2;
  wire [0:0] u_csamul_pg_rca24_fa11_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_2_or0;
  wire [0:0] u_csamul_pg_rca24_and12_2;
  wire [0:0] u_csamul_pg_rca24_fa12_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_2_or0;
  wire [0:0] u_csamul_pg_rca24_and13_2;
  wire [0:0] u_csamul_pg_rca24_fa13_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_2_or0;
  wire [0:0] u_csamul_pg_rca24_and14_2;
  wire [0:0] u_csamul_pg_rca24_fa14_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_2_or0;
  wire [0:0] u_csamul_pg_rca24_and15_2;
  wire [0:0] u_csamul_pg_rca24_fa15_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_2_or0;
  wire [0:0] u_csamul_pg_rca24_and16_2;
  wire [0:0] u_csamul_pg_rca24_fa16_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_2_or0;
  wire [0:0] u_csamul_pg_rca24_and17_2;
  wire [0:0] u_csamul_pg_rca24_fa17_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_2_or0;
  wire [0:0] u_csamul_pg_rca24_and18_2;
  wire [0:0] u_csamul_pg_rca24_fa18_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_2_or0;
  wire [0:0] u_csamul_pg_rca24_and19_2;
  wire [0:0] u_csamul_pg_rca24_fa19_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_2_or0;
  wire [0:0] u_csamul_pg_rca24_and20_2;
  wire [0:0] u_csamul_pg_rca24_fa20_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_2_or0;
  wire [0:0] u_csamul_pg_rca24_and21_2;
  wire [0:0] u_csamul_pg_rca24_fa21_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_2_or0;
  wire [0:0] u_csamul_pg_rca24_and22_2;
  wire [0:0] u_csamul_pg_rca24_fa22_2_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_2_or0;
  wire [0:0] u_csamul_pg_rca24_and23_2;
  wire [0:0] u_csamul_pg_rca24_and0_3;
  wire [0:0] u_csamul_pg_rca24_fa0_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_3_or0;
  wire [0:0] u_csamul_pg_rca24_and1_3;
  wire [0:0] u_csamul_pg_rca24_fa1_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_3_or0;
  wire [0:0] u_csamul_pg_rca24_and2_3;
  wire [0:0] u_csamul_pg_rca24_fa2_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_3_or0;
  wire [0:0] u_csamul_pg_rca24_and3_3;
  wire [0:0] u_csamul_pg_rca24_fa3_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_3_or0;
  wire [0:0] u_csamul_pg_rca24_and4_3;
  wire [0:0] u_csamul_pg_rca24_fa4_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_3_or0;
  wire [0:0] u_csamul_pg_rca24_and5_3;
  wire [0:0] u_csamul_pg_rca24_fa5_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_3_or0;
  wire [0:0] u_csamul_pg_rca24_and6_3;
  wire [0:0] u_csamul_pg_rca24_fa6_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_3_or0;
  wire [0:0] u_csamul_pg_rca24_and7_3;
  wire [0:0] u_csamul_pg_rca24_fa7_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_3_or0;
  wire [0:0] u_csamul_pg_rca24_and8_3;
  wire [0:0] u_csamul_pg_rca24_fa8_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_3_or0;
  wire [0:0] u_csamul_pg_rca24_and9_3;
  wire [0:0] u_csamul_pg_rca24_fa9_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_3_or0;
  wire [0:0] u_csamul_pg_rca24_and10_3;
  wire [0:0] u_csamul_pg_rca24_fa10_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_3_or0;
  wire [0:0] u_csamul_pg_rca24_and11_3;
  wire [0:0] u_csamul_pg_rca24_fa11_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_3_or0;
  wire [0:0] u_csamul_pg_rca24_and12_3;
  wire [0:0] u_csamul_pg_rca24_fa12_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_3_or0;
  wire [0:0] u_csamul_pg_rca24_and13_3;
  wire [0:0] u_csamul_pg_rca24_fa13_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_3_or0;
  wire [0:0] u_csamul_pg_rca24_and14_3;
  wire [0:0] u_csamul_pg_rca24_fa14_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_3_or0;
  wire [0:0] u_csamul_pg_rca24_and15_3;
  wire [0:0] u_csamul_pg_rca24_fa15_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_3_or0;
  wire [0:0] u_csamul_pg_rca24_and16_3;
  wire [0:0] u_csamul_pg_rca24_fa16_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_3_or0;
  wire [0:0] u_csamul_pg_rca24_and17_3;
  wire [0:0] u_csamul_pg_rca24_fa17_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_3_or0;
  wire [0:0] u_csamul_pg_rca24_and18_3;
  wire [0:0] u_csamul_pg_rca24_fa18_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_3_or0;
  wire [0:0] u_csamul_pg_rca24_and19_3;
  wire [0:0] u_csamul_pg_rca24_fa19_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_3_or0;
  wire [0:0] u_csamul_pg_rca24_and20_3;
  wire [0:0] u_csamul_pg_rca24_fa20_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_3_or0;
  wire [0:0] u_csamul_pg_rca24_and21_3;
  wire [0:0] u_csamul_pg_rca24_fa21_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_3_or0;
  wire [0:0] u_csamul_pg_rca24_and22_3;
  wire [0:0] u_csamul_pg_rca24_fa22_3_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_3_or0;
  wire [0:0] u_csamul_pg_rca24_and23_3;
  wire [0:0] u_csamul_pg_rca24_and0_4;
  wire [0:0] u_csamul_pg_rca24_fa0_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_4_or0;
  wire [0:0] u_csamul_pg_rca24_and1_4;
  wire [0:0] u_csamul_pg_rca24_fa1_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_4_or0;
  wire [0:0] u_csamul_pg_rca24_and2_4;
  wire [0:0] u_csamul_pg_rca24_fa2_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_4_or0;
  wire [0:0] u_csamul_pg_rca24_and3_4;
  wire [0:0] u_csamul_pg_rca24_fa3_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_4_or0;
  wire [0:0] u_csamul_pg_rca24_and4_4;
  wire [0:0] u_csamul_pg_rca24_fa4_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_4_or0;
  wire [0:0] u_csamul_pg_rca24_and5_4;
  wire [0:0] u_csamul_pg_rca24_fa5_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_4_or0;
  wire [0:0] u_csamul_pg_rca24_and6_4;
  wire [0:0] u_csamul_pg_rca24_fa6_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_4_or0;
  wire [0:0] u_csamul_pg_rca24_and7_4;
  wire [0:0] u_csamul_pg_rca24_fa7_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_4_or0;
  wire [0:0] u_csamul_pg_rca24_and8_4;
  wire [0:0] u_csamul_pg_rca24_fa8_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_4_or0;
  wire [0:0] u_csamul_pg_rca24_and9_4;
  wire [0:0] u_csamul_pg_rca24_fa9_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_4_or0;
  wire [0:0] u_csamul_pg_rca24_and10_4;
  wire [0:0] u_csamul_pg_rca24_fa10_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_4_or0;
  wire [0:0] u_csamul_pg_rca24_and11_4;
  wire [0:0] u_csamul_pg_rca24_fa11_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_4_or0;
  wire [0:0] u_csamul_pg_rca24_and12_4;
  wire [0:0] u_csamul_pg_rca24_fa12_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_4_or0;
  wire [0:0] u_csamul_pg_rca24_and13_4;
  wire [0:0] u_csamul_pg_rca24_fa13_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_4_or0;
  wire [0:0] u_csamul_pg_rca24_and14_4;
  wire [0:0] u_csamul_pg_rca24_fa14_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_4_or0;
  wire [0:0] u_csamul_pg_rca24_and15_4;
  wire [0:0] u_csamul_pg_rca24_fa15_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_4_or0;
  wire [0:0] u_csamul_pg_rca24_and16_4;
  wire [0:0] u_csamul_pg_rca24_fa16_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_4_or0;
  wire [0:0] u_csamul_pg_rca24_and17_4;
  wire [0:0] u_csamul_pg_rca24_fa17_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_4_or0;
  wire [0:0] u_csamul_pg_rca24_and18_4;
  wire [0:0] u_csamul_pg_rca24_fa18_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_4_or0;
  wire [0:0] u_csamul_pg_rca24_and19_4;
  wire [0:0] u_csamul_pg_rca24_fa19_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_4_or0;
  wire [0:0] u_csamul_pg_rca24_and20_4;
  wire [0:0] u_csamul_pg_rca24_fa20_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_4_or0;
  wire [0:0] u_csamul_pg_rca24_and21_4;
  wire [0:0] u_csamul_pg_rca24_fa21_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_4_or0;
  wire [0:0] u_csamul_pg_rca24_and22_4;
  wire [0:0] u_csamul_pg_rca24_fa22_4_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_4_or0;
  wire [0:0] u_csamul_pg_rca24_and23_4;
  wire [0:0] u_csamul_pg_rca24_and0_5;
  wire [0:0] u_csamul_pg_rca24_fa0_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_5_or0;
  wire [0:0] u_csamul_pg_rca24_and1_5;
  wire [0:0] u_csamul_pg_rca24_fa1_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_5_or0;
  wire [0:0] u_csamul_pg_rca24_and2_5;
  wire [0:0] u_csamul_pg_rca24_fa2_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_5_or0;
  wire [0:0] u_csamul_pg_rca24_and3_5;
  wire [0:0] u_csamul_pg_rca24_fa3_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_5_or0;
  wire [0:0] u_csamul_pg_rca24_and4_5;
  wire [0:0] u_csamul_pg_rca24_fa4_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_5_or0;
  wire [0:0] u_csamul_pg_rca24_and5_5;
  wire [0:0] u_csamul_pg_rca24_fa5_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_5_or0;
  wire [0:0] u_csamul_pg_rca24_and6_5;
  wire [0:0] u_csamul_pg_rca24_fa6_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_5_or0;
  wire [0:0] u_csamul_pg_rca24_and7_5;
  wire [0:0] u_csamul_pg_rca24_fa7_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_5_or0;
  wire [0:0] u_csamul_pg_rca24_and8_5;
  wire [0:0] u_csamul_pg_rca24_fa8_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_5_or0;
  wire [0:0] u_csamul_pg_rca24_and9_5;
  wire [0:0] u_csamul_pg_rca24_fa9_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_5_or0;
  wire [0:0] u_csamul_pg_rca24_and10_5;
  wire [0:0] u_csamul_pg_rca24_fa10_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_5_or0;
  wire [0:0] u_csamul_pg_rca24_and11_5;
  wire [0:0] u_csamul_pg_rca24_fa11_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_5_or0;
  wire [0:0] u_csamul_pg_rca24_and12_5;
  wire [0:0] u_csamul_pg_rca24_fa12_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_5_or0;
  wire [0:0] u_csamul_pg_rca24_and13_5;
  wire [0:0] u_csamul_pg_rca24_fa13_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_5_or0;
  wire [0:0] u_csamul_pg_rca24_and14_5;
  wire [0:0] u_csamul_pg_rca24_fa14_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_5_or0;
  wire [0:0] u_csamul_pg_rca24_and15_5;
  wire [0:0] u_csamul_pg_rca24_fa15_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_5_or0;
  wire [0:0] u_csamul_pg_rca24_and16_5;
  wire [0:0] u_csamul_pg_rca24_fa16_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_5_or0;
  wire [0:0] u_csamul_pg_rca24_and17_5;
  wire [0:0] u_csamul_pg_rca24_fa17_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_5_or0;
  wire [0:0] u_csamul_pg_rca24_and18_5;
  wire [0:0] u_csamul_pg_rca24_fa18_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_5_or0;
  wire [0:0] u_csamul_pg_rca24_and19_5;
  wire [0:0] u_csamul_pg_rca24_fa19_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_5_or0;
  wire [0:0] u_csamul_pg_rca24_and20_5;
  wire [0:0] u_csamul_pg_rca24_fa20_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_5_or0;
  wire [0:0] u_csamul_pg_rca24_and21_5;
  wire [0:0] u_csamul_pg_rca24_fa21_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_5_or0;
  wire [0:0] u_csamul_pg_rca24_and22_5;
  wire [0:0] u_csamul_pg_rca24_fa22_5_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_5_or0;
  wire [0:0] u_csamul_pg_rca24_and23_5;
  wire [0:0] u_csamul_pg_rca24_and0_6;
  wire [0:0] u_csamul_pg_rca24_fa0_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_6_or0;
  wire [0:0] u_csamul_pg_rca24_and1_6;
  wire [0:0] u_csamul_pg_rca24_fa1_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_6_or0;
  wire [0:0] u_csamul_pg_rca24_and2_6;
  wire [0:0] u_csamul_pg_rca24_fa2_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_6_or0;
  wire [0:0] u_csamul_pg_rca24_and3_6;
  wire [0:0] u_csamul_pg_rca24_fa3_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_6_or0;
  wire [0:0] u_csamul_pg_rca24_and4_6;
  wire [0:0] u_csamul_pg_rca24_fa4_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_6_or0;
  wire [0:0] u_csamul_pg_rca24_and5_6;
  wire [0:0] u_csamul_pg_rca24_fa5_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_6_or0;
  wire [0:0] u_csamul_pg_rca24_and6_6;
  wire [0:0] u_csamul_pg_rca24_fa6_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_6_or0;
  wire [0:0] u_csamul_pg_rca24_and7_6;
  wire [0:0] u_csamul_pg_rca24_fa7_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_6_or0;
  wire [0:0] u_csamul_pg_rca24_and8_6;
  wire [0:0] u_csamul_pg_rca24_fa8_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_6_or0;
  wire [0:0] u_csamul_pg_rca24_and9_6;
  wire [0:0] u_csamul_pg_rca24_fa9_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_6_or0;
  wire [0:0] u_csamul_pg_rca24_and10_6;
  wire [0:0] u_csamul_pg_rca24_fa10_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_6_or0;
  wire [0:0] u_csamul_pg_rca24_and11_6;
  wire [0:0] u_csamul_pg_rca24_fa11_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_6_or0;
  wire [0:0] u_csamul_pg_rca24_and12_6;
  wire [0:0] u_csamul_pg_rca24_fa12_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_6_or0;
  wire [0:0] u_csamul_pg_rca24_and13_6;
  wire [0:0] u_csamul_pg_rca24_fa13_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_6_or0;
  wire [0:0] u_csamul_pg_rca24_and14_6;
  wire [0:0] u_csamul_pg_rca24_fa14_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_6_or0;
  wire [0:0] u_csamul_pg_rca24_and15_6;
  wire [0:0] u_csamul_pg_rca24_fa15_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_6_or0;
  wire [0:0] u_csamul_pg_rca24_and16_6;
  wire [0:0] u_csamul_pg_rca24_fa16_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_6_or0;
  wire [0:0] u_csamul_pg_rca24_and17_6;
  wire [0:0] u_csamul_pg_rca24_fa17_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_6_or0;
  wire [0:0] u_csamul_pg_rca24_and18_6;
  wire [0:0] u_csamul_pg_rca24_fa18_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_6_or0;
  wire [0:0] u_csamul_pg_rca24_and19_6;
  wire [0:0] u_csamul_pg_rca24_fa19_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_6_or0;
  wire [0:0] u_csamul_pg_rca24_and20_6;
  wire [0:0] u_csamul_pg_rca24_fa20_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_6_or0;
  wire [0:0] u_csamul_pg_rca24_and21_6;
  wire [0:0] u_csamul_pg_rca24_fa21_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_6_or0;
  wire [0:0] u_csamul_pg_rca24_and22_6;
  wire [0:0] u_csamul_pg_rca24_fa22_6_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_6_or0;
  wire [0:0] u_csamul_pg_rca24_and23_6;
  wire [0:0] u_csamul_pg_rca24_and0_7;
  wire [0:0] u_csamul_pg_rca24_fa0_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_7_or0;
  wire [0:0] u_csamul_pg_rca24_and1_7;
  wire [0:0] u_csamul_pg_rca24_fa1_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_7_or0;
  wire [0:0] u_csamul_pg_rca24_and2_7;
  wire [0:0] u_csamul_pg_rca24_fa2_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_7_or0;
  wire [0:0] u_csamul_pg_rca24_and3_7;
  wire [0:0] u_csamul_pg_rca24_fa3_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_7_or0;
  wire [0:0] u_csamul_pg_rca24_and4_7;
  wire [0:0] u_csamul_pg_rca24_fa4_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_7_or0;
  wire [0:0] u_csamul_pg_rca24_and5_7;
  wire [0:0] u_csamul_pg_rca24_fa5_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_7_or0;
  wire [0:0] u_csamul_pg_rca24_and6_7;
  wire [0:0] u_csamul_pg_rca24_fa6_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_7_or0;
  wire [0:0] u_csamul_pg_rca24_and7_7;
  wire [0:0] u_csamul_pg_rca24_fa7_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_7_or0;
  wire [0:0] u_csamul_pg_rca24_and8_7;
  wire [0:0] u_csamul_pg_rca24_fa8_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_7_or0;
  wire [0:0] u_csamul_pg_rca24_and9_7;
  wire [0:0] u_csamul_pg_rca24_fa9_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_7_or0;
  wire [0:0] u_csamul_pg_rca24_and10_7;
  wire [0:0] u_csamul_pg_rca24_fa10_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_7_or0;
  wire [0:0] u_csamul_pg_rca24_and11_7;
  wire [0:0] u_csamul_pg_rca24_fa11_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_7_or0;
  wire [0:0] u_csamul_pg_rca24_and12_7;
  wire [0:0] u_csamul_pg_rca24_fa12_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_7_or0;
  wire [0:0] u_csamul_pg_rca24_and13_7;
  wire [0:0] u_csamul_pg_rca24_fa13_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_7_or0;
  wire [0:0] u_csamul_pg_rca24_and14_7;
  wire [0:0] u_csamul_pg_rca24_fa14_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_7_or0;
  wire [0:0] u_csamul_pg_rca24_and15_7;
  wire [0:0] u_csamul_pg_rca24_fa15_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_7_or0;
  wire [0:0] u_csamul_pg_rca24_and16_7;
  wire [0:0] u_csamul_pg_rca24_fa16_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_7_or0;
  wire [0:0] u_csamul_pg_rca24_and17_7;
  wire [0:0] u_csamul_pg_rca24_fa17_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_7_or0;
  wire [0:0] u_csamul_pg_rca24_and18_7;
  wire [0:0] u_csamul_pg_rca24_fa18_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_7_or0;
  wire [0:0] u_csamul_pg_rca24_and19_7;
  wire [0:0] u_csamul_pg_rca24_fa19_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_7_or0;
  wire [0:0] u_csamul_pg_rca24_and20_7;
  wire [0:0] u_csamul_pg_rca24_fa20_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_7_or0;
  wire [0:0] u_csamul_pg_rca24_and21_7;
  wire [0:0] u_csamul_pg_rca24_fa21_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_7_or0;
  wire [0:0] u_csamul_pg_rca24_and22_7;
  wire [0:0] u_csamul_pg_rca24_fa22_7_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_7_or0;
  wire [0:0] u_csamul_pg_rca24_and23_7;
  wire [0:0] u_csamul_pg_rca24_and0_8;
  wire [0:0] u_csamul_pg_rca24_fa0_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_8_or0;
  wire [0:0] u_csamul_pg_rca24_and1_8;
  wire [0:0] u_csamul_pg_rca24_fa1_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_8_or0;
  wire [0:0] u_csamul_pg_rca24_and2_8;
  wire [0:0] u_csamul_pg_rca24_fa2_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_8_or0;
  wire [0:0] u_csamul_pg_rca24_and3_8;
  wire [0:0] u_csamul_pg_rca24_fa3_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_8_or0;
  wire [0:0] u_csamul_pg_rca24_and4_8;
  wire [0:0] u_csamul_pg_rca24_fa4_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_8_or0;
  wire [0:0] u_csamul_pg_rca24_and5_8;
  wire [0:0] u_csamul_pg_rca24_fa5_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_8_or0;
  wire [0:0] u_csamul_pg_rca24_and6_8;
  wire [0:0] u_csamul_pg_rca24_fa6_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_8_or0;
  wire [0:0] u_csamul_pg_rca24_and7_8;
  wire [0:0] u_csamul_pg_rca24_fa7_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_8_or0;
  wire [0:0] u_csamul_pg_rca24_and8_8;
  wire [0:0] u_csamul_pg_rca24_fa8_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_8_or0;
  wire [0:0] u_csamul_pg_rca24_and9_8;
  wire [0:0] u_csamul_pg_rca24_fa9_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_8_or0;
  wire [0:0] u_csamul_pg_rca24_and10_8;
  wire [0:0] u_csamul_pg_rca24_fa10_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_8_or0;
  wire [0:0] u_csamul_pg_rca24_and11_8;
  wire [0:0] u_csamul_pg_rca24_fa11_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_8_or0;
  wire [0:0] u_csamul_pg_rca24_and12_8;
  wire [0:0] u_csamul_pg_rca24_fa12_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_8_or0;
  wire [0:0] u_csamul_pg_rca24_and13_8;
  wire [0:0] u_csamul_pg_rca24_fa13_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_8_or0;
  wire [0:0] u_csamul_pg_rca24_and14_8;
  wire [0:0] u_csamul_pg_rca24_fa14_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_8_or0;
  wire [0:0] u_csamul_pg_rca24_and15_8;
  wire [0:0] u_csamul_pg_rca24_fa15_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_8_or0;
  wire [0:0] u_csamul_pg_rca24_and16_8;
  wire [0:0] u_csamul_pg_rca24_fa16_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_8_or0;
  wire [0:0] u_csamul_pg_rca24_and17_8;
  wire [0:0] u_csamul_pg_rca24_fa17_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_8_or0;
  wire [0:0] u_csamul_pg_rca24_and18_8;
  wire [0:0] u_csamul_pg_rca24_fa18_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_8_or0;
  wire [0:0] u_csamul_pg_rca24_and19_8;
  wire [0:0] u_csamul_pg_rca24_fa19_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_8_or0;
  wire [0:0] u_csamul_pg_rca24_and20_8;
  wire [0:0] u_csamul_pg_rca24_fa20_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_8_or0;
  wire [0:0] u_csamul_pg_rca24_and21_8;
  wire [0:0] u_csamul_pg_rca24_fa21_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_8_or0;
  wire [0:0] u_csamul_pg_rca24_and22_8;
  wire [0:0] u_csamul_pg_rca24_fa22_8_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_8_or0;
  wire [0:0] u_csamul_pg_rca24_and23_8;
  wire [0:0] u_csamul_pg_rca24_and0_9;
  wire [0:0] u_csamul_pg_rca24_fa0_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_9_or0;
  wire [0:0] u_csamul_pg_rca24_and1_9;
  wire [0:0] u_csamul_pg_rca24_fa1_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_9_or0;
  wire [0:0] u_csamul_pg_rca24_and2_9;
  wire [0:0] u_csamul_pg_rca24_fa2_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_9_or0;
  wire [0:0] u_csamul_pg_rca24_and3_9;
  wire [0:0] u_csamul_pg_rca24_fa3_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_9_or0;
  wire [0:0] u_csamul_pg_rca24_and4_9;
  wire [0:0] u_csamul_pg_rca24_fa4_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_9_or0;
  wire [0:0] u_csamul_pg_rca24_and5_9;
  wire [0:0] u_csamul_pg_rca24_fa5_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_9_or0;
  wire [0:0] u_csamul_pg_rca24_and6_9;
  wire [0:0] u_csamul_pg_rca24_fa6_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_9_or0;
  wire [0:0] u_csamul_pg_rca24_and7_9;
  wire [0:0] u_csamul_pg_rca24_fa7_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_9_or0;
  wire [0:0] u_csamul_pg_rca24_and8_9;
  wire [0:0] u_csamul_pg_rca24_fa8_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_9_or0;
  wire [0:0] u_csamul_pg_rca24_and9_9;
  wire [0:0] u_csamul_pg_rca24_fa9_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_9_or0;
  wire [0:0] u_csamul_pg_rca24_and10_9;
  wire [0:0] u_csamul_pg_rca24_fa10_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_9_or0;
  wire [0:0] u_csamul_pg_rca24_and11_9;
  wire [0:0] u_csamul_pg_rca24_fa11_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_9_or0;
  wire [0:0] u_csamul_pg_rca24_and12_9;
  wire [0:0] u_csamul_pg_rca24_fa12_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_9_or0;
  wire [0:0] u_csamul_pg_rca24_and13_9;
  wire [0:0] u_csamul_pg_rca24_fa13_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_9_or0;
  wire [0:0] u_csamul_pg_rca24_and14_9;
  wire [0:0] u_csamul_pg_rca24_fa14_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_9_or0;
  wire [0:0] u_csamul_pg_rca24_and15_9;
  wire [0:0] u_csamul_pg_rca24_fa15_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_9_or0;
  wire [0:0] u_csamul_pg_rca24_and16_9;
  wire [0:0] u_csamul_pg_rca24_fa16_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_9_or0;
  wire [0:0] u_csamul_pg_rca24_and17_9;
  wire [0:0] u_csamul_pg_rca24_fa17_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_9_or0;
  wire [0:0] u_csamul_pg_rca24_and18_9;
  wire [0:0] u_csamul_pg_rca24_fa18_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_9_or0;
  wire [0:0] u_csamul_pg_rca24_and19_9;
  wire [0:0] u_csamul_pg_rca24_fa19_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_9_or0;
  wire [0:0] u_csamul_pg_rca24_and20_9;
  wire [0:0] u_csamul_pg_rca24_fa20_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_9_or0;
  wire [0:0] u_csamul_pg_rca24_and21_9;
  wire [0:0] u_csamul_pg_rca24_fa21_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_9_or0;
  wire [0:0] u_csamul_pg_rca24_and22_9;
  wire [0:0] u_csamul_pg_rca24_fa22_9_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_9_or0;
  wire [0:0] u_csamul_pg_rca24_and23_9;
  wire [0:0] u_csamul_pg_rca24_and0_10;
  wire [0:0] u_csamul_pg_rca24_fa0_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_10_or0;
  wire [0:0] u_csamul_pg_rca24_and1_10;
  wire [0:0] u_csamul_pg_rca24_fa1_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_10_or0;
  wire [0:0] u_csamul_pg_rca24_and2_10;
  wire [0:0] u_csamul_pg_rca24_fa2_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_10_or0;
  wire [0:0] u_csamul_pg_rca24_and3_10;
  wire [0:0] u_csamul_pg_rca24_fa3_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_10_or0;
  wire [0:0] u_csamul_pg_rca24_and4_10;
  wire [0:0] u_csamul_pg_rca24_fa4_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_10_or0;
  wire [0:0] u_csamul_pg_rca24_and5_10;
  wire [0:0] u_csamul_pg_rca24_fa5_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_10_or0;
  wire [0:0] u_csamul_pg_rca24_and6_10;
  wire [0:0] u_csamul_pg_rca24_fa6_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_10_or0;
  wire [0:0] u_csamul_pg_rca24_and7_10;
  wire [0:0] u_csamul_pg_rca24_fa7_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_10_or0;
  wire [0:0] u_csamul_pg_rca24_and8_10;
  wire [0:0] u_csamul_pg_rca24_fa8_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_10_or0;
  wire [0:0] u_csamul_pg_rca24_and9_10;
  wire [0:0] u_csamul_pg_rca24_fa9_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_10_or0;
  wire [0:0] u_csamul_pg_rca24_and10_10;
  wire [0:0] u_csamul_pg_rca24_fa10_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_10_or0;
  wire [0:0] u_csamul_pg_rca24_and11_10;
  wire [0:0] u_csamul_pg_rca24_fa11_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_10_or0;
  wire [0:0] u_csamul_pg_rca24_and12_10;
  wire [0:0] u_csamul_pg_rca24_fa12_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_10_or0;
  wire [0:0] u_csamul_pg_rca24_and13_10;
  wire [0:0] u_csamul_pg_rca24_fa13_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_10_or0;
  wire [0:0] u_csamul_pg_rca24_and14_10;
  wire [0:0] u_csamul_pg_rca24_fa14_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_10_or0;
  wire [0:0] u_csamul_pg_rca24_and15_10;
  wire [0:0] u_csamul_pg_rca24_fa15_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_10_or0;
  wire [0:0] u_csamul_pg_rca24_and16_10;
  wire [0:0] u_csamul_pg_rca24_fa16_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_10_or0;
  wire [0:0] u_csamul_pg_rca24_and17_10;
  wire [0:0] u_csamul_pg_rca24_fa17_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_10_or0;
  wire [0:0] u_csamul_pg_rca24_and18_10;
  wire [0:0] u_csamul_pg_rca24_fa18_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_10_or0;
  wire [0:0] u_csamul_pg_rca24_and19_10;
  wire [0:0] u_csamul_pg_rca24_fa19_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_10_or0;
  wire [0:0] u_csamul_pg_rca24_and20_10;
  wire [0:0] u_csamul_pg_rca24_fa20_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_10_or0;
  wire [0:0] u_csamul_pg_rca24_and21_10;
  wire [0:0] u_csamul_pg_rca24_fa21_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_10_or0;
  wire [0:0] u_csamul_pg_rca24_and22_10;
  wire [0:0] u_csamul_pg_rca24_fa22_10_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_10_or0;
  wire [0:0] u_csamul_pg_rca24_and23_10;
  wire [0:0] u_csamul_pg_rca24_and0_11;
  wire [0:0] u_csamul_pg_rca24_fa0_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_11_or0;
  wire [0:0] u_csamul_pg_rca24_and1_11;
  wire [0:0] u_csamul_pg_rca24_fa1_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_11_or0;
  wire [0:0] u_csamul_pg_rca24_and2_11;
  wire [0:0] u_csamul_pg_rca24_fa2_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_11_or0;
  wire [0:0] u_csamul_pg_rca24_and3_11;
  wire [0:0] u_csamul_pg_rca24_fa3_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_11_or0;
  wire [0:0] u_csamul_pg_rca24_and4_11;
  wire [0:0] u_csamul_pg_rca24_fa4_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_11_or0;
  wire [0:0] u_csamul_pg_rca24_and5_11;
  wire [0:0] u_csamul_pg_rca24_fa5_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_11_or0;
  wire [0:0] u_csamul_pg_rca24_and6_11;
  wire [0:0] u_csamul_pg_rca24_fa6_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_11_or0;
  wire [0:0] u_csamul_pg_rca24_and7_11;
  wire [0:0] u_csamul_pg_rca24_fa7_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_11_or0;
  wire [0:0] u_csamul_pg_rca24_and8_11;
  wire [0:0] u_csamul_pg_rca24_fa8_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_11_or0;
  wire [0:0] u_csamul_pg_rca24_and9_11;
  wire [0:0] u_csamul_pg_rca24_fa9_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_11_or0;
  wire [0:0] u_csamul_pg_rca24_and10_11;
  wire [0:0] u_csamul_pg_rca24_fa10_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_11_or0;
  wire [0:0] u_csamul_pg_rca24_and11_11;
  wire [0:0] u_csamul_pg_rca24_fa11_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_11_or0;
  wire [0:0] u_csamul_pg_rca24_and12_11;
  wire [0:0] u_csamul_pg_rca24_fa12_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_11_or0;
  wire [0:0] u_csamul_pg_rca24_and13_11;
  wire [0:0] u_csamul_pg_rca24_fa13_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_11_or0;
  wire [0:0] u_csamul_pg_rca24_and14_11;
  wire [0:0] u_csamul_pg_rca24_fa14_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_11_or0;
  wire [0:0] u_csamul_pg_rca24_and15_11;
  wire [0:0] u_csamul_pg_rca24_fa15_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_11_or0;
  wire [0:0] u_csamul_pg_rca24_and16_11;
  wire [0:0] u_csamul_pg_rca24_fa16_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_11_or0;
  wire [0:0] u_csamul_pg_rca24_and17_11;
  wire [0:0] u_csamul_pg_rca24_fa17_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_11_or0;
  wire [0:0] u_csamul_pg_rca24_and18_11;
  wire [0:0] u_csamul_pg_rca24_fa18_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_11_or0;
  wire [0:0] u_csamul_pg_rca24_and19_11;
  wire [0:0] u_csamul_pg_rca24_fa19_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_11_or0;
  wire [0:0] u_csamul_pg_rca24_and20_11;
  wire [0:0] u_csamul_pg_rca24_fa20_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_11_or0;
  wire [0:0] u_csamul_pg_rca24_and21_11;
  wire [0:0] u_csamul_pg_rca24_fa21_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_11_or0;
  wire [0:0] u_csamul_pg_rca24_and22_11;
  wire [0:0] u_csamul_pg_rca24_fa22_11_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_11_or0;
  wire [0:0] u_csamul_pg_rca24_and23_11;
  wire [0:0] u_csamul_pg_rca24_and0_12;
  wire [0:0] u_csamul_pg_rca24_fa0_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_12_or0;
  wire [0:0] u_csamul_pg_rca24_and1_12;
  wire [0:0] u_csamul_pg_rca24_fa1_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_12_or0;
  wire [0:0] u_csamul_pg_rca24_and2_12;
  wire [0:0] u_csamul_pg_rca24_fa2_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_12_or0;
  wire [0:0] u_csamul_pg_rca24_and3_12;
  wire [0:0] u_csamul_pg_rca24_fa3_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_12_or0;
  wire [0:0] u_csamul_pg_rca24_and4_12;
  wire [0:0] u_csamul_pg_rca24_fa4_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_12_or0;
  wire [0:0] u_csamul_pg_rca24_and5_12;
  wire [0:0] u_csamul_pg_rca24_fa5_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_12_or0;
  wire [0:0] u_csamul_pg_rca24_and6_12;
  wire [0:0] u_csamul_pg_rca24_fa6_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_12_or0;
  wire [0:0] u_csamul_pg_rca24_and7_12;
  wire [0:0] u_csamul_pg_rca24_fa7_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_12_or0;
  wire [0:0] u_csamul_pg_rca24_and8_12;
  wire [0:0] u_csamul_pg_rca24_fa8_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_12_or0;
  wire [0:0] u_csamul_pg_rca24_and9_12;
  wire [0:0] u_csamul_pg_rca24_fa9_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_12_or0;
  wire [0:0] u_csamul_pg_rca24_and10_12;
  wire [0:0] u_csamul_pg_rca24_fa10_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_12_or0;
  wire [0:0] u_csamul_pg_rca24_and11_12;
  wire [0:0] u_csamul_pg_rca24_fa11_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_12_or0;
  wire [0:0] u_csamul_pg_rca24_and12_12;
  wire [0:0] u_csamul_pg_rca24_fa12_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_12_or0;
  wire [0:0] u_csamul_pg_rca24_and13_12;
  wire [0:0] u_csamul_pg_rca24_fa13_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_12_or0;
  wire [0:0] u_csamul_pg_rca24_and14_12;
  wire [0:0] u_csamul_pg_rca24_fa14_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_12_or0;
  wire [0:0] u_csamul_pg_rca24_and15_12;
  wire [0:0] u_csamul_pg_rca24_fa15_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_12_or0;
  wire [0:0] u_csamul_pg_rca24_and16_12;
  wire [0:0] u_csamul_pg_rca24_fa16_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_12_or0;
  wire [0:0] u_csamul_pg_rca24_and17_12;
  wire [0:0] u_csamul_pg_rca24_fa17_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_12_or0;
  wire [0:0] u_csamul_pg_rca24_and18_12;
  wire [0:0] u_csamul_pg_rca24_fa18_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_12_or0;
  wire [0:0] u_csamul_pg_rca24_and19_12;
  wire [0:0] u_csamul_pg_rca24_fa19_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_12_or0;
  wire [0:0] u_csamul_pg_rca24_and20_12;
  wire [0:0] u_csamul_pg_rca24_fa20_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_12_or0;
  wire [0:0] u_csamul_pg_rca24_and21_12;
  wire [0:0] u_csamul_pg_rca24_fa21_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_12_or0;
  wire [0:0] u_csamul_pg_rca24_and22_12;
  wire [0:0] u_csamul_pg_rca24_fa22_12_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_12_or0;
  wire [0:0] u_csamul_pg_rca24_and23_12;
  wire [0:0] u_csamul_pg_rca24_and0_13;
  wire [0:0] u_csamul_pg_rca24_fa0_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_13_or0;
  wire [0:0] u_csamul_pg_rca24_and1_13;
  wire [0:0] u_csamul_pg_rca24_fa1_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_13_or0;
  wire [0:0] u_csamul_pg_rca24_and2_13;
  wire [0:0] u_csamul_pg_rca24_fa2_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_13_or0;
  wire [0:0] u_csamul_pg_rca24_and3_13;
  wire [0:0] u_csamul_pg_rca24_fa3_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_13_or0;
  wire [0:0] u_csamul_pg_rca24_and4_13;
  wire [0:0] u_csamul_pg_rca24_fa4_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_13_or0;
  wire [0:0] u_csamul_pg_rca24_and5_13;
  wire [0:0] u_csamul_pg_rca24_fa5_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_13_or0;
  wire [0:0] u_csamul_pg_rca24_and6_13;
  wire [0:0] u_csamul_pg_rca24_fa6_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_13_or0;
  wire [0:0] u_csamul_pg_rca24_and7_13;
  wire [0:0] u_csamul_pg_rca24_fa7_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_13_or0;
  wire [0:0] u_csamul_pg_rca24_and8_13;
  wire [0:0] u_csamul_pg_rca24_fa8_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_13_or0;
  wire [0:0] u_csamul_pg_rca24_and9_13;
  wire [0:0] u_csamul_pg_rca24_fa9_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_13_or0;
  wire [0:0] u_csamul_pg_rca24_and10_13;
  wire [0:0] u_csamul_pg_rca24_fa10_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_13_or0;
  wire [0:0] u_csamul_pg_rca24_and11_13;
  wire [0:0] u_csamul_pg_rca24_fa11_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_13_or0;
  wire [0:0] u_csamul_pg_rca24_and12_13;
  wire [0:0] u_csamul_pg_rca24_fa12_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_13_or0;
  wire [0:0] u_csamul_pg_rca24_and13_13;
  wire [0:0] u_csamul_pg_rca24_fa13_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_13_or0;
  wire [0:0] u_csamul_pg_rca24_and14_13;
  wire [0:0] u_csamul_pg_rca24_fa14_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_13_or0;
  wire [0:0] u_csamul_pg_rca24_and15_13;
  wire [0:0] u_csamul_pg_rca24_fa15_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_13_or0;
  wire [0:0] u_csamul_pg_rca24_and16_13;
  wire [0:0] u_csamul_pg_rca24_fa16_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_13_or0;
  wire [0:0] u_csamul_pg_rca24_and17_13;
  wire [0:0] u_csamul_pg_rca24_fa17_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_13_or0;
  wire [0:0] u_csamul_pg_rca24_and18_13;
  wire [0:0] u_csamul_pg_rca24_fa18_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_13_or0;
  wire [0:0] u_csamul_pg_rca24_and19_13;
  wire [0:0] u_csamul_pg_rca24_fa19_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_13_or0;
  wire [0:0] u_csamul_pg_rca24_and20_13;
  wire [0:0] u_csamul_pg_rca24_fa20_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_13_or0;
  wire [0:0] u_csamul_pg_rca24_and21_13;
  wire [0:0] u_csamul_pg_rca24_fa21_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_13_or0;
  wire [0:0] u_csamul_pg_rca24_and22_13;
  wire [0:0] u_csamul_pg_rca24_fa22_13_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_13_or0;
  wire [0:0] u_csamul_pg_rca24_and23_13;
  wire [0:0] u_csamul_pg_rca24_and0_14;
  wire [0:0] u_csamul_pg_rca24_fa0_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_14_or0;
  wire [0:0] u_csamul_pg_rca24_and1_14;
  wire [0:0] u_csamul_pg_rca24_fa1_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_14_or0;
  wire [0:0] u_csamul_pg_rca24_and2_14;
  wire [0:0] u_csamul_pg_rca24_fa2_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_14_or0;
  wire [0:0] u_csamul_pg_rca24_and3_14;
  wire [0:0] u_csamul_pg_rca24_fa3_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_14_or0;
  wire [0:0] u_csamul_pg_rca24_and4_14;
  wire [0:0] u_csamul_pg_rca24_fa4_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_14_or0;
  wire [0:0] u_csamul_pg_rca24_and5_14;
  wire [0:0] u_csamul_pg_rca24_fa5_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_14_or0;
  wire [0:0] u_csamul_pg_rca24_and6_14;
  wire [0:0] u_csamul_pg_rca24_fa6_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_14_or0;
  wire [0:0] u_csamul_pg_rca24_and7_14;
  wire [0:0] u_csamul_pg_rca24_fa7_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_14_or0;
  wire [0:0] u_csamul_pg_rca24_and8_14;
  wire [0:0] u_csamul_pg_rca24_fa8_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_14_or0;
  wire [0:0] u_csamul_pg_rca24_and9_14;
  wire [0:0] u_csamul_pg_rca24_fa9_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_14_or0;
  wire [0:0] u_csamul_pg_rca24_and10_14;
  wire [0:0] u_csamul_pg_rca24_fa10_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_14_or0;
  wire [0:0] u_csamul_pg_rca24_and11_14;
  wire [0:0] u_csamul_pg_rca24_fa11_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_14_or0;
  wire [0:0] u_csamul_pg_rca24_and12_14;
  wire [0:0] u_csamul_pg_rca24_fa12_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_14_or0;
  wire [0:0] u_csamul_pg_rca24_and13_14;
  wire [0:0] u_csamul_pg_rca24_fa13_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_14_or0;
  wire [0:0] u_csamul_pg_rca24_and14_14;
  wire [0:0] u_csamul_pg_rca24_fa14_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_14_or0;
  wire [0:0] u_csamul_pg_rca24_and15_14;
  wire [0:0] u_csamul_pg_rca24_fa15_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_14_or0;
  wire [0:0] u_csamul_pg_rca24_and16_14;
  wire [0:0] u_csamul_pg_rca24_fa16_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_14_or0;
  wire [0:0] u_csamul_pg_rca24_and17_14;
  wire [0:0] u_csamul_pg_rca24_fa17_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_14_or0;
  wire [0:0] u_csamul_pg_rca24_and18_14;
  wire [0:0] u_csamul_pg_rca24_fa18_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_14_or0;
  wire [0:0] u_csamul_pg_rca24_and19_14;
  wire [0:0] u_csamul_pg_rca24_fa19_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_14_or0;
  wire [0:0] u_csamul_pg_rca24_and20_14;
  wire [0:0] u_csamul_pg_rca24_fa20_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_14_or0;
  wire [0:0] u_csamul_pg_rca24_and21_14;
  wire [0:0] u_csamul_pg_rca24_fa21_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_14_or0;
  wire [0:0] u_csamul_pg_rca24_and22_14;
  wire [0:0] u_csamul_pg_rca24_fa22_14_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_14_or0;
  wire [0:0] u_csamul_pg_rca24_and23_14;
  wire [0:0] u_csamul_pg_rca24_and0_15;
  wire [0:0] u_csamul_pg_rca24_fa0_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_15_or0;
  wire [0:0] u_csamul_pg_rca24_and1_15;
  wire [0:0] u_csamul_pg_rca24_fa1_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_15_or0;
  wire [0:0] u_csamul_pg_rca24_and2_15;
  wire [0:0] u_csamul_pg_rca24_fa2_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_15_or0;
  wire [0:0] u_csamul_pg_rca24_and3_15;
  wire [0:0] u_csamul_pg_rca24_fa3_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_15_or0;
  wire [0:0] u_csamul_pg_rca24_and4_15;
  wire [0:0] u_csamul_pg_rca24_fa4_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_15_or0;
  wire [0:0] u_csamul_pg_rca24_and5_15;
  wire [0:0] u_csamul_pg_rca24_fa5_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_15_or0;
  wire [0:0] u_csamul_pg_rca24_and6_15;
  wire [0:0] u_csamul_pg_rca24_fa6_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_15_or0;
  wire [0:0] u_csamul_pg_rca24_and7_15;
  wire [0:0] u_csamul_pg_rca24_fa7_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_15_or0;
  wire [0:0] u_csamul_pg_rca24_and8_15;
  wire [0:0] u_csamul_pg_rca24_fa8_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_15_or0;
  wire [0:0] u_csamul_pg_rca24_and9_15;
  wire [0:0] u_csamul_pg_rca24_fa9_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_15_or0;
  wire [0:0] u_csamul_pg_rca24_and10_15;
  wire [0:0] u_csamul_pg_rca24_fa10_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_15_or0;
  wire [0:0] u_csamul_pg_rca24_and11_15;
  wire [0:0] u_csamul_pg_rca24_fa11_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_15_or0;
  wire [0:0] u_csamul_pg_rca24_and12_15;
  wire [0:0] u_csamul_pg_rca24_fa12_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_15_or0;
  wire [0:0] u_csamul_pg_rca24_and13_15;
  wire [0:0] u_csamul_pg_rca24_fa13_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_15_or0;
  wire [0:0] u_csamul_pg_rca24_and14_15;
  wire [0:0] u_csamul_pg_rca24_fa14_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_15_or0;
  wire [0:0] u_csamul_pg_rca24_and15_15;
  wire [0:0] u_csamul_pg_rca24_fa15_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_15_or0;
  wire [0:0] u_csamul_pg_rca24_and16_15;
  wire [0:0] u_csamul_pg_rca24_fa16_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_15_or0;
  wire [0:0] u_csamul_pg_rca24_and17_15;
  wire [0:0] u_csamul_pg_rca24_fa17_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_15_or0;
  wire [0:0] u_csamul_pg_rca24_and18_15;
  wire [0:0] u_csamul_pg_rca24_fa18_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_15_or0;
  wire [0:0] u_csamul_pg_rca24_and19_15;
  wire [0:0] u_csamul_pg_rca24_fa19_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_15_or0;
  wire [0:0] u_csamul_pg_rca24_and20_15;
  wire [0:0] u_csamul_pg_rca24_fa20_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_15_or0;
  wire [0:0] u_csamul_pg_rca24_and21_15;
  wire [0:0] u_csamul_pg_rca24_fa21_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_15_or0;
  wire [0:0] u_csamul_pg_rca24_and22_15;
  wire [0:0] u_csamul_pg_rca24_fa22_15_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_15_or0;
  wire [0:0] u_csamul_pg_rca24_and23_15;
  wire [0:0] u_csamul_pg_rca24_and0_16;
  wire [0:0] u_csamul_pg_rca24_fa0_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_16_or0;
  wire [0:0] u_csamul_pg_rca24_and1_16;
  wire [0:0] u_csamul_pg_rca24_fa1_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_16_or0;
  wire [0:0] u_csamul_pg_rca24_and2_16;
  wire [0:0] u_csamul_pg_rca24_fa2_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_16_or0;
  wire [0:0] u_csamul_pg_rca24_and3_16;
  wire [0:0] u_csamul_pg_rca24_fa3_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_16_or0;
  wire [0:0] u_csamul_pg_rca24_and4_16;
  wire [0:0] u_csamul_pg_rca24_fa4_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_16_or0;
  wire [0:0] u_csamul_pg_rca24_and5_16;
  wire [0:0] u_csamul_pg_rca24_fa5_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_16_or0;
  wire [0:0] u_csamul_pg_rca24_and6_16;
  wire [0:0] u_csamul_pg_rca24_fa6_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_16_or0;
  wire [0:0] u_csamul_pg_rca24_and7_16;
  wire [0:0] u_csamul_pg_rca24_fa7_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_16_or0;
  wire [0:0] u_csamul_pg_rca24_and8_16;
  wire [0:0] u_csamul_pg_rca24_fa8_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_16_or0;
  wire [0:0] u_csamul_pg_rca24_and9_16;
  wire [0:0] u_csamul_pg_rca24_fa9_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_16_or0;
  wire [0:0] u_csamul_pg_rca24_and10_16;
  wire [0:0] u_csamul_pg_rca24_fa10_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_16_or0;
  wire [0:0] u_csamul_pg_rca24_and11_16;
  wire [0:0] u_csamul_pg_rca24_fa11_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_16_or0;
  wire [0:0] u_csamul_pg_rca24_and12_16;
  wire [0:0] u_csamul_pg_rca24_fa12_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_16_or0;
  wire [0:0] u_csamul_pg_rca24_and13_16;
  wire [0:0] u_csamul_pg_rca24_fa13_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_16_or0;
  wire [0:0] u_csamul_pg_rca24_and14_16;
  wire [0:0] u_csamul_pg_rca24_fa14_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_16_or0;
  wire [0:0] u_csamul_pg_rca24_and15_16;
  wire [0:0] u_csamul_pg_rca24_fa15_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_16_or0;
  wire [0:0] u_csamul_pg_rca24_and16_16;
  wire [0:0] u_csamul_pg_rca24_fa16_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_16_or0;
  wire [0:0] u_csamul_pg_rca24_and17_16;
  wire [0:0] u_csamul_pg_rca24_fa17_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_16_or0;
  wire [0:0] u_csamul_pg_rca24_and18_16;
  wire [0:0] u_csamul_pg_rca24_fa18_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_16_or0;
  wire [0:0] u_csamul_pg_rca24_and19_16;
  wire [0:0] u_csamul_pg_rca24_fa19_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_16_or0;
  wire [0:0] u_csamul_pg_rca24_and20_16;
  wire [0:0] u_csamul_pg_rca24_fa20_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_16_or0;
  wire [0:0] u_csamul_pg_rca24_and21_16;
  wire [0:0] u_csamul_pg_rca24_fa21_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_16_or0;
  wire [0:0] u_csamul_pg_rca24_and22_16;
  wire [0:0] u_csamul_pg_rca24_fa22_16_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_16_or0;
  wire [0:0] u_csamul_pg_rca24_and23_16;
  wire [0:0] u_csamul_pg_rca24_and0_17;
  wire [0:0] u_csamul_pg_rca24_fa0_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_17_or0;
  wire [0:0] u_csamul_pg_rca24_and1_17;
  wire [0:0] u_csamul_pg_rca24_fa1_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_17_or0;
  wire [0:0] u_csamul_pg_rca24_and2_17;
  wire [0:0] u_csamul_pg_rca24_fa2_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_17_or0;
  wire [0:0] u_csamul_pg_rca24_and3_17;
  wire [0:0] u_csamul_pg_rca24_fa3_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_17_or0;
  wire [0:0] u_csamul_pg_rca24_and4_17;
  wire [0:0] u_csamul_pg_rca24_fa4_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_17_or0;
  wire [0:0] u_csamul_pg_rca24_and5_17;
  wire [0:0] u_csamul_pg_rca24_fa5_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_17_or0;
  wire [0:0] u_csamul_pg_rca24_and6_17;
  wire [0:0] u_csamul_pg_rca24_fa6_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_17_or0;
  wire [0:0] u_csamul_pg_rca24_and7_17;
  wire [0:0] u_csamul_pg_rca24_fa7_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_17_or0;
  wire [0:0] u_csamul_pg_rca24_and8_17;
  wire [0:0] u_csamul_pg_rca24_fa8_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_17_or0;
  wire [0:0] u_csamul_pg_rca24_and9_17;
  wire [0:0] u_csamul_pg_rca24_fa9_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_17_or0;
  wire [0:0] u_csamul_pg_rca24_and10_17;
  wire [0:0] u_csamul_pg_rca24_fa10_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_17_or0;
  wire [0:0] u_csamul_pg_rca24_and11_17;
  wire [0:0] u_csamul_pg_rca24_fa11_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_17_or0;
  wire [0:0] u_csamul_pg_rca24_and12_17;
  wire [0:0] u_csamul_pg_rca24_fa12_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_17_or0;
  wire [0:0] u_csamul_pg_rca24_and13_17;
  wire [0:0] u_csamul_pg_rca24_fa13_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_17_or0;
  wire [0:0] u_csamul_pg_rca24_and14_17;
  wire [0:0] u_csamul_pg_rca24_fa14_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_17_or0;
  wire [0:0] u_csamul_pg_rca24_and15_17;
  wire [0:0] u_csamul_pg_rca24_fa15_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_17_or0;
  wire [0:0] u_csamul_pg_rca24_and16_17;
  wire [0:0] u_csamul_pg_rca24_fa16_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_17_or0;
  wire [0:0] u_csamul_pg_rca24_and17_17;
  wire [0:0] u_csamul_pg_rca24_fa17_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_17_or0;
  wire [0:0] u_csamul_pg_rca24_and18_17;
  wire [0:0] u_csamul_pg_rca24_fa18_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_17_or0;
  wire [0:0] u_csamul_pg_rca24_and19_17;
  wire [0:0] u_csamul_pg_rca24_fa19_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_17_or0;
  wire [0:0] u_csamul_pg_rca24_and20_17;
  wire [0:0] u_csamul_pg_rca24_fa20_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_17_or0;
  wire [0:0] u_csamul_pg_rca24_and21_17;
  wire [0:0] u_csamul_pg_rca24_fa21_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_17_or0;
  wire [0:0] u_csamul_pg_rca24_and22_17;
  wire [0:0] u_csamul_pg_rca24_fa22_17_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_17_or0;
  wire [0:0] u_csamul_pg_rca24_and23_17;
  wire [0:0] u_csamul_pg_rca24_and0_18;
  wire [0:0] u_csamul_pg_rca24_fa0_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_18_or0;
  wire [0:0] u_csamul_pg_rca24_and1_18;
  wire [0:0] u_csamul_pg_rca24_fa1_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_18_or0;
  wire [0:0] u_csamul_pg_rca24_and2_18;
  wire [0:0] u_csamul_pg_rca24_fa2_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_18_or0;
  wire [0:0] u_csamul_pg_rca24_and3_18;
  wire [0:0] u_csamul_pg_rca24_fa3_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_18_or0;
  wire [0:0] u_csamul_pg_rca24_and4_18;
  wire [0:0] u_csamul_pg_rca24_fa4_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_18_or0;
  wire [0:0] u_csamul_pg_rca24_and5_18;
  wire [0:0] u_csamul_pg_rca24_fa5_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_18_or0;
  wire [0:0] u_csamul_pg_rca24_and6_18;
  wire [0:0] u_csamul_pg_rca24_fa6_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_18_or0;
  wire [0:0] u_csamul_pg_rca24_and7_18;
  wire [0:0] u_csamul_pg_rca24_fa7_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_18_or0;
  wire [0:0] u_csamul_pg_rca24_and8_18;
  wire [0:0] u_csamul_pg_rca24_fa8_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_18_or0;
  wire [0:0] u_csamul_pg_rca24_and9_18;
  wire [0:0] u_csamul_pg_rca24_fa9_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_18_or0;
  wire [0:0] u_csamul_pg_rca24_and10_18;
  wire [0:0] u_csamul_pg_rca24_fa10_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_18_or0;
  wire [0:0] u_csamul_pg_rca24_and11_18;
  wire [0:0] u_csamul_pg_rca24_fa11_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_18_or0;
  wire [0:0] u_csamul_pg_rca24_and12_18;
  wire [0:0] u_csamul_pg_rca24_fa12_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_18_or0;
  wire [0:0] u_csamul_pg_rca24_and13_18;
  wire [0:0] u_csamul_pg_rca24_fa13_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_18_or0;
  wire [0:0] u_csamul_pg_rca24_and14_18;
  wire [0:0] u_csamul_pg_rca24_fa14_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_18_or0;
  wire [0:0] u_csamul_pg_rca24_and15_18;
  wire [0:0] u_csamul_pg_rca24_fa15_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_18_or0;
  wire [0:0] u_csamul_pg_rca24_and16_18;
  wire [0:0] u_csamul_pg_rca24_fa16_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_18_or0;
  wire [0:0] u_csamul_pg_rca24_and17_18;
  wire [0:0] u_csamul_pg_rca24_fa17_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_18_or0;
  wire [0:0] u_csamul_pg_rca24_and18_18;
  wire [0:0] u_csamul_pg_rca24_fa18_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_18_or0;
  wire [0:0] u_csamul_pg_rca24_and19_18;
  wire [0:0] u_csamul_pg_rca24_fa19_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_18_or0;
  wire [0:0] u_csamul_pg_rca24_and20_18;
  wire [0:0] u_csamul_pg_rca24_fa20_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_18_or0;
  wire [0:0] u_csamul_pg_rca24_and21_18;
  wire [0:0] u_csamul_pg_rca24_fa21_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_18_or0;
  wire [0:0] u_csamul_pg_rca24_and22_18;
  wire [0:0] u_csamul_pg_rca24_fa22_18_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_18_or0;
  wire [0:0] u_csamul_pg_rca24_and23_18;
  wire [0:0] u_csamul_pg_rca24_and0_19;
  wire [0:0] u_csamul_pg_rca24_fa0_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_19_or0;
  wire [0:0] u_csamul_pg_rca24_and1_19;
  wire [0:0] u_csamul_pg_rca24_fa1_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_19_or0;
  wire [0:0] u_csamul_pg_rca24_and2_19;
  wire [0:0] u_csamul_pg_rca24_fa2_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_19_or0;
  wire [0:0] u_csamul_pg_rca24_and3_19;
  wire [0:0] u_csamul_pg_rca24_fa3_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_19_or0;
  wire [0:0] u_csamul_pg_rca24_and4_19;
  wire [0:0] u_csamul_pg_rca24_fa4_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_19_or0;
  wire [0:0] u_csamul_pg_rca24_and5_19;
  wire [0:0] u_csamul_pg_rca24_fa5_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_19_or0;
  wire [0:0] u_csamul_pg_rca24_and6_19;
  wire [0:0] u_csamul_pg_rca24_fa6_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_19_or0;
  wire [0:0] u_csamul_pg_rca24_and7_19;
  wire [0:0] u_csamul_pg_rca24_fa7_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_19_or0;
  wire [0:0] u_csamul_pg_rca24_and8_19;
  wire [0:0] u_csamul_pg_rca24_fa8_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_19_or0;
  wire [0:0] u_csamul_pg_rca24_and9_19;
  wire [0:0] u_csamul_pg_rca24_fa9_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_19_or0;
  wire [0:0] u_csamul_pg_rca24_and10_19;
  wire [0:0] u_csamul_pg_rca24_fa10_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_19_or0;
  wire [0:0] u_csamul_pg_rca24_and11_19;
  wire [0:0] u_csamul_pg_rca24_fa11_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_19_or0;
  wire [0:0] u_csamul_pg_rca24_and12_19;
  wire [0:0] u_csamul_pg_rca24_fa12_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_19_or0;
  wire [0:0] u_csamul_pg_rca24_and13_19;
  wire [0:0] u_csamul_pg_rca24_fa13_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_19_or0;
  wire [0:0] u_csamul_pg_rca24_and14_19;
  wire [0:0] u_csamul_pg_rca24_fa14_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_19_or0;
  wire [0:0] u_csamul_pg_rca24_and15_19;
  wire [0:0] u_csamul_pg_rca24_fa15_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_19_or0;
  wire [0:0] u_csamul_pg_rca24_and16_19;
  wire [0:0] u_csamul_pg_rca24_fa16_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_19_or0;
  wire [0:0] u_csamul_pg_rca24_and17_19;
  wire [0:0] u_csamul_pg_rca24_fa17_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_19_or0;
  wire [0:0] u_csamul_pg_rca24_and18_19;
  wire [0:0] u_csamul_pg_rca24_fa18_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_19_or0;
  wire [0:0] u_csamul_pg_rca24_and19_19;
  wire [0:0] u_csamul_pg_rca24_fa19_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_19_or0;
  wire [0:0] u_csamul_pg_rca24_and20_19;
  wire [0:0] u_csamul_pg_rca24_fa20_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_19_or0;
  wire [0:0] u_csamul_pg_rca24_and21_19;
  wire [0:0] u_csamul_pg_rca24_fa21_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_19_or0;
  wire [0:0] u_csamul_pg_rca24_and22_19;
  wire [0:0] u_csamul_pg_rca24_fa22_19_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_19_or0;
  wire [0:0] u_csamul_pg_rca24_and23_19;
  wire [0:0] u_csamul_pg_rca24_and0_20;
  wire [0:0] u_csamul_pg_rca24_fa0_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_20_or0;
  wire [0:0] u_csamul_pg_rca24_and1_20;
  wire [0:0] u_csamul_pg_rca24_fa1_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_20_or0;
  wire [0:0] u_csamul_pg_rca24_and2_20;
  wire [0:0] u_csamul_pg_rca24_fa2_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_20_or0;
  wire [0:0] u_csamul_pg_rca24_and3_20;
  wire [0:0] u_csamul_pg_rca24_fa3_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_20_or0;
  wire [0:0] u_csamul_pg_rca24_and4_20;
  wire [0:0] u_csamul_pg_rca24_fa4_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_20_or0;
  wire [0:0] u_csamul_pg_rca24_and5_20;
  wire [0:0] u_csamul_pg_rca24_fa5_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_20_or0;
  wire [0:0] u_csamul_pg_rca24_and6_20;
  wire [0:0] u_csamul_pg_rca24_fa6_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_20_or0;
  wire [0:0] u_csamul_pg_rca24_and7_20;
  wire [0:0] u_csamul_pg_rca24_fa7_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_20_or0;
  wire [0:0] u_csamul_pg_rca24_and8_20;
  wire [0:0] u_csamul_pg_rca24_fa8_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_20_or0;
  wire [0:0] u_csamul_pg_rca24_and9_20;
  wire [0:0] u_csamul_pg_rca24_fa9_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_20_or0;
  wire [0:0] u_csamul_pg_rca24_and10_20;
  wire [0:0] u_csamul_pg_rca24_fa10_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_20_or0;
  wire [0:0] u_csamul_pg_rca24_and11_20;
  wire [0:0] u_csamul_pg_rca24_fa11_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_20_or0;
  wire [0:0] u_csamul_pg_rca24_and12_20;
  wire [0:0] u_csamul_pg_rca24_fa12_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_20_or0;
  wire [0:0] u_csamul_pg_rca24_and13_20;
  wire [0:0] u_csamul_pg_rca24_fa13_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_20_or0;
  wire [0:0] u_csamul_pg_rca24_and14_20;
  wire [0:0] u_csamul_pg_rca24_fa14_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_20_or0;
  wire [0:0] u_csamul_pg_rca24_and15_20;
  wire [0:0] u_csamul_pg_rca24_fa15_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_20_or0;
  wire [0:0] u_csamul_pg_rca24_and16_20;
  wire [0:0] u_csamul_pg_rca24_fa16_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_20_or0;
  wire [0:0] u_csamul_pg_rca24_and17_20;
  wire [0:0] u_csamul_pg_rca24_fa17_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_20_or0;
  wire [0:0] u_csamul_pg_rca24_and18_20;
  wire [0:0] u_csamul_pg_rca24_fa18_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_20_or0;
  wire [0:0] u_csamul_pg_rca24_and19_20;
  wire [0:0] u_csamul_pg_rca24_fa19_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_20_or0;
  wire [0:0] u_csamul_pg_rca24_and20_20;
  wire [0:0] u_csamul_pg_rca24_fa20_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_20_or0;
  wire [0:0] u_csamul_pg_rca24_and21_20;
  wire [0:0] u_csamul_pg_rca24_fa21_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_20_or0;
  wire [0:0] u_csamul_pg_rca24_and22_20;
  wire [0:0] u_csamul_pg_rca24_fa22_20_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_20_or0;
  wire [0:0] u_csamul_pg_rca24_and23_20;
  wire [0:0] u_csamul_pg_rca24_and0_21;
  wire [0:0] u_csamul_pg_rca24_fa0_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_21_or0;
  wire [0:0] u_csamul_pg_rca24_and1_21;
  wire [0:0] u_csamul_pg_rca24_fa1_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_21_or0;
  wire [0:0] u_csamul_pg_rca24_and2_21;
  wire [0:0] u_csamul_pg_rca24_fa2_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_21_or0;
  wire [0:0] u_csamul_pg_rca24_and3_21;
  wire [0:0] u_csamul_pg_rca24_fa3_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_21_or0;
  wire [0:0] u_csamul_pg_rca24_and4_21;
  wire [0:0] u_csamul_pg_rca24_fa4_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_21_or0;
  wire [0:0] u_csamul_pg_rca24_and5_21;
  wire [0:0] u_csamul_pg_rca24_fa5_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_21_or0;
  wire [0:0] u_csamul_pg_rca24_and6_21;
  wire [0:0] u_csamul_pg_rca24_fa6_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_21_or0;
  wire [0:0] u_csamul_pg_rca24_and7_21;
  wire [0:0] u_csamul_pg_rca24_fa7_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_21_or0;
  wire [0:0] u_csamul_pg_rca24_and8_21;
  wire [0:0] u_csamul_pg_rca24_fa8_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_21_or0;
  wire [0:0] u_csamul_pg_rca24_and9_21;
  wire [0:0] u_csamul_pg_rca24_fa9_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_21_or0;
  wire [0:0] u_csamul_pg_rca24_and10_21;
  wire [0:0] u_csamul_pg_rca24_fa10_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_21_or0;
  wire [0:0] u_csamul_pg_rca24_and11_21;
  wire [0:0] u_csamul_pg_rca24_fa11_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_21_or0;
  wire [0:0] u_csamul_pg_rca24_and12_21;
  wire [0:0] u_csamul_pg_rca24_fa12_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_21_or0;
  wire [0:0] u_csamul_pg_rca24_and13_21;
  wire [0:0] u_csamul_pg_rca24_fa13_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_21_or0;
  wire [0:0] u_csamul_pg_rca24_and14_21;
  wire [0:0] u_csamul_pg_rca24_fa14_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_21_or0;
  wire [0:0] u_csamul_pg_rca24_and15_21;
  wire [0:0] u_csamul_pg_rca24_fa15_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_21_or0;
  wire [0:0] u_csamul_pg_rca24_and16_21;
  wire [0:0] u_csamul_pg_rca24_fa16_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_21_or0;
  wire [0:0] u_csamul_pg_rca24_and17_21;
  wire [0:0] u_csamul_pg_rca24_fa17_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_21_or0;
  wire [0:0] u_csamul_pg_rca24_and18_21;
  wire [0:0] u_csamul_pg_rca24_fa18_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_21_or0;
  wire [0:0] u_csamul_pg_rca24_and19_21;
  wire [0:0] u_csamul_pg_rca24_fa19_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_21_or0;
  wire [0:0] u_csamul_pg_rca24_and20_21;
  wire [0:0] u_csamul_pg_rca24_fa20_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_21_or0;
  wire [0:0] u_csamul_pg_rca24_and21_21;
  wire [0:0] u_csamul_pg_rca24_fa21_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_21_or0;
  wire [0:0] u_csamul_pg_rca24_and22_21;
  wire [0:0] u_csamul_pg_rca24_fa22_21_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_21_or0;
  wire [0:0] u_csamul_pg_rca24_and23_21;
  wire [0:0] u_csamul_pg_rca24_and0_22;
  wire [0:0] u_csamul_pg_rca24_fa0_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_22_or0;
  wire [0:0] u_csamul_pg_rca24_and1_22;
  wire [0:0] u_csamul_pg_rca24_fa1_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_22_or0;
  wire [0:0] u_csamul_pg_rca24_and2_22;
  wire [0:0] u_csamul_pg_rca24_fa2_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_22_or0;
  wire [0:0] u_csamul_pg_rca24_and3_22;
  wire [0:0] u_csamul_pg_rca24_fa3_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_22_or0;
  wire [0:0] u_csamul_pg_rca24_and4_22;
  wire [0:0] u_csamul_pg_rca24_fa4_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_22_or0;
  wire [0:0] u_csamul_pg_rca24_and5_22;
  wire [0:0] u_csamul_pg_rca24_fa5_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_22_or0;
  wire [0:0] u_csamul_pg_rca24_and6_22;
  wire [0:0] u_csamul_pg_rca24_fa6_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_22_or0;
  wire [0:0] u_csamul_pg_rca24_and7_22;
  wire [0:0] u_csamul_pg_rca24_fa7_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_22_or0;
  wire [0:0] u_csamul_pg_rca24_and8_22;
  wire [0:0] u_csamul_pg_rca24_fa8_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_22_or0;
  wire [0:0] u_csamul_pg_rca24_and9_22;
  wire [0:0] u_csamul_pg_rca24_fa9_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_22_or0;
  wire [0:0] u_csamul_pg_rca24_and10_22;
  wire [0:0] u_csamul_pg_rca24_fa10_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_22_or0;
  wire [0:0] u_csamul_pg_rca24_and11_22;
  wire [0:0] u_csamul_pg_rca24_fa11_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_22_or0;
  wire [0:0] u_csamul_pg_rca24_and12_22;
  wire [0:0] u_csamul_pg_rca24_fa12_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_22_or0;
  wire [0:0] u_csamul_pg_rca24_and13_22;
  wire [0:0] u_csamul_pg_rca24_fa13_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_22_or0;
  wire [0:0] u_csamul_pg_rca24_and14_22;
  wire [0:0] u_csamul_pg_rca24_fa14_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_22_or0;
  wire [0:0] u_csamul_pg_rca24_and15_22;
  wire [0:0] u_csamul_pg_rca24_fa15_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_22_or0;
  wire [0:0] u_csamul_pg_rca24_and16_22;
  wire [0:0] u_csamul_pg_rca24_fa16_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_22_or0;
  wire [0:0] u_csamul_pg_rca24_and17_22;
  wire [0:0] u_csamul_pg_rca24_fa17_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_22_or0;
  wire [0:0] u_csamul_pg_rca24_and18_22;
  wire [0:0] u_csamul_pg_rca24_fa18_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_22_or0;
  wire [0:0] u_csamul_pg_rca24_and19_22;
  wire [0:0] u_csamul_pg_rca24_fa19_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_22_or0;
  wire [0:0] u_csamul_pg_rca24_and20_22;
  wire [0:0] u_csamul_pg_rca24_fa20_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_22_or0;
  wire [0:0] u_csamul_pg_rca24_and21_22;
  wire [0:0] u_csamul_pg_rca24_fa21_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_22_or0;
  wire [0:0] u_csamul_pg_rca24_and22_22;
  wire [0:0] u_csamul_pg_rca24_fa22_22_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_22_or0;
  wire [0:0] u_csamul_pg_rca24_and23_22;
  wire [0:0] u_csamul_pg_rca24_and0_23;
  wire [0:0] u_csamul_pg_rca24_fa0_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa0_23_or0;
  wire [0:0] u_csamul_pg_rca24_and1_23;
  wire [0:0] u_csamul_pg_rca24_fa1_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa1_23_or0;
  wire [0:0] u_csamul_pg_rca24_and2_23;
  wire [0:0] u_csamul_pg_rca24_fa2_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa2_23_or0;
  wire [0:0] u_csamul_pg_rca24_and3_23;
  wire [0:0] u_csamul_pg_rca24_fa3_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa3_23_or0;
  wire [0:0] u_csamul_pg_rca24_and4_23;
  wire [0:0] u_csamul_pg_rca24_fa4_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa4_23_or0;
  wire [0:0] u_csamul_pg_rca24_and5_23;
  wire [0:0] u_csamul_pg_rca24_fa5_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa5_23_or0;
  wire [0:0] u_csamul_pg_rca24_and6_23;
  wire [0:0] u_csamul_pg_rca24_fa6_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa6_23_or0;
  wire [0:0] u_csamul_pg_rca24_and7_23;
  wire [0:0] u_csamul_pg_rca24_fa7_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa7_23_or0;
  wire [0:0] u_csamul_pg_rca24_and8_23;
  wire [0:0] u_csamul_pg_rca24_fa8_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa8_23_or0;
  wire [0:0] u_csamul_pg_rca24_and9_23;
  wire [0:0] u_csamul_pg_rca24_fa9_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa9_23_or0;
  wire [0:0] u_csamul_pg_rca24_and10_23;
  wire [0:0] u_csamul_pg_rca24_fa10_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa10_23_or0;
  wire [0:0] u_csamul_pg_rca24_and11_23;
  wire [0:0] u_csamul_pg_rca24_fa11_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa11_23_or0;
  wire [0:0] u_csamul_pg_rca24_and12_23;
  wire [0:0] u_csamul_pg_rca24_fa12_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa12_23_or0;
  wire [0:0] u_csamul_pg_rca24_and13_23;
  wire [0:0] u_csamul_pg_rca24_fa13_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa13_23_or0;
  wire [0:0] u_csamul_pg_rca24_and14_23;
  wire [0:0] u_csamul_pg_rca24_fa14_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa14_23_or0;
  wire [0:0] u_csamul_pg_rca24_and15_23;
  wire [0:0] u_csamul_pg_rca24_fa15_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa15_23_or0;
  wire [0:0] u_csamul_pg_rca24_and16_23;
  wire [0:0] u_csamul_pg_rca24_fa16_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa16_23_or0;
  wire [0:0] u_csamul_pg_rca24_and17_23;
  wire [0:0] u_csamul_pg_rca24_fa17_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa17_23_or0;
  wire [0:0] u_csamul_pg_rca24_and18_23;
  wire [0:0] u_csamul_pg_rca24_fa18_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa18_23_or0;
  wire [0:0] u_csamul_pg_rca24_and19_23;
  wire [0:0] u_csamul_pg_rca24_fa19_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa19_23_or0;
  wire [0:0] u_csamul_pg_rca24_and20_23;
  wire [0:0] u_csamul_pg_rca24_fa20_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa20_23_or0;
  wire [0:0] u_csamul_pg_rca24_and21_23;
  wire [0:0] u_csamul_pg_rca24_fa21_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa21_23_or0;
  wire [0:0] u_csamul_pg_rca24_and22_23;
  wire [0:0] u_csamul_pg_rca24_fa22_23_xor1;
  wire [0:0] u_csamul_pg_rca24_fa22_23_or0;
  wire [0:0] u_csamul_pg_rca24_and23_23;
  wire [23:0] u_csamul_pg_rca24_u_pg_rca24_a;
  wire [23:0] u_csamul_pg_rca24_u_pg_rca24_b;
  wire [24:0] u_csamul_pg_rca24_u_pg_rca24_out;

  and_gate and_gate_u_csamul_pg_rca24_and0_0(.a(a[0]), .b(b[0]), .out(u_csamul_pg_rca24_and0_0));
  and_gate and_gate_u_csamul_pg_rca24_and1_0(.a(a[1]), .b(b[0]), .out(u_csamul_pg_rca24_and1_0));
  and_gate and_gate_u_csamul_pg_rca24_and2_0(.a(a[2]), .b(b[0]), .out(u_csamul_pg_rca24_and2_0));
  and_gate and_gate_u_csamul_pg_rca24_and3_0(.a(a[3]), .b(b[0]), .out(u_csamul_pg_rca24_and3_0));
  and_gate and_gate_u_csamul_pg_rca24_and4_0(.a(a[4]), .b(b[0]), .out(u_csamul_pg_rca24_and4_0));
  and_gate and_gate_u_csamul_pg_rca24_and5_0(.a(a[5]), .b(b[0]), .out(u_csamul_pg_rca24_and5_0));
  and_gate and_gate_u_csamul_pg_rca24_and6_0(.a(a[6]), .b(b[0]), .out(u_csamul_pg_rca24_and6_0));
  and_gate and_gate_u_csamul_pg_rca24_and7_0(.a(a[7]), .b(b[0]), .out(u_csamul_pg_rca24_and7_0));
  and_gate and_gate_u_csamul_pg_rca24_and8_0(.a(a[8]), .b(b[0]), .out(u_csamul_pg_rca24_and8_0));
  and_gate and_gate_u_csamul_pg_rca24_and9_0(.a(a[9]), .b(b[0]), .out(u_csamul_pg_rca24_and9_0));
  and_gate and_gate_u_csamul_pg_rca24_and10_0(.a(a[10]), .b(b[0]), .out(u_csamul_pg_rca24_and10_0));
  and_gate and_gate_u_csamul_pg_rca24_and11_0(.a(a[11]), .b(b[0]), .out(u_csamul_pg_rca24_and11_0));
  and_gate and_gate_u_csamul_pg_rca24_and12_0(.a(a[12]), .b(b[0]), .out(u_csamul_pg_rca24_and12_0));
  and_gate and_gate_u_csamul_pg_rca24_and13_0(.a(a[13]), .b(b[0]), .out(u_csamul_pg_rca24_and13_0));
  and_gate and_gate_u_csamul_pg_rca24_and14_0(.a(a[14]), .b(b[0]), .out(u_csamul_pg_rca24_and14_0));
  and_gate and_gate_u_csamul_pg_rca24_and15_0(.a(a[15]), .b(b[0]), .out(u_csamul_pg_rca24_and15_0));
  and_gate and_gate_u_csamul_pg_rca24_and16_0(.a(a[16]), .b(b[0]), .out(u_csamul_pg_rca24_and16_0));
  and_gate and_gate_u_csamul_pg_rca24_and17_0(.a(a[17]), .b(b[0]), .out(u_csamul_pg_rca24_and17_0));
  and_gate and_gate_u_csamul_pg_rca24_and18_0(.a(a[18]), .b(b[0]), .out(u_csamul_pg_rca24_and18_0));
  and_gate and_gate_u_csamul_pg_rca24_and19_0(.a(a[19]), .b(b[0]), .out(u_csamul_pg_rca24_and19_0));
  and_gate and_gate_u_csamul_pg_rca24_and20_0(.a(a[20]), .b(b[0]), .out(u_csamul_pg_rca24_and20_0));
  and_gate and_gate_u_csamul_pg_rca24_and21_0(.a(a[21]), .b(b[0]), .out(u_csamul_pg_rca24_and21_0));
  and_gate and_gate_u_csamul_pg_rca24_and22_0(.a(a[22]), .b(b[0]), .out(u_csamul_pg_rca24_and22_0));
  and_gate and_gate_u_csamul_pg_rca24_and23_0(.a(a[23]), .b(b[0]), .out(u_csamul_pg_rca24_and23_0));
  and_gate and_gate_u_csamul_pg_rca24_and0_1(.a(a[0]), .b(b[1]), .out(u_csamul_pg_rca24_and0_1));
  ha ha_u_csamul_pg_rca24_ha0_1_out(.a(u_csamul_pg_rca24_and0_1[0]), .b(u_csamul_pg_rca24_and1_0[0]), .ha_xor0(u_csamul_pg_rca24_ha0_1_xor0), .ha_and0(u_csamul_pg_rca24_ha0_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and1_1(.a(a[1]), .b(b[1]), .out(u_csamul_pg_rca24_and1_1));
  ha ha_u_csamul_pg_rca24_ha1_1_out(.a(u_csamul_pg_rca24_and1_1[0]), .b(u_csamul_pg_rca24_and2_0[0]), .ha_xor0(u_csamul_pg_rca24_ha1_1_xor0), .ha_and0(u_csamul_pg_rca24_ha1_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and2_1(.a(a[2]), .b(b[1]), .out(u_csamul_pg_rca24_and2_1));
  ha ha_u_csamul_pg_rca24_ha2_1_out(.a(u_csamul_pg_rca24_and2_1[0]), .b(u_csamul_pg_rca24_and3_0[0]), .ha_xor0(u_csamul_pg_rca24_ha2_1_xor0), .ha_and0(u_csamul_pg_rca24_ha2_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and3_1(.a(a[3]), .b(b[1]), .out(u_csamul_pg_rca24_and3_1));
  ha ha_u_csamul_pg_rca24_ha3_1_out(.a(u_csamul_pg_rca24_and3_1[0]), .b(u_csamul_pg_rca24_and4_0[0]), .ha_xor0(u_csamul_pg_rca24_ha3_1_xor0), .ha_and0(u_csamul_pg_rca24_ha3_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and4_1(.a(a[4]), .b(b[1]), .out(u_csamul_pg_rca24_and4_1));
  ha ha_u_csamul_pg_rca24_ha4_1_out(.a(u_csamul_pg_rca24_and4_1[0]), .b(u_csamul_pg_rca24_and5_0[0]), .ha_xor0(u_csamul_pg_rca24_ha4_1_xor0), .ha_and0(u_csamul_pg_rca24_ha4_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and5_1(.a(a[5]), .b(b[1]), .out(u_csamul_pg_rca24_and5_1));
  ha ha_u_csamul_pg_rca24_ha5_1_out(.a(u_csamul_pg_rca24_and5_1[0]), .b(u_csamul_pg_rca24_and6_0[0]), .ha_xor0(u_csamul_pg_rca24_ha5_1_xor0), .ha_and0(u_csamul_pg_rca24_ha5_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and6_1(.a(a[6]), .b(b[1]), .out(u_csamul_pg_rca24_and6_1));
  ha ha_u_csamul_pg_rca24_ha6_1_out(.a(u_csamul_pg_rca24_and6_1[0]), .b(u_csamul_pg_rca24_and7_0[0]), .ha_xor0(u_csamul_pg_rca24_ha6_1_xor0), .ha_and0(u_csamul_pg_rca24_ha6_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and7_1(.a(a[7]), .b(b[1]), .out(u_csamul_pg_rca24_and7_1));
  ha ha_u_csamul_pg_rca24_ha7_1_out(.a(u_csamul_pg_rca24_and7_1[0]), .b(u_csamul_pg_rca24_and8_0[0]), .ha_xor0(u_csamul_pg_rca24_ha7_1_xor0), .ha_and0(u_csamul_pg_rca24_ha7_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and8_1(.a(a[8]), .b(b[1]), .out(u_csamul_pg_rca24_and8_1));
  ha ha_u_csamul_pg_rca24_ha8_1_out(.a(u_csamul_pg_rca24_and8_1[0]), .b(u_csamul_pg_rca24_and9_0[0]), .ha_xor0(u_csamul_pg_rca24_ha8_1_xor0), .ha_and0(u_csamul_pg_rca24_ha8_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and9_1(.a(a[9]), .b(b[1]), .out(u_csamul_pg_rca24_and9_1));
  ha ha_u_csamul_pg_rca24_ha9_1_out(.a(u_csamul_pg_rca24_and9_1[0]), .b(u_csamul_pg_rca24_and10_0[0]), .ha_xor0(u_csamul_pg_rca24_ha9_1_xor0), .ha_and0(u_csamul_pg_rca24_ha9_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and10_1(.a(a[10]), .b(b[1]), .out(u_csamul_pg_rca24_and10_1));
  ha ha_u_csamul_pg_rca24_ha10_1_out(.a(u_csamul_pg_rca24_and10_1[0]), .b(u_csamul_pg_rca24_and11_0[0]), .ha_xor0(u_csamul_pg_rca24_ha10_1_xor0), .ha_and0(u_csamul_pg_rca24_ha10_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and11_1(.a(a[11]), .b(b[1]), .out(u_csamul_pg_rca24_and11_1));
  ha ha_u_csamul_pg_rca24_ha11_1_out(.a(u_csamul_pg_rca24_and11_1[0]), .b(u_csamul_pg_rca24_and12_0[0]), .ha_xor0(u_csamul_pg_rca24_ha11_1_xor0), .ha_and0(u_csamul_pg_rca24_ha11_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and12_1(.a(a[12]), .b(b[1]), .out(u_csamul_pg_rca24_and12_1));
  ha ha_u_csamul_pg_rca24_ha12_1_out(.a(u_csamul_pg_rca24_and12_1[0]), .b(u_csamul_pg_rca24_and13_0[0]), .ha_xor0(u_csamul_pg_rca24_ha12_1_xor0), .ha_and0(u_csamul_pg_rca24_ha12_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and13_1(.a(a[13]), .b(b[1]), .out(u_csamul_pg_rca24_and13_1));
  ha ha_u_csamul_pg_rca24_ha13_1_out(.a(u_csamul_pg_rca24_and13_1[0]), .b(u_csamul_pg_rca24_and14_0[0]), .ha_xor0(u_csamul_pg_rca24_ha13_1_xor0), .ha_and0(u_csamul_pg_rca24_ha13_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and14_1(.a(a[14]), .b(b[1]), .out(u_csamul_pg_rca24_and14_1));
  ha ha_u_csamul_pg_rca24_ha14_1_out(.a(u_csamul_pg_rca24_and14_1[0]), .b(u_csamul_pg_rca24_and15_0[0]), .ha_xor0(u_csamul_pg_rca24_ha14_1_xor0), .ha_and0(u_csamul_pg_rca24_ha14_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and15_1(.a(a[15]), .b(b[1]), .out(u_csamul_pg_rca24_and15_1));
  ha ha_u_csamul_pg_rca24_ha15_1_out(.a(u_csamul_pg_rca24_and15_1[0]), .b(u_csamul_pg_rca24_and16_0[0]), .ha_xor0(u_csamul_pg_rca24_ha15_1_xor0), .ha_and0(u_csamul_pg_rca24_ha15_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and16_1(.a(a[16]), .b(b[1]), .out(u_csamul_pg_rca24_and16_1));
  ha ha_u_csamul_pg_rca24_ha16_1_out(.a(u_csamul_pg_rca24_and16_1[0]), .b(u_csamul_pg_rca24_and17_0[0]), .ha_xor0(u_csamul_pg_rca24_ha16_1_xor0), .ha_and0(u_csamul_pg_rca24_ha16_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and17_1(.a(a[17]), .b(b[1]), .out(u_csamul_pg_rca24_and17_1));
  ha ha_u_csamul_pg_rca24_ha17_1_out(.a(u_csamul_pg_rca24_and17_1[0]), .b(u_csamul_pg_rca24_and18_0[0]), .ha_xor0(u_csamul_pg_rca24_ha17_1_xor0), .ha_and0(u_csamul_pg_rca24_ha17_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and18_1(.a(a[18]), .b(b[1]), .out(u_csamul_pg_rca24_and18_1));
  ha ha_u_csamul_pg_rca24_ha18_1_out(.a(u_csamul_pg_rca24_and18_1[0]), .b(u_csamul_pg_rca24_and19_0[0]), .ha_xor0(u_csamul_pg_rca24_ha18_1_xor0), .ha_and0(u_csamul_pg_rca24_ha18_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and19_1(.a(a[19]), .b(b[1]), .out(u_csamul_pg_rca24_and19_1));
  ha ha_u_csamul_pg_rca24_ha19_1_out(.a(u_csamul_pg_rca24_and19_1[0]), .b(u_csamul_pg_rca24_and20_0[0]), .ha_xor0(u_csamul_pg_rca24_ha19_1_xor0), .ha_and0(u_csamul_pg_rca24_ha19_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and20_1(.a(a[20]), .b(b[1]), .out(u_csamul_pg_rca24_and20_1));
  ha ha_u_csamul_pg_rca24_ha20_1_out(.a(u_csamul_pg_rca24_and20_1[0]), .b(u_csamul_pg_rca24_and21_0[0]), .ha_xor0(u_csamul_pg_rca24_ha20_1_xor0), .ha_and0(u_csamul_pg_rca24_ha20_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and21_1(.a(a[21]), .b(b[1]), .out(u_csamul_pg_rca24_and21_1));
  ha ha_u_csamul_pg_rca24_ha21_1_out(.a(u_csamul_pg_rca24_and21_1[0]), .b(u_csamul_pg_rca24_and22_0[0]), .ha_xor0(u_csamul_pg_rca24_ha21_1_xor0), .ha_and0(u_csamul_pg_rca24_ha21_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and22_1(.a(a[22]), .b(b[1]), .out(u_csamul_pg_rca24_and22_1));
  ha ha_u_csamul_pg_rca24_ha22_1_out(.a(u_csamul_pg_rca24_and22_1[0]), .b(u_csamul_pg_rca24_and23_0[0]), .ha_xor0(u_csamul_pg_rca24_ha22_1_xor0), .ha_and0(u_csamul_pg_rca24_ha22_1_and0));
  and_gate and_gate_u_csamul_pg_rca24_and23_1(.a(a[23]), .b(b[1]), .out(u_csamul_pg_rca24_and23_1));
  and_gate and_gate_u_csamul_pg_rca24_and0_2(.a(a[0]), .b(b[2]), .out(u_csamul_pg_rca24_and0_2));
  fa fa_u_csamul_pg_rca24_fa0_2_out(.a(u_csamul_pg_rca24_and0_2[0]), .b(u_csamul_pg_rca24_ha1_1_xor0[0]), .cin(u_csamul_pg_rca24_ha0_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_2_xor1), .fa_or0(u_csamul_pg_rca24_fa0_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_2(.a(a[1]), .b(b[2]), .out(u_csamul_pg_rca24_and1_2));
  fa fa_u_csamul_pg_rca24_fa1_2_out(.a(u_csamul_pg_rca24_and1_2[0]), .b(u_csamul_pg_rca24_ha2_1_xor0[0]), .cin(u_csamul_pg_rca24_ha1_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_2_xor1), .fa_or0(u_csamul_pg_rca24_fa1_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_2(.a(a[2]), .b(b[2]), .out(u_csamul_pg_rca24_and2_2));
  fa fa_u_csamul_pg_rca24_fa2_2_out(.a(u_csamul_pg_rca24_and2_2[0]), .b(u_csamul_pg_rca24_ha3_1_xor0[0]), .cin(u_csamul_pg_rca24_ha2_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_2_xor1), .fa_or0(u_csamul_pg_rca24_fa2_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_2(.a(a[3]), .b(b[2]), .out(u_csamul_pg_rca24_and3_2));
  fa fa_u_csamul_pg_rca24_fa3_2_out(.a(u_csamul_pg_rca24_and3_2[0]), .b(u_csamul_pg_rca24_ha4_1_xor0[0]), .cin(u_csamul_pg_rca24_ha3_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_2_xor1), .fa_or0(u_csamul_pg_rca24_fa3_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_2(.a(a[4]), .b(b[2]), .out(u_csamul_pg_rca24_and4_2));
  fa fa_u_csamul_pg_rca24_fa4_2_out(.a(u_csamul_pg_rca24_and4_2[0]), .b(u_csamul_pg_rca24_ha5_1_xor0[0]), .cin(u_csamul_pg_rca24_ha4_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_2_xor1), .fa_or0(u_csamul_pg_rca24_fa4_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_2(.a(a[5]), .b(b[2]), .out(u_csamul_pg_rca24_and5_2));
  fa fa_u_csamul_pg_rca24_fa5_2_out(.a(u_csamul_pg_rca24_and5_2[0]), .b(u_csamul_pg_rca24_ha6_1_xor0[0]), .cin(u_csamul_pg_rca24_ha5_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_2_xor1), .fa_or0(u_csamul_pg_rca24_fa5_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_2(.a(a[6]), .b(b[2]), .out(u_csamul_pg_rca24_and6_2));
  fa fa_u_csamul_pg_rca24_fa6_2_out(.a(u_csamul_pg_rca24_and6_2[0]), .b(u_csamul_pg_rca24_ha7_1_xor0[0]), .cin(u_csamul_pg_rca24_ha6_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_2_xor1), .fa_or0(u_csamul_pg_rca24_fa6_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_2(.a(a[7]), .b(b[2]), .out(u_csamul_pg_rca24_and7_2));
  fa fa_u_csamul_pg_rca24_fa7_2_out(.a(u_csamul_pg_rca24_and7_2[0]), .b(u_csamul_pg_rca24_ha8_1_xor0[0]), .cin(u_csamul_pg_rca24_ha7_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_2_xor1), .fa_or0(u_csamul_pg_rca24_fa7_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_2(.a(a[8]), .b(b[2]), .out(u_csamul_pg_rca24_and8_2));
  fa fa_u_csamul_pg_rca24_fa8_2_out(.a(u_csamul_pg_rca24_and8_2[0]), .b(u_csamul_pg_rca24_ha9_1_xor0[0]), .cin(u_csamul_pg_rca24_ha8_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_2_xor1), .fa_or0(u_csamul_pg_rca24_fa8_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_2(.a(a[9]), .b(b[2]), .out(u_csamul_pg_rca24_and9_2));
  fa fa_u_csamul_pg_rca24_fa9_2_out(.a(u_csamul_pg_rca24_and9_2[0]), .b(u_csamul_pg_rca24_ha10_1_xor0[0]), .cin(u_csamul_pg_rca24_ha9_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_2_xor1), .fa_or0(u_csamul_pg_rca24_fa9_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_2(.a(a[10]), .b(b[2]), .out(u_csamul_pg_rca24_and10_2));
  fa fa_u_csamul_pg_rca24_fa10_2_out(.a(u_csamul_pg_rca24_and10_2[0]), .b(u_csamul_pg_rca24_ha11_1_xor0[0]), .cin(u_csamul_pg_rca24_ha10_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_2_xor1), .fa_or0(u_csamul_pg_rca24_fa10_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_2(.a(a[11]), .b(b[2]), .out(u_csamul_pg_rca24_and11_2));
  fa fa_u_csamul_pg_rca24_fa11_2_out(.a(u_csamul_pg_rca24_and11_2[0]), .b(u_csamul_pg_rca24_ha12_1_xor0[0]), .cin(u_csamul_pg_rca24_ha11_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_2_xor1), .fa_or0(u_csamul_pg_rca24_fa11_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_2(.a(a[12]), .b(b[2]), .out(u_csamul_pg_rca24_and12_2));
  fa fa_u_csamul_pg_rca24_fa12_2_out(.a(u_csamul_pg_rca24_and12_2[0]), .b(u_csamul_pg_rca24_ha13_1_xor0[0]), .cin(u_csamul_pg_rca24_ha12_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_2_xor1), .fa_or0(u_csamul_pg_rca24_fa12_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_2(.a(a[13]), .b(b[2]), .out(u_csamul_pg_rca24_and13_2));
  fa fa_u_csamul_pg_rca24_fa13_2_out(.a(u_csamul_pg_rca24_and13_2[0]), .b(u_csamul_pg_rca24_ha14_1_xor0[0]), .cin(u_csamul_pg_rca24_ha13_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_2_xor1), .fa_or0(u_csamul_pg_rca24_fa13_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_2(.a(a[14]), .b(b[2]), .out(u_csamul_pg_rca24_and14_2));
  fa fa_u_csamul_pg_rca24_fa14_2_out(.a(u_csamul_pg_rca24_and14_2[0]), .b(u_csamul_pg_rca24_ha15_1_xor0[0]), .cin(u_csamul_pg_rca24_ha14_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_2_xor1), .fa_or0(u_csamul_pg_rca24_fa14_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_2(.a(a[15]), .b(b[2]), .out(u_csamul_pg_rca24_and15_2));
  fa fa_u_csamul_pg_rca24_fa15_2_out(.a(u_csamul_pg_rca24_and15_2[0]), .b(u_csamul_pg_rca24_ha16_1_xor0[0]), .cin(u_csamul_pg_rca24_ha15_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_2_xor1), .fa_or0(u_csamul_pg_rca24_fa15_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_2(.a(a[16]), .b(b[2]), .out(u_csamul_pg_rca24_and16_2));
  fa fa_u_csamul_pg_rca24_fa16_2_out(.a(u_csamul_pg_rca24_and16_2[0]), .b(u_csamul_pg_rca24_ha17_1_xor0[0]), .cin(u_csamul_pg_rca24_ha16_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_2_xor1), .fa_or0(u_csamul_pg_rca24_fa16_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_2(.a(a[17]), .b(b[2]), .out(u_csamul_pg_rca24_and17_2));
  fa fa_u_csamul_pg_rca24_fa17_2_out(.a(u_csamul_pg_rca24_and17_2[0]), .b(u_csamul_pg_rca24_ha18_1_xor0[0]), .cin(u_csamul_pg_rca24_ha17_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_2_xor1), .fa_or0(u_csamul_pg_rca24_fa17_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_2(.a(a[18]), .b(b[2]), .out(u_csamul_pg_rca24_and18_2));
  fa fa_u_csamul_pg_rca24_fa18_2_out(.a(u_csamul_pg_rca24_and18_2[0]), .b(u_csamul_pg_rca24_ha19_1_xor0[0]), .cin(u_csamul_pg_rca24_ha18_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_2_xor1), .fa_or0(u_csamul_pg_rca24_fa18_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_2(.a(a[19]), .b(b[2]), .out(u_csamul_pg_rca24_and19_2));
  fa fa_u_csamul_pg_rca24_fa19_2_out(.a(u_csamul_pg_rca24_and19_2[0]), .b(u_csamul_pg_rca24_ha20_1_xor0[0]), .cin(u_csamul_pg_rca24_ha19_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_2_xor1), .fa_or0(u_csamul_pg_rca24_fa19_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_2(.a(a[20]), .b(b[2]), .out(u_csamul_pg_rca24_and20_2));
  fa fa_u_csamul_pg_rca24_fa20_2_out(.a(u_csamul_pg_rca24_and20_2[0]), .b(u_csamul_pg_rca24_ha21_1_xor0[0]), .cin(u_csamul_pg_rca24_ha20_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_2_xor1), .fa_or0(u_csamul_pg_rca24_fa20_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_2(.a(a[21]), .b(b[2]), .out(u_csamul_pg_rca24_and21_2));
  fa fa_u_csamul_pg_rca24_fa21_2_out(.a(u_csamul_pg_rca24_and21_2[0]), .b(u_csamul_pg_rca24_ha22_1_xor0[0]), .cin(u_csamul_pg_rca24_ha21_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_2_xor1), .fa_or0(u_csamul_pg_rca24_fa21_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_2(.a(a[22]), .b(b[2]), .out(u_csamul_pg_rca24_and22_2));
  fa fa_u_csamul_pg_rca24_fa22_2_out(.a(u_csamul_pg_rca24_and22_2[0]), .b(u_csamul_pg_rca24_and23_1[0]), .cin(u_csamul_pg_rca24_ha22_1_and0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_2_xor1), .fa_or0(u_csamul_pg_rca24_fa22_2_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_2(.a(a[23]), .b(b[2]), .out(u_csamul_pg_rca24_and23_2));
  and_gate and_gate_u_csamul_pg_rca24_and0_3(.a(a[0]), .b(b[3]), .out(u_csamul_pg_rca24_and0_3));
  fa fa_u_csamul_pg_rca24_fa0_3_out(.a(u_csamul_pg_rca24_and0_3[0]), .b(u_csamul_pg_rca24_fa1_2_xor1[0]), .cin(u_csamul_pg_rca24_fa0_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_3_xor1), .fa_or0(u_csamul_pg_rca24_fa0_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_3(.a(a[1]), .b(b[3]), .out(u_csamul_pg_rca24_and1_3));
  fa fa_u_csamul_pg_rca24_fa1_3_out(.a(u_csamul_pg_rca24_and1_3[0]), .b(u_csamul_pg_rca24_fa2_2_xor1[0]), .cin(u_csamul_pg_rca24_fa1_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_3_xor1), .fa_or0(u_csamul_pg_rca24_fa1_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_3(.a(a[2]), .b(b[3]), .out(u_csamul_pg_rca24_and2_3));
  fa fa_u_csamul_pg_rca24_fa2_3_out(.a(u_csamul_pg_rca24_and2_3[0]), .b(u_csamul_pg_rca24_fa3_2_xor1[0]), .cin(u_csamul_pg_rca24_fa2_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_3_xor1), .fa_or0(u_csamul_pg_rca24_fa2_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_3(.a(a[3]), .b(b[3]), .out(u_csamul_pg_rca24_and3_3));
  fa fa_u_csamul_pg_rca24_fa3_3_out(.a(u_csamul_pg_rca24_and3_3[0]), .b(u_csamul_pg_rca24_fa4_2_xor1[0]), .cin(u_csamul_pg_rca24_fa3_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_3_xor1), .fa_or0(u_csamul_pg_rca24_fa3_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_3(.a(a[4]), .b(b[3]), .out(u_csamul_pg_rca24_and4_3));
  fa fa_u_csamul_pg_rca24_fa4_3_out(.a(u_csamul_pg_rca24_and4_3[0]), .b(u_csamul_pg_rca24_fa5_2_xor1[0]), .cin(u_csamul_pg_rca24_fa4_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_3_xor1), .fa_or0(u_csamul_pg_rca24_fa4_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_3(.a(a[5]), .b(b[3]), .out(u_csamul_pg_rca24_and5_3));
  fa fa_u_csamul_pg_rca24_fa5_3_out(.a(u_csamul_pg_rca24_and5_3[0]), .b(u_csamul_pg_rca24_fa6_2_xor1[0]), .cin(u_csamul_pg_rca24_fa5_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_3_xor1), .fa_or0(u_csamul_pg_rca24_fa5_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_3(.a(a[6]), .b(b[3]), .out(u_csamul_pg_rca24_and6_3));
  fa fa_u_csamul_pg_rca24_fa6_3_out(.a(u_csamul_pg_rca24_and6_3[0]), .b(u_csamul_pg_rca24_fa7_2_xor1[0]), .cin(u_csamul_pg_rca24_fa6_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_3_xor1), .fa_or0(u_csamul_pg_rca24_fa6_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_3(.a(a[7]), .b(b[3]), .out(u_csamul_pg_rca24_and7_3));
  fa fa_u_csamul_pg_rca24_fa7_3_out(.a(u_csamul_pg_rca24_and7_3[0]), .b(u_csamul_pg_rca24_fa8_2_xor1[0]), .cin(u_csamul_pg_rca24_fa7_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_3_xor1), .fa_or0(u_csamul_pg_rca24_fa7_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_3(.a(a[8]), .b(b[3]), .out(u_csamul_pg_rca24_and8_3));
  fa fa_u_csamul_pg_rca24_fa8_3_out(.a(u_csamul_pg_rca24_and8_3[0]), .b(u_csamul_pg_rca24_fa9_2_xor1[0]), .cin(u_csamul_pg_rca24_fa8_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_3_xor1), .fa_or0(u_csamul_pg_rca24_fa8_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_3(.a(a[9]), .b(b[3]), .out(u_csamul_pg_rca24_and9_3));
  fa fa_u_csamul_pg_rca24_fa9_3_out(.a(u_csamul_pg_rca24_and9_3[0]), .b(u_csamul_pg_rca24_fa10_2_xor1[0]), .cin(u_csamul_pg_rca24_fa9_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_3_xor1), .fa_or0(u_csamul_pg_rca24_fa9_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_3(.a(a[10]), .b(b[3]), .out(u_csamul_pg_rca24_and10_3));
  fa fa_u_csamul_pg_rca24_fa10_3_out(.a(u_csamul_pg_rca24_and10_3[0]), .b(u_csamul_pg_rca24_fa11_2_xor1[0]), .cin(u_csamul_pg_rca24_fa10_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_3_xor1), .fa_or0(u_csamul_pg_rca24_fa10_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_3(.a(a[11]), .b(b[3]), .out(u_csamul_pg_rca24_and11_3));
  fa fa_u_csamul_pg_rca24_fa11_3_out(.a(u_csamul_pg_rca24_and11_3[0]), .b(u_csamul_pg_rca24_fa12_2_xor1[0]), .cin(u_csamul_pg_rca24_fa11_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_3_xor1), .fa_or0(u_csamul_pg_rca24_fa11_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_3(.a(a[12]), .b(b[3]), .out(u_csamul_pg_rca24_and12_3));
  fa fa_u_csamul_pg_rca24_fa12_3_out(.a(u_csamul_pg_rca24_and12_3[0]), .b(u_csamul_pg_rca24_fa13_2_xor1[0]), .cin(u_csamul_pg_rca24_fa12_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_3_xor1), .fa_or0(u_csamul_pg_rca24_fa12_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_3(.a(a[13]), .b(b[3]), .out(u_csamul_pg_rca24_and13_3));
  fa fa_u_csamul_pg_rca24_fa13_3_out(.a(u_csamul_pg_rca24_and13_3[0]), .b(u_csamul_pg_rca24_fa14_2_xor1[0]), .cin(u_csamul_pg_rca24_fa13_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_3_xor1), .fa_or0(u_csamul_pg_rca24_fa13_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_3(.a(a[14]), .b(b[3]), .out(u_csamul_pg_rca24_and14_3));
  fa fa_u_csamul_pg_rca24_fa14_3_out(.a(u_csamul_pg_rca24_and14_3[0]), .b(u_csamul_pg_rca24_fa15_2_xor1[0]), .cin(u_csamul_pg_rca24_fa14_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_3_xor1), .fa_or0(u_csamul_pg_rca24_fa14_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_3(.a(a[15]), .b(b[3]), .out(u_csamul_pg_rca24_and15_3));
  fa fa_u_csamul_pg_rca24_fa15_3_out(.a(u_csamul_pg_rca24_and15_3[0]), .b(u_csamul_pg_rca24_fa16_2_xor1[0]), .cin(u_csamul_pg_rca24_fa15_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_3_xor1), .fa_or0(u_csamul_pg_rca24_fa15_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_3(.a(a[16]), .b(b[3]), .out(u_csamul_pg_rca24_and16_3));
  fa fa_u_csamul_pg_rca24_fa16_3_out(.a(u_csamul_pg_rca24_and16_3[0]), .b(u_csamul_pg_rca24_fa17_2_xor1[0]), .cin(u_csamul_pg_rca24_fa16_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_3_xor1), .fa_or0(u_csamul_pg_rca24_fa16_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_3(.a(a[17]), .b(b[3]), .out(u_csamul_pg_rca24_and17_3));
  fa fa_u_csamul_pg_rca24_fa17_3_out(.a(u_csamul_pg_rca24_and17_3[0]), .b(u_csamul_pg_rca24_fa18_2_xor1[0]), .cin(u_csamul_pg_rca24_fa17_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_3_xor1), .fa_or0(u_csamul_pg_rca24_fa17_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_3(.a(a[18]), .b(b[3]), .out(u_csamul_pg_rca24_and18_3));
  fa fa_u_csamul_pg_rca24_fa18_3_out(.a(u_csamul_pg_rca24_and18_3[0]), .b(u_csamul_pg_rca24_fa19_2_xor1[0]), .cin(u_csamul_pg_rca24_fa18_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_3_xor1), .fa_or0(u_csamul_pg_rca24_fa18_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_3(.a(a[19]), .b(b[3]), .out(u_csamul_pg_rca24_and19_3));
  fa fa_u_csamul_pg_rca24_fa19_3_out(.a(u_csamul_pg_rca24_and19_3[0]), .b(u_csamul_pg_rca24_fa20_2_xor1[0]), .cin(u_csamul_pg_rca24_fa19_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_3_xor1), .fa_or0(u_csamul_pg_rca24_fa19_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_3(.a(a[20]), .b(b[3]), .out(u_csamul_pg_rca24_and20_3));
  fa fa_u_csamul_pg_rca24_fa20_3_out(.a(u_csamul_pg_rca24_and20_3[0]), .b(u_csamul_pg_rca24_fa21_2_xor1[0]), .cin(u_csamul_pg_rca24_fa20_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_3_xor1), .fa_or0(u_csamul_pg_rca24_fa20_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_3(.a(a[21]), .b(b[3]), .out(u_csamul_pg_rca24_and21_3));
  fa fa_u_csamul_pg_rca24_fa21_3_out(.a(u_csamul_pg_rca24_and21_3[0]), .b(u_csamul_pg_rca24_fa22_2_xor1[0]), .cin(u_csamul_pg_rca24_fa21_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_3_xor1), .fa_or0(u_csamul_pg_rca24_fa21_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_3(.a(a[22]), .b(b[3]), .out(u_csamul_pg_rca24_and22_3));
  fa fa_u_csamul_pg_rca24_fa22_3_out(.a(u_csamul_pg_rca24_and22_3[0]), .b(u_csamul_pg_rca24_and23_2[0]), .cin(u_csamul_pg_rca24_fa22_2_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_3_xor1), .fa_or0(u_csamul_pg_rca24_fa22_3_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_3(.a(a[23]), .b(b[3]), .out(u_csamul_pg_rca24_and23_3));
  and_gate and_gate_u_csamul_pg_rca24_and0_4(.a(a[0]), .b(b[4]), .out(u_csamul_pg_rca24_and0_4));
  fa fa_u_csamul_pg_rca24_fa0_4_out(.a(u_csamul_pg_rca24_and0_4[0]), .b(u_csamul_pg_rca24_fa1_3_xor1[0]), .cin(u_csamul_pg_rca24_fa0_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_4_xor1), .fa_or0(u_csamul_pg_rca24_fa0_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_4(.a(a[1]), .b(b[4]), .out(u_csamul_pg_rca24_and1_4));
  fa fa_u_csamul_pg_rca24_fa1_4_out(.a(u_csamul_pg_rca24_and1_4[0]), .b(u_csamul_pg_rca24_fa2_3_xor1[0]), .cin(u_csamul_pg_rca24_fa1_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_4_xor1), .fa_or0(u_csamul_pg_rca24_fa1_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_4(.a(a[2]), .b(b[4]), .out(u_csamul_pg_rca24_and2_4));
  fa fa_u_csamul_pg_rca24_fa2_4_out(.a(u_csamul_pg_rca24_and2_4[0]), .b(u_csamul_pg_rca24_fa3_3_xor1[0]), .cin(u_csamul_pg_rca24_fa2_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_4_xor1), .fa_or0(u_csamul_pg_rca24_fa2_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_4(.a(a[3]), .b(b[4]), .out(u_csamul_pg_rca24_and3_4));
  fa fa_u_csamul_pg_rca24_fa3_4_out(.a(u_csamul_pg_rca24_and3_4[0]), .b(u_csamul_pg_rca24_fa4_3_xor1[0]), .cin(u_csamul_pg_rca24_fa3_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_4_xor1), .fa_or0(u_csamul_pg_rca24_fa3_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_4(.a(a[4]), .b(b[4]), .out(u_csamul_pg_rca24_and4_4));
  fa fa_u_csamul_pg_rca24_fa4_4_out(.a(u_csamul_pg_rca24_and4_4[0]), .b(u_csamul_pg_rca24_fa5_3_xor1[0]), .cin(u_csamul_pg_rca24_fa4_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_4_xor1), .fa_or0(u_csamul_pg_rca24_fa4_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_4(.a(a[5]), .b(b[4]), .out(u_csamul_pg_rca24_and5_4));
  fa fa_u_csamul_pg_rca24_fa5_4_out(.a(u_csamul_pg_rca24_and5_4[0]), .b(u_csamul_pg_rca24_fa6_3_xor1[0]), .cin(u_csamul_pg_rca24_fa5_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_4_xor1), .fa_or0(u_csamul_pg_rca24_fa5_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_4(.a(a[6]), .b(b[4]), .out(u_csamul_pg_rca24_and6_4));
  fa fa_u_csamul_pg_rca24_fa6_4_out(.a(u_csamul_pg_rca24_and6_4[0]), .b(u_csamul_pg_rca24_fa7_3_xor1[0]), .cin(u_csamul_pg_rca24_fa6_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_4_xor1), .fa_or0(u_csamul_pg_rca24_fa6_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_4(.a(a[7]), .b(b[4]), .out(u_csamul_pg_rca24_and7_4));
  fa fa_u_csamul_pg_rca24_fa7_4_out(.a(u_csamul_pg_rca24_and7_4[0]), .b(u_csamul_pg_rca24_fa8_3_xor1[0]), .cin(u_csamul_pg_rca24_fa7_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_4_xor1), .fa_or0(u_csamul_pg_rca24_fa7_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_4(.a(a[8]), .b(b[4]), .out(u_csamul_pg_rca24_and8_4));
  fa fa_u_csamul_pg_rca24_fa8_4_out(.a(u_csamul_pg_rca24_and8_4[0]), .b(u_csamul_pg_rca24_fa9_3_xor1[0]), .cin(u_csamul_pg_rca24_fa8_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_4_xor1), .fa_or0(u_csamul_pg_rca24_fa8_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_4(.a(a[9]), .b(b[4]), .out(u_csamul_pg_rca24_and9_4));
  fa fa_u_csamul_pg_rca24_fa9_4_out(.a(u_csamul_pg_rca24_and9_4[0]), .b(u_csamul_pg_rca24_fa10_3_xor1[0]), .cin(u_csamul_pg_rca24_fa9_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_4_xor1), .fa_or0(u_csamul_pg_rca24_fa9_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_4(.a(a[10]), .b(b[4]), .out(u_csamul_pg_rca24_and10_4));
  fa fa_u_csamul_pg_rca24_fa10_4_out(.a(u_csamul_pg_rca24_and10_4[0]), .b(u_csamul_pg_rca24_fa11_3_xor1[0]), .cin(u_csamul_pg_rca24_fa10_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_4_xor1), .fa_or0(u_csamul_pg_rca24_fa10_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_4(.a(a[11]), .b(b[4]), .out(u_csamul_pg_rca24_and11_4));
  fa fa_u_csamul_pg_rca24_fa11_4_out(.a(u_csamul_pg_rca24_and11_4[0]), .b(u_csamul_pg_rca24_fa12_3_xor1[0]), .cin(u_csamul_pg_rca24_fa11_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_4_xor1), .fa_or0(u_csamul_pg_rca24_fa11_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_4(.a(a[12]), .b(b[4]), .out(u_csamul_pg_rca24_and12_4));
  fa fa_u_csamul_pg_rca24_fa12_4_out(.a(u_csamul_pg_rca24_and12_4[0]), .b(u_csamul_pg_rca24_fa13_3_xor1[0]), .cin(u_csamul_pg_rca24_fa12_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_4_xor1), .fa_or0(u_csamul_pg_rca24_fa12_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_4(.a(a[13]), .b(b[4]), .out(u_csamul_pg_rca24_and13_4));
  fa fa_u_csamul_pg_rca24_fa13_4_out(.a(u_csamul_pg_rca24_and13_4[0]), .b(u_csamul_pg_rca24_fa14_3_xor1[0]), .cin(u_csamul_pg_rca24_fa13_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_4_xor1), .fa_or0(u_csamul_pg_rca24_fa13_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_4(.a(a[14]), .b(b[4]), .out(u_csamul_pg_rca24_and14_4));
  fa fa_u_csamul_pg_rca24_fa14_4_out(.a(u_csamul_pg_rca24_and14_4[0]), .b(u_csamul_pg_rca24_fa15_3_xor1[0]), .cin(u_csamul_pg_rca24_fa14_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_4_xor1), .fa_or0(u_csamul_pg_rca24_fa14_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_4(.a(a[15]), .b(b[4]), .out(u_csamul_pg_rca24_and15_4));
  fa fa_u_csamul_pg_rca24_fa15_4_out(.a(u_csamul_pg_rca24_and15_4[0]), .b(u_csamul_pg_rca24_fa16_3_xor1[0]), .cin(u_csamul_pg_rca24_fa15_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_4_xor1), .fa_or0(u_csamul_pg_rca24_fa15_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_4(.a(a[16]), .b(b[4]), .out(u_csamul_pg_rca24_and16_4));
  fa fa_u_csamul_pg_rca24_fa16_4_out(.a(u_csamul_pg_rca24_and16_4[0]), .b(u_csamul_pg_rca24_fa17_3_xor1[0]), .cin(u_csamul_pg_rca24_fa16_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_4_xor1), .fa_or0(u_csamul_pg_rca24_fa16_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_4(.a(a[17]), .b(b[4]), .out(u_csamul_pg_rca24_and17_4));
  fa fa_u_csamul_pg_rca24_fa17_4_out(.a(u_csamul_pg_rca24_and17_4[0]), .b(u_csamul_pg_rca24_fa18_3_xor1[0]), .cin(u_csamul_pg_rca24_fa17_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_4_xor1), .fa_or0(u_csamul_pg_rca24_fa17_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_4(.a(a[18]), .b(b[4]), .out(u_csamul_pg_rca24_and18_4));
  fa fa_u_csamul_pg_rca24_fa18_4_out(.a(u_csamul_pg_rca24_and18_4[0]), .b(u_csamul_pg_rca24_fa19_3_xor1[0]), .cin(u_csamul_pg_rca24_fa18_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_4_xor1), .fa_or0(u_csamul_pg_rca24_fa18_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_4(.a(a[19]), .b(b[4]), .out(u_csamul_pg_rca24_and19_4));
  fa fa_u_csamul_pg_rca24_fa19_4_out(.a(u_csamul_pg_rca24_and19_4[0]), .b(u_csamul_pg_rca24_fa20_3_xor1[0]), .cin(u_csamul_pg_rca24_fa19_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_4_xor1), .fa_or0(u_csamul_pg_rca24_fa19_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_4(.a(a[20]), .b(b[4]), .out(u_csamul_pg_rca24_and20_4));
  fa fa_u_csamul_pg_rca24_fa20_4_out(.a(u_csamul_pg_rca24_and20_4[0]), .b(u_csamul_pg_rca24_fa21_3_xor1[0]), .cin(u_csamul_pg_rca24_fa20_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_4_xor1), .fa_or0(u_csamul_pg_rca24_fa20_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_4(.a(a[21]), .b(b[4]), .out(u_csamul_pg_rca24_and21_4));
  fa fa_u_csamul_pg_rca24_fa21_4_out(.a(u_csamul_pg_rca24_and21_4[0]), .b(u_csamul_pg_rca24_fa22_3_xor1[0]), .cin(u_csamul_pg_rca24_fa21_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_4_xor1), .fa_or0(u_csamul_pg_rca24_fa21_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_4(.a(a[22]), .b(b[4]), .out(u_csamul_pg_rca24_and22_4));
  fa fa_u_csamul_pg_rca24_fa22_4_out(.a(u_csamul_pg_rca24_and22_4[0]), .b(u_csamul_pg_rca24_and23_3[0]), .cin(u_csamul_pg_rca24_fa22_3_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_4_xor1), .fa_or0(u_csamul_pg_rca24_fa22_4_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_4(.a(a[23]), .b(b[4]), .out(u_csamul_pg_rca24_and23_4));
  and_gate and_gate_u_csamul_pg_rca24_and0_5(.a(a[0]), .b(b[5]), .out(u_csamul_pg_rca24_and0_5));
  fa fa_u_csamul_pg_rca24_fa0_5_out(.a(u_csamul_pg_rca24_and0_5[0]), .b(u_csamul_pg_rca24_fa1_4_xor1[0]), .cin(u_csamul_pg_rca24_fa0_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_5_xor1), .fa_or0(u_csamul_pg_rca24_fa0_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_5(.a(a[1]), .b(b[5]), .out(u_csamul_pg_rca24_and1_5));
  fa fa_u_csamul_pg_rca24_fa1_5_out(.a(u_csamul_pg_rca24_and1_5[0]), .b(u_csamul_pg_rca24_fa2_4_xor1[0]), .cin(u_csamul_pg_rca24_fa1_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_5_xor1), .fa_or0(u_csamul_pg_rca24_fa1_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_5(.a(a[2]), .b(b[5]), .out(u_csamul_pg_rca24_and2_5));
  fa fa_u_csamul_pg_rca24_fa2_5_out(.a(u_csamul_pg_rca24_and2_5[0]), .b(u_csamul_pg_rca24_fa3_4_xor1[0]), .cin(u_csamul_pg_rca24_fa2_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_5_xor1), .fa_or0(u_csamul_pg_rca24_fa2_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_5(.a(a[3]), .b(b[5]), .out(u_csamul_pg_rca24_and3_5));
  fa fa_u_csamul_pg_rca24_fa3_5_out(.a(u_csamul_pg_rca24_and3_5[0]), .b(u_csamul_pg_rca24_fa4_4_xor1[0]), .cin(u_csamul_pg_rca24_fa3_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_5_xor1), .fa_or0(u_csamul_pg_rca24_fa3_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_5(.a(a[4]), .b(b[5]), .out(u_csamul_pg_rca24_and4_5));
  fa fa_u_csamul_pg_rca24_fa4_5_out(.a(u_csamul_pg_rca24_and4_5[0]), .b(u_csamul_pg_rca24_fa5_4_xor1[0]), .cin(u_csamul_pg_rca24_fa4_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_5_xor1), .fa_or0(u_csamul_pg_rca24_fa4_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_5(.a(a[5]), .b(b[5]), .out(u_csamul_pg_rca24_and5_5));
  fa fa_u_csamul_pg_rca24_fa5_5_out(.a(u_csamul_pg_rca24_and5_5[0]), .b(u_csamul_pg_rca24_fa6_4_xor1[0]), .cin(u_csamul_pg_rca24_fa5_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_5_xor1), .fa_or0(u_csamul_pg_rca24_fa5_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_5(.a(a[6]), .b(b[5]), .out(u_csamul_pg_rca24_and6_5));
  fa fa_u_csamul_pg_rca24_fa6_5_out(.a(u_csamul_pg_rca24_and6_5[0]), .b(u_csamul_pg_rca24_fa7_4_xor1[0]), .cin(u_csamul_pg_rca24_fa6_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_5_xor1), .fa_or0(u_csamul_pg_rca24_fa6_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_5(.a(a[7]), .b(b[5]), .out(u_csamul_pg_rca24_and7_5));
  fa fa_u_csamul_pg_rca24_fa7_5_out(.a(u_csamul_pg_rca24_and7_5[0]), .b(u_csamul_pg_rca24_fa8_4_xor1[0]), .cin(u_csamul_pg_rca24_fa7_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_5_xor1), .fa_or0(u_csamul_pg_rca24_fa7_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_5(.a(a[8]), .b(b[5]), .out(u_csamul_pg_rca24_and8_5));
  fa fa_u_csamul_pg_rca24_fa8_5_out(.a(u_csamul_pg_rca24_and8_5[0]), .b(u_csamul_pg_rca24_fa9_4_xor1[0]), .cin(u_csamul_pg_rca24_fa8_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_5_xor1), .fa_or0(u_csamul_pg_rca24_fa8_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_5(.a(a[9]), .b(b[5]), .out(u_csamul_pg_rca24_and9_5));
  fa fa_u_csamul_pg_rca24_fa9_5_out(.a(u_csamul_pg_rca24_and9_5[0]), .b(u_csamul_pg_rca24_fa10_4_xor1[0]), .cin(u_csamul_pg_rca24_fa9_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_5_xor1), .fa_or0(u_csamul_pg_rca24_fa9_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_5(.a(a[10]), .b(b[5]), .out(u_csamul_pg_rca24_and10_5));
  fa fa_u_csamul_pg_rca24_fa10_5_out(.a(u_csamul_pg_rca24_and10_5[0]), .b(u_csamul_pg_rca24_fa11_4_xor1[0]), .cin(u_csamul_pg_rca24_fa10_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_5_xor1), .fa_or0(u_csamul_pg_rca24_fa10_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_5(.a(a[11]), .b(b[5]), .out(u_csamul_pg_rca24_and11_5));
  fa fa_u_csamul_pg_rca24_fa11_5_out(.a(u_csamul_pg_rca24_and11_5[0]), .b(u_csamul_pg_rca24_fa12_4_xor1[0]), .cin(u_csamul_pg_rca24_fa11_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_5_xor1), .fa_or0(u_csamul_pg_rca24_fa11_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_5(.a(a[12]), .b(b[5]), .out(u_csamul_pg_rca24_and12_5));
  fa fa_u_csamul_pg_rca24_fa12_5_out(.a(u_csamul_pg_rca24_and12_5[0]), .b(u_csamul_pg_rca24_fa13_4_xor1[0]), .cin(u_csamul_pg_rca24_fa12_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_5_xor1), .fa_or0(u_csamul_pg_rca24_fa12_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_5(.a(a[13]), .b(b[5]), .out(u_csamul_pg_rca24_and13_5));
  fa fa_u_csamul_pg_rca24_fa13_5_out(.a(u_csamul_pg_rca24_and13_5[0]), .b(u_csamul_pg_rca24_fa14_4_xor1[0]), .cin(u_csamul_pg_rca24_fa13_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_5_xor1), .fa_or0(u_csamul_pg_rca24_fa13_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_5(.a(a[14]), .b(b[5]), .out(u_csamul_pg_rca24_and14_5));
  fa fa_u_csamul_pg_rca24_fa14_5_out(.a(u_csamul_pg_rca24_and14_5[0]), .b(u_csamul_pg_rca24_fa15_4_xor1[0]), .cin(u_csamul_pg_rca24_fa14_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_5_xor1), .fa_or0(u_csamul_pg_rca24_fa14_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_5(.a(a[15]), .b(b[5]), .out(u_csamul_pg_rca24_and15_5));
  fa fa_u_csamul_pg_rca24_fa15_5_out(.a(u_csamul_pg_rca24_and15_5[0]), .b(u_csamul_pg_rca24_fa16_4_xor1[0]), .cin(u_csamul_pg_rca24_fa15_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_5_xor1), .fa_or0(u_csamul_pg_rca24_fa15_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_5(.a(a[16]), .b(b[5]), .out(u_csamul_pg_rca24_and16_5));
  fa fa_u_csamul_pg_rca24_fa16_5_out(.a(u_csamul_pg_rca24_and16_5[0]), .b(u_csamul_pg_rca24_fa17_4_xor1[0]), .cin(u_csamul_pg_rca24_fa16_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_5_xor1), .fa_or0(u_csamul_pg_rca24_fa16_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_5(.a(a[17]), .b(b[5]), .out(u_csamul_pg_rca24_and17_5));
  fa fa_u_csamul_pg_rca24_fa17_5_out(.a(u_csamul_pg_rca24_and17_5[0]), .b(u_csamul_pg_rca24_fa18_4_xor1[0]), .cin(u_csamul_pg_rca24_fa17_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_5_xor1), .fa_or0(u_csamul_pg_rca24_fa17_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_5(.a(a[18]), .b(b[5]), .out(u_csamul_pg_rca24_and18_5));
  fa fa_u_csamul_pg_rca24_fa18_5_out(.a(u_csamul_pg_rca24_and18_5[0]), .b(u_csamul_pg_rca24_fa19_4_xor1[0]), .cin(u_csamul_pg_rca24_fa18_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_5_xor1), .fa_or0(u_csamul_pg_rca24_fa18_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_5(.a(a[19]), .b(b[5]), .out(u_csamul_pg_rca24_and19_5));
  fa fa_u_csamul_pg_rca24_fa19_5_out(.a(u_csamul_pg_rca24_and19_5[0]), .b(u_csamul_pg_rca24_fa20_4_xor1[0]), .cin(u_csamul_pg_rca24_fa19_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_5_xor1), .fa_or0(u_csamul_pg_rca24_fa19_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_5(.a(a[20]), .b(b[5]), .out(u_csamul_pg_rca24_and20_5));
  fa fa_u_csamul_pg_rca24_fa20_5_out(.a(u_csamul_pg_rca24_and20_5[0]), .b(u_csamul_pg_rca24_fa21_4_xor1[0]), .cin(u_csamul_pg_rca24_fa20_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_5_xor1), .fa_or0(u_csamul_pg_rca24_fa20_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_5(.a(a[21]), .b(b[5]), .out(u_csamul_pg_rca24_and21_5));
  fa fa_u_csamul_pg_rca24_fa21_5_out(.a(u_csamul_pg_rca24_and21_5[0]), .b(u_csamul_pg_rca24_fa22_4_xor1[0]), .cin(u_csamul_pg_rca24_fa21_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_5_xor1), .fa_or0(u_csamul_pg_rca24_fa21_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_5(.a(a[22]), .b(b[5]), .out(u_csamul_pg_rca24_and22_5));
  fa fa_u_csamul_pg_rca24_fa22_5_out(.a(u_csamul_pg_rca24_and22_5[0]), .b(u_csamul_pg_rca24_and23_4[0]), .cin(u_csamul_pg_rca24_fa22_4_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_5_xor1), .fa_or0(u_csamul_pg_rca24_fa22_5_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_5(.a(a[23]), .b(b[5]), .out(u_csamul_pg_rca24_and23_5));
  and_gate and_gate_u_csamul_pg_rca24_and0_6(.a(a[0]), .b(b[6]), .out(u_csamul_pg_rca24_and0_6));
  fa fa_u_csamul_pg_rca24_fa0_6_out(.a(u_csamul_pg_rca24_and0_6[0]), .b(u_csamul_pg_rca24_fa1_5_xor1[0]), .cin(u_csamul_pg_rca24_fa0_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_6_xor1), .fa_or0(u_csamul_pg_rca24_fa0_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_6(.a(a[1]), .b(b[6]), .out(u_csamul_pg_rca24_and1_6));
  fa fa_u_csamul_pg_rca24_fa1_6_out(.a(u_csamul_pg_rca24_and1_6[0]), .b(u_csamul_pg_rca24_fa2_5_xor1[0]), .cin(u_csamul_pg_rca24_fa1_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_6_xor1), .fa_or0(u_csamul_pg_rca24_fa1_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_6(.a(a[2]), .b(b[6]), .out(u_csamul_pg_rca24_and2_6));
  fa fa_u_csamul_pg_rca24_fa2_6_out(.a(u_csamul_pg_rca24_and2_6[0]), .b(u_csamul_pg_rca24_fa3_5_xor1[0]), .cin(u_csamul_pg_rca24_fa2_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_6_xor1), .fa_or0(u_csamul_pg_rca24_fa2_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_6(.a(a[3]), .b(b[6]), .out(u_csamul_pg_rca24_and3_6));
  fa fa_u_csamul_pg_rca24_fa3_6_out(.a(u_csamul_pg_rca24_and3_6[0]), .b(u_csamul_pg_rca24_fa4_5_xor1[0]), .cin(u_csamul_pg_rca24_fa3_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_6_xor1), .fa_or0(u_csamul_pg_rca24_fa3_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_6(.a(a[4]), .b(b[6]), .out(u_csamul_pg_rca24_and4_6));
  fa fa_u_csamul_pg_rca24_fa4_6_out(.a(u_csamul_pg_rca24_and4_6[0]), .b(u_csamul_pg_rca24_fa5_5_xor1[0]), .cin(u_csamul_pg_rca24_fa4_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_6_xor1), .fa_or0(u_csamul_pg_rca24_fa4_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_6(.a(a[5]), .b(b[6]), .out(u_csamul_pg_rca24_and5_6));
  fa fa_u_csamul_pg_rca24_fa5_6_out(.a(u_csamul_pg_rca24_and5_6[0]), .b(u_csamul_pg_rca24_fa6_5_xor1[0]), .cin(u_csamul_pg_rca24_fa5_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_6_xor1), .fa_or0(u_csamul_pg_rca24_fa5_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_6(.a(a[6]), .b(b[6]), .out(u_csamul_pg_rca24_and6_6));
  fa fa_u_csamul_pg_rca24_fa6_6_out(.a(u_csamul_pg_rca24_and6_6[0]), .b(u_csamul_pg_rca24_fa7_5_xor1[0]), .cin(u_csamul_pg_rca24_fa6_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_6_xor1), .fa_or0(u_csamul_pg_rca24_fa6_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_6(.a(a[7]), .b(b[6]), .out(u_csamul_pg_rca24_and7_6));
  fa fa_u_csamul_pg_rca24_fa7_6_out(.a(u_csamul_pg_rca24_and7_6[0]), .b(u_csamul_pg_rca24_fa8_5_xor1[0]), .cin(u_csamul_pg_rca24_fa7_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_6_xor1), .fa_or0(u_csamul_pg_rca24_fa7_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_6(.a(a[8]), .b(b[6]), .out(u_csamul_pg_rca24_and8_6));
  fa fa_u_csamul_pg_rca24_fa8_6_out(.a(u_csamul_pg_rca24_and8_6[0]), .b(u_csamul_pg_rca24_fa9_5_xor1[0]), .cin(u_csamul_pg_rca24_fa8_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_6_xor1), .fa_or0(u_csamul_pg_rca24_fa8_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_6(.a(a[9]), .b(b[6]), .out(u_csamul_pg_rca24_and9_6));
  fa fa_u_csamul_pg_rca24_fa9_6_out(.a(u_csamul_pg_rca24_and9_6[0]), .b(u_csamul_pg_rca24_fa10_5_xor1[0]), .cin(u_csamul_pg_rca24_fa9_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_6_xor1), .fa_or0(u_csamul_pg_rca24_fa9_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_6(.a(a[10]), .b(b[6]), .out(u_csamul_pg_rca24_and10_6));
  fa fa_u_csamul_pg_rca24_fa10_6_out(.a(u_csamul_pg_rca24_and10_6[0]), .b(u_csamul_pg_rca24_fa11_5_xor1[0]), .cin(u_csamul_pg_rca24_fa10_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_6_xor1), .fa_or0(u_csamul_pg_rca24_fa10_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_6(.a(a[11]), .b(b[6]), .out(u_csamul_pg_rca24_and11_6));
  fa fa_u_csamul_pg_rca24_fa11_6_out(.a(u_csamul_pg_rca24_and11_6[0]), .b(u_csamul_pg_rca24_fa12_5_xor1[0]), .cin(u_csamul_pg_rca24_fa11_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_6_xor1), .fa_or0(u_csamul_pg_rca24_fa11_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_6(.a(a[12]), .b(b[6]), .out(u_csamul_pg_rca24_and12_6));
  fa fa_u_csamul_pg_rca24_fa12_6_out(.a(u_csamul_pg_rca24_and12_6[0]), .b(u_csamul_pg_rca24_fa13_5_xor1[0]), .cin(u_csamul_pg_rca24_fa12_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_6_xor1), .fa_or0(u_csamul_pg_rca24_fa12_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_6(.a(a[13]), .b(b[6]), .out(u_csamul_pg_rca24_and13_6));
  fa fa_u_csamul_pg_rca24_fa13_6_out(.a(u_csamul_pg_rca24_and13_6[0]), .b(u_csamul_pg_rca24_fa14_5_xor1[0]), .cin(u_csamul_pg_rca24_fa13_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_6_xor1), .fa_or0(u_csamul_pg_rca24_fa13_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_6(.a(a[14]), .b(b[6]), .out(u_csamul_pg_rca24_and14_6));
  fa fa_u_csamul_pg_rca24_fa14_6_out(.a(u_csamul_pg_rca24_and14_6[0]), .b(u_csamul_pg_rca24_fa15_5_xor1[0]), .cin(u_csamul_pg_rca24_fa14_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_6_xor1), .fa_or0(u_csamul_pg_rca24_fa14_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_6(.a(a[15]), .b(b[6]), .out(u_csamul_pg_rca24_and15_6));
  fa fa_u_csamul_pg_rca24_fa15_6_out(.a(u_csamul_pg_rca24_and15_6[0]), .b(u_csamul_pg_rca24_fa16_5_xor1[0]), .cin(u_csamul_pg_rca24_fa15_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_6_xor1), .fa_or0(u_csamul_pg_rca24_fa15_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_6(.a(a[16]), .b(b[6]), .out(u_csamul_pg_rca24_and16_6));
  fa fa_u_csamul_pg_rca24_fa16_6_out(.a(u_csamul_pg_rca24_and16_6[0]), .b(u_csamul_pg_rca24_fa17_5_xor1[0]), .cin(u_csamul_pg_rca24_fa16_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_6_xor1), .fa_or0(u_csamul_pg_rca24_fa16_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_6(.a(a[17]), .b(b[6]), .out(u_csamul_pg_rca24_and17_6));
  fa fa_u_csamul_pg_rca24_fa17_6_out(.a(u_csamul_pg_rca24_and17_6[0]), .b(u_csamul_pg_rca24_fa18_5_xor1[0]), .cin(u_csamul_pg_rca24_fa17_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_6_xor1), .fa_or0(u_csamul_pg_rca24_fa17_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_6(.a(a[18]), .b(b[6]), .out(u_csamul_pg_rca24_and18_6));
  fa fa_u_csamul_pg_rca24_fa18_6_out(.a(u_csamul_pg_rca24_and18_6[0]), .b(u_csamul_pg_rca24_fa19_5_xor1[0]), .cin(u_csamul_pg_rca24_fa18_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_6_xor1), .fa_or0(u_csamul_pg_rca24_fa18_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_6(.a(a[19]), .b(b[6]), .out(u_csamul_pg_rca24_and19_6));
  fa fa_u_csamul_pg_rca24_fa19_6_out(.a(u_csamul_pg_rca24_and19_6[0]), .b(u_csamul_pg_rca24_fa20_5_xor1[0]), .cin(u_csamul_pg_rca24_fa19_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_6_xor1), .fa_or0(u_csamul_pg_rca24_fa19_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_6(.a(a[20]), .b(b[6]), .out(u_csamul_pg_rca24_and20_6));
  fa fa_u_csamul_pg_rca24_fa20_6_out(.a(u_csamul_pg_rca24_and20_6[0]), .b(u_csamul_pg_rca24_fa21_5_xor1[0]), .cin(u_csamul_pg_rca24_fa20_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_6_xor1), .fa_or0(u_csamul_pg_rca24_fa20_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_6(.a(a[21]), .b(b[6]), .out(u_csamul_pg_rca24_and21_6));
  fa fa_u_csamul_pg_rca24_fa21_6_out(.a(u_csamul_pg_rca24_and21_6[0]), .b(u_csamul_pg_rca24_fa22_5_xor1[0]), .cin(u_csamul_pg_rca24_fa21_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_6_xor1), .fa_or0(u_csamul_pg_rca24_fa21_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_6(.a(a[22]), .b(b[6]), .out(u_csamul_pg_rca24_and22_6));
  fa fa_u_csamul_pg_rca24_fa22_6_out(.a(u_csamul_pg_rca24_and22_6[0]), .b(u_csamul_pg_rca24_and23_5[0]), .cin(u_csamul_pg_rca24_fa22_5_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_6_xor1), .fa_or0(u_csamul_pg_rca24_fa22_6_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_6(.a(a[23]), .b(b[6]), .out(u_csamul_pg_rca24_and23_6));
  and_gate and_gate_u_csamul_pg_rca24_and0_7(.a(a[0]), .b(b[7]), .out(u_csamul_pg_rca24_and0_7));
  fa fa_u_csamul_pg_rca24_fa0_7_out(.a(u_csamul_pg_rca24_and0_7[0]), .b(u_csamul_pg_rca24_fa1_6_xor1[0]), .cin(u_csamul_pg_rca24_fa0_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_7_xor1), .fa_or0(u_csamul_pg_rca24_fa0_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_7(.a(a[1]), .b(b[7]), .out(u_csamul_pg_rca24_and1_7));
  fa fa_u_csamul_pg_rca24_fa1_7_out(.a(u_csamul_pg_rca24_and1_7[0]), .b(u_csamul_pg_rca24_fa2_6_xor1[0]), .cin(u_csamul_pg_rca24_fa1_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_7_xor1), .fa_or0(u_csamul_pg_rca24_fa1_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_7(.a(a[2]), .b(b[7]), .out(u_csamul_pg_rca24_and2_7));
  fa fa_u_csamul_pg_rca24_fa2_7_out(.a(u_csamul_pg_rca24_and2_7[0]), .b(u_csamul_pg_rca24_fa3_6_xor1[0]), .cin(u_csamul_pg_rca24_fa2_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_7_xor1), .fa_or0(u_csamul_pg_rca24_fa2_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_7(.a(a[3]), .b(b[7]), .out(u_csamul_pg_rca24_and3_7));
  fa fa_u_csamul_pg_rca24_fa3_7_out(.a(u_csamul_pg_rca24_and3_7[0]), .b(u_csamul_pg_rca24_fa4_6_xor1[0]), .cin(u_csamul_pg_rca24_fa3_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_7_xor1), .fa_or0(u_csamul_pg_rca24_fa3_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_7(.a(a[4]), .b(b[7]), .out(u_csamul_pg_rca24_and4_7));
  fa fa_u_csamul_pg_rca24_fa4_7_out(.a(u_csamul_pg_rca24_and4_7[0]), .b(u_csamul_pg_rca24_fa5_6_xor1[0]), .cin(u_csamul_pg_rca24_fa4_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_7_xor1), .fa_or0(u_csamul_pg_rca24_fa4_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_7(.a(a[5]), .b(b[7]), .out(u_csamul_pg_rca24_and5_7));
  fa fa_u_csamul_pg_rca24_fa5_7_out(.a(u_csamul_pg_rca24_and5_7[0]), .b(u_csamul_pg_rca24_fa6_6_xor1[0]), .cin(u_csamul_pg_rca24_fa5_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_7_xor1), .fa_or0(u_csamul_pg_rca24_fa5_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_7(.a(a[6]), .b(b[7]), .out(u_csamul_pg_rca24_and6_7));
  fa fa_u_csamul_pg_rca24_fa6_7_out(.a(u_csamul_pg_rca24_and6_7[0]), .b(u_csamul_pg_rca24_fa7_6_xor1[0]), .cin(u_csamul_pg_rca24_fa6_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_7_xor1), .fa_or0(u_csamul_pg_rca24_fa6_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_7(.a(a[7]), .b(b[7]), .out(u_csamul_pg_rca24_and7_7));
  fa fa_u_csamul_pg_rca24_fa7_7_out(.a(u_csamul_pg_rca24_and7_7[0]), .b(u_csamul_pg_rca24_fa8_6_xor1[0]), .cin(u_csamul_pg_rca24_fa7_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_7_xor1), .fa_or0(u_csamul_pg_rca24_fa7_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_7(.a(a[8]), .b(b[7]), .out(u_csamul_pg_rca24_and8_7));
  fa fa_u_csamul_pg_rca24_fa8_7_out(.a(u_csamul_pg_rca24_and8_7[0]), .b(u_csamul_pg_rca24_fa9_6_xor1[0]), .cin(u_csamul_pg_rca24_fa8_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_7_xor1), .fa_or0(u_csamul_pg_rca24_fa8_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_7(.a(a[9]), .b(b[7]), .out(u_csamul_pg_rca24_and9_7));
  fa fa_u_csamul_pg_rca24_fa9_7_out(.a(u_csamul_pg_rca24_and9_7[0]), .b(u_csamul_pg_rca24_fa10_6_xor1[0]), .cin(u_csamul_pg_rca24_fa9_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_7_xor1), .fa_or0(u_csamul_pg_rca24_fa9_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_7(.a(a[10]), .b(b[7]), .out(u_csamul_pg_rca24_and10_7));
  fa fa_u_csamul_pg_rca24_fa10_7_out(.a(u_csamul_pg_rca24_and10_7[0]), .b(u_csamul_pg_rca24_fa11_6_xor1[0]), .cin(u_csamul_pg_rca24_fa10_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_7_xor1), .fa_or0(u_csamul_pg_rca24_fa10_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_7(.a(a[11]), .b(b[7]), .out(u_csamul_pg_rca24_and11_7));
  fa fa_u_csamul_pg_rca24_fa11_7_out(.a(u_csamul_pg_rca24_and11_7[0]), .b(u_csamul_pg_rca24_fa12_6_xor1[0]), .cin(u_csamul_pg_rca24_fa11_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_7_xor1), .fa_or0(u_csamul_pg_rca24_fa11_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_7(.a(a[12]), .b(b[7]), .out(u_csamul_pg_rca24_and12_7));
  fa fa_u_csamul_pg_rca24_fa12_7_out(.a(u_csamul_pg_rca24_and12_7[0]), .b(u_csamul_pg_rca24_fa13_6_xor1[0]), .cin(u_csamul_pg_rca24_fa12_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_7_xor1), .fa_or0(u_csamul_pg_rca24_fa12_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_7(.a(a[13]), .b(b[7]), .out(u_csamul_pg_rca24_and13_7));
  fa fa_u_csamul_pg_rca24_fa13_7_out(.a(u_csamul_pg_rca24_and13_7[0]), .b(u_csamul_pg_rca24_fa14_6_xor1[0]), .cin(u_csamul_pg_rca24_fa13_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_7_xor1), .fa_or0(u_csamul_pg_rca24_fa13_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_7(.a(a[14]), .b(b[7]), .out(u_csamul_pg_rca24_and14_7));
  fa fa_u_csamul_pg_rca24_fa14_7_out(.a(u_csamul_pg_rca24_and14_7[0]), .b(u_csamul_pg_rca24_fa15_6_xor1[0]), .cin(u_csamul_pg_rca24_fa14_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_7_xor1), .fa_or0(u_csamul_pg_rca24_fa14_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_7(.a(a[15]), .b(b[7]), .out(u_csamul_pg_rca24_and15_7));
  fa fa_u_csamul_pg_rca24_fa15_7_out(.a(u_csamul_pg_rca24_and15_7[0]), .b(u_csamul_pg_rca24_fa16_6_xor1[0]), .cin(u_csamul_pg_rca24_fa15_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_7_xor1), .fa_or0(u_csamul_pg_rca24_fa15_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_7(.a(a[16]), .b(b[7]), .out(u_csamul_pg_rca24_and16_7));
  fa fa_u_csamul_pg_rca24_fa16_7_out(.a(u_csamul_pg_rca24_and16_7[0]), .b(u_csamul_pg_rca24_fa17_6_xor1[0]), .cin(u_csamul_pg_rca24_fa16_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_7_xor1), .fa_or0(u_csamul_pg_rca24_fa16_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_7(.a(a[17]), .b(b[7]), .out(u_csamul_pg_rca24_and17_7));
  fa fa_u_csamul_pg_rca24_fa17_7_out(.a(u_csamul_pg_rca24_and17_7[0]), .b(u_csamul_pg_rca24_fa18_6_xor1[0]), .cin(u_csamul_pg_rca24_fa17_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_7_xor1), .fa_or0(u_csamul_pg_rca24_fa17_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_7(.a(a[18]), .b(b[7]), .out(u_csamul_pg_rca24_and18_7));
  fa fa_u_csamul_pg_rca24_fa18_7_out(.a(u_csamul_pg_rca24_and18_7[0]), .b(u_csamul_pg_rca24_fa19_6_xor1[0]), .cin(u_csamul_pg_rca24_fa18_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_7_xor1), .fa_or0(u_csamul_pg_rca24_fa18_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_7(.a(a[19]), .b(b[7]), .out(u_csamul_pg_rca24_and19_7));
  fa fa_u_csamul_pg_rca24_fa19_7_out(.a(u_csamul_pg_rca24_and19_7[0]), .b(u_csamul_pg_rca24_fa20_6_xor1[0]), .cin(u_csamul_pg_rca24_fa19_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_7_xor1), .fa_or0(u_csamul_pg_rca24_fa19_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_7(.a(a[20]), .b(b[7]), .out(u_csamul_pg_rca24_and20_7));
  fa fa_u_csamul_pg_rca24_fa20_7_out(.a(u_csamul_pg_rca24_and20_7[0]), .b(u_csamul_pg_rca24_fa21_6_xor1[0]), .cin(u_csamul_pg_rca24_fa20_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_7_xor1), .fa_or0(u_csamul_pg_rca24_fa20_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_7(.a(a[21]), .b(b[7]), .out(u_csamul_pg_rca24_and21_7));
  fa fa_u_csamul_pg_rca24_fa21_7_out(.a(u_csamul_pg_rca24_and21_7[0]), .b(u_csamul_pg_rca24_fa22_6_xor1[0]), .cin(u_csamul_pg_rca24_fa21_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_7_xor1), .fa_or0(u_csamul_pg_rca24_fa21_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_7(.a(a[22]), .b(b[7]), .out(u_csamul_pg_rca24_and22_7));
  fa fa_u_csamul_pg_rca24_fa22_7_out(.a(u_csamul_pg_rca24_and22_7[0]), .b(u_csamul_pg_rca24_and23_6[0]), .cin(u_csamul_pg_rca24_fa22_6_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_7_xor1), .fa_or0(u_csamul_pg_rca24_fa22_7_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_7(.a(a[23]), .b(b[7]), .out(u_csamul_pg_rca24_and23_7));
  and_gate and_gate_u_csamul_pg_rca24_and0_8(.a(a[0]), .b(b[8]), .out(u_csamul_pg_rca24_and0_8));
  fa fa_u_csamul_pg_rca24_fa0_8_out(.a(u_csamul_pg_rca24_and0_8[0]), .b(u_csamul_pg_rca24_fa1_7_xor1[0]), .cin(u_csamul_pg_rca24_fa0_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_8_xor1), .fa_or0(u_csamul_pg_rca24_fa0_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_8(.a(a[1]), .b(b[8]), .out(u_csamul_pg_rca24_and1_8));
  fa fa_u_csamul_pg_rca24_fa1_8_out(.a(u_csamul_pg_rca24_and1_8[0]), .b(u_csamul_pg_rca24_fa2_7_xor1[0]), .cin(u_csamul_pg_rca24_fa1_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_8_xor1), .fa_or0(u_csamul_pg_rca24_fa1_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_8(.a(a[2]), .b(b[8]), .out(u_csamul_pg_rca24_and2_8));
  fa fa_u_csamul_pg_rca24_fa2_8_out(.a(u_csamul_pg_rca24_and2_8[0]), .b(u_csamul_pg_rca24_fa3_7_xor1[0]), .cin(u_csamul_pg_rca24_fa2_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_8_xor1), .fa_or0(u_csamul_pg_rca24_fa2_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_8(.a(a[3]), .b(b[8]), .out(u_csamul_pg_rca24_and3_8));
  fa fa_u_csamul_pg_rca24_fa3_8_out(.a(u_csamul_pg_rca24_and3_8[0]), .b(u_csamul_pg_rca24_fa4_7_xor1[0]), .cin(u_csamul_pg_rca24_fa3_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_8_xor1), .fa_or0(u_csamul_pg_rca24_fa3_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_8(.a(a[4]), .b(b[8]), .out(u_csamul_pg_rca24_and4_8));
  fa fa_u_csamul_pg_rca24_fa4_8_out(.a(u_csamul_pg_rca24_and4_8[0]), .b(u_csamul_pg_rca24_fa5_7_xor1[0]), .cin(u_csamul_pg_rca24_fa4_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_8_xor1), .fa_or0(u_csamul_pg_rca24_fa4_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_8(.a(a[5]), .b(b[8]), .out(u_csamul_pg_rca24_and5_8));
  fa fa_u_csamul_pg_rca24_fa5_8_out(.a(u_csamul_pg_rca24_and5_8[0]), .b(u_csamul_pg_rca24_fa6_7_xor1[0]), .cin(u_csamul_pg_rca24_fa5_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_8_xor1), .fa_or0(u_csamul_pg_rca24_fa5_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_8(.a(a[6]), .b(b[8]), .out(u_csamul_pg_rca24_and6_8));
  fa fa_u_csamul_pg_rca24_fa6_8_out(.a(u_csamul_pg_rca24_and6_8[0]), .b(u_csamul_pg_rca24_fa7_7_xor1[0]), .cin(u_csamul_pg_rca24_fa6_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_8_xor1), .fa_or0(u_csamul_pg_rca24_fa6_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_8(.a(a[7]), .b(b[8]), .out(u_csamul_pg_rca24_and7_8));
  fa fa_u_csamul_pg_rca24_fa7_8_out(.a(u_csamul_pg_rca24_and7_8[0]), .b(u_csamul_pg_rca24_fa8_7_xor1[0]), .cin(u_csamul_pg_rca24_fa7_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_8_xor1), .fa_or0(u_csamul_pg_rca24_fa7_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_8(.a(a[8]), .b(b[8]), .out(u_csamul_pg_rca24_and8_8));
  fa fa_u_csamul_pg_rca24_fa8_8_out(.a(u_csamul_pg_rca24_and8_8[0]), .b(u_csamul_pg_rca24_fa9_7_xor1[0]), .cin(u_csamul_pg_rca24_fa8_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_8_xor1), .fa_or0(u_csamul_pg_rca24_fa8_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_8(.a(a[9]), .b(b[8]), .out(u_csamul_pg_rca24_and9_8));
  fa fa_u_csamul_pg_rca24_fa9_8_out(.a(u_csamul_pg_rca24_and9_8[0]), .b(u_csamul_pg_rca24_fa10_7_xor1[0]), .cin(u_csamul_pg_rca24_fa9_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_8_xor1), .fa_or0(u_csamul_pg_rca24_fa9_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_8(.a(a[10]), .b(b[8]), .out(u_csamul_pg_rca24_and10_8));
  fa fa_u_csamul_pg_rca24_fa10_8_out(.a(u_csamul_pg_rca24_and10_8[0]), .b(u_csamul_pg_rca24_fa11_7_xor1[0]), .cin(u_csamul_pg_rca24_fa10_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_8_xor1), .fa_or0(u_csamul_pg_rca24_fa10_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_8(.a(a[11]), .b(b[8]), .out(u_csamul_pg_rca24_and11_8));
  fa fa_u_csamul_pg_rca24_fa11_8_out(.a(u_csamul_pg_rca24_and11_8[0]), .b(u_csamul_pg_rca24_fa12_7_xor1[0]), .cin(u_csamul_pg_rca24_fa11_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_8_xor1), .fa_or0(u_csamul_pg_rca24_fa11_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_8(.a(a[12]), .b(b[8]), .out(u_csamul_pg_rca24_and12_8));
  fa fa_u_csamul_pg_rca24_fa12_8_out(.a(u_csamul_pg_rca24_and12_8[0]), .b(u_csamul_pg_rca24_fa13_7_xor1[0]), .cin(u_csamul_pg_rca24_fa12_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_8_xor1), .fa_or0(u_csamul_pg_rca24_fa12_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_8(.a(a[13]), .b(b[8]), .out(u_csamul_pg_rca24_and13_8));
  fa fa_u_csamul_pg_rca24_fa13_8_out(.a(u_csamul_pg_rca24_and13_8[0]), .b(u_csamul_pg_rca24_fa14_7_xor1[0]), .cin(u_csamul_pg_rca24_fa13_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_8_xor1), .fa_or0(u_csamul_pg_rca24_fa13_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_8(.a(a[14]), .b(b[8]), .out(u_csamul_pg_rca24_and14_8));
  fa fa_u_csamul_pg_rca24_fa14_8_out(.a(u_csamul_pg_rca24_and14_8[0]), .b(u_csamul_pg_rca24_fa15_7_xor1[0]), .cin(u_csamul_pg_rca24_fa14_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_8_xor1), .fa_or0(u_csamul_pg_rca24_fa14_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_8(.a(a[15]), .b(b[8]), .out(u_csamul_pg_rca24_and15_8));
  fa fa_u_csamul_pg_rca24_fa15_8_out(.a(u_csamul_pg_rca24_and15_8[0]), .b(u_csamul_pg_rca24_fa16_7_xor1[0]), .cin(u_csamul_pg_rca24_fa15_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_8_xor1), .fa_or0(u_csamul_pg_rca24_fa15_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_8(.a(a[16]), .b(b[8]), .out(u_csamul_pg_rca24_and16_8));
  fa fa_u_csamul_pg_rca24_fa16_8_out(.a(u_csamul_pg_rca24_and16_8[0]), .b(u_csamul_pg_rca24_fa17_7_xor1[0]), .cin(u_csamul_pg_rca24_fa16_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_8_xor1), .fa_or0(u_csamul_pg_rca24_fa16_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_8(.a(a[17]), .b(b[8]), .out(u_csamul_pg_rca24_and17_8));
  fa fa_u_csamul_pg_rca24_fa17_8_out(.a(u_csamul_pg_rca24_and17_8[0]), .b(u_csamul_pg_rca24_fa18_7_xor1[0]), .cin(u_csamul_pg_rca24_fa17_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_8_xor1), .fa_or0(u_csamul_pg_rca24_fa17_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_8(.a(a[18]), .b(b[8]), .out(u_csamul_pg_rca24_and18_8));
  fa fa_u_csamul_pg_rca24_fa18_8_out(.a(u_csamul_pg_rca24_and18_8[0]), .b(u_csamul_pg_rca24_fa19_7_xor1[0]), .cin(u_csamul_pg_rca24_fa18_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_8_xor1), .fa_or0(u_csamul_pg_rca24_fa18_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_8(.a(a[19]), .b(b[8]), .out(u_csamul_pg_rca24_and19_8));
  fa fa_u_csamul_pg_rca24_fa19_8_out(.a(u_csamul_pg_rca24_and19_8[0]), .b(u_csamul_pg_rca24_fa20_7_xor1[0]), .cin(u_csamul_pg_rca24_fa19_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_8_xor1), .fa_or0(u_csamul_pg_rca24_fa19_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_8(.a(a[20]), .b(b[8]), .out(u_csamul_pg_rca24_and20_8));
  fa fa_u_csamul_pg_rca24_fa20_8_out(.a(u_csamul_pg_rca24_and20_8[0]), .b(u_csamul_pg_rca24_fa21_7_xor1[0]), .cin(u_csamul_pg_rca24_fa20_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_8_xor1), .fa_or0(u_csamul_pg_rca24_fa20_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_8(.a(a[21]), .b(b[8]), .out(u_csamul_pg_rca24_and21_8));
  fa fa_u_csamul_pg_rca24_fa21_8_out(.a(u_csamul_pg_rca24_and21_8[0]), .b(u_csamul_pg_rca24_fa22_7_xor1[0]), .cin(u_csamul_pg_rca24_fa21_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_8_xor1), .fa_or0(u_csamul_pg_rca24_fa21_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_8(.a(a[22]), .b(b[8]), .out(u_csamul_pg_rca24_and22_8));
  fa fa_u_csamul_pg_rca24_fa22_8_out(.a(u_csamul_pg_rca24_and22_8[0]), .b(u_csamul_pg_rca24_and23_7[0]), .cin(u_csamul_pg_rca24_fa22_7_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_8_xor1), .fa_or0(u_csamul_pg_rca24_fa22_8_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_8(.a(a[23]), .b(b[8]), .out(u_csamul_pg_rca24_and23_8));
  and_gate and_gate_u_csamul_pg_rca24_and0_9(.a(a[0]), .b(b[9]), .out(u_csamul_pg_rca24_and0_9));
  fa fa_u_csamul_pg_rca24_fa0_9_out(.a(u_csamul_pg_rca24_and0_9[0]), .b(u_csamul_pg_rca24_fa1_8_xor1[0]), .cin(u_csamul_pg_rca24_fa0_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_9_xor1), .fa_or0(u_csamul_pg_rca24_fa0_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_9(.a(a[1]), .b(b[9]), .out(u_csamul_pg_rca24_and1_9));
  fa fa_u_csamul_pg_rca24_fa1_9_out(.a(u_csamul_pg_rca24_and1_9[0]), .b(u_csamul_pg_rca24_fa2_8_xor1[0]), .cin(u_csamul_pg_rca24_fa1_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_9_xor1), .fa_or0(u_csamul_pg_rca24_fa1_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_9(.a(a[2]), .b(b[9]), .out(u_csamul_pg_rca24_and2_9));
  fa fa_u_csamul_pg_rca24_fa2_9_out(.a(u_csamul_pg_rca24_and2_9[0]), .b(u_csamul_pg_rca24_fa3_8_xor1[0]), .cin(u_csamul_pg_rca24_fa2_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_9_xor1), .fa_or0(u_csamul_pg_rca24_fa2_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_9(.a(a[3]), .b(b[9]), .out(u_csamul_pg_rca24_and3_9));
  fa fa_u_csamul_pg_rca24_fa3_9_out(.a(u_csamul_pg_rca24_and3_9[0]), .b(u_csamul_pg_rca24_fa4_8_xor1[0]), .cin(u_csamul_pg_rca24_fa3_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_9_xor1), .fa_or0(u_csamul_pg_rca24_fa3_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_9(.a(a[4]), .b(b[9]), .out(u_csamul_pg_rca24_and4_9));
  fa fa_u_csamul_pg_rca24_fa4_9_out(.a(u_csamul_pg_rca24_and4_9[0]), .b(u_csamul_pg_rca24_fa5_8_xor1[0]), .cin(u_csamul_pg_rca24_fa4_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_9_xor1), .fa_or0(u_csamul_pg_rca24_fa4_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_9(.a(a[5]), .b(b[9]), .out(u_csamul_pg_rca24_and5_9));
  fa fa_u_csamul_pg_rca24_fa5_9_out(.a(u_csamul_pg_rca24_and5_9[0]), .b(u_csamul_pg_rca24_fa6_8_xor1[0]), .cin(u_csamul_pg_rca24_fa5_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_9_xor1), .fa_or0(u_csamul_pg_rca24_fa5_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_9(.a(a[6]), .b(b[9]), .out(u_csamul_pg_rca24_and6_9));
  fa fa_u_csamul_pg_rca24_fa6_9_out(.a(u_csamul_pg_rca24_and6_9[0]), .b(u_csamul_pg_rca24_fa7_8_xor1[0]), .cin(u_csamul_pg_rca24_fa6_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_9_xor1), .fa_or0(u_csamul_pg_rca24_fa6_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_9(.a(a[7]), .b(b[9]), .out(u_csamul_pg_rca24_and7_9));
  fa fa_u_csamul_pg_rca24_fa7_9_out(.a(u_csamul_pg_rca24_and7_9[0]), .b(u_csamul_pg_rca24_fa8_8_xor1[0]), .cin(u_csamul_pg_rca24_fa7_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_9_xor1), .fa_or0(u_csamul_pg_rca24_fa7_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_9(.a(a[8]), .b(b[9]), .out(u_csamul_pg_rca24_and8_9));
  fa fa_u_csamul_pg_rca24_fa8_9_out(.a(u_csamul_pg_rca24_and8_9[0]), .b(u_csamul_pg_rca24_fa9_8_xor1[0]), .cin(u_csamul_pg_rca24_fa8_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_9_xor1), .fa_or0(u_csamul_pg_rca24_fa8_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_9(.a(a[9]), .b(b[9]), .out(u_csamul_pg_rca24_and9_9));
  fa fa_u_csamul_pg_rca24_fa9_9_out(.a(u_csamul_pg_rca24_and9_9[0]), .b(u_csamul_pg_rca24_fa10_8_xor1[0]), .cin(u_csamul_pg_rca24_fa9_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_9_xor1), .fa_or0(u_csamul_pg_rca24_fa9_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_9(.a(a[10]), .b(b[9]), .out(u_csamul_pg_rca24_and10_9));
  fa fa_u_csamul_pg_rca24_fa10_9_out(.a(u_csamul_pg_rca24_and10_9[0]), .b(u_csamul_pg_rca24_fa11_8_xor1[0]), .cin(u_csamul_pg_rca24_fa10_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_9_xor1), .fa_or0(u_csamul_pg_rca24_fa10_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_9(.a(a[11]), .b(b[9]), .out(u_csamul_pg_rca24_and11_9));
  fa fa_u_csamul_pg_rca24_fa11_9_out(.a(u_csamul_pg_rca24_and11_9[0]), .b(u_csamul_pg_rca24_fa12_8_xor1[0]), .cin(u_csamul_pg_rca24_fa11_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_9_xor1), .fa_or0(u_csamul_pg_rca24_fa11_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_9(.a(a[12]), .b(b[9]), .out(u_csamul_pg_rca24_and12_9));
  fa fa_u_csamul_pg_rca24_fa12_9_out(.a(u_csamul_pg_rca24_and12_9[0]), .b(u_csamul_pg_rca24_fa13_8_xor1[0]), .cin(u_csamul_pg_rca24_fa12_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_9_xor1), .fa_or0(u_csamul_pg_rca24_fa12_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_9(.a(a[13]), .b(b[9]), .out(u_csamul_pg_rca24_and13_9));
  fa fa_u_csamul_pg_rca24_fa13_9_out(.a(u_csamul_pg_rca24_and13_9[0]), .b(u_csamul_pg_rca24_fa14_8_xor1[0]), .cin(u_csamul_pg_rca24_fa13_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_9_xor1), .fa_or0(u_csamul_pg_rca24_fa13_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_9(.a(a[14]), .b(b[9]), .out(u_csamul_pg_rca24_and14_9));
  fa fa_u_csamul_pg_rca24_fa14_9_out(.a(u_csamul_pg_rca24_and14_9[0]), .b(u_csamul_pg_rca24_fa15_8_xor1[0]), .cin(u_csamul_pg_rca24_fa14_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_9_xor1), .fa_or0(u_csamul_pg_rca24_fa14_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_9(.a(a[15]), .b(b[9]), .out(u_csamul_pg_rca24_and15_9));
  fa fa_u_csamul_pg_rca24_fa15_9_out(.a(u_csamul_pg_rca24_and15_9[0]), .b(u_csamul_pg_rca24_fa16_8_xor1[0]), .cin(u_csamul_pg_rca24_fa15_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_9_xor1), .fa_or0(u_csamul_pg_rca24_fa15_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_9(.a(a[16]), .b(b[9]), .out(u_csamul_pg_rca24_and16_9));
  fa fa_u_csamul_pg_rca24_fa16_9_out(.a(u_csamul_pg_rca24_and16_9[0]), .b(u_csamul_pg_rca24_fa17_8_xor1[0]), .cin(u_csamul_pg_rca24_fa16_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_9_xor1), .fa_or0(u_csamul_pg_rca24_fa16_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_9(.a(a[17]), .b(b[9]), .out(u_csamul_pg_rca24_and17_9));
  fa fa_u_csamul_pg_rca24_fa17_9_out(.a(u_csamul_pg_rca24_and17_9[0]), .b(u_csamul_pg_rca24_fa18_8_xor1[0]), .cin(u_csamul_pg_rca24_fa17_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_9_xor1), .fa_or0(u_csamul_pg_rca24_fa17_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_9(.a(a[18]), .b(b[9]), .out(u_csamul_pg_rca24_and18_9));
  fa fa_u_csamul_pg_rca24_fa18_9_out(.a(u_csamul_pg_rca24_and18_9[0]), .b(u_csamul_pg_rca24_fa19_8_xor1[0]), .cin(u_csamul_pg_rca24_fa18_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_9_xor1), .fa_or0(u_csamul_pg_rca24_fa18_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_9(.a(a[19]), .b(b[9]), .out(u_csamul_pg_rca24_and19_9));
  fa fa_u_csamul_pg_rca24_fa19_9_out(.a(u_csamul_pg_rca24_and19_9[0]), .b(u_csamul_pg_rca24_fa20_8_xor1[0]), .cin(u_csamul_pg_rca24_fa19_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_9_xor1), .fa_or0(u_csamul_pg_rca24_fa19_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_9(.a(a[20]), .b(b[9]), .out(u_csamul_pg_rca24_and20_9));
  fa fa_u_csamul_pg_rca24_fa20_9_out(.a(u_csamul_pg_rca24_and20_9[0]), .b(u_csamul_pg_rca24_fa21_8_xor1[0]), .cin(u_csamul_pg_rca24_fa20_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_9_xor1), .fa_or0(u_csamul_pg_rca24_fa20_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_9(.a(a[21]), .b(b[9]), .out(u_csamul_pg_rca24_and21_9));
  fa fa_u_csamul_pg_rca24_fa21_9_out(.a(u_csamul_pg_rca24_and21_9[0]), .b(u_csamul_pg_rca24_fa22_8_xor1[0]), .cin(u_csamul_pg_rca24_fa21_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_9_xor1), .fa_or0(u_csamul_pg_rca24_fa21_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_9(.a(a[22]), .b(b[9]), .out(u_csamul_pg_rca24_and22_9));
  fa fa_u_csamul_pg_rca24_fa22_9_out(.a(u_csamul_pg_rca24_and22_9[0]), .b(u_csamul_pg_rca24_and23_8[0]), .cin(u_csamul_pg_rca24_fa22_8_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_9_xor1), .fa_or0(u_csamul_pg_rca24_fa22_9_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_9(.a(a[23]), .b(b[9]), .out(u_csamul_pg_rca24_and23_9));
  and_gate and_gate_u_csamul_pg_rca24_and0_10(.a(a[0]), .b(b[10]), .out(u_csamul_pg_rca24_and0_10));
  fa fa_u_csamul_pg_rca24_fa0_10_out(.a(u_csamul_pg_rca24_and0_10[0]), .b(u_csamul_pg_rca24_fa1_9_xor1[0]), .cin(u_csamul_pg_rca24_fa0_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_10_xor1), .fa_or0(u_csamul_pg_rca24_fa0_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_10(.a(a[1]), .b(b[10]), .out(u_csamul_pg_rca24_and1_10));
  fa fa_u_csamul_pg_rca24_fa1_10_out(.a(u_csamul_pg_rca24_and1_10[0]), .b(u_csamul_pg_rca24_fa2_9_xor1[0]), .cin(u_csamul_pg_rca24_fa1_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_10_xor1), .fa_or0(u_csamul_pg_rca24_fa1_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_10(.a(a[2]), .b(b[10]), .out(u_csamul_pg_rca24_and2_10));
  fa fa_u_csamul_pg_rca24_fa2_10_out(.a(u_csamul_pg_rca24_and2_10[0]), .b(u_csamul_pg_rca24_fa3_9_xor1[0]), .cin(u_csamul_pg_rca24_fa2_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_10_xor1), .fa_or0(u_csamul_pg_rca24_fa2_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_10(.a(a[3]), .b(b[10]), .out(u_csamul_pg_rca24_and3_10));
  fa fa_u_csamul_pg_rca24_fa3_10_out(.a(u_csamul_pg_rca24_and3_10[0]), .b(u_csamul_pg_rca24_fa4_9_xor1[0]), .cin(u_csamul_pg_rca24_fa3_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_10_xor1), .fa_or0(u_csamul_pg_rca24_fa3_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_10(.a(a[4]), .b(b[10]), .out(u_csamul_pg_rca24_and4_10));
  fa fa_u_csamul_pg_rca24_fa4_10_out(.a(u_csamul_pg_rca24_and4_10[0]), .b(u_csamul_pg_rca24_fa5_9_xor1[0]), .cin(u_csamul_pg_rca24_fa4_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_10_xor1), .fa_or0(u_csamul_pg_rca24_fa4_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_10(.a(a[5]), .b(b[10]), .out(u_csamul_pg_rca24_and5_10));
  fa fa_u_csamul_pg_rca24_fa5_10_out(.a(u_csamul_pg_rca24_and5_10[0]), .b(u_csamul_pg_rca24_fa6_9_xor1[0]), .cin(u_csamul_pg_rca24_fa5_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_10_xor1), .fa_or0(u_csamul_pg_rca24_fa5_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_10(.a(a[6]), .b(b[10]), .out(u_csamul_pg_rca24_and6_10));
  fa fa_u_csamul_pg_rca24_fa6_10_out(.a(u_csamul_pg_rca24_and6_10[0]), .b(u_csamul_pg_rca24_fa7_9_xor1[0]), .cin(u_csamul_pg_rca24_fa6_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_10_xor1), .fa_or0(u_csamul_pg_rca24_fa6_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_10(.a(a[7]), .b(b[10]), .out(u_csamul_pg_rca24_and7_10));
  fa fa_u_csamul_pg_rca24_fa7_10_out(.a(u_csamul_pg_rca24_and7_10[0]), .b(u_csamul_pg_rca24_fa8_9_xor1[0]), .cin(u_csamul_pg_rca24_fa7_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_10_xor1), .fa_or0(u_csamul_pg_rca24_fa7_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_10(.a(a[8]), .b(b[10]), .out(u_csamul_pg_rca24_and8_10));
  fa fa_u_csamul_pg_rca24_fa8_10_out(.a(u_csamul_pg_rca24_and8_10[0]), .b(u_csamul_pg_rca24_fa9_9_xor1[0]), .cin(u_csamul_pg_rca24_fa8_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_10_xor1), .fa_or0(u_csamul_pg_rca24_fa8_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_10(.a(a[9]), .b(b[10]), .out(u_csamul_pg_rca24_and9_10));
  fa fa_u_csamul_pg_rca24_fa9_10_out(.a(u_csamul_pg_rca24_and9_10[0]), .b(u_csamul_pg_rca24_fa10_9_xor1[0]), .cin(u_csamul_pg_rca24_fa9_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_10_xor1), .fa_or0(u_csamul_pg_rca24_fa9_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_10(.a(a[10]), .b(b[10]), .out(u_csamul_pg_rca24_and10_10));
  fa fa_u_csamul_pg_rca24_fa10_10_out(.a(u_csamul_pg_rca24_and10_10[0]), .b(u_csamul_pg_rca24_fa11_9_xor1[0]), .cin(u_csamul_pg_rca24_fa10_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_10_xor1), .fa_or0(u_csamul_pg_rca24_fa10_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_10(.a(a[11]), .b(b[10]), .out(u_csamul_pg_rca24_and11_10));
  fa fa_u_csamul_pg_rca24_fa11_10_out(.a(u_csamul_pg_rca24_and11_10[0]), .b(u_csamul_pg_rca24_fa12_9_xor1[0]), .cin(u_csamul_pg_rca24_fa11_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_10_xor1), .fa_or0(u_csamul_pg_rca24_fa11_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_10(.a(a[12]), .b(b[10]), .out(u_csamul_pg_rca24_and12_10));
  fa fa_u_csamul_pg_rca24_fa12_10_out(.a(u_csamul_pg_rca24_and12_10[0]), .b(u_csamul_pg_rca24_fa13_9_xor1[0]), .cin(u_csamul_pg_rca24_fa12_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_10_xor1), .fa_or0(u_csamul_pg_rca24_fa12_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_10(.a(a[13]), .b(b[10]), .out(u_csamul_pg_rca24_and13_10));
  fa fa_u_csamul_pg_rca24_fa13_10_out(.a(u_csamul_pg_rca24_and13_10[0]), .b(u_csamul_pg_rca24_fa14_9_xor1[0]), .cin(u_csamul_pg_rca24_fa13_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_10_xor1), .fa_or0(u_csamul_pg_rca24_fa13_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_10(.a(a[14]), .b(b[10]), .out(u_csamul_pg_rca24_and14_10));
  fa fa_u_csamul_pg_rca24_fa14_10_out(.a(u_csamul_pg_rca24_and14_10[0]), .b(u_csamul_pg_rca24_fa15_9_xor1[0]), .cin(u_csamul_pg_rca24_fa14_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_10_xor1), .fa_or0(u_csamul_pg_rca24_fa14_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_10(.a(a[15]), .b(b[10]), .out(u_csamul_pg_rca24_and15_10));
  fa fa_u_csamul_pg_rca24_fa15_10_out(.a(u_csamul_pg_rca24_and15_10[0]), .b(u_csamul_pg_rca24_fa16_9_xor1[0]), .cin(u_csamul_pg_rca24_fa15_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_10_xor1), .fa_or0(u_csamul_pg_rca24_fa15_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_10(.a(a[16]), .b(b[10]), .out(u_csamul_pg_rca24_and16_10));
  fa fa_u_csamul_pg_rca24_fa16_10_out(.a(u_csamul_pg_rca24_and16_10[0]), .b(u_csamul_pg_rca24_fa17_9_xor1[0]), .cin(u_csamul_pg_rca24_fa16_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_10_xor1), .fa_or0(u_csamul_pg_rca24_fa16_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_10(.a(a[17]), .b(b[10]), .out(u_csamul_pg_rca24_and17_10));
  fa fa_u_csamul_pg_rca24_fa17_10_out(.a(u_csamul_pg_rca24_and17_10[0]), .b(u_csamul_pg_rca24_fa18_9_xor1[0]), .cin(u_csamul_pg_rca24_fa17_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_10_xor1), .fa_or0(u_csamul_pg_rca24_fa17_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_10(.a(a[18]), .b(b[10]), .out(u_csamul_pg_rca24_and18_10));
  fa fa_u_csamul_pg_rca24_fa18_10_out(.a(u_csamul_pg_rca24_and18_10[0]), .b(u_csamul_pg_rca24_fa19_9_xor1[0]), .cin(u_csamul_pg_rca24_fa18_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_10_xor1), .fa_or0(u_csamul_pg_rca24_fa18_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_10(.a(a[19]), .b(b[10]), .out(u_csamul_pg_rca24_and19_10));
  fa fa_u_csamul_pg_rca24_fa19_10_out(.a(u_csamul_pg_rca24_and19_10[0]), .b(u_csamul_pg_rca24_fa20_9_xor1[0]), .cin(u_csamul_pg_rca24_fa19_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_10_xor1), .fa_or0(u_csamul_pg_rca24_fa19_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_10(.a(a[20]), .b(b[10]), .out(u_csamul_pg_rca24_and20_10));
  fa fa_u_csamul_pg_rca24_fa20_10_out(.a(u_csamul_pg_rca24_and20_10[0]), .b(u_csamul_pg_rca24_fa21_9_xor1[0]), .cin(u_csamul_pg_rca24_fa20_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_10_xor1), .fa_or0(u_csamul_pg_rca24_fa20_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_10(.a(a[21]), .b(b[10]), .out(u_csamul_pg_rca24_and21_10));
  fa fa_u_csamul_pg_rca24_fa21_10_out(.a(u_csamul_pg_rca24_and21_10[0]), .b(u_csamul_pg_rca24_fa22_9_xor1[0]), .cin(u_csamul_pg_rca24_fa21_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_10_xor1), .fa_or0(u_csamul_pg_rca24_fa21_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_10(.a(a[22]), .b(b[10]), .out(u_csamul_pg_rca24_and22_10));
  fa fa_u_csamul_pg_rca24_fa22_10_out(.a(u_csamul_pg_rca24_and22_10[0]), .b(u_csamul_pg_rca24_and23_9[0]), .cin(u_csamul_pg_rca24_fa22_9_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_10_xor1), .fa_or0(u_csamul_pg_rca24_fa22_10_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_10(.a(a[23]), .b(b[10]), .out(u_csamul_pg_rca24_and23_10));
  and_gate and_gate_u_csamul_pg_rca24_and0_11(.a(a[0]), .b(b[11]), .out(u_csamul_pg_rca24_and0_11));
  fa fa_u_csamul_pg_rca24_fa0_11_out(.a(u_csamul_pg_rca24_and0_11[0]), .b(u_csamul_pg_rca24_fa1_10_xor1[0]), .cin(u_csamul_pg_rca24_fa0_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_11_xor1), .fa_or0(u_csamul_pg_rca24_fa0_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_11(.a(a[1]), .b(b[11]), .out(u_csamul_pg_rca24_and1_11));
  fa fa_u_csamul_pg_rca24_fa1_11_out(.a(u_csamul_pg_rca24_and1_11[0]), .b(u_csamul_pg_rca24_fa2_10_xor1[0]), .cin(u_csamul_pg_rca24_fa1_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_11_xor1), .fa_or0(u_csamul_pg_rca24_fa1_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_11(.a(a[2]), .b(b[11]), .out(u_csamul_pg_rca24_and2_11));
  fa fa_u_csamul_pg_rca24_fa2_11_out(.a(u_csamul_pg_rca24_and2_11[0]), .b(u_csamul_pg_rca24_fa3_10_xor1[0]), .cin(u_csamul_pg_rca24_fa2_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_11_xor1), .fa_or0(u_csamul_pg_rca24_fa2_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_11(.a(a[3]), .b(b[11]), .out(u_csamul_pg_rca24_and3_11));
  fa fa_u_csamul_pg_rca24_fa3_11_out(.a(u_csamul_pg_rca24_and3_11[0]), .b(u_csamul_pg_rca24_fa4_10_xor1[0]), .cin(u_csamul_pg_rca24_fa3_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_11_xor1), .fa_or0(u_csamul_pg_rca24_fa3_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_11(.a(a[4]), .b(b[11]), .out(u_csamul_pg_rca24_and4_11));
  fa fa_u_csamul_pg_rca24_fa4_11_out(.a(u_csamul_pg_rca24_and4_11[0]), .b(u_csamul_pg_rca24_fa5_10_xor1[0]), .cin(u_csamul_pg_rca24_fa4_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_11_xor1), .fa_or0(u_csamul_pg_rca24_fa4_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_11(.a(a[5]), .b(b[11]), .out(u_csamul_pg_rca24_and5_11));
  fa fa_u_csamul_pg_rca24_fa5_11_out(.a(u_csamul_pg_rca24_and5_11[0]), .b(u_csamul_pg_rca24_fa6_10_xor1[0]), .cin(u_csamul_pg_rca24_fa5_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_11_xor1), .fa_or0(u_csamul_pg_rca24_fa5_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_11(.a(a[6]), .b(b[11]), .out(u_csamul_pg_rca24_and6_11));
  fa fa_u_csamul_pg_rca24_fa6_11_out(.a(u_csamul_pg_rca24_and6_11[0]), .b(u_csamul_pg_rca24_fa7_10_xor1[0]), .cin(u_csamul_pg_rca24_fa6_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_11_xor1), .fa_or0(u_csamul_pg_rca24_fa6_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_11(.a(a[7]), .b(b[11]), .out(u_csamul_pg_rca24_and7_11));
  fa fa_u_csamul_pg_rca24_fa7_11_out(.a(u_csamul_pg_rca24_and7_11[0]), .b(u_csamul_pg_rca24_fa8_10_xor1[0]), .cin(u_csamul_pg_rca24_fa7_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_11_xor1), .fa_or0(u_csamul_pg_rca24_fa7_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_11(.a(a[8]), .b(b[11]), .out(u_csamul_pg_rca24_and8_11));
  fa fa_u_csamul_pg_rca24_fa8_11_out(.a(u_csamul_pg_rca24_and8_11[0]), .b(u_csamul_pg_rca24_fa9_10_xor1[0]), .cin(u_csamul_pg_rca24_fa8_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_11_xor1), .fa_or0(u_csamul_pg_rca24_fa8_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_11(.a(a[9]), .b(b[11]), .out(u_csamul_pg_rca24_and9_11));
  fa fa_u_csamul_pg_rca24_fa9_11_out(.a(u_csamul_pg_rca24_and9_11[0]), .b(u_csamul_pg_rca24_fa10_10_xor1[0]), .cin(u_csamul_pg_rca24_fa9_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_11_xor1), .fa_or0(u_csamul_pg_rca24_fa9_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_11(.a(a[10]), .b(b[11]), .out(u_csamul_pg_rca24_and10_11));
  fa fa_u_csamul_pg_rca24_fa10_11_out(.a(u_csamul_pg_rca24_and10_11[0]), .b(u_csamul_pg_rca24_fa11_10_xor1[0]), .cin(u_csamul_pg_rca24_fa10_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_11_xor1), .fa_or0(u_csamul_pg_rca24_fa10_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_11(.a(a[11]), .b(b[11]), .out(u_csamul_pg_rca24_and11_11));
  fa fa_u_csamul_pg_rca24_fa11_11_out(.a(u_csamul_pg_rca24_and11_11[0]), .b(u_csamul_pg_rca24_fa12_10_xor1[0]), .cin(u_csamul_pg_rca24_fa11_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_11_xor1), .fa_or0(u_csamul_pg_rca24_fa11_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_11(.a(a[12]), .b(b[11]), .out(u_csamul_pg_rca24_and12_11));
  fa fa_u_csamul_pg_rca24_fa12_11_out(.a(u_csamul_pg_rca24_and12_11[0]), .b(u_csamul_pg_rca24_fa13_10_xor1[0]), .cin(u_csamul_pg_rca24_fa12_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_11_xor1), .fa_or0(u_csamul_pg_rca24_fa12_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_11(.a(a[13]), .b(b[11]), .out(u_csamul_pg_rca24_and13_11));
  fa fa_u_csamul_pg_rca24_fa13_11_out(.a(u_csamul_pg_rca24_and13_11[0]), .b(u_csamul_pg_rca24_fa14_10_xor1[0]), .cin(u_csamul_pg_rca24_fa13_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_11_xor1), .fa_or0(u_csamul_pg_rca24_fa13_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_11(.a(a[14]), .b(b[11]), .out(u_csamul_pg_rca24_and14_11));
  fa fa_u_csamul_pg_rca24_fa14_11_out(.a(u_csamul_pg_rca24_and14_11[0]), .b(u_csamul_pg_rca24_fa15_10_xor1[0]), .cin(u_csamul_pg_rca24_fa14_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_11_xor1), .fa_or0(u_csamul_pg_rca24_fa14_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_11(.a(a[15]), .b(b[11]), .out(u_csamul_pg_rca24_and15_11));
  fa fa_u_csamul_pg_rca24_fa15_11_out(.a(u_csamul_pg_rca24_and15_11[0]), .b(u_csamul_pg_rca24_fa16_10_xor1[0]), .cin(u_csamul_pg_rca24_fa15_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_11_xor1), .fa_or0(u_csamul_pg_rca24_fa15_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_11(.a(a[16]), .b(b[11]), .out(u_csamul_pg_rca24_and16_11));
  fa fa_u_csamul_pg_rca24_fa16_11_out(.a(u_csamul_pg_rca24_and16_11[0]), .b(u_csamul_pg_rca24_fa17_10_xor1[0]), .cin(u_csamul_pg_rca24_fa16_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_11_xor1), .fa_or0(u_csamul_pg_rca24_fa16_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_11(.a(a[17]), .b(b[11]), .out(u_csamul_pg_rca24_and17_11));
  fa fa_u_csamul_pg_rca24_fa17_11_out(.a(u_csamul_pg_rca24_and17_11[0]), .b(u_csamul_pg_rca24_fa18_10_xor1[0]), .cin(u_csamul_pg_rca24_fa17_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_11_xor1), .fa_or0(u_csamul_pg_rca24_fa17_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_11(.a(a[18]), .b(b[11]), .out(u_csamul_pg_rca24_and18_11));
  fa fa_u_csamul_pg_rca24_fa18_11_out(.a(u_csamul_pg_rca24_and18_11[0]), .b(u_csamul_pg_rca24_fa19_10_xor1[0]), .cin(u_csamul_pg_rca24_fa18_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_11_xor1), .fa_or0(u_csamul_pg_rca24_fa18_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_11(.a(a[19]), .b(b[11]), .out(u_csamul_pg_rca24_and19_11));
  fa fa_u_csamul_pg_rca24_fa19_11_out(.a(u_csamul_pg_rca24_and19_11[0]), .b(u_csamul_pg_rca24_fa20_10_xor1[0]), .cin(u_csamul_pg_rca24_fa19_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_11_xor1), .fa_or0(u_csamul_pg_rca24_fa19_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_11(.a(a[20]), .b(b[11]), .out(u_csamul_pg_rca24_and20_11));
  fa fa_u_csamul_pg_rca24_fa20_11_out(.a(u_csamul_pg_rca24_and20_11[0]), .b(u_csamul_pg_rca24_fa21_10_xor1[0]), .cin(u_csamul_pg_rca24_fa20_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_11_xor1), .fa_or0(u_csamul_pg_rca24_fa20_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_11(.a(a[21]), .b(b[11]), .out(u_csamul_pg_rca24_and21_11));
  fa fa_u_csamul_pg_rca24_fa21_11_out(.a(u_csamul_pg_rca24_and21_11[0]), .b(u_csamul_pg_rca24_fa22_10_xor1[0]), .cin(u_csamul_pg_rca24_fa21_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_11_xor1), .fa_or0(u_csamul_pg_rca24_fa21_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_11(.a(a[22]), .b(b[11]), .out(u_csamul_pg_rca24_and22_11));
  fa fa_u_csamul_pg_rca24_fa22_11_out(.a(u_csamul_pg_rca24_and22_11[0]), .b(u_csamul_pg_rca24_and23_10[0]), .cin(u_csamul_pg_rca24_fa22_10_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_11_xor1), .fa_or0(u_csamul_pg_rca24_fa22_11_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_11(.a(a[23]), .b(b[11]), .out(u_csamul_pg_rca24_and23_11));
  and_gate and_gate_u_csamul_pg_rca24_and0_12(.a(a[0]), .b(b[12]), .out(u_csamul_pg_rca24_and0_12));
  fa fa_u_csamul_pg_rca24_fa0_12_out(.a(u_csamul_pg_rca24_and0_12[0]), .b(u_csamul_pg_rca24_fa1_11_xor1[0]), .cin(u_csamul_pg_rca24_fa0_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_12_xor1), .fa_or0(u_csamul_pg_rca24_fa0_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_12(.a(a[1]), .b(b[12]), .out(u_csamul_pg_rca24_and1_12));
  fa fa_u_csamul_pg_rca24_fa1_12_out(.a(u_csamul_pg_rca24_and1_12[0]), .b(u_csamul_pg_rca24_fa2_11_xor1[0]), .cin(u_csamul_pg_rca24_fa1_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_12_xor1), .fa_or0(u_csamul_pg_rca24_fa1_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_12(.a(a[2]), .b(b[12]), .out(u_csamul_pg_rca24_and2_12));
  fa fa_u_csamul_pg_rca24_fa2_12_out(.a(u_csamul_pg_rca24_and2_12[0]), .b(u_csamul_pg_rca24_fa3_11_xor1[0]), .cin(u_csamul_pg_rca24_fa2_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_12_xor1), .fa_or0(u_csamul_pg_rca24_fa2_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_12(.a(a[3]), .b(b[12]), .out(u_csamul_pg_rca24_and3_12));
  fa fa_u_csamul_pg_rca24_fa3_12_out(.a(u_csamul_pg_rca24_and3_12[0]), .b(u_csamul_pg_rca24_fa4_11_xor1[0]), .cin(u_csamul_pg_rca24_fa3_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_12_xor1), .fa_or0(u_csamul_pg_rca24_fa3_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_12(.a(a[4]), .b(b[12]), .out(u_csamul_pg_rca24_and4_12));
  fa fa_u_csamul_pg_rca24_fa4_12_out(.a(u_csamul_pg_rca24_and4_12[0]), .b(u_csamul_pg_rca24_fa5_11_xor1[0]), .cin(u_csamul_pg_rca24_fa4_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_12_xor1), .fa_or0(u_csamul_pg_rca24_fa4_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_12(.a(a[5]), .b(b[12]), .out(u_csamul_pg_rca24_and5_12));
  fa fa_u_csamul_pg_rca24_fa5_12_out(.a(u_csamul_pg_rca24_and5_12[0]), .b(u_csamul_pg_rca24_fa6_11_xor1[0]), .cin(u_csamul_pg_rca24_fa5_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_12_xor1), .fa_or0(u_csamul_pg_rca24_fa5_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_12(.a(a[6]), .b(b[12]), .out(u_csamul_pg_rca24_and6_12));
  fa fa_u_csamul_pg_rca24_fa6_12_out(.a(u_csamul_pg_rca24_and6_12[0]), .b(u_csamul_pg_rca24_fa7_11_xor1[0]), .cin(u_csamul_pg_rca24_fa6_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_12_xor1), .fa_or0(u_csamul_pg_rca24_fa6_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_12(.a(a[7]), .b(b[12]), .out(u_csamul_pg_rca24_and7_12));
  fa fa_u_csamul_pg_rca24_fa7_12_out(.a(u_csamul_pg_rca24_and7_12[0]), .b(u_csamul_pg_rca24_fa8_11_xor1[0]), .cin(u_csamul_pg_rca24_fa7_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_12_xor1), .fa_or0(u_csamul_pg_rca24_fa7_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_12(.a(a[8]), .b(b[12]), .out(u_csamul_pg_rca24_and8_12));
  fa fa_u_csamul_pg_rca24_fa8_12_out(.a(u_csamul_pg_rca24_and8_12[0]), .b(u_csamul_pg_rca24_fa9_11_xor1[0]), .cin(u_csamul_pg_rca24_fa8_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_12_xor1), .fa_or0(u_csamul_pg_rca24_fa8_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_12(.a(a[9]), .b(b[12]), .out(u_csamul_pg_rca24_and9_12));
  fa fa_u_csamul_pg_rca24_fa9_12_out(.a(u_csamul_pg_rca24_and9_12[0]), .b(u_csamul_pg_rca24_fa10_11_xor1[0]), .cin(u_csamul_pg_rca24_fa9_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_12_xor1), .fa_or0(u_csamul_pg_rca24_fa9_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_12(.a(a[10]), .b(b[12]), .out(u_csamul_pg_rca24_and10_12));
  fa fa_u_csamul_pg_rca24_fa10_12_out(.a(u_csamul_pg_rca24_and10_12[0]), .b(u_csamul_pg_rca24_fa11_11_xor1[0]), .cin(u_csamul_pg_rca24_fa10_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_12_xor1), .fa_or0(u_csamul_pg_rca24_fa10_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_12(.a(a[11]), .b(b[12]), .out(u_csamul_pg_rca24_and11_12));
  fa fa_u_csamul_pg_rca24_fa11_12_out(.a(u_csamul_pg_rca24_and11_12[0]), .b(u_csamul_pg_rca24_fa12_11_xor1[0]), .cin(u_csamul_pg_rca24_fa11_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_12_xor1), .fa_or0(u_csamul_pg_rca24_fa11_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_12(.a(a[12]), .b(b[12]), .out(u_csamul_pg_rca24_and12_12));
  fa fa_u_csamul_pg_rca24_fa12_12_out(.a(u_csamul_pg_rca24_and12_12[0]), .b(u_csamul_pg_rca24_fa13_11_xor1[0]), .cin(u_csamul_pg_rca24_fa12_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_12_xor1), .fa_or0(u_csamul_pg_rca24_fa12_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_12(.a(a[13]), .b(b[12]), .out(u_csamul_pg_rca24_and13_12));
  fa fa_u_csamul_pg_rca24_fa13_12_out(.a(u_csamul_pg_rca24_and13_12[0]), .b(u_csamul_pg_rca24_fa14_11_xor1[0]), .cin(u_csamul_pg_rca24_fa13_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_12_xor1), .fa_or0(u_csamul_pg_rca24_fa13_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_12(.a(a[14]), .b(b[12]), .out(u_csamul_pg_rca24_and14_12));
  fa fa_u_csamul_pg_rca24_fa14_12_out(.a(u_csamul_pg_rca24_and14_12[0]), .b(u_csamul_pg_rca24_fa15_11_xor1[0]), .cin(u_csamul_pg_rca24_fa14_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_12_xor1), .fa_or0(u_csamul_pg_rca24_fa14_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_12(.a(a[15]), .b(b[12]), .out(u_csamul_pg_rca24_and15_12));
  fa fa_u_csamul_pg_rca24_fa15_12_out(.a(u_csamul_pg_rca24_and15_12[0]), .b(u_csamul_pg_rca24_fa16_11_xor1[0]), .cin(u_csamul_pg_rca24_fa15_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_12_xor1), .fa_or0(u_csamul_pg_rca24_fa15_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_12(.a(a[16]), .b(b[12]), .out(u_csamul_pg_rca24_and16_12));
  fa fa_u_csamul_pg_rca24_fa16_12_out(.a(u_csamul_pg_rca24_and16_12[0]), .b(u_csamul_pg_rca24_fa17_11_xor1[0]), .cin(u_csamul_pg_rca24_fa16_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_12_xor1), .fa_or0(u_csamul_pg_rca24_fa16_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_12(.a(a[17]), .b(b[12]), .out(u_csamul_pg_rca24_and17_12));
  fa fa_u_csamul_pg_rca24_fa17_12_out(.a(u_csamul_pg_rca24_and17_12[0]), .b(u_csamul_pg_rca24_fa18_11_xor1[0]), .cin(u_csamul_pg_rca24_fa17_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_12_xor1), .fa_or0(u_csamul_pg_rca24_fa17_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_12(.a(a[18]), .b(b[12]), .out(u_csamul_pg_rca24_and18_12));
  fa fa_u_csamul_pg_rca24_fa18_12_out(.a(u_csamul_pg_rca24_and18_12[0]), .b(u_csamul_pg_rca24_fa19_11_xor1[0]), .cin(u_csamul_pg_rca24_fa18_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_12_xor1), .fa_or0(u_csamul_pg_rca24_fa18_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_12(.a(a[19]), .b(b[12]), .out(u_csamul_pg_rca24_and19_12));
  fa fa_u_csamul_pg_rca24_fa19_12_out(.a(u_csamul_pg_rca24_and19_12[0]), .b(u_csamul_pg_rca24_fa20_11_xor1[0]), .cin(u_csamul_pg_rca24_fa19_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_12_xor1), .fa_or0(u_csamul_pg_rca24_fa19_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_12(.a(a[20]), .b(b[12]), .out(u_csamul_pg_rca24_and20_12));
  fa fa_u_csamul_pg_rca24_fa20_12_out(.a(u_csamul_pg_rca24_and20_12[0]), .b(u_csamul_pg_rca24_fa21_11_xor1[0]), .cin(u_csamul_pg_rca24_fa20_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_12_xor1), .fa_or0(u_csamul_pg_rca24_fa20_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_12(.a(a[21]), .b(b[12]), .out(u_csamul_pg_rca24_and21_12));
  fa fa_u_csamul_pg_rca24_fa21_12_out(.a(u_csamul_pg_rca24_and21_12[0]), .b(u_csamul_pg_rca24_fa22_11_xor1[0]), .cin(u_csamul_pg_rca24_fa21_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_12_xor1), .fa_or0(u_csamul_pg_rca24_fa21_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_12(.a(a[22]), .b(b[12]), .out(u_csamul_pg_rca24_and22_12));
  fa fa_u_csamul_pg_rca24_fa22_12_out(.a(u_csamul_pg_rca24_and22_12[0]), .b(u_csamul_pg_rca24_and23_11[0]), .cin(u_csamul_pg_rca24_fa22_11_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_12_xor1), .fa_or0(u_csamul_pg_rca24_fa22_12_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_12(.a(a[23]), .b(b[12]), .out(u_csamul_pg_rca24_and23_12));
  and_gate and_gate_u_csamul_pg_rca24_and0_13(.a(a[0]), .b(b[13]), .out(u_csamul_pg_rca24_and0_13));
  fa fa_u_csamul_pg_rca24_fa0_13_out(.a(u_csamul_pg_rca24_and0_13[0]), .b(u_csamul_pg_rca24_fa1_12_xor1[0]), .cin(u_csamul_pg_rca24_fa0_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_13_xor1), .fa_or0(u_csamul_pg_rca24_fa0_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_13(.a(a[1]), .b(b[13]), .out(u_csamul_pg_rca24_and1_13));
  fa fa_u_csamul_pg_rca24_fa1_13_out(.a(u_csamul_pg_rca24_and1_13[0]), .b(u_csamul_pg_rca24_fa2_12_xor1[0]), .cin(u_csamul_pg_rca24_fa1_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_13_xor1), .fa_or0(u_csamul_pg_rca24_fa1_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_13(.a(a[2]), .b(b[13]), .out(u_csamul_pg_rca24_and2_13));
  fa fa_u_csamul_pg_rca24_fa2_13_out(.a(u_csamul_pg_rca24_and2_13[0]), .b(u_csamul_pg_rca24_fa3_12_xor1[0]), .cin(u_csamul_pg_rca24_fa2_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_13_xor1), .fa_or0(u_csamul_pg_rca24_fa2_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_13(.a(a[3]), .b(b[13]), .out(u_csamul_pg_rca24_and3_13));
  fa fa_u_csamul_pg_rca24_fa3_13_out(.a(u_csamul_pg_rca24_and3_13[0]), .b(u_csamul_pg_rca24_fa4_12_xor1[0]), .cin(u_csamul_pg_rca24_fa3_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_13_xor1), .fa_or0(u_csamul_pg_rca24_fa3_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_13(.a(a[4]), .b(b[13]), .out(u_csamul_pg_rca24_and4_13));
  fa fa_u_csamul_pg_rca24_fa4_13_out(.a(u_csamul_pg_rca24_and4_13[0]), .b(u_csamul_pg_rca24_fa5_12_xor1[0]), .cin(u_csamul_pg_rca24_fa4_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_13_xor1), .fa_or0(u_csamul_pg_rca24_fa4_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_13(.a(a[5]), .b(b[13]), .out(u_csamul_pg_rca24_and5_13));
  fa fa_u_csamul_pg_rca24_fa5_13_out(.a(u_csamul_pg_rca24_and5_13[0]), .b(u_csamul_pg_rca24_fa6_12_xor1[0]), .cin(u_csamul_pg_rca24_fa5_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_13_xor1), .fa_or0(u_csamul_pg_rca24_fa5_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_13(.a(a[6]), .b(b[13]), .out(u_csamul_pg_rca24_and6_13));
  fa fa_u_csamul_pg_rca24_fa6_13_out(.a(u_csamul_pg_rca24_and6_13[0]), .b(u_csamul_pg_rca24_fa7_12_xor1[0]), .cin(u_csamul_pg_rca24_fa6_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_13_xor1), .fa_or0(u_csamul_pg_rca24_fa6_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_13(.a(a[7]), .b(b[13]), .out(u_csamul_pg_rca24_and7_13));
  fa fa_u_csamul_pg_rca24_fa7_13_out(.a(u_csamul_pg_rca24_and7_13[0]), .b(u_csamul_pg_rca24_fa8_12_xor1[0]), .cin(u_csamul_pg_rca24_fa7_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_13_xor1), .fa_or0(u_csamul_pg_rca24_fa7_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_13(.a(a[8]), .b(b[13]), .out(u_csamul_pg_rca24_and8_13));
  fa fa_u_csamul_pg_rca24_fa8_13_out(.a(u_csamul_pg_rca24_and8_13[0]), .b(u_csamul_pg_rca24_fa9_12_xor1[0]), .cin(u_csamul_pg_rca24_fa8_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_13_xor1), .fa_or0(u_csamul_pg_rca24_fa8_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_13(.a(a[9]), .b(b[13]), .out(u_csamul_pg_rca24_and9_13));
  fa fa_u_csamul_pg_rca24_fa9_13_out(.a(u_csamul_pg_rca24_and9_13[0]), .b(u_csamul_pg_rca24_fa10_12_xor1[0]), .cin(u_csamul_pg_rca24_fa9_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_13_xor1), .fa_or0(u_csamul_pg_rca24_fa9_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_13(.a(a[10]), .b(b[13]), .out(u_csamul_pg_rca24_and10_13));
  fa fa_u_csamul_pg_rca24_fa10_13_out(.a(u_csamul_pg_rca24_and10_13[0]), .b(u_csamul_pg_rca24_fa11_12_xor1[0]), .cin(u_csamul_pg_rca24_fa10_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_13_xor1), .fa_or0(u_csamul_pg_rca24_fa10_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_13(.a(a[11]), .b(b[13]), .out(u_csamul_pg_rca24_and11_13));
  fa fa_u_csamul_pg_rca24_fa11_13_out(.a(u_csamul_pg_rca24_and11_13[0]), .b(u_csamul_pg_rca24_fa12_12_xor1[0]), .cin(u_csamul_pg_rca24_fa11_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_13_xor1), .fa_or0(u_csamul_pg_rca24_fa11_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_13(.a(a[12]), .b(b[13]), .out(u_csamul_pg_rca24_and12_13));
  fa fa_u_csamul_pg_rca24_fa12_13_out(.a(u_csamul_pg_rca24_and12_13[0]), .b(u_csamul_pg_rca24_fa13_12_xor1[0]), .cin(u_csamul_pg_rca24_fa12_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_13_xor1), .fa_or0(u_csamul_pg_rca24_fa12_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_13(.a(a[13]), .b(b[13]), .out(u_csamul_pg_rca24_and13_13));
  fa fa_u_csamul_pg_rca24_fa13_13_out(.a(u_csamul_pg_rca24_and13_13[0]), .b(u_csamul_pg_rca24_fa14_12_xor1[0]), .cin(u_csamul_pg_rca24_fa13_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_13_xor1), .fa_or0(u_csamul_pg_rca24_fa13_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_13(.a(a[14]), .b(b[13]), .out(u_csamul_pg_rca24_and14_13));
  fa fa_u_csamul_pg_rca24_fa14_13_out(.a(u_csamul_pg_rca24_and14_13[0]), .b(u_csamul_pg_rca24_fa15_12_xor1[0]), .cin(u_csamul_pg_rca24_fa14_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_13_xor1), .fa_or0(u_csamul_pg_rca24_fa14_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_13(.a(a[15]), .b(b[13]), .out(u_csamul_pg_rca24_and15_13));
  fa fa_u_csamul_pg_rca24_fa15_13_out(.a(u_csamul_pg_rca24_and15_13[0]), .b(u_csamul_pg_rca24_fa16_12_xor1[0]), .cin(u_csamul_pg_rca24_fa15_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_13_xor1), .fa_or0(u_csamul_pg_rca24_fa15_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_13(.a(a[16]), .b(b[13]), .out(u_csamul_pg_rca24_and16_13));
  fa fa_u_csamul_pg_rca24_fa16_13_out(.a(u_csamul_pg_rca24_and16_13[0]), .b(u_csamul_pg_rca24_fa17_12_xor1[0]), .cin(u_csamul_pg_rca24_fa16_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_13_xor1), .fa_or0(u_csamul_pg_rca24_fa16_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_13(.a(a[17]), .b(b[13]), .out(u_csamul_pg_rca24_and17_13));
  fa fa_u_csamul_pg_rca24_fa17_13_out(.a(u_csamul_pg_rca24_and17_13[0]), .b(u_csamul_pg_rca24_fa18_12_xor1[0]), .cin(u_csamul_pg_rca24_fa17_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_13_xor1), .fa_or0(u_csamul_pg_rca24_fa17_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_13(.a(a[18]), .b(b[13]), .out(u_csamul_pg_rca24_and18_13));
  fa fa_u_csamul_pg_rca24_fa18_13_out(.a(u_csamul_pg_rca24_and18_13[0]), .b(u_csamul_pg_rca24_fa19_12_xor1[0]), .cin(u_csamul_pg_rca24_fa18_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_13_xor1), .fa_or0(u_csamul_pg_rca24_fa18_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_13(.a(a[19]), .b(b[13]), .out(u_csamul_pg_rca24_and19_13));
  fa fa_u_csamul_pg_rca24_fa19_13_out(.a(u_csamul_pg_rca24_and19_13[0]), .b(u_csamul_pg_rca24_fa20_12_xor1[0]), .cin(u_csamul_pg_rca24_fa19_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_13_xor1), .fa_or0(u_csamul_pg_rca24_fa19_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_13(.a(a[20]), .b(b[13]), .out(u_csamul_pg_rca24_and20_13));
  fa fa_u_csamul_pg_rca24_fa20_13_out(.a(u_csamul_pg_rca24_and20_13[0]), .b(u_csamul_pg_rca24_fa21_12_xor1[0]), .cin(u_csamul_pg_rca24_fa20_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_13_xor1), .fa_or0(u_csamul_pg_rca24_fa20_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_13(.a(a[21]), .b(b[13]), .out(u_csamul_pg_rca24_and21_13));
  fa fa_u_csamul_pg_rca24_fa21_13_out(.a(u_csamul_pg_rca24_and21_13[0]), .b(u_csamul_pg_rca24_fa22_12_xor1[0]), .cin(u_csamul_pg_rca24_fa21_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_13_xor1), .fa_or0(u_csamul_pg_rca24_fa21_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_13(.a(a[22]), .b(b[13]), .out(u_csamul_pg_rca24_and22_13));
  fa fa_u_csamul_pg_rca24_fa22_13_out(.a(u_csamul_pg_rca24_and22_13[0]), .b(u_csamul_pg_rca24_and23_12[0]), .cin(u_csamul_pg_rca24_fa22_12_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_13_xor1), .fa_or0(u_csamul_pg_rca24_fa22_13_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_13(.a(a[23]), .b(b[13]), .out(u_csamul_pg_rca24_and23_13));
  and_gate and_gate_u_csamul_pg_rca24_and0_14(.a(a[0]), .b(b[14]), .out(u_csamul_pg_rca24_and0_14));
  fa fa_u_csamul_pg_rca24_fa0_14_out(.a(u_csamul_pg_rca24_and0_14[0]), .b(u_csamul_pg_rca24_fa1_13_xor1[0]), .cin(u_csamul_pg_rca24_fa0_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_14_xor1), .fa_or0(u_csamul_pg_rca24_fa0_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_14(.a(a[1]), .b(b[14]), .out(u_csamul_pg_rca24_and1_14));
  fa fa_u_csamul_pg_rca24_fa1_14_out(.a(u_csamul_pg_rca24_and1_14[0]), .b(u_csamul_pg_rca24_fa2_13_xor1[0]), .cin(u_csamul_pg_rca24_fa1_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_14_xor1), .fa_or0(u_csamul_pg_rca24_fa1_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_14(.a(a[2]), .b(b[14]), .out(u_csamul_pg_rca24_and2_14));
  fa fa_u_csamul_pg_rca24_fa2_14_out(.a(u_csamul_pg_rca24_and2_14[0]), .b(u_csamul_pg_rca24_fa3_13_xor1[0]), .cin(u_csamul_pg_rca24_fa2_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_14_xor1), .fa_or0(u_csamul_pg_rca24_fa2_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_14(.a(a[3]), .b(b[14]), .out(u_csamul_pg_rca24_and3_14));
  fa fa_u_csamul_pg_rca24_fa3_14_out(.a(u_csamul_pg_rca24_and3_14[0]), .b(u_csamul_pg_rca24_fa4_13_xor1[0]), .cin(u_csamul_pg_rca24_fa3_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_14_xor1), .fa_or0(u_csamul_pg_rca24_fa3_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_14(.a(a[4]), .b(b[14]), .out(u_csamul_pg_rca24_and4_14));
  fa fa_u_csamul_pg_rca24_fa4_14_out(.a(u_csamul_pg_rca24_and4_14[0]), .b(u_csamul_pg_rca24_fa5_13_xor1[0]), .cin(u_csamul_pg_rca24_fa4_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_14_xor1), .fa_or0(u_csamul_pg_rca24_fa4_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_14(.a(a[5]), .b(b[14]), .out(u_csamul_pg_rca24_and5_14));
  fa fa_u_csamul_pg_rca24_fa5_14_out(.a(u_csamul_pg_rca24_and5_14[0]), .b(u_csamul_pg_rca24_fa6_13_xor1[0]), .cin(u_csamul_pg_rca24_fa5_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_14_xor1), .fa_or0(u_csamul_pg_rca24_fa5_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_14(.a(a[6]), .b(b[14]), .out(u_csamul_pg_rca24_and6_14));
  fa fa_u_csamul_pg_rca24_fa6_14_out(.a(u_csamul_pg_rca24_and6_14[0]), .b(u_csamul_pg_rca24_fa7_13_xor1[0]), .cin(u_csamul_pg_rca24_fa6_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_14_xor1), .fa_or0(u_csamul_pg_rca24_fa6_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_14(.a(a[7]), .b(b[14]), .out(u_csamul_pg_rca24_and7_14));
  fa fa_u_csamul_pg_rca24_fa7_14_out(.a(u_csamul_pg_rca24_and7_14[0]), .b(u_csamul_pg_rca24_fa8_13_xor1[0]), .cin(u_csamul_pg_rca24_fa7_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_14_xor1), .fa_or0(u_csamul_pg_rca24_fa7_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_14(.a(a[8]), .b(b[14]), .out(u_csamul_pg_rca24_and8_14));
  fa fa_u_csamul_pg_rca24_fa8_14_out(.a(u_csamul_pg_rca24_and8_14[0]), .b(u_csamul_pg_rca24_fa9_13_xor1[0]), .cin(u_csamul_pg_rca24_fa8_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_14_xor1), .fa_or0(u_csamul_pg_rca24_fa8_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_14(.a(a[9]), .b(b[14]), .out(u_csamul_pg_rca24_and9_14));
  fa fa_u_csamul_pg_rca24_fa9_14_out(.a(u_csamul_pg_rca24_and9_14[0]), .b(u_csamul_pg_rca24_fa10_13_xor1[0]), .cin(u_csamul_pg_rca24_fa9_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_14_xor1), .fa_or0(u_csamul_pg_rca24_fa9_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_14(.a(a[10]), .b(b[14]), .out(u_csamul_pg_rca24_and10_14));
  fa fa_u_csamul_pg_rca24_fa10_14_out(.a(u_csamul_pg_rca24_and10_14[0]), .b(u_csamul_pg_rca24_fa11_13_xor1[0]), .cin(u_csamul_pg_rca24_fa10_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_14_xor1), .fa_or0(u_csamul_pg_rca24_fa10_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_14(.a(a[11]), .b(b[14]), .out(u_csamul_pg_rca24_and11_14));
  fa fa_u_csamul_pg_rca24_fa11_14_out(.a(u_csamul_pg_rca24_and11_14[0]), .b(u_csamul_pg_rca24_fa12_13_xor1[0]), .cin(u_csamul_pg_rca24_fa11_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_14_xor1), .fa_or0(u_csamul_pg_rca24_fa11_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_14(.a(a[12]), .b(b[14]), .out(u_csamul_pg_rca24_and12_14));
  fa fa_u_csamul_pg_rca24_fa12_14_out(.a(u_csamul_pg_rca24_and12_14[0]), .b(u_csamul_pg_rca24_fa13_13_xor1[0]), .cin(u_csamul_pg_rca24_fa12_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_14_xor1), .fa_or0(u_csamul_pg_rca24_fa12_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_14(.a(a[13]), .b(b[14]), .out(u_csamul_pg_rca24_and13_14));
  fa fa_u_csamul_pg_rca24_fa13_14_out(.a(u_csamul_pg_rca24_and13_14[0]), .b(u_csamul_pg_rca24_fa14_13_xor1[0]), .cin(u_csamul_pg_rca24_fa13_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_14_xor1), .fa_or0(u_csamul_pg_rca24_fa13_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_14(.a(a[14]), .b(b[14]), .out(u_csamul_pg_rca24_and14_14));
  fa fa_u_csamul_pg_rca24_fa14_14_out(.a(u_csamul_pg_rca24_and14_14[0]), .b(u_csamul_pg_rca24_fa15_13_xor1[0]), .cin(u_csamul_pg_rca24_fa14_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_14_xor1), .fa_or0(u_csamul_pg_rca24_fa14_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_14(.a(a[15]), .b(b[14]), .out(u_csamul_pg_rca24_and15_14));
  fa fa_u_csamul_pg_rca24_fa15_14_out(.a(u_csamul_pg_rca24_and15_14[0]), .b(u_csamul_pg_rca24_fa16_13_xor1[0]), .cin(u_csamul_pg_rca24_fa15_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_14_xor1), .fa_or0(u_csamul_pg_rca24_fa15_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_14(.a(a[16]), .b(b[14]), .out(u_csamul_pg_rca24_and16_14));
  fa fa_u_csamul_pg_rca24_fa16_14_out(.a(u_csamul_pg_rca24_and16_14[0]), .b(u_csamul_pg_rca24_fa17_13_xor1[0]), .cin(u_csamul_pg_rca24_fa16_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_14_xor1), .fa_or0(u_csamul_pg_rca24_fa16_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_14(.a(a[17]), .b(b[14]), .out(u_csamul_pg_rca24_and17_14));
  fa fa_u_csamul_pg_rca24_fa17_14_out(.a(u_csamul_pg_rca24_and17_14[0]), .b(u_csamul_pg_rca24_fa18_13_xor1[0]), .cin(u_csamul_pg_rca24_fa17_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_14_xor1), .fa_or0(u_csamul_pg_rca24_fa17_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_14(.a(a[18]), .b(b[14]), .out(u_csamul_pg_rca24_and18_14));
  fa fa_u_csamul_pg_rca24_fa18_14_out(.a(u_csamul_pg_rca24_and18_14[0]), .b(u_csamul_pg_rca24_fa19_13_xor1[0]), .cin(u_csamul_pg_rca24_fa18_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_14_xor1), .fa_or0(u_csamul_pg_rca24_fa18_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_14(.a(a[19]), .b(b[14]), .out(u_csamul_pg_rca24_and19_14));
  fa fa_u_csamul_pg_rca24_fa19_14_out(.a(u_csamul_pg_rca24_and19_14[0]), .b(u_csamul_pg_rca24_fa20_13_xor1[0]), .cin(u_csamul_pg_rca24_fa19_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_14_xor1), .fa_or0(u_csamul_pg_rca24_fa19_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_14(.a(a[20]), .b(b[14]), .out(u_csamul_pg_rca24_and20_14));
  fa fa_u_csamul_pg_rca24_fa20_14_out(.a(u_csamul_pg_rca24_and20_14[0]), .b(u_csamul_pg_rca24_fa21_13_xor1[0]), .cin(u_csamul_pg_rca24_fa20_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_14_xor1), .fa_or0(u_csamul_pg_rca24_fa20_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_14(.a(a[21]), .b(b[14]), .out(u_csamul_pg_rca24_and21_14));
  fa fa_u_csamul_pg_rca24_fa21_14_out(.a(u_csamul_pg_rca24_and21_14[0]), .b(u_csamul_pg_rca24_fa22_13_xor1[0]), .cin(u_csamul_pg_rca24_fa21_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_14_xor1), .fa_or0(u_csamul_pg_rca24_fa21_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_14(.a(a[22]), .b(b[14]), .out(u_csamul_pg_rca24_and22_14));
  fa fa_u_csamul_pg_rca24_fa22_14_out(.a(u_csamul_pg_rca24_and22_14[0]), .b(u_csamul_pg_rca24_and23_13[0]), .cin(u_csamul_pg_rca24_fa22_13_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_14_xor1), .fa_or0(u_csamul_pg_rca24_fa22_14_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_14(.a(a[23]), .b(b[14]), .out(u_csamul_pg_rca24_and23_14));
  and_gate and_gate_u_csamul_pg_rca24_and0_15(.a(a[0]), .b(b[15]), .out(u_csamul_pg_rca24_and0_15));
  fa fa_u_csamul_pg_rca24_fa0_15_out(.a(u_csamul_pg_rca24_and0_15[0]), .b(u_csamul_pg_rca24_fa1_14_xor1[0]), .cin(u_csamul_pg_rca24_fa0_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_15_xor1), .fa_or0(u_csamul_pg_rca24_fa0_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_15(.a(a[1]), .b(b[15]), .out(u_csamul_pg_rca24_and1_15));
  fa fa_u_csamul_pg_rca24_fa1_15_out(.a(u_csamul_pg_rca24_and1_15[0]), .b(u_csamul_pg_rca24_fa2_14_xor1[0]), .cin(u_csamul_pg_rca24_fa1_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_15_xor1), .fa_or0(u_csamul_pg_rca24_fa1_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_15(.a(a[2]), .b(b[15]), .out(u_csamul_pg_rca24_and2_15));
  fa fa_u_csamul_pg_rca24_fa2_15_out(.a(u_csamul_pg_rca24_and2_15[0]), .b(u_csamul_pg_rca24_fa3_14_xor1[0]), .cin(u_csamul_pg_rca24_fa2_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_15_xor1), .fa_or0(u_csamul_pg_rca24_fa2_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_15(.a(a[3]), .b(b[15]), .out(u_csamul_pg_rca24_and3_15));
  fa fa_u_csamul_pg_rca24_fa3_15_out(.a(u_csamul_pg_rca24_and3_15[0]), .b(u_csamul_pg_rca24_fa4_14_xor1[0]), .cin(u_csamul_pg_rca24_fa3_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_15_xor1), .fa_or0(u_csamul_pg_rca24_fa3_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_15(.a(a[4]), .b(b[15]), .out(u_csamul_pg_rca24_and4_15));
  fa fa_u_csamul_pg_rca24_fa4_15_out(.a(u_csamul_pg_rca24_and4_15[0]), .b(u_csamul_pg_rca24_fa5_14_xor1[0]), .cin(u_csamul_pg_rca24_fa4_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_15_xor1), .fa_or0(u_csamul_pg_rca24_fa4_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_15(.a(a[5]), .b(b[15]), .out(u_csamul_pg_rca24_and5_15));
  fa fa_u_csamul_pg_rca24_fa5_15_out(.a(u_csamul_pg_rca24_and5_15[0]), .b(u_csamul_pg_rca24_fa6_14_xor1[0]), .cin(u_csamul_pg_rca24_fa5_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_15_xor1), .fa_or0(u_csamul_pg_rca24_fa5_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_15(.a(a[6]), .b(b[15]), .out(u_csamul_pg_rca24_and6_15));
  fa fa_u_csamul_pg_rca24_fa6_15_out(.a(u_csamul_pg_rca24_and6_15[0]), .b(u_csamul_pg_rca24_fa7_14_xor1[0]), .cin(u_csamul_pg_rca24_fa6_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_15_xor1), .fa_or0(u_csamul_pg_rca24_fa6_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_15(.a(a[7]), .b(b[15]), .out(u_csamul_pg_rca24_and7_15));
  fa fa_u_csamul_pg_rca24_fa7_15_out(.a(u_csamul_pg_rca24_and7_15[0]), .b(u_csamul_pg_rca24_fa8_14_xor1[0]), .cin(u_csamul_pg_rca24_fa7_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_15_xor1), .fa_or0(u_csamul_pg_rca24_fa7_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_15(.a(a[8]), .b(b[15]), .out(u_csamul_pg_rca24_and8_15));
  fa fa_u_csamul_pg_rca24_fa8_15_out(.a(u_csamul_pg_rca24_and8_15[0]), .b(u_csamul_pg_rca24_fa9_14_xor1[0]), .cin(u_csamul_pg_rca24_fa8_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_15_xor1), .fa_or0(u_csamul_pg_rca24_fa8_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_15(.a(a[9]), .b(b[15]), .out(u_csamul_pg_rca24_and9_15));
  fa fa_u_csamul_pg_rca24_fa9_15_out(.a(u_csamul_pg_rca24_and9_15[0]), .b(u_csamul_pg_rca24_fa10_14_xor1[0]), .cin(u_csamul_pg_rca24_fa9_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_15_xor1), .fa_or0(u_csamul_pg_rca24_fa9_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_15(.a(a[10]), .b(b[15]), .out(u_csamul_pg_rca24_and10_15));
  fa fa_u_csamul_pg_rca24_fa10_15_out(.a(u_csamul_pg_rca24_and10_15[0]), .b(u_csamul_pg_rca24_fa11_14_xor1[0]), .cin(u_csamul_pg_rca24_fa10_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_15_xor1), .fa_or0(u_csamul_pg_rca24_fa10_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_15(.a(a[11]), .b(b[15]), .out(u_csamul_pg_rca24_and11_15));
  fa fa_u_csamul_pg_rca24_fa11_15_out(.a(u_csamul_pg_rca24_and11_15[0]), .b(u_csamul_pg_rca24_fa12_14_xor1[0]), .cin(u_csamul_pg_rca24_fa11_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_15_xor1), .fa_or0(u_csamul_pg_rca24_fa11_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_15(.a(a[12]), .b(b[15]), .out(u_csamul_pg_rca24_and12_15));
  fa fa_u_csamul_pg_rca24_fa12_15_out(.a(u_csamul_pg_rca24_and12_15[0]), .b(u_csamul_pg_rca24_fa13_14_xor1[0]), .cin(u_csamul_pg_rca24_fa12_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_15_xor1), .fa_or0(u_csamul_pg_rca24_fa12_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_15(.a(a[13]), .b(b[15]), .out(u_csamul_pg_rca24_and13_15));
  fa fa_u_csamul_pg_rca24_fa13_15_out(.a(u_csamul_pg_rca24_and13_15[0]), .b(u_csamul_pg_rca24_fa14_14_xor1[0]), .cin(u_csamul_pg_rca24_fa13_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_15_xor1), .fa_or0(u_csamul_pg_rca24_fa13_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_15(.a(a[14]), .b(b[15]), .out(u_csamul_pg_rca24_and14_15));
  fa fa_u_csamul_pg_rca24_fa14_15_out(.a(u_csamul_pg_rca24_and14_15[0]), .b(u_csamul_pg_rca24_fa15_14_xor1[0]), .cin(u_csamul_pg_rca24_fa14_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_15_xor1), .fa_or0(u_csamul_pg_rca24_fa14_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_15(.a(a[15]), .b(b[15]), .out(u_csamul_pg_rca24_and15_15));
  fa fa_u_csamul_pg_rca24_fa15_15_out(.a(u_csamul_pg_rca24_and15_15[0]), .b(u_csamul_pg_rca24_fa16_14_xor1[0]), .cin(u_csamul_pg_rca24_fa15_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_15_xor1), .fa_or0(u_csamul_pg_rca24_fa15_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_15(.a(a[16]), .b(b[15]), .out(u_csamul_pg_rca24_and16_15));
  fa fa_u_csamul_pg_rca24_fa16_15_out(.a(u_csamul_pg_rca24_and16_15[0]), .b(u_csamul_pg_rca24_fa17_14_xor1[0]), .cin(u_csamul_pg_rca24_fa16_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_15_xor1), .fa_or0(u_csamul_pg_rca24_fa16_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_15(.a(a[17]), .b(b[15]), .out(u_csamul_pg_rca24_and17_15));
  fa fa_u_csamul_pg_rca24_fa17_15_out(.a(u_csamul_pg_rca24_and17_15[0]), .b(u_csamul_pg_rca24_fa18_14_xor1[0]), .cin(u_csamul_pg_rca24_fa17_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_15_xor1), .fa_or0(u_csamul_pg_rca24_fa17_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_15(.a(a[18]), .b(b[15]), .out(u_csamul_pg_rca24_and18_15));
  fa fa_u_csamul_pg_rca24_fa18_15_out(.a(u_csamul_pg_rca24_and18_15[0]), .b(u_csamul_pg_rca24_fa19_14_xor1[0]), .cin(u_csamul_pg_rca24_fa18_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_15_xor1), .fa_or0(u_csamul_pg_rca24_fa18_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_15(.a(a[19]), .b(b[15]), .out(u_csamul_pg_rca24_and19_15));
  fa fa_u_csamul_pg_rca24_fa19_15_out(.a(u_csamul_pg_rca24_and19_15[0]), .b(u_csamul_pg_rca24_fa20_14_xor1[0]), .cin(u_csamul_pg_rca24_fa19_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_15_xor1), .fa_or0(u_csamul_pg_rca24_fa19_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_15(.a(a[20]), .b(b[15]), .out(u_csamul_pg_rca24_and20_15));
  fa fa_u_csamul_pg_rca24_fa20_15_out(.a(u_csamul_pg_rca24_and20_15[0]), .b(u_csamul_pg_rca24_fa21_14_xor1[0]), .cin(u_csamul_pg_rca24_fa20_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_15_xor1), .fa_or0(u_csamul_pg_rca24_fa20_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_15(.a(a[21]), .b(b[15]), .out(u_csamul_pg_rca24_and21_15));
  fa fa_u_csamul_pg_rca24_fa21_15_out(.a(u_csamul_pg_rca24_and21_15[0]), .b(u_csamul_pg_rca24_fa22_14_xor1[0]), .cin(u_csamul_pg_rca24_fa21_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_15_xor1), .fa_or0(u_csamul_pg_rca24_fa21_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_15(.a(a[22]), .b(b[15]), .out(u_csamul_pg_rca24_and22_15));
  fa fa_u_csamul_pg_rca24_fa22_15_out(.a(u_csamul_pg_rca24_and22_15[0]), .b(u_csamul_pg_rca24_and23_14[0]), .cin(u_csamul_pg_rca24_fa22_14_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_15_xor1), .fa_or0(u_csamul_pg_rca24_fa22_15_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_15(.a(a[23]), .b(b[15]), .out(u_csamul_pg_rca24_and23_15));
  and_gate and_gate_u_csamul_pg_rca24_and0_16(.a(a[0]), .b(b[16]), .out(u_csamul_pg_rca24_and0_16));
  fa fa_u_csamul_pg_rca24_fa0_16_out(.a(u_csamul_pg_rca24_and0_16[0]), .b(u_csamul_pg_rca24_fa1_15_xor1[0]), .cin(u_csamul_pg_rca24_fa0_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_16_xor1), .fa_or0(u_csamul_pg_rca24_fa0_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_16(.a(a[1]), .b(b[16]), .out(u_csamul_pg_rca24_and1_16));
  fa fa_u_csamul_pg_rca24_fa1_16_out(.a(u_csamul_pg_rca24_and1_16[0]), .b(u_csamul_pg_rca24_fa2_15_xor1[0]), .cin(u_csamul_pg_rca24_fa1_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_16_xor1), .fa_or0(u_csamul_pg_rca24_fa1_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_16(.a(a[2]), .b(b[16]), .out(u_csamul_pg_rca24_and2_16));
  fa fa_u_csamul_pg_rca24_fa2_16_out(.a(u_csamul_pg_rca24_and2_16[0]), .b(u_csamul_pg_rca24_fa3_15_xor1[0]), .cin(u_csamul_pg_rca24_fa2_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_16_xor1), .fa_or0(u_csamul_pg_rca24_fa2_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_16(.a(a[3]), .b(b[16]), .out(u_csamul_pg_rca24_and3_16));
  fa fa_u_csamul_pg_rca24_fa3_16_out(.a(u_csamul_pg_rca24_and3_16[0]), .b(u_csamul_pg_rca24_fa4_15_xor1[0]), .cin(u_csamul_pg_rca24_fa3_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_16_xor1), .fa_or0(u_csamul_pg_rca24_fa3_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_16(.a(a[4]), .b(b[16]), .out(u_csamul_pg_rca24_and4_16));
  fa fa_u_csamul_pg_rca24_fa4_16_out(.a(u_csamul_pg_rca24_and4_16[0]), .b(u_csamul_pg_rca24_fa5_15_xor1[0]), .cin(u_csamul_pg_rca24_fa4_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_16_xor1), .fa_or0(u_csamul_pg_rca24_fa4_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_16(.a(a[5]), .b(b[16]), .out(u_csamul_pg_rca24_and5_16));
  fa fa_u_csamul_pg_rca24_fa5_16_out(.a(u_csamul_pg_rca24_and5_16[0]), .b(u_csamul_pg_rca24_fa6_15_xor1[0]), .cin(u_csamul_pg_rca24_fa5_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_16_xor1), .fa_or0(u_csamul_pg_rca24_fa5_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_16(.a(a[6]), .b(b[16]), .out(u_csamul_pg_rca24_and6_16));
  fa fa_u_csamul_pg_rca24_fa6_16_out(.a(u_csamul_pg_rca24_and6_16[0]), .b(u_csamul_pg_rca24_fa7_15_xor1[0]), .cin(u_csamul_pg_rca24_fa6_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_16_xor1), .fa_or0(u_csamul_pg_rca24_fa6_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_16(.a(a[7]), .b(b[16]), .out(u_csamul_pg_rca24_and7_16));
  fa fa_u_csamul_pg_rca24_fa7_16_out(.a(u_csamul_pg_rca24_and7_16[0]), .b(u_csamul_pg_rca24_fa8_15_xor1[0]), .cin(u_csamul_pg_rca24_fa7_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_16_xor1), .fa_or0(u_csamul_pg_rca24_fa7_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_16(.a(a[8]), .b(b[16]), .out(u_csamul_pg_rca24_and8_16));
  fa fa_u_csamul_pg_rca24_fa8_16_out(.a(u_csamul_pg_rca24_and8_16[0]), .b(u_csamul_pg_rca24_fa9_15_xor1[0]), .cin(u_csamul_pg_rca24_fa8_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_16_xor1), .fa_or0(u_csamul_pg_rca24_fa8_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_16(.a(a[9]), .b(b[16]), .out(u_csamul_pg_rca24_and9_16));
  fa fa_u_csamul_pg_rca24_fa9_16_out(.a(u_csamul_pg_rca24_and9_16[0]), .b(u_csamul_pg_rca24_fa10_15_xor1[0]), .cin(u_csamul_pg_rca24_fa9_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_16_xor1), .fa_or0(u_csamul_pg_rca24_fa9_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_16(.a(a[10]), .b(b[16]), .out(u_csamul_pg_rca24_and10_16));
  fa fa_u_csamul_pg_rca24_fa10_16_out(.a(u_csamul_pg_rca24_and10_16[0]), .b(u_csamul_pg_rca24_fa11_15_xor1[0]), .cin(u_csamul_pg_rca24_fa10_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_16_xor1), .fa_or0(u_csamul_pg_rca24_fa10_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_16(.a(a[11]), .b(b[16]), .out(u_csamul_pg_rca24_and11_16));
  fa fa_u_csamul_pg_rca24_fa11_16_out(.a(u_csamul_pg_rca24_and11_16[0]), .b(u_csamul_pg_rca24_fa12_15_xor1[0]), .cin(u_csamul_pg_rca24_fa11_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_16_xor1), .fa_or0(u_csamul_pg_rca24_fa11_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_16(.a(a[12]), .b(b[16]), .out(u_csamul_pg_rca24_and12_16));
  fa fa_u_csamul_pg_rca24_fa12_16_out(.a(u_csamul_pg_rca24_and12_16[0]), .b(u_csamul_pg_rca24_fa13_15_xor1[0]), .cin(u_csamul_pg_rca24_fa12_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_16_xor1), .fa_or0(u_csamul_pg_rca24_fa12_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_16(.a(a[13]), .b(b[16]), .out(u_csamul_pg_rca24_and13_16));
  fa fa_u_csamul_pg_rca24_fa13_16_out(.a(u_csamul_pg_rca24_and13_16[0]), .b(u_csamul_pg_rca24_fa14_15_xor1[0]), .cin(u_csamul_pg_rca24_fa13_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_16_xor1), .fa_or0(u_csamul_pg_rca24_fa13_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_16(.a(a[14]), .b(b[16]), .out(u_csamul_pg_rca24_and14_16));
  fa fa_u_csamul_pg_rca24_fa14_16_out(.a(u_csamul_pg_rca24_and14_16[0]), .b(u_csamul_pg_rca24_fa15_15_xor1[0]), .cin(u_csamul_pg_rca24_fa14_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_16_xor1), .fa_or0(u_csamul_pg_rca24_fa14_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_16(.a(a[15]), .b(b[16]), .out(u_csamul_pg_rca24_and15_16));
  fa fa_u_csamul_pg_rca24_fa15_16_out(.a(u_csamul_pg_rca24_and15_16[0]), .b(u_csamul_pg_rca24_fa16_15_xor1[0]), .cin(u_csamul_pg_rca24_fa15_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_16_xor1), .fa_or0(u_csamul_pg_rca24_fa15_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_16(.a(a[16]), .b(b[16]), .out(u_csamul_pg_rca24_and16_16));
  fa fa_u_csamul_pg_rca24_fa16_16_out(.a(u_csamul_pg_rca24_and16_16[0]), .b(u_csamul_pg_rca24_fa17_15_xor1[0]), .cin(u_csamul_pg_rca24_fa16_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_16_xor1), .fa_or0(u_csamul_pg_rca24_fa16_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_16(.a(a[17]), .b(b[16]), .out(u_csamul_pg_rca24_and17_16));
  fa fa_u_csamul_pg_rca24_fa17_16_out(.a(u_csamul_pg_rca24_and17_16[0]), .b(u_csamul_pg_rca24_fa18_15_xor1[0]), .cin(u_csamul_pg_rca24_fa17_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_16_xor1), .fa_or0(u_csamul_pg_rca24_fa17_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_16(.a(a[18]), .b(b[16]), .out(u_csamul_pg_rca24_and18_16));
  fa fa_u_csamul_pg_rca24_fa18_16_out(.a(u_csamul_pg_rca24_and18_16[0]), .b(u_csamul_pg_rca24_fa19_15_xor1[0]), .cin(u_csamul_pg_rca24_fa18_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_16_xor1), .fa_or0(u_csamul_pg_rca24_fa18_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_16(.a(a[19]), .b(b[16]), .out(u_csamul_pg_rca24_and19_16));
  fa fa_u_csamul_pg_rca24_fa19_16_out(.a(u_csamul_pg_rca24_and19_16[0]), .b(u_csamul_pg_rca24_fa20_15_xor1[0]), .cin(u_csamul_pg_rca24_fa19_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_16_xor1), .fa_or0(u_csamul_pg_rca24_fa19_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_16(.a(a[20]), .b(b[16]), .out(u_csamul_pg_rca24_and20_16));
  fa fa_u_csamul_pg_rca24_fa20_16_out(.a(u_csamul_pg_rca24_and20_16[0]), .b(u_csamul_pg_rca24_fa21_15_xor1[0]), .cin(u_csamul_pg_rca24_fa20_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_16_xor1), .fa_or0(u_csamul_pg_rca24_fa20_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_16(.a(a[21]), .b(b[16]), .out(u_csamul_pg_rca24_and21_16));
  fa fa_u_csamul_pg_rca24_fa21_16_out(.a(u_csamul_pg_rca24_and21_16[0]), .b(u_csamul_pg_rca24_fa22_15_xor1[0]), .cin(u_csamul_pg_rca24_fa21_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_16_xor1), .fa_or0(u_csamul_pg_rca24_fa21_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_16(.a(a[22]), .b(b[16]), .out(u_csamul_pg_rca24_and22_16));
  fa fa_u_csamul_pg_rca24_fa22_16_out(.a(u_csamul_pg_rca24_and22_16[0]), .b(u_csamul_pg_rca24_and23_15[0]), .cin(u_csamul_pg_rca24_fa22_15_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_16_xor1), .fa_or0(u_csamul_pg_rca24_fa22_16_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_16(.a(a[23]), .b(b[16]), .out(u_csamul_pg_rca24_and23_16));
  and_gate and_gate_u_csamul_pg_rca24_and0_17(.a(a[0]), .b(b[17]), .out(u_csamul_pg_rca24_and0_17));
  fa fa_u_csamul_pg_rca24_fa0_17_out(.a(u_csamul_pg_rca24_and0_17[0]), .b(u_csamul_pg_rca24_fa1_16_xor1[0]), .cin(u_csamul_pg_rca24_fa0_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_17_xor1), .fa_or0(u_csamul_pg_rca24_fa0_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_17(.a(a[1]), .b(b[17]), .out(u_csamul_pg_rca24_and1_17));
  fa fa_u_csamul_pg_rca24_fa1_17_out(.a(u_csamul_pg_rca24_and1_17[0]), .b(u_csamul_pg_rca24_fa2_16_xor1[0]), .cin(u_csamul_pg_rca24_fa1_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_17_xor1), .fa_or0(u_csamul_pg_rca24_fa1_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_17(.a(a[2]), .b(b[17]), .out(u_csamul_pg_rca24_and2_17));
  fa fa_u_csamul_pg_rca24_fa2_17_out(.a(u_csamul_pg_rca24_and2_17[0]), .b(u_csamul_pg_rca24_fa3_16_xor1[0]), .cin(u_csamul_pg_rca24_fa2_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_17_xor1), .fa_or0(u_csamul_pg_rca24_fa2_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_17(.a(a[3]), .b(b[17]), .out(u_csamul_pg_rca24_and3_17));
  fa fa_u_csamul_pg_rca24_fa3_17_out(.a(u_csamul_pg_rca24_and3_17[0]), .b(u_csamul_pg_rca24_fa4_16_xor1[0]), .cin(u_csamul_pg_rca24_fa3_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_17_xor1), .fa_or0(u_csamul_pg_rca24_fa3_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_17(.a(a[4]), .b(b[17]), .out(u_csamul_pg_rca24_and4_17));
  fa fa_u_csamul_pg_rca24_fa4_17_out(.a(u_csamul_pg_rca24_and4_17[0]), .b(u_csamul_pg_rca24_fa5_16_xor1[0]), .cin(u_csamul_pg_rca24_fa4_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_17_xor1), .fa_or0(u_csamul_pg_rca24_fa4_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_17(.a(a[5]), .b(b[17]), .out(u_csamul_pg_rca24_and5_17));
  fa fa_u_csamul_pg_rca24_fa5_17_out(.a(u_csamul_pg_rca24_and5_17[0]), .b(u_csamul_pg_rca24_fa6_16_xor1[0]), .cin(u_csamul_pg_rca24_fa5_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_17_xor1), .fa_or0(u_csamul_pg_rca24_fa5_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_17(.a(a[6]), .b(b[17]), .out(u_csamul_pg_rca24_and6_17));
  fa fa_u_csamul_pg_rca24_fa6_17_out(.a(u_csamul_pg_rca24_and6_17[0]), .b(u_csamul_pg_rca24_fa7_16_xor1[0]), .cin(u_csamul_pg_rca24_fa6_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_17_xor1), .fa_or0(u_csamul_pg_rca24_fa6_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_17(.a(a[7]), .b(b[17]), .out(u_csamul_pg_rca24_and7_17));
  fa fa_u_csamul_pg_rca24_fa7_17_out(.a(u_csamul_pg_rca24_and7_17[0]), .b(u_csamul_pg_rca24_fa8_16_xor1[0]), .cin(u_csamul_pg_rca24_fa7_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_17_xor1), .fa_or0(u_csamul_pg_rca24_fa7_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_17(.a(a[8]), .b(b[17]), .out(u_csamul_pg_rca24_and8_17));
  fa fa_u_csamul_pg_rca24_fa8_17_out(.a(u_csamul_pg_rca24_and8_17[0]), .b(u_csamul_pg_rca24_fa9_16_xor1[0]), .cin(u_csamul_pg_rca24_fa8_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_17_xor1), .fa_or0(u_csamul_pg_rca24_fa8_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_17(.a(a[9]), .b(b[17]), .out(u_csamul_pg_rca24_and9_17));
  fa fa_u_csamul_pg_rca24_fa9_17_out(.a(u_csamul_pg_rca24_and9_17[0]), .b(u_csamul_pg_rca24_fa10_16_xor1[0]), .cin(u_csamul_pg_rca24_fa9_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_17_xor1), .fa_or0(u_csamul_pg_rca24_fa9_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_17(.a(a[10]), .b(b[17]), .out(u_csamul_pg_rca24_and10_17));
  fa fa_u_csamul_pg_rca24_fa10_17_out(.a(u_csamul_pg_rca24_and10_17[0]), .b(u_csamul_pg_rca24_fa11_16_xor1[0]), .cin(u_csamul_pg_rca24_fa10_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_17_xor1), .fa_or0(u_csamul_pg_rca24_fa10_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_17(.a(a[11]), .b(b[17]), .out(u_csamul_pg_rca24_and11_17));
  fa fa_u_csamul_pg_rca24_fa11_17_out(.a(u_csamul_pg_rca24_and11_17[0]), .b(u_csamul_pg_rca24_fa12_16_xor1[0]), .cin(u_csamul_pg_rca24_fa11_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_17_xor1), .fa_or0(u_csamul_pg_rca24_fa11_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_17(.a(a[12]), .b(b[17]), .out(u_csamul_pg_rca24_and12_17));
  fa fa_u_csamul_pg_rca24_fa12_17_out(.a(u_csamul_pg_rca24_and12_17[0]), .b(u_csamul_pg_rca24_fa13_16_xor1[0]), .cin(u_csamul_pg_rca24_fa12_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_17_xor1), .fa_or0(u_csamul_pg_rca24_fa12_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_17(.a(a[13]), .b(b[17]), .out(u_csamul_pg_rca24_and13_17));
  fa fa_u_csamul_pg_rca24_fa13_17_out(.a(u_csamul_pg_rca24_and13_17[0]), .b(u_csamul_pg_rca24_fa14_16_xor1[0]), .cin(u_csamul_pg_rca24_fa13_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_17_xor1), .fa_or0(u_csamul_pg_rca24_fa13_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_17(.a(a[14]), .b(b[17]), .out(u_csamul_pg_rca24_and14_17));
  fa fa_u_csamul_pg_rca24_fa14_17_out(.a(u_csamul_pg_rca24_and14_17[0]), .b(u_csamul_pg_rca24_fa15_16_xor1[0]), .cin(u_csamul_pg_rca24_fa14_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_17_xor1), .fa_or0(u_csamul_pg_rca24_fa14_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_17(.a(a[15]), .b(b[17]), .out(u_csamul_pg_rca24_and15_17));
  fa fa_u_csamul_pg_rca24_fa15_17_out(.a(u_csamul_pg_rca24_and15_17[0]), .b(u_csamul_pg_rca24_fa16_16_xor1[0]), .cin(u_csamul_pg_rca24_fa15_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_17_xor1), .fa_or0(u_csamul_pg_rca24_fa15_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_17(.a(a[16]), .b(b[17]), .out(u_csamul_pg_rca24_and16_17));
  fa fa_u_csamul_pg_rca24_fa16_17_out(.a(u_csamul_pg_rca24_and16_17[0]), .b(u_csamul_pg_rca24_fa17_16_xor1[0]), .cin(u_csamul_pg_rca24_fa16_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_17_xor1), .fa_or0(u_csamul_pg_rca24_fa16_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_17(.a(a[17]), .b(b[17]), .out(u_csamul_pg_rca24_and17_17));
  fa fa_u_csamul_pg_rca24_fa17_17_out(.a(u_csamul_pg_rca24_and17_17[0]), .b(u_csamul_pg_rca24_fa18_16_xor1[0]), .cin(u_csamul_pg_rca24_fa17_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_17_xor1), .fa_or0(u_csamul_pg_rca24_fa17_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_17(.a(a[18]), .b(b[17]), .out(u_csamul_pg_rca24_and18_17));
  fa fa_u_csamul_pg_rca24_fa18_17_out(.a(u_csamul_pg_rca24_and18_17[0]), .b(u_csamul_pg_rca24_fa19_16_xor1[0]), .cin(u_csamul_pg_rca24_fa18_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_17_xor1), .fa_or0(u_csamul_pg_rca24_fa18_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_17(.a(a[19]), .b(b[17]), .out(u_csamul_pg_rca24_and19_17));
  fa fa_u_csamul_pg_rca24_fa19_17_out(.a(u_csamul_pg_rca24_and19_17[0]), .b(u_csamul_pg_rca24_fa20_16_xor1[0]), .cin(u_csamul_pg_rca24_fa19_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_17_xor1), .fa_or0(u_csamul_pg_rca24_fa19_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_17(.a(a[20]), .b(b[17]), .out(u_csamul_pg_rca24_and20_17));
  fa fa_u_csamul_pg_rca24_fa20_17_out(.a(u_csamul_pg_rca24_and20_17[0]), .b(u_csamul_pg_rca24_fa21_16_xor1[0]), .cin(u_csamul_pg_rca24_fa20_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_17_xor1), .fa_or0(u_csamul_pg_rca24_fa20_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_17(.a(a[21]), .b(b[17]), .out(u_csamul_pg_rca24_and21_17));
  fa fa_u_csamul_pg_rca24_fa21_17_out(.a(u_csamul_pg_rca24_and21_17[0]), .b(u_csamul_pg_rca24_fa22_16_xor1[0]), .cin(u_csamul_pg_rca24_fa21_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_17_xor1), .fa_or0(u_csamul_pg_rca24_fa21_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_17(.a(a[22]), .b(b[17]), .out(u_csamul_pg_rca24_and22_17));
  fa fa_u_csamul_pg_rca24_fa22_17_out(.a(u_csamul_pg_rca24_and22_17[0]), .b(u_csamul_pg_rca24_and23_16[0]), .cin(u_csamul_pg_rca24_fa22_16_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_17_xor1), .fa_or0(u_csamul_pg_rca24_fa22_17_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_17(.a(a[23]), .b(b[17]), .out(u_csamul_pg_rca24_and23_17));
  and_gate and_gate_u_csamul_pg_rca24_and0_18(.a(a[0]), .b(b[18]), .out(u_csamul_pg_rca24_and0_18));
  fa fa_u_csamul_pg_rca24_fa0_18_out(.a(u_csamul_pg_rca24_and0_18[0]), .b(u_csamul_pg_rca24_fa1_17_xor1[0]), .cin(u_csamul_pg_rca24_fa0_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_18_xor1), .fa_or0(u_csamul_pg_rca24_fa0_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_18(.a(a[1]), .b(b[18]), .out(u_csamul_pg_rca24_and1_18));
  fa fa_u_csamul_pg_rca24_fa1_18_out(.a(u_csamul_pg_rca24_and1_18[0]), .b(u_csamul_pg_rca24_fa2_17_xor1[0]), .cin(u_csamul_pg_rca24_fa1_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_18_xor1), .fa_or0(u_csamul_pg_rca24_fa1_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_18(.a(a[2]), .b(b[18]), .out(u_csamul_pg_rca24_and2_18));
  fa fa_u_csamul_pg_rca24_fa2_18_out(.a(u_csamul_pg_rca24_and2_18[0]), .b(u_csamul_pg_rca24_fa3_17_xor1[0]), .cin(u_csamul_pg_rca24_fa2_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_18_xor1), .fa_or0(u_csamul_pg_rca24_fa2_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_18(.a(a[3]), .b(b[18]), .out(u_csamul_pg_rca24_and3_18));
  fa fa_u_csamul_pg_rca24_fa3_18_out(.a(u_csamul_pg_rca24_and3_18[0]), .b(u_csamul_pg_rca24_fa4_17_xor1[0]), .cin(u_csamul_pg_rca24_fa3_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_18_xor1), .fa_or0(u_csamul_pg_rca24_fa3_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_18(.a(a[4]), .b(b[18]), .out(u_csamul_pg_rca24_and4_18));
  fa fa_u_csamul_pg_rca24_fa4_18_out(.a(u_csamul_pg_rca24_and4_18[0]), .b(u_csamul_pg_rca24_fa5_17_xor1[0]), .cin(u_csamul_pg_rca24_fa4_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_18_xor1), .fa_or0(u_csamul_pg_rca24_fa4_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_18(.a(a[5]), .b(b[18]), .out(u_csamul_pg_rca24_and5_18));
  fa fa_u_csamul_pg_rca24_fa5_18_out(.a(u_csamul_pg_rca24_and5_18[0]), .b(u_csamul_pg_rca24_fa6_17_xor1[0]), .cin(u_csamul_pg_rca24_fa5_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_18_xor1), .fa_or0(u_csamul_pg_rca24_fa5_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_18(.a(a[6]), .b(b[18]), .out(u_csamul_pg_rca24_and6_18));
  fa fa_u_csamul_pg_rca24_fa6_18_out(.a(u_csamul_pg_rca24_and6_18[0]), .b(u_csamul_pg_rca24_fa7_17_xor1[0]), .cin(u_csamul_pg_rca24_fa6_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_18_xor1), .fa_or0(u_csamul_pg_rca24_fa6_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_18(.a(a[7]), .b(b[18]), .out(u_csamul_pg_rca24_and7_18));
  fa fa_u_csamul_pg_rca24_fa7_18_out(.a(u_csamul_pg_rca24_and7_18[0]), .b(u_csamul_pg_rca24_fa8_17_xor1[0]), .cin(u_csamul_pg_rca24_fa7_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_18_xor1), .fa_or0(u_csamul_pg_rca24_fa7_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_18(.a(a[8]), .b(b[18]), .out(u_csamul_pg_rca24_and8_18));
  fa fa_u_csamul_pg_rca24_fa8_18_out(.a(u_csamul_pg_rca24_and8_18[0]), .b(u_csamul_pg_rca24_fa9_17_xor1[0]), .cin(u_csamul_pg_rca24_fa8_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_18_xor1), .fa_or0(u_csamul_pg_rca24_fa8_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_18(.a(a[9]), .b(b[18]), .out(u_csamul_pg_rca24_and9_18));
  fa fa_u_csamul_pg_rca24_fa9_18_out(.a(u_csamul_pg_rca24_and9_18[0]), .b(u_csamul_pg_rca24_fa10_17_xor1[0]), .cin(u_csamul_pg_rca24_fa9_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_18_xor1), .fa_or0(u_csamul_pg_rca24_fa9_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_18(.a(a[10]), .b(b[18]), .out(u_csamul_pg_rca24_and10_18));
  fa fa_u_csamul_pg_rca24_fa10_18_out(.a(u_csamul_pg_rca24_and10_18[0]), .b(u_csamul_pg_rca24_fa11_17_xor1[0]), .cin(u_csamul_pg_rca24_fa10_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_18_xor1), .fa_or0(u_csamul_pg_rca24_fa10_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_18(.a(a[11]), .b(b[18]), .out(u_csamul_pg_rca24_and11_18));
  fa fa_u_csamul_pg_rca24_fa11_18_out(.a(u_csamul_pg_rca24_and11_18[0]), .b(u_csamul_pg_rca24_fa12_17_xor1[0]), .cin(u_csamul_pg_rca24_fa11_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_18_xor1), .fa_or0(u_csamul_pg_rca24_fa11_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_18(.a(a[12]), .b(b[18]), .out(u_csamul_pg_rca24_and12_18));
  fa fa_u_csamul_pg_rca24_fa12_18_out(.a(u_csamul_pg_rca24_and12_18[0]), .b(u_csamul_pg_rca24_fa13_17_xor1[0]), .cin(u_csamul_pg_rca24_fa12_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_18_xor1), .fa_or0(u_csamul_pg_rca24_fa12_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_18(.a(a[13]), .b(b[18]), .out(u_csamul_pg_rca24_and13_18));
  fa fa_u_csamul_pg_rca24_fa13_18_out(.a(u_csamul_pg_rca24_and13_18[0]), .b(u_csamul_pg_rca24_fa14_17_xor1[0]), .cin(u_csamul_pg_rca24_fa13_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_18_xor1), .fa_or0(u_csamul_pg_rca24_fa13_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_18(.a(a[14]), .b(b[18]), .out(u_csamul_pg_rca24_and14_18));
  fa fa_u_csamul_pg_rca24_fa14_18_out(.a(u_csamul_pg_rca24_and14_18[0]), .b(u_csamul_pg_rca24_fa15_17_xor1[0]), .cin(u_csamul_pg_rca24_fa14_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_18_xor1), .fa_or0(u_csamul_pg_rca24_fa14_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_18(.a(a[15]), .b(b[18]), .out(u_csamul_pg_rca24_and15_18));
  fa fa_u_csamul_pg_rca24_fa15_18_out(.a(u_csamul_pg_rca24_and15_18[0]), .b(u_csamul_pg_rca24_fa16_17_xor1[0]), .cin(u_csamul_pg_rca24_fa15_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_18_xor1), .fa_or0(u_csamul_pg_rca24_fa15_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_18(.a(a[16]), .b(b[18]), .out(u_csamul_pg_rca24_and16_18));
  fa fa_u_csamul_pg_rca24_fa16_18_out(.a(u_csamul_pg_rca24_and16_18[0]), .b(u_csamul_pg_rca24_fa17_17_xor1[0]), .cin(u_csamul_pg_rca24_fa16_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_18_xor1), .fa_or0(u_csamul_pg_rca24_fa16_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_18(.a(a[17]), .b(b[18]), .out(u_csamul_pg_rca24_and17_18));
  fa fa_u_csamul_pg_rca24_fa17_18_out(.a(u_csamul_pg_rca24_and17_18[0]), .b(u_csamul_pg_rca24_fa18_17_xor1[0]), .cin(u_csamul_pg_rca24_fa17_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_18_xor1), .fa_or0(u_csamul_pg_rca24_fa17_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_18(.a(a[18]), .b(b[18]), .out(u_csamul_pg_rca24_and18_18));
  fa fa_u_csamul_pg_rca24_fa18_18_out(.a(u_csamul_pg_rca24_and18_18[0]), .b(u_csamul_pg_rca24_fa19_17_xor1[0]), .cin(u_csamul_pg_rca24_fa18_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_18_xor1), .fa_or0(u_csamul_pg_rca24_fa18_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_18(.a(a[19]), .b(b[18]), .out(u_csamul_pg_rca24_and19_18));
  fa fa_u_csamul_pg_rca24_fa19_18_out(.a(u_csamul_pg_rca24_and19_18[0]), .b(u_csamul_pg_rca24_fa20_17_xor1[0]), .cin(u_csamul_pg_rca24_fa19_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_18_xor1), .fa_or0(u_csamul_pg_rca24_fa19_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_18(.a(a[20]), .b(b[18]), .out(u_csamul_pg_rca24_and20_18));
  fa fa_u_csamul_pg_rca24_fa20_18_out(.a(u_csamul_pg_rca24_and20_18[0]), .b(u_csamul_pg_rca24_fa21_17_xor1[0]), .cin(u_csamul_pg_rca24_fa20_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_18_xor1), .fa_or0(u_csamul_pg_rca24_fa20_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_18(.a(a[21]), .b(b[18]), .out(u_csamul_pg_rca24_and21_18));
  fa fa_u_csamul_pg_rca24_fa21_18_out(.a(u_csamul_pg_rca24_and21_18[0]), .b(u_csamul_pg_rca24_fa22_17_xor1[0]), .cin(u_csamul_pg_rca24_fa21_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_18_xor1), .fa_or0(u_csamul_pg_rca24_fa21_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_18(.a(a[22]), .b(b[18]), .out(u_csamul_pg_rca24_and22_18));
  fa fa_u_csamul_pg_rca24_fa22_18_out(.a(u_csamul_pg_rca24_and22_18[0]), .b(u_csamul_pg_rca24_and23_17[0]), .cin(u_csamul_pg_rca24_fa22_17_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_18_xor1), .fa_or0(u_csamul_pg_rca24_fa22_18_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_18(.a(a[23]), .b(b[18]), .out(u_csamul_pg_rca24_and23_18));
  and_gate and_gate_u_csamul_pg_rca24_and0_19(.a(a[0]), .b(b[19]), .out(u_csamul_pg_rca24_and0_19));
  fa fa_u_csamul_pg_rca24_fa0_19_out(.a(u_csamul_pg_rca24_and0_19[0]), .b(u_csamul_pg_rca24_fa1_18_xor1[0]), .cin(u_csamul_pg_rca24_fa0_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_19_xor1), .fa_or0(u_csamul_pg_rca24_fa0_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_19(.a(a[1]), .b(b[19]), .out(u_csamul_pg_rca24_and1_19));
  fa fa_u_csamul_pg_rca24_fa1_19_out(.a(u_csamul_pg_rca24_and1_19[0]), .b(u_csamul_pg_rca24_fa2_18_xor1[0]), .cin(u_csamul_pg_rca24_fa1_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_19_xor1), .fa_or0(u_csamul_pg_rca24_fa1_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_19(.a(a[2]), .b(b[19]), .out(u_csamul_pg_rca24_and2_19));
  fa fa_u_csamul_pg_rca24_fa2_19_out(.a(u_csamul_pg_rca24_and2_19[0]), .b(u_csamul_pg_rca24_fa3_18_xor1[0]), .cin(u_csamul_pg_rca24_fa2_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_19_xor1), .fa_or0(u_csamul_pg_rca24_fa2_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_19(.a(a[3]), .b(b[19]), .out(u_csamul_pg_rca24_and3_19));
  fa fa_u_csamul_pg_rca24_fa3_19_out(.a(u_csamul_pg_rca24_and3_19[0]), .b(u_csamul_pg_rca24_fa4_18_xor1[0]), .cin(u_csamul_pg_rca24_fa3_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_19_xor1), .fa_or0(u_csamul_pg_rca24_fa3_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_19(.a(a[4]), .b(b[19]), .out(u_csamul_pg_rca24_and4_19));
  fa fa_u_csamul_pg_rca24_fa4_19_out(.a(u_csamul_pg_rca24_and4_19[0]), .b(u_csamul_pg_rca24_fa5_18_xor1[0]), .cin(u_csamul_pg_rca24_fa4_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_19_xor1), .fa_or0(u_csamul_pg_rca24_fa4_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_19(.a(a[5]), .b(b[19]), .out(u_csamul_pg_rca24_and5_19));
  fa fa_u_csamul_pg_rca24_fa5_19_out(.a(u_csamul_pg_rca24_and5_19[0]), .b(u_csamul_pg_rca24_fa6_18_xor1[0]), .cin(u_csamul_pg_rca24_fa5_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_19_xor1), .fa_or0(u_csamul_pg_rca24_fa5_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_19(.a(a[6]), .b(b[19]), .out(u_csamul_pg_rca24_and6_19));
  fa fa_u_csamul_pg_rca24_fa6_19_out(.a(u_csamul_pg_rca24_and6_19[0]), .b(u_csamul_pg_rca24_fa7_18_xor1[0]), .cin(u_csamul_pg_rca24_fa6_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_19_xor1), .fa_or0(u_csamul_pg_rca24_fa6_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_19(.a(a[7]), .b(b[19]), .out(u_csamul_pg_rca24_and7_19));
  fa fa_u_csamul_pg_rca24_fa7_19_out(.a(u_csamul_pg_rca24_and7_19[0]), .b(u_csamul_pg_rca24_fa8_18_xor1[0]), .cin(u_csamul_pg_rca24_fa7_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_19_xor1), .fa_or0(u_csamul_pg_rca24_fa7_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_19(.a(a[8]), .b(b[19]), .out(u_csamul_pg_rca24_and8_19));
  fa fa_u_csamul_pg_rca24_fa8_19_out(.a(u_csamul_pg_rca24_and8_19[0]), .b(u_csamul_pg_rca24_fa9_18_xor1[0]), .cin(u_csamul_pg_rca24_fa8_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_19_xor1), .fa_or0(u_csamul_pg_rca24_fa8_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_19(.a(a[9]), .b(b[19]), .out(u_csamul_pg_rca24_and9_19));
  fa fa_u_csamul_pg_rca24_fa9_19_out(.a(u_csamul_pg_rca24_and9_19[0]), .b(u_csamul_pg_rca24_fa10_18_xor1[0]), .cin(u_csamul_pg_rca24_fa9_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_19_xor1), .fa_or0(u_csamul_pg_rca24_fa9_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_19(.a(a[10]), .b(b[19]), .out(u_csamul_pg_rca24_and10_19));
  fa fa_u_csamul_pg_rca24_fa10_19_out(.a(u_csamul_pg_rca24_and10_19[0]), .b(u_csamul_pg_rca24_fa11_18_xor1[0]), .cin(u_csamul_pg_rca24_fa10_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_19_xor1), .fa_or0(u_csamul_pg_rca24_fa10_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_19(.a(a[11]), .b(b[19]), .out(u_csamul_pg_rca24_and11_19));
  fa fa_u_csamul_pg_rca24_fa11_19_out(.a(u_csamul_pg_rca24_and11_19[0]), .b(u_csamul_pg_rca24_fa12_18_xor1[0]), .cin(u_csamul_pg_rca24_fa11_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_19_xor1), .fa_or0(u_csamul_pg_rca24_fa11_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_19(.a(a[12]), .b(b[19]), .out(u_csamul_pg_rca24_and12_19));
  fa fa_u_csamul_pg_rca24_fa12_19_out(.a(u_csamul_pg_rca24_and12_19[0]), .b(u_csamul_pg_rca24_fa13_18_xor1[0]), .cin(u_csamul_pg_rca24_fa12_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_19_xor1), .fa_or0(u_csamul_pg_rca24_fa12_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_19(.a(a[13]), .b(b[19]), .out(u_csamul_pg_rca24_and13_19));
  fa fa_u_csamul_pg_rca24_fa13_19_out(.a(u_csamul_pg_rca24_and13_19[0]), .b(u_csamul_pg_rca24_fa14_18_xor1[0]), .cin(u_csamul_pg_rca24_fa13_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_19_xor1), .fa_or0(u_csamul_pg_rca24_fa13_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_19(.a(a[14]), .b(b[19]), .out(u_csamul_pg_rca24_and14_19));
  fa fa_u_csamul_pg_rca24_fa14_19_out(.a(u_csamul_pg_rca24_and14_19[0]), .b(u_csamul_pg_rca24_fa15_18_xor1[0]), .cin(u_csamul_pg_rca24_fa14_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_19_xor1), .fa_or0(u_csamul_pg_rca24_fa14_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_19(.a(a[15]), .b(b[19]), .out(u_csamul_pg_rca24_and15_19));
  fa fa_u_csamul_pg_rca24_fa15_19_out(.a(u_csamul_pg_rca24_and15_19[0]), .b(u_csamul_pg_rca24_fa16_18_xor1[0]), .cin(u_csamul_pg_rca24_fa15_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_19_xor1), .fa_or0(u_csamul_pg_rca24_fa15_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_19(.a(a[16]), .b(b[19]), .out(u_csamul_pg_rca24_and16_19));
  fa fa_u_csamul_pg_rca24_fa16_19_out(.a(u_csamul_pg_rca24_and16_19[0]), .b(u_csamul_pg_rca24_fa17_18_xor1[0]), .cin(u_csamul_pg_rca24_fa16_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_19_xor1), .fa_or0(u_csamul_pg_rca24_fa16_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_19(.a(a[17]), .b(b[19]), .out(u_csamul_pg_rca24_and17_19));
  fa fa_u_csamul_pg_rca24_fa17_19_out(.a(u_csamul_pg_rca24_and17_19[0]), .b(u_csamul_pg_rca24_fa18_18_xor1[0]), .cin(u_csamul_pg_rca24_fa17_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_19_xor1), .fa_or0(u_csamul_pg_rca24_fa17_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_19(.a(a[18]), .b(b[19]), .out(u_csamul_pg_rca24_and18_19));
  fa fa_u_csamul_pg_rca24_fa18_19_out(.a(u_csamul_pg_rca24_and18_19[0]), .b(u_csamul_pg_rca24_fa19_18_xor1[0]), .cin(u_csamul_pg_rca24_fa18_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_19_xor1), .fa_or0(u_csamul_pg_rca24_fa18_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_19(.a(a[19]), .b(b[19]), .out(u_csamul_pg_rca24_and19_19));
  fa fa_u_csamul_pg_rca24_fa19_19_out(.a(u_csamul_pg_rca24_and19_19[0]), .b(u_csamul_pg_rca24_fa20_18_xor1[0]), .cin(u_csamul_pg_rca24_fa19_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_19_xor1), .fa_or0(u_csamul_pg_rca24_fa19_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_19(.a(a[20]), .b(b[19]), .out(u_csamul_pg_rca24_and20_19));
  fa fa_u_csamul_pg_rca24_fa20_19_out(.a(u_csamul_pg_rca24_and20_19[0]), .b(u_csamul_pg_rca24_fa21_18_xor1[0]), .cin(u_csamul_pg_rca24_fa20_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_19_xor1), .fa_or0(u_csamul_pg_rca24_fa20_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_19(.a(a[21]), .b(b[19]), .out(u_csamul_pg_rca24_and21_19));
  fa fa_u_csamul_pg_rca24_fa21_19_out(.a(u_csamul_pg_rca24_and21_19[0]), .b(u_csamul_pg_rca24_fa22_18_xor1[0]), .cin(u_csamul_pg_rca24_fa21_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_19_xor1), .fa_or0(u_csamul_pg_rca24_fa21_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_19(.a(a[22]), .b(b[19]), .out(u_csamul_pg_rca24_and22_19));
  fa fa_u_csamul_pg_rca24_fa22_19_out(.a(u_csamul_pg_rca24_and22_19[0]), .b(u_csamul_pg_rca24_and23_18[0]), .cin(u_csamul_pg_rca24_fa22_18_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_19_xor1), .fa_or0(u_csamul_pg_rca24_fa22_19_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_19(.a(a[23]), .b(b[19]), .out(u_csamul_pg_rca24_and23_19));
  and_gate and_gate_u_csamul_pg_rca24_and0_20(.a(a[0]), .b(b[20]), .out(u_csamul_pg_rca24_and0_20));
  fa fa_u_csamul_pg_rca24_fa0_20_out(.a(u_csamul_pg_rca24_and0_20[0]), .b(u_csamul_pg_rca24_fa1_19_xor1[0]), .cin(u_csamul_pg_rca24_fa0_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_20_xor1), .fa_or0(u_csamul_pg_rca24_fa0_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_20(.a(a[1]), .b(b[20]), .out(u_csamul_pg_rca24_and1_20));
  fa fa_u_csamul_pg_rca24_fa1_20_out(.a(u_csamul_pg_rca24_and1_20[0]), .b(u_csamul_pg_rca24_fa2_19_xor1[0]), .cin(u_csamul_pg_rca24_fa1_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_20_xor1), .fa_or0(u_csamul_pg_rca24_fa1_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_20(.a(a[2]), .b(b[20]), .out(u_csamul_pg_rca24_and2_20));
  fa fa_u_csamul_pg_rca24_fa2_20_out(.a(u_csamul_pg_rca24_and2_20[0]), .b(u_csamul_pg_rca24_fa3_19_xor1[0]), .cin(u_csamul_pg_rca24_fa2_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_20_xor1), .fa_or0(u_csamul_pg_rca24_fa2_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_20(.a(a[3]), .b(b[20]), .out(u_csamul_pg_rca24_and3_20));
  fa fa_u_csamul_pg_rca24_fa3_20_out(.a(u_csamul_pg_rca24_and3_20[0]), .b(u_csamul_pg_rca24_fa4_19_xor1[0]), .cin(u_csamul_pg_rca24_fa3_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_20_xor1), .fa_or0(u_csamul_pg_rca24_fa3_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_20(.a(a[4]), .b(b[20]), .out(u_csamul_pg_rca24_and4_20));
  fa fa_u_csamul_pg_rca24_fa4_20_out(.a(u_csamul_pg_rca24_and4_20[0]), .b(u_csamul_pg_rca24_fa5_19_xor1[0]), .cin(u_csamul_pg_rca24_fa4_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_20_xor1), .fa_or0(u_csamul_pg_rca24_fa4_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_20(.a(a[5]), .b(b[20]), .out(u_csamul_pg_rca24_and5_20));
  fa fa_u_csamul_pg_rca24_fa5_20_out(.a(u_csamul_pg_rca24_and5_20[0]), .b(u_csamul_pg_rca24_fa6_19_xor1[0]), .cin(u_csamul_pg_rca24_fa5_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_20_xor1), .fa_or0(u_csamul_pg_rca24_fa5_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_20(.a(a[6]), .b(b[20]), .out(u_csamul_pg_rca24_and6_20));
  fa fa_u_csamul_pg_rca24_fa6_20_out(.a(u_csamul_pg_rca24_and6_20[0]), .b(u_csamul_pg_rca24_fa7_19_xor1[0]), .cin(u_csamul_pg_rca24_fa6_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_20_xor1), .fa_or0(u_csamul_pg_rca24_fa6_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_20(.a(a[7]), .b(b[20]), .out(u_csamul_pg_rca24_and7_20));
  fa fa_u_csamul_pg_rca24_fa7_20_out(.a(u_csamul_pg_rca24_and7_20[0]), .b(u_csamul_pg_rca24_fa8_19_xor1[0]), .cin(u_csamul_pg_rca24_fa7_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_20_xor1), .fa_or0(u_csamul_pg_rca24_fa7_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_20(.a(a[8]), .b(b[20]), .out(u_csamul_pg_rca24_and8_20));
  fa fa_u_csamul_pg_rca24_fa8_20_out(.a(u_csamul_pg_rca24_and8_20[0]), .b(u_csamul_pg_rca24_fa9_19_xor1[0]), .cin(u_csamul_pg_rca24_fa8_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_20_xor1), .fa_or0(u_csamul_pg_rca24_fa8_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_20(.a(a[9]), .b(b[20]), .out(u_csamul_pg_rca24_and9_20));
  fa fa_u_csamul_pg_rca24_fa9_20_out(.a(u_csamul_pg_rca24_and9_20[0]), .b(u_csamul_pg_rca24_fa10_19_xor1[0]), .cin(u_csamul_pg_rca24_fa9_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_20_xor1), .fa_or0(u_csamul_pg_rca24_fa9_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_20(.a(a[10]), .b(b[20]), .out(u_csamul_pg_rca24_and10_20));
  fa fa_u_csamul_pg_rca24_fa10_20_out(.a(u_csamul_pg_rca24_and10_20[0]), .b(u_csamul_pg_rca24_fa11_19_xor1[0]), .cin(u_csamul_pg_rca24_fa10_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_20_xor1), .fa_or0(u_csamul_pg_rca24_fa10_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_20(.a(a[11]), .b(b[20]), .out(u_csamul_pg_rca24_and11_20));
  fa fa_u_csamul_pg_rca24_fa11_20_out(.a(u_csamul_pg_rca24_and11_20[0]), .b(u_csamul_pg_rca24_fa12_19_xor1[0]), .cin(u_csamul_pg_rca24_fa11_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_20_xor1), .fa_or0(u_csamul_pg_rca24_fa11_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_20(.a(a[12]), .b(b[20]), .out(u_csamul_pg_rca24_and12_20));
  fa fa_u_csamul_pg_rca24_fa12_20_out(.a(u_csamul_pg_rca24_and12_20[0]), .b(u_csamul_pg_rca24_fa13_19_xor1[0]), .cin(u_csamul_pg_rca24_fa12_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_20_xor1), .fa_or0(u_csamul_pg_rca24_fa12_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_20(.a(a[13]), .b(b[20]), .out(u_csamul_pg_rca24_and13_20));
  fa fa_u_csamul_pg_rca24_fa13_20_out(.a(u_csamul_pg_rca24_and13_20[0]), .b(u_csamul_pg_rca24_fa14_19_xor1[0]), .cin(u_csamul_pg_rca24_fa13_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_20_xor1), .fa_or0(u_csamul_pg_rca24_fa13_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_20(.a(a[14]), .b(b[20]), .out(u_csamul_pg_rca24_and14_20));
  fa fa_u_csamul_pg_rca24_fa14_20_out(.a(u_csamul_pg_rca24_and14_20[0]), .b(u_csamul_pg_rca24_fa15_19_xor1[0]), .cin(u_csamul_pg_rca24_fa14_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_20_xor1), .fa_or0(u_csamul_pg_rca24_fa14_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_20(.a(a[15]), .b(b[20]), .out(u_csamul_pg_rca24_and15_20));
  fa fa_u_csamul_pg_rca24_fa15_20_out(.a(u_csamul_pg_rca24_and15_20[0]), .b(u_csamul_pg_rca24_fa16_19_xor1[0]), .cin(u_csamul_pg_rca24_fa15_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_20_xor1), .fa_or0(u_csamul_pg_rca24_fa15_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_20(.a(a[16]), .b(b[20]), .out(u_csamul_pg_rca24_and16_20));
  fa fa_u_csamul_pg_rca24_fa16_20_out(.a(u_csamul_pg_rca24_and16_20[0]), .b(u_csamul_pg_rca24_fa17_19_xor1[0]), .cin(u_csamul_pg_rca24_fa16_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_20_xor1), .fa_or0(u_csamul_pg_rca24_fa16_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_20(.a(a[17]), .b(b[20]), .out(u_csamul_pg_rca24_and17_20));
  fa fa_u_csamul_pg_rca24_fa17_20_out(.a(u_csamul_pg_rca24_and17_20[0]), .b(u_csamul_pg_rca24_fa18_19_xor1[0]), .cin(u_csamul_pg_rca24_fa17_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_20_xor1), .fa_or0(u_csamul_pg_rca24_fa17_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_20(.a(a[18]), .b(b[20]), .out(u_csamul_pg_rca24_and18_20));
  fa fa_u_csamul_pg_rca24_fa18_20_out(.a(u_csamul_pg_rca24_and18_20[0]), .b(u_csamul_pg_rca24_fa19_19_xor1[0]), .cin(u_csamul_pg_rca24_fa18_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_20_xor1), .fa_or0(u_csamul_pg_rca24_fa18_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_20(.a(a[19]), .b(b[20]), .out(u_csamul_pg_rca24_and19_20));
  fa fa_u_csamul_pg_rca24_fa19_20_out(.a(u_csamul_pg_rca24_and19_20[0]), .b(u_csamul_pg_rca24_fa20_19_xor1[0]), .cin(u_csamul_pg_rca24_fa19_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_20_xor1), .fa_or0(u_csamul_pg_rca24_fa19_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_20(.a(a[20]), .b(b[20]), .out(u_csamul_pg_rca24_and20_20));
  fa fa_u_csamul_pg_rca24_fa20_20_out(.a(u_csamul_pg_rca24_and20_20[0]), .b(u_csamul_pg_rca24_fa21_19_xor1[0]), .cin(u_csamul_pg_rca24_fa20_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_20_xor1), .fa_or0(u_csamul_pg_rca24_fa20_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_20(.a(a[21]), .b(b[20]), .out(u_csamul_pg_rca24_and21_20));
  fa fa_u_csamul_pg_rca24_fa21_20_out(.a(u_csamul_pg_rca24_and21_20[0]), .b(u_csamul_pg_rca24_fa22_19_xor1[0]), .cin(u_csamul_pg_rca24_fa21_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_20_xor1), .fa_or0(u_csamul_pg_rca24_fa21_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_20(.a(a[22]), .b(b[20]), .out(u_csamul_pg_rca24_and22_20));
  fa fa_u_csamul_pg_rca24_fa22_20_out(.a(u_csamul_pg_rca24_and22_20[0]), .b(u_csamul_pg_rca24_and23_19[0]), .cin(u_csamul_pg_rca24_fa22_19_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_20_xor1), .fa_or0(u_csamul_pg_rca24_fa22_20_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_20(.a(a[23]), .b(b[20]), .out(u_csamul_pg_rca24_and23_20));
  and_gate and_gate_u_csamul_pg_rca24_and0_21(.a(a[0]), .b(b[21]), .out(u_csamul_pg_rca24_and0_21));
  fa fa_u_csamul_pg_rca24_fa0_21_out(.a(u_csamul_pg_rca24_and0_21[0]), .b(u_csamul_pg_rca24_fa1_20_xor1[0]), .cin(u_csamul_pg_rca24_fa0_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_21_xor1), .fa_or0(u_csamul_pg_rca24_fa0_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_21(.a(a[1]), .b(b[21]), .out(u_csamul_pg_rca24_and1_21));
  fa fa_u_csamul_pg_rca24_fa1_21_out(.a(u_csamul_pg_rca24_and1_21[0]), .b(u_csamul_pg_rca24_fa2_20_xor1[0]), .cin(u_csamul_pg_rca24_fa1_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_21_xor1), .fa_or0(u_csamul_pg_rca24_fa1_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_21(.a(a[2]), .b(b[21]), .out(u_csamul_pg_rca24_and2_21));
  fa fa_u_csamul_pg_rca24_fa2_21_out(.a(u_csamul_pg_rca24_and2_21[0]), .b(u_csamul_pg_rca24_fa3_20_xor1[0]), .cin(u_csamul_pg_rca24_fa2_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_21_xor1), .fa_or0(u_csamul_pg_rca24_fa2_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_21(.a(a[3]), .b(b[21]), .out(u_csamul_pg_rca24_and3_21));
  fa fa_u_csamul_pg_rca24_fa3_21_out(.a(u_csamul_pg_rca24_and3_21[0]), .b(u_csamul_pg_rca24_fa4_20_xor1[0]), .cin(u_csamul_pg_rca24_fa3_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_21_xor1), .fa_or0(u_csamul_pg_rca24_fa3_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_21(.a(a[4]), .b(b[21]), .out(u_csamul_pg_rca24_and4_21));
  fa fa_u_csamul_pg_rca24_fa4_21_out(.a(u_csamul_pg_rca24_and4_21[0]), .b(u_csamul_pg_rca24_fa5_20_xor1[0]), .cin(u_csamul_pg_rca24_fa4_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_21_xor1), .fa_or0(u_csamul_pg_rca24_fa4_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_21(.a(a[5]), .b(b[21]), .out(u_csamul_pg_rca24_and5_21));
  fa fa_u_csamul_pg_rca24_fa5_21_out(.a(u_csamul_pg_rca24_and5_21[0]), .b(u_csamul_pg_rca24_fa6_20_xor1[0]), .cin(u_csamul_pg_rca24_fa5_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_21_xor1), .fa_or0(u_csamul_pg_rca24_fa5_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_21(.a(a[6]), .b(b[21]), .out(u_csamul_pg_rca24_and6_21));
  fa fa_u_csamul_pg_rca24_fa6_21_out(.a(u_csamul_pg_rca24_and6_21[0]), .b(u_csamul_pg_rca24_fa7_20_xor1[0]), .cin(u_csamul_pg_rca24_fa6_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_21_xor1), .fa_or0(u_csamul_pg_rca24_fa6_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_21(.a(a[7]), .b(b[21]), .out(u_csamul_pg_rca24_and7_21));
  fa fa_u_csamul_pg_rca24_fa7_21_out(.a(u_csamul_pg_rca24_and7_21[0]), .b(u_csamul_pg_rca24_fa8_20_xor1[0]), .cin(u_csamul_pg_rca24_fa7_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_21_xor1), .fa_or0(u_csamul_pg_rca24_fa7_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_21(.a(a[8]), .b(b[21]), .out(u_csamul_pg_rca24_and8_21));
  fa fa_u_csamul_pg_rca24_fa8_21_out(.a(u_csamul_pg_rca24_and8_21[0]), .b(u_csamul_pg_rca24_fa9_20_xor1[0]), .cin(u_csamul_pg_rca24_fa8_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_21_xor1), .fa_or0(u_csamul_pg_rca24_fa8_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_21(.a(a[9]), .b(b[21]), .out(u_csamul_pg_rca24_and9_21));
  fa fa_u_csamul_pg_rca24_fa9_21_out(.a(u_csamul_pg_rca24_and9_21[0]), .b(u_csamul_pg_rca24_fa10_20_xor1[0]), .cin(u_csamul_pg_rca24_fa9_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_21_xor1), .fa_or0(u_csamul_pg_rca24_fa9_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_21(.a(a[10]), .b(b[21]), .out(u_csamul_pg_rca24_and10_21));
  fa fa_u_csamul_pg_rca24_fa10_21_out(.a(u_csamul_pg_rca24_and10_21[0]), .b(u_csamul_pg_rca24_fa11_20_xor1[0]), .cin(u_csamul_pg_rca24_fa10_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_21_xor1), .fa_or0(u_csamul_pg_rca24_fa10_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_21(.a(a[11]), .b(b[21]), .out(u_csamul_pg_rca24_and11_21));
  fa fa_u_csamul_pg_rca24_fa11_21_out(.a(u_csamul_pg_rca24_and11_21[0]), .b(u_csamul_pg_rca24_fa12_20_xor1[0]), .cin(u_csamul_pg_rca24_fa11_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_21_xor1), .fa_or0(u_csamul_pg_rca24_fa11_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_21(.a(a[12]), .b(b[21]), .out(u_csamul_pg_rca24_and12_21));
  fa fa_u_csamul_pg_rca24_fa12_21_out(.a(u_csamul_pg_rca24_and12_21[0]), .b(u_csamul_pg_rca24_fa13_20_xor1[0]), .cin(u_csamul_pg_rca24_fa12_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_21_xor1), .fa_or0(u_csamul_pg_rca24_fa12_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_21(.a(a[13]), .b(b[21]), .out(u_csamul_pg_rca24_and13_21));
  fa fa_u_csamul_pg_rca24_fa13_21_out(.a(u_csamul_pg_rca24_and13_21[0]), .b(u_csamul_pg_rca24_fa14_20_xor1[0]), .cin(u_csamul_pg_rca24_fa13_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_21_xor1), .fa_or0(u_csamul_pg_rca24_fa13_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_21(.a(a[14]), .b(b[21]), .out(u_csamul_pg_rca24_and14_21));
  fa fa_u_csamul_pg_rca24_fa14_21_out(.a(u_csamul_pg_rca24_and14_21[0]), .b(u_csamul_pg_rca24_fa15_20_xor1[0]), .cin(u_csamul_pg_rca24_fa14_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_21_xor1), .fa_or0(u_csamul_pg_rca24_fa14_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_21(.a(a[15]), .b(b[21]), .out(u_csamul_pg_rca24_and15_21));
  fa fa_u_csamul_pg_rca24_fa15_21_out(.a(u_csamul_pg_rca24_and15_21[0]), .b(u_csamul_pg_rca24_fa16_20_xor1[0]), .cin(u_csamul_pg_rca24_fa15_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_21_xor1), .fa_or0(u_csamul_pg_rca24_fa15_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_21(.a(a[16]), .b(b[21]), .out(u_csamul_pg_rca24_and16_21));
  fa fa_u_csamul_pg_rca24_fa16_21_out(.a(u_csamul_pg_rca24_and16_21[0]), .b(u_csamul_pg_rca24_fa17_20_xor1[0]), .cin(u_csamul_pg_rca24_fa16_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_21_xor1), .fa_or0(u_csamul_pg_rca24_fa16_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_21(.a(a[17]), .b(b[21]), .out(u_csamul_pg_rca24_and17_21));
  fa fa_u_csamul_pg_rca24_fa17_21_out(.a(u_csamul_pg_rca24_and17_21[0]), .b(u_csamul_pg_rca24_fa18_20_xor1[0]), .cin(u_csamul_pg_rca24_fa17_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_21_xor1), .fa_or0(u_csamul_pg_rca24_fa17_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_21(.a(a[18]), .b(b[21]), .out(u_csamul_pg_rca24_and18_21));
  fa fa_u_csamul_pg_rca24_fa18_21_out(.a(u_csamul_pg_rca24_and18_21[0]), .b(u_csamul_pg_rca24_fa19_20_xor1[0]), .cin(u_csamul_pg_rca24_fa18_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_21_xor1), .fa_or0(u_csamul_pg_rca24_fa18_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_21(.a(a[19]), .b(b[21]), .out(u_csamul_pg_rca24_and19_21));
  fa fa_u_csamul_pg_rca24_fa19_21_out(.a(u_csamul_pg_rca24_and19_21[0]), .b(u_csamul_pg_rca24_fa20_20_xor1[0]), .cin(u_csamul_pg_rca24_fa19_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_21_xor1), .fa_or0(u_csamul_pg_rca24_fa19_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_21(.a(a[20]), .b(b[21]), .out(u_csamul_pg_rca24_and20_21));
  fa fa_u_csamul_pg_rca24_fa20_21_out(.a(u_csamul_pg_rca24_and20_21[0]), .b(u_csamul_pg_rca24_fa21_20_xor1[0]), .cin(u_csamul_pg_rca24_fa20_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_21_xor1), .fa_or0(u_csamul_pg_rca24_fa20_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_21(.a(a[21]), .b(b[21]), .out(u_csamul_pg_rca24_and21_21));
  fa fa_u_csamul_pg_rca24_fa21_21_out(.a(u_csamul_pg_rca24_and21_21[0]), .b(u_csamul_pg_rca24_fa22_20_xor1[0]), .cin(u_csamul_pg_rca24_fa21_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_21_xor1), .fa_or0(u_csamul_pg_rca24_fa21_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_21(.a(a[22]), .b(b[21]), .out(u_csamul_pg_rca24_and22_21));
  fa fa_u_csamul_pg_rca24_fa22_21_out(.a(u_csamul_pg_rca24_and22_21[0]), .b(u_csamul_pg_rca24_and23_20[0]), .cin(u_csamul_pg_rca24_fa22_20_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_21_xor1), .fa_or0(u_csamul_pg_rca24_fa22_21_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_21(.a(a[23]), .b(b[21]), .out(u_csamul_pg_rca24_and23_21));
  and_gate and_gate_u_csamul_pg_rca24_and0_22(.a(a[0]), .b(b[22]), .out(u_csamul_pg_rca24_and0_22));
  fa fa_u_csamul_pg_rca24_fa0_22_out(.a(u_csamul_pg_rca24_and0_22[0]), .b(u_csamul_pg_rca24_fa1_21_xor1[0]), .cin(u_csamul_pg_rca24_fa0_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_22_xor1), .fa_or0(u_csamul_pg_rca24_fa0_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_22(.a(a[1]), .b(b[22]), .out(u_csamul_pg_rca24_and1_22));
  fa fa_u_csamul_pg_rca24_fa1_22_out(.a(u_csamul_pg_rca24_and1_22[0]), .b(u_csamul_pg_rca24_fa2_21_xor1[0]), .cin(u_csamul_pg_rca24_fa1_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_22_xor1), .fa_or0(u_csamul_pg_rca24_fa1_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_22(.a(a[2]), .b(b[22]), .out(u_csamul_pg_rca24_and2_22));
  fa fa_u_csamul_pg_rca24_fa2_22_out(.a(u_csamul_pg_rca24_and2_22[0]), .b(u_csamul_pg_rca24_fa3_21_xor1[0]), .cin(u_csamul_pg_rca24_fa2_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_22_xor1), .fa_or0(u_csamul_pg_rca24_fa2_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_22(.a(a[3]), .b(b[22]), .out(u_csamul_pg_rca24_and3_22));
  fa fa_u_csamul_pg_rca24_fa3_22_out(.a(u_csamul_pg_rca24_and3_22[0]), .b(u_csamul_pg_rca24_fa4_21_xor1[0]), .cin(u_csamul_pg_rca24_fa3_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_22_xor1), .fa_or0(u_csamul_pg_rca24_fa3_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_22(.a(a[4]), .b(b[22]), .out(u_csamul_pg_rca24_and4_22));
  fa fa_u_csamul_pg_rca24_fa4_22_out(.a(u_csamul_pg_rca24_and4_22[0]), .b(u_csamul_pg_rca24_fa5_21_xor1[0]), .cin(u_csamul_pg_rca24_fa4_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_22_xor1), .fa_or0(u_csamul_pg_rca24_fa4_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_22(.a(a[5]), .b(b[22]), .out(u_csamul_pg_rca24_and5_22));
  fa fa_u_csamul_pg_rca24_fa5_22_out(.a(u_csamul_pg_rca24_and5_22[0]), .b(u_csamul_pg_rca24_fa6_21_xor1[0]), .cin(u_csamul_pg_rca24_fa5_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_22_xor1), .fa_or0(u_csamul_pg_rca24_fa5_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_22(.a(a[6]), .b(b[22]), .out(u_csamul_pg_rca24_and6_22));
  fa fa_u_csamul_pg_rca24_fa6_22_out(.a(u_csamul_pg_rca24_and6_22[0]), .b(u_csamul_pg_rca24_fa7_21_xor1[0]), .cin(u_csamul_pg_rca24_fa6_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_22_xor1), .fa_or0(u_csamul_pg_rca24_fa6_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_22(.a(a[7]), .b(b[22]), .out(u_csamul_pg_rca24_and7_22));
  fa fa_u_csamul_pg_rca24_fa7_22_out(.a(u_csamul_pg_rca24_and7_22[0]), .b(u_csamul_pg_rca24_fa8_21_xor1[0]), .cin(u_csamul_pg_rca24_fa7_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_22_xor1), .fa_or0(u_csamul_pg_rca24_fa7_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_22(.a(a[8]), .b(b[22]), .out(u_csamul_pg_rca24_and8_22));
  fa fa_u_csamul_pg_rca24_fa8_22_out(.a(u_csamul_pg_rca24_and8_22[0]), .b(u_csamul_pg_rca24_fa9_21_xor1[0]), .cin(u_csamul_pg_rca24_fa8_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_22_xor1), .fa_or0(u_csamul_pg_rca24_fa8_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_22(.a(a[9]), .b(b[22]), .out(u_csamul_pg_rca24_and9_22));
  fa fa_u_csamul_pg_rca24_fa9_22_out(.a(u_csamul_pg_rca24_and9_22[0]), .b(u_csamul_pg_rca24_fa10_21_xor1[0]), .cin(u_csamul_pg_rca24_fa9_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_22_xor1), .fa_or0(u_csamul_pg_rca24_fa9_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_22(.a(a[10]), .b(b[22]), .out(u_csamul_pg_rca24_and10_22));
  fa fa_u_csamul_pg_rca24_fa10_22_out(.a(u_csamul_pg_rca24_and10_22[0]), .b(u_csamul_pg_rca24_fa11_21_xor1[0]), .cin(u_csamul_pg_rca24_fa10_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_22_xor1), .fa_or0(u_csamul_pg_rca24_fa10_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_22(.a(a[11]), .b(b[22]), .out(u_csamul_pg_rca24_and11_22));
  fa fa_u_csamul_pg_rca24_fa11_22_out(.a(u_csamul_pg_rca24_and11_22[0]), .b(u_csamul_pg_rca24_fa12_21_xor1[0]), .cin(u_csamul_pg_rca24_fa11_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_22_xor1), .fa_or0(u_csamul_pg_rca24_fa11_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_22(.a(a[12]), .b(b[22]), .out(u_csamul_pg_rca24_and12_22));
  fa fa_u_csamul_pg_rca24_fa12_22_out(.a(u_csamul_pg_rca24_and12_22[0]), .b(u_csamul_pg_rca24_fa13_21_xor1[0]), .cin(u_csamul_pg_rca24_fa12_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_22_xor1), .fa_or0(u_csamul_pg_rca24_fa12_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_22(.a(a[13]), .b(b[22]), .out(u_csamul_pg_rca24_and13_22));
  fa fa_u_csamul_pg_rca24_fa13_22_out(.a(u_csamul_pg_rca24_and13_22[0]), .b(u_csamul_pg_rca24_fa14_21_xor1[0]), .cin(u_csamul_pg_rca24_fa13_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_22_xor1), .fa_or0(u_csamul_pg_rca24_fa13_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_22(.a(a[14]), .b(b[22]), .out(u_csamul_pg_rca24_and14_22));
  fa fa_u_csamul_pg_rca24_fa14_22_out(.a(u_csamul_pg_rca24_and14_22[0]), .b(u_csamul_pg_rca24_fa15_21_xor1[0]), .cin(u_csamul_pg_rca24_fa14_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_22_xor1), .fa_or0(u_csamul_pg_rca24_fa14_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_22(.a(a[15]), .b(b[22]), .out(u_csamul_pg_rca24_and15_22));
  fa fa_u_csamul_pg_rca24_fa15_22_out(.a(u_csamul_pg_rca24_and15_22[0]), .b(u_csamul_pg_rca24_fa16_21_xor1[0]), .cin(u_csamul_pg_rca24_fa15_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_22_xor1), .fa_or0(u_csamul_pg_rca24_fa15_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_22(.a(a[16]), .b(b[22]), .out(u_csamul_pg_rca24_and16_22));
  fa fa_u_csamul_pg_rca24_fa16_22_out(.a(u_csamul_pg_rca24_and16_22[0]), .b(u_csamul_pg_rca24_fa17_21_xor1[0]), .cin(u_csamul_pg_rca24_fa16_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_22_xor1), .fa_or0(u_csamul_pg_rca24_fa16_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_22(.a(a[17]), .b(b[22]), .out(u_csamul_pg_rca24_and17_22));
  fa fa_u_csamul_pg_rca24_fa17_22_out(.a(u_csamul_pg_rca24_and17_22[0]), .b(u_csamul_pg_rca24_fa18_21_xor1[0]), .cin(u_csamul_pg_rca24_fa17_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_22_xor1), .fa_or0(u_csamul_pg_rca24_fa17_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_22(.a(a[18]), .b(b[22]), .out(u_csamul_pg_rca24_and18_22));
  fa fa_u_csamul_pg_rca24_fa18_22_out(.a(u_csamul_pg_rca24_and18_22[0]), .b(u_csamul_pg_rca24_fa19_21_xor1[0]), .cin(u_csamul_pg_rca24_fa18_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_22_xor1), .fa_or0(u_csamul_pg_rca24_fa18_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_22(.a(a[19]), .b(b[22]), .out(u_csamul_pg_rca24_and19_22));
  fa fa_u_csamul_pg_rca24_fa19_22_out(.a(u_csamul_pg_rca24_and19_22[0]), .b(u_csamul_pg_rca24_fa20_21_xor1[0]), .cin(u_csamul_pg_rca24_fa19_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_22_xor1), .fa_or0(u_csamul_pg_rca24_fa19_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_22(.a(a[20]), .b(b[22]), .out(u_csamul_pg_rca24_and20_22));
  fa fa_u_csamul_pg_rca24_fa20_22_out(.a(u_csamul_pg_rca24_and20_22[0]), .b(u_csamul_pg_rca24_fa21_21_xor1[0]), .cin(u_csamul_pg_rca24_fa20_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_22_xor1), .fa_or0(u_csamul_pg_rca24_fa20_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_22(.a(a[21]), .b(b[22]), .out(u_csamul_pg_rca24_and21_22));
  fa fa_u_csamul_pg_rca24_fa21_22_out(.a(u_csamul_pg_rca24_and21_22[0]), .b(u_csamul_pg_rca24_fa22_21_xor1[0]), .cin(u_csamul_pg_rca24_fa21_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_22_xor1), .fa_or0(u_csamul_pg_rca24_fa21_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_22(.a(a[22]), .b(b[22]), .out(u_csamul_pg_rca24_and22_22));
  fa fa_u_csamul_pg_rca24_fa22_22_out(.a(u_csamul_pg_rca24_and22_22[0]), .b(u_csamul_pg_rca24_and23_21[0]), .cin(u_csamul_pg_rca24_fa22_21_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_22_xor1), .fa_or0(u_csamul_pg_rca24_fa22_22_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_22(.a(a[23]), .b(b[22]), .out(u_csamul_pg_rca24_and23_22));
  and_gate and_gate_u_csamul_pg_rca24_and0_23(.a(a[0]), .b(b[23]), .out(u_csamul_pg_rca24_and0_23));
  fa fa_u_csamul_pg_rca24_fa0_23_out(.a(u_csamul_pg_rca24_and0_23[0]), .b(u_csamul_pg_rca24_fa1_22_xor1[0]), .cin(u_csamul_pg_rca24_fa0_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa0_23_xor1), .fa_or0(u_csamul_pg_rca24_fa0_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and1_23(.a(a[1]), .b(b[23]), .out(u_csamul_pg_rca24_and1_23));
  fa fa_u_csamul_pg_rca24_fa1_23_out(.a(u_csamul_pg_rca24_and1_23[0]), .b(u_csamul_pg_rca24_fa2_22_xor1[0]), .cin(u_csamul_pg_rca24_fa1_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa1_23_xor1), .fa_or0(u_csamul_pg_rca24_fa1_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and2_23(.a(a[2]), .b(b[23]), .out(u_csamul_pg_rca24_and2_23));
  fa fa_u_csamul_pg_rca24_fa2_23_out(.a(u_csamul_pg_rca24_and2_23[0]), .b(u_csamul_pg_rca24_fa3_22_xor1[0]), .cin(u_csamul_pg_rca24_fa2_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa2_23_xor1), .fa_or0(u_csamul_pg_rca24_fa2_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and3_23(.a(a[3]), .b(b[23]), .out(u_csamul_pg_rca24_and3_23));
  fa fa_u_csamul_pg_rca24_fa3_23_out(.a(u_csamul_pg_rca24_and3_23[0]), .b(u_csamul_pg_rca24_fa4_22_xor1[0]), .cin(u_csamul_pg_rca24_fa3_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa3_23_xor1), .fa_or0(u_csamul_pg_rca24_fa3_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and4_23(.a(a[4]), .b(b[23]), .out(u_csamul_pg_rca24_and4_23));
  fa fa_u_csamul_pg_rca24_fa4_23_out(.a(u_csamul_pg_rca24_and4_23[0]), .b(u_csamul_pg_rca24_fa5_22_xor1[0]), .cin(u_csamul_pg_rca24_fa4_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa4_23_xor1), .fa_or0(u_csamul_pg_rca24_fa4_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and5_23(.a(a[5]), .b(b[23]), .out(u_csamul_pg_rca24_and5_23));
  fa fa_u_csamul_pg_rca24_fa5_23_out(.a(u_csamul_pg_rca24_and5_23[0]), .b(u_csamul_pg_rca24_fa6_22_xor1[0]), .cin(u_csamul_pg_rca24_fa5_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa5_23_xor1), .fa_or0(u_csamul_pg_rca24_fa5_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and6_23(.a(a[6]), .b(b[23]), .out(u_csamul_pg_rca24_and6_23));
  fa fa_u_csamul_pg_rca24_fa6_23_out(.a(u_csamul_pg_rca24_and6_23[0]), .b(u_csamul_pg_rca24_fa7_22_xor1[0]), .cin(u_csamul_pg_rca24_fa6_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa6_23_xor1), .fa_or0(u_csamul_pg_rca24_fa6_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and7_23(.a(a[7]), .b(b[23]), .out(u_csamul_pg_rca24_and7_23));
  fa fa_u_csamul_pg_rca24_fa7_23_out(.a(u_csamul_pg_rca24_and7_23[0]), .b(u_csamul_pg_rca24_fa8_22_xor1[0]), .cin(u_csamul_pg_rca24_fa7_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa7_23_xor1), .fa_or0(u_csamul_pg_rca24_fa7_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and8_23(.a(a[8]), .b(b[23]), .out(u_csamul_pg_rca24_and8_23));
  fa fa_u_csamul_pg_rca24_fa8_23_out(.a(u_csamul_pg_rca24_and8_23[0]), .b(u_csamul_pg_rca24_fa9_22_xor1[0]), .cin(u_csamul_pg_rca24_fa8_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa8_23_xor1), .fa_or0(u_csamul_pg_rca24_fa8_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and9_23(.a(a[9]), .b(b[23]), .out(u_csamul_pg_rca24_and9_23));
  fa fa_u_csamul_pg_rca24_fa9_23_out(.a(u_csamul_pg_rca24_and9_23[0]), .b(u_csamul_pg_rca24_fa10_22_xor1[0]), .cin(u_csamul_pg_rca24_fa9_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa9_23_xor1), .fa_or0(u_csamul_pg_rca24_fa9_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and10_23(.a(a[10]), .b(b[23]), .out(u_csamul_pg_rca24_and10_23));
  fa fa_u_csamul_pg_rca24_fa10_23_out(.a(u_csamul_pg_rca24_and10_23[0]), .b(u_csamul_pg_rca24_fa11_22_xor1[0]), .cin(u_csamul_pg_rca24_fa10_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa10_23_xor1), .fa_or0(u_csamul_pg_rca24_fa10_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and11_23(.a(a[11]), .b(b[23]), .out(u_csamul_pg_rca24_and11_23));
  fa fa_u_csamul_pg_rca24_fa11_23_out(.a(u_csamul_pg_rca24_and11_23[0]), .b(u_csamul_pg_rca24_fa12_22_xor1[0]), .cin(u_csamul_pg_rca24_fa11_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa11_23_xor1), .fa_or0(u_csamul_pg_rca24_fa11_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and12_23(.a(a[12]), .b(b[23]), .out(u_csamul_pg_rca24_and12_23));
  fa fa_u_csamul_pg_rca24_fa12_23_out(.a(u_csamul_pg_rca24_and12_23[0]), .b(u_csamul_pg_rca24_fa13_22_xor1[0]), .cin(u_csamul_pg_rca24_fa12_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa12_23_xor1), .fa_or0(u_csamul_pg_rca24_fa12_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and13_23(.a(a[13]), .b(b[23]), .out(u_csamul_pg_rca24_and13_23));
  fa fa_u_csamul_pg_rca24_fa13_23_out(.a(u_csamul_pg_rca24_and13_23[0]), .b(u_csamul_pg_rca24_fa14_22_xor1[0]), .cin(u_csamul_pg_rca24_fa13_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa13_23_xor1), .fa_or0(u_csamul_pg_rca24_fa13_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and14_23(.a(a[14]), .b(b[23]), .out(u_csamul_pg_rca24_and14_23));
  fa fa_u_csamul_pg_rca24_fa14_23_out(.a(u_csamul_pg_rca24_and14_23[0]), .b(u_csamul_pg_rca24_fa15_22_xor1[0]), .cin(u_csamul_pg_rca24_fa14_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa14_23_xor1), .fa_or0(u_csamul_pg_rca24_fa14_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and15_23(.a(a[15]), .b(b[23]), .out(u_csamul_pg_rca24_and15_23));
  fa fa_u_csamul_pg_rca24_fa15_23_out(.a(u_csamul_pg_rca24_and15_23[0]), .b(u_csamul_pg_rca24_fa16_22_xor1[0]), .cin(u_csamul_pg_rca24_fa15_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa15_23_xor1), .fa_or0(u_csamul_pg_rca24_fa15_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and16_23(.a(a[16]), .b(b[23]), .out(u_csamul_pg_rca24_and16_23));
  fa fa_u_csamul_pg_rca24_fa16_23_out(.a(u_csamul_pg_rca24_and16_23[0]), .b(u_csamul_pg_rca24_fa17_22_xor1[0]), .cin(u_csamul_pg_rca24_fa16_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa16_23_xor1), .fa_or0(u_csamul_pg_rca24_fa16_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and17_23(.a(a[17]), .b(b[23]), .out(u_csamul_pg_rca24_and17_23));
  fa fa_u_csamul_pg_rca24_fa17_23_out(.a(u_csamul_pg_rca24_and17_23[0]), .b(u_csamul_pg_rca24_fa18_22_xor1[0]), .cin(u_csamul_pg_rca24_fa17_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa17_23_xor1), .fa_or0(u_csamul_pg_rca24_fa17_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and18_23(.a(a[18]), .b(b[23]), .out(u_csamul_pg_rca24_and18_23));
  fa fa_u_csamul_pg_rca24_fa18_23_out(.a(u_csamul_pg_rca24_and18_23[0]), .b(u_csamul_pg_rca24_fa19_22_xor1[0]), .cin(u_csamul_pg_rca24_fa18_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa18_23_xor1), .fa_or0(u_csamul_pg_rca24_fa18_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and19_23(.a(a[19]), .b(b[23]), .out(u_csamul_pg_rca24_and19_23));
  fa fa_u_csamul_pg_rca24_fa19_23_out(.a(u_csamul_pg_rca24_and19_23[0]), .b(u_csamul_pg_rca24_fa20_22_xor1[0]), .cin(u_csamul_pg_rca24_fa19_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa19_23_xor1), .fa_or0(u_csamul_pg_rca24_fa19_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and20_23(.a(a[20]), .b(b[23]), .out(u_csamul_pg_rca24_and20_23));
  fa fa_u_csamul_pg_rca24_fa20_23_out(.a(u_csamul_pg_rca24_and20_23[0]), .b(u_csamul_pg_rca24_fa21_22_xor1[0]), .cin(u_csamul_pg_rca24_fa20_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa20_23_xor1), .fa_or0(u_csamul_pg_rca24_fa20_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and21_23(.a(a[21]), .b(b[23]), .out(u_csamul_pg_rca24_and21_23));
  fa fa_u_csamul_pg_rca24_fa21_23_out(.a(u_csamul_pg_rca24_and21_23[0]), .b(u_csamul_pg_rca24_fa22_22_xor1[0]), .cin(u_csamul_pg_rca24_fa21_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa21_23_xor1), .fa_or0(u_csamul_pg_rca24_fa21_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and22_23(.a(a[22]), .b(b[23]), .out(u_csamul_pg_rca24_and22_23));
  fa fa_u_csamul_pg_rca24_fa22_23_out(.a(u_csamul_pg_rca24_and22_23[0]), .b(u_csamul_pg_rca24_and23_22[0]), .cin(u_csamul_pg_rca24_fa22_22_or0[0]), .fa_xor1(u_csamul_pg_rca24_fa22_23_xor1), .fa_or0(u_csamul_pg_rca24_fa22_23_or0));
  and_gate and_gate_u_csamul_pg_rca24_and23_23(.a(a[23]), .b(b[23]), .out(u_csamul_pg_rca24_and23_23));
  assign u_csamul_pg_rca24_u_pg_rca24_a[0] = u_csamul_pg_rca24_fa1_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[1] = u_csamul_pg_rca24_fa2_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[2] = u_csamul_pg_rca24_fa3_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[3] = u_csamul_pg_rca24_fa4_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[4] = u_csamul_pg_rca24_fa5_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[5] = u_csamul_pg_rca24_fa6_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[6] = u_csamul_pg_rca24_fa7_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[7] = u_csamul_pg_rca24_fa8_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[8] = u_csamul_pg_rca24_fa9_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[9] = u_csamul_pg_rca24_fa10_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[10] = u_csamul_pg_rca24_fa11_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[11] = u_csamul_pg_rca24_fa12_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[12] = u_csamul_pg_rca24_fa13_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[13] = u_csamul_pg_rca24_fa14_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[14] = u_csamul_pg_rca24_fa15_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[15] = u_csamul_pg_rca24_fa16_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[16] = u_csamul_pg_rca24_fa17_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[17] = u_csamul_pg_rca24_fa18_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[18] = u_csamul_pg_rca24_fa19_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[19] = u_csamul_pg_rca24_fa20_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[20] = u_csamul_pg_rca24_fa21_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[21] = u_csamul_pg_rca24_fa22_23_xor1[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[22] = u_csamul_pg_rca24_and23_23[0];
  assign u_csamul_pg_rca24_u_pg_rca24_a[23] = 1'b0;
  assign u_csamul_pg_rca24_u_pg_rca24_b[0] = u_csamul_pg_rca24_fa0_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[1] = u_csamul_pg_rca24_fa1_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[2] = u_csamul_pg_rca24_fa2_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[3] = u_csamul_pg_rca24_fa3_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[4] = u_csamul_pg_rca24_fa4_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[5] = u_csamul_pg_rca24_fa5_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[6] = u_csamul_pg_rca24_fa6_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[7] = u_csamul_pg_rca24_fa7_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[8] = u_csamul_pg_rca24_fa8_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[9] = u_csamul_pg_rca24_fa9_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[10] = u_csamul_pg_rca24_fa10_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[11] = u_csamul_pg_rca24_fa11_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[12] = u_csamul_pg_rca24_fa12_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[13] = u_csamul_pg_rca24_fa13_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[14] = u_csamul_pg_rca24_fa14_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[15] = u_csamul_pg_rca24_fa15_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[16] = u_csamul_pg_rca24_fa16_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[17] = u_csamul_pg_rca24_fa17_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[18] = u_csamul_pg_rca24_fa18_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[19] = u_csamul_pg_rca24_fa19_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[20] = u_csamul_pg_rca24_fa20_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[21] = u_csamul_pg_rca24_fa21_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[22] = u_csamul_pg_rca24_fa22_23_or0[0];
  assign u_csamul_pg_rca24_u_pg_rca24_b[23] = 1'b0;
  u_pg_rca24 u_pg_rca24_u_csamul_pg_rca24_u_pg_rca24_out(.a(u_csamul_pg_rca24_u_pg_rca24_a), .b(u_csamul_pg_rca24_u_pg_rca24_b), .u_pg_rca24_out(u_csamul_pg_rca24_u_pg_rca24_out));

  assign u_csamul_pg_rca24_out[0] = u_csamul_pg_rca24_and0_0[0];
  assign u_csamul_pg_rca24_out[1] = u_csamul_pg_rca24_ha0_1_xor0[0];
  assign u_csamul_pg_rca24_out[2] = u_csamul_pg_rca24_fa0_2_xor1[0];
  assign u_csamul_pg_rca24_out[3] = u_csamul_pg_rca24_fa0_3_xor1[0];
  assign u_csamul_pg_rca24_out[4] = u_csamul_pg_rca24_fa0_4_xor1[0];
  assign u_csamul_pg_rca24_out[5] = u_csamul_pg_rca24_fa0_5_xor1[0];
  assign u_csamul_pg_rca24_out[6] = u_csamul_pg_rca24_fa0_6_xor1[0];
  assign u_csamul_pg_rca24_out[7] = u_csamul_pg_rca24_fa0_7_xor1[0];
  assign u_csamul_pg_rca24_out[8] = u_csamul_pg_rca24_fa0_8_xor1[0];
  assign u_csamul_pg_rca24_out[9] = u_csamul_pg_rca24_fa0_9_xor1[0];
  assign u_csamul_pg_rca24_out[10] = u_csamul_pg_rca24_fa0_10_xor1[0];
  assign u_csamul_pg_rca24_out[11] = u_csamul_pg_rca24_fa0_11_xor1[0];
  assign u_csamul_pg_rca24_out[12] = u_csamul_pg_rca24_fa0_12_xor1[0];
  assign u_csamul_pg_rca24_out[13] = u_csamul_pg_rca24_fa0_13_xor1[0];
  assign u_csamul_pg_rca24_out[14] = u_csamul_pg_rca24_fa0_14_xor1[0];
  assign u_csamul_pg_rca24_out[15] = u_csamul_pg_rca24_fa0_15_xor1[0];
  assign u_csamul_pg_rca24_out[16] = u_csamul_pg_rca24_fa0_16_xor1[0];
  assign u_csamul_pg_rca24_out[17] = u_csamul_pg_rca24_fa0_17_xor1[0];
  assign u_csamul_pg_rca24_out[18] = u_csamul_pg_rca24_fa0_18_xor1[0];
  assign u_csamul_pg_rca24_out[19] = u_csamul_pg_rca24_fa0_19_xor1[0];
  assign u_csamul_pg_rca24_out[20] = u_csamul_pg_rca24_fa0_20_xor1[0];
  assign u_csamul_pg_rca24_out[21] = u_csamul_pg_rca24_fa0_21_xor1[0];
  assign u_csamul_pg_rca24_out[22] = u_csamul_pg_rca24_fa0_22_xor1[0];
  assign u_csamul_pg_rca24_out[23] = u_csamul_pg_rca24_fa0_23_xor1[0];
  assign u_csamul_pg_rca24_out[24] = u_csamul_pg_rca24_u_pg_rca24_out[0];
  assign u_csamul_pg_rca24_out[25] = u_csamul_pg_rca24_u_pg_rca24_out[1];
  assign u_csamul_pg_rca24_out[26] = u_csamul_pg_rca24_u_pg_rca24_out[2];
  assign u_csamul_pg_rca24_out[27] = u_csamul_pg_rca24_u_pg_rca24_out[3];
  assign u_csamul_pg_rca24_out[28] = u_csamul_pg_rca24_u_pg_rca24_out[4];
  assign u_csamul_pg_rca24_out[29] = u_csamul_pg_rca24_u_pg_rca24_out[5];
  assign u_csamul_pg_rca24_out[30] = u_csamul_pg_rca24_u_pg_rca24_out[6];
  assign u_csamul_pg_rca24_out[31] = u_csamul_pg_rca24_u_pg_rca24_out[7];
  assign u_csamul_pg_rca24_out[32] = u_csamul_pg_rca24_u_pg_rca24_out[8];
  assign u_csamul_pg_rca24_out[33] = u_csamul_pg_rca24_u_pg_rca24_out[9];
  assign u_csamul_pg_rca24_out[34] = u_csamul_pg_rca24_u_pg_rca24_out[10];
  assign u_csamul_pg_rca24_out[35] = u_csamul_pg_rca24_u_pg_rca24_out[11];
  assign u_csamul_pg_rca24_out[36] = u_csamul_pg_rca24_u_pg_rca24_out[12];
  assign u_csamul_pg_rca24_out[37] = u_csamul_pg_rca24_u_pg_rca24_out[13];
  assign u_csamul_pg_rca24_out[38] = u_csamul_pg_rca24_u_pg_rca24_out[14];
  assign u_csamul_pg_rca24_out[39] = u_csamul_pg_rca24_u_pg_rca24_out[15];
  assign u_csamul_pg_rca24_out[40] = u_csamul_pg_rca24_u_pg_rca24_out[16];
  assign u_csamul_pg_rca24_out[41] = u_csamul_pg_rca24_u_pg_rca24_out[17];
  assign u_csamul_pg_rca24_out[42] = u_csamul_pg_rca24_u_pg_rca24_out[18];
  assign u_csamul_pg_rca24_out[43] = u_csamul_pg_rca24_u_pg_rca24_out[19];
  assign u_csamul_pg_rca24_out[44] = u_csamul_pg_rca24_u_pg_rca24_out[20];
  assign u_csamul_pg_rca24_out[45] = u_csamul_pg_rca24_u_pg_rca24_out[21];
  assign u_csamul_pg_rca24_out[46] = u_csamul_pg_rca24_u_pg_rca24_out[22];
  assign u_csamul_pg_rca24_out[47] = u_csamul_pg_rca24_u_pg_rca24_out[23];
endmodule