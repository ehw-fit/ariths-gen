module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module u_rca12(input [11:0] a, input [11:0] b, output [12:0] u_rca12_out);
  wire [0:0] u_rca12_ha_xor0;
  wire [0:0] u_rca12_ha_and0;
  wire [0:0] u_rca12_fa1_xor1;
  wire [0:0] u_rca12_fa1_or0;
  wire [0:0] u_rca12_fa2_xor1;
  wire [0:0] u_rca12_fa2_or0;
  wire [0:0] u_rca12_fa3_xor1;
  wire [0:0] u_rca12_fa3_or0;
  wire [0:0] u_rca12_fa4_xor1;
  wire [0:0] u_rca12_fa4_or0;
  wire [0:0] u_rca12_fa5_xor1;
  wire [0:0] u_rca12_fa5_or0;
  wire [0:0] u_rca12_fa6_xor1;
  wire [0:0] u_rca12_fa6_or0;
  wire [0:0] u_rca12_fa7_xor1;
  wire [0:0] u_rca12_fa7_or0;
  wire [0:0] u_rca12_fa8_xor1;
  wire [0:0] u_rca12_fa8_or0;
  wire [0:0] u_rca12_fa9_xor1;
  wire [0:0] u_rca12_fa9_or0;
  wire [0:0] u_rca12_fa10_xor1;
  wire [0:0] u_rca12_fa10_or0;
  wire [0:0] u_rca12_fa11_xor1;
  wire [0:0] u_rca12_fa11_or0;

  ha ha_u_rca12_ha_out(.a(a[0]), .b(b[0]), .ha_xor0(u_rca12_ha_xor0), .ha_and0(u_rca12_ha_and0));
  fa fa_u_rca12_fa1_out(.a(a[1]), .b(b[1]), .cin(u_rca12_ha_and0[0]), .fa_xor1(u_rca12_fa1_xor1), .fa_or0(u_rca12_fa1_or0));
  fa fa_u_rca12_fa2_out(.a(a[2]), .b(b[2]), .cin(u_rca12_fa1_or0[0]), .fa_xor1(u_rca12_fa2_xor1), .fa_or0(u_rca12_fa2_or0));
  fa fa_u_rca12_fa3_out(.a(a[3]), .b(b[3]), .cin(u_rca12_fa2_or0[0]), .fa_xor1(u_rca12_fa3_xor1), .fa_or0(u_rca12_fa3_or0));
  fa fa_u_rca12_fa4_out(.a(a[4]), .b(b[4]), .cin(u_rca12_fa3_or0[0]), .fa_xor1(u_rca12_fa4_xor1), .fa_or0(u_rca12_fa4_or0));
  fa fa_u_rca12_fa5_out(.a(a[5]), .b(b[5]), .cin(u_rca12_fa4_or0[0]), .fa_xor1(u_rca12_fa5_xor1), .fa_or0(u_rca12_fa5_or0));
  fa fa_u_rca12_fa6_out(.a(a[6]), .b(b[6]), .cin(u_rca12_fa5_or0[0]), .fa_xor1(u_rca12_fa6_xor1), .fa_or0(u_rca12_fa6_or0));
  fa fa_u_rca12_fa7_out(.a(a[7]), .b(b[7]), .cin(u_rca12_fa6_or0[0]), .fa_xor1(u_rca12_fa7_xor1), .fa_or0(u_rca12_fa7_or0));
  fa fa_u_rca12_fa8_out(.a(a[8]), .b(b[8]), .cin(u_rca12_fa7_or0[0]), .fa_xor1(u_rca12_fa8_xor1), .fa_or0(u_rca12_fa8_or0));
  fa fa_u_rca12_fa9_out(.a(a[9]), .b(b[9]), .cin(u_rca12_fa8_or0[0]), .fa_xor1(u_rca12_fa9_xor1), .fa_or0(u_rca12_fa9_or0));
  fa fa_u_rca12_fa10_out(.a(a[10]), .b(b[10]), .cin(u_rca12_fa9_or0[0]), .fa_xor1(u_rca12_fa10_xor1), .fa_or0(u_rca12_fa10_or0));
  fa fa_u_rca12_fa11_out(.a(a[11]), .b(b[11]), .cin(u_rca12_fa10_or0[0]), .fa_xor1(u_rca12_fa11_xor1), .fa_or0(u_rca12_fa11_or0));

  assign u_rca12_out[0] = u_rca12_ha_xor0[0];
  assign u_rca12_out[1] = u_rca12_fa1_xor1[0];
  assign u_rca12_out[2] = u_rca12_fa2_xor1[0];
  assign u_rca12_out[3] = u_rca12_fa3_xor1[0];
  assign u_rca12_out[4] = u_rca12_fa4_xor1[0];
  assign u_rca12_out[5] = u_rca12_fa5_xor1[0];
  assign u_rca12_out[6] = u_rca12_fa6_xor1[0];
  assign u_rca12_out[7] = u_rca12_fa7_xor1[0];
  assign u_rca12_out[8] = u_rca12_fa8_xor1[0];
  assign u_rca12_out[9] = u_rca12_fa9_xor1[0];
  assign u_rca12_out[10] = u_rca12_fa10_xor1[0];
  assign u_rca12_out[11] = u_rca12_fa11_xor1[0];
  assign u_rca12_out[12] = u_rca12_fa11_or0[0];
endmodule

module s_csamul_rca12(input [11:0] a, input [11:0] b, output [23:0] s_csamul_rca12_out);
  wire [0:0] s_csamul_rca12_and0_0;
  wire [0:0] s_csamul_rca12_and1_0;
  wire [0:0] s_csamul_rca12_and2_0;
  wire [0:0] s_csamul_rca12_and3_0;
  wire [0:0] s_csamul_rca12_and4_0;
  wire [0:0] s_csamul_rca12_and5_0;
  wire [0:0] s_csamul_rca12_and6_0;
  wire [0:0] s_csamul_rca12_and7_0;
  wire [0:0] s_csamul_rca12_and8_0;
  wire [0:0] s_csamul_rca12_and9_0;
  wire [0:0] s_csamul_rca12_and10_0;
  wire [0:0] s_csamul_rca12_nand11_0;
  wire [0:0] s_csamul_rca12_and0_1;
  wire [0:0] s_csamul_rca12_ha0_1_xor0;
  wire [0:0] s_csamul_rca12_ha0_1_and0;
  wire [0:0] s_csamul_rca12_and1_1;
  wire [0:0] s_csamul_rca12_ha1_1_xor0;
  wire [0:0] s_csamul_rca12_ha1_1_and0;
  wire [0:0] s_csamul_rca12_and2_1;
  wire [0:0] s_csamul_rca12_ha2_1_xor0;
  wire [0:0] s_csamul_rca12_ha2_1_and0;
  wire [0:0] s_csamul_rca12_and3_1;
  wire [0:0] s_csamul_rca12_ha3_1_xor0;
  wire [0:0] s_csamul_rca12_ha3_1_and0;
  wire [0:0] s_csamul_rca12_and4_1;
  wire [0:0] s_csamul_rca12_ha4_1_xor0;
  wire [0:0] s_csamul_rca12_ha4_1_and0;
  wire [0:0] s_csamul_rca12_and5_1;
  wire [0:0] s_csamul_rca12_ha5_1_xor0;
  wire [0:0] s_csamul_rca12_ha5_1_and0;
  wire [0:0] s_csamul_rca12_and6_1;
  wire [0:0] s_csamul_rca12_ha6_1_xor0;
  wire [0:0] s_csamul_rca12_ha6_1_and0;
  wire [0:0] s_csamul_rca12_and7_1;
  wire [0:0] s_csamul_rca12_ha7_1_xor0;
  wire [0:0] s_csamul_rca12_ha7_1_and0;
  wire [0:0] s_csamul_rca12_and8_1;
  wire [0:0] s_csamul_rca12_ha8_1_xor0;
  wire [0:0] s_csamul_rca12_ha8_1_and0;
  wire [0:0] s_csamul_rca12_and9_1;
  wire [0:0] s_csamul_rca12_ha9_1_xor0;
  wire [0:0] s_csamul_rca12_ha9_1_and0;
  wire [0:0] s_csamul_rca12_and10_1;
  wire [0:0] s_csamul_rca12_ha10_1_xor0;
  wire [0:0] s_csamul_rca12_ha10_1_and0;
  wire [0:0] s_csamul_rca12_nand11_1;
  wire [0:0] s_csamul_rca12_ha11_1_xor0;
  wire [0:0] s_csamul_rca12_and0_2;
  wire [0:0] s_csamul_rca12_fa0_2_xor1;
  wire [0:0] s_csamul_rca12_fa0_2_or0;
  wire [0:0] s_csamul_rca12_and1_2;
  wire [0:0] s_csamul_rca12_fa1_2_xor1;
  wire [0:0] s_csamul_rca12_fa1_2_or0;
  wire [0:0] s_csamul_rca12_and2_2;
  wire [0:0] s_csamul_rca12_fa2_2_xor1;
  wire [0:0] s_csamul_rca12_fa2_2_or0;
  wire [0:0] s_csamul_rca12_and3_2;
  wire [0:0] s_csamul_rca12_fa3_2_xor1;
  wire [0:0] s_csamul_rca12_fa3_2_or0;
  wire [0:0] s_csamul_rca12_and4_2;
  wire [0:0] s_csamul_rca12_fa4_2_xor1;
  wire [0:0] s_csamul_rca12_fa4_2_or0;
  wire [0:0] s_csamul_rca12_and5_2;
  wire [0:0] s_csamul_rca12_fa5_2_xor1;
  wire [0:0] s_csamul_rca12_fa5_2_or0;
  wire [0:0] s_csamul_rca12_and6_2;
  wire [0:0] s_csamul_rca12_fa6_2_xor1;
  wire [0:0] s_csamul_rca12_fa6_2_or0;
  wire [0:0] s_csamul_rca12_and7_2;
  wire [0:0] s_csamul_rca12_fa7_2_xor1;
  wire [0:0] s_csamul_rca12_fa7_2_or0;
  wire [0:0] s_csamul_rca12_and8_2;
  wire [0:0] s_csamul_rca12_fa8_2_xor1;
  wire [0:0] s_csamul_rca12_fa8_2_or0;
  wire [0:0] s_csamul_rca12_and9_2;
  wire [0:0] s_csamul_rca12_fa9_2_xor1;
  wire [0:0] s_csamul_rca12_fa9_2_or0;
  wire [0:0] s_csamul_rca12_and10_2;
  wire [0:0] s_csamul_rca12_fa10_2_xor1;
  wire [0:0] s_csamul_rca12_fa10_2_or0;
  wire [0:0] s_csamul_rca12_nand11_2;
  wire [0:0] s_csamul_rca12_ha11_2_xor0;
  wire [0:0] s_csamul_rca12_ha11_2_and0;
  wire [0:0] s_csamul_rca12_and0_3;
  wire [0:0] s_csamul_rca12_fa0_3_xor1;
  wire [0:0] s_csamul_rca12_fa0_3_or0;
  wire [0:0] s_csamul_rca12_and1_3;
  wire [0:0] s_csamul_rca12_fa1_3_xor1;
  wire [0:0] s_csamul_rca12_fa1_3_or0;
  wire [0:0] s_csamul_rca12_and2_3;
  wire [0:0] s_csamul_rca12_fa2_3_xor1;
  wire [0:0] s_csamul_rca12_fa2_3_or0;
  wire [0:0] s_csamul_rca12_and3_3;
  wire [0:0] s_csamul_rca12_fa3_3_xor1;
  wire [0:0] s_csamul_rca12_fa3_3_or0;
  wire [0:0] s_csamul_rca12_and4_3;
  wire [0:0] s_csamul_rca12_fa4_3_xor1;
  wire [0:0] s_csamul_rca12_fa4_3_or0;
  wire [0:0] s_csamul_rca12_and5_3;
  wire [0:0] s_csamul_rca12_fa5_3_xor1;
  wire [0:0] s_csamul_rca12_fa5_3_or0;
  wire [0:0] s_csamul_rca12_and6_3;
  wire [0:0] s_csamul_rca12_fa6_3_xor1;
  wire [0:0] s_csamul_rca12_fa6_3_or0;
  wire [0:0] s_csamul_rca12_and7_3;
  wire [0:0] s_csamul_rca12_fa7_3_xor1;
  wire [0:0] s_csamul_rca12_fa7_3_or0;
  wire [0:0] s_csamul_rca12_and8_3;
  wire [0:0] s_csamul_rca12_fa8_3_xor1;
  wire [0:0] s_csamul_rca12_fa8_3_or0;
  wire [0:0] s_csamul_rca12_and9_3;
  wire [0:0] s_csamul_rca12_fa9_3_xor1;
  wire [0:0] s_csamul_rca12_fa9_3_or0;
  wire [0:0] s_csamul_rca12_and10_3;
  wire [0:0] s_csamul_rca12_fa10_3_xor1;
  wire [0:0] s_csamul_rca12_fa10_3_or0;
  wire [0:0] s_csamul_rca12_nand11_3;
  wire [0:0] s_csamul_rca12_ha11_3_xor0;
  wire [0:0] s_csamul_rca12_ha11_3_and0;
  wire [0:0] s_csamul_rca12_and0_4;
  wire [0:0] s_csamul_rca12_fa0_4_xor1;
  wire [0:0] s_csamul_rca12_fa0_4_or0;
  wire [0:0] s_csamul_rca12_and1_4;
  wire [0:0] s_csamul_rca12_fa1_4_xor1;
  wire [0:0] s_csamul_rca12_fa1_4_or0;
  wire [0:0] s_csamul_rca12_and2_4;
  wire [0:0] s_csamul_rca12_fa2_4_xor1;
  wire [0:0] s_csamul_rca12_fa2_4_or0;
  wire [0:0] s_csamul_rca12_and3_4;
  wire [0:0] s_csamul_rca12_fa3_4_xor1;
  wire [0:0] s_csamul_rca12_fa3_4_or0;
  wire [0:0] s_csamul_rca12_and4_4;
  wire [0:0] s_csamul_rca12_fa4_4_xor1;
  wire [0:0] s_csamul_rca12_fa4_4_or0;
  wire [0:0] s_csamul_rca12_and5_4;
  wire [0:0] s_csamul_rca12_fa5_4_xor1;
  wire [0:0] s_csamul_rca12_fa5_4_or0;
  wire [0:0] s_csamul_rca12_and6_4;
  wire [0:0] s_csamul_rca12_fa6_4_xor1;
  wire [0:0] s_csamul_rca12_fa6_4_or0;
  wire [0:0] s_csamul_rca12_and7_4;
  wire [0:0] s_csamul_rca12_fa7_4_xor1;
  wire [0:0] s_csamul_rca12_fa7_4_or0;
  wire [0:0] s_csamul_rca12_and8_4;
  wire [0:0] s_csamul_rca12_fa8_4_xor1;
  wire [0:0] s_csamul_rca12_fa8_4_or0;
  wire [0:0] s_csamul_rca12_and9_4;
  wire [0:0] s_csamul_rca12_fa9_4_xor1;
  wire [0:0] s_csamul_rca12_fa9_4_or0;
  wire [0:0] s_csamul_rca12_and10_4;
  wire [0:0] s_csamul_rca12_fa10_4_xor1;
  wire [0:0] s_csamul_rca12_fa10_4_or0;
  wire [0:0] s_csamul_rca12_nand11_4;
  wire [0:0] s_csamul_rca12_ha11_4_xor0;
  wire [0:0] s_csamul_rca12_ha11_4_and0;
  wire [0:0] s_csamul_rca12_and0_5;
  wire [0:0] s_csamul_rca12_fa0_5_xor1;
  wire [0:0] s_csamul_rca12_fa0_5_or0;
  wire [0:0] s_csamul_rca12_and1_5;
  wire [0:0] s_csamul_rca12_fa1_5_xor1;
  wire [0:0] s_csamul_rca12_fa1_5_or0;
  wire [0:0] s_csamul_rca12_and2_5;
  wire [0:0] s_csamul_rca12_fa2_5_xor1;
  wire [0:0] s_csamul_rca12_fa2_5_or0;
  wire [0:0] s_csamul_rca12_and3_5;
  wire [0:0] s_csamul_rca12_fa3_5_xor1;
  wire [0:0] s_csamul_rca12_fa3_5_or0;
  wire [0:0] s_csamul_rca12_and4_5;
  wire [0:0] s_csamul_rca12_fa4_5_xor1;
  wire [0:0] s_csamul_rca12_fa4_5_or0;
  wire [0:0] s_csamul_rca12_and5_5;
  wire [0:0] s_csamul_rca12_fa5_5_xor1;
  wire [0:0] s_csamul_rca12_fa5_5_or0;
  wire [0:0] s_csamul_rca12_and6_5;
  wire [0:0] s_csamul_rca12_fa6_5_xor1;
  wire [0:0] s_csamul_rca12_fa6_5_or0;
  wire [0:0] s_csamul_rca12_and7_5;
  wire [0:0] s_csamul_rca12_fa7_5_xor1;
  wire [0:0] s_csamul_rca12_fa7_5_or0;
  wire [0:0] s_csamul_rca12_and8_5;
  wire [0:0] s_csamul_rca12_fa8_5_xor1;
  wire [0:0] s_csamul_rca12_fa8_5_or0;
  wire [0:0] s_csamul_rca12_and9_5;
  wire [0:0] s_csamul_rca12_fa9_5_xor1;
  wire [0:0] s_csamul_rca12_fa9_5_or0;
  wire [0:0] s_csamul_rca12_and10_5;
  wire [0:0] s_csamul_rca12_fa10_5_xor1;
  wire [0:0] s_csamul_rca12_fa10_5_or0;
  wire [0:0] s_csamul_rca12_nand11_5;
  wire [0:0] s_csamul_rca12_ha11_5_xor0;
  wire [0:0] s_csamul_rca12_ha11_5_and0;
  wire [0:0] s_csamul_rca12_and0_6;
  wire [0:0] s_csamul_rca12_fa0_6_xor1;
  wire [0:0] s_csamul_rca12_fa0_6_or0;
  wire [0:0] s_csamul_rca12_and1_6;
  wire [0:0] s_csamul_rca12_fa1_6_xor1;
  wire [0:0] s_csamul_rca12_fa1_6_or0;
  wire [0:0] s_csamul_rca12_and2_6;
  wire [0:0] s_csamul_rca12_fa2_6_xor1;
  wire [0:0] s_csamul_rca12_fa2_6_or0;
  wire [0:0] s_csamul_rca12_and3_6;
  wire [0:0] s_csamul_rca12_fa3_6_xor1;
  wire [0:0] s_csamul_rca12_fa3_6_or0;
  wire [0:0] s_csamul_rca12_and4_6;
  wire [0:0] s_csamul_rca12_fa4_6_xor1;
  wire [0:0] s_csamul_rca12_fa4_6_or0;
  wire [0:0] s_csamul_rca12_and5_6;
  wire [0:0] s_csamul_rca12_fa5_6_xor1;
  wire [0:0] s_csamul_rca12_fa5_6_or0;
  wire [0:0] s_csamul_rca12_and6_6;
  wire [0:0] s_csamul_rca12_fa6_6_xor1;
  wire [0:0] s_csamul_rca12_fa6_6_or0;
  wire [0:0] s_csamul_rca12_and7_6;
  wire [0:0] s_csamul_rca12_fa7_6_xor1;
  wire [0:0] s_csamul_rca12_fa7_6_or0;
  wire [0:0] s_csamul_rca12_and8_6;
  wire [0:0] s_csamul_rca12_fa8_6_xor1;
  wire [0:0] s_csamul_rca12_fa8_6_or0;
  wire [0:0] s_csamul_rca12_and9_6;
  wire [0:0] s_csamul_rca12_fa9_6_xor1;
  wire [0:0] s_csamul_rca12_fa9_6_or0;
  wire [0:0] s_csamul_rca12_and10_6;
  wire [0:0] s_csamul_rca12_fa10_6_xor1;
  wire [0:0] s_csamul_rca12_fa10_6_or0;
  wire [0:0] s_csamul_rca12_nand11_6;
  wire [0:0] s_csamul_rca12_ha11_6_xor0;
  wire [0:0] s_csamul_rca12_ha11_6_and0;
  wire [0:0] s_csamul_rca12_and0_7;
  wire [0:0] s_csamul_rca12_fa0_7_xor1;
  wire [0:0] s_csamul_rca12_fa0_7_or0;
  wire [0:0] s_csamul_rca12_and1_7;
  wire [0:0] s_csamul_rca12_fa1_7_xor1;
  wire [0:0] s_csamul_rca12_fa1_7_or0;
  wire [0:0] s_csamul_rca12_and2_7;
  wire [0:0] s_csamul_rca12_fa2_7_xor1;
  wire [0:0] s_csamul_rca12_fa2_7_or0;
  wire [0:0] s_csamul_rca12_and3_7;
  wire [0:0] s_csamul_rca12_fa3_7_xor1;
  wire [0:0] s_csamul_rca12_fa3_7_or0;
  wire [0:0] s_csamul_rca12_and4_7;
  wire [0:0] s_csamul_rca12_fa4_7_xor1;
  wire [0:0] s_csamul_rca12_fa4_7_or0;
  wire [0:0] s_csamul_rca12_and5_7;
  wire [0:0] s_csamul_rca12_fa5_7_xor1;
  wire [0:0] s_csamul_rca12_fa5_7_or0;
  wire [0:0] s_csamul_rca12_and6_7;
  wire [0:0] s_csamul_rca12_fa6_7_xor1;
  wire [0:0] s_csamul_rca12_fa6_7_or0;
  wire [0:0] s_csamul_rca12_and7_7;
  wire [0:0] s_csamul_rca12_fa7_7_xor1;
  wire [0:0] s_csamul_rca12_fa7_7_or0;
  wire [0:0] s_csamul_rca12_and8_7;
  wire [0:0] s_csamul_rca12_fa8_7_xor1;
  wire [0:0] s_csamul_rca12_fa8_7_or0;
  wire [0:0] s_csamul_rca12_and9_7;
  wire [0:0] s_csamul_rca12_fa9_7_xor1;
  wire [0:0] s_csamul_rca12_fa9_7_or0;
  wire [0:0] s_csamul_rca12_and10_7;
  wire [0:0] s_csamul_rca12_fa10_7_xor1;
  wire [0:0] s_csamul_rca12_fa10_7_or0;
  wire [0:0] s_csamul_rca12_nand11_7;
  wire [0:0] s_csamul_rca12_ha11_7_xor0;
  wire [0:0] s_csamul_rca12_ha11_7_and0;
  wire [0:0] s_csamul_rca12_and0_8;
  wire [0:0] s_csamul_rca12_fa0_8_xor1;
  wire [0:0] s_csamul_rca12_fa0_8_or0;
  wire [0:0] s_csamul_rca12_and1_8;
  wire [0:0] s_csamul_rca12_fa1_8_xor1;
  wire [0:0] s_csamul_rca12_fa1_8_or0;
  wire [0:0] s_csamul_rca12_and2_8;
  wire [0:0] s_csamul_rca12_fa2_8_xor1;
  wire [0:0] s_csamul_rca12_fa2_8_or0;
  wire [0:0] s_csamul_rca12_and3_8;
  wire [0:0] s_csamul_rca12_fa3_8_xor1;
  wire [0:0] s_csamul_rca12_fa3_8_or0;
  wire [0:0] s_csamul_rca12_and4_8;
  wire [0:0] s_csamul_rca12_fa4_8_xor1;
  wire [0:0] s_csamul_rca12_fa4_8_or0;
  wire [0:0] s_csamul_rca12_and5_8;
  wire [0:0] s_csamul_rca12_fa5_8_xor1;
  wire [0:0] s_csamul_rca12_fa5_8_or0;
  wire [0:0] s_csamul_rca12_and6_8;
  wire [0:0] s_csamul_rca12_fa6_8_xor1;
  wire [0:0] s_csamul_rca12_fa6_8_or0;
  wire [0:0] s_csamul_rca12_and7_8;
  wire [0:0] s_csamul_rca12_fa7_8_xor1;
  wire [0:0] s_csamul_rca12_fa7_8_or0;
  wire [0:0] s_csamul_rca12_and8_8;
  wire [0:0] s_csamul_rca12_fa8_8_xor1;
  wire [0:0] s_csamul_rca12_fa8_8_or0;
  wire [0:0] s_csamul_rca12_and9_8;
  wire [0:0] s_csamul_rca12_fa9_8_xor1;
  wire [0:0] s_csamul_rca12_fa9_8_or0;
  wire [0:0] s_csamul_rca12_and10_8;
  wire [0:0] s_csamul_rca12_fa10_8_xor1;
  wire [0:0] s_csamul_rca12_fa10_8_or0;
  wire [0:0] s_csamul_rca12_nand11_8;
  wire [0:0] s_csamul_rca12_ha11_8_xor0;
  wire [0:0] s_csamul_rca12_ha11_8_and0;
  wire [0:0] s_csamul_rca12_and0_9;
  wire [0:0] s_csamul_rca12_fa0_9_xor1;
  wire [0:0] s_csamul_rca12_fa0_9_or0;
  wire [0:0] s_csamul_rca12_and1_9;
  wire [0:0] s_csamul_rca12_fa1_9_xor1;
  wire [0:0] s_csamul_rca12_fa1_9_or0;
  wire [0:0] s_csamul_rca12_and2_9;
  wire [0:0] s_csamul_rca12_fa2_9_xor1;
  wire [0:0] s_csamul_rca12_fa2_9_or0;
  wire [0:0] s_csamul_rca12_and3_9;
  wire [0:0] s_csamul_rca12_fa3_9_xor1;
  wire [0:0] s_csamul_rca12_fa3_9_or0;
  wire [0:0] s_csamul_rca12_and4_9;
  wire [0:0] s_csamul_rca12_fa4_9_xor1;
  wire [0:0] s_csamul_rca12_fa4_9_or0;
  wire [0:0] s_csamul_rca12_and5_9;
  wire [0:0] s_csamul_rca12_fa5_9_xor1;
  wire [0:0] s_csamul_rca12_fa5_9_or0;
  wire [0:0] s_csamul_rca12_and6_9;
  wire [0:0] s_csamul_rca12_fa6_9_xor1;
  wire [0:0] s_csamul_rca12_fa6_9_or0;
  wire [0:0] s_csamul_rca12_and7_9;
  wire [0:0] s_csamul_rca12_fa7_9_xor1;
  wire [0:0] s_csamul_rca12_fa7_9_or0;
  wire [0:0] s_csamul_rca12_and8_9;
  wire [0:0] s_csamul_rca12_fa8_9_xor1;
  wire [0:0] s_csamul_rca12_fa8_9_or0;
  wire [0:0] s_csamul_rca12_and9_9;
  wire [0:0] s_csamul_rca12_fa9_9_xor1;
  wire [0:0] s_csamul_rca12_fa9_9_or0;
  wire [0:0] s_csamul_rca12_and10_9;
  wire [0:0] s_csamul_rca12_fa10_9_xor1;
  wire [0:0] s_csamul_rca12_fa10_9_or0;
  wire [0:0] s_csamul_rca12_nand11_9;
  wire [0:0] s_csamul_rca12_ha11_9_xor0;
  wire [0:0] s_csamul_rca12_ha11_9_and0;
  wire [0:0] s_csamul_rca12_and0_10;
  wire [0:0] s_csamul_rca12_fa0_10_xor1;
  wire [0:0] s_csamul_rca12_fa0_10_or0;
  wire [0:0] s_csamul_rca12_and1_10;
  wire [0:0] s_csamul_rca12_fa1_10_xor1;
  wire [0:0] s_csamul_rca12_fa1_10_or0;
  wire [0:0] s_csamul_rca12_and2_10;
  wire [0:0] s_csamul_rca12_fa2_10_xor1;
  wire [0:0] s_csamul_rca12_fa2_10_or0;
  wire [0:0] s_csamul_rca12_and3_10;
  wire [0:0] s_csamul_rca12_fa3_10_xor1;
  wire [0:0] s_csamul_rca12_fa3_10_or0;
  wire [0:0] s_csamul_rca12_and4_10;
  wire [0:0] s_csamul_rca12_fa4_10_xor1;
  wire [0:0] s_csamul_rca12_fa4_10_or0;
  wire [0:0] s_csamul_rca12_and5_10;
  wire [0:0] s_csamul_rca12_fa5_10_xor1;
  wire [0:0] s_csamul_rca12_fa5_10_or0;
  wire [0:0] s_csamul_rca12_and6_10;
  wire [0:0] s_csamul_rca12_fa6_10_xor1;
  wire [0:0] s_csamul_rca12_fa6_10_or0;
  wire [0:0] s_csamul_rca12_and7_10;
  wire [0:0] s_csamul_rca12_fa7_10_xor1;
  wire [0:0] s_csamul_rca12_fa7_10_or0;
  wire [0:0] s_csamul_rca12_and8_10;
  wire [0:0] s_csamul_rca12_fa8_10_xor1;
  wire [0:0] s_csamul_rca12_fa8_10_or0;
  wire [0:0] s_csamul_rca12_and9_10;
  wire [0:0] s_csamul_rca12_fa9_10_xor1;
  wire [0:0] s_csamul_rca12_fa9_10_or0;
  wire [0:0] s_csamul_rca12_and10_10;
  wire [0:0] s_csamul_rca12_fa10_10_xor1;
  wire [0:0] s_csamul_rca12_fa10_10_or0;
  wire [0:0] s_csamul_rca12_nand11_10;
  wire [0:0] s_csamul_rca12_ha11_10_xor0;
  wire [0:0] s_csamul_rca12_ha11_10_and0;
  wire [0:0] s_csamul_rca12_nand0_11;
  wire [0:0] s_csamul_rca12_fa0_11_xor1;
  wire [0:0] s_csamul_rca12_fa0_11_or0;
  wire [0:0] s_csamul_rca12_nand1_11;
  wire [0:0] s_csamul_rca12_fa1_11_xor1;
  wire [0:0] s_csamul_rca12_fa1_11_or0;
  wire [0:0] s_csamul_rca12_nand2_11;
  wire [0:0] s_csamul_rca12_fa2_11_xor1;
  wire [0:0] s_csamul_rca12_fa2_11_or0;
  wire [0:0] s_csamul_rca12_nand3_11;
  wire [0:0] s_csamul_rca12_fa3_11_xor1;
  wire [0:0] s_csamul_rca12_fa3_11_or0;
  wire [0:0] s_csamul_rca12_nand4_11;
  wire [0:0] s_csamul_rca12_fa4_11_xor1;
  wire [0:0] s_csamul_rca12_fa4_11_or0;
  wire [0:0] s_csamul_rca12_nand5_11;
  wire [0:0] s_csamul_rca12_fa5_11_xor1;
  wire [0:0] s_csamul_rca12_fa5_11_or0;
  wire [0:0] s_csamul_rca12_nand6_11;
  wire [0:0] s_csamul_rca12_fa6_11_xor1;
  wire [0:0] s_csamul_rca12_fa6_11_or0;
  wire [0:0] s_csamul_rca12_nand7_11;
  wire [0:0] s_csamul_rca12_fa7_11_xor1;
  wire [0:0] s_csamul_rca12_fa7_11_or0;
  wire [0:0] s_csamul_rca12_nand8_11;
  wire [0:0] s_csamul_rca12_fa8_11_xor1;
  wire [0:0] s_csamul_rca12_fa8_11_or0;
  wire [0:0] s_csamul_rca12_nand9_11;
  wire [0:0] s_csamul_rca12_fa9_11_xor1;
  wire [0:0] s_csamul_rca12_fa9_11_or0;
  wire [0:0] s_csamul_rca12_nand10_11;
  wire [0:0] s_csamul_rca12_fa10_11_xor1;
  wire [0:0] s_csamul_rca12_fa10_11_or0;
  wire [0:0] s_csamul_rca12_and11_11;
  wire [0:0] s_csamul_rca12_ha11_11_xor0;
  wire [0:0] s_csamul_rca12_ha11_11_and0;
  wire [11:0] s_csamul_rca12_u_rca12_a;
  wire [11:0] s_csamul_rca12_u_rca12_b;
  wire [12:0] s_csamul_rca12_u_rca12_out;

  and_gate and_gate_s_csamul_rca12_and0_0(.a(a[0]), .b(b[0]), .out(s_csamul_rca12_and0_0));
  and_gate and_gate_s_csamul_rca12_and1_0(.a(a[1]), .b(b[0]), .out(s_csamul_rca12_and1_0));
  and_gate and_gate_s_csamul_rca12_and2_0(.a(a[2]), .b(b[0]), .out(s_csamul_rca12_and2_0));
  and_gate and_gate_s_csamul_rca12_and3_0(.a(a[3]), .b(b[0]), .out(s_csamul_rca12_and3_0));
  and_gate and_gate_s_csamul_rca12_and4_0(.a(a[4]), .b(b[0]), .out(s_csamul_rca12_and4_0));
  and_gate and_gate_s_csamul_rca12_and5_0(.a(a[5]), .b(b[0]), .out(s_csamul_rca12_and5_0));
  and_gate and_gate_s_csamul_rca12_and6_0(.a(a[6]), .b(b[0]), .out(s_csamul_rca12_and6_0));
  and_gate and_gate_s_csamul_rca12_and7_0(.a(a[7]), .b(b[0]), .out(s_csamul_rca12_and7_0));
  and_gate and_gate_s_csamul_rca12_and8_0(.a(a[8]), .b(b[0]), .out(s_csamul_rca12_and8_0));
  and_gate and_gate_s_csamul_rca12_and9_0(.a(a[9]), .b(b[0]), .out(s_csamul_rca12_and9_0));
  and_gate and_gate_s_csamul_rca12_and10_0(.a(a[10]), .b(b[0]), .out(s_csamul_rca12_and10_0));
  nand_gate nand_gate_s_csamul_rca12_nand11_0(.a(a[11]), .b(b[0]), .out(s_csamul_rca12_nand11_0));
  and_gate and_gate_s_csamul_rca12_and0_1(.a(a[0]), .b(b[1]), .out(s_csamul_rca12_and0_1));
  ha ha_s_csamul_rca12_ha0_1_out(.a(s_csamul_rca12_and0_1[0]), .b(s_csamul_rca12_and1_0[0]), .ha_xor0(s_csamul_rca12_ha0_1_xor0), .ha_and0(s_csamul_rca12_ha0_1_and0));
  and_gate and_gate_s_csamul_rca12_and1_1(.a(a[1]), .b(b[1]), .out(s_csamul_rca12_and1_1));
  ha ha_s_csamul_rca12_ha1_1_out(.a(s_csamul_rca12_and1_1[0]), .b(s_csamul_rca12_and2_0[0]), .ha_xor0(s_csamul_rca12_ha1_1_xor0), .ha_and0(s_csamul_rca12_ha1_1_and0));
  and_gate and_gate_s_csamul_rca12_and2_1(.a(a[2]), .b(b[1]), .out(s_csamul_rca12_and2_1));
  ha ha_s_csamul_rca12_ha2_1_out(.a(s_csamul_rca12_and2_1[0]), .b(s_csamul_rca12_and3_0[0]), .ha_xor0(s_csamul_rca12_ha2_1_xor0), .ha_and0(s_csamul_rca12_ha2_1_and0));
  and_gate and_gate_s_csamul_rca12_and3_1(.a(a[3]), .b(b[1]), .out(s_csamul_rca12_and3_1));
  ha ha_s_csamul_rca12_ha3_1_out(.a(s_csamul_rca12_and3_1[0]), .b(s_csamul_rca12_and4_0[0]), .ha_xor0(s_csamul_rca12_ha3_1_xor0), .ha_and0(s_csamul_rca12_ha3_1_and0));
  and_gate and_gate_s_csamul_rca12_and4_1(.a(a[4]), .b(b[1]), .out(s_csamul_rca12_and4_1));
  ha ha_s_csamul_rca12_ha4_1_out(.a(s_csamul_rca12_and4_1[0]), .b(s_csamul_rca12_and5_0[0]), .ha_xor0(s_csamul_rca12_ha4_1_xor0), .ha_and0(s_csamul_rca12_ha4_1_and0));
  and_gate and_gate_s_csamul_rca12_and5_1(.a(a[5]), .b(b[1]), .out(s_csamul_rca12_and5_1));
  ha ha_s_csamul_rca12_ha5_1_out(.a(s_csamul_rca12_and5_1[0]), .b(s_csamul_rca12_and6_0[0]), .ha_xor0(s_csamul_rca12_ha5_1_xor0), .ha_and0(s_csamul_rca12_ha5_1_and0));
  and_gate and_gate_s_csamul_rca12_and6_1(.a(a[6]), .b(b[1]), .out(s_csamul_rca12_and6_1));
  ha ha_s_csamul_rca12_ha6_1_out(.a(s_csamul_rca12_and6_1[0]), .b(s_csamul_rca12_and7_0[0]), .ha_xor0(s_csamul_rca12_ha6_1_xor0), .ha_and0(s_csamul_rca12_ha6_1_and0));
  and_gate and_gate_s_csamul_rca12_and7_1(.a(a[7]), .b(b[1]), .out(s_csamul_rca12_and7_1));
  ha ha_s_csamul_rca12_ha7_1_out(.a(s_csamul_rca12_and7_1[0]), .b(s_csamul_rca12_and8_0[0]), .ha_xor0(s_csamul_rca12_ha7_1_xor0), .ha_and0(s_csamul_rca12_ha7_1_and0));
  and_gate and_gate_s_csamul_rca12_and8_1(.a(a[8]), .b(b[1]), .out(s_csamul_rca12_and8_1));
  ha ha_s_csamul_rca12_ha8_1_out(.a(s_csamul_rca12_and8_1[0]), .b(s_csamul_rca12_and9_0[0]), .ha_xor0(s_csamul_rca12_ha8_1_xor0), .ha_and0(s_csamul_rca12_ha8_1_and0));
  and_gate and_gate_s_csamul_rca12_and9_1(.a(a[9]), .b(b[1]), .out(s_csamul_rca12_and9_1));
  ha ha_s_csamul_rca12_ha9_1_out(.a(s_csamul_rca12_and9_1[0]), .b(s_csamul_rca12_and10_0[0]), .ha_xor0(s_csamul_rca12_ha9_1_xor0), .ha_and0(s_csamul_rca12_ha9_1_and0));
  and_gate and_gate_s_csamul_rca12_and10_1(.a(a[10]), .b(b[1]), .out(s_csamul_rca12_and10_1));
  ha ha_s_csamul_rca12_ha10_1_out(.a(s_csamul_rca12_and10_1[0]), .b(s_csamul_rca12_nand11_0[0]), .ha_xor0(s_csamul_rca12_ha10_1_xor0), .ha_and0(s_csamul_rca12_ha10_1_and0));
  nand_gate nand_gate_s_csamul_rca12_nand11_1(.a(a[11]), .b(b[1]), .out(s_csamul_rca12_nand11_1));
  ha ha_s_csamul_rca12_ha11_1_out(.a(s_csamul_rca12_nand11_1[0]), .b(1'b1), .ha_xor0(s_csamul_rca12_ha11_1_xor0), .ha_and0(s_csamul_rca12_nand11_1));
  and_gate and_gate_s_csamul_rca12_and0_2(.a(a[0]), .b(b[2]), .out(s_csamul_rca12_and0_2));
  fa fa_s_csamul_rca12_fa0_2_out(.a(s_csamul_rca12_and0_2[0]), .b(s_csamul_rca12_ha1_1_xor0[0]), .cin(s_csamul_rca12_ha0_1_and0[0]), .fa_xor1(s_csamul_rca12_fa0_2_xor1), .fa_or0(s_csamul_rca12_fa0_2_or0));
  and_gate and_gate_s_csamul_rca12_and1_2(.a(a[1]), .b(b[2]), .out(s_csamul_rca12_and1_2));
  fa fa_s_csamul_rca12_fa1_2_out(.a(s_csamul_rca12_and1_2[0]), .b(s_csamul_rca12_ha2_1_xor0[0]), .cin(s_csamul_rca12_ha1_1_and0[0]), .fa_xor1(s_csamul_rca12_fa1_2_xor1), .fa_or0(s_csamul_rca12_fa1_2_or0));
  and_gate and_gate_s_csamul_rca12_and2_2(.a(a[2]), .b(b[2]), .out(s_csamul_rca12_and2_2));
  fa fa_s_csamul_rca12_fa2_2_out(.a(s_csamul_rca12_and2_2[0]), .b(s_csamul_rca12_ha3_1_xor0[0]), .cin(s_csamul_rca12_ha2_1_and0[0]), .fa_xor1(s_csamul_rca12_fa2_2_xor1), .fa_or0(s_csamul_rca12_fa2_2_or0));
  and_gate and_gate_s_csamul_rca12_and3_2(.a(a[3]), .b(b[2]), .out(s_csamul_rca12_and3_2));
  fa fa_s_csamul_rca12_fa3_2_out(.a(s_csamul_rca12_and3_2[0]), .b(s_csamul_rca12_ha4_1_xor0[0]), .cin(s_csamul_rca12_ha3_1_and0[0]), .fa_xor1(s_csamul_rca12_fa3_2_xor1), .fa_or0(s_csamul_rca12_fa3_2_or0));
  and_gate and_gate_s_csamul_rca12_and4_2(.a(a[4]), .b(b[2]), .out(s_csamul_rca12_and4_2));
  fa fa_s_csamul_rca12_fa4_2_out(.a(s_csamul_rca12_and4_2[0]), .b(s_csamul_rca12_ha5_1_xor0[0]), .cin(s_csamul_rca12_ha4_1_and0[0]), .fa_xor1(s_csamul_rca12_fa4_2_xor1), .fa_or0(s_csamul_rca12_fa4_2_or0));
  and_gate and_gate_s_csamul_rca12_and5_2(.a(a[5]), .b(b[2]), .out(s_csamul_rca12_and5_2));
  fa fa_s_csamul_rca12_fa5_2_out(.a(s_csamul_rca12_and5_2[0]), .b(s_csamul_rca12_ha6_1_xor0[0]), .cin(s_csamul_rca12_ha5_1_and0[0]), .fa_xor1(s_csamul_rca12_fa5_2_xor1), .fa_or0(s_csamul_rca12_fa5_2_or0));
  and_gate and_gate_s_csamul_rca12_and6_2(.a(a[6]), .b(b[2]), .out(s_csamul_rca12_and6_2));
  fa fa_s_csamul_rca12_fa6_2_out(.a(s_csamul_rca12_and6_2[0]), .b(s_csamul_rca12_ha7_1_xor0[0]), .cin(s_csamul_rca12_ha6_1_and0[0]), .fa_xor1(s_csamul_rca12_fa6_2_xor1), .fa_or0(s_csamul_rca12_fa6_2_or0));
  and_gate and_gate_s_csamul_rca12_and7_2(.a(a[7]), .b(b[2]), .out(s_csamul_rca12_and7_2));
  fa fa_s_csamul_rca12_fa7_2_out(.a(s_csamul_rca12_and7_2[0]), .b(s_csamul_rca12_ha8_1_xor0[0]), .cin(s_csamul_rca12_ha7_1_and0[0]), .fa_xor1(s_csamul_rca12_fa7_2_xor1), .fa_or0(s_csamul_rca12_fa7_2_or0));
  and_gate and_gate_s_csamul_rca12_and8_2(.a(a[8]), .b(b[2]), .out(s_csamul_rca12_and8_2));
  fa fa_s_csamul_rca12_fa8_2_out(.a(s_csamul_rca12_and8_2[0]), .b(s_csamul_rca12_ha9_1_xor0[0]), .cin(s_csamul_rca12_ha8_1_and0[0]), .fa_xor1(s_csamul_rca12_fa8_2_xor1), .fa_or0(s_csamul_rca12_fa8_2_or0));
  and_gate and_gate_s_csamul_rca12_and9_2(.a(a[9]), .b(b[2]), .out(s_csamul_rca12_and9_2));
  fa fa_s_csamul_rca12_fa9_2_out(.a(s_csamul_rca12_and9_2[0]), .b(s_csamul_rca12_ha10_1_xor0[0]), .cin(s_csamul_rca12_ha9_1_and0[0]), .fa_xor1(s_csamul_rca12_fa9_2_xor1), .fa_or0(s_csamul_rca12_fa9_2_or0));
  and_gate and_gate_s_csamul_rca12_and10_2(.a(a[10]), .b(b[2]), .out(s_csamul_rca12_and10_2));
  fa fa_s_csamul_rca12_fa10_2_out(.a(s_csamul_rca12_and10_2[0]), .b(s_csamul_rca12_ha11_1_xor0[0]), .cin(s_csamul_rca12_ha10_1_and0[0]), .fa_xor1(s_csamul_rca12_fa10_2_xor1), .fa_or0(s_csamul_rca12_fa10_2_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_2(.a(a[11]), .b(b[2]), .out(s_csamul_rca12_nand11_2));
  ha ha_s_csamul_rca12_ha11_2_out(.a(s_csamul_rca12_nand11_2[0]), .b(s_csamul_rca12_nand11_1[0]), .ha_xor0(s_csamul_rca12_ha11_2_xor0), .ha_and0(s_csamul_rca12_ha11_2_and0));
  and_gate and_gate_s_csamul_rca12_and0_3(.a(a[0]), .b(b[3]), .out(s_csamul_rca12_and0_3));
  fa fa_s_csamul_rca12_fa0_3_out(.a(s_csamul_rca12_and0_3[0]), .b(s_csamul_rca12_fa1_2_xor1[0]), .cin(s_csamul_rca12_fa0_2_or0[0]), .fa_xor1(s_csamul_rca12_fa0_3_xor1), .fa_or0(s_csamul_rca12_fa0_3_or0));
  and_gate and_gate_s_csamul_rca12_and1_3(.a(a[1]), .b(b[3]), .out(s_csamul_rca12_and1_3));
  fa fa_s_csamul_rca12_fa1_3_out(.a(s_csamul_rca12_and1_3[0]), .b(s_csamul_rca12_fa2_2_xor1[0]), .cin(s_csamul_rca12_fa1_2_or0[0]), .fa_xor1(s_csamul_rca12_fa1_3_xor1), .fa_or0(s_csamul_rca12_fa1_3_or0));
  and_gate and_gate_s_csamul_rca12_and2_3(.a(a[2]), .b(b[3]), .out(s_csamul_rca12_and2_3));
  fa fa_s_csamul_rca12_fa2_3_out(.a(s_csamul_rca12_and2_3[0]), .b(s_csamul_rca12_fa3_2_xor1[0]), .cin(s_csamul_rca12_fa2_2_or0[0]), .fa_xor1(s_csamul_rca12_fa2_3_xor1), .fa_or0(s_csamul_rca12_fa2_3_or0));
  and_gate and_gate_s_csamul_rca12_and3_3(.a(a[3]), .b(b[3]), .out(s_csamul_rca12_and3_3));
  fa fa_s_csamul_rca12_fa3_3_out(.a(s_csamul_rca12_and3_3[0]), .b(s_csamul_rca12_fa4_2_xor1[0]), .cin(s_csamul_rca12_fa3_2_or0[0]), .fa_xor1(s_csamul_rca12_fa3_3_xor1), .fa_or0(s_csamul_rca12_fa3_3_or0));
  and_gate and_gate_s_csamul_rca12_and4_3(.a(a[4]), .b(b[3]), .out(s_csamul_rca12_and4_3));
  fa fa_s_csamul_rca12_fa4_3_out(.a(s_csamul_rca12_and4_3[0]), .b(s_csamul_rca12_fa5_2_xor1[0]), .cin(s_csamul_rca12_fa4_2_or0[0]), .fa_xor1(s_csamul_rca12_fa4_3_xor1), .fa_or0(s_csamul_rca12_fa4_3_or0));
  and_gate and_gate_s_csamul_rca12_and5_3(.a(a[5]), .b(b[3]), .out(s_csamul_rca12_and5_3));
  fa fa_s_csamul_rca12_fa5_3_out(.a(s_csamul_rca12_and5_3[0]), .b(s_csamul_rca12_fa6_2_xor1[0]), .cin(s_csamul_rca12_fa5_2_or0[0]), .fa_xor1(s_csamul_rca12_fa5_3_xor1), .fa_or0(s_csamul_rca12_fa5_3_or0));
  and_gate and_gate_s_csamul_rca12_and6_3(.a(a[6]), .b(b[3]), .out(s_csamul_rca12_and6_3));
  fa fa_s_csamul_rca12_fa6_3_out(.a(s_csamul_rca12_and6_3[0]), .b(s_csamul_rca12_fa7_2_xor1[0]), .cin(s_csamul_rca12_fa6_2_or0[0]), .fa_xor1(s_csamul_rca12_fa6_3_xor1), .fa_or0(s_csamul_rca12_fa6_3_or0));
  and_gate and_gate_s_csamul_rca12_and7_3(.a(a[7]), .b(b[3]), .out(s_csamul_rca12_and7_3));
  fa fa_s_csamul_rca12_fa7_3_out(.a(s_csamul_rca12_and7_3[0]), .b(s_csamul_rca12_fa8_2_xor1[0]), .cin(s_csamul_rca12_fa7_2_or0[0]), .fa_xor1(s_csamul_rca12_fa7_3_xor1), .fa_or0(s_csamul_rca12_fa7_3_or0));
  and_gate and_gate_s_csamul_rca12_and8_3(.a(a[8]), .b(b[3]), .out(s_csamul_rca12_and8_3));
  fa fa_s_csamul_rca12_fa8_3_out(.a(s_csamul_rca12_and8_3[0]), .b(s_csamul_rca12_fa9_2_xor1[0]), .cin(s_csamul_rca12_fa8_2_or0[0]), .fa_xor1(s_csamul_rca12_fa8_3_xor1), .fa_or0(s_csamul_rca12_fa8_3_or0));
  and_gate and_gate_s_csamul_rca12_and9_3(.a(a[9]), .b(b[3]), .out(s_csamul_rca12_and9_3));
  fa fa_s_csamul_rca12_fa9_3_out(.a(s_csamul_rca12_and9_3[0]), .b(s_csamul_rca12_fa10_2_xor1[0]), .cin(s_csamul_rca12_fa9_2_or0[0]), .fa_xor1(s_csamul_rca12_fa9_3_xor1), .fa_or0(s_csamul_rca12_fa9_3_or0));
  and_gate and_gate_s_csamul_rca12_and10_3(.a(a[10]), .b(b[3]), .out(s_csamul_rca12_and10_3));
  fa fa_s_csamul_rca12_fa10_3_out(.a(s_csamul_rca12_and10_3[0]), .b(s_csamul_rca12_ha11_2_xor0[0]), .cin(s_csamul_rca12_fa10_2_or0[0]), .fa_xor1(s_csamul_rca12_fa10_3_xor1), .fa_or0(s_csamul_rca12_fa10_3_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_3(.a(a[11]), .b(b[3]), .out(s_csamul_rca12_nand11_3));
  ha ha_s_csamul_rca12_ha11_3_out(.a(s_csamul_rca12_nand11_3[0]), .b(s_csamul_rca12_ha11_2_and0[0]), .ha_xor0(s_csamul_rca12_ha11_3_xor0), .ha_and0(s_csamul_rca12_ha11_3_and0));
  and_gate and_gate_s_csamul_rca12_and0_4(.a(a[0]), .b(b[4]), .out(s_csamul_rca12_and0_4));
  fa fa_s_csamul_rca12_fa0_4_out(.a(s_csamul_rca12_and0_4[0]), .b(s_csamul_rca12_fa1_3_xor1[0]), .cin(s_csamul_rca12_fa0_3_or0[0]), .fa_xor1(s_csamul_rca12_fa0_4_xor1), .fa_or0(s_csamul_rca12_fa0_4_or0));
  and_gate and_gate_s_csamul_rca12_and1_4(.a(a[1]), .b(b[4]), .out(s_csamul_rca12_and1_4));
  fa fa_s_csamul_rca12_fa1_4_out(.a(s_csamul_rca12_and1_4[0]), .b(s_csamul_rca12_fa2_3_xor1[0]), .cin(s_csamul_rca12_fa1_3_or0[0]), .fa_xor1(s_csamul_rca12_fa1_4_xor1), .fa_or0(s_csamul_rca12_fa1_4_or0));
  and_gate and_gate_s_csamul_rca12_and2_4(.a(a[2]), .b(b[4]), .out(s_csamul_rca12_and2_4));
  fa fa_s_csamul_rca12_fa2_4_out(.a(s_csamul_rca12_and2_4[0]), .b(s_csamul_rca12_fa3_3_xor1[0]), .cin(s_csamul_rca12_fa2_3_or0[0]), .fa_xor1(s_csamul_rca12_fa2_4_xor1), .fa_or0(s_csamul_rca12_fa2_4_or0));
  and_gate and_gate_s_csamul_rca12_and3_4(.a(a[3]), .b(b[4]), .out(s_csamul_rca12_and3_4));
  fa fa_s_csamul_rca12_fa3_4_out(.a(s_csamul_rca12_and3_4[0]), .b(s_csamul_rca12_fa4_3_xor1[0]), .cin(s_csamul_rca12_fa3_3_or0[0]), .fa_xor1(s_csamul_rca12_fa3_4_xor1), .fa_or0(s_csamul_rca12_fa3_4_or0));
  and_gate and_gate_s_csamul_rca12_and4_4(.a(a[4]), .b(b[4]), .out(s_csamul_rca12_and4_4));
  fa fa_s_csamul_rca12_fa4_4_out(.a(s_csamul_rca12_and4_4[0]), .b(s_csamul_rca12_fa5_3_xor1[0]), .cin(s_csamul_rca12_fa4_3_or0[0]), .fa_xor1(s_csamul_rca12_fa4_4_xor1), .fa_or0(s_csamul_rca12_fa4_4_or0));
  and_gate and_gate_s_csamul_rca12_and5_4(.a(a[5]), .b(b[4]), .out(s_csamul_rca12_and5_4));
  fa fa_s_csamul_rca12_fa5_4_out(.a(s_csamul_rca12_and5_4[0]), .b(s_csamul_rca12_fa6_3_xor1[0]), .cin(s_csamul_rca12_fa5_3_or0[0]), .fa_xor1(s_csamul_rca12_fa5_4_xor1), .fa_or0(s_csamul_rca12_fa5_4_or0));
  and_gate and_gate_s_csamul_rca12_and6_4(.a(a[6]), .b(b[4]), .out(s_csamul_rca12_and6_4));
  fa fa_s_csamul_rca12_fa6_4_out(.a(s_csamul_rca12_and6_4[0]), .b(s_csamul_rca12_fa7_3_xor1[0]), .cin(s_csamul_rca12_fa6_3_or0[0]), .fa_xor1(s_csamul_rca12_fa6_4_xor1), .fa_or0(s_csamul_rca12_fa6_4_or0));
  and_gate and_gate_s_csamul_rca12_and7_4(.a(a[7]), .b(b[4]), .out(s_csamul_rca12_and7_4));
  fa fa_s_csamul_rca12_fa7_4_out(.a(s_csamul_rca12_and7_4[0]), .b(s_csamul_rca12_fa8_3_xor1[0]), .cin(s_csamul_rca12_fa7_3_or0[0]), .fa_xor1(s_csamul_rca12_fa7_4_xor1), .fa_or0(s_csamul_rca12_fa7_4_or0));
  and_gate and_gate_s_csamul_rca12_and8_4(.a(a[8]), .b(b[4]), .out(s_csamul_rca12_and8_4));
  fa fa_s_csamul_rca12_fa8_4_out(.a(s_csamul_rca12_and8_4[0]), .b(s_csamul_rca12_fa9_3_xor1[0]), .cin(s_csamul_rca12_fa8_3_or0[0]), .fa_xor1(s_csamul_rca12_fa8_4_xor1), .fa_or0(s_csamul_rca12_fa8_4_or0));
  and_gate and_gate_s_csamul_rca12_and9_4(.a(a[9]), .b(b[4]), .out(s_csamul_rca12_and9_4));
  fa fa_s_csamul_rca12_fa9_4_out(.a(s_csamul_rca12_and9_4[0]), .b(s_csamul_rca12_fa10_3_xor1[0]), .cin(s_csamul_rca12_fa9_3_or0[0]), .fa_xor1(s_csamul_rca12_fa9_4_xor1), .fa_or0(s_csamul_rca12_fa9_4_or0));
  and_gate and_gate_s_csamul_rca12_and10_4(.a(a[10]), .b(b[4]), .out(s_csamul_rca12_and10_4));
  fa fa_s_csamul_rca12_fa10_4_out(.a(s_csamul_rca12_and10_4[0]), .b(s_csamul_rca12_ha11_3_xor0[0]), .cin(s_csamul_rca12_fa10_3_or0[0]), .fa_xor1(s_csamul_rca12_fa10_4_xor1), .fa_or0(s_csamul_rca12_fa10_4_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_4(.a(a[11]), .b(b[4]), .out(s_csamul_rca12_nand11_4));
  ha ha_s_csamul_rca12_ha11_4_out(.a(s_csamul_rca12_nand11_4[0]), .b(s_csamul_rca12_ha11_3_and0[0]), .ha_xor0(s_csamul_rca12_ha11_4_xor0), .ha_and0(s_csamul_rca12_ha11_4_and0));
  and_gate and_gate_s_csamul_rca12_and0_5(.a(a[0]), .b(b[5]), .out(s_csamul_rca12_and0_5));
  fa fa_s_csamul_rca12_fa0_5_out(.a(s_csamul_rca12_and0_5[0]), .b(s_csamul_rca12_fa1_4_xor1[0]), .cin(s_csamul_rca12_fa0_4_or0[0]), .fa_xor1(s_csamul_rca12_fa0_5_xor1), .fa_or0(s_csamul_rca12_fa0_5_or0));
  and_gate and_gate_s_csamul_rca12_and1_5(.a(a[1]), .b(b[5]), .out(s_csamul_rca12_and1_5));
  fa fa_s_csamul_rca12_fa1_5_out(.a(s_csamul_rca12_and1_5[0]), .b(s_csamul_rca12_fa2_4_xor1[0]), .cin(s_csamul_rca12_fa1_4_or0[0]), .fa_xor1(s_csamul_rca12_fa1_5_xor1), .fa_or0(s_csamul_rca12_fa1_5_or0));
  and_gate and_gate_s_csamul_rca12_and2_5(.a(a[2]), .b(b[5]), .out(s_csamul_rca12_and2_5));
  fa fa_s_csamul_rca12_fa2_5_out(.a(s_csamul_rca12_and2_5[0]), .b(s_csamul_rca12_fa3_4_xor1[0]), .cin(s_csamul_rca12_fa2_4_or0[0]), .fa_xor1(s_csamul_rca12_fa2_5_xor1), .fa_or0(s_csamul_rca12_fa2_5_or0));
  and_gate and_gate_s_csamul_rca12_and3_5(.a(a[3]), .b(b[5]), .out(s_csamul_rca12_and3_5));
  fa fa_s_csamul_rca12_fa3_5_out(.a(s_csamul_rca12_and3_5[0]), .b(s_csamul_rca12_fa4_4_xor1[0]), .cin(s_csamul_rca12_fa3_4_or0[0]), .fa_xor1(s_csamul_rca12_fa3_5_xor1), .fa_or0(s_csamul_rca12_fa3_5_or0));
  and_gate and_gate_s_csamul_rca12_and4_5(.a(a[4]), .b(b[5]), .out(s_csamul_rca12_and4_5));
  fa fa_s_csamul_rca12_fa4_5_out(.a(s_csamul_rca12_and4_5[0]), .b(s_csamul_rca12_fa5_4_xor1[0]), .cin(s_csamul_rca12_fa4_4_or0[0]), .fa_xor1(s_csamul_rca12_fa4_5_xor1), .fa_or0(s_csamul_rca12_fa4_5_or0));
  and_gate and_gate_s_csamul_rca12_and5_5(.a(a[5]), .b(b[5]), .out(s_csamul_rca12_and5_5));
  fa fa_s_csamul_rca12_fa5_5_out(.a(s_csamul_rca12_and5_5[0]), .b(s_csamul_rca12_fa6_4_xor1[0]), .cin(s_csamul_rca12_fa5_4_or0[0]), .fa_xor1(s_csamul_rca12_fa5_5_xor1), .fa_or0(s_csamul_rca12_fa5_5_or0));
  and_gate and_gate_s_csamul_rca12_and6_5(.a(a[6]), .b(b[5]), .out(s_csamul_rca12_and6_5));
  fa fa_s_csamul_rca12_fa6_5_out(.a(s_csamul_rca12_and6_5[0]), .b(s_csamul_rca12_fa7_4_xor1[0]), .cin(s_csamul_rca12_fa6_4_or0[0]), .fa_xor1(s_csamul_rca12_fa6_5_xor1), .fa_or0(s_csamul_rca12_fa6_5_or0));
  and_gate and_gate_s_csamul_rca12_and7_5(.a(a[7]), .b(b[5]), .out(s_csamul_rca12_and7_5));
  fa fa_s_csamul_rca12_fa7_5_out(.a(s_csamul_rca12_and7_5[0]), .b(s_csamul_rca12_fa8_4_xor1[0]), .cin(s_csamul_rca12_fa7_4_or0[0]), .fa_xor1(s_csamul_rca12_fa7_5_xor1), .fa_or0(s_csamul_rca12_fa7_5_or0));
  and_gate and_gate_s_csamul_rca12_and8_5(.a(a[8]), .b(b[5]), .out(s_csamul_rca12_and8_5));
  fa fa_s_csamul_rca12_fa8_5_out(.a(s_csamul_rca12_and8_5[0]), .b(s_csamul_rca12_fa9_4_xor1[0]), .cin(s_csamul_rca12_fa8_4_or0[0]), .fa_xor1(s_csamul_rca12_fa8_5_xor1), .fa_or0(s_csamul_rca12_fa8_5_or0));
  and_gate and_gate_s_csamul_rca12_and9_5(.a(a[9]), .b(b[5]), .out(s_csamul_rca12_and9_5));
  fa fa_s_csamul_rca12_fa9_5_out(.a(s_csamul_rca12_and9_5[0]), .b(s_csamul_rca12_fa10_4_xor1[0]), .cin(s_csamul_rca12_fa9_4_or0[0]), .fa_xor1(s_csamul_rca12_fa9_5_xor1), .fa_or0(s_csamul_rca12_fa9_5_or0));
  and_gate and_gate_s_csamul_rca12_and10_5(.a(a[10]), .b(b[5]), .out(s_csamul_rca12_and10_5));
  fa fa_s_csamul_rca12_fa10_5_out(.a(s_csamul_rca12_and10_5[0]), .b(s_csamul_rca12_ha11_4_xor0[0]), .cin(s_csamul_rca12_fa10_4_or0[0]), .fa_xor1(s_csamul_rca12_fa10_5_xor1), .fa_or0(s_csamul_rca12_fa10_5_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_5(.a(a[11]), .b(b[5]), .out(s_csamul_rca12_nand11_5));
  ha ha_s_csamul_rca12_ha11_5_out(.a(s_csamul_rca12_nand11_5[0]), .b(s_csamul_rca12_ha11_4_and0[0]), .ha_xor0(s_csamul_rca12_ha11_5_xor0), .ha_and0(s_csamul_rca12_ha11_5_and0));
  and_gate and_gate_s_csamul_rca12_and0_6(.a(a[0]), .b(b[6]), .out(s_csamul_rca12_and0_6));
  fa fa_s_csamul_rca12_fa0_6_out(.a(s_csamul_rca12_and0_6[0]), .b(s_csamul_rca12_fa1_5_xor1[0]), .cin(s_csamul_rca12_fa0_5_or0[0]), .fa_xor1(s_csamul_rca12_fa0_6_xor1), .fa_or0(s_csamul_rca12_fa0_6_or0));
  and_gate and_gate_s_csamul_rca12_and1_6(.a(a[1]), .b(b[6]), .out(s_csamul_rca12_and1_6));
  fa fa_s_csamul_rca12_fa1_6_out(.a(s_csamul_rca12_and1_6[0]), .b(s_csamul_rca12_fa2_5_xor1[0]), .cin(s_csamul_rca12_fa1_5_or0[0]), .fa_xor1(s_csamul_rca12_fa1_6_xor1), .fa_or0(s_csamul_rca12_fa1_6_or0));
  and_gate and_gate_s_csamul_rca12_and2_6(.a(a[2]), .b(b[6]), .out(s_csamul_rca12_and2_6));
  fa fa_s_csamul_rca12_fa2_6_out(.a(s_csamul_rca12_and2_6[0]), .b(s_csamul_rca12_fa3_5_xor1[0]), .cin(s_csamul_rca12_fa2_5_or0[0]), .fa_xor1(s_csamul_rca12_fa2_6_xor1), .fa_or0(s_csamul_rca12_fa2_6_or0));
  and_gate and_gate_s_csamul_rca12_and3_6(.a(a[3]), .b(b[6]), .out(s_csamul_rca12_and3_6));
  fa fa_s_csamul_rca12_fa3_6_out(.a(s_csamul_rca12_and3_6[0]), .b(s_csamul_rca12_fa4_5_xor1[0]), .cin(s_csamul_rca12_fa3_5_or0[0]), .fa_xor1(s_csamul_rca12_fa3_6_xor1), .fa_or0(s_csamul_rca12_fa3_6_or0));
  and_gate and_gate_s_csamul_rca12_and4_6(.a(a[4]), .b(b[6]), .out(s_csamul_rca12_and4_6));
  fa fa_s_csamul_rca12_fa4_6_out(.a(s_csamul_rca12_and4_6[0]), .b(s_csamul_rca12_fa5_5_xor1[0]), .cin(s_csamul_rca12_fa4_5_or0[0]), .fa_xor1(s_csamul_rca12_fa4_6_xor1), .fa_or0(s_csamul_rca12_fa4_6_or0));
  and_gate and_gate_s_csamul_rca12_and5_6(.a(a[5]), .b(b[6]), .out(s_csamul_rca12_and5_6));
  fa fa_s_csamul_rca12_fa5_6_out(.a(s_csamul_rca12_and5_6[0]), .b(s_csamul_rca12_fa6_5_xor1[0]), .cin(s_csamul_rca12_fa5_5_or0[0]), .fa_xor1(s_csamul_rca12_fa5_6_xor1), .fa_or0(s_csamul_rca12_fa5_6_or0));
  and_gate and_gate_s_csamul_rca12_and6_6(.a(a[6]), .b(b[6]), .out(s_csamul_rca12_and6_6));
  fa fa_s_csamul_rca12_fa6_6_out(.a(s_csamul_rca12_and6_6[0]), .b(s_csamul_rca12_fa7_5_xor1[0]), .cin(s_csamul_rca12_fa6_5_or0[0]), .fa_xor1(s_csamul_rca12_fa6_6_xor1), .fa_or0(s_csamul_rca12_fa6_6_or0));
  and_gate and_gate_s_csamul_rca12_and7_6(.a(a[7]), .b(b[6]), .out(s_csamul_rca12_and7_6));
  fa fa_s_csamul_rca12_fa7_6_out(.a(s_csamul_rca12_and7_6[0]), .b(s_csamul_rca12_fa8_5_xor1[0]), .cin(s_csamul_rca12_fa7_5_or0[0]), .fa_xor1(s_csamul_rca12_fa7_6_xor1), .fa_or0(s_csamul_rca12_fa7_6_or0));
  and_gate and_gate_s_csamul_rca12_and8_6(.a(a[8]), .b(b[6]), .out(s_csamul_rca12_and8_6));
  fa fa_s_csamul_rca12_fa8_6_out(.a(s_csamul_rca12_and8_6[0]), .b(s_csamul_rca12_fa9_5_xor1[0]), .cin(s_csamul_rca12_fa8_5_or0[0]), .fa_xor1(s_csamul_rca12_fa8_6_xor1), .fa_or0(s_csamul_rca12_fa8_6_or0));
  and_gate and_gate_s_csamul_rca12_and9_6(.a(a[9]), .b(b[6]), .out(s_csamul_rca12_and9_6));
  fa fa_s_csamul_rca12_fa9_6_out(.a(s_csamul_rca12_and9_6[0]), .b(s_csamul_rca12_fa10_5_xor1[0]), .cin(s_csamul_rca12_fa9_5_or0[0]), .fa_xor1(s_csamul_rca12_fa9_6_xor1), .fa_or0(s_csamul_rca12_fa9_6_or0));
  and_gate and_gate_s_csamul_rca12_and10_6(.a(a[10]), .b(b[6]), .out(s_csamul_rca12_and10_6));
  fa fa_s_csamul_rca12_fa10_6_out(.a(s_csamul_rca12_and10_6[0]), .b(s_csamul_rca12_ha11_5_xor0[0]), .cin(s_csamul_rca12_fa10_5_or0[0]), .fa_xor1(s_csamul_rca12_fa10_6_xor1), .fa_or0(s_csamul_rca12_fa10_6_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_6(.a(a[11]), .b(b[6]), .out(s_csamul_rca12_nand11_6));
  ha ha_s_csamul_rca12_ha11_6_out(.a(s_csamul_rca12_nand11_6[0]), .b(s_csamul_rca12_ha11_5_and0[0]), .ha_xor0(s_csamul_rca12_ha11_6_xor0), .ha_and0(s_csamul_rca12_ha11_6_and0));
  and_gate and_gate_s_csamul_rca12_and0_7(.a(a[0]), .b(b[7]), .out(s_csamul_rca12_and0_7));
  fa fa_s_csamul_rca12_fa0_7_out(.a(s_csamul_rca12_and0_7[0]), .b(s_csamul_rca12_fa1_6_xor1[0]), .cin(s_csamul_rca12_fa0_6_or0[0]), .fa_xor1(s_csamul_rca12_fa0_7_xor1), .fa_or0(s_csamul_rca12_fa0_7_or0));
  and_gate and_gate_s_csamul_rca12_and1_7(.a(a[1]), .b(b[7]), .out(s_csamul_rca12_and1_7));
  fa fa_s_csamul_rca12_fa1_7_out(.a(s_csamul_rca12_and1_7[0]), .b(s_csamul_rca12_fa2_6_xor1[0]), .cin(s_csamul_rca12_fa1_6_or0[0]), .fa_xor1(s_csamul_rca12_fa1_7_xor1), .fa_or0(s_csamul_rca12_fa1_7_or0));
  and_gate and_gate_s_csamul_rca12_and2_7(.a(a[2]), .b(b[7]), .out(s_csamul_rca12_and2_7));
  fa fa_s_csamul_rca12_fa2_7_out(.a(s_csamul_rca12_and2_7[0]), .b(s_csamul_rca12_fa3_6_xor1[0]), .cin(s_csamul_rca12_fa2_6_or0[0]), .fa_xor1(s_csamul_rca12_fa2_7_xor1), .fa_or0(s_csamul_rca12_fa2_7_or0));
  and_gate and_gate_s_csamul_rca12_and3_7(.a(a[3]), .b(b[7]), .out(s_csamul_rca12_and3_7));
  fa fa_s_csamul_rca12_fa3_7_out(.a(s_csamul_rca12_and3_7[0]), .b(s_csamul_rca12_fa4_6_xor1[0]), .cin(s_csamul_rca12_fa3_6_or0[0]), .fa_xor1(s_csamul_rca12_fa3_7_xor1), .fa_or0(s_csamul_rca12_fa3_7_or0));
  and_gate and_gate_s_csamul_rca12_and4_7(.a(a[4]), .b(b[7]), .out(s_csamul_rca12_and4_7));
  fa fa_s_csamul_rca12_fa4_7_out(.a(s_csamul_rca12_and4_7[0]), .b(s_csamul_rca12_fa5_6_xor1[0]), .cin(s_csamul_rca12_fa4_6_or0[0]), .fa_xor1(s_csamul_rca12_fa4_7_xor1), .fa_or0(s_csamul_rca12_fa4_7_or0));
  and_gate and_gate_s_csamul_rca12_and5_7(.a(a[5]), .b(b[7]), .out(s_csamul_rca12_and5_7));
  fa fa_s_csamul_rca12_fa5_7_out(.a(s_csamul_rca12_and5_7[0]), .b(s_csamul_rca12_fa6_6_xor1[0]), .cin(s_csamul_rca12_fa5_6_or0[0]), .fa_xor1(s_csamul_rca12_fa5_7_xor1), .fa_or0(s_csamul_rca12_fa5_7_or0));
  and_gate and_gate_s_csamul_rca12_and6_7(.a(a[6]), .b(b[7]), .out(s_csamul_rca12_and6_7));
  fa fa_s_csamul_rca12_fa6_7_out(.a(s_csamul_rca12_and6_7[0]), .b(s_csamul_rca12_fa7_6_xor1[0]), .cin(s_csamul_rca12_fa6_6_or0[0]), .fa_xor1(s_csamul_rca12_fa6_7_xor1), .fa_or0(s_csamul_rca12_fa6_7_or0));
  and_gate and_gate_s_csamul_rca12_and7_7(.a(a[7]), .b(b[7]), .out(s_csamul_rca12_and7_7));
  fa fa_s_csamul_rca12_fa7_7_out(.a(s_csamul_rca12_and7_7[0]), .b(s_csamul_rca12_fa8_6_xor1[0]), .cin(s_csamul_rca12_fa7_6_or0[0]), .fa_xor1(s_csamul_rca12_fa7_7_xor1), .fa_or0(s_csamul_rca12_fa7_7_or0));
  and_gate and_gate_s_csamul_rca12_and8_7(.a(a[8]), .b(b[7]), .out(s_csamul_rca12_and8_7));
  fa fa_s_csamul_rca12_fa8_7_out(.a(s_csamul_rca12_and8_7[0]), .b(s_csamul_rca12_fa9_6_xor1[0]), .cin(s_csamul_rca12_fa8_6_or0[0]), .fa_xor1(s_csamul_rca12_fa8_7_xor1), .fa_or0(s_csamul_rca12_fa8_7_or0));
  and_gate and_gate_s_csamul_rca12_and9_7(.a(a[9]), .b(b[7]), .out(s_csamul_rca12_and9_7));
  fa fa_s_csamul_rca12_fa9_7_out(.a(s_csamul_rca12_and9_7[0]), .b(s_csamul_rca12_fa10_6_xor1[0]), .cin(s_csamul_rca12_fa9_6_or0[0]), .fa_xor1(s_csamul_rca12_fa9_7_xor1), .fa_or0(s_csamul_rca12_fa9_7_or0));
  and_gate and_gate_s_csamul_rca12_and10_7(.a(a[10]), .b(b[7]), .out(s_csamul_rca12_and10_7));
  fa fa_s_csamul_rca12_fa10_7_out(.a(s_csamul_rca12_and10_7[0]), .b(s_csamul_rca12_ha11_6_xor0[0]), .cin(s_csamul_rca12_fa10_6_or0[0]), .fa_xor1(s_csamul_rca12_fa10_7_xor1), .fa_or0(s_csamul_rca12_fa10_7_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_7(.a(a[11]), .b(b[7]), .out(s_csamul_rca12_nand11_7));
  ha ha_s_csamul_rca12_ha11_7_out(.a(s_csamul_rca12_nand11_7[0]), .b(s_csamul_rca12_ha11_6_and0[0]), .ha_xor0(s_csamul_rca12_ha11_7_xor0), .ha_and0(s_csamul_rca12_ha11_7_and0));
  and_gate and_gate_s_csamul_rca12_and0_8(.a(a[0]), .b(b[8]), .out(s_csamul_rca12_and0_8));
  fa fa_s_csamul_rca12_fa0_8_out(.a(s_csamul_rca12_and0_8[0]), .b(s_csamul_rca12_fa1_7_xor1[0]), .cin(s_csamul_rca12_fa0_7_or0[0]), .fa_xor1(s_csamul_rca12_fa0_8_xor1), .fa_or0(s_csamul_rca12_fa0_8_or0));
  and_gate and_gate_s_csamul_rca12_and1_8(.a(a[1]), .b(b[8]), .out(s_csamul_rca12_and1_8));
  fa fa_s_csamul_rca12_fa1_8_out(.a(s_csamul_rca12_and1_8[0]), .b(s_csamul_rca12_fa2_7_xor1[0]), .cin(s_csamul_rca12_fa1_7_or0[0]), .fa_xor1(s_csamul_rca12_fa1_8_xor1), .fa_or0(s_csamul_rca12_fa1_8_or0));
  and_gate and_gate_s_csamul_rca12_and2_8(.a(a[2]), .b(b[8]), .out(s_csamul_rca12_and2_8));
  fa fa_s_csamul_rca12_fa2_8_out(.a(s_csamul_rca12_and2_8[0]), .b(s_csamul_rca12_fa3_7_xor1[0]), .cin(s_csamul_rca12_fa2_7_or0[0]), .fa_xor1(s_csamul_rca12_fa2_8_xor1), .fa_or0(s_csamul_rca12_fa2_8_or0));
  and_gate and_gate_s_csamul_rca12_and3_8(.a(a[3]), .b(b[8]), .out(s_csamul_rca12_and3_8));
  fa fa_s_csamul_rca12_fa3_8_out(.a(s_csamul_rca12_and3_8[0]), .b(s_csamul_rca12_fa4_7_xor1[0]), .cin(s_csamul_rca12_fa3_7_or0[0]), .fa_xor1(s_csamul_rca12_fa3_8_xor1), .fa_or0(s_csamul_rca12_fa3_8_or0));
  and_gate and_gate_s_csamul_rca12_and4_8(.a(a[4]), .b(b[8]), .out(s_csamul_rca12_and4_8));
  fa fa_s_csamul_rca12_fa4_8_out(.a(s_csamul_rca12_and4_8[0]), .b(s_csamul_rca12_fa5_7_xor1[0]), .cin(s_csamul_rca12_fa4_7_or0[0]), .fa_xor1(s_csamul_rca12_fa4_8_xor1), .fa_or0(s_csamul_rca12_fa4_8_or0));
  and_gate and_gate_s_csamul_rca12_and5_8(.a(a[5]), .b(b[8]), .out(s_csamul_rca12_and5_8));
  fa fa_s_csamul_rca12_fa5_8_out(.a(s_csamul_rca12_and5_8[0]), .b(s_csamul_rca12_fa6_7_xor1[0]), .cin(s_csamul_rca12_fa5_7_or0[0]), .fa_xor1(s_csamul_rca12_fa5_8_xor1), .fa_or0(s_csamul_rca12_fa5_8_or0));
  and_gate and_gate_s_csamul_rca12_and6_8(.a(a[6]), .b(b[8]), .out(s_csamul_rca12_and6_8));
  fa fa_s_csamul_rca12_fa6_8_out(.a(s_csamul_rca12_and6_8[0]), .b(s_csamul_rca12_fa7_7_xor1[0]), .cin(s_csamul_rca12_fa6_7_or0[0]), .fa_xor1(s_csamul_rca12_fa6_8_xor1), .fa_or0(s_csamul_rca12_fa6_8_or0));
  and_gate and_gate_s_csamul_rca12_and7_8(.a(a[7]), .b(b[8]), .out(s_csamul_rca12_and7_8));
  fa fa_s_csamul_rca12_fa7_8_out(.a(s_csamul_rca12_and7_8[0]), .b(s_csamul_rca12_fa8_7_xor1[0]), .cin(s_csamul_rca12_fa7_7_or0[0]), .fa_xor1(s_csamul_rca12_fa7_8_xor1), .fa_or0(s_csamul_rca12_fa7_8_or0));
  and_gate and_gate_s_csamul_rca12_and8_8(.a(a[8]), .b(b[8]), .out(s_csamul_rca12_and8_8));
  fa fa_s_csamul_rca12_fa8_8_out(.a(s_csamul_rca12_and8_8[0]), .b(s_csamul_rca12_fa9_7_xor1[0]), .cin(s_csamul_rca12_fa8_7_or0[0]), .fa_xor1(s_csamul_rca12_fa8_8_xor1), .fa_or0(s_csamul_rca12_fa8_8_or0));
  and_gate and_gate_s_csamul_rca12_and9_8(.a(a[9]), .b(b[8]), .out(s_csamul_rca12_and9_8));
  fa fa_s_csamul_rca12_fa9_8_out(.a(s_csamul_rca12_and9_8[0]), .b(s_csamul_rca12_fa10_7_xor1[0]), .cin(s_csamul_rca12_fa9_7_or0[0]), .fa_xor1(s_csamul_rca12_fa9_8_xor1), .fa_or0(s_csamul_rca12_fa9_8_or0));
  and_gate and_gate_s_csamul_rca12_and10_8(.a(a[10]), .b(b[8]), .out(s_csamul_rca12_and10_8));
  fa fa_s_csamul_rca12_fa10_8_out(.a(s_csamul_rca12_and10_8[0]), .b(s_csamul_rca12_ha11_7_xor0[0]), .cin(s_csamul_rca12_fa10_7_or0[0]), .fa_xor1(s_csamul_rca12_fa10_8_xor1), .fa_or0(s_csamul_rca12_fa10_8_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_8(.a(a[11]), .b(b[8]), .out(s_csamul_rca12_nand11_8));
  ha ha_s_csamul_rca12_ha11_8_out(.a(s_csamul_rca12_nand11_8[0]), .b(s_csamul_rca12_ha11_7_and0[0]), .ha_xor0(s_csamul_rca12_ha11_8_xor0), .ha_and0(s_csamul_rca12_ha11_8_and0));
  and_gate and_gate_s_csamul_rca12_and0_9(.a(a[0]), .b(b[9]), .out(s_csamul_rca12_and0_9));
  fa fa_s_csamul_rca12_fa0_9_out(.a(s_csamul_rca12_and0_9[0]), .b(s_csamul_rca12_fa1_8_xor1[0]), .cin(s_csamul_rca12_fa0_8_or0[0]), .fa_xor1(s_csamul_rca12_fa0_9_xor1), .fa_or0(s_csamul_rca12_fa0_9_or0));
  and_gate and_gate_s_csamul_rca12_and1_9(.a(a[1]), .b(b[9]), .out(s_csamul_rca12_and1_9));
  fa fa_s_csamul_rca12_fa1_9_out(.a(s_csamul_rca12_and1_9[0]), .b(s_csamul_rca12_fa2_8_xor1[0]), .cin(s_csamul_rca12_fa1_8_or0[0]), .fa_xor1(s_csamul_rca12_fa1_9_xor1), .fa_or0(s_csamul_rca12_fa1_9_or0));
  and_gate and_gate_s_csamul_rca12_and2_9(.a(a[2]), .b(b[9]), .out(s_csamul_rca12_and2_9));
  fa fa_s_csamul_rca12_fa2_9_out(.a(s_csamul_rca12_and2_9[0]), .b(s_csamul_rca12_fa3_8_xor1[0]), .cin(s_csamul_rca12_fa2_8_or0[0]), .fa_xor1(s_csamul_rca12_fa2_9_xor1), .fa_or0(s_csamul_rca12_fa2_9_or0));
  and_gate and_gate_s_csamul_rca12_and3_9(.a(a[3]), .b(b[9]), .out(s_csamul_rca12_and3_9));
  fa fa_s_csamul_rca12_fa3_9_out(.a(s_csamul_rca12_and3_9[0]), .b(s_csamul_rca12_fa4_8_xor1[0]), .cin(s_csamul_rca12_fa3_8_or0[0]), .fa_xor1(s_csamul_rca12_fa3_9_xor1), .fa_or0(s_csamul_rca12_fa3_9_or0));
  and_gate and_gate_s_csamul_rca12_and4_9(.a(a[4]), .b(b[9]), .out(s_csamul_rca12_and4_9));
  fa fa_s_csamul_rca12_fa4_9_out(.a(s_csamul_rca12_and4_9[0]), .b(s_csamul_rca12_fa5_8_xor1[0]), .cin(s_csamul_rca12_fa4_8_or0[0]), .fa_xor1(s_csamul_rca12_fa4_9_xor1), .fa_or0(s_csamul_rca12_fa4_9_or0));
  and_gate and_gate_s_csamul_rca12_and5_9(.a(a[5]), .b(b[9]), .out(s_csamul_rca12_and5_9));
  fa fa_s_csamul_rca12_fa5_9_out(.a(s_csamul_rca12_and5_9[0]), .b(s_csamul_rca12_fa6_8_xor1[0]), .cin(s_csamul_rca12_fa5_8_or0[0]), .fa_xor1(s_csamul_rca12_fa5_9_xor1), .fa_or0(s_csamul_rca12_fa5_9_or0));
  and_gate and_gate_s_csamul_rca12_and6_9(.a(a[6]), .b(b[9]), .out(s_csamul_rca12_and6_9));
  fa fa_s_csamul_rca12_fa6_9_out(.a(s_csamul_rca12_and6_9[0]), .b(s_csamul_rca12_fa7_8_xor1[0]), .cin(s_csamul_rca12_fa6_8_or0[0]), .fa_xor1(s_csamul_rca12_fa6_9_xor1), .fa_or0(s_csamul_rca12_fa6_9_or0));
  and_gate and_gate_s_csamul_rca12_and7_9(.a(a[7]), .b(b[9]), .out(s_csamul_rca12_and7_9));
  fa fa_s_csamul_rca12_fa7_9_out(.a(s_csamul_rca12_and7_9[0]), .b(s_csamul_rca12_fa8_8_xor1[0]), .cin(s_csamul_rca12_fa7_8_or0[0]), .fa_xor1(s_csamul_rca12_fa7_9_xor1), .fa_or0(s_csamul_rca12_fa7_9_or0));
  and_gate and_gate_s_csamul_rca12_and8_9(.a(a[8]), .b(b[9]), .out(s_csamul_rca12_and8_9));
  fa fa_s_csamul_rca12_fa8_9_out(.a(s_csamul_rca12_and8_9[0]), .b(s_csamul_rca12_fa9_8_xor1[0]), .cin(s_csamul_rca12_fa8_8_or0[0]), .fa_xor1(s_csamul_rca12_fa8_9_xor1), .fa_or0(s_csamul_rca12_fa8_9_or0));
  and_gate and_gate_s_csamul_rca12_and9_9(.a(a[9]), .b(b[9]), .out(s_csamul_rca12_and9_9));
  fa fa_s_csamul_rca12_fa9_9_out(.a(s_csamul_rca12_and9_9[0]), .b(s_csamul_rca12_fa10_8_xor1[0]), .cin(s_csamul_rca12_fa9_8_or0[0]), .fa_xor1(s_csamul_rca12_fa9_9_xor1), .fa_or0(s_csamul_rca12_fa9_9_or0));
  and_gate and_gate_s_csamul_rca12_and10_9(.a(a[10]), .b(b[9]), .out(s_csamul_rca12_and10_9));
  fa fa_s_csamul_rca12_fa10_9_out(.a(s_csamul_rca12_and10_9[0]), .b(s_csamul_rca12_ha11_8_xor0[0]), .cin(s_csamul_rca12_fa10_8_or0[0]), .fa_xor1(s_csamul_rca12_fa10_9_xor1), .fa_or0(s_csamul_rca12_fa10_9_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_9(.a(a[11]), .b(b[9]), .out(s_csamul_rca12_nand11_9));
  ha ha_s_csamul_rca12_ha11_9_out(.a(s_csamul_rca12_nand11_9[0]), .b(s_csamul_rca12_ha11_8_and0[0]), .ha_xor0(s_csamul_rca12_ha11_9_xor0), .ha_and0(s_csamul_rca12_ha11_9_and0));
  and_gate and_gate_s_csamul_rca12_and0_10(.a(a[0]), .b(b[10]), .out(s_csamul_rca12_and0_10));
  fa fa_s_csamul_rca12_fa0_10_out(.a(s_csamul_rca12_and0_10[0]), .b(s_csamul_rca12_fa1_9_xor1[0]), .cin(s_csamul_rca12_fa0_9_or0[0]), .fa_xor1(s_csamul_rca12_fa0_10_xor1), .fa_or0(s_csamul_rca12_fa0_10_or0));
  and_gate and_gate_s_csamul_rca12_and1_10(.a(a[1]), .b(b[10]), .out(s_csamul_rca12_and1_10));
  fa fa_s_csamul_rca12_fa1_10_out(.a(s_csamul_rca12_and1_10[0]), .b(s_csamul_rca12_fa2_9_xor1[0]), .cin(s_csamul_rca12_fa1_9_or0[0]), .fa_xor1(s_csamul_rca12_fa1_10_xor1), .fa_or0(s_csamul_rca12_fa1_10_or0));
  and_gate and_gate_s_csamul_rca12_and2_10(.a(a[2]), .b(b[10]), .out(s_csamul_rca12_and2_10));
  fa fa_s_csamul_rca12_fa2_10_out(.a(s_csamul_rca12_and2_10[0]), .b(s_csamul_rca12_fa3_9_xor1[0]), .cin(s_csamul_rca12_fa2_9_or0[0]), .fa_xor1(s_csamul_rca12_fa2_10_xor1), .fa_or0(s_csamul_rca12_fa2_10_or0));
  and_gate and_gate_s_csamul_rca12_and3_10(.a(a[3]), .b(b[10]), .out(s_csamul_rca12_and3_10));
  fa fa_s_csamul_rca12_fa3_10_out(.a(s_csamul_rca12_and3_10[0]), .b(s_csamul_rca12_fa4_9_xor1[0]), .cin(s_csamul_rca12_fa3_9_or0[0]), .fa_xor1(s_csamul_rca12_fa3_10_xor1), .fa_or0(s_csamul_rca12_fa3_10_or0));
  and_gate and_gate_s_csamul_rca12_and4_10(.a(a[4]), .b(b[10]), .out(s_csamul_rca12_and4_10));
  fa fa_s_csamul_rca12_fa4_10_out(.a(s_csamul_rca12_and4_10[0]), .b(s_csamul_rca12_fa5_9_xor1[0]), .cin(s_csamul_rca12_fa4_9_or0[0]), .fa_xor1(s_csamul_rca12_fa4_10_xor1), .fa_or0(s_csamul_rca12_fa4_10_or0));
  and_gate and_gate_s_csamul_rca12_and5_10(.a(a[5]), .b(b[10]), .out(s_csamul_rca12_and5_10));
  fa fa_s_csamul_rca12_fa5_10_out(.a(s_csamul_rca12_and5_10[0]), .b(s_csamul_rca12_fa6_9_xor1[0]), .cin(s_csamul_rca12_fa5_9_or0[0]), .fa_xor1(s_csamul_rca12_fa5_10_xor1), .fa_or0(s_csamul_rca12_fa5_10_or0));
  and_gate and_gate_s_csamul_rca12_and6_10(.a(a[6]), .b(b[10]), .out(s_csamul_rca12_and6_10));
  fa fa_s_csamul_rca12_fa6_10_out(.a(s_csamul_rca12_and6_10[0]), .b(s_csamul_rca12_fa7_9_xor1[0]), .cin(s_csamul_rca12_fa6_9_or0[0]), .fa_xor1(s_csamul_rca12_fa6_10_xor1), .fa_or0(s_csamul_rca12_fa6_10_or0));
  and_gate and_gate_s_csamul_rca12_and7_10(.a(a[7]), .b(b[10]), .out(s_csamul_rca12_and7_10));
  fa fa_s_csamul_rca12_fa7_10_out(.a(s_csamul_rca12_and7_10[0]), .b(s_csamul_rca12_fa8_9_xor1[0]), .cin(s_csamul_rca12_fa7_9_or0[0]), .fa_xor1(s_csamul_rca12_fa7_10_xor1), .fa_or0(s_csamul_rca12_fa7_10_or0));
  and_gate and_gate_s_csamul_rca12_and8_10(.a(a[8]), .b(b[10]), .out(s_csamul_rca12_and8_10));
  fa fa_s_csamul_rca12_fa8_10_out(.a(s_csamul_rca12_and8_10[0]), .b(s_csamul_rca12_fa9_9_xor1[0]), .cin(s_csamul_rca12_fa8_9_or0[0]), .fa_xor1(s_csamul_rca12_fa8_10_xor1), .fa_or0(s_csamul_rca12_fa8_10_or0));
  and_gate and_gate_s_csamul_rca12_and9_10(.a(a[9]), .b(b[10]), .out(s_csamul_rca12_and9_10));
  fa fa_s_csamul_rca12_fa9_10_out(.a(s_csamul_rca12_and9_10[0]), .b(s_csamul_rca12_fa10_9_xor1[0]), .cin(s_csamul_rca12_fa9_9_or0[0]), .fa_xor1(s_csamul_rca12_fa9_10_xor1), .fa_or0(s_csamul_rca12_fa9_10_or0));
  and_gate and_gate_s_csamul_rca12_and10_10(.a(a[10]), .b(b[10]), .out(s_csamul_rca12_and10_10));
  fa fa_s_csamul_rca12_fa10_10_out(.a(s_csamul_rca12_and10_10[0]), .b(s_csamul_rca12_ha11_9_xor0[0]), .cin(s_csamul_rca12_fa10_9_or0[0]), .fa_xor1(s_csamul_rca12_fa10_10_xor1), .fa_or0(s_csamul_rca12_fa10_10_or0));
  nand_gate nand_gate_s_csamul_rca12_nand11_10(.a(a[11]), .b(b[10]), .out(s_csamul_rca12_nand11_10));
  ha ha_s_csamul_rca12_ha11_10_out(.a(s_csamul_rca12_nand11_10[0]), .b(s_csamul_rca12_ha11_9_and0[0]), .ha_xor0(s_csamul_rca12_ha11_10_xor0), .ha_and0(s_csamul_rca12_ha11_10_and0));
  nand_gate nand_gate_s_csamul_rca12_nand0_11(.a(a[0]), .b(b[11]), .out(s_csamul_rca12_nand0_11));
  fa fa_s_csamul_rca12_fa0_11_out(.a(s_csamul_rca12_nand0_11[0]), .b(s_csamul_rca12_fa1_10_xor1[0]), .cin(s_csamul_rca12_fa0_10_or0[0]), .fa_xor1(s_csamul_rca12_fa0_11_xor1), .fa_or0(s_csamul_rca12_fa0_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand1_11(.a(a[1]), .b(b[11]), .out(s_csamul_rca12_nand1_11));
  fa fa_s_csamul_rca12_fa1_11_out(.a(s_csamul_rca12_nand1_11[0]), .b(s_csamul_rca12_fa2_10_xor1[0]), .cin(s_csamul_rca12_fa1_10_or0[0]), .fa_xor1(s_csamul_rca12_fa1_11_xor1), .fa_or0(s_csamul_rca12_fa1_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand2_11(.a(a[2]), .b(b[11]), .out(s_csamul_rca12_nand2_11));
  fa fa_s_csamul_rca12_fa2_11_out(.a(s_csamul_rca12_nand2_11[0]), .b(s_csamul_rca12_fa3_10_xor1[0]), .cin(s_csamul_rca12_fa2_10_or0[0]), .fa_xor1(s_csamul_rca12_fa2_11_xor1), .fa_or0(s_csamul_rca12_fa2_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand3_11(.a(a[3]), .b(b[11]), .out(s_csamul_rca12_nand3_11));
  fa fa_s_csamul_rca12_fa3_11_out(.a(s_csamul_rca12_nand3_11[0]), .b(s_csamul_rca12_fa4_10_xor1[0]), .cin(s_csamul_rca12_fa3_10_or0[0]), .fa_xor1(s_csamul_rca12_fa3_11_xor1), .fa_or0(s_csamul_rca12_fa3_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand4_11(.a(a[4]), .b(b[11]), .out(s_csamul_rca12_nand4_11));
  fa fa_s_csamul_rca12_fa4_11_out(.a(s_csamul_rca12_nand4_11[0]), .b(s_csamul_rca12_fa5_10_xor1[0]), .cin(s_csamul_rca12_fa4_10_or0[0]), .fa_xor1(s_csamul_rca12_fa4_11_xor1), .fa_or0(s_csamul_rca12_fa4_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand5_11(.a(a[5]), .b(b[11]), .out(s_csamul_rca12_nand5_11));
  fa fa_s_csamul_rca12_fa5_11_out(.a(s_csamul_rca12_nand5_11[0]), .b(s_csamul_rca12_fa6_10_xor1[0]), .cin(s_csamul_rca12_fa5_10_or0[0]), .fa_xor1(s_csamul_rca12_fa5_11_xor1), .fa_or0(s_csamul_rca12_fa5_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand6_11(.a(a[6]), .b(b[11]), .out(s_csamul_rca12_nand6_11));
  fa fa_s_csamul_rca12_fa6_11_out(.a(s_csamul_rca12_nand6_11[0]), .b(s_csamul_rca12_fa7_10_xor1[0]), .cin(s_csamul_rca12_fa6_10_or0[0]), .fa_xor1(s_csamul_rca12_fa6_11_xor1), .fa_or0(s_csamul_rca12_fa6_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand7_11(.a(a[7]), .b(b[11]), .out(s_csamul_rca12_nand7_11));
  fa fa_s_csamul_rca12_fa7_11_out(.a(s_csamul_rca12_nand7_11[0]), .b(s_csamul_rca12_fa8_10_xor1[0]), .cin(s_csamul_rca12_fa7_10_or0[0]), .fa_xor1(s_csamul_rca12_fa7_11_xor1), .fa_or0(s_csamul_rca12_fa7_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand8_11(.a(a[8]), .b(b[11]), .out(s_csamul_rca12_nand8_11));
  fa fa_s_csamul_rca12_fa8_11_out(.a(s_csamul_rca12_nand8_11[0]), .b(s_csamul_rca12_fa9_10_xor1[0]), .cin(s_csamul_rca12_fa8_10_or0[0]), .fa_xor1(s_csamul_rca12_fa8_11_xor1), .fa_or0(s_csamul_rca12_fa8_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand9_11(.a(a[9]), .b(b[11]), .out(s_csamul_rca12_nand9_11));
  fa fa_s_csamul_rca12_fa9_11_out(.a(s_csamul_rca12_nand9_11[0]), .b(s_csamul_rca12_fa10_10_xor1[0]), .cin(s_csamul_rca12_fa9_10_or0[0]), .fa_xor1(s_csamul_rca12_fa9_11_xor1), .fa_or0(s_csamul_rca12_fa9_11_or0));
  nand_gate nand_gate_s_csamul_rca12_nand10_11(.a(a[10]), .b(b[11]), .out(s_csamul_rca12_nand10_11));
  fa fa_s_csamul_rca12_fa10_11_out(.a(s_csamul_rca12_nand10_11[0]), .b(s_csamul_rca12_ha11_10_xor0[0]), .cin(s_csamul_rca12_fa10_10_or0[0]), .fa_xor1(s_csamul_rca12_fa10_11_xor1), .fa_or0(s_csamul_rca12_fa10_11_or0));
  and_gate and_gate_s_csamul_rca12_and11_11(.a(a[11]), .b(b[11]), .out(s_csamul_rca12_and11_11));
  ha ha_s_csamul_rca12_ha11_11_out(.a(s_csamul_rca12_and11_11[0]), .b(s_csamul_rca12_ha11_10_and0[0]), .ha_xor0(s_csamul_rca12_ha11_11_xor0), .ha_and0(s_csamul_rca12_ha11_11_and0));
  assign s_csamul_rca12_u_rca12_a[0] = s_csamul_rca12_fa1_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[1] = s_csamul_rca12_fa2_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[2] = s_csamul_rca12_fa3_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[3] = s_csamul_rca12_fa4_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[4] = s_csamul_rca12_fa5_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[5] = s_csamul_rca12_fa6_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[6] = s_csamul_rca12_fa7_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[7] = s_csamul_rca12_fa8_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[8] = s_csamul_rca12_fa9_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[9] = s_csamul_rca12_fa10_11_xor1[0];
  assign s_csamul_rca12_u_rca12_a[10] = s_csamul_rca12_ha11_11_xor0[0];
  assign s_csamul_rca12_u_rca12_a[11] = 1'b1;
  assign s_csamul_rca12_u_rca12_b[0] = s_csamul_rca12_fa0_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[1] = s_csamul_rca12_fa1_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[2] = s_csamul_rca12_fa2_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[3] = s_csamul_rca12_fa3_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[4] = s_csamul_rca12_fa4_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[5] = s_csamul_rca12_fa5_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[6] = s_csamul_rca12_fa6_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[7] = s_csamul_rca12_fa7_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[8] = s_csamul_rca12_fa8_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[9] = s_csamul_rca12_fa9_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[10] = s_csamul_rca12_fa10_11_or0[0];
  assign s_csamul_rca12_u_rca12_b[11] = s_csamul_rca12_ha11_11_and0[0];
  u_rca12 u_rca12_s_csamul_rca12_u_rca12_out(.a(s_csamul_rca12_u_rca12_a), .b(s_csamul_rca12_u_rca12_b), .u_rca12_out(s_csamul_rca12_u_rca12_out));

  assign s_csamul_rca12_out[0] = s_csamul_rca12_and0_0[0];
  assign s_csamul_rca12_out[1] = s_csamul_rca12_ha0_1_xor0[0];
  assign s_csamul_rca12_out[2] = s_csamul_rca12_fa0_2_xor1[0];
  assign s_csamul_rca12_out[3] = s_csamul_rca12_fa0_3_xor1[0];
  assign s_csamul_rca12_out[4] = s_csamul_rca12_fa0_4_xor1[0];
  assign s_csamul_rca12_out[5] = s_csamul_rca12_fa0_5_xor1[0];
  assign s_csamul_rca12_out[6] = s_csamul_rca12_fa0_6_xor1[0];
  assign s_csamul_rca12_out[7] = s_csamul_rca12_fa0_7_xor1[0];
  assign s_csamul_rca12_out[8] = s_csamul_rca12_fa0_8_xor1[0];
  assign s_csamul_rca12_out[9] = s_csamul_rca12_fa0_9_xor1[0];
  assign s_csamul_rca12_out[10] = s_csamul_rca12_fa0_10_xor1[0];
  assign s_csamul_rca12_out[11] = s_csamul_rca12_fa0_11_xor1[0];
  assign s_csamul_rca12_out[12] = s_csamul_rca12_u_rca12_out[0];
  assign s_csamul_rca12_out[13] = s_csamul_rca12_u_rca12_out[1];
  assign s_csamul_rca12_out[14] = s_csamul_rca12_u_rca12_out[2];
  assign s_csamul_rca12_out[15] = s_csamul_rca12_u_rca12_out[3];
  assign s_csamul_rca12_out[16] = s_csamul_rca12_u_rca12_out[4];
  assign s_csamul_rca12_out[17] = s_csamul_rca12_u_rca12_out[5];
  assign s_csamul_rca12_out[18] = s_csamul_rca12_u_rca12_out[6];
  assign s_csamul_rca12_out[19] = s_csamul_rca12_u_rca12_out[7];
  assign s_csamul_rca12_out[20] = s_csamul_rca12_u_rca12_out[8];
  assign s_csamul_rca12_out[21] = s_csamul_rca12_u_rca12_out[9];
  assign s_csamul_rca12_out[22] = s_csamul_rca12_u_rca12_out[10];
  assign s_csamul_rca12_out[23] = s_csamul_rca12_u_rca12_out[11];
endmodule