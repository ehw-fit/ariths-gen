module s_cla4(input [3:0] a, input [3:0] b, output [4:0] s_cla4_out);
  wire s_cla4_pg_logic0_or0;
  wire s_cla4_pg_logic0_and0;
  wire s_cla4_pg_logic0_xor0;
  wire s_cla4_pg_logic1_or0;
  wire s_cla4_pg_logic1_and0;
  wire s_cla4_pg_logic1_xor0;
  wire s_cla4_xor1;
  wire s_cla4_and0;
  wire s_cla4_or0;
  wire s_cla4_pg_logic2_or0;
  wire s_cla4_pg_logic2_and0;
  wire s_cla4_pg_logic2_xor0;
  wire s_cla4_xor2;
  wire s_cla4_and1;
  wire s_cla4_and2;
  wire s_cla4_and3;
  wire s_cla4_and4;
  wire s_cla4_or1;
  wire s_cla4_or2;
  wire s_cla4_pg_logic3_or0;
  wire s_cla4_pg_logic3_and0;
  wire s_cla4_pg_logic3_xor0;
  wire s_cla4_xor3;
  wire s_cla4_and5;
  wire s_cla4_and6;
  wire s_cla4_and7;
  wire s_cla4_and8;
  wire s_cla4_and9;
  wire s_cla4_and10;
  wire s_cla4_and11;
  wire s_cla4_or3;
  wire s_cla4_or4;
  wire s_cla4_or5;
  wire s_cla4_xor4;
  wire s_cla4_xor5;

  assign s_cla4_pg_logic0_or0 = a[0] | b[0];
  assign s_cla4_pg_logic0_and0 = a[0] & b[0];
  assign s_cla4_pg_logic0_xor0 = a[0] ^ b[0];
  assign s_cla4_pg_logic1_or0 = a[1] | b[1];
  assign s_cla4_pg_logic1_and0 = a[1] & b[1];
  assign s_cla4_pg_logic1_xor0 = a[1] ^ b[1];
  assign s_cla4_xor1 = s_cla4_pg_logic1_xor0 ^ s_cla4_pg_logic0_and0;
  assign s_cla4_and0 = s_cla4_pg_logic0_and0 & s_cla4_pg_logic1_or0;
  assign s_cla4_or0 = s_cla4_pg_logic1_and0 | s_cla4_and0;
  assign s_cla4_pg_logic2_or0 = a[2] | b[2];
  assign s_cla4_pg_logic2_and0 = a[2] & b[2];
  assign s_cla4_pg_logic2_xor0 = a[2] ^ b[2];
  assign s_cla4_xor2 = s_cla4_pg_logic2_xor0 ^ s_cla4_or0;
  assign s_cla4_and1 = s_cla4_pg_logic2_or0 & s_cla4_pg_logic0_or0;
  assign s_cla4_and2 = s_cla4_pg_logic0_and0 & s_cla4_pg_logic2_or0;
  assign s_cla4_and3 = s_cla4_and2 & s_cla4_pg_logic1_or0;
  assign s_cla4_and4 = s_cla4_pg_logic1_and0 & s_cla4_pg_logic2_or0;
  assign s_cla4_or1 = s_cla4_and3 | s_cla4_and4;
  assign s_cla4_or2 = s_cla4_pg_logic2_and0 | s_cla4_or1;
  assign s_cla4_pg_logic3_or0 = a[3] | b[3];
  assign s_cla4_pg_logic3_and0 = a[3] & b[3];
  assign s_cla4_pg_logic3_xor0 = a[3] ^ b[3];
  assign s_cla4_xor3 = s_cla4_pg_logic3_xor0 ^ s_cla4_or2;
  assign s_cla4_and5 = s_cla4_pg_logic3_or0 & s_cla4_pg_logic1_or0;
  assign s_cla4_and6 = s_cla4_pg_logic0_and0 & s_cla4_pg_logic2_or0;
  assign s_cla4_and7 = s_cla4_pg_logic3_or0 & s_cla4_pg_logic1_or0;
  assign s_cla4_and8 = s_cla4_and6 & s_cla4_and7;
  assign s_cla4_and9 = s_cla4_pg_logic1_and0 & s_cla4_pg_logic3_or0;
  assign s_cla4_and10 = s_cla4_and9 & s_cla4_pg_logic2_or0;
  assign s_cla4_and11 = s_cla4_pg_logic2_and0 & s_cla4_pg_logic3_or0;
  assign s_cla4_or3 = s_cla4_and8 | s_cla4_and11;
  assign s_cla4_or4 = s_cla4_and10 | s_cla4_or3;
  assign s_cla4_or5 = s_cla4_pg_logic3_and0 | s_cla4_or4;
  assign s_cla4_xor4 = a[3] ^ b[3];
  assign s_cla4_xor5 = s_cla4_xor4 ^ s_cla4_or5;

  assign s_cla4_out[0] = s_cla4_pg_logic0_xor0;
  assign s_cla4_out[1] = s_cla4_xor1;
  assign s_cla4_out[2] = s_cla4_xor2;
  assign s_cla4_out[3] = s_cla4_xor3;
  assign s_cla4_out[4] = s_cla4_xor5;
endmodule