module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module csa_component26(input [25:0] a, input [25:0] b, input [25:0] c, output [53:0] csa_component26_out);
  wire [0:0] csa_component26_fa0_xor1;
  wire [0:0] csa_component26_fa0_or0;
  wire [0:0] csa_component26_fa1_xor1;
  wire [0:0] csa_component26_fa1_or0;
  wire [0:0] csa_component26_fa2_xor1;
  wire [0:0] csa_component26_fa2_or0;
  wire [0:0] csa_component26_fa3_xor1;
  wire [0:0] csa_component26_fa3_or0;
  wire [0:0] csa_component26_fa4_xor1;
  wire [0:0] csa_component26_fa4_or0;
  wire [0:0] csa_component26_fa5_xor1;
  wire [0:0] csa_component26_fa5_or0;
  wire [0:0] csa_component26_fa6_xor1;
  wire [0:0] csa_component26_fa6_or0;
  wire [0:0] csa_component26_fa7_xor1;
  wire [0:0] csa_component26_fa7_or0;
  wire [0:0] csa_component26_fa8_xor1;
  wire [0:0] csa_component26_fa8_or0;
  wire [0:0] csa_component26_fa9_xor1;
  wire [0:0] csa_component26_fa9_or0;
  wire [0:0] csa_component26_fa10_xor1;
  wire [0:0] csa_component26_fa10_or0;
  wire [0:0] csa_component26_fa11_xor1;
  wire [0:0] csa_component26_fa11_or0;
  wire [0:0] csa_component26_fa12_xor1;
  wire [0:0] csa_component26_fa12_or0;
  wire [0:0] csa_component26_fa13_xor1;
  wire [0:0] csa_component26_fa13_or0;
  wire [0:0] csa_component26_fa14_xor1;
  wire [0:0] csa_component26_fa14_or0;
  wire [0:0] csa_component26_fa15_xor1;
  wire [0:0] csa_component26_fa15_or0;
  wire [0:0] csa_component26_fa16_xor1;
  wire [0:0] csa_component26_fa16_or0;
  wire [0:0] csa_component26_fa17_xor1;
  wire [0:0] csa_component26_fa17_or0;
  wire [0:0] csa_component26_fa18_xor1;
  wire [0:0] csa_component26_fa18_or0;
  wire [0:0] csa_component26_fa19_xor1;
  wire [0:0] csa_component26_fa19_or0;
  wire [0:0] csa_component26_fa20_xor1;
  wire [0:0] csa_component26_fa20_or0;
  wire [0:0] csa_component26_fa21_xor1;
  wire [0:0] csa_component26_fa21_or0;
  wire [0:0] csa_component26_fa22_xor1;
  wire [0:0] csa_component26_fa22_or0;
  wire [0:0] csa_component26_fa23_xor1;
  wire [0:0] csa_component26_fa23_or0;
  wire [0:0] csa_component26_fa24_xor1;
  wire [0:0] csa_component26_fa24_or0;
  wire [0:0] csa_component26_fa25_xor1;
  wire [0:0] csa_component26_fa25_or0;

  fa fa_csa_component26_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component26_fa0_xor1), .fa_or0(csa_component26_fa0_or0));
  fa fa_csa_component26_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component26_fa1_xor1), .fa_or0(csa_component26_fa1_or0));
  fa fa_csa_component26_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component26_fa2_xor1), .fa_or0(csa_component26_fa2_or0));
  fa fa_csa_component26_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component26_fa3_xor1), .fa_or0(csa_component26_fa3_or0));
  fa fa_csa_component26_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component26_fa4_xor1), .fa_or0(csa_component26_fa4_or0));
  fa fa_csa_component26_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component26_fa5_xor1), .fa_or0(csa_component26_fa5_or0));
  fa fa_csa_component26_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component26_fa6_xor1), .fa_or0(csa_component26_fa6_or0));
  fa fa_csa_component26_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component26_fa7_xor1), .fa_or0(csa_component26_fa7_or0));
  fa fa_csa_component26_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component26_fa8_xor1), .fa_or0(csa_component26_fa8_or0));
  fa fa_csa_component26_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component26_fa9_xor1), .fa_or0(csa_component26_fa9_or0));
  fa fa_csa_component26_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component26_fa10_xor1), .fa_or0(csa_component26_fa10_or0));
  fa fa_csa_component26_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component26_fa11_xor1), .fa_or0(csa_component26_fa11_or0));
  fa fa_csa_component26_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component26_fa12_xor1), .fa_or0(csa_component26_fa12_or0));
  fa fa_csa_component26_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component26_fa13_xor1), .fa_or0(csa_component26_fa13_or0));
  fa fa_csa_component26_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component26_fa14_xor1), .fa_or0(csa_component26_fa14_or0));
  fa fa_csa_component26_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component26_fa15_xor1), .fa_or0(csa_component26_fa15_or0));
  fa fa_csa_component26_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component26_fa16_xor1), .fa_or0(csa_component26_fa16_or0));
  fa fa_csa_component26_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component26_fa17_xor1), .fa_or0(csa_component26_fa17_or0));
  fa fa_csa_component26_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component26_fa18_xor1), .fa_or0(csa_component26_fa18_or0));
  fa fa_csa_component26_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component26_fa19_xor1), .fa_or0(csa_component26_fa19_or0));
  fa fa_csa_component26_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component26_fa20_xor1), .fa_or0(csa_component26_fa20_or0));
  fa fa_csa_component26_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component26_fa21_xor1), .fa_or0(csa_component26_fa21_or0));
  fa fa_csa_component26_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component26_fa22_xor1), .fa_or0(csa_component26_fa22_or0));
  fa fa_csa_component26_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component26_fa23_xor1), .fa_or0(csa_component26_fa23_or0));
  fa fa_csa_component26_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component26_fa24_xor1), .fa_or0(csa_component26_fa24_or0));
  fa fa_csa_component26_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component26_fa25_xor1), .fa_or0(csa_component26_fa25_or0));

  assign csa_component26_out[0] = csa_component26_fa0_xor1[0];
  assign csa_component26_out[1] = csa_component26_fa1_xor1[0];
  assign csa_component26_out[2] = csa_component26_fa2_xor1[0];
  assign csa_component26_out[3] = csa_component26_fa3_xor1[0];
  assign csa_component26_out[4] = csa_component26_fa4_xor1[0];
  assign csa_component26_out[5] = csa_component26_fa5_xor1[0];
  assign csa_component26_out[6] = csa_component26_fa6_xor1[0];
  assign csa_component26_out[7] = csa_component26_fa7_xor1[0];
  assign csa_component26_out[8] = csa_component26_fa8_xor1[0];
  assign csa_component26_out[9] = csa_component26_fa9_xor1[0];
  assign csa_component26_out[10] = csa_component26_fa10_xor1[0];
  assign csa_component26_out[11] = csa_component26_fa11_xor1[0];
  assign csa_component26_out[12] = csa_component26_fa12_xor1[0];
  assign csa_component26_out[13] = csa_component26_fa13_xor1[0];
  assign csa_component26_out[14] = csa_component26_fa14_xor1[0];
  assign csa_component26_out[15] = csa_component26_fa15_xor1[0];
  assign csa_component26_out[16] = csa_component26_fa16_xor1[0];
  assign csa_component26_out[17] = csa_component26_fa17_xor1[0];
  assign csa_component26_out[18] = csa_component26_fa18_xor1[0];
  assign csa_component26_out[19] = csa_component26_fa19_xor1[0];
  assign csa_component26_out[20] = csa_component26_fa20_xor1[0];
  assign csa_component26_out[21] = csa_component26_fa21_xor1[0];
  assign csa_component26_out[22] = csa_component26_fa22_xor1[0];
  assign csa_component26_out[23] = csa_component26_fa23_xor1[0];
  assign csa_component26_out[24] = csa_component26_fa24_xor1[0];
  assign csa_component26_out[25] = csa_component26_fa25_xor1[0];
  assign csa_component26_out[26] = 1'b0;
  assign csa_component26_out[27] = 1'b0;
  assign csa_component26_out[28] = csa_component26_fa0_or0[0];
  assign csa_component26_out[29] = csa_component26_fa1_or0[0];
  assign csa_component26_out[30] = csa_component26_fa2_or0[0];
  assign csa_component26_out[31] = csa_component26_fa3_or0[0];
  assign csa_component26_out[32] = csa_component26_fa4_or0[0];
  assign csa_component26_out[33] = csa_component26_fa5_or0[0];
  assign csa_component26_out[34] = csa_component26_fa6_or0[0];
  assign csa_component26_out[35] = csa_component26_fa7_or0[0];
  assign csa_component26_out[36] = csa_component26_fa8_or0[0];
  assign csa_component26_out[37] = csa_component26_fa9_or0[0];
  assign csa_component26_out[38] = csa_component26_fa10_or0[0];
  assign csa_component26_out[39] = csa_component26_fa11_or0[0];
  assign csa_component26_out[40] = csa_component26_fa12_or0[0];
  assign csa_component26_out[41] = csa_component26_fa13_or0[0];
  assign csa_component26_out[42] = csa_component26_fa14_or0[0];
  assign csa_component26_out[43] = csa_component26_fa15_or0[0];
  assign csa_component26_out[44] = csa_component26_fa16_or0[0];
  assign csa_component26_out[45] = csa_component26_fa17_or0[0];
  assign csa_component26_out[46] = csa_component26_fa18_or0[0];
  assign csa_component26_out[47] = csa_component26_fa19_or0[0];
  assign csa_component26_out[48] = csa_component26_fa20_or0[0];
  assign csa_component26_out[49] = csa_component26_fa21_or0[0];
  assign csa_component26_out[50] = csa_component26_fa22_or0[0];
  assign csa_component26_out[51] = csa_component26_fa23_or0[0];
  assign csa_component26_out[52] = csa_component26_fa24_or0[0];
  assign csa_component26_out[53] = csa_component26_fa25_or0[0];
endmodule

module csa_component29(input [28:0] a, input [28:0] b, input [28:0] c, output [59:0] csa_component29_out);
  wire [0:0] csa_component29_fa0_xor1;
  wire [0:0] csa_component29_fa0_or0;
  wire [0:0] csa_component29_fa1_xor1;
  wire [0:0] csa_component29_fa1_or0;
  wire [0:0] csa_component29_fa2_xor1;
  wire [0:0] csa_component29_fa2_or0;
  wire [0:0] csa_component29_fa3_xor1;
  wire [0:0] csa_component29_fa3_or0;
  wire [0:0] csa_component29_fa4_xor1;
  wire [0:0] csa_component29_fa4_or0;
  wire [0:0] csa_component29_fa5_xor1;
  wire [0:0] csa_component29_fa5_or0;
  wire [0:0] csa_component29_fa6_xor1;
  wire [0:0] csa_component29_fa6_or0;
  wire [0:0] csa_component29_fa7_xor1;
  wire [0:0] csa_component29_fa7_or0;
  wire [0:0] csa_component29_fa8_xor1;
  wire [0:0] csa_component29_fa8_or0;
  wire [0:0] csa_component29_fa9_xor1;
  wire [0:0] csa_component29_fa9_or0;
  wire [0:0] csa_component29_fa10_xor1;
  wire [0:0] csa_component29_fa10_or0;
  wire [0:0] csa_component29_fa11_xor1;
  wire [0:0] csa_component29_fa11_or0;
  wire [0:0] csa_component29_fa12_xor1;
  wire [0:0] csa_component29_fa12_or0;
  wire [0:0] csa_component29_fa13_xor1;
  wire [0:0] csa_component29_fa13_or0;
  wire [0:0] csa_component29_fa14_xor1;
  wire [0:0] csa_component29_fa14_or0;
  wire [0:0] csa_component29_fa15_xor1;
  wire [0:0] csa_component29_fa15_or0;
  wire [0:0] csa_component29_fa16_xor1;
  wire [0:0] csa_component29_fa16_or0;
  wire [0:0] csa_component29_fa17_xor1;
  wire [0:0] csa_component29_fa17_or0;
  wire [0:0] csa_component29_fa18_xor1;
  wire [0:0] csa_component29_fa18_or0;
  wire [0:0] csa_component29_fa19_xor1;
  wire [0:0] csa_component29_fa19_or0;
  wire [0:0] csa_component29_fa20_xor1;
  wire [0:0] csa_component29_fa20_or0;
  wire [0:0] csa_component29_fa21_xor1;
  wire [0:0] csa_component29_fa21_or0;
  wire [0:0] csa_component29_fa22_xor1;
  wire [0:0] csa_component29_fa22_or0;
  wire [0:0] csa_component29_fa23_xor1;
  wire [0:0] csa_component29_fa23_or0;
  wire [0:0] csa_component29_fa24_xor1;
  wire [0:0] csa_component29_fa24_or0;
  wire [0:0] csa_component29_fa25_xor1;
  wire [0:0] csa_component29_fa25_or0;
  wire [0:0] csa_component29_fa26_xor1;
  wire [0:0] csa_component29_fa26_or0;
  wire [0:0] csa_component29_fa27_xor1;
  wire [0:0] csa_component29_fa27_or0;
  wire [0:0] csa_component29_fa28_xor1;
  wire [0:0] csa_component29_fa28_or0;

  fa fa_csa_component29_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component29_fa0_xor1), .fa_or0(csa_component29_fa0_or0));
  fa fa_csa_component29_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component29_fa1_xor1), .fa_or0(csa_component29_fa1_or0));
  fa fa_csa_component29_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component29_fa2_xor1), .fa_or0(csa_component29_fa2_or0));
  fa fa_csa_component29_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component29_fa3_xor1), .fa_or0(csa_component29_fa3_or0));
  fa fa_csa_component29_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component29_fa4_xor1), .fa_or0(csa_component29_fa4_or0));
  fa fa_csa_component29_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component29_fa5_xor1), .fa_or0(csa_component29_fa5_or0));
  fa fa_csa_component29_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component29_fa6_xor1), .fa_or0(csa_component29_fa6_or0));
  fa fa_csa_component29_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component29_fa7_xor1), .fa_or0(csa_component29_fa7_or0));
  fa fa_csa_component29_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component29_fa8_xor1), .fa_or0(csa_component29_fa8_or0));
  fa fa_csa_component29_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component29_fa9_xor1), .fa_or0(csa_component29_fa9_or0));
  fa fa_csa_component29_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component29_fa10_xor1), .fa_or0(csa_component29_fa10_or0));
  fa fa_csa_component29_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component29_fa11_xor1), .fa_or0(csa_component29_fa11_or0));
  fa fa_csa_component29_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component29_fa12_xor1), .fa_or0(csa_component29_fa12_or0));
  fa fa_csa_component29_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component29_fa13_xor1), .fa_or0(csa_component29_fa13_or0));
  fa fa_csa_component29_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component29_fa14_xor1), .fa_or0(csa_component29_fa14_or0));
  fa fa_csa_component29_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component29_fa15_xor1), .fa_or0(csa_component29_fa15_or0));
  fa fa_csa_component29_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component29_fa16_xor1), .fa_or0(csa_component29_fa16_or0));
  fa fa_csa_component29_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component29_fa17_xor1), .fa_or0(csa_component29_fa17_or0));
  fa fa_csa_component29_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component29_fa18_xor1), .fa_or0(csa_component29_fa18_or0));
  fa fa_csa_component29_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component29_fa19_xor1), .fa_or0(csa_component29_fa19_or0));
  fa fa_csa_component29_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component29_fa20_xor1), .fa_or0(csa_component29_fa20_or0));
  fa fa_csa_component29_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component29_fa21_xor1), .fa_or0(csa_component29_fa21_or0));
  fa fa_csa_component29_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component29_fa22_xor1), .fa_or0(csa_component29_fa22_or0));
  fa fa_csa_component29_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component29_fa23_xor1), .fa_or0(csa_component29_fa23_or0));
  fa fa_csa_component29_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component29_fa24_xor1), .fa_or0(csa_component29_fa24_or0));
  fa fa_csa_component29_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component29_fa25_xor1), .fa_or0(csa_component29_fa25_or0));
  fa fa_csa_component29_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component29_fa26_xor1), .fa_or0(csa_component29_fa26_or0));
  fa fa_csa_component29_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component29_fa27_xor1), .fa_or0(csa_component29_fa27_or0));
  fa fa_csa_component29_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component29_fa28_xor1), .fa_or0(csa_component29_fa28_or0));

  assign csa_component29_out[0] = csa_component29_fa0_xor1[0];
  assign csa_component29_out[1] = csa_component29_fa1_xor1[0];
  assign csa_component29_out[2] = csa_component29_fa2_xor1[0];
  assign csa_component29_out[3] = csa_component29_fa3_xor1[0];
  assign csa_component29_out[4] = csa_component29_fa4_xor1[0];
  assign csa_component29_out[5] = csa_component29_fa5_xor1[0];
  assign csa_component29_out[6] = csa_component29_fa6_xor1[0];
  assign csa_component29_out[7] = csa_component29_fa7_xor1[0];
  assign csa_component29_out[8] = csa_component29_fa8_xor1[0];
  assign csa_component29_out[9] = csa_component29_fa9_xor1[0];
  assign csa_component29_out[10] = csa_component29_fa10_xor1[0];
  assign csa_component29_out[11] = csa_component29_fa11_xor1[0];
  assign csa_component29_out[12] = csa_component29_fa12_xor1[0];
  assign csa_component29_out[13] = csa_component29_fa13_xor1[0];
  assign csa_component29_out[14] = csa_component29_fa14_xor1[0];
  assign csa_component29_out[15] = csa_component29_fa15_xor1[0];
  assign csa_component29_out[16] = csa_component29_fa16_xor1[0];
  assign csa_component29_out[17] = csa_component29_fa17_xor1[0];
  assign csa_component29_out[18] = csa_component29_fa18_xor1[0];
  assign csa_component29_out[19] = csa_component29_fa19_xor1[0];
  assign csa_component29_out[20] = csa_component29_fa20_xor1[0];
  assign csa_component29_out[21] = csa_component29_fa21_xor1[0];
  assign csa_component29_out[22] = csa_component29_fa22_xor1[0];
  assign csa_component29_out[23] = csa_component29_fa23_xor1[0];
  assign csa_component29_out[24] = csa_component29_fa24_xor1[0];
  assign csa_component29_out[25] = csa_component29_fa25_xor1[0];
  assign csa_component29_out[26] = csa_component29_fa26_xor1[0];
  assign csa_component29_out[27] = csa_component29_fa27_xor1[0];
  assign csa_component29_out[28] = csa_component29_fa28_xor1[0];
  assign csa_component29_out[29] = 1'b0;
  assign csa_component29_out[30] = 1'b0;
  assign csa_component29_out[31] = csa_component29_fa0_or0[0];
  assign csa_component29_out[32] = csa_component29_fa1_or0[0];
  assign csa_component29_out[33] = csa_component29_fa2_or0[0];
  assign csa_component29_out[34] = csa_component29_fa3_or0[0];
  assign csa_component29_out[35] = csa_component29_fa4_or0[0];
  assign csa_component29_out[36] = csa_component29_fa5_or0[0];
  assign csa_component29_out[37] = csa_component29_fa6_or0[0];
  assign csa_component29_out[38] = csa_component29_fa7_or0[0];
  assign csa_component29_out[39] = csa_component29_fa8_or0[0];
  assign csa_component29_out[40] = csa_component29_fa9_or0[0];
  assign csa_component29_out[41] = csa_component29_fa10_or0[0];
  assign csa_component29_out[42] = csa_component29_fa11_or0[0];
  assign csa_component29_out[43] = csa_component29_fa12_or0[0];
  assign csa_component29_out[44] = csa_component29_fa13_or0[0];
  assign csa_component29_out[45] = csa_component29_fa14_or0[0];
  assign csa_component29_out[46] = csa_component29_fa15_or0[0];
  assign csa_component29_out[47] = csa_component29_fa16_or0[0];
  assign csa_component29_out[48] = csa_component29_fa17_or0[0];
  assign csa_component29_out[49] = csa_component29_fa18_or0[0];
  assign csa_component29_out[50] = csa_component29_fa19_or0[0];
  assign csa_component29_out[51] = csa_component29_fa20_or0[0];
  assign csa_component29_out[52] = csa_component29_fa21_or0[0];
  assign csa_component29_out[53] = csa_component29_fa22_or0[0];
  assign csa_component29_out[54] = csa_component29_fa23_or0[0];
  assign csa_component29_out[55] = csa_component29_fa24_or0[0];
  assign csa_component29_out[56] = csa_component29_fa25_or0[0];
  assign csa_component29_out[57] = csa_component29_fa26_or0[0];
  assign csa_component29_out[58] = csa_component29_fa27_or0[0];
  assign csa_component29_out[59] = csa_component29_fa28_or0[0];
endmodule

module csa_component32(input [31:0] a, input [31:0] b, input [31:0] c, output [65:0] csa_component32_out);
  wire [0:0] csa_component32_fa0_xor1;
  wire [0:0] csa_component32_fa0_or0;
  wire [0:0] csa_component32_fa1_xor1;
  wire [0:0] csa_component32_fa1_or0;
  wire [0:0] csa_component32_fa2_xor1;
  wire [0:0] csa_component32_fa2_or0;
  wire [0:0] csa_component32_fa3_xor1;
  wire [0:0] csa_component32_fa3_or0;
  wire [0:0] csa_component32_fa4_xor1;
  wire [0:0] csa_component32_fa4_or0;
  wire [0:0] csa_component32_fa5_xor1;
  wire [0:0] csa_component32_fa5_or0;
  wire [0:0] csa_component32_fa6_xor1;
  wire [0:0] csa_component32_fa6_or0;
  wire [0:0] csa_component32_fa7_xor1;
  wire [0:0] csa_component32_fa7_or0;
  wire [0:0] csa_component32_fa8_xor1;
  wire [0:0] csa_component32_fa8_or0;
  wire [0:0] csa_component32_fa9_xor1;
  wire [0:0] csa_component32_fa9_or0;
  wire [0:0] csa_component32_fa10_xor1;
  wire [0:0] csa_component32_fa10_or0;
  wire [0:0] csa_component32_fa11_xor1;
  wire [0:0] csa_component32_fa11_or0;
  wire [0:0] csa_component32_fa12_xor1;
  wire [0:0] csa_component32_fa12_or0;
  wire [0:0] csa_component32_fa13_xor1;
  wire [0:0] csa_component32_fa13_or0;
  wire [0:0] csa_component32_fa14_xor1;
  wire [0:0] csa_component32_fa14_or0;
  wire [0:0] csa_component32_fa15_xor1;
  wire [0:0] csa_component32_fa15_or0;
  wire [0:0] csa_component32_fa16_xor1;
  wire [0:0] csa_component32_fa16_or0;
  wire [0:0] csa_component32_fa17_xor1;
  wire [0:0] csa_component32_fa17_or0;
  wire [0:0] csa_component32_fa18_xor1;
  wire [0:0] csa_component32_fa18_or0;
  wire [0:0] csa_component32_fa19_xor1;
  wire [0:0] csa_component32_fa19_or0;
  wire [0:0] csa_component32_fa20_xor1;
  wire [0:0] csa_component32_fa20_or0;
  wire [0:0] csa_component32_fa21_xor1;
  wire [0:0] csa_component32_fa21_or0;
  wire [0:0] csa_component32_fa22_xor1;
  wire [0:0] csa_component32_fa22_or0;
  wire [0:0] csa_component32_fa23_xor1;
  wire [0:0] csa_component32_fa23_or0;
  wire [0:0] csa_component32_fa24_xor1;
  wire [0:0] csa_component32_fa24_or0;
  wire [0:0] csa_component32_fa25_xor1;
  wire [0:0] csa_component32_fa25_or0;
  wire [0:0] csa_component32_fa26_xor1;
  wire [0:0] csa_component32_fa26_or0;
  wire [0:0] csa_component32_fa27_xor1;
  wire [0:0] csa_component32_fa27_or0;
  wire [0:0] csa_component32_fa28_xor1;
  wire [0:0] csa_component32_fa28_or0;
  wire [0:0] csa_component32_fa29_xor1;
  wire [0:0] csa_component32_fa29_or0;
  wire [0:0] csa_component32_fa30_xor1;
  wire [0:0] csa_component32_fa30_or0;
  wire [0:0] csa_component32_fa31_xor1;
  wire [0:0] csa_component32_fa31_or0;

  fa fa_csa_component32_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component32_fa0_xor1), .fa_or0(csa_component32_fa0_or0));
  fa fa_csa_component32_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component32_fa1_xor1), .fa_or0(csa_component32_fa1_or0));
  fa fa_csa_component32_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component32_fa2_xor1), .fa_or0(csa_component32_fa2_or0));
  fa fa_csa_component32_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component32_fa3_xor1), .fa_or0(csa_component32_fa3_or0));
  fa fa_csa_component32_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component32_fa4_xor1), .fa_or0(csa_component32_fa4_or0));
  fa fa_csa_component32_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component32_fa5_xor1), .fa_or0(csa_component32_fa5_or0));
  fa fa_csa_component32_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component32_fa6_xor1), .fa_or0(csa_component32_fa6_or0));
  fa fa_csa_component32_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component32_fa7_xor1), .fa_or0(csa_component32_fa7_or0));
  fa fa_csa_component32_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component32_fa8_xor1), .fa_or0(csa_component32_fa8_or0));
  fa fa_csa_component32_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component32_fa9_xor1), .fa_or0(csa_component32_fa9_or0));
  fa fa_csa_component32_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component32_fa10_xor1), .fa_or0(csa_component32_fa10_or0));
  fa fa_csa_component32_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component32_fa11_xor1), .fa_or0(csa_component32_fa11_or0));
  fa fa_csa_component32_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component32_fa12_xor1), .fa_or0(csa_component32_fa12_or0));
  fa fa_csa_component32_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component32_fa13_xor1), .fa_or0(csa_component32_fa13_or0));
  fa fa_csa_component32_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component32_fa14_xor1), .fa_or0(csa_component32_fa14_or0));
  fa fa_csa_component32_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component32_fa15_xor1), .fa_or0(csa_component32_fa15_or0));
  fa fa_csa_component32_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component32_fa16_xor1), .fa_or0(csa_component32_fa16_or0));
  fa fa_csa_component32_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component32_fa17_xor1), .fa_or0(csa_component32_fa17_or0));
  fa fa_csa_component32_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component32_fa18_xor1), .fa_or0(csa_component32_fa18_or0));
  fa fa_csa_component32_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component32_fa19_xor1), .fa_or0(csa_component32_fa19_or0));
  fa fa_csa_component32_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component32_fa20_xor1), .fa_or0(csa_component32_fa20_or0));
  fa fa_csa_component32_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component32_fa21_xor1), .fa_or0(csa_component32_fa21_or0));
  fa fa_csa_component32_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component32_fa22_xor1), .fa_or0(csa_component32_fa22_or0));
  fa fa_csa_component32_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component32_fa23_xor1), .fa_or0(csa_component32_fa23_or0));
  fa fa_csa_component32_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component32_fa24_xor1), .fa_or0(csa_component32_fa24_or0));
  fa fa_csa_component32_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component32_fa25_xor1), .fa_or0(csa_component32_fa25_or0));
  fa fa_csa_component32_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component32_fa26_xor1), .fa_or0(csa_component32_fa26_or0));
  fa fa_csa_component32_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component32_fa27_xor1), .fa_or0(csa_component32_fa27_or0));
  fa fa_csa_component32_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component32_fa28_xor1), .fa_or0(csa_component32_fa28_or0));
  fa fa_csa_component32_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component32_fa29_xor1), .fa_or0(csa_component32_fa29_or0));
  fa fa_csa_component32_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component32_fa30_xor1), .fa_or0(csa_component32_fa30_or0));
  fa fa_csa_component32_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component32_fa31_xor1), .fa_or0(csa_component32_fa31_or0));

  assign csa_component32_out[0] = csa_component32_fa0_xor1[0];
  assign csa_component32_out[1] = csa_component32_fa1_xor1[0];
  assign csa_component32_out[2] = csa_component32_fa2_xor1[0];
  assign csa_component32_out[3] = csa_component32_fa3_xor1[0];
  assign csa_component32_out[4] = csa_component32_fa4_xor1[0];
  assign csa_component32_out[5] = csa_component32_fa5_xor1[0];
  assign csa_component32_out[6] = csa_component32_fa6_xor1[0];
  assign csa_component32_out[7] = csa_component32_fa7_xor1[0];
  assign csa_component32_out[8] = csa_component32_fa8_xor1[0];
  assign csa_component32_out[9] = csa_component32_fa9_xor1[0];
  assign csa_component32_out[10] = csa_component32_fa10_xor1[0];
  assign csa_component32_out[11] = csa_component32_fa11_xor1[0];
  assign csa_component32_out[12] = csa_component32_fa12_xor1[0];
  assign csa_component32_out[13] = csa_component32_fa13_xor1[0];
  assign csa_component32_out[14] = csa_component32_fa14_xor1[0];
  assign csa_component32_out[15] = csa_component32_fa15_xor1[0];
  assign csa_component32_out[16] = csa_component32_fa16_xor1[0];
  assign csa_component32_out[17] = csa_component32_fa17_xor1[0];
  assign csa_component32_out[18] = csa_component32_fa18_xor1[0];
  assign csa_component32_out[19] = csa_component32_fa19_xor1[0];
  assign csa_component32_out[20] = csa_component32_fa20_xor1[0];
  assign csa_component32_out[21] = csa_component32_fa21_xor1[0];
  assign csa_component32_out[22] = csa_component32_fa22_xor1[0];
  assign csa_component32_out[23] = csa_component32_fa23_xor1[0];
  assign csa_component32_out[24] = csa_component32_fa24_xor1[0];
  assign csa_component32_out[25] = csa_component32_fa25_xor1[0];
  assign csa_component32_out[26] = csa_component32_fa26_xor1[0];
  assign csa_component32_out[27] = csa_component32_fa27_xor1[0];
  assign csa_component32_out[28] = csa_component32_fa28_xor1[0];
  assign csa_component32_out[29] = csa_component32_fa29_xor1[0];
  assign csa_component32_out[30] = csa_component32_fa30_xor1[0];
  assign csa_component32_out[31] = csa_component32_fa31_xor1[0];
  assign csa_component32_out[32] = 1'b0;
  assign csa_component32_out[33] = 1'b0;
  assign csa_component32_out[34] = csa_component32_fa0_or0[0];
  assign csa_component32_out[35] = csa_component32_fa1_or0[0];
  assign csa_component32_out[36] = csa_component32_fa2_or0[0];
  assign csa_component32_out[37] = csa_component32_fa3_or0[0];
  assign csa_component32_out[38] = csa_component32_fa4_or0[0];
  assign csa_component32_out[39] = csa_component32_fa5_or0[0];
  assign csa_component32_out[40] = csa_component32_fa6_or0[0];
  assign csa_component32_out[41] = csa_component32_fa7_or0[0];
  assign csa_component32_out[42] = csa_component32_fa8_or0[0];
  assign csa_component32_out[43] = csa_component32_fa9_or0[0];
  assign csa_component32_out[44] = csa_component32_fa10_or0[0];
  assign csa_component32_out[45] = csa_component32_fa11_or0[0];
  assign csa_component32_out[46] = csa_component32_fa12_or0[0];
  assign csa_component32_out[47] = csa_component32_fa13_or0[0];
  assign csa_component32_out[48] = csa_component32_fa14_or0[0];
  assign csa_component32_out[49] = csa_component32_fa15_or0[0];
  assign csa_component32_out[50] = csa_component32_fa16_or0[0];
  assign csa_component32_out[51] = csa_component32_fa17_or0[0];
  assign csa_component32_out[52] = csa_component32_fa18_or0[0];
  assign csa_component32_out[53] = csa_component32_fa19_or0[0];
  assign csa_component32_out[54] = csa_component32_fa20_or0[0];
  assign csa_component32_out[55] = csa_component32_fa21_or0[0];
  assign csa_component32_out[56] = csa_component32_fa22_or0[0];
  assign csa_component32_out[57] = csa_component32_fa23_or0[0];
  assign csa_component32_out[58] = csa_component32_fa24_or0[0];
  assign csa_component32_out[59] = csa_component32_fa25_or0[0];
  assign csa_component32_out[60] = csa_component32_fa26_or0[0];
  assign csa_component32_out[61] = csa_component32_fa27_or0[0];
  assign csa_component32_out[62] = csa_component32_fa28_or0[0];
  assign csa_component32_out[63] = csa_component32_fa29_or0[0];
  assign csa_component32_out[64] = csa_component32_fa30_or0[0];
  assign csa_component32_out[65] = csa_component32_fa31_or0[0];
endmodule

module csa_component35(input [34:0] a, input [34:0] b, input [34:0] c, output [71:0] csa_component35_out);
  wire [0:0] csa_component35_fa0_xor1;
  wire [0:0] csa_component35_fa0_or0;
  wire [0:0] csa_component35_fa1_xor1;
  wire [0:0] csa_component35_fa1_or0;
  wire [0:0] csa_component35_fa2_xor1;
  wire [0:0] csa_component35_fa2_or0;
  wire [0:0] csa_component35_fa3_xor1;
  wire [0:0] csa_component35_fa3_or0;
  wire [0:0] csa_component35_fa4_xor1;
  wire [0:0] csa_component35_fa4_or0;
  wire [0:0] csa_component35_fa5_xor1;
  wire [0:0] csa_component35_fa5_or0;
  wire [0:0] csa_component35_fa6_xor1;
  wire [0:0] csa_component35_fa6_or0;
  wire [0:0] csa_component35_fa7_xor1;
  wire [0:0] csa_component35_fa7_or0;
  wire [0:0] csa_component35_fa8_xor1;
  wire [0:0] csa_component35_fa8_or0;
  wire [0:0] csa_component35_fa9_xor1;
  wire [0:0] csa_component35_fa9_or0;
  wire [0:0] csa_component35_fa10_xor1;
  wire [0:0] csa_component35_fa10_or0;
  wire [0:0] csa_component35_fa11_xor1;
  wire [0:0] csa_component35_fa11_or0;
  wire [0:0] csa_component35_fa12_xor1;
  wire [0:0] csa_component35_fa12_or0;
  wire [0:0] csa_component35_fa13_xor1;
  wire [0:0] csa_component35_fa13_or0;
  wire [0:0] csa_component35_fa14_xor1;
  wire [0:0] csa_component35_fa14_or0;
  wire [0:0] csa_component35_fa15_xor1;
  wire [0:0] csa_component35_fa15_or0;
  wire [0:0] csa_component35_fa16_xor1;
  wire [0:0] csa_component35_fa16_or0;
  wire [0:0] csa_component35_fa17_xor1;
  wire [0:0] csa_component35_fa17_or0;
  wire [0:0] csa_component35_fa18_xor1;
  wire [0:0] csa_component35_fa18_or0;
  wire [0:0] csa_component35_fa19_xor1;
  wire [0:0] csa_component35_fa19_or0;
  wire [0:0] csa_component35_fa20_xor1;
  wire [0:0] csa_component35_fa20_or0;
  wire [0:0] csa_component35_fa21_xor1;
  wire [0:0] csa_component35_fa21_or0;
  wire [0:0] csa_component35_fa22_xor1;
  wire [0:0] csa_component35_fa22_or0;
  wire [0:0] csa_component35_fa23_xor1;
  wire [0:0] csa_component35_fa23_or0;
  wire [0:0] csa_component35_fa24_xor1;
  wire [0:0] csa_component35_fa24_or0;
  wire [0:0] csa_component35_fa25_xor1;
  wire [0:0] csa_component35_fa25_or0;
  wire [0:0] csa_component35_fa26_xor1;
  wire [0:0] csa_component35_fa26_or0;
  wire [0:0] csa_component35_fa27_xor1;
  wire [0:0] csa_component35_fa27_or0;
  wire [0:0] csa_component35_fa28_xor1;
  wire [0:0] csa_component35_fa28_or0;
  wire [0:0] csa_component35_fa29_xor1;
  wire [0:0] csa_component35_fa29_or0;
  wire [0:0] csa_component35_fa30_xor1;
  wire [0:0] csa_component35_fa30_or0;
  wire [0:0] csa_component35_fa31_xor1;
  wire [0:0] csa_component35_fa31_or0;
  wire [0:0] csa_component35_fa32_xor1;
  wire [0:0] csa_component35_fa32_or0;
  wire [0:0] csa_component35_fa33_xor1;
  wire [0:0] csa_component35_fa33_or0;
  wire [0:0] csa_component35_fa34_xor1;
  wire [0:0] csa_component35_fa34_or0;

  fa fa_csa_component35_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component35_fa0_xor1), .fa_or0(csa_component35_fa0_or0));
  fa fa_csa_component35_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component35_fa1_xor1), .fa_or0(csa_component35_fa1_or0));
  fa fa_csa_component35_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component35_fa2_xor1), .fa_or0(csa_component35_fa2_or0));
  fa fa_csa_component35_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component35_fa3_xor1), .fa_or0(csa_component35_fa3_or0));
  fa fa_csa_component35_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component35_fa4_xor1), .fa_or0(csa_component35_fa4_or0));
  fa fa_csa_component35_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component35_fa5_xor1), .fa_or0(csa_component35_fa5_or0));
  fa fa_csa_component35_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component35_fa6_xor1), .fa_or0(csa_component35_fa6_or0));
  fa fa_csa_component35_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component35_fa7_xor1), .fa_or0(csa_component35_fa7_or0));
  fa fa_csa_component35_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component35_fa8_xor1), .fa_or0(csa_component35_fa8_or0));
  fa fa_csa_component35_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component35_fa9_xor1), .fa_or0(csa_component35_fa9_or0));
  fa fa_csa_component35_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component35_fa10_xor1), .fa_or0(csa_component35_fa10_or0));
  fa fa_csa_component35_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component35_fa11_xor1), .fa_or0(csa_component35_fa11_or0));
  fa fa_csa_component35_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component35_fa12_xor1), .fa_or0(csa_component35_fa12_or0));
  fa fa_csa_component35_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component35_fa13_xor1), .fa_or0(csa_component35_fa13_or0));
  fa fa_csa_component35_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component35_fa14_xor1), .fa_or0(csa_component35_fa14_or0));
  fa fa_csa_component35_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component35_fa15_xor1), .fa_or0(csa_component35_fa15_or0));
  fa fa_csa_component35_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component35_fa16_xor1), .fa_or0(csa_component35_fa16_or0));
  fa fa_csa_component35_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component35_fa17_xor1), .fa_or0(csa_component35_fa17_or0));
  fa fa_csa_component35_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component35_fa18_xor1), .fa_or0(csa_component35_fa18_or0));
  fa fa_csa_component35_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component35_fa19_xor1), .fa_or0(csa_component35_fa19_or0));
  fa fa_csa_component35_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component35_fa20_xor1), .fa_or0(csa_component35_fa20_or0));
  fa fa_csa_component35_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component35_fa21_xor1), .fa_or0(csa_component35_fa21_or0));
  fa fa_csa_component35_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component35_fa22_xor1), .fa_or0(csa_component35_fa22_or0));
  fa fa_csa_component35_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component35_fa23_xor1), .fa_or0(csa_component35_fa23_or0));
  fa fa_csa_component35_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component35_fa24_xor1), .fa_or0(csa_component35_fa24_or0));
  fa fa_csa_component35_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component35_fa25_xor1), .fa_or0(csa_component35_fa25_or0));
  fa fa_csa_component35_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component35_fa26_xor1), .fa_or0(csa_component35_fa26_or0));
  fa fa_csa_component35_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component35_fa27_xor1), .fa_or0(csa_component35_fa27_or0));
  fa fa_csa_component35_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component35_fa28_xor1), .fa_or0(csa_component35_fa28_or0));
  fa fa_csa_component35_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component35_fa29_xor1), .fa_or0(csa_component35_fa29_or0));
  fa fa_csa_component35_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component35_fa30_xor1), .fa_or0(csa_component35_fa30_or0));
  fa fa_csa_component35_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component35_fa31_xor1), .fa_or0(csa_component35_fa31_or0));
  fa fa_csa_component35_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component35_fa32_xor1), .fa_or0(csa_component35_fa32_or0));
  fa fa_csa_component35_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component35_fa33_xor1), .fa_or0(csa_component35_fa33_or0));
  fa fa_csa_component35_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component35_fa34_xor1), .fa_or0(csa_component35_fa34_or0));

  assign csa_component35_out[0] = csa_component35_fa0_xor1[0];
  assign csa_component35_out[1] = csa_component35_fa1_xor1[0];
  assign csa_component35_out[2] = csa_component35_fa2_xor1[0];
  assign csa_component35_out[3] = csa_component35_fa3_xor1[0];
  assign csa_component35_out[4] = csa_component35_fa4_xor1[0];
  assign csa_component35_out[5] = csa_component35_fa5_xor1[0];
  assign csa_component35_out[6] = csa_component35_fa6_xor1[0];
  assign csa_component35_out[7] = csa_component35_fa7_xor1[0];
  assign csa_component35_out[8] = csa_component35_fa8_xor1[0];
  assign csa_component35_out[9] = csa_component35_fa9_xor1[0];
  assign csa_component35_out[10] = csa_component35_fa10_xor1[0];
  assign csa_component35_out[11] = csa_component35_fa11_xor1[0];
  assign csa_component35_out[12] = csa_component35_fa12_xor1[0];
  assign csa_component35_out[13] = csa_component35_fa13_xor1[0];
  assign csa_component35_out[14] = csa_component35_fa14_xor1[0];
  assign csa_component35_out[15] = csa_component35_fa15_xor1[0];
  assign csa_component35_out[16] = csa_component35_fa16_xor1[0];
  assign csa_component35_out[17] = csa_component35_fa17_xor1[0];
  assign csa_component35_out[18] = csa_component35_fa18_xor1[0];
  assign csa_component35_out[19] = csa_component35_fa19_xor1[0];
  assign csa_component35_out[20] = csa_component35_fa20_xor1[0];
  assign csa_component35_out[21] = csa_component35_fa21_xor1[0];
  assign csa_component35_out[22] = csa_component35_fa22_xor1[0];
  assign csa_component35_out[23] = csa_component35_fa23_xor1[0];
  assign csa_component35_out[24] = csa_component35_fa24_xor1[0];
  assign csa_component35_out[25] = csa_component35_fa25_xor1[0];
  assign csa_component35_out[26] = csa_component35_fa26_xor1[0];
  assign csa_component35_out[27] = csa_component35_fa27_xor1[0];
  assign csa_component35_out[28] = csa_component35_fa28_xor1[0];
  assign csa_component35_out[29] = csa_component35_fa29_xor1[0];
  assign csa_component35_out[30] = csa_component35_fa30_xor1[0];
  assign csa_component35_out[31] = csa_component35_fa31_xor1[0];
  assign csa_component35_out[32] = csa_component35_fa32_xor1[0];
  assign csa_component35_out[33] = csa_component35_fa33_xor1[0];
  assign csa_component35_out[34] = csa_component35_fa34_xor1[0];
  assign csa_component35_out[35] = 1'b0;
  assign csa_component35_out[36] = 1'b0;
  assign csa_component35_out[37] = csa_component35_fa0_or0[0];
  assign csa_component35_out[38] = csa_component35_fa1_or0[0];
  assign csa_component35_out[39] = csa_component35_fa2_or0[0];
  assign csa_component35_out[40] = csa_component35_fa3_or0[0];
  assign csa_component35_out[41] = csa_component35_fa4_or0[0];
  assign csa_component35_out[42] = csa_component35_fa5_or0[0];
  assign csa_component35_out[43] = csa_component35_fa6_or0[0];
  assign csa_component35_out[44] = csa_component35_fa7_or0[0];
  assign csa_component35_out[45] = csa_component35_fa8_or0[0];
  assign csa_component35_out[46] = csa_component35_fa9_or0[0];
  assign csa_component35_out[47] = csa_component35_fa10_or0[0];
  assign csa_component35_out[48] = csa_component35_fa11_or0[0];
  assign csa_component35_out[49] = csa_component35_fa12_or0[0];
  assign csa_component35_out[50] = csa_component35_fa13_or0[0];
  assign csa_component35_out[51] = csa_component35_fa14_or0[0];
  assign csa_component35_out[52] = csa_component35_fa15_or0[0];
  assign csa_component35_out[53] = csa_component35_fa16_or0[0];
  assign csa_component35_out[54] = csa_component35_fa17_or0[0];
  assign csa_component35_out[55] = csa_component35_fa18_or0[0];
  assign csa_component35_out[56] = csa_component35_fa19_or0[0];
  assign csa_component35_out[57] = csa_component35_fa20_or0[0];
  assign csa_component35_out[58] = csa_component35_fa21_or0[0];
  assign csa_component35_out[59] = csa_component35_fa22_or0[0];
  assign csa_component35_out[60] = csa_component35_fa23_or0[0];
  assign csa_component35_out[61] = csa_component35_fa24_or0[0];
  assign csa_component35_out[62] = csa_component35_fa25_or0[0];
  assign csa_component35_out[63] = csa_component35_fa26_or0[0];
  assign csa_component35_out[64] = csa_component35_fa27_or0[0];
  assign csa_component35_out[65] = csa_component35_fa28_or0[0];
  assign csa_component35_out[66] = csa_component35_fa29_or0[0];
  assign csa_component35_out[67] = csa_component35_fa30_or0[0];
  assign csa_component35_out[68] = csa_component35_fa31_or0[0];
  assign csa_component35_out[69] = csa_component35_fa32_or0[0];
  assign csa_component35_out[70] = csa_component35_fa33_or0[0];
  assign csa_component35_out[71] = csa_component35_fa34_or0[0];
endmodule

module csa_component38(input [37:0] a, input [37:0] b, input [37:0] c, output [77:0] csa_component38_out);
  wire [0:0] csa_component38_fa0_xor1;
  wire [0:0] csa_component38_fa0_or0;
  wire [0:0] csa_component38_fa1_xor1;
  wire [0:0] csa_component38_fa1_or0;
  wire [0:0] csa_component38_fa2_xor1;
  wire [0:0] csa_component38_fa2_or0;
  wire [0:0] csa_component38_fa3_xor1;
  wire [0:0] csa_component38_fa3_or0;
  wire [0:0] csa_component38_fa4_xor1;
  wire [0:0] csa_component38_fa4_or0;
  wire [0:0] csa_component38_fa5_xor1;
  wire [0:0] csa_component38_fa5_or0;
  wire [0:0] csa_component38_fa6_xor1;
  wire [0:0] csa_component38_fa6_or0;
  wire [0:0] csa_component38_fa7_xor1;
  wire [0:0] csa_component38_fa7_or0;
  wire [0:0] csa_component38_fa8_xor1;
  wire [0:0] csa_component38_fa8_or0;
  wire [0:0] csa_component38_fa9_xor1;
  wire [0:0] csa_component38_fa9_or0;
  wire [0:0] csa_component38_fa10_xor1;
  wire [0:0] csa_component38_fa10_or0;
  wire [0:0] csa_component38_fa11_xor1;
  wire [0:0] csa_component38_fa11_or0;
  wire [0:0] csa_component38_fa12_xor1;
  wire [0:0] csa_component38_fa12_or0;
  wire [0:0] csa_component38_fa13_xor1;
  wire [0:0] csa_component38_fa13_or0;
  wire [0:0] csa_component38_fa14_xor1;
  wire [0:0] csa_component38_fa14_or0;
  wire [0:0] csa_component38_fa15_xor1;
  wire [0:0] csa_component38_fa15_or0;
  wire [0:0] csa_component38_fa16_xor1;
  wire [0:0] csa_component38_fa16_or0;
  wire [0:0] csa_component38_fa17_xor1;
  wire [0:0] csa_component38_fa17_or0;
  wire [0:0] csa_component38_fa18_xor1;
  wire [0:0] csa_component38_fa18_or0;
  wire [0:0] csa_component38_fa19_xor1;
  wire [0:0] csa_component38_fa19_or0;
  wire [0:0] csa_component38_fa20_xor1;
  wire [0:0] csa_component38_fa20_or0;
  wire [0:0] csa_component38_fa21_xor1;
  wire [0:0] csa_component38_fa21_or0;
  wire [0:0] csa_component38_fa22_xor1;
  wire [0:0] csa_component38_fa22_or0;
  wire [0:0] csa_component38_fa23_xor1;
  wire [0:0] csa_component38_fa23_or0;
  wire [0:0] csa_component38_fa24_xor1;
  wire [0:0] csa_component38_fa24_or0;
  wire [0:0] csa_component38_fa25_xor1;
  wire [0:0] csa_component38_fa25_or0;
  wire [0:0] csa_component38_fa26_xor1;
  wire [0:0] csa_component38_fa26_or0;
  wire [0:0] csa_component38_fa27_xor1;
  wire [0:0] csa_component38_fa27_or0;
  wire [0:0] csa_component38_fa28_xor1;
  wire [0:0] csa_component38_fa28_or0;
  wire [0:0] csa_component38_fa29_xor1;
  wire [0:0] csa_component38_fa29_or0;
  wire [0:0] csa_component38_fa30_xor1;
  wire [0:0] csa_component38_fa30_or0;
  wire [0:0] csa_component38_fa31_xor1;
  wire [0:0] csa_component38_fa31_or0;
  wire [0:0] csa_component38_fa32_xor1;
  wire [0:0] csa_component38_fa32_or0;
  wire [0:0] csa_component38_fa33_xor1;
  wire [0:0] csa_component38_fa33_or0;
  wire [0:0] csa_component38_fa34_xor1;
  wire [0:0] csa_component38_fa34_or0;
  wire [0:0] csa_component38_fa35_xor1;
  wire [0:0] csa_component38_fa35_or0;
  wire [0:0] csa_component38_fa36_xor1;
  wire [0:0] csa_component38_fa36_or0;
  wire [0:0] csa_component38_fa37_xor1;
  wire [0:0] csa_component38_fa37_or0;

  fa fa_csa_component38_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component38_fa0_xor1), .fa_or0(csa_component38_fa0_or0));
  fa fa_csa_component38_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component38_fa1_xor1), .fa_or0(csa_component38_fa1_or0));
  fa fa_csa_component38_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component38_fa2_xor1), .fa_or0(csa_component38_fa2_or0));
  fa fa_csa_component38_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component38_fa3_xor1), .fa_or0(csa_component38_fa3_or0));
  fa fa_csa_component38_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component38_fa4_xor1), .fa_or0(csa_component38_fa4_or0));
  fa fa_csa_component38_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component38_fa5_xor1), .fa_or0(csa_component38_fa5_or0));
  fa fa_csa_component38_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component38_fa6_xor1), .fa_or0(csa_component38_fa6_or0));
  fa fa_csa_component38_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component38_fa7_xor1), .fa_or0(csa_component38_fa7_or0));
  fa fa_csa_component38_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component38_fa8_xor1), .fa_or0(csa_component38_fa8_or0));
  fa fa_csa_component38_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component38_fa9_xor1), .fa_or0(csa_component38_fa9_or0));
  fa fa_csa_component38_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component38_fa10_xor1), .fa_or0(csa_component38_fa10_or0));
  fa fa_csa_component38_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component38_fa11_xor1), .fa_or0(csa_component38_fa11_or0));
  fa fa_csa_component38_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component38_fa12_xor1), .fa_or0(csa_component38_fa12_or0));
  fa fa_csa_component38_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component38_fa13_xor1), .fa_or0(csa_component38_fa13_or0));
  fa fa_csa_component38_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component38_fa14_xor1), .fa_or0(csa_component38_fa14_or0));
  fa fa_csa_component38_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component38_fa15_xor1), .fa_or0(csa_component38_fa15_or0));
  fa fa_csa_component38_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component38_fa16_xor1), .fa_or0(csa_component38_fa16_or0));
  fa fa_csa_component38_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component38_fa17_xor1), .fa_or0(csa_component38_fa17_or0));
  fa fa_csa_component38_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component38_fa18_xor1), .fa_or0(csa_component38_fa18_or0));
  fa fa_csa_component38_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component38_fa19_xor1), .fa_or0(csa_component38_fa19_or0));
  fa fa_csa_component38_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component38_fa20_xor1), .fa_or0(csa_component38_fa20_or0));
  fa fa_csa_component38_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component38_fa21_xor1), .fa_or0(csa_component38_fa21_or0));
  fa fa_csa_component38_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component38_fa22_xor1), .fa_or0(csa_component38_fa22_or0));
  fa fa_csa_component38_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component38_fa23_xor1), .fa_or0(csa_component38_fa23_or0));
  fa fa_csa_component38_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component38_fa24_xor1), .fa_or0(csa_component38_fa24_or0));
  fa fa_csa_component38_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component38_fa25_xor1), .fa_or0(csa_component38_fa25_or0));
  fa fa_csa_component38_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component38_fa26_xor1), .fa_or0(csa_component38_fa26_or0));
  fa fa_csa_component38_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component38_fa27_xor1), .fa_or0(csa_component38_fa27_or0));
  fa fa_csa_component38_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component38_fa28_xor1), .fa_or0(csa_component38_fa28_or0));
  fa fa_csa_component38_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component38_fa29_xor1), .fa_or0(csa_component38_fa29_or0));
  fa fa_csa_component38_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component38_fa30_xor1), .fa_or0(csa_component38_fa30_or0));
  fa fa_csa_component38_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component38_fa31_xor1), .fa_or0(csa_component38_fa31_or0));
  fa fa_csa_component38_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component38_fa32_xor1), .fa_or0(csa_component38_fa32_or0));
  fa fa_csa_component38_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component38_fa33_xor1), .fa_or0(csa_component38_fa33_or0));
  fa fa_csa_component38_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component38_fa34_xor1), .fa_or0(csa_component38_fa34_or0));
  fa fa_csa_component38_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component38_fa35_xor1), .fa_or0(csa_component38_fa35_or0));
  fa fa_csa_component38_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component38_fa36_xor1), .fa_or0(csa_component38_fa36_or0));
  fa fa_csa_component38_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component38_fa37_xor1), .fa_or0(csa_component38_fa37_or0));

  assign csa_component38_out[0] = csa_component38_fa0_xor1[0];
  assign csa_component38_out[1] = csa_component38_fa1_xor1[0];
  assign csa_component38_out[2] = csa_component38_fa2_xor1[0];
  assign csa_component38_out[3] = csa_component38_fa3_xor1[0];
  assign csa_component38_out[4] = csa_component38_fa4_xor1[0];
  assign csa_component38_out[5] = csa_component38_fa5_xor1[0];
  assign csa_component38_out[6] = csa_component38_fa6_xor1[0];
  assign csa_component38_out[7] = csa_component38_fa7_xor1[0];
  assign csa_component38_out[8] = csa_component38_fa8_xor1[0];
  assign csa_component38_out[9] = csa_component38_fa9_xor1[0];
  assign csa_component38_out[10] = csa_component38_fa10_xor1[0];
  assign csa_component38_out[11] = csa_component38_fa11_xor1[0];
  assign csa_component38_out[12] = csa_component38_fa12_xor1[0];
  assign csa_component38_out[13] = csa_component38_fa13_xor1[0];
  assign csa_component38_out[14] = csa_component38_fa14_xor1[0];
  assign csa_component38_out[15] = csa_component38_fa15_xor1[0];
  assign csa_component38_out[16] = csa_component38_fa16_xor1[0];
  assign csa_component38_out[17] = csa_component38_fa17_xor1[0];
  assign csa_component38_out[18] = csa_component38_fa18_xor1[0];
  assign csa_component38_out[19] = csa_component38_fa19_xor1[0];
  assign csa_component38_out[20] = csa_component38_fa20_xor1[0];
  assign csa_component38_out[21] = csa_component38_fa21_xor1[0];
  assign csa_component38_out[22] = csa_component38_fa22_xor1[0];
  assign csa_component38_out[23] = csa_component38_fa23_xor1[0];
  assign csa_component38_out[24] = csa_component38_fa24_xor1[0];
  assign csa_component38_out[25] = csa_component38_fa25_xor1[0];
  assign csa_component38_out[26] = csa_component38_fa26_xor1[0];
  assign csa_component38_out[27] = csa_component38_fa27_xor1[0];
  assign csa_component38_out[28] = csa_component38_fa28_xor1[0];
  assign csa_component38_out[29] = csa_component38_fa29_xor1[0];
  assign csa_component38_out[30] = csa_component38_fa30_xor1[0];
  assign csa_component38_out[31] = csa_component38_fa31_xor1[0];
  assign csa_component38_out[32] = csa_component38_fa32_xor1[0];
  assign csa_component38_out[33] = csa_component38_fa33_xor1[0];
  assign csa_component38_out[34] = csa_component38_fa34_xor1[0];
  assign csa_component38_out[35] = csa_component38_fa35_xor1[0];
  assign csa_component38_out[36] = csa_component38_fa36_xor1[0];
  assign csa_component38_out[37] = csa_component38_fa37_xor1[0];
  assign csa_component38_out[38] = 1'b0;
  assign csa_component38_out[39] = 1'b0;
  assign csa_component38_out[40] = csa_component38_fa0_or0[0];
  assign csa_component38_out[41] = csa_component38_fa1_or0[0];
  assign csa_component38_out[42] = csa_component38_fa2_or0[0];
  assign csa_component38_out[43] = csa_component38_fa3_or0[0];
  assign csa_component38_out[44] = csa_component38_fa4_or0[0];
  assign csa_component38_out[45] = csa_component38_fa5_or0[0];
  assign csa_component38_out[46] = csa_component38_fa6_or0[0];
  assign csa_component38_out[47] = csa_component38_fa7_or0[0];
  assign csa_component38_out[48] = csa_component38_fa8_or0[0];
  assign csa_component38_out[49] = csa_component38_fa9_or0[0];
  assign csa_component38_out[50] = csa_component38_fa10_or0[0];
  assign csa_component38_out[51] = csa_component38_fa11_or0[0];
  assign csa_component38_out[52] = csa_component38_fa12_or0[0];
  assign csa_component38_out[53] = csa_component38_fa13_or0[0];
  assign csa_component38_out[54] = csa_component38_fa14_or0[0];
  assign csa_component38_out[55] = csa_component38_fa15_or0[0];
  assign csa_component38_out[56] = csa_component38_fa16_or0[0];
  assign csa_component38_out[57] = csa_component38_fa17_or0[0];
  assign csa_component38_out[58] = csa_component38_fa18_or0[0];
  assign csa_component38_out[59] = csa_component38_fa19_or0[0];
  assign csa_component38_out[60] = csa_component38_fa20_or0[0];
  assign csa_component38_out[61] = csa_component38_fa21_or0[0];
  assign csa_component38_out[62] = csa_component38_fa22_or0[0];
  assign csa_component38_out[63] = csa_component38_fa23_or0[0];
  assign csa_component38_out[64] = csa_component38_fa24_or0[0];
  assign csa_component38_out[65] = csa_component38_fa25_or0[0];
  assign csa_component38_out[66] = csa_component38_fa26_or0[0];
  assign csa_component38_out[67] = csa_component38_fa27_or0[0];
  assign csa_component38_out[68] = csa_component38_fa28_or0[0];
  assign csa_component38_out[69] = csa_component38_fa29_or0[0];
  assign csa_component38_out[70] = csa_component38_fa30_or0[0];
  assign csa_component38_out[71] = csa_component38_fa31_or0[0];
  assign csa_component38_out[72] = csa_component38_fa32_or0[0];
  assign csa_component38_out[73] = csa_component38_fa33_or0[0];
  assign csa_component38_out[74] = csa_component38_fa34_or0[0];
  assign csa_component38_out[75] = csa_component38_fa35_or0[0];
  assign csa_component38_out[76] = csa_component38_fa36_or0[0];
  assign csa_component38_out[77] = csa_component38_fa37_or0[0];
endmodule

module csa_component41(input [40:0] a, input [40:0] b, input [40:0] c, output [83:0] csa_component41_out);
  wire [0:0] csa_component41_fa0_xor1;
  wire [0:0] csa_component41_fa0_or0;
  wire [0:0] csa_component41_fa1_xor1;
  wire [0:0] csa_component41_fa1_or0;
  wire [0:0] csa_component41_fa2_xor1;
  wire [0:0] csa_component41_fa2_or0;
  wire [0:0] csa_component41_fa3_xor1;
  wire [0:0] csa_component41_fa3_or0;
  wire [0:0] csa_component41_fa4_xor1;
  wire [0:0] csa_component41_fa4_or0;
  wire [0:0] csa_component41_fa5_xor1;
  wire [0:0] csa_component41_fa5_or0;
  wire [0:0] csa_component41_fa6_xor1;
  wire [0:0] csa_component41_fa6_or0;
  wire [0:0] csa_component41_fa7_xor1;
  wire [0:0] csa_component41_fa7_or0;
  wire [0:0] csa_component41_fa8_xor1;
  wire [0:0] csa_component41_fa8_or0;
  wire [0:0] csa_component41_fa9_xor1;
  wire [0:0] csa_component41_fa9_or0;
  wire [0:0] csa_component41_fa10_xor1;
  wire [0:0] csa_component41_fa10_or0;
  wire [0:0] csa_component41_fa11_xor1;
  wire [0:0] csa_component41_fa11_or0;
  wire [0:0] csa_component41_fa12_xor1;
  wire [0:0] csa_component41_fa12_or0;
  wire [0:0] csa_component41_fa13_xor1;
  wire [0:0] csa_component41_fa13_or0;
  wire [0:0] csa_component41_fa14_xor1;
  wire [0:0] csa_component41_fa14_or0;
  wire [0:0] csa_component41_fa15_xor1;
  wire [0:0] csa_component41_fa15_or0;
  wire [0:0] csa_component41_fa16_xor1;
  wire [0:0] csa_component41_fa16_or0;
  wire [0:0] csa_component41_fa17_xor1;
  wire [0:0] csa_component41_fa17_or0;
  wire [0:0] csa_component41_fa18_xor1;
  wire [0:0] csa_component41_fa18_or0;
  wire [0:0] csa_component41_fa19_xor1;
  wire [0:0] csa_component41_fa19_or0;
  wire [0:0] csa_component41_fa20_xor1;
  wire [0:0] csa_component41_fa20_or0;
  wire [0:0] csa_component41_fa21_xor1;
  wire [0:0] csa_component41_fa21_or0;
  wire [0:0] csa_component41_fa22_xor1;
  wire [0:0] csa_component41_fa22_or0;
  wire [0:0] csa_component41_fa23_xor1;
  wire [0:0] csa_component41_fa23_or0;
  wire [0:0] csa_component41_fa24_xor1;
  wire [0:0] csa_component41_fa24_or0;
  wire [0:0] csa_component41_fa25_xor1;
  wire [0:0] csa_component41_fa25_or0;
  wire [0:0] csa_component41_fa26_xor1;
  wire [0:0] csa_component41_fa26_or0;
  wire [0:0] csa_component41_fa27_xor1;
  wire [0:0] csa_component41_fa27_or0;
  wire [0:0] csa_component41_fa28_xor1;
  wire [0:0] csa_component41_fa28_or0;
  wire [0:0] csa_component41_fa29_xor1;
  wire [0:0] csa_component41_fa29_or0;
  wire [0:0] csa_component41_fa30_xor1;
  wire [0:0] csa_component41_fa30_or0;
  wire [0:0] csa_component41_fa31_xor1;
  wire [0:0] csa_component41_fa31_or0;
  wire [0:0] csa_component41_fa32_xor1;
  wire [0:0] csa_component41_fa32_or0;
  wire [0:0] csa_component41_fa33_xor1;
  wire [0:0] csa_component41_fa33_or0;
  wire [0:0] csa_component41_fa34_xor1;
  wire [0:0] csa_component41_fa34_or0;
  wire [0:0] csa_component41_fa35_xor1;
  wire [0:0] csa_component41_fa35_or0;
  wire [0:0] csa_component41_fa36_xor1;
  wire [0:0] csa_component41_fa36_or0;
  wire [0:0] csa_component41_fa37_xor1;
  wire [0:0] csa_component41_fa37_or0;
  wire [0:0] csa_component41_fa38_xor1;
  wire [0:0] csa_component41_fa38_or0;
  wire [0:0] csa_component41_fa39_xor1;
  wire [0:0] csa_component41_fa39_or0;
  wire [0:0] csa_component41_fa40_xor1;
  wire [0:0] csa_component41_fa40_or0;

  fa fa_csa_component41_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component41_fa0_xor1), .fa_or0(csa_component41_fa0_or0));
  fa fa_csa_component41_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component41_fa1_xor1), .fa_or0(csa_component41_fa1_or0));
  fa fa_csa_component41_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component41_fa2_xor1), .fa_or0(csa_component41_fa2_or0));
  fa fa_csa_component41_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component41_fa3_xor1), .fa_or0(csa_component41_fa3_or0));
  fa fa_csa_component41_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component41_fa4_xor1), .fa_or0(csa_component41_fa4_or0));
  fa fa_csa_component41_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component41_fa5_xor1), .fa_or0(csa_component41_fa5_or0));
  fa fa_csa_component41_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component41_fa6_xor1), .fa_or0(csa_component41_fa6_or0));
  fa fa_csa_component41_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component41_fa7_xor1), .fa_or0(csa_component41_fa7_or0));
  fa fa_csa_component41_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component41_fa8_xor1), .fa_or0(csa_component41_fa8_or0));
  fa fa_csa_component41_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component41_fa9_xor1), .fa_or0(csa_component41_fa9_or0));
  fa fa_csa_component41_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component41_fa10_xor1), .fa_or0(csa_component41_fa10_or0));
  fa fa_csa_component41_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component41_fa11_xor1), .fa_or0(csa_component41_fa11_or0));
  fa fa_csa_component41_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component41_fa12_xor1), .fa_or0(csa_component41_fa12_or0));
  fa fa_csa_component41_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component41_fa13_xor1), .fa_or0(csa_component41_fa13_or0));
  fa fa_csa_component41_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component41_fa14_xor1), .fa_or0(csa_component41_fa14_or0));
  fa fa_csa_component41_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component41_fa15_xor1), .fa_or0(csa_component41_fa15_or0));
  fa fa_csa_component41_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component41_fa16_xor1), .fa_or0(csa_component41_fa16_or0));
  fa fa_csa_component41_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component41_fa17_xor1), .fa_or0(csa_component41_fa17_or0));
  fa fa_csa_component41_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component41_fa18_xor1), .fa_or0(csa_component41_fa18_or0));
  fa fa_csa_component41_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component41_fa19_xor1), .fa_or0(csa_component41_fa19_or0));
  fa fa_csa_component41_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component41_fa20_xor1), .fa_or0(csa_component41_fa20_or0));
  fa fa_csa_component41_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component41_fa21_xor1), .fa_or0(csa_component41_fa21_or0));
  fa fa_csa_component41_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component41_fa22_xor1), .fa_or0(csa_component41_fa22_or0));
  fa fa_csa_component41_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component41_fa23_xor1), .fa_or0(csa_component41_fa23_or0));
  fa fa_csa_component41_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component41_fa24_xor1), .fa_or0(csa_component41_fa24_or0));
  fa fa_csa_component41_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component41_fa25_xor1), .fa_or0(csa_component41_fa25_or0));
  fa fa_csa_component41_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component41_fa26_xor1), .fa_or0(csa_component41_fa26_or0));
  fa fa_csa_component41_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component41_fa27_xor1), .fa_or0(csa_component41_fa27_or0));
  fa fa_csa_component41_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component41_fa28_xor1), .fa_or0(csa_component41_fa28_or0));
  fa fa_csa_component41_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component41_fa29_xor1), .fa_or0(csa_component41_fa29_or0));
  fa fa_csa_component41_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component41_fa30_xor1), .fa_or0(csa_component41_fa30_or0));
  fa fa_csa_component41_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component41_fa31_xor1), .fa_or0(csa_component41_fa31_or0));
  fa fa_csa_component41_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component41_fa32_xor1), .fa_or0(csa_component41_fa32_or0));
  fa fa_csa_component41_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component41_fa33_xor1), .fa_or0(csa_component41_fa33_or0));
  fa fa_csa_component41_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component41_fa34_xor1), .fa_or0(csa_component41_fa34_or0));
  fa fa_csa_component41_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component41_fa35_xor1), .fa_or0(csa_component41_fa35_or0));
  fa fa_csa_component41_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component41_fa36_xor1), .fa_or0(csa_component41_fa36_or0));
  fa fa_csa_component41_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component41_fa37_xor1), .fa_or0(csa_component41_fa37_or0));
  fa fa_csa_component41_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component41_fa38_xor1), .fa_or0(csa_component41_fa38_or0));
  fa fa_csa_component41_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component41_fa39_xor1), .fa_or0(csa_component41_fa39_or0));
  fa fa_csa_component41_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component41_fa40_xor1), .fa_or0(csa_component41_fa40_or0));

  assign csa_component41_out[0] = csa_component41_fa0_xor1[0];
  assign csa_component41_out[1] = csa_component41_fa1_xor1[0];
  assign csa_component41_out[2] = csa_component41_fa2_xor1[0];
  assign csa_component41_out[3] = csa_component41_fa3_xor1[0];
  assign csa_component41_out[4] = csa_component41_fa4_xor1[0];
  assign csa_component41_out[5] = csa_component41_fa5_xor1[0];
  assign csa_component41_out[6] = csa_component41_fa6_xor1[0];
  assign csa_component41_out[7] = csa_component41_fa7_xor1[0];
  assign csa_component41_out[8] = csa_component41_fa8_xor1[0];
  assign csa_component41_out[9] = csa_component41_fa9_xor1[0];
  assign csa_component41_out[10] = csa_component41_fa10_xor1[0];
  assign csa_component41_out[11] = csa_component41_fa11_xor1[0];
  assign csa_component41_out[12] = csa_component41_fa12_xor1[0];
  assign csa_component41_out[13] = csa_component41_fa13_xor1[0];
  assign csa_component41_out[14] = csa_component41_fa14_xor1[0];
  assign csa_component41_out[15] = csa_component41_fa15_xor1[0];
  assign csa_component41_out[16] = csa_component41_fa16_xor1[0];
  assign csa_component41_out[17] = csa_component41_fa17_xor1[0];
  assign csa_component41_out[18] = csa_component41_fa18_xor1[0];
  assign csa_component41_out[19] = csa_component41_fa19_xor1[0];
  assign csa_component41_out[20] = csa_component41_fa20_xor1[0];
  assign csa_component41_out[21] = csa_component41_fa21_xor1[0];
  assign csa_component41_out[22] = csa_component41_fa22_xor1[0];
  assign csa_component41_out[23] = csa_component41_fa23_xor1[0];
  assign csa_component41_out[24] = csa_component41_fa24_xor1[0];
  assign csa_component41_out[25] = csa_component41_fa25_xor1[0];
  assign csa_component41_out[26] = csa_component41_fa26_xor1[0];
  assign csa_component41_out[27] = csa_component41_fa27_xor1[0];
  assign csa_component41_out[28] = csa_component41_fa28_xor1[0];
  assign csa_component41_out[29] = csa_component41_fa29_xor1[0];
  assign csa_component41_out[30] = csa_component41_fa30_xor1[0];
  assign csa_component41_out[31] = csa_component41_fa31_xor1[0];
  assign csa_component41_out[32] = csa_component41_fa32_xor1[0];
  assign csa_component41_out[33] = csa_component41_fa33_xor1[0];
  assign csa_component41_out[34] = csa_component41_fa34_xor1[0];
  assign csa_component41_out[35] = csa_component41_fa35_xor1[0];
  assign csa_component41_out[36] = csa_component41_fa36_xor1[0];
  assign csa_component41_out[37] = csa_component41_fa37_xor1[0];
  assign csa_component41_out[38] = csa_component41_fa38_xor1[0];
  assign csa_component41_out[39] = csa_component41_fa39_xor1[0];
  assign csa_component41_out[40] = csa_component41_fa40_xor1[0];
  assign csa_component41_out[41] = 1'b0;
  assign csa_component41_out[42] = 1'b0;
  assign csa_component41_out[43] = csa_component41_fa0_or0[0];
  assign csa_component41_out[44] = csa_component41_fa1_or0[0];
  assign csa_component41_out[45] = csa_component41_fa2_or0[0];
  assign csa_component41_out[46] = csa_component41_fa3_or0[0];
  assign csa_component41_out[47] = csa_component41_fa4_or0[0];
  assign csa_component41_out[48] = csa_component41_fa5_or0[0];
  assign csa_component41_out[49] = csa_component41_fa6_or0[0];
  assign csa_component41_out[50] = csa_component41_fa7_or0[0];
  assign csa_component41_out[51] = csa_component41_fa8_or0[0];
  assign csa_component41_out[52] = csa_component41_fa9_or0[0];
  assign csa_component41_out[53] = csa_component41_fa10_or0[0];
  assign csa_component41_out[54] = csa_component41_fa11_or0[0];
  assign csa_component41_out[55] = csa_component41_fa12_or0[0];
  assign csa_component41_out[56] = csa_component41_fa13_or0[0];
  assign csa_component41_out[57] = csa_component41_fa14_or0[0];
  assign csa_component41_out[58] = csa_component41_fa15_or0[0];
  assign csa_component41_out[59] = csa_component41_fa16_or0[0];
  assign csa_component41_out[60] = csa_component41_fa17_or0[0];
  assign csa_component41_out[61] = csa_component41_fa18_or0[0];
  assign csa_component41_out[62] = csa_component41_fa19_or0[0];
  assign csa_component41_out[63] = csa_component41_fa20_or0[0];
  assign csa_component41_out[64] = csa_component41_fa21_or0[0];
  assign csa_component41_out[65] = csa_component41_fa22_or0[0];
  assign csa_component41_out[66] = csa_component41_fa23_or0[0];
  assign csa_component41_out[67] = csa_component41_fa24_or0[0];
  assign csa_component41_out[68] = csa_component41_fa25_or0[0];
  assign csa_component41_out[69] = csa_component41_fa26_or0[0];
  assign csa_component41_out[70] = csa_component41_fa27_or0[0];
  assign csa_component41_out[71] = csa_component41_fa28_or0[0];
  assign csa_component41_out[72] = csa_component41_fa29_or0[0];
  assign csa_component41_out[73] = csa_component41_fa30_or0[0];
  assign csa_component41_out[74] = csa_component41_fa31_or0[0];
  assign csa_component41_out[75] = csa_component41_fa32_or0[0];
  assign csa_component41_out[76] = csa_component41_fa33_or0[0];
  assign csa_component41_out[77] = csa_component41_fa34_or0[0];
  assign csa_component41_out[78] = csa_component41_fa35_or0[0];
  assign csa_component41_out[79] = csa_component41_fa36_or0[0];
  assign csa_component41_out[80] = csa_component41_fa37_or0[0];
  assign csa_component41_out[81] = csa_component41_fa38_or0[0];
  assign csa_component41_out[82] = csa_component41_fa39_or0[0];
  assign csa_component41_out[83] = csa_component41_fa40_or0[0];
endmodule

module csa_component44(input [43:0] a, input [43:0] b, input [43:0] c, output [89:0] csa_component44_out);
  wire [0:0] csa_component44_fa0_xor1;
  wire [0:0] csa_component44_fa0_or0;
  wire [0:0] csa_component44_fa1_xor1;
  wire [0:0] csa_component44_fa1_or0;
  wire [0:0] csa_component44_fa2_xor1;
  wire [0:0] csa_component44_fa2_or0;
  wire [0:0] csa_component44_fa3_xor1;
  wire [0:0] csa_component44_fa3_or0;
  wire [0:0] csa_component44_fa4_xor1;
  wire [0:0] csa_component44_fa4_or0;
  wire [0:0] csa_component44_fa5_xor1;
  wire [0:0] csa_component44_fa5_or0;
  wire [0:0] csa_component44_fa6_xor1;
  wire [0:0] csa_component44_fa6_or0;
  wire [0:0] csa_component44_fa7_xor1;
  wire [0:0] csa_component44_fa7_or0;
  wire [0:0] csa_component44_fa8_xor1;
  wire [0:0] csa_component44_fa8_or0;
  wire [0:0] csa_component44_fa9_xor1;
  wire [0:0] csa_component44_fa9_or0;
  wire [0:0] csa_component44_fa10_xor1;
  wire [0:0] csa_component44_fa10_or0;
  wire [0:0] csa_component44_fa11_xor1;
  wire [0:0] csa_component44_fa11_or0;
  wire [0:0] csa_component44_fa12_xor1;
  wire [0:0] csa_component44_fa12_or0;
  wire [0:0] csa_component44_fa13_xor1;
  wire [0:0] csa_component44_fa13_or0;
  wire [0:0] csa_component44_fa14_xor1;
  wire [0:0] csa_component44_fa14_or0;
  wire [0:0] csa_component44_fa15_xor1;
  wire [0:0] csa_component44_fa15_or0;
  wire [0:0] csa_component44_fa16_xor1;
  wire [0:0] csa_component44_fa16_or0;
  wire [0:0] csa_component44_fa17_xor1;
  wire [0:0] csa_component44_fa17_or0;
  wire [0:0] csa_component44_fa18_xor1;
  wire [0:0] csa_component44_fa18_or0;
  wire [0:0] csa_component44_fa19_xor1;
  wire [0:0] csa_component44_fa19_or0;
  wire [0:0] csa_component44_fa20_xor1;
  wire [0:0] csa_component44_fa20_or0;
  wire [0:0] csa_component44_fa21_xor1;
  wire [0:0] csa_component44_fa21_or0;
  wire [0:0] csa_component44_fa22_xor1;
  wire [0:0] csa_component44_fa22_or0;
  wire [0:0] csa_component44_fa23_xor1;
  wire [0:0] csa_component44_fa23_or0;
  wire [0:0] csa_component44_fa24_xor1;
  wire [0:0] csa_component44_fa24_or0;
  wire [0:0] csa_component44_fa25_xor1;
  wire [0:0] csa_component44_fa25_or0;
  wire [0:0] csa_component44_fa26_xor1;
  wire [0:0] csa_component44_fa26_or0;
  wire [0:0] csa_component44_fa27_xor1;
  wire [0:0] csa_component44_fa27_or0;
  wire [0:0] csa_component44_fa28_xor1;
  wire [0:0] csa_component44_fa28_or0;
  wire [0:0] csa_component44_fa29_xor1;
  wire [0:0] csa_component44_fa29_or0;
  wire [0:0] csa_component44_fa30_xor1;
  wire [0:0] csa_component44_fa30_or0;
  wire [0:0] csa_component44_fa31_xor1;
  wire [0:0] csa_component44_fa31_or0;
  wire [0:0] csa_component44_fa32_xor1;
  wire [0:0] csa_component44_fa32_or0;
  wire [0:0] csa_component44_fa33_xor1;
  wire [0:0] csa_component44_fa33_or0;
  wire [0:0] csa_component44_fa34_xor1;
  wire [0:0] csa_component44_fa34_or0;
  wire [0:0] csa_component44_fa35_xor1;
  wire [0:0] csa_component44_fa35_or0;
  wire [0:0] csa_component44_fa36_xor1;
  wire [0:0] csa_component44_fa36_or0;
  wire [0:0] csa_component44_fa37_xor1;
  wire [0:0] csa_component44_fa37_or0;
  wire [0:0] csa_component44_fa38_xor1;
  wire [0:0] csa_component44_fa38_or0;
  wire [0:0] csa_component44_fa39_xor1;
  wire [0:0] csa_component44_fa39_or0;
  wire [0:0] csa_component44_fa40_xor1;
  wire [0:0] csa_component44_fa40_or0;
  wire [0:0] csa_component44_fa41_xor1;
  wire [0:0] csa_component44_fa41_or0;
  wire [0:0] csa_component44_fa42_xor1;
  wire [0:0] csa_component44_fa42_or0;
  wire [0:0] csa_component44_fa43_xor1;
  wire [0:0] csa_component44_fa43_or0;

  fa fa_csa_component44_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component44_fa0_xor1), .fa_or0(csa_component44_fa0_or0));
  fa fa_csa_component44_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component44_fa1_xor1), .fa_or0(csa_component44_fa1_or0));
  fa fa_csa_component44_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component44_fa2_xor1), .fa_or0(csa_component44_fa2_or0));
  fa fa_csa_component44_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component44_fa3_xor1), .fa_or0(csa_component44_fa3_or0));
  fa fa_csa_component44_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component44_fa4_xor1), .fa_or0(csa_component44_fa4_or0));
  fa fa_csa_component44_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component44_fa5_xor1), .fa_or0(csa_component44_fa5_or0));
  fa fa_csa_component44_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component44_fa6_xor1), .fa_or0(csa_component44_fa6_or0));
  fa fa_csa_component44_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component44_fa7_xor1), .fa_or0(csa_component44_fa7_or0));
  fa fa_csa_component44_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component44_fa8_xor1), .fa_or0(csa_component44_fa8_or0));
  fa fa_csa_component44_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component44_fa9_xor1), .fa_or0(csa_component44_fa9_or0));
  fa fa_csa_component44_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component44_fa10_xor1), .fa_or0(csa_component44_fa10_or0));
  fa fa_csa_component44_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component44_fa11_xor1), .fa_or0(csa_component44_fa11_or0));
  fa fa_csa_component44_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component44_fa12_xor1), .fa_or0(csa_component44_fa12_or0));
  fa fa_csa_component44_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component44_fa13_xor1), .fa_or0(csa_component44_fa13_or0));
  fa fa_csa_component44_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component44_fa14_xor1), .fa_or0(csa_component44_fa14_or0));
  fa fa_csa_component44_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component44_fa15_xor1), .fa_or0(csa_component44_fa15_or0));
  fa fa_csa_component44_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component44_fa16_xor1), .fa_or0(csa_component44_fa16_or0));
  fa fa_csa_component44_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component44_fa17_xor1), .fa_or0(csa_component44_fa17_or0));
  fa fa_csa_component44_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component44_fa18_xor1), .fa_or0(csa_component44_fa18_or0));
  fa fa_csa_component44_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component44_fa19_xor1), .fa_or0(csa_component44_fa19_or0));
  fa fa_csa_component44_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component44_fa20_xor1), .fa_or0(csa_component44_fa20_or0));
  fa fa_csa_component44_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component44_fa21_xor1), .fa_or0(csa_component44_fa21_or0));
  fa fa_csa_component44_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component44_fa22_xor1), .fa_or0(csa_component44_fa22_or0));
  fa fa_csa_component44_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component44_fa23_xor1), .fa_or0(csa_component44_fa23_or0));
  fa fa_csa_component44_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component44_fa24_xor1), .fa_or0(csa_component44_fa24_or0));
  fa fa_csa_component44_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component44_fa25_xor1), .fa_or0(csa_component44_fa25_or0));
  fa fa_csa_component44_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component44_fa26_xor1), .fa_or0(csa_component44_fa26_or0));
  fa fa_csa_component44_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component44_fa27_xor1), .fa_or0(csa_component44_fa27_or0));
  fa fa_csa_component44_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component44_fa28_xor1), .fa_or0(csa_component44_fa28_or0));
  fa fa_csa_component44_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component44_fa29_xor1), .fa_or0(csa_component44_fa29_or0));
  fa fa_csa_component44_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component44_fa30_xor1), .fa_or0(csa_component44_fa30_or0));
  fa fa_csa_component44_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component44_fa31_xor1), .fa_or0(csa_component44_fa31_or0));
  fa fa_csa_component44_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component44_fa32_xor1), .fa_or0(csa_component44_fa32_or0));
  fa fa_csa_component44_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component44_fa33_xor1), .fa_or0(csa_component44_fa33_or0));
  fa fa_csa_component44_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component44_fa34_xor1), .fa_or0(csa_component44_fa34_or0));
  fa fa_csa_component44_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component44_fa35_xor1), .fa_or0(csa_component44_fa35_or0));
  fa fa_csa_component44_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component44_fa36_xor1), .fa_or0(csa_component44_fa36_or0));
  fa fa_csa_component44_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component44_fa37_xor1), .fa_or0(csa_component44_fa37_or0));
  fa fa_csa_component44_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component44_fa38_xor1), .fa_or0(csa_component44_fa38_or0));
  fa fa_csa_component44_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component44_fa39_xor1), .fa_or0(csa_component44_fa39_or0));
  fa fa_csa_component44_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component44_fa40_xor1), .fa_or0(csa_component44_fa40_or0));
  fa fa_csa_component44_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component44_fa41_xor1), .fa_or0(csa_component44_fa41_or0));
  fa fa_csa_component44_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component44_fa42_xor1), .fa_or0(csa_component44_fa42_or0));
  fa fa_csa_component44_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component44_fa43_xor1), .fa_or0(csa_component44_fa43_or0));

  assign csa_component44_out[0] = csa_component44_fa0_xor1[0];
  assign csa_component44_out[1] = csa_component44_fa1_xor1[0];
  assign csa_component44_out[2] = csa_component44_fa2_xor1[0];
  assign csa_component44_out[3] = csa_component44_fa3_xor1[0];
  assign csa_component44_out[4] = csa_component44_fa4_xor1[0];
  assign csa_component44_out[5] = csa_component44_fa5_xor1[0];
  assign csa_component44_out[6] = csa_component44_fa6_xor1[0];
  assign csa_component44_out[7] = csa_component44_fa7_xor1[0];
  assign csa_component44_out[8] = csa_component44_fa8_xor1[0];
  assign csa_component44_out[9] = csa_component44_fa9_xor1[0];
  assign csa_component44_out[10] = csa_component44_fa10_xor1[0];
  assign csa_component44_out[11] = csa_component44_fa11_xor1[0];
  assign csa_component44_out[12] = csa_component44_fa12_xor1[0];
  assign csa_component44_out[13] = csa_component44_fa13_xor1[0];
  assign csa_component44_out[14] = csa_component44_fa14_xor1[0];
  assign csa_component44_out[15] = csa_component44_fa15_xor1[0];
  assign csa_component44_out[16] = csa_component44_fa16_xor1[0];
  assign csa_component44_out[17] = csa_component44_fa17_xor1[0];
  assign csa_component44_out[18] = csa_component44_fa18_xor1[0];
  assign csa_component44_out[19] = csa_component44_fa19_xor1[0];
  assign csa_component44_out[20] = csa_component44_fa20_xor1[0];
  assign csa_component44_out[21] = csa_component44_fa21_xor1[0];
  assign csa_component44_out[22] = csa_component44_fa22_xor1[0];
  assign csa_component44_out[23] = csa_component44_fa23_xor1[0];
  assign csa_component44_out[24] = csa_component44_fa24_xor1[0];
  assign csa_component44_out[25] = csa_component44_fa25_xor1[0];
  assign csa_component44_out[26] = csa_component44_fa26_xor1[0];
  assign csa_component44_out[27] = csa_component44_fa27_xor1[0];
  assign csa_component44_out[28] = csa_component44_fa28_xor1[0];
  assign csa_component44_out[29] = csa_component44_fa29_xor1[0];
  assign csa_component44_out[30] = csa_component44_fa30_xor1[0];
  assign csa_component44_out[31] = csa_component44_fa31_xor1[0];
  assign csa_component44_out[32] = csa_component44_fa32_xor1[0];
  assign csa_component44_out[33] = csa_component44_fa33_xor1[0];
  assign csa_component44_out[34] = csa_component44_fa34_xor1[0];
  assign csa_component44_out[35] = csa_component44_fa35_xor1[0];
  assign csa_component44_out[36] = csa_component44_fa36_xor1[0];
  assign csa_component44_out[37] = csa_component44_fa37_xor1[0];
  assign csa_component44_out[38] = csa_component44_fa38_xor1[0];
  assign csa_component44_out[39] = csa_component44_fa39_xor1[0];
  assign csa_component44_out[40] = csa_component44_fa40_xor1[0];
  assign csa_component44_out[41] = csa_component44_fa41_xor1[0];
  assign csa_component44_out[42] = csa_component44_fa42_xor1[0];
  assign csa_component44_out[43] = csa_component44_fa43_xor1[0];
  assign csa_component44_out[44] = 1'b0;
  assign csa_component44_out[45] = 1'b0;
  assign csa_component44_out[46] = csa_component44_fa0_or0[0];
  assign csa_component44_out[47] = csa_component44_fa1_or0[0];
  assign csa_component44_out[48] = csa_component44_fa2_or0[0];
  assign csa_component44_out[49] = csa_component44_fa3_or0[0];
  assign csa_component44_out[50] = csa_component44_fa4_or0[0];
  assign csa_component44_out[51] = csa_component44_fa5_or0[0];
  assign csa_component44_out[52] = csa_component44_fa6_or0[0];
  assign csa_component44_out[53] = csa_component44_fa7_or0[0];
  assign csa_component44_out[54] = csa_component44_fa8_or0[0];
  assign csa_component44_out[55] = csa_component44_fa9_or0[0];
  assign csa_component44_out[56] = csa_component44_fa10_or0[0];
  assign csa_component44_out[57] = csa_component44_fa11_or0[0];
  assign csa_component44_out[58] = csa_component44_fa12_or0[0];
  assign csa_component44_out[59] = csa_component44_fa13_or0[0];
  assign csa_component44_out[60] = csa_component44_fa14_or0[0];
  assign csa_component44_out[61] = csa_component44_fa15_or0[0];
  assign csa_component44_out[62] = csa_component44_fa16_or0[0];
  assign csa_component44_out[63] = csa_component44_fa17_or0[0];
  assign csa_component44_out[64] = csa_component44_fa18_or0[0];
  assign csa_component44_out[65] = csa_component44_fa19_or0[0];
  assign csa_component44_out[66] = csa_component44_fa20_or0[0];
  assign csa_component44_out[67] = csa_component44_fa21_or0[0];
  assign csa_component44_out[68] = csa_component44_fa22_or0[0];
  assign csa_component44_out[69] = csa_component44_fa23_or0[0];
  assign csa_component44_out[70] = csa_component44_fa24_or0[0];
  assign csa_component44_out[71] = csa_component44_fa25_or0[0];
  assign csa_component44_out[72] = csa_component44_fa26_or0[0];
  assign csa_component44_out[73] = csa_component44_fa27_or0[0];
  assign csa_component44_out[74] = csa_component44_fa28_or0[0];
  assign csa_component44_out[75] = csa_component44_fa29_or0[0];
  assign csa_component44_out[76] = csa_component44_fa30_or0[0];
  assign csa_component44_out[77] = csa_component44_fa31_or0[0];
  assign csa_component44_out[78] = csa_component44_fa32_or0[0];
  assign csa_component44_out[79] = csa_component44_fa33_or0[0];
  assign csa_component44_out[80] = csa_component44_fa34_or0[0];
  assign csa_component44_out[81] = csa_component44_fa35_or0[0];
  assign csa_component44_out[82] = csa_component44_fa36_or0[0];
  assign csa_component44_out[83] = csa_component44_fa37_or0[0];
  assign csa_component44_out[84] = csa_component44_fa38_or0[0];
  assign csa_component44_out[85] = csa_component44_fa39_or0[0];
  assign csa_component44_out[86] = csa_component44_fa40_or0[0];
  assign csa_component44_out[87] = csa_component44_fa41_or0[0];
  assign csa_component44_out[88] = csa_component44_fa42_or0[0];
  assign csa_component44_out[89] = csa_component44_fa43_or0[0];
endmodule

module csa_component47(input [46:0] a, input [46:0] b, input [46:0] c, output [95:0] csa_component47_out);
  wire [0:0] csa_component47_fa0_xor1;
  wire [0:0] csa_component47_fa0_or0;
  wire [0:0] csa_component47_fa1_xor1;
  wire [0:0] csa_component47_fa1_or0;
  wire [0:0] csa_component47_fa2_xor1;
  wire [0:0] csa_component47_fa2_or0;
  wire [0:0] csa_component47_fa3_xor1;
  wire [0:0] csa_component47_fa3_or0;
  wire [0:0] csa_component47_fa4_xor1;
  wire [0:0] csa_component47_fa4_or0;
  wire [0:0] csa_component47_fa5_xor1;
  wire [0:0] csa_component47_fa5_or0;
  wire [0:0] csa_component47_fa6_xor1;
  wire [0:0] csa_component47_fa6_or0;
  wire [0:0] csa_component47_fa7_xor1;
  wire [0:0] csa_component47_fa7_or0;
  wire [0:0] csa_component47_fa8_xor1;
  wire [0:0] csa_component47_fa8_or0;
  wire [0:0] csa_component47_fa9_xor1;
  wire [0:0] csa_component47_fa9_or0;
  wire [0:0] csa_component47_fa10_xor1;
  wire [0:0] csa_component47_fa10_or0;
  wire [0:0] csa_component47_fa11_xor1;
  wire [0:0] csa_component47_fa11_or0;
  wire [0:0] csa_component47_fa12_xor1;
  wire [0:0] csa_component47_fa12_or0;
  wire [0:0] csa_component47_fa13_xor1;
  wire [0:0] csa_component47_fa13_or0;
  wire [0:0] csa_component47_fa14_xor1;
  wire [0:0] csa_component47_fa14_or0;
  wire [0:0] csa_component47_fa15_xor1;
  wire [0:0] csa_component47_fa15_or0;
  wire [0:0] csa_component47_fa16_xor1;
  wire [0:0] csa_component47_fa16_or0;
  wire [0:0] csa_component47_fa17_xor1;
  wire [0:0] csa_component47_fa17_or0;
  wire [0:0] csa_component47_fa18_xor1;
  wire [0:0] csa_component47_fa18_or0;
  wire [0:0] csa_component47_fa19_xor1;
  wire [0:0] csa_component47_fa19_or0;
  wire [0:0] csa_component47_fa20_xor1;
  wire [0:0] csa_component47_fa20_or0;
  wire [0:0] csa_component47_fa21_xor1;
  wire [0:0] csa_component47_fa21_or0;
  wire [0:0] csa_component47_fa22_xor1;
  wire [0:0] csa_component47_fa22_or0;
  wire [0:0] csa_component47_fa23_xor1;
  wire [0:0] csa_component47_fa23_or0;
  wire [0:0] csa_component47_fa24_xor1;
  wire [0:0] csa_component47_fa24_or0;
  wire [0:0] csa_component47_fa25_xor1;
  wire [0:0] csa_component47_fa25_or0;
  wire [0:0] csa_component47_fa26_xor1;
  wire [0:0] csa_component47_fa26_or0;
  wire [0:0] csa_component47_fa27_xor1;
  wire [0:0] csa_component47_fa27_or0;
  wire [0:0] csa_component47_fa28_xor1;
  wire [0:0] csa_component47_fa28_or0;
  wire [0:0] csa_component47_fa29_xor1;
  wire [0:0] csa_component47_fa29_or0;
  wire [0:0] csa_component47_fa30_xor1;
  wire [0:0] csa_component47_fa30_or0;
  wire [0:0] csa_component47_fa31_xor1;
  wire [0:0] csa_component47_fa31_or0;
  wire [0:0] csa_component47_fa32_xor1;
  wire [0:0] csa_component47_fa32_or0;
  wire [0:0] csa_component47_fa33_xor1;
  wire [0:0] csa_component47_fa33_or0;
  wire [0:0] csa_component47_fa34_xor1;
  wire [0:0] csa_component47_fa34_or0;
  wire [0:0] csa_component47_fa35_xor1;
  wire [0:0] csa_component47_fa35_or0;
  wire [0:0] csa_component47_fa36_xor1;
  wire [0:0] csa_component47_fa36_or0;
  wire [0:0] csa_component47_fa37_xor1;
  wire [0:0] csa_component47_fa37_or0;
  wire [0:0] csa_component47_fa38_xor1;
  wire [0:0] csa_component47_fa38_or0;
  wire [0:0] csa_component47_fa39_xor1;
  wire [0:0] csa_component47_fa39_or0;
  wire [0:0] csa_component47_fa40_xor1;
  wire [0:0] csa_component47_fa40_or0;
  wire [0:0] csa_component47_fa41_xor1;
  wire [0:0] csa_component47_fa41_or0;
  wire [0:0] csa_component47_fa42_xor1;
  wire [0:0] csa_component47_fa42_or0;
  wire [0:0] csa_component47_fa43_xor1;
  wire [0:0] csa_component47_fa43_or0;
  wire [0:0] csa_component47_fa44_xor1;
  wire [0:0] csa_component47_fa44_or0;
  wire [0:0] csa_component47_fa45_xor1;
  wire [0:0] csa_component47_fa45_or0;
  wire [0:0] csa_component47_fa46_xor1;
  wire [0:0] csa_component47_fa46_or0;

  fa fa_csa_component47_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component47_fa0_xor1), .fa_or0(csa_component47_fa0_or0));
  fa fa_csa_component47_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component47_fa1_xor1), .fa_or0(csa_component47_fa1_or0));
  fa fa_csa_component47_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component47_fa2_xor1), .fa_or0(csa_component47_fa2_or0));
  fa fa_csa_component47_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component47_fa3_xor1), .fa_or0(csa_component47_fa3_or0));
  fa fa_csa_component47_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component47_fa4_xor1), .fa_or0(csa_component47_fa4_or0));
  fa fa_csa_component47_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component47_fa5_xor1), .fa_or0(csa_component47_fa5_or0));
  fa fa_csa_component47_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component47_fa6_xor1), .fa_or0(csa_component47_fa6_or0));
  fa fa_csa_component47_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component47_fa7_xor1), .fa_or0(csa_component47_fa7_or0));
  fa fa_csa_component47_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component47_fa8_xor1), .fa_or0(csa_component47_fa8_or0));
  fa fa_csa_component47_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component47_fa9_xor1), .fa_or0(csa_component47_fa9_or0));
  fa fa_csa_component47_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component47_fa10_xor1), .fa_or0(csa_component47_fa10_or0));
  fa fa_csa_component47_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component47_fa11_xor1), .fa_or0(csa_component47_fa11_or0));
  fa fa_csa_component47_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component47_fa12_xor1), .fa_or0(csa_component47_fa12_or0));
  fa fa_csa_component47_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component47_fa13_xor1), .fa_or0(csa_component47_fa13_or0));
  fa fa_csa_component47_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component47_fa14_xor1), .fa_or0(csa_component47_fa14_or0));
  fa fa_csa_component47_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component47_fa15_xor1), .fa_or0(csa_component47_fa15_or0));
  fa fa_csa_component47_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component47_fa16_xor1), .fa_or0(csa_component47_fa16_or0));
  fa fa_csa_component47_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component47_fa17_xor1), .fa_or0(csa_component47_fa17_or0));
  fa fa_csa_component47_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component47_fa18_xor1), .fa_or0(csa_component47_fa18_or0));
  fa fa_csa_component47_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component47_fa19_xor1), .fa_or0(csa_component47_fa19_or0));
  fa fa_csa_component47_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component47_fa20_xor1), .fa_or0(csa_component47_fa20_or0));
  fa fa_csa_component47_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component47_fa21_xor1), .fa_or0(csa_component47_fa21_or0));
  fa fa_csa_component47_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component47_fa22_xor1), .fa_or0(csa_component47_fa22_or0));
  fa fa_csa_component47_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component47_fa23_xor1), .fa_or0(csa_component47_fa23_or0));
  fa fa_csa_component47_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component47_fa24_xor1), .fa_or0(csa_component47_fa24_or0));
  fa fa_csa_component47_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component47_fa25_xor1), .fa_or0(csa_component47_fa25_or0));
  fa fa_csa_component47_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component47_fa26_xor1), .fa_or0(csa_component47_fa26_or0));
  fa fa_csa_component47_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component47_fa27_xor1), .fa_or0(csa_component47_fa27_or0));
  fa fa_csa_component47_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component47_fa28_xor1), .fa_or0(csa_component47_fa28_or0));
  fa fa_csa_component47_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component47_fa29_xor1), .fa_or0(csa_component47_fa29_or0));
  fa fa_csa_component47_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component47_fa30_xor1), .fa_or0(csa_component47_fa30_or0));
  fa fa_csa_component47_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component47_fa31_xor1), .fa_or0(csa_component47_fa31_or0));
  fa fa_csa_component47_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component47_fa32_xor1), .fa_or0(csa_component47_fa32_or0));
  fa fa_csa_component47_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component47_fa33_xor1), .fa_or0(csa_component47_fa33_or0));
  fa fa_csa_component47_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component47_fa34_xor1), .fa_or0(csa_component47_fa34_or0));
  fa fa_csa_component47_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component47_fa35_xor1), .fa_or0(csa_component47_fa35_or0));
  fa fa_csa_component47_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component47_fa36_xor1), .fa_or0(csa_component47_fa36_or0));
  fa fa_csa_component47_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component47_fa37_xor1), .fa_or0(csa_component47_fa37_or0));
  fa fa_csa_component47_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component47_fa38_xor1), .fa_or0(csa_component47_fa38_or0));
  fa fa_csa_component47_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component47_fa39_xor1), .fa_or0(csa_component47_fa39_or0));
  fa fa_csa_component47_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component47_fa40_xor1), .fa_or0(csa_component47_fa40_or0));
  fa fa_csa_component47_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component47_fa41_xor1), .fa_or0(csa_component47_fa41_or0));
  fa fa_csa_component47_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component47_fa42_xor1), .fa_or0(csa_component47_fa42_or0));
  fa fa_csa_component47_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component47_fa43_xor1), .fa_or0(csa_component47_fa43_or0));
  fa fa_csa_component47_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component47_fa44_xor1), .fa_or0(csa_component47_fa44_or0));
  fa fa_csa_component47_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component47_fa45_xor1), .fa_or0(csa_component47_fa45_or0));
  fa fa_csa_component47_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component47_fa46_xor1), .fa_or0(csa_component47_fa46_or0));

  assign csa_component47_out[0] = csa_component47_fa0_xor1[0];
  assign csa_component47_out[1] = csa_component47_fa1_xor1[0];
  assign csa_component47_out[2] = csa_component47_fa2_xor1[0];
  assign csa_component47_out[3] = csa_component47_fa3_xor1[0];
  assign csa_component47_out[4] = csa_component47_fa4_xor1[0];
  assign csa_component47_out[5] = csa_component47_fa5_xor1[0];
  assign csa_component47_out[6] = csa_component47_fa6_xor1[0];
  assign csa_component47_out[7] = csa_component47_fa7_xor1[0];
  assign csa_component47_out[8] = csa_component47_fa8_xor1[0];
  assign csa_component47_out[9] = csa_component47_fa9_xor1[0];
  assign csa_component47_out[10] = csa_component47_fa10_xor1[0];
  assign csa_component47_out[11] = csa_component47_fa11_xor1[0];
  assign csa_component47_out[12] = csa_component47_fa12_xor1[0];
  assign csa_component47_out[13] = csa_component47_fa13_xor1[0];
  assign csa_component47_out[14] = csa_component47_fa14_xor1[0];
  assign csa_component47_out[15] = csa_component47_fa15_xor1[0];
  assign csa_component47_out[16] = csa_component47_fa16_xor1[0];
  assign csa_component47_out[17] = csa_component47_fa17_xor1[0];
  assign csa_component47_out[18] = csa_component47_fa18_xor1[0];
  assign csa_component47_out[19] = csa_component47_fa19_xor1[0];
  assign csa_component47_out[20] = csa_component47_fa20_xor1[0];
  assign csa_component47_out[21] = csa_component47_fa21_xor1[0];
  assign csa_component47_out[22] = csa_component47_fa22_xor1[0];
  assign csa_component47_out[23] = csa_component47_fa23_xor1[0];
  assign csa_component47_out[24] = csa_component47_fa24_xor1[0];
  assign csa_component47_out[25] = csa_component47_fa25_xor1[0];
  assign csa_component47_out[26] = csa_component47_fa26_xor1[0];
  assign csa_component47_out[27] = csa_component47_fa27_xor1[0];
  assign csa_component47_out[28] = csa_component47_fa28_xor1[0];
  assign csa_component47_out[29] = csa_component47_fa29_xor1[0];
  assign csa_component47_out[30] = csa_component47_fa30_xor1[0];
  assign csa_component47_out[31] = csa_component47_fa31_xor1[0];
  assign csa_component47_out[32] = csa_component47_fa32_xor1[0];
  assign csa_component47_out[33] = csa_component47_fa33_xor1[0];
  assign csa_component47_out[34] = csa_component47_fa34_xor1[0];
  assign csa_component47_out[35] = csa_component47_fa35_xor1[0];
  assign csa_component47_out[36] = csa_component47_fa36_xor1[0];
  assign csa_component47_out[37] = csa_component47_fa37_xor1[0];
  assign csa_component47_out[38] = csa_component47_fa38_xor1[0];
  assign csa_component47_out[39] = csa_component47_fa39_xor1[0];
  assign csa_component47_out[40] = csa_component47_fa40_xor1[0];
  assign csa_component47_out[41] = csa_component47_fa41_xor1[0];
  assign csa_component47_out[42] = csa_component47_fa42_xor1[0];
  assign csa_component47_out[43] = csa_component47_fa43_xor1[0];
  assign csa_component47_out[44] = csa_component47_fa44_xor1[0];
  assign csa_component47_out[45] = csa_component47_fa45_xor1[0];
  assign csa_component47_out[46] = csa_component47_fa46_xor1[0];
  assign csa_component47_out[47] = 1'b0;
  assign csa_component47_out[48] = 1'b0;
  assign csa_component47_out[49] = csa_component47_fa0_or0[0];
  assign csa_component47_out[50] = csa_component47_fa1_or0[0];
  assign csa_component47_out[51] = csa_component47_fa2_or0[0];
  assign csa_component47_out[52] = csa_component47_fa3_or0[0];
  assign csa_component47_out[53] = csa_component47_fa4_or0[0];
  assign csa_component47_out[54] = csa_component47_fa5_or0[0];
  assign csa_component47_out[55] = csa_component47_fa6_or0[0];
  assign csa_component47_out[56] = csa_component47_fa7_or0[0];
  assign csa_component47_out[57] = csa_component47_fa8_or0[0];
  assign csa_component47_out[58] = csa_component47_fa9_or0[0];
  assign csa_component47_out[59] = csa_component47_fa10_or0[0];
  assign csa_component47_out[60] = csa_component47_fa11_or0[0];
  assign csa_component47_out[61] = csa_component47_fa12_or0[0];
  assign csa_component47_out[62] = csa_component47_fa13_or0[0];
  assign csa_component47_out[63] = csa_component47_fa14_or0[0];
  assign csa_component47_out[64] = csa_component47_fa15_or0[0];
  assign csa_component47_out[65] = csa_component47_fa16_or0[0];
  assign csa_component47_out[66] = csa_component47_fa17_or0[0];
  assign csa_component47_out[67] = csa_component47_fa18_or0[0];
  assign csa_component47_out[68] = csa_component47_fa19_or0[0];
  assign csa_component47_out[69] = csa_component47_fa20_or0[0];
  assign csa_component47_out[70] = csa_component47_fa21_or0[0];
  assign csa_component47_out[71] = csa_component47_fa22_or0[0];
  assign csa_component47_out[72] = csa_component47_fa23_or0[0];
  assign csa_component47_out[73] = csa_component47_fa24_or0[0];
  assign csa_component47_out[74] = csa_component47_fa25_or0[0];
  assign csa_component47_out[75] = csa_component47_fa26_or0[0];
  assign csa_component47_out[76] = csa_component47_fa27_or0[0];
  assign csa_component47_out[77] = csa_component47_fa28_or0[0];
  assign csa_component47_out[78] = csa_component47_fa29_or0[0];
  assign csa_component47_out[79] = csa_component47_fa30_or0[0];
  assign csa_component47_out[80] = csa_component47_fa31_or0[0];
  assign csa_component47_out[81] = csa_component47_fa32_or0[0];
  assign csa_component47_out[82] = csa_component47_fa33_or0[0];
  assign csa_component47_out[83] = csa_component47_fa34_or0[0];
  assign csa_component47_out[84] = csa_component47_fa35_or0[0];
  assign csa_component47_out[85] = csa_component47_fa36_or0[0];
  assign csa_component47_out[86] = csa_component47_fa37_or0[0];
  assign csa_component47_out[87] = csa_component47_fa38_or0[0];
  assign csa_component47_out[88] = csa_component47_fa39_or0[0];
  assign csa_component47_out[89] = csa_component47_fa40_or0[0];
  assign csa_component47_out[90] = csa_component47_fa41_or0[0];
  assign csa_component47_out[91] = csa_component47_fa42_or0[0];
  assign csa_component47_out[92] = csa_component47_fa43_or0[0];
  assign csa_component47_out[93] = csa_component47_fa44_or0[0];
  assign csa_component47_out[94] = csa_component47_fa45_or0[0];
  assign csa_component47_out[95] = csa_component47_fa46_or0[0];
endmodule

module csa_component30(input [29:0] a, input [29:0] b, input [29:0] c, output [61:0] csa_component30_out);
  wire [0:0] csa_component30_fa0_xor1;
  wire [0:0] csa_component30_fa0_or0;
  wire [0:0] csa_component30_fa1_xor1;
  wire [0:0] csa_component30_fa1_or0;
  wire [0:0] csa_component30_fa2_xor1;
  wire [0:0] csa_component30_fa2_or0;
  wire [0:0] csa_component30_fa3_xor1;
  wire [0:0] csa_component30_fa3_or0;
  wire [0:0] csa_component30_fa4_xor1;
  wire [0:0] csa_component30_fa4_or0;
  wire [0:0] csa_component30_fa5_xor1;
  wire [0:0] csa_component30_fa5_or0;
  wire [0:0] csa_component30_fa6_xor1;
  wire [0:0] csa_component30_fa6_or0;
  wire [0:0] csa_component30_fa7_xor1;
  wire [0:0] csa_component30_fa7_or0;
  wire [0:0] csa_component30_fa8_xor1;
  wire [0:0] csa_component30_fa8_or0;
  wire [0:0] csa_component30_fa9_xor1;
  wire [0:0] csa_component30_fa9_or0;
  wire [0:0] csa_component30_fa10_xor1;
  wire [0:0] csa_component30_fa10_or0;
  wire [0:0] csa_component30_fa11_xor1;
  wire [0:0] csa_component30_fa11_or0;
  wire [0:0] csa_component30_fa12_xor1;
  wire [0:0] csa_component30_fa12_or0;
  wire [0:0] csa_component30_fa13_xor1;
  wire [0:0] csa_component30_fa13_or0;
  wire [0:0] csa_component30_fa14_xor1;
  wire [0:0] csa_component30_fa14_or0;
  wire [0:0] csa_component30_fa15_xor1;
  wire [0:0] csa_component30_fa15_or0;
  wire [0:0] csa_component30_fa16_xor1;
  wire [0:0] csa_component30_fa16_or0;
  wire [0:0] csa_component30_fa17_xor1;
  wire [0:0] csa_component30_fa17_or0;
  wire [0:0] csa_component30_fa18_xor1;
  wire [0:0] csa_component30_fa18_or0;
  wire [0:0] csa_component30_fa19_xor1;
  wire [0:0] csa_component30_fa19_or0;
  wire [0:0] csa_component30_fa20_xor1;
  wire [0:0] csa_component30_fa20_or0;
  wire [0:0] csa_component30_fa21_xor1;
  wire [0:0] csa_component30_fa21_or0;
  wire [0:0] csa_component30_fa22_xor1;
  wire [0:0] csa_component30_fa22_or0;
  wire [0:0] csa_component30_fa23_xor1;
  wire [0:0] csa_component30_fa23_or0;
  wire [0:0] csa_component30_fa24_xor1;
  wire [0:0] csa_component30_fa24_or0;
  wire [0:0] csa_component30_fa25_xor1;
  wire [0:0] csa_component30_fa25_or0;
  wire [0:0] csa_component30_fa26_xor1;
  wire [0:0] csa_component30_fa26_or0;
  wire [0:0] csa_component30_fa27_xor1;
  wire [0:0] csa_component30_fa27_or0;
  wire [0:0] csa_component30_fa28_xor1;
  wire [0:0] csa_component30_fa28_or0;
  wire [0:0] csa_component30_fa29_xor1;
  wire [0:0] csa_component30_fa29_or0;

  fa fa_csa_component30_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component30_fa0_xor1), .fa_or0(csa_component30_fa0_or0));
  fa fa_csa_component30_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component30_fa1_xor1), .fa_or0(csa_component30_fa1_or0));
  fa fa_csa_component30_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component30_fa2_xor1), .fa_or0(csa_component30_fa2_or0));
  fa fa_csa_component30_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component30_fa3_xor1), .fa_or0(csa_component30_fa3_or0));
  fa fa_csa_component30_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component30_fa4_xor1), .fa_or0(csa_component30_fa4_or0));
  fa fa_csa_component30_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component30_fa5_xor1), .fa_or0(csa_component30_fa5_or0));
  fa fa_csa_component30_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component30_fa6_xor1), .fa_or0(csa_component30_fa6_or0));
  fa fa_csa_component30_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component30_fa7_xor1), .fa_or0(csa_component30_fa7_or0));
  fa fa_csa_component30_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component30_fa8_xor1), .fa_or0(csa_component30_fa8_or0));
  fa fa_csa_component30_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component30_fa9_xor1), .fa_or0(csa_component30_fa9_or0));
  fa fa_csa_component30_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component30_fa10_xor1), .fa_or0(csa_component30_fa10_or0));
  fa fa_csa_component30_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component30_fa11_xor1), .fa_or0(csa_component30_fa11_or0));
  fa fa_csa_component30_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component30_fa12_xor1), .fa_or0(csa_component30_fa12_or0));
  fa fa_csa_component30_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component30_fa13_xor1), .fa_or0(csa_component30_fa13_or0));
  fa fa_csa_component30_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component30_fa14_xor1), .fa_or0(csa_component30_fa14_or0));
  fa fa_csa_component30_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component30_fa15_xor1), .fa_or0(csa_component30_fa15_or0));
  fa fa_csa_component30_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component30_fa16_xor1), .fa_or0(csa_component30_fa16_or0));
  fa fa_csa_component30_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component30_fa17_xor1), .fa_or0(csa_component30_fa17_or0));
  fa fa_csa_component30_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component30_fa18_xor1), .fa_or0(csa_component30_fa18_or0));
  fa fa_csa_component30_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component30_fa19_xor1), .fa_or0(csa_component30_fa19_or0));
  fa fa_csa_component30_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component30_fa20_xor1), .fa_or0(csa_component30_fa20_or0));
  fa fa_csa_component30_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component30_fa21_xor1), .fa_or0(csa_component30_fa21_or0));
  fa fa_csa_component30_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component30_fa22_xor1), .fa_or0(csa_component30_fa22_or0));
  fa fa_csa_component30_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component30_fa23_xor1), .fa_or0(csa_component30_fa23_or0));
  fa fa_csa_component30_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component30_fa24_xor1), .fa_or0(csa_component30_fa24_or0));
  fa fa_csa_component30_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component30_fa25_xor1), .fa_or0(csa_component30_fa25_or0));
  fa fa_csa_component30_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component30_fa26_xor1), .fa_or0(csa_component30_fa26_or0));
  fa fa_csa_component30_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component30_fa27_xor1), .fa_or0(csa_component30_fa27_or0));
  fa fa_csa_component30_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component30_fa28_xor1), .fa_or0(csa_component30_fa28_or0));
  fa fa_csa_component30_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component30_fa29_xor1), .fa_or0(csa_component30_fa29_or0));

  assign csa_component30_out[0] = csa_component30_fa0_xor1[0];
  assign csa_component30_out[1] = csa_component30_fa1_xor1[0];
  assign csa_component30_out[2] = csa_component30_fa2_xor1[0];
  assign csa_component30_out[3] = csa_component30_fa3_xor1[0];
  assign csa_component30_out[4] = csa_component30_fa4_xor1[0];
  assign csa_component30_out[5] = csa_component30_fa5_xor1[0];
  assign csa_component30_out[6] = csa_component30_fa6_xor1[0];
  assign csa_component30_out[7] = csa_component30_fa7_xor1[0];
  assign csa_component30_out[8] = csa_component30_fa8_xor1[0];
  assign csa_component30_out[9] = csa_component30_fa9_xor1[0];
  assign csa_component30_out[10] = csa_component30_fa10_xor1[0];
  assign csa_component30_out[11] = csa_component30_fa11_xor1[0];
  assign csa_component30_out[12] = csa_component30_fa12_xor1[0];
  assign csa_component30_out[13] = csa_component30_fa13_xor1[0];
  assign csa_component30_out[14] = csa_component30_fa14_xor1[0];
  assign csa_component30_out[15] = csa_component30_fa15_xor1[0];
  assign csa_component30_out[16] = csa_component30_fa16_xor1[0];
  assign csa_component30_out[17] = csa_component30_fa17_xor1[0];
  assign csa_component30_out[18] = csa_component30_fa18_xor1[0];
  assign csa_component30_out[19] = csa_component30_fa19_xor1[0];
  assign csa_component30_out[20] = csa_component30_fa20_xor1[0];
  assign csa_component30_out[21] = csa_component30_fa21_xor1[0];
  assign csa_component30_out[22] = csa_component30_fa22_xor1[0];
  assign csa_component30_out[23] = csa_component30_fa23_xor1[0];
  assign csa_component30_out[24] = csa_component30_fa24_xor1[0];
  assign csa_component30_out[25] = csa_component30_fa25_xor1[0];
  assign csa_component30_out[26] = csa_component30_fa26_xor1[0];
  assign csa_component30_out[27] = csa_component30_fa27_xor1[0];
  assign csa_component30_out[28] = csa_component30_fa28_xor1[0];
  assign csa_component30_out[29] = csa_component30_fa29_xor1[0];
  assign csa_component30_out[30] = 1'b0;
  assign csa_component30_out[31] = 1'b0;
  assign csa_component30_out[32] = csa_component30_fa0_or0[0];
  assign csa_component30_out[33] = csa_component30_fa1_or0[0];
  assign csa_component30_out[34] = csa_component30_fa2_or0[0];
  assign csa_component30_out[35] = csa_component30_fa3_or0[0];
  assign csa_component30_out[36] = csa_component30_fa4_or0[0];
  assign csa_component30_out[37] = csa_component30_fa5_or0[0];
  assign csa_component30_out[38] = csa_component30_fa6_or0[0];
  assign csa_component30_out[39] = csa_component30_fa7_or0[0];
  assign csa_component30_out[40] = csa_component30_fa8_or0[0];
  assign csa_component30_out[41] = csa_component30_fa9_or0[0];
  assign csa_component30_out[42] = csa_component30_fa10_or0[0];
  assign csa_component30_out[43] = csa_component30_fa11_or0[0];
  assign csa_component30_out[44] = csa_component30_fa12_or0[0];
  assign csa_component30_out[45] = csa_component30_fa13_or0[0];
  assign csa_component30_out[46] = csa_component30_fa14_or0[0];
  assign csa_component30_out[47] = csa_component30_fa15_or0[0];
  assign csa_component30_out[48] = csa_component30_fa16_or0[0];
  assign csa_component30_out[49] = csa_component30_fa17_or0[0];
  assign csa_component30_out[50] = csa_component30_fa18_or0[0];
  assign csa_component30_out[51] = csa_component30_fa19_or0[0];
  assign csa_component30_out[52] = csa_component30_fa20_or0[0];
  assign csa_component30_out[53] = csa_component30_fa21_or0[0];
  assign csa_component30_out[54] = csa_component30_fa22_or0[0];
  assign csa_component30_out[55] = csa_component30_fa23_or0[0];
  assign csa_component30_out[56] = csa_component30_fa24_or0[0];
  assign csa_component30_out[57] = csa_component30_fa25_or0[0];
  assign csa_component30_out[58] = csa_component30_fa26_or0[0];
  assign csa_component30_out[59] = csa_component30_fa27_or0[0];
  assign csa_component30_out[60] = csa_component30_fa28_or0[0];
  assign csa_component30_out[61] = csa_component30_fa29_or0[0];
endmodule

module csa_component33(input [32:0] a, input [32:0] b, input [32:0] c, output [67:0] csa_component33_out);
  wire [0:0] csa_component33_fa0_xor1;
  wire [0:0] csa_component33_fa0_or0;
  wire [0:0] csa_component33_fa1_xor1;
  wire [0:0] csa_component33_fa1_or0;
  wire [0:0] csa_component33_fa2_xor1;
  wire [0:0] csa_component33_fa2_or0;
  wire [0:0] csa_component33_fa3_xor1;
  wire [0:0] csa_component33_fa3_or0;
  wire [0:0] csa_component33_fa4_xor1;
  wire [0:0] csa_component33_fa4_or0;
  wire [0:0] csa_component33_fa5_xor1;
  wire [0:0] csa_component33_fa5_or0;
  wire [0:0] csa_component33_fa6_xor1;
  wire [0:0] csa_component33_fa6_or0;
  wire [0:0] csa_component33_fa7_xor1;
  wire [0:0] csa_component33_fa7_or0;
  wire [0:0] csa_component33_fa8_xor1;
  wire [0:0] csa_component33_fa8_or0;
  wire [0:0] csa_component33_fa9_xor1;
  wire [0:0] csa_component33_fa9_or0;
  wire [0:0] csa_component33_fa10_xor1;
  wire [0:0] csa_component33_fa10_or0;
  wire [0:0] csa_component33_fa11_xor1;
  wire [0:0] csa_component33_fa11_or0;
  wire [0:0] csa_component33_fa12_xor1;
  wire [0:0] csa_component33_fa12_or0;
  wire [0:0] csa_component33_fa13_xor1;
  wire [0:0] csa_component33_fa13_or0;
  wire [0:0] csa_component33_fa14_xor1;
  wire [0:0] csa_component33_fa14_or0;
  wire [0:0] csa_component33_fa15_xor1;
  wire [0:0] csa_component33_fa15_or0;
  wire [0:0] csa_component33_fa16_xor1;
  wire [0:0] csa_component33_fa16_or0;
  wire [0:0] csa_component33_fa17_xor1;
  wire [0:0] csa_component33_fa17_or0;
  wire [0:0] csa_component33_fa18_xor1;
  wire [0:0] csa_component33_fa18_or0;
  wire [0:0] csa_component33_fa19_xor1;
  wire [0:0] csa_component33_fa19_or0;
  wire [0:0] csa_component33_fa20_xor1;
  wire [0:0] csa_component33_fa20_or0;
  wire [0:0] csa_component33_fa21_xor1;
  wire [0:0] csa_component33_fa21_or0;
  wire [0:0] csa_component33_fa22_xor1;
  wire [0:0] csa_component33_fa22_or0;
  wire [0:0] csa_component33_fa23_xor1;
  wire [0:0] csa_component33_fa23_or0;
  wire [0:0] csa_component33_fa24_xor1;
  wire [0:0] csa_component33_fa24_or0;
  wire [0:0] csa_component33_fa25_xor1;
  wire [0:0] csa_component33_fa25_or0;
  wire [0:0] csa_component33_fa26_xor1;
  wire [0:0] csa_component33_fa26_or0;
  wire [0:0] csa_component33_fa27_xor1;
  wire [0:0] csa_component33_fa27_or0;
  wire [0:0] csa_component33_fa28_xor1;
  wire [0:0] csa_component33_fa28_or0;
  wire [0:0] csa_component33_fa29_xor1;
  wire [0:0] csa_component33_fa29_or0;
  wire [0:0] csa_component33_fa30_xor1;
  wire [0:0] csa_component33_fa30_or0;
  wire [0:0] csa_component33_fa31_xor1;
  wire [0:0] csa_component33_fa31_or0;
  wire [0:0] csa_component33_fa32_xor1;
  wire [0:0] csa_component33_fa32_or0;

  fa fa_csa_component33_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component33_fa0_xor1), .fa_or0(csa_component33_fa0_or0));
  fa fa_csa_component33_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component33_fa1_xor1), .fa_or0(csa_component33_fa1_or0));
  fa fa_csa_component33_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component33_fa2_xor1), .fa_or0(csa_component33_fa2_or0));
  fa fa_csa_component33_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component33_fa3_xor1), .fa_or0(csa_component33_fa3_or0));
  fa fa_csa_component33_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component33_fa4_xor1), .fa_or0(csa_component33_fa4_or0));
  fa fa_csa_component33_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component33_fa5_xor1), .fa_or0(csa_component33_fa5_or0));
  fa fa_csa_component33_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component33_fa6_xor1), .fa_or0(csa_component33_fa6_or0));
  fa fa_csa_component33_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component33_fa7_xor1), .fa_or0(csa_component33_fa7_or0));
  fa fa_csa_component33_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component33_fa8_xor1), .fa_or0(csa_component33_fa8_or0));
  fa fa_csa_component33_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component33_fa9_xor1), .fa_or0(csa_component33_fa9_or0));
  fa fa_csa_component33_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component33_fa10_xor1), .fa_or0(csa_component33_fa10_or0));
  fa fa_csa_component33_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component33_fa11_xor1), .fa_or0(csa_component33_fa11_or0));
  fa fa_csa_component33_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component33_fa12_xor1), .fa_or0(csa_component33_fa12_or0));
  fa fa_csa_component33_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component33_fa13_xor1), .fa_or0(csa_component33_fa13_or0));
  fa fa_csa_component33_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component33_fa14_xor1), .fa_or0(csa_component33_fa14_or0));
  fa fa_csa_component33_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component33_fa15_xor1), .fa_or0(csa_component33_fa15_or0));
  fa fa_csa_component33_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component33_fa16_xor1), .fa_or0(csa_component33_fa16_or0));
  fa fa_csa_component33_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component33_fa17_xor1), .fa_or0(csa_component33_fa17_or0));
  fa fa_csa_component33_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component33_fa18_xor1), .fa_or0(csa_component33_fa18_or0));
  fa fa_csa_component33_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component33_fa19_xor1), .fa_or0(csa_component33_fa19_or0));
  fa fa_csa_component33_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component33_fa20_xor1), .fa_or0(csa_component33_fa20_or0));
  fa fa_csa_component33_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component33_fa21_xor1), .fa_or0(csa_component33_fa21_or0));
  fa fa_csa_component33_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component33_fa22_xor1), .fa_or0(csa_component33_fa22_or0));
  fa fa_csa_component33_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component33_fa23_xor1), .fa_or0(csa_component33_fa23_or0));
  fa fa_csa_component33_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component33_fa24_xor1), .fa_or0(csa_component33_fa24_or0));
  fa fa_csa_component33_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component33_fa25_xor1), .fa_or0(csa_component33_fa25_or0));
  fa fa_csa_component33_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component33_fa26_xor1), .fa_or0(csa_component33_fa26_or0));
  fa fa_csa_component33_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component33_fa27_xor1), .fa_or0(csa_component33_fa27_or0));
  fa fa_csa_component33_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component33_fa28_xor1), .fa_or0(csa_component33_fa28_or0));
  fa fa_csa_component33_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component33_fa29_xor1), .fa_or0(csa_component33_fa29_or0));
  fa fa_csa_component33_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component33_fa30_xor1), .fa_or0(csa_component33_fa30_or0));
  fa fa_csa_component33_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component33_fa31_xor1), .fa_or0(csa_component33_fa31_or0));
  fa fa_csa_component33_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component33_fa32_xor1), .fa_or0(csa_component33_fa32_or0));

  assign csa_component33_out[0] = csa_component33_fa0_xor1[0];
  assign csa_component33_out[1] = csa_component33_fa1_xor1[0];
  assign csa_component33_out[2] = csa_component33_fa2_xor1[0];
  assign csa_component33_out[3] = csa_component33_fa3_xor1[0];
  assign csa_component33_out[4] = csa_component33_fa4_xor1[0];
  assign csa_component33_out[5] = csa_component33_fa5_xor1[0];
  assign csa_component33_out[6] = csa_component33_fa6_xor1[0];
  assign csa_component33_out[7] = csa_component33_fa7_xor1[0];
  assign csa_component33_out[8] = csa_component33_fa8_xor1[0];
  assign csa_component33_out[9] = csa_component33_fa9_xor1[0];
  assign csa_component33_out[10] = csa_component33_fa10_xor1[0];
  assign csa_component33_out[11] = csa_component33_fa11_xor1[0];
  assign csa_component33_out[12] = csa_component33_fa12_xor1[0];
  assign csa_component33_out[13] = csa_component33_fa13_xor1[0];
  assign csa_component33_out[14] = csa_component33_fa14_xor1[0];
  assign csa_component33_out[15] = csa_component33_fa15_xor1[0];
  assign csa_component33_out[16] = csa_component33_fa16_xor1[0];
  assign csa_component33_out[17] = csa_component33_fa17_xor1[0];
  assign csa_component33_out[18] = csa_component33_fa18_xor1[0];
  assign csa_component33_out[19] = csa_component33_fa19_xor1[0];
  assign csa_component33_out[20] = csa_component33_fa20_xor1[0];
  assign csa_component33_out[21] = csa_component33_fa21_xor1[0];
  assign csa_component33_out[22] = csa_component33_fa22_xor1[0];
  assign csa_component33_out[23] = csa_component33_fa23_xor1[0];
  assign csa_component33_out[24] = csa_component33_fa24_xor1[0];
  assign csa_component33_out[25] = csa_component33_fa25_xor1[0];
  assign csa_component33_out[26] = csa_component33_fa26_xor1[0];
  assign csa_component33_out[27] = csa_component33_fa27_xor1[0];
  assign csa_component33_out[28] = csa_component33_fa28_xor1[0];
  assign csa_component33_out[29] = csa_component33_fa29_xor1[0];
  assign csa_component33_out[30] = csa_component33_fa30_xor1[0];
  assign csa_component33_out[31] = csa_component33_fa31_xor1[0];
  assign csa_component33_out[32] = csa_component33_fa32_xor1[0];
  assign csa_component33_out[33] = 1'b0;
  assign csa_component33_out[34] = 1'b0;
  assign csa_component33_out[35] = csa_component33_fa0_or0[0];
  assign csa_component33_out[36] = csa_component33_fa1_or0[0];
  assign csa_component33_out[37] = csa_component33_fa2_or0[0];
  assign csa_component33_out[38] = csa_component33_fa3_or0[0];
  assign csa_component33_out[39] = csa_component33_fa4_or0[0];
  assign csa_component33_out[40] = csa_component33_fa5_or0[0];
  assign csa_component33_out[41] = csa_component33_fa6_or0[0];
  assign csa_component33_out[42] = csa_component33_fa7_or0[0];
  assign csa_component33_out[43] = csa_component33_fa8_or0[0];
  assign csa_component33_out[44] = csa_component33_fa9_or0[0];
  assign csa_component33_out[45] = csa_component33_fa10_or0[0];
  assign csa_component33_out[46] = csa_component33_fa11_or0[0];
  assign csa_component33_out[47] = csa_component33_fa12_or0[0];
  assign csa_component33_out[48] = csa_component33_fa13_or0[0];
  assign csa_component33_out[49] = csa_component33_fa14_or0[0];
  assign csa_component33_out[50] = csa_component33_fa15_or0[0];
  assign csa_component33_out[51] = csa_component33_fa16_or0[0];
  assign csa_component33_out[52] = csa_component33_fa17_or0[0];
  assign csa_component33_out[53] = csa_component33_fa18_or0[0];
  assign csa_component33_out[54] = csa_component33_fa19_or0[0];
  assign csa_component33_out[55] = csa_component33_fa20_or0[0];
  assign csa_component33_out[56] = csa_component33_fa21_or0[0];
  assign csa_component33_out[57] = csa_component33_fa22_or0[0];
  assign csa_component33_out[58] = csa_component33_fa23_or0[0];
  assign csa_component33_out[59] = csa_component33_fa24_or0[0];
  assign csa_component33_out[60] = csa_component33_fa25_or0[0];
  assign csa_component33_out[61] = csa_component33_fa26_or0[0];
  assign csa_component33_out[62] = csa_component33_fa27_or0[0];
  assign csa_component33_out[63] = csa_component33_fa28_or0[0];
  assign csa_component33_out[64] = csa_component33_fa29_or0[0];
  assign csa_component33_out[65] = csa_component33_fa30_or0[0];
  assign csa_component33_out[66] = csa_component33_fa31_or0[0];
  assign csa_component33_out[67] = csa_component33_fa32_or0[0];
endmodule

module csa_component39(input [38:0] a, input [38:0] b, input [38:0] c, output [79:0] csa_component39_out);
  wire [0:0] csa_component39_fa0_xor1;
  wire [0:0] csa_component39_fa0_or0;
  wire [0:0] csa_component39_fa1_xor1;
  wire [0:0] csa_component39_fa1_or0;
  wire [0:0] csa_component39_fa2_xor1;
  wire [0:0] csa_component39_fa2_or0;
  wire [0:0] csa_component39_fa3_xor1;
  wire [0:0] csa_component39_fa3_or0;
  wire [0:0] csa_component39_fa4_xor1;
  wire [0:0] csa_component39_fa4_or0;
  wire [0:0] csa_component39_fa5_xor1;
  wire [0:0] csa_component39_fa5_or0;
  wire [0:0] csa_component39_fa6_xor1;
  wire [0:0] csa_component39_fa6_or0;
  wire [0:0] csa_component39_fa7_xor1;
  wire [0:0] csa_component39_fa7_or0;
  wire [0:0] csa_component39_fa8_xor1;
  wire [0:0] csa_component39_fa8_or0;
  wire [0:0] csa_component39_fa9_xor1;
  wire [0:0] csa_component39_fa9_or0;
  wire [0:0] csa_component39_fa10_xor1;
  wire [0:0] csa_component39_fa10_or0;
  wire [0:0] csa_component39_fa11_xor1;
  wire [0:0] csa_component39_fa11_or0;
  wire [0:0] csa_component39_fa12_xor1;
  wire [0:0] csa_component39_fa12_or0;
  wire [0:0] csa_component39_fa13_xor1;
  wire [0:0] csa_component39_fa13_or0;
  wire [0:0] csa_component39_fa14_xor1;
  wire [0:0] csa_component39_fa14_or0;
  wire [0:0] csa_component39_fa15_xor1;
  wire [0:0] csa_component39_fa15_or0;
  wire [0:0] csa_component39_fa16_xor1;
  wire [0:0] csa_component39_fa16_or0;
  wire [0:0] csa_component39_fa17_xor1;
  wire [0:0] csa_component39_fa17_or0;
  wire [0:0] csa_component39_fa18_xor1;
  wire [0:0] csa_component39_fa18_or0;
  wire [0:0] csa_component39_fa19_xor1;
  wire [0:0] csa_component39_fa19_or0;
  wire [0:0] csa_component39_fa20_xor1;
  wire [0:0] csa_component39_fa20_or0;
  wire [0:0] csa_component39_fa21_xor1;
  wire [0:0] csa_component39_fa21_or0;
  wire [0:0] csa_component39_fa22_xor1;
  wire [0:0] csa_component39_fa22_or0;
  wire [0:0] csa_component39_fa23_xor1;
  wire [0:0] csa_component39_fa23_or0;
  wire [0:0] csa_component39_fa24_xor1;
  wire [0:0] csa_component39_fa24_or0;
  wire [0:0] csa_component39_fa25_xor1;
  wire [0:0] csa_component39_fa25_or0;
  wire [0:0] csa_component39_fa26_xor1;
  wire [0:0] csa_component39_fa26_or0;
  wire [0:0] csa_component39_fa27_xor1;
  wire [0:0] csa_component39_fa27_or0;
  wire [0:0] csa_component39_fa28_xor1;
  wire [0:0] csa_component39_fa28_or0;
  wire [0:0] csa_component39_fa29_xor1;
  wire [0:0] csa_component39_fa29_or0;
  wire [0:0] csa_component39_fa30_xor1;
  wire [0:0] csa_component39_fa30_or0;
  wire [0:0] csa_component39_fa31_xor1;
  wire [0:0] csa_component39_fa31_or0;
  wire [0:0] csa_component39_fa32_xor1;
  wire [0:0] csa_component39_fa32_or0;
  wire [0:0] csa_component39_fa33_xor1;
  wire [0:0] csa_component39_fa33_or0;
  wire [0:0] csa_component39_fa34_xor1;
  wire [0:0] csa_component39_fa34_or0;
  wire [0:0] csa_component39_fa35_xor1;
  wire [0:0] csa_component39_fa35_or0;
  wire [0:0] csa_component39_fa36_xor1;
  wire [0:0] csa_component39_fa36_or0;
  wire [0:0] csa_component39_fa37_xor1;
  wire [0:0] csa_component39_fa37_or0;
  wire [0:0] csa_component39_fa38_xor1;
  wire [0:0] csa_component39_fa38_or0;

  fa fa_csa_component39_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component39_fa0_xor1), .fa_or0(csa_component39_fa0_or0));
  fa fa_csa_component39_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component39_fa1_xor1), .fa_or0(csa_component39_fa1_or0));
  fa fa_csa_component39_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component39_fa2_xor1), .fa_or0(csa_component39_fa2_or0));
  fa fa_csa_component39_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component39_fa3_xor1), .fa_or0(csa_component39_fa3_or0));
  fa fa_csa_component39_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component39_fa4_xor1), .fa_or0(csa_component39_fa4_or0));
  fa fa_csa_component39_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component39_fa5_xor1), .fa_or0(csa_component39_fa5_or0));
  fa fa_csa_component39_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component39_fa6_xor1), .fa_or0(csa_component39_fa6_or0));
  fa fa_csa_component39_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component39_fa7_xor1), .fa_or0(csa_component39_fa7_or0));
  fa fa_csa_component39_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component39_fa8_xor1), .fa_or0(csa_component39_fa8_or0));
  fa fa_csa_component39_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component39_fa9_xor1), .fa_or0(csa_component39_fa9_or0));
  fa fa_csa_component39_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component39_fa10_xor1), .fa_or0(csa_component39_fa10_or0));
  fa fa_csa_component39_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component39_fa11_xor1), .fa_or0(csa_component39_fa11_or0));
  fa fa_csa_component39_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component39_fa12_xor1), .fa_or0(csa_component39_fa12_or0));
  fa fa_csa_component39_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component39_fa13_xor1), .fa_or0(csa_component39_fa13_or0));
  fa fa_csa_component39_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component39_fa14_xor1), .fa_or0(csa_component39_fa14_or0));
  fa fa_csa_component39_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component39_fa15_xor1), .fa_or0(csa_component39_fa15_or0));
  fa fa_csa_component39_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component39_fa16_xor1), .fa_or0(csa_component39_fa16_or0));
  fa fa_csa_component39_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component39_fa17_xor1), .fa_or0(csa_component39_fa17_or0));
  fa fa_csa_component39_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component39_fa18_xor1), .fa_or0(csa_component39_fa18_or0));
  fa fa_csa_component39_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component39_fa19_xor1), .fa_or0(csa_component39_fa19_or0));
  fa fa_csa_component39_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component39_fa20_xor1), .fa_or0(csa_component39_fa20_or0));
  fa fa_csa_component39_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component39_fa21_xor1), .fa_or0(csa_component39_fa21_or0));
  fa fa_csa_component39_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component39_fa22_xor1), .fa_or0(csa_component39_fa22_or0));
  fa fa_csa_component39_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component39_fa23_xor1), .fa_or0(csa_component39_fa23_or0));
  fa fa_csa_component39_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component39_fa24_xor1), .fa_or0(csa_component39_fa24_or0));
  fa fa_csa_component39_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component39_fa25_xor1), .fa_or0(csa_component39_fa25_or0));
  fa fa_csa_component39_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component39_fa26_xor1), .fa_or0(csa_component39_fa26_or0));
  fa fa_csa_component39_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component39_fa27_xor1), .fa_or0(csa_component39_fa27_or0));
  fa fa_csa_component39_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component39_fa28_xor1), .fa_or0(csa_component39_fa28_or0));
  fa fa_csa_component39_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component39_fa29_xor1), .fa_or0(csa_component39_fa29_or0));
  fa fa_csa_component39_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component39_fa30_xor1), .fa_or0(csa_component39_fa30_or0));
  fa fa_csa_component39_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component39_fa31_xor1), .fa_or0(csa_component39_fa31_or0));
  fa fa_csa_component39_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component39_fa32_xor1), .fa_or0(csa_component39_fa32_or0));
  fa fa_csa_component39_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component39_fa33_xor1), .fa_or0(csa_component39_fa33_or0));
  fa fa_csa_component39_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component39_fa34_xor1), .fa_or0(csa_component39_fa34_or0));
  fa fa_csa_component39_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component39_fa35_xor1), .fa_or0(csa_component39_fa35_or0));
  fa fa_csa_component39_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component39_fa36_xor1), .fa_or0(csa_component39_fa36_or0));
  fa fa_csa_component39_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component39_fa37_xor1), .fa_or0(csa_component39_fa37_or0));
  fa fa_csa_component39_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component39_fa38_xor1), .fa_or0(csa_component39_fa38_or0));

  assign csa_component39_out[0] = csa_component39_fa0_xor1[0];
  assign csa_component39_out[1] = csa_component39_fa1_xor1[0];
  assign csa_component39_out[2] = csa_component39_fa2_xor1[0];
  assign csa_component39_out[3] = csa_component39_fa3_xor1[0];
  assign csa_component39_out[4] = csa_component39_fa4_xor1[0];
  assign csa_component39_out[5] = csa_component39_fa5_xor1[0];
  assign csa_component39_out[6] = csa_component39_fa6_xor1[0];
  assign csa_component39_out[7] = csa_component39_fa7_xor1[0];
  assign csa_component39_out[8] = csa_component39_fa8_xor1[0];
  assign csa_component39_out[9] = csa_component39_fa9_xor1[0];
  assign csa_component39_out[10] = csa_component39_fa10_xor1[0];
  assign csa_component39_out[11] = csa_component39_fa11_xor1[0];
  assign csa_component39_out[12] = csa_component39_fa12_xor1[0];
  assign csa_component39_out[13] = csa_component39_fa13_xor1[0];
  assign csa_component39_out[14] = csa_component39_fa14_xor1[0];
  assign csa_component39_out[15] = csa_component39_fa15_xor1[0];
  assign csa_component39_out[16] = csa_component39_fa16_xor1[0];
  assign csa_component39_out[17] = csa_component39_fa17_xor1[0];
  assign csa_component39_out[18] = csa_component39_fa18_xor1[0];
  assign csa_component39_out[19] = csa_component39_fa19_xor1[0];
  assign csa_component39_out[20] = csa_component39_fa20_xor1[0];
  assign csa_component39_out[21] = csa_component39_fa21_xor1[0];
  assign csa_component39_out[22] = csa_component39_fa22_xor1[0];
  assign csa_component39_out[23] = csa_component39_fa23_xor1[0];
  assign csa_component39_out[24] = csa_component39_fa24_xor1[0];
  assign csa_component39_out[25] = csa_component39_fa25_xor1[0];
  assign csa_component39_out[26] = csa_component39_fa26_xor1[0];
  assign csa_component39_out[27] = csa_component39_fa27_xor1[0];
  assign csa_component39_out[28] = csa_component39_fa28_xor1[0];
  assign csa_component39_out[29] = csa_component39_fa29_xor1[0];
  assign csa_component39_out[30] = csa_component39_fa30_xor1[0];
  assign csa_component39_out[31] = csa_component39_fa31_xor1[0];
  assign csa_component39_out[32] = csa_component39_fa32_xor1[0];
  assign csa_component39_out[33] = csa_component39_fa33_xor1[0];
  assign csa_component39_out[34] = csa_component39_fa34_xor1[0];
  assign csa_component39_out[35] = csa_component39_fa35_xor1[0];
  assign csa_component39_out[36] = csa_component39_fa36_xor1[0];
  assign csa_component39_out[37] = csa_component39_fa37_xor1[0];
  assign csa_component39_out[38] = csa_component39_fa38_xor1[0];
  assign csa_component39_out[39] = 1'b0;
  assign csa_component39_out[40] = 1'b0;
  assign csa_component39_out[41] = csa_component39_fa0_or0[0];
  assign csa_component39_out[42] = csa_component39_fa1_or0[0];
  assign csa_component39_out[43] = csa_component39_fa2_or0[0];
  assign csa_component39_out[44] = csa_component39_fa3_or0[0];
  assign csa_component39_out[45] = csa_component39_fa4_or0[0];
  assign csa_component39_out[46] = csa_component39_fa5_or0[0];
  assign csa_component39_out[47] = csa_component39_fa6_or0[0];
  assign csa_component39_out[48] = csa_component39_fa7_or0[0];
  assign csa_component39_out[49] = csa_component39_fa8_or0[0];
  assign csa_component39_out[50] = csa_component39_fa9_or0[0];
  assign csa_component39_out[51] = csa_component39_fa10_or0[0];
  assign csa_component39_out[52] = csa_component39_fa11_or0[0];
  assign csa_component39_out[53] = csa_component39_fa12_or0[0];
  assign csa_component39_out[54] = csa_component39_fa13_or0[0];
  assign csa_component39_out[55] = csa_component39_fa14_or0[0];
  assign csa_component39_out[56] = csa_component39_fa15_or0[0];
  assign csa_component39_out[57] = csa_component39_fa16_or0[0];
  assign csa_component39_out[58] = csa_component39_fa17_or0[0];
  assign csa_component39_out[59] = csa_component39_fa18_or0[0];
  assign csa_component39_out[60] = csa_component39_fa19_or0[0];
  assign csa_component39_out[61] = csa_component39_fa20_or0[0];
  assign csa_component39_out[62] = csa_component39_fa21_or0[0];
  assign csa_component39_out[63] = csa_component39_fa22_or0[0];
  assign csa_component39_out[64] = csa_component39_fa23_or0[0];
  assign csa_component39_out[65] = csa_component39_fa24_or0[0];
  assign csa_component39_out[66] = csa_component39_fa25_or0[0];
  assign csa_component39_out[67] = csa_component39_fa26_or0[0];
  assign csa_component39_out[68] = csa_component39_fa27_or0[0];
  assign csa_component39_out[69] = csa_component39_fa28_or0[0];
  assign csa_component39_out[70] = csa_component39_fa29_or0[0];
  assign csa_component39_out[71] = csa_component39_fa30_or0[0];
  assign csa_component39_out[72] = csa_component39_fa31_or0[0];
  assign csa_component39_out[73] = csa_component39_fa32_or0[0];
  assign csa_component39_out[74] = csa_component39_fa33_or0[0];
  assign csa_component39_out[75] = csa_component39_fa34_or0[0];
  assign csa_component39_out[76] = csa_component39_fa35_or0[0];
  assign csa_component39_out[77] = csa_component39_fa36_or0[0];
  assign csa_component39_out[78] = csa_component39_fa37_or0[0];
  assign csa_component39_out[79] = csa_component39_fa38_or0[0];
endmodule

module csa_component42(input [41:0] a, input [41:0] b, input [41:0] c, output [85:0] csa_component42_out);
  wire [0:0] csa_component42_fa0_xor1;
  wire [0:0] csa_component42_fa0_or0;
  wire [0:0] csa_component42_fa1_xor1;
  wire [0:0] csa_component42_fa1_or0;
  wire [0:0] csa_component42_fa2_xor1;
  wire [0:0] csa_component42_fa2_or0;
  wire [0:0] csa_component42_fa3_xor1;
  wire [0:0] csa_component42_fa3_or0;
  wire [0:0] csa_component42_fa4_xor1;
  wire [0:0] csa_component42_fa4_or0;
  wire [0:0] csa_component42_fa5_xor1;
  wire [0:0] csa_component42_fa5_or0;
  wire [0:0] csa_component42_fa6_xor1;
  wire [0:0] csa_component42_fa6_or0;
  wire [0:0] csa_component42_fa7_xor1;
  wire [0:0] csa_component42_fa7_or0;
  wire [0:0] csa_component42_fa8_xor1;
  wire [0:0] csa_component42_fa8_or0;
  wire [0:0] csa_component42_fa9_xor1;
  wire [0:0] csa_component42_fa9_or0;
  wire [0:0] csa_component42_fa10_xor1;
  wire [0:0] csa_component42_fa10_or0;
  wire [0:0] csa_component42_fa11_xor1;
  wire [0:0] csa_component42_fa11_or0;
  wire [0:0] csa_component42_fa12_xor1;
  wire [0:0] csa_component42_fa12_or0;
  wire [0:0] csa_component42_fa13_xor1;
  wire [0:0] csa_component42_fa13_or0;
  wire [0:0] csa_component42_fa14_xor1;
  wire [0:0] csa_component42_fa14_or0;
  wire [0:0] csa_component42_fa15_xor1;
  wire [0:0] csa_component42_fa15_or0;
  wire [0:0] csa_component42_fa16_xor1;
  wire [0:0] csa_component42_fa16_or0;
  wire [0:0] csa_component42_fa17_xor1;
  wire [0:0] csa_component42_fa17_or0;
  wire [0:0] csa_component42_fa18_xor1;
  wire [0:0] csa_component42_fa18_or0;
  wire [0:0] csa_component42_fa19_xor1;
  wire [0:0] csa_component42_fa19_or0;
  wire [0:0] csa_component42_fa20_xor1;
  wire [0:0] csa_component42_fa20_or0;
  wire [0:0] csa_component42_fa21_xor1;
  wire [0:0] csa_component42_fa21_or0;
  wire [0:0] csa_component42_fa22_xor1;
  wire [0:0] csa_component42_fa22_or0;
  wire [0:0] csa_component42_fa23_xor1;
  wire [0:0] csa_component42_fa23_or0;
  wire [0:0] csa_component42_fa24_xor1;
  wire [0:0] csa_component42_fa24_or0;
  wire [0:0] csa_component42_fa25_xor1;
  wire [0:0] csa_component42_fa25_or0;
  wire [0:0] csa_component42_fa26_xor1;
  wire [0:0] csa_component42_fa26_or0;
  wire [0:0] csa_component42_fa27_xor1;
  wire [0:0] csa_component42_fa27_or0;
  wire [0:0] csa_component42_fa28_xor1;
  wire [0:0] csa_component42_fa28_or0;
  wire [0:0] csa_component42_fa29_xor1;
  wire [0:0] csa_component42_fa29_or0;
  wire [0:0] csa_component42_fa30_xor1;
  wire [0:0] csa_component42_fa30_or0;
  wire [0:0] csa_component42_fa31_xor1;
  wire [0:0] csa_component42_fa31_or0;
  wire [0:0] csa_component42_fa32_xor1;
  wire [0:0] csa_component42_fa32_or0;
  wire [0:0] csa_component42_fa33_xor1;
  wire [0:0] csa_component42_fa33_or0;
  wire [0:0] csa_component42_fa34_xor1;
  wire [0:0] csa_component42_fa34_or0;
  wire [0:0] csa_component42_fa35_xor1;
  wire [0:0] csa_component42_fa35_or0;
  wire [0:0] csa_component42_fa36_xor1;
  wire [0:0] csa_component42_fa36_or0;
  wire [0:0] csa_component42_fa37_xor1;
  wire [0:0] csa_component42_fa37_or0;
  wire [0:0] csa_component42_fa38_xor1;
  wire [0:0] csa_component42_fa38_or0;
  wire [0:0] csa_component42_fa39_xor1;
  wire [0:0] csa_component42_fa39_or0;
  wire [0:0] csa_component42_fa40_xor1;
  wire [0:0] csa_component42_fa40_or0;
  wire [0:0] csa_component42_fa41_xor1;
  wire [0:0] csa_component42_fa41_or0;

  fa fa_csa_component42_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component42_fa0_xor1), .fa_or0(csa_component42_fa0_or0));
  fa fa_csa_component42_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component42_fa1_xor1), .fa_or0(csa_component42_fa1_or0));
  fa fa_csa_component42_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component42_fa2_xor1), .fa_or0(csa_component42_fa2_or0));
  fa fa_csa_component42_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component42_fa3_xor1), .fa_or0(csa_component42_fa3_or0));
  fa fa_csa_component42_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component42_fa4_xor1), .fa_or0(csa_component42_fa4_or0));
  fa fa_csa_component42_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component42_fa5_xor1), .fa_or0(csa_component42_fa5_or0));
  fa fa_csa_component42_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component42_fa6_xor1), .fa_or0(csa_component42_fa6_or0));
  fa fa_csa_component42_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component42_fa7_xor1), .fa_or0(csa_component42_fa7_or0));
  fa fa_csa_component42_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component42_fa8_xor1), .fa_or0(csa_component42_fa8_or0));
  fa fa_csa_component42_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component42_fa9_xor1), .fa_or0(csa_component42_fa9_or0));
  fa fa_csa_component42_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component42_fa10_xor1), .fa_or0(csa_component42_fa10_or0));
  fa fa_csa_component42_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component42_fa11_xor1), .fa_or0(csa_component42_fa11_or0));
  fa fa_csa_component42_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component42_fa12_xor1), .fa_or0(csa_component42_fa12_or0));
  fa fa_csa_component42_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component42_fa13_xor1), .fa_or0(csa_component42_fa13_or0));
  fa fa_csa_component42_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component42_fa14_xor1), .fa_or0(csa_component42_fa14_or0));
  fa fa_csa_component42_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component42_fa15_xor1), .fa_or0(csa_component42_fa15_or0));
  fa fa_csa_component42_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component42_fa16_xor1), .fa_or0(csa_component42_fa16_or0));
  fa fa_csa_component42_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component42_fa17_xor1), .fa_or0(csa_component42_fa17_or0));
  fa fa_csa_component42_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component42_fa18_xor1), .fa_or0(csa_component42_fa18_or0));
  fa fa_csa_component42_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component42_fa19_xor1), .fa_or0(csa_component42_fa19_or0));
  fa fa_csa_component42_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component42_fa20_xor1), .fa_or0(csa_component42_fa20_or0));
  fa fa_csa_component42_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component42_fa21_xor1), .fa_or0(csa_component42_fa21_or0));
  fa fa_csa_component42_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component42_fa22_xor1), .fa_or0(csa_component42_fa22_or0));
  fa fa_csa_component42_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component42_fa23_xor1), .fa_or0(csa_component42_fa23_or0));
  fa fa_csa_component42_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component42_fa24_xor1), .fa_or0(csa_component42_fa24_or0));
  fa fa_csa_component42_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component42_fa25_xor1), .fa_or0(csa_component42_fa25_or0));
  fa fa_csa_component42_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component42_fa26_xor1), .fa_or0(csa_component42_fa26_or0));
  fa fa_csa_component42_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component42_fa27_xor1), .fa_or0(csa_component42_fa27_or0));
  fa fa_csa_component42_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component42_fa28_xor1), .fa_or0(csa_component42_fa28_or0));
  fa fa_csa_component42_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component42_fa29_xor1), .fa_or0(csa_component42_fa29_or0));
  fa fa_csa_component42_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component42_fa30_xor1), .fa_or0(csa_component42_fa30_or0));
  fa fa_csa_component42_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component42_fa31_xor1), .fa_or0(csa_component42_fa31_or0));
  fa fa_csa_component42_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component42_fa32_xor1), .fa_or0(csa_component42_fa32_or0));
  fa fa_csa_component42_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component42_fa33_xor1), .fa_or0(csa_component42_fa33_or0));
  fa fa_csa_component42_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component42_fa34_xor1), .fa_or0(csa_component42_fa34_or0));
  fa fa_csa_component42_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component42_fa35_xor1), .fa_or0(csa_component42_fa35_or0));
  fa fa_csa_component42_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component42_fa36_xor1), .fa_or0(csa_component42_fa36_or0));
  fa fa_csa_component42_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component42_fa37_xor1), .fa_or0(csa_component42_fa37_or0));
  fa fa_csa_component42_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component42_fa38_xor1), .fa_or0(csa_component42_fa38_or0));
  fa fa_csa_component42_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component42_fa39_xor1), .fa_or0(csa_component42_fa39_or0));
  fa fa_csa_component42_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component42_fa40_xor1), .fa_or0(csa_component42_fa40_or0));
  fa fa_csa_component42_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component42_fa41_xor1), .fa_or0(csa_component42_fa41_or0));

  assign csa_component42_out[0] = csa_component42_fa0_xor1[0];
  assign csa_component42_out[1] = csa_component42_fa1_xor1[0];
  assign csa_component42_out[2] = csa_component42_fa2_xor1[0];
  assign csa_component42_out[3] = csa_component42_fa3_xor1[0];
  assign csa_component42_out[4] = csa_component42_fa4_xor1[0];
  assign csa_component42_out[5] = csa_component42_fa5_xor1[0];
  assign csa_component42_out[6] = csa_component42_fa6_xor1[0];
  assign csa_component42_out[7] = csa_component42_fa7_xor1[0];
  assign csa_component42_out[8] = csa_component42_fa8_xor1[0];
  assign csa_component42_out[9] = csa_component42_fa9_xor1[0];
  assign csa_component42_out[10] = csa_component42_fa10_xor1[0];
  assign csa_component42_out[11] = csa_component42_fa11_xor1[0];
  assign csa_component42_out[12] = csa_component42_fa12_xor1[0];
  assign csa_component42_out[13] = csa_component42_fa13_xor1[0];
  assign csa_component42_out[14] = csa_component42_fa14_xor1[0];
  assign csa_component42_out[15] = csa_component42_fa15_xor1[0];
  assign csa_component42_out[16] = csa_component42_fa16_xor1[0];
  assign csa_component42_out[17] = csa_component42_fa17_xor1[0];
  assign csa_component42_out[18] = csa_component42_fa18_xor1[0];
  assign csa_component42_out[19] = csa_component42_fa19_xor1[0];
  assign csa_component42_out[20] = csa_component42_fa20_xor1[0];
  assign csa_component42_out[21] = csa_component42_fa21_xor1[0];
  assign csa_component42_out[22] = csa_component42_fa22_xor1[0];
  assign csa_component42_out[23] = csa_component42_fa23_xor1[0];
  assign csa_component42_out[24] = csa_component42_fa24_xor1[0];
  assign csa_component42_out[25] = csa_component42_fa25_xor1[0];
  assign csa_component42_out[26] = csa_component42_fa26_xor1[0];
  assign csa_component42_out[27] = csa_component42_fa27_xor1[0];
  assign csa_component42_out[28] = csa_component42_fa28_xor1[0];
  assign csa_component42_out[29] = csa_component42_fa29_xor1[0];
  assign csa_component42_out[30] = csa_component42_fa30_xor1[0];
  assign csa_component42_out[31] = csa_component42_fa31_xor1[0];
  assign csa_component42_out[32] = csa_component42_fa32_xor1[0];
  assign csa_component42_out[33] = csa_component42_fa33_xor1[0];
  assign csa_component42_out[34] = csa_component42_fa34_xor1[0];
  assign csa_component42_out[35] = csa_component42_fa35_xor1[0];
  assign csa_component42_out[36] = csa_component42_fa36_xor1[0];
  assign csa_component42_out[37] = csa_component42_fa37_xor1[0];
  assign csa_component42_out[38] = csa_component42_fa38_xor1[0];
  assign csa_component42_out[39] = csa_component42_fa39_xor1[0];
  assign csa_component42_out[40] = csa_component42_fa40_xor1[0];
  assign csa_component42_out[41] = csa_component42_fa41_xor1[0];
  assign csa_component42_out[42] = 1'b0;
  assign csa_component42_out[43] = 1'b0;
  assign csa_component42_out[44] = csa_component42_fa0_or0[0];
  assign csa_component42_out[45] = csa_component42_fa1_or0[0];
  assign csa_component42_out[46] = csa_component42_fa2_or0[0];
  assign csa_component42_out[47] = csa_component42_fa3_or0[0];
  assign csa_component42_out[48] = csa_component42_fa4_or0[0];
  assign csa_component42_out[49] = csa_component42_fa5_or0[0];
  assign csa_component42_out[50] = csa_component42_fa6_or0[0];
  assign csa_component42_out[51] = csa_component42_fa7_or0[0];
  assign csa_component42_out[52] = csa_component42_fa8_or0[0];
  assign csa_component42_out[53] = csa_component42_fa9_or0[0];
  assign csa_component42_out[54] = csa_component42_fa10_or0[0];
  assign csa_component42_out[55] = csa_component42_fa11_or0[0];
  assign csa_component42_out[56] = csa_component42_fa12_or0[0];
  assign csa_component42_out[57] = csa_component42_fa13_or0[0];
  assign csa_component42_out[58] = csa_component42_fa14_or0[0];
  assign csa_component42_out[59] = csa_component42_fa15_or0[0];
  assign csa_component42_out[60] = csa_component42_fa16_or0[0];
  assign csa_component42_out[61] = csa_component42_fa17_or0[0];
  assign csa_component42_out[62] = csa_component42_fa18_or0[0];
  assign csa_component42_out[63] = csa_component42_fa19_or0[0];
  assign csa_component42_out[64] = csa_component42_fa20_or0[0];
  assign csa_component42_out[65] = csa_component42_fa21_or0[0];
  assign csa_component42_out[66] = csa_component42_fa22_or0[0];
  assign csa_component42_out[67] = csa_component42_fa23_or0[0];
  assign csa_component42_out[68] = csa_component42_fa24_or0[0];
  assign csa_component42_out[69] = csa_component42_fa25_or0[0];
  assign csa_component42_out[70] = csa_component42_fa26_or0[0];
  assign csa_component42_out[71] = csa_component42_fa27_or0[0];
  assign csa_component42_out[72] = csa_component42_fa28_or0[0];
  assign csa_component42_out[73] = csa_component42_fa29_or0[0];
  assign csa_component42_out[74] = csa_component42_fa30_or0[0];
  assign csa_component42_out[75] = csa_component42_fa31_or0[0];
  assign csa_component42_out[76] = csa_component42_fa32_or0[0];
  assign csa_component42_out[77] = csa_component42_fa33_or0[0];
  assign csa_component42_out[78] = csa_component42_fa34_or0[0];
  assign csa_component42_out[79] = csa_component42_fa35_or0[0];
  assign csa_component42_out[80] = csa_component42_fa36_or0[0];
  assign csa_component42_out[81] = csa_component42_fa37_or0[0];
  assign csa_component42_out[82] = csa_component42_fa38_or0[0];
  assign csa_component42_out[83] = csa_component42_fa39_or0[0];
  assign csa_component42_out[84] = csa_component42_fa40_or0[0];
  assign csa_component42_out[85] = csa_component42_fa41_or0[0];
endmodule

module csa_component48(input [47:0] a, input [47:0] b, input [47:0] c, output [97:0] csa_component48_out);
  wire [0:0] csa_component48_fa0_xor1;
  wire [0:0] csa_component48_fa0_or0;
  wire [0:0] csa_component48_fa1_xor1;
  wire [0:0] csa_component48_fa1_or0;
  wire [0:0] csa_component48_fa2_xor1;
  wire [0:0] csa_component48_fa2_or0;
  wire [0:0] csa_component48_fa3_xor1;
  wire [0:0] csa_component48_fa3_or0;
  wire [0:0] csa_component48_fa4_xor1;
  wire [0:0] csa_component48_fa4_or0;
  wire [0:0] csa_component48_fa5_xor1;
  wire [0:0] csa_component48_fa5_or0;
  wire [0:0] csa_component48_fa6_xor1;
  wire [0:0] csa_component48_fa6_or0;
  wire [0:0] csa_component48_fa7_xor1;
  wire [0:0] csa_component48_fa7_or0;
  wire [0:0] csa_component48_fa8_xor1;
  wire [0:0] csa_component48_fa8_or0;
  wire [0:0] csa_component48_fa9_xor1;
  wire [0:0] csa_component48_fa9_or0;
  wire [0:0] csa_component48_fa10_xor1;
  wire [0:0] csa_component48_fa10_or0;
  wire [0:0] csa_component48_fa11_xor1;
  wire [0:0] csa_component48_fa11_or0;
  wire [0:0] csa_component48_fa12_xor1;
  wire [0:0] csa_component48_fa12_or0;
  wire [0:0] csa_component48_fa13_xor1;
  wire [0:0] csa_component48_fa13_or0;
  wire [0:0] csa_component48_fa14_xor1;
  wire [0:0] csa_component48_fa14_or0;
  wire [0:0] csa_component48_fa15_xor1;
  wire [0:0] csa_component48_fa15_or0;
  wire [0:0] csa_component48_fa16_xor1;
  wire [0:0] csa_component48_fa16_or0;
  wire [0:0] csa_component48_fa17_xor1;
  wire [0:0] csa_component48_fa17_or0;
  wire [0:0] csa_component48_fa18_xor1;
  wire [0:0] csa_component48_fa18_or0;
  wire [0:0] csa_component48_fa19_xor1;
  wire [0:0] csa_component48_fa19_or0;
  wire [0:0] csa_component48_fa20_xor1;
  wire [0:0] csa_component48_fa20_or0;
  wire [0:0] csa_component48_fa21_xor1;
  wire [0:0] csa_component48_fa21_or0;
  wire [0:0] csa_component48_fa22_xor1;
  wire [0:0] csa_component48_fa22_or0;
  wire [0:0] csa_component48_fa23_xor1;
  wire [0:0] csa_component48_fa23_or0;
  wire [0:0] csa_component48_fa24_xor1;
  wire [0:0] csa_component48_fa24_or0;
  wire [0:0] csa_component48_fa25_xor1;
  wire [0:0] csa_component48_fa25_or0;
  wire [0:0] csa_component48_fa26_xor1;
  wire [0:0] csa_component48_fa26_or0;
  wire [0:0] csa_component48_fa27_xor1;
  wire [0:0] csa_component48_fa27_or0;
  wire [0:0] csa_component48_fa28_xor1;
  wire [0:0] csa_component48_fa28_or0;
  wire [0:0] csa_component48_fa29_xor1;
  wire [0:0] csa_component48_fa29_or0;
  wire [0:0] csa_component48_fa30_xor1;
  wire [0:0] csa_component48_fa30_or0;
  wire [0:0] csa_component48_fa31_xor1;
  wire [0:0] csa_component48_fa31_or0;
  wire [0:0] csa_component48_fa32_xor1;
  wire [0:0] csa_component48_fa32_or0;
  wire [0:0] csa_component48_fa33_xor1;
  wire [0:0] csa_component48_fa33_or0;
  wire [0:0] csa_component48_fa34_xor1;
  wire [0:0] csa_component48_fa34_or0;
  wire [0:0] csa_component48_fa35_xor1;
  wire [0:0] csa_component48_fa35_or0;
  wire [0:0] csa_component48_fa36_xor1;
  wire [0:0] csa_component48_fa36_or0;
  wire [0:0] csa_component48_fa37_xor1;
  wire [0:0] csa_component48_fa37_or0;
  wire [0:0] csa_component48_fa38_xor1;
  wire [0:0] csa_component48_fa38_or0;
  wire [0:0] csa_component48_fa39_xor1;
  wire [0:0] csa_component48_fa39_or0;
  wire [0:0] csa_component48_fa40_xor1;
  wire [0:0] csa_component48_fa40_or0;
  wire [0:0] csa_component48_fa41_xor1;
  wire [0:0] csa_component48_fa41_or0;
  wire [0:0] csa_component48_fa42_xor1;
  wire [0:0] csa_component48_fa42_or0;
  wire [0:0] csa_component48_fa43_xor1;
  wire [0:0] csa_component48_fa43_or0;
  wire [0:0] csa_component48_fa44_xor1;
  wire [0:0] csa_component48_fa44_or0;
  wire [0:0] csa_component48_fa45_xor1;
  wire [0:0] csa_component48_fa45_or0;
  wire [0:0] csa_component48_fa46_xor1;
  wire [0:0] csa_component48_fa46_or0;
  wire [0:0] csa_component48_fa47_xor1;
  wire [0:0] csa_component48_fa47_or0;

  fa fa_csa_component48_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component48_fa0_xor1), .fa_or0(csa_component48_fa0_or0));
  fa fa_csa_component48_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component48_fa1_xor1), .fa_or0(csa_component48_fa1_or0));
  fa fa_csa_component48_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component48_fa2_xor1), .fa_or0(csa_component48_fa2_or0));
  fa fa_csa_component48_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component48_fa3_xor1), .fa_or0(csa_component48_fa3_or0));
  fa fa_csa_component48_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component48_fa4_xor1), .fa_or0(csa_component48_fa4_or0));
  fa fa_csa_component48_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component48_fa5_xor1), .fa_or0(csa_component48_fa5_or0));
  fa fa_csa_component48_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component48_fa6_xor1), .fa_or0(csa_component48_fa6_or0));
  fa fa_csa_component48_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component48_fa7_xor1), .fa_or0(csa_component48_fa7_or0));
  fa fa_csa_component48_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component48_fa8_xor1), .fa_or0(csa_component48_fa8_or0));
  fa fa_csa_component48_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component48_fa9_xor1), .fa_or0(csa_component48_fa9_or0));
  fa fa_csa_component48_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component48_fa10_xor1), .fa_or0(csa_component48_fa10_or0));
  fa fa_csa_component48_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component48_fa11_xor1), .fa_or0(csa_component48_fa11_or0));
  fa fa_csa_component48_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component48_fa12_xor1), .fa_or0(csa_component48_fa12_or0));
  fa fa_csa_component48_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component48_fa13_xor1), .fa_or0(csa_component48_fa13_or0));
  fa fa_csa_component48_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component48_fa14_xor1), .fa_or0(csa_component48_fa14_or0));
  fa fa_csa_component48_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component48_fa15_xor1), .fa_or0(csa_component48_fa15_or0));
  fa fa_csa_component48_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component48_fa16_xor1), .fa_or0(csa_component48_fa16_or0));
  fa fa_csa_component48_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component48_fa17_xor1), .fa_or0(csa_component48_fa17_or0));
  fa fa_csa_component48_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component48_fa18_xor1), .fa_or0(csa_component48_fa18_or0));
  fa fa_csa_component48_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component48_fa19_xor1), .fa_or0(csa_component48_fa19_or0));
  fa fa_csa_component48_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component48_fa20_xor1), .fa_or0(csa_component48_fa20_or0));
  fa fa_csa_component48_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component48_fa21_xor1), .fa_or0(csa_component48_fa21_or0));
  fa fa_csa_component48_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component48_fa22_xor1), .fa_or0(csa_component48_fa22_or0));
  fa fa_csa_component48_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component48_fa23_xor1), .fa_or0(csa_component48_fa23_or0));
  fa fa_csa_component48_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component48_fa24_xor1), .fa_or0(csa_component48_fa24_or0));
  fa fa_csa_component48_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component48_fa25_xor1), .fa_or0(csa_component48_fa25_or0));
  fa fa_csa_component48_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component48_fa26_xor1), .fa_or0(csa_component48_fa26_or0));
  fa fa_csa_component48_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component48_fa27_xor1), .fa_or0(csa_component48_fa27_or0));
  fa fa_csa_component48_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component48_fa28_xor1), .fa_or0(csa_component48_fa28_or0));
  fa fa_csa_component48_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component48_fa29_xor1), .fa_or0(csa_component48_fa29_or0));
  fa fa_csa_component48_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component48_fa30_xor1), .fa_or0(csa_component48_fa30_or0));
  fa fa_csa_component48_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component48_fa31_xor1), .fa_or0(csa_component48_fa31_or0));
  fa fa_csa_component48_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component48_fa32_xor1), .fa_or0(csa_component48_fa32_or0));
  fa fa_csa_component48_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component48_fa33_xor1), .fa_or0(csa_component48_fa33_or0));
  fa fa_csa_component48_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component48_fa34_xor1), .fa_or0(csa_component48_fa34_or0));
  fa fa_csa_component48_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component48_fa35_xor1), .fa_or0(csa_component48_fa35_or0));
  fa fa_csa_component48_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component48_fa36_xor1), .fa_or0(csa_component48_fa36_or0));
  fa fa_csa_component48_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component48_fa37_xor1), .fa_or0(csa_component48_fa37_or0));
  fa fa_csa_component48_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component48_fa38_xor1), .fa_or0(csa_component48_fa38_or0));
  fa fa_csa_component48_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component48_fa39_xor1), .fa_or0(csa_component48_fa39_or0));
  fa fa_csa_component48_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component48_fa40_xor1), .fa_or0(csa_component48_fa40_or0));
  fa fa_csa_component48_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component48_fa41_xor1), .fa_or0(csa_component48_fa41_or0));
  fa fa_csa_component48_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component48_fa42_xor1), .fa_or0(csa_component48_fa42_or0));
  fa fa_csa_component48_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component48_fa43_xor1), .fa_or0(csa_component48_fa43_or0));
  fa fa_csa_component48_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component48_fa44_xor1), .fa_or0(csa_component48_fa44_or0));
  fa fa_csa_component48_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component48_fa45_xor1), .fa_or0(csa_component48_fa45_or0));
  fa fa_csa_component48_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component48_fa46_xor1), .fa_or0(csa_component48_fa46_or0));
  fa fa_csa_component48_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component48_fa47_xor1), .fa_or0(csa_component48_fa47_or0));

  assign csa_component48_out[0] = csa_component48_fa0_xor1[0];
  assign csa_component48_out[1] = csa_component48_fa1_xor1[0];
  assign csa_component48_out[2] = csa_component48_fa2_xor1[0];
  assign csa_component48_out[3] = csa_component48_fa3_xor1[0];
  assign csa_component48_out[4] = csa_component48_fa4_xor1[0];
  assign csa_component48_out[5] = csa_component48_fa5_xor1[0];
  assign csa_component48_out[6] = csa_component48_fa6_xor1[0];
  assign csa_component48_out[7] = csa_component48_fa7_xor1[0];
  assign csa_component48_out[8] = csa_component48_fa8_xor1[0];
  assign csa_component48_out[9] = csa_component48_fa9_xor1[0];
  assign csa_component48_out[10] = csa_component48_fa10_xor1[0];
  assign csa_component48_out[11] = csa_component48_fa11_xor1[0];
  assign csa_component48_out[12] = csa_component48_fa12_xor1[0];
  assign csa_component48_out[13] = csa_component48_fa13_xor1[0];
  assign csa_component48_out[14] = csa_component48_fa14_xor1[0];
  assign csa_component48_out[15] = csa_component48_fa15_xor1[0];
  assign csa_component48_out[16] = csa_component48_fa16_xor1[0];
  assign csa_component48_out[17] = csa_component48_fa17_xor1[0];
  assign csa_component48_out[18] = csa_component48_fa18_xor1[0];
  assign csa_component48_out[19] = csa_component48_fa19_xor1[0];
  assign csa_component48_out[20] = csa_component48_fa20_xor1[0];
  assign csa_component48_out[21] = csa_component48_fa21_xor1[0];
  assign csa_component48_out[22] = csa_component48_fa22_xor1[0];
  assign csa_component48_out[23] = csa_component48_fa23_xor1[0];
  assign csa_component48_out[24] = csa_component48_fa24_xor1[0];
  assign csa_component48_out[25] = csa_component48_fa25_xor1[0];
  assign csa_component48_out[26] = csa_component48_fa26_xor1[0];
  assign csa_component48_out[27] = csa_component48_fa27_xor1[0];
  assign csa_component48_out[28] = csa_component48_fa28_xor1[0];
  assign csa_component48_out[29] = csa_component48_fa29_xor1[0];
  assign csa_component48_out[30] = csa_component48_fa30_xor1[0];
  assign csa_component48_out[31] = csa_component48_fa31_xor1[0];
  assign csa_component48_out[32] = csa_component48_fa32_xor1[0];
  assign csa_component48_out[33] = csa_component48_fa33_xor1[0];
  assign csa_component48_out[34] = csa_component48_fa34_xor1[0];
  assign csa_component48_out[35] = csa_component48_fa35_xor1[0];
  assign csa_component48_out[36] = csa_component48_fa36_xor1[0];
  assign csa_component48_out[37] = csa_component48_fa37_xor1[0];
  assign csa_component48_out[38] = csa_component48_fa38_xor1[0];
  assign csa_component48_out[39] = csa_component48_fa39_xor1[0];
  assign csa_component48_out[40] = csa_component48_fa40_xor1[0];
  assign csa_component48_out[41] = csa_component48_fa41_xor1[0];
  assign csa_component48_out[42] = csa_component48_fa42_xor1[0];
  assign csa_component48_out[43] = csa_component48_fa43_xor1[0];
  assign csa_component48_out[44] = csa_component48_fa44_xor1[0];
  assign csa_component48_out[45] = csa_component48_fa45_xor1[0];
  assign csa_component48_out[46] = csa_component48_fa46_xor1[0];
  assign csa_component48_out[47] = csa_component48_fa47_xor1[0];
  assign csa_component48_out[48] = 1'b0;
  assign csa_component48_out[49] = 1'b0;
  assign csa_component48_out[50] = csa_component48_fa0_or0[0];
  assign csa_component48_out[51] = csa_component48_fa1_or0[0];
  assign csa_component48_out[52] = csa_component48_fa2_or0[0];
  assign csa_component48_out[53] = csa_component48_fa3_or0[0];
  assign csa_component48_out[54] = csa_component48_fa4_or0[0];
  assign csa_component48_out[55] = csa_component48_fa5_or0[0];
  assign csa_component48_out[56] = csa_component48_fa6_or0[0];
  assign csa_component48_out[57] = csa_component48_fa7_or0[0];
  assign csa_component48_out[58] = csa_component48_fa8_or0[0];
  assign csa_component48_out[59] = csa_component48_fa9_or0[0];
  assign csa_component48_out[60] = csa_component48_fa10_or0[0];
  assign csa_component48_out[61] = csa_component48_fa11_or0[0];
  assign csa_component48_out[62] = csa_component48_fa12_or0[0];
  assign csa_component48_out[63] = csa_component48_fa13_or0[0];
  assign csa_component48_out[64] = csa_component48_fa14_or0[0];
  assign csa_component48_out[65] = csa_component48_fa15_or0[0];
  assign csa_component48_out[66] = csa_component48_fa16_or0[0];
  assign csa_component48_out[67] = csa_component48_fa17_or0[0];
  assign csa_component48_out[68] = csa_component48_fa18_or0[0];
  assign csa_component48_out[69] = csa_component48_fa19_or0[0];
  assign csa_component48_out[70] = csa_component48_fa20_or0[0];
  assign csa_component48_out[71] = csa_component48_fa21_or0[0];
  assign csa_component48_out[72] = csa_component48_fa22_or0[0];
  assign csa_component48_out[73] = csa_component48_fa23_or0[0];
  assign csa_component48_out[74] = csa_component48_fa24_or0[0];
  assign csa_component48_out[75] = csa_component48_fa25_or0[0];
  assign csa_component48_out[76] = csa_component48_fa26_or0[0];
  assign csa_component48_out[77] = csa_component48_fa27_or0[0];
  assign csa_component48_out[78] = csa_component48_fa28_or0[0];
  assign csa_component48_out[79] = csa_component48_fa29_or0[0];
  assign csa_component48_out[80] = csa_component48_fa30_or0[0];
  assign csa_component48_out[81] = csa_component48_fa31_or0[0];
  assign csa_component48_out[82] = csa_component48_fa32_or0[0];
  assign csa_component48_out[83] = csa_component48_fa33_or0[0];
  assign csa_component48_out[84] = csa_component48_fa34_or0[0];
  assign csa_component48_out[85] = csa_component48_fa35_or0[0];
  assign csa_component48_out[86] = csa_component48_fa36_or0[0];
  assign csa_component48_out[87] = csa_component48_fa37_or0[0];
  assign csa_component48_out[88] = csa_component48_fa38_or0[0];
  assign csa_component48_out[89] = csa_component48_fa39_or0[0];
  assign csa_component48_out[90] = csa_component48_fa40_or0[0];
  assign csa_component48_out[91] = csa_component48_fa41_or0[0];
  assign csa_component48_out[92] = csa_component48_fa42_or0[0];
  assign csa_component48_out[93] = csa_component48_fa43_or0[0];
  assign csa_component48_out[94] = csa_component48_fa44_or0[0];
  assign csa_component48_out[95] = csa_component48_fa45_or0[0];
  assign csa_component48_out[96] = csa_component48_fa46_or0[0];
  assign csa_component48_out[97] = csa_component48_fa47_or0[0];
endmodule

module csa_component34(input [33:0] a, input [33:0] b, input [33:0] c, output [69:0] csa_component34_out);
  wire [0:0] csa_component34_fa0_xor1;
  wire [0:0] csa_component34_fa0_or0;
  wire [0:0] csa_component34_fa1_xor1;
  wire [0:0] csa_component34_fa1_or0;
  wire [0:0] csa_component34_fa2_xor1;
  wire [0:0] csa_component34_fa2_or0;
  wire [0:0] csa_component34_fa3_xor1;
  wire [0:0] csa_component34_fa3_or0;
  wire [0:0] csa_component34_fa4_xor1;
  wire [0:0] csa_component34_fa4_or0;
  wire [0:0] csa_component34_fa5_xor1;
  wire [0:0] csa_component34_fa5_or0;
  wire [0:0] csa_component34_fa6_xor1;
  wire [0:0] csa_component34_fa6_or0;
  wire [0:0] csa_component34_fa7_xor1;
  wire [0:0] csa_component34_fa7_or0;
  wire [0:0] csa_component34_fa8_xor1;
  wire [0:0] csa_component34_fa8_or0;
  wire [0:0] csa_component34_fa9_xor1;
  wire [0:0] csa_component34_fa9_or0;
  wire [0:0] csa_component34_fa10_xor1;
  wire [0:0] csa_component34_fa10_or0;
  wire [0:0] csa_component34_fa11_xor1;
  wire [0:0] csa_component34_fa11_or0;
  wire [0:0] csa_component34_fa12_xor1;
  wire [0:0] csa_component34_fa12_or0;
  wire [0:0] csa_component34_fa13_xor1;
  wire [0:0] csa_component34_fa13_or0;
  wire [0:0] csa_component34_fa14_xor1;
  wire [0:0] csa_component34_fa14_or0;
  wire [0:0] csa_component34_fa15_xor1;
  wire [0:0] csa_component34_fa15_or0;
  wire [0:0] csa_component34_fa16_xor1;
  wire [0:0] csa_component34_fa16_or0;
  wire [0:0] csa_component34_fa17_xor1;
  wire [0:0] csa_component34_fa17_or0;
  wire [0:0] csa_component34_fa18_xor1;
  wire [0:0] csa_component34_fa18_or0;
  wire [0:0] csa_component34_fa19_xor1;
  wire [0:0] csa_component34_fa19_or0;
  wire [0:0] csa_component34_fa20_xor1;
  wire [0:0] csa_component34_fa20_or0;
  wire [0:0] csa_component34_fa21_xor1;
  wire [0:0] csa_component34_fa21_or0;
  wire [0:0] csa_component34_fa22_xor1;
  wire [0:0] csa_component34_fa22_or0;
  wire [0:0] csa_component34_fa23_xor1;
  wire [0:0] csa_component34_fa23_or0;
  wire [0:0] csa_component34_fa24_xor1;
  wire [0:0] csa_component34_fa24_or0;
  wire [0:0] csa_component34_fa25_xor1;
  wire [0:0] csa_component34_fa25_or0;
  wire [0:0] csa_component34_fa26_xor1;
  wire [0:0] csa_component34_fa26_or0;
  wire [0:0] csa_component34_fa27_xor1;
  wire [0:0] csa_component34_fa27_or0;
  wire [0:0] csa_component34_fa28_xor1;
  wire [0:0] csa_component34_fa28_or0;
  wire [0:0] csa_component34_fa29_xor1;
  wire [0:0] csa_component34_fa29_or0;
  wire [0:0] csa_component34_fa30_xor1;
  wire [0:0] csa_component34_fa30_or0;
  wire [0:0] csa_component34_fa31_xor1;
  wire [0:0] csa_component34_fa31_or0;
  wire [0:0] csa_component34_fa32_xor1;
  wire [0:0] csa_component34_fa32_or0;
  wire [0:0] csa_component34_fa33_xor1;
  wire [0:0] csa_component34_fa33_or0;

  fa fa_csa_component34_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component34_fa0_xor1), .fa_or0(csa_component34_fa0_or0));
  fa fa_csa_component34_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component34_fa1_xor1), .fa_or0(csa_component34_fa1_or0));
  fa fa_csa_component34_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component34_fa2_xor1), .fa_or0(csa_component34_fa2_or0));
  fa fa_csa_component34_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component34_fa3_xor1), .fa_or0(csa_component34_fa3_or0));
  fa fa_csa_component34_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component34_fa4_xor1), .fa_or0(csa_component34_fa4_or0));
  fa fa_csa_component34_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component34_fa5_xor1), .fa_or0(csa_component34_fa5_or0));
  fa fa_csa_component34_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component34_fa6_xor1), .fa_or0(csa_component34_fa6_or0));
  fa fa_csa_component34_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component34_fa7_xor1), .fa_or0(csa_component34_fa7_or0));
  fa fa_csa_component34_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component34_fa8_xor1), .fa_or0(csa_component34_fa8_or0));
  fa fa_csa_component34_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component34_fa9_xor1), .fa_or0(csa_component34_fa9_or0));
  fa fa_csa_component34_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component34_fa10_xor1), .fa_or0(csa_component34_fa10_or0));
  fa fa_csa_component34_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component34_fa11_xor1), .fa_or0(csa_component34_fa11_or0));
  fa fa_csa_component34_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component34_fa12_xor1), .fa_or0(csa_component34_fa12_or0));
  fa fa_csa_component34_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component34_fa13_xor1), .fa_or0(csa_component34_fa13_or0));
  fa fa_csa_component34_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component34_fa14_xor1), .fa_or0(csa_component34_fa14_or0));
  fa fa_csa_component34_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component34_fa15_xor1), .fa_or0(csa_component34_fa15_or0));
  fa fa_csa_component34_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component34_fa16_xor1), .fa_or0(csa_component34_fa16_or0));
  fa fa_csa_component34_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component34_fa17_xor1), .fa_or0(csa_component34_fa17_or0));
  fa fa_csa_component34_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component34_fa18_xor1), .fa_or0(csa_component34_fa18_or0));
  fa fa_csa_component34_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component34_fa19_xor1), .fa_or0(csa_component34_fa19_or0));
  fa fa_csa_component34_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component34_fa20_xor1), .fa_or0(csa_component34_fa20_or0));
  fa fa_csa_component34_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component34_fa21_xor1), .fa_or0(csa_component34_fa21_or0));
  fa fa_csa_component34_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component34_fa22_xor1), .fa_or0(csa_component34_fa22_or0));
  fa fa_csa_component34_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component34_fa23_xor1), .fa_or0(csa_component34_fa23_or0));
  fa fa_csa_component34_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component34_fa24_xor1), .fa_or0(csa_component34_fa24_or0));
  fa fa_csa_component34_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component34_fa25_xor1), .fa_or0(csa_component34_fa25_or0));
  fa fa_csa_component34_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component34_fa26_xor1), .fa_or0(csa_component34_fa26_or0));
  fa fa_csa_component34_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component34_fa27_xor1), .fa_or0(csa_component34_fa27_or0));
  fa fa_csa_component34_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component34_fa28_xor1), .fa_or0(csa_component34_fa28_or0));
  fa fa_csa_component34_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component34_fa29_xor1), .fa_or0(csa_component34_fa29_or0));
  fa fa_csa_component34_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component34_fa30_xor1), .fa_or0(csa_component34_fa30_or0));
  fa fa_csa_component34_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component34_fa31_xor1), .fa_or0(csa_component34_fa31_or0));
  fa fa_csa_component34_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component34_fa32_xor1), .fa_or0(csa_component34_fa32_or0));
  fa fa_csa_component34_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component34_fa33_xor1), .fa_or0(csa_component34_fa33_or0));

  assign csa_component34_out[0] = csa_component34_fa0_xor1[0];
  assign csa_component34_out[1] = csa_component34_fa1_xor1[0];
  assign csa_component34_out[2] = csa_component34_fa2_xor1[0];
  assign csa_component34_out[3] = csa_component34_fa3_xor1[0];
  assign csa_component34_out[4] = csa_component34_fa4_xor1[0];
  assign csa_component34_out[5] = csa_component34_fa5_xor1[0];
  assign csa_component34_out[6] = csa_component34_fa6_xor1[0];
  assign csa_component34_out[7] = csa_component34_fa7_xor1[0];
  assign csa_component34_out[8] = csa_component34_fa8_xor1[0];
  assign csa_component34_out[9] = csa_component34_fa9_xor1[0];
  assign csa_component34_out[10] = csa_component34_fa10_xor1[0];
  assign csa_component34_out[11] = csa_component34_fa11_xor1[0];
  assign csa_component34_out[12] = csa_component34_fa12_xor1[0];
  assign csa_component34_out[13] = csa_component34_fa13_xor1[0];
  assign csa_component34_out[14] = csa_component34_fa14_xor1[0];
  assign csa_component34_out[15] = csa_component34_fa15_xor1[0];
  assign csa_component34_out[16] = csa_component34_fa16_xor1[0];
  assign csa_component34_out[17] = csa_component34_fa17_xor1[0];
  assign csa_component34_out[18] = csa_component34_fa18_xor1[0];
  assign csa_component34_out[19] = csa_component34_fa19_xor1[0];
  assign csa_component34_out[20] = csa_component34_fa20_xor1[0];
  assign csa_component34_out[21] = csa_component34_fa21_xor1[0];
  assign csa_component34_out[22] = csa_component34_fa22_xor1[0];
  assign csa_component34_out[23] = csa_component34_fa23_xor1[0];
  assign csa_component34_out[24] = csa_component34_fa24_xor1[0];
  assign csa_component34_out[25] = csa_component34_fa25_xor1[0];
  assign csa_component34_out[26] = csa_component34_fa26_xor1[0];
  assign csa_component34_out[27] = csa_component34_fa27_xor1[0];
  assign csa_component34_out[28] = csa_component34_fa28_xor1[0];
  assign csa_component34_out[29] = csa_component34_fa29_xor1[0];
  assign csa_component34_out[30] = csa_component34_fa30_xor1[0];
  assign csa_component34_out[31] = csa_component34_fa31_xor1[0];
  assign csa_component34_out[32] = csa_component34_fa32_xor1[0];
  assign csa_component34_out[33] = csa_component34_fa33_xor1[0];
  assign csa_component34_out[34] = 1'b0;
  assign csa_component34_out[35] = 1'b0;
  assign csa_component34_out[36] = csa_component34_fa0_or0[0];
  assign csa_component34_out[37] = csa_component34_fa1_or0[0];
  assign csa_component34_out[38] = csa_component34_fa2_or0[0];
  assign csa_component34_out[39] = csa_component34_fa3_or0[0];
  assign csa_component34_out[40] = csa_component34_fa4_or0[0];
  assign csa_component34_out[41] = csa_component34_fa5_or0[0];
  assign csa_component34_out[42] = csa_component34_fa6_or0[0];
  assign csa_component34_out[43] = csa_component34_fa7_or0[0];
  assign csa_component34_out[44] = csa_component34_fa8_or0[0];
  assign csa_component34_out[45] = csa_component34_fa9_or0[0];
  assign csa_component34_out[46] = csa_component34_fa10_or0[0];
  assign csa_component34_out[47] = csa_component34_fa11_or0[0];
  assign csa_component34_out[48] = csa_component34_fa12_or0[0];
  assign csa_component34_out[49] = csa_component34_fa13_or0[0];
  assign csa_component34_out[50] = csa_component34_fa14_or0[0];
  assign csa_component34_out[51] = csa_component34_fa15_or0[0];
  assign csa_component34_out[52] = csa_component34_fa16_or0[0];
  assign csa_component34_out[53] = csa_component34_fa17_or0[0];
  assign csa_component34_out[54] = csa_component34_fa18_or0[0];
  assign csa_component34_out[55] = csa_component34_fa19_or0[0];
  assign csa_component34_out[56] = csa_component34_fa20_or0[0];
  assign csa_component34_out[57] = csa_component34_fa21_or0[0];
  assign csa_component34_out[58] = csa_component34_fa22_or0[0];
  assign csa_component34_out[59] = csa_component34_fa23_or0[0];
  assign csa_component34_out[60] = csa_component34_fa24_or0[0];
  assign csa_component34_out[61] = csa_component34_fa25_or0[0];
  assign csa_component34_out[62] = csa_component34_fa26_or0[0];
  assign csa_component34_out[63] = csa_component34_fa27_or0[0];
  assign csa_component34_out[64] = csa_component34_fa28_or0[0];
  assign csa_component34_out[65] = csa_component34_fa29_or0[0];
  assign csa_component34_out[66] = csa_component34_fa30_or0[0];
  assign csa_component34_out[67] = csa_component34_fa31_or0[0];
  assign csa_component34_out[68] = csa_component34_fa32_or0[0];
  assign csa_component34_out[69] = csa_component34_fa33_or0[0];
endmodule

module csa_component40(input [39:0] a, input [39:0] b, input [39:0] c, output [81:0] csa_component40_out);
  wire [0:0] csa_component40_fa0_xor1;
  wire [0:0] csa_component40_fa0_or0;
  wire [0:0] csa_component40_fa1_xor1;
  wire [0:0] csa_component40_fa1_or0;
  wire [0:0] csa_component40_fa2_xor1;
  wire [0:0] csa_component40_fa2_or0;
  wire [0:0] csa_component40_fa3_xor1;
  wire [0:0] csa_component40_fa3_or0;
  wire [0:0] csa_component40_fa4_xor1;
  wire [0:0] csa_component40_fa4_or0;
  wire [0:0] csa_component40_fa5_xor1;
  wire [0:0] csa_component40_fa5_or0;
  wire [0:0] csa_component40_fa6_xor1;
  wire [0:0] csa_component40_fa6_or0;
  wire [0:0] csa_component40_fa7_xor1;
  wire [0:0] csa_component40_fa7_or0;
  wire [0:0] csa_component40_fa8_xor1;
  wire [0:0] csa_component40_fa8_or0;
  wire [0:0] csa_component40_fa9_xor1;
  wire [0:0] csa_component40_fa9_or0;
  wire [0:0] csa_component40_fa10_xor1;
  wire [0:0] csa_component40_fa10_or0;
  wire [0:0] csa_component40_fa11_xor1;
  wire [0:0] csa_component40_fa11_or0;
  wire [0:0] csa_component40_fa12_xor1;
  wire [0:0] csa_component40_fa12_or0;
  wire [0:0] csa_component40_fa13_xor1;
  wire [0:0] csa_component40_fa13_or0;
  wire [0:0] csa_component40_fa14_xor1;
  wire [0:0] csa_component40_fa14_or0;
  wire [0:0] csa_component40_fa15_xor1;
  wire [0:0] csa_component40_fa15_or0;
  wire [0:0] csa_component40_fa16_xor1;
  wire [0:0] csa_component40_fa16_or0;
  wire [0:0] csa_component40_fa17_xor1;
  wire [0:0] csa_component40_fa17_or0;
  wire [0:0] csa_component40_fa18_xor1;
  wire [0:0] csa_component40_fa18_or0;
  wire [0:0] csa_component40_fa19_xor1;
  wire [0:0] csa_component40_fa19_or0;
  wire [0:0] csa_component40_fa20_xor1;
  wire [0:0] csa_component40_fa20_or0;
  wire [0:0] csa_component40_fa21_xor1;
  wire [0:0] csa_component40_fa21_or0;
  wire [0:0] csa_component40_fa22_xor1;
  wire [0:0] csa_component40_fa22_or0;
  wire [0:0] csa_component40_fa23_xor1;
  wire [0:0] csa_component40_fa23_or0;
  wire [0:0] csa_component40_fa24_xor1;
  wire [0:0] csa_component40_fa24_or0;
  wire [0:0] csa_component40_fa25_xor1;
  wire [0:0] csa_component40_fa25_or0;
  wire [0:0] csa_component40_fa26_xor1;
  wire [0:0] csa_component40_fa26_or0;
  wire [0:0] csa_component40_fa27_xor1;
  wire [0:0] csa_component40_fa27_or0;
  wire [0:0] csa_component40_fa28_xor1;
  wire [0:0] csa_component40_fa28_or0;
  wire [0:0] csa_component40_fa29_xor1;
  wire [0:0] csa_component40_fa29_or0;
  wire [0:0] csa_component40_fa30_xor1;
  wire [0:0] csa_component40_fa30_or0;
  wire [0:0] csa_component40_fa31_xor1;
  wire [0:0] csa_component40_fa31_or0;
  wire [0:0] csa_component40_fa32_xor1;
  wire [0:0] csa_component40_fa32_or0;
  wire [0:0] csa_component40_fa33_xor1;
  wire [0:0] csa_component40_fa33_or0;
  wire [0:0] csa_component40_fa34_xor1;
  wire [0:0] csa_component40_fa34_or0;
  wire [0:0] csa_component40_fa35_xor1;
  wire [0:0] csa_component40_fa35_or0;
  wire [0:0] csa_component40_fa36_xor1;
  wire [0:0] csa_component40_fa36_or0;
  wire [0:0] csa_component40_fa37_xor1;
  wire [0:0] csa_component40_fa37_or0;
  wire [0:0] csa_component40_fa38_xor1;
  wire [0:0] csa_component40_fa38_or0;
  wire [0:0] csa_component40_fa39_xor1;
  wire [0:0] csa_component40_fa39_or0;

  fa fa_csa_component40_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component40_fa0_xor1), .fa_or0(csa_component40_fa0_or0));
  fa fa_csa_component40_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component40_fa1_xor1), .fa_or0(csa_component40_fa1_or0));
  fa fa_csa_component40_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component40_fa2_xor1), .fa_or0(csa_component40_fa2_or0));
  fa fa_csa_component40_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component40_fa3_xor1), .fa_or0(csa_component40_fa3_or0));
  fa fa_csa_component40_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component40_fa4_xor1), .fa_or0(csa_component40_fa4_or0));
  fa fa_csa_component40_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component40_fa5_xor1), .fa_or0(csa_component40_fa5_or0));
  fa fa_csa_component40_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component40_fa6_xor1), .fa_or0(csa_component40_fa6_or0));
  fa fa_csa_component40_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component40_fa7_xor1), .fa_or0(csa_component40_fa7_or0));
  fa fa_csa_component40_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component40_fa8_xor1), .fa_or0(csa_component40_fa8_or0));
  fa fa_csa_component40_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component40_fa9_xor1), .fa_or0(csa_component40_fa9_or0));
  fa fa_csa_component40_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component40_fa10_xor1), .fa_or0(csa_component40_fa10_or0));
  fa fa_csa_component40_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component40_fa11_xor1), .fa_or0(csa_component40_fa11_or0));
  fa fa_csa_component40_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component40_fa12_xor1), .fa_or0(csa_component40_fa12_or0));
  fa fa_csa_component40_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component40_fa13_xor1), .fa_or0(csa_component40_fa13_or0));
  fa fa_csa_component40_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component40_fa14_xor1), .fa_or0(csa_component40_fa14_or0));
  fa fa_csa_component40_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component40_fa15_xor1), .fa_or0(csa_component40_fa15_or0));
  fa fa_csa_component40_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component40_fa16_xor1), .fa_or0(csa_component40_fa16_or0));
  fa fa_csa_component40_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component40_fa17_xor1), .fa_or0(csa_component40_fa17_or0));
  fa fa_csa_component40_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component40_fa18_xor1), .fa_or0(csa_component40_fa18_or0));
  fa fa_csa_component40_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component40_fa19_xor1), .fa_or0(csa_component40_fa19_or0));
  fa fa_csa_component40_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component40_fa20_xor1), .fa_or0(csa_component40_fa20_or0));
  fa fa_csa_component40_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component40_fa21_xor1), .fa_or0(csa_component40_fa21_or0));
  fa fa_csa_component40_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component40_fa22_xor1), .fa_or0(csa_component40_fa22_or0));
  fa fa_csa_component40_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component40_fa23_xor1), .fa_or0(csa_component40_fa23_or0));
  fa fa_csa_component40_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component40_fa24_xor1), .fa_or0(csa_component40_fa24_or0));
  fa fa_csa_component40_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component40_fa25_xor1), .fa_or0(csa_component40_fa25_or0));
  fa fa_csa_component40_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component40_fa26_xor1), .fa_or0(csa_component40_fa26_or0));
  fa fa_csa_component40_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component40_fa27_xor1), .fa_or0(csa_component40_fa27_or0));
  fa fa_csa_component40_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component40_fa28_xor1), .fa_or0(csa_component40_fa28_or0));
  fa fa_csa_component40_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component40_fa29_xor1), .fa_or0(csa_component40_fa29_or0));
  fa fa_csa_component40_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component40_fa30_xor1), .fa_or0(csa_component40_fa30_or0));
  fa fa_csa_component40_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component40_fa31_xor1), .fa_or0(csa_component40_fa31_or0));
  fa fa_csa_component40_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component40_fa32_xor1), .fa_or0(csa_component40_fa32_or0));
  fa fa_csa_component40_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component40_fa33_xor1), .fa_or0(csa_component40_fa33_or0));
  fa fa_csa_component40_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component40_fa34_xor1), .fa_or0(csa_component40_fa34_or0));
  fa fa_csa_component40_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component40_fa35_xor1), .fa_or0(csa_component40_fa35_or0));
  fa fa_csa_component40_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component40_fa36_xor1), .fa_or0(csa_component40_fa36_or0));
  fa fa_csa_component40_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component40_fa37_xor1), .fa_or0(csa_component40_fa37_or0));
  fa fa_csa_component40_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component40_fa38_xor1), .fa_or0(csa_component40_fa38_or0));
  fa fa_csa_component40_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component40_fa39_xor1), .fa_or0(csa_component40_fa39_or0));

  assign csa_component40_out[0] = csa_component40_fa0_xor1[0];
  assign csa_component40_out[1] = csa_component40_fa1_xor1[0];
  assign csa_component40_out[2] = csa_component40_fa2_xor1[0];
  assign csa_component40_out[3] = csa_component40_fa3_xor1[0];
  assign csa_component40_out[4] = csa_component40_fa4_xor1[0];
  assign csa_component40_out[5] = csa_component40_fa5_xor1[0];
  assign csa_component40_out[6] = csa_component40_fa6_xor1[0];
  assign csa_component40_out[7] = csa_component40_fa7_xor1[0];
  assign csa_component40_out[8] = csa_component40_fa8_xor1[0];
  assign csa_component40_out[9] = csa_component40_fa9_xor1[0];
  assign csa_component40_out[10] = csa_component40_fa10_xor1[0];
  assign csa_component40_out[11] = csa_component40_fa11_xor1[0];
  assign csa_component40_out[12] = csa_component40_fa12_xor1[0];
  assign csa_component40_out[13] = csa_component40_fa13_xor1[0];
  assign csa_component40_out[14] = csa_component40_fa14_xor1[0];
  assign csa_component40_out[15] = csa_component40_fa15_xor1[0];
  assign csa_component40_out[16] = csa_component40_fa16_xor1[0];
  assign csa_component40_out[17] = csa_component40_fa17_xor1[0];
  assign csa_component40_out[18] = csa_component40_fa18_xor1[0];
  assign csa_component40_out[19] = csa_component40_fa19_xor1[0];
  assign csa_component40_out[20] = csa_component40_fa20_xor1[0];
  assign csa_component40_out[21] = csa_component40_fa21_xor1[0];
  assign csa_component40_out[22] = csa_component40_fa22_xor1[0];
  assign csa_component40_out[23] = csa_component40_fa23_xor1[0];
  assign csa_component40_out[24] = csa_component40_fa24_xor1[0];
  assign csa_component40_out[25] = csa_component40_fa25_xor1[0];
  assign csa_component40_out[26] = csa_component40_fa26_xor1[0];
  assign csa_component40_out[27] = csa_component40_fa27_xor1[0];
  assign csa_component40_out[28] = csa_component40_fa28_xor1[0];
  assign csa_component40_out[29] = csa_component40_fa29_xor1[0];
  assign csa_component40_out[30] = csa_component40_fa30_xor1[0];
  assign csa_component40_out[31] = csa_component40_fa31_xor1[0];
  assign csa_component40_out[32] = csa_component40_fa32_xor1[0];
  assign csa_component40_out[33] = csa_component40_fa33_xor1[0];
  assign csa_component40_out[34] = csa_component40_fa34_xor1[0];
  assign csa_component40_out[35] = csa_component40_fa35_xor1[0];
  assign csa_component40_out[36] = csa_component40_fa36_xor1[0];
  assign csa_component40_out[37] = csa_component40_fa37_xor1[0];
  assign csa_component40_out[38] = csa_component40_fa38_xor1[0];
  assign csa_component40_out[39] = csa_component40_fa39_xor1[0];
  assign csa_component40_out[40] = 1'b0;
  assign csa_component40_out[41] = 1'b0;
  assign csa_component40_out[42] = csa_component40_fa0_or0[0];
  assign csa_component40_out[43] = csa_component40_fa1_or0[0];
  assign csa_component40_out[44] = csa_component40_fa2_or0[0];
  assign csa_component40_out[45] = csa_component40_fa3_or0[0];
  assign csa_component40_out[46] = csa_component40_fa4_or0[0];
  assign csa_component40_out[47] = csa_component40_fa5_or0[0];
  assign csa_component40_out[48] = csa_component40_fa6_or0[0];
  assign csa_component40_out[49] = csa_component40_fa7_or0[0];
  assign csa_component40_out[50] = csa_component40_fa8_or0[0];
  assign csa_component40_out[51] = csa_component40_fa9_or0[0];
  assign csa_component40_out[52] = csa_component40_fa10_or0[0];
  assign csa_component40_out[53] = csa_component40_fa11_or0[0];
  assign csa_component40_out[54] = csa_component40_fa12_or0[0];
  assign csa_component40_out[55] = csa_component40_fa13_or0[0];
  assign csa_component40_out[56] = csa_component40_fa14_or0[0];
  assign csa_component40_out[57] = csa_component40_fa15_or0[0];
  assign csa_component40_out[58] = csa_component40_fa16_or0[0];
  assign csa_component40_out[59] = csa_component40_fa17_or0[0];
  assign csa_component40_out[60] = csa_component40_fa18_or0[0];
  assign csa_component40_out[61] = csa_component40_fa19_or0[0];
  assign csa_component40_out[62] = csa_component40_fa20_or0[0];
  assign csa_component40_out[63] = csa_component40_fa21_or0[0];
  assign csa_component40_out[64] = csa_component40_fa22_or0[0];
  assign csa_component40_out[65] = csa_component40_fa23_or0[0];
  assign csa_component40_out[66] = csa_component40_fa24_or0[0];
  assign csa_component40_out[67] = csa_component40_fa25_or0[0];
  assign csa_component40_out[68] = csa_component40_fa26_or0[0];
  assign csa_component40_out[69] = csa_component40_fa27_or0[0];
  assign csa_component40_out[70] = csa_component40_fa28_or0[0];
  assign csa_component40_out[71] = csa_component40_fa29_or0[0];
  assign csa_component40_out[72] = csa_component40_fa30_or0[0];
  assign csa_component40_out[73] = csa_component40_fa31_or0[0];
  assign csa_component40_out[74] = csa_component40_fa32_or0[0];
  assign csa_component40_out[75] = csa_component40_fa33_or0[0];
  assign csa_component40_out[76] = csa_component40_fa34_or0[0];
  assign csa_component40_out[77] = csa_component40_fa35_or0[0];
  assign csa_component40_out[78] = csa_component40_fa36_or0[0];
  assign csa_component40_out[79] = csa_component40_fa37_or0[0];
  assign csa_component40_out[80] = csa_component40_fa38_or0[0];
  assign csa_component40_out[81] = csa_component40_fa39_or0[0];
endmodule

module u_cska48(input [47:0] a, input [47:0] b, output [48:0] u_cska48_out);
  wire [0:0] u_cska48_xor0;
  wire [0:0] u_cska48_ha0_xor0;
  wire [0:0] u_cska48_ha0_and0;
  wire [0:0] u_cska48_xor1;
  wire [0:0] u_cska48_fa0_xor1;
  wire [0:0] u_cska48_fa0_or0;
  wire [0:0] u_cska48_xor2;
  wire [0:0] u_cska48_fa1_xor1;
  wire [0:0] u_cska48_fa1_or0;
  wire [0:0] u_cska48_xor3;
  wire [0:0] u_cska48_fa2_xor1;
  wire [0:0] u_cska48_fa2_or0;
  wire [0:0] u_cska48_and_propagate00;
  wire [0:0] u_cska48_and_propagate01;
  wire [0:0] u_cska48_and_propagate02;
  wire [0:0] u_cska48_mux2to10_and1;
  wire [0:0] u_cska48_xor4;
  wire [0:0] u_cska48_fa3_xor1;
  wire [0:0] u_cska48_fa3_or0;
  wire [0:0] u_cska48_xor5;
  wire [0:0] u_cska48_fa4_xor1;
  wire [0:0] u_cska48_fa4_or0;
  wire [0:0] u_cska48_xor6;
  wire [0:0] u_cska48_fa5_xor1;
  wire [0:0] u_cska48_fa5_or0;
  wire [0:0] u_cska48_xor7;
  wire [0:0] u_cska48_fa6_xor1;
  wire [0:0] u_cska48_fa6_or0;
  wire [0:0] u_cska48_and_propagate13;
  wire [0:0] u_cska48_and_propagate14;
  wire [0:0] u_cska48_and_propagate15;
  wire [0:0] u_cska48_mux2to11_xor0;
  wire [0:0] u_cska48_xor8;
  wire [0:0] u_cska48_fa7_xor1;
  wire [0:0] u_cska48_fa7_or0;
  wire [0:0] u_cska48_xor9;
  wire [0:0] u_cska48_fa8_xor1;
  wire [0:0] u_cska48_fa8_or0;
  wire [0:0] u_cska48_xor10;
  wire [0:0] u_cska48_fa9_xor1;
  wire [0:0] u_cska48_fa9_or0;
  wire [0:0] u_cska48_xor11;
  wire [0:0] u_cska48_fa10_xor1;
  wire [0:0] u_cska48_fa10_or0;
  wire [0:0] u_cska48_and_propagate26;
  wire [0:0] u_cska48_and_propagate27;
  wire [0:0] u_cska48_and_propagate28;
  wire [0:0] u_cska48_mux2to12_xor0;
  wire [0:0] u_cska48_xor12;
  wire [0:0] u_cska48_fa11_xor1;
  wire [0:0] u_cska48_fa11_or0;
  wire [0:0] u_cska48_xor13;
  wire [0:0] u_cska48_fa12_xor1;
  wire [0:0] u_cska48_fa12_or0;
  wire [0:0] u_cska48_xor14;
  wire [0:0] u_cska48_fa13_xor1;
  wire [0:0] u_cska48_fa13_or0;
  wire [0:0] u_cska48_xor15;
  wire [0:0] u_cska48_fa14_xor1;
  wire [0:0] u_cska48_fa14_or0;
  wire [0:0] u_cska48_and_propagate39;
  wire [0:0] u_cska48_and_propagate310;
  wire [0:0] u_cska48_and_propagate311;
  wire [0:0] u_cska48_mux2to13_xor0;
  wire [0:0] u_cska48_xor16;
  wire [0:0] u_cska48_fa15_xor1;
  wire [0:0] u_cska48_fa15_or0;
  wire [0:0] u_cska48_xor17;
  wire [0:0] u_cska48_fa16_xor1;
  wire [0:0] u_cska48_fa16_or0;
  wire [0:0] u_cska48_xor18;
  wire [0:0] u_cska48_fa17_xor1;
  wire [0:0] u_cska48_fa17_or0;
  wire [0:0] u_cska48_xor19;
  wire [0:0] u_cska48_fa18_xor1;
  wire [0:0] u_cska48_fa18_or0;
  wire [0:0] u_cska48_and_propagate412;
  wire [0:0] u_cska48_and_propagate413;
  wire [0:0] u_cska48_and_propagate414;
  wire [0:0] u_cska48_mux2to14_xor0;
  wire [0:0] u_cska48_xor20;
  wire [0:0] u_cska48_fa19_xor1;
  wire [0:0] u_cska48_fa19_or0;
  wire [0:0] u_cska48_xor21;
  wire [0:0] u_cska48_fa20_xor1;
  wire [0:0] u_cska48_fa20_or0;
  wire [0:0] u_cska48_xor22;
  wire [0:0] u_cska48_fa21_xor1;
  wire [0:0] u_cska48_fa21_or0;
  wire [0:0] u_cska48_xor23;
  wire [0:0] u_cska48_fa22_xor1;
  wire [0:0] u_cska48_fa22_or0;
  wire [0:0] u_cska48_and_propagate515;
  wire [0:0] u_cska48_and_propagate516;
  wire [0:0] u_cska48_and_propagate517;
  wire [0:0] u_cska48_mux2to15_xor0;
  wire [0:0] u_cska48_xor24;
  wire [0:0] u_cska48_fa23_xor1;
  wire [0:0] u_cska48_fa23_or0;
  wire [0:0] u_cska48_xor25;
  wire [0:0] u_cska48_fa24_xor1;
  wire [0:0] u_cska48_fa24_or0;
  wire [0:0] u_cska48_xor26;
  wire [0:0] u_cska48_fa25_xor1;
  wire [0:0] u_cska48_fa25_or0;
  wire [0:0] u_cska48_xor27;
  wire [0:0] u_cska48_fa26_xor1;
  wire [0:0] u_cska48_fa26_or0;
  wire [0:0] u_cska48_and_propagate618;
  wire [0:0] u_cska48_and_propagate619;
  wire [0:0] u_cska48_and_propagate620;
  wire [0:0] u_cska48_mux2to16_xor0;
  wire [0:0] u_cska48_xor28;
  wire [0:0] u_cska48_fa27_xor1;
  wire [0:0] u_cska48_fa27_or0;
  wire [0:0] u_cska48_xor29;
  wire [0:0] u_cska48_fa28_xor1;
  wire [0:0] u_cska48_fa28_or0;
  wire [0:0] u_cska48_xor30;
  wire [0:0] u_cska48_fa29_xor1;
  wire [0:0] u_cska48_fa29_or0;
  wire [0:0] u_cska48_xor31;
  wire [0:0] u_cska48_fa30_xor1;
  wire [0:0] u_cska48_fa30_or0;
  wire [0:0] u_cska48_and_propagate721;
  wire [0:0] u_cska48_and_propagate722;
  wire [0:0] u_cska48_and_propagate723;
  wire [0:0] u_cska48_mux2to17_xor0;
  wire [0:0] u_cska48_xor32;
  wire [0:0] u_cska48_fa31_xor1;
  wire [0:0] u_cska48_fa31_or0;
  wire [0:0] u_cska48_xor33;
  wire [0:0] u_cska48_fa32_xor1;
  wire [0:0] u_cska48_fa32_or0;
  wire [0:0] u_cska48_xor34;
  wire [0:0] u_cska48_fa33_xor1;
  wire [0:0] u_cska48_fa33_or0;
  wire [0:0] u_cska48_xor35;
  wire [0:0] u_cska48_fa34_xor1;
  wire [0:0] u_cska48_fa34_or0;
  wire [0:0] u_cska48_and_propagate824;
  wire [0:0] u_cska48_and_propagate825;
  wire [0:0] u_cska48_and_propagate826;
  wire [0:0] u_cska48_mux2to18_xor0;
  wire [0:0] u_cska48_xor36;
  wire [0:0] u_cska48_fa35_xor1;
  wire [0:0] u_cska48_fa35_or0;
  wire [0:0] u_cska48_xor37;
  wire [0:0] u_cska48_fa36_xor1;
  wire [0:0] u_cska48_fa36_or0;
  wire [0:0] u_cska48_xor38;
  wire [0:0] u_cska48_fa37_xor1;
  wire [0:0] u_cska48_fa37_or0;
  wire [0:0] u_cska48_xor39;
  wire [0:0] u_cska48_fa38_xor1;
  wire [0:0] u_cska48_fa38_or0;
  wire [0:0] u_cska48_and_propagate927;
  wire [0:0] u_cska48_and_propagate928;
  wire [0:0] u_cska48_and_propagate929;
  wire [0:0] u_cska48_mux2to19_xor0;
  wire [0:0] u_cska48_xor40;
  wire [0:0] u_cska48_fa39_xor1;
  wire [0:0] u_cska48_fa39_or0;
  wire [0:0] u_cska48_xor41;
  wire [0:0] u_cska48_fa40_xor1;
  wire [0:0] u_cska48_fa40_or0;
  wire [0:0] u_cska48_xor42;
  wire [0:0] u_cska48_fa41_xor1;
  wire [0:0] u_cska48_fa41_or0;
  wire [0:0] u_cska48_xor43;
  wire [0:0] u_cska48_fa42_xor1;
  wire [0:0] u_cska48_fa42_or0;
  wire [0:0] u_cska48_and_propagate1030;
  wire [0:0] u_cska48_and_propagate1031;
  wire [0:0] u_cska48_and_propagate1032;
  wire [0:0] u_cska48_mux2to110_xor0;
  wire [0:0] u_cska48_xor44;
  wire [0:0] u_cska48_fa43_xor1;
  wire [0:0] u_cska48_fa43_or0;
  wire [0:0] u_cska48_xor45;
  wire [0:0] u_cska48_fa44_xor1;
  wire [0:0] u_cska48_fa44_or0;
  wire [0:0] u_cska48_xor46;
  wire [0:0] u_cska48_fa45_xor1;
  wire [0:0] u_cska48_fa45_or0;
  wire [0:0] u_cska48_xor47;
  wire [0:0] u_cska48_fa46_xor1;
  wire [0:0] u_cska48_fa46_or0;
  wire [0:0] u_cska48_and_propagate1133;
  wire [0:0] u_cska48_and_propagate1134;
  wire [0:0] u_cska48_and_propagate1135;
  wire [0:0] u_cska48_mux2to111_xor0;

  xor_gate xor_gate_u_cska48_xor0(.a(a[0]), .b(b[0]), .out(u_cska48_xor0));
  ha ha_u_cska48_ha0_out(.a(a[0]), .b(b[0]), .ha_xor0(u_cska48_ha0_xor0), .ha_and0(u_cska48_ha0_and0));
  xor_gate xor_gate_u_cska48_xor1(.a(a[1]), .b(b[1]), .out(u_cska48_xor1));
  fa fa_u_cska48_fa0_out(.a(a[1]), .b(b[1]), .cin(u_cska48_ha0_and0[0]), .fa_xor1(u_cska48_fa0_xor1), .fa_or0(u_cska48_fa0_or0));
  xor_gate xor_gate_u_cska48_xor2(.a(a[2]), .b(b[2]), .out(u_cska48_xor2));
  fa fa_u_cska48_fa1_out(.a(a[2]), .b(b[2]), .cin(u_cska48_fa0_or0[0]), .fa_xor1(u_cska48_fa1_xor1), .fa_or0(u_cska48_fa1_or0));
  xor_gate xor_gate_u_cska48_xor3(.a(a[3]), .b(b[3]), .out(u_cska48_xor3));
  fa fa_u_cska48_fa2_out(.a(a[3]), .b(b[3]), .cin(u_cska48_fa1_or0[0]), .fa_xor1(u_cska48_fa2_xor1), .fa_or0(u_cska48_fa2_or0));
  and_gate and_gate_u_cska48_and_propagate00(.a(u_cska48_xor0[0]), .b(u_cska48_xor2[0]), .out(u_cska48_and_propagate00));
  and_gate and_gate_u_cska48_and_propagate01(.a(u_cska48_xor1[0]), .b(u_cska48_xor3[0]), .out(u_cska48_and_propagate01));
  and_gate and_gate_u_cska48_and_propagate02(.a(u_cska48_and_propagate00[0]), .b(u_cska48_and_propagate01[0]), .out(u_cska48_and_propagate02));
  mux2to1 mux2to1_u_cska48_mux2to10_out(.d0(u_cska48_fa2_or0[0]), .d1(1'b0), .sel(u_cska48_and_propagate02[0]), .mux2to1_xor0(u_cska48_mux2to10_and1));
  xor_gate xor_gate_u_cska48_xor4(.a(a[4]), .b(b[4]), .out(u_cska48_xor4));
  fa fa_u_cska48_fa3_out(.a(a[4]), .b(b[4]), .cin(u_cska48_mux2to10_and1[0]), .fa_xor1(u_cska48_fa3_xor1), .fa_or0(u_cska48_fa3_or0));
  xor_gate xor_gate_u_cska48_xor5(.a(a[5]), .b(b[5]), .out(u_cska48_xor5));
  fa fa_u_cska48_fa4_out(.a(a[5]), .b(b[5]), .cin(u_cska48_fa3_or0[0]), .fa_xor1(u_cska48_fa4_xor1), .fa_or0(u_cska48_fa4_or0));
  xor_gate xor_gate_u_cska48_xor6(.a(a[6]), .b(b[6]), .out(u_cska48_xor6));
  fa fa_u_cska48_fa5_out(.a(a[6]), .b(b[6]), .cin(u_cska48_fa4_or0[0]), .fa_xor1(u_cska48_fa5_xor1), .fa_or0(u_cska48_fa5_or0));
  xor_gate xor_gate_u_cska48_xor7(.a(a[7]), .b(b[7]), .out(u_cska48_xor7));
  fa fa_u_cska48_fa6_out(.a(a[7]), .b(b[7]), .cin(u_cska48_fa5_or0[0]), .fa_xor1(u_cska48_fa6_xor1), .fa_or0(u_cska48_fa6_or0));
  and_gate and_gate_u_cska48_and_propagate13(.a(u_cska48_xor4[0]), .b(u_cska48_xor6[0]), .out(u_cska48_and_propagate13));
  and_gate and_gate_u_cska48_and_propagate14(.a(u_cska48_xor5[0]), .b(u_cska48_xor7[0]), .out(u_cska48_and_propagate14));
  and_gate and_gate_u_cska48_and_propagate15(.a(u_cska48_and_propagate13[0]), .b(u_cska48_and_propagate14[0]), .out(u_cska48_and_propagate15));
  mux2to1 mux2to1_u_cska48_mux2to11_out(.d0(u_cska48_fa6_or0[0]), .d1(u_cska48_mux2to10_and1[0]), .sel(u_cska48_and_propagate15[0]), .mux2to1_xor0(u_cska48_mux2to11_xor0));
  xor_gate xor_gate_u_cska48_xor8(.a(a[8]), .b(b[8]), .out(u_cska48_xor8));
  fa fa_u_cska48_fa7_out(.a(a[8]), .b(b[8]), .cin(u_cska48_mux2to11_xor0[0]), .fa_xor1(u_cska48_fa7_xor1), .fa_or0(u_cska48_fa7_or0));
  xor_gate xor_gate_u_cska48_xor9(.a(a[9]), .b(b[9]), .out(u_cska48_xor9));
  fa fa_u_cska48_fa8_out(.a(a[9]), .b(b[9]), .cin(u_cska48_fa7_or0[0]), .fa_xor1(u_cska48_fa8_xor1), .fa_or0(u_cska48_fa8_or0));
  xor_gate xor_gate_u_cska48_xor10(.a(a[10]), .b(b[10]), .out(u_cska48_xor10));
  fa fa_u_cska48_fa9_out(.a(a[10]), .b(b[10]), .cin(u_cska48_fa8_or0[0]), .fa_xor1(u_cska48_fa9_xor1), .fa_or0(u_cska48_fa9_or0));
  xor_gate xor_gate_u_cska48_xor11(.a(a[11]), .b(b[11]), .out(u_cska48_xor11));
  fa fa_u_cska48_fa10_out(.a(a[11]), .b(b[11]), .cin(u_cska48_fa9_or0[0]), .fa_xor1(u_cska48_fa10_xor1), .fa_or0(u_cska48_fa10_or0));
  and_gate and_gate_u_cska48_and_propagate26(.a(u_cska48_xor8[0]), .b(u_cska48_xor10[0]), .out(u_cska48_and_propagate26));
  and_gate and_gate_u_cska48_and_propagate27(.a(u_cska48_xor9[0]), .b(u_cska48_xor11[0]), .out(u_cska48_and_propagate27));
  and_gate and_gate_u_cska48_and_propagate28(.a(u_cska48_and_propagate26[0]), .b(u_cska48_and_propagate27[0]), .out(u_cska48_and_propagate28));
  mux2to1 mux2to1_u_cska48_mux2to12_out(.d0(u_cska48_fa10_or0[0]), .d1(u_cska48_mux2to11_xor0[0]), .sel(u_cska48_and_propagate28[0]), .mux2to1_xor0(u_cska48_mux2to12_xor0));
  xor_gate xor_gate_u_cska48_xor12(.a(a[12]), .b(b[12]), .out(u_cska48_xor12));
  fa fa_u_cska48_fa11_out(.a(a[12]), .b(b[12]), .cin(u_cska48_mux2to12_xor0[0]), .fa_xor1(u_cska48_fa11_xor1), .fa_or0(u_cska48_fa11_or0));
  xor_gate xor_gate_u_cska48_xor13(.a(a[13]), .b(b[13]), .out(u_cska48_xor13));
  fa fa_u_cska48_fa12_out(.a(a[13]), .b(b[13]), .cin(u_cska48_fa11_or0[0]), .fa_xor1(u_cska48_fa12_xor1), .fa_or0(u_cska48_fa12_or0));
  xor_gate xor_gate_u_cska48_xor14(.a(a[14]), .b(b[14]), .out(u_cska48_xor14));
  fa fa_u_cska48_fa13_out(.a(a[14]), .b(b[14]), .cin(u_cska48_fa12_or0[0]), .fa_xor1(u_cska48_fa13_xor1), .fa_or0(u_cska48_fa13_or0));
  xor_gate xor_gate_u_cska48_xor15(.a(a[15]), .b(b[15]), .out(u_cska48_xor15));
  fa fa_u_cska48_fa14_out(.a(a[15]), .b(b[15]), .cin(u_cska48_fa13_or0[0]), .fa_xor1(u_cska48_fa14_xor1), .fa_or0(u_cska48_fa14_or0));
  and_gate and_gate_u_cska48_and_propagate39(.a(u_cska48_xor12[0]), .b(u_cska48_xor14[0]), .out(u_cska48_and_propagate39));
  and_gate and_gate_u_cska48_and_propagate310(.a(u_cska48_xor13[0]), .b(u_cska48_xor15[0]), .out(u_cska48_and_propagate310));
  and_gate and_gate_u_cska48_and_propagate311(.a(u_cska48_and_propagate39[0]), .b(u_cska48_and_propagate310[0]), .out(u_cska48_and_propagate311));
  mux2to1 mux2to1_u_cska48_mux2to13_out(.d0(u_cska48_fa14_or0[0]), .d1(u_cska48_mux2to12_xor0[0]), .sel(u_cska48_and_propagate311[0]), .mux2to1_xor0(u_cska48_mux2to13_xor0));
  xor_gate xor_gate_u_cska48_xor16(.a(a[16]), .b(b[16]), .out(u_cska48_xor16));
  fa fa_u_cska48_fa15_out(.a(a[16]), .b(b[16]), .cin(u_cska48_mux2to13_xor0[0]), .fa_xor1(u_cska48_fa15_xor1), .fa_or0(u_cska48_fa15_or0));
  xor_gate xor_gate_u_cska48_xor17(.a(a[17]), .b(b[17]), .out(u_cska48_xor17));
  fa fa_u_cska48_fa16_out(.a(a[17]), .b(b[17]), .cin(u_cska48_fa15_or0[0]), .fa_xor1(u_cska48_fa16_xor1), .fa_or0(u_cska48_fa16_or0));
  xor_gate xor_gate_u_cska48_xor18(.a(a[18]), .b(b[18]), .out(u_cska48_xor18));
  fa fa_u_cska48_fa17_out(.a(a[18]), .b(b[18]), .cin(u_cska48_fa16_or0[0]), .fa_xor1(u_cska48_fa17_xor1), .fa_or0(u_cska48_fa17_or0));
  xor_gate xor_gate_u_cska48_xor19(.a(a[19]), .b(b[19]), .out(u_cska48_xor19));
  fa fa_u_cska48_fa18_out(.a(a[19]), .b(b[19]), .cin(u_cska48_fa17_or0[0]), .fa_xor1(u_cska48_fa18_xor1), .fa_or0(u_cska48_fa18_or0));
  and_gate and_gate_u_cska48_and_propagate412(.a(u_cska48_xor16[0]), .b(u_cska48_xor18[0]), .out(u_cska48_and_propagate412));
  and_gate and_gate_u_cska48_and_propagate413(.a(u_cska48_xor17[0]), .b(u_cska48_xor19[0]), .out(u_cska48_and_propagate413));
  and_gate and_gate_u_cska48_and_propagate414(.a(u_cska48_and_propagate412[0]), .b(u_cska48_and_propagate413[0]), .out(u_cska48_and_propagate414));
  mux2to1 mux2to1_u_cska48_mux2to14_out(.d0(u_cska48_fa18_or0[0]), .d1(u_cska48_mux2to13_xor0[0]), .sel(u_cska48_and_propagate414[0]), .mux2to1_xor0(u_cska48_mux2to14_xor0));
  xor_gate xor_gate_u_cska48_xor20(.a(a[20]), .b(b[20]), .out(u_cska48_xor20));
  fa fa_u_cska48_fa19_out(.a(a[20]), .b(b[20]), .cin(u_cska48_mux2to14_xor0[0]), .fa_xor1(u_cska48_fa19_xor1), .fa_or0(u_cska48_fa19_or0));
  xor_gate xor_gate_u_cska48_xor21(.a(a[21]), .b(b[21]), .out(u_cska48_xor21));
  fa fa_u_cska48_fa20_out(.a(a[21]), .b(b[21]), .cin(u_cska48_fa19_or0[0]), .fa_xor1(u_cska48_fa20_xor1), .fa_or0(u_cska48_fa20_or0));
  xor_gate xor_gate_u_cska48_xor22(.a(a[22]), .b(b[22]), .out(u_cska48_xor22));
  fa fa_u_cska48_fa21_out(.a(a[22]), .b(b[22]), .cin(u_cska48_fa20_or0[0]), .fa_xor1(u_cska48_fa21_xor1), .fa_or0(u_cska48_fa21_or0));
  xor_gate xor_gate_u_cska48_xor23(.a(a[23]), .b(b[23]), .out(u_cska48_xor23));
  fa fa_u_cska48_fa22_out(.a(a[23]), .b(b[23]), .cin(u_cska48_fa21_or0[0]), .fa_xor1(u_cska48_fa22_xor1), .fa_or0(u_cska48_fa22_or0));
  and_gate and_gate_u_cska48_and_propagate515(.a(u_cska48_xor20[0]), .b(u_cska48_xor22[0]), .out(u_cska48_and_propagate515));
  and_gate and_gate_u_cska48_and_propagate516(.a(u_cska48_xor21[0]), .b(u_cska48_xor23[0]), .out(u_cska48_and_propagate516));
  and_gate and_gate_u_cska48_and_propagate517(.a(u_cska48_and_propagate515[0]), .b(u_cska48_and_propagate516[0]), .out(u_cska48_and_propagate517));
  mux2to1 mux2to1_u_cska48_mux2to15_out(.d0(u_cska48_fa22_or0[0]), .d1(u_cska48_mux2to14_xor0[0]), .sel(u_cska48_and_propagate517[0]), .mux2to1_xor0(u_cska48_mux2to15_xor0));
  xor_gate xor_gate_u_cska48_xor24(.a(a[24]), .b(b[24]), .out(u_cska48_xor24));
  fa fa_u_cska48_fa23_out(.a(a[24]), .b(b[24]), .cin(u_cska48_mux2to15_xor0[0]), .fa_xor1(u_cska48_fa23_xor1), .fa_or0(u_cska48_fa23_or0));
  xor_gate xor_gate_u_cska48_xor25(.a(a[25]), .b(b[25]), .out(u_cska48_xor25));
  fa fa_u_cska48_fa24_out(.a(a[25]), .b(b[25]), .cin(u_cska48_fa23_or0[0]), .fa_xor1(u_cska48_fa24_xor1), .fa_or0(u_cska48_fa24_or0));
  xor_gate xor_gate_u_cska48_xor26(.a(a[26]), .b(b[26]), .out(u_cska48_xor26));
  fa fa_u_cska48_fa25_out(.a(a[26]), .b(b[26]), .cin(u_cska48_fa24_or0[0]), .fa_xor1(u_cska48_fa25_xor1), .fa_or0(u_cska48_fa25_or0));
  xor_gate xor_gate_u_cska48_xor27(.a(a[27]), .b(b[27]), .out(u_cska48_xor27));
  fa fa_u_cska48_fa26_out(.a(a[27]), .b(b[27]), .cin(u_cska48_fa25_or0[0]), .fa_xor1(u_cska48_fa26_xor1), .fa_or0(u_cska48_fa26_or0));
  and_gate and_gate_u_cska48_and_propagate618(.a(u_cska48_xor24[0]), .b(u_cska48_xor26[0]), .out(u_cska48_and_propagate618));
  and_gate and_gate_u_cska48_and_propagate619(.a(u_cska48_xor25[0]), .b(u_cska48_xor27[0]), .out(u_cska48_and_propagate619));
  and_gate and_gate_u_cska48_and_propagate620(.a(u_cska48_and_propagate618[0]), .b(u_cska48_and_propagate619[0]), .out(u_cska48_and_propagate620));
  mux2to1 mux2to1_u_cska48_mux2to16_out(.d0(u_cska48_fa26_or0[0]), .d1(u_cska48_mux2to15_xor0[0]), .sel(u_cska48_and_propagate620[0]), .mux2to1_xor0(u_cska48_mux2to16_xor0));
  xor_gate xor_gate_u_cska48_xor28(.a(a[28]), .b(b[28]), .out(u_cska48_xor28));
  fa fa_u_cska48_fa27_out(.a(a[28]), .b(b[28]), .cin(u_cska48_mux2to16_xor0[0]), .fa_xor1(u_cska48_fa27_xor1), .fa_or0(u_cska48_fa27_or0));
  xor_gate xor_gate_u_cska48_xor29(.a(a[29]), .b(b[29]), .out(u_cska48_xor29));
  fa fa_u_cska48_fa28_out(.a(a[29]), .b(b[29]), .cin(u_cska48_fa27_or0[0]), .fa_xor1(u_cska48_fa28_xor1), .fa_or0(u_cska48_fa28_or0));
  xor_gate xor_gate_u_cska48_xor30(.a(a[30]), .b(b[30]), .out(u_cska48_xor30));
  fa fa_u_cska48_fa29_out(.a(a[30]), .b(b[30]), .cin(u_cska48_fa28_or0[0]), .fa_xor1(u_cska48_fa29_xor1), .fa_or0(u_cska48_fa29_or0));
  xor_gate xor_gate_u_cska48_xor31(.a(a[31]), .b(b[31]), .out(u_cska48_xor31));
  fa fa_u_cska48_fa30_out(.a(a[31]), .b(b[31]), .cin(u_cska48_fa29_or0[0]), .fa_xor1(u_cska48_fa30_xor1), .fa_or0(u_cska48_fa30_or0));
  and_gate and_gate_u_cska48_and_propagate721(.a(u_cska48_xor28[0]), .b(u_cska48_xor30[0]), .out(u_cska48_and_propagate721));
  and_gate and_gate_u_cska48_and_propagate722(.a(u_cska48_xor29[0]), .b(u_cska48_xor31[0]), .out(u_cska48_and_propagate722));
  and_gate and_gate_u_cska48_and_propagate723(.a(u_cska48_and_propagate721[0]), .b(u_cska48_and_propagate722[0]), .out(u_cska48_and_propagate723));
  mux2to1 mux2to1_u_cska48_mux2to17_out(.d0(u_cska48_fa30_or0[0]), .d1(u_cska48_mux2to16_xor0[0]), .sel(u_cska48_and_propagate723[0]), .mux2to1_xor0(u_cska48_mux2to17_xor0));
  xor_gate xor_gate_u_cska48_xor32(.a(a[32]), .b(b[32]), .out(u_cska48_xor32));
  fa fa_u_cska48_fa31_out(.a(a[32]), .b(b[32]), .cin(u_cska48_mux2to17_xor0[0]), .fa_xor1(u_cska48_fa31_xor1), .fa_or0(u_cska48_fa31_or0));
  xor_gate xor_gate_u_cska48_xor33(.a(a[33]), .b(b[33]), .out(u_cska48_xor33));
  fa fa_u_cska48_fa32_out(.a(a[33]), .b(b[33]), .cin(u_cska48_fa31_or0[0]), .fa_xor1(u_cska48_fa32_xor1), .fa_or0(u_cska48_fa32_or0));
  xor_gate xor_gate_u_cska48_xor34(.a(a[34]), .b(b[34]), .out(u_cska48_xor34));
  fa fa_u_cska48_fa33_out(.a(a[34]), .b(b[34]), .cin(u_cska48_fa32_or0[0]), .fa_xor1(u_cska48_fa33_xor1), .fa_or0(u_cska48_fa33_or0));
  xor_gate xor_gate_u_cska48_xor35(.a(a[35]), .b(b[35]), .out(u_cska48_xor35));
  fa fa_u_cska48_fa34_out(.a(a[35]), .b(b[35]), .cin(u_cska48_fa33_or0[0]), .fa_xor1(u_cska48_fa34_xor1), .fa_or0(u_cska48_fa34_or0));
  and_gate and_gate_u_cska48_and_propagate824(.a(u_cska48_xor32[0]), .b(u_cska48_xor34[0]), .out(u_cska48_and_propagate824));
  and_gate and_gate_u_cska48_and_propagate825(.a(u_cska48_xor33[0]), .b(u_cska48_xor35[0]), .out(u_cska48_and_propagate825));
  and_gate and_gate_u_cska48_and_propagate826(.a(u_cska48_and_propagate824[0]), .b(u_cska48_and_propagate825[0]), .out(u_cska48_and_propagate826));
  mux2to1 mux2to1_u_cska48_mux2to18_out(.d0(u_cska48_fa34_or0[0]), .d1(u_cska48_mux2to17_xor0[0]), .sel(u_cska48_and_propagate826[0]), .mux2to1_xor0(u_cska48_mux2to18_xor0));
  xor_gate xor_gate_u_cska48_xor36(.a(a[36]), .b(b[36]), .out(u_cska48_xor36));
  fa fa_u_cska48_fa35_out(.a(a[36]), .b(b[36]), .cin(u_cska48_mux2to18_xor0[0]), .fa_xor1(u_cska48_fa35_xor1), .fa_or0(u_cska48_fa35_or0));
  xor_gate xor_gate_u_cska48_xor37(.a(a[37]), .b(b[37]), .out(u_cska48_xor37));
  fa fa_u_cska48_fa36_out(.a(a[37]), .b(b[37]), .cin(u_cska48_fa35_or0[0]), .fa_xor1(u_cska48_fa36_xor1), .fa_or0(u_cska48_fa36_or0));
  xor_gate xor_gate_u_cska48_xor38(.a(a[38]), .b(b[38]), .out(u_cska48_xor38));
  fa fa_u_cska48_fa37_out(.a(a[38]), .b(b[38]), .cin(u_cska48_fa36_or0[0]), .fa_xor1(u_cska48_fa37_xor1), .fa_or0(u_cska48_fa37_or0));
  xor_gate xor_gate_u_cska48_xor39(.a(a[39]), .b(b[39]), .out(u_cska48_xor39));
  fa fa_u_cska48_fa38_out(.a(a[39]), .b(b[39]), .cin(u_cska48_fa37_or0[0]), .fa_xor1(u_cska48_fa38_xor1), .fa_or0(u_cska48_fa38_or0));
  and_gate and_gate_u_cska48_and_propagate927(.a(u_cska48_xor36[0]), .b(u_cska48_xor38[0]), .out(u_cska48_and_propagate927));
  and_gate and_gate_u_cska48_and_propagate928(.a(u_cska48_xor37[0]), .b(u_cska48_xor39[0]), .out(u_cska48_and_propagate928));
  and_gate and_gate_u_cska48_and_propagate929(.a(u_cska48_and_propagate927[0]), .b(u_cska48_and_propagate928[0]), .out(u_cska48_and_propagate929));
  mux2to1 mux2to1_u_cska48_mux2to19_out(.d0(u_cska48_fa38_or0[0]), .d1(u_cska48_mux2to18_xor0[0]), .sel(u_cska48_and_propagate929[0]), .mux2to1_xor0(u_cska48_mux2to19_xor0));
  xor_gate xor_gate_u_cska48_xor40(.a(a[40]), .b(b[40]), .out(u_cska48_xor40));
  fa fa_u_cska48_fa39_out(.a(a[40]), .b(b[40]), .cin(u_cska48_mux2to19_xor0[0]), .fa_xor1(u_cska48_fa39_xor1), .fa_or0(u_cska48_fa39_or0));
  xor_gate xor_gate_u_cska48_xor41(.a(a[41]), .b(b[41]), .out(u_cska48_xor41));
  fa fa_u_cska48_fa40_out(.a(a[41]), .b(b[41]), .cin(u_cska48_fa39_or0[0]), .fa_xor1(u_cska48_fa40_xor1), .fa_or0(u_cska48_fa40_or0));
  xor_gate xor_gate_u_cska48_xor42(.a(a[42]), .b(b[42]), .out(u_cska48_xor42));
  fa fa_u_cska48_fa41_out(.a(a[42]), .b(b[42]), .cin(u_cska48_fa40_or0[0]), .fa_xor1(u_cska48_fa41_xor1), .fa_or0(u_cska48_fa41_or0));
  xor_gate xor_gate_u_cska48_xor43(.a(a[43]), .b(b[43]), .out(u_cska48_xor43));
  fa fa_u_cska48_fa42_out(.a(a[43]), .b(b[43]), .cin(u_cska48_fa41_or0[0]), .fa_xor1(u_cska48_fa42_xor1), .fa_or0(u_cska48_fa42_or0));
  and_gate and_gate_u_cska48_and_propagate1030(.a(u_cska48_xor40[0]), .b(u_cska48_xor42[0]), .out(u_cska48_and_propagate1030));
  and_gate and_gate_u_cska48_and_propagate1031(.a(u_cska48_xor41[0]), .b(u_cska48_xor43[0]), .out(u_cska48_and_propagate1031));
  and_gate and_gate_u_cska48_and_propagate1032(.a(u_cska48_and_propagate1030[0]), .b(u_cska48_and_propagate1031[0]), .out(u_cska48_and_propagate1032));
  mux2to1 mux2to1_u_cska48_mux2to110_out(.d0(u_cska48_fa42_or0[0]), .d1(u_cska48_mux2to19_xor0[0]), .sel(u_cska48_and_propagate1032[0]), .mux2to1_xor0(u_cska48_mux2to110_xor0));
  xor_gate xor_gate_u_cska48_xor44(.a(a[44]), .b(b[44]), .out(u_cska48_xor44));
  fa fa_u_cska48_fa43_out(.a(a[44]), .b(b[44]), .cin(u_cska48_mux2to110_xor0[0]), .fa_xor1(u_cska48_fa43_xor1), .fa_or0(u_cska48_fa43_or0));
  xor_gate xor_gate_u_cska48_xor45(.a(a[45]), .b(b[45]), .out(u_cska48_xor45));
  fa fa_u_cska48_fa44_out(.a(a[45]), .b(b[45]), .cin(u_cska48_fa43_or0[0]), .fa_xor1(u_cska48_fa44_xor1), .fa_or0(u_cska48_fa44_or0));
  xor_gate xor_gate_u_cska48_xor46(.a(a[46]), .b(b[46]), .out(u_cska48_xor46));
  fa fa_u_cska48_fa45_out(.a(a[46]), .b(b[46]), .cin(u_cska48_fa44_or0[0]), .fa_xor1(u_cska48_fa45_xor1), .fa_or0(u_cska48_fa45_or0));
  xor_gate xor_gate_u_cska48_xor47(.a(a[47]), .b(b[47]), .out(u_cska48_xor47));
  fa fa_u_cska48_fa46_out(.a(a[47]), .b(b[47]), .cin(u_cska48_fa45_or0[0]), .fa_xor1(u_cska48_fa46_xor1), .fa_or0(u_cska48_fa46_or0));
  and_gate and_gate_u_cska48_and_propagate1133(.a(u_cska48_xor44[0]), .b(u_cska48_xor46[0]), .out(u_cska48_and_propagate1133));
  and_gate and_gate_u_cska48_and_propagate1134(.a(u_cska48_xor45[0]), .b(u_cska48_xor47[0]), .out(u_cska48_and_propagate1134));
  and_gate and_gate_u_cska48_and_propagate1135(.a(u_cska48_and_propagate1133[0]), .b(u_cska48_and_propagate1134[0]), .out(u_cska48_and_propagate1135));
  mux2to1 mux2to1_u_cska48_mux2to111_out(.d0(u_cska48_fa46_or0[0]), .d1(u_cska48_mux2to110_xor0[0]), .sel(u_cska48_and_propagate1135[0]), .mux2to1_xor0(u_cska48_mux2to111_xor0));

  assign u_cska48_out[0] = u_cska48_ha0_xor0[0];
  assign u_cska48_out[1] = u_cska48_fa0_xor1[0];
  assign u_cska48_out[2] = u_cska48_fa1_xor1[0];
  assign u_cska48_out[3] = u_cska48_fa2_xor1[0];
  assign u_cska48_out[4] = u_cska48_fa3_xor1[0];
  assign u_cska48_out[5] = u_cska48_fa4_xor1[0];
  assign u_cska48_out[6] = u_cska48_fa5_xor1[0];
  assign u_cska48_out[7] = u_cska48_fa6_xor1[0];
  assign u_cska48_out[8] = u_cska48_fa7_xor1[0];
  assign u_cska48_out[9] = u_cska48_fa8_xor1[0];
  assign u_cska48_out[10] = u_cska48_fa9_xor1[0];
  assign u_cska48_out[11] = u_cska48_fa10_xor1[0];
  assign u_cska48_out[12] = u_cska48_fa11_xor1[0];
  assign u_cska48_out[13] = u_cska48_fa12_xor1[0];
  assign u_cska48_out[14] = u_cska48_fa13_xor1[0];
  assign u_cska48_out[15] = u_cska48_fa14_xor1[0];
  assign u_cska48_out[16] = u_cska48_fa15_xor1[0];
  assign u_cska48_out[17] = u_cska48_fa16_xor1[0];
  assign u_cska48_out[18] = u_cska48_fa17_xor1[0];
  assign u_cska48_out[19] = u_cska48_fa18_xor1[0];
  assign u_cska48_out[20] = u_cska48_fa19_xor1[0];
  assign u_cska48_out[21] = u_cska48_fa20_xor1[0];
  assign u_cska48_out[22] = u_cska48_fa21_xor1[0];
  assign u_cska48_out[23] = u_cska48_fa22_xor1[0];
  assign u_cska48_out[24] = u_cska48_fa23_xor1[0];
  assign u_cska48_out[25] = u_cska48_fa24_xor1[0];
  assign u_cska48_out[26] = u_cska48_fa25_xor1[0];
  assign u_cska48_out[27] = u_cska48_fa26_xor1[0];
  assign u_cska48_out[28] = u_cska48_fa27_xor1[0];
  assign u_cska48_out[29] = u_cska48_fa28_xor1[0];
  assign u_cska48_out[30] = u_cska48_fa29_xor1[0];
  assign u_cska48_out[31] = u_cska48_fa30_xor1[0];
  assign u_cska48_out[32] = u_cska48_fa31_xor1[0];
  assign u_cska48_out[33] = u_cska48_fa32_xor1[0];
  assign u_cska48_out[34] = u_cska48_fa33_xor1[0];
  assign u_cska48_out[35] = u_cska48_fa34_xor1[0];
  assign u_cska48_out[36] = u_cska48_fa35_xor1[0];
  assign u_cska48_out[37] = u_cska48_fa36_xor1[0];
  assign u_cska48_out[38] = u_cska48_fa37_xor1[0];
  assign u_cska48_out[39] = u_cska48_fa38_xor1[0];
  assign u_cska48_out[40] = u_cska48_fa39_xor1[0];
  assign u_cska48_out[41] = u_cska48_fa40_xor1[0];
  assign u_cska48_out[42] = u_cska48_fa41_xor1[0];
  assign u_cska48_out[43] = u_cska48_fa42_xor1[0];
  assign u_cska48_out[44] = u_cska48_fa43_xor1[0];
  assign u_cska48_out[45] = u_cska48_fa44_xor1[0];
  assign u_cska48_out[46] = u_cska48_fa45_xor1[0];
  assign u_cska48_out[47] = u_cska48_fa46_xor1[0];
  assign u_cska48_out[48] = u_cska48_mux2to111_xor0[0];
endmodule

module s_CSAwallace_cska24(input [23:0] a, input [23:0] b, output [47:0] s_CSAwallace_cska24_out);
  wire [0:0] s_CSAwallace_cska24_and_0_0;
  wire [0:0] s_CSAwallace_cska24_and_1_0;
  wire [0:0] s_CSAwallace_cska24_and_2_0;
  wire [0:0] s_CSAwallace_cska24_and_3_0;
  wire [0:0] s_CSAwallace_cska24_and_4_0;
  wire [0:0] s_CSAwallace_cska24_and_5_0;
  wire [0:0] s_CSAwallace_cska24_and_6_0;
  wire [0:0] s_CSAwallace_cska24_and_7_0;
  wire [0:0] s_CSAwallace_cska24_and_8_0;
  wire [0:0] s_CSAwallace_cska24_and_9_0;
  wire [0:0] s_CSAwallace_cska24_and_10_0;
  wire [0:0] s_CSAwallace_cska24_and_11_0;
  wire [0:0] s_CSAwallace_cska24_and_12_0;
  wire [0:0] s_CSAwallace_cska24_and_13_0;
  wire [0:0] s_CSAwallace_cska24_and_14_0;
  wire [0:0] s_CSAwallace_cska24_and_15_0;
  wire [0:0] s_CSAwallace_cska24_and_16_0;
  wire [0:0] s_CSAwallace_cska24_and_17_0;
  wire [0:0] s_CSAwallace_cska24_and_18_0;
  wire [0:0] s_CSAwallace_cska24_and_19_0;
  wire [0:0] s_CSAwallace_cska24_and_20_0;
  wire [0:0] s_CSAwallace_cska24_and_21_0;
  wire [0:0] s_CSAwallace_cska24_and_22_0;
  wire [0:0] s_CSAwallace_cska24_nand_23_0;
  wire [0:0] s_CSAwallace_cska24_and_0_1;
  wire [0:0] s_CSAwallace_cska24_and_1_1;
  wire [0:0] s_CSAwallace_cska24_and_2_1;
  wire [0:0] s_CSAwallace_cska24_and_3_1;
  wire [0:0] s_CSAwallace_cska24_and_4_1;
  wire [0:0] s_CSAwallace_cska24_and_5_1;
  wire [0:0] s_CSAwallace_cska24_and_6_1;
  wire [0:0] s_CSAwallace_cska24_and_7_1;
  wire [0:0] s_CSAwallace_cska24_and_8_1;
  wire [0:0] s_CSAwallace_cska24_and_9_1;
  wire [0:0] s_CSAwallace_cska24_and_10_1;
  wire [0:0] s_CSAwallace_cska24_and_11_1;
  wire [0:0] s_CSAwallace_cska24_and_12_1;
  wire [0:0] s_CSAwallace_cska24_and_13_1;
  wire [0:0] s_CSAwallace_cska24_and_14_1;
  wire [0:0] s_CSAwallace_cska24_and_15_1;
  wire [0:0] s_CSAwallace_cska24_and_16_1;
  wire [0:0] s_CSAwallace_cska24_and_17_1;
  wire [0:0] s_CSAwallace_cska24_and_18_1;
  wire [0:0] s_CSAwallace_cska24_and_19_1;
  wire [0:0] s_CSAwallace_cska24_and_20_1;
  wire [0:0] s_CSAwallace_cska24_and_21_1;
  wire [0:0] s_CSAwallace_cska24_and_22_1;
  wire [0:0] s_CSAwallace_cska24_nand_23_1;
  wire [0:0] s_CSAwallace_cska24_and_0_2;
  wire [0:0] s_CSAwallace_cska24_and_1_2;
  wire [0:0] s_CSAwallace_cska24_and_2_2;
  wire [0:0] s_CSAwallace_cska24_and_3_2;
  wire [0:0] s_CSAwallace_cska24_and_4_2;
  wire [0:0] s_CSAwallace_cska24_and_5_2;
  wire [0:0] s_CSAwallace_cska24_and_6_2;
  wire [0:0] s_CSAwallace_cska24_and_7_2;
  wire [0:0] s_CSAwallace_cska24_and_8_2;
  wire [0:0] s_CSAwallace_cska24_and_9_2;
  wire [0:0] s_CSAwallace_cska24_and_10_2;
  wire [0:0] s_CSAwallace_cska24_and_11_2;
  wire [0:0] s_CSAwallace_cska24_and_12_2;
  wire [0:0] s_CSAwallace_cska24_and_13_2;
  wire [0:0] s_CSAwallace_cska24_and_14_2;
  wire [0:0] s_CSAwallace_cska24_and_15_2;
  wire [0:0] s_CSAwallace_cska24_and_16_2;
  wire [0:0] s_CSAwallace_cska24_and_17_2;
  wire [0:0] s_CSAwallace_cska24_and_18_2;
  wire [0:0] s_CSAwallace_cska24_and_19_2;
  wire [0:0] s_CSAwallace_cska24_and_20_2;
  wire [0:0] s_CSAwallace_cska24_and_21_2;
  wire [0:0] s_CSAwallace_cska24_and_22_2;
  wire [0:0] s_CSAwallace_cska24_nand_23_2;
  wire [0:0] s_CSAwallace_cska24_and_0_3;
  wire [0:0] s_CSAwallace_cska24_and_1_3;
  wire [0:0] s_CSAwallace_cska24_and_2_3;
  wire [0:0] s_CSAwallace_cska24_and_3_3;
  wire [0:0] s_CSAwallace_cska24_and_4_3;
  wire [0:0] s_CSAwallace_cska24_and_5_3;
  wire [0:0] s_CSAwallace_cska24_and_6_3;
  wire [0:0] s_CSAwallace_cska24_and_7_3;
  wire [0:0] s_CSAwallace_cska24_and_8_3;
  wire [0:0] s_CSAwallace_cska24_and_9_3;
  wire [0:0] s_CSAwallace_cska24_and_10_3;
  wire [0:0] s_CSAwallace_cska24_and_11_3;
  wire [0:0] s_CSAwallace_cska24_and_12_3;
  wire [0:0] s_CSAwallace_cska24_and_13_3;
  wire [0:0] s_CSAwallace_cska24_and_14_3;
  wire [0:0] s_CSAwallace_cska24_and_15_3;
  wire [0:0] s_CSAwallace_cska24_and_16_3;
  wire [0:0] s_CSAwallace_cska24_and_17_3;
  wire [0:0] s_CSAwallace_cska24_and_18_3;
  wire [0:0] s_CSAwallace_cska24_and_19_3;
  wire [0:0] s_CSAwallace_cska24_and_20_3;
  wire [0:0] s_CSAwallace_cska24_and_21_3;
  wire [0:0] s_CSAwallace_cska24_and_22_3;
  wire [0:0] s_CSAwallace_cska24_nand_23_3;
  wire [0:0] s_CSAwallace_cska24_and_0_4;
  wire [0:0] s_CSAwallace_cska24_and_1_4;
  wire [0:0] s_CSAwallace_cska24_and_2_4;
  wire [0:0] s_CSAwallace_cska24_and_3_4;
  wire [0:0] s_CSAwallace_cska24_and_4_4;
  wire [0:0] s_CSAwallace_cska24_and_5_4;
  wire [0:0] s_CSAwallace_cska24_and_6_4;
  wire [0:0] s_CSAwallace_cska24_and_7_4;
  wire [0:0] s_CSAwallace_cska24_and_8_4;
  wire [0:0] s_CSAwallace_cska24_and_9_4;
  wire [0:0] s_CSAwallace_cska24_and_10_4;
  wire [0:0] s_CSAwallace_cska24_and_11_4;
  wire [0:0] s_CSAwallace_cska24_and_12_4;
  wire [0:0] s_CSAwallace_cska24_and_13_4;
  wire [0:0] s_CSAwallace_cska24_and_14_4;
  wire [0:0] s_CSAwallace_cska24_and_15_4;
  wire [0:0] s_CSAwallace_cska24_and_16_4;
  wire [0:0] s_CSAwallace_cska24_and_17_4;
  wire [0:0] s_CSAwallace_cska24_and_18_4;
  wire [0:0] s_CSAwallace_cska24_and_19_4;
  wire [0:0] s_CSAwallace_cska24_and_20_4;
  wire [0:0] s_CSAwallace_cska24_and_21_4;
  wire [0:0] s_CSAwallace_cska24_and_22_4;
  wire [0:0] s_CSAwallace_cska24_nand_23_4;
  wire [0:0] s_CSAwallace_cska24_and_0_5;
  wire [0:0] s_CSAwallace_cska24_and_1_5;
  wire [0:0] s_CSAwallace_cska24_and_2_5;
  wire [0:0] s_CSAwallace_cska24_and_3_5;
  wire [0:0] s_CSAwallace_cska24_and_4_5;
  wire [0:0] s_CSAwallace_cska24_and_5_5;
  wire [0:0] s_CSAwallace_cska24_and_6_5;
  wire [0:0] s_CSAwallace_cska24_and_7_5;
  wire [0:0] s_CSAwallace_cska24_and_8_5;
  wire [0:0] s_CSAwallace_cska24_and_9_5;
  wire [0:0] s_CSAwallace_cska24_and_10_5;
  wire [0:0] s_CSAwallace_cska24_and_11_5;
  wire [0:0] s_CSAwallace_cska24_and_12_5;
  wire [0:0] s_CSAwallace_cska24_and_13_5;
  wire [0:0] s_CSAwallace_cska24_and_14_5;
  wire [0:0] s_CSAwallace_cska24_and_15_5;
  wire [0:0] s_CSAwallace_cska24_and_16_5;
  wire [0:0] s_CSAwallace_cska24_and_17_5;
  wire [0:0] s_CSAwallace_cska24_and_18_5;
  wire [0:0] s_CSAwallace_cska24_and_19_5;
  wire [0:0] s_CSAwallace_cska24_and_20_5;
  wire [0:0] s_CSAwallace_cska24_and_21_5;
  wire [0:0] s_CSAwallace_cska24_and_22_5;
  wire [0:0] s_CSAwallace_cska24_nand_23_5;
  wire [0:0] s_CSAwallace_cska24_and_0_6;
  wire [0:0] s_CSAwallace_cska24_and_1_6;
  wire [0:0] s_CSAwallace_cska24_and_2_6;
  wire [0:0] s_CSAwallace_cska24_and_3_6;
  wire [0:0] s_CSAwallace_cska24_and_4_6;
  wire [0:0] s_CSAwallace_cska24_and_5_6;
  wire [0:0] s_CSAwallace_cska24_and_6_6;
  wire [0:0] s_CSAwallace_cska24_and_7_6;
  wire [0:0] s_CSAwallace_cska24_and_8_6;
  wire [0:0] s_CSAwallace_cska24_and_9_6;
  wire [0:0] s_CSAwallace_cska24_and_10_6;
  wire [0:0] s_CSAwallace_cska24_and_11_6;
  wire [0:0] s_CSAwallace_cska24_and_12_6;
  wire [0:0] s_CSAwallace_cska24_and_13_6;
  wire [0:0] s_CSAwallace_cska24_and_14_6;
  wire [0:0] s_CSAwallace_cska24_and_15_6;
  wire [0:0] s_CSAwallace_cska24_and_16_6;
  wire [0:0] s_CSAwallace_cska24_and_17_6;
  wire [0:0] s_CSAwallace_cska24_and_18_6;
  wire [0:0] s_CSAwallace_cska24_and_19_6;
  wire [0:0] s_CSAwallace_cska24_and_20_6;
  wire [0:0] s_CSAwallace_cska24_and_21_6;
  wire [0:0] s_CSAwallace_cska24_and_22_6;
  wire [0:0] s_CSAwallace_cska24_nand_23_6;
  wire [0:0] s_CSAwallace_cska24_and_0_7;
  wire [0:0] s_CSAwallace_cska24_and_1_7;
  wire [0:0] s_CSAwallace_cska24_and_2_7;
  wire [0:0] s_CSAwallace_cska24_and_3_7;
  wire [0:0] s_CSAwallace_cska24_and_4_7;
  wire [0:0] s_CSAwallace_cska24_and_5_7;
  wire [0:0] s_CSAwallace_cska24_and_6_7;
  wire [0:0] s_CSAwallace_cska24_and_7_7;
  wire [0:0] s_CSAwallace_cska24_and_8_7;
  wire [0:0] s_CSAwallace_cska24_and_9_7;
  wire [0:0] s_CSAwallace_cska24_and_10_7;
  wire [0:0] s_CSAwallace_cska24_and_11_7;
  wire [0:0] s_CSAwallace_cska24_and_12_7;
  wire [0:0] s_CSAwallace_cska24_and_13_7;
  wire [0:0] s_CSAwallace_cska24_and_14_7;
  wire [0:0] s_CSAwallace_cska24_and_15_7;
  wire [0:0] s_CSAwallace_cska24_and_16_7;
  wire [0:0] s_CSAwallace_cska24_and_17_7;
  wire [0:0] s_CSAwallace_cska24_and_18_7;
  wire [0:0] s_CSAwallace_cska24_and_19_7;
  wire [0:0] s_CSAwallace_cska24_and_20_7;
  wire [0:0] s_CSAwallace_cska24_and_21_7;
  wire [0:0] s_CSAwallace_cska24_and_22_7;
  wire [0:0] s_CSAwallace_cska24_nand_23_7;
  wire [0:0] s_CSAwallace_cska24_and_0_8;
  wire [0:0] s_CSAwallace_cska24_and_1_8;
  wire [0:0] s_CSAwallace_cska24_and_2_8;
  wire [0:0] s_CSAwallace_cska24_and_3_8;
  wire [0:0] s_CSAwallace_cska24_and_4_8;
  wire [0:0] s_CSAwallace_cska24_and_5_8;
  wire [0:0] s_CSAwallace_cska24_and_6_8;
  wire [0:0] s_CSAwallace_cska24_and_7_8;
  wire [0:0] s_CSAwallace_cska24_and_8_8;
  wire [0:0] s_CSAwallace_cska24_and_9_8;
  wire [0:0] s_CSAwallace_cska24_and_10_8;
  wire [0:0] s_CSAwallace_cska24_and_11_8;
  wire [0:0] s_CSAwallace_cska24_and_12_8;
  wire [0:0] s_CSAwallace_cska24_and_13_8;
  wire [0:0] s_CSAwallace_cska24_and_14_8;
  wire [0:0] s_CSAwallace_cska24_and_15_8;
  wire [0:0] s_CSAwallace_cska24_and_16_8;
  wire [0:0] s_CSAwallace_cska24_and_17_8;
  wire [0:0] s_CSAwallace_cska24_and_18_8;
  wire [0:0] s_CSAwallace_cska24_and_19_8;
  wire [0:0] s_CSAwallace_cska24_and_20_8;
  wire [0:0] s_CSAwallace_cska24_and_21_8;
  wire [0:0] s_CSAwallace_cska24_and_22_8;
  wire [0:0] s_CSAwallace_cska24_nand_23_8;
  wire [0:0] s_CSAwallace_cska24_and_0_9;
  wire [0:0] s_CSAwallace_cska24_and_1_9;
  wire [0:0] s_CSAwallace_cska24_and_2_9;
  wire [0:0] s_CSAwallace_cska24_and_3_9;
  wire [0:0] s_CSAwallace_cska24_and_4_9;
  wire [0:0] s_CSAwallace_cska24_and_5_9;
  wire [0:0] s_CSAwallace_cska24_and_6_9;
  wire [0:0] s_CSAwallace_cska24_and_7_9;
  wire [0:0] s_CSAwallace_cska24_and_8_9;
  wire [0:0] s_CSAwallace_cska24_and_9_9;
  wire [0:0] s_CSAwallace_cska24_and_10_9;
  wire [0:0] s_CSAwallace_cska24_and_11_9;
  wire [0:0] s_CSAwallace_cska24_and_12_9;
  wire [0:0] s_CSAwallace_cska24_and_13_9;
  wire [0:0] s_CSAwallace_cska24_and_14_9;
  wire [0:0] s_CSAwallace_cska24_and_15_9;
  wire [0:0] s_CSAwallace_cska24_and_16_9;
  wire [0:0] s_CSAwallace_cska24_and_17_9;
  wire [0:0] s_CSAwallace_cska24_and_18_9;
  wire [0:0] s_CSAwallace_cska24_and_19_9;
  wire [0:0] s_CSAwallace_cska24_and_20_9;
  wire [0:0] s_CSAwallace_cska24_and_21_9;
  wire [0:0] s_CSAwallace_cska24_and_22_9;
  wire [0:0] s_CSAwallace_cska24_nand_23_9;
  wire [0:0] s_CSAwallace_cska24_and_0_10;
  wire [0:0] s_CSAwallace_cska24_and_1_10;
  wire [0:0] s_CSAwallace_cska24_and_2_10;
  wire [0:0] s_CSAwallace_cska24_and_3_10;
  wire [0:0] s_CSAwallace_cska24_and_4_10;
  wire [0:0] s_CSAwallace_cska24_and_5_10;
  wire [0:0] s_CSAwallace_cska24_and_6_10;
  wire [0:0] s_CSAwallace_cska24_and_7_10;
  wire [0:0] s_CSAwallace_cska24_and_8_10;
  wire [0:0] s_CSAwallace_cska24_and_9_10;
  wire [0:0] s_CSAwallace_cska24_and_10_10;
  wire [0:0] s_CSAwallace_cska24_and_11_10;
  wire [0:0] s_CSAwallace_cska24_and_12_10;
  wire [0:0] s_CSAwallace_cska24_and_13_10;
  wire [0:0] s_CSAwallace_cska24_and_14_10;
  wire [0:0] s_CSAwallace_cska24_and_15_10;
  wire [0:0] s_CSAwallace_cska24_and_16_10;
  wire [0:0] s_CSAwallace_cska24_and_17_10;
  wire [0:0] s_CSAwallace_cska24_and_18_10;
  wire [0:0] s_CSAwallace_cska24_and_19_10;
  wire [0:0] s_CSAwallace_cska24_and_20_10;
  wire [0:0] s_CSAwallace_cska24_and_21_10;
  wire [0:0] s_CSAwallace_cska24_and_22_10;
  wire [0:0] s_CSAwallace_cska24_nand_23_10;
  wire [0:0] s_CSAwallace_cska24_and_0_11;
  wire [0:0] s_CSAwallace_cska24_and_1_11;
  wire [0:0] s_CSAwallace_cska24_and_2_11;
  wire [0:0] s_CSAwallace_cska24_and_3_11;
  wire [0:0] s_CSAwallace_cska24_and_4_11;
  wire [0:0] s_CSAwallace_cska24_and_5_11;
  wire [0:0] s_CSAwallace_cska24_and_6_11;
  wire [0:0] s_CSAwallace_cska24_and_7_11;
  wire [0:0] s_CSAwallace_cska24_and_8_11;
  wire [0:0] s_CSAwallace_cska24_and_9_11;
  wire [0:0] s_CSAwallace_cska24_and_10_11;
  wire [0:0] s_CSAwallace_cska24_and_11_11;
  wire [0:0] s_CSAwallace_cska24_and_12_11;
  wire [0:0] s_CSAwallace_cska24_and_13_11;
  wire [0:0] s_CSAwallace_cska24_and_14_11;
  wire [0:0] s_CSAwallace_cska24_and_15_11;
  wire [0:0] s_CSAwallace_cska24_and_16_11;
  wire [0:0] s_CSAwallace_cska24_and_17_11;
  wire [0:0] s_CSAwallace_cska24_and_18_11;
  wire [0:0] s_CSAwallace_cska24_and_19_11;
  wire [0:0] s_CSAwallace_cska24_and_20_11;
  wire [0:0] s_CSAwallace_cska24_and_21_11;
  wire [0:0] s_CSAwallace_cska24_and_22_11;
  wire [0:0] s_CSAwallace_cska24_nand_23_11;
  wire [0:0] s_CSAwallace_cska24_and_0_12;
  wire [0:0] s_CSAwallace_cska24_and_1_12;
  wire [0:0] s_CSAwallace_cska24_and_2_12;
  wire [0:0] s_CSAwallace_cska24_and_3_12;
  wire [0:0] s_CSAwallace_cska24_and_4_12;
  wire [0:0] s_CSAwallace_cska24_and_5_12;
  wire [0:0] s_CSAwallace_cska24_and_6_12;
  wire [0:0] s_CSAwallace_cska24_and_7_12;
  wire [0:0] s_CSAwallace_cska24_and_8_12;
  wire [0:0] s_CSAwallace_cska24_and_9_12;
  wire [0:0] s_CSAwallace_cska24_and_10_12;
  wire [0:0] s_CSAwallace_cska24_and_11_12;
  wire [0:0] s_CSAwallace_cska24_and_12_12;
  wire [0:0] s_CSAwallace_cska24_and_13_12;
  wire [0:0] s_CSAwallace_cska24_and_14_12;
  wire [0:0] s_CSAwallace_cska24_and_15_12;
  wire [0:0] s_CSAwallace_cska24_and_16_12;
  wire [0:0] s_CSAwallace_cska24_and_17_12;
  wire [0:0] s_CSAwallace_cska24_and_18_12;
  wire [0:0] s_CSAwallace_cska24_and_19_12;
  wire [0:0] s_CSAwallace_cska24_and_20_12;
  wire [0:0] s_CSAwallace_cska24_and_21_12;
  wire [0:0] s_CSAwallace_cska24_and_22_12;
  wire [0:0] s_CSAwallace_cska24_nand_23_12;
  wire [0:0] s_CSAwallace_cska24_and_0_13;
  wire [0:0] s_CSAwallace_cska24_and_1_13;
  wire [0:0] s_CSAwallace_cska24_and_2_13;
  wire [0:0] s_CSAwallace_cska24_and_3_13;
  wire [0:0] s_CSAwallace_cska24_and_4_13;
  wire [0:0] s_CSAwallace_cska24_and_5_13;
  wire [0:0] s_CSAwallace_cska24_and_6_13;
  wire [0:0] s_CSAwallace_cska24_and_7_13;
  wire [0:0] s_CSAwallace_cska24_and_8_13;
  wire [0:0] s_CSAwallace_cska24_and_9_13;
  wire [0:0] s_CSAwallace_cska24_and_10_13;
  wire [0:0] s_CSAwallace_cska24_and_11_13;
  wire [0:0] s_CSAwallace_cska24_and_12_13;
  wire [0:0] s_CSAwallace_cska24_and_13_13;
  wire [0:0] s_CSAwallace_cska24_and_14_13;
  wire [0:0] s_CSAwallace_cska24_and_15_13;
  wire [0:0] s_CSAwallace_cska24_and_16_13;
  wire [0:0] s_CSAwallace_cska24_and_17_13;
  wire [0:0] s_CSAwallace_cska24_and_18_13;
  wire [0:0] s_CSAwallace_cska24_and_19_13;
  wire [0:0] s_CSAwallace_cska24_and_20_13;
  wire [0:0] s_CSAwallace_cska24_and_21_13;
  wire [0:0] s_CSAwallace_cska24_and_22_13;
  wire [0:0] s_CSAwallace_cska24_nand_23_13;
  wire [0:0] s_CSAwallace_cska24_and_0_14;
  wire [0:0] s_CSAwallace_cska24_and_1_14;
  wire [0:0] s_CSAwallace_cska24_and_2_14;
  wire [0:0] s_CSAwallace_cska24_and_3_14;
  wire [0:0] s_CSAwallace_cska24_and_4_14;
  wire [0:0] s_CSAwallace_cska24_and_5_14;
  wire [0:0] s_CSAwallace_cska24_and_6_14;
  wire [0:0] s_CSAwallace_cska24_and_7_14;
  wire [0:0] s_CSAwallace_cska24_and_8_14;
  wire [0:0] s_CSAwallace_cska24_and_9_14;
  wire [0:0] s_CSAwallace_cska24_and_10_14;
  wire [0:0] s_CSAwallace_cska24_and_11_14;
  wire [0:0] s_CSAwallace_cska24_and_12_14;
  wire [0:0] s_CSAwallace_cska24_and_13_14;
  wire [0:0] s_CSAwallace_cska24_and_14_14;
  wire [0:0] s_CSAwallace_cska24_and_15_14;
  wire [0:0] s_CSAwallace_cska24_and_16_14;
  wire [0:0] s_CSAwallace_cska24_and_17_14;
  wire [0:0] s_CSAwallace_cska24_and_18_14;
  wire [0:0] s_CSAwallace_cska24_and_19_14;
  wire [0:0] s_CSAwallace_cska24_and_20_14;
  wire [0:0] s_CSAwallace_cska24_and_21_14;
  wire [0:0] s_CSAwallace_cska24_and_22_14;
  wire [0:0] s_CSAwallace_cska24_nand_23_14;
  wire [0:0] s_CSAwallace_cska24_and_0_15;
  wire [0:0] s_CSAwallace_cska24_and_1_15;
  wire [0:0] s_CSAwallace_cska24_and_2_15;
  wire [0:0] s_CSAwallace_cska24_and_3_15;
  wire [0:0] s_CSAwallace_cska24_and_4_15;
  wire [0:0] s_CSAwallace_cska24_and_5_15;
  wire [0:0] s_CSAwallace_cska24_and_6_15;
  wire [0:0] s_CSAwallace_cska24_and_7_15;
  wire [0:0] s_CSAwallace_cska24_and_8_15;
  wire [0:0] s_CSAwallace_cska24_and_9_15;
  wire [0:0] s_CSAwallace_cska24_and_10_15;
  wire [0:0] s_CSAwallace_cska24_and_11_15;
  wire [0:0] s_CSAwallace_cska24_and_12_15;
  wire [0:0] s_CSAwallace_cska24_and_13_15;
  wire [0:0] s_CSAwallace_cska24_and_14_15;
  wire [0:0] s_CSAwallace_cska24_and_15_15;
  wire [0:0] s_CSAwallace_cska24_and_16_15;
  wire [0:0] s_CSAwallace_cska24_and_17_15;
  wire [0:0] s_CSAwallace_cska24_and_18_15;
  wire [0:0] s_CSAwallace_cska24_and_19_15;
  wire [0:0] s_CSAwallace_cska24_and_20_15;
  wire [0:0] s_CSAwallace_cska24_and_21_15;
  wire [0:0] s_CSAwallace_cska24_and_22_15;
  wire [0:0] s_CSAwallace_cska24_nand_23_15;
  wire [0:0] s_CSAwallace_cska24_and_0_16;
  wire [0:0] s_CSAwallace_cska24_and_1_16;
  wire [0:0] s_CSAwallace_cska24_and_2_16;
  wire [0:0] s_CSAwallace_cska24_and_3_16;
  wire [0:0] s_CSAwallace_cska24_and_4_16;
  wire [0:0] s_CSAwallace_cska24_and_5_16;
  wire [0:0] s_CSAwallace_cska24_and_6_16;
  wire [0:0] s_CSAwallace_cska24_and_7_16;
  wire [0:0] s_CSAwallace_cska24_and_8_16;
  wire [0:0] s_CSAwallace_cska24_and_9_16;
  wire [0:0] s_CSAwallace_cska24_and_10_16;
  wire [0:0] s_CSAwallace_cska24_and_11_16;
  wire [0:0] s_CSAwallace_cska24_and_12_16;
  wire [0:0] s_CSAwallace_cska24_and_13_16;
  wire [0:0] s_CSAwallace_cska24_and_14_16;
  wire [0:0] s_CSAwallace_cska24_and_15_16;
  wire [0:0] s_CSAwallace_cska24_and_16_16;
  wire [0:0] s_CSAwallace_cska24_and_17_16;
  wire [0:0] s_CSAwallace_cska24_and_18_16;
  wire [0:0] s_CSAwallace_cska24_and_19_16;
  wire [0:0] s_CSAwallace_cska24_and_20_16;
  wire [0:0] s_CSAwallace_cska24_and_21_16;
  wire [0:0] s_CSAwallace_cska24_and_22_16;
  wire [0:0] s_CSAwallace_cska24_nand_23_16;
  wire [0:0] s_CSAwallace_cska24_and_0_17;
  wire [0:0] s_CSAwallace_cska24_and_1_17;
  wire [0:0] s_CSAwallace_cska24_and_2_17;
  wire [0:0] s_CSAwallace_cska24_and_3_17;
  wire [0:0] s_CSAwallace_cska24_and_4_17;
  wire [0:0] s_CSAwallace_cska24_and_5_17;
  wire [0:0] s_CSAwallace_cska24_and_6_17;
  wire [0:0] s_CSAwallace_cska24_and_7_17;
  wire [0:0] s_CSAwallace_cska24_and_8_17;
  wire [0:0] s_CSAwallace_cska24_and_9_17;
  wire [0:0] s_CSAwallace_cska24_and_10_17;
  wire [0:0] s_CSAwallace_cska24_and_11_17;
  wire [0:0] s_CSAwallace_cska24_and_12_17;
  wire [0:0] s_CSAwallace_cska24_and_13_17;
  wire [0:0] s_CSAwallace_cska24_and_14_17;
  wire [0:0] s_CSAwallace_cska24_and_15_17;
  wire [0:0] s_CSAwallace_cska24_and_16_17;
  wire [0:0] s_CSAwallace_cska24_and_17_17;
  wire [0:0] s_CSAwallace_cska24_and_18_17;
  wire [0:0] s_CSAwallace_cska24_and_19_17;
  wire [0:0] s_CSAwallace_cska24_and_20_17;
  wire [0:0] s_CSAwallace_cska24_and_21_17;
  wire [0:0] s_CSAwallace_cska24_and_22_17;
  wire [0:0] s_CSAwallace_cska24_nand_23_17;
  wire [0:0] s_CSAwallace_cska24_and_0_18;
  wire [0:0] s_CSAwallace_cska24_and_1_18;
  wire [0:0] s_CSAwallace_cska24_and_2_18;
  wire [0:0] s_CSAwallace_cska24_and_3_18;
  wire [0:0] s_CSAwallace_cska24_and_4_18;
  wire [0:0] s_CSAwallace_cska24_and_5_18;
  wire [0:0] s_CSAwallace_cska24_and_6_18;
  wire [0:0] s_CSAwallace_cska24_and_7_18;
  wire [0:0] s_CSAwallace_cska24_and_8_18;
  wire [0:0] s_CSAwallace_cska24_and_9_18;
  wire [0:0] s_CSAwallace_cska24_and_10_18;
  wire [0:0] s_CSAwallace_cska24_and_11_18;
  wire [0:0] s_CSAwallace_cska24_and_12_18;
  wire [0:0] s_CSAwallace_cska24_and_13_18;
  wire [0:0] s_CSAwallace_cska24_and_14_18;
  wire [0:0] s_CSAwallace_cska24_and_15_18;
  wire [0:0] s_CSAwallace_cska24_and_16_18;
  wire [0:0] s_CSAwallace_cska24_and_17_18;
  wire [0:0] s_CSAwallace_cska24_and_18_18;
  wire [0:0] s_CSAwallace_cska24_and_19_18;
  wire [0:0] s_CSAwallace_cska24_and_20_18;
  wire [0:0] s_CSAwallace_cska24_and_21_18;
  wire [0:0] s_CSAwallace_cska24_and_22_18;
  wire [0:0] s_CSAwallace_cska24_nand_23_18;
  wire [0:0] s_CSAwallace_cska24_and_0_19;
  wire [0:0] s_CSAwallace_cska24_and_1_19;
  wire [0:0] s_CSAwallace_cska24_and_2_19;
  wire [0:0] s_CSAwallace_cska24_and_3_19;
  wire [0:0] s_CSAwallace_cska24_and_4_19;
  wire [0:0] s_CSAwallace_cska24_and_5_19;
  wire [0:0] s_CSAwallace_cska24_and_6_19;
  wire [0:0] s_CSAwallace_cska24_and_7_19;
  wire [0:0] s_CSAwallace_cska24_and_8_19;
  wire [0:0] s_CSAwallace_cska24_and_9_19;
  wire [0:0] s_CSAwallace_cska24_and_10_19;
  wire [0:0] s_CSAwallace_cska24_and_11_19;
  wire [0:0] s_CSAwallace_cska24_and_12_19;
  wire [0:0] s_CSAwallace_cska24_and_13_19;
  wire [0:0] s_CSAwallace_cska24_and_14_19;
  wire [0:0] s_CSAwallace_cska24_and_15_19;
  wire [0:0] s_CSAwallace_cska24_and_16_19;
  wire [0:0] s_CSAwallace_cska24_and_17_19;
  wire [0:0] s_CSAwallace_cska24_and_18_19;
  wire [0:0] s_CSAwallace_cska24_and_19_19;
  wire [0:0] s_CSAwallace_cska24_and_20_19;
  wire [0:0] s_CSAwallace_cska24_and_21_19;
  wire [0:0] s_CSAwallace_cska24_and_22_19;
  wire [0:0] s_CSAwallace_cska24_nand_23_19;
  wire [0:0] s_CSAwallace_cska24_and_0_20;
  wire [0:0] s_CSAwallace_cska24_and_1_20;
  wire [0:0] s_CSAwallace_cska24_and_2_20;
  wire [0:0] s_CSAwallace_cska24_and_3_20;
  wire [0:0] s_CSAwallace_cska24_and_4_20;
  wire [0:0] s_CSAwallace_cska24_and_5_20;
  wire [0:0] s_CSAwallace_cska24_and_6_20;
  wire [0:0] s_CSAwallace_cska24_and_7_20;
  wire [0:0] s_CSAwallace_cska24_and_8_20;
  wire [0:0] s_CSAwallace_cska24_and_9_20;
  wire [0:0] s_CSAwallace_cska24_and_10_20;
  wire [0:0] s_CSAwallace_cska24_and_11_20;
  wire [0:0] s_CSAwallace_cska24_and_12_20;
  wire [0:0] s_CSAwallace_cska24_and_13_20;
  wire [0:0] s_CSAwallace_cska24_and_14_20;
  wire [0:0] s_CSAwallace_cska24_and_15_20;
  wire [0:0] s_CSAwallace_cska24_and_16_20;
  wire [0:0] s_CSAwallace_cska24_and_17_20;
  wire [0:0] s_CSAwallace_cska24_and_18_20;
  wire [0:0] s_CSAwallace_cska24_and_19_20;
  wire [0:0] s_CSAwallace_cska24_and_20_20;
  wire [0:0] s_CSAwallace_cska24_and_21_20;
  wire [0:0] s_CSAwallace_cska24_and_22_20;
  wire [0:0] s_CSAwallace_cska24_nand_23_20;
  wire [0:0] s_CSAwallace_cska24_and_0_21;
  wire [0:0] s_CSAwallace_cska24_and_1_21;
  wire [0:0] s_CSAwallace_cska24_and_2_21;
  wire [0:0] s_CSAwallace_cska24_and_3_21;
  wire [0:0] s_CSAwallace_cska24_and_4_21;
  wire [0:0] s_CSAwallace_cska24_and_5_21;
  wire [0:0] s_CSAwallace_cska24_and_6_21;
  wire [0:0] s_CSAwallace_cska24_and_7_21;
  wire [0:0] s_CSAwallace_cska24_and_8_21;
  wire [0:0] s_CSAwallace_cska24_and_9_21;
  wire [0:0] s_CSAwallace_cska24_and_10_21;
  wire [0:0] s_CSAwallace_cska24_and_11_21;
  wire [0:0] s_CSAwallace_cska24_and_12_21;
  wire [0:0] s_CSAwallace_cska24_and_13_21;
  wire [0:0] s_CSAwallace_cska24_and_14_21;
  wire [0:0] s_CSAwallace_cska24_and_15_21;
  wire [0:0] s_CSAwallace_cska24_and_16_21;
  wire [0:0] s_CSAwallace_cska24_and_17_21;
  wire [0:0] s_CSAwallace_cska24_and_18_21;
  wire [0:0] s_CSAwallace_cska24_and_19_21;
  wire [0:0] s_CSAwallace_cska24_and_20_21;
  wire [0:0] s_CSAwallace_cska24_and_21_21;
  wire [0:0] s_CSAwallace_cska24_and_22_21;
  wire [0:0] s_CSAwallace_cska24_nand_23_21;
  wire [0:0] s_CSAwallace_cska24_and_0_22;
  wire [0:0] s_CSAwallace_cska24_and_1_22;
  wire [0:0] s_CSAwallace_cska24_and_2_22;
  wire [0:0] s_CSAwallace_cska24_and_3_22;
  wire [0:0] s_CSAwallace_cska24_and_4_22;
  wire [0:0] s_CSAwallace_cska24_and_5_22;
  wire [0:0] s_CSAwallace_cska24_and_6_22;
  wire [0:0] s_CSAwallace_cska24_and_7_22;
  wire [0:0] s_CSAwallace_cska24_and_8_22;
  wire [0:0] s_CSAwallace_cska24_and_9_22;
  wire [0:0] s_CSAwallace_cska24_and_10_22;
  wire [0:0] s_CSAwallace_cska24_and_11_22;
  wire [0:0] s_CSAwallace_cska24_and_12_22;
  wire [0:0] s_CSAwallace_cska24_and_13_22;
  wire [0:0] s_CSAwallace_cska24_and_14_22;
  wire [0:0] s_CSAwallace_cska24_and_15_22;
  wire [0:0] s_CSAwallace_cska24_and_16_22;
  wire [0:0] s_CSAwallace_cska24_and_17_22;
  wire [0:0] s_CSAwallace_cska24_and_18_22;
  wire [0:0] s_CSAwallace_cska24_and_19_22;
  wire [0:0] s_CSAwallace_cska24_and_20_22;
  wire [0:0] s_CSAwallace_cska24_and_21_22;
  wire [0:0] s_CSAwallace_cska24_and_22_22;
  wire [0:0] s_CSAwallace_cska24_nand_23_22;
  wire [0:0] s_CSAwallace_cska24_nand_0_23;
  wire [0:0] s_CSAwallace_cska24_nand_1_23;
  wire [0:0] s_CSAwallace_cska24_nand_2_23;
  wire [0:0] s_CSAwallace_cska24_nand_3_23;
  wire [0:0] s_CSAwallace_cska24_nand_4_23;
  wire [0:0] s_CSAwallace_cska24_nand_5_23;
  wire [0:0] s_CSAwallace_cska24_nand_6_23;
  wire [0:0] s_CSAwallace_cska24_nand_7_23;
  wire [0:0] s_CSAwallace_cska24_nand_8_23;
  wire [0:0] s_CSAwallace_cska24_nand_9_23;
  wire [0:0] s_CSAwallace_cska24_nand_10_23;
  wire [0:0] s_CSAwallace_cska24_nand_11_23;
  wire [0:0] s_CSAwallace_cska24_nand_12_23;
  wire [0:0] s_CSAwallace_cska24_nand_13_23;
  wire [0:0] s_CSAwallace_cska24_nand_14_23;
  wire [0:0] s_CSAwallace_cska24_nand_15_23;
  wire [0:0] s_CSAwallace_cska24_nand_16_23;
  wire [0:0] s_CSAwallace_cska24_nand_17_23;
  wire [0:0] s_CSAwallace_cska24_nand_18_23;
  wire [0:0] s_CSAwallace_cska24_nand_19_23;
  wire [0:0] s_CSAwallace_cska24_nand_20_23;
  wire [0:0] s_CSAwallace_cska24_nand_21_23;
  wire [0:0] s_CSAwallace_cska24_nand_22_23;
  wire [0:0] s_CSAwallace_cska24_and_23_23;
  wire [25:0] s_CSAwallace_cska24_csa0_csa_component_pp_row0;
  wire [25:0] s_CSAwallace_cska24_csa0_csa_component_pp_row1;
  wire [25:0] s_CSAwallace_cska24_csa0_csa_component_pp_row2;
  wire [53:0] s_CSAwallace_cska24_csa0_csa_component_out;
  wire [28:0] s_CSAwallace_cska24_csa1_csa_component_pp_row3;
  wire [28:0] s_CSAwallace_cska24_csa1_csa_component_pp_row4;
  wire [28:0] s_CSAwallace_cska24_csa1_csa_component_pp_row5;
  wire [59:0] s_CSAwallace_cska24_csa1_csa_component_out;
  wire [31:0] s_CSAwallace_cska24_csa2_csa_component_pp_row6;
  wire [31:0] s_CSAwallace_cska24_csa2_csa_component_pp_row7;
  wire [31:0] s_CSAwallace_cska24_csa2_csa_component_pp_row8;
  wire [65:0] s_CSAwallace_cska24_csa2_csa_component_out;
  wire [34:0] s_CSAwallace_cska24_csa3_csa_component_pp_row9;
  wire [34:0] s_CSAwallace_cska24_csa3_csa_component_pp_row10;
  wire [34:0] s_CSAwallace_cska24_csa3_csa_component_pp_row11;
  wire [71:0] s_CSAwallace_cska24_csa3_csa_component_out;
  wire [37:0] s_CSAwallace_cska24_csa4_csa_component_pp_row12;
  wire [37:0] s_CSAwallace_cska24_csa4_csa_component_pp_row13;
  wire [37:0] s_CSAwallace_cska24_csa4_csa_component_pp_row14;
  wire [77:0] s_CSAwallace_cska24_csa4_csa_component_out;
  wire [40:0] s_CSAwallace_cska24_csa5_csa_component_pp_row15;
  wire [40:0] s_CSAwallace_cska24_csa5_csa_component_pp_row16;
  wire [40:0] s_CSAwallace_cska24_csa5_csa_component_pp_row17;
  wire [83:0] s_CSAwallace_cska24_csa5_csa_component_out;
  wire [43:0] s_CSAwallace_cska24_csa6_csa_component_pp_row18;
  wire [43:0] s_CSAwallace_cska24_csa6_csa_component_pp_row19;
  wire [43:0] s_CSAwallace_cska24_csa6_csa_component_pp_row20;
  wire [89:0] s_CSAwallace_cska24_csa6_csa_component_out;
  wire [46:0] s_CSAwallace_cska24_csa7_csa_component_pp_row21;
  wire [46:0] s_CSAwallace_cska24_csa7_csa_component_pp_row22;
  wire [46:0] s_CSAwallace_cska24_csa7_csa_component_pp_row23;
  wire [95:0] s_CSAwallace_cska24_csa7_csa_component_out;
  wire [29:0] s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1;
  wire [29:0] s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1;
  wire [29:0] s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2;
  wire [61:0] s_CSAwallace_cska24_csa8_csa_component_out;
  wire [32:0] s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2;
  wire [32:0] s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3;
  wire [32:0] s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3;
  wire [67:0] s_CSAwallace_cska24_csa9_csa_component_out;
  wire [38:0] s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4;
  wire [38:0] s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4;
  wire [38:0] s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5;
  wire [79:0] s_CSAwallace_cska24_csa10_csa_component_out;
  wire [41:0] s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5;
  wire [41:0] s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6;
  wire [41:0] s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6;
  wire [85:0] s_CSAwallace_cska24_csa11_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7;
  wire [47:0] s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7;
  wire [47:0] s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8;
  wire [97:0] s_CSAwallace_cska24_csa12_csa_component_out;
  wire [33:0] s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9;
  wire [33:0] s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9;
  wire [33:0] s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10;
  wire [69:0] s_CSAwallace_cska24_csa13_csa_component_out;
  wire [39:0] s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10;
  wire [39:0] s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11;
  wire [39:0] s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11;
  wire [81:0] s_CSAwallace_cska24_csa14_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12;
  wire [47:0] s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12;
  wire [47:0] s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13;
  wire [97:0] s_CSAwallace_cska24_csa15_csa_component_out;
  wire [40:0] s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14;
  wire [40:0] s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14;
  wire [40:0] s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15;
  wire [83:0] s_CSAwallace_cska24_csa16_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15;
  wire [47:0] s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16;
  wire [47:0] s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16;
  wire [97:0] s_CSAwallace_cska24_csa17_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17;
  wire [47:0] s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17;
  wire [47:0] s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18;
  wire [97:0] s_CSAwallace_cska24_csa18_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18;
  wire [47:0] s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13;
  wire [47:0] s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8;
  wire [97:0] s_CSAwallace_cska24_csa19_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19;
  wire [47:0] s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19;
  wire [47:0] s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20;
  wire [97:0] s_CSAwallace_cska24_csa20_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21;
  wire [47:0] s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21;
  wire [47:0] s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20;
  wire [97:0] s_CSAwallace_cska24_csa21_csa_component_out;
  wire [47:0] s_CSAwallace_cska24_u_cska48_a;
  wire [47:0] s_CSAwallace_cska24_u_cska48_b;
  wire [48:0] s_CSAwallace_cska24_u_cska48_out;
  wire [0:0] s_CSAwallace_cska24_xor0;

  and_gate and_gate_s_CSAwallace_cska24_and_0_0(.a(a[0]), .b(b[0]), .out(s_CSAwallace_cska24_and_0_0));
  and_gate and_gate_s_CSAwallace_cska24_and_1_0(.a(a[1]), .b(b[0]), .out(s_CSAwallace_cska24_and_1_0));
  and_gate and_gate_s_CSAwallace_cska24_and_2_0(.a(a[2]), .b(b[0]), .out(s_CSAwallace_cska24_and_2_0));
  and_gate and_gate_s_CSAwallace_cska24_and_3_0(.a(a[3]), .b(b[0]), .out(s_CSAwallace_cska24_and_3_0));
  and_gate and_gate_s_CSAwallace_cska24_and_4_0(.a(a[4]), .b(b[0]), .out(s_CSAwallace_cska24_and_4_0));
  and_gate and_gate_s_CSAwallace_cska24_and_5_0(.a(a[5]), .b(b[0]), .out(s_CSAwallace_cska24_and_5_0));
  and_gate and_gate_s_CSAwallace_cska24_and_6_0(.a(a[6]), .b(b[0]), .out(s_CSAwallace_cska24_and_6_0));
  and_gate and_gate_s_CSAwallace_cska24_and_7_0(.a(a[7]), .b(b[0]), .out(s_CSAwallace_cska24_and_7_0));
  and_gate and_gate_s_CSAwallace_cska24_and_8_0(.a(a[8]), .b(b[0]), .out(s_CSAwallace_cska24_and_8_0));
  and_gate and_gate_s_CSAwallace_cska24_and_9_0(.a(a[9]), .b(b[0]), .out(s_CSAwallace_cska24_and_9_0));
  and_gate and_gate_s_CSAwallace_cska24_and_10_0(.a(a[10]), .b(b[0]), .out(s_CSAwallace_cska24_and_10_0));
  and_gate and_gate_s_CSAwallace_cska24_and_11_0(.a(a[11]), .b(b[0]), .out(s_CSAwallace_cska24_and_11_0));
  and_gate and_gate_s_CSAwallace_cska24_and_12_0(.a(a[12]), .b(b[0]), .out(s_CSAwallace_cska24_and_12_0));
  and_gate and_gate_s_CSAwallace_cska24_and_13_0(.a(a[13]), .b(b[0]), .out(s_CSAwallace_cska24_and_13_0));
  and_gate and_gate_s_CSAwallace_cska24_and_14_0(.a(a[14]), .b(b[0]), .out(s_CSAwallace_cska24_and_14_0));
  and_gate and_gate_s_CSAwallace_cska24_and_15_0(.a(a[15]), .b(b[0]), .out(s_CSAwallace_cska24_and_15_0));
  and_gate and_gate_s_CSAwallace_cska24_and_16_0(.a(a[16]), .b(b[0]), .out(s_CSAwallace_cska24_and_16_0));
  and_gate and_gate_s_CSAwallace_cska24_and_17_0(.a(a[17]), .b(b[0]), .out(s_CSAwallace_cska24_and_17_0));
  and_gate and_gate_s_CSAwallace_cska24_and_18_0(.a(a[18]), .b(b[0]), .out(s_CSAwallace_cska24_and_18_0));
  and_gate and_gate_s_CSAwallace_cska24_and_19_0(.a(a[19]), .b(b[0]), .out(s_CSAwallace_cska24_and_19_0));
  and_gate and_gate_s_CSAwallace_cska24_and_20_0(.a(a[20]), .b(b[0]), .out(s_CSAwallace_cska24_and_20_0));
  and_gate and_gate_s_CSAwallace_cska24_and_21_0(.a(a[21]), .b(b[0]), .out(s_CSAwallace_cska24_and_21_0));
  and_gate and_gate_s_CSAwallace_cska24_and_22_0(.a(a[22]), .b(b[0]), .out(s_CSAwallace_cska24_and_22_0));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_0(.a(a[23]), .b(b[0]), .out(s_CSAwallace_cska24_nand_23_0));
  and_gate and_gate_s_CSAwallace_cska24_and_0_1(.a(a[0]), .b(b[1]), .out(s_CSAwallace_cska24_and_0_1));
  and_gate and_gate_s_CSAwallace_cska24_and_1_1(.a(a[1]), .b(b[1]), .out(s_CSAwallace_cska24_and_1_1));
  and_gate and_gate_s_CSAwallace_cska24_and_2_1(.a(a[2]), .b(b[1]), .out(s_CSAwallace_cska24_and_2_1));
  and_gate and_gate_s_CSAwallace_cska24_and_3_1(.a(a[3]), .b(b[1]), .out(s_CSAwallace_cska24_and_3_1));
  and_gate and_gate_s_CSAwallace_cska24_and_4_1(.a(a[4]), .b(b[1]), .out(s_CSAwallace_cska24_and_4_1));
  and_gate and_gate_s_CSAwallace_cska24_and_5_1(.a(a[5]), .b(b[1]), .out(s_CSAwallace_cska24_and_5_1));
  and_gate and_gate_s_CSAwallace_cska24_and_6_1(.a(a[6]), .b(b[1]), .out(s_CSAwallace_cska24_and_6_1));
  and_gate and_gate_s_CSAwallace_cska24_and_7_1(.a(a[7]), .b(b[1]), .out(s_CSAwallace_cska24_and_7_1));
  and_gate and_gate_s_CSAwallace_cska24_and_8_1(.a(a[8]), .b(b[1]), .out(s_CSAwallace_cska24_and_8_1));
  and_gate and_gate_s_CSAwallace_cska24_and_9_1(.a(a[9]), .b(b[1]), .out(s_CSAwallace_cska24_and_9_1));
  and_gate and_gate_s_CSAwallace_cska24_and_10_1(.a(a[10]), .b(b[1]), .out(s_CSAwallace_cska24_and_10_1));
  and_gate and_gate_s_CSAwallace_cska24_and_11_1(.a(a[11]), .b(b[1]), .out(s_CSAwallace_cska24_and_11_1));
  and_gate and_gate_s_CSAwallace_cska24_and_12_1(.a(a[12]), .b(b[1]), .out(s_CSAwallace_cska24_and_12_1));
  and_gate and_gate_s_CSAwallace_cska24_and_13_1(.a(a[13]), .b(b[1]), .out(s_CSAwallace_cska24_and_13_1));
  and_gate and_gate_s_CSAwallace_cska24_and_14_1(.a(a[14]), .b(b[1]), .out(s_CSAwallace_cska24_and_14_1));
  and_gate and_gate_s_CSAwallace_cska24_and_15_1(.a(a[15]), .b(b[1]), .out(s_CSAwallace_cska24_and_15_1));
  and_gate and_gate_s_CSAwallace_cska24_and_16_1(.a(a[16]), .b(b[1]), .out(s_CSAwallace_cska24_and_16_1));
  and_gate and_gate_s_CSAwallace_cska24_and_17_1(.a(a[17]), .b(b[1]), .out(s_CSAwallace_cska24_and_17_1));
  and_gate and_gate_s_CSAwallace_cska24_and_18_1(.a(a[18]), .b(b[1]), .out(s_CSAwallace_cska24_and_18_1));
  and_gate and_gate_s_CSAwallace_cska24_and_19_1(.a(a[19]), .b(b[1]), .out(s_CSAwallace_cska24_and_19_1));
  and_gate and_gate_s_CSAwallace_cska24_and_20_1(.a(a[20]), .b(b[1]), .out(s_CSAwallace_cska24_and_20_1));
  and_gate and_gate_s_CSAwallace_cska24_and_21_1(.a(a[21]), .b(b[1]), .out(s_CSAwallace_cska24_and_21_1));
  and_gate and_gate_s_CSAwallace_cska24_and_22_1(.a(a[22]), .b(b[1]), .out(s_CSAwallace_cska24_and_22_1));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_1(.a(a[23]), .b(b[1]), .out(s_CSAwallace_cska24_nand_23_1));
  and_gate and_gate_s_CSAwallace_cska24_and_0_2(.a(a[0]), .b(b[2]), .out(s_CSAwallace_cska24_and_0_2));
  and_gate and_gate_s_CSAwallace_cska24_and_1_2(.a(a[1]), .b(b[2]), .out(s_CSAwallace_cska24_and_1_2));
  and_gate and_gate_s_CSAwallace_cska24_and_2_2(.a(a[2]), .b(b[2]), .out(s_CSAwallace_cska24_and_2_2));
  and_gate and_gate_s_CSAwallace_cska24_and_3_2(.a(a[3]), .b(b[2]), .out(s_CSAwallace_cska24_and_3_2));
  and_gate and_gate_s_CSAwallace_cska24_and_4_2(.a(a[4]), .b(b[2]), .out(s_CSAwallace_cska24_and_4_2));
  and_gate and_gate_s_CSAwallace_cska24_and_5_2(.a(a[5]), .b(b[2]), .out(s_CSAwallace_cska24_and_5_2));
  and_gate and_gate_s_CSAwallace_cska24_and_6_2(.a(a[6]), .b(b[2]), .out(s_CSAwallace_cska24_and_6_2));
  and_gate and_gate_s_CSAwallace_cska24_and_7_2(.a(a[7]), .b(b[2]), .out(s_CSAwallace_cska24_and_7_2));
  and_gate and_gate_s_CSAwallace_cska24_and_8_2(.a(a[8]), .b(b[2]), .out(s_CSAwallace_cska24_and_8_2));
  and_gate and_gate_s_CSAwallace_cska24_and_9_2(.a(a[9]), .b(b[2]), .out(s_CSAwallace_cska24_and_9_2));
  and_gate and_gate_s_CSAwallace_cska24_and_10_2(.a(a[10]), .b(b[2]), .out(s_CSAwallace_cska24_and_10_2));
  and_gate and_gate_s_CSAwallace_cska24_and_11_2(.a(a[11]), .b(b[2]), .out(s_CSAwallace_cska24_and_11_2));
  and_gate and_gate_s_CSAwallace_cska24_and_12_2(.a(a[12]), .b(b[2]), .out(s_CSAwallace_cska24_and_12_2));
  and_gate and_gate_s_CSAwallace_cska24_and_13_2(.a(a[13]), .b(b[2]), .out(s_CSAwallace_cska24_and_13_2));
  and_gate and_gate_s_CSAwallace_cska24_and_14_2(.a(a[14]), .b(b[2]), .out(s_CSAwallace_cska24_and_14_2));
  and_gate and_gate_s_CSAwallace_cska24_and_15_2(.a(a[15]), .b(b[2]), .out(s_CSAwallace_cska24_and_15_2));
  and_gate and_gate_s_CSAwallace_cska24_and_16_2(.a(a[16]), .b(b[2]), .out(s_CSAwallace_cska24_and_16_2));
  and_gate and_gate_s_CSAwallace_cska24_and_17_2(.a(a[17]), .b(b[2]), .out(s_CSAwallace_cska24_and_17_2));
  and_gate and_gate_s_CSAwallace_cska24_and_18_2(.a(a[18]), .b(b[2]), .out(s_CSAwallace_cska24_and_18_2));
  and_gate and_gate_s_CSAwallace_cska24_and_19_2(.a(a[19]), .b(b[2]), .out(s_CSAwallace_cska24_and_19_2));
  and_gate and_gate_s_CSAwallace_cska24_and_20_2(.a(a[20]), .b(b[2]), .out(s_CSAwallace_cska24_and_20_2));
  and_gate and_gate_s_CSAwallace_cska24_and_21_2(.a(a[21]), .b(b[2]), .out(s_CSAwallace_cska24_and_21_2));
  and_gate and_gate_s_CSAwallace_cska24_and_22_2(.a(a[22]), .b(b[2]), .out(s_CSAwallace_cska24_and_22_2));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_2(.a(a[23]), .b(b[2]), .out(s_CSAwallace_cska24_nand_23_2));
  and_gate and_gate_s_CSAwallace_cska24_and_0_3(.a(a[0]), .b(b[3]), .out(s_CSAwallace_cska24_and_0_3));
  and_gate and_gate_s_CSAwallace_cska24_and_1_3(.a(a[1]), .b(b[3]), .out(s_CSAwallace_cska24_and_1_3));
  and_gate and_gate_s_CSAwallace_cska24_and_2_3(.a(a[2]), .b(b[3]), .out(s_CSAwallace_cska24_and_2_3));
  and_gate and_gate_s_CSAwallace_cska24_and_3_3(.a(a[3]), .b(b[3]), .out(s_CSAwallace_cska24_and_3_3));
  and_gate and_gate_s_CSAwallace_cska24_and_4_3(.a(a[4]), .b(b[3]), .out(s_CSAwallace_cska24_and_4_3));
  and_gate and_gate_s_CSAwallace_cska24_and_5_3(.a(a[5]), .b(b[3]), .out(s_CSAwallace_cska24_and_5_3));
  and_gate and_gate_s_CSAwallace_cska24_and_6_3(.a(a[6]), .b(b[3]), .out(s_CSAwallace_cska24_and_6_3));
  and_gate and_gate_s_CSAwallace_cska24_and_7_3(.a(a[7]), .b(b[3]), .out(s_CSAwallace_cska24_and_7_3));
  and_gate and_gate_s_CSAwallace_cska24_and_8_3(.a(a[8]), .b(b[3]), .out(s_CSAwallace_cska24_and_8_3));
  and_gate and_gate_s_CSAwallace_cska24_and_9_3(.a(a[9]), .b(b[3]), .out(s_CSAwallace_cska24_and_9_3));
  and_gate and_gate_s_CSAwallace_cska24_and_10_3(.a(a[10]), .b(b[3]), .out(s_CSAwallace_cska24_and_10_3));
  and_gate and_gate_s_CSAwallace_cska24_and_11_3(.a(a[11]), .b(b[3]), .out(s_CSAwallace_cska24_and_11_3));
  and_gate and_gate_s_CSAwallace_cska24_and_12_3(.a(a[12]), .b(b[3]), .out(s_CSAwallace_cska24_and_12_3));
  and_gate and_gate_s_CSAwallace_cska24_and_13_3(.a(a[13]), .b(b[3]), .out(s_CSAwallace_cska24_and_13_3));
  and_gate and_gate_s_CSAwallace_cska24_and_14_3(.a(a[14]), .b(b[3]), .out(s_CSAwallace_cska24_and_14_3));
  and_gate and_gate_s_CSAwallace_cska24_and_15_3(.a(a[15]), .b(b[3]), .out(s_CSAwallace_cska24_and_15_3));
  and_gate and_gate_s_CSAwallace_cska24_and_16_3(.a(a[16]), .b(b[3]), .out(s_CSAwallace_cska24_and_16_3));
  and_gate and_gate_s_CSAwallace_cska24_and_17_3(.a(a[17]), .b(b[3]), .out(s_CSAwallace_cska24_and_17_3));
  and_gate and_gate_s_CSAwallace_cska24_and_18_3(.a(a[18]), .b(b[3]), .out(s_CSAwallace_cska24_and_18_3));
  and_gate and_gate_s_CSAwallace_cska24_and_19_3(.a(a[19]), .b(b[3]), .out(s_CSAwallace_cska24_and_19_3));
  and_gate and_gate_s_CSAwallace_cska24_and_20_3(.a(a[20]), .b(b[3]), .out(s_CSAwallace_cska24_and_20_3));
  and_gate and_gate_s_CSAwallace_cska24_and_21_3(.a(a[21]), .b(b[3]), .out(s_CSAwallace_cska24_and_21_3));
  and_gate and_gate_s_CSAwallace_cska24_and_22_3(.a(a[22]), .b(b[3]), .out(s_CSAwallace_cska24_and_22_3));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_3(.a(a[23]), .b(b[3]), .out(s_CSAwallace_cska24_nand_23_3));
  and_gate and_gate_s_CSAwallace_cska24_and_0_4(.a(a[0]), .b(b[4]), .out(s_CSAwallace_cska24_and_0_4));
  and_gate and_gate_s_CSAwallace_cska24_and_1_4(.a(a[1]), .b(b[4]), .out(s_CSAwallace_cska24_and_1_4));
  and_gate and_gate_s_CSAwallace_cska24_and_2_4(.a(a[2]), .b(b[4]), .out(s_CSAwallace_cska24_and_2_4));
  and_gate and_gate_s_CSAwallace_cska24_and_3_4(.a(a[3]), .b(b[4]), .out(s_CSAwallace_cska24_and_3_4));
  and_gate and_gate_s_CSAwallace_cska24_and_4_4(.a(a[4]), .b(b[4]), .out(s_CSAwallace_cska24_and_4_4));
  and_gate and_gate_s_CSAwallace_cska24_and_5_4(.a(a[5]), .b(b[4]), .out(s_CSAwallace_cska24_and_5_4));
  and_gate and_gate_s_CSAwallace_cska24_and_6_4(.a(a[6]), .b(b[4]), .out(s_CSAwallace_cska24_and_6_4));
  and_gate and_gate_s_CSAwallace_cska24_and_7_4(.a(a[7]), .b(b[4]), .out(s_CSAwallace_cska24_and_7_4));
  and_gate and_gate_s_CSAwallace_cska24_and_8_4(.a(a[8]), .b(b[4]), .out(s_CSAwallace_cska24_and_8_4));
  and_gate and_gate_s_CSAwallace_cska24_and_9_4(.a(a[9]), .b(b[4]), .out(s_CSAwallace_cska24_and_9_4));
  and_gate and_gate_s_CSAwallace_cska24_and_10_4(.a(a[10]), .b(b[4]), .out(s_CSAwallace_cska24_and_10_4));
  and_gate and_gate_s_CSAwallace_cska24_and_11_4(.a(a[11]), .b(b[4]), .out(s_CSAwallace_cska24_and_11_4));
  and_gate and_gate_s_CSAwallace_cska24_and_12_4(.a(a[12]), .b(b[4]), .out(s_CSAwallace_cska24_and_12_4));
  and_gate and_gate_s_CSAwallace_cska24_and_13_4(.a(a[13]), .b(b[4]), .out(s_CSAwallace_cska24_and_13_4));
  and_gate and_gate_s_CSAwallace_cska24_and_14_4(.a(a[14]), .b(b[4]), .out(s_CSAwallace_cska24_and_14_4));
  and_gate and_gate_s_CSAwallace_cska24_and_15_4(.a(a[15]), .b(b[4]), .out(s_CSAwallace_cska24_and_15_4));
  and_gate and_gate_s_CSAwallace_cska24_and_16_4(.a(a[16]), .b(b[4]), .out(s_CSAwallace_cska24_and_16_4));
  and_gate and_gate_s_CSAwallace_cska24_and_17_4(.a(a[17]), .b(b[4]), .out(s_CSAwallace_cska24_and_17_4));
  and_gate and_gate_s_CSAwallace_cska24_and_18_4(.a(a[18]), .b(b[4]), .out(s_CSAwallace_cska24_and_18_4));
  and_gate and_gate_s_CSAwallace_cska24_and_19_4(.a(a[19]), .b(b[4]), .out(s_CSAwallace_cska24_and_19_4));
  and_gate and_gate_s_CSAwallace_cska24_and_20_4(.a(a[20]), .b(b[4]), .out(s_CSAwallace_cska24_and_20_4));
  and_gate and_gate_s_CSAwallace_cska24_and_21_4(.a(a[21]), .b(b[4]), .out(s_CSAwallace_cska24_and_21_4));
  and_gate and_gate_s_CSAwallace_cska24_and_22_4(.a(a[22]), .b(b[4]), .out(s_CSAwallace_cska24_and_22_4));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_4(.a(a[23]), .b(b[4]), .out(s_CSAwallace_cska24_nand_23_4));
  and_gate and_gate_s_CSAwallace_cska24_and_0_5(.a(a[0]), .b(b[5]), .out(s_CSAwallace_cska24_and_0_5));
  and_gate and_gate_s_CSAwallace_cska24_and_1_5(.a(a[1]), .b(b[5]), .out(s_CSAwallace_cska24_and_1_5));
  and_gate and_gate_s_CSAwallace_cska24_and_2_5(.a(a[2]), .b(b[5]), .out(s_CSAwallace_cska24_and_2_5));
  and_gate and_gate_s_CSAwallace_cska24_and_3_5(.a(a[3]), .b(b[5]), .out(s_CSAwallace_cska24_and_3_5));
  and_gate and_gate_s_CSAwallace_cska24_and_4_5(.a(a[4]), .b(b[5]), .out(s_CSAwallace_cska24_and_4_5));
  and_gate and_gate_s_CSAwallace_cska24_and_5_5(.a(a[5]), .b(b[5]), .out(s_CSAwallace_cska24_and_5_5));
  and_gate and_gate_s_CSAwallace_cska24_and_6_5(.a(a[6]), .b(b[5]), .out(s_CSAwallace_cska24_and_6_5));
  and_gate and_gate_s_CSAwallace_cska24_and_7_5(.a(a[7]), .b(b[5]), .out(s_CSAwallace_cska24_and_7_5));
  and_gate and_gate_s_CSAwallace_cska24_and_8_5(.a(a[8]), .b(b[5]), .out(s_CSAwallace_cska24_and_8_5));
  and_gate and_gate_s_CSAwallace_cska24_and_9_5(.a(a[9]), .b(b[5]), .out(s_CSAwallace_cska24_and_9_5));
  and_gate and_gate_s_CSAwallace_cska24_and_10_5(.a(a[10]), .b(b[5]), .out(s_CSAwallace_cska24_and_10_5));
  and_gate and_gate_s_CSAwallace_cska24_and_11_5(.a(a[11]), .b(b[5]), .out(s_CSAwallace_cska24_and_11_5));
  and_gate and_gate_s_CSAwallace_cska24_and_12_5(.a(a[12]), .b(b[5]), .out(s_CSAwallace_cska24_and_12_5));
  and_gate and_gate_s_CSAwallace_cska24_and_13_5(.a(a[13]), .b(b[5]), .out(s_CSAwallace_cska24_and_13_5));
  and_gate and_gate_s_CSAwallace_cska24_and_14_5(.a(a[14]), .b(b[5]), .out(s_CSAwallace_cska24_and_14_5));
  and_gate and_gate_s_CSAwallace_cska24_and_15_5(.a(a[15]), .b(b[5]), .out(s_CSAwallace_cska24_and_15_5));
  and_gate and_gate_s_CSAwallace_cska24_and_16_5(.a(a[16]), .b(b[5]), .out(s_CSAwallace_cska24_and_16_5));
  and_gate and_gate_s_CSAwallace_cska24_and_17_5(.a(a[17]), .b(b[5]), .out(s_CSAwallace_cska24_and_17_5));
  and_gate and_gate_s_CSAwallace_cska24_and_18_5(.a(a[18]), .b(b[5]), .out(s_CSAwallace_cska24_and_18_5));
  and_gate and_gate_s_CSAwallace_cska24_and_19_5(.a(a[19]), .b(b[5]), .out(s_CSAwallace_cska24_and_19_5));
  and_gate and_gate_s_CSAwallace_cska24_and_20_5(.a(a[20]), .b(b[5]), .out(s_CSAwallace_cska24_and_20_5));
  and_gate and_gate_s_CSAwallace_cska24_and_21_5(.a(a[21]), .b(b[5]), .out(s_CSAwallace_cska24_and_21_5));
  and_gate and_gate_s_CSAwallace_cska24_and_22_5(.a(a[22]), .b(b[5]), .out(s_CSAwallace_cska24_and_22_5));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_5(.a(a[23]), .b(b[5]), .out(s_CSAwallace_cska24_nand_23_5));
  and_gate and_gate_s_CSAwallace_cska24_and_0_6(.a(a[0]), .b(b[6]), .out(s_CSAwallace_cska24_and_0_6));
  and_gate and_gate_s_CSAwallace_cska24_and_1_6(.a(a[1]), .b(b[6]), .out(s_CSAwallace_cska24_and_1_6));
  and_gate and_gate_s_CSAwallace_cska24_and_2_6(.a(a[2]), .b(b[6]), .out(s_CSAwallace_cska24_and_2_6));
  and_gate and_gate_s_CSAwallace_cska24_and_3_6(.a(a[3]), .b(b[6]), .out(s_CSAwallace_cska24_and_3_6));
  and_gate and_gate_s_CSAwallace_cska24_and_4_6(.a(a[4]), .b(b[6]), .out(s_CSAwallace_cska24_and_4_6));
  and_gate and_gate_s_CSAwallace_cska24_and_5_6(.a(a[5]), .b(b[6]), .out(s_CSAwallace_cska24_and_5_6));
  and_gate and_gate_s_CSAwallace_cska24_and_6_6(.a(a[6]), .b(b[6]), .out(s_CSAwallace_cska24_and_6_6));
  and_gate and_gate_s_CSAwallace_cska24_and_7_6(.a(a[7]), .b(b[6]), .out(s_CSAwallace_cska24_and_7_6));
  and_gate and_gate_s_CSAwallace_cska24_and_8_6(.a(a[8]), .b(b[6]), .out(s_CSAwallace_cska24_and_8_6));
  and_gate and_gate_s_CSAwallace_cska24_and_9_6(.a(a[9]), .b(b[6]), .out(s_CSAwallace_cska24_and_9_6));
  and_gate and_gate_s_CSAwallace_cska24_and_10_6(.a(a[10]), .b(b[6]), .out(s_CSAwallace_cska24_and_10_6));
  and_gate and_gate_s_CSAwallace_cska24_and_11_6(.a(a[11]), .b(b[6]), .out(s_CSAwallace_cska24_and_11_6));
  and_gate and_gate_s_CSAwallace_cska24_and_12_6(.a(a[12]), .b(b[6]), .out(s_CSAwallace_cska24_and_12_6));
  and_gate and_gate_s_CSAwallace_cska24_and_13_6(.a(a[13]), .b(b[6]), .out(s_CSAwallace_cska24_and_13_6));
  and_gate and_gate_s_CSAwallace_cska24_and_14_6(.a(a[14]), .b(b[6]), .out(s_CSAwallace_cska24_and_14_6));
  and_gate and_gate_s_CSAwallace_cska24_and_15_6(.a(a[15]), .b(b[6]), .out(s_CSAwallace_cska24_and_15_6));
  and_gate and_gate_s_CSAwallace_cska24_and_16_6(.a(a[16]), .b(b[6]), .out(s_CSAwallace_cska24_and_16_6));
  and_gate and_gate_s_CSAwallace_cska24_and_17_6(.a(a[17]), .b(b[6]), .out(s_CSAwallace_cska24_and_17_6));
  and_gate and_gate_s_CSAwallace_cska24_and_18_6(.a(a[18]), .b(b[6]), .out(s_CSAwallace_cska24_and_18_6));
  and_gate and_gate_s_CSAwallace_cska24_and_19_6(.a(a[19]), .b(b[6]), .out(s_CSAwallace_cska24_and_19_6));
  and_gate and_gate_s_CSAwallace_cska24_and_20_6(.a(a[20]), .b(b[6]), .out(s_CSAwallace_cska24_and_20_6));
  and_gate and_gate_s_CSAwallace_cska24_and_21_6(.a(a[21]), .b(b[6]), .out(s_CSAwallace_cska24_and_21_6));
  and_gate and_gate_s_CSAwallace_cska24_and_22_6(.a(a[22]), .b(b[6]), .out(s_CSAwallace_cska24_and_22_6));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_6(.a(a[23]), .b(b[6]), .out(s_CSAwallace_cska24_nand_23_6));
  and_gate and_gate_s_CSAwallace_cska24_and_0_7(.a(a[0]), .b(b[7]), .out(s_CSAwallace_cska24_and_0_7));
  and_gate and_gate_s_CSAwallace_cska24_and_1_7(.a(a[1]), .b(b[7]), .out(s_CSAwallace_cska24_and_1_7));
  and_gate and_gate_s_CSAwallace_cska24_and_2_7(.a(a[2]), .b(b[7]), .out(s_CSAwallace_cska24_and_2_7));
  and_gate and_gate_s_CSAwallace_cska24_and_3_7(.a(a[3]), .b(b[7]), .out(s_CSAwallace_cska24_and_3_7));
  and_gate and_gate_s_CSAwallace_cska24_and_4_7(.a(a[4]), .b(b[7]), .out(s_CSAwallace_cska24_and_4_7));
  and_gate and_gate_s_CSAwallace_cska24_and_5_7(.a(a[5]), .b(b[7]), .out(s_CSAwallace_cska24_and_5_7));
  and_gate and_gate_s_CSAwallace_cska24_and_6_7(.a(a[6]), .b(b[7]), .out(s_CSAwallace_cska24_and_6_7));
  and_gate and_gate_s_CSAwallace_cska24_and_7_7(.a(a[7]), .b(b[7]), .out(s_CSAwallace_cska24_and_7_7));
  and_gate and_gate_s_CSAwallace_cska24_and_8_7(.a(a[8]), .b(b[7]), .out(s_CSAwallace_cska24_and_8_7));
  and_gate and_gate_s_CSAwallace_cska24_and_9_7(.a(a[9]), .b(b[7]), .out(s_CSAwallace_cska24_and_9_7));
  and_gate and_gate_s_CSAwallace_cska24_and_10_7(.a(a[10]), .b(b[7]), .out(s_CSAwallace_cska24_and_10_7));
  and_gate and_gate_s_CSAwallace_cska24_and_11_7(.a(a[11]), .b(b[7]), .out(s_CSAwallace_cska24_and_11_7));
  and_gate and_gate_s_CSAwallace_cska24_and_12_7(.a(a[12]), .b(b[7]), .out(s_CSAwallace_cska24_and_12_7));
  and_gate and_gate_s_CSAwallace_cska24_and_13_7(.a(a[13]), .b(b[7]), .out(s_CSAwallace_cska24_and_13_7));
  and_gate and_gate_s_CSAwallace_cska24_and_14_7(.a(a[14]), .b(b[7]), .out(s_CSAwallace_cska24_and_14_7));
  and_gate and_gate_s_CSAwallace_cska24_and_15_7(.a(a[15]), .b(b[7]), .out(s_CSAwallace_cska24_and_15_7));
  and_gate and_gate_s_CSAwallace_cska24_and_16_7(.a(a[16]), .b(b[7]), .out(s_CSAwallace_cska24_and_16_7));
  and_gate and_gate_s_CSAwallace_cska24_and_17_7(.a(a[17]), .b(b[7]), .out(s_CSAwallace_cska24_and_17_7));
  and_gate and_gate_s_CSAwallace_cska24_and_18_7(.a(a[18]), .b(b[7]), .out(s_CSAwallace_cska24_and_18_7));
  and_gate and_gate_s_CSAwallace_cska24_and_19_7(.a(a[19]), .b(b[7]), .out(s_CSAwallace_cska24_and_19_7));
  and_gate and_gate_s_CSAwallace_cska24_and_20_7(.a(a[20]), .b(b[7]), .out(s_CSAwallace_cska24_and_20_7));
  and_gate and_gate_s_CSAwallace_cska24_and_21_7(.a(a[21]), .b(b[7]), .out(s_CSAwallace_cska24_and_21_7));
  and_gate and_gate_s_CSAwallace_cska24_and_22_7(.a(a[22]), .b(b[7]), .out(s_CSAwallace_cska24_and_22_7));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_7(.a(a[23]), .b(b[7]), .out(s_CSAwallace_cska24_nand_23_7));
  and_gate and_gate_s_CSAwallace_cska24_and_0_8(.a(a[0]), .b(b[8]), .out(s_CSAwallace_cska24_and_0_8));
  and_gate and_gate_s_CSAwallace_cska24_and_1_8(.a(a[1]), .b(b[8]), .out(s_CSAwallace_cska24_and_1_8));
  and_gate and_gate_s_CSAwallace_cska24_and_2_8(.a(a[2]), .b(b[8]), .out(s_CSAwallace_cska24_and_2_8));
  and_gate and_gate_s_CSAwallace_cska24_and_3_8(.a(a[3]), .b(b[8]), .out(s_CSAwallace_cska24_and_3_8));
  and_gate and_gate_s_CSAwallace_cska24_and_4_8(.a(a[4]), .b(b[8]), .out(s_CSAwallace_cska24_and_4_8));
  and_gate and_gate_s_CSAwallace_cska24_and_5_8(.a(a[5]), .b(b[8]), .out(s_CSAwallace_cska24_and_5_8));
  and_gate and_gate_s_CSAwallace_cska24_and_6_8(.a(a[6]), .b(b[8]), .out(s_CSAwallace_cska24_and_6_8));
  and_gate and_gate_s_CSAwallace_cska24_and_7_8(.a(a[7]), .b(b[8]), .out(s_CSAwallace_cska24_and_7_8));
  and_gate and_gate_s_CSAwallace_cska24_and_8_8(.a(a[8]), .b(b[8]), .out(s_CSAwallace_cska24_and_8_8));
  and_gate and_gate_s_CSAwallace_cska24_and_9_8(.a(a[9]), .b(b[8]), .out(s_CSAwallace_cska24_and_9_8));
  and_gate and_gate_s_CSAwallace_cska24_and_10_8(.a(a[10]), .b(b[8]), .out(s_CSAwallace_cska24_and_10_8));
  and_gate and_gate_s_CSAwallace_cska24_and_11_8(.a(a[11]), .b(b[8]), .out(s_CSAwallace_cska24_and_11_8));
  and_gate and_gate_s_CSAwallace_cska24_and_12_8(.a(a[12]), .b(b[8]), .out(s_CSAwallace_cska24_and_12_8));
  and_gate and_gate_s_CSAwallace_cska24_and_13_8(.a(a[13]), .b(b[8]), .out(s_CSAwallace_cska24_and_13_8));
  and_gate and_gate_s_CSAwallace_cska24_and_14_8(.a(a[14]), .b(b[8]), .out(s_CSAwallace_cska24_and_14_8));
  and_gate and_gate_s_CSAwallace_cska24_and_15_8(.a(a[15]), .b(b[8]), .out(s_CSAwallace_cska24_and_15_8));
  and_gate and_gate_s_CSAwallace_cska24_and_16_8(.a(a[16]), .b(b[8]), .out(s_CSAwallace_cska24_and_16_8));
  and_gate and_gate_s_CSAwallace_cska24_and_17_8(.a(a[17]), .b(b[8]), .out(s_CSAwallace_cska24_and_17_8));
  and_gate and_gate_s_CSAwallace_cska24_and_18_8(.a(a[18]), .b(b[8]), .out(s_CSAwallace_cska24_and_18_8));
  and_gate and_gate_s_CSAwallace_cska24_and_19_8(.a(a[19]), .b(b[8]), .out(s_CSAwallace_cska24_and_19_8));
  and_gate and_gate_s_CSAwallace_cska24_and_20_8(.a(a[20]), .b(b[8]), .out(s_CSAwallace_cska24_and_20_8));
  and_gate and_gate_s_CSAwallace_cska24_and_21_8(.a(a[21]), .b(b[8]), .out(s_CSAwallace_cska24_and_21_8));
  and_gate and_gate_s_CSAwallace_cska24_and_22_8(.a(a[22]), .b(b[8]), .out(s_CSAwallace_cska24_and_22_8));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_8(.a(a[23]), .b(b[8]), .out(s_CSAwallace_cska24_nand_23_8));
  and_gate and_gate_s_CSAwallace_cska24_and_0_9(.a(a[0]), .b(b[9]), .out(s_CSAwallace_cska24_and_0_9));
  and_gate and_gate_s_CSAwallace_cska24_and_1_9(.a(a[1]), .b(b[9]), .out(s_CSAwallace_cska24_and_1_9));
  and_gate and_gate_s_CSAwallace_cska24_and_2_9(.a(a[2]), .b(b[9]), .out(s_CSAwallace_cska24_and_2_9));
  and_gate and_gate_s_CSAwallace_cska24_and_3_9(.a(a[3]), .b(b[9]), .out(s_CSAwallace_cska24_and_3_9));
  and_gate and_gate_s_CSAwallace_cska24_and_4_9(.a(a[4]), .b(b[9]), .out(s_CSAwallace_cska24_and_4_9));
  and_gate and_gate_s_CSAwallace_cska24_and_5_9(.a(a[5]), .b(b[9]), .out(s_CSAwallace_cska24_and_5_9));
  and_gate and_gate_s_CSAwallace_cska24_and_6_9(.a(a[6]), .b(b[9]), .out(s_CSAwallace_cska24_and_6_9));
  and_gate and_gate_s_CSAwallace_cska24_and_7_9(.a(a[7]), .b(b[9]), .out(s_CSAwallace_cska24_and_7_9));
  and_gate and_gate_s_CSAwallace_cska24_and_8_9(.a(a[8]), .b(b[9]), .out(s_CSAwallace_cska24_and_8_9));
  and_gate and_gate_s_CSAwallace_cska24_and_9_9(.a(a[9]), .b(b[9]), .out(s_CSAwallace_cska24_and_9_9));
  and_gate and_gate_s_CSAwallace_cska24_and_10_9(.a(a[10]), .b(b[9]), .out(s_CSAwallace_cska24_and_10_9));
  and_gate and_gate_s_CSAwallace_cska24_and_11_9(.a(a[11]), .b(b[9]), .out(s_CSAwallace_cska24_and_11_9));
  and_gate and_gate_s_CSAwallace_cska24_and_12_9(.a(a[12]), .b(b[9]), .out(s_CSAwallace_cska24_and_12_9));
  and_gate and_gate_s_CSAwallace_cska24_and_13_9(.a(a[13]), .b(b[9]), .out(s_CSAwallace_cska24_and_13_9));
  and_gate and_gate_s_CSAwallace_cska24_and_14_9(.a(a[14]), .b(b[9]), .out(s_CSAwallace_cska24_and_14_9));
  and_gate and_gate_s_CSAwallace_cska24_and_15_9(.a(a[15]), .b(b[9]), .out(s_CSAwallace_cska24_and_15_9));
  and_gate and_gate_s_CSAwallace_cska24_and_16_9(.a(a[16]), .b(b[9]), .out(s_CSAwallace_cska24_and_16_9));
  and_gate and_gate_s_CSAwallace_cska24_and_17_9(.a(a[17]), .b(b[9]), .out(s_CSAwallace_cska24_and_17_9));
  and_gate and_gate_s_CSAwallace_cska24_and_18_9(.a(a[18]), .b(b[9]), .out(s_CSAwallace_cska24_and_18_9));
  and_gate and_gate_s_CSAwallace_cska24_and_19_9(.a(a[19]), .b(b[9]), .out(s_CSAwallace_cska24_and_19_9));
  and_gate and_gate_s_CSAwallace_cska24_and_20_9(.a(a[20]), .b(b[9]), .out(s_CSAwallace_cska24_and_20_9));
  and_gate and_gate_s_CSAwallace_cska24_and_21_9(.a(a[21]), .b(b[9]), .out(s_CSAwallace_cska24_and_21_9));
  and_gate and_gate_s_CSAwallace_cska24_and_22_9(.a(a[22]), .b(b[9]), .out(s_CSAwallace_cska24_and_22_9));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_9(.a(a[23]), .b(b[9]), .out(s_CSAwallace_cska24_nand_23_9));
  and_gate and_gate_s_CSAwallace_cska24_and_0_10(.a(a[0]), .b(b[10]), .out(s_CSAwallace_cska24_and_0_10));
  and_gate and_gate_s_CSAwallace_cska24_and_1_10(.a(a[1]), .b(b[10]), .out(s_CSAwallace_cska24_and_1_10));
  and_gate and_gate_s_CSAwallace_cska24_and_2_10(.a(a[2]), .b(b[10]), .out(s_CSAwallace_cska24_and_2_10));
  and_gate and_gate_s_CSAwallace_cska24_and_3_10(.a(a[3]), .b(b[10]), .out(s_CSAwallace_cska24_and_3_10));
  and_gate and_gate_s_CSAwallace_cska24_and_4_10(.a(a[4]), .b(b[10]), .out(s_CSAwallace_cska24_and_4_10));
  and_gate and_gate_s_CSAwallace_cska24_and_5_10(.a(a[5]), .b(b[10]), .out(s_CSAwallace_cska24_and_5_10));
  and_gate and_gate_s_CSAwallace_cska24_and_6_10(.a(a[6]), .b(b[10]), .out(s_CSAwallace_cska24_and_6_10));
  and_gate and_gate_s_CSAwallace_cska24_and_7_10(.a(a[7]), .b(b[10]), .out(s_CSAwallace_cska24_and_7_10));
  and_gate and_gate_s_CSAwallace_cska24_and_8_10(.a(a[8]), .b(b[10]), .out(s_CSAwallace_cska24_and_8_10));
  and_gate and_gate_s_CSAwallace_cska24_and_9_10(.a(a[9]), .b(b[10]), .out(s_CSAwallace_cska24_and_9_10));
  and_gate and_gate_s_CSAwallace_cska24_and_10_10(.a(a[10]), .b(b[10]), .out(s_CSAwallace_cska24_and_10_10));
  and_gate and_gate_s_CSAwallace_cska24_and_11_10(.a(a[11]), .b(b[10]), .out(s_CSAwallace_cska24_and_11_10));
  and_gate and_gate_s_CSAwallace_cska24_and_12_10(.a(a[12]), .b(b[10]), .out(s_CSAwallace_cska24_and_12_10));
  and_gate and_gate_s_CSAwallace_cska24_and_13_10(.a(a[13]), .b(b[10]), .out(s_CSAwallace_cska24_and_13_10));
  and_gate and_gate_s_CSAwallace_cska24_and_14_10(.a(a[14]), .b(b[10]), .out(s_CSAwallace_cska24_and_14_10));
  and_gate and_gate_s_CSAwallace_cska24_and_15_10(.a(a[15]), .b(b[10]), .out(s_CSAwallace_cska24_and_15_10));
  and_gate and_gate_s_CSAwallace_cska24_and_16_10(.a(a[16]), .b(b[10]), .out(s_CSAwallace_cska24_and_16_10));
  and_gate and_gate_s_CSAwallace_cska24_and_17_10(.a(a[17]), .b(b[10]), .out(s_CSAwallace_cska24_and_17_10));
  and_gate and_gate_s_CSAwallace_cska24_and_18_10(.a(a[18]), .b(b[10]), .out(s_CSAwallace_cska24_and_18_10));
  and_gate and_gate_s_CSAwallace_cska24_and_19_10(.a(a[19]), .b(b[10]), .out(s_CSAwallace_cska24_and_19_10));
  and_gate and_gate_s_CSAwallace_cska24_and_20_10(.a(a[20]), .b(b[10]), .out(s_CSAwallace_cska24_and_20_10));
  and_gate and_gate_s_CSAwallace_cska24_and_21_10(.a(a[21]), .b(b[10]), .out(s_CSAwallace_cska24_and_21_10));
  and_gate and_gate_s_CSAwallace_cska24_and_22_10(.a(a[22]), .b(b[10]), .out(s_CSAwallace_cska24_and_22_10));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_10(.a(a[23]), .b(b[10]), .out(s_CSAwallace_cska24_nand_23_10));
  and_gate and_gate_s_CSAwallace_cska24_and_0_11(.a(a[0]), .b(b[11]), .out(s_CSAwallace_cska24_and_0_11));
  and_gate and_gate_s_CSAwallace_cska24_and_1_11(.a(a[1]), .b(b[11]), .out(s_CSAwallace_cska24_and_1_11));
  and_gate and_gate_s_CSAwallace_cska24_and_2_11(.a(a[2]), .b(b[11]), .out(s_CSAwallace_cska24_and_2_11));
  and_gate and_gate_s_CSAwallace_cska24_and_3_11(.a(a[3]), .b(b[11]), .out(s_CSAwallace_cska24_and_3_11));
  and_gate and_gate_s_CSAwallace_cska24_and_4_11(.a(a[4]), .b(b[11]), .out(s_CSAwallace_cska24_and_4_11));
  and_gate and_gate_s_CSAwallace_cska24_and_5_11(.a(a[5]), .b(b[11]), .out(s_CSAwallace_cska24_and_5_11));
  and_gate and_gate_s_CSAwallace_cska24_and_6_11(.a(a[6]), .b(b[11]), .out(s_CSAwallace_cska24_and_6_11));
  and_gate and_gate_s_CSAwallace_cska24_and_7_11(.a(a[7]), .b(b[11]), .out(s_CSAwallace_cska24_and_7_11));
  and_gate and_gate_s_CSAwallace_cska24_and_8_11(.a(a[8]), .b(b[11]), .out(s_CSAwallace_cska24_and_8_11));
  and_gate and_gate_s_CSAwallace_cska24_and_9_11(.a(a[9]), .b(b[11]), .out(s_CSAwallace_cska24_and_9_11));
  and_gate and_gate_s_CSAwallace_cska24_and_10_11(.a(a[10]), .b(b[11]), .out(s_CSAwallace_cska24_and_10_11));
  and_gate and_gate_s_CSAwallace_cska24_and_11_11(.a(a[11]), .b(b[11]), .out(s_CSAwallace_cska24_and_11_11));
  and_gate and_gate_s_CSAwallace_cska24_and_12_11(.a(a[12]), .b(b[11]), .out(s_CSAwallace_cska24_and_12_11));
  and_gate and_gate_s_CSAwallace_cska24_and_13_11(.a(a[13]), .b(b[11]), .out(s_CSAwallace_cska24_and_13_11));
  and_gate and_gate_s_CSAwallace_cska24_and_14_11(.a(a[14]), .b(b[11]), .out(s_CSAwallace_cska24_and_14_11));
  and_gate and_gate_s_CSAwallace_cska24_and_15_11(.a(a[15]), .b(b[11]), .out(s_CSAwallace_cska24_and_15_11));
  and_gate and_gate_s_CSAwallace_cska24_and_16_11(.a(a[16]), .b(b[11]), .out(s_CSAwallace_cska24_and_16_11));
  and_gate and_gate_s_CSAwallace_cska24_and_17_11(.a(a[17]), .b(b[11]), .out(s_CSAwallace_cska24_and_17_11));
  and_gate and_gate_s_CSAwallace_cska24_and_18_11(.a(a[18]), .b(b[11]), .out(s_CSAwallace_cska24_and_18_11));
  and_gate and_gate_s_CSAwallace_cska24_and_19_11(.a(a[19]), .b(b[11]), .out(s_CSAwallace_cska24_and_19_11));
  and_gate and_gate_s_CSAwallace_cska24_and_20_11(.a(a[20]), .b(b[11]), .out(s_CSAwallace_cska24_and_20_11));
  and_gate and_gate_s_CSAwallace_cska24_and_21_11(.a(a[21]), .b(b[11]), .out(s_CSAwallace_cska24_and_21_11));
  and_gate and_gate_s_CSAwallace_cska24_and_22_11(.a(a[22]), .b(b[11]), .out(s_CSAwallace_cska24_and_22_11));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_11(.a(a[23]), .b(b[11]), .out(s_CSAwallace_cska24_nand_23_11));
  and_gate and_gate_s_CSAwallace_cska24_and_0_12(.a(a[0]), .b(b[12]), .out(s_CSAwallace_cska24_and_0_12));
  and_gate and_gate_s_CSAwallace_cska24_and_1_12(.a(a[1]), .b(b[12]), .out(s_CSAwallace_cska24_and_1_12));
  and_gate and_gate_s_CSAwallace_cska24_and_2_12(.a(a[2]), .b(b[12]), .out(s_CSAwallace_cska24_and_2_12));
  and_gate and_gate_s_CSAwallace_cska24_and_3_12(.a(a[3]), .b(b[12]), .out(s_CSAwallace_cska24_and_3_12));
  and_gate and_gate_s_CSAwallace_cska24_and_4_12(.a(a[4]), .b(b[12]), .out(s_CSAwallace_cska24_and_4_12));
  and_gate and_gate_s_CSAwallace_cska24_and_5_12(.a(a[5]), .b(b[12]), .out(s_CSAwallace_cska24_and_5_12));
  and_gate and_gate_s_CSAwallace_cska24_and_6_12(.a(a[6]), .b(b[12]), .out(s_CSAwallace_cska24_and_6_12));
  and_gate and_gate_s_CSAwallace_cska24_and_7_12(.a(a[7]), .b(b[12]), .out(s_CSAwallace_cska24_and_7_12));
  and_gate and_gate_s_CSAwallace_cska24_and_8_12(.a(a[8]), .b(b[12]), .out(s_CSAwallace_cska24_and_8_12));
  and_gate and_gate_s_CSAwallace_cska24_and_9_12(.a(a[9]), .b(b[12]), .out(s_CSAwallace_cska24_and_9_12));
  and_gate and_gate_s_CSAwallace_cska24_and_10_12(.a(a[10]), .b(b[12]), .out(s_CSAwallace_cska24_and_10_12));
  and_gate and_gate_s_CSAwallace_cska24_and_11_12(.a(a[11]), .b(b[12]), .out(s_CSAwallace_cska24_and_11_12));
  and_gate and_gate_s_CSAwallace_cska24_and_12_12(.a(a[12]), .b(b[12]), .out(s_CSAwallace_cska24_and_12_12));
  and_gate and_gate_s_CSAwallace_cska24_and_13_12(.a(a[13]), .b(b[12]), .out(s_CSAwallace_cska24_and_13_12));
  and_gate and_gate_s_CSAwallace_cska24_and_14_12(.a(a[14]), .b(b[12]), .out(s_CSAwallace_cska24_and_14_12));
  and_gate and_gate_s_CSAwallace_cska24_and_15_12(.a(a[15]), .b(b[12]), .out(s_CSAwallace_cska24_and_15_12));
  and_gate and_gate_s_CSAwallace_cska24_and_16_12(.a(a[16]), .b(b[12]), .out(s_CSAwallace_cska24_and_16_12));
  and_gate and_gate_s_CSAwallace_cska24_and_17_12(.a(a[17]), .b(b[12]), .out(s_CSAwallace_cska24_and_17_12));
  and_gate and_gate_s_CSAwallace_cska24_and_18_12(.a(a[18]), .b(b[12]), .out(s_CSAwallace_cska24_and_18_12));
  and_gate and_gate_s_CSAwallace_cska24_and_19_12(.a(a[19]), .b(b[12]), .out(s_CSAwallace_cska24_and_19_12));
  and_gate and_gate_s_CSAwallace_cska24_and_20_12(.a(a[20]), .b(b[12]), .out(s_CSAwallace_cska24_and_20_12));
  and_gate and_gate_s_CSAwallace_cska24_and_21_12(.a(a[21]), .b(b[12]), .out(s_CSAwallace_cska24_and_21_12));
  and_gate and_gate_s_CSAwallace_cska24_and_22_12(.a(a[22]), .b(b[12]), .out(s_CSAwallace_cska24_and_22_12));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_12(.a(a[23]), .b(b[12]), .out(s_CSAwallace_cska24_nand_23_12));
  and_gate and_gate_s_CSAwallace_cska24_and_0_13(.a(a[0]), .b(b[13]), .out(s_CSAwallace_cska24_and_0_13));
  and_gate and_gate_s_CSAwallace_cska24_and_1_13(.a(a[1]), .b(b[13]), .out(s_CSAwallace_cska24_and_1_13));
  and_gate and_gate_s_CSAwallace_cska24_and_2_13(.a(a[2]), .b(b[13]), .out(s_CSAwallace_cska24_and_2_13));
  and_gate and_gate_s_CSAwallace_cska24_and_3_13(.a(a[3]), .b(b[13]), .out(s_CSAwallace_cska24_and_3_13));
  and_gate and_gate_s_CSAwallace_cska24_and_4_13(.a(a[4]), .b(b[13]), .out(s_CSAwallace_cska24_and_4_13));
  and_gate and_gate_s_CSAwallace_cska24_and_5_13(.a(a[5]), .b(b[13]), .out(s_CSAwallace_cska24_and_5_13));
  and_gate and_gate_s_CSAwallace_cska24_and_6_13(.a(a[6]), .b(b[13]), .out(s_CSAwallace_cska24_and_6_13));
  and_gate and_gate_s_CSAwallace_cska24_and_7_13(.a(a[7]), .b(b[13]), .out(s_CSAwallace_cska24_and_7_13));
  and_gate and_gate_s_CSAwallace_cska24_and_8_13(.a(a[8]), .b(b[13]), .out(s_CSAwallace_cska24_and_8_13));
  and_gate and_gate_s_CSAwallace_cska24_and_9_13(.a(a[9]), .b(b[13]), .out(s_CSAwallace_cska24_and_9_13));
  and_gate and_gate_s_CSAwallace_cska24_and_10_13(.a(a[10]), .b(b[13]), .out(s_CSAwallace_cska24_and_10_13));
  and_gate and_gate_s_CSAwallace_cska24_and_11_13(.a(a[11]), .b(b[13]), .out(s_CSAwallace_cska24_and_11_13));
  and_gate and_gate_s_CSAwallace_cska24_and_12_13(.a(a[12]), .b(b[13]), .out(s_CSAwallace_cska24_and_12_13));
  and_gate and_gate_s_CSAwallace_cska24_and_13_13(.a(a[13]), .b(b[13]), .out(s_CSAwallace_cska24_and_13_13));
  and_gate and_gate_s_CSAwallace_cska24_and_14_13(.a(a[14]), .b(b[13]), .out(s_CSAwallace_cska24_and_14_13));
  and_gate and_gate_s_CSAwallace_cska24_and_15_13(.a(a[15]), .b(b[13]), .out(s_CSAwallace_cska24_and_15_13));
  and_gate and_gate_s_CSAwallace_cska24_and_16_13(.a(a[16]), .b(b[13]), .out(s_CSAwallace_cska24_and_16_13));
  and_gate and_gate_s_CSAwallace_cska24_and_17_13(.a(a[17]), .b(b[13]), .out(s_CSAwallace_cska24_and_17_13));
  and_gate and_gate_s_CSAwallace_cska24_and_18_13(.a(a[18]), .b(b[13]), .out(s_CSAwallace_cska24_and_18_13));
  and_gate and_gate_s_CSAwallace_cska24_and_19_13(.a(a[19]), .b(b[13]), .out(s_CSAwallace_cska24_and_19_13));
  and_gate and_gate_s_CSAwallace_cska24_and_20_13(.a(a[20]), .b(b[13]), .out(s_CSAwallace_cska24_and_20_13));
  and_gate and_gate_s_CSAwallace_cska24_and_21_13(.a(a[21]), .b(b[13]), .out(s_CSAwallace_cska24_and_21_13));
  and_gate and_gate_s_CSAwallace_cska24_and_22_13(.a(a[22]), .b(b[13]), .out(s_CSAwallace_cska24_and_22_13));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_13(.a(a[23]), .b(b[13]), .out(s_CSAwallace_cska24_nand_23_13));
  and_gate and_gate_s_CSAwallace_cska24_and_0_14(.a(a[0]), .b(b[14]), .out(s_CSAwallace_cska24_and_0_14));
  and_gate and_gate_s_CSAwallace_cska24_and_1_14(.a(a[1]), .b(b[14]), .out(s_CSAwallace_cska24_and_1_14));
  and_gate and_gate_s_CSAwallace_cska24_and_2_14(.a(a[2]), .b(b[14]), .out(s_CSAwallace_cska24_and_2_14));
  and_gate and_gate_s_CSAwallace_cska24_and_3_14(.a(a[3]), .b(b[14]), .out(s_CSAwallace_cska24_and_3_14));
  and_gate and_gate_s_CSAwallace_cska24_and_4_14(.a(a[4]), .b(b[14]), .out(s_CSAwallace_cska24_and_4_14));
  and_gate and_gate_s_CSAwallace_cska24_and_5_14(.a(a[5]), .b(b[14]), .out(s_CSAwallace_cska24_and_5_14));
  and_gate and_gate_s_CSAwallace_cska24_and_6_14(.a(a[6]), .b(b[14]), .out(s_CSAwallace_cska24_and_6_14));
  and_gate and_gate_s_CSAwallace_cska24_and_7_14(.a(a[7]), .b(b[14]), .out(s_CSAwallace_cska24_and_7_14));
  and_gate and_gate_s_CSAwallace_cska24_and_8_14(.a(a[8]), .b(b[14]), .out(s_CSAwallace_cska24_and_8_14));
  and_gate and_gate_s_CSAwallace_cska24_and_9_14(.a(a[9]), .b(b[14]), .out(s_CSAwallace_cska24_and_9_14));
  and_gate and_gate_s_CSAwallace_cska24_and_10_14(.a(a[10]), .b(b[14]), .out(s_CSAwallace_cska24_and_10_14));
  and_gate and_gate_s_CSAwallace_cska24_and_11_14(.a(a[11]), .b(b[14]), .out(s_CSAwallace_cska24_and_11_14));
  and_gate and_gate_s_CSAwallace_cska24_and_12_14(.a(a[12]), .b(b[14]), .out(s_CSAwallace_cska24_and_12_14));
  and_gate and_gate_s_CSAwallace_cska24_and_13_14(.a(a[13]), .b(b[14]), .out(s_CSAwallace_cska24_and_13_14));
  and_gate and_gate_s_CSAwallace_cska24_and_14_14(.a(a[14]), .b(b[14]), .out(s_CSAwallace_cska24_and_14_14));
  and_gate and_gate_s_CSAwallace_cska24_and_15_14(.a(a[15]), .b(b[14]), .out(s_CSAwallace_cska24_and_15_14));
  and_gate and_gate_s_CSAwallace_cska24_and_16_14(.a(a[16]), .b(b[14]), .out(s_CSAwallace_cska24_and_16_14));
  and_gate and_gate_s_CSAwallace_cska24_and_17_14(.a(a[17]), .b(b[14]), .out(s_CSAwallace_cska24_and_17_14));
  and_gate and_gate_s_CSAwallace_cska24_and_18_14(.a(a[18]), .b(b[14]), .out(s_CSAwallace_cska24_and_18_14));
  and_gate and_gate_s_CSAwallace_cska24_and_19_14(.a(a[19]), .b(b[14]), .out(s_CSAwallace_cska24_and_19_14));
  and_gate and_gate_s_CSAwallace_cska24_and_20_14(.a(a[20]), .b(b[14]), .out(s_CSAwallace_cska24_and_20_14));
  and_gate and_gate_s_CSAwallace_cska24_and_21_14(.a(a[21]), .b(b[14]), .out(s_CSAwallace_cska24_and_21_14));
  and_gate and_gate_s_CSAwallace_cska24_and_22_14(.a(a[22]), .b(b[14]), .out(s_CSAwallace_cska24_and_22_14));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_14(.a(a[23]), .b(b[14]), .out(s_CSAwallace_cska24_nand_23_14));
  and_gate and_gate_s_CSAwallace_cska24_and_0_15(.a(a[0]), .b(b[15]), .out(s_CSAwallace_cska24_and_0_15));
  and_gate and_gate_s_CSAwallace_cska24_and_1_15(.a(a[1]), .b(b[15]), .out(s_CSAwallace_cska24_and_1_15));
  and_gate and_gate_s_CSAwallace_cska24_and_2_15(.a(a[2]), .b(b[15]), .out(s_CSAwallace_cska24_and_2_15));
  and_gate and_gate_s_CSAwallace_cska24_and_3_15(.a(a[3]), .b(b[15]), .out(s_CSAwallace_cska24_and_3_15));
  and_gate and_gate_s_CSAwallace_cska24_and_4_15(.a(a[4]), .b(b[15]), .out(s_CSAwallace_cska24_and_4_15));
  and_gate and_gate_s_CSAwallace_cska24_and_5_15(.a(a[5]), .b(b[15]), .out(s_CSAwallace_cska24_and_5_15));
  and_gate and_gate_s_CSAwallace_cska24_and_6_15(.a(a[6]), .b(b[15]), .out(s_CSAwallace_cska24_and_6_15));
  and_gate and_gate_s_CSAwallace_cska24_and_7_15(.a(a[7]), .b(b[15]), .out(s_CSAwallace_cska24_and_7_15));
  and_gate and_gate_s_CSAwallace_cska24_and_8_15(.a(a[8]), .b(b[15]), .out(s_CSAwallace_cska24_and_8_15));
  and_gate and_gate_s_CSAwallace_cska24_and_9_15(.a(a[9]), .b(b[15]), .out(s_CSAwallace_cska24_and_9_15));
  and_gate and_gate_s_CSAwallace_cska24_and_10_15(.a(a[10]), .b(b[15]), .out(s_CSAwallace_cska24_and_10_15));
  and_gate and_gate_s_CSAwallace_cska24_and_11_15(.a(a[11]), .b(b[15]), .out(s_CSAwallace_cska24_and_11_15));
  and_gate and_gate_s_CSAwallace_cska24_and_12_15(.a(a[12]), .b(b[15]), .out(s_CSAwallace_cska24_and_12_15));
  and_gate and_gate_s_CSAwallace_cska24_and_13_15(.a(a[13]), .b(b[15]), .out(s_CSAwallace_cska24_and_13_15));
  and_gate and_gate_s_CSAwallace_cska24_and_14_15(.a(a[14]), .b(b[15]), .out(s_CSAwallace_cska24_and_14_15));
  and_gate and_gate_s_CSAwallace_cska24_and_15_15(.a(a[15]), .b(b[15]), .out(s_CSAwallace_cska24_and_15_15));
  and_gate and_gate_s_CSAwallace_cska24_and_16_15(.a(a[16]), .b(b[15]), .out(s_CSAwallace_cska24_and_16_15));
  and_gate and_gate_s_CSAwallace_cska24_and_17_15(.a(a[17]), .b(b[15]), .out(s_CSAwallace_cska24_and_17_15));
  and_gate and_gate_s_CSAwallace_cska24_and_18_15(.a(a[18]), .b(b[15]), .out(s_CSAwallace_cska24_and_18_15));
  and_gate and_gate_s_CSAwallace_cska24_and_19_15(.a(a[19]), .b(b[15]), .out(s_CSAwallace_cska24_and_19_15));
  and_gate and_gate_s_CSAwallace_cska24_and_20_15(.a(a[20]), .b(b[15]), .out(s_CSAwallace_cska24_and_20_15));
  and_gate and_gate_s_CSAwallace_cska24_and_21_15(.a(a[21]), .b(b[15]), .out(s_CSAwallace_cska24_and_21_15));
  and_gate and_gate_s_CSAwallace_cska24_and_22_15(.a(a[22]), .b(b[15]), .out(s_CSAwallace_cska24_and_22_15));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_15(.a(a[23]), .b(b[15]), .out(s_CSAwallace_cska24_nand_23_15));
  and_gate and_gate_s_CSAwallace_cska24_and_0_16(.a(a[0]), .b(b[16]), .out(s_CSAwallace_cska24_and_0_16));
  and_gate and_gate_s_CSAwallace_cska24_and_1_16(.a(a[1]), .b(b[16]), .out(s_CSAwallace_cska24_and_1_16));
  and_gate and_gate_s_CSAwallace_cska24_and_2_16(.a(a[2]), .b(b[16]), .out(s_CSAwallace_cska24_and_2_16));
  and_gate and_gate_s_CSAwallace_cska24_and_3_16(.a(a[3]), .b(b[16]), .out(s_CSAwallace_cska24_and_3_16));
  and_gate and_gate_s_CSAwallace_cska24_and_4_16(.a(a[4]), .b(b[16]), .out(s_CSAwallace_cska24_and_4_16));
  and_gate and_gate_s_CSAwallace_cska24_and_5_16(.a(a[5]), .b(b[16]), .out(s_CSAwallace_cska24_and_5_16));
  and_gate and_gate_s_CSAwallace_cska24_and_6_16(.a(a[6]), .b(b[16]), .out(s_CSAwallace_cska24_and_6_16));
  and_gate and_gate_s_CSAwallace_cska24_and_7_16(.a(a[7]), .b(b[16]), .out(s_CSAwallace_cska24_and_7_16));
  and_gate and_gate_s_CSAwallace_cska24_and_8_16(.a(a[8]), .b(b[16]), .out(s_CSAwallace_cska24_and_8_16));
  and_gate and_gate_s_CSAwallace_cska24_and_9_16(.a(a[9]), .b(b[16]), .out(s_CSAwallace_cska24_and_9_16));
  and_gate and_gate_s_CSAwallace_cska24_and_10_16(.a(a[10]), .b(b[16]), .out(s_CSAwallace_cska24_and_10_16));
  and_gate and_gate_s_CSAwallace_cska24_and_11_16(.a(a[11]), .b(b[16]), .out(s_CSAwallace_cska24_and_11_16));
  and_gate and_gate_s_CSAwallace_cska24_and_12_16(.a(a[12]), .b(b[16]), .out(s_CSAwallace_cska24_and_12_16));
  and_gate and_gate_s_CSAwallace_cska24_and_13_16(.a(a[13]), .b(b[16]), .out(s_CSAwallace_cska24_and_13_16));
  and_gate and_gate_s_CSAwallace_cska24_and_14_16(.a(a[14]), .b(b[16]), .out(s_CSAwallace_cska24_and_14_16));
  and_gate and_gate_s_CSAwallace_cska24_and_15_16(.a(a[15]), .b(b[16]), .out(s_CSAwallace_cska24_and_15_16));
  and_gate and_gate_s_CSAwallace_cska24_and_16_16(.a(a[16]), .b(b[16]), .out(s_CSAwallace_cska24_and_16_16));
  and_gate and_gate_s_CSAwallace_cska24_and_17_16(.a(a[17]), .b(b[16]), .out(s_CSAwallace_cska24_and_17_16));
  and_gate and_gate_s_CSAwallace_cska24_and_18_16(.a(a[18]), .b(b[16]), .out(s_CSAwallace_cska24_and_18_16));
  and_gate and_gate_s_CSAwallace_cska24_and_19_16(.a(a[19]), .b(b[16]), .out(s_CSAwallace_cska24_and_19_16));
  and_gate and_gate_s_CSAwallace_cska24_and_20_16(.a(a[20]), .b(b[16]), .out(s_CSAwallace_cska24_and_20_16));
  and_gate and_gate_s_CSAwallace_cska24_and_21_16(.a(a[21]), .b(b[16]), .out(s_CSAwallace_cska24_and_21_16));
  and_gate and_gate_s_CSAwallace_cska24_and_22_16(.a(a[22]), .b(b[16]), .out(s_CSAwallace_cska24_and_22_16));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_16(.a(a[23]), .b(b[16]), .out(s_CSAwallace_cska24_nand_23_16));
  and_gate and_gate_s_CSAwallace_cska24_and_0_17(.a(a[0]), .b(b[17]), .out(s_CSAwallace_cska24_and_0_17));
  and_gate and_gate_s_CSAwallace_cska24_and_1_17(.a(a[1]), .b(b[17]), .out(s_CSAwallace_cska24_and_1_17));
  and_gate and_gate_s_CSAwallace_cska24_and_2_17(.a(a[2]), .b(b[17]), .out(s_CSAwallace_cska24_and_2_17));
  and_gate and_gate_s_CSAwallace_cska24_and_3_17(.a(a[3]), .b(b[17]), .out(s_CSAwallace_cska24_and_3_17));
  and_gate and_gate_s_CSAwallace_cska24_and_4_17(.a(a[4]), .b(b[17]), .out(s_CSAwallace_cska24_and_4_17));
  and_gate and_gate_s_CSAwallace_cska24_and_5_17(.a(a[5]), .b(b[17]), .out(s_CSAwallace_cska24_and_5_17));
  and_gate and_gate_s_CSAwallace_cska24_and_6_17(.a(a[6]), .b(b[17]), .out(s_CSAwallace_cska24_and_6_17));
  and_gate and_gate_s_CSAwallace_cska24_and_7_17(.a(a[7]), .b(b[17]), .out(s_CSAwallace_cska24_and_7_17));
  and_gate and_gate_s_CSAwallace_cska24_and_8_17(.a(a[8]), .b(b[17]), .out(s_CSAwallace_cska24_and_8_17));
  and_gate and_gate_s_CSAwallace_cska24_and_9_17(.a(a[9]), .b(b[17]), .out(s_CSAwallace_cska24_and_9_17));
  and_gate and_gate_s_CSAwallace_cska24_and_10_17(.a(a[10]), .b(b[17]), .out(s_CSAwallace_cska24_and_10_17));
  and_gate and_gate_s_CSAwallace_cska24_and_11_17(.a(a[11]), .b(b[17]), .out(s_CSAwallace_cska24_and_11_17));
  and_gate and_gate_s_CSAwallace_cska24_and_12_17(.a(a[12]), .b(b[17]), .out(s_CSAwallace_cska24_and_12_17));
  and_gate and_gate_s_CSAwallace_cska24_and_13_17(.a(a[13]), .b(b[17]), .out(s_CSAwallace_cska24_and_13_17));
  and_gate and_gate_s_CSAwallace_cska24_and_14_17(.a(a[14]), .b(b[17]), .out(s_CSAwallace_cska24_and_14_17));
  and_gate and_gate_s_CSAwallace_cska24_and_15_17(.a(a[15]), .b(b[17]), .out(s_CSAwallace_cska24_and_15_17));
  and_gate and_gate_s_CSAwallace_cska24_and_16_17(.a(a[16]), .b(b[17]), .out(s_CSAwallace_cska24_and_16_17));
  and_gate and_gate_s_CSAwallace_cska24_and_17_17(.a(a[17]), .b(b[17]), .out(s_CSAwallace_cska24_and_17_17));
  and_gate and_gate_s_CSAwallace_cska24_and_18_17(.a(a[18]), .b(b[17]), .out(s_CSAwallace_cska24_and_18_17));
  and_gate and_gate_s_CSAwallace_cska24_and_19_17(.a(a[19]), .b(b[17]), .out(s_CSAwallace_cska24_and_19_17));
  and_gate and_gate_s_CSAwallace_cska24_and_20_17(.a(a[20]), .b(b[17]), .out(s_CSAwallace_cska24_and_20_17));
  and_gate and_gate_s_CSAwallace_cska24_and_21_17(.a(a[21]), .b(b[17]), .out(s_CSAwallace_cska24_and_21_17));
  and_gate and_gate_s_CSAwallace_cska24_and_22_17(.a(a[22]), .b(b[17]), .out(s_CSAwallace_cska24_and_22_17));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_17(.a(a[23]), .b(b[17]), .out(s_CSAwallace_cska24_nand_23_17));
  and_gate and_gate_s_CSAwallace_cska24_and_0_18(.a(a[0]), .b(b[18]), .out(s_CSAwallace_cska24_and_0_18));
  and_gate and_gate_s_CSAwallace_cska24_and_1_18(.a(a[1]), .b(b[18]), .out(s_CSAwallace_cska24_and_1_18));
  and_gate and_gate_s_CSAwallace_cska24_and_2_18(.a(a[2]), .b(b[18]), .out(s_CSAwallace_cska24_and_2_18));
  and_gate and_gate_s_CSAwallace_cska24_and_3_18(.a(a[3]), .b(b[18]), .out(s_CSAwallace_cska24_and_3_18));
  and_gate and_gate_s_CSAwallace_cska24_and_4_18(.a(a[4]), .b(b[18]), .out(s_CSAwallace_cska24_and_4_18));
  and_gate and_gate_s_CSAwallace_cska24_and_5_18(.a(a[5]), .b(b[18]), .out(s_CSAwallace_cska24_and_5_18));
  and_gate and_gate_s_CSAwallace_cska24_and_6_18(.a(a[6]), .b(b[18]), .out(s_CSAwallace_cska24_and_6_18));
  and_gate and_gate_s_CSAwallace_cska24_and_7_18(.a(a[7]), .b(b[18]), .out(s_CSAwallace_cska24_and_7_18));
  and_gate and_gate_s_CSAwallace_cska24_and_8_18(.a(a[8]), .b(b[18]), .out(s_CSAwallace_cska24_and_8_18));
  and_gate and_gate_s_CSAwallace_cska24_and_9_18(.a(a[9]), .b(b[18]), .out(s_CSAwallace_cska24_and_9_18));
  and_gate and_gate_s_CSAwallace_cska24_and_10_18(.a(a[10]), .b(b[18]), .out(s_CSAwallace_cska24_and_10_18));
  and_gate and_gate_s_CSAwallace_cska24_and_11_18(.a(a[11]), .b(b[18]), .out(s_CSAwallace_cska24_and_11_18));
  and_gate and_gate_s_CSAwallace_cska24_and_12_18(.a(a[12]), .b(b[18]), .out(s_CSAwallace_cska24_and_12_18));
  and_gate and_gate_s_CSAwallace_cska24_and_13_18(.a(a[13]), .b(b[18]), .out(s_CSAwallace_cska24_and_13_18));
  and_gate and_gate_s_CSAwallace_cska24_and_14_18(.a(a[14]), .b(b[18]), .out(s_CSAwallace_cska24_and_14_18));
  and_gate and_gate_s_CSAwallace_cska24_and_15_18(.a(a[15]), .b(b[18]), .out(s_CSAwallace_cska24_and_15_18));
  and_gate and_gate_s_CSAwallace_cska24_and_16_18(.a(a[16]), .b(b[18]), .out(s_CSAwallace_cska24_and_16_18));
  and_gate and_gate_s_CSAwallace_cska24_and_17_18(.a(a[17]), .b(b[18]), .out(s_CSAwallace_cska24_and_17_18));
  and_gate and_gate_s_CSAwallace_cska24_and_18_18(.a(a[18]), .b(b[18]), .out(s_CSAwallace_cska24_and_18_18));
  and_gate and_gate_s_CSAwallace_cska24_and_19_18(.a(a[19]), .b(b[18]), .out(s_CSAwallace_cska24_and_19_18));
  and_gate and_gate_s_CSAwallace_cska24_and_20_18(.a(a[20]), .b(b[18]), .out(s_CSAwallace_cska24_and_20_18));
  and_gate and_gate_s_CSAwallace_cska24_and_21_18(.a(a[21]), .b(b[18]), .out(s_CSAwallace_cska24_and_21_18));
  and_gate and_gate_s_CSAwallace_cska24_and_22_18(.a(a[22]), .b(b[18]), .out(s_CSAwallace_cska24_and_22_18));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_18(.a(a[23]), .b(b[18]), .out(s_CSAwallace_cska24_nand_23_18));
  and_gate and_gate_s_CSAwallace_cska24_and_0_19(.a(a[0]), .b(b[19]), .out(s_CSAwallace_cska24_and_0_19));
  and_gate and_gate_s_CSAwallace_cska24_and_1_19(.a(a[1]), .b(b[19]), .out(s_CSAwallace_cska24_and_1_19));
  and_gate and_gate_s_CSAwallace_cska24_and_2_19(.a(a[2]), .b(b[19]), .out(s_CSAwallace_cska24_and_2_19));
  and_gate and_gate_s_CSAwallace_cska24_and_3_19(.a(a[3]), .b(b[19]), .out(s_CSAwallace_cska24_and_3_19));
  and_gate and_gate_s_CSAwallace_cska24_and_4_19(.a(a[4]), .b(b[19]), .out(s_CSAwallace_cska24_and_4_19));
  and_gate and_gate_s_CSAwallace_cska24_and_5_19(.a(a[5]), .b(b[19]), .out(s_CSAwallace_cska24_and_5_19));
  and_gate and_gate_s_CSAwallace_cska24_and_6_19(.a(a[6]), .b(b[19]), .out(s_CSAwallace_cska24_and_6_19));
  and_gate and_gate_s_CSAwallace_cska24_and_7_19(.a(a[7]), .b(b[19]), .out(s_CSAwallace_cska24_and_7_19));
  and_gate and_gate_s_CSAwallace_cska24_and_8_19(.a(a[8]), .b(b[19]), .out(s_CSAwallace_cska24_and_8_19));
  and_gate and_gate_s_CSAwallace_cska24_and_9_19(.a(a[9]), .b(b[19]), .out(s_CSAwallace_cska24_and_9_19));
  and_gate and_gate_s_CSAwallace_cska24_and_10_19(.a(a[10]), .b(b[19]), .out(s_CSAwallace_cska24_and_10_19));
  and_gate and_gate_s_CSAwallace_cska24_and_11_19(.a(a[11]), .b(b[19]), .out(s_CSAwallace_cska24_and_11_19));
  and_gate and_gate_s_CSAwallace_cska24_and_12_19(.a(a[12]), .b(b[19]), .out(s_CSAwallace_cska24_and_12_19));
  and_gate and_gate_s_CSAwallace_cska24_and_13_19(.a(a[13]), .b(b[19]), .out(s_CSAwallace_cska24_and_13_19));
  and_gate and_gate_s_CSAwallace_cska24_and_14_19(.a(a[14]), .b(b[19]), .out(s_CSAwallace_cska24_and_14_19));
  and_gate and_gate_s_CSAwallace_cska24_and_15_19(.a(a[15]), .b(b[19]), .out(s_CSAwallace_cska24_and_15_19));
  and_gate and_gate_s_CSAwallace_cska24_and_16_19(.a(a[16]), .b(b[19]), .out(s_CSAwallace_cska24_and_16_19));
  and_gate and_gate_s_CSAwallace_cska24_and_17_19(.a(a[17]), .b(b[19]), .out(s_CSAwallace_cska24_and_17_19));
  and_gate and_gate_s_CSAwallace_cska24_and_18_19(.a(a[18]), .b(b[19]), .out(s_CSAwallace_cska24_and_18_19));
  and_gate and_gate_s_CSAwallace_cska24_and_19_19(.a(a[19]), .b(b[19]), .out(s_CSAwallace_cska24_and_19_19));
  and_gate and_gate_s_CSAwallace_cska24_and_20_19(.a(a[20]), .b(b[19]), .out(s_CSAwallace_cska24_and_20_19));
  and_gate and_gate_s_CSAwallace_cska24_and_21_19(.a(a[21]), .b(b[19]), .out(s_CSAwallace_cska24_and_21_19));
  and_gate and_gate_s_CSAwallace_cska24_and_22_19(.a(a[22]), .b(b[19]), .out(s_CSAwallace_cska24_and_22_19));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_19(.a(a[23]), .b(b[19]), .out(s_CSAwallace_cska24_nand_23_19));
  and_gate and_gate_s_CSAwallace_cska24_and_0_20(.a(a[0]), .b(b[20]), .out(s_CSAwallace_cska24_and_0_20));
  and_gate and_gate_s_CSAwallace_cska24_and_1_20(.a(a[1]), .b(b[20]), .out(s_CSAwallace_cska24_and_1_20));
  and_gate and_gate_s_CSAwallace_cska24_and_2_20(.a(a[2]), .b(b[20]), .out(s_CSAwallace_cska24_and_2_20));
  and_gate and_gate_s_CSAwallace_cska24_and_3_20(.a(a[3]), .b(b[20]), .out(s_CSAwallace_cska24_and_3_20));
  and_gate and_gate_s_CSAwallace_cska24_and_4_20(.a(a[4]), .b(b[20]), .out(s_CSAwallace_cska24_and_4_20));
  and_gate and_gate_s_CSAwallace_cska24_and_5_20(.a(a[5]), .b(b[20]), .out(s_CSAwallace_cska24_and_5_20));
  and_gate and_gate_s_CSAwallace_cska24_and_6_20(.a(a[6]), .b(b[20]), .out(s_CSAwallace_cska24_and_6_20));
  and_gate and_gate_s_CSAwallace_cska24_and_7_20(.a(a[7]), .b(b[20]), .out(s_CSAwallace_cska24_and_7_20));
  and_gate and_gate_s_CSAwallace_cska24_and_8_20(.a(a[8]), .b(b[20]), .out(s_CSAwallace_cska24_and_8_20));
  and_gate and_gate_s_CSAwallace_cska24_and_9_20(.a(a[9]), .b(b[20]), .out(s_CSAwallace_cska24_and_9_20));
  and_gate and_gate_s_CSAwallace_cska24_and_10_20(.a(a[10]), .b(b[20]), .out(s_CSAwallace_cska24_and_10_20));
  and_gate and_gate_s_CSAwallace_cska24_and_11_20(.a(a[11]), .b(b[20]), .out(s_CSAwallace_cska24_and_11_20));
  and_gate and_gate_s_CSAwallace_cska24_and_12_20(.a(a[12]), .b(b[20]), .out(s_CSAwallace_cska24_and_12_20));
  and_gate and_gate_s_CSAwallace_cska24_and_13_20(.a(a[13]), .b(b[20]), .out(s_CSAwallace_cska24_and_13_20));
  and_gate and_gate_s_CSAwallace_cska24_and_14_20(.a(a[14]), .b(b[20]), .out(s_CSAwallace_cska24_and_14_20));
  and_gate and_gate_s_CSAwallace_cska24_and_15_20(.a(a[15]), .b(b[20]), .out(s_CSAwallace_cska24_and_15_20));
  and_gate and_gate_s_CSAwallace_cska24_and_16_20(.a(a[16]), .b(b[20]), .out(s_CSAwallace_cska24_and_16_20));
  and_gate and_gate_s_CSAwallace_cska24_and_17_20(.a(a[17]), .b(b[20]), .out(s_CSAwallace_cska24_and_17_20));
  and_gate and_gate_s_CSAwallace_cska24_and_18_20(.a(a[18]), .b(b[20]), .out(s_CSAwallace_cska24_and_18_20));
  and_gate and_gate_s_CSAwallace_cska24_and_19_20(.a(a[19]), .b(b[20]), .out(s_CSAwallace_cska24_and_19_20));
  and_gate and_gate_s_CSAwallace_cska24_and_20_20(.a(a[20]), .b(b[20]), .out(s_CSAwallace_cska24_and_20_20));
  and_gate and_gate_s_CSAwallace_cska24_and_21_20(.a(a[21]), .b(b[20]), .out(s_CSAwallace_cska24_and_21_20));
  and_gate and_gate_s_CSAwallace_cska24_and_22_20(.a(a[22]), .b(b[20]), .out(s_CSAwallace_cska24_and_22_20));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_20(.a(a[23]), .b(b[20]), .out(s_CSAwallace_cska24_nand_23_20));
  and_gate and_gate_s_CSAwallace_cska24_and_0_21(.a(a[0]), .b(b[21]), .out(s_CSAwallace_cska24_and_0_21));
  and_gate and_gate_s_CSAwallace_cska24_and_1_21(.a(a[1]), .b(b[21]), .out(s_CSAwallace_cska24_and_1_21));
  and_gate and_gate_s_CSAwallace_cska24_and_2_21(.a(a[2]), .b(b[21]), .out(s_CSAwallace_cska24_and_2_21));
  and_gate and_gate_s_CSAwallace_cska24_and_3_21(.a(a[3]), .b(b[21]), .out(s_CSAwallace_cska24_and_3_21));
  and_gate and_gate_s_CSAwallace_cska24_and_4_21(.a(a[4]), .b(b[21]), .out(s_CSAwallace_cska24_and_4_21));
  and_gate and_gate_s_CSAwallace_cska24_and_5_21(.a(a[5]), .b(b[21]), .out(s_CSAwallace_cska24_and_5_21));
  and_gate and_gate_s_CSAwallace_cska24_and_6_21(.a(a[6]), .b(b[21]), .out(s_CSAwallace_cska24_and_6_21));
  and_gate and_gate_s_CSAwallace_cska24_and_7_21(.a(a[7]), .b(b[21]), .out(s_CSAwallace_cska24_and_7_21));
  and_gate and_gate_s_CSAwallace_cska24_and_8_21(.a(a[8]), .b(b[21]), .out(s_CSAwallace_cska24_and_8_21));
  and_gate and_gate_s_CSAwallace_cska24_and_9_21(.a(a[9]), .b(b[21]), .out(s_CSAwallace_cska24_and_9_21));
  and_gate and_gate_s_CSAwallace_cska24_and_10_21(.a(a[10]), .b(b[21]), .out(s_CSAwallace_cska24_and_10_21));
  and_gate and_gate_s_CSAwallace_cska24_and_11_21(.a(a[11]), .b(b[21]), .out(s_CSAwallace_cska24_and_11_21));
  and_gate and_gate_s_CSAwallace_cska24_and_12_21(.a(a[12]), .b(b[21]), .out(s_CSAwallace_cska24_and_12_21));
  and_gate and_gate_s_CSAwallace_cska24_and_13_21(.a(a[13]), .b(b[21]), .out(s_CSAwallace_cska24_and_13_21));
  and_gate and_gate_s_CSAwallace_cska24_and_14_21(.a(a[14]), .b(b[21]), .out(s_CSAwallace_cska24_and_14_21));
  and_gate and_gate_s_CSAwallace_cska24_and_15_21(.a(a[15]), .b(b[21]), .out(s_CSAwallace_cska24_and_15_21));
  and_gate and_gate_s_CSAwallace_cska24_and_16_21(.a(a[16]), .b(b[21]), .out(s_CSAwallace_cska24_and_16_21));
  and_gate and_gate_s_CSAwallace_cska24_and_17_21(.a(a[17]), .b(b[21]), .out(s_CSAwallace_cska24_and_17_21));
  and_gate and_gate_s_CSAwallace_cska24_and_18_21(.a(a[18]), .b(b[21]), .out(s_CSAwallace_cska24_and_18_21));
  and_gate and_gate_s_CSAwallace_cska24_and_19_21(.a(a[19]), .b(b[21]), .out(s_CSAwallace_cska24_and_19_21));
  and_gate and_gate_s_CSAwallace_cska24_and_20_21(.a(a[20]), .b(b[21]), .out(s_CSAwallace_cska24_and_20_21));
  and_gate and_gate_s_CSAwallace_cska24_and_21_21(.a(a[21]), .b(b[21]), .out(s_CSAwallace_cska24_and_21_21));
  and_gate and_gate_s_CSAwallace_cska24_and_22_21(.a(a[22]), .b(b[21]), .out(s_CSAwallace_cska24_and_22_21));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_21(.a(a[23]), .b(b[21]), .out(s_CSAwallace_cska24_nand_23_21));
  and_gate and_gate_s_CSAwallace_cska24_and_0_22(.a(a[0]), .b(b[22]), .out(s_CSAwallace_cska24_and_0_22));
  and_gate and_gate_s_CSAwallace_cska24_and_1_22(.a(a[1]), .b(b[22]), .out(s_CSAwallace_cska24_and_1_22));
  and_gate and_gate_s_CSAwallace_cska24_and_2_22(.a(a[2]), .b(b[22]), .out(s_CSAwallace_cska24_and_2_22));
  and_gate and_gate_s_CSAwallace_cska24_and_3_22(.a(a[3]), .b(b[22]), .out(s_CSAwallace_cska24_and_3_22));
  and_gate and_gate_s_CSAwallace_cska24_and_4_22(.a(a[4]), .b(b[22]), .out(s_CSAwallace_cska24_and_4_22));
  and_gate and_gate_s_CSAwallace_cska24_and_5_22(.a(a[5]), .b(b[22]), .out(s_CSAwallace_cska24_and_5_22));
  and_gate and_gate_s_CSAwallace_cska24_and_6_22(.a(a[6]), .b(b[22]), .out(s_CSAwallace_cska24_and_6_22));
  and_gate and_gate_s_CSAwallace_cska24_and_7_22(.a(a[7]), .b(b[22]), .out(s_CSAwallace_cska24_and_7_22));
  and_gate and_gate_s_CSAwallace_cska24_and_8_22(.a(a[8]), .b(b[22]), .out(s_CSAwallace_cska24_and_8_22));
  and_gate and_gate_s_CSAwallace_cska24_and_9_22(.a(a[9]), .b(b[22]), .out(s_CSAwallace_cska24_and_9_22));
  and_gate and_gate_s_CSAwallace_cska24_and_10_22(.a(a[10]), .b(b[22]), .out(s_CSAwallace_cska24_and_10_22));
  and_gate and_gate_s_CSAwallace_cska24_and_11_22(.a(a[11]), .b(b[22]), .out(s_CSAwallace_cska24_and_11_22));
  and_gate and_gate_s_CSAwallace_cska24_and_12_22(.a(a[12]), .b(b[22]), .out(s_CSAwallace_cska24_and_12_22));
  and_gate and_gate_s_CSAwallace_cska24_and_13_22(.a(a[13]), .b(b[22]), .out(s_CSAwallace_cska24_and_13_22));
  and_gate and_gate_s_CSAwallace_cska24_and_14_22(.a(a[14]), .b(b[22]), .out(s_CSAwallace_cska24_and_14_22));
  and_gate and_gate_s_CSAwallace_cska24_and_15_22(.a(a[15]), .b(b[22]), .out(s_CSAwallace_cska24_and_15_22));
  and_gate and_gate_s_CSAwallace_cska24_and_16_22(.a(a[16]), .b(b[22]), .out(s_CSAwallace_cska24_and_16_22));
  and_gate and_gate_s_CSAwallace_cska24_and_17_22(.a(a[17]), .b(b[22]), .out(s_CSAwallace_cska24_and_17_22));
  and_gate and_gate_s_CSAwallace_cska24_and_18_22(.a(a[18]), .b(b[22]), .out(s_CSAwallace_cska24_and_18_22));
  and_gate and_gate_s_CSAwallace_cska24_and_19_22(.a(a[19]), .b(b[22]), .out(s_CSAwallace_cska24_and_19_22));
  and_gate and_gate_s_CSAwallace_cska24_and_20_22(.a(a[20]), .b(b[22]), .out(s_CSAwallace_cska24_and_20_22));
  and_gate and_gate_s_CSAwallace_cska24_and_21_22(.a(a[21]), .b(b[22]), .out(s_CSAwallace_cska24_and_21_22));
  and_gate and_gate_s_CSAwallace_cska24_and_22_22(.a(a[22]), .b(b[22]), .out(s_CSAwallace_cska24_and_22_22));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_23_22(.a(a[23]), .b(b[22]), .out(s_CSAwallace_cska24_nand_23_22));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_0_23(.a(a[0]), .b(b[23]), .out(s_CSAwallace_cska24_nand_0_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_1_23(.a(a[1]), .b(b[23]), .out(s_CSAwallace_cska24_nand_1_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_2_23(.a(a[2]), .b(b[23]), .out(s_CSAwallace_cska24_nand_2_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_3_23(.a(a[3]), .b(b[23]), .out(s_CSAwallace_cska24_nand_3_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_4_23(.a(a[4]), .b(b[23]), .out(s_CSAwallace_cska24_nand_4_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_5_23(.a(a[5]), .b(b[23]), .out(s_CSAwallace_cska24_nand_5_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_6_23(.a(a[6]), .b(b[23]), .out(s_CSAwallace_cska24_nand_6_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_7_23(.a(a[7]), .b(b[23]), .out(s_CSAwallace_cska24_nand_7_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_8_23(.a(a[8]), .b(b[23]), .out(s_CSAwallace_cska24_nand_8_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_9_23(.a(a[9]), .b(b[23]), .out(s_CSAwallace_cska24_nand_9_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_10_23(.a(a[10]), .b(b[23]), .out(s_CSAwallace_cska24_nand_10_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_11_23(.a(a[11]), .b(b[23]), .out(s_CSAwallace_cska24_nand_11_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_12_23(.a(a[12]), .b(b[23]), .out(s_CSAwallace_cska24_nand_12_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_13_23(.a(a[13]), .b(b[23]), .out(s_CSAwallace_cska24_nand_13_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_14_23(.a(a[14]), .b(b[23]), .out(s_CSAwallace_cska24_nand_14_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_15_23(.a(a[15]), .b(b[23]), .out(s_CSAwallace_cska24_nand_15_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_16_23(.a(a[16]), .b(b[23]), .out(s_CSAwallace_cska24_nand_16_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_17_23(.a(a[17]), .b(b[23]), .out(s_CSAwallace_cska24_nand_17_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_18_23(.a(a[18]), .b(b[23]), .out(s_CSAwallace_cska24_nand_18_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_19_23(.a(a[19]), .b(b[23]), .out(s_CSAwallace_cska24_nand_19_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_20_23(.a(a[20]), .b(b[23]), .out(s_CSAwallace_cska24_nand_20_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_21_23(.a(a[21]), .b(b[23]), .out(s_CSAwallace_cska24_nand_21_23));
  nand_gate nand_gate_s_CSAwallace_cska24_nand_22_23(.a(a[22]), .b(b[23]), .out(s_CSAwallace_cska24_nand_22_23));
  and_gate and_gate_s_CSAwallace_cska24_and_23_23(.a(a[23]), .b(b[23]), .out(s_CSAwallace_cska24_and_23_23));
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[0] = s_CSAwallace_cska24_and_0_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[1] = s_CSAwallace_cska24_and_1_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[2] = s_CSAwallace_cska24_and_2_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[3] = s_CSAwallace_cska24_and_3_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[4] = s_CSAwallace_cska24_and_4_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[5] = s_CSAwallace_cska24_and_5_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[6] = s_CSAwallace_cska24_and_6_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[7] = s_CSAwallace_cska24_and_7_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[8] = s_CSAwallace_cska24_and_8_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[9] = s_CSAwallace_cska24_and_9_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[10] = s_CSAwallace_cska24_and_10_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[11] = s_CSAwallace_cska24_and_11_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[12] = s_CSAwallace_cska24_and_12_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[13] = s_CSAwallace_cska24_and_13_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[14] = s_CSAwallace_cska24_and_14_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[15] = s_CSAwallace_cska24_and_15_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[16] = s_CSAwallace_cska24_and_16_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[17] = s_CSAwallace_cska24_and_17_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[18] = s_CSAwallace_cska24_and_18_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[19] = s_CSAwallace_cska24_and_19_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[20] = s_CSAwallace_cska24_and_20_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[21] = s_CSAwallace_cska24_and_21_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[22] = s_CSAwallace_cska24_and_22_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[23] = s_CSAwallace_cska24_nand_23_0[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[24] = 1'b1;
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row0[25] = 1'b1;
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[0] = 1'b0;
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[1] = s_CSAwallace_cska24_and_0_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[2] = s_CSAwallace_cska24_and_1_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[3] = s_CSAwallace_cska24_and_2_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[4] = s_CSAwallace_cska24_and_3_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[5] = s_CSAwallace_cska24_and_4_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[6] = s_CSAwallace_cska24_and_5_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[7] = s_CSAwallace_cska24_and_6_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[8] = s_CSAwallace_cska24_and_7_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[9] = s_CSAwallace_cska24_and_8_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[10] = s_CSAwallace_cska24_and_9_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[11] = s_CSAwallace_cska24_and_10_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[12] = s_CSAwallace_cska24_and_11_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[13] = s_CSAwallace_cska24_and_12_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[14] = s_CSAwallace_cska24_and_13_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[15] = s_CSAwallace_cska24_and_14_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[16] = s_CSAwallace_cska24_and_15_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[17] = s_CSAwallace_cska24_and_16_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[18] = s_CSAwallace_cska24_and_17_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[19] = s_CSAwallace_cska24_and_18_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[20] = s_CSAwallace_cska24_and_19_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[21] = s_CSAwallace_cska24_and_20_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[22] = s_CSAwallace_cska24_and_21_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[23] = s_CSAwallace_cska24_and_22_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[24] = s_CSAwallace_cska24_nand_23_1[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row1[25] = 1'b1;
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[0] = 1'b0;
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[1] = 1'b0;
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[2] = s_CSAwallace_cska24_and_0_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[3] = s_CSAwallace_cska24_and_1_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[4] = s_CSAwallace_cska24_and_2_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[5] = s_CSAwallace_cska24_and_3_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[6] = s_CSAwallace_cska24_and_4_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[7] = s_CSAwallace_cska24_and_5_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[8] = s_CSAwallace_cska24_and_6_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[9] = s_CSAwallace_cska24_and_7_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[10] = s_CSAwallace_cska24_and_8_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[11] = s_CSAwallace_cska24_and_9_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[12] = s_CSAwallace_cska24_and_10_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[13] = s_CSAwallace_cska24_and_11_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[14] = s_CSAwallace_cska24_and_12_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[15] = s_CSAwallace_cska24_and_13_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[16] = s_CSAwallace_cska24_and_14_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[17] = s_CSAwallace_cska24_and_15_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[18] = s_CSAwallace_cska24_and_16_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[19] = s_CSAwallace_cska24_and_17_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[20] = s_CSAwallace_cska24_and_18_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[21] = s_CSAwallace_cska24_and_19_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[22] = s_CSAwallace_cska24_and_20_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[23] = s_CSAwallace_cska24_and_21_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[24] = s_CSAwallace_cska24_and_22_2[0];
  assign s_CSAwallace_cska24_csa0_csa_component_pp_row2[25] = s_CSAwallace_cska24_nand_23_2[0];
  csa_component26 csa_component26_s_CSAwallace_cska24_csa0_csa_component_out(.a(s_CSAwallace_cska24_csa0_csa_component_pp_row0), .b(s_CSAwallace_cska24_csa0_csa_component_pp_row1), .c(s_CSAwallace_cska24_csa0_csa_component_pp_row2), .csa_component26_out(s_CSAwallace_cska24_csa0_csa_component_out));
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[0] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[1] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[2] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[3] = s_CSAwallace_cska24_and_0_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[4] = s_CSAwallace_cska24_and_1_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[5] = s_CSAwallace_cska24_and_2_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[6] = s_CSAwallace_cska24_and_3_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[7] = s_CSAwallace_cska24_and_4_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[8] = s_CSAwallace_cska24_and_5_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[9] = s_CSAwallace_cska24_and_6_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[10] = s_CSAwallace_cska24_and_7_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[11] = s_CSAwallace_cska24_and_8_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[12] = s_CSAwallace_cska24_and_9_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[13] = s_CSAwallace_cska24_and_10_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[14] = s_CSAwallace_cska24_and_11_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[15] = s_CSAwallace_cska24_and_12_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[16] = s_CSAwallace_cska24_and_13_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[17] = s_CSAwallace_cska24_and_14_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[18] = s_CSAwallace_cska24_and_15_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[19] = s_CSAwallace_cska24_and_16_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[20] = s_CSAwallace_cska24_and_17_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[21] = s_CSAwallace_cska24_and_18_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[22] = s_CSAwallace_cska24_and_19_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[23] = s_CSAwallace_cska24_and_20_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[24] = s_CSAwallace_cska24_and_21_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[25] = s_CSAwallace_cska24_and_22_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[26] = s_CSAwallace_cska24_nand_23_3[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[27] = 1'b1;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row3[28] = 1'b1;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[0] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[1] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[2] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[3] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[4] = s_CSAwallace_cska24_and_0_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[5] = s_CSAwallace_cska24_and_1_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[6] = s_CSAwallace_cska24_and_2_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[7] = s_CSAwallace_cska24_and_3_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[8] = s_CSAwallace_cska24_and_4_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[9] = s_CSAwallace_cska24_and_5_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[10] = s_CSAwallace_cska24_and_6_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[11] = s_CSAwallace_cska24_and_7_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[12] = s_CSAwallace_cska24_and_8_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[13] = s_CSAwallace_cska24_and_9_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[14] = s_CSAwallace_cska24_and_10_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[15] = s_CSAwallace_cska24_and_11_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[16] = s_CSAwallace_cska24_and_12_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[17] = s_CSAwallace_cska24_and_13_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[18] = s_CSAwallace_cska24_and_14_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[19] = s_CSAwallace_cska24_and_15_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[20] = s_CSAwallace_cska24_and_16_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[21] = s_CSAwallace_cska24_and_17_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[22] = s_CSAwallace_cska24_and_18_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[23] = s_CSAwallace_cska24_and_19_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[24] = s_CSAwallace_cska24_and_20_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[25] = s_CSAwallace_cska24_and_21_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[26] = s_CSAwallace_cska24_and_22_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[27] = s_CSAwallace_cska24_nand_23_4[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row4[28] = 1'b1;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[0] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[1] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[2] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[3] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[4] = 1'b0;
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[5] = s_CSAwallace_cska24_and_0_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[6] = s_CSAwallace_cska24_and_1_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[7] = s_CSAwallace_cska24_and_2_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[8] = s_CSAwallace_cska24_and_3_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[9] = s_CSAwallace_cska24_and_4_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[10] = s_CSAwallace_cska24_and_5_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[11] = s_CSAwallace_cska24_and_6_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[12] = s_CSAwallace_cska24_and_7_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[13] = s_CSAwallace_cska24_and_8_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[14] = s_CSAwallace_cska24_and_9_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[15] = s_CSAwallace_cska24_and_10_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[16] = s_CSAwallace_cska24_and_11_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[17] = s_CSAwallace_cska24_and_12_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[18] = s_CSAwallace_cska24_and_13_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[19] = s_CSAwallace_cska24_and_14_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[20] = s_CSAwallace_cska24_and_15_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[21] = s_CSAwallace_cska24_and_16_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[22] = s_CSAwallace_cska24_and_17_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[23] = s_CSAwallace_cska24_and_18_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[24] = s_CSAwallace_cska24_and_19_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[25] = s_CSAwallace_cska24_and_20_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[26] = s_CSAwallace_cska24_and_21_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[27] = s_CSAwallace_cska24_and_22_5[0];
  assign s_CSAwallace_cska24_csa1_csa_component_pp_row5[28] = s_CSAwallace_cska24_nand_23_5[0];
  csa_component29 csa_component29_s_CSAwallace_cska24_csa1_csa_component_out(.a(s_CSAwallace_cska24_csa1_csa_component_pp_row3), .b(s_CSAwallace_cska24_csa1_csa_component_pp_row4), .c(s_CSAwallace_cska24_csa1_csa_component_pp_row5), .csa_component29_out(s_CSAwallace_cska24_csa1_csa_component_out));
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[0] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[1] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[2] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[3] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[4] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[5] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[6] = s_CSAwallace_cska24_and_0_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[7] = s_CSAwallace_cska24_and_1_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[8] = s_CSAwallace_cska24_and_2_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[9] = s_CSAwallace_cska24_and_3_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[10] = s_CSAwallace_cska24_and_4_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[11] = s_CSAwallace_cska24_and_5_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[12] = s_CSAwallace_cska24_and_6_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[13] = s_CSAwallace_cska24_and_7_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[14] = s_CSAwallace_cska24_and_8_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[15] = s_CSAwallace_cska24_and_9_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[16] = s_CSAwallace_cska24_and_10_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[17] = s_CSAwallace_cska24_and_11_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[18] = s_CSAwallace_cska24_and_12_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[19] = s_CSAwallace_cska24_and_13_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[20] = s_CSAwallace_cska24_and_14_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[21] = s_CSAwallace_cska24_and_15_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[22] = s_CSAwallace_cska24_and_16_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[23] = s_CSAwallace_cska24_and_17_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[24] = s_CSAwallace_cska24_and_18_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[25] = s_CSAwallace_cska24_and_19_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[26] = s_CSAwallace_cska24_and_20_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[27] = s_CSAwallace_cska24_and_21_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[28] = s_CSAwallace_cska24_and_22_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[29] = s_CSAwallace_cska24_nand_23_6[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[30] = 1'b1;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row6[31] = 1'b1;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[0] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[1] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[2] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[3] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[4] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[5] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[6] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[7] = s_CSAwallace_cska24_and_0_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[8] = s_CSAwallace_cska24_and_1_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[9] = s_CSAwallace_cska24_and_2_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[10] = s_CSAwallace_cska24_and_3_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[11] = s_CSAwallace_cska24_and_4_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[12] = s_CSAwallace_cska24_and_5_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[13] = s_CSAwallace_cska24_and_6_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[14] = s_CSAwallace_cska24_and_7_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[15] = s_CSAwallace_cska24_and_8_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[16] = s_CSAwallace_cska24_and_9_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[17] = s_CSAwallace_cska24_and_10_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[18] = s_CSAwallace_cska24_and_11_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[19] = s_CSAwallace_cska24_and_12_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[20] = s_CSAwallace_cska24_and_13_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[21] = s_CSAwallace_cska24_and_14_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[22] = s_CSAwallace_cska24_and_15_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[23] = s_CSAwallace_cska24_and_16_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[24] = s_CSAwallace_cska24_and_17_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[25] = s_CSAwallace_cska24_and_18_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[26] = s_CSAwallace_cska24_and_19_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[27] = s_CSAwallace_cska24_and_20_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[28] = s_CSAwallace_cska24_and_21_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[29] = s_CSAwallace_cska24_and_22_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[30] = s_CSAwallace_cska24_nand_23_7[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row7[31] = 1'b1;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[0] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[1] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[2] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[3] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[4] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[5] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[6] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[7] = 1'b0;
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[8] = s_CSAwallace_cska24_and_0_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[9] = s_CSAwallace_cska24_and_1_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[10] = s_CSAwallace_cska24_and_2_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[11] = s_CSAwallace_cska24_and_3_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[12] = s_CSAwallace_cska24_and_4_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[13] = s_CSAwallace_cska24_and_5_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[14] = s_CSAwallace_cska24_and_6_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[15] = s_CSAwallace_cska24_and_7_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[16] = s_CSAwallace_cska24_and_8_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[17] = s_CSAwallace_cska24_and_9_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[18] = s_CSAwallace_cska24_and_10_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[19] = s_CSAwallace_cska24_and_11_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[20] = s_CSAwallace_cska24_and_12_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[21] = s_CSAwallace_cska24_and_13_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[22] = s_CSAwallace_cska24_and_14_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[23] = s_CSAwallace_cska24_and_15_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[24] = s_CSAwallace_cska24_and_16_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[25] = s_CSAwallace_cska24_and_17_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[26] = s_CSAwallace_cska24_and_18_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[27] = s_CSAwallace_cska24_and_19_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[28] = s_CSAwallace_cska24_and_20_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[29] = s_CSAwallace_cska24_and_21_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[30] = s_CSAwallace_cska24_and_22_8[0];
  assign s_CSAwallace_cska24_csa2_csa_component_pp_row8[31] = s_CSAwallace_cska24_nand_23_8[0];
  csa_component32 csa_component32_s_CSAwallace_cska24_csa2_csa_component_out(.a(s_CSAwallace_cska24_csa2_csa_component_pp_row6), .b(s_CSAwallace_cska24_csa2_csa_component_pp_row7), .c(s_CSAwallace_cska24_csa2_csa_component_pp_row8), .csa_component32_out(s_CSAwallace_cska24_csa2_csa_component_out));
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[0] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[1] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[2] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[3] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[4] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[5] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[6] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[7] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[8] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[9] = s_CSAwallace_cska24_and_0_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[10] = s_CSAwallace_cska24_and_1_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[11] = s_CSAwallace_cska24_and_2_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[12] = s_CSAwallace_cska24_and_3_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[13] = s_CSAwallace_cska24_and_4_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[14] = s_CSAwallace_cska24_and_5_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[15] = s_CSAwallace_cska24_and_6_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[16] = s_CSAwallace_cska24_and_7_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[17] = s_CSAwallace_cska24_and_8_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[18] = s_CSAwallace_cska24_and_9_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[19] = s_CSAwallace_cska24_and_10_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[20] = s_CSAwallace_cska24_and_11_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[21] = s_CSAwallace_cska24_and_12_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[22] = s_CSAwallace_cska24_and_13_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[23] = s_CSAwallace_cska24_and_14_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[24] = s_CSAwallace_cska24_and_15_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[25] = s_CSAwallace_cska24_and_16_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[26] = s_CSAwallace_cska24_and_17_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[27] = s_CSAwallace_cska24_and_18_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[28] = s_CSAwallace_cska24_and_19_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[29] = s_CSAwallace_cska24_and_20_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[30] = s_CSAwallace_cska24_and_21_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[31] = s_CSAwallace_cska24_and_22_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[32] = s_CSAwallace_cska24_nand_23_9[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[33] = 1'b1;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row9[34] = 1'b1;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[0] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[1] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[2] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[3] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[4] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[5] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[6] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[7] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[8] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[9] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[10] = s_CSAwallace_cska24_and_0_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[11] = s_CSAwallace_cska24_and_1_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[12] = s_CSAwallace_cska24_and_2_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[13] = s_CSAwallace_cska24_and_3_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[14] = s_CSAwallace_cska24_and_4_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[15] = s_CSAwallace_cska24_and_5_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[16] = s_CSAwallace_cska24_and_6_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[17] = s_CSAwallace_cska24_and_7_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[18] = s_CSAwallace_cska24_and_8_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[19] = s_CSAwallace_cska24_and_9_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[20] = s_CSAwallace_cska24_and_10_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[21] = s_CSAwallace_cska24_and_11_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[22] = s_CSAwallace_cska24_and_12_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[23] = s_CSAwallace_cska24_and_13_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[24] = s_CSAwallace_cska24_and_14_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[25] = s_CSAwallace_cska24_and_15_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[26] = s_CSAwallace_cska24_and_16_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[27] = s_CSAwallace_cska24_and_17_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[28] = s_CSAwallace_cska24_and_18_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[29] = s_CSAwallace_cska24_and_19_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[30] = s_CSAwallace_cska24_and_20_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[31] = s_CSAwallace_cska24_and_21_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[32] = s_CSAwallace_cska24_and_22_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[33] = s_CSAwallace_cska24_nand_23_10[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row10[34] = 1'b1;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[0] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[1] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[2] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[3] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[4] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[5] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[6] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[7] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[8] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[9] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[10] = 1'b0;
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[11] = s_CSAwallace_cska24_and_0_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[12] = s_CSAwallace_cska24_and_1_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[13] = s_CSAwallace_cska24_and_2_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[14] = s_CSAwallace_cska24_and_3_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[15] = s_CSAwallace_cska24_and_4_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[16] = s_CSAwallace_cska24_and_5_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[17] = s_CSAwallace_cska24_and_6_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[18] = s_CSAwallace_cska24_and_7_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[19] = s_CSAwallace_cska24_and_8_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[20] = s_CSAwallace_cska24_and_9_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[21] = s_CSAwallace_cska24_and_10_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[22] = s_CSAwallace_cska24_and_11_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[23] = s_CSAwallace_cska24_and_12_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[24] = s_CSAwallace_cska24_and_13_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[25] = s_CSAwallace_cska24_and_14_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[26] = s_CSAwallace_cska24_and_15_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[27] = s_CSAwallace_cska24_and_16_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[28] = s_CSAwallace_cska24_and_17_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[29] = s_CSAwallace_cska24_and_18_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[30] = s_CSAwallace_cska24_and_19_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[31] = s_CSAwallace_cska24_and_20_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[32] = s_CSAwallace_cska24_and_21_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[33] = s_CSAwallace_cska24_and_22_11[0];
  assign s_CSAwallace_cska24_csa3_csa_component_pp_row11[34] = s_CSAwallace_cska24_nand_23_11[0];
  csa_component35 csa_component35_s_CSAwallace_cska24_csa3_csa_component_out(.a(s_CSAwallace_cska24_csa3_csa_component_pp_row9), .b(s_CSAwallace_cska24_csa3_csa_component_pp_row10), .c(s_CSAwallace_cska24_csa3_csa_component_pp_row11), .csa_component35_out(s_CSAwallace_cska24_csa3_csa_component_out));
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[0] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[1] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[2] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[3] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[4] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[5] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[6] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[7] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[8] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[9] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[10] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[11] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[12] = s_CSAwallace_cska24_and_0_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[13] = s_CSAwallace_cska24_and_1_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[14] = s_CSAwallace_cska24_and_2_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[15] = s_CSAwallace_cska24_and_3_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[16] = s_CSAwallace_cska24_and_4_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[17] = s_CSAwallace_cska24_and_5_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[18] = s_CSAwallace_cska24_and_6_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[19] = s_CSAwallace_cska24_and_7_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[20] = s_CSAwallace_cska24_and_8_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[21] = s_CSAwallace_cska24_and_9_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[22] = s_CSAwallace_cska24_and_10_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[23] = s_CSAwallace_cska24_and_11_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[24] = s_CSAwallace_cska24_and_12_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[25] = s_CSAwallace_cska24_and_13_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[26] = s_CSAwallace_cska24_and_14_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[27] = s_CSAwallace_cska24_and_15_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[28] = s_CSAwallace_cska24_and_16_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[29] = s_CSAwallace_cska24_and_17_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[30] = s_CSAwallace_cska24_and_18_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[31] = s_CSAwallace_cska24_and_19_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[32] = s_CSAwallace_cska24_and_20_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[33] = s_CSAwallace_cska24_and_21_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[34] = s_CSAwallace_cska24_and_22_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[35] = s_CSAwallace_cska24_nand_23_12[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[36] = 1'b1;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row12[37] = 1'b1;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[0] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[1] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[2] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[3] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[4] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[5] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[6] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[7] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[8] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[9] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[10] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[11] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[12] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[13] = s_CSAwallace_cska24_and_0_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[14] = s_CSAwallace_cska24_and_1_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[15] = s_CSAwallace_cska24_and_2_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[16] = s_CSAwallace_cska24_and_3_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[17] = s_CSAwallace_cska24_and_4_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[18] = s_CSAwallace_cska24_and_5_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[19] = s_CSAwallace_cska24_and_6_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[20] = s_CSAwallace_cska24_and_7_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[21] = s_CSAwallace_cska24_and_8_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[22] = s_CSAwallace_cska24_and_9_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[23] = s_CSAwallace_cska24_and_10_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[24] = s_CSAwallace_cska24_and_11_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[25] = s_CSAwallace_cska24_and_12_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[26] = s_CSAwallace_cska24_and_13_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[27] = s_CSAwallace_cska24_and_14_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[28] = s_CSAwallace_cska24_and_15_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[29] = s_CSAwallace_cska24_and_16_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[30] = s_CSAwallace_cska24_and_17_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[31] = s_CSAwallace_cska24_and_18_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[32] = s_CSAwallace_cska24_and_19_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[33] = s_CSAwallace_cska24_and_20_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[34] = s_CSAwallace_cska24_and_21_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[35] = s_CSAwallace_cska24_and_22_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[36] = s_CSAwallace_cska24_nand_23_13[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row13[37] = 1'b1;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[0] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[1] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[2] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[3] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[4] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[5] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[6] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[7] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[8] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[9] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[10] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[11] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[12] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[13] = 1'b0;
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[14] = s_CSAwallace_cska24_and_0_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[15] = s_CSAwallace_cska24_and_1_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[16] = s_CSAwallace_cska24_and_2_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[17] = s_CSAwallace_cska24_and_3_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[18] = s_CSAwallace_cska24_and_4_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[19] = s_CSAwallace_cska24_and_5_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[20] = s_CSAwallace_cska24_and_6_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[21] = s_CSAwallace_cska24_and_7_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[22] = s_CSAwallace_cska24_and_8_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[23] = s_CSAwallace_cska24_and_9_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[24] = s_CSAwallace_cska24_and_10_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[25] = s_CSAwallace_cska24_and_11_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[26] = s_CSAwallace_cska24_and_12_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[27] = s_CSAwallace_cska24_and_13_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[28] = s_CSAwallace_cska24_and_14_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[29] = s_CSAwallace_cska24_and_15_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[30] = s_CSAwallace_cska24_and_16_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[31] = s_CSAwallace_cska24_and_17_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[32] = s_CSAwallace_cska24_and_18_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[33] = s_CSAwallace_cska24_and_19_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[34] = s_CSAwallace_cska24_and_20_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[35] = s_CSAwallace_cska24_and_21_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[36] = s_CSAwallace_cska24_and_22_14[0];
  assign s_CSAwallace_cska24_csa4_csa_component_pp_row14[37] = s_CSAwallace_cska24_nand_23_14[0];
  csa_component38 csa_component38_s_CSAwallace_cska24_csa4_csa_component_out(.a(s_CSAwallace_cska24_csa4_csa_component_pp_row12), .b(s_CSAwallace_cska24_csa4_csa_component_pp_row13), .c(s_CSAwallace_cska24_csa4_csa_component_pp_row14), .csa_component38_out(s_CSAwallace_cska24_csa4_csa_component_out));
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[0] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[1] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[2] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[3] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[4] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[5] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[6] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[7] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[8] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[9] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[10] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[11] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[12] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[13] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[14] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[15] = s_CSAwallace_cska24_and_0_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[16] = s_CSAwallace_cska24_and_1_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[17] = s_CSAwallace_cska24_and_2_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[18] = s_CSAwallace_cska24_and_3_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[19] = s_CSAwallace_cska24_and_4_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[20] = s_CSAwallace_cska24_and_5_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[21] = s_CSAwallace_cska24_and_6_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[22] = s_CSAwallace_cska24_and_7_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[23] = s_CSAwallace_cska24_and_8_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[24] = s_CSAwallace_cska24_and_9_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[25] = s_CSAwallace_cska24_and_10_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[26] = s_CSAwallace_cska24_and_11_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[27] = s_CSAwallace_cska24_and_12_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[28] = s_CSAwallace_cska24_and_13_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[29] = s_CSAwallace_cska24_and_14_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[30] = s_CSAwallace_cska24_and_15_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[31] = s_CSAwallace_cska24_and_16_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[32] = s_CSAwallace_cska24_and_17_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[33] = s_CSAwallace_cska24_and_18_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[34] = s_CSAwallace_cska24_and_19_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[35] = s_CSAwallace_cska24_and_20_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[36] = s_CSAwallace_cska24_and_21_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[37] = s_CSAwallace_cska24_and_22_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[38] = s_CSAwallace_cska24_nand_23_15[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[39] = 1'b1;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row15[40] = 1'b1;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[0] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[1] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[2] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[3] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[4] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[5] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[6] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[7] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[8] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[9] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[10] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[11] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[12] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[13] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[14] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[15] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[16] = s_CSAwallace_cska24_and_0_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[17] = s_CSAwallace_cska24_and_1_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[18] = s_CSAwallace_cska24_and_2_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[19] = s_CSAwallace_cska24_and_3_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[20] = s_CSAwallace_cska24_and_4_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[21] = s_CSAwallace_cska24_and_5_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[22] = s_CSAwallace_cska24_and_6_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[23] = s_CSAwallace_cska24_and_7_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[24] = s_CSAwallace_cska24_and_8_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[25] = s_CSAwallace_cska24_and_9_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[26] = s_CSAwallace_cska24_and_10_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[27] = s_CSAwallace_cska24_and_11_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[28] = s_CSAwallace_cska24_and_12_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[29] = s_CSAwallace_cska24_and_13_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[30] = s_CSAwallace_cska24_and_14_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[31] = s_CSAwallace_cska24_and_15_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[32] = s_CSAwallace_cska24_and_16_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[33] = s_CSAwallace_cska24_and_17_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[34] = s_CSAwallace_cska24_and_18_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[35] = s_CSAwallace_cska24_and_19_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[36] = s_CSAwallace_cska24_and_20_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[37] = s_CSAwallace_cska24_and_21_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[38] = s_CSAwallace_cska24_and_22_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[39] = s_CSAwallace_cska24_nand_23_16[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row16[40] = 1'b1;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[0] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[1] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[2] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[3] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[4] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[5] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[6] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[7] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[8] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[9] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[10] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[11] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[12] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[13] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[14] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[15] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[16] = 1'b0;
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[17] = s_CSAwallace_cska24_and_0_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[18] = s_CSAwallace_cska24_and_1_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[19] = s_CSAwallace_cska24_and_2_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[20] = s_CSAwallace_cska24_and_3_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[21] = s_CSAwallace_cska24_and_4_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[22] = s_CSAwallace_cska24_and_5_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[23] = s_CSAwallace_cska24_and_6_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[24] = s_CSAwallace_cska24_and_7_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[25] = s_CSAwallace_cska24_and_8_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[26] = s_CSAwallace_cska24_and_9_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[27] = s_CSAwallace_cska24_and_10_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[28] = s_CSAwallace_cska24_and_11_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[29] = s_CSAwallace_cska24_and_12_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[30] = s_CSAwallace_cska24_and_13_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[31] = s_CSAwallace_cska24_and_14_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[32] = s_CSAwallace_cska24_and_15_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[33] = s_CSAwallace_cska24_and_16_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[34] = s_CSAwallace_cska24_and_17_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[35] = s_CSAwallace_cska24_and_18_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[36] = s_CSAwallace_cska24_and_19_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[37] = s_CSAwallace_cska24_and_20_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[38] = s_CSAwallace_cska24_and_21_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[39] = s_CSAwallace_cska24_and_22_17[0];
  assign s_CSAwallace_cska24_csa5_csa_component_pp_row17[40] = s_CSAwallace_cska24_nand_23_17[0];
  csa_component41 csa_component41_s_CSAwallace_cska24_csa5_csa_component_out(.a(s_CSAwallace_cska24_csa5_csa_component_pp_row15), .b(s_CSAwallace_cska24_csa5_csa_component_pp_row16), .c(s_CSAwallace_cska24_csa5_csa_component_pp_row17), .csa_component41_out(s_CSAwallace_cska24_csa5_csa_component_out));
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[0] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[1] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[2] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[3] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[4] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[5] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[6] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[7] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[8] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[9] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[10] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[11] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[12] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[13] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[14] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[15] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[16] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[17] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[18] = s_CSAwallace_cska24_and_0_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[19] = s_CSAwallace_cska24_and_1_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[20] = s_CSAwallace_cska24_and_2_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[21] = s_CSAwallace_cska24_and_3_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[22] = s_CSAwallace_cska24_and_4_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[23] = s_CSAwallace_cska24_and_5_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[24] = s_CSAwallace_cska24_and_6_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[25] = s_CSAwallace_cska24_and_7_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[26] = s_CSAwallace_cska24_and_8_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[27] = s_CSAwallace_cska24_and_9_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[28] = s_CSAwallace_cska24_and_10_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[29] = s_CSAwallace_cska24_and_11_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[30] = s_CSAwallace_cska24_and_12_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[31] = s_CSAwallace_cska24_and_13_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[32] = s_CSAwallace_cska24_and_14_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[33] = s_CSAwallace_cska24_and_15_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[34] = s_CSAwallace_cska24_and_16_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[35] = s_CSAwallace_cska24_and_17_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[36] = s_CSAwallace_cska24_and_18_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[37] = s_CSAwallace_cska24_and_19_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[38] = s_CSAwallace_cska24_and_20_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[39] = s_CSAwallace_cska24_and_21_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[40] = s_CSAwallace_cska24_and_22_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[41] = s_CSAwallace_cska24_nand_23_18[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[42] = 1'b1;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row18[43] = 1'b1;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[0] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[1] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[2] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[3] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[4] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[5] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[6] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[7] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[8] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[9] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[10] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[11] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[12] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[13] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[14] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[15] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[16] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[17] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[18] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[19] = s_CSAwallace_cska24_and_0_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[20] = s_CSAwallace_cska24_and_1_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[21] = s_CSAwallace_cska24_and_2_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[22] = s_CSAwallace_cska24_and_3_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[23] = s_CSAwallace_cska24_and_4_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[24] = s_CSAwallace_cska24_and_5_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[25] = s_CSAwallace_cska24_and_6_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[26] = s_CSAwallace_cska24_and_7_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[27] = s_CSAwallace_cska24_and_8_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[28] = s_CSAwallace_cska24_and_9_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[29] = s_CSAwallace_cska24_and_10_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[30] = s_CSAwallace_cska24_and_11_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[31] = s_CSAwallace_cska24_and_12_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[32] = s_CSAwallace_cska24_and_13_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[33] = s_CSAwallace_cska24_and_14_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[34] = s_CSAwallace_cska24_and_15_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[35] = s_CSAwallace_cska24_and_16_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[36] = s_CSAwallace_cska24_and_17_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[37] = s_CSAwallace_cska24_and_18_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[38] = s_CSAwallace_cska24_and_19_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[39] = s_CSAwallace_cska24_and_20_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[40] = s_CSAwallace_cska24_and_21_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[41] = s_CSAwallace_cska24_and_22_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[42] = s_CSAwallace_cska24_nand_23_19[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row19[43] = 1'b1;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[0] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[1] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[2] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[3] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[4] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[5] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[6] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[7] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[8] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[9] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[10] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[11] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[12] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[13] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[14] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[15] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[16] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[17] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[18] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[19] = 1'b0;
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[20] = s_CSAwallace_cska24_and_0_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[21] = s_CSAwallace_cska24_and_1_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[22] = s_CSAwallace_cska24_and_2_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[23] = s_CSAwallace_cska24_and_3_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[24] = s_CSAwallace_cska24_and_4_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[25] = s_CSAwallace_cska24_and_5_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[26] = s_CSAwallace_cska24_and_6_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[27] = s_CSAwallace_cska24_and_7_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[28] = s_CSAwallace_cska24_and_8_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[29] = s_CSAwallace_cska24_and_9_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[30] = s_CSAwallace_cska24_and_10_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[31] = s_CSAwallace_cska24_and_11_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[32] = s_CSAwallace_cska24_and_12_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[33] = s_CSAwallace_cska24_and_13_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[34] = s_CSAwallace_cska24_and_14_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[35] = s_CSAwallace_cska24_and_15_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[36] = s_CSAwallace_cska24_and_16_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[37] = s_CSAwallace_cska24_and_17_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[38] = s_CSAwallace_cska24_and_18_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[39] = s_CSAwallace_cska24_and_19_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[40] = s_CSAwallace_cska24_and_20_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[41] = s_CSAwallace_cska24_and_21_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[42] = s_CSAwallace_cska24_and_22_20[0];
  assign s_CSAwallace_cska24_csa6_csa_component_pp_row20[43] = s_CSAwallace_cska24_nand_23_20[0];
  csa_component44 csa_component44_s_CSAwallace_cska24_csa6_csa_component_out(.a(s_CSAwallace_cska24_csa6_csa_component_pp_row18), .b(s_CSAwallace_cska24_csa6_csa_component_pp_row19), .c(s_CSAwallace_cska24_csa6_csa_component_pp_row20), .csa_component44_out(s_CSAwallace_cska24_csa6_csa_component_out));
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[0] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[1] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[2] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[3] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[4] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[5] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[6] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[7] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[8] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[9] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[10] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[11] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[12] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[13] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[14] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[15] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[16] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[17] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[18] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[19] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[20] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[21] = s_CSAwallace_cska24_and_0_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[22] = s_CSAwallace_cska24_and_1_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[23] = s_CSAwallace_cska24_and_2_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[24] = s_CSAwallace_cska24_and_3_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[25] = s_CSAwallace_cska24_and_4_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[26] = s_CSAwallace_cska24_and_5_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[27] = s_CSAwallace_cska24_and_6_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[28] = s_CSAwallace_cska24_and_7_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[29] = s_CSAwallace_cska24_and_8_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[30] = s_CSAwallace_cska24_and_9_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[31] = s_CSAwallace_cska24_and_10_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[32] = s_CSAwallace_cska24_and_11_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[33] = s_CSAwallace_cska24_and_12_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[34] = s_CSAwallace_cska24_and_13_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[35] = s_CSAwallace_cska24_and_14_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[36] = s_CSAwallace_cska24_and_15_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[37] = s_CSAwallace_cska24_and_16_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[38] = s_CSAwallace_cska24_and_17_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[39] = s_CSAwallace_cska24_and_18_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[40] = s_CSAwallace_cska24_and_19_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[41] = s_CSAwallace_cska24_and_20_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[42] = s_CSAwallace_cska24_and_21_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[43] = s_CSAwallace_cska24_and_22_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[44] = s_CSAwallace_cska24_nand_23_21[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[45] = 1'b1;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row21[46] = 1'b1;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[0] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[1] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[2] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[3] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[4] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[5] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[6] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[7] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[8] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[9] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[10] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[11] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[12] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[13] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[14] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[15] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[16] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[17] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[18] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[19] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[20] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[21] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[22] = s_CSAwallace_cska24_and_0_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[23] = s_CSAwallace_cska24_and_1_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[24] = s_CSAwallace_cska24_and_2_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[25] = s_CSAwallace_cska24_and_3_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[26] = s_CSAwallace_cska24_and_4_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[27] = s_CSAwallace_cska24_and_5_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[28] = s_CSAwallace_cska24_and_6_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[29] = s_CSAwallace_cska24_and_7_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[30] = s_CSAwallace_cska24_and_8_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[31] = s_CSAwallace_cska24_and_9_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[32] = s_CSAwallace_cska24_and_10_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[33] = s_CSAwallace_cska24_and_11_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[34] = s_CSAwallace_cska24_and_12_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[35] = s_CSAwallace_cska24_and_13_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[36] = s_CSAwallace_cska24_and_14_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[37] = s_CSAwallace_cska24_and_15_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[38] = s_CSAwallace_cska24_and_16_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[39] = s_CSAwallace_cska24_and_17_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[40] = s_CSAwallace_cska24_and_18_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[41] = s_CSAwallace_cska24_and_19_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[42] = s_CSAwallace_cska24_and_20_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[43] = s_CSAwallace_cska24_and_21_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[44] = s_CSAwallace_cska24_and_22_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[45] = s_CSAwallace_cska24_nand_23_22[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row22[46] = 1'b1;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[0] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[1] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[2] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[3] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[4] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[5] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[6] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[7] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[8] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[9] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[10] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[11] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[12] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[13] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[14] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[15] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[16] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[17] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[18] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[19] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[20] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[21] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[22] = 1'b0;
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[23] = s_CSAwallace_cska24_nand_0_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[24] = s_CSAwallace_cska24_nand_1_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[25] = s_CSAwallace_cska24_nand_2_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[26] = s_CSAwallace_cska24_nand_3_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[27] = s_CSAwallace_cska24_nand_4_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[28] = s_CSAwallace_cska24_nand_5_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[29] = s_CSAwallace_cska24_nand_6_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[30] = s_CSAwallace_cska24_nand_7_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[31] = s_CSAwallace_cska24_nand_8_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[32] = s_CSAwallace_cska24_nand_9_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[33] = s_CSAwallace_cska24_nand_10_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[34] = s_CSAwallace_cska24_nand_11_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[35] = s_CSAwallace_cska24_nand_12_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[36] = s_CSAwallace_cska24_nand_13_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[37] = s_CSAwallace_cska24_nand_14_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[38] = s_CSAwallace_cska24_nand_15_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[39] = s_CSAwallace_cska24_nand_16_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[40] = s_CSAwallace_cska24_nand_17_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[41] = s_CSAwallace_cska24_nand_18_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[42] = s_CSAwallace_cska24_nand_19_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[43] = s_CSAwallace_cska24_nand_20_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[44] = s_CSAwallace_cska24_nand_21_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[45] = s_CSAwallace_cska24_nand_22_23[0];
  assign s_CSAwallace_cska24_csa7_csa_component_pp_row23[46] = s_CSAwallace_cska24_and_23_23[0];
  csa_component47 csa_component47_s_CSAwallace_cska24_csa7_csa_component_out(.a(s_CSAwallace_cska24_csa7_csa_component_pp_row21), .b(s_CSAwallace_cska24_csa7_csa_component_pp_row22), .c(s_CSAwallace_cska24_csa7_csa_component_pp_row23), .csa_component47_out(s_CSAwallace_cska24_csa7_csa_component_out));
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[0] = s_CSAwallace_cska24_csa0_csa_component_out[0];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[1] = s_CSAwallace_cska24_csa0_csa_component_out[1];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[2] = s_CSAwallace_cska24_csa0_csa_component_out[2];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[3] = s_CSAwallace_cska24_csa0_csa_component_out[3];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[4] = s_CSAwallace_cska24_csa0_csa_component_out[4];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[5] = s_CSAwallace_cska24_csa0_csa_component_out[5];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[6] = s_CSAwallace_cska24_csa0_csa_component_out[6];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[7] = s_CSAwallace_cska24_csa0_csa_component_out[7];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[8] = s_CSAwallace_cska24_csa0_csa_component_out[8];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[9] = s_CSAwallace_cska24_csa0_csa_component_out[9];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[10] = s_CSAwallace_cska24_csa0_csa_component_out[10];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[11] = s_CSAwallace_cska24_csa0_csa_component_out[11];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[12] = s_CSAwallace_cska24_csa0_csa_component_out[12];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[13] = s_CSAwallace_cska24_csa0_csa_component_out[13];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[14] = s_CSAwallace_cska24_csa0_csa_component_out[14];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[15] = s_CSAwallace_cska24_csa0_csa_component_out[15];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[16] = s_CSAwallace_cska24_csa0_csa_component_out[16];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[17] = s_CSAwallace_cska24_csa0_csa_component_out[17];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[18] = s_CSAwallace_cska24_csa0_csa_component_out[18];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[19] = s_CSAwallace_cska24_csa0_csa_component_out[19];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[20] = s_CSAwallace_cska24_csa0_csa_component_out[20];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[21] = s_CSAwallace_cska24_csa0_csa_component_out[21];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[22] = s_CSAwallace_cska24_csa0_csa_component_out[22];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[23] = s_CSAwallace_cska24_csa0_csa_component_out[23];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[24] = s_CSAwallace_cska24_csa0_csa_component_out[24];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[25] = s_CSAwallace_cska24_csa0_csa_component_out[25];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[26] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[27] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[28] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1[29] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[0] = 1'b0;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[1] = 1'b0;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[2] = s_CSAwallace_cska24_csa0_csa_component_out[29];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[3] = s_CSAwallace_cska24_csa0_csa_component_out[30];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[4] = s_CSAwallace_cska24_csa0_csa_component_out[31];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[5] = s_CSAwallace_cska24_csa0_csa_component_out[32];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[6] = s_CSAwallace_cska24_csa0_csa_component_out[33];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[7] = s_CSAwallace_cska24_csa0_csa_component_out[34];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[8] = s_CSAwallace_cska24_csa0_csa_component_out[35];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[9] = s_CSAwallace_cska24_csa0_csa_component_out[36];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[10] = s_CSAwallace_cska24_csa0_csa_component_out[37];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[11] = s_CSAwallace_cska24_csa0_csa_component_out[38];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[12] = s_CSAwallace_cska24_csa0_csa_component_out[39];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[13] = s_CSAwallace_cska24_csa0_csa_component_out[40];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[14] = s_CSAwallace_cska24_csa0_csa_component_out[41];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[15] = s_CSAwallace_cska24_csa0_csa_component_out[42];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[16] = s_CSAwallace_cska24_csa0_csa_component_out[43];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[17] = s_CSAwallace_cska24_csa0_csa_component_out[44];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[18] = s_CSAwallace_cska24_csa0_csa_component_out[45];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[19] = s_CSAwallace_cska24_csa0_csa_component_out[46];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[20] = s_CSAwallace_cska24_csa0_csa_component_out[47];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[21] = s_CSAwallace_cska24_csa0_csa_component_out[48];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[22] = s_CSAwallace_cska24_csa0_csa_component_out[49];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[23] = s_CSAwallace_cska24_csa0_csa_component_out[50];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[24] = s_CSAwallace_cska24_csa0_csa_component_out[51];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[25] = s_CSAwallace_cska24_csa0_csa_component_out[52];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[26] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[27] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[28] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1[29] = 1'b1;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[0] = 1'b0;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[1] = 1'b0;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[2] = 1'b0;
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[3] = s_CSAwallace_cska24_csa1_csa_component_out[3];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[4] = s_CSAwallace_cska24_csa1_csa_component_out[4];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[5] = s_CSAwallace_cska24_csa1_csa_component_out[5];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[6] = s_CSAwallace_cska24_csa1_csa_component_out[6];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[7] = s_CSAwallace_cska24_csa1_csa_component_out[7];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[8] = s_CSAwallace_cska24_csa1_csa_component_out[8];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[9] = s_CSAwallace_cska24_csa1_csa_component_out[9];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[10] = s_CSAwallace_cska24_csa1_csa_component_out[10];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[11] = s_CSAwallace_cska24_csa1_csa_component_out[11];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[12] = s_CSAwallace_cska24_csa1_csa_component_out[12];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[13] = s_CSAwallace_cska24_csa1_csa_component_out[13];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[14] = s_CSAwallace_cska24_csa1_csa_component_out[14];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[15] = s_CSAwallace_cska24_csa1_csa_component_out[15];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[16] = s_CSAwallace_cska24_csa1_csa_component_out[16];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[17] = s_CSAwallace_cska24_csa1_csa_component_out[17];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[18] = s_CSAwallace_cska24_csa1_csa_component_out[18];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[19] = s_CSAwallace_cska24_csa1_csa_component_out[19];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[20] = s_CSAwallace_cska24_csa1_csa_component_out[20];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[21] = s_CSAwallace_cska24_csa1_csa_component_out[21];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[22] = s_CSAwallace_cska24_csa1_csa_component_out[22];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[23] = s_CSAwallace_cska24_csa1_csa_component_out[23];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[24] = s_CSAwallace_cska24_csa1_csa_component_out[24];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[25] = s_CSAwallace_cska24_csa1_csa_component_out[25];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[26] = s_CSAwallace_cska24_csa1_csa_component_out[26];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[27] = s_CSAwallace_cska24_csa1_csa_component_out[27];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[28] = s_CSAwallace_cska24_csa1_csa_component_out[28];
  assign s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2[29] = 1'b1;
  csa_component30 csa_component30_s_CSAwallace_cska24_csa8_csa_component_out(.a(s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s1), .b(s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_c1), .c(s_CSAwallace_cska24_csa8_csa_component_s_CSAwallace_cska24_csa_s2), .csa_component30_out(s_CSAwallace_cska24_csa8_csa_component_out));
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[0] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[1] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[2] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[3] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[4] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[5] = s_CSAwallace_cska24_csa1_csa_component_out[35];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[6] = s_CSAwallace_cska24_csa1_csa_component_out[36];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[7] = s_CSAwallace_cska24_csa1_csa_component_out[37];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[8] = s_CSAwallace_cska24_csa1_csa_component_out[38];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[9] = s_CSAwallace_cska24_csa1_csa_component_out[39];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[10] = s_CSAwallace_cska24_csa1_csa_component_out[40];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[11] = s_CSAwallace_cska24_csa1_csa_component_out[41];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[12] = s_CSAwallace_cska24_csa1_csa_component_out[42];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[13] = s_CSAwallace_cska24_csa1_csa_component_out[43];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[14] = s_CSAwallace_cska24_csa1_csa_component_out[44];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[15] = s_CSAwallace_cska24_csa1_csa_component_out[45];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[16] = s_CSAwallace_cska24_csa1_csa_component_out[46];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[17] = s_CSAwallace_cska24_csa1_csa_component_out[47];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[18] = s_CSAwallace_cska24_csa1_csa_component_out[48];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[19] = s_CSAwallace_cska24_csa1_csa_component_out[49];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[20] = s_CSAwallace_cska24_csa1_csa_component_out[50];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[21] = s_CSAwallace_cska24_csa1_csa_component_out[51];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[22] = s_CSAwallace_cska24_csa1_csa_component_out[52];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[23] = s_CSAwallace_cska24_csa1_csa_component_out[53];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[24] = s_CSAwallace_cska24_csa1_csa_component_out[54];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[25] = s_CSAwallace_cska24_csa1_csa_component_out[55];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[26] = s_CSAwallace_cska24_csa1_csa_component_out[56];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[27] = s_CSAwallace_cska24_csa1_csa_component_out[57];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[28] = s_CSAwallace_cska24_csa1_csa_component_out[58];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[29] = 1'b1;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[30] = 1'b1;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[31] = 1'b1;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2[32] = 1'b1;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[0] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[1] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[2] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[3] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[4] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[5] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[6] = s_CSAwallace_cska24_csa2_csa_component_out[6];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[7] = s_CSAwallace_cska24_csa2_csa_component_out[7];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[8] = s_CSAwallace_cska24_csa2_csa_component_out[8];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[9] = s_CSAwallace_cska24_csa2_csa_component_out[9];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[10] = s_CSAwallace_cska24_csa2_csa_component_out[10];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[11] = s_CSAwallace_cska24_csa2_csa_component_out[11];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[12] = s_CSAwallace_cska24_csa2_csa_component_out[12];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[13] = s_CSAwallace_cska24_csa2_csa_component_out[13];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[14] = s_CSAwallace_cska24_csa2_csa_component_out[14];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[15] = s_CSAwallace_cska24_csa2_csa_component_out[15];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[16] = s_CSAwallace_cska24_csa2_csa_component_out[16];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[17] = s_CSAwallace_cska24_csa2_csa_component_out[17];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[18] = s_CSAwallace_cska24_csa2_csa_component_out[18];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[19] = s_CSAwallace_cska24_csa2_csa_component_out[19];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[20] = s_CSAwallace_cska24_csa2_csa_component_out[20];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[21] = s_CSAwallace_cska24_csa2_csa_component_out[21];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[22] = s_CSAwallace_cska24_csa2_csa_component_out[22];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[23] = s_CSAwallace_cska24_csa2_csa_component_out[23];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[24] = s_CSAwallace_cska24_csa2_csa_component_out[24];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[25] = s_CSAwallace_cska24_csa2_csa_component_out[25];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[26] = s_CSAwallace_cska24_csa2_csa_component_out[26];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[27] = s_CSAwallace_cska24_csa2_csa_component_out[27];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[28] = s_CSAwallace_cska24_csa2_csa_component_out[28];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[29] = s_CSAwallace_cska24_csa2_csa_component_out[29];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[30] = s_CSAwallace_cska24_csa2_csa_component_out[30];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[31] = s_CSAwallace_cska24_csa2_csa_component_out[31];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3[32] = 1'b1;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[0] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[1] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[2] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[3] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[4] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[5] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[6] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[7] = 1'b0;
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[8] = s_CSAwallace_cska24_csa2_csa_component_out[41];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[9] = s_CSAwallace_cska24_csa2_csa_component_out[42];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[10] = s_CSAwallace_cska24_csa2_csa_component_out[43];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[11] = s_CSAwallace_cska24_csa2_csa_component_out[44];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[12] = s_CSAwallace_cska24_csa2_csa_component_out[45];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[13] = s_CSAwallace_cska24_csa2_csa_component_out[46];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[14] = s_CSAwallace_cska24_csa2_csa_component_out[47];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[15] = s_CSAwallace_cska24_csa2_csa_component_out[48];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[16] = s_CSAwallace_cska24_csa2_csa_component_out[49];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[17] = s_CSAwallace_cska24_csa2_csa_component_out[50];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[18] = s_CSAwallace_cska24_csa2_csa_component_out[51];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[19] = s_CSAwallace_cska24_csa2_csa_component_out[52];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[20] = s_CSAwallace_cska24_csa2_csa_component_out[53];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[21] = s_CSAwallace_cska24_csa2_csa_component_out[54];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[22] = s_CSAwallace_cska24_csa2_csa_component_out[55];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[23] = s_CSAwallace_cska24_csa2_csa_component_out[56];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[24] = s_CSAwallace_cska24_csa2_csa_component_out[57];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[25] = s_CSAwallace_cska24_csa2_csa_component_out[58];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[26] = s_CSAwallace_cska24_csa2_csa_component_out[59];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[27] = s_CSAwallace_cska24_csa2_csa_component_out[60];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[28] = s_CSAwallace_cska24_csa2_csa_component_out[61];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[29] = s_CSAwallace_cska24_csa2_csa_component_out[62];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[30] = s_CSAwallace_cska24_csa2_csa_component_out[63];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[31] = s_CSAwallace_cska24_csa2_csa_component_out[64];
  assign s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3[32] = 1'b1;
  csa_component33 csa_component33_s_CSAwallace_cska24_csa9_csa_component_out(.a(s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c2), .b(s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_s3), .c(s_CSAwallace_cska24_csa9_csa_component_s_CSAwallace_cska24_csa_c3), .csa_component33_out(s_CSAwallace_cska24_csa9_csa_component_out));
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[0] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[1] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[2] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[3] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[4] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[5] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[6] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[7] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[8] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[9] = s_CSAwallace_cska24_csa3_csa_component_out[9];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[10] = s_CSAwallace_cska24_csa3_csa_component_out[10];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[11] = s_CSAwallace_cska24_csa3_csa_component_out[11];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[12] = s_CSAwallace_cska24_csa3_csa_component_out[12];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[13] = s_CSAwallace_cska24_csa3_csa_component_out[13];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[14] = s_CSAwallace_cska24_csa3_csa_component_out[14];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[15] = s_CSAwallace_cska24_csa3_csa_component_out[15];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[16] = s_CSAwallace_cska24_csa3_csa_component_out[16];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[17] = s_CSAwallace_cska24_csa3_csa_component_out[17];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[18] = s_CSAwallace_cska24_csa3_csa_component_out[18];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[19] = s_CSAwallace_cska24_csa3_csa_component_out[19];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[20] = s_CSAwallace_cska24_csa3_csa_component_out[20];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[21] = s_CSAwallace_cska24_csa3_csa_component_out[21];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[22] = s_CSAwallace_cska24_csa3_csa_component_out[22];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[23] = s_CSAwallace_cska24_csa3_csa_component_out[23];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[24] = s_CSAwallace_cska24_csa3_csa_component_out[24];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[25] = s_CSAwallace_cska24_csa3_csa_component_out[25];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[26] = s_CSAwallace_cska24_csa3_csa_component_out[26];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[27] = s_CSAwallace_cska24_csa3_csa_component_out[27];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[28] = s_CSAwallace_cska24_csa3_csa_component_out[28];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[29] = s_CSAwallace_cska24_csa3_csa_component_out[29];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[30] = s_CSAwallace_cska24_csa3_csa_component_out[30];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[31] = s_CSAwallace_cska24_csa3_csa_component_out[31];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[32] = s_CSAwallace_cska24_csa3_csa_component_out[32];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[33] = s_CSAwallace_cska24_csa3_csa_component_out[33];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[34] = s_CSAwallace_cska24_csa3_csa_component_out[34];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[35] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[36] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[37] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4[38] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[0] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[1] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[2] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[3] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[4] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[5] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[6] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[7] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[8] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[9] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[10] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[11] = s_CSAwallace_cska24_csa3_csa_component_out[47];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[12] = s_CSAwallace_cska24_csa3_csa_component_out[48];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[13] = s_CSAwallace_cska24_csa3_csa_component_out[49];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[14] = s_CSAwallace_cska24_csa3_csa_component_out[50];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[15] = s_CSAwallace_cska24_csa3_csa_component_out[51];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[16] = s_CSAwallace_cska24_csa3_csa_component_out[52];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[17] = s_CSAwallace_cska24_csa3_csa_component_out[53];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[18] = s_CSAwallace_cska24_csa3_csa_component_out[54];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[19] = s_CSAwallace_cska24_csa3_csa_component_out[55];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[20] = s_CSAwallace_cska24_csa3_csa_component_out[56];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[21] = s_CSAwallace_cska24_csa3_csa_component_out[57];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[22] = s_CSAwallace_cska24_csa3_csa_component_out[58];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[23] = s_CSAwallace_cska24_csa3_csa_component_out[59];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[24] = s_CSAwallace_cska24_csa3_csa_component_out[60];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[25] = s_CSAwallace_cska24_csa3_csa_component_out[61];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[26] = s_CSAwallace_cska24_csa3_csa_component_out[62];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[27] = s_CSAwallace_cska24_csa3_csa_component_out[63];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[28] = s_CSAwallace_cska24_csa3_csa_component_out[64];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[29] = s_CSAwallace_cska24_csa3_csa_component_out[65];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[30] = s_CSAwallace_cska24_csa3_csa_component_out[66];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[31] = s_CSAwallace_cska24_csa3_csa_component_out[67];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[32] = s_CSAwallace_cska24_csa3_csa_component_out[68];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[33] = s_CSAwallace_cska24_csa3_csa_component_out[69];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[34] = s_CSAwallace_cska24_csa3_csa_component_out[70];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[35] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[36] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[37] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4[38] = 1'b1;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[0] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[1] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[2] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[3] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[4] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[5] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[6] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[7] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[8] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[9] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[10] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[11] = 1'b0;
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[12] = s_CSAwallace_cska24_csa4_csa_component_out[12];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[13] = s_CSAwallace_cska24_csa4_csa_component_out[13];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[14] = s_CSAwallace_cska24_csa4_csa_component_out[14];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[15] = s_CSAwallace_cska24_csa4_csa_component_out[15];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[16] = s_CSAwallace_cska24_csa4_csa_component_out[16];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[17] = s_CSAwallace_cska24_csa4_csa_component_out[17];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[18] = s_CSAwallace_cska24_csa4_csa_component_out[18];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[19] = s_CSAwallace_cska24_csa4_csa_component_out[19];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[20] = s_CSAwallace_cska24_csa4_csa_component_out[20];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[21] = s_CSAwallace_cska24_csa4_csa_component_out[21];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[22] = s_CSAwallace_cska24_csa4_csa_component_out[22];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[23] = s_CSAwallace_cska24_csa4_csa_component_out[23];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[24] = s_CSAwallace_cska24_csa4_csa_component_out[24];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[25] = s_CSAwallace_cska24_csa4_csa_component_out[25];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[26] = s_CSAwallace_cska24_csa4_csa_component_out[26];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[27] = s_CSAwallace_cska24_csa4_csa_component_out[27];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[28] = s_CSAwallace_cska24_csa4_csa_component_out[28];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[29] = s_CSAwallace_cska24_csa4_csa_component_out[29];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[30] = s_CSAwallace_cska24_csa4_csa_component_out[30];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[31] = s_CSAwallace_cska24_csa4_csa_component_out[31];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[32] = s_CSAwallace_cska24_csa4_csa_component_out[32];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[33] = s_CSAwallace_cska24_csa4_csa_component_out[33];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[34] = s_CSAwallace_cska24_csa4_csa_component_out[34];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[35] = s_CSAwallace_cska24_csa4_csa_component_out[35];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[36] = s_CSAwallace_cska24_csa4_csa_component_out[36];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[37] = s_CSAwallace_cska24_csa4_csa_component_out[37];
  assign s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5[38] = 1'b1;
  csa_component39 csa_component39_s_CSAwallace_cska24_csa10_csa_component_out(.a(s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s4), .b(s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_c4), .c(s_CSAwallace_cska24_csa10_csa_component_s_CSAwallace_cska24_csa_s5), .csa_component39_out(s_CSAwallace_cska24_csa10_csa_component_out));
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[0] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[1] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[2] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[3] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[4] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[5] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[6] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[7] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[8] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[9] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[10] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[11] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[12] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[13] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[14] = s_CSAwallace_cska24_csa4_csa_component_out[53];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[15] = s_CSAwallace_cska24_csa4_csa_component_out[54];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[16] = s_CSAwallace_cska24_csa4_csa_component_out[55];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[17] = s_CSAwallace_cska24_csa4_csa_component_out[56];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[18] = s_CSAwallace_cska24_csa4_csa_component_out[57];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[19] = s_CSAwallace_cska24_csa4_csa_component_out[58];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[20] = s_CSAwallace_cska24_csa4_csa_component_out[59];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[21] = s_CSAwallace_cska24_csa4_csa_component_out[60];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[22] = s_CSAwallace_cska24_csa4_csa_component_out[61];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[23] = s_CSAwallace_cska24_csa4_csa_component_out[62];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[24] = s_CSAwallace_cska24_csa4_csa_component_out[63];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[25] = s_CSAwallace_cska24_csa4_csa_component_out[64];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[26] = s_CSAwallace_cska24_csa4_csa_component_out[65];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[27] = s_CSAwallace_cska24_csa4_csa_component_out[66];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[28] = s_CSAwallace_cska24_csa4_csa_component_out[67];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[29] = s_CSAwallace_cska24_csa4_csa_component_out[68];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[30] = s_CSAwallace_cska24_csa4_csa_component_out[69];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[31] = s_CSAwallace_cska24_csa4_csa_component_out[70];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[32] = s_CSAwallace_cska24_csa4_csa_component_out[71];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[33] = s_CSAwallace_cska24_csa4_csa_component_out[72];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[34] = s_CSAwallace_cska24_csa4_csa_component_out[73];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[35] = s_CSAwallace_cska24_csa4_csa_component_out[74];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[36] = s_CSAwallace_cska24_csa4_csa_component_out[75];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[37] = s_CSAwallace_cska24_csa4_csa_component_out[76];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[38] = 1'b1;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[39] = 1'b1;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[40] = 1'b1;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5[41] = 1'b1;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[0] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[1] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[2] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[3] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[4] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[5] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[6] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[7] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[8] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[9] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[10] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[11] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[12] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[13] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[14] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[15] = s_CSAwallace_cska24_csa5_csa_component_out[15];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[16] = s_CSAwallace_cska24_csa5_csa_component_out[16];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[17] = s_CSAwallace_cska24_csa5_csa_component_out[17];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[18] = s_CSAwallace_cska24_csa5_csa_component_out[18];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[19] = s_CSAwallace_cska24_csa5_csa_component_out[19];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[20] = s_CSAwallace_cska24_csa5_csa_component_out[20];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[21] = s_CSAwallace_cska24_csa5_csa_component_out[21];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[22] = s_CSAwallace_cska24_csa5_csa_component_out[22];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[23] = s_CSAwallace_cska24_csa5_csa_component_out[23];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[24] = s_CSAwallace_cska24_csa5_csa_component_out[24];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[25] = s_CSAwallace_cska24_csa5_csa_component_out[25];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[26] = s_CSAwallace_cska24_csa5_csa_component_out[26];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[27] = s_CSAwallace_cska24_csa5_csa_component_out[27];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[28] = s_CSAwallace_cska24_csa5_csa_component_out[28];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[29] = s_CSAwallace_cska24_csa5_csa_component_out[29];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[30] = s_CSAwallace_cska24_csa5_csa_component_out[30];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[31] = s_CSAwallace_cska24_csa5_csa_component_out[31];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[32] = s_CSAwallace_cska24_csa5_csa_component_out[32];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[33] = s_CSAwallace_cska24_csa5_csa_component_out[33];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[34] = s_CSAwallace_cska24_csa5_csa_component_out[34];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[35] = s_CSAwallace_cska24_csa5_csa_component_out[35];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[36] = s_CSAwallace_cska24_csa5_csa_component_out[36];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[37] = s_CSAwallace_cska24_csa5_csa_component_out[37];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[38] = s_CSAwallace_cska24_csa5_csa_component_out[38];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[39] = s_CSAwallace_cska24_csa5_csa_component_out[39];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[40] = s_CSAwallace_cska24_csa5_csa_component_out[40];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6[41] = 1'b1;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[0] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[1] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[2] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[3] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[4] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[5] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[6] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[7] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[8] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[9] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[10] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[11] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[12] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[13] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[14] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[15] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[16] = 1'b0;
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[17] = s_CSAwallace_cska24_csa5_csa_component_out[59];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[18] = s_CSAwallace_cska24_csa5_csa_component_out[60];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[19] = s_CSAwallace_cska24_csa5_csa_component_out[61];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[20] = s_CSAwallace_cska24_csa5_csa_component_out[62];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[21] = s_CSAwallace_cska24_csa5_csa_component_out[63];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[22] = s_CSAwallace_cska24_csa5_csa_component_out[64];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[23] = s_CSAwallace_cska24_csa5_csa_component_out[65];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[24] = s_CSAwallace_cska24_csa5_csa_component_out[66];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[25] = s_CSAwallace_cska24_csa5_csa_component_out[67];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[26] = s_CSAwallace_cska24_csa5_csa_component_out[68];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[27] = s_CSAwallace_cska24_csa5_csa_component_out[69];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[28] = s_CSAwallace_cska24_csa5_csa_component_out[70];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[29] = s_CSAwallace_cska24_csa5_csa_component_out[71];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[30] = s_CSAwallace_cska24_csa5_csa_component_out[72];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[31] = s_CSAwallace_cska24_csa5_csa_component_out[73];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[32] = s_CSAwallace_cska24_csa5_csa_component_out[74];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[33] = s_CSAwallace_cska24_csa5_csa_component_out[75];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[34] = s_CSAwallace_cska24_csa5_csa_component_out[76];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[35] = s_CSAwallace_cska24_csa5_csa_component_out[77];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[36] = s_CSAwallace_cska24_csa5_csa_component_out[78];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[37] = s_CSAwallace_cska24_csa5_csa_component_out[79];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[38] = s_CSAwallace_cska24_csa5_csa_component_out[80];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[39] = s_CSAwallace_cska24_csa5_csa_component_out[81];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[40] = s_CSAwallace_cska24_csa5_csa_component_out[82];
  assign s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6[41] = 1'b1;
  csa_component42 csa_component42_s_CSAwallace_cska24_csa11_csa_component_out(.a(s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c5), .b(s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_s6), .c(s_CSAwallace_cska24_csa11_csa_component_s_CSAwallace_cska24_csa_c6), .csa_component42_out(s_CSAwallace_cska24_csa11_csa_component_out));
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[0] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[1] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[2] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[3] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[4] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[5] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[6] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[7] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[8] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[9] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[10] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[11] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[12] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[13] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[14] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[15] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[16] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[17] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[18] = s_CSAwallace_cska24_csa6_csa_component_out[18];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[19] = s_CSAwallace_cska24_csa6_csa_component_out[19];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[20] = s_CSAwallace_cska24_csa6_csa_component_out[20];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[21] = s_CSAwallace_cska24_csa6_csa_component_out[21];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[22] = s_CSAwallace_cska24_csa6_csa_component_out[22];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[23] = s_CSAwallace_cska24_csa6_csa_component_out[23];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[24] = s_CSAwallace_cska24_csa6_csa_component_out[24];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[25] = s_CSAwallace_cska24_csa6_csa_component_out[25];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[26] = s_CSAwallace_cska24_csa6_csa_component_out[26];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[27] = s_CSAwallace_cska24_csa6_csa_component_out[27];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[28] = s_CSAwallace_cska24_csa6_csa_component_out[28];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[29] = s_CSAwallace_cska24_csa6_csa_component_out[29];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[30] = s_CSAwallace_cska24_csa6_csa_component_out[30];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[31] = s_CSAwallace_cska24_csa6_csa_component_out[31];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[32] = s_CSAwallace_cska24_csa6_csa_component_out[32];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[33] = s_CSAwallace_cska24_csa6_csa_component_out[33];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[34] = s_CSAwallace_cska24_csa6_csa_component_out[34];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[35] = s_CSAwallace_cska24_csa6_csa_component_out[35];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[36] = s_CSAwallace_cska24_csa6_csa_component_out[36];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[37] = s_CSAwallace_cska24_csa6_csa_component_out[37];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[38] = s_CSAwallace_cska24_csa6_csa_component_out[38];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[39] = s_CSAwallace_cska24_csa6_csa_component_out[39];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[40] = s_CSAwallace_cska24_csa6_csa_component_out[40];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[41] = s_CSAwallace_cska24_csa6_csa_component_out[41];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[42] = s_CSAwallace_cska24_csa6_csa_component_out[42];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[43] = s_CSAwallace_cska24_csa6_csa_component_out[43];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[44] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[45] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[46] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7[47] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[0] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[1] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[2] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[3] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[4] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[5] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[6] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[7] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[8] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[9] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[10] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[11] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[12] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[13] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[14] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[15] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[16] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[17] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[18] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[19] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[20] = s_CSAwallace_cska24_csa6_csa_component_out[65];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[21] = s_CSAwallace_cska24_csa6_csa_component_out[66];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[22] = s_CSAwallace_cska24_csa6_csa_component_out[67];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[23] = s_CSAwallace_cska24_csa6_csa_component_out[68];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[24] = s_CSAwallace_cska24_csa6_csa_component_out[69];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[25] = s_CSAwallace_cska24_csa6_csa_component_out[70];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[26] = s_CSAwallace_cska24_csa6_csa_component_out[71];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[27] = s_CSAwallace_cska24_csa6_csa_component_out[72];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[28] = s_CSAwallace_cska24_csa6_csa_component_out[73];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[29] = s_CSAwallace_cska24_csa6_csa_component_out[74];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[30] = s_CSAwallace_cska24_csa6_csa_component_out[75];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[31] = s_CSAwallace_cska24_csa6_csa_component_out[76];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[32] = s_CSAwallace_cska24_csa6_csa_component_out[77];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[33] = s_CSAwallace_cska24_csa6_csa_component_out[78];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[34] = s_CSAwallace_cska24_csa6_csa_component_out[79];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[35] = s_CSAwallace_cska24_csa6_csa_component_out[80];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[36] = s_CSAwallace_cska24_csa6_csa_component_out[81];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[37] = s_CSAwallace_cska24_csa6_csa_component_out[82];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[38] = s_CSAwallace_cska24_csa6_csa_component_out[83];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[39] = s_CSAwallace_cska24_csa6_csa_component_out[84];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[40] = s_CSAwallace_cska24_csa6_csa_component_out[85];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[41] = s_CSAwallace_cska24_csa6_csa_component_out[86];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[42] = s_CSAwallace_cska24_csa6_csa_component_out[87];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[43] = s_CSAwallace_cska24_csa6_csa_component_out[88];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[44] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[45] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[46] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7[47] = 1'b1;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[0] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[1] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[2] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[3] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[4] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[5] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[6] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[7] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[8] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[9] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[10] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[11] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[12] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[13] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[14] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[15] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[16] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[17] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[18] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[19] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[20] = 1'b0;
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[21] = s_CSAwallace_cska24_csa7_csa_component_out[21];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[22] = s_CSAwallace_cska24_csa7_csa_component_out[22];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[23] = s_CSAwallace_cska24_csa7_csa_component_out[23];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[24] = s_CSAwallace_cska24_csa7_csa_component_out[24];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[25] = s_CSAwallace_cska24_csa7_csa_component_out[25];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[26] = s_CSAwallace_cska24_csa7_csa_component_out[26];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[27] = s_CSAwallace_cska24_csa7_csa_component_out[27];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[28] = s_CSAwallace_cska24_csa7_csa_component_out[28];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[29] = s_CSAwallace_cska24_csa7_csa_component_out[29];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[30] = s_CSAwallace_cska24_csa7_csa_component_out[30];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[31] = s_CSAwallace_cska24_csa7_csa_component_out[31];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[32] = s_CSAwallace_cska24_csa7_csa_component_out[32];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[33] = s_CSAwallace_cska24_csa7_csa_component_out[33];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[34] = s_CSAwallace_cska24_csa7_csa_component_out[34];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[35] = s_CSAwallace_cska24_csa7_csa_component_out[35];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[36] = s_CSAwallace_cska24_csa7_csa_component_out[36];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[37] = s_CSAwallace_cska24_csa7_csa_component_out[37];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[38] = s_CSAwallace_cska24_csa7_csa_component_out[38];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[39] = s_CSAwallace_cska24_csa7_csa_component_out[39];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[40] = s_CSAwallace_cska24_csa7_csa_component_out[40];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[41] = s_CSAwallace_cska24_csa7_csa_component_out[41];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[42] = s_CSAwallace_cska24_csa7_csa_component_out[42];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[43] = s_CSAwallace_cska24_csa7_csa_component_out[43];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[44] = s_CSAwallace_cska24_csa7_csa_component_out[44];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[45] = s_CSAwallace_cska24_csa7_csa_component_out[45];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[46] = s_CSAwallace_cska24_csa7_csa_component_out[46];
  assign s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8[47] = 1'b1;
  csa_component48 csa_component48_s_CSAwallace_cska24_csa12_csa_component_out(.a(s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s7), .b(s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_c7), .c(s_CSAwallace_cska24_csa12_csa_component_s_CSAwallace_cska24_csa_s8), .csa_component48_out(s_CSAwallace_cska24_csa12_csa_component_out));
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[0] = s_CSAwallace_cska24_csa8_csa_component_out[0];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[1] = s_CSAwallace_cska24_csa8_csa_component_out[1];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[2] = s_CSAwallace_cska24_csa8_csa_component_out[2];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[3] = s_CSAwallace_cska24_csa8_csa_component_out[3];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[4] = s_CSAwallace_cska24_csa8_csa_component_out[4];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[5] = s_CSAwallace_cska24_csa8_csa_component_out[5];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[6] = s_CSAwallace_cska24_csa8_csa_component_out[6];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[7] = s_CSAwallace_cska24_csa8_csa_component_out[7];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[8] = s_CSAwallace_cska24_csa8_csa_component_out[8];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[9] = s_CSAwallace_cska24_csa8_csa_component_out[9];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[10] = s_CSAwallace_cska24_csa8_csa_component_out[10];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[11] = s_CSAwallace_cska24_csa8_csa_component_out[11];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[12] = s_CSAwallace_cska24_csa8_csa_component_out[12];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[13] = s_CSAwallace_cska24_csa8_csa_component_out[13];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[14] = s_CSAwallace_cska24_csa8_csa_component_out[14];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[15] = s_CSAwallace_cska24_csa8_csa_component_out[15];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[16] = s_CSAwallace_cska24_csa8_csa_component_out[16];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[17] = s_CSAwallace_cska24_csa8_csa_component_out[17];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[18] = s_CSAwallace_cska24_csa8_csa_component_out[18];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[19] = s_CSAwallace_cska24_csa8_csa_component_out[19];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[20] = s_CSAwallace_cska24_csa8_csa_component_out[20];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[21] = s_CSAwallace_cska24_csa8_csa_component_out[21];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[22] = s_CSAwallace_cska24_csa8_csa_component_out[22];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[23] = s_CSAwallace_cska24_csa8_csa_component_out[23];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[24] = s_CSAwallace_cska24_csa8_csa_component_out[24];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[25] = s_CSAwallace_cska24_csa8_csa_component_out[25];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[26] = s_CSAwallace_cska24_csa8_csa_component_out[26];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[27] = s_CSAwallace_cska24_csa8_csa_component_out[27];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[28] = s_CSAwallace_cska24_csa8_csa_component_out[28];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[29] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[30] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[31] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[32] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9[33] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[0] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[1] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[2] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[3] = s_CSAwallace_cska24_csa8_csa_component_out[34];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[4] = s_CSAwallace_cska24_csa8_csa_component_out[35];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[5] = s_CSAwallace_cska24_csa8_csa_component_out[36];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[6] = s_CSAwallace_cska24_csa8_csa_component_out[37];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[7] = s_CSAwallace_cska24_csa8_csa_component_out[38];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[8] = s_CSAwallace_cska24_csa8_csa_component_out[39];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[9] = s_CSAwallace_cska24_csa8_csa_component_out[40];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[10] = s_CSAwallace_cska24_csa8_csa_component_out[41];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[11] = s_CSAwallace_cska24_csa8_csa_component_out[42];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[12] = s_CSAwallace_cska24_csa8_csa_component_out[43];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[13] = s_CSAwallace_cska24_csa8_csa_component_out[44];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[14] = s_CSAwallace_cska24_csa8_csa_component_out[45];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[15] = s_CSAwallace_cska24_csa8_csa_component_out[46];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[16] = s_CSAwallace_cska24_csa8_csa_component_out[47];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[17] = s_CSAwallace_cska24_csa8_csa_component_out[48];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[18] = s_CSAwallace_cska24_csa8_csa_component_out[49];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[19] = s_CSAwallace_cska24_csa8_csa_component_out[50];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[20] = s_CSAwallace_cska24_csa8_csa_component_out[51];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[21] = s_CSAwallace_cska24_csa8_csa_component_out[52];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[22] = s_CSAwallace_cska24_csa8_csa_component_out[53];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[23] = s_CSAwallace_cska24_csa8_csa_component_out[54];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[24] = s_CSAwallace_cska24_csa8_csa_component_out[55];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[25] = s_CSAwallace_cska24_csa8_csa_component_out[56];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[26] = s_CSAwallace_cska24_csa8_csa_component_out[57];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[27] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[28] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[29] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[30] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[31] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[32] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9[33] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[0] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[1] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[2] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[3] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[4] = 1'b0;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[5] = s_CSAwallace_cska24_csa9_csa_component_out[5];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[6] = s_CSAwallace_cska24_csa9_csa_component_out[6];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[7] = s_CSAwallace_cska24_csa9_csa_component_out[7];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[8] = s_CSAwallace_cska24_csa9_csa_component_out[8];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[9] = s_CSAwallace_cska24_csa9_csa_component_out[9];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[10] = s_CSAwallace_cska24_csa9_csa_component_out[10];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[11] = s_CSAwallace_cska24_csa9_csa_component_out[11];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[12] = s_CSAwallace_cska24_csa9_csa_component_out[12];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[13] = s_CSAwallace_cska24_csa9_csa_component_out[13];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[14] = s_CSAwallace_cska24_csa9_csa_component_out[14];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[15] = s_CSAwallace_cska24_csa9_csa_component_out[15];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[16] = s_CSAwallace_cska24_csa9_csa_component_out[16];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[17] = s_CSAwallace_cska24_csa9_csa_component_out[17];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[18] = s_CSAwallace_cska24_csa9_csa_component_out[18];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[19] = s_CSAwallace_cska24_csa9_csa_component_out[19];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[20] = s_CSAwallace_cska24_csa9_csa_component_out[20];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[21] = s_CSAwallace_cska24_csa9_csa_component_out[21];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[22] = s_CSAwallace_cska24_csa9_csa_component_out[22];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[23] = s_CSAwallace_cska24_csa9_csa_component_out[23];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[24] = s_CSAwallace_cska24_csa9_csa_component_out[24];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[25] = s_CSAwallace_cska24_csa9_csa_component_out[25];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[26] = s_CSAwallace_cska24_csa9_csa_component_out[26];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[27] = s_CSAwallace_cska24_csa9_csa_component_out[27];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[28] = s_CSAwallace_cska24_csa9_csa_component_out[28];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[29] = s_CSAwallace_cska24_csa9_csa_component_out[29];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[30] = s_CSAwallace_cska24_csa9_csa_component_out[30];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[31] = s_CSAwallace_cska24_csa9_csa_component_out[31];
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[32] = 1'b1;
  assign s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10[33] = 1'b1;
  csa_component34 csa_component34_s_CSAwallace_cska24_csa13_csa_component_out(.a(s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s9), .b(s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_c9), .c(s_CSAwallace_cska24_csa13_csa_component_s_CSAwallace_cska24_csa_s10), .csa_component34_out(s_CSAwallace_cska24_csa13_csa_component_out));
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[0] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[1] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[2] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[3] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[4] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[5] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[6] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[7] = s_CSAwallace_cska24_csa9_csa_component_out[41];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[8] = s_CSAwallace_cska24_csa9_csa_component_out[42];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[9] = s_CSAwallace_cska24_csa9_csa_component_out[43];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[10] = s_CSAwallace_cska24_csa9_csa_component_out[44];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[11] = s_CSAwallace_cska24_csa9_csa_component_out[45];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[12] = s_CSAwallace_cska24_csa9_csa_component_out[46];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[13] = s_CSAwallace_cska24_csa9_csa_component_out[47];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[14] = s_CSAwallace_cska24_csa9_csa_component_out[48];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[15] = s_CSAwallace_cska24_csa9_csa_component_out[49];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[16] = s_CSAwallace_cska24_csa9_csa_component_out[50];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[17] = s_CSAwallace_cska24_csa9_csa_component_out[51];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[18] = s_CSAwallace_cska24_csa9_csa_component_out[52];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[19] = s_CSAwallace_cska24_csa9_csa_component_out[53];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[20] = s_CSAwallace_cska24_csa9_csa_component_out[54];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[21] = s_CSAwallace_cska24_csa9_csa_component_out[55];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[22] = s_CSAwallace_cska24_csa9_csa_component_out[56];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[23] = s_CSAwallace_cska24_csa9_csa_component_out[57];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[24] = s_CSAwallace_cska24_csa9_csa_component_out[58];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[25] = s_CSAwallace_cska24_csa9_csa_component_out[59];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[26] = s_CSAwallace_cska24_csa9_csa_component_out[60];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[27] = s_CSAwallace_cska24_csa9_csa_component_out[61];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[28] = s_CSAwallace_cska24_csa9_csa_component_out[62];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[29] = s_CSAwallace_cska24_csa9_csa_component_out[63];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[30] = s_CSAwallace_cska24_csa9_csa_component_out[64];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[31] = s_CSAwallace_cska24_csa9_csa_component_out[65];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[32] = s_CSAwallace_cska24_csa9_csa_component_out[66];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[33] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[34] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[35] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[36] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[37] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[38] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10[39] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[0] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[1] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[2] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[3] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[4] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[5] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[6] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[7] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[8] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[9] = s_CSAwallace_cska24_csa10_csa_component_out[9];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[10] = s_CSAwallace_cska24_csa10_csa_component_out[10];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[11] = s_CSAwallace_cska24_csa10_csa_component_out[11];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[12] = s_CSAwallace_cska24_csa10_csa_component_out[12];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[13] = s_CSAwallace_cska24_csa10_csa_component_out[13];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[14] = s_CSAwallace_cska24_csa10_csa_component_out[14];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[15] = s_CSAwallace_cska24_csa10_csa_component_out[15];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[16] = s_CSAwallace_cska24_csa10_csa_component_out[16];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[17] = s_CSAwallace_cska24_csa10_csa_component_out[17];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[18] = s_CSAwallace_cska24_csa10_csa_component_out[18];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[19] = s_CSAwallace_cska24_csa10_csa_component_out[19];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[20] = s_CSAwallace_cska24_csa10_csa_component_out[20];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[21] = s_CSAwallace_cska24_csa10_csa_component_out[21];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[22] = s_CSAwallace_cska24_csa10_csa_component_out[22];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[23] = s_CSAwallace_cska24_csa10_csa_component_out[23];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[24] = s_CSAwallace_cska24_csa10_csa_component_out[24];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[25] = s_CSAwallace_cska24_csa10_csa_component_out[25];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[26] = s_CSAwallace_cska24_csa10_csa_component_out[26];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[27] = s_CSAwallace_cska24_csa10_csa_component_out[27];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[28] = s_CSAwallace_cska24_csa10_csa_component_out[28];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[29] = s_CSAwallace_cska24_csa10_csa_component_out[29];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[30] = s_CSAwallace_cska24_csa10_csa_component_out[30];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[31] = s_CSAwallace_cska24_csa10_csa_component_out[31];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[32] = s_CSAwallace_cska24_csa10_csa_component_out[32];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[33] = s_CSAwallace_cska24_csa10_csa_component_out[33];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[34] = s_CSAwallace_cska24_csa10_csa_component_out[34];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[35] = s_CSAwallace_cska24_csa10_csa_component_out[35];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[36] = s_CSAwallace_cska24_csa10_csa_component_out[36];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[37] = s_CSAwallace_cska24_csa10_csa_component_out[37];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[38] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11[39] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[0] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[1] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[2] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[3] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[4] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[5] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[6] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[7] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[8] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[9] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[10] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[11] = 1'b0;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[12] = s_CSAwallace_cska24_csa10_csa_component_out[52];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[13] = s_CSAwallace_cska24_csa10_csa_component_out[53];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[14] = s_CSAwallace_cska24_csa10_csa_component_out[54];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[15] = s_CSAwallace_cska24_csa10_csa_component_out[55];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[16] = s_CSAwallace_cska24_csa10_csa_component_out[56];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[17] = s_CSAwallace_cska24_csa10_csa_component_out[57];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[18] = s_CSAwallace_cska24_csa10_csa_component_out[58];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[19] = s_CSAwallace_cska24_csa10_csa_component_out[59];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[20] = s_CSAwallace_cska24_csa10_csa_component_out[60];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[21] = s_CSAwallace_cska24_csa10_csa_component_out[61];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[22] = s_CSAwallace_cska24_csa10_csa_component_out[62];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[23] = s_CSAwallace_cska24_csa10_csa_component_out[63];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[24] = s_CSAwallace_cska24_csa10_csa_component_out[64];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[25] = s_CSAwallace_cska24_csa10_csa_component_out[65];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[26] = s_CSAwallace_cska24_csa10_csa_component_out[66];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[27] = s_CSAwallace_cska24_csa10_csa_component_out[67];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[28] = s_CSAwallace_cska24_csa10_csa_component_out[68];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[29] = s_CSAwallace_cska24_csa10_csa_component_out[69];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[30] = s_CSAwallace_cska24_csa10_csa_component_out[70];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[31] = s_CSAwallace_cska24_csa10_csa_component_out[71];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[32] = s_CSAwallace_cska24_csa10_csa_component_out[72];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[33] = s_CSAwallace_cska24_csa10_csa_component_out[73];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[34] = s_CSAwallace_cska24_csa10_csa_component_out[74];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[35] = s_CSAwallace_cska24_csa10_csa_component_out[75];
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[36] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[37] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[38] = 1'b1;
  assign s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11[39] = 1'b1;
  csa_component40 csa_component40_s_CSAwallace_cska24_csa14_csa_component_out(.a(s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c10), .b(s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_s11), .c(s_CSAwallace_cska24_csa14_csa_component_s_CSAwallace_cska24_csa_c11), .csa_component40_out(s_CSAwallace_cska24_csa14_csa_component_out));
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[0] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[1] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[2] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[3] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[4] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[5] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[6] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[7] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[8] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[9] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[10] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[11] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[12] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[13] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[14] = s_CSAwallace_cska24_csa11_csa_component_out[14];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[15] = s_CSAwallace_cska24_csa11_csa_component_out[15];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[16] = s_CSAwallace_cska24_csa11_csa_component_out[16];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[17] = s_CSAwallace_cska24_csa11_csa_component_out[17];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[18] = s_CSAwallace_cska24_csa11_csa_component_out[18];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[19] = s_CSAwallace_cska24_csa11_csa_component_out[19];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[20] = s_CSAwallace_cska24_csa11_csa_component_out[20];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[21] = s_CSAwallace_cska24_csa11_csa_component_out[21];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[22] = s_CSAwallace_cska24_csa11_csa_component_out[22];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[23] = s_CSAwallace_cska24_csa11_csa_component_out[23];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[24] = s_CSAwallace_cska24_csa11_csa_component_out[24];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[25] = s_CSAwallace_cska24_csa11_csa_component_out[25];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[26] = s_CSAwallace_cska24_csa11_csa_component_out[26];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[27] = s_CSAwallace_cska24_csa11_csa_component_out[27];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[28] = s_CSAwallace_cska24_csa11_csa_component_out[28];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[29] = s_CSAwallace_cska24_csa11_csa_component_out[29];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[30] = s_CSAwallace_cska24_csa11_csa_component_out[30];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[31] = s_CSAwallace_cska24_csa11_csa_component_out[31];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[32] = s_CSAwallace_cska24_csa11_csa_component_out[32];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[33] = s_CSAwallace_cska24_csa11_csa_component_out[33];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[34] = s_CSAwallace_cska24_csa11_csa_component_out[34];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[35] = s_CSAwallace_cska24_csa11_csa_component_out[35];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[36] = s_CSAwallace_cska24_csa11_csa_component_out[36];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[37] = s_CSAwallace_cska24_csa11_csa_component_out[37];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[38] = s_CSAwallace_cska24_csa11_csa_component_out[38];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[39] = s_CSAwallace_cska24_csa11_csa_component_out[39];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[40] = s_CSAwallace_cska24_csa11_csa_component_out[40];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[41] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[42] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[43] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[44] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[45] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[46] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12[47] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[0] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[1] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[2] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[3] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[4] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[5] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[6] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[7] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[8] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[9] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[10] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[11] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[12] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[13] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[14] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[15] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[16] = s_CSAwallace_cska24_csa11_csa_component_out[59];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[17] = s_CSAwallace_cska24_csa11_csa_component_out[60];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[18] = s_CSAwallace_cska24_csa11_csa_component_out[61];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[19] = s_CSAwallace_cska24_csa11_csa_component_out[62];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[20] = s_CSAwallace_cska24_csa11_csa_component_out[63];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[21] = s_CSAwallace_cska24_csa11_csa_component_out[64];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[22] = s_CSAwallace_cska24_csa11_csa_component_out[65];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[23] = s_CSAwallace_cska24_csa11_csa_component_out[66];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[24] = s_CSAwallace_cska24_csa11_csa_component_out[67];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[25] = s_CSAwallace_cska24_csa11_csa_component_out[68];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[26] = s_CSAwallace_cska24_csa11_csa_component_out[69];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[27] = s_CSAwallace_cska24_csa11_csa_component_out[70];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[28] = s_CSAwallace_cska24_csa11_csa_component_out[71];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[29] = s_CSAwallace_cska24_csa11_csa_component_out[72];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[30] = s_CSAwallace_cska24_csa11_csa_component_out[73];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[31] = s_CSAwallace_cska24_csa11_csa_component_out[74];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[32] = s_CSAwallace_cska24_csa11_csa_component_out[75];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[33] = s_CSAwallace_cska24_csa11_csa_component_out[76];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[34] = s_CSAwallace_cska24_csa11_csa_component_out[77];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[35] = s_CSAwallace_cska24_csa11_csa_component_out[78];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[36] = s_CSAwallace_cska24_csa11_csa_component_out[79];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[37] = s_CSAwallace_cska24_csa11_csa_component_out[80];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[38] = s_CSAwallace_cska24_csa11_csa_component_out[81];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[39] = s_CSAwallace_cska24_csa11_csa_component_out[82];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[40] = s_CSAwallace_cska24_csa11_csa_component_out[83];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[41] = s_CSAwallace_cska24_csa11_csa_component_out[84];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[42] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[43] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[44] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[45] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[46] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12[47] = 1'b1;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[0] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[1] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[2] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[3] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[4] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[5] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[6] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[7] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[8] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[9] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[10] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[11] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[12] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[13] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[14] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[15] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[16] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[17] = 1'b0;
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[18] = s_CSAwallace_cska24_csa12_csa_component_out[18];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[19] = s_CSAwallace_cska24_csa12_csa_component_out[19];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[20] = s_CSAwallace_cska24_csa12_csa_component_out[20];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[21] = s_CSAwallace_cska24_csa12_csa_component_out[21];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[22] = s_CSAwallace_cska24_csa12_csa_component_out[22];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[23] = s_CSAwallace_cska24_csa12_csa_component_out[23];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[24] = s_CSAwallace_cska24_csa12_csa_component_out[24];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[25] = s_CSAwallace_cska24_csa12_csa_component_out[25];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[26] = s_CSAwallace_cska24_csa12_csa_component_out[26];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[27] = s_CSAwallace_cska24_csa12_csa_component_out[27];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[28] = s_CSAwallace_cska24_csa12_csa_component_out[28];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[29] = s_CSAwallace_cska24_csa12_csa_component_out[29];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[30] = s_CSAwallace_cska24_csa12_csa_component_out[30];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[31] = s_CSAwallace_cska24_csa12_csa_component_out[31];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[32] = s_CSAwallace_cska24_csa12_csa_component_out[32];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[33] = s_CSAwallace_cska24_csa12_csa_component_out[33];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[34] = s_CSAwallace_cska24_csa12_csa_component_out[34];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[35] = s_CSAwallace_cska24_csa12_csa_component_out[35];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[36] = s_CSAwallace_cska24_csa12_csa_component_out[36];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[37] = s_CSAwallace_cska24_csa12_csa_component_out[37];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[38] = s_CSAwallace_cska24_csa12_csa_component_out[38];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[39] = s_CSAwallace_cska24_csa12_csa_component_out[39];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[40] = s_CSAwallace_cska24_csa12_csa_component_out[40];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[41] = s_CSAwallace_cska24_csa12_csa_component_out[41];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[42] = s_CSAwallace_cska24_csa12_csa_component_out[42];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[43] = s_CSAwallace_cska24_csa12_csa_component_out[43];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[44] = s_CSAwallace_cska24_csa12_csa_component_out[44];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[45] = s_CSAwallace_cska24_csa12_csa_component_out[45];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[46] = s_CSAwallace_cska24_csa12_csa_component_out[46];
  assign s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13[47] = 1'b1;
  csa_component48 csa_component48_s_CSAwallace_cska24_csa15_csa_component_out(.a(s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s12), .b(s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_c12), .c(s_CSAwallace_cska24_csa15_csa_component_s_CSAwallace_cska24_csa_s13), .csa_component48_out(s_CSAwallace_cska24_csa15_csa_component_out));
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[0] = s_CSAwallace_cska24_csa13_csa_component_out[0];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[1] = s_CSAwallace_cska24_csa13_csa_component_out[1];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[2] = s_CSAwallace_cska24_csa13_csa_component_out[2];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[3] = s_CSAwallace_cska24_csa13_csa_component_out[3];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[4] = s_CSAwallace_cska24_csa13_csa_component_out[4];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[5] = s_CSAwallace_cska24_csa13_csa_component_out[5];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[6] = s_CSAwallace_cska24_csa13_csa_component_out[6];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[7] = s_CSAwallace_cska24_csa13_csa_component_out[7];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[8] = s_CSAwallace_cska24_csa13_csa_component_out[8];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[9] = s_CSAwallace_cska24_csa13_csa_component_out[9];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[10] = s_CSAwallace_cska24_csa13_csa_component_out[10];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[11] = s_CSAwallace_cska24_csa13_csa_component_out[11];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[12] = s_CSAwallace_cska24_csa13_csa_component_out[12];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[13] = s_CSAwallace_cska24_csa13_csa_component_out[13];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[14] = s_CSAwallace_cska24_csa13_csa_component_out[14];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[15] = s_CSAwallace_cska24_csa13_csa_component_out[15];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[16] = s_CSAwallace_cska24_csa13_csa_component_out[16];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[17] = s_CSAwallace_cska24_csa13_csa_component_out[17];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[18] = s_CSAwallace_cska24_csa13_csa_component_out[18];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[19] = s_CSAwallace_cska24_csa13_csa_component_out[19];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[20] = s_CSAwallace_cska24_csa13_csa_component_out[20];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[21] = s_CSAwallace_cska24_csa13_csa_component_out[21];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[22] = s_CSAwallace_cska24_csa13_csa_component_out[22];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[23] = s_CSAwallace_cska24_csa13_csa_component_out[23];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[24] = s_CSAwallace_cska24_csa13_csa_component_out[24];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[25] = s_CSAwallace_cska24_csa13_csa_component_out[25];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[26] = s_CSAwallace_cska24_csa13_csa_component_out[26];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[27] = s_CSAwallace_cska24_csa13_csa_component_out[27];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[28] = s_CSAwallace_cska24_csa13_csa_component_out[28];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[29] = s_CSAwallace_cska24_csa13_csa_component_out[29];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[30] = s_CSAwallace_cska24_csa13_csa_component_out[30];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[31] = s_CSAwallace_cska24_csa13_csa_component_out[31];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[32] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[33] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[34] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[35] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[36] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[37] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[38] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[39] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14[40] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[0] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[1] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[2] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[3] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[4] = s_CSAwallace_cska24_csa13_csa_component_out[39];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[5] = s_CSAwallace_cska24_csa13_csa_component_out[40];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[6] = s_CSAwallace_cska24_csa13_csa_component_out[41];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[7] = s_CSAwallace_cska24_csa13_csa_component_out[42];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[8] = s_CSAwallace_cska24_csa13_csa_component_out[43];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[9] = s_CSAwallace_cska24_csa13_csa_component_out[44];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[10] = s_CSAwallace_cska24_csa13_csa_component_out[45];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[11] = s_CSAwallace_cska24_csa13_csa_component_out[46];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[12] = s_CSAwallace_cska24_csa13_csa_component_out[47];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[13] = s_CSAwallace_cska24_csa13_csa_component_out[48];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[14] = s_CSAwallace_cska24_csa13_csa_component_out[49];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[15] = s_CSAwallace_cska24_csa13_csa_component_out[50];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[16] = s_CSAwallace_cska24_csa13_csa_component_out[51];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[17] = s_CSAwallace_cska24_csa13_csa_component_out[52];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[18] = s_CSAwallace_cska24_csa13_csa_component_out[53];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[19] = s_CSAwallace_cska24_csa13_csa_component_out[54];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[20] = s_CSAwallace_cska24_csa13_csa_component_out[55];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[21] = s_CSAwallace_cska24_csa13_csa_component_out[56];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[22] = s_CSAwallace_cska24_csa13_csa_component_out[57];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[23] = s_CSAwallace_cska24_csa13_csa_component_out[58];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[24] = s_CSAwallace_cska24_csa13_csa_component_out[59];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[25] = s_CSAwallace_cska24_csa13_csa_component_out[60];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[26] = s_CSAwallace_cska24_csa13_csa_component_out[61];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[27] = s_CSAwallace_cska24_csa13_csa_component_out[62];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[28] = s_CSAwallace_cska24_csa13_csa_component_out[63];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[29] = s_CSAwallace_cska24_csa13_csa_component_out[64];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[30] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[31] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[32] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[33] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[34] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[35] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[36] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[37] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[38] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[39] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14[40] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[0] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[1] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[2] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[3] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[4] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[5] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[6] = 1'b0;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[7] = s_CSAwallace_cska24_csa14_csa_component_out[7];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[8] = s_CSAwallace_cska24_csa14_csa_component_out[8];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[9] = s_CSAwallace_cska24_csa14_csa_component_out[9];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[10] = s_CSAwallace_cska24_csa14_csa_component_out[10];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[11] = s_CSAwallace_cska24_csa14_csa_component_out[11];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[12] = s_CSAwallace_cska24_csa14_csa_component_out[12];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[13] = s_CSAwallace_cska24_csa14_csa_component_out[13];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[14] = s_CSAwallace_cska24_csa14_csa_component_out[14];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[15] = s_CSAwallace_cska24_csa14_csa_component_out[15];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[16] = s_CSAwallace_cska24_csa14_csa_component_out[16];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[17] = s_CSAwallace_cska24_csa14_csa_component_out[17];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[18] = s_CSAwallace_cska24_csa14_csa_component_out[18];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[19] = s_CSAwallace_cska24_csa14_csa_component_out[19];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[20] = s_CSAwallace_cska24_csa14_csa_component_out[20];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[21] = s_CSAwallace_cska24_csa14_csa_component_out[21];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[22] = s_CSAwallace_cska24_csa14_csa_component_out[22];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[23] = s_CSAwallace_cska24_csa14_csa_component_out[23];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[24] = s_CSAwallace_cska24_csa14_csa_component_out[24];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[25] = s_CSAwallace_cska24_csa14_csa_component_out[25];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[26] = s_CSAwallace_cska24_csa14_csa_component_out[26];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[27] = s_CSAwallace_cska24_csa14_csa_component_out[27];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[28] = s_CSAwallace_cska24_csa14_csa_component_out[28];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[29] = s_CSAwallace_cska24_csa14_csa_component_out[29];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[30] = s_CSAwallace_cska24_csa14_csa_component_out[30];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[31] = s_CSAwallace_cska24_csa14_csa_component_out[31];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[32] = s_CSAwallace_cska24_csa14_csa_component_out[32];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[33] = s_CSAwallace_cska24_csa14_csa_component_out[33];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[34] = s_CSAwallace_cska24_csa14_csa_component_out[34];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[35] = s_CSAwallace_cska24_csa14_csa_component_out[35];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[36] = s_CSAwallace_cska24_csa14_csa_component_out[36];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[37] = s_CSAwallace_cska24_csa14_csa_component_out[37];
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[38] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[39] = 1'b1;
  assign s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15[40] = 1'b1;
  csa_component41 csa_component41_s_CSAwallace_cska24_csa16_csa_component_out(.a(s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s14), .b(s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_c14), .c(s_CSAwallace_cska24_csa16_csa_component_s_CSAwallace_cska24_csa_s15), .csa_component41_out(s_CSAwallace_cska24_csa16_csa_component_out));
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[0] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[1] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[2] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[3] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[4] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[5] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[6] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[7] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[8] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[9] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[10] = s_CSAwallace_cska24_csa14_csa_component_out[51];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[11] = s_CSAwallace_cska24_csa14_csa_component_out[52];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[12] = s_CSAwallace_cska24_csa14_csa_component_out[53];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[13] = s_CSAwallace_cska24_csa14_csa_component_out[54];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[14] = s_CSAwallace_cska24_csa14_csa_component_out[55];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[15] = s_CSAwallace_cska24_csa14_csa_component_out[56];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[16] = s_CSAwallace_cska24_csa14_csa_component_out[57];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[17] = s_CSAwallace_cska24_csa14_csa_component_out[58];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[18] = s_CSAwallace_cska24_csa14_csa_component_out[59];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[19] = s_CSAwallace_cska24_csa14_csa_component_out[60];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[20] = s_CSAwallace_cska24_csa14_csa_component_out[61];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[21] = s_CSAwallace_cska24_csa14_csa_component_out[62];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[22] = s_CSAwallace_cska24_csa14_csa_component_out[63];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[23] = s_CSAwallace_cska24_csa14_csa_component_out[64];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[24] = s_CSAwallace_cska24_csa14_csa_component_out[65];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[25] = s_CSAwallace_cska24_csa14_csa_component_out[66];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[26] = s_CSAwallace_cska24_csa14_csa_component_out[67];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[27] = s_CSAwallace_cska24_csa14_csa_component_out[68];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[28] = s_CSAwallace_cska24_csa14_csa_component_out[69];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[29] = s_CSAwallace_cska24_csa14_csa_component_out[70];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[30] = s_CSAwallace_cska24_csa14_csa_component_out[71];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[31] = s_CSAwallace_cska24_csa14_csa_component_out[72];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[32] = s_CSAwallace_cska24_csa14_csa_component_out[73];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[33] = s_CSAwallace_cska24_csa14_csa_component_out[74];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[34] = s_CSAwallace_cska24_csa14_csa_component_out[75];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[35] = s_CSAwallace_cska24_csa14_csa_component_out[76];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[36] = s_CSAwallace_cska24_csa14_csa_component_out[77];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[37] = s_CSAwallace_cska24_csa14_csa_component_out[78];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[38] = s_CSAwallace_cska24_csa14_csa_component_out[79];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[39] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[40] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[41] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[42] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[43] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[44] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[45] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[46] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15[47] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[0] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[1] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[2] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[3] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[4] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[5] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[6] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[7] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[8] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[9] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[10] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[11] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[12] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[13] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[14] = s_CSAwallace_cska24_csa15_csa_component_out[14];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[15] = s_CSAwallace_cska24_csa15_csa_component_out[15];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[16] = s_CSAwallace_cska24_csa15_csa_component_out[16];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[17] = s_CSAwallace_cska24_csa15_csa_component_out[17];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[18] = s_CSAwallace_cska24_csa15_csa_component_out[18];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[19] = s_CSAwallace_cska24_csa15_csa_component_out[19];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[20] = s_CSAwallace_cska24_csa15_csa_component_out[20];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[21] = s_CSAwallace_cska24_csa15_csa_component_out[21];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[22] = s_CSAwallace_cska24_csa15_csa_component_out[22];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[23] = s_CSAwallace_cska24_csa15_csa_component_out[23];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[24] = s_CSAwallace_cska24_csa15_csa_component_out[24];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[25] = s_CSAwallace_cska24_csa15_csa_component_out[25];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[26] = s_CSAwallace_cska24_csa15_csa_component_out[26];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[27] = s_CSAwallace_cska24_csa15_csa_component_out[27];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[28] = s_CSAwallace_cska24_csa15_csa_component_out[28];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[29] = s_CSAwallace_cska24_csa15_csa_component_out[29];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[30] = s_CSAwallace_cska24_csa15_csa_component_out[30];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[31] = s_CSAwallace_cska24_csa15_csa_component_out[31];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[32] = s_CSAwallace_cska24_csa15_csa_component_out[32];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[33] = s_CSAwallace_cska24_csa15_csa_component_out[33];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[34] = s_CSAwallace_cska24_csa15_csa_component_out[34];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[35] = s_CSAwallace_cska24_csa15_csa_component_out[35];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[36] = s_CSAwallace_cska24_csa15_csa_component_out[36];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[37] = s_CSAwallace_cska24_csa15_csa_component_out[37];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[38] = s_CSAwallace_cska24_csa15_csa_component_out[38];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[39] = s_CSAwallace_cska24_csa15_csa_component_out[39];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[40] = s_CSAwallace_cska24_csa15_csa_component_out[40];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[41] = s_CSAwallace_cska24_csa15_csa_component_out[41];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[42] = s_CSAwallace_cska24_csa15_csa_component_out[42];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[43] = s_CSAwallace_cska24_csa15_csa_component_out[43];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[44] = s_CSAwallace_cska24_csa15_csa_component_out[44];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[45] = s_CSAwallace_cska24_csa15_csa_component_out[45];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[46] = s_CSAwallace_cska24_csa15_csa_component_out[46];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16[47] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[0] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[1] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[2] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[3] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[4] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[5] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[6] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[7] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[8] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[9] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[10] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[11] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[12] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[13] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[14] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[15] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[16] = 1'b0;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[17] = s_CSAwallace_cska24_csa15_csa_component_out[66];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[18] = s_CSAwallace_cska24_csa15_csa_component_out[67];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[19] = s_CSAwallace_cska24_csa15_csa_component_out[68];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[20] = s_CSAwallace_cska24_csa15_csa_component_out[69];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[21] = s_CSAwallace_cska24_csa15_csa_component_out[70];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[22] = s_CSAwallace_cska24_csa15_csa_component_out[71];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[23] = s_CSAwallace_cska24_csa15_csa_component_out[72];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[24] = s_CSAwallace_cska24_csa15_csa_component_out[73];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[25] = s_CSAwallace_cska24_csa15_csa_component_out[74];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[26] = s_CSAwallace_cska24_csa15_csa_component_out[75];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[27] = s_CSAwallace_cska24_csa15_csa_component_out[76];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[28] = s_CSAwallace_cska24_csa15_csa_component_out[77];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[29] = s_CSAwallace_cska24_csa15_csa_component_out[78];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[30] = s_CSAwallace_cska24_csa15_csa_component_out[79];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[31] = s_CSAwallace_cska24_csa15_csa_component_out[80];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[32] = s_CSAwallace_cska24_csa15_csa_component_out[81];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[33] = s_CSAwallace_cska24_csa15_csa_component_out[82];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[34] = s_CSAwallace_cska24_csa15_csa_component_out[83];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[35] = s_CSAwallace_cska24_csa15_csa_component_out[84];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[36] = s_CSAwallace_cska24_csa15_csa_component_out[85];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[37] = s_CSAwallace_cska24_csa15_csa_component_out[86];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[38] = s_CSAwallace_cska24_csa15_csa_component_out[87];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[39] = s_CSAwallace_cska24_csa15_csa_component_out[88];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[40] = s_CSAwallace_cska24_csa15_csa_component_out[89];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[41] = s_CSAwallace_cska24_csa15_csa_component_out[90];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[42] = s_CSAwallace_cska24_csa15_csa_component_out[91];
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[43] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[44] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[45] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[46] = 1'b1;
  assign s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16[47] = 1'b1;
  csa_component48 csa_component48_s_CSAwallace_cska24_csa17_csa_component_out(.a(s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c15), .b(s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_s16), .c(s_CSAwallace_cska24_csa17_csa_component_s_CSAwallace_cska24_csa_c16), .csa_component48_out(s_CSAwallace_cska24_csa17_csa_component_out));
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[0] = s_CSAwallace_cska24_csa16_csa_component_out[0];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[1] = s_CSAwallace_cska24_csa16_csa_component_out[1];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[2] = s_CSAwallace_cska24_csa16_csa_component_out[2];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[3] = s_CSAwallace_cska24_csa16_csa_component_out[3];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[4] = s_CSAwallace_cska24_csa16_csa_component_out[4];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[5] = s_CSAwallace_cska24_csa16_csa_component_out[5];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[6] = s_CSAwallace_cska24_csa16_csa_component_out[6];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[7] = s_CSAwallace_cska24_csa16_csa_component_out[7];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[8] = s_CSAwallace_cska24_csa16_csa_component_out[8];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[9] = s_CSAwallace_cska24_csa16_csa_component_out[9];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[10] = s_CSAwallace_cska24_csa16_csa_component_out[10];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[11] = s_CSAwallace_cska24_csa16_csa_component_out[11];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[12] = s_CSAwallace_cska24_csa16_csa_component_out[12];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[13] = s_CSAwallace_cska24_csa16_csa_component_out[13];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[14] = s_CSAwallace_cska24_csa16_csa_component_out[14];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[15] = s_CSAwallace_cska24_csa16_csa_component_out[15];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[16] = s_CSAwallace_cska24_csa16_csa_component_out[16];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[17] = s_CSAwallace_cska24_csa16_csa_component_out[17];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[18] = s_CSAwallace_cska24_csa16_csa_component_out[18];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[19] = s_CSAwallace_cska24_csa16_csa_component_out[19];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[20] = s_CSAwallace_cska24_csa16_csa_component_out[20];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[21] = s_CSAwallace_cska24_csa16_csa_component_out[21];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[22] = s_CSAwallace_cska24_csa16_csa_component_out[22];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[23] = s_CSAwallace_cska24_csa16_csa_component_out[23];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[24] = s_CSAwallace_cska24_csa16_csa_component_out[24];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[25] = s_CSAwallace_cska24_csa16_csa_component_out[25];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[26] = s_CSAwallace_cska24_csa16_csa_component_out[26];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[27] = s_CSAwallace_cska24_csa16_csa_component_out[27];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[28] = s_CSAwallace_cska24_csa16_csa_component_out[28];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[29] = s_CSAwallace_cska24_csa16_csa_component_out[29];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[30] = s_CSAwallace_cska24_csa16_csa_component_out[30];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[31] = s_CSAwallace_cska24_csa16_csa_component_out[31];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[32] = s_CSAwallace_cska24_csa16_csa_component_out[32];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[33] = s_CSAwallace_cska24_csa16_csa_component_out[33];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[34] = s_CSAwallace_cska24_csa16_csa_component_out[34];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[35] = s_CSAwallace_cska24_csa16_csa_component_out[35];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[36] = s_CSAwallace_cska24_csa16_csa_component_out[36];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[37] = s_CSAwallace_cska24_csa16_csa_component_out[37];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[38] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[39] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[40] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[41] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[42] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[43] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[44] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[45] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[46] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17[47] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[0] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[1] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[2] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[3] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[4] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[5] = s_CSAwallace_cska24_csa16_csa_component_out[47];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[6] = s_CSAwallace_cska24_csa16_csa_component_out[48];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[7] = s_CSAwallace_cska24_csa16_csa_component_out[49];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[8] = s_CSAwallace_cska24_csa16_csa_component_out[50];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[9] = s_CSAwallace_cska24_csa16_csa_component_out[51];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[10] = s_CSAwallace_cska24_csa16_csa_component_out[52];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[11] = s_CSAwallace_cska24_csa16_csa_component_out[53];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[12] = s_CSAwallace_cska24_csa16_csa_component_out[54];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[13] = s_CSAwallace_cska24_csa16_csa_component_out[55];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[14] = s_CSAwallace_cska24_csa16_csa_component_out[56];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[15] = s_CSAwallace_cska24_csa16_csa_component_out[57];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[16] = s_CSAwallace_cska24_csa16_csa_component_out[58];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[17] = s_CSAwallace_cska24_csa16_csa_component_out[59];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[18] = s_CSAwallace_cska24_csa16_csa_component_out[60];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[19] = s_CSAwallace_cska24_csa16_csa_component_out[61];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[20] = s_CSAwallace_cska24_csa16_csa_component_out[62];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[21] = s_CSAwallace_cska24_csa16_csa_component_out[63];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[22] = s_CSAwallace_cska24_csa16_csa_component_out[64];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[23] = s_CSAwallace_cska24_csa16_csa_component_out[65];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[24] = s_CSAwallace_cska24_csa16_csa_component_out[66];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[25] = s_CSAwallace_cska24_csa16_csa_component_out[67];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[26] = s_CSAwallace_cska24_csa16_csa_component_out[68];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[27] = s_CSAwallace_cska24_csa16_csa_component_out[69];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[28] = s_CSAwallace_cska24_csa16_csa_component_out[70];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[29] = s_CSAwallace_cska24_csa16_csa_component_out[71];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[30] = s_CSAwallace_cska24_csa16_csa_component_out[72];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[31] = s_CSAwallace_cska24_csa16_csa_component_out[73];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[32] = s_CSAwallace_cska24_csa16_csa_component_out[74];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[33] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[34] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[35] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[36] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[37] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[38] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[39] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[40] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[41] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[42] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[43] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[44] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[45] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[46] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17[47] = 1'b1;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[0] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[1] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[2] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[3] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[4] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[5] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[6] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[7] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[8] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[9] = 1'b0;
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[10] = s_CSAwallace_cska24_csa17_csa_component_out[10];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[11] = s_CSAwallace_cska24_csa17_csa_component_out[11];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[12] = s_CSAwallace_cska24_csa17_csa_component_out[12];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[13] = s_CSAwallace_cska24_csa17_csa_component_out[13];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[14] = s_CSAwallace_cska24_csa17_csa_component_out[14];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[15] = s_CSAwallace_cska24_csa17_csa_component_out[15];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[16] = s_CSAwallace_cska24_csa17_csa_component_out[16];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[17] = s_CSAwallace_cska24_csa17_csa_component_out[17];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[18] = s_CSAwallace_cska24_csa17_csa_component_out[18];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[19] = s_CSAwallace_cska24_csa17_csa_component_out[19];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[20] = s_CSAwallace_cska24_csa17_csa_component_out[20];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[21] = s_CSAwallace_cska24_csa17_csa_component_out[21];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[22] = s_CSAwallace_cska24_csa17_csa_component_out[22];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[23] = s_CSAwallace_cska24_csa17_csa_component_out[23];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[24] = s_CSAwallace_cska24_csa17_csa_component_out[24];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[25] = s_CSAwallace_cska24_csa17_csa_component_out[25];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[26] = s_CSAwallace_cska24_csa17_csa_component_out[26];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[27] = s_CSAwallace_cska24_csa17_csa_component_out[27];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[28] = s_CSAwallace_cska24_csa17_csa_component_out[28];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[29] = s_CSAwallace_cska24_csa17_csa_component_out[29];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[30] = s_CSAwallace_cska24_csa17_csa_component_out[30];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[31] = s_CSAwallace_cska24_csa17_csa_component_out[31];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[32] = s_CSAwallace_cska24_csa17_csa_component_out[32];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[33] = s_CSAwallace_cska24_csa17_csa_component_out[33];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[34] = s_CSAwallace_cska24_csa17_csa_component_out[34];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[35] = s_CSAwallace_cska24_csa17_csa_component_out[35];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[36] = s_CSAwallace_cska24_csa17_csa_component_out[36];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[37] = s_CSAwallace_cska24_csa17_csa_component_out[37];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[38] = s_CSAwallace_cska24_csa17_csa_component_out[38];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[39] = s_CSAwallace_cska24_csa17_csa_component_out[39];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[40] = s_CSAwallace_cska24_csa17_csa_component_out[40];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[41] = s_CSAwallace_cska24_csa17_csa_component_out[41];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[42] = s_CSAwallace_cska24_csa17_csa_component_out[42];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[43] = s_CSAwallace_cska24_csa17_csa_component_out[43];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[44] = s_CSAwallace_cska24_csa17_csa_component_out[44];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[45] = s_CSAwallace_cska24_csa17_csa_component_out[45];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[46] = s_CSAwallace_cska24_csa17_csa_component_out[46];
  assign s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18[47] = 1'b1;
  csa_component48 csa_component48_s_CSAwallace_cska24_csa18_csa_component_out(.a(s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s17), .b(s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_c17), .c(s_CSAwallace_cska24_csa18_csa_component_s_CSAwallace_cska24_csa_s18), .csa_component48_out(s_CSAwallace_cska24_csa18_csa_component_out));
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[0] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[1] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[2] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[3] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[4] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[5] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[6] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[7] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[8] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[9] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[10] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[11] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[12] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[13] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[14] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[15] = s_CSAwallace_cska24_csa17_csa_component_out[64];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[16] = s_CSAwallace_cska24_csa17_csa_component_out[65];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[17] = s_CSAwallace_cska24_csa17_csa_component_out[66];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[18] = s_CSAwallace_cska24_csa17_csa_component_out[67];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[19] = s_CSAwallace_cska24_csa17_csa_component_out[68];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[20] = s_CSAwallace_cska24_csa17_csa_component_out[69];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[21] = s_CSAwallace_cska24_csa17_csa_component_out[70];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[22] = s_CSAwallace_cska24_csa17_csa_component_out[71];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[23] = s_CSAwallace_cska24_csa17_csa_component_out[72];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[24] = s_CSAwallace_cska24_csa17_csa_component_out[73];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[25] = s_CSAwallace_cska24_csa17_csa_component_out[74];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[26] = s_CSAwallace_cska24_csa17_csa_component_out[75];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[27] = s_CSAwallace_cska24_csa17_csa_component_out[76];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[28] = s_CSAwallace_cska24_csa17_csa_component_out[77];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[29] = s_CSAwallace_cska24_csa17_csa_component_out[78];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[30] = s_CSAwallace_cska24_csa17_csa_component_out[79];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[31] = s_CSAwallace_cska24_csa17_csa_component_out[80];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[32] = s_CSAwallace_cska24_csa17_csa_component_out[81];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[33] = s_CSAwallace_cska24_csa17_csa_component_out[82];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[34] = s_CSAwallace_cska24_csa17_csa_component_out[83];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[35] = s_CSAwallace_cska24_csa17_csa_component_out[84];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[36] = s_CSAwallace_cska24_csa17_csa_component_out[85];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[37] = s_CSAwallace_cska24_csa17_csa_component_out[86];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[38] = s_CSAwallace_cska24_csa17_csa_component_out[87];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[39] = s_CSAwallace_cska24_csa17_csa_component_out[88];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[40] = s_CSAwallace_cska24_csa17_csa_component_out[89];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[41] = s_CSAwallace_cska24_csa17_csa_component_out[90];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[42] = s_CSAwallace_cska24_csa17_csa_component_out[91];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[43] = s_CSAwallace_cska24_csa17_csa_component_out[92];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[44] = s_CSAwallace_cska24_csa17_csa_component_out[93];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[45] = s_CSAwallace_cska24_csa17_csa_component_out[94];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[46] = s_CSAwallace_cska24_csa17_csa_component_out[95];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18[47] = s_CSAwallace_cska24_csa17_csa_component_out[96];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[0] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[1] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[2] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[3] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[4] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[5] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[6] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[7] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[8] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[9] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[10] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[11] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[12] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[13] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[14] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[15] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[16] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[17] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[18] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[19] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[20] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[21] = s_CSAwallace_cska24_csa12_csa_component_out[70];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[22] = s_CSAwallace_cska24_csa12_csa_component_out[71];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[23] = s_CSAwallace_cska24_csa12_csa_component_out[72];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[24] = s_CSAwallace_cska24_csa12_csa_component_out[73];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[25] = s_CSAwallace_cska24_csa12_csa_component_out[74];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[26] = s_CSAwallace_cska24_csa12_csa_component_out[75];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[27] = s_CSAwallace_cska24_csa12_csa_component_out[76];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[28] = s_CSAwallace_cska24_csa12_csa_component_out[77];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[29] = s_CSAwallace_cska24_csa12_csa_component_out[78];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[30] = s_CSAwallace_cska24_csa12_csa_component_out[79];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[31] = s_CSAwallace_cska24_csa12_csa_component_out[80];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[32] = s_CSAwallace_cska24_csa12_csa_component_out[81];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[33] = s_CSAwallace_cska24_csa12_csa_component_out[82];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[34] = s_CSAwallace_cska24_csa12_csa_component_out[83];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[35] = s_CSAwallace_cska24_csa12_csa_component_out[84];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[36] = s_CSAwallace_cska24_csa12_csa_component_out[85];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[37] = s_CSAwallace_cska24_csa12_csa_component_out[86];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[38] = s_CSAwallace_cska24_csa12_csa_component_out[87];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[39] = s_CSAwallace_cska24_csa12_csa_component_out[88];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[40] = s_CSAwallace_cska24_csa12_csa_component_out[89];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[41] = s_CSAwallace_cska24_csa12_csa_component_out[90];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[42] = s_CSAwallace_cska24_csa12_csa_component_out[91];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[43] = s_CSAwallace_cska24_csa12_csa_component_out[92];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[44] = s_CSAwallace_cska24_csa12_csa_component_out[93];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[45] = 1'b1;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[46] = 1'b1;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13[47] = 1'b1;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[0] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[1] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[2] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[3] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[4] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[5] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[6] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[7] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[8] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[9] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[10] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[11] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[12] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[13] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[14] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[15] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[16] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[17] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[18] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[19] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[20] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[21] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[22] = 1'b0;
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[23] = s_CSAwallace_cska24_csa7_csa_component_out[71];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[24] = s_CSAwallace_cska24_csa7_csa_component_out[72];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[25] = s_CSAwallace_cska24_csa7_csa_component_out[73];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[26] = s_CSAwallace_cska24_csa7_csa_component_out[74];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[27] = s_CSAwallace_cska24_csa7_csa_component_out[75];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[28] = s_CSAwallace_cska24_csa7_csa_component_out[76];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[29] = s_CSAwallace_cska24_csa7_csa_component_out[77];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[30] = s_CSAwallace_cska24_csa7_csa_component_out[78];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[31] = s_CSAwallace_cska24_csa7_csa_component_out[79];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[32] = s_CSAwallace_cska24_csa7_csa_component_out[80];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[33] = s_CSAwallace_cska24_csa7_csa_component_out[81];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[34] = s_CSAwallace_cska24_csa7_csa_component_out[82];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[35] = s_CSAwallace_cska24_csa7_csa_component_out[83];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[36] = s_CSAwallace_cska24_csa7_csa_component_out[84];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[37] = s_CSAwallace_cska24_csa7_csa_component_out[85];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[38] = s_CSAwallace_cska24_csa7_csa_component_out[86];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[39] = s_CSAwallace_cska24_csa7_csa_component_out[87];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[40] = s_CSAwallace_cska24_csa7_csa_component_out[88];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[41] = s_CSAwallace_cska24_csa7_csa_component_out[89];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[42] = s_CSAwallace_cska24_csa7_csa_component_out[90];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[43] = s_CSAwallace_cska24_csa7_csa_component_out[91];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[44] = s_CSAwallace_cska24_csa7_csa_component_out[92];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[45] = s_CSAwallace_cska24_csa7_csa_component_out[93];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[46] = s_CSAwallace_cska24_csa7_csa_component_out[94];
  assign s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8[47] = 1'b1;
  csa_component48 csa_component48_s_CSAwallace_cska24_csa19_csa_component_out(.a(s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c18), .b(s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c13), .c(s_CSAwallace_cska24_csa19_csa_component_s_CSAwallace_cska24_csa_c8), .csa_component48_out(s_CSAwallace_cska24_csa19_csa_component_out));
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[0] = s_CSAwallace_cska24_csa18_csa_component_out[0];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[1] = s_CSAwallace_cska24_csa18_csa_component_out[1];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[2] = s_CSAwallace_cska24_csa18_csa_component_out[2];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[3] = s_CSAwallace_cska24_csa18_csa_component_out[3];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[4] = s_CSAwallace_cska24_csa18_csa_component_out[4];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[5] = s_CSAwallace_cska24_csa18_csa_component_out[5];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[6] = s_CSAwallace_cska24_csa18_csa_component_out[6];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[7] = s_CSAwallace_cska24_csa18_csa_component_out[7];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[8] = s_CSAwallace_cska24_csa18_csa_component_out[8];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[9] = s_CSAwallace_cska24_csa18_csa_component_out[9];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[10] = s_CSAwallace_cska24_csa18_csa_component_out[10];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[11] = s_CSAwallace_cska24_csa18_csa_component_out[11];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[12] = s_CSAwallace_cska24_csa18_csa_component_out[12];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[13] = s_CSAwallace_cska24_csa18_csa_component_out[13];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[14] = s_CSAwallace_cska24_csa18_csa_component_out[14];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[15] = s_CSAwallace_cska24_csa18_csa_component_out[15];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[16] = s_CSAwallace_cska24_csa18_csa_component_out[16];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[17] = s_CSAwallace_cska24_csa18_csa_component_out[17];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[18] = s_CSAwallace_cska24_csa18_csa_component_out[18];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[19] = s_CSAwallace_cska24_csa18_csa_component_out[19];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[20] = s_CSAwallace_cska24_csa18_csa_component_out[20];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[21] = s_CSAwallace_cska24_csa18_csa_component_out[21];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[22] = s_CSAwallace_cska24_csa18_csa_component_out[22];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[23] = s_CSAwallace_cska24_csa18_csa_component_out[23];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[24] = s_CSAwallace_cska24_csa18_csa_component_out[24];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[25] = s_CSAwallace_cska24_csa18_csa_component_out[25];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[26] = s_CSAwallace_cska24_csa18_csa_component_out[26];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[27] = s_CSAwallace_cska24_csa18_csa_component_out[27];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[28] = s_CSAwallace_cska24_csa18_csa_component_out[28];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[29] = s_CSAwallace_cska24_csa18_csa_component_out[29];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[30] = s_CSAwallace_cska24_csa18_csa_component_out[30];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[31] = s_CSAwallace_cska24_csa18_csa_component_out[31];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[32] = s_CSAwallace_cska24_csa18_csa_component_out[32];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[33] = s_CSAwallace_cska24_csa18_csa_component_out[33];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[34] = s_CSAwallace_cska24_csa18_csa_component_out[34];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[35] = s_CSAwallace_cska24_csa18_csa_component_out[35];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[36] = s_CSAwallace_cska24_csa18_csa_component_out[36];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[37] = s_CSAwallace_cska24_csa18_csa_component_out[37];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[38] = s_CSAwallace_cska24_csa18_csa_component_out[38];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[39] = s_CSAwallace_cska24_csa18_csa_component_out[39];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[40] = s_CSAwallace_cska24_csa18_csa_component_out[40];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[41] = s_CSAwallace_cska24_csa18_csa_component_out[41];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[42] = s_CSAwallace_cska24_csa18_csa_component_out[42];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[43] = s_CSAwallace_cska24_csa18_csa_component_out[43];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[44] = s_CSAwallace_cska24_csa18_csa_component_out[44];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[45] = s_CSAwallace_cska24_csa18_csa_component_out[45];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[46] = s_CSAwallace_cska24_csa18_csa_component_out[46];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19[47] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[0] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[1] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[2] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[3] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[4] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[5] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[6] = s_CSAwallace_cska24_csa18_csa_component_out[55];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[7] = s_CSAwallace_cska24_csa18_csa_component_out[56];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[8] = s_CSAwallace_cska24_csa18_csa_component_out[57];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[9] = s_CSAwallace_cska24_csa18_csa_component_out[58];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[10] = s_CSAwallace_cska24_csa18_csa_component_out[59];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[11] = s_CSAwallace_cska24_csa18_csa_component_out[60];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[12] = s_CSAwallace_cska24_csa18_csa_component_out[61];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[13] = s_CSAwallace_cska24_csa18_csa_component_out[62];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[14] = s_CSAwallace_cska24_csa18_csa_component_out[63];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[15] = s_CSAwallace_cska24_csa18_csa_component_out[64];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[16] = s_CSAwallace_cska24_csa18_csa_component_out[65];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[17] = s_CSAwallace_cska24_csa18_csa_component_out[66];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[18] = s_CSAwallace_cska24_csa18_csa_component_out[67];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[19] = s_CSAwallace_cska24_csa18_csa_component_out[68];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[20] = s_CSAwallace_cska24_csa18_csa_component_out[69];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[21] = s_CSAwallace_cska24_csa18_csa_component_out[70];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[22] = s_CSAwallace_cska24_csa18_csa_component_out[71];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[23] = s_CSAwallace_cska24_csa18_csa_component_out[72];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[24] = s_CSAwallace_cska24_csa18_csa_component_out[73];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[25] = s_CSAwallace_cska24_csa18_csa_component_out[74];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[26] = s_CSAwallace_cska24_csa18_csa_component_out[75];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[27] = s_CSAwallace_cska24_csa18_csa_component_out[76];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[28] = s_CSAwallace_cska24_csa18_csa_component_out[77];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[29] = s_CSAwallace_cska24_csa18_csa_component_out[78];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[30] = s_CSAwallace_cska24_csa18_csa_component_out[79];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[31] = s_CSAwallace_cska24_csa18_csa_component_out[80];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[32] = s_CSAwallace_cska24_csa18_csa_component_out[81];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[33] = s_CSAwallace_cska24_csa18_csa_component_out[82];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[34] = s_CSAwallace_cska24_csa18_csa_component_out[83];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[35] = s_CSAwallace_cska24_csa18_csa_component_out[84];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[36] = s_CSAwallace_cska24_csa18_csa_component_out[85];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[37] = s_CSAwallace_cska24_csa18_csa_component_out[86];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[38] = s_CSAwallace_cska24_csa18_csa_component_out[87];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[39] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[40] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[41] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[42] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[43] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[44] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[45] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[46] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19[47] = 1'b1;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[0] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[1] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[2] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[3] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[4] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[5] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[6] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[7] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[8] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[9] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[10] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[11] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[12] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[13] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[14] = 1'b0;
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[15] = s_CSAwallace_cska24_csa19_csa_component_out[15];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[16] = s_CSAwallace_cska24_csa19_csa_component_out[16];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[17] = s_CSAwallace_cska24_csa19_csa_component_out[17];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[18] = s_CSAwallace_cska24_csa19_csa_component_out[18];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[19] = s_CSAwallace_cska24_csa19_csa_component_out[19];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[20] = s_CSAwallace_cska24_csa19_csa_component_out[20];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[21] = s_CSAwallace_cska24_csa19_csa_component_out[21];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[22] = s_CSAwallace_cska24_csa19_csa_component_out[22];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[23] = s_CSAwallace_cska24_csa19_csa_component_out[23];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[24] = s_CSAwallace_cska24_csa19_csa_component_out[24];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[25] = s_CSAwallace_cska24_csa19_csa_component_out[25];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[26] = s_CSAwallace_cska24_csa19_csa_component_out[26];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[27] = s_CSAwallace_cska24_csa19_csa_component_out[27];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[28] = s_CSAwallace_cska24_csa19_csa_component_out[28];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[29] = s_CSAwallace_cska24_csa19_csa_component_out[29];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[30] = s_CSAwallace_cska24_csa19_csa_component_out[30];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[31] = s_CSAwallace_cska24_csa19_csa_component_out[31];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[32] = s_CSAwallace_cska24_csa19_csa_component_out[32];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[33] = s_CSAwallace_cska24_csa19_csa_component_out[33];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[34] = s_CSAwallace_cska24_csa19_csa_component_out[34];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[35] = s_CSAwallace_cska24_csa19_csa_component_out[35];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[36] = s_CSAwallace_cska24_csa19_csa_component_out[36];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[37] = s_CSAwallace_cska24_csa19_csa_component_out[37];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[38] = s_CSAwallace_cska24_csa19_csa_component_out[38];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[39] = s_CSAwallace_cska24_csa19_csa_component_out[39];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[40] = s_CSAwallace_cska24_csa19_csa_component_out[40];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[41] = s_CSAwallace_cska24_csa19_csa_component_out[41];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[42] = s_CSAwallace_cska24_csa19_csa_component_out[42];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[43] = s_CSAwallace_cska24_csa19_csa_component_out[43];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[44] = s_CSAwallace_cska24_csa19_csa_component_out[44];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[45] = s_CSAwallace_cska24_csa19_csa_component_out[45];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[46] = s_CSAwallace_cska24_csa19_csa_component_out[46];
  assign s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20[47] = s_CSAwallace_cska24_csa19_csa_component_out[47];
  csa_component48 csa_component48_s_CSAwallace_cska24_csa20_csa_component_out(.a(s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s19), .b(s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_c19), .c(s_CSAwallace_cska24_csa20_csa_component_s_CSAwallace_cska24_csa_s20), .csa_component48_out(s_CSAwallace_cska24_csa20_csa_component_out));
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[0] = s_CSAwallace_cska24_csa20_csa_component_out[0];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[1] = s_CSAwallace_cska24_csa20_csa_component_out[1];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[2] = s_CSAwallace_cska24_csa20_csa_component_out[2];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[3] = s_CSAwallace_cska24_csa20_csa_component_out[3];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[4] = s_CSAwallace_cska24_csa20_csa_component_out[4];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[5] = s_CSAwallace_cska24_csa20_csa_component_out[5];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[6] = s_CSAwallace_cska24_csa20_csa_component_out[6];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[7] = s_CSAwallace_cska24_csa20_csa_component_out[7];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[8] = s_CSAwallace_cska24_csa20_csa_component_out[8];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[9] = s_CSAwallace_cska24_csa20_csa_component_out[9];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[10] = s_CSAwallace_cska24_csa20_csa_component_out[10];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[11] = s_CSAwallace_cska24_csa20_csa_component_out[11];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[12] = s_CSAwallace_cska24_csa20_csa_component_out[12];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[13] = s_CSAwallace_cska24_csa20_csa_component_out[13];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[14] = s_CSAwallace_cska24_csa20_csa_component_out[14];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[15] = s_CSAwallace_cska24_csa20_csa_component_out[15];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[16] = s_CSAwallace_cska24_csa20_csa_component_out[16];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[17] = s_CSAwallace_cska24_csa20_csa_component_out[17];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[18] = s_CSAwallace_cska24_csa20_csa_component_out[18];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[19] = s_CSAwallace_cska24_csa20_csa_component_out[19];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[20] = s_CSAwallace_cska24_csa20_csa_component_out[20];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[21] = s_CSAwallace_cska24_csa20_csa_component_out[21];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[22] = s_CSAwallace_cska24_csa20_csa_component_out[22];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[23] = s_CSAwallace_cska24_csa20_csa_component_out[23];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[24] = s_CSAwallace_cska24_csa20_csa_component_out[24];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[25] = s_CSAwallace_cska24_csa20_csa_component_out[25];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[26] = s_CSAwallace_cska24_csa20_csa_component_out[26];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[27] = s_CSAwallace_cska24_csa20_csa_component_out[27];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[28] = s_CSAwallace_cska24_csa20_csa_component_out[28];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[29] = s_CSAwallace_cska24_csa20_csa_component_out[29];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[30] = s_CSAwallace_cska24_csa20_csa_component_out[30];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[31] = s_CSAwallace_cska24_csa20_csa_component_out[31];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[32] = s_CSAwallace_cska24_csa20_csa_component_out[32];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[33] = s_CSAwallace_cska24_csa20_csa_component_out[33];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[34] = s_CSAwallace_cska24_csa20_csa_component_out[34];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[35] = s_CSAwallace_cska24_csa20_csa_component_out[35];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[36] = s_CSAwallace_cska24_csa20_csa_component_out[36];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[37] = s_CSAwallace_cska24_csa20_csa_component_out[37];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[38] = s_CSAwallace_cska24_csa20_csa_component_out[38];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[39] = s_CSAwallace_cska24_csa20_csa_component_out[39];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[40] = s_CSAwallace_cska24_csa20_csa_component_out[40];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[41] = s_CSAwallace_cska24_csa20_csa_component_out[41];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[42] = s_CSAwallace_cska24_csa20_csa_component_out[42];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[43] = s_CSAwallace_cska24_csa20_csa_component_out[43];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[44] = s_CSAwallace_cska24_csa20_csa_component_out[44];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[45] = s_CSAwallace_cska24_csa20_csa_component_out[45];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[46] = s_CSAwallace_cska24_csa20_csa_component_out[46];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21[47] = s_CSAwallace_cska24_csa20_csa_component_out[47];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[0] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[1] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[2] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[3] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[4] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[5] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[6] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[7] = s_CSAwallace_cska24_csa20_csa_component_out[56];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[8] = s_CSAwallace_cska24_csa20_csa_component_out[57];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[9] = s_CSAwallace_cska24_csa20_csa_component_out[58];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[10] = s_CSAwallace_cska24_csa20_csa_component_out[59];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[11] = s_CSAwallace_cska24_csa20_csa_component_out[60];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[12] = s_CSAwallace_cska24_csa20_csa_component_out[61];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[13] = s_CSAwallace_cska24_csa20_csa_component_out[62];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[14] = s_CSAwallace_cska24_csa20_csa_component_out[63];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[15] = s_CSAwallace_cska24_csa20_csa_component_out[64];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[16] = s_CSAwallace_cska24_csa20_csa_component_out[65];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[17] = s_CSAwallace_cska24_csa20_csa_component_out[66];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[18] = s_CSAwallace_cska24_csa20_csa_component_out[67];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[19] = s_CSAwallace_cska24_csa20_csa_component_out[68];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[20] = s_CSAwallace_cska24_csa20_csa_component_out[69];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[21] = s_CSAwallace_cska24_csa20_csa_component_out[70];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[22] = s_CSAwallace_cska24_csa20_csa_component_out[71];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[23] = s_CSAwallace_cska24_csa20_csa_component_out[72];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[24] = s_CSAwallace_cska24_csa20_csa_component_out[73];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[25] = s_CSAwallace_cska24_csa20_csa_component_out[74];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[26] = s_CSAwallace_cska24_csa20_csa_component_out[75];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[27] = s_CSAwallace_cska24_csa20_csa_component_out[76];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[28] = s_CSAwallace_cska24_csa20_csa_component_out[77];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[29] = s_CSAwallace_cska24_csa20_csa_component_out[78];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[30] = s_CSAwallace_cska24_csa20_csa_component_out[79];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[31] = s_CSAwallace_cska24_csa20_csa_component_out[80];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[32] = s_CSAwallace_cska24_csa20_csa_component_out[81];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[33] = s_CSAwallace_cska24_csa20_csa_component_out[82];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[34] = s_CSAwallace_cska24_csa20_csa_component_out[83];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[35] = s_CSAwallace_cska24_csa20_csa_component_out[84];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[36] = s_CSAwallace_cska24_csa20_csa_component_out[85];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[37] = s_CSAwallace_cska24_csa20_csa_component_out[86];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[38] = s_CSAwallace_cska24_csa20_csa_component_out[87];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[39] = s_CSAwallace_cska24_csa20_csa_component_out[88];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[40] = s_CSAwallace_cska24_csa20_csa_component_out[89];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[41] = s_CSAwallace_cska24_csa20_csa_component_out[90];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[42] = s_CSAwallace_cska24_csa20_csa_component_out[91];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[43] = s_CSAwallace_cska24_csa20_csa_component_out[92];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[44] = s_CSAwallace_cska24_csa20_csa_component_out[93];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[45] = s_CSAwallace_cska24_csa20_csa_component_out[94];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[46] = s_CSAwallace_cska24_csa20_csa_component_out[95];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21[47] = s_CSAwallace_cska24_csa20_csa_component_out[96];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[0] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[1] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[2] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[3] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[4] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[5] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[6] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[7] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[8] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[9] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[10] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[11] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[12] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[13] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[14] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[15] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[16] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[17] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[18] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[19] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[20] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[21] = 1'b0;
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[22] = s_CSAwallace_cska24_csa19_csa_component_out[71];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[23] = s_CSAwallace_cska24_csa19_csa_component_out[72];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[24] = s_CSAwallace_cska24_csa19_csa_component_out[73];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[25] = s_CSAwallace_cska24_csa19_csa_component_out[74];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[26] = s_CSAwallace_cska24_csa19_csa_component_out[75];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[27] = s_CSAwallace_cska24_csa19_csa_component_out[76];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[28] = s_CSAwallace_cska24_csa19_csa_component_out[77];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[29] = s_CSAwallace_cska24_csa19_csa_component_out[78];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[30] = s_CSAwallace_cska24_csa19_csa_component_out[79];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[31] = s_CSAwallace_cska24_csa19_csa_component_out[80];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[32] = s_CSAwallace_cska24_csa19_csa_component_out[81];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[33] = s_CSAwallace_cska24_csa19_csa_component_out[82];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[34] = s_CSAwallace_cska24_csa19_csa_component_out[83];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[35] = s_CSAwallace_cska24_csa19_csa_component_out[84];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[36] = s_CSAwallace_cska24_csa19_csa_component_out[85];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[37] = s_CSAwallace_cska24_csa19_csa_component_out[86];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[38] = s_CSAwallace_cska24_csa19_csa_component_out[87];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[39] = s_CSAwallace_cska24_csa19_csa_component_out[88];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[40] = s_CSAwallace_cska24_csa19_csa_component_out[89];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[41] = s_CSAwallace_cska24_csa19_csa_component_out[90];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[42] = s_CSAwallace_cska24_csa19_csa_component_out[91];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[43] = s_CSAwallace_cska24_csa19_csa_component_out[92];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[44] = s_CSAwallace_cska24_csa19_csa_component_out[93];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[45] = s_CSAwallace_cska24_csa19_csa_component_out[94];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[46] = s_CSAwallace_cska24_csa19_csa_component_out[95];
  assign s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20[47] = s_CSAwallace_cska24_csa19_csa_component_out[96];
  csa_component48 csa_component48_s_CSAwallace_cska24_csa21_csa_component_out(.a(s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_s21), .b(s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c21), .c(s_CSAwallace_cska24_csa21_csa_component_s_CSAwallace_cska24_csa_c20), .csa_component48_out(s_CSAwallace_cska24_csa21_csa_component_out));
  assign s_CSAwallace_cska24_u_cska48_a[0] = s_CSAwallace_cska24_csa21_csa_component_out[0];
  assign s_CSAwallace_cska24_u_cska48_a[1] = s_CSAwallace_cska24_csa21_csa_component_out[1];
  assign s_CSAwallace_cska24_u_cska48_a[2] = s_CSAwallace_cska24_csa21_csa_component_out[2];
  assign s_CSAwallace_cska24_u_cska48_a[3] = s_CSAwallace_cska24_csa21_csa_component_out[3];
  assign s_CSAwallace_cska24_u_cska48_a[4] = s_CSAwallace_cska24_csa21_csa_component_out[4];
  assign s_CSAwallace_cska24_u_cska48_a[5] = s_CSAwallace_cska24_csa21_csa_component_out[5];
  assign s_CSAwallace_cska24_u_cska48_a[6] = s_CSAwallace_cska24_csa21_csa_component_out[6];
  assign s_CSAwallace_cska24_u_cska48_a[7] = s_CSAwallace_cska24_csa21_csa_component_out[7];
  assign s_CSAwallace_cska24_u_cska48_a[8] = s_CSAwallace_cska24_csa21_csa_component_out[8];
  assign s_CSAwallace_cska24_u_cska48_a[9] = s_CSAwallace_cska24_csa21_csa_component_out[9];
  assign s_CSAwallace_cska24_u_cska48_a[10] = s_CSAwallace_cska24_csa21_csa_component_out[10];
  assign s_CSAwallace_cska24_u_cska48_a[11] = s_CSAwallace_cska24_csa21_csa_component_out[11];
  assign s_CSAwallace_cska24_u_cska48_a[12] = s_CSAwallace_cska24_csa21_csa_component_out[12];
  assign s_CSAwallace_cska24_u_cska48_a[13] = s_CSAwallace_cska24_csa21_csa_component_out[13];
  assign s_CSAwallace_cska24_u_cska48_a[14] = s_CSAwallace_cska24_csa21_csa_component_out[14];
  assign s_CSAwallace_cska24_u_cska48_a[15] = s_CSAwallace_cska24_csa21_csa_component_out[15];
  assign s_CSAwallace_cska24_u_cska48_a[16] = s_CSAwallace_cska24_csa21_csa_component_out[16];
  assign s_CSAwallace_cska24_u_cska48_a[17] = s_CSAwallace_cska24_csa21_csa_component_out[17];
  assign s_CSAwallace_cska24_u_cska48_a[18] = s_CSAwallace_cska24_csa21_csa_component_out[18];
  assign s_CSAwallace_cska24_u_cska48_a[19] = s_CSAwallace_cska24_csa21_csa_component_out[19];
  assign s_CSAwallace_cska24_u_cska48_a[20] = s_CSAwallace_cska24_csa21_csa_component_out[20];
  assign s_CSAwallace_cska24_u_cska48_a[21] = s_CSAwallace_cska24_csa21_csa_component_out[21];
  assign s_CSAwallace_cska24_u_cska48_a[22] = s_CSAwallace_cska24_csa21_csa_component_out[22];
  assign s_CSAwallace_cska24_u_cska48_a[23] = s_CSAwallace_cska24_csa21_csa_component_out[23];
  assign s_CSAwallace_cska24_u_cska48_a[24] = s_CSAwallace_cska24_csa21_csa_component_out[24];
  assign s_CSAwallace_cska24_u_cska48_a[25] = s_CSAwallace_cska24_csa21_csa_component_out[25];
  assign s_CSAwallace_cska24_u_cska48_a[26] = s_CSAwallace_cska24_csa21_csa_component_out[26];
  assign s_CSAwallace_cska24_u_cska48_a[27] = s_CSAwallace_cska24_csa21_csa_component_out[27];
  assign s_CSAwallace_cska24_u_cska48_a[28] = s_CSAwallace_cska24_csa21_csa_component_out[28];
  assign s_CSAwallace_cska24_u_cska48_a[29] = s_CSAwallace_cska24_csa21_csa_component_out[29];
  assign s_CSAwallace_cska24_u_cska48_a[30] = s_CSAwallace_cska24_csa21_csa_component_out[30];
  assign s_CSAwallace_cska24_u_cska48_a[31] = s_CSAwallace_cska24_csa21_csa_component_out[31];
  assign s_CSAwallace_cska24_u_cska48_a[32] = s_CSAwallace_cska24_csa21_csa_component_out[32];
  assign s_CSAwallace_cska24_u_cska48_a[33] = s_CSAwallace_cska24_csa21_csa_component_out[33];
  assign s_CSAwallace_cska24_u_cska48_a[34] = s_CSAwallace_cska24_csa21_csa_component_out[34];
  assign s_CSAwallace_cska24_u_cska48_a[35] = s_CSAwallace_cska24_csa21_csa_component_out[35];
  assign s_CSAwallace_cska24_u_cska48_a[36] = s_CSAwallace_cska24_csa21_csa_component_out[36];
  assign s_CSAwallace_cska24_u_cska48_a[37] = s_CSAwallace_cska24_csa21_csa_component_out[37];
  assign s_CSAwallace_cska24_u_cska48_a[38] = s_CSAwallace_cska24_csa21_csa_component_out[38];
  assign s_CSAwallace_cska24_u_cska48_a[39] = s_CSAwallace_cska24_csa21_csa_component_out[39];
  assign s_CSAwallace_cska24_u_cska48_a[40] = s_CSAwallace_cska24_csa21_csa_component_out[40];
  assign s_CSAwallace_cska24_u_cska48_a[41] = s_CSAwallace_cska24_csa21_csa_component_out[41];
  assign s_CSAwallace_cska24_u_cska48_a[42] = s_CSAwallace_cska24_csa21_csa_component_out[42];
  assign s_CSAwallace_cska24_u_cska48_a[43] = s_CSAwallace_cska24_csa21_csa_component_out[43];
  assign s_CSAwallace_cska24_u_cska48_a[44] = s_CSAwallace_cska24_csa21_csa_component_out[44];
  assign s_CSAwallace_cska24_u_cska48_a[45] = s_CSAwallace_cska24_csa21_csa_component_out[45];
  assign s_CSAwallace_cska24_u_cska48_a[46] = s_CSAwallace_cska24_csa21_csa_component_out[46];
  assign s_CSAwallace_cska24_u_cska48_a[47] = s_CSAwallace_cska24_csa21_csa_component_out[47];
  assign s_CSAwallace_cska24_u_cska48_b[0] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[1] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[2] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[3] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[4] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[5] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[6] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[7] = 1'b0;
  assign s_CSAwallace_cska24_u_cska48_b[8] = s_CSAwallace_cska24_csa21_csa_component_out[57];
  assign s_CSAwallace_cska24_u_cska48_b[9] = s_CSAwallace_cska24_csa21_csa_component_out[58];
  assign s_CSAwallace_cska24_u_cska48_b[10] = s_CSAwallace_cska24_csa21_csa_component_out[59];
  assign s_CSAwallace_cska24_u_cska48_b[11] = s_CSAwallace_cska24_csa21_csa_component_out[60];
  assign s_CSAwallace_cska24_u_cska48_b[12] = s_CSAwallace_cska24_csa21_csa_component_out[61];
  assign s_CSAwallace_cska24_u_cska48_b[13] = s_CSAwallace_cska24_csa21_csa_component_out[62];
  assign s_CSAwallace_cska24_u_cska48_b[14] = s_CSAwallace_cska24_csa21_csa_component_out[63];
  assign s_CSAwallace_cska24_u_cska48_b[15] = s_CSAwallace_cska24_csa21_csa_component_out[64];
  assign s_CSAwallace_cska24_u_cska48_b[16] = s_CSAwallace_cska24_csa21_csa_component_out[65];
  assign s_CSAwallace_cska24_u_cska48_b[17] = s_CSAwallace_cska24_csa21_csa_component_out[66];
  assign s_CSAwallace_cska24_u_cska48_b[18] = s_CSAwallace_cska24_csa21_csa_component_out[67];
  assign s_CSAwallace_cska24_u_cska48_b[19] = s_CSAwallace_cska24_csa21_csa_component_out[68];
  assign s_CSAwallace_cska24_u_cska48_b[20] = s_CSAwallace_cska24_csa21_csa_component_out[69];
  assign s_CSAwallace_cska24_u_cska48_b[21] = s_CSAwallace_cska24_csa21_csa_component_out[70];
  assign s_CSAwallace_cska24_u_cska48_b[22] = s_CSAwallace_cska24_csa21_csa_component_out[71];
  assign s_CSAwallace_cska24_u_cska48_b[23] = s_CSAwallace_cska24_csa21_csa_component_out[72];
  assign s_CSAwallace_cska24_u_cska48_b[24] = s_CSAwallace_cska24_csa21_csa_component_out[73];
  assign s_CSAwallace_cska24_u_cska48_b[25] = s_CSAwallace_cska24_csa21_csa_component_out[74];
  assign s_CSAwallace_cska24_u_cska48_b[26] = s_CSAwallace_cska24_csa21_csa_component_out[75];
  assign s_CSAwallace_cska24_u_cska48_b[27] = s_CSAwallace_cska24_csa21_csa_component_out[76];
  assign s_CSAwallace_cska24_u_cska48_b[28] = s_CSAwallace_cska24_csa21_csa_component_out[77];
  assign s_CSAwallace_cska24_u_cska48_b[29] = s_CSAwallace_cska24_csa21_csa_component_out[78];
  assign s_CSAwallace_cska24_u_cska48_b[30] = s_CSAwallace_cska24_csa21_csa_component_out[79];
  assign s_CSAwallace_cska24_u_cska48_b[31] = s_CSAwallace_cska24_csa21_csa_component_out[80];
  assign s_CSAwallace_cska24_u_cska48_b[32] = s_CSAwallace_cska24_csa21_csa_component_out[81];
  assign s_CSAwallace_cska24_u_cska48_b[33] = s_CSAwallace_cska24_csa21_csa_component_out[82];
  assign s_CSAwallace_cska24_u_cska48_b[34] = s_CSAwallace_cska24_csa21_csa_component_out[83];
  assign s_CSAwallace_cska24_u_cska48_b[35] = s_CSAwallace_cska24_csa21_csa_component_out[84];
  assign s_CSAwallace_cska24_u_cska48_b[36] = s_CSAwallace_cska24_csa21_csa_component_out[85];
  assign s_CSAwallace_cska24_u_cska48_b[37] = s_CSAwallace_cska24_csa21_csa_component_out[86];
  assign s_CSAwallace_cska24_u_cska48_b[38] = s_CSAwallace_cska24_csa21_csa_component_out[87];
  assign s_CSAwallace_cska24_u_cska48_b[39] = s_CSAwallace_cska24_csa21_csa_component_out[88];
  assign s_CSAwallace_cska24_u_cska48_b[40] = s_CSAwallace_cska24_csa21_csa_component_out[89];
  assign s_CSAwallace_cska24_u_cska48_b[41] = s_CSAwallace_cska24_csa21_csa_component_out[90];
  assign s_CSAwallace_cska24_u_cska48_b[42] = s_CSAwallace_cska24_csa21_csa_component_out[91];
  assign s_CSAwallace_cska24_u_cska48_b[43] = s_CSAwallace_cska24_csa21_csa_component_out[92];
  assign s_CSAwallace_cska24_u_cska48_b[44] = s_CSAwallace_cska24_csa21_csa_component_out[93];
  assign s_CSAwallace_cska24_u_cska48_b[45] = s_CSAwallace_cska24_csa21_csa_component_out[94];
  assign s_CSAwallace_cska24_u_cska48_b[46] = s_CSAwallace_cska24_csa21_csa_component_out[95];
  assign s_CSAwallace_cska24_u_cska48_b[47] = s_CSAwallace_cska24_csa21_csa_component_out[96];
  u_cska48 u_cska48_s_CSAwallace_cska24_u_cska48_out(.a(s_CSAwallace_cska24_u_cska48_a), .b(s_CSAwallace_cska24_u_cska48_b), .u_cska48_out(s_CSAwallace_cska24_u_cska48_out));
  not_gate not_gate_s_CSAwallace_cska24_xor0(.a(s_CSAwallace_cska24_u_cska48_out[47]), .out(s_CSAwallace_cska24_xor0));

  assign s_CSAwallace_cska24_out[0] = s_CSAwallace_cska24_u_cska48_out[0];
  assign s_CSAwallace_cska24_out[1] = s_CSAwallace_cska24_u_cska48_out[1];
  assign s_CSAwallace_cska24_out[2] = s_CSAwallace_cska24_u_cska48_out[2];
  assign s_CSAwallace_cska24_out[3] = s_CSAwallace_cska24_u_cska48_out[3];
  assign s_CSAwallace_cska24_out[4] = s_CSAwallace_cska24_u_cska48_out[4];
  assign s_CSAwallace_cska24_out[5] = s_CSAwallace_cska24_u_cska48_out[5];
  assign s_CSAwallace_cska24_out[6] = s_CSAwallace_cska24_u_cska48_out[6];
  assign s_CSAwallace_cska24_out[7] = s_CSAwallace_cska24_u_cska48_out[7];
  assign s_CSAwallace_cska24_out[8] = s_CSAwallace_cska24_u_cska48_out[8];
  assign s_CSAwallace_cska24_out[9] = s_CSAwallace_cska24_u_cska48_out[9];
  assign s_CSAwallace_cska24_out[10] = s_CSAwallace_cska24_u_cska48_out[10];
  assign s_CSAwallace_cska24_out[11] = s_CSAwallace_cska24_u_cska48_out[11];
  assign s_CSAwallace_cska24_out[12] = s_CSAwallace_cska24_u_cska48_out[12];
  assign s_CSAwallace_cska24_out[13] = s_CSAwallace_cska24_u_cska48_out[13];
  assign s_CSAwallace_cska24_out[14] = s_CSAwallace_cska24_u_cska48_out[14];
  assign s_CSAwallace_cska24_out[15] = s_CSAwallace_cska24_u_cska48_out[15];
  assign s_CSAwallace_cska24_out[16] = s_CSAwallace_cska24_u_cska48_out[16];
  assign s_CSAwallace_cska24_out[17] = s_CSAwallace_cska24_u_cska48_out[17];
  assign s_CSAwallace_cska24_out[18] = s_CSAwallace_cska24_u_cska48_out[18];
  assign s_CSAwallace_cska24_out[19] = s_CSAwallace_cska24_u_cska48_out[19];
  assign s_CSAwallace_cska24_out[20] = s_CSAwallace_cska24_u_cska48_out[20];
  assign s_CSAwallace_cska24_out[21] = s_CSAwallace_cska24_u_cska48_out[21];
  assign s_CSAwallace_cska24_out[22] = s_CSAwallace_cska24_u_cska48_out[22];
  assign s_CSAwallace_cska24_out[23] = s_CSAwallace_cska24_u_cska48_out[23];
  assign s_CSAwallace_cska24_out[24] = s_CSAwallace_cska24_u_cska48_out[24];
  assign s_CSAwallace_cska24_out[25] = s_CSAwallace_cska24_u_cska48_out[25];
  assign s_CSAwallace_cska24_out[26] = s_CSAwallace_cska24_u_cska48_out[26];
  assign s_CSAwallace_cska24_out[27] = s_CSAwallace_cska24_u_cska48_out[27];
  assign s_CSAwallace_cska24_out[28] = s_CSAwallace_cska24_u_cska48_out[28];
  assign s_CSAwallace_cska24_out[29] = s_CSAwallace_cska24_u_cska48_out[29];
  assign s_CSAwallace_cska24_out[30] = s_CSAwallace_cska24_u_cska48_out[30];
  assign s_CSAwallace_cska24_out[31] = s_CSAwallace_cska24_u_cska48_out[31];
  assign s_CSAwallace_cska24_out[32] = s_CSAwallace_cska24_u_cska48_out[32];
  assign s_CSAwallace_cska24_out[33] = s_CSAwallace_cska24_u_cska48_out[33];
  assign s_CSAwallace_cska24_out[34] = s_CSAwallace_cska24_u_cska48_out[34];
  assign s_CSAwallace_cska24_out[35] = s_CSAwallace_cska24_u_cska48_out[35];
  assign s_CSAwallace_cska24_out[36] = s_CSAwallace_cska24_u_cska48_out[36];
  assign s_CSAwallace_cska24_out[37] = s_CSAwallace_cska24_u_cska48_out[37];
  assign s_CSAwallace_cska24_out[38] = s_CSAwallace_cska24_u_cska48_out[38];
  assign s_CSAwallace_cska24_out[39] = s_CSAwallace_cska24_u_cska48_out[39];
  assign s_CSAwallace_cska24_out[40] = s_CSAwallace_cska24_u_cska48_out[40];
  assign s_CSAwallace_cska24_out[41] = s_CSAwallace_cska24_u_cska48_out[41];
  assign s_CSAwallace_cska24_out[42] = s_CSAwallace_cska24_u_cska48_out[42];
  assign s_CSAwallace_cska24_out[43] = s_CSAwallace_cska24_u_cska48_out[43];
  assign s_CSAwallace_cska24_out[44] = s_CSAwallace_cska24_u_cska48_out[44];
  assign s_CSAwallace_cska24_out[45] = s_CSAwallace_cska24_u_cska48_out[45];
  assign s_CSAwallace_cska24_out[46] = s_CSAwallace_cska24_u_cska48_out[46];
  assign s_CSAwallace_cska24_out[47] = s_CSAwallace_cska24_xor0[0];
endmodule