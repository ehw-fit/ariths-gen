module f_s_cla24(input [23:0] a, input [23:0] b, output [24:0] f_s_cla24_out);
  wire f_s_cla24_pg_logic0_or0;
  wire f_s_cla24_pg_logic0_and0;
  wire f_s_cla24_pg_logic0_xor0;
  wire f_s_cla24_pg_logic1_or0;
  wire f_s_cla24_pg_logic1_and0;
  wire f_s_cla24_pg_logic1_xor0;
  wire f_s_cla24_xor1;
  wire f_s_cla24_and0;
  wire f_s_cla24_or0;
  wire f_s_cla24_pg_logic2_or0;
  wire f_s_cla24_pg_logic2_and0;
  wire f_s_cla24_pg_logic2_xor0;
  wire f_s_cla24_xor2;
  wire f_s_cla24_and1;
  wire f_s_cla24_and2;
  wire f_s_cla24_and3;
  wire f_s_cla24_and4;
  wire f_s_cla24_or1;
  wire f_s_cla24_or2;
  wire f_s_cla24_pg_logic3_or0;
  wire f_s_cla24_pg_logic3_and0;
  wire f_s_cla24_pg_logic3_xor0;
  wire f_s_cla24_xor3;
  wire f_s_cla24_and5;
  wire f_s_cla24_and6;
  wire f_s_cla24_and7;
  wire f_s_cla24_and8;
  wire f_s_cla24_and9;
  wire f_s_cla24_and10;
  wire f_s_cla24_and11;
  wire f_s_cla24_or3;
  wire f_s_cla24_or4;
  wire f_s_cla24_or5;
  wire f_s_cla24_pg_logic4_or0;
  wire f_s_cla24_pg_logic4_and0;
  wire f_s_cla24_pg_logic4_xor0;
  wire f_s_cla24_xor4;
  wire f_s_cla24_and12;
  wire f_s_cla24_or6;
  wire f_s_cla24_pg_logic5_or0;
  wire f_s_cla24_pg_logic5_and0;
  wire f_s_cla24_pg_logic5_xor0;
  wire f_s_cla24_xor5;
  wire f_s_cla24_and13;
  wire f_s_cla24_and14;
  wire f_s_cla24_and15;
  wire f_s_cla24_or7;
  wire f_s_cla24_or8;
  wire f_s_cla24_pg_logic6_or0;
  wire f_s_cla24_pg_logic6_and0;
  wire f_s_cla24_pg_logic6_xor0;
  wire f_s_cla24_xor6;
  wire f_s_cla24_and16;
  wire f_s_cla24_and17;
  wire f_s_cla24_and18;
  wire f_s_cla24_and19;
  wire f_s_cla24_and20;
  wire f_s_cla24_and21;
  wire f_s_cla24_or9;
  wire f_s_cla24_or10;
  wire f_s_cla24_or11;
  wire f_s_cla24_pg_logic7_or0;
  wire f_s_cla24_pg_logic7_and0;
  wire f_s_cla24_pg_logic7_xor0;
  wire f_s_cla24_xor7;
  wire f_s_cla24_and22;
  wire f_s_cla24_and23;
  wire f_s_cla24_and24;
  wire f_s_cla24_and25;
  wire f_s_cla24_and26;
  wire f_s_cla24_and27;
  wire f_s_cla24_and28;
  wire f_s_cla24_and29;
  wire f_s_cla24_and30;
  wire f_s_cla24_and31;
  wire f_s_cla24_or12;
  wire f_s_cla24_or13;
  wire f_s_cla24_or14;
  wire f_s_cla24_or15;
  wire f_s_cla24_pg_logic8_or0;
  wire f_s_cla24_pg_logic8_and0;
  wire f_s_cla24_pg_logic8_xor0;
  wire f_s_cla24_xor8;
  wire f_s_cla24_and32;
  wire f_s_cla24_or16;
  wire f_s_cla24_pg_logic9_or0;
  wire f_s_cla24_pg_logic9_and0;
  wire f_s_cla24_pg_logic9_xor0;
  wire f_s_cla24_xor9;
  wire f_s_cla24_and33;
  wire f_s_cla24_and34;
  wire f_s_cla24_and35;
  wire f_s_cla24_or17;
  wire f_s_cla24_or18;
  wire f_s_cla24_pg_logic10_or0;
  wire f_s_cla24_pg_logic10_and0;
  wire f_s_cla24_pg_logic10_xor0;
  wire f_s_cla24_xor10;
  wire f_s_cla24_and36;
  wire f_s_cla24_and37;
  wire f_s_cla24_and38;
  wire f_s_cla24_and39;
  wire f_s_cla24_and40;
  wire f_s_cla24_and41;
  wire f_s_cla24_or19;
  wire f_s_cla24_or20;
  wire f_s_cla24_or21;
  wire f_s_cla24_pg_logic11_or0;
  wire f_s_cla24_pg_logic11_and0;
  wire f_s_cla24_pg_logic11_xor0;
  wire f_s_cla24_xor11;
  wire f_s_cla24_and42;
  wire f_s_cla24_and43;
  wire f_s_cla24_and44;
  wire f_s_cla24_and45;
  wire f_s_cla24_and46;
  wire f_s_cla24_and47;
  wire f_s_cla24_and48;
  wire f_s_cla24_and49;
  wire f_s_cla24_and50;
  wire f_s_cla24_and51;
  wire f_s_cla24_or22;
  wire f_s_cla24_or23;
  wire f_s_cla24_or24;
  wire f_s_cla24_or25;
  wire f_s_cla24_pg_logic12_or0;
  wire f_s_cla24_pg_logic12_and0;
  wire f_s_cla24_pg_logic12_xor0;
  wire f_s_cla24_xor12;
  wire f_s_cla24_and52;
  wire f_s_cla24_or26;
  wire f_s_cla24_pg_logic13_or0;
  wire f_s_cla24_pg_logic13_and0;
  wire f_s_cla24_pg_logic13_xor0;
  wire f_s_cla24_xor13;
  wire f_s_cla24_and53;
  wire f_s_cla24_and54;
  wire f_s_cla24_and55;
  wire f_s_cla24_or27;
  wire f_s_cla24_or28;
  wire f_s_cla24_pg_logic14_or0;
  wire f_s_cla24_pg_logic14_and0;
  wire f_s_cla24_pg_logic14_xor0;
  wire f_s_cla24_xor14;
  wire f_s_cla24_and56;
  wire f_s_cla24_and57;
  wire f_s_cla24_and58;
  wire f_s_cla24_and59;
  wire f_s_cla24_and60;
  wire f_s_cla24_and61;
  wire f_s_cla24_or29;
  wire f_s_cla24_or30;
  wire f_s_cla24_or31;
  wire f_s_cla24_pg_logic15_or0;
  wire f_s_cla24_pg_logic15_and0;
  wire f_s_cla24_pg_logic15_xor0;
  wire f_s_cla24_xor15;
  wire f_s_cla24_and62;
  wire f_s_cla24_and63;
  wire f_s_cla24_and64;
  wire f_s_cla24_and65;
  wire f_s_cla24_and66;
  wire f_s_cla24_and67;
  wire f_s_cla24_and68;
  wire f_s_cla24_and69;
  wire f_s_cla24_and70;
  wire f_s_cla24_and71;
  wire f_s_cla24_or32;
  wire f_s_cla24_or33;
  wire f_s_cla24_or34;
  wire f_s_cla24_or35;
  wire f_s_cla24_pg_logic16_or0;
  wire f_s_cla24_pg_logic16_and0;
  wire f_s_cla24_pg_logic16_xor0;
  wire f_s_cla24_xor16;
  wire f_s_cla24_and72;
  wire f_s_cla24_or36;
  wire f_s_cla24_pg_logic17_or0;
  wire f_s_cla24_pg_logic17_and0;
  wire f_s_cla24_pg_logic17_xor0;
  wire f_s_cla24_xor17;
  wire f_s_cla24_and73;
  wire f_s_cla24_and74;
  wire f_s_cla24_and75;
  wire f_s_cla24_or37;
  wire f_s_cla24_or38;
  wire f_s_cla24_pg_logic18_or0;
  wire f_s_cla24_pg_logic18_and0;
  wire f_s_cla24_pg_logic18_xor0;
  wire f_s_cla24_xor18;
  wire f_s_cla24_and76;
  wire f_s_cla24_and77;
  wire f_s_cla24_and78;
  wire f_s_cla24_and79;
  wire f_s_cla24_and80;
  wire f_s_cla24_and81;
  wire f_s_cla24_or39;
  wire f_s_cla24_or40;
  wire f_s_cla24_or41;
  wire f_s_cla24_pg_logic19_or0;
  wire f_s_cla24_pg_logic19_and0;
  wire f_s_cla24_pg_logic19_xor0;
  wire f_s_cla24_xor19;
  wire f_s_cla24_and82;
  wire f_s_cla24_and83;
  wire f_s_cla24_and84;
  wire f_s_cla24_and85;
  wire f_s_cla24_and86;
  wire f_s_cla24_and87;
  wire f_s_cla24_and88;
  wire f_s_cla24_and89;
  wire f_s_cla24_and90;
  wire f_s_cla24_and91;
  wire f_s_cla24_or42;
  wire f_s_cla24_or43;
  wire f_s_cla24_or44;
  wire f_s_cla24_or45;
  wire f_s_cla24_pg_logic20_or0;
  wire f_s_cla24_pg_logic20_and0;
  wire f_s_cla24_pg_logic20_xor0;
  wire f_s_cla24_xor20;
  wire f_s_cla24_and92;
  wire f_s_cla24_or46;
  wire f_s_cla24_pg_logic21_or0;
  wire f_s_cla24_pg_logic21_and0;
  wire f_s_cla24_pg_logic21_xor0;
  wire f_s_cla24_xor21;
  wire f_s_cla24_and93;
  wire f_s_cla24_and94;
  wire f_s_cla24_and95;
  wire f_s_cla24_or47;
  wire f_s_cla24_or48;
  wire f_s_cla24_pg_logic22_or0;
  wire f_s_cla24_pg_logic22_and0;
  wire f_s_cla24_pg_logic22_xor0;
  wire f_s_cla24_xor22;
  wire f_s_cla24_and96;
  wire f_s_cla24_and97;
  wire f_s_cla24_and98;
  wire f_s_cla24_and99;
  wire f_s_cla24_and100;
  wire f_s_cla24_and101;
  wire f_s_cla24_or49;
  wire f_s_cla24_or50;
  wire f_s_cla24_or51;
  wire f_s_cla24_pg_logic23_or0;
  wire f_s_cla24_pg_logic23_and0;
  wire f_s_cla24_pg_logic23_xor0;
  wire f_s_cla24_xor23;
  wire f_s_cla24_and102;
  wire f_s_cla24_and103;
  wire f_s_cla24_and104;
  wire f_s_cla24_and105;
  wire f_s_cla24_and106;
  wire f_s_cla24_and107;
  wire f_s_cla24_and108;
  wire f_s_cla24_and109;
  wire f_s_cla24_and110;
  wire f_s_cla24_and111;
  wire f_s_cla24_or52;
  wire f_s_cla24_or53;
  wire f_s_cla24_or54;
  wire f_s_cla24_or55;
  wire f_s_cla24_xor24;
  wire f_s_cla24_xor25;

  assign f_s_cla24_pg_logic0_or0 = a[0] | b[0];
  assign f_s_cla24_pg_logic0_and0 = a[0] & b[0];
  assign f_s_cla24_pg_logic0_xor0 = a[0] ^ b[0];
  assign f_s_cla24_pg_logic1_or0 = a[1] | b[1];
  assign f_s_cla24_pg_logic1_and0 = a[1] & b[1];
  assign f_s_cla24_pg_logic1_xor0 = a[1] ^ b[1];
  assign f_s_cla24_xor1 = f_s_cla24_pg_logic1_xor0 ^ f_s_cla24_pg_logic0_and0;
  assign f_s_cla24_and0 = f_s_cla24_pg_logic0_and0 & f_s_cla24_pg_logic1_or0;
  assign f_s_cla24_or0 = f_s_cla24_pg_logic1_and0 | f_s_cla24_and0;
  assign f_s_cla24_pg_logic2_or0 = a[2] | b[2];
  assign f_s_cla24_pg_logic2_and0 = a[2] & b[2];
  assign f_s_cla24_pg_logic2_xor0 = a[2] ^ b[2];
  assign f_s_cla24_xor2 = f_s_cla24_pg_logic2_xor0 ^ f_s_cla24_or0;
  assign f_s_cla24_and1 = f_s_cla24_pg_logic2_or0 & f_s_cla24_pg_logic0_or0;
  assign f_s_cla24_and2 = f_s_cla24_pg_logic0_and0 & f_s_cla24_pg_logic2_or0;
  assign f_s_cla24_and3 = f_s_cla24_and2 & f_s_cla24_pg_logic1_or0;
  assign f_s_cla24_and4 = f_s_cla24_pg_logic1_and0 & f_s_cla24_pg_logic2_or0;
  assign f_s_cla24_or1 = f_s_cla24_and3 | f_s_cla24_and4;
  assign f_s_cla24_or2 = f_s_cla24_pg_logic2_and0 | f_s_cla24_or1;
  assign f_s_cla24_pg_logic3_or0 = a[3] | b[3];
  assign f_s_cla24_pg_logic3_and0 = a[3] & b[3];
  assign f_s_cla24_pg_logic3_xor0 = a[3] ^ b[3];
  assign f_s_cla24_xor3 = f_s_cla24_pg_logic3_xor0 ^ f_s_cla24_or2;
  assign f_s_cla24_and5 = f_s_cla24_pg_logic3_or0 & f_s_cla24_pg_logic1_or0;
  assign f_s_cla24_and6 = f_s_cla24_pg_logic0_and0 & f_s_cla24_pg_logic2_or0;
  assign f_s_cla24_and7 = f_s_cla24_pg_logic3_or0 & f_s_cla24_pg_logic1_or0;
  assign f_s_cla24_and8 = f_s_cla24_and6 & f_s_cla24_and7;
  assign f_s_cla24_and9 = f_s_cla24_pg_logic1_and0 & f_s_cla24_pg_logic3_or0;
  assign f_s_cla24_and10 = f_s_cla24_and9 & f_s_cla24_pg_logic2_or0;
  assign f_s_cla24_and11 = f_s_cla24_pg_logic2_and0 & f_s_cla24_pg_logic3_or0;
  assign f_s_cla24_or3 = f_s_cla24_and8 | f_s_cla24_and11;
  assign f_s_cla24_or4 = f_s_cla24_and10 | f_s_cla24_or3;
  assign f_s_cla24_or5 = f_s_cla24_pg_logic3_and0 | f_s_cla24_or4;
  assign f_s_cla24_pg_logic4_or0 = a[4] | b[4];
  assign f_s_cla24_pg_logic4_and0 = a[4] & b[4];
  assign f_s_cla24_pg_logic4_xor0 = a[4] ^ b[4];
  assign f_s_cla24_xor4 = f_s_cla24_pg_logic4_xor0 ^ f_s_cla24_or5;
  assign f_s_cla24_and12 = f_s_cla24_or5 & f_s_cla24_pg_logic4_or0;
  assign f_s_cla24_or6 = f_s_cla24_pg_logic4_and0 | f_s_cla24_and12;
  assign f_s_cla24_pg_logic5_or0 = a[5] | b[5];
  assign f_s_cla24_pg_logic5_and0 = a[5] & b[5];
  assign f_s_cla24_pg_logic5_xor0 = a[5] ^ b[5];
  assign f_s_cla24_xor5 = f_s_cla24_pg_logic5_xor0 ^ f_s_cla24_or6;
  assign f_s_cla24_and13 = f_s_cla24_or5 & f_s_cla24_pg_logic5_or0;
  assign f_s_cla24_and14 = f_s_cla24_and13 & f_s_cla24_pg_logic4_or0;
  assign f_s_cla24_and15 = f_s_cla24_pg_logic4_and0 & f_s_cla24_pg_logic5_or0;
  assign f_s_cla24_or7 = f_s_cla24_and14 | f_s_cla24_and15;
  assign f_s_cla24_or8 = f_s_cla24_pg_logic5_and0 | f_s_cla24_or7;
  assign f_s_cla24_pg_logic6_or0 = a[6] | b[6];
  assign f_s_cla24_pg_logic6_and0 = a[6] & b[6];
  assign f_s_cla24_pg_logic6_xor0 = a[6] ^ b[6];
  assign f_s_cla24_xor6 = f_s_cla24_pg_logic6_xor0 ^ f_s_cla24_or8;
  assign f_s_cla24_and16 = f_s_cla24_or5 & f_s_cla24_pg_logic5_or0;
  assign f_s_cla24_and17 = f_s_cla24_pg_logic6_or0 & f_s_cla24_pg_logic4_or0;
  assign f_s_cla24_and18 = f_s_cla24_and16 & f_s_cla24_and17;
  assign f_s_cla24_and19 = f_s_cla24_pg_logic4_and0 & f_s_cla24_pg_logic6_or0;
  assign f_s_cla24_and20 = f_s_cla24_and19 & f_s_cla24_pg_logic5_or0;
  assign f_s_cla24_and21 = f_s_cla24_pg_logic5_and0 & f_s_cla24_pg_logic6_or0;
  assign f_s_cla24_or9 = f_s_cla24_and18 | f_s_cla24_and20;
  assign f_s_cla24_or10 = f_s_cla24_or9 | f_s_cla24_and21;
  assign f_s_cla24_or11 = f_s_cla24_pg_logic6_and0 | f_s_cla24_or10;
  assign f_s_cla24_pg_logic7_or0 = a[7] | b[7];
  assign f_s_cla24_pg_logic7_and0 = a[7] & b[7];
  assign f_s_cla24_pg_logic7_xor0 = a[7] ^ b[7];
  assign f_s_cla24_xor7 = f_s_cla24_pg_logic7_xor0 ^ f_s_cla24_or11;
  assign f_s_cla24_and22 = f_s_cla24_or5 & f_s_cla24_pg_logic6_or0;
  assign f_s_cla24_and23 = f_s_cla24_pg_logic7_or0 & f_s_cla24_pg_logic5_or0;
  assign f_s_cla24_and24 = f_s_cla24_and22 & f_s_cla24_and23;
  assign f_s_cla24_and25 = f_s_cla24_and24 & f_s_cla24_pg_logic4_or0;
  assign f_s_cla24_and26 = f_s_cla24_pg_logic4_and0 & f_s_cla24_pg_logic6_or0;
  assign f_s_cla24_and27 = f_s_cla24_pg_logic7_or0 & f_s_cla24_pg_logic5_or0;
  assign f_s_cla24_and28 = f_s_cla24_and26 & f_s_cla24_and27;
  assign f_s_cla24_and29 = f_s_cla24_pg_logic5_and0 & f_s_cla24_pg_logic7_or0;
  assign f_s_cla24_and30 = f_s_cla24_and29 & f_s_cla24_pg_logic6_or0;
  assign f_s_cla24_and31 = f_s_cla24_pg_logic6_and0 & f_s_cla24_pg_logic7_or0;
  assign f_s_cla24_or12 = f_s_cla24_and25 | f_s_cla24_and30;
  assign f_s_cla24_or13 = f_s_cla24_and28 | f_s_cla24_and31;
  assign f_s_cla24_or14 = f_s_cla24_or12 | f_s_cla24_or13;
  assign f_s_cla24_or15 = f_s_cla24_pg_logic7_and0 | f_s_cla24_or14;
  assign f_s_cla24_pg_logic8_or0 = a[8] | b[8];
  assign f_s_cla24_pg_logic8_and0 = a[8] & b[8];
  assign f_s_cla24_pg_logic8_xor0 = a[8] ^ b[8];
  assign f_s_cla24_xor8 = f_s_cla24_pg_logic8_xor0 ^ f_s_cla24_or15;
  assign f_s_cla24_and32 = f_s_cla24_or15 & f_s_cla24_pg_logic8_or0;
  assign f_s_cla24_or16 = f_s_cla24_pg_logic8_and0 | f_s_cla24_and32;
  assign f_s_cla24_pg_logic9_or0 = a[9] | b[9];
  assign f_s_cla24_pg_logic9_and0 = a[9] & b[9];
  assign f_s_cla24_pg_logic9_xor0 = a[9] ^ b[9];
  assign f_s_cla24_xor9 = f_s_cla24_pg_logic9_xor0 ^ f_s_cla24_or16;
  assign f_s_cla24_and33 = f_s_cla24_or15 & f_s_cla24_pg_logic9_or0;
  assign f_s_cla24_and34 = f_s_cla24_and33 & f_s_cla24_pg_logic8_or0;
  assign f_s_cla24_and35 = f_s_cla24_pg_logic8_and0 & f_s_cla24_pg_logic9_or0;
  assign f_s_cla24_or17 = f_s_cla24_and34 | f_s_cla24_and35;
  assign f_s_cla24_or18 = f_s_cla24_pg_logic9_and0 | f_s_cla24_or17;
  assign f_s_cla24_pg_logic10_or0 = a[10] | b[10];
  assign f_s_cla24_pg_logic10_and0 = a[10] & b[10];
  assign f_s_cla24_pg_logic10_xor0 = a[10] ^ b[10];
  assign f_s_cla24_xor10 = f_s_cla24_pg_logic10_xor0 ^ f_s_cla24_or18;
  assign f_s_cla24_and36 = f_s_cla24_or15 & f_s_cla24_pg_logic9_or0;
  assign f_s_cla24_and37 = f_s_cla24_pg_logic10_or0 & f_s_cla24_pg_logic8_or0;
  assign f_s_cla24_and38 = f_s_cla24_and36 & f_s_cla24_and37;
  assign f_s_cla24_and39 = f_s_cla24_pg_logic8_and0 & f_s_cla24_pg_logic10_or0;
  assign f_s_cla24_and40 = f_s_cla24_and39 & f_s_cla24_pg_logic9_or0;
  assign f_s_cla24_and41 = f_s_cla24_pg_logic9_and0 & f_s_cla24_pg_logic10_or0;
  assign f_s_cla24_or19 = f_s_cla24_and38 | f_s_cla24_and40;
  assign f_s_cla24_or20 = f_s_cla24_or19 | f_s_cla24_and41;
  assign f_s_cla24_or21 = f_s_cla24_pg_logic10_and0 | f_s_cla24_or20;
  assign f_s_cla24_pg_logic11_or0 = a[11] | b[11];
  assign f_s_cla24_pg_logic11_and0 = a[11] & b[11];
  assign f_s_cla24_pg_logic11_xor0 = a[11] ^ b[11];
  assign f_s_cla24_xor11 = f_s_cla24_pg_logic11_xor0 ^ f_s_cla24_or21;
  assign f_s_cla24_and42 = f_s_cla24_or15 & f_s_cla24_pg_logic10_or0;
  assign f_s_cla24_and43 = f_s_cla24_pg_logic11_or0 & f_s_cla24_pg_logic9_or0;
  assign f_s_cla24_and44 = f_s_cla24_and42 & f_s_cla24_and43;
  assign f_s_cla24_and45 = f_s_cla24_and44 & f_s_cla24_pg_logic8_or0;
  assign f_s_cla24_and46 = f_s_cla24_pg_logic8_and0 & f_s_cla24_pg_logic10_or0;
  assign f_s_cla24_and47 = f_s_cla24_pg_logic11_or0 & f_s_cla24_pg_logic9_or0;
  assign f_s_cla24_and48 = f_s_cla24_and46 & f_s_cla24_and47;
  assign f_s_cla24_and49 = f_s_cla24_pg_logic9_and0 & f_s_cla24_pg_logic11_or0;
  assign f_s_cla24_and50 = f_s_cla24_and49 & f_s_cla24_pg_logic10_or0;
  assign f_s_cla24_and51 = f_s_cla24_pg_logic10_and0 & f_s_cla24_pg_logic11_or0;
  assign f_s_cla24_or22 = f_s_cla24_and45 | f_s_cla24_and50;
  assign f_s_cla24_or23 = f_s_cla24_and48 | f_s_cla24_and51;
  assign f_s_cla24_or24 = f_s_cla24_or22 | f_s_cla24_or23;
  assign f_s_cla24_or25 = f_s_cla24_pg_logic11_and0 | f_s_cla24_or24;
  assign f_s_cla24_pg_logic12_or0 = a[12] | b[12];
  assign f_s_cla24_pg_logic12_and0 = a[12] & b[12];
  assign f_s_cla24_pg_logic12_xor0 = a[12] ^ b[12];
  assign f_s_cla24_xor12 = f_s_cla24_pg_logic12_xor0 ^ f_s_cla24_or25;
  assign f_s_cla24_and52 = f_s_cla24_or25 & f_s_cla24_pg_logic12_or0;
  assign f_s_cla24_or26 = f_s_cla24_pg_logic12_and0 | f_s_cla24_and52;
  assign f_s_cla24_pg_logic13_or0 = a[13] | b[13];
  assign f_s_cla24_pg_logic13_and0 = a[13] & b[13];
  assign f_s_cla24_pg_logic13_xor0 = a[13] ^ b[13];
  assign f_s_cla24_xor13 = f_s_cla24_pg_logic13_xor0 ^ f_s_cla24_or26;
  assign f_s_cla24_and53 = f_s_cla24_or25 & f_s_cla24_pg_logic13_or0;
  assign f_s_cla24_and54 = f_s_cla24_and53 & f_s_cla24_pg_logic12_or0;
  assign f_s_cla24_and55 = f_s_cla24_pg_logic12_and0 & f_s_cla24_pg_logic13_or0;
  assign f_s_cla24_or27 = f_s_cla24_and54 | f_s_cla24_and55;
  assign f_s_cla24_or28 = f_s_cla24_pg_logic13_and0 | f_s_cla24_or27;
  assign f_s_cla24_pg_logic14_or0 = a[14] | b[14];
  assign f_s_cla24_pg_logic14_and0 = a[14] & b[14];
  assign f_s_cla24_pg_logic14_xor0 = a[14] ^ b[14];
  assign f_s_cla24_xor14 = f_s_cla24_pg_logic14_xor0 ^ f_s_cla24_or28;
  assign f_s_cla24_and56 = f_s_cla24_or25 & f_s_cla24_pg_logic13_or0;
  assign f_s_cla24_and57 = f_s_cla24_pg_logic14_or0 & f_s_cla24_pg_logic12_or0;
  assign f_s_cla24_and58 = f_s_cla24_and56 & f_s_cla24_and57;
  assign f_s_cla24_and59 = f_s_cla24_pg_logic12_and0 & f_s_cla24_pg_logic14_or0;
  assign f_s_cla24_and60 = f_s_cla24_and59 & f_s_cla24_pg_logic13_or0;
  assign f_s_cla24_and61 = f_s_cla24_pg_logic13_and0 & f_s_cla24_pg_logic14_or0;
  assign f_s_cla24_or29 = f_s_cla24_and58 | f_s_cla24_and60;
  assign f_s_cla24_or30 = f_s_cla24_or29 | f_s_cla24_and61;
  assign f_s_cla24_or31 = f_s_cla24_pg_logic14_and0 | f_s_cla24_or30;
  assign f_s_cla24_pg_logic15_or0 = a[15] | b[15];
  assign f_s_cla24_pg_logic15_and0 = a[15] & b[15];
  assign f_s_cla24_pg_logic15_xor0 = a[15] ^ b[15];
  assign f_s_cla24_xor15 = f_s_cla24_pg_logic15_xor0 ^ f_s_cla24_or31;
  assign f_s_cla24_and62 = f_s_cla24_or25 & f_s_cla24_pg_logic14_or0;
  assign f_s_cla24_and63 = f_s_cla24_pg_logic15_or0 & f_s_cla24_pg_logic13_or0;
  assign f_s_cla24_and64 = f_s_cla24_and62 & f_s_cla24_and63;
  assign f_s_cla24_and65 = f_s_cla24_and64 & f_s_cla24_pg_logic12_or0;
  assign f_s_cla24_and66 = f_s_cla24_pg_logic12_and0 & f_s_cla24_pg_logic14_or0;
  assign f_s_cla24_and67 = f_s_cla24_pg_logic15_or0 & f_s_cla24_pg_logic13_or0;
  assign f_s_cla24_and68 = f_s_cla24_and66 & f_s_cla24_and67;
  assign f_s_cla24_and69 = f_s_cla24_pg_logic13_and0 & f_s_cla24_pg_logic15_or0;
  assign f_s_cla24_and70 = f_s_cla24_and69 & f_s_cla24_pg_logic14_or0;
  assign f_s_cla24_and71 = f_s_cla24_pg_logic14_and0 & f_s_cla24_pg_logic15_or0;
  assign f_s_cla24_or32 = f_s_cla24_and65 | f_s_cla24_and70;
  assign f_s_cla24_or33 = f_s_cla24_and68 | f_s_cla24_and71;
  assign f_s_cla24_or34 = f_s_cla24_or32 | f_s_cla24_or33;
  assign f_s_cla24_or35 = f_s_cla24_pg_logic15_and0 | f_s_cla24_or34;
  assign f_s_cla24_pg_logic16_or0 = a[16] | b[16];
  assign f_s_cla24_pg_logic16_and0 = a[16] & b[16];
  assign f_s_cla24_pg_logic16_xor0 = a[16] ^ b[16];
  assign f_s_cla24_xor16 = f_s_cla24_pg_logic16_xor0 ^ f_s_cla24_or35;
  assign f_s_cla24_and72 = f_s_cla24_or35 & f_s_cla24_pg_logic16_or0;
  assign f_s_cla24_or36 = f_s_cla24_pg_logic16_and0 | f_s_cla24_and72;
  assign f_s_cla24_pg_logic17_or0 = a[17] | b[17];
  assign f_s_cla24_pg_logic17_and0 = a[17] & b[17];
  assign f_s_cla24_pg_logic17_xor0 = a[17] ^ b[17];
  assign f_s_cla24_xor17 = f_s_cla24_pg_logic17_xor0 ^ f_s_cla24_or36;
  assign f_s_cla24_and73 = f_s_cla24_or35 & f_s_cla24_pg_logic17_or0;
  assign f_s_cla24_and74 = f_s_cla24_and73 & f_s_cla24_pg_logic16_or0;
  assign f_s_cla24_and75 = f_s_cla24_pg_logic16_and0 & f_s_cla24_pg_logic17_or0;
  assign f_s_cla24_or37 = f_s_cla24_and74 | f_s_cla24_and75;
  assign f_s_cla24_or38 = f_s_cla24_pg_logic17_and0 | f_s_cla24_or37;
  assign f_s_cla24_pg_logic18_or0 = a[18] | b[18];
  assign f_s_cla24_pg_logic18_and0 = a[18] & b[18];
  assign f_s_cla24_pg_logic18_xor0 = a[18] ^ b[18];
  assign f_s_cla24_xor18 = f_s_cla24_pg_logic18_xor0 ^ f_s_cla24_or38;
  assign f_s_cla24_and76 = f_s_cla24_or35 & f_s_cla24_pg_logic17_or0;
  assign f_s_cla24_and77 = f_s_cla24_pg_logic18_or0 & f_s_cla24_pg_logic16_or0;
  assign f_s_cla24_and78 = f_s_cla24_and76 & f_s_cla24_and77;
  assign f_s_cla24_and79 = f_s_cla24_pg_logic16_and0 & f_s_cla24_pg_logic18_or0;
  assign f_s_cla24_and80 = f_s_cla24_and79 & f_s_cla24_pg_logic17_or0;
  assign f_s_cla24_and81 = f_s_cla24_pg_logic17_and0 & f_s_cla24_pg_logic18_or0;
  assign f_s_cla24_or39 = f_s_cla24_and78 | f_s_cla24_and80;
  assign f_s_cla24_or40 = f_s_cla24_or39 | f_s_cla24_and81;
  assign f_s_cla24_or41 = f_s_cla24_pg_logic18_and0 | f_s_cla24_or40;
  assign f_s_cla24_pg_logic19_or0 = a[19] | b[19];
  assign f_s_cla24_pg_logic19_and0 = a[19] & b[19];
  assign f_s_cla24_pg_logic19_xor0 = a[19] ^ b[19];
  assign f_s_cla24_xor19 = f_s_cla24_pg_logic19_xor0 ^ f_s_cla24_or41;
  assign f_s_cla24_and82 = f_s_cla24_or35 & f_s_cla24_pg_logic18_or0;
  assign f_s_cla24_and83 = f_s_cla24_pg_logic19_or0 & f_s_cla24_pg_logic17_or0;
  assign f_s_cla24_and84 = f_s_cla24_and82 & f_s_cla24_and83;
  assign f_s_cla24_and85 = f_s_cla24_and84 & f_s_cla24_pg_logic16_or0;
  assign f_s_cla24_and86 = f_s_cla24_pg_logic16_and0 & f_s_cla24_pg_logic18_or0;
  assign f_s_cla24_and87 = f_s_cla24_pg_logic19_or0 & f_s_cla24_pg_logic17_or0;
  assign f_s_cla24_and88 = f_s_cla24_and86 & f_s_cla24_and87;
  assign f_s_cla24_and89 = f_s_cla24_pg_logic17_and0 & f_s_cla24_pg_logic19_or0;
  assign f_s_cla24_and90 = f_s_cla24_and89 & f_s_cla24_pg_logic18_or0;
  assign f_s_cla24_and91 = f_s_cla24_pg_logic18_and0 & f_s_cla24_pg_logic19_or0;
  assign f_s_cla24_or42 = f_s_cla24_and85 | f_s_cla24_and90;
  assign f_s_cla24_or43 = f_s_cla24_and88 | f_s_cla24_and91;
  assign f_s_cla24_or44 = f_s_cla24_or42 | f_s_cla24_or43;
  assign f_s_cla24_or45 = f_s_cla24_pg_logic19_and0 | f_s_cla24_or44;
  assign f_s_cla24_pg_logic20_or0 = a[20] | b[20];
  assign f_s_cla24_pg_logic20_and0 = a[20] & b[20];
  assign f_s_cla24_pg_logic20_xor0 = a[20] ^ b[20];
  assign f_s_cla24_xor20 = f_s_cla24_pg_logic20_xor0 ^ f_s_cla24_or45;
  assign f_s_cla24_and92 = f_s_cla24_or45 & f_s_cla24_pg_logic20_or0;
  assign f_s_cla24_or46 = f_s_cla24_pg_logic20_and0 | f_s_cla24_and92;
  assign f_s_cla24_pg_logic21_or0 = a[21] | b[21];
  assign f_s_cla24_pg_logic21_and0 = a[21] & b[21];
  assign f_s_cla24_pg_logic21_xor0 = a[21] ^ b[21];
  assign f_s_cla24_xor21 = f_s_cla24_pg_logic21_xor0 ^ f_s_cla24_or46;
  assign f_s_cla24_and93 = f_s_cla24_or45 & f_s_cla24_pg_logic21_or0;
  assign f_s_cla24_and94 = f_s_cla24_and93 & f_s_cla24_pg_logic20_or0;
  assign f_s_cla24_and95 = f_s_cla24_pg_logic20_and0 & f_s_cla24_pg_logic21_or0;
  assign f_s_cla24_or47 = f_s_cla24_and94 | f_s_cla24_and95;
  assign f_s_cla24_or48 = f_s_cla24_pg_logic21_and0 | f_s_cla24_or47;
  assign f_s_cla24_pg_logic22_or0 = a[22] | b[22];
  assign f_s_cla24_pg_logic22_and0 = a[22] & b[22];
  assign f_s_cla24_pg_logic22_xor0 = a[22] ^ b[22];
  assign f_s_cla24_xor22 = f_s_cla24_pg_logic22_xor0 ^ f_s_cla24_or48;
  assign f_s_cla24_and96 = f_s_cla24_or45 & f_s_cla24_pg_logic21_or0;
  assign f_s_cla24_and97 = f_s_cla24_pg_logic22_or0 & f_s_cla24_pg_logic20_or0;
  assign f_s_cla24_and98 = f_s_cla24_and96 & f_s_cla24_and97;
  assign f_s_cla24_and99 = f_s_cla24_pg_logic20_and0 & f_s_cla24_pg_logic22_or0;
  assign f_s_cla24_and100 = f_s_cla24_and99 & f_s_cla24_pg_logic21_or0;
  assign f_s_cla24_and101 = f_s_cla24_pg_logic21_and0 & f_s_cla24_pg_logic22_or0;
  assign f_s_cla24_or49 = f_s_cla24_and98 | f_s_cla24_and100;
  assign f_s_cla24_or50 = f_s_cla24_or49 | f_s_cla24_and101;
  assign f_s_cla24_or51 = f_s_cla24_pg_logic22_and0 | f_s_cla24_or50;
  assign f_s_cla24_pg_logic23_or0 = a[23] | b[23];
  assign f_s_cla24_pg_logic23_and0 = a[23] & b[23];
  assign f_s_cla24_pg_logic23_xor0 = a[23] ^ b[23];
  assign f_s_cla24_xor23 = f_s_cla24_pg_logic23_xor0 ^ f_s_cla24_or51;
  assign f_s_cla24_and102 = f_s_cla24_or45 & f_s_cla24_pg_logic22_or0;
  assign f_s_cla24_and103 = f_s_cla24_pg_logic23_or0 & f_s_cla24_pg_logic21_or0;
  assign f_s_cla24_and104 = f_s_cla24_and102 & f_s_cla24_and103;
  assign f_s_cla24_and105 = f_s_cla24_and104 & f_s_cla24_pg_logic20_or0;
  assign f_s_cla24_and106 = f_s_cla24_pg_logic20_and0 & f_s_cla24_pg_logic22_or0;
  assign f_s_cla24_and107 = f_s_cla24_pg_logic23_or0 & f_s_cla24_pg_logic21_or0;
  assign f_s_cla24_and108 = f_s_cla24_and106 & f_s_cla24_and107;
  assign f_s_cla24_and109 = f_s_cla24_pg_logic21_and0 & f_s_cla24_pg_logic23_or0;
  assign f_s_cla24_and110 = f_s_cla24_and109 & f_s_cla24_pg_logic22_or0;
  assign f_s_cla24_and111 = f_s_cla24_pg_logic22_and0 & f_s_cla24_pg_logic23_or0;
  assign f_s_cla24_or52 = f_s_cla24_and105 | f_s_cla24_and110;
  assign f_s_cla24_or53 = f_s_cla24_and108 | f_s_cla24_and111;
  assign f_s_cla24_or54 = f_s_cla24_or52 | f_s_cla24_or53;
  assign f_s_cla24_or55 = f_s_cla24_pg_logic23_and0 | f_s_cla24_or54;
  assign f_s_cla24_xor24 = a[23] ^ b[23];
  assign f_s_cla24_xor25 = f_s_cla24_xor24 ^ f_s_cla24_or55;

  assign f_s_cla24_out[0] = f_s_cla24_pg_logic0_xor0;
  assign f_s_cla24_out[1] = f_s_cla24_xor1;
  assign f_s_cla24_out[2] = f_s_cla24_xor2;
  assign f_s_cla24_out[3] = f_s_cla24_xor3;
  assign f_s_cla24_out[4] = f_s_cla24_xor4;
  assign f_s_cla24_out[5] = f_s_cla24_xor5;
  assign f_s_cla24_out[6] = f_s_cla24_xor6;
  assign f_s_cla24_out[7] = f_s_cla24_xor7;
  assign f_s_cla24_out[8] = f_s_cla24_xor8;
  assign f_s_cla24_out[9] = f_s_cla24_xor9;
  assign f_s_cla24_out[10] = f_s_cla24_xor10;
  assign f_s_cla24_out[11] = f_s_cla24_xor11;
  assign f_s_cla24_out[12] = f_s_cla24_xor12;
  assign f_s_cla24_out[13] = f_s_cla24_xor13;
  assign f_s_cla24_out[14] = f_s_cla24_xor14;
  assign f_s_cla24_out[15] = f_s_cla24_xor15;
  assign f_s_cla24_out[16] = f_s_cla24_xor16;
  assign f_s_cla24_out[17] = f_s_cla24_xor17;
  assign f_s_cla24_out[18] = f_s_cla24_xor18;
  assign f_s_cla24_out[19] = f_s_cla24_xor19;
  assign f_s_cla24_out[20] = f_s_cla24_xor20;
  assign f_s_cla24_out[21] = f_s_cla24_xor21;
  assign f_s_cla24_out[22] = f_s_cla24_xor22;
  assign f_s_cla24_out[23] = f_s_cla24_xor23;
  assign f_s_cla24_out[24] = f_s_cla24_xor25;
endmodule