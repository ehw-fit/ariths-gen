module f_s_rca32(input [31:0] a, input [31:0] b, output [32:0] f_s_rca32_out);
  wire f_s_rca32_ha_xor0;
  wire f_s_rca32_ha_and0;
  wire f_s_rca32_fa1_xor0;
  wire f_s_rca32_fa1_and0;
  wire f_s_rca32_fa1_xor1;
  wire f_s_rca32_fa1_and1;
  wire f_s_rca32_fa1_or0;
  wire f_s_rca32_fa2_xor0;
  wire f_s_rca32_fa2_and0;
  wire f_s_rca32_fa2_xor1;
  wire f_s_rca32_fa2_and1;
  wire f_s_rca32_fa2_or0;
  wire f_s_rca32_fa3_xor0;
  wire f_s_rca32_fa3_and0;
  wire f_s_rca32_fa3_xor1;
  wire f_s_rca32_fa3_and1;
  wire f_s_rca32_fa3_or0;
  wire f_s_rca32_fa4_xor0;
  wire f_s_rca32_fa4_and0;
  wire f_s_rca32_fa4_xor1;
  wire f_s_rca32_fa4_and1;
  wire f_s_rca32_fa4_or0;
  wire f_s_rca32_fa5_xor0;
  wire f_s_rca32_fa5_and0;
  wire f_s_rca32_fa5_xor1;
  wire f_s_rca32_fa5_and1;
  wire f_s_rca32_fa5_or0;
  wire f_s_rca32_fa6_xor0;
  wire f_s_rca32_fa6_and0;
  wire f_s_rca32_fa6_xor1;
  wire f_s_rca32_fa6_and1;
  wire f_s_rca32_fa6_or0;
  wire f_s_rca32_fa7_xor0;
  wire f_s_rca32_fa7_and0;
  wire f_s_rca32_fa7_xor1;
  wire f_s_rca32_fa7_and1;
  wire f_s_rca32_fa7_or0;
  wire f_s_rca32_fa8_xor0;
  wire f_s_rca32_fa8_and0;
  wire f_s_rca32_fa8_xor1;
  wire f_s_rca32_fa8_and1;
  wire f_s_rca32_fa8_or0;
  wire f_s_rca32_fa9_xor0;
  wire f_s_rca32_fa9_and0;
  wire f_s_rca32_fa9_xor1;
  wire f_s_rca32_fa9_and1;
  wire f_s_rca32_fa9_or0;
  wire f_s_rca32_fa10_xor0;
  wire f_s_rca32_fa10_and0;
  wire f_s_rca32_fa10_xor1;
  wire f_s_rca32_fa10_and1;
  wire f_s_rca32_fa10_or0;
  wire f_s_rca32_fa11_xor0;
  wire f_s_rca32_fa11_and0;
  wire f_s_rca32_fa11_xor1;
  wire f_s_rca32_fa11_and1;
  wire f_s_rca32_fa11_or0;
  wire f_s_rca32_fa12_xor0;
  wire f_s_rca32_fa12_and0;
  wire f_s_rca32_fa12_xor1;
  wire f_s_rca32_fa12_and1;
  wire f_s_rca32_fa12_or0;
  wire f_s_rca32_fa13_xor0;
  wire f_s_rca32_fa13_and0;
  wire f_s_rca32_fa13_xor1;
  wire f_s_rca32_fa13_and1;
  wire f_s_rca32_fa13_or0;
  wire f_s_rca32_fa14_xor0;
  wire f_s_rca32_fa14_and0;
  wire f_s_rca32_fa14_xor1;
  wire f_s_rca32_fa14_and1;
  wire f_s_rca32_fa14_or0;
  wire f_s_rca32_fa15_xor0;
  wire f_s_rca32_fa15_and0;
  wire f_s_rca32_fa15_xor1;
  wire f_s_rca32_fa15_and1;
  wire f_s_rca32_fa15_or0;
  wire f_s_rca32_fa16_xor0;
  wire f_s_rca32_fa16_and0;
  wire f_s_rca32_fa16_xor1;
  wire f_s_rca32_fa16_and1;
  wire f_s_rca32_fa16_or0;
  wire f_s_rca32_fa17_xor0;
  wire f_s_rca32_fa17_and0;
  wire f_s_rca32_fa17_xor1;
  wire f_s_rca32_fa17_and1;
  wire f_s_rca32_fa17_or0;
  wire f_s_rca32_fa18_xor0;
  wire f_s_rca32_fa18_and0;
  wire f_s_rca32_fa18_xor1;
  wire f_s_rca32_fa18_and1;
  wire f_s_rca32_fa18_or0;
  wire f_s_rca32_fa19_xor0;
  wire f_s_rca32_fa19_and0;
  wire f_s_rca32_fa19_xor1;
  wire f_s_rca32_fa19_and1;
  wire f_s_rca32_fa19_or0;
  wire f_s_rca32_fa20_xor0;
  wire f_s_rca32_fa20_and0;
  wire f_s_rca32_fa20_xor1;
  wire f_s_rca32_fa20_and1;
  wire f_s_rca32_fa20_or0;
  wire f_s_rca32_fa21_xor0;
  wire f_s_rca32_fa21_and0;
  wire f_s_rca32_fa21_xor1;
  wire f_s_rca32_fa21_and1;
  wire f_s_rca32_fa21_or0;
  wire f_s_rca32_fa22_xor0;
  wire f_s_rca32_fa22_and0;
  wire f_s_rca32_fa22_xor1;
  wire f_s_rca32_fa22_and1;
  wire f_s_rca32_fa22_or0;
  wire f_s_rca32_fa23_xor0;
  wire f_s_rca32_fa23_and0;
  wire f_s_rca32_fa23_xor1;
  wire f_s_rca32_fa23_and1;
  wire f_s_rca32_fa23_or0;
  wire f_s_rca32_fa24_xor0;
  wire f_s_rca32_fa24_and0;
  wire f_s_rca32_fa24_xor1;
  wire f_s_rca32_fa24_and1;
  wire f_s_rca32_fa24_or0;
  wire f_s_rca32_fa25_xor0;
  wire f_s_rca32_fa25_and0;
  wire f_s_rca32_fa25_xor1;
  wire f_s_rca32_fa25_and1;
  wire f_s_rca32_fa25_or0;
  wire f_s_rca32_fa26_xor0;
  wire f_s_rca32_fa26_and0;
  wire f_s_rca32_fa26_xor1;
  wire f_s_rca32_fa26_and1;
  wire f_s_rca32_fa26_or0;
  wire f_s_rca32_fa27_xor0;
  wire f_s_rca32_fa27_and0;
  wire f_s_rca32_fa27_xor1;
  wire f_s_rca32_fa27_and1;
  wire f_s_rca32_fa27_or0;
  wire f_s_rca32_fa28_xor0;
  wire f_s_rca32_fa28_and0;
  wire f_s_rca32_fa28_xor1;
  wire f_s_rca32_fa28_and1;
  wire f_s_rca32_fa28_or0;
  wire f_s_rca32_fa29_xor0;
  wire f_s_rca32_fa29_and0;
  wire f_s_rca32_fa29_xor1;
  wire f_s_rca32_fa29_and1;
  wire f_s_rca32_fa29_or0;
  wire f_s_rca32_fa30_xor0;
  wire f_s_rca32_fa30_and0;
  wire f_s_rca32_fa30_xor1;
  wire f_s_rca32_fa30_and1;
  wire f_s_rca32_fa30_or0;
  wire f_s_rca32_fa31_xor0;
  wire f_s_rca32_fa31_and0;
  wire f_s_rca32_fa31_xor1;
  wire f_s_rca32_fa31_and1;
  wire f_s_rca32_fa31_or0;
  wire f_s_rca32_xor0;
  wire f_s_rca32_xor1;

  assign f_s_rca32_ha_xor0 = a[0] ^ b[0];
  assign f_s_rca32_ha_and0 = a[0] & b[0];
  assign f_s_rca32_fa1_xor0 = a[1] ^ b[1];
  assign f_s_rca32_fa1_and0 = a[1] & b[1];
  assign f_s_rca32_fa1_xor1 = f_s_rca32_fa1_xor0 ^ f_s_rca32_ha_and0;
  assign f_s_rca32_fa1_and1 = f_s_rca32_fa1_xor0 & f_s_rca32_ha_and0;
  assign f_s_rca32_fa1_or0 = f_s_rca32_fa1_and0 | f_s_rca32_fa1_and1;
  assign f_s_rca32_fa2_xor0 = a[2] ^ b[2];
  assign f_s_rca32_fa2_and0 = a[2] & b[2];
  assign f_s_rca32_fa2_xor1 = f_s_rca32_fa2_xor0 ^ f_s_rca32_fa1_or0;
  assign f_s_rca32_fa2_and1 = f_s_rca32_fa2_xor0 & f_s_rca32_fa1_or0;
  assign f_s_rca32_fa2_or0 = f_s_rca32_fa2_and0 | f_s_rca32_fa2_and1;
  assign f_s_rca32_fa3_xor0 = a[3] ^ b[3];
  assign f_s_rca32_fa3_and0 = a[3] & b[3];
  assign f_s_rca32_fa3_xor1 = f_s_rca32_fa3_xor0 ^ f_s_rca32_fa2_or0;
  assign f_s_rca32_fa3_and1 = f_s_rca32_fa3_xor0 & f_s_rca32_fa2_or0;
  assign f_s_rca32_fa3_or0 = f_s_rca32_fa3_and0 | f_s_rca32_fa3_and1;
  assign f_s_rca32_fa4_xor0 = a[4] ^ b[4];
  assign f_s_rca32_fa4_and0 = a[4] & b[4];
  assign f_s_rca32_fa4_xor1 = f_s_rca32_fa4_xor0 ^ f_s_rca32_fa3_or0;
  assign f_s_rca32_fa4_and1 = f_s_rca32_fa4_xor0 & f_s_rca32_fa3_or0;
  assign f_s_rca32_fa4_or0 = f_s_rca32_fa4_and0 | f_s_rca32_fa4_and1;
  assign f_s_rca32_fa5_xor0 = a[5] ^ b[5];
  assign f_s_rca32_fa5_and0 = a[5] & b[5];
  assign f_s_rca32_fa5_xor1 = f_s_rca32_fa5_xor0 ^ f_s_rca32_fa4_or0;
  assign f_s_rca32_fa5_and1 = f_s_rca32_fa5_xor0 & f_s_rca32_fa4_or0;
  assign f_s_rca32_fa5_or0 = f_s_rca32_fa5_and0 | f_s_rca32_fa5_and1;
  assign f_s_rca32_fa6_xor0 = a[6] ^ b[6];
  assign f_s_rca32_fa6_and0 = a[6] & b[6];
  assign f_s_rca32_fa6_xor1 = f_s_rca32_fa6_xor0 ^ f_s_rca32_fa5_or0;
  assign f_s_rca32_fa6_and1 = f_s_rca32_fa6_xor0 & f_s_rca32_fa5_or0;
  assign f_s_rca32_fa6_or0 = f_s_rca32_fa6_and0 | f_s_rca32_fa6_and1;
  assign f_s_rca32_fa7_xor0 = a[7] ^ b[7];
  assign f_s_rca32_fa7_and0 = a[7] & b[7];
  assign f_s_rca32_fa7_xor1 = f_s_rca32_fa7_xor0 ^ f_s_rca32_fa6_or0;
  assign f_s_rca32_fa7_and1 = f_s_rca32_fa7_xor0 & f_s_rca32_fa6_or0;
  assign f_s_rca32_fa7_or0 = f_s_rca32_fa7_and0 | f_s_rca32_fa7_and1;
  assign f_s_rca32_fa8_xor0 = a[8] ^ b[8];
  assign f_s_rca32_fa8_and0 = a[8] & b[8];
  assign f_s_rca32_fa8_xor1 = f_s_rca32_fa8_xor0 ^ f_s_rca32_fa7_or0;
  assign f_s_rca32_fa8_and1 = f_s_rca32_fa8_xor0 & f_s_rca32_fa7_or0;
  assign f_s_rca32_fa8_or0 = f_s_rca32_fa8_and0 | f_s_rca32_fa8_and1;
  assign f_s_rca32_fa9_xor0 = a[9] ^ b[9];
  assign f_s_rca32_fa9_and0 = a[9] & b[9];
  assign f_s_rca32_fa9_xor1 = f_s_rca32_fa9_xor0 ^ f_s_rca32_fa8_or0;
  assign f_s_rca32_fa9_and1 = f_s_rca32_fa9_xor0 & f_s_rca32_fa8_or0;
  assign f_s_rca32_fa9_or0 = f_s_rca32_fa9_and0 | f_s_rca32_fa9_and1;
  assign f_s_rca32_fa10_xor0 = a[10] ^ b[10];
  assign f_s_rca32_fa10_and0 = a[10] & b[10];
  assign f_s_rca32_fa10_xor1 = f_s_rca32_fa10_xor0 ^ f_s_rca32_fa9_or0;
  assign f_s_rca32_fa10_and1 = f_s_rca32_fa10_xor0 & f_s_rca32_fa9_or0;
  assign f_s_rca32_fa10_or0 = f_s_rca32_fa10_and0 | f_s_rca32_fa10_and1;
  assign f_s_rca32_fa11_xor0 = a[11] ^ b[11];
  assign f_s_rca32_fa11_and0 = a[11] & b[11];
  assign f_s_rca32_fa11_xor1 = f_s_rca32_fa11_xor0 ^ f_s_rca32_fa10_or0;
  assign f_s_rca32_fa11_and1 = f_s_rca32_fa11_xor0 & f_s_rca32_fa10_or0;
  assign f_s_rca32_fa11_or0 = f_s_rca32_fa11_and0 | f_s_rca32_fa11_and1;
  assign f_s_rca32_fa12_xor0 = a[12] ^ b[12];
  assign f_s_rca32_fa12_and0 = a[12] & b[12];
  assign f_s_rca32_fa12_xor1 = f_s_rca32_fa12_xor0 ^ f_s_rca32_fa11_or0;
  assign f_s_rca32_fa12_and1 = f_s_rca32_fa12_xor0 & f_s_rca32_fa11_or0;
  assign f_s_rca32_fa12_or0 = f_s_rca32_fa12_and0 | f_s_rca32_fa12_and1;
  assign f_s_rca32_fa13_xor0 = a[13] ^ b[13];
  assign f_s_rca32_fa13_and0 = a[13] & b[13];
  assign f_s_rca32_fa13_xor1 = f_s_rca32_fa13_xor0 ^ f_s_rca32_fa12_or0;
  assign f_s_rca32_fa13_and1 = f_s_rca32_fa13_xor0 & f_s_rca32_fa12_or0;
  assign f_s_rca32_fa13_or0 = f_s_rca32_fa13_and0 | f_s_rca32_fa13_and1;
  assign f_s_rca32_fa14_xor0 = a[14] ^ b[14];
  assign f_s_rca32_fa14_and0 = a[14] & b[14];
  assign f_s_rca32_fa14_xor1 = f_s_rca32_fa14_xor0 ^ f_s_rca32_fa13_or0;
  assign f_s_rca32_fa14_and1 = f_s_rca32_fa14_xor0 & f_s_rca32_fa13_or0;
  assign f_s_rca32_fa14_or0 = f_s_rca32_fa14_and0 | f_s_rca32_fa14_and1;
  assign f_s_rca32_fa15_xor0 = a[15] ^ b[15];
  assign f_s_rca32_fa15_and0 = a[15] & b[15];
  assign f_s_rca32_fa15_xor1 = f_s_rca32_fa15_xor0 ^ f_s_rca32_fa14_or0;
  assign f_s_rca32_fa15_and1 = f_s_rca32_fa15_xor0 & f_s_rca32_fa14_or0;
  assign f_s_rca32_fa15_or0 = f_s_rca32_fa15_and0 | f_s_rca32_fa15_and1;
  assign f_s_rca32_fa16_xor0 = a[16] ^ b[16];
  assign f_s_rca32_fa16_and0 = a[16] & b[16];
  assign f_s_rca32_fa16_xor1 = f_s_rca32_fa16_xor0 ^ f_s_rca32_fa15_or0;
  assign f_s_rca32_fa16_and1 = f_s_rca32_fa16_xor0 & f_s_rca32_fa15_or0;
  assign f_s_rca32_fa16_or0 = f_s_rca32_fa16_and0 | f_s_rca32_fa16_and1;
  assign f_s_rca32_fa17_xor0 = a[17] ^ b[17];
  assign f_s_rca32_fa17_and0 = a[17] & b[17];
  assign f_s_rca32_fa17_xor1 = f_s_rca32_fa17_xor0 ^ f_s_rca32_fa16_or0;
  assign f_s_rca32_fa17_and1 = f_s_rca32_fa17_xor0 & f_s_rca32_fa16_or0;
  assign f_s_rca32_fa17_or0 = f_s_rca32_fa17_and0 | f_s_rca32_fa17_and1;
  assign f_s_rca32_fa18_xor0 = a[18] ^ b[18];
  assign f_s_rca32_fa18_and0 = a[18] & b[18];
  assign f_s_rca32_fa18_xor1 = f_s_rca32_fa18_xor0 ^ f_s_rca32_fa17_or0;
  assign f_s_rca32_fa18_and1 = f_s_rca32_fa18_xor0 & f_s_rca32_fa17_or0;
  assign f_s_rca32_fa18_or0 = f_s_rca32_fa18_and0 | f_s_rca32_fa18_and1;
  assign f_s_rca32_fa19_xor0 = a[19] ^ b[19];
  assign f_s_rca32_fa19_and0 = a[19] & b[19];
  assign f_s_rca32_fa19_xor1 = f_s_rca32_fa19_xor0 ^ f_s_rca32_fa18_or0;
  assign f_s_rca32_fa19_and1 = f_s_rca32_fa19_xor0 & f_s_rca32_fa18_or0;
  assign f_s_rca32_fa19_or0 = f_s_rca32_fa19_and0 | f_s_rca32_fa19_and1;
  assign f_s_rca32_fa20_xor0 = a[20] ^ b[20];
  assign f_s_rca32_fa20_and0 = a[20] & b[20];
  assign f_s_rca32_fa20_xor1 = f_s_rca32_fa20_xor0 ^ f_s_rca32_fa19_or0;
  assign f_s_rca32_fa20_and1 = f_s_rca32_fa20_xor0 & f_s_rca32_fa19_or0;
  assign f_s_rca32_fa20_or0 = f_s_rca32_fa20_and0 | f_s_rca32_fa20_and1;
  assign f_s_rca32_fa21_xor0 = a[21] ^ b[21];
  assign f_s_rca32_fa21_and0 = a[21] & b[21];
  assign f_s_rca32_fa21_xor1 = f_s_rca32_fa21_xor0 ^ f_s_rca32_fa20_or0;
  assign f_s_rca32_fa21_and1 = f_s_rca32_fa21_xor0 & f_s_rca32_fa20_or0;
  assign f_s_rca32_fa21_or0 = f_s_rca32_fa21_and0 | f_s_rca32_fa21_and1;
  assign f_s_rca32_fa22_xor0 = a[22] ^ b[22];
  assign f_s_rca32_fa22_and0 = a[22] & b[22];
  assign f_s_rca32_fa22_xor1 = f_s_rca32_fa22_xor0 ^ f_s_rca32_fa21_or0;
  assign f_s_rca32_fa22_and1 = f_s_rca32_fa22_xor0 & f_s_rca32_fa21_or0;
  assign f_s_rca32_fa22_or0 = f_s_rca32_fa22_and0 | f_s_rca32_fa22_and1;
  assign f_s_rca32_fa23_xor0 = a[23] ^ b[23];
  assign f_s_rca32_fa23_and0 = a[23] & b[23];
  assign f_s_rca32_fa23_xor1 = f_s_rca32_fa23_xor0 ^ f_s_rca32_fa22_or0;
  assign f_s_rca32_fa23_and1 = f_s_rca32_fa23_xor0 & f_s_rca32_fa22_or0;
  assign f_s_rca32_fa23_or0 = f_s_rca32_fa23_and0 | f_s_rca32_fa23_and1;
  assign f_s_rca32_fa24_xor0 = a[24] ^ b[24];
  assign f_s_rca32_fa24_and0 = a[24] & b[24];
  assign f_s_rca32_fa24_xor1 = f_s_rca32_fa24_xor0 ^ f_s_rca32_fa23_or0;
  assign f_s_rca32_fa24_and1 = f_s_rca32_fa24_xor0 & f_s_rca32_fa23_or0;
  assign f_s_rca32_fa24_or0 = f_s_rca32_fa24_and0 | f_s_rca32_fa24_and1;
  assign f_s_rca32_fa25_xor0 = a[25] ^ b[25];
  assign f_s_rca32_fa25_and0 = a[25] & b[25];
  assign f_s_rca32_fa25_xor1 = f_s_rca32_fa25_xor0 ^ f_s_rca32_fa24_or0;
  assign f_s_rca32_fa25_and1 = f_s_rca32_fa25_xor0 & f_s_rca32_fa24_or0;
  assign f_s_rca32_fa25_or0 = f_s_rca32_fa25_and0 | f_s_rca32_fa25_and1;
  assign f_s_rca32_fa26_xor0 = a[26] ^ b[26];
  assign f_s_rca32_fa26_and0 = a[26] & b[26];
  assign f_s_rca32_fa26_xor1 = f_s_rca32_fa26_xor0 ^ f_s_rca32_fa25_or0;
  assign f_s_rca32_fa26_and1 = f_s_rca32_fa26_xor0 & f_s_rca32_fa25_or0;
  assign f_s_rca32_fa26_or0 = f_s_rca32_fa26_and0 | f_s_rca32_fa26_and1;
  assign f_s_rca32_fa27_xor0 = a[27] ^ b[27];
  assign f_s_rca32_fa27_and0 = a[27] & b[27];
  assign f_s_rca32_fa27_xor1 = f_s_rca32_fa27_xor0 ^ f_s_rca32_fa26_or0;
  assign f_s_rca32_fa27_and1 = f_s_rca32_fa27_xor0 & f_s_rca32_fa26_or0;
  assign f_s_rca32_fa27_or0 = f_s_rca32_fa27_and0 | f_s_rca32_fa27_and1;
  assign f_s_rca32_fa28_xor0 = a[28] ^ b[28];
  assign f_s_rca32_fa28_and0 = a[28] & b[28];
  assign f_s_rca32_fa28_xor1 = f_s_rca32_fa28_xor0 ^ f_s_rca32_fa27_or0;
  assign f_s_rca32_fa28_and1 = f_s_rca32_fa28_xor0 & f_s_rca32_fa27_or0;
  assign f_s_rca32_fa28_or0 = f_s_rca32_fa28_and0 | f_s_rca32_fa28_and1;
  assign f_s_rca32_fa29_xor0 = a[29] ^ b[29];
  assign f_s_rca32_fa29_and0 = a[29] & b[29];
  assign f_s_rca32_fa29_xor1 = f_s_rca32_fa29_xor0 ^ f_s_rca32_fa28_or0;
  assign f_s_rca32_fa29_and1 = f_s_rca32_fa29_xor0 & f_s_rca32_fa28_or0;
  assign f_s_rca32_fa29_or0 = f_s_rca32_fa29_and0 | f_s_rca32_fa29_and1;
  assign f_s_rca32_fa30_xor0 = a[30] ^ b[30];
  assign f_s_rca32_fa30_and0 = a[30] & b[30];
  assign f_s_rca32_fa30_xor1 = f_s_rca32_fa30_xor0 ^ f_s_rca32_fa29_or0;
  assign f_s_rca32_fa30_and1 = f_s_rca32_fa30_xor0 & f_s_rca32_fa29_or0;
  assign f_s_rca32_fa30_or0 = f_s_rca32_fa30_and0 | f_s_rca32_fa30_and1;
  assign f_s_rca32_fa31_xor0 = a[31] ^ b[31];
  assign f_s_rca32_fa31_and0 = a[31] & b[31];
  assign f_s_rca32_fa31_xor1 = f_s_rca32_fa31_xor0 ^ f_s_rca32_fa30_or0;
  assign f_s_rca32_fa31_and1 = f_s_rca32_fa31_xor0 & f_s_rca32_fa30_or0;
  assign f_s_rca32_fa31_or0 = f_s_rca32_fa31_and0 | f_s_rca32_fa31_and1;
  assign f_s_rca32_xor0 = a[31] ^ b[31];
  assign f_s_rca32_xor1 = f_s_rca32_xor0 ^ f_s_rca32_fa31_or0;

  assign f_s_rca32_out[0] = f_s_rca32_ha_xor0;
  assign f_s_rca32_out[1] = f_s_rca32_fa1_xor1;
  assign f_s_rca32_out[2] = f_s_rca32_fa2_xor1;
  assign f_s_rca32_out[3] = f_s_rca32_fa3_xor1;
  assign f_s_rca32_out[4] = f_s_rca32_fa4_xor1;
  assign f_s_rca32_out[5] = f_s_rca32_fa5_xor1;
  assign f_s_rca32_out[6] = f_s_rca32_fa6_xor1;
  assign f_s_rca32_out[7] = f_s_rca32_fa7_xor1;
  assign f_s_rca32_out[8] = f_s_rca32_fa8_xor1;
  assign f_s_rca32_out[9] = f_s_rca32_fa9_xor1;
  assign f_s_rca32_out[10] = f_s_rca32_fa10_xor1;
  assign f_s_rca32_out[11] = f_s_rca32_fa11_xor1;
  assign f_s_rca32_out[12] = f_s_rca32_fa12_xor1;
  assign f_s_rca32_out[13] = f_s_rca32_fa13_xor1;
  assign f_s_rca32_out[14] = f_s_rca32_fa14_xor1;
  assign f_s_rca32_out[15] = f_s_rca32_fa15_xor1;
  assign f_s_rca32_out[16] = f_s_rca32_fa16_xor1;
  assign f_s_rca32_out[17] = f_s_rca32_fa17_xor1;
  assign f_s_rca32_out[18] = f_s_rca32_fa18_xor1;
  assign f_s_rca32_out[19] = f_s_rca32_fa19_xor1;
  assign f_s_rca32_out[20] = f_s_rca32_fa20_xor1;
  assign f_s_rca32_out[21] = f_s_rca32_fa21_xor1;
  assign f_s_rca32_out[22] = f_s_rca32_fa22_xor1;
  assign f_s_rca32_out[23] = f_s_rca32_fa23_xor1;
  assign f_s_rca32_out[24] = f_s_rca32_fa24_xor1;
  assign f_s_rca32_out[25] = f_s_rca32_fa25_xor1;
  assign f_s_rca32_out[26] = f_s_rca32_fa26_xor1;
  assign f_s_rca32_out[27] = f_s_rca32_fa27_xor1;
  assign f_s_rca32_out[28] = f_s_rca32_fa28_xor1;
  assign f_s_rca32_out[29] = f_s_rca32_fa29_xor1;
  assign f_s_rca32_out[30] = f_s_rca32_fa30_xor1;
  assign f_s_rca32_out[31] = f_s_rca32_fa31_xor1;
  assign f_s_rca32_out[32] = f_s_rca32_xor1;
endmodule