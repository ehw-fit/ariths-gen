module s_dadda_cla12(input [11:0] a, input [11:0] b, output [23:0] s_dadda_cla12_out);
  wire s_dadda_cla12_and_9_0;
  wire s_dadda_cla12_and_8_1;
  wire s_dadda_cla12_ha0_xor0;
  wire s_dadda_cla12_ha0_and0;
  wire s_dadda_cla12_and_10_0;
  wire s_dadda_cla12_and_9_1;
  wire s_dadda_cla12_fa0_xor0;
  wire s_dadda_cla12_fa0_and0;
  wire s_dadda_cla12_fa0_xor1;
  wire s_dadda_cla12_fa0_and1;
  wire s_dadda_cla12_fa0_or0;
  wire s_dadda_cla12_and_8_2;
  wire s_dadda_cla12_and_7_3;
  wire s_dadda_cla12_ha1_xor0;
  wire s_dadda_cla12_ha1_and0;
  wire s_dadda_cla12_nand_11_0;
  wire s_dadda_cla12_fa1_xor0;
  wire s_dadda_cla12_fa1_and0;
  wire s_dadda_cla12_fa1_xor1;
  wire s_dadda_cla12_fa1_and1;
  wire s_dadda_cla12_fa1_or0;
  wire s_dadda_cla12_and_10_1;
  wire s_dadda_cla12_and_9_2;
  wire s_dadda_cla12_and_8_3;
  wire s_dadda_cla12_fa2_xor0;
  wire s_dadda_cla12_fa2_and0;
  wire s_dadda_cla12_fa2_xor1;
  wire s_dadda_cla12_fa2_and1;
  wire s_dadda_cla12_fa2_or0;
  wire s_dadda_cla12_and_7_4;
  wire s_dadda_cla12_and_6_5;
  wire s_dadda_cla12_ha2_xor0;
  wire s_dadda_cla12_ha2_and0;
  wire s_dadda_cla12_fa3_xor0;
  wire s_dadda_cla12_fa3_and0;
  wire s_dadda_cla12_fa3_xor1;
  wire s_dadda_cla12_fa3_and1;
  wire s_dadda_cla12_fa3_or0;
  wire s_dadda_cla12_nand_11_1;
  wire s_dadda_cla12_and_10_2;
  wire s_dadda_cla12_fa4_xor0;
  wire s_dadda_cla12_fa4_xor1;
  wire s_dadda_cla12_fa4_and1;
  wire s_dadda_cla12_fa4_or0;
  wire s_dadda_cla12_and_9_3;
  wire s_dadda_cla12_and_8_4;
  wire s_dadda_cla12_and_7_5;
  wire s_dadda_cla12_fa5_xor0;
  wire s_dadda_cla12_fa5_and0;
  wire s_dadda_cla12_fa5_xor1;
  wire s_dadda_cla12_fa5_and1;
  wire s_dadda_cla12_fa5_or0;
  wire s_dadda_cla12_fa6_xor0;
  wire s_dadda_cla12_fa6_and0;
  wire s_dadda_cla12_fa6_xor1;
  wire s_dadda_cla12_fa6_and1;
  wire s_dadda_cla12_fa6_or0;
  wire s_dadda_cla12_nand_11_2;
  wire s_dadda_cla12_and_10_3;
  wire s_dadda_cla12_and_9_4;
  wire s_dadda_cla12_fa7_xor0;
  wire s_dadda_cla12_fa7_and0;
  wire s_dadda_cla12_fa7_xor1;
  wire s_dadda_cla12_fa7_and1;
  wire s_dadda_cla12_fa7_or0;
  wire s_dadda_cla12_nand_11_3;
  wire s_dadda_cla12_fa8_xor0;
  wire s_dadda_cla12_fa8_and0;
  wire s_dadda_cla12_fa8_xor1;
  wire s_dadda_cla12_fa8_and1;
  wire s_dadda_cla12_fa8_or0;
  wire s_dadda_cla12_and_4_0;
  wire s_dadda_cla12_and_3_1;
  wire s_dadda_cla12_ha3_xor0;
  wire s_dadda_cla12_ha3_and0;
  wire s_dadda_cla12_and_5_0;
  wire s_dadda_cla12_and_4_1;
  wire s_dadda_cla12_fa9_xor0;
  wire s_dadda_cla12_fa9_and0;
  wire s_dadda_cla12_fa9_xor1;
  wire s_dadda_cla12_fa9_and1;
  wire s_dadda_cla12_fa9_or0;
  wire s_dadda_cla12_and_3_2;
  wire s_dadda_cla12_and_2_3;
  wire s_dadda_cla12_ha4_xor0;
  wire s_dadda_cla12_ha4_and0;
  wire s_dadda_cla12_and_6_0;
  wire s_dadda_cla12_fa10_xor0;
  wire s_dadda_cla12_fa10_and0;
  wire s_dadda_cla12_fa10_xor1;
  wire s_dadda_cla12_fa10_and1;
  wire s_dadda_cla12_fa10_or0;
  wire s_dadda_cla12_and_5_1;
  wire s_dadda_cla12_and_4_2;
  wire s_dadda_cla12_and_3_3;
  wire s_dadda_cla12_fa11_xor0;
  wire s_dadda_cla12_fa11_and0;
  wire s_dadda_cla12_fa11_xor1;
  wire s_dadda_cla12_fa11_and1;
  wire s_dadda_cla12_fa11_or0;
  wire s_dadda_cla12_and_2_4;
  wire s_dadda_cla12_and_1_5;
  wire s_dadda_cla12_ha5_xor0;
  wire s_dadda_cla12_ha5_and0;
  wire s_dadda_cla12_fa12_xor0;
  wire s_dadda_cla12_fa12_and0;
  wire s_dadda_cla12_fa12_xor1;
  wire s_dadda_cla12_fa12_and1;
  wire s_dadda_cla12_fa12_or0;
  wire s_dadda_cla12_and_7_0;
  wire s_dadda_cla12_and_6_1;
  wire s_dadda_cla12_and_5_2;
  wire s_dadda_cla12_fa13_xor0;
  wire s_dadda_cla12_fa13_and0;
  wire s_dadda_cla12_fa13_xor1;
  wire s_dadda_cla12_fa13_and1;
  wire s_dadda_cla12_fa13_or0;
  wire s_dadda_cla12_and_4_3;
  wire s_dadda_cla12_and_3_4;
  wire s_dadda_cla12_and_2_5;
  wire s_dadda_cla12_fa14_xor0;
  wire s_dadda_cla12_fa14_and0;
  wire s_dadda_cla12_fa14_xor1;
  wire s_dadda_cla12_fa14_and1;
  wire s_dadda_cla12_fa14_or0;
  wire s_dadda_cla12_and_1_6;
  wire s_dadda_cla12_and_0_7;
  wire s_dadda_cla12_ha6_xor0;
  wire s_dadda_cla12_ha6_and0;
  wire s_dadda_cla12_fa15_xor0;
  wire s_dadda_cla12_fa15_and0;
  wire s_dadda_cla12_fa15_xor1;
  wire s_dadda_cla12_fa15_and1;
  wire s_dadda_cla12_fa15_or0;
  wire s_dadda_cla12_and_8_0;
  wire s_dadda_cla12_and_7_1;
  wire s_dadda_cla12_fa16_xor0;
  wire s_dadda_cla12_fa16_and0;
  wire s_dadda_cla12_fa16_xor1;
  wire s_dadda_cla12_fa16_and1;
  wire s_dadda_cla12_fa16_or0;
  wire s_dadda_cla12_and_6_2;
  wire s_dadda_cla12_and_5_3;
  wire s_dadda_cla12_and_4_4;
  wire s_dadda_cla12_fa17_xor0;
  wire s_dadda_cla12_fa17_and0;
  wire s_dadda_cla12_fa17_xor1;
  wire s_dadda_cla12_fa17_and1;
  wire s_dadda_cla12_fa17_or0;
  wire s_dadda_cla12_and_3_5;
  wire s_dadda_cla12_and_2_6;
  wire s_dadda_cla12_and_1_7;
  wire s_dadda_cla12_fa18_xor0;
  wire s_dadda_cla12_fa18_and0;
  wire s_dadda_cla12_fa18_xor1;
  wire s_dadda_cla12_fa18_and1;
  wire s_dadda_cla12_fa18_or0;
  wire s_dadda_cla12_and_0_8;
  wire s_dadda_cla12_ha7_xor0;
  wire s_dadda_cla12_ha7_and0;
  wire s_dadda_cla12_fa19_xor0;
  wire s_dadda_cla12_fa19_and0;
  wire s_dadda_cla12_fa19_xor1;
  wire s_dadda_cla12_fa19_and1;
  wire s_dadda_cla12_fa19_or0;
  wire s_dadda_cla12_and_7_2;
  wire s_dadda_cla12_fa20_xor0;
  wire s_dadda_cla12_fa20_and0;
  wire s_dadda_cla12_fa20_xor1;
  wire s_dadda_cla12_fa20_and1;
  wire s_dadda_cla12_fa20_or0;
  wire s_dadda_cla12_and_6_3;
  wire s_dadda_cla12_and_5_4;
  wire s_dadda_cla12_and_4_5;
  wire s_dadda_cla12_fa21_xor0;
  wire s_dadda_cla12_fa21_and0;
  wire s_dadda_cla12_fa21_xor1;
  wire s_dadda_cla12_fa21_and1;
  wire s_dadda_cla12_fa21_or0;
  wire s_dadda_cla12_and_3_6;
  wire s_dadda_cla12_and_2_7;
  wire s_dadda_cla12_and_1_8;
  wire s_dadda_cla12_fa22_xor0;
  wire s_dadda_cla12_fa22_and0;
  wire s_dadda_cla12_fa22_xor1;
  wire s_dadda_cla12_fa22_and1;
  wire s_dadda_cla12_fa22_or0;
  wire s_dadda_cla12_and_0_9;
  wire s_dadda_cla12_fa23_xor0;
  wire s_dadda_cla12_fa23_and0;
  wire s_dadda_cla12_fa23_xor1;
  wire s_dadda_cla12_fa23_and1;
  wire s_dadda_cla12_fa23_or0;
  wire s_dadda_cla12_fa24_xor0;
  wire s_dadda_cla12_fa24_and0;
  wire s_dadda_cla12_fa24_xor1;
  wire s_dadda_cla12_fa24_and1;
  wire s_dadda_cla12_fa24_or0;
  wire s_dadda_cla12_and_6_4;
  wire s_dadda_cla12_fa25_xor0;
  wire s_dadda_cla12_fa25_and0;
  wire s_dadda_cla12_fa25_xor1;
  wire s_dadda_cla12_fa25_and1;
  wire s_dadda_cla12_fa25_or0;
  wire s_dadda_cla12_and_5_5;
  wire s_dadda_cla12_and_4_6;
  wire s_dadda_cla12_and_3_7;
  wire s_dadda_cla12_fa26_xor0;
  wire s_dadda_cla12_fa26_and0;
  wire s_dadda_cla12_fa26_xor1;
  wire s_dadda_cla12_fa26_and1;
  wire s_dadda_cla12_fa26_or0;
  wire s_dadda_cla12_and_2_8;
  wire s_dadda_cla12_and_1_9;
  wire s_dadda_cla12_and_0_10;
  wire s_dadda_cla12_fa27_xor0;
  wire s_dadda_cla12_fa27_and0;
  wire s_dadda_cla12_fa27_xor1;
  wire s_dadda_cla12_fa27_and1;
  wire s_dadda_cla12_fa27_or0;
  wire s_dadda_cla12_fa28_xor0;
  wire s_dadda_cla12_fa28_and0;
  wire s_dadda_cla12_fa28_xor1;
  wire s_dadda_cla12_fa28_and1;
  wire s_dadda_cla12_fa28_or0;
  wire s_dadda_cla12_fa29_xor0;
  wire s_dadda_cla12_fa29_and0;
  wire s_dadda_cla12_fa29_xor1;
  wire s_dadda_cla12_fa29_and1;
  wire s_dadda_cla12_fa29_or0;
  wire s_dadda_cla12_and_5_6;
  wire s_dadda_cla12_fa30_xor0;
  wire s_dadda_cla12_fa30_and0;
  wire s_dadda_cla12_fa30_xor1;
  wire s_dadda_cla12_fa30_and1;
  wire s_dadda_cla12_fa30_or0;
  wire s_dadda_cla12_and_4_7;
  wire s_dadda_cla12_and_3_8;
  wire s_dadda_cla12_and_2_9;
  wire s_dadda_cla12_fa31_xor0;
  wire s_dadda_cla12_fa31_and0;
  wire s_dadda_cla12_fa31_xor1;
  wire s_dadda_cla12_fa31_and1;
  wire s_dadda_cla12_fa31_or0;
  wire s_dadda_cla12_and_1_10;
  wire s_dadda_cla12_nand_0_11;
  wire s_dadda_cla12_fa32_xor0;
  wire s_dadda_cla12_fa32_and0;
  wire s_dadda_cla12_fa32_xor1;
  wire s_dadda_cla12_fa32_and1;
  wire s_dadda_cla12_fa32_or0;
  wire s_dadda_cla12_fa33_xor0;
  wire s_dadda_cla12_fa33_and0;
  wire s_dadda_cla12_fa33_xor1;
  wire s_dadda_cla12_fa33_and1;
  wire s_dadda_cla12_fa33_or0;
  wire s_dadda_cla12_fa34_xor0;
  wire s_dadda_cla12_fa34_and0;
  wire s_dadda_cla12_fa34_xor1;
  wire s_dadda_cla12_fa34_and1;
  wire s_dadda_cla12_fa34_or0;
  wire s_dadda_cla12_and_6_6;
  wire s_dadda_cla12_fa35_xor0;
  wire s_dadda_cla12_fa35_and0;
  wire s_dadda_cla12_fa35_xor1;
  wire s_dadda_cla12_fa35_and1;
  wire s_dadda_cla12_fa35_or0;
  wire s_dadda_cla12_and_5_7;
  wire s_dadda_cla12_and_4_8;
  wire s_dadda_cla12_and_3_9;
  wire s_dadda_cla12_fa36_xor0;
  wire s_dadda_cla12_fa36_and0;
  wire s_dadda_cla12_fa36_xor1;
  wire s_dadda_cla12_fa36_and1;
  wire s_dadda_cla12_fa36_or0;
  wire s_dadda_cla12_and_2_10;
  wire s_dadda_cla12_nand_1_11;
  wire s_dadda_cla12_fa37_xor0;
  wire s_dadda_cla12_fa37_and0;
  wire s_dadda_cla12_fa37_xor1;
  wire s_dadda_cla12_fa37_and1;
  wire s_dadda_cla12_fa37_or0;
  wire s_dadda_cla12_fa38_xor0;
  wire s_dadda_cla12_fa38_and0;
  wire s_dadda_cla12_fa38_xor1;
  wire s_dadda_cla12_fa38_and1;
  wire s_dadda_cla12_fa38_or0;
  wire s_dadda_cla12_fa39_xor0;
  wire s_dadda_cla12_fa39_and0;
  wire s_dadda_cla12_fa39_xor1;
  wire s_dadda_cla12_fa39_and1;
  wire s_dadda_cla12_fa39_or0;
  wire s_dadda_cla12_and_8_5;
  wire s_dadda_cla12_fa40_xor0;
  wire s_dadda_cla12_fa40_and0;
  wire s_dadda_cla12_fa40_xor1;
  wire s_dadda_cla12_fa40_and1;
  wire s_dadda_cla12_fa40_or0;
  wire s_dadda_cla12_and_7_6;
  wire s_dadda_cla12_and_6_7;
  wire s_dadda_cla12_and_5_8;
  wire s_dadda_cla12_fa41_xor0;
  wire s_dadda_cla12_fa41_and0;
  wire s_dadda_cla12_fa41_xor1;
  wire s_dadda_cla12_fa41_and1;
  wire s_dadda_cla12_fa41_or0;
  wire s_dadda_cla12_and_4_9;
  wire s_dadda_cla12_and_3_10;
  wire s_dadda_cla12_nand_2_11;
  wire s_dadda_cla12_fa42_xor0;
  wire s_dadda_cla12_fa42_and0;
  wire s_dadda_cla12_fa42_xor1;
  wire s_dadda_cla12_fa42_and1;
  wire s_dadda_cla12_fa42_or0;
  wire s_dadda_cla12_fa43_xor0;
  wire s_dadda_cla12_fa43_and0;
  wire s_dadda_cla12_fa43_xor1;
  wire s_dadda_cla12_fa43_and1;
  wire s_dadda_cla12_fa43_or0;
  wire s_dadda_cla12_fa44_xor0;
  wire s_dadda_cla12_fa44_and0;
  wire s_dadda_cla12_fa44_xor1;
  wire s_dadda_cla12_fa44_and1;
  wire s_dadda_cla12_fa44_or0;
  wire s_dadda_cla12_and_10_4;
  wire s_dadda_cla12_fa45_xor0;
  wire s_dadda_cla12_fa45_and0;
  wire s_dadda_cla12_fa45_xor1;
  wire s_dadda_cla12_fa45_and1;
  wire s_dadda_cla12_fa45_or0;
  wire s_dadda_cla12_and_9_5;
  wire s_dadda_cla12_and_8_6;
  wire s_dadda_cla12_and_7_7;
  wire s_dadda_cla12_fa46_xor0;
  wire s_dadda_cla12_fa46_and0;
  wire s_dadda_cla12_fa46_xor1;
  wire s_dadda_cla12_fa46_and1;
  wire s_dadda_cla12_fa46_or0;
  wire s_dadda_cla12_and_6_8;
  wire s_dadda_cla12_and_5_9;
  wire s_dadda_cla12_and_4_10;
  wire s_dadda_cla12_fa47_xor0;
  wire s_dadda_cla12_fa47_and0;
  wire s_dadda_cla12_fa47_xor1;
  wire s_dadda_cla12_fa47_and1;
  wire s_dadda_cla12_fa47_or0;
  wire s_dadda_cla12_nand_3_11;
  wire s_dadda_cla12_fa48_xor0;
  wire s_dadda_cla12_fa48_and0;
  wire s_dadda_cla12_fa48_xor1;
  wire s_dadda_cla12_fa48_and1;
  wire s_dadda_cla12_fa48_or0;
  wire s_dadda_cla12_fa49_xor0;
  wire s_dadda_cla12_fa49_and0;
  wire s_dadda_cla12_fa49_xor1;
  wire s_dadda_cla12_fa49_and1;
  wire s_dadda_cla12_fa49_or0;
  wire s_dadda_cla12_fa50_xor0;
  wire s_dadda_cla12_fa50_and0;
  wire s_dadda_cla12_fa50_xor1;
  wire s_dadda_cla12_fa50_and1;
  wire s_dadda_cla12_fa50_or0;
  wire s_dadda_cla12_nand_11_4;
  wire s_dadda_cla12_and_10_5;
  wire s_dadda_cla12_and_9_6;
  wire s_dadda_cla12_fa51_xor0;
  wire s_dadda_cla12_fa51_and0;
  wire s_dadda_cla12_fa51_xor1;
  wire s_dadda_cla12_fa51_and1;
  wire s_dadda_cla12_fa51_or0;
  wire s_dadda_cla12_and_8_7;
  wire s_dadda_cla12_and_7_8;
  wire s_dadda_cla12_and_6_9;
  wire s_dadda_cla12_fa52_xor0;
  wire s_dadda_cla12_fa52_and0;
  wire s_dadda_cla12_fa52_xor1;
  wire s_dadda_cla12_fa52_and1;
  wire s_dadda_cla12_fa52_or0;
  wire s_dadda_cla12_and_5_10;
  wire s_dadda_cla12_nand_4_11;
  wire s_dadda_cla12_fa53_xor0;
  wire s_dadda_cla12_fa53_and0;
  wire s_dadda_cla12_fa53_xor1;
  wire s_dadda_cla12_fa53_and1;
  wire s_dadda_cla12_fa53_or0;
  wire s_dadda_cla12_fa54_xor0;
  wire s_dadda_cla12_fa54_and0;
  wire s_dadda_cla12_fa54_xor1;
  wire s_dadda_cla12_fa54_and1;
  wire s_dadda_cla12_fa54_or0;
  wire s_dadda_cla12_nand_11_5;
  wire s_dadda_cla12_fa55_xor0;
  wire s_dadda_cla12_fa55_and0;
  wire s_dadda_cla12_fa55_xor1;
  wire s_dadda_cla12_fa55_and1;
  wire s_dadda_cla12_fa55_or0;
  wire s_dadda_cla12_and_10_6;
  wire s_dadda_cla12_and_9_7;
  wire s_dadda_cla12_and_8_8;
  wire s_dadda_cla12_fa56_xor0;
  wire s_dadda_cla12_fa56_and0;
  wire s_dadda_cla12_fa56_xor1;
  wire s_dadda_cla12_fa56_and1;
  wire s_dadda_cla12_fa56_or0;
  wire s_dadda_cla12_and_7_9;
  wire s_dadda_cla12_and_6_10;
  wire s_dadda_cla12_nand_5_11;
  wire s_dadda_cla12_fa57_xor0;
  wire s_dadda_cla12_fa57_and0;
  wire s_dadda_cla12_fa57_xor1;
  wire s_dadda_cla12_fa57_and1;
  wire s_dadda_cla12_fa57_or0;
  wire s_dadda_cla12_fa58_xor0;
  wire s_dadda_cla12_fa58_and0;
  wire s_dadda_cla12_fa58_xor1;
  wire s_dadda_cla12_fa58_and1;
  wire s_dadda_cla12_fa58_or0;
  wire s_dadda_cla12_nand_11_6;
  wire s_dadda_cla12_and_10_7;
  wire s_dadda_cla12_fa59_xor0;
  wire s_dadda_cla12_fa59_and0;
  wire s_dadda_cla12_fa59_xor1;
  wire s_dadda_cla12_fa59_and1;
  wire s_dadda_cla12_fa59_or0;
  wire s_dadda_cla12_and_9_8;
  wire s_dadda_cla12_and_8_9;
  wire s_dadda_cla12_and_7_10;
  wire s_dadda_cla12_fa60_xor0;
  wire s_dadda_cla12_fa60_and0;
  wire s_dadda_cla12_fa60_xor1;
  wire s_dadda_cla12_fa60_and1;
  wire s_dadda_cla12_fa60_or0;
  wire s_dadda_cla12_fa61_xor0;
  wire s_dadda_cla12_fa61_and0;
  wire s_dadda_cla12_fa61_xor1;
  wire s_dadda_cla12_fa61_and1;
  wire s_dadda_cla12_fa61_or0;
  wire s_dadda_cla12_nand_11_7;
  wire s_dadda_cla12_and_10_8;
  wire s_dadda_cla12_and_9_9;
  wire s_dadda_cla12_fa62_xor0;
  wire s_dadda_cla12_fa62_and0;
  wire s_dadda_cla12_fa62_xor1;
  wire s_dadda_cla12_fa62_and1;
  wire s_dadda_cla12_fa62_or0;
  wire s_dadda_cla12_nand_11_8;
  wire s_dadda_cla12_fa63_xor0;
  wire s_dadda_cla12_fa63_and0;
  wire s_dadda_cla12_fa63_xor1;
  wire s_dadda_cla12_fa63_and1;
  wire s_dadda_cla12_fa63_or0;
  wire s_dadda_cla12_and_3_0;
  wire s_dadda_cla12_and_2_1;
  wire s_dadda_cla12_ha8_xor0;
  wire s_dadda_cla12_ha8_and0;
  wire s_dadda_cla12_and_2_2;
  wire s_dadda_cla12_and_1_3;
  wire s_dadda_cla12_fa64_xor0;
  wire s_dadda_cla12_fa64_and0;
  wire s_dadda_cla12_fa64_xor1;
  wire s_dadda_cla12_fa64_and1;
  wire s_dadda_cla12_fa64_or0;
  wire s_dadda_cla12_and_1_4;
  wire s_dadda_cla12_and_0_5;
  wire s_dadda_cla12_fa65_xor0;
  wire s_dadda_cla12_fa65_and0;
  wire s_dadda_cla12_fa65_xor1;
  wire s_dadda_cla12_fa65_and1;
  wire s_dadda_cla12_fa65_or0;
  wire s_dadda_cla12_and_0_6;
  wire s_dadda_cla12_fa66_xor0;
  wire s_dadda_cla12_fa66_and0;
  wire s_dadda_cla12_fa66_xor1;
  wire s_dadda_cla12_fa66_and1;
  wire s_dadda_cla12_fa66_or0;
  wire s_dadda_cla12_fa67_xor0;
  wire s_dadda_cla12_fa67_and0;
  wire s_dadda_cla12_fa67_xor1;
  wire s_dadda_cla12_fa67_and1;
  wire s_dadda_cla12_fa67_or0;
  wire s_dadda_cla12_fa68_xor0;
  wire s_dadda_cla12_fa68_and0;
  wire s_dadda_cla12_fa68_xor1;
  wire s_dadda_cla12_fa68_and1;
  wire s_dadda_cla12_fa68_or0;
  wire s_dadda_cla12_fa69_xor0;
  wire s_dadda_cla12_fa69_and0;
  wire s_dadda_cla12_fa69_xor1;
  wire s_dadda_cla12_fa69_and1;
  wire s_dadda_cla12_fa69_or0;
  wire s_dadda_cla12_fa70_xor0;
  wire s_dadda_cla12_fa70_and0;
  wire s_dadda_cla12_fa70_xor1;
  wire s_dadda_cla12_fa70_and1;
  wire s_dadda_cla12_fa70_or0;
  wire s_dadda_cla12_fa71_xor0;
  wire s_dadda_cla12_fa71_and0;
  wire s_dadda_cla12_fa71_xor1;
  wire s_dadda_cla12_fa71_and1;
  wire s_dadda_cla12_fa71_or0;
  wire s_dadda_cla12_fa72_xor0;
  wire s_dadda_cla12_fa72_and0;
  wire s_dadda_cla12_fa72_xor1;
  wire s_dadda_cla12_fa72_and1;
  wire s_dadda_cla12_fa72_or0;
  wire s_dadda_cla12_fa73_xor0;
  wire s_dadda_cla12_fa73_and0;
  wire s_dadda_cla12_fa73_xor1;
  wire s_dadda_cla12_fa73_and1;
  wire s_dadda_cla12_fa73_or0;
  wire s_dadda_cla12_fa74_xor0;
  wire s_dadda_cla12_fa74_and0;
  wire s_dadda_cla12_fa74_xor1;
  wire s_dadda_cla12_fa74_and1;
  wire s_dadda_cla12_fa74_or0;
  wire s_dadda_cla12_fa75_xor0;
  wire s_dadda_cla12_fa75_and0;
  wire s_dadda_cla12_fa75_xor1;
  wire s_dadda_cla12_fa75_and1;
  wire s_dadda_cla12_fa75_or0;
  wire s_dadda_cla12_fa76_xor0;
  wire s_dadda_cla12_fa76_and0;
  wire s_dadda_cla12_fa76_xor1;
  wire s_dadda_cla12_fa76_and1;
  wire s_dadda_cla12_fa76_or0;
  wire s_dadda_cla12_nand_6_11;
  wire s_dadda_cla12_fa77_xor0;
  wire s_dadda_cla12_fa77_and0;
  wire s_dadda_cla12_fa77_xor1;
  wire s_dadda_cla12_fa77_and1;
  wire s_dadda_cla12_fa77_or0;
  wire s_dadda_cla12_and_8_10;
  wire s_dadda_cla12_nand_7_11;
  wire s_dadda_cla12_fa78_xor0;
  wire s_dadda_cla12_fa78_and0;
  wire s_dadda_cla12_fa78_xor1;
  wire s_dadda_cla12_fa78_and1;
  wire s_dadda_cla12_fa78_or0;
  wire s_dadda_cla12_and_10_9;
  wire s_dadda_cla12_and_9_10;
  wire s_dadda_cla12_fa79_xor0;
  wire s_dadda_cla12_fa79_and0;
  wire s_dadda_cla12_fa79_xor1;
  wire s_dadda_cla12_fa79_and1;
  wire s_dadda_cla12_fa79_or0;
  wire s_dadda_cla12_nand_11_9;
  wire s_dadda_cla12_fa80_xor0;
  wire s_dadda_cla12_fa80_and0;
  wire s_dadda_cla12_fa80_xor1;
  wire s_dadda_cla12_fa80_and1;
  wire s_dadda_cla12_fa80_or0;
  wire s_dadda_cla12_and_2_0;
  wire s_dadda_cla12_and_1_1;
  wire s_dadda_cla12_ha9_xor0;
  wire s_dadda_cla12_ha9_and0;
  wire s_dadda_cla12_and_1_2;
  wire s_dadda_cla12_and_0_3;
  wire s_dadda_cla12_fa81_xor0;
  wire s_dadda_cla12_fa81_and0;
  wire s_dadda_cla12_fa81_xor1;
  wire s_dadda_cla12_fa81_and1;
  wire s_dadda_cla12_fa81_or0;
  wire s_dadda_cla12_and_0_4;
  wire s_dadda_cla12_fa82_xor0;
  wire s_dadda_cla12_fa82_and0;
  wire s_dadda_cla12_fa82_xor1;
  wire s_dadda_cla12_fa82_and1;
  wire s_dadda_cla12_fa82_or0;
  wire s_dadda_cla12_fa83_xor0;
  wire s_dadda_cla12_fa83_and0;
  wire s_dadda_cla12_fa83_xor1;
  wire s_dadda_cla12_fa83_and1;
  wire s_dadda_cla12_fa83_or0;
  wire s_dadda_cla12_fa84_xor0;
  wire s_dadda_cla12_fa84_and0;
  wire s_dadda_cla12_fa84_xor1;
  wire s_dadda_cla12_fa84_and1;
  wire s_dadda_cla12_fa84_or0;
  wire s_dadda_cla12_fa85_xor0;
  wire s_dadda_cla12_fa85_and0;
  wire s_dadda_cla12_fa85_xor1;
  wire s_dadda_cla12_fa85_and1;
  wire s_dadda_cla12_fa85_or0;
  wire s_dadda_cla12_fa86_xor0;
  wire s_dadda_cla12_fa86_and0;
  wire s_dadda_cla12_fa86_xor1;
  wire s_dadda_cla12_fa86_and1;
  wire s_dadda_cla12_fa86_or0;
  wire s_dadda_cla12_fa87_xor0;
  wire s_dadda_cla12_fa87_and0;
  wire s_dadda_cla12_fa87_xor1;
  wire s_dadda_cla12_fa87_and1;
  wire s_dadda_cla12_fa87_or0;
  wire s_dadda_cla12_fa88_xor0;
  wire s_dadda_cla12_fa88_and0;
  wire s_dadda_cla12_fa88_xor1;
  wire s_dadda_cla12_fa88_and1;
  wire s_dadda_cla12_fa88_or0;
  wire s_dadda_cla12_fa89_xor0;
  wire s_dadda_cla12_fa89_and0;
  wire s_dadda_cla12_fa89_xor1;
  wire s_dadda_cla12_fa89_and1;
  wire s_dadda_cla12_fa89_or0;
  wire s_dadda_cla12_fa90_xor0;
  wire s_dadda_cla12_fa90_and0;
  wire s_dadda_cla12_fa90_xor1;
  wire s_dadda_cla12_fa90_and1;
  wire s_dadda_cla12_fa90_or0;
  wire s_dadda_cla12_fa91_xor0;
  wire s_dadda_cla12_fa91_and0;
  wire s_dadda_cla12_fa91_xor1;
  wire s_dadda_cla12_fa91_and1;
  wire s_dadda_cla12_fa91_or0;
  wire s_dadda_cla12_fa92_xor0;
  wire s_dadda_cla12_fa92_and0;
  wire s_dadda_cla12_fa92_xor1;
  wire s_dadda_cla12_fa92_and1;
  wire s_dadda_cla12_fa92_or0;
  wire s_dadda_cla12_fa93_xor0;
  wire s_dadda_cla12_fa93_and0;
  wire s_dadda_cla12_fa93_xor1;
  wire s_dadda_cla12_fa93_and1;
  wire s_dadda_cla12_fa93_or0;
  wire s_dadda_cla12_fa94_xor0;
  wire s_dadda_cla12_fa94_and0;
  wire s_dadda_cla12_fa94_xor1;
  wire s_dadda_cla12_fa94_and1;
  wire s_dadda_cla12_fa94_or0;
  wire s_dadda_cla12_fa95_xor0;
  wire s_dadda_cla12_fa95_and0;
  wire s_dadda_cla12_fa95_xor1;
  wire s_dadda_cla12_fa95_and1;
  wire s_dadda_cla12_fa95_or0;
  wire s_dadda_cla12_fa96_xor0;
  wire s_dadda_cla12_fa96_and0;
  wire s_dadda_cla12_fa96_xor1;
  wire s_dadda_cla12_fa96_and1;
  wire s_dadda_cla12_fa96_or0;
  wire s_dadda_cla12_nand_8_11;
  wire s_dadda_cla12_fa97_xor0;
  wire s_dadda_cla12_fa97_and0;
  wire s_dadda_cla12_fa97_xor1;
  wire s_dadda_cla12_fa97_and1;
  wire s_dadda_cla12_fa97_or0;
  wire s_dadda_cla12_and_10_10;
  wire s_dadda_cla12_nand_9_11;
  wire s_dadda_cla12_fa98_xor0;
  wire s_dadda_cla12_fa98_and0;
  wire s_dadda_cla12_fa98_xor1;
  wire s_dadda_cla12_fa98_and1;
  wire s_dadda_cla12_fa98_or0;
  wire s_dadda_cla12_nand_11_10;
  wire s_dadda_cla12_fa99_xor0;
  wire s_dadda_cla12_fa99_and0;
  wire s_dadda_cla12_fa99_xor1;
  wire s_dadda_cla12_fa99_and1;
  wire s_dadda_cla12_fa99_or0;
  wire s_dadda_cla12_and_0_0;
  wire s_dadda_cla12_and_1_0;
  wire s_dadda_cla12_and_0_2;
  wire s_dadda_cla12_nand_10_11;
  wire s_dadda_cla12_and_0_1;
  wire s_dadda_cla12_and_11_11;
  wire s_dadda_cla12_u_cla22_pg_logic0_or0;
  wire s_dadda_cla12_u_cla22_pg_logic0_and0;
  wire s_dadda_cla12_u_cla22_pg_logic0_xor0;
  wire s_dadda_cla12_u_cla22_pg_logic1_or0;
  wire s_dadda_cla12_u_cla22_pg_logic1_and0;
  wire s_dadda_cla12_u_cla22_pg_logic1_xor0;
  wire s_dadda_cla12_u_cla22_xor1;
  wire s_dadda_cla12_u_cla22_and0;
  wire s_dadda_cla12_u_cla22_or0;
  wire s_dadda_cla12_u_cla22_pg_logic2_or0;
  wire s_dadda_cla12_u_cla22_pg_logic2_and0;
  wire s_dadda_cla12_u_cla22_pg_logic2_xor0;
  wire s_dadda_cla12_u_cla22_xor2;
  wire s_dadda_cla12_u_cla22_and1;
  wire s_dadda_cla12_u_cla22_and2;
  wire s_dadda_cla12_u_cla22_and3;
  wire s_dadda_cla12_u_cla22_and4;
  wire s_dadda_cla12_u_cla22_or1;
  wire s_dadda_cla12_u_cla22_or2;
  wire s_dadda_cla12_u_cla22_pg_logic3_or0;
  wire s_dadda_cla12_u_cla22_pg_logic3_and0;
  wire s_dadda_cla12_u_cla22_pg_logic3_xor0;
  wire s_dadda_cla12_u_cla22_xor3;
  wire s_dadda_cla12_u_cla22_and5;
  wire s_dadda_cla12_u_cla22_and6;
  wire s_dadda_cla12_u_cla22_and7;
  wire s_dadda_cla12_u_cla22_and8;
  wire s_dadda_cla12_u_cla22_and9;
  wire s_dadda_cla12_u_cla22_and10;
  wire s_dadda_cla12_u_cla22_and11;
  wire s_dadda_cla12_u_cla22_or3;
  wire s_dadda_cla12_u_cla22_or4;
  wire s_dadda_cla12_u_cla22_or5;
  wire s_dadda_cla12_u_cla22_pg_logic4_or0;
  wire s_dadda_cla12_u_cla22_pg_logic4_and0;
  wire s_dadda_cla12_u_cla22_pg_logic4_xor0;
  wire s_dadda_cla12_u_cla22_xor4;
  wire s_dadda_cla12_u_cla22_and12;
  wire s_dadda_cla12_u_cla22_or6;
  wire s_dadda_cla12_u_cla22_pg_logic5_or0;
  wire s_dadda_cla12_u_cla22_pg_logic5_and0;
  wire s_dadda_cla12_u_cla22_pg_logic5_xor0;
  wire s_dadda_cla12_u_cla22_xor5;
  wire s_dadda_cla12_u_cla22_and13;
  wire s_dadda_cla12_u_cla22_and14;
  wire s_dadda_cla12_u_cla22_and15;
  wire s_dadda_cla12_u_cla22_or7;
  wire s_dadda_cla12_u_cla22_or8;
  wire s_dadda_cla12_u_cla22_pg_logic6_or0;
  wire s_dadda_cla12_u_cla22_pg_logic6_and0;
  wire s_dadda_cla12_u_cla22_pg_logic6_xor0;
  wire s_dadda_cla12_u_cla22_xor6;
  wire s_dadda_cla12_u_cla22_and16;
  wire s_dadda_cla12_u_cla22_and17;
  wire s_dadda_cla12_u_cla22_and18;
  wire s_dadda_cla12_u_cla22_and19;
  wire s_dadda_cla12_u_cla22_and20;
  wire s_dadda_cla12_u_cla22_and21;
  wire s_dadda_cla12_u_cla22_or9;
  wire s_dadda_cla12_u_cla22_or10;
  wire s_dadda_cla12_u_cla22_or11;
  wire s_dadda_cla12_u_cla22_pg_logic7_or0;
  wire s_dadda_cla12_u_cla22_pg_logic7_and0;
  wire s_dadda_cla12_u_cla22_pg_logic7_xor0;
  wire s_dadda_cla12_u_cla22_xor7;
  wire s_dadda_cla12_u_cla22_and22;
  wire s_dadda_cla12_u_cla22_and23;
  wire s_dadda_cla12_u_cla22_and24;
  wire s_dadda_cla12_u_cla22_and25;
  wire s_dadda_cla12_u_cla22_and26;
  wire s_dadda_cla12_u_cla22_and27;
  wire s_dadda_cla12_u_cla22_and28;
  wire s_dadda_cla12_u_cla22_and29;
  wire s_dadda_cla12_u_cla22_and30;
  wire s_dadda_cla12_u_cla22_and31;
  wire s_dadda_cla12_u_cla22_or12;
  wire s_dadda_cla12_u_cla22_or13;
  wire s_dadda_cla12_u_cla22_or14;
  wire s_dadda_cla12_u_cla22_or15;
  wire s_dadda_cla12_u_cla22_pg_logic8_or0;
  wire s_dadda_cla12_u_cla22_pg_logic8_and0;
  wire s_dadda_cla12_u_cla22_pg_logic8_xor0;
  wire s_dadda_cla12_u_cla22_xor8;
  wire s_dadda_cla12_u_cla22_and32;
  wire s_dadda_cla12_u_cla22_or16;
  wire s_dadda_cla12_u_cla22_pg_logic9_or0;
  wire s_dadda_cla12_u_cla22_pg_logic9_and0;
  wire s_dadda_cla12_u_cla22_pg_logic9_xor0;
  wire s_dadda_cla12_u_cla22_xor9;
  wire s_dadda_cla12_u_cla22_and33;
  wire s_dadda_cla12_u_cla22_and34;
  wire s_dadda_cla12_u_cla22_and35;
  wire s_dadda_cla12_u_cla22_or17;
  wire s_dadda_cla12_u_cla22_or18;
  wire s_dadda_cla12_u_cla22_pg_logic10_or0;
  wire s_dadda_cla12_u_cla22_pg_logic10_and0;
  wire s_dadda_cla12_u_cla22_pg_logic10_xor0;
  wire s_dadda_cla12_u_cla22_xor10;
  wire s_dadda_cla12_u_cla22_and36;
  wire s_dadda_cla12_u_cla22_and37;
  wire s_dadda_cla12_u_cla22_and38;
  wire s_dadda_cla12_u_cla22_and39;
  wire s_dadda_cla12_u_cla22_and40;
  wire s_dadda_cla12_u_cla22_and41;
  wire s_dadda_cla12_u_cla22_or19;
  wire s_dadda_cla12_u_cla22_or20;
  wire s_dadda_cla12_u_cla22_or21;
  wire s_dadda_cla12_u_cla22_pg_logic11_or0;
  wire s_dadda_cla12_u_cla22_pg_logic11_and0;
  wire s_dadda_cla12_u_cla22_pg_logic11_xor0;
  wire s_dadda_cla12_u_cla22_xor11;
  wire s_dadda_cla12_u_cla22_and42;
  wire s_dadda_cla12_u_cla22_and43;
  wire s_dadda_cla12_u_cla22_and44;
  wire s_dadda_cla12_u_cla22_and45;
  wire s_dadda_cla12_u_cla22_and46;
  wire s_dadda_cla12_u_cla22_and47;
  wire s_dadda_cla12_u_cla22_and48;
  wire s_dadda_cla12_u_cla22_and49;
  wire s_dadda_cla12_u_cla22_and50;
  wire s_dadda_cla12_u_cla22_and51;
  wire s_dadda_cla12_u_cla22_or22;
  wire s_dadda_cla12_u_cla22_or23;
  wire s_dadda_cla12_u_cla22_or24;
  wire s_dadda_cla12_u_cla22_or25;
  wire s_dadda_cla12_u_cla22_pg_logic12_or0;
  wire s_dadda_cla12_u_cla22_pg_logic12_and0;
  wire s_dadda_cla12_u_cla22_pg_logic12_xor0;
  wire s_dadda_cla12_u_cla22_xor12;
  wire s_dadda_cla12_u_cla22_and52;
  wire s_dadda_cla12_u_cla22_or26;
  wire s_dadda_cla12_u_cla22_pg_logic13_or0;
  wire s_dadda_cla12_u_cla22_pg_logic13_and0;
  wire s_dadda_cla12_u_cla22_pg_logic13_xor0;
  wire s_dadda_cla12_u_cla22_xor13;
  wire s_dadda_cla12_u_cla22_and53;
  wire s_dadda_cla12_u_cla22_and54;
  wire s_dadda_cla12_u_cla22_and55;
  wire s_dadda_cla12_u_cla22_or27;
  wire s_dadda_cla12_u_cla22_or28;
  wire s_dadda_cla12_u_cla22_pg_logic14_or0;
  wire s_dadda_cla12_u_cla22_pg_logic14_and0;
  wire s_dadda_cla12_u_cla22_pg_logic14_xor0;
  wire s_dadda_cla12_u_cla22_xor14;
  wire s_dadda_cla12_u_cla22_and56;
  wire s_dadda_cla12_u_cla22_and57;
  wire s_dadda_cla12_u_cla22_and58;
  wire s_dadda_cla12_u_cla22_and59;
  wire s_dadda_cla12_u_cla22_and60;
  wire s_dadda_cla12_u_cla22_and61;
  wire s_dadda_cla12_u_cla22_or29;
  wire s_dadda_cla12_u_cla22_or30;
  wire s_dadda_cla12_u_cla22_or31;
  wire s_dadda_cla12_u_cla22_pg_logic15_or0;
  wire s_dadda_cla12_u_cla22_pg_logic15_and0;
  wire s_dadda_cla12_u_cla22_pg_logic15_xor0;
  wire s_dadda_cla12_u_cla22_xor15;
  wire s_dadda_cla12_u_cla22_and62;
  wire s_dadda_cla12_u_cla22_and63;
  wire s_dadda_cla12_u_cla22_and64;
  wire s_dadda_cla12_u_cla22_and65;
  wire s_dadda_cla12_u_cla22_and66;
  wire s_dadda_cla12_u_cla22_and67;
  wire s_dadda_cla12_u_cla22_and68;
  wire s_dadda_cla12_u_cla22_and69;
  wire s_dadda_cla12_u_cla22_and70;
  wire s_dadda_cla12_u_cla22_and71;
  wire s_dadda_cla12_u_cla22_or32;
  wire s_dadda_cla12_u_cla22_or33;
  wire s_dadda_cla12_u_cla22_or34;
  wire s_dadda_cla12_u_cla22_or35;
  wire s_dadda_cla12_u_cla22_pg_logic16_or0;
  wire s_dadda_cla12_u_cla22_pg_logic16_and0;
  wire s_dadda_cla12_u_cla22_pg_logic16_xor0;
  wire s_dadda_cla12_u_cla22_xor16;
  wire s_dadda_cla12_u_cla22_and72;
  wire s_dadda_cla12_u_cla22_or36;
  wire s_dadda_cla12_u_cla22_pg_logic17_or0;
  wire s_dadda_cla12_u_cla22_pg_logic17_and0;
  wire s_dadda_cla12_u_cla22_pg_logic17_xor0;
  wire s_dadda_cla12_u_cla22_xor17;
  wire s_dadda_cla12_u_cla22_and73;
  wire s_dadda_cla12_u_cla22_and74;
  wire s_dadda_cla12_u_cla22_and75;
  wire s_dadda_cla12_u_cla22_or37;
  wire s_dadda_cla12_u_cla22_or38;
  wire s_dadda_cla12_u_cla22_pg_logic18_or0;
  wire s_dadda_cla12_u_cla22_pg_logic18_and0;
  wire s_dadda_cla12_u_cla22_pg_logic18_xor0;
  wire s_dadda_cla12_u_cla22_xor18;
  wire s_dadda_cla12_u_cla22_and76;
  wire s_dadda_cla12_u_cla22_and77;
  wire s_dadda_cla12_u_cla22_and78;
  wire s_dadda_cla12_u_cla22_and79;
  wire s_dadda_cla12_u_cla22_and80;
  wire s_dadda_cla12_u_cla22_and81;
  wire s_dadda_cla12_u_cla22_or39;
  wire s_dadda_cla12_u_cla22_or40;
  wire s_dadda_cla12_u_cla22_or41;
  wire s_dadda_cla12_u_cla22_pg_logic19_or0;
  wire s_dadda_cla12_u_cla22_pg_logic19_and0;
  wire s_dadda_cla12_u_cla22_pg_logic19_xor0;
  wire s_dadda_cla12_u_cla22_xor19;
  wire s_dadda_cla12_u_cla22_and82;
  wire s_dadda_cla12_u_cla22_and83;
  wire s_dadda_cla12_u_cla22_and84;
  wire s_dadda_cla12_u_cla22_and85;
  wire s_dadda_cla12_u_cla22_and86;
  wire s_dadda_cla12_u_cla22_and87;
  wire s_dadda_cla12_u_cla22_and88;
  wire s_dadda_cla12_u_cla22_and89;
  wire s_dadda_cla12_u_cla22_and90;
  wire s_dadda_cla12_u_cla22_and91;
  wire s_dadda_cla12_u_cla22_or42;
  wire s_dadda_cla12_u_cla22_or43;
  wire s_dadda_cla12_u_cla22_or44;
  wire s_dadda_cla12_u_cla22_or45;
  wire s_dadda_cla12_u_cla22_pg_logic20_or0;
  wire s_dadda_cla12_u_cla22_pg_logic20_and0;
  wire s_dadda_cla12_u_cla22_pg_logic20_xor0;
  wire s_dadda_cla12_u_cla22_xor20;
  wire s_dadda_cla12_u_cla22_and92;
  wire s_dadda_cla12_u_cla22_or46;
  wire s_dadda_cla12_u_cla22_pg_logic21_or0;
  wire s_dadda_cla12_u_cla22_pg_logic21_and0;
  wire s_dadda_cla12_u_cla22_pg_logic21_xor0;
  wire s_dadda_cla12_u_cla22_xor21;
  wire s_dadda_cla12_u_cla22_and93;
  wire s_dadda_cla12_u_cla22_and94;
  wire s_dadda_cla12_u_cla22_and95;
  wire s_dadda_cla12_u_cla22_or47;
  wire s_dadda_cla12_u_cla22_or48;
  wire s_dadda_cla12_xor0;

  assign s_dadda_cla12_and_9_0 = a[9] & b[0];
  assign s_dadda_cla12_and_8_1 = a[8] & b[1];
  assign s_dadda_cla12_ha0_xor0 = s_dadda_cla12_and_9_0 ^ s_dadda_cla12_and_8_1;
  assign s_dadda_cla12_ha0_and0 = s_dadda_cla12_and_9_0 & s_dadda_cla12_and_8_1;
  assign s_dadda_cla12_and_10_0 = a[10] & b[0];
  assign s_dadda_cla12_and_9_1 = a[9] & b[1];
  assign s_dadda_cla12_fa0_xor0 = s_dadda_cla12_ha0_and0 ^ s_dadda_cla12_and_10_0;
  assign s_dadda_cla12_fa0_and0 = s_dadda_cla12_ha0_and0 & s_dadda_cla12_and_10_0;
  assign s_dadda_cla12_fa0_xor1 = s_dadda_cla12_fa0_xor0 ^ s_dadda_cla12_and_9_1;
  assign s_dadda_cla12_fa0_and1 = s_dadda_cla12_fa0_xor0 & s_dadda_cla12_and_9_1;
  assign s_dadda_cla12_fa0_or0 = s_dadda_cla12_fa0_and0 | s_dadda_cla12_fa0_and1;
  assign s_dadda_cla12_and_8_2 = a[8] & b[2];
  assign s_dadda_cla12_and_7_3 = a[7] & b[3];
  assign s_dadda_cla12_ha1_xor0 = s_dadda_cla12_and_8_2 ^ s_dadda_cla12_and_7_3;
  assign s_dadda_cla12_ha1_and0 = s_dadda_cla12_and_8_2 & s_dadda_cla12_and_7_3;
  assign s_dadda_cla12_nand_11_0 = ~(a[11] & b[0]);
  assign s_dadda_cla12_fa1_xor0 = s_dadda_cla12_ha1_and0 ^ s_dadda_cla12_fa0_or0;
  assign s_dadda_cla12_fa1_and0 = s_dadda_cla12_ha1_and0 & s_dadda_cla12_fa0_or0;
  assign s_dadda_cla12_fa1_xor1 = s_dadda_cla12_fa1_xor0 ^ s_dadda_cla12_nand_11_0;
  assign s_dadda_cla12_fa1_and1 = s_dadda_cla12_fa1_xor0 & s_dadda_cla12_nand_11_0;
  assign s_dadda_cla12_fa1_or0 = s_dadda_cla12_fa1_and0 | s_dadda_cla12_fa1_and1;
  assign s_dadda_cla12_and_10_1 = a[10] & b[1];
  assign s_dadda_cla12_and_9_2 = a[9] & b[2];
  assign s_dadda_cla12_and_8_3 = a[8] & b[3];
  assign s_dadda_cla12_fa2_xor0 = s_dadda_cla12_and_10_1 ^ s_dadda_cla12_and_9_2;
  assign s_dadda_cla12_fa2_and0 = s_dadda_cla12_and_10_1 & s_dadda_cla12_and_9_2;
  assign s_dadda_cla12_fa2_xor1 = s_dadda_cla12_fa2_xor0 ^ s_dadda_cla12_and_8_3;
  assign s_dadda_cla12_fa2_and1 = s_dadda_cla12_fa2_xor0 & s_dadda_cla12_and_8_3;
  assign s_dadda_cla12_fa2_or0 = s_dadda_cla12_fa2_and0 | s_dadda_cla12_fa2_and1;
  assign s_dadda_cla12_and_7_4 = a[7] & b[4];
  assign s_dadda_cla12_and_6_5 = a[6] & b[5];
  assign s_dadda_cla12_ha2_xor0 = s_dadda_cla12_and_7_4 ^ s_dadda_cla12_and_6_5;
  assign s_dadda_cla12_ha2_and0 = s_dadda_cla12_and_7_4 & s_dadda_cla12_and_6_5;
  assign s_dadda_cla12_fa3_xor0 = s_dadda_cla12_ha2_and0 ^ s_dadda_cla12_fa2_or0;
  assign s_dadda_cla12_fa3_and0 = s_dadda_cla12_ha2_and0 & s_dadda_cla12_fa2_or0;
  assign s_dadda_cla12_fa3_xor1 = s_dadda_cla12_fa3_xor0 ^ s_dadda_cla12_fa1_or0;
  assign s_dadda_cla12_fa3_and1 = s_dadda_cla12_fa3_xor0 & s_dadda_cla12_fa1_or0;
  assign s_dadda_cla12_fa3_or0 = s_dadda_cla12_fa3_and0 | s_dadda_cla12_fa3_and1;
  assign s_dadda_cla12_nand_11_1 = ~(a[11] & b[1]);
  assign s_dadda_cla12_and_10_2 = a[10] & b[2];
  assign s_dadda_cla12_fa4_xor0 = ~s_dadda_cla12_nand_11_1;
  assign s_dadda_cla12_fa4_xor1 = s_dadda_cla12_fa4_xor0 ^ s_dadda_cla12_and_10_2;
  assign s_dadda_cla12_fa4_and1 = s_dadda_cla12_fa4_xor0 & s_dadda_cla12_and_10_2;
  assign s_dadda_cla12_fa4_or0 = s_dadda_cla12_nand_11_1 | s_dadda_cla12_fa4_and1;
  assign s_dadda_cla12_and_9_3 = a[9] & b[3];
  assign s_dadda_cla12_and_8_4 = a[8] & b[4];
  assign s_dadda_cla12_and_7_5 = a[7] & b[5];
  assign s_dadda_cla12_fa5_xor0 = s_dadda_cla12_and_9_3 ^ s_dadda_cla12_and_8_4;
  assign s_dadda_cla12_fa5_and0 = s_dadda_cla12_and_9_3 & s_dadda_cla12_and_8_4;
  assign s_dadda_cla12_fa5_xor1 = s_dadda_cla12_fa5_xor0 ^ s_dadda_cla12_and_7_5;
  assign s_dadda_cla12_fa5_and1 = s_dadda_cla12_fa5_xor0 & s_dadda_cla12_and_7_5;
  assign s_dadda_cla12_fa5_or0 = s_dadda_cla12_fa5_and0 | s_dadda_cla12_fa5_and1;
  assign s_dadda_cla12_fa6_xor0 = s_dadda_cla12_fa5_or0 ^ s_dadda_cla12_fa4_or0;
  assign s_dadda_cla12_fa6_and0 = s_dadda_cla12_fa5_or0 & s_dadda_cla12_fa4_or0;
  assign s_dadda_cla12_fa6_xor1 = s_dadda_cla12_fa6_xor0 ^ s_dadda_cla12_fa3_or0;
  assign s_dadda_cla12_fa6_and1 = s_dadda_cla12_fa6_xor0 & s_dadda_cla12_fa3_or0;
  assign s_dadda_cla12_fa6_or0 = s_dadda_cla12_fa6_and0 | s_dadda_cla12_fa6_and1;
  assign s_dadda_cla12_nand_11_2 = ~(a[11] & b[2]);
  assign s_dadda_cla12_and_10_3 = a[10] & b[3];
  assign s_dadda_cla12_and_9_4 = a[9] & b[4];
  assign s_dadda_cla12_fa7_xor0 = s_dadda_cla12_nand_11_2 ^ s_dadda_cla12_and_10_3;
  assign s_dadda_cla12_fa7_and0 = s_dadda_cla12_nand_11_2 & s_dadda_cla12_and_10_3;
  assign s_dadda_cla12_fa7_xor1 = s_dadda_cla12_fa7_xor0 ^ s_dadda_cla12_and_9_4;
  assign s_dadda_cla12_fa7_and1 = s_dadda_cla12_fa7_xor0 & s_dadda_cla12_and_9_4;
  assign s_dadda_cla12_fa7_or0 = s_dadda_cla12_fa7_and0 | s_dadda_cla12_fa7_and1;
  assign s_dadda_cla12_nand_11_3 = ~(a[11] & b[3]);
  assign s_dadda_cla12_fa8_xor0 = s_dadda_cla12_fa7_or0 ^ s_dadda_cla12_fa6_or0;
  assign s_dadda_cla12_fa8_and0 = s_dadda_cla12_fa7_or0 & s_dadda_cla12_fa6_or0;
  assign s_dadda_cla12_fa8_xor1 = s_dadda_cla12_fa8_xor0 ^ s_dadda_cla12_nand_11_3;
  assign s_dadda_cla12_fa8_and1 = s_dadda_cla12_fa8_xor0 & s_dadda_cla12_nand_11_3;
  assign s_dadda_cla12_fa8_or0 = s_dadda_cla12_fa8_and0 | s_dadda_cla12_fa8_and1;
  assign s_dadda_cla12_and_4_0 = a[4] & b[0];
  assign s_dadda_cla12_and_3_1 = a[3] & b[1];
  assign s_dadda_cla12_ha3_xor0 = s_dadda_cla12_and_4_0 ^ s_dadda_cla12_and_3_1;
  assign s_dadda_cla12_ha3_and0 = s_dadda_cla12_and_4_0 & s_dadda_cla12_and_3_1;
  assign s_dadda_cla12_and_5_0 = a[5] & b[0];
  assign s_dadda_cla12_and_4_1 = a[4] & b[1];
  assign s_dadda_cla12_fa9_xor0 = s_dadda_cla12_ha3_and0 ^ s_dadda_cla12_and_5_0;
  assign s_dadda_cla12_fa9_and0 = s_dadda_cla12_ha3_and0 & s_dadda_cla12_and_5_0;
  assign s_dadda_cla12_fa9_xor1 = s_dadda_cla12_fa9_xor0 ^ s_dadda_cla12_and_4_1;
  assign s_dadda_cla12_fa9_and1 = s_dadda_cla12_fa9_xor0 & s_dadda_cla12_and_4_1;
  assign s_dadda_cla12_fa9_or0 = s_dadda_cla12_fa9_and0 | s_dadda_cla12_fa9_and1;
  assign s_dadda_cla12_and_3_2 = a[3] & b[2];
  assign s_dadda_cla12_and_2_3 = a[2] & b[3];
  assign s_dadda_cla12_ha4_xor0 = s_dadda_cla12_and_3_2 ^ s_dadda_cla12_and_2_3;
  assign s_dadda_cla12_ha4_and0 = s_dadda_cla12_and_3_2 & s_dadda_cla12_and_2_3;
  assign s_dadda_cla12_and_6_0 = a[6] & b[0];
  assign s_dadda_cla12_fa10_xor0 = s_dadda_cla12_ha4_and0 ^ s_dadda_cla12_fa9_or0;
  assign s_dadda_cla12_fa10_and0 = s_dadda_cla12_ha4_and0 & s_dadda_cla12_fa9_or0;
  assign s_dadda_cla12_fa10_xor1 = s_dadda_cla12_fa10_xor0 ^ s_dadda_cla12_and_6_0;
  assign s_dadda_cla12_fa10_and1 = s_dadda_cla12_fa10_xor0 & s_dadda_cla12_and_6_0;
  assign s_dadda_cla12_fa10_or0 = s_dadda_cla12_fa10_and0 | s_dadda_cla12_fa10_and1;
  assign s_dadda_cla12_and_5_1 = a[5] & b[1];
  assign s_dadda_cla12_and_4_2 = a[4] & b[2];
  assign s_dadda_cla12_and_3_3 = a[3] & b[3];
  assign s_dadda_cla12_fa11_xor0 = s_dadda_cla12_and_5_1 ^ s_dadda_cla12_and_4_2;
  assign s_dadda_cla12_fa11_and0 = s_dadda_cla12_and_5_1 & s_dadda_cla12_and_4_2;
  assign s_dadda_cla12_fa11_xor1 = s_dadda_cla12_fa11_xor0 ^ s_dadda_cla12_and_3_3;
  assign s_dadda_cla12_fa11_and1 = s_dadda_cla12_fa11_xor0 & s_dadda_cla12_and_3_3;
  assign s_dadda_cla12_fa11_or0 = s_dadda_cla12_fa11_and0 | s_dadda_cla12_fa11_and1;
  assign s_dadda_cla12_and_2_4 = a[2] & b[4];
  assign s_dadda_cla12_and_1_5 = a[1] & b[5];
  assign s_dadda_cla12_ha5_xor0 = s_dadda_cla12_and_2_4 ^ s_dadda_cla12_and_1_5;
  assign s_dadda_cla12_ha5_and0 = s_dadda_cla12_and_2_4 & s_dadda_cla12_and_1_5;
  assign s_dadda_cla12_fa12_xor0 = s_dadda_cla12_ha5_and0 ^ s_dadda_cla12_fa11_or0;
  assign s_dadda_cla12_fa12_and0 = s_dadda_cla12_ha5_and0 & s_dadda_cla12_fa11_or0;
  assign s_dadda_cla12_fa12_xor1 = s_dadda_cla12_fa12_xor0 ^ s_dadda_cla12_fa10_or0;
  assign s_dadda_cla12_fa12_and1 = s_dadda_cla12_fa12_xor0 & s_dadda_cla12_fa10_or0;
  assign s_dadda_cla12_fa12_or0 = s_dadda_cla12_fa12_and0 | s_dadda_cla12_fa12_and1;
  assign s_dadda_cla12_and_7_0 = a[7] & b[0];
  assign s_dadda_cla12_and_6_1 = a[6] & b[1];
  assign s_dadda_cla12_and_5_2 = a[5] & b[2];
  assign s_dadda_cla12_fa13_xor0 = s_dadda_cla12_and_7_0 ^ s_dadda_cla12_and_6_1;
  assign s_dadda_cla12_fa13_and0 = s_dadda_cla12_and_7_0 & s_dadda_cla12_and_6_1;
  assign s_dadda_cla12_fa13_xor1 = s_dadda_cla12_fa13_xor0 ^ s_dadda_cla12_and_5_2;
  assign s_dadda_cla12_fa13_and1 = s_dadda_cla12_fa13_xor0 & s_dadda_cla12_and_5_2;
  assign s_dadda_cla12_fa13_or0 = s_dadda_cla12_fa13_and0 | s_dadda_cla12_fa13_and1;
  assign s_dadda_cla12_and_4_3 = a[4] & b[3];
  assign s_dadda_cla12_and_3_4 = a[3] & b[4];
  assign s_dadda_cla12_and_2_5 = a[2] & b[5];
  assign s_dadda_cla12_fa14_xor0 = s_dadda_cla12_and_4_3 ^ s_dadda_cla12_and_3_4;
  assign s_dadda_cla12_fa14_and0 = s_dadda_cla12_and_4_3 & s_dadda_cla12_and_3_4;
  assign s_dadda_cla12_fa14_xor1 = s_dadda_cla12_fa14_xor0 ^ s_dadda_cla12_and_2_5;
  assign s_dadda_cla12_fa14_and1 = s_dadda_cla12_fa14_xor0 & s_dadda_cla12_and_2_5;
  assign s_dadda_cla12_fa14_or0 = s_dadda_cla12_fa14_and0 | s_dadda_cla12_fa14_and1;
  assign s_dadda_cla12_and_1_6 = a[1] & b[6];
  assign s_dadda_cla12_and_0_7 = a[0] & b[7];
  assign s_dadda_cla12_ha6_xor0 = s_dadda_cla12_and_1_6 ^ s_dadda_cla12_and_0_7;
  assign s_dadda_cla12_ha6_and0 = s_dadda_cla12_and_1_6 & s_dadda_cla12_and_0_7;
  assign s_dadda_cla12_fa15_xor0 = s_dadda_cla12_ha6_and0 ^ s_dadda_cla12_fa14_or0;
  assign s_dadda_cla12_fa15_and0 = s_dadda_cla12_ha6_and0 & s_dadda_cla12_fa14_or0;
  assign s_dadda_cla12_fa15_xor1 = s_dadda_cla12_fa15_xor0 ^ s_dadda_cla12_fa13_or0;
  assign s_dadda_cla12_fa15_and1 = s_dadda_cla12_fa15_xor0 & s_dadda_cla12_fa13_or0;
  assign s_dadda_cla12_fa15_or0 = s_dadda_cla12_fa15_and0 | s_dadda_cla12_fa15_and1;
  assign s_dadda_cla12_and_8_0 = a[8] & b[0];
  assign s_dadda_cla12_and_7_1 = a[7] & b[1];
  assign s_dadda_cla12_fa16_xor0 = s_dadda_cla12_fa12_or0 ^ s_dadda_cla12_and_8_0;
  assign s_dadda_cla12_fa16_and0 = s_dadda_cla12_fa12_or0 & s_dadda_cla12_and_8_0;
  assign s_dadda_cla12_fa16_xor1 = s_dadda_cla12_fa16_xor0 ^ s_dadda_cla12_and_7_1;
  assign s_dadda_cla12_fa16_and1 = s_dadda_cla12_fa16_xor0 & s_dadda_cla12_and_7_1;
  assign s_dadda_cla12_fa16_or0 = s_dadda_cla12_fa16_and0 | s_dadda_cla12_fa16_and1;
  assign s_dadda_cla12_and_6_2 = a[6] & b[2];
  assign s_dadda_cla12_and_5_3 = a[5] & b[3];
  assign s_dadda_cla12_and_4_4 = a[4] & b[4];
  assign s_dadda_cla12_fa17_xor0 = s_dadda_cla12_and_6_2 ^ s_dadda_cla12_and_5_3;
  assign s_dadda_cla12_fa17_and0 = s_dadda_cla12_and_6_2 & s_dadda_cla12_and_5_3;
  assign s_dadda_cla12_fa17_xor1 = s_dadda_cla12_fa17_xor0 ^ s_dadda_cla12_and_4_4;
  assign s_dadda_cla12_fa17_and1 = s_dadda_cla12_fa17_xor0 & s_dadda_cla12_and_4_4;
  assign s_dadda_cla12_fa17_or0 = s_dadda_cla12_fa17_and0 | s_dadda_cla12_fa17_and1;
  assign s_dadda_cla12_and_3_5 = a[3] & b[5];
  assign s_dadda_cla12_and_2_6 = a[2] & b[6];
  assign s_dadda_cla12_and_1_7 = a[1] & b[7];
  assign s_dadda_cla12_fa18_xor0 = s_dadda_cla12_and_3_5 ^ s_dadda_cla12_and_2_6;
  assign s_dadda_cla12_fa18_and0 = s_dadda_cla12_and_3_5 & s_dadda_cla12_and_2_6;
  assign s_dadda_cla12_fa18_xor1 = s_dadda_cla12_fa18_xor0 ^ s_dadda_cla12_and_1_7;
  assign s_dadda_cla12_fa18_and1 = s_dadda_cla12_fa18_xor0 & s_dadda_cla12_and_1_7;
  assign s_dadda_cla12_fa18_or0 = s_dadda_cla12_fa18_and0 | s_dadda_cla12_fa18_and1;
  assign s_dadda_cla12_and_0_8 = a[0] & b[8];
  assign s_dadda_cla12_ha7_xor0 = s_dadda_cla12_and_0_8 ^ s_dadda_cla12_fa15_xor1;
  assign s_dadda_cla12_ha7_and0 = s_dadda_cla12_and_0_8 & s_dadda_cla12_fa15_xor1;
  assign s_dadda_cla12_fa19_xor0 = s_dadda_cla12_ha7_and0 ^ s_dadda_cla12_fa18_or0;
  assign s_dadda_cla12_fa19_and0 = s_dadda_cla12_ha7_and0 & s_dadda_cla12_fa18_or0;
  assign s_dadda_cla12_fa19_xor1 = s_dadda_cla12_fa19_xor0 ^ s_dadda_cla12_fa17_or0;
  assign s_dadda_cla12_fa19_and1 = s_dadda_cla12_fa19_xor0 & s_dadda_cla12_fa17_or0;
  assign s_dadda_cla12_fa19_or0 = s_dadda_cla12_fa19_and0 | s_dadda_cla12_fa19_and1;
  assign s_dadda_cla12_and_7_2 = a[7] & b[2];
  assign s_dadda_cla12_fa20_xor0 = s_dadda_cla12_fa16_or0 ^ s_dadda_cla12_fa15_or0;
  assign s_dadda_cla12_fa20_and0 = s_dadda_cla12_fa16_or0 & s_dadda_cla12_fa15_or0;
  assign s_dadda_cla12_fa20_xor1 = s_dadda_cla12_fa20_xor0 ^ s_dadda_cla12_and_7_2;
  assign s_dadda_cla12_fa20_and1 = s_dadda_cla12_fa20_xor0 & s_dadda_cla12_and_7_2;
  assign s_dadda_cla12_fa20_or0 = s_dadda_cla12_fa20_and0 | s_dadda_cla12_fa20_and1;
  assign s_dadda_cla12_and_6_3 = a[6] & b[3];
  assign s_dadda_cla12_and_5_4 = a[5] & b[4];
  assign s_dadda_cla12_and_4_5 = a[4] & b[5];
  assign s_dadda_cla12_fa21_xor0 = s_dadda_cla12_and_6_3 ^ s_dadda_cla12_and_5_4;
  assign s_dadda_cla12_fa21_and0 = s_dadda_cla12_and_6_3 & s_dadda_cla12_and_5_4;
  assign s_dadda_cla12_fa21_xor1 = s_dadda_cla12_fa21_xor0 ^ s_dadda_cla12_and_4_5;
  assign s_dadda_cla12_fa21_and1 = s_dadda_cla12_fa21_xor0 & s_dadda_cla12_and_4_5;
  assign s_dadda_cla12_fa21_or0 = s_dadda_cla12_fa21_and0 | s_dadda_cla12_fa21_and1;
  assign s_dadda_cla12_and_3_6 = a[3] & b[6];
  assign s_dadda_cla12_and_2_7 = a[2] & b[7];
  assign s_dadda_cla12_and_1_8 = a[1] & b[8];
  assign s_dadda_cla12_fa22_xor0 = s_dadda_cla12_and_3_6 ^ s_dadda_cla12_and_2_7;
  assign s_dadda_cla12_fa22_and0 = s_dadda_cla12_and_3_6 & s_dadda_cla12_and_2_7;
  assign s_dadda_cla12_fa22_xor1 = s_dadda_cla12_fa22_xor0 ^ s_dadda_cla12_and_1_8;
  assign s_dadda_cla12_fa22_and1 = s_dadda_cla12_fa22_xor0 & s_dadda_cla12_and_1_8;
  assign s_dadda_cla12_fa22_or0 = s_dadda_cla12_fa22_and0 | s_dadda_cla12_fa22_and1;
  assign s_dadda_cla12_and_0_9 = a[0] & b[9];
  assign s_dadda_cla12_fa23_xor0 = s_dadda_cla12_and_0_9 ^ s_dadda_cla12_ha0_xor0;
  assign s_dadda_cla12_fa23_and0 = s_dadda_cla12_and_0_9 & s_dadda_cla12_ha0_xor0;
  assign s_dadda_cla12_fa23_xor1 = s_dadda_cla12_fa23_xor0 ^ s_dadda_cla12_fa19_xor1;
  assign s_dadda_cla12_fa23_and1 = s_dadda_cla12_fa23_xor0 & s_dadda_cla12_fa19_xor1;
  assign s_dadda_cla12_fa23_or0 = s_dadda_cla12_fa23_and0 | s_dadda_cla12_fa23_and1;
  assign s_dadda_cla12_fa24_xor0 = s_dadda_cla12_fa23_or0 ^ s_dadda_cla12_fa22_or0;
  assign s_dadda_cla12_fa24_and0 = s_dadda_cla12_fa23_or0 & s_dadda_cla12_fa22_or0;
  assign s_dadda_cla12_fa24_xor1 = s_dadda_cla12_fa24_xor0 ^ s_dadda_cla12_fa21_or0;
  assign s_dadda_cla12_fa24_and1 = s_dadda_cla12_fa24_xor0 & s_dadda_cla12_fa21_or0;
  assign s_dadda_cla12_fa24_or0 = s_dadda_cla12_fa24_and0 | s_dadda_cla12_fa24_and1;
  assign s_dadda_cla12_and_6_4 = a[6] & b[4];
  assign s_dadda_cla12_fa25_xor0 = s_dadda_cla12_fa20_or0 ^ s_dadda_cla12_fa19_or0;
  assign s_dadda_cla12_fa25_and0 = s_dadda_cla12_fa20_or0 & s_dadda_cla12_fa19_or0;
  assign s_dadda_cla12_fa25_xor1 = s_dadda_cla12_fa25_xor0 ^ s_dadda_cla12_and_6_4;
  assign s_dadda_cla12_fa25_and1 = s_dadda_cla12_fa25_xor0 & s_dadda_cla12_and_6_4;
  assign s_dadda_cla12_fa25_or0 = s_dadda_cla12_fa25_and0 | s_dadda_cla12_fa25_and1;
  assign s_dadda_cla12_and_5_5 = a[5] & b[5];
  assign s_dadda_cla12_and_4_6 = a[4] & b[6];
  assign s_dadda_cla12_and_3_7 = a[3] & b[7];
  assign s_dadda_cla12_fa26_xor0 = s_dadda_cla12_and_5_5 ^ s_dadda_cla12_and_4_6;
  assign s_dadda_cla12_fa26_and0 = s_dadda_cla12_and_5_5 & s_dadda_cla12_and_4_6;
  assign s_dadda_cla12_fa26_xor1 = s_dadda_cla12_fa26_xor0 ^ s_dadda_cla12_and_3_7;
  assign s_dadda_cla12_fa26_and1 = s_dadda_cla12_fa26_xor0 & s_dadda_cla12_and_3_7;
  assign s_dadda_cla12_fa26_or0 = s_dadda_cla12_fa26_and0 | s_dadda_cla12_fa26_and1;
  assign s_dadda_cla12_and_2_8 = a[2] & b[8];
  assign s_dadda_cla12_and_1_9 = a[1] & b[9];
  assign s_dadda_cla12_and_0_10 = a[0] & b[10];
  assign s_dadda_cla12_fa27_xor0 = s_dadda_cla12_and_2_8 ^ s_dadda_cla12_and_1_9;
  assign s_dadda_cla12_fa27_and0 = s_dadda_cla12_and_2_8 & s_dadda_cla12_and_1_9;
  assign s_dadda_cla12_fa27_xor1 = s_dadda_cla12_fa27_xor0 ^ s_dadda_cla12_and_0_10;
  assign s_dadda_cla12_fa27_and1 = s_dadda_cla12_fa27_xor0 & s_dadda_cla12_and_0_10;
  assign s_dadda_cla12_fa27_or0 = s_dadda_cla12_fa27_and0 | s_dadda_cla12_fa27_and1;
  assign s_dadda_cla12_fa28_xor0 = s_dadda_cla12_fa0_xor1 ^ s_dadda_cla12_ha1_xor0;
  assign s_dadda_cla12_fa28_and0 = s_dadda_cla12_fa0_xor1 & s_dadda_cla12_ha1_xor0;
  assign s_dadda_cla12_fa28_xor1 = s_dadda_cla12_fa28_xor0 ^ s_dadda_cla12_fa24_xor1;
  assign s_dadda_cla12_fa28_and1 = s_dadda_cla12_fa28_xor0 & s_dadda_cla12_fa24_xor1;
  assign s_dadda_cla12_fa28_or0 = s_dadda_cla12_fa28_and0 | s_dadda_cla12_fa28_and1;
  assign s_dadda_cla12_fa29_xor0 = s_dadda_cla12_fa28_or0 ^ s_dadda_cla12_fa27_or0;
  assign s_dadda_cla12_fa29_and0 = s_dadda_cla12_fa28_or0 & s_dadda_cla12_fa27_or0;
  assign s_dadda_cla12_fa29_xor1 = s_dadda_cla12_fa29_xor0 ^ s_dadda_cla12_fa26_or0;
  assign s_dadda_cla12_fa29_and1 = s_dadda_cla12_fa29_xor0 & s_dadda_cla12_fa26_or0;
  assign s_dadda_cla12_fa29_or0 = s_dadda_cla12_fa29_and0 | s_dadda_cla12_fa29_and1;
  assign s_dadda_cla12_and_5_6 = a[5] & b[6];
  assign s_dadda_cla12_fa30_xor0 = s_dadda_cla12_fa25_or0 ^ s_dadda_cla12_fa24_or0;
  assign s_dadda_cla12_fa30_and0 = s_dadda_cla12_fa25_or0 & s_dadda_cla12_fa24_or0;
  assign s_dadda_cla12_fa30_xor1 = s_dadda_cla12_fa30_xor0 ^ s_dadda_cla12_and_5_6;
  assign s_dadda_cla12_fa30_and1 = s_dadda_cla12_fa30_xor0 & s_dadda_cla12_and_5_6;
  assign s_dadda_cla12_fa30_or0 = s_dadda_cla12_fa30_and0 | s_dadda_cla12_fa30_and1;
  assign s_dadda_cla12_and_4_7 = a[4] & b[7];
  assign s_dadda_cla12_and_3_8 = a[3] & b[8];
  assign s_dadda_cla12_and_2_9 = a[2] & b[9];
  assign s_dadda_cla12_fa31_xor0 = s_dadda_cla12_and_4_7 ^ s_dadda_cla12_and_3_8;
  assign s_dadda_cla12_fa31_and0 = s_dadda_cla12_and_4_7 & s_dadda_cla12_and_3_8;
  assign s_dadda_cla12_fa31_xor1 = s_dadda_cla12_fa31_xor0 ^ s_dadda_cla12_and_2_9;
  assign s_dadda_cla12_fa31_and1 = s_dadda_cla12_fa31_xor0 & s_dadda_cla12_and_2_9;
  assign s_dadda_cla12_fa31_or0 = s_dadda_cla12_fa31_and0 | s_dadda_cla12_fa31_and1;
  assign s_dadda_cla12_and_1_10 = a[1] & b[10];
  assign s_dadda_cla12_nand_0_11 = ~(a[0] & b[11]);
  assign s_dadda_cla12_fa32_xor0 = s_dadda_cla12_and_1_10 ^ s_dadda_cla12_nand_0_11;
  assign s_dadda_cla12_fa32_and0 = s_dadda_cla12_and_1_10 & s_dadda_cla12_nand_0_11;
  assign s_dadda_cla12_fa32_xor1 = s_dadda_cla12_fa32_xor0 ^ s_dadda_cla12_fa1_xor1;
  assign s_dadda_cla12_fa32_and1 = s_dadda_cla12_fa32_xor0 & s_dadda_cla12_fa1_xor1;
  assign s_dadda_cla12_fa32_or0 = s_dadda_cla12_fa32_and0 | s_dadda_cla12_fa32_and1;
  assign s_dadda_cla12_fa33_xor0 = s_dadda_cla12_fa2_xor1 ^ s_dadda_cla12_ha2_xor0;
  assign s_dadda_cla12_fa33_and0 = s_dadda_cla12_fa2_xor1 & s_dadda_cla12_ha2_xor0;
  assign s_dadda_cla12_fa33_xor1 = s_dadda_cla12_fa33_xor0 ^ s_dadda_cla12_fa29_xor1;
  assign s_dadda_cla12_fa33_and1 = s_dadda_cla12_fa33_xor0 & s_dadda_cla12_fa29_xor1;
  assign s_dadda_cla12_fa33_or0 = s_dadda_cla12_fa33_and0 | s_dadda_cla12_fa33_and1;
  assign s_dadda_cla12_fa34_xor0 = s_dadda_cla12_fa33_or0 ^ s_dadda_cla12_fa32_or0;
  assign s_dadda_cla12_fa34_and0 = s_dadda_cla12_fa33_or0 & s_dadda_cla12_fa32_or0;
  assign s_dadda_cla12_fa34_xor1 = s_dadda_cla12_fa34_xor0 ^ s_dadda_cla12_fa31_or0;
  assign s_dadda_cla12_fa34_and1 = s_dadda_cla12_fa34_xor0 & s_dadda_cla12_fa31_or0;
  assign s_dadda_cla12_fa34_or0 = s_dadda_cla12_fa34_and0 | s_dadda_cla12_fa34_and1;
  assign s_dadda_cla12_and_6_6 = a[6] & b[6];
  assign s_dadda_cla12_fa35_xor0 = s_dadda_cla12_fa30_or0 ^ s_dadda_cla12_fa29_or0;
  assign s_dadda_cla12_fa35_and0 = s_dadda_cla12_fa30_or0 & s_dadda_cla12_fa29_or0;
  assign s_dadda_cla12_fa35_xor1 = s_dadda_cla12_fa35_xor0 ^ s_dadda_cla12_and_6_6;
  assign s_dadda_cla12_fa35_and1 = s_dadda_cla12_fa35_xor0 & s_dadda_cla12_and_6_6;
  assign s_dadda_cla12_fa35_or0 = s_dadda_cla12_fa35_and0 | s_dadda_cla12_fa35_and1;
  assign s_dadda_cla12_and_5_7 = a[5] & b[7];
  assign s_dadda_cla12_and_4_8 = a[4] & b[8];
  assign s_dadda_cla12_and_3_9 = a[3] & b[9];
  assign s_dadda_cla12_fa36_xor0 = s_dadda_cla12_and_5_7 ^ s_dadda_cla12_and_4_8;
  assign s_dadda_cla12_fa36_and0 = s_dadda_cla12_and_5_7 & s_dadda_cla12_and_4_8;
  assign s_dadda_cla12_fa36_xor1 = s_dadda_cla12_fa36_xor0 ^ s_dadda_cla12_and_3_9;
  assign s_dadda_cla12_fa36_and1 = s_dadda_cla12_fa36_xor0 & s_dadda_cla12_and_3_9;
  assign s_dadda_cla12_fa36_or0 = s_dadda_cla12_fa36_and0 | s_dadda_cla12_fa36_and1;
  assign s_dadda_cla12_and_2_10 = a[2] & b[10];
  assign s_dadda_cla12_nand_1_11 = ~(a[1] & b[11]);
  assign s_dadda_cla12_fa37_xor0 = s_dadda_cla12_and_2_10 ^ s_dadda_cla12_nand_1_11;
  assign s_dadda_cla12_fa37_and0 = s_dadda_cla12_and_2_10 & s_dadda_cla12_nand_1_11;
  assign s_dadda_cla12_fa37_xor1 = s_dadda_cla12_fa37_xor0 ^ s_dadda_cla12_fa3_xor1;
  assign s_dadda_cla12_fa37_and1 = s_dadda_cla12_fa37_xor0 & s_dadda_cla12_fa3_xor1;
  assign s_dadda_cla12_fa37_or0 = s_dadda_cla12_fa37_and0 | s_dadda_cla12_fa37_and1;
  assign s_dadda_cla12_fa38_xor0 = s_dadda_cla12_fa4_xor1 ^ s_dadda_cla12_fa5_xor1;
  assign s_dadda_cla12_fa38_and0 = s_dadda_cla12_fa4_xor1 & s_dadda_cla12_fa5_xor1;
  assign s_dadda_cla12_fa38_xor1 = s_dadda_cla12_fa38_xor0 ^ s_dadda_cla12_fa34_xor1;
  assign s_dadda_cla12_fa38_and1 = s_dadda_cla12_fa38_xor0 & s_dadda_cla12_fa34_xor1;
  assign s_dadda_cla12_fa38_or0 = s_dadda_cla12_fa38_and0 | s_dadda_cla12_fa38_and1;
  assign s_dadda_cla12_fa39_xor0 = s_dadda_cla12_fa38_or0 ^ s_dadda_cla12_fa37_or0;
  assign s_dadda_cla12_fa39_and0 = s_dadda_cla12_fa38_or0 & s_dadda_cla12_fa37_or0;
  assign s_dadda_cla12_fa39_xor1 = s_dadda_cla12_fa39_xor0 ^ s_dadda_cla12_fa36_or0;
  assign s_dadda_cla12_fa39_and1 = s_dadda_cla12_fa39_xor0 & s_dadda_cla12_fa36_or0;
  assign s_dadda_cla12_fa39_or0 = s_dadda_cla12_fa39_and0 | s_dadda_cla12_fa39_and1;
  assign s_dadda_cla12_and_8_5 = a[8] & b[5];
  assign s_dadda_cla12_fa40_xor0 = s_dadda_cla12_fa35_or0 ^ s_dadda_cla12_fa34_or0;
  assign s_dadda_cla12_fa40_and0 = s_dadda_cla12_fa35_or0 & s_dadda_cla12_fa34_or0;
  assign s_dadda_cla12_fa40_xor1 = s_dadda_cla12_fa40_xor0 ^ s_dadda_cla12_and_8_5;
  assign s_dadda_cla12_fa40_and1 = s_dadda_cla12_fa40_xor0 & s_dadda_cla12_and_8_5;
  assign s_dadda_cla12_fa40_or0 = s_dadda_cla12_fa40_and0 | s_dadda_cla12_fa40_and1;
  assign s_dadda_cla12_and_7_6 = a[7] & b[6];
  assign s_dadda_cla12_and_6_7 = a[6] & b[7];
  assign s_dadda_cla12_and_5_8 = a[5] & b[8];
  assign s_dadda_cla12_fa41_xor0 = s_dadda_cla12_and_7_6 ^ s_dadda_cla12_and_6_7;
  assign s_dadda_cla12_fa41_and0 = s_dadda_cla12_and_7_6 & s_dadda_cla12_and_6_7;
  assign s_dadda_cla12_fa41_xor1 = s_dadda_cla12_fa41_xor0 ^ s_dadda_cla12_and_5_8;
  assign s_dadda_cla12_fa41_and1 = s_dadda_cla12_fa41_xor0 & s_dadda_cla12_and_5_8;
  assign s_dadda_cla12_fa41_or0 = s_dadda_cla12_fa41_and0 | s_dadda_cla12_fa41_and1;
  assign s_dadda_cla12_and_4_9 = a[4] & b[9];
  assign s_dadda_cla12_and_3_10 = a[3] & b[10];
  assign s_dadda_cla12_nand_2_11 = ~(a[2] & b[11]);
  assign s_dadda_cla12_fa42_xor0 = s_dadda_cla12_and_4_9 ^ s_dadda_cla12_and_3_10;
  assign s_dadda_cla12_fa42_and0 = s_dadda_cla12_and_4_9 & s_dadda_cla12_and_3_10;
  assign s_dadda_cla12_fa42_xor1 = s_dadda_cla12_fa42_xor0 ^ s_dadda_cla12_nand_2_11;
  assign s_dadda_cla12_fa42_and1 = s_dadda_cla12_fa42_xor0 & s_dadda_cla12_nand_2_11;
  assign s_dadda_cla12_fa42_or0 = s_dadda_cla12_fa42_and0 | s_dadda_cla12_fa42_and1;
  assign s_dadda_cla12_fa43_xor0 = s_dadda_cla12_fa6_xor1 ^ s_dadda_cla12_fa7_xor1;
  assign s_dadda_cla12_fa43_and0 = s_dadda_cla12_fa6_xor1 & s_dadda_cla12_fa7_xor1;
  assign s_dadda_cla12_fa43_xor1 = s_dadda_cla12_fa43_xor0 ^ s_dadda_cla12_fa39_xor1;
  assign s_dadda_cla12_fa43_and1 = s_dadda_cla12_fa43_xor0 & s_dadda_cla12_fa39_xor1;
  assign s_dadda_cla12_fa43_or0 = s_dadda_cla12_fa43_and0 | s_dadda_cla12_fa43_and1;
  assign s_dadda_cla12_fa44_xor0 = s_dadda_cla12_fa43_or0 ^ s_dadda_cla12_fa42_or0;
  assign s_dadda_cla12_fa44_and0 = s_dadda_cla12_fa43_or0 & s_dadda_cla12_fa42_or0;
  assign s_dadda_cla12_fa44_xor1 = s_dadda_cla12_fa44_xor0 ^ s_dadda_cla12_fa41_or0;
  assign s_dadda_cla12_fa44_and1 = s_dadda_cla12_fa44_xor0 & s_dadda_cla12_fa41_or0;
  assign s_dadda_cla12_fa44_or0 = s_dadda_cla12_fa44_and0 | s_dadda_cla12_fa44_and1;
  assign s_dadda_cla12_and_10_4 = a[10] & b[4];
  assign s_dadda_cla12_fa45_xor0 = s_dadda_cla12_fa40_or0 ^ s_dadda_cla12_fa39_or0;
  assign s_dadda_cla12_fa45_and0 = s_dadda_cla12_fa40_or0 & s_dadda_cla12_fa39_or0;
  assign s_dadda_cla12_fa45_xor1 = s_dadda_cla12_fa45_xor0 ^ s_dadda_cla12_and_10_4;
  assign s_dadda_cla12_fa45_and1 = s_dadda_cla12_fa45_xor0 & s_dadda_cla12_and_10_4;
  assign s_dadda_cla12_fa45_or0 = s_dadda_cla12_fa45_and0 | s_dadda_cla12_fa45_and1;
  assign s_dadda_cla12_and_9_5 = a[9] & b[5];
  assign s_dadda_cla12_and_8_6 = a[8] & b[6];
  assign s_dadda_cla12_and_7_7 = a[7] & b[7];
  assign s_dadda_cla12_fa46_xor0 = s_dadda_cla12_and_9_5 ^ s_dadda_cla12_and_8_6;
  assign s_dadda_cla12_fa46_and0 = s_dadda_cla12_and_9_5 & s_dadda_cla12_and_8_6;
  assign s_dadda_cla12_fa46_xor1 = s_dadda_cla12_fa46_xor0 ^ s_dadda_cla12_and_7_7;
  assign s_dadda_cla12_fa46_and1 = s_dadda_cla12_fa46_xor0 & s_dadda_cla12_and_7_7;
  assign s_dadda_cla12_fa46_or0 = s_dadda_cla12_fa46_and0 | s_dadda_cla12_fa46_and1;
  assign s_dadda_cla12_and_6_8 = a[6] & b[8];
  assign s_dadda_cla12_and_5_9 = a[5] & b[9];
  assign s_dadda_cla12_and_4_10 = a[4] & b[10];
  assign s_dadda_cla12_fa47_xor0 = s_dadda_cla12_and_6_8 ^ s_dadda_cla12_and_5_9;
  assign s_dadda_cla12_fa47_and0 = s_dadda_cla12_and_6_8 & s_dadda_cla12_and_5_9;
  assign s_dadda_cla12_fa47_xor1 = s_dadda_cla12_fa47_xor0 ^ s_dadda_cla12_and_4_10;
  assign s_dadda_cla12_fa47_and1 = s_dadda_cla12_fa47_xor0 & s_dadda_cla12_and_4_10;
  assign s_dadda_cla12_fa47_or0 = s_dadda_cla12_fa47_and0 | s_dadda_cla12_fa47_and1;
  assign s_dadda_cla12_nand_3_11 = ~(a[3] & b[11]);
  assign s_dadda_cla12_fa48_xor0 = s_dadda_cla12_nand_3_11 ^ s_dadda_cla12_fa8_xor1;
  assign s_dadda_cla12_fa48_and0 = s_dadda_cla12_nand_3_11 & s_dadda_cla12_fa8_xor1;
  assign s_dadda_cla12_fa48_xor1 = s_dadda_cla12_fa48_xor0 ^ s_dadda_cla12_fa44_xor1;
  assign s_dadda_cla12_fa48_and1 = s_dadda_cla12_fa48_xor0 & s_dadda_cla12_fa44_xor1;
  assign s_dadda_cla12_fa48_or0 = s_dadda_cla12_fa48_and0 | s_dadda_cla12_fa48_and1;
  assign s_dadda_cla12_fa49_xor0 = s_dadda_cla12_fa48_or0 ^ s_dadda_cla12_fa47_or0;
  assign s_dadda_cla12_fa49_and0 = s_dadda_cla12_fa48_or0 & s_dadda_cla12_fa47_or0;
  assign s_dadda_cla12_fa49_xor1 = s_dadda_cla12_fa49_xor0 ^ s_dadda_cla12_fa46_or0;
  assign s_dadda_cla12_fa49_and1 = s_dadda_cla12_fa49_xor0 & s_dadda_cla12_fa46_or0;
  assign s_dadda_cla12_fa49_or0 = s_dadda_cla12_fa49_and0 | s_dadda_cla12_fa49_and1;
  assign s_dadda_cla12_fa50_xor0 = s_dadda_cla12_fa45_or0 ^ s_dadda_cla12_fa44_or0;
  assign s_dadda_cla12_fa50_and0 = s_dadda_cla12_fa45_or0 & s_dadda_cla12_fa44_or0;
  assign s_dadda_cla12_fa50_xor1 = s_dadda_cla12_fa50_xor0 ^ s_dadda_cla12_fa8_or0;
  assign s_dadda_cla12_fa50_and1 = s_dadda_cla12_fa50_xor0 & s_dadda_cla12_fa8_or0;
  assign s_dadda_cla12_fa50_or0 = s_dadda_cla12_fa50_and0 | s_dadda_cla12_fa50_and1;
  assign s_dadda_cla12_nand_11_4 = ~(a[11] & b[4]);
  assign s_dadda_cla12_and_10_5 = a[10] & b[5];
  assign s_dadda_cla12_and_9_6 = a[9] & b[6];
  assign s_dadda_cla12_fa51_xor0 = s_dadda_cla12_nand_11_4 ^ s_dadda_cla12_and_10_5;
  assign s_dadda_cla12_fa51_and0 = s_dadda_cla12_nand_11_4 & s_dadda_cla12_and_10_5;
  assign s_dadda_cla12_fa51_xor1 = s_dadda_cla12_fa51_xor0 ^ s_dadda_cla12_and_9_6;
  assign s_dadda_cla12_fa51_and1 = s_dadda_cla12_fa51_xor0 & s_dadda_cla12_and_9_6;
  assign s_dadda_cla12_fa51_or0 = s_dadda_cla12_fa51_and0 | s_dadda_cla12_fa51_and1;
  assign s_dadda_cla12_and_8_7 = a[8] & b[7];
  assign s_dadda_cla12_and_7_8 = a[7] & b[8];
  assign s_dadda_cla12_and_6_9 = a[6] & b[9];
  assign s_dadda_cla12_fa52_xor0 = s_dadda_cla12_and_8_7 ^ s_dadda_cla12_and_7_8;
  assign s_dadda_cla12_fa52_and0 = s_dadda_cla12_and_8_7 & s_dadda_cla12_and_7_8;
  assign s_dadda_cla12_fa52_xor1 = s_dadda_cla12_fa52_xor0 ^ s_dadda_cla12_and_6_9;
  assign s_dadda_cla12_fa52_and1 = s_dadda_cla12_fa52_xor0 & s_dadda_cla12_and_6_9;
  assign s_dadda_cla12_fa52_or0 = s_dadda_cla12_fa52_and0 | s_dadda_cla12_fa52_and1;
  assign s_dadda_cla12_and_5_10 = a[5] & b[10];
  assign s_dadda_cla12_nand_4_11 = ~(a[4] & b[11]);
  assign s_dadda_cla12_fa53_xor0 = s_dadda_cla12_and_5_10 ^ s_dadda_cla12_nand_4_11;
  assign s_dadda_cla12_fa53_and0 = s_dadda_cla12_and_5_10 & s_dadda_cla12_nand_4_11;
  assign s_dadda_cla12_fa53_xor1 = s_dadda_cla12_fa53_xor0 ^ s_dadda_cla12_fa49_xor1;
  assign s_dadda_cla12_fa53_and1 = s_dadda_cla12_fa53_xor0 & s_dadda_cla12_fa49_xor1;
  assign s_dadda_cla12_fa53_or0 = s_dadda_cla12_fa53_and0 | s_dadda_cla12_fa53_and1;
  assign s_dadda_cla12_fa54_xor0 = s_dadda_cla12_fa53_or0 ^ s_dadda_cla12_fa52_or0;
  assign s_dadda_cla12_fa54_and0 = s_dadda_cla12_fa53_or0 & s_dadda_cla12_fa52_or0;
  assign s_dadda_cla12_fa54_xor1 = s_dadda_cla12_fa54_xor0 ^ s_dadda_cla12_fa51_or0;
  assign s_dadda_cla12_fa54_and1 = s_dadda_cla12_fa54_xor0 & s_dadda_cla12_fa51_or0;
  assign s_dadda_cla12_fa54_or0 = s_dadda_cla12_fa54_and0 | s_dadda_cla12_fa54_and1;
  assign s_dadda_cla12_nand_11_5 = ~(a[11] & b[5]);
  assign s_dadda_cla12_fa55_xor0 = s_dadda_cla12_fa50_or0 ^ s_dadda_cla12_fa49_or0;
  assign s_dadda_cla12_fa55_and0 = s_dadda_cla12_fa50_or0 & s_dadda_cla12_fa49_or0;
  assign s_dadda_cla12_fa55_xor1 = s_dadda_cla12_fa55_xor0 ^ s_dadda_cla12_nand_11_5;
  assign s_dadda_cla12_fa55_and1 = s_dadda_cla12_fa55_xor0 & s_dadda_cla12_nand_11_5;
  assign s_dadda_cla12_fa55_or0 = s_dadda_cla12_fa55_and0 | s_dadda_cla12_fa55_and1;
  assign s_dadda_cla12_and_10_6 = a[10] & b[6];
  assign s_dadda_cla12_and_9_7 = a[9] & b[7];
  assign s_dadda_cla12_and_8_8 = a[8] & b[8];
  assign s_dadda_cla12_fa56_xor0 = s_dadda_cla12_and_10_6 ^ s_dadda_cla12_and_9_7;
  assign s_dadda_cla12_fa56_and0 = s_dadda_cla12_and_10_6 & s_dadda_cla12_and_9_7;
  assign s_dadda_cla12_fa56_xor1 = s_dadda_cla12_fa56_xor0 ^ s_dadda_cla12_and_8_8;
  assign s_dadda_cla12_fa56_and1 = s_dadda_cla12_fa56_xor0 & s_dadda_cla12_and_8_8;
  assign s_dadda_cla12_fa56_or0 = s_dadda_cla12_fa56_and0 | s_dadda_cla12_fa56_and1;
  assign s_dadda_cla12_and_7_9 = a[7] & b[9];
  assign s_dadda_cla12_and_6_10 = a[6] & b[10];
  assign s_dadda_cla12_nand_5_11 = ~(a[5] & b[11]);
  assign s_dadda_cla12_fa57_xor0 = s_dadda_cla12_and_7_9 ^ s_dadda_cla12_and_6_10;
  assign s_dadda_cla12_fa57_and0 = s_dadda_cla12_and_7_9 & s_dadda_cla12_and_6_10;
  assign s_dadda_cla12_fa57_xor1 = s_dadda_cla12_fa57_xor0 ^ s_dadda_cla12_nand_5_11;
  assign s_dadda_cla12_fa57_and1 = s_dadda_cla12_fa57_xor0 & s_dadda_cla12_nand_5_11;
  assign s_dadda_cla12_fa57_or0 = s_dadda_cla12_fa57_and0 | s_dadda_cla12_fa57_and1;
  assign s_dadda_cla12_fa58_xor0 = s_dadda_cla12_fa57_or0 ^ s_dadda_cla12_fa56_or0;
  assign s_dadda_cla12_fa58_and0 = s_dadda_cla12_fa57_or0 & s_dadda_cla12_fa56_or0;
  assign s_dadda_cla12_fa58_xor1 = s_dadda_cla12_fa58_xor0 ^ s_dadda_cla12_fa55_or0;
  assign s_dadda_cla12_fa58_and1 = s_dadda_cla12_fa58_xor0 & s_dadda_cla12_fa55_or0;
  assign s_dadda_cla12_fa58_or0 = s_dadda_cla12_fa58_and0 | s_dadda_cla12_fa58_and1;
  assign s_dadda_cla12_nand_11_6 = ~(a[11] & b[6]);
  assign s_dadda_cla12_and_10_7 = a[10] & b[7];
  assign s_dadda_cla12_fa59_xor0 = s_dadda_cla12_fa54_or0 ^ s_dadda_cla12_nand_11_6;
  assign s_dadda_cla12_fa59_and0 = s_dadda_cla12_fa54_or0 & s_dadda_cla12_nand_11_6;
  assign s_dadda_cla12_fa59_xor1 = s_dadda_cla12_fa59_xor0 ^ s_dadda_cla12_and_10_7;
  assign s_dadda_cla12_fa59_and1 = s_dadda_cla12_fa59_xor0 & s_dadda_cla12_and_10_7;
  assign s_dadda_cla12_fa59_or0 = s_dadda_cla12_fa59_and0 | s_dadda_cla12_fa59_and1;
  assign s_dadda_cla12_and_9_8 = a[9] & b[8];
  assign s_dadda_cla12_and_8_9 = a[8] & b[9];
  assign s_dadda_cla12_and_7_10 = a[7] & b[10];
  assign s_dadda_cla12_fa60_xor0 = s_dadda_cla12_and_9_8 ^ s_dadda_cla12_and_8_9;
  assign s_dadda_cla12_fa60_and0 = s_dadda_cla12_and_9_8 & s_dadda_cla12_and_8_9;
  assign s_dadda_cla12_fa60_xor1 = s_dadda_cla12_fa60_xor0 ^ s_dadda_cla12_and_7_10;
  assign s_dadda_cla12_fa60_and1 = s_dadda_cla12_fa60_xor0 & s_dadda_cla12_and_7_10;
  assign s_dadda_cla12_fa60_or0 = s_dadda_cla12_fa60_and0 | s_dadda_cla12_fa60_and1;
  assign s_dadda_cla12_fa61_xor0 = s_dadda_cla12_fa60_or0 ^ s_dadda_cla12_fa59_or0;
  assign s_dadda_cla12_fa61_and0 = s_dadda_cla12_fa60_or0 & s_dadda_cla12_fa59_or0;
  assign s_dadda_cla12_fa61_xor1 = s_dadda_cla12_fa61_xor0 ^ s_dadda_cla12_fa58_or0;
  assign s_dadda_cla12_fa61_and1 = s_dadda_cla12_fa61_xor0 & s_dadda_cla12_fa58_or0;
  assign s_dadda_cla12_fa61_or0 = s_dadda_cla12_fa61_and0 | s_dadda_cla12_fa61_and1;
  assign s_dadda_cla12_nand_11_7 = ~(a[11] & b[7]);
  assign s_dadda_cla12_and_10_8 = a[10] & b[8];
  assign s_dadda_cla12_and_9_9 = a[9] & b[9];
  assign s_dadda_cla12_fa62_xor0 = s_dadda_cla12_nand_11_7 ^ s_dadda_cla12_and_10_8;
  assign s_dadda_cla12_fa62_and0 = s_dadda_cla12_nand_11_7 & s_dadda_cla12_and_10_8;
  assign s_dadda_cla12_fa62_xor1 = s_dadda_cla12_fa62_xor0 ^ s_dadda_cla12_and_9_9;
  assign s_dadda_cla12_fa62_and1 = s_dadda_cla12_fa62_xor0 & s_dadda_cla12_and_9_9;
  assign s_dadda_cla12_fa62_or0 = s_dadda_cla12_fa62_and0 | s_dadda_cla12_fa62_and1;
  assign s_dadda_cla12_nand_11_8 = ~(a[11] & b[8]);
  assign s_dadda_cla12_fa63_xor0 = s_dadda_cla12_fa62_or0 ^ s_dadda_cla12_fa61_or0;
  assign s_dadda_cla12_fa63_and0 = s_dadda_cla12_fa62_or0 & s_dadda_cla12_fa61_or0;
  assign s_dadda_cla12_fa63_xor1 = s_dadda_cla12_fa63_xor0 ^ s_dadda_cla12_nand_11_8;
  assign s_dadda_cla12_fa63_and1 = s_dadda_cla12_fa63_xor0 & s_dadda_cla12_nand_11_8;
  assign s_dadda_cla12_fa63_or0 = s_dadda_cla12_fa63_and0 | s_dadda_cla12_fa63_and1;
  assign s_dadda_cla12_and_3_0 = a[3] & b[0];
  assign s_dadda_cla12_and_2_1 = a[2] & b[1];
  assign s_dadda_cla12_ha8_xor0 = s_dadda_cla12_and_3_0 ^ s_dadda_cla12_and_2_1;
  assign s_dadda_cla12_ha8_and0 = s_dadda_cla12_and_3_0 & s_dadda_cla12_and_2_1;
  assign s_dadda_cla12_and_2_2 = a[2] & b[2];
  assign s_dadda_cla12_and_1_3 = a[1] & b[3];
  assign s_dadda_cla12_fa64_xor0 = s_dadda_cla12_ha8_and0 ^ s_dadda_cla12_and_2_2;
  assign s_dadda_cla12_fa64_and0 = s_dadda_cla12_ha8_and0 & s_dadda_cla12_and_2_2;
  assign s_dadda_cla12_fa64_xor1 = s_dadda_cla12_fa64_xor0 ^ s_dadda_cla12_and_1_3;
  assign s_dadda_cla12_fa64_and1 = s_dadda_cla12_fa64_xor0 & s_dadda_cla12_and_1_3;
  assign s_dadda_cla12_fa64_or0 = s_dadda_cla12_fa64_and0 | s_dadda_cla12_fa64_and1;
  assign s_dadda_cla12_and_1_4 = a[1] & b[4];
  assign s_dadda_cla12_and_0_5 = a[0] & b[5];
  assign s_dadda_cla12_fa65_xor0 = s_dadda_cla12_fa64_or0 ^ s_dadda_cla12_and_1_4;
  assign s_dadda_cla12_fa65_and0 = s_dadda_cla12_fa64_or0 & s_dadda_cla12_and_1_4;
  assign s_dadda_cla12_fa65_xor1 = s_dadda_cla12_fa65_xor0 ^ s_dadda_cla12_and_0_5;
  assign s_dadda_cla12_fa65_and1 = s_dadda_cla12_fa65_xor0 & s_dadda_cla12_and_0_5;
  assign s_dadda_cla12_fa65_or0 = s_dadda_cla12_fa65_and0 | s_dadda_cla12_fa65_and1;
  assign s_dadda_cla12_and_0_6 = a[0] & b[6];
  assign s_dadda_cla12_fa66_xor0 = s_dadda_cla12_fa65_or0 ^ s_dadda_cla12_and_0_6;
  assign s_dadda_cla12_fa66_and0 = s_dadda_cla12_fa65_or0 & s_dadda_cla12_and_0_6;
  assign s_dadda_cla12_fa66_xor1 = s_dadda_cla12_fa66_xor0 ^ s_dadda_cla12_fa10_xor1;
  assign s_dadda_cla12_fa66_and1 = s_dadda_cla12_fa66_xor0 & s_dadda_cla12_fa10_xor1;
  assign s_dadda_cla12_fa66_or0 = s_dadda_cla12_fa66_and0 | s_dadda_cla12_fa66_and1;
  assign s_dadda_cla12_fa67_xor0 = s_dadda_cla12_fa66_or0 ^ s_dadda_cla12_fa12_xor1;
  assign s_dadda_cla12_fa67_and0 = s_dadda_cla12_fa66_or0 & s_dadda_cla12_fa12_xor1;
  assign s_dadda_cla12_fa67_xor1 = s_dadda_cla12_fa67_xor0 ^ s_dadda_cla12_fa13_xor1;
  assign s_dadda_cla12_fa67_and1 = s_dadda_cla12_fa67_xor0 & s_dadda_cla12_fa13_xor1;
  assign s_dadda_cla12_fa67_or0 = s_dadda_cla12_fa67_and0 | s_dadda_cla12_fa67_and1;
  assign s_dadda_cla12_fa68_xor0 = s_dadda_cla12_fa67_or0 ^ s_dadda_cla12_fa16_xor1;
  assign s_dadda_cla12_fa68_and0 = s_dadda_cla12_fa67_or0 & s_dadda_cla12_fa16_xor1;
  assign s_dadda_cla12_fa68_xor1 = s_dadda_cla12_fa68_xor0 ^ s_dadda_cla12_fa17_xor1;
  assign s_dadda_cla12_fa68_and1 = s_dadda_cla12_fa68_xor0 & s_dadda_cla12_fa17_xor1;
  assign s_dadda_cla12_fa68_or0 = s_dadda_cla12_fa68_and0 | s_dadda_cla12_fa68_and1;
  assign s_dadda_cla12_fa69_xor0 = s_dadda_cla12_fa68_or0 ^ s_dadda_cla12_fa20_xor1;
  assign s_dadda_cla12_fa69_and0 = s_dadda_cla12_fa68_or0 & s_dadda_cla12_fa20_xor1;
  assign s_dadda_cla12_fa69_xor1 = s_dadda_cla12_fa69_xor0 ^ s_dadda_cla12_fa21_xor1;
  assign s_dadda_cla12_fa69_and1 = s_dadda_cla12_fa69_xor0 & s_dadda_cla12_fa21_xor1;
  assign s_dadda_cla12_fa69_or0 = s_dadda_cla12_fa69_and0 | s_dadda_cla12_fa69_and1;
  assign s_dadda_cla12_fa70_xor0 = s_dadda_cla12_fa69_or0 ^ s_dadda_cla12_fa25_xor1;
  assign s_dadda_cla12_fa70_and0 = s_dadda_cla12_fa69_or0 & s_dadda_cla12_fa25_xor1;
  assign s_dadda_cla12_fa70_xor1 = s_dadda_cla12_fa70_xor0 ^ s_dadda_cla12_fa26_xor1;
  assign s_dadda_cla12_fa70_and1 = s_dadda_cla12_fa70_xor0 & s_dadda_cla12_fa26_xor1;
  assign s_dadda_cla12_fa70_or0 = s_dadda_cla12_fa70_and0 | s_dadda_cla12_fa70_and1;
  assign s_dadda_cla12_fa71_xor0 = s_dadda_cla12_fa70_or0 ^ s_dadda_cla12_fa30_xor1;
  assign s_dadda_cla12_fa71_and0 = s_dadda_cla12_fa70_or0 & s_dadda_cla12_fa30_xor1;
  assign s_dadda_cla12_fa71_xor1 = s_dadda_cla12_fa71_xor0 ^ s_dadda_cla12_fa31_xor1;
  assign s_dadda_cla12_fa71_and1 = s_dadda_cla12_fa71_xor0 & s_dadda_cla12_fa31_xor1;
  assign s_dadda_cla12_fa71_or0 = s_dadda_cla12_fa71_and0 | s_dadda_cla12_fa71_and1;
  assign s_dadda_cla12_fa72_xor0 = s_dadda_cla12_fa71_or0 ^ s_dadda_cla12_fa35_xor1;
  assign s_dadda_cla12_fa72_and0 = s_dadda_cla12_fa71_or0 & s_dadda_cla12_fa35_xor1;
  assign s_dadda_cla12_fa72_xor1 = s_dadda_cla12_fa72_xor0 ^ s_dadda_cla12_fa36_xor1;
  assign s_dadda_cla12_fa72_and1 = s_dadda_cla12_fa72_xor0 & s_dadda_cla12_fa36_xor1;
  assign s_dadda_cla12_fa72_or0 = s_dadda_cla12_fa72_and0 | s_dadda_cla12_fa72_and1;
  assign s_dadda_cla12_fa73_xor0 = s_dadda_cla12_fa72_or0 ^ s_dadda_cla12_fa40_xor1;
  assign s_dadda_cla12_fa73_and0 = s_dadda_cla12_fa72_or0 & s_dadda_cla12_fa40_xor1;
  assign s_dadda_cla12_fa73_xor1 = s_dadda_cla12_fa73_xor0 ^ s_dadda_cla12_fa41_xor1;
  assign s_dadda_cla12_fa73_and1 = s_dadda_cla12_fa73_xor0 & s_dadda_cla12_fa41_xor1;
  assign s_dadda_cla12_fa73_or0 = s_dadda_cla12_fa73_and0 | s_dadda_cla12_fa73_and1;
  assign s_dadda_cla12_fa74_xor0 = s_dadda_cla12_fa73_or0 ^ s_dadda_cla12_fa45_xor1;
  assign s_dadda_cla12_fa74_and0 = s_dadda_cla12_fa73_or0 & s_dadda_cla12_fa45_xor1;
  assign s_dadda_cla12_fa74_xor1 = s_dadda_cla12_fa74_xor0 ^ s_dadda_cla12_fa46_xor1;
  assign s_dadda_cla12_fa74_and1 = s_dadda_cla12_fa74_xor0 & s_dadda_cla12_fa46_xor1;
  assign s_dadda_cla12_fa74_or0 = s_dadda_cla12_fa74_and0 | s_dadda_cla12_fa74_and1;
  assign s_dadda_cla12_fa75_xor0 = s_dadda_cla12_fa74_or0 ^ s_dadda_cla12_fa50_xor1;
  assign s_dadda_cla12_fa75_and0 = s_dadda_cla12_fa74_or0 & s_dadda_cla12_fa50_xor1;
  assign s_dadda_cla12_fa75_xor1 = s_dadda_cla12_fa75_xor0 ^ s_dadda_cla12_fa51_xor1;
  assign s_dadda_cla12_fa75_and1 = s_dadda_cla12_fa75_xor0 & s_dadda_cla12_fa51_xor1;
  assign s_dadda_cla12_fa75_or0 = s_dadda_cla12_fa75_and0 | s_dadda_cla12_fa75_and1;
  assign s_dadda_cla12_fa76_xor0 = s_dadda_cla12_fa75_or0 ^ s_dadda_cla12_fa54_xor1;
  assign s_dadda_cla12_fa76_and0 = s_dadda_cla12_fa75_or0 & s_dadda_cla12_fa54_xor1;
  assign s_dadda_cla12_fa76_xor1 = s_dadda_cla12_fa76_xor0 ^ s_dadda_cla12_fa55_xor1;
  assign s_dadda_cla12_fa76_and1 = s_dadda_cla12_fa76_xor0 & s_dadda_cla12_fa55_xor1;
  assign s_dadda_cla12_fa76_or0 = s_dadda_cla12_fa76_and0 | s_dadda_cla12_fa76_and1;
  assign s_dadda_cla12_nand_6_11 = ~(a[6] & b[11]);
  assign s_dadda_cla12_fa77_xor0 = s_dadda_cla12_fa76_or0 ^ s_dadda_cla12_nand_6_11;
  assign s_dadda_cla12_fa77_and0 = s_dadda_cla12_fa76_or0 & s_dadda_cla12_nand_6_11;
  assign s_dadda_cla12_fa77_xor1 = s_dadda_cla12_fa77_xor0 ^ s_dadda_cla12_fa58_xor1;
  assign s_dadda_cla12_fa77_and1 = s_dadda_cla12_fa77_xor0 & s_dadda_cla12_fa58_xor1;
  assign s_dadda_cla12_fa77_or0 = s_dadda_cla12_fa77_and0 | s_dadda_cla12_fa77_and1;
  assign s_dadda_cla12_and_8_10 = a[8] & b[10];
  assign s_dadda_cla12_nand_7_11 = ~(a[7] & b[11]);
  assign s_dadda_cla12_fa78_xor0 = s_dadda_cla12_fa77_or0 ^ s_dadda_cla12_and_8_10;
  assign s_dadda_cla12_fa78_and0 = s_dadda_cla12_fa77_or0 & s_dadda_cla12_and_8_10;
  assign s_dadda_cla12_fa78_xor1 = s_dadda_cla12_fa78_xor0 ^ s_dadda_cla12_nand_7_11;
  assign s_dadda_cla12_fa78_and1 = s_dadda_cla12_fa78_xor0 & s_dadda_cla12_nand_7_11;
  assign s_dadda_cla12_fa78_or0 = s_dadda_cla12_fa78_and0 | s_dadda_cla12_fa78_and1;
  assign s_dadda_cla12_and_10_9 = a[10] & b[9];
  assign s_dadda_cla12_and_9_10 = a[9] & b[10];
  assign s_dadda_cla12_fa79_xor0 = s_dadda_cla12_fa78_or0 ^ s_dadda_cla12_and_10_9;
  assign s_dadda_cla12_fa79_and0 = s_dadda_cla12_fa78_or0 & s_dadda_cla12_and_10_9;
  assign s_dadda_cla12_fa79_xor1 = s_dadda_cla12_fa79_xor0 ^ s_dadda_cla12_and_9_10;
  assign s_dadda_cla12_fa79_and1 = s_dadda_cla12_fa79_xor0 & s_dadda_cla12_and_9_10;
  assign s_dadda_cla12_fa79_or0 = s_dadda_cla12_fa79_and0 | s_dadda_cla12_fa79_and1;
  assign s_dadda_cla12_nand_11_9 = ~(a[11] & b[9]);
  assign s_dadda_cla12_fa80_xor0 = s_dadda_cla12_fa79_or0 ^ s_dadda_cla12_fa63_or0;
  assign s_dadda_cla12_fa80_and0 = s_dadda_cla12_fa79_or0 & s_dadda_cla12_fa63_or0;
  assign s_dadda_cla12_fa80_xor1 = s_dadda_cla12_fa80_xor0 ^ s_dadda_cla12_nand_11_9;
  assign s_dadda_cla12_fa80_and1 = s_dadda_cla12_fa80_xor0 & s_dadda_cla12_nand_11_9;
  assign s_dadda_cla12_fa80_or0 = s_dadda_cla12_fa80_and0 | s_dadda_cla12_fa80_and1;
  assign s_dadda_cla12_and_2_0 = a[2] & b[0];
  assign s_dadda_cla12_and_1_1 = a[1] & b[1];
  assign s_dadda_cla12_ha9_xor0 = s_dadda_cla12_and_2_0 ^ s_dadda_cla12_and_1_1;
  assign s_dadda_cla12_ha9_and0 = s_dadda_cla12_and_2_0 & s_dadda_cla12_and_1_1;
  assign s_dadda_cla12_and_1_2 = a[1] & b[2];
  assign s_dadda_cla12_and_0_3 = a[0] & b[3];
  assign s_dadda_cla12_fa81_xor0 = s_dadda_cla12_ha9_and0 ^ s_dadda_cla12_and_1_2;
  assign s_dadda_cla12_fa81_and0 = s_dadda_cla12_ha9_and0 & s_dadda_cla12_and_1_2;
  assign s_dadda_cla12_fa81_xor1 = s_dadda_cla12_fa81_xor0 ^ s_dadda_cla12_and_0_3;
  assign s_dadda_cla12_fa81_and1 = s_dadda_cla12_fa81_xor0 & s_dadda_cla12_and_0_3;
  assign s_dadda_cla12_fa81_or0 = s_dadda_cla12_fa81_and0 | s_dadda_cla12_fa81_and1;
  assign s_dadda_cla12_and_0_4 = a[0] & b[4];
  assign s_dadda_cla12_fa82_xor0 = s_dadda_cla12_fa81_or0 ^ s_dadda_cla12_and_0_4;
  assign s_dadda_cla12_fa82_and0 = s_dadda_cla12_fa81_or0 & s_dadda_cla12_and_0_4;
  assign s_dadda_cla12_fa82_xor1 = s_dadda_cla12_fa82_xor0 ^ s_dadda_cla12_ha3_xor0;
  assign s_dadda_cla12_fa82_and1 = s_dadda_cla12_fa82_xor0 & s_dadda_cla12_ha3_xor0;
  assign s_dadda_cla12_fa82_or0 = s_dadda_cla12_fa82_and0 | s_dadda_cla12_fa82_and1;
  assign s_dadda_cla12_fa83_xor0 = s_dadda_cla12_fa82_or0 ^ s_dadda_cla12_fa9_xor1;
  assign s_dadda_cla12_fa83_and0 = s_dadda_cla12_fa82_or0 & s_dadda_cla12_fa9_xor1;
  assign s_dadda_cla12_fa83_xor1 = s_dadda_cla12_fa83_xor0 ^ s_dadda_cla12_ha4_xor0;
  assign s_dadda_cla12_fa83_and1 = s_dadda_cla12_fa83_xor0 & s_dadda_cla12_ha4_xor0;
  assign s_dadda_cla12_fa83_or0 = s_dadda_cla12_fa83_and0 | s_dadda_cla12_fa83_and1;
  assign s_dadda_cla12_fa84_xor0 = s_dadda_cla12_fa83_or0 ^ s_dadda_cla12_fa11_xor1;
  assign s_dadda_cla12_fa84_and0 = s_dadda_cla12_fa83_or0 & s_dadda_cla12_fa11_xor1;
  assign s_dadda_cla12_fa84_xor1 = s_dadda_cla12_fa84_xor0 ^ s_dadda_cla12_ha5_xor0;
  assign s_dadda_cla12_fa84_and1 = s_dadda_cla12_fa84_xor0 & s_dadda_cla12_ha5_xor0;
  assign s_dadda_cla12_fa84_or0 = s_dadda_cla12_fa84_and0 | s_dadda_cla12_fa84_and1;
  assign s_dadda_cla12_fa85_xor0 = s_dadda_cla12_fa84_or0 ^ s_dadda_cla12_fa14_xor1;
  assign s_dadda_cla12_fa85_and0 = s_dadda_cla12_fa84_or0 & s_dadda_cla12_fa14_xor1;
  assign s_dadda_cla12_fa85_xor1 = s_dadda_cla12_fa85_xor0 ^ s_dadda_cla12_ha6_xor0;
  assign s_dadda_cla12_fa85_and1 = s_dadda_cla12_fa85_xor0 & s_dadda_cla12_ha6_xor0;
  assign s_dadda_cla12_fa85_or0 = s_dadda_cla12_fa85_and0 | s_dadda_cla12_fa85_and1;
  assign s_dadda_cla12_fa86_xor0 = s_dadda_cla12_fa85_or0 ^ s_dadda_cla12_fa18_xor1;
  assign s_dadda_cla12_fa86_and0 = s_dadda_cla12_fa85_or0 & s_dadda_cla12_fa18_xor1;
  assign s_dadda_cla12_fa86_xor1 = s_dadda_cla12_fa86_xor0 ^ s_dadda_cla12_ha7_xor0;
  assign s_dadda_cla12_fa86_and1 = s_dadda_cla12_fa86_xor0 & s_dadda_cla12_ha7_xor0;
  assign s_dadda_cla12_fa86_or0 = s_dadda_cla12_fa86_and0 | s_dadda_cla12_fa86_and1;
  assign s_dadda_cla12_fa87_xor0 = s_dadda_cla12_fa86_or0 ^ s_dadda_cla12_fa22_xor1;
  assign s_dadda_cla12_fa87_and0 = s_dadda_cla12_fa86_or0 & s_dadda_cla12_fa22_xor1;
  assign s_dadda_cla12_fa87_xor1 = s_dadda_cla12_fa87_xor0 ^ s_dadda_cla12_fa23_xor1;
  assign s_dadda_cla12_fa87_and1 = s_dadda_cla12_fa87_xor0 & s_dadda_cla12_fa23_xor1;
  assign s_dadda_cla12_fa87_or0 = s_dadda_cla12_fa87_and0 | s_dadda_cla12_fa87_and1;
  assign s_dadda_cla12_fa88_xor0 = s_dadda_cla12_fa87_or0 ^ s_dadda_cla12_fa27_xor1;
  assign s_dadda_cla12_fa88_and0 = s_dadda_cla12_fa87_or0 & s_dadda_cla12_fa27_xor1;
  assign s_dadda_cla12_fa88_xor1 = s_dadda_cla12_fa88_xor0 ^ s_dadda_cla12_fa28_xor1;
  assign s_dadda_cla12_fa88_and1 = s_dadda_cla12_fa88_xor0 & s_dadda_cla12_fa28_xor1;
  assign s_dadda_cla12_fa88_or0 = s_dadda_cla12_fa88_and0 | s_dadda_cla12_fa88_and1;
  assign s_dadda_cla12_fa89_xor0 = s_dadda_cla12_fa88_or0 ^ s_dadda_cla12_fa32_xor1;
  assign s_dadda_cla12_fa89_and0 = s_dadda_cla12_fa88_or0 & s_dadda_cla12_fa32_xor1;
  assign s_dadda_cla12_fa89_xor1 = s_dadda_cla12_fa89_xor0 ^ s_dadda_cla12_fa33_xor1;
  assign s_dadda_cla12_fa89_and1 = s_dadda_cla12_fa89_xor0 & s_dadda_cla12_fa33_xor1;
  assign s_dadda_cla12_fa89_or0 = s_dadda_cla12_fa89_and0 | s_dadda_cla12_fa89_and1;
  assign s_dadda_cla12_fa90_xor0 = s_dadda_cla12_fa89_or0 ^ s_dadda_cla12_fa37_xor1;
  assign s_dadda_cla12_fa90_and0 = s_dadda_cla12_fa89_or0 & s_dadda_cla12_fa37_xor1;
  assign s_dadda_cla12_fa90_xor1 = s_dadda_cla12_fa90_xor0 ^ s_dadda_cla12_fa38_xor1;
  assign s_dadda_cla12_fa90_and1 = s_dadda_cla12_fa90_xor0 & s_dadda_cla12_fa38_xor1;
  assign s_dadda_cla12_fa90_or0 = s_dadda_cla12_fa90_and0 | s_dadda_cla12_fa90_and1;
  assign s_dadda_cla12_fa91_xor0 = s_dadda_cla12_fa90_or0 ^ s_dadda_cla12_fa42_xor1;
  assign s_dadda_cla12_fa91_and0 = s_dadda_cla12_fa90_or0 & s_dadda_cla12_fa42_xor1;
  assign s_dadda_cla12_fa91_xor1 = s_dadda_cla12_fa91_xor0 ^ s_dadda_cla12_fa43_xor1;
  assign s_dadda_cla12_fa91_and1 = s_dadda_cla12_fa91_xor0 & s_dadda_cla12_fa43_xor1;
  assign s_dadda_cla12_fa91_or0 = s_dadda_cla12_fa91_and0 | s_dadda_cla12_fa91_and1;
  assign s_dadda_cla12_fa92_xor0 = s_dadda_cla12_fa91_or0 ^ s_dadda_cla12_fa47_xor1;
  assign s_dadda_cla12_fa92_and0 = s_dadda_cla12_fa91_or0 & s_dadda_cla12_fa47_xor1;
  assign s_dadda_cla12_fa92_xor1 = s_dadda_cla12_fa92_xor0 ^ s_dadda_cla12_fa48_xor1;
  assign s_dadda_cla12_fa92_and1 = s_dadda_cla12_fa92_xor0 & s_dadda_cla12_fa48_xor1;
  assign s_dadda_cla12_fa92_or0 = s_dadda_cla12_fa92_and0 | s_dadda_cla12_fa92_and1;
  assign s_dadda_cla12_fa93_xor0 = s_dadda_cla12_fa92_or0 ^ s_dadda_cla12_fa52_xor1;
  assign s_dadda_cla12_fa93_and0 = s_dadda_cla12_fa92_or0 & s_dadda_cla12_fa52_xor1;
  assign s_dadda_cla12_fa93_xor1 = s_dadda_cla12_fa93_xor0 ^ s_dadda_cla12_fa53_xor1;
  assign s_dadda_cla12_fa93_and1 = s_dadda_cla12_fa93_xor0 & s_dadda_cla12_fa53_xor1;
  assign s_dadda_cla12_fa93_or0 = s_dadda_cla12_fa93_and0 | s_dadda_cla12_fa93_and1;
  assign s_dadda_cla12_fa94_xor0 = s_dadda_cla12_fa93_or0 ^ s_dadda_cla12_fa56_xor1;
  assign s_dadda_cla12_fa94_and0 = s_dadda_cla12_fa93_or0 & s_dadda_cla12_fa56_xor1;
  assign s_dadda_cla12_fa94_xor1 = s_dadda_cla12_fa94_xor0 ^ s_dadda_cla12_fa57_xor1;
  assign s_dadda_cla12_fa94_and1 = s_dadda_cla12_fa94_xor0 & s_dadda_cla12_fa57_xor1;
  assign s_dadda_cla12_fa94_or0 = s_dadda_cla12_fa94_and0 | s_dadda_cla12_fa94_and1;
  assign s_dadda_cla12_fa95_xor0 = s_dadda_cla12_fa94_or0 ^ s_dadda_cla12_fa59_xor1;
  assign s_dadda_cla12_fa95_and0 = s_dadda_cla12_fa94_or0 & s_dadda_cla12_fa59_xor1;
  assign s_dadda_cla12_fa95_xor1 = s_dadda_cla12_fa95_xor0 ^ s_dadda_cla12_fa60_xor1;
  assign s_dadda_cla12_fa95_and1 = s_dadda_cla12_fa95_xor0 & s_dadda_cla12_fa60_xor1;
  assign s_dadda_cla12_fa95_or0 = s_dadda_cla12_fa95_and0 | s_dadda_cla12_fa95_and1;
  assign s_dadda_cla12_fa96_xor0 = s_dadda_cla12_fa95_or0 ^ s_dadda_cla12_fa61_xor1;
  assign s_dadda_cla12_fa96_and0 = s_dadda_cla12_fa95_or0 & s_dadda_cla12_fa61_xor1;
  assign s_dadda_cla12_fa96_xor1 = s_dadda_cla12_fa96_xor0 ^ s_dadda_cla12_fa62_xor1;
  assign s_dadda_cla12_fa96_and1 = s_dadda_cla12_fa96_xor0 & s_dadda_cla12_fa62_xor1;
  assign s_dadda_cla12_fa96_or0 = s_dadda_cla12_fa96_and0 | s_dadda_cla12_fa96_and1;
  assign s_dadda_cla12_nand_8_11 = ~(a[8] & b[11]);
  assign s_dadda_cla12_fa97_xor0 = s_dadda_cla12_fa96_or0 ^ s_dadda_cla12_nand_8_11;
  assign s_dadda_cla12_fa97_and0 = s_dadda_cla12_fa96_or0 & s_dadda_cla12_nand_8_11;
  assign s_dadda_cla12_fa97_xor1 = s_dadda_cla12_fa97_xor0 ^ s_dadda_cla12_fa63_xor1;
  assign s_dadda_cla12_fa97_and1 = s_dadda_cla12_fa97_xor0 & s_dadda_cla12_fa63_xor1;
  assign s_dadda_cla12_fa97_or0 = s_dadda_cla12_fa97_and0 | s_dadda_cla12_fa97_and1;
  assign s_dadda_cla12_and_10_10 = a[10] & b[10];
  assign s_dadda_cla12_nand_9_11 = ~(a[9] & b[11]);
  assign s_dadda_cla12_fa98_xor0 = s_dadda_cla12_fa97_or0 ^ s_dadda_cla12_and_10_10;
  assign s_dadda_cla12_fa98_and0 = s_dadda_cla12_fa97_or0 & s_dadda_cla12_and_10_10;
  assign s_dadda_cla12_fa98_xor1 = s_dadda_cla12_fa98_xor0 ^ s_dadda_cla12_nand_9_11;
  assign s_dadda_cla12_fa98_and1 = s_dadda_cla12_fa98_xor0 & s_dadda_cla12_nand_9_11;
  assign s_dadda_cla12_fa98_or0 = s_dadda_cla12_fa98_and0 | s_dadda_cla12_fa98_and1;
  assign s_dadda_cla12_nand_11_10 = ~(a[11] & b[10]);
  assign s_dadda_cla12_fa99_xor0 = s_dadda_cla12_fa98_or0 ^ s_dadda_cla12_fa80_or0;
  assign s_dadda_cla12_fa99_and0 = s_dadda_cla12_fa98_or0 & s_dadda_cla12_fa80_or0;
  assign s_dadda_cla12_fa99_xor1 = s_dadda_cla12_fa99_xor0 ^ s_dadda_cla12_nand_11_10;
  assign s_dadda_cla12_fa99_and1 = s_dadda_cla12_fa99_xor0 & s_dadda_cla12_nand_11_10;
  assign s_dadda_cla12_fa99_or0 = s_dadda_cla12_fa99_and0 | s_dadda_cla12_fa99_and1;
  assign s_dadda_cla12_and_0_0 = a[0] & b[0];
  assign s_dadda_cla12_and_1_0 = a[1] & b[0];
  assign s_dadda_cla12_and_0_2 = a[0] & b[2];
  assign s_dadda_cla12_nand_10_11 = ~(a[10] & b[11]);
  assign s_dadda_cla12_and_0_1 = a[0] & b[1];
  assign s_dadda_cla12_and_11_11 = a[11] & b[11];
  assign s_dadda_cla12_u_cla22_pg_logic0_or0 = s_dadda_cla12_and_1_0 | s_dadda_cla12_and_0_1;
  assign s_dadda_cla12_u_cla22_pg_logic0_and0 = s_dadda_cla12_and_1_0 & s_dadda_cla12_and_0_1;
  assign s_dadda_cla12_u_cla22_pg_logic0_xor0 = s_dadda_cla12_and_1_0 ^ s_dadda_cla12_and_0_1;
  assign s_dadda_cla12_u_cla22_pg_logic1_or0 = s_dadda_cla12_and_0_2 | s_dadda_cla12_ha9_xor0;
  assign s_dadda_cla12_u_cla22_pg_logic1_and0 = s_dadda_cla12_and_0_2 & s_dadda_cla12_ha9_xor0;
  assign s_dadda_cla12_u_cla22_pg_logic1_xor0 = s_dadda_cla12_and_0_2 ^ s_dadda_cla12_ha9_xor0;
  assign s_dadda_cla12_u_cla22_xor1 = s_dadda_cla12_u_cla22_pg_logic1_xor0 ^ s_dadda_cla12_u_cla22_pg_logic0_and0;
  assign s_dadda_cla12_u_cla22_and0 = s_dadda_cla12_u_cla22_pg_logic0_and0 & s_dadda_cla12_u_cla22_pg_logic1_or0;
  assign s_dadda_cla12_u_cla22_or0 = s_dadda_cla12_u_cla22_pg_logic1_and0 | s_dadda_cla12_u_cla22_and0;
  assign s_dadda_cla12_u_cla22_pg_logic2_or0 = s_dadda_cla12_ha8_xor0 | s_dadda_cla12_fa81_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic2_and0 = s_dadda_cla12_ha8_xor0 & s_dadda_cla12_fa81_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic2_xor0 = s_dadda_cla12_ha8_xor0 ^ s_dadda_cla12_fa81_xor1;
  assign s_dadda_cla12_u_cla22_xor2 = s_dadda_cla12_u_cla22_pg_logic2_xor0 ^ s_dadda_cla12_u_cla22_or0;
  assign s_dadda_cla12_u_cla22_and1 = s_dadda_cla12_u_cla22_pg_logic2_or0 & s_dadda_cla12_u_cla22_pg_logic0_or0;
  assign s_dadda_cla12_u_cla22_and2 = s_dadda_cla12_u_cla22_pg_logic0_and0 & s_dadda_cla12_u_cla22_pg_logic2_or0;
  assign s_dadda_cla12_u_cla22_and3 = s_dadda_cla12_u_cla22_and2 & s_dadda_cla12_u_cla22_pg_logic1_or0;
  assign s_dadda_cla12_u_cla22_and4 = s_dadda_cla12_u_cla22_pg_logic1_and0 & s_dadda_cla12_u_cla22_pg_logic2_or0;
  assign s_dadda_cla12_u_cla22_or1 = s_dadda_cla12_u_cla22_and3 | s_dadda_cla12_u_cla22_and4;
  assign s_dadda_cla12_u_cla22_or2 = s_dadda_cla12_u_cla22_pg_logic2_and0 | s_dadda_cla12_u_cla22_or1;
  assign s_dadda_cla12_u_cla22_pg_logic3_or0 = s_dadda_cla12_fa64_xor1 | s_dadda_cla12_fa82_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic3_and0 = s_dadda_cla12_fa64_xor1 & s_dadda_cla12_fa82_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic3_xor0 = s_dadda_cla12_fa64_xor1 ^ s_dadda_cla12_fa82_xor1;
  assign s_dadda_cla12_u_cla22_xor3 = s_dadda_cla12_u_cla22_pg_logic3_xor0 ^ s_dadda_cla12_u_cla22_or2;
  assign s_dadda_cla12_u_cla22_and5 = s_dadda_cla12_u_cla22_pg_logic3_or0 & s_dadda_cla12_u_cla22_pg_logic1_or0;
  assign s_dadda_cla12_u_cla22_and6 = s_dadda_cla12_u_cla22_pg_logic0_and0 & s_dadda_cla12_u_cla22_pg_logic2_or0;
  assign s_dadda_cla12_u_cla22_and7 = s_dadda_cla12_u_cla22_pg_logic3_or0 & s_dadda_cla12_u_cla22_pg_logic1_or0;
  assign s_dadda_cla12_u_cla22_and8 = s_dadda_cla12_u_cla22_and6 & s_dadda_cla12_u_cla22_and7;
  assign s_dadda_cla12_u_cla22_and9 = s_dadda_cla12_u_cla22_pg_logic1_and0 & s_dadda_cla12_u_cla22_pg_logic3_or0;
  assign s_dadda_cla12_u_cla22_and10 = s_dadda_cla12_u_cla22_and9 & s_dadda_cla12_u_cla22_pg_logic2_or0;
  assign s_dadda_cla12_u_cla22_and11 = s_dadda_cla12_u_cla22_pg_logic2_and0 & s_dadda_cla12_u_cla22_pg_logic3_or0;
  assign s_dadda_cla12_u_cla22_or3 = s_dadda_cla12_u_cla22_and8 | s_dadda_cla12_u_cla22_and11;
  assign s_dadda_cla12_u_cla22_or4 = s_dadda_cla12_u_cla22_and10 | s_dadda_cla12_u_cla22_or3;
  assign s_dadda_cla12_u_cla22_or5 = s_dadda_cla12_u_cla22_pg_logic3_and0 | s_dadda_cla12_u_cla22_or4;
  assign s_dadda_cla12_u_cla22_pg_logic4_or0 = s_dadda_cla12_fa65_xor1 | s_dadda_cla12_fa83_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic4_and0 = s_dadda_cla12_fa65_xor1 & s_dadda_cla12_fa83_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic4_xor0 = s_dadda_cla12_fa65_xor1 ^ s_dadda_cla12_fa83_xor1;
  assign s_dadda_cla12_u_cla22_xor4 = s_dadda_cla12_u_cla22_pg_logic4_xor0 ^ s_dadda_cla12_u_cla22_or5;
  assign s_dadda_cla12_u_cla22_and12 = s_dadda_cla12_u_cla22_or5 & s_dadda_cla12_u_cla22_pg_logic4_or0;
  assign s_dadda_cla12_u_cla22_or6 = s_dadda_cla12_u_cla22_pg_logic4_and0 | s_dadda_cla12_u_cla22_and12;
  assign s_dadda_cla12_u_cla22_pg_logic5_or0 = s_dadda_cla12_fa66_xor1 | s_dadda_cla12_fa84_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic5_and0 = s_dadda_cla12_fa66_xor1 & s_dadda_cla12_fa84_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic5_xor0 = s_dadda_cla12_fa66_xor1 ^ s_dadda_cla12_fa84_xor1;
  assign s_dadda_cla12_u_cla22_xor5 = s_dadda_cla12_u_cla22_pg_logic5_xor0 ^ s_dadda_cla12_u_cla22_or6;
  assign s_dadda_cla12_u_cla22_and13 = s_dadda_cla12_u_cla22_or5 & s_dadda_cla12_u_cla22_pg_logic5_or0;
  assign s_dadda_cla12_u_cla22_and14 = s_dadda_cla12_u_cla22_and13 & s_dadda_cla12_u_cla22_pg_logic4_or0;
  assign s_dadda_cla12_u_cla22_and15 = s_dadda_cla12_u_cla22_pg_logic4_and0 & s_dadda_cla12_u_cla22_pg_logic5_or0;
  assign s_dadda_cla12_u_cla22_or7 = s_dadda_cla12_u_cla22_and14 | s_dadda_cla12_u_cla22_and15;
  assign s_dadda_cla12_u_cla22_or8 = s_dadda_cla12_u_cla22_pg_logic5_and0 | s_dadda_cla12_u_cla22_or7;
  assign s_dadda_cla12_u_cla22_pg_logic6_or0 = s_dadda_cla12_fa67_xor1 | s_dadda_cla12_fa85_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic6_and0 = s_dadda_cla12_fa67_xor1 & s_dadda_cla12_fa85_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic6_xor0 = s_dadda_cla12_fa67_xor1 ^ s_dadda_cla12_fa85_xor1;
  assign s_dadda_cla12_u_cla22_xor6 = s_dadda_cla12_u_cla22_pg_logic6_xor0 ^ s_dadda_cla12_u_cla22_or8;
  assign s_dadda_cla12_u_cla22_and16 = s_dadda_cla12_u_cla22_or5 & s_dadda_cla12_u_cla22_pg_logic5_or0;
  assign s_dadda_cla12_u_cla22_and17 = s_dadda_cla12_u_cla22_pg_logic6_or0 & s_dadda_cla12_u_cla22_pg_logic4_or0;
  assign s_dadda_cla12_u_cla22_and18 = s_dadda_cla12_u_cla22_and16 & s_dadda_cla12_u_cla22_and17;
  assign s_dadda_cla12_u_cla22_and19 = s_dadda_cla12_u_cla22_pg_logic4_and0 & s_dadda_cla12_u_cla22_pg_logic6_or0;
  assign s_dadda_cla12_u_cla22_and20 = s_dadda_cla12_u_cla22_and19 & s_dadda_cla12_u_cla22_pg_logic5_or0;
  assign s_dadda_cla12_u_cla22_and21 = s_dadda_cla12_u_cla22_pg_logic5_and0 & s_dadda_cla12_u_cla22_pg_logic6_or0;
  assign s_dadda_cla12_u_cla22_or9 = s_dadda_cla12_u_cla22_and18 | s_dadda_cla12_u_cla22_and20;
  assign s_dadda_cla12_u_cla22_or10 = s_dadda_cla12_u_cla22_or9 | s_dadda_cla12_u_cla22_and21;
  assign s_dadda_cla12_u_cla22_or11 = s_dadda_cla12_u_cla22_pg_logic6_and0 | s_dadda_cla12_u_cla22_or10;
  assign s_dadda_cla12_u_cla22_pg_logic7_or0 = s_dadda_cla12_fa68_xor1 | s_dadda_cla12_fa86_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic7_and0 = s_dadda_cla12_fa68_xor1 & s_dadda_cla12_fa86_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic7_xor0 = s_dadda_cla12_fa68_xor1 ^ s_dadda_cla12_fa86_xor1;
  assign s_dadda_cla12_u_cla22_xor7 = s_dadda_cla12_u_cla22_pg_logic7_xor0 ^ s_dadda_cla12_u_cla22_or11;
  assign s_dadda_cla12_u_cla22_and22 = s_dadda_cla12_u_cla22_or5 & s_dadda_cla12_u_cla22_pg_logic6_or0;
  assign s_dadda_cla12_u_cla22_and23 = s_dadda_cla12_u_cla22_pg_logic7_or0 & s_dadda_cla12_u_cla22_pg_logic5_or0;
  assign s_dadda_cla12_u_cla22_and24 = s_dadda_cla12_u_cla22_and22 & s_dadda_cla12_u_cla22_and23;
  assign s_dadda_cla12_u_cla22_and25 = s_dadda_cla12_u_cla22_and24 & s_dadda_cla12_u_cla22_pg_logic4_or0;
  assign s_dadda_cla12_u_cla22_and26 = s_dadda_cla12_u_cla22_pg_logic4_and0 & s_dadda_cla12_u_cla22_pg_logic6_or0;
  assign s_dadda_cla12_u_cla22_and27 = s_dadda_cla12_u_cla22_pg_logic7_or0 & s_dadda_cla12_u_cla22_pg_logic5_or0;
  assign s_dadda_cla12_u_cla22_and28 = s_dadda_cla12_u_cla22_and26 & s_dadda_cla12_u_cla22_and27;
  assign s_dadda_cla12_u_cla22_and29 = s_dadda_cla12_u_cla22_pg_logic5_and0 & s_dadda_cla12_u_cla22_pg_logic7_or0;
  assign s_dadda_cla12_u_cla22_and30 = s_dadda_cla12_u_cla22_and29 & s_dadda_cla12_u_cla22_pg_logic6_or0;
  assign s_dadda_cla12_u_cla22_and31 = s_dadda_cla12_u_cla22_pg_logic6_and0 & s_dadda_cla12_u_cla22_pg_logic7_or0;
  assign s_dadda_cla12_u_cla22_or12 = s_dadda_cla12_u_cla22_and25 | s_dadda_cla12_u_cla22_and30;
  assign s_dadda_cla12_u_cla22_or13 = s_dadda_cla12_u_cla22_and28 | s_dadda_cla12_u_cla22_and31;
  assign s_dadda_cla12_u_cla22_or14 = s_dadda_cla12_u_cla22_or12 | s_dadda_cla12_u_cla22_or13;
  assign s_dadda_cla12_u_cla22_or15 = s_dadda_cla12_u_cla22_pg_logic7_and0 | s_dadda_cla12_u_cla22_or14;
  assign s_dadda_cla12_u_cla22_pg_logic8_or0 = s_dadda_cla12_fa69_xor1 | s_dadda_cla12_fa87_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic8_and0 = s_dadda_cla12_fa69_xor1 & s_dadda_cla12_fa87_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic8_xor0 = s_dadda_cla12_fa69_xor1 ^ s_dadda_cla12_fa87_xor1;
  assign s_dadda_cla12_u_cla22_xor8 = s_dadda_cla12_u_cla22_pg_logic8_xor0 ^ s_dadda_cla12_u_cla22_or15;
  assign s_dadda_cla12_u_cla22_and32 = s_dadda_cla12_u_cla22_or15 & s_dadda_cla12_u_cla22_pg_logic8_or0;
  assign s_dadda_cla12_u_cla22_or16 = s_dadda_cla12_u_cla22_pg_logic8_and0 | s_dadda_cla12_u_cla22_and32;
  assign s_dadda_cla12_u_cla22_pg_logic9_or0 = s_dadda_cla12_fa70_xor1 | s_dadda_cla12_fa88_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic9_and0 = s_dadda_cla12_fa70_xor1 & s_dadda_cla12_fa88_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic9_xor0 = s_dadda_cla12_fa70_xor1 ^ s_dadda_cla12_fa88_xor1;
  assign s_dadda_cla12_u_cla22_xor9 = s_dadda_cla12_u_cla22_pg_logic9_xor0 ^ s_dadda_cla12_u_cla22_or16;
  assign s_dadda_cla12_u_cla22_and33 = s_dadda_cla12_u_cla22_or15 & s_dadda_cla12_u_cla22_pg_logic9_or0;
  assign s_dadda_cla12_u_cla22_and34 = s_dadda_cla12_u_cla22_and33 & s_dadda_cla12_u_cla22_pg_logic8_or0;
  assign s_dadda_cla12_u_cla22_and35 = s_dadda_cla12_u_cla22_pg_logic8_and0 & s_dadda_cla12_u_cla22_pg_logic9_or0;
  assign s_dadda_cla12_u_cla22_or17 = s_dadda_cla12_u_cla22_and34 | s_dadda_cla12_u_cla22_and35;
  assign s_dadda_cla12_u_cla22_or18 = s_dadda_cla12_u_cla22_pg_logic9_and0 | s_dadda_cla12_u_cla22_or17;
  assign s_dadda_cla12_u_cla22_pg_logic10_or0 = s_dadda_cla12_fa71_xor1 | s_dadda_cla12_fa89_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic10_and0 = s_dadda_cla12_fa71_xor1 & s_dadda_cla12_fa89_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic10_xor0 = s_dadda_cla12_fa71_xor1 ^ s_dadda_cla12_fa89_xor1;
  assign s_dadda_cla12_u_cla22_xor10 = s_dadda_cla12_u_cla22_pg_logic10_xor0 ^ s_dadda_cla12_u_cla22_or18;
  assign s_dadda_cla12_u_cla22_and36 = s_dadda_cla12_u_cla22_or15 & s_dadda_cla12_u_cla22_pg_logic9_or0;
  assign s_dadda_cla12_u_cla22_and37 = s_dadda_cla12_u_cla22_pg_logic10_or0 & s_dadda_cla12_u_cla22_pg_logic8_or0;
  assign s_dadda_cla12_u_cla22_and38 = s_dadda_cla12_u_cla22_and36 & s_dadda_cla12_u_cla22_and37;
  assign s_dadda_cla12_u_cla22_and39 = s_dadda_cla12_u_cla22_pg_logic8_and0 & s_dadda_cla12_u_cla22_pg_logic10_or0;
  assign s_dadda_cla12_u_cla22_and40 = s_dadda_cla12_u_cla22_and39 & s_dadda_cla12_u_cla22_pg_logic9_or0;
  assign s_dadda_cla12_u_cla22_and41 = s_dadda_cla12_u_cla22_pg_logic9_and0 & s_dadda_cla12_u_cla22_pg_logic10_or0;
  assign s_dadda_cla12_u_cla22_or19 = s_dadda_cla12_u_cla22_and38 | s_dadda_cla12_u_cla22_and40;
  assign s_dadda_cla12_u_cla22_or20 = s_dadda_cla12_u_cla22_or19 | s_dadda_cla12_u_cla22_and41;
  assign s_dadda_cla12_u_cla22_or21 = s_dadda_cla12_u_cla22_pg_logic10_and0 | s_dadda_cla12_u_cla22_or20;
  assign s_dadda_cla12_u_cla22_pg_logic11_or0 = s_dadda_cla12_fa72_xor1 | s_dadda_cla12_fa90_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic11_and0 = s_dadda_cla12_fa72_xor1 & s_dadda_cla12_fa90_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic11_xor0 = s_dadda_cla12_fa72_xor1 ^ s_dadda_cla12_fa90_xor1;
  assign s_dadda_cla12_u_cla22_xor11 = s_dadda_cla12_u_cla22_pg_logic11_xor0 ^ s_dadda_cla12_u_cla22_or21;
  assign s_dadda_cla12_u_cla22_and42 = s_dadda_cla12_u_cla22_or15 & s_dadda_cla12_u_cla22_pg_logic10_or0;
  assign s_dadda_cla12_u_cla22_and43 = s_dadda_cla12_u_cla22_pg_logic11_or0 & s_dadda_cla12_u_cla22_pg_logic9_or0;
  assign s_dadda_cla12_u_cla22_and44 = s_dadda_cla12_u_cla22_and42 & s_dadda_cla12_u_cla22_and43;
  assign s_dadda_cla12_u_cla22_and45 = s_dadda_cla12_u_cla22_and44 & s_dadda_cla12_u_cla22_pg_logic8_or0;
  assign s_dadda_cla12_u_cla22_and46 = s_dadda_cla12_u_cla22_pg_logic8_and0 & s_dadda_cla12_u_cla22_pg_logic10_or0;
  assign s_dadda_cla12_u_cla22_and47 = s_dadda_cla12_u_cla22_pg_logic11_or0 & s_dadda_cla12_u_cla22_pg_logic9_or0;
  assign s_dadda_cla12_u_cla22_and48 = s_dadda_cla12_u_cla22_and46 & s_dadda_cla12_u_cla22_and47;
  assign s_dadda_cla12_u_cla22_and49 = s_dadda_cla12_u_cla22_pg_logic9_and0 & s_dadda_cla12_u_cla22_pg_logic11_or0;
  assign s_dadda_cla12_u_cla22_and50 = s_dadda_cla12_u_cla22_and49 & s_dadda_cla12_u_cla22_pg_logic10_or0;
  assign s_dadda_cla12_u_cla22_and51 = s_dadda_cla12_u_cla22_pg_logic10_and0 & s_dadda_cla12_u_cla22_pg_logic11_or0;
  assign s_dadda_cla12_u_cla22_or22 = s_dadda_cla12_u_cla22_and45 | s_dadda_cla12_u_cla22_and50;
  assign s_dadda_cla12_u_cla22_or23 = s_dadda_cla12_u_cla22_and48 | s_dadda_cla12_u_cla22_and51;
  assign s_dadda_cla12_u_cla22_or24 = s_dadda_cla12_u_cla22_or22 | s_dadda_cla12_u_cla22_or23;
  assign s_dadda_cla12_u_cla22_or25 = s_dadda_cla12_u_cla22_pg_logic11_and0 | s_dadda_cla12_u_cla22_or24;
  assign s_dadda_cla12_u_cla22_pg_logic12_or0 = s_dadda_cla12_fa73_xor1 | s_dadda_cla12_fa91_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic12_and0 = s_dadda_cla12_fa73_xor1 & s_dadda_cla12_fa91_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic12_xor0 = s_dadda_cla12_fa73_xor1 ^ s_dadda_cla12_fa91_xor1;
  assign s_dadda_cla12_u_cla22_xor12 = s_dadda_cla12_u_cla22_pg_logic12_xor0 ^ s_dadda_cla12_u_cla22_or25;
  assign s_dadda_cla12_u_cla22_and52 = s_dadda_cla12_u_cla22_or25 & s_dadda_cla12_u_cla22_pg_logic12_or0;
  assign s_dadda_cla12_u_cla22_or26 = s_dadda_cla12_u_cla22_pg_logic12_and0 | s_dadda_cla12_u_cla22_and52;
  assign s_dadda_cla12_u_cla22_pg_logic13_or0 = s_dadda_cla12_fa74_xor1 | s_dadda_cla12_fa92_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic13_and0 = s_dadda_cla12_fa74_xor1 & s_dadda_cla12_fa92_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic13_xor0 = s_dadda_cla12_fa74_xor1 ^ s_dadda_cla12_fa92_xor1;
  assign s_dadda_cla12_u_cla22_xor13 = s_dadda_cla12_u_cla22_pg_logic13_xor0 ^ s_dadda_cla12_u_cla22_or26;
  assign s_dadda_cla12_u_cla22_and53 = s_dadda_cla12_u_cla22_or25 & s_dadda_cla12_u_cla22_pg_logic13_or0;
  assign s_dadda_cla12_u_cla22_and54 = s_dadda_cla12_u_cla22_and53 & s_dadda_cla12_u_cla22_pg_logic12_or0;
  assign s_dadda_cla12_u_cla22_and55 = s_dadda_cla12_u_cla22_pg_logic12_and0 & s_dadda_cla12_u_cla22_pg_logic13_or0;
  assign s_dadda_cla12_u_cla22_or27 = s_dadda_cla12_u_cla22_and54 | s_dadda_cla12_u_cla22_and55;
  assign s_dadda_cla12_u_cla22_or28 = s_dadda_cla12_u_cla22_pg_logic13_and0 | s_dadda_cla12_u_cla22_or27;
  assign s_dadda_cla12_u_cla22_pg_logic14_or0 = s_dadda_cla12_fa75_xor1 | s_dadda_cla12_fa93_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic14_and0 = s_dadda_cla12_fa75_xor1 & s_dadda_cla12_fa93_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic14_xor0 = s_dadda_cla12_fa75_xor1 ^ s_dadda_cla12_fa93_xor1;
  assign s_dadda_cla12_u_cla22_xor14 = s_dadda_cla12_u_cla22_pg_logic14_xor0 ^ s_dadda_cla12_u_cla22_or28;
  assign s_dadda_cla12_u_cla22_and56 = s_dadda_cla12_u_cla22_or25 & s_dadda_cla12_u_cla22_pg_logic13_or0;
  assign s_dadda_cla12_u_cla22_and57 = s_dadda_cla12_u_cla22_pg_logic14_or0 & s_dadda_cla12_u_cla22_pg_logic12_or0;
  assign s_dadda_cla12_u_cla22_and58 = s_dadda_cla12_u_cla22_and56 & s_dadda_cla12_u_cla22_and57;
  assign s_dadda_cla12_u_cla22_and59 = s_dadda_cla12_u_cla22_pg_logic12_and0 & s_dadda_cla12_u_cla22_pg_logic14_or0;
  assign s_dadda_cla12_u_cla22_and60 = s_dadda_cla12_u_cla22_and59 & s_dadda_cla12_u_cla22_pg_logic13_or0;
  assign s_dadda_cla12_u_cla22_and61 = s_dadda_cla12_u_cla22_pg_logic13_and0 & s_dadda_cla12_u_cla22_pg_logic14_or0;
  assign s_dadda_cla12_u_cla22_or29 = s_dadda_cla12_u_cla22_and58 | s_dadda_cla12_u_cla22_and60;
  assign s_dadda_cla12_u_cla22_or30 = s_dadda_cla12_u_cla22_or29 | s_dadda_cla12_u_cla22_and61;
  assign s_dadda_cla12_u_cla22_or31 = s_dadda_cla12_u_cla22_pg_logic14_and0 | s_dadda_cla12_u_cla22_or30;
  assign s_dadda_cla12_u_cla22_pg_logic15_or0 = s_dadda_cla12_fa76_xor1 | s_dadda_cla12_fa94_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic15_and0 = s_dadda_cla12_fa76_xor1 & s_dadda_cla12_fa94_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic15_xor0 = s_dadda_cla12_fa76_xor1 ^ s_dadda_cla12_fa94_xor1;
  assign s_dadda_cla12_u_cla22_xor15 = s_dadda_cla12_u_cla22_pg_logic15_xor0 ^ s_dadda_cla12_u_cla22_or31;
  assign s_dadda_cla12_u_cla22_and62 = s_dadda_cla12_u_cla22_or25 & s_dadda_cla12_u_cla22_pg_logic14_or0;
  assign s_dadda_cla12_u_cla22_and63 = s_dadda_cla12_u_cla22_pg_logic15_or0 & s_dadda_cla12_u_cla22_pg_logic13_or0;
  assign s_dadda_cla12_u_cla22_and64 = s_dadda_cla12_u_cla22_and62 & s_dadda_cla12_u_cla22_and63;
  assign s_dadda_cla12_u_cla22_and65 = s_dadda_cla12_u_cla22_and64 & s_dadda_cla12_u_cla22_pg_logic12_or0;
  assign s_dadda_cla12_u_cla22_and66 = s_dadda_cla12_u_cla22_pg_logic12_and0 & s_dadda_cla12_u_cla22_pg_logic14_or0;
  assign s_dadda_cla12_u_cla22_and67 = s_dadda_cla12_u_cla22_pg_logic15_or0 & s_dadda_cla12_u_cla22_pg_logic13_or0;
  assign s_dadda_cla12_u_cla22_and68 = s_dadda_cla12_u_cla22_and66 & s_dadda_cla12_u_cla22_and67;
  assign s_dadda_cla12_u_cla22_and69 = s_dadda_cla12_u_cla22_pg_logic13_and0 & s_dadda_cla12_u_cla22_pg_logic15_or0;
  assign s_dadda_cla12_u_cla22_and70 = s_dadda_cla12_u_cla22_and69 & s_dadda_cla12_u_cla22_pg_logic14_or0;
  assign s_dadda_cla12_u_cla22_and71 = s_dadda_cla12_u_cla22_pg_logic14_and0 & s_dadda_cla12_u_cla22_pg_logic15_or0;
  assign s_dadda_cla12_u_cla22_or32 = s_dadda_cla12_u_cla22_and65 | s_dadda_cla12_u_cla22_and70;
  assign s_dadda_cla12_u_cla22_or33 = s_dadda_cla12_u_cla22_and68 | s_dadda_cla12_u_cla22_and71;
  assign s_dadda_cla12_u_cla22_or34 = s_dadda_cla12_u_cla22_or32 | s_dadda_cla12_u_cla22_or33;
  assign s_dadda_cla12_u_cla22_or35 = s_dadda_cla12_u_cla22_pg_logic15_and0 | s_dadda_cla12_u_cla22_or34;
  assign s_dadda_cla12_u_cla22_pg_logic16_or0 = s_dadda_cla12_fa77_xor1 | s_dadda_cla12_fa95_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic16_and0 = s_dadda_cla12_fa77_xor1 & s_dadda_cla12_fa95_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic16_xor0 = s_dadda_cla12_fa77_xor1 ^ s_dadda_cla12_fa95_xor1;
  assign s_dadda_cla12_u_cla22_xor16 = s_dadda_cla12_u_cla22_pg_logic16_xor0 ^ s_dadda_cla12_u_cla22_or35;
  assign s_dadda_cla12_u_cla22_and72 = s_dadda_cla12_u_cla22_or35 & s_dadda_cla12_u_cla22_pg_logic16_or0;
  assign s_dadda_cla12_u_cla22_or36 = s_dadda_cla12_u_cla22_pg_logic16_and0 | s_dadda_cla12_u_cla22_and72;
  assign s_dadda_cla12_u_cla22_pg_logic17_or0 = s_dadda_cla12_fa78_xor1 | s_dadda_cla12_fa96_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic17_and0 = s_dadda_cla12_fa78_xor1 & s_dadda_cla12_fa96_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic17_xor0 = s_dadda_cla12_fa78_xor1 ^ s_dadda_cla12_fa96_xor1;
  assign s_dadda_cla12_u_cla22_xor17 = s_dadda_cla12_u_cla22_pg_logic17_xor0 ^ s_dadda_cla12_u_cla22_or36;
  assign s_dadda_cla12_u_cla22_and73 = s_dadda_cla12_u_cla22_or35 & s_dadda_cla12_u_cla22_pg_logic17_or0;
  assign s_dadda_cla12_u_cla22_and74 = s_dadda_cla12_u_cla22_and73 & s_dadda_cla12_u_cla22_pg_logic16_or0;
  assign s_dadda_cla12_u_cla22_and75 = s_dadda_cla12_u_cla22_pg_logic16_and0 & s_dadda_cla12_u_cla22_pg_logic17_or0;
  assign s_dadda_cla12_u_cla22_or37 = s_dadda_cla12_u_cla22_and74 | s_dadda_cla12_u_cla22_and75;
  assign s_dadda_cla12_u_cla22_or38 = s_dadda_cla12_u_cla22_pg_logic17_and0 | s_dadda_cla12_u_cla22_or37;
  assign s_dadda_cla12_u_cla22_pg_logic18_or0 = s_dadda_cla12_fa79_xor1 | s_dadda_cla12_fa97_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic18_and0 = s_dadda_cla12_fa79_xor1 & s_dadda_cla12_fa97_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic18_xor0 = s_dadda_cla12_fa79_xor1 ^ s_dadda_cla12_fa97_xor1;
  assign s_dadda_cla12_u_cla22_xor18 = s_dadda_cla12_u_cla22_pg_logic18_xor0 ^ s_dadda_cla12_u_cla22_or38;
  assign s_dadda_cla12_u_cla22_and76 = s_dadda_cla12_u_cla22_or35 & s_dadda_cla12_u_cla22_pg_logic17_or0;
  assign s_dadda_cla12_u_cla22_and77 = s_dadda_cla12_u_cla22_pg_logic18_or0 & s_dadda_cla12_u_cla22_pg_logic16_or0;
  assign s_dadda_cla12_u_cla22_and78 = s_dadda_cla12_u_cla22_and76 & s_dadda_cla12_u_cla22_and77;
  assign s_dadda_cla12_u_cla22_and79 = s_dadda_cla12_u_cla22_pg_logic16_and0 & s_dadda_cla12_u_cla22_pg_logic18_or0;
  assign s_dadda_cla12_u_cla22_and80 = s_dadda_cla12_u_cla22_and79 & s_dadda_cla12_u_cla22_pg_logic17_or0;
  assign s_dadda_cla12_u_cla22_and81 = s_dadda_cla12_u_cla22_pg_logic17_and0 & s_dadda_cla12_u_cla22_pg_logic18_or0;
  assign s_dadda_cla12_u_cla22_or39 = s_dadda_cla12_u_cla22_and78 | s_dadda_cla12_u_cla22_and80;
  assign s_dadda_cla12_u_cla22_or40 = s_dadda_cla12_u_cla22_or39 | s_dadda_cla12_u_cla22_and81;
  assign s_dadda_cla12_u_cla22_or41 = s_dadda_cla12_u_cla22_pg_logic18_and0 | s_dadda_cla12_u_cla22_or40;
  assign s_dadda_cla12_u_cla22_pg_logic19_or0 = s_dadda_cla12_fa80_xor1 | s_dadda_cla12_fa98_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic19_and0 = s_dadda_cla12_fa80_xor1 & s_dadda_cla12_fa98_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic19_xor0 = s_dadda_cla12_fa80_xor1 ^ s_dadda_cla12_fa98_xor1;
  assign s_dadda_cla12_u_cla22_xor19 = s_dadda_cla12_u_cla22_pg_logic19_xor0 ^ s_dadda_cla12_u_cla22_or41;
  assign s_dadda_cla12_u_cla22_and82 = s_dadda_cla12_u_cla22_or35 & s_dadda_cla12_u_cla22_pg_logic18_or0;
  assign s_dadda_cla12_u_cla22_and83 = s_dadda_cla12_u_cla22_pg_logic19_or0 & s_dadda_cla12_u_cla22_pg_logic17_or0;
  assign s_dadda_cla12_u_cla22_and84 = s_dadda_cla12_u_cla22_and82 & s_dadda_cla12_u_cla22_and83;
  assign s_dadda_cla12_u_cla22_and85 = s_dadda_cla12_u_cla22_and84 & s_dadda_cla12_u_cla22_pg_logic16_or0;
  assign s_dadda_cla12_u_cla22_and86 = s_dadda_cla12_u_cla22_pg_logic16_and0 & s_dadda_cla12_u_cla22_pg_logic18_or0;
  assign s_dadda_cla12_u_cla22_and87 = s_dadda_cla12_u_cla22_pg_logic19_or0 & s_dadda_cla12_u_cla22_pg_logic17_or0;
  assign s_dadda_cla12_u_cla22_and88 = s_dadda_cla12_u_cla22_and86 & s_dadda_cla12_u_cla22_and87;
  assign s_dadda_cla12_u_cla22_and89 = s_dadda_cla12_u_cla22_pg_logic17_and0 & s_dadda_cla12_u_cla22_pg_logic19_or0;
  assign s_dadda_cla12_u_cla22_and90 = s_dadda_cla12_u_cla22_and89 & s_dadda_cla12_u_cla22_pg_logic18_or0;
  assign s_dadda_cla12_u_cla22_and91 = s_dadda_cla12_u_cla22_pg_logic18_and0 & s_dadda_cla12_u_cla22_pg_logic19_or0;
  assign s_dadda_cla12_u_cla22_or42 = s_dadda_cla12_u_cla22_and85 | s_dadda_cla12_u_cla22_and90;
  assign s_dadda_cla12_u_cla22_or43 = s_dadda_cla12_u_cla22_and88 | s_dadda_cla12_u_cla22_and91;
  assign s_dadda_cla12_u_cla22_or44 = s_dadda_cla12_u_cla22_or42 | s_dadda_cla12_u_cla22_or43;
  assign s_dadda_cla12_u_cla22_or45 = s_dadda_cla12_u_cla22_pg_logic19_and0 | s_dadda_cla12_u_cla22_or44;
  assign s_dadda_cla12_u_cla22_pg_logic20_or0 = s_dadda_cla12_nand_10_11 | s_dadda_cla12_fa99_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic20_and0 = s_dadda_cla12_nand_10_11 & s_dadda_cla12_fa99_xor1;
  assign s_dadda_cla12_u_cla22_pg_logic20_xor0 = s_dadda_cla12_nand_10_11 ^ s_dadda_cla12_fa99_xor1;
  assign s_dadda_cla12_u_cla22_xor20 = s_dadda_cla12_u_cla22_pg_logic20_xor0 ^ s_dadda_cla12_u_cla22_or45;
  assign s_dadda_cla12_u_cla22_and92 = s_dadda_cla12_u_cla22_or45 & s_dadda_cla12_u_cla22_pg_logic20_or0;
  assign s_dadda_cla12_u_cla22_or46 = s_dadda_cla12_u_cla22_pg_logic20_and0 | s_dadda_cla12_u_cla22_and92;
  assign s_dadda_cla12_u_cla22_pg_logic21_or0 = s_dadda_cla12_fa99_or0 | s_dadda_cla12_and_11_11;
  assign s_dadda_cla12_u_cla22_pg_logic21_and0 = s_dadda_cla12_fa99_or0 & s_dadda_cla12_and_11_11;
  assign s_dadda_cla12_u_cla22_pg_logic21_xor0 = s_dadda_cla12_fa99_or0 ^ s_dadda_cla12_and_11_11;
  assign s_dadda_cla12_u_cla22_xor21 = s_dadda_cla12_u_cla22_pg_logic21_xor0 ^ s_dadda_cla12_u_cla22_or46;
  assign s_dadda_cla12_u_cla22_and93 = s_dadda_cla12_u_cla22_or45 & s_dadda_cla12_u_cla22_pg_logic21_or0;
  assign s_dadda_cla12_u_cla22_and94 = s_dadda_cla12_u_cla22_and93 & s_dadda_cla12_u_cla22_pg_logic20_or0;
  assign s_dadda_cla12_u_cla22_and95 = s_dadda_cla12_u_cla22_pg_logic20_and0 & s_dadda_cla12_u_cla22_pg_logic21_or0;
  assign s_dadda_cla12_u_cla22_or47 = s_dadda_cla12_u_cla22_and94 | s_dadda_cla12_u_cla22_and95;
  assign s_dadda_cla12_u_cla22_or48 = s_dadda_cla12_u_cla22_pg_logic21_and0 | s_dadda_cla12_u_cla22_or47;
  assign s_dadda_cla12_xor0 = ~s_dadda_cla12_u_cla22_or48;

  assign s_dadda_cla12_out[0] = s_dadda_cla12_and_0_0;
  assign s_dadda_cla12_out[1] = s_dadda_cla12_u_cla22_pg_logic0_xor0;
  assign s_dadda_cla12_out[2] = s_dadda_cla12_u_cla22_xor1;
  assign s_dadda_cla12_out[3] = s_dadda_cla12_u_cla22_xor2;
  assign s_dadda_cla12_out[4] = s_dadda_cla12_u_cla22_xor3;
  assign s_dadda_cla12_out[5] = s_dadda_cla12_u_cla22_xor4;
  assign s_dadda_cla12_out[6] = s_dadda_cla12_u_cla22_xor5;
  assign s_dadda_cla12_out[7] = s_dadda_cla12_u_cla22_xor6;
  assign s_dadda_cla12_out[8] = s_dadda_cla12_u_cla22_xor7;
  assign s_dadda_cla12_out[9] = s_dadda_cla12_u_cla22_xor8;
  assign s_dadda_cla12_out[10] = s_dadda_cla12_u_cla22_xor9;
  assign s_dadda_cla12_out[11] = s_dadda_cla12_u_cla22_xor10;
  assign s_dadda_cla12_out[12] = s_dadda_cla12_u_cla22_xor11;
  assign s_dadda_cla12_out[13] = s_dadda_cla12_u_cla22_xor12;
  assign s_dadda_cla12_out[14] = s_dadda_cla12_u_cla22_xor13;
  assign s_dadda_cla12_out[15] = s_dadda_cla12_u_cla22_xor14;
  assign s_dadda_cla12_out[16] = s_dadda_cla12_u_cla22_xor15;
  assign s_dadda_cla12_out[17] = s_dadda_cla12_u_cla22_xor16;
  assign s_dadda_cla12_out[18] = s_dadda_cla12_u_cla22_xor17;
  assign s_dadda_cla12_out[19] = s_dadda_cla12_u_cla22_xor18;
  assign s_dadda_cla12_out[20] = s_dadda_cla12_u_cla22_xor19;
  assign s_dadda_cla12_out[21] = s_dadda_cla12_u_cla22_xor20;
  assign s_dadda_cla12_out[22] = s_dadda_cla12_u_cla22_xor21;
  assign s_dadda_cla12_out[23] = s_dadda_cla12_xor0;
endmodule