module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] pg_fa_xor0, output [0:0] pg_fa_and0, output [0:0] pg_fa_xor1);
  xor_gate xor_gate_pg_fa_xor0(.a(a[0]), .b(b[0]), .out(pg_fa_xor0));
  and_gate and_gate_pg_fa_and0(.a(a[0]), .b(b[0]), .out(pg_fa_and0));
  xor_gate xor_gate_pg_fa_xor1(.a(pg_fa_xor0[0]), .b(cin[0]), .out(pg_fa_xor1));
endmodule

module csa_component18(input [17:0] a, input [17:0] b, input [17:0] c, output [37:0] csa_component18_out);
  wire [0:0] csa_component18_fa0_xor1;
  wire [0:0] csa_component18_fa0_or0;
  wire [0:0] csa_component18_fa1_xor1;
  wire [0:0] csa_component18_fa1_or0;
  wire [0:0] csa_component18_fa2_xor1;
  wire [0:0] csa_component18_fa2_or0;
  wire [0:0] csa_component18_fa3_xor1;
  wire [0:0] csa_component18_fa3_or0;
  wire [0:0] csa_component18_fa4_xor1;
  wire [0:0] csa_component18_fa4_or0;
  wire [0:0] csa_component18_fa5_xor1;
  wire [0:0] csa_component18_fa5_or0;
  wire [0:0] csa_component18_fa6_xor1;
  wire [0:0] csa_component18_fa6_or0;
  wire [0:0] csa_component18_fa7_xor1;
  wire [0:0] csa_component18_fa7_or0;
  wire [0:0] csa_component18_fa8_xor1;
  wire [0:0] csa_component18_fa8_or0;
  wire [0:0] csa_component18_fa9_xor1;
  wire [0:0] csa_component18_fa9_or0;
  wire [0:0] csa_component18_fa10_xor1;
  wire [0:0] csa_component18_fa10_or0;
  wire [0:0] csa_component18_fa11_xor1;
  wire [0:0] csa_component18_fa11_or0;
  wire [0:0] csa_component18_fa12_xor1;
  wire [0:0] csa_component18_fa12_or0;
  wire [0:0] csa_component18_fa13_xor1;
  wire [0:0] csa_component18_fa13_or0;
  wire [0:0] csa_component18_fa14_xor1;
  wire [0:0] csa_component18_fa14_or0;
  wire [0:0] csa_component18_fa15_xor1;
  wire [0:0] csa_component18_fa15_or0;
  wire [0:0] csa_component18_fa16_xor1;
  wire [0:0] csa_component18_fa16_or0;
  wire [0:0] csa_component18_fa17_xor1;
  wire [0:0] csa_component18_fa17_or0;

  fa fa_csa_component18_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component18_fa0_xor1), .fa_or0(csa_component18_fa0_or0));
  fa fa_csa_component18_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component18_fa1_xor1), .fa_or0(csa_component18_fa1_or0));
  fa fa_csa_component18_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component18_fa2_xor1), .fa_or0(csa_component18_fa2_or0));
  fa fa_csa_component18_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component18_fa3_xor1), .fa_or0(csa_component18_fa3_or0));
  fa fa_csa_component18_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component18_fa4_xor1), .fa_or0(csa_component18_fa4_or0));
  fa fa_csa_component18_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component18_fa5_xor1), .fa_or0(csa_component18_fa5_or0));
  fa fa_csa_component18_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component18_fa6_xor1), .fa_or0(csa_component18_fa6_or0));
  fa fa_csa_component18_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component18_fa7_xor1), .fa_or0(csa_component18_fa7_or0));
  fa fa_csa_component18_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component18_fa8_xor1), .fa_or0(csa_component18_fa8_or0));
  fa fa_csa_component18_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component18_fa9_xor1), .fa_or0(csa_component18_fa9_or0));
  fa fa_csa_component18_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component18_fa10_xor1), .fa_or0(csa_component18_fa10_or0));
  fa fa_csa_component18_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component18_fa11_xor1), .fa_or0(csa_component18_fa11_or0));
  fa fa_csa_component18_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component18_fa12_xor1), .fa_or0(csa_component18_fa12_or0));
  fa fa_csa_component18_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component18_fa13_xor1), .fa_or0(csa_component18_fa13_or0));
  fa fa_csa_component18_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component18_fa14_xor1), .fa_or0(csa_component18_fa14_or0));
  fa fa_csa_component18_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component18_fa15_xor1), .fa_or0(csa_component18_fa15_or0));
  fa fa_csa_component18_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component18_fa16_xor1), .fa_or0(csa_component18_fa16_or0));
  fa fa_csa_component18_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component18_fa17_xor1), .fa_or0(csa_component18_fa17_or0));

  assign csa_component18_out[0] = csa_component18_fa0_xor1[0];
  assign csa_component18_out[1] = csa_component18_fa1_xor1[0];
  assign csa_component18_out[2] = csa_component18_fa2_xor1[0];
  assign csa_component18_out[3] = csa_component18_fa3_xor1[0];
  assign csa_component18_out[4] = csa_component18_fa4_xor1[0];
  assign csa_component18_out[5] = csa_component18_fa5_xor1[0];
  assign csa_component18_out[6] = csa_component18_fa6_xor1[0];
  assign csa_component18_out[7] = csa_component18_fa7_xor1[0];
  assign csa_component18_out[8] = csa_component18_fa8_xor1[0];
  assign csa_component18_out[9] = csa_component18_fa9_xor1[0];
  assign csa_component18_out[10] = csa_component18_fa10_xor1[0];
  assign csa_component18_out[11] = csa_component18_fa11_xor1[0];
  assign csa_component18_out[12] = csa_component18_fa12_xor1[0];
  assign csa_component18_out[13] = csa_component18_fa13_xor1[0];
  assign csa_component18_out[14] = csa_component18_fa14_xor1[0];
  assign csa_component18_out[15] = csa_component18_fa15_xor1[0];
  assign csa_component18_out[16] = csa_component18_fa16_xor1[0];
  assign csa_component18_out[17] = csa_component18_fa17_xor1[0];
  assign csa_component18_out[18] = 1'b0;
  assign csa_component18_out[19] = 1'b0;
  assign csa_component18_out[20] = csa_component18_fa0_or0[0];
  assign csa_component18_out[21] = csa_component18_fa1_or0[0];
  assign csa_component18_out[22] = csa_component18_fa2_or0[0];
  assign csa_component18_out[23] = csa_component18_fa3_or0[0];
  assign csa_component18_out[24] = csa_component18_fa4_or0[0];
  assign csa_component18_out[25] = csa_component18_fa5_or0[0];
  assign csa_component18_out[26] = csa_component18_fa6_or0[0];
  assign csa_component18_out[27] = csa_component18_fa7_or0[0];
  assign csa_component18_out[28] = csa_component18_fa8_or0[0];
  assign csa_component18_out[29] = csa_component18_fa9_or0[0];
  assign csa_component18_out[30] = csa_component18_fa10_or0[0];
  assign csa_component18_out[31] = csa_component18_fa11_or0[0];
  assign csa_component18_out[32] = csa_component18_fa12_or0[0];
  assign csa_component18_out[33] = csa_component18_fa13_or0[0];
  assign csa_component18_out[34] = csa_component18_fa14_or0[0];
  assign csa_component18_out[35] = csa_component18_fa15_or0[0];
  assign csa_component18_out[36] = csa_component18_fa16_or0[0];
  assign csa_component18_out[37] = csa_component18_fa17_or0[0];
endmodule

module csa_component21(input [20:0] a, input [20:0] b, input [20:0] c, output [43:0] csa_component21_out);
  wire [0:0] csa_component21_fa0_xor1;
  wire [0:0] csa_component21_fa0_or0;
  wire [0:0] csa_component21_fa1_xor1;
  wire [0:0] csa_component21_fa1_or0;
  wire [0:0] csa_component21_fa2_xor1;
  wire [0:0] csa_component21_fa2_or0;
  wire [0:0] csa_component21_fa3_xor1;
  wire [0:0] csa_component21_fa3_or0;
  wire [0:0] csa_component21_fa4_xor1;
  wire [0:0] csa_component21_fa4_or0;
  wire [0:0] csa_component21_fa5_xor1;
  wire [0:0] csa_component21_fa5_or0;
  wire [0:0] csa_component21_fa6_xor1;
  wire [0:0] csa_component21_fa6_or0;
  wire [0:0] csa_component21_fa7_xor1;
  wire [0:0] csa_component21_fa7_or0;
  wire [0:0] csa_component21_fa8_xor1;
  wire [0:0] csa_component21_fa8_or0;
  wire [0:0] csa_component21_fa9_xor1;
  wire [0:0] csa_component21_fa9_or0;
  wire [0:0] csa_component21_fa10_xor1;
  wire [0:0] csa_component21_fa10_or0;
  wire [0:0] csa_component21_fa11_xor1;
  wire [0:0] csa_component21_fa11_or0;
  wire [0:0] csa_component21_fa12_xor1;
  wire [0:0] csa_component21_fa12_or0;
  wire [0:0] csa_component21_fa13_xor1;
  wire [0:0] csa_component21_fa13_or0;
  wire [0:0] csa_component21_fa14_xor1;
  wire [0:0] csa_component21_fa14_or0;
  wire [0:0] csa_component21_fa15_xor1;
  wire [0:0] csa_component21_fa15_or0;
  wire [0:0] csa_component21_fa16_xor1;
  wire [0:0] csa_component21_fa16_or0;
  wire [0:0] csa_component21_fa17_xor1;
  wire [0:0] csa_component21_fa17_or0;
  wire [0:0] csa_component21_fa18_xor1;
  wire [0:0] csa_component21_fa18_or0;
  wire [0:0] csa_component21_fa19_xor1;
  wire [0:0] csa_component21_fa19_or0;
  wire [0:0] csa_component21_fa20_xor1;
  wire [0:0] csa_component21_fa20_or0;

  fa fa_csa_component21_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component21_fa0_xor1), .fa_or0(csa_component21_fa0_or0));
  fa fa_csa_component21_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component21_fa1_xor1), .fa_or0(csa_component21_fa1_or0));
  fa fa_csa_component21_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component21_fa2_xor1), .fa_or0(csa_component21_fa2_or0));
  fa fa_csa_component21_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component21_fa3_xor1), .fa_or0(csa_component21_fa3_or0));
  fa fa_csa_component21_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component21_fa4_xor1), .fa_or0(csa_component21_fa4_or0));
  fa fa_csa_component21_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component21_fa5_xor1), .fa_or0(csa_component21_fa5_or0));
  fa fa_csa_component21_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component21_fa6_xor1), .fa_or0(csa_component21_fa6_or0));
  fa fa_csa_component21_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component21_fa7_xor1), .fa_or0(csa_component21_fa7_or0));
  fa fa_csa_component21_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component21_fa8_xor1), .fa_or0(csa_component21_fa8_or0));
  fa fa_csa_component21_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component21_fa9_xor1), .fa_or0(csa_component21_fa9_or0));
  fa fa_csa_component21_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component21_fa10_xor1), .fa_or0(csa_component21_fa10_or0));
  fa fa_csa_component21_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component21_fa11_xor1), .fa_or0(csa_component21_fa11_or0));
  fa fa_csa_component21_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component21_fa12_xor1), .fa_or0(csa_component21_fa12_or0));
  fa fa_csa_component21_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component21_fa13_xor1), .fa_or0(csa_component21_fa13_or0));
  fa fa_csa_component21_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component21_fa14_xor1), .fa_or0(csa_component21_fa14_or0));
  fa fa_csa_component21_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component21_fa15_xor1), .fa_or0(csa_component21_fa15_or0));
  fa fa_csa_component21_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component21_fa16_xor1), .fa_or0(csa_component21_fa16_or0));
  fa fa_csa_component21_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component21_fa17_xor1), .fa_or0(csa_component21_fa17_or0));
  fa fa_csa_component21_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component21_fa18_xor1), .fa_or0(csa_component21_fa18_or0));
  fa fa_csa_component21_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component21_fa19_xor1), .fa_or0(csa_component21_fa19_or0));
  fa fa_csa_component21_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component21_fa20_xor1), .fa_or0(csa_component21_fa20_or0));

  assign csa_component21_out[0] = csa_component21_fa0_xor1[0];
  assign csa_component21_out[1] = csa_component21_fa1_xor1[0];
  assign csa_component21_out[2] = csa_component21_fa2_xor1[0];
  assign csa_component21_out[3] = csa_component21_fa3_xor1[0];
  assign csa_component21_out[4] = csa_component21_fa4_xor1[0];
  assign csa_component21_out[5] = csa_component21_fa5_xor1[0];
  assign csa_component21_out[6] = csa_component21_fa6_xor1[0];
  assign csa_component21_out[7] = csa_component21_fa7_xor1[0];
  assign csa_component21_out[8] = csa_component21_fa8_xor1[0];
  assign csa_component21_out[9] = csa_component21_fa9_xor1[0];
  assign csa_component21_out[10] = csa_component21_fa10_xor1[0];
  assign csa_component21_out[11] = csa_component21_fa11_xor1[0];
  assign csa_component21_out[12] = csa_component21_fa12_xor1[0];
  assign csa_component21_out[13] = csa_component21_fa13_xor1[0];
  assign csa_component21_out[14] = csa_component21_fa14_xor1[0];
  assign csa_component21_out[15] = csa_component21_fa15_xor1[0];
  assign csa_component21_out[16] = csa_component21_fa16_xor1[0];
  assign csa_component21_out[17] = csa_component21_fa17_xor1[0];
  assign csa_component21_out[18] = csa_component21_fa18_xor1[0];
  assign csa_component21_out[19] = csa_component21_fa19_xor1[0];
  assign csa_component21_out[20] = csa_component21_fa20_xor1[0];
  assign csa_component21_out[21] = 1'b0;
  assign csa_component21_out[22] = 1'b0;
  assign csa_component21_out[23] = csa_component21_fa0_or0[0];
  assign csa_component21_out[24] = csa_component21_fa1_or0[0];
  assign csa_component21_out[25] = csa_component21_fa2_or0[0];
  assign csa_component21_out[26] = csa_component21_fa3_or0[0];
  assign csa_component21_out[27] = csa_component21_fa4_or0[0];
  assign csa_component21_out[28] = csa_component21_fa5_or0[0];
  assign csa_component21_out[29] = csa_component21_fa6_or0[0];
  assign csa_component21_out[30] = csa_component21_fa7_or0[0];
  assign csa_component21_out[31] = csa_component21_fa8_or0[0];
  assign csa_component21_out[32] = csa_component21_fa9_or0[0];
  assign csa_component21_out[33] = csa_component21_fa10_or0[0];
  assign csa_component21_out[34] = csa_component21_fa11_or0[0];
  assign csa_component21_out[35] = csa_component21_fa12_or0[0];
  assign csa_component21_out[36] = csa_component21_fa13_or0[0];
  assign csa_component21_out[37] = csa_component21_fa14_or0[0];
  assign csa_component21_out[38] = csa_component21_fa15_or0[0];
  assign csa_component21_out[39] = csa_component21_fa16_or0[0];
  assign csa_component21_out[40] = csa_component21_fa17_or0[0];
  assign csa_component21_out[41] = csa_component21_fa18_or0[0];
  assign csa_component21_out[42] = csa_component21_fa19_or0[0];
  assign csa_component21_out[43] = csa_component21_fa20_or0[0];
endmodule

module csa_component24(input [23:0] a, input [23:0] b, input [23:0] c, output [49:0] csa_component24_out);
  wire [0:0] csa_component24_fa0_xor1;
  wire [0:0] csa_component24_fa0_or0;
  wire [0:0] csa_component24_fa1_xor1;
  wire [0:0] csa_component24_fa1_or0;
  wire [0:0] csa_component24_fa2_xor1;
  wire [0:0] csa_component24_fa2_or0;
  wire [0:0] csa_component24_fa3_xor1;
  wire [0:0] csa_component24_fa3_or0;
  wire [0:0] csa_component24_fa4_xor1;
  wire [0:0] csa_component24_fa4_or0;
  wire [0:0] csa_component24_fa5_xor1;
  wire [0:0] csa_component24_fa5_or0;
  wire [0:0] csa_component24_fa6_xor1;
  wire [0:0] csa_component24_fa6_or0;
  wire [0:0] csa_component24_fa7_xor1;
  wire [0:0] csa_component24_fa7_or0;
  wire [0:0] csa_component24_fa8_xor1;
  wire [0:0] csa_component24_fa8_or0;
  wire [0:0] csa_component24_fa9_xor1;
  wire [0:0] csa_component24_fa9_or0;
  wire [0:0] csa_component24_fa10_xor1;
  wire [0:0] csa_component24_fa10_or0;
  wire [0:0] csa_component24_fa11_xor1;
  wire [0:0] csa_component24_fa11_or0;
  wire [0:0] csa_component24_fa12_xor1;
  wire [0:0] csa_component24_fa12_or0;
  wire [0:0] csa_component24_fa13_xor1;
  wire [0:0] csa_component24_fa13_or0;
  wire [0:0] csa_component24_fa14_xor1;
  wire [0:0] csa_component24_fa14_or0;
  wire [0:0] csa_component24_fa15_xor1;
  wire [0:0] csa_component24_fa15_or0;
  wire [0:0] csa_component24_fa16_xor1;
  wire [0:0] csa_component24_fa16_or0;
  wire [0:0] csa_component24_fa17_xor1;
  wire [0:0] csa_component24_fa17_or0;
  wire [0:0] csa_component24_fa18_xor1;
  wire [0:0] csa_component24_fa18_or0;
  wire [0:0] csa_component24_fa19_xor1;
  wire [0:0] csa_component24_fa19_or0;
  wire [0:0] csa_component24_fa20_xor1;
  wire [0:0] csa_component24_fa20_or0;
  wire [0:0] csa_component24_fa21_xor1;
  wire [0:0] csa_component24_fa21_or0;
  wire [0:0] csa_component24_fa22_xor1;
  wire [0:0] csa_component24_fa22_or0;
  wire [0:0] csa_component24_fa23_xor1;
  wire [0:0] csa_component24_fa23_or0;

  fa fa_csa_component24_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component24_fa0_xor1), .fa_or0(csa_component24_fa0_or0));
  fa fa_csa_component24_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component24_fa1_xor1), .fa_or0(csa_component24_fa1_or0));
  fa fa_csa_component24_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component24_fa2_xor1), .fa_or0(csa_component24_fa2_or0));
  fa fa_csa_component24_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component24_fa3_xor1), .fa_or0(csa_component24_fa3_or0));
  fa fa_csa_component24_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component24_fa4_xor1), .fa_or0(csa_component24_fa4_or0));
  fa fa_csa_component24_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component24_fa5_xor1), .fa_or0(csa_component24_fa5_or0));
  fa fa_csa_component24_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component24_fa6_xor1), .fa_or0(csa_component24_fa6_or0));
  fa fa_csa_component24_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component24_fa7_xor1), .fa_or0(csa_component24_fa7_or0));
  fa fa_csa_component24_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component24_fa8_xor1), .fa_or0(csa_component24_fa8_or0));
  fa fa_csa_component24_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component24_fa9_xor1), .fa_or0(csa_component24_fa9_or0));
  fa fa_csa_component24_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component24_fa10_xor1), .fa_or0(csa_component24_fa10_or0));
  fa fa_csa_component24_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component24_fa11_xor1), .fa_or0(csa_component24_fa11_or0));
  fa fa_csa_component24_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component24_fa12_xor1), .fa_or0(csa_component24_fa12_or0));
  fa fa_csa_component24_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component24_fa13_xor1), .fa_or0(csa_component24_fa13_or0));
  fa fa_csa_component24_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component24_fa14_xor1), .fa_or0(csa_component24_fa14_or0));
  fa fa_csa_component24_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component24_fa15_xor1), .fa_or0(csa_component24_fa15_or0));
  fa fa_csa_component24_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component24_fa16_xor1), .fa_or0(csa_component24_fa16_or0));
  fa fa_csa_component24_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component24_fa17_xor1), .fa_or0(csa_component24_fa17_or0));
  fa fa_csa_component24_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component24_fa18_xor1), .fa_or0(csa_component24_fa18_or0));
  fa fa_csa_component24_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component24_fa19_xor1), .fa_or0(csa_component24_fa19_or0));
  fa fa_csa_component24_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component24_fa20_xor1), .fa_or0(csa_component24_fa20_or0));
  fa fa_csa_component24_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component24_fa21_xor1), .fa_or0(csa_component24_fa21_or0));
  fa fa_csa_component24_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component24_fa22_xor1), .fa_or0(csa_component24_fa22_or0));
  fa fa_csa_component24_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component24_fa23_xor1), .fa_or0(csa_component24_fa23_or0));

  assign csa_component24_out[0] = csa_component24_fa0_xor1[0];
  assign csa_component24_out[1] = csa_component24_fa1_xor1[0];
  assign csa_component24_out[2] = csa_component24_fa2_xor1[0];
  assign csa_component24_out[3] = csa_component24_fa3_xor1[0];
  assign csa_component24_out[4] = csa_component24_fa4_xor1[0];
  assign csa_component24_out[5] = csa_component24_fa5_xor1[0];
  assign csa_component24_out[6] = csa_component24_fa6_xor1[0];
  assign csa_component24_out[7] = csa_component24_fa7_xor1[0];
  assign csa_component24_out[8] = csa_component24_fa8_xor1[0];
  assign csa_component24_out[9] = csa_component24_fa9_xor1[0];
  assign csa_component24_out[10] = csa_component24_fa10_xor1[0];
  assign csa_component24_out[11] = csa_component24_fa11_xor1[0];
  assign csa_component24_out[12] = csa_component24_fa12_xor1[0];
  assign csa_component24_out[13] = csa_component24_fa13_xor1[0];
  assign csa_component24_out[14] = csa_component24_fa14_xor1[0];
  assign csa_component24_out[15] = csa_component24_fa15_xor1[0];
  assign csa_component24_out[16] = csa_component24_fa16_xor1[0];
  assign csa_component24_out[17] = csa_component24_fa17_xor1[0];
  assign csa_component24_out[18] = csa_component24_fa18_xor1[0];
  assign csa_component24_out[19] = csa_component24_fa19_xor1[0];
  assign csa_component24_out[20] = csa_component24_fa20_xor1[0];
  assign csa_component24_out[21] = csa_component24_fa21_xor1[0];
  assign csa_component24_out[22] = csa_component24_fa22_xor1[0];
  assign csa_component24_out[23] = csa_component24_fa23_xor1[0];
  assign csa_component24_out[24] = 1'b0;
  assign csa_component24_out[25] = 1'b0;
  assign csa_component24_out[26] = csa_component24_fa0_or0[0];
  assign csa_component24_out[27] = csa_component24_fa1_or0[0];
  assign csa_component24_out[28] = csa_component24_fa2_or0[0];
  assign csa_component24_out[29] = csa_component24_fa3_or0[0];
  assign csa_component24_out[30] = csa_component24_fa4_or0[0];
  assign csa_component24_out[31] = csa_component24_fa5_or0[0];
  assign csa_component24_out[32] = csa_component24_fa6_or0[0];
  assign csa_component24_out[33] = csa_component24_fa7_or0[0];
  assign csa_component24_out[34] = csa_component24_fa8_or0[0];
  assign csa_component24_out[35] = csa_component24_fa9_or0[0];
  assign csa_component24_out[36] = csa_component24_fa10_or0[0];
  assign csa_component24_out[37] = csa_component24_fa11_or0[0];
  assign csa_component24_out[38] = csa_component24_fa12_or0[0];
  assign csa_component24_out[39] = csa_component24_fa13_or0[0];
  assign csa_component24_out[40] = csa_component24_fa14_or0[0];
  assign csa_component24_out[41] = csa_component24_fa15_or0[0];
  assign csa_component24_out[42] = csa_component24_fa16_or0[0];
  assign csa_component24_out[43] = csa_component24_fa17_or0[0];
  assign csa_component24_out[44] = csa_component24_fa18_or0[0];
  assign csa_component24_out[45] = csa_component24_fa19_or0[0];
  assign csa_component24_out[46] = csa_component24_fa20_or0[0];
  assign csa_component24_out[47] = csa_component24_fa21_or0[0];
  assign csa_component24_out[48] = csa_component24_fa22_or0[0];
  assign csa_component24_out[49] = csa_component24_fa23_or0[0];
endmodule

module csa_component27(input [26:0] a, input [26:0] b, input [26:0] c, output [55:0] csa_component27_out);
  wire [0:0] csa_component27_fa0_xor1;
  wire [0:0] csa_component27_fa0_or0;
  wire [0:0] csa_component27_fa1_xor1;
  wire [0:0] csa_component27_fa1_or0;
  wire [0:0] csa_component27_fa2_xor1;
  wire [0:0] csa_component27_fa2_or0;
  wire [0:0] csa_component27_fa3_xor1;
  wire [0:0] csa_component27_fa3_or0;
  wire [0:0] csa_component27_fa4_xor1;
  wire [0:0] csa_component27_fa4_or0;
  wire [0:0] csa_component27_fa5_xor1;
  wire [0:0] csa_component27_fa5_or0;
  wire [0:0] csa_component27_fa6_xor1;
  wire [0:0] csa_component27_fa6_or0;
  wire [0:0] csa_component27_fa7_xor1;
  wire [0:0] csa_component27_fa7_or0;
  wire [0:0] csa_component27_fa8_xor1;
  wire [0:0] csa_component27_fa8_or0;
  wire [0:0] csa_component27_fa9_xor1;
  wire [0:0] csa_component27_fa9_or0;
  wire [0:0] csa_component27_fa10_xor1;
  wire [0:0] csa_component27_fa10_or0;
  wire [0:0] csa_component27_fa11_xor1;
  wire [0:0] csa_component27_fa11_or0;
  wire [0:0] csa_component27_fa12_xor1;
  wire [0:0] csa_component27_fa12_or0;
  wire [0:0] csa_component27_fa13_xor1;
  wire [0:0] csa_component27_fa13_or0;
  wire [0:0] csa_component27_fa14_xor1;
  wire [0:0] csa_component27_fa14_or0;
  wire [0:0] csa_component27_fa15_xor1;
  wire [0:0] csa_component27_fa15_or0;
  wire [0:0] csa_component27_fa16_xor1;
  wire [0:0] csa_component27_fa16_or0;
  wire [0:0] csa_component27_fa17_xor1;
  wire [0:0] csa_component27_fa17_or0;
  wire [0:0] csa_component27_fa18_xor1;
  wire [0:0] csa_component27_fa18_or0;
  wire [0:0] csa_component27_fa19_xor1;
  wire [0:0] csa_component27_fa19_or0;
  wire [0:0] csa_component27_fa20_xor1;
  wire [0:0] csa_component27_fa20_or0;
  wire [0:0] csa_component27_fa21_xor1;
  wire [0:0] csa_component27_fa21_or0;
  wire [0:0] csa_component27_fa22_xor1;
  wire [0:0] csa_component27_fa22_or0;
  wire [0:0] csa_component27_fa23_xor1;
  wire [0:0] csa_component27_fa23_or0;
  wire [0:0] csa_component27_fa24_xor1;
  wire [0:0] csa_component27_fa24_or0;
  wire [0:0] csa_component27_fa25_xor1;
  wire [0:0] csa_component27_fa25_or0;
  wire [0:0] csa_component27_fa26_xor1;
  wire [0:0] csa_component27_fa26_or0;

  fa fa_csa_component27_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component27_fa0_xor1), .fa_or0(csa_component27_fa0_or0));
  fa fa_csa_component27_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component27_fa1_xor1), .fa_or0(csa_component27_fa1_or0));
  fa fa_csa_component27_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component27_fa2_xor1), .fa_or0(csa_component27_fa2_or0));
  fa fa_csa_component27_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component27_fa3_xor1), .fa_or0(csa_component27_fa3_or0));
  fa fa_csa_component27_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component27_fa4_xor1), .fa_or0(csa_component27_fa4_or0));
  fa fa_csa_component27_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component27_fa5_xor1), .fa_or0(csa_component27_fa5_or0));
  fa fa_csa_component27_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component27_fa6_xor1), .fa_or0(csa_component27_fa6_or0));
  fa fa_csa_component27_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component27_fa7_xor1), .fa_or0(csa_component27_fa7_or0));
  fa fa_csa_component27_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component27_fa8_xor1), .fa_or0(csa_component27_fa8_or0));
  fa fa_csa_component27_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component27_fa9_xor1), .fa_or0(csa_component27_fa9_or0));
  fa fa_csa_component27_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component27_fa10_xor1), .fa_or0(csa_component27_fa10_or0));
  fa fa_csa_component27_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component27_fa11_xor1), .fa_or0(csa_component27_fa11_or0));
  fa fa_csa_component27_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component27_fa12_xor1), .fa_or0(csa_component27_fa12_or0));
  fa fa_csa_component27_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component27_fa13_xor1), .fa_or0(csa_component27_fa13_or0));
  fa fa_csa_component27_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component27_fa14_xor1), .fa_or0(csa_component27_fa14_or0));
  fa fa_csa_component27_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component27_fa15_xor1), .fa_or0(csa_component27_fa15_or0));
  fa fa_csa_component27_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component27_fa16_xor1), .fa_or0(csa_component27_fa16_or0));
  fa fa_csa_component27_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component27_fa17_xor1), .fa_or0(csa_component27_fa17_or0));
  fa fa_csa_component27_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component27_fa18_xor1), .fa_or0(csa_component27_fa18_or0));
  fa fa_csa_component27_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component27_fa19_xor1), .fa_or0(csa_component27_fa19_or0));
  fa fa_csa_component27_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component27_fa20_xor1), .fa_or0(csa_component27_fa20_or0));
  fa fa_csa_component27_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component27_fa21_xor1), .fa_or0(csa_component27_fa21_or0));
  fa fa_csa_component27_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component27_fa22_xor1), .fa_or0(csa_component27_fa22_or0));
  fa fa_csa_component27_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component27_fa23_xor1), .fa_or0(csa_component27_fa23_or0));
  fa fa_csa_component27_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component27_fa24_xor1), .fa_or0(csa_component27_fa24_or0));
  fa fa_csa_component27_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component27_fa25_xor1), .fa_or0(csa_component27_fa25_or0));
  fa fa_csa_component27_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component27_fa26_xor1), .fa_or0(csa_component27_fa26_or0));

  assign csa_component27_out[0] = csa_component27_fa0_xor1[0];
  assign csa_component27_out[1] = csa_component27_fa1_xor1[0];
  assign csa_component27_out[2] = csa_component27_fa2_xor1[0];
  assign csa_component27_out[3] = csa_component27_fa3_xor1[0];
  assign csa_component27_out[4] = csa_component27_fa4_xor1[0];
  assign csa_component27_out[5] = csa_component27_fa5_xor1[0];
  assign csa_component27_out[6] = csa_component27_fa6_xor1[0];
  assign csa_component27_out[7] = csa_component27_fa7_xor1[0];
  assign csa_component27_out[8] = csa_component27_fa8_xor1[0];
  assign csa_component27_out[9] = csa_component27_fa9_xor1[0];
  assign csa_component27_out[10] = csa_component27_fa10_xor1[0];
  assign csa_component27_out[11] = csa_component27_fa11_xor1[0];
  assign csa_component27_out[12] = csa_component27_fa12_xor1[0];
  assign csa_component27_out[13] = csa_component27_fa13_xor1[0];
  assign csa_component27_out[14] = csa_component27_fa14_xor1[0];
  assign csa_component27_out[15] = csa_component27_fa15_xor1[0];
  assign csa_component27_out[16] = csa_component27_fa16_xor1[0];
  assign csa_component27_out[17] = csa_component27_fa17_xor1[0];
  assign csa_component27_out[18] = csa_component27_fa18_xor1[0];
  assign csa_component27_out[19] = csa_component27_fa19_xor1[0];
  assign csa_component27_out[20] = csa_component27_fa20_xor1[0];
  assign csa_component27_out[21] = csa_component27_fa21_xor1[0];
  assign csa_component27_out[22] = csa_component27_fa22_xor1[0];
  assign csa_component27_out[23] = csa_component27_fa23_xor1[0];
  assign csa_component27_out[24] = csa_component27_fa24_xor1[0];
  assign csa_component27_out[25] = csa_component27_fa25_xor1[0];
  assign csa_component27_out[26] = csa_component27_fa26_xor1[0];
  assign csa_component27_out[27] = 1'b0;
  assign csa_component27_out[28] = 1'b0;
  assign csa_component27_out[29] = csa_component27_fa0_or0[0];
  assign csa_component27_out[30] = csa_component27_fa1_or0[0];
  assign csa_component27_out[31] = csa_component27_fa2_or0[0];
  assign csa_component27_out[32] = csa_component27_fa3_or0[0];
  assign csa_component27_out[33] = csa_component27_fa4_or0[0];
  assign csa_component27_out[34] = csa_component27_fa5_or0[0];
  assign csa_component27_out[35] = csa_component27_fa6_or0[0];
  assign csa_component27_out[36] = csa_component27_fa7_or0[0];
  assign csa_component27_out[37] = csa_component27_fa8_or0[0];
  assign csa_component27_out[38] = csa_component27_fa9_or0[0];
  assign csa_component27_out[39] = csa_component27_fa10_or0[0];
  assign csa_component27_out[40] = csa_component27_fa11_or0[0];
  assign csa_component27_out[41] = csa_component27_fa12_or0[0];
  assign csa_component27_out[42] = csa_component27_fa13_or0[0];
  assign csa_component27_out[43] = csa_component27_fa14_or0[0];
  assign csa_component27_out[44] = csa_component27_fa15_or0[0];
  assign csa_component27_out[45] = csa_component27_fa16_or0[0];
  assign csa_component27_out[46] = csa_component27_fa17_or0[0];
  assign csa_component27_out[47] = csa_component27_fa18_or0[0];
  assign csa_component27_out[48] = csa_component27_fa19_or0[0];
  assign csa_component27_out[49] = csa_component27_fa20_or0[0];
  assign csa_component27_out[50] = csa_component27_fa21_or0[0];
  assign csa_component27_out[51] = csa_component27_fa22_or0[0];
  assign csa_component27_out[52] = csa_component27_fa23_or0[0];
  assign csa_component27_out[53] = csa_component27_fa24_or0[0];
  assign csa_component27_out[54] = csa_component27_fa25_or0[0];
  assign csa_component27_out[55] = csa_component27_fa26_or0[0];
endmodule

module csa_component30(input [29:0] a, input [29:0] b, input [29:0] c, output [61:0] csa_component30_out);
  wire [0:0] csa_component30_fa0_xor1;
  wire [0:0] csa_component30_fa0_or0;
  wire [0:0] csa_component30_fa1_xor1;
  wire [0:0] csa_component30_fa1_or0;
  wire [0:0] csa_component30_fa2_xor1;
  wire [0:0] csa_component30_fa2_or0;
  wire [0:0] csa_component30_fa3_xor1;
  wire [0:0] csa_component30_fa3_or0;
  wire [0:0] csa_component30_fa4_xor1;
  wire [0:0] csa_component30_fa4_or0;
  wire [0:0] csa_component30_fa5_xor1;
  wire [0:0] csa_component30_fa5_or0;
  wire [0:0] csa_component30_fa6_xor1;
  wire [0:0] csa_component30_fa6_or0;
  wire [0:0] csa_component30_fa7_xor1;
  wire [0:0] csa_component30_fa7_or0;
  wire [0:0] csa_component30_fa8_xor1;
  wire [0:0] csa_component30_fa8_or0;
  wire [0:0] csa_component30_fa9_xor1;
  wire [0:0] csa_component30_fa9_or0;
  wire [0:0] csa_component30_fa10_xor1;
  wire [0:0] csa_component30_fa10_or0;
  wire [0:0] csa_component30_fa11_xor1;
  wire [0:0] csa_component30_fa11_or0;
  wire [0:0] csa_component30_fa12_xor1;
  wire [0:0] csa_component30_fa12_or0;
  wire [0:0] csa_component30_fa13_xor1;
  wire [0:0] csa_component30_fa13_or0;
  wire [0:0] csa_component30_fa14_xor1;
  wire [0:0] csa_component30_fa14_or0;
  wire [0:0] csa_component30_fa15_xor1;
  wire [0:0] csa_component30_fa15_or0;
  wire [0:0] csa_component30_fa16_xor1;
  wire [0:0] csa_component30_fa16_or0;
  wire [0:0] csa_component30_fa17_xor1;
  wire [0:0] csa_component30_fa17_or0;
  wire [0:0] csa_component30_fa18_xor1;
  wire [0:0] csa_component30_fa18_or0;
  wire [0:0] csa_component30_fa19_xor1;
  wire [0:0] csa_component30_fa19_or0;
  wire [0:0] csa_component30_fa20_xor1;
  wire [0:0] csa_component30_fa20_or0;
  wire [0:0] csa_component30_fa21_xor1;
  wire [0:0] csa_component30_fa21_or0;
  wire [0:0] csa_component30_fa22_xor1;
  wire [0:0] csa_component30_fa22_or0;
  wire [0:0] csa_component30_fa23_xor1;
  wire [0:0] csa_component30_fa23_or0;
  wire [0:0] csa_component30_fa24_xor1;
  wire [0:0] csa_component30_fa24_or0;
  wire [0:0] csa_component30_fa25_xor1;
  wire [0:0] csa_component30_fa25_or0;
  wire [0:0] csa_component30_fa26_xor1;
  wire [0:0] csa_component30_fa26_or0;
  wire [0:0] csa_component30_fa27_xor1;
  wire [0:0] csa_component30_fa27_or0;
  wire [0:0] csa_component30_fa28_xor1;
  wire [0:0] csa_component30_fa28_or0;
  wire [0:0] csa_component30_fa29_xor1;
  wire [0:0] csa_component30_fa29_or0;

  fa fa_csa_component30_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component30_fa0_xor1), .fa_or0(csa_component30_fa0_or0));
  fa fa_csa_component30_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component30_fa1_xor1), .fa_or0(csa_component30_fa1_or0));
  fa fa_csa_component30_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component30_fa2_xor1), .fa_or0(csa_component30_fa2_or0));
  fa fa_csa_component30_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component30_fa3_xor1), .fa_or0(csa_component30_fa3_or0));
  fa fa_csa_component30_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component30_fa4_xor1), .fa_or0(csa_component30_fa4_or0));
  fa fa_csa_component30_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component30_fa5_xor1), .fa_or0(csa_component30_fa5_or0));
  fa fa_csa_component30_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component30_fa6_xor1), .fa_or0(csa_component30_fa6_or0));
  fa fa_csa_component30_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component30_fa7_xor1), .fa_or0(csa_component30_fa7_or0));
  fa fa_csa_component30_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component30_fa8_xor1), .fa_or0(csa_component30_fa8_or0));
  fa fa_csa_component30_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component30_fa9_xor1), .fa_or0(csa_component30_fa9_or0));
  fa fa_csa_component30_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component30_fa10_xor1), .fa_or0(csa_component30_fa10_or0));
  fa fa_csa_component30_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component30_fa11_xor1), .fa_or0(csa_component30_fa11_or0));
  fa fa_csa_component30_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component30_fa12_xor1), .fa_or0(csa_component30_fa12_or0));
  fa fa_csa_component30_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component30_fa13_xor1), .fa_or0(csa_component30_fa13_or0));
  fa fa_csa_component30_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component30_fa14_xor1), .fa_or0(csa_component30_fa14_or0));
  fa fa_csa_component30_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component30_fa15_xor1), .fa_or0(csa_component30_fa15_or0));
  fa fa_csa_component30_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component30_fa16_xor1), .fa_or0(csa_component30_fa16_or0));
  fa fa_csa_component30_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component30_fa17_xor1), .fa_or0(csa_component30_fa17_or0));
  fa fa_csa_component30_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component30_fa18_xor1), .fa_or0(csa_component30_fa18_or0));
  fa fa_csa_component30_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component30_fa19_xor1), .fa_or0(csa_component30_fa19_or0));
  fa fa_csa_component30_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component30_fa20_xor1), .fa_or0(csa_component30_fa20_or0));
  fa fa_csa_component30_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component30_fa21_xor1), .fa_or0(csa_component30_fa21_or0));
  fa fa_csa_component30_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component30_fa22_xor1), .fa_or0(csa_component30_fa22_or0));
  fa fa_csa_component30_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component30_fa23_xor1), .fa_or0(csa_component30_fa23_or0));
  fa fa_csa_component30_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component30_fa24_xor1), .fa_or0(csa_component30_fa24_or0));
  fa fa_csa_component30_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component30_fa25_xor1), .fa_or0(csa_component30_fa25_or0));
  fa fa_csa_component30_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component30_fa26_xor1), .fa_or0(csa_component30_fa26_or0));
  fa fa_csa_component30_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component30_fa27_xor1), .fa_or0(csa_component30_fa27_or0));
  fa fa_csa_component30_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component30_fa28_xor1), .fa_or0(csa_component30_fa28_or0));
  fa fa_csa_component30_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component30_fa29_xor1), .fa_or0(csa_component30_fa29_or0));

  assign csa_component30_out[0] = csa_component30_fa0_xor1[0];
  assign csa_component30_out[1] = csa_component30_fa1_xor1[0];
  assign csa_component30_out[2] = csa_component30_fa2_xor1[0];
  assign csa_component30_out[3] = csa_component30_fa3_xor1[0];
  assign csa_component30_out[4] = csa_component30_fa4_xor1[0];
  assign csa_component30_out[5] = csa_component30_fa5_xor1[0];
  assign csa_component30_out[6] = csa_component30_fa6_xor1[0];
  assign csa_component30_out[7] = csa_component30_fa7_xor1[0];
  assign csa_component30_out[8] = csa_component30_fa8_xor1[0];
  assign csa_component30_out[9] = csa_component30_fa9_xor1[0];
  assign csa_component30_out[10] = csa_component30_fa10_xor1[0];
  assign csa_component30_out[11] = csa_component30_fa11_xor1[0];
  assign csa_component30_out[12] = csa_component30_fa12_xor1[0];
  assign csa_component30_out[13] = csa_component30_fa13_xor1[0];
  assign csa_component30_out[14] = csa_component30_fa14_xor1[0];
  assign csa_component30_out[15] = csa_component30_fa15_xor1[0];
  assign csa_component30_out[16] = csa_component30_fa16_xor1[0];
  assign csa_component30_out[17] = csa_component30_fa17_xor1[0];
  assign csa_component30_out[18] = csa_component30_fa18_xor1[0];
  assign csa_component30_out[19] = csa_component30_fa19_xor1[0];
  assign csa_component30_out[20] = csa_component30_fa20_xor1[0];
  assign csa_component30_out[21] = csa_component30_fa21_xor1[0];
  assign csa_component30_out[22] = csa_component30_fa22_xor1[0];
  assign csa_component30_out[23] = csa_component30_fa23_xor1[0];
  assign csa_component30_out[24] = csa_component30_fa24_xor1[0];
  assign csa_component30_out[25] = csa_component30_fa25_xor1[0];
  assign csa_component30_out[26] = csa_component30_fa26_xor1[0];
  assign csa_component30_out[27] = csa_component30_fa27_xor1[0];
  assign csa_component30_out[28] = csa_component30_fa28_xor1[0];
  assign csa_component30_out[29] = csa_component30_fa29_xor1[0];
  assign csa_component30_out[30] = 1'b0;
  assign csa_component30_out[31] = 1'b0;
  assign csa_component30_out[32] = csa_component30_fa0_or0[0];
  assign csa_component30_out[33] = csa_component30_fa1_or0[0];
  assign csa_component30_out[34] = csa_component30_fa2_or0[0];
  assign csa_component30_out[35] = csa_component30_fa3_or0[0];
  assign csa_component30_out[36] = csa_component30_fa4_or0[0];
  assign csa_component30_out[37] = csa_component30_fa5_or0[0];
  assign csa_component30_out[38] = csa_component30_fa6_or0[0];
  assign csa_component30_out[39] = csa_component30_fa7_or0[0];
  assign csa_component30_out[40] = csa_component30_fa8_or0[0];
  assign csa_component30_out[41] = csa_component30_fa9_or0[0];
  assign csa_component30_out[42] = csa_component30_fa10_or0[0];
  assign csa_component30_out[43] = csa_component30_fa11_or0[0];
  assign csa_component30_out[44] = csa_component30_fa12_or0[0];
  assign csa_component30_out[45] = csa_component30_fa13_or0[0];
  assign csa_component30_out[46] = csa_component30_fa14_or0[0];
  assign csa_component30_out[47] = csa_component30_fa15_or0[0];
  assign csa_component30_out[48] = csa_component30_fa16_or0[0];
  assign csa_component30_out[49] = csa_component30_fa17_or0[0];
  assign csa_component30_out[50] = csa_component30_fa18_or0[0];
  assign csa_component30_out[51] = csa_component30_fa19_or0[0];
  assign csa_component30_out[52] = csa_component30_fa20_or0[0];
  assign csa_component30_out[53] = csa_component30_fa21_or0[0];
  assign csa_component30_out[54] = csa_component30_fa22_or0[0];
  assign csa_component30_out[55] = csa_component30_fa23_or0[0];
  assign csa_component30_out[56] = csa_component30_fa24_or0[0];
  assign csa_component30_out[57] = csa_component30_fa25_or0[0];
  assign csa_component30_out[58] = csa_component30_fa26_or0[0];
  assign csa_component30_out[59] = csa_component30_fa27_or0[0];
  assign csa_component30_out[60] = csa_component30_fa28_or0[0];
  assign csa_component30_out[61] = csa_component30_fa29_or0[0];
endmodule

module csa_component22(input [21:0] a, input [21:0] b, input [21:0] c, output [45:0] csa_component22_out);
  wire [0:0] csa_component22_fa0_xor1;
  wire [0:0] csa_component22_fa0_or0;
  wire [0:0] csa_component22_fa1_xor1;
  wire [0:0] csa_component22_fa1_or0;
  wire [0:0] csa_component22_fa2_xor1;
  wire [0:0] csa_component22_fa2_or0;
  wire [0:0] csa_component22_fa3_xor1;
  wire [0:0] csa_component22_fa3_or0;
  wire [0:0] csa_component22_fa4_xor1;
  wire [0:0] csa_component22_fa4_or0;
  wire [0:0] csa_component22_fa5_xor1;
  wire [0:0] csa_component22_fa5_or0;
  wire [0:0] csa_component22_fa6_xor1;
  wire [0:0] csa_component22_fa6_or0;
  wire [0:0] csa_component22_fa7_xor1;
  wire [0:0] csa_component22_fa7_or0;
  wire [0:0] csa_component22_fa8_xor1;
  wire [0:0] csa_component22_fa8_or0;
  wire [0:0] csa_component22_fa9_xor1;
  wire [0:0] csa_component22_fa9_or0;
  wire [0:0] csa_component22_fa10_xor1;
  wire [0:0] csa_component22_fa10_or0;
  wire [0:0] csa_component22_fa11_xor1;
  wire [0:0] csa_component22_fa11_or0;
  wire [0:0] csa_component22_fa12_xor1;
  wire [0:0] csa_component22_fa12_or0;
  wire [0:0] csa_component22_fa13_xor1;
  wire [0:0] csa_component22_fa13_or0;
  wire [0:0] csa_component22_fa14_xor1;
  wire [0:0] csa_component22_fa14_or0;
  wire [0:0] csa_component22_fa15_xor1;
  wire [0:0] csa_component22_fa15_or0;
  wire [0:0] csa_component22_fa16_xor1;
  wire [0:0] csa_component22_fa16_or0;
  wire [0:0] csa_component22_fa17_xor1;
  wire [0:0] csa_component22_fa17_or0;
  wire [0:0] csa_component22_fa18_xor1;
  wire [0:0] csa_component22_fa18_or0;
  wire [0:0] csa_component22_fa19_xor1;
  wire [0:0] csa_component22_fa19_or0;
  wire [0:0] csa_component22_fa20_xor1;
  wire [0:0] csa_component22_fa20_or0;
  wire [0:0] csa_component22_fa21_xor1;
  wire [0:0] csa_component22_fa21_or0;

  fa fa_csa_component22_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component22_fa0_xor1), .fa_or0(csa_component22_fa0_or0));
  fa fa_csa_component22_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component22_fa1_xor1), .fa_or0(csa_component22_fa1_or0));
  fa fa_csa_component22_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component22_fa2_xor1), .fa_or0(csa_component22_fa2_or0));
  fa fa_csa_component22_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component22_fa3_xor1), .fa_or0(csa_component22_fa3_or0));
  fa fa_csa_component22_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component22_fa4_xor1), .fa_or0(csa_component22_fa4_or0));
  fa fa_csa_component22_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component22_fa5_xor1), .fa_or0(csa_component22_fa5_or0));
  fa fa_csa_component22_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component22_fa6_xor1), .fa_or0(csa_component22_fa6_or0));
  fa fa_csa_component22_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component22_fa7_xor1), .fa_or0(csa_component22_fa7_or0));
  fa fa_csa_component22_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component22_fa8_xor1), .fa_or0(csa_component22_fa8_or0));
  fa fa_csa_component22_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component22_fa9_xor1), .fa_or0(csa_component22_fa9_or0));
  fa fa_csa_component22_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component22_fa10_xor1), .fa_or0(csa_component22_fa10_or0));
  fa fa_csa_component22_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component22_fa11_xor1), .fa_or0(csa_component22_fa11_or0));
  fa fa_csa_component22_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component22_fa12_xor1), .fa_or0(csa_component22_fa12_or0));
  fa fa_csa_component22_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component22_fa13_xor1), .fa_or0(csa_component22_fa13_or0));
  fa fa_csa_component22_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component22_fa14_xor1), .fa_or0(csa_component22_fa14_or0));
  fa fa_csa_component22_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component22_fa15_xor1), .fa_or0(csa_component22_fa15_or0));
  fa fa_csa_component22_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component22_fa16_xor1), .fa_or0(csa_component22_fa16_or0));
  fa fa_csa_component22_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component22_fa17_xor1), .fa_or0(csa_component22_fa17_or0));
  fa fa_csa_component22_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component22_fa18_xor1), .fa_or0(csa_component22_fa18_or0));
  fa fa_csa_component22_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component22_fa19_xor1), .fa_or0(csa_component22_fa19_or0));
  fa fa_csa_component22_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component22_fa20_xor1), .fa_or0(csa_component22_fa20_or0));
  fa fa_csa_component22_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component22_fa21_xor1), .fa_or0(csa_component22_fa21_or0));

  assign csa_component22_out[0] = csa_component22_fa0_xor1[0];
  assign csa_component22_out[1] = csa_component22_fa1_xor1[0];
  assign csa_component22_out[2] = csa_component22_fa2_xor1[0];
  assign csa_component22_out[3] = csa_component22_fa3_xor1[0];
  assign csa_component22_out[4] = csa_component22_fa4_xor1[0];
  assign csa_component22_out[5] = csa_component22_fa5_xor1[0];
  assign csa_component22_out[6] = csa_component22_fa6_xor1[0];
  assign csa_component22_out[7] = csa_component22_fa7_xor1[0];
  assign csa_component22_out[8] = csa_component22_fa8_xor1[0];
  assign csa_component22_out[9] = csa_component22_fa9_xor1[0];
  assign csa_component22_out[10] = csa_component22_fa10_xor1[0];
  assign csa_component22_out[11] = csa_component22_fa11_xor1[0];
  assign csa_component22_out[12] = csa_component22_fa12_xor1[0];
  assign csa_component22_out[13] = csa_component22_fa13_xor1[0];
  assign csa_component22_out[14] = csa_component22_fa14_xor1[0];
  assign csa_component22_out[15] = csa_component22_fa15_xor1[0];
  assign csa_component22_out[16] = csa_component22_fa16_xor1[0];
  assign csa_component22_out[17] = csa_component22_fa17_xor1[0];
  assign csa_component22_out[18] = csa_component22_fa18_xor1[0];
  assign csa_component22_out[19] = csa_component22_fa19_xor1[0];
  assign csa_component22_out[20] = csa_component22_fa20_xor1[0];
  assign csa_component22_out[21] = csa_component22_fa21_xor1[0];
  assign csa_component22_out[22] = 1'b0;
  assign csa_component22_out[23] = 1'b0;
  assign csa_component22_out[24] = csa_component22_fa0_or0[0];
  assign csa_component22_out[25] = csa_component22_fa1_or0[0];
  assign csa_component22_out[26] = csa_component22_fa2_or0[0];
  assign csa_component22_out[27] = csa_component22_fa3_or0[0];
  assign csa_component22_out[28] = csa_component22_fa4_or0[0];
  assign csa_component22_out[29] = csa_component22_fa5_or0[0];
  assign csa_component22_out[30] = csa_component22_fa6_or0[0];
  assign csa_component22_out[31] = csa_component22_fa7_or0[0];
  assign csa_component22_out[32] = csa_component22_fa8_or0[0];
  assign csa_component22_out[33] = csa_component22_fa9_or0[0];
  assign csa_component22_out[34] = csa_component22_fa10_or0[0];
  assign csa_component22_out[35] = csa_component22_fa11_or0[0];
  assign csa_component22_out[36] = csa_component22_fa12_or0[0];
  assign csa_component22_out[37] = csa_component22_fa13_or0[0];
  assign csa_component22_out[38] = csa_component22_fa14_or0[0];
  assign csa_component22_out[39] = csa_component22_fa15_or0[0];
  assign csa_component22_out[40] = csa_component22_fa16_or0[0];
  assign csa_component22_out[41] = csa_component22_fa17_or0[0];
  assign csa_component22_out[42] = csa_component22_fa18_or0[0];
  assign csa_component22_out[43] = csa_component22_fa19_or0[0];
  assign csa_component22_out[44] = csa_component22_fa20_or0[0];
  assign csa_component22_out[45] = csa_component22_fa21_or0[0];
endmodule

module csa_component25(input [24:0] a, input [24:0] b, input [24:0] c, output [51:0] csa_component25_out);
  wire [0:0] csa_component25_fa0_xor1;
  wire [0:0] csa_component25_fa0_or0;
  wire [0:0] csa_component25_fa1_xor1;
  wire [0:0] csa_component25_fa1_or0;
  wire [0:0] csa_component25_fa2_xor1;
  wire [0:0] csa_component25_fa2_or0;
  wire [0:0] csa_component25_fa3_xor1;
  wire [0:0] csa_component25_fa3_or0;
  wire [0:0] csa_component25_fa4_xor1;
  wire [0:0] csa_component25_fa4_or0;
  wire [0:0] csa_component25_fa5_xor1;
  wire [0:0] csa_component25_fa5_or0;
  wire [0:0] csa_component25_fa6_xor1;
  wire [0:0] csa_component25_fa6_or0;
  wire [0:0] csa_component25_fa7_xor1;
  wire [0:0] csa_component25_fa7_or0;
  wire [0:0] csa_component25_fa8_xor1;
  wire [0:0] csa_component25_fa8_or0;
  wire [0:0] csa_component25_fa9_xor1;
  wire [0:0] csa_component25_fa9_or0;
  wire [0:0] csa_component25_fa10_xor1;
  wire [0:0] csa_component25_fa10_or0;
  wire [0:0] csa_component25_fa11_xor1;
  wire [0:0] csa_component25_fa11_or0;
  wire [0:0] csa_component25_fa12_xor1;
  wire [0:0] csa_component25_fa12_or0;
  wire [0:0] csa_component25_fa13_xor1;
  wire [0:0] csa_component25_fa13_or0;
  wire [0:0] csa_component25_fa14_xor1;
  wire [0:0] csa_component25_fa14_or0;
  wire [0:0] csa_component25_fa15_xor1;
  wire [0:0] csa_component25_fa15_or0;
  wire [0:0] csa_component25_fa16_xor1;
  wire [0:0] csa_component25_fa16_or0;
  wire [0:0] csa_component25_fa17_xor1;
  wire [0:0] csa_component25_fa17_or0;
  wire [0:0] csa_component25_fa18_xor1;
  wire [0:0] csa_component25_fa18_or0;
  wire [0:0] csa_component25_fa19_xor1;
  wire [0:0] csa_component25_fa19_or0;
  wire [0:0] csa_component25_fa20_xor1;
  wire [0:0] csa_component25_fa20_or0;
  wire [0:0] csa_component25_fa21_xor1;
  wire [0:0] csa_component25_fa21_or0;
  wire [0:0] csa_component25_fa22_xor1;
  wire [0:0] csa_component25_fa22_or0;
  wire [0:0] csa_component25_fa23_xor1;
  wire [0:0] csa_component25_fa23_or0;
  wire [0:0] csa_component25_fa24_xor1;
  wire [0:0] csa_component25_fa24_or0;

  fa fa_csa_component25_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component25_fa0_xor1), .fa_or0(csa_component25_fa0_or0));
  fa fa_csa_component25_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component25_fa1_xor1), .fa_or0(csa_component25_fa1_or0));
  fa fa_csa_component25_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component25_fa2_xor1), .fa_or0(csa_component25_fa2_or0));
  fa fa_csa_component25_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component25_fa3_xor1), .fa_or0(csa_component25_fa3_or0));
  fa fa_csa_component25_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component25_fa4_xor1), .fa_or0(csa_component25_fa4_or0));
  fa fa_csa_component25_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component25_fa5_xor1), .fa_or0(csa_component25_fa5_or0));
  fa fa_csa_component25_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component25_fa6_xor1), .fa_or0(csa_component25_fa6_or0));
  fa fa_csa_component25_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component25_fa7_xor1), .fa_or0(csa_component25_fa7_or0));
  fa fa_csa_component25_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component25_fa8_xor1), .fa_or0(csa_component25_fa8_or0));
  fa fa_csa_component25_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component25_fa9_xor1), .fa_or0(csa_component25_fa9_or0));
  fa fa_csa_component25_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component25_fa10_xor1), .fa_or0(csa_component25_fa10_or0));
  fa fa_csa_component25_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component25_fa11_xor1), .fa_or0(csa_component25_fa11_or0));
  fa fa_csa_component25_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component25_fa12_xor1), .fa_or0(csa_component25_fa12_or0));
  fa fa_csa_component25_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component25_fa13_xor1), .fa_or0(csa_component25_fa13_or0));
  fa fa_csa_component25_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component25_fa14_xor1), .fa_or0(csa_component25_fa14_or0));
  fa fa_csa_component25_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component25_fa15_xor1), .fa_or0(csa_component25_fa15_or0));
  fa fa_csa_component25_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component25_fa16_xor1), .fa_or0(csa_component25_fa16_or0));
  fa fa_csa_component25_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component25_fa17_xor1), .fa_or0(csa_component25_fa17_or0));
  fa fa_csa_component25_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component25_fa18_xor1), .fa_or0(csa_component25_fa18_or0));
  fa fa_csa_component25_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component25_fa19_xor1), .fa_or0(csa_component25_fa19_or0));
  fa fa_csa_component25_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component25_fa20_xor1), .fa_or0(csa_component25_fa20_or0));
  fa fa_csa_component25_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component25_fa21_xor1), .fa_or0(csa_component25_fa21_or0));
  fa fa_csa_component25_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component25_fa22_xor1), .fa_or0(csa_component25_fa22_or0));
  fa fa_csa_component25_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component25_fa23_xor1), .fa_or0(csa_component25_fa23_or0));
  fa fa_csa_component25_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component25_fa24_xor1), .fa_or0(csa_component25_fa24_or0));

  assign csa_component25_out[0] = csa_component25_fa0_xor1[0];
  assign csa_component25_out[1] = csa_component25_fa1_xor1[0];
  assign csa_component25_out[2] = csa_component25_fa2_xor1[0];
  assign csa_component25_out[3] = csa_component25_fa3_xor1[0];
  assign csa_component25_out[4] = csa_component25_fa4_xor1[0];
  assign csa_component25_out[5] = csa_component25_fa5_xor1[0];
  assign csa_component25_out[6] = csa_component25_fa6_xor1[0];
  assign csa_component25_out[7] = csa_component25_fa7_xor1[0];
  assign csa_component25_out[8] = csa_component25_fa8_xor1[0];
  assign csa_component25_out[9] = csa_component25_fa9_xor1[0];
  assign csa_component25_out[10] = csa_component25_fa10_xor1[0];
  assign csa_component25_out[11] = csa_component25_fa11_xor1[0];
  assign csa_component25_out[12] = csa_component25_fa12_xor1[0];
  assign csa_component25_out[13] = csa_component25_fa13_xor1[0];
  assign csa_component25_out[14] = csa_component25_fa14_xor1[0];
  assign csa_component25_out[15] = csa_component25_fa15_xor1[0];
  assign csa_component25_out[16] = csa_component25_fa16_xor1[0];
  assign csa_component25_out[17] = csa_component25_fa17_xor1[0];
  assign csa_component25_out[18] = csa_component25_fa18_xor1[0];
  assign csa_component25_out[19] = csa_component25_fa19_xor1[0];
  assign csa_component25_out[20] = csa_component25_fa20_xor1[0];
  assign csa_component25_out[21] = csa_component25_fa21_xor1[0];
  assign csa_component25_out[22] = csa_component25_fa22_xor1[0];
  assign csa_component25_out[23] = csa_component25_fa23_xor1[0];
  assign csa_component25_out[24] = csa_component25_fa24_xor1[0];
  assign csa_component25_out[25] = 1'b0;
  assign csa_component25_out[26] = 1'b0;
  assign csa_component25_out[27] = csa_component25_fa0_or0[0];
  assign csa_component25_out[28] = csa_component25_fa1_or0[0];
  assign csa_component25_out[29] = csa_component25_fa2_or0[0];
  assign csa_component25_out[30] = csa_component25_fa3_or0[0];
  assign csa_component25_out[31] = csa_component25_fa4_or0[0];
  assign csa_component25_out[32] = csa_component25_fa5_or0[0];
  assign csa_component25_out[33] = csa_component25_fa6_or0[0];
  assign csa_component25_out[34] = csa_component25_fa7_or0[0];
  assign csa_component25_out[35] = csa_component25_fa8_or0[0];
  assign csa_component25_out[36] = csa_component25_fa9_or0[0];
  assign csa_component25_out[37] = csa_component25_fa10_or0[0];
  assign csa_component25_out[38] = csa_component25_fa11_or0[0];
  assign csa_component25_out[39] = csa_component25_fa12_or0[0];
  assign csa_component25_out[40] = csa_component25_fa13_or0[0];
  assign csa_component25_out[41] = csa_component25_fa14_or0[0];
  assign csa_component25_out[42] = csa_component25_fa15_or0[0];
  assign csa_component25_out[43] = csa_component25_fa16_or0[0];
  assign csa_component25_out[44] = csa_component25_fa17_or0[0];
  assign csa_component25_out[45] = csa_component25_fa18_or0[0];
  assign csa_component25_out[46] = csa_component25_fa19_or0[0];
  assign csa_component25_out[47] = csa_component25_fa20_or0[0];
  assign csa_component25_out[48] = csa_component25_fa21_or0[0];
  assign csa_component25_out[49] = csa_component25_fa22_or0[0];
  assign csa_component25_out[50] = csa_component25_fa23_or0[0];
  assign csa_component25_out[51] = csa_component25_fa24_or0[0];
endmodule

module csa_component31(input [30:0] a, input [30:0] b, input [30:0] c, output [63:0] csa_component31_out);
  wire [0:0] csa_component31_fa0_xor1;
  wire [0:0] csa_component31_fa0_or0;
  wire [0:0] csa_component31_fa1_xor1;
  wire [0:0] csa_component31_fa1_or0;
  wire [0:0] csa_component31_fa2_xor1;
  wire [0:0] csa_component31_fa2_or0;
  wire [0:0] csa_component31_fa3_xor1;
  wire [0:0] csa_component31_fa3_or0;
  wire [0:0] csa_component31_fa4_xor1;
  wire [0:0] csa_component31_fa4_or0;
  wire [0:0] csa_component31_fa5_xor1;
  wire [0:0] csa_component31_fa5_or0;
  wire [0:0] csa_component31_fa6_xor1;
  wire [0:0] csa_component31_fa6_or0;
  wire [0:0] csa_component31_fa7_xor1;
  wire [0:0] csa_component31_fa7_or0;
  wire [0:0] csa_component31_fa8_xor1;
  wire [0:0] csa_component31_fa8_or0;
  wire [0:0] csa_component31_fa9_xor1;
  wire [0:0] csa_component31_fa9_or0;
  wire [0:0] csa_component31_fa10_xor1;
  wire [0:0] csa_component31_fa10_or0;
  wire [0:0] csa_component31_fa11_xor1;
  wire [0:0] csa_component31_fa11_or0;
  wire [0:0] csa_component31_fa12_xor1;
  wire [0:0] csa_component31_fa12_or0;
  wire [0:0] csa_component31_fa13_xor1;
  wire [0:0] csa_component31_fa13_or0;
  wire [0:0] csa_component31_fa14_xor1;
  wire [0:0] csa_component31_fa14_or0;
  wire [0:0] csa_component31_fa15_xor1;
  wire [0:0] csa_component31_fa15_or0;
  wire [0:0] csa_component31_fa16_xor1;
  wire [0:0] csa_component31_fa16_or0;
  wire [0:0] csa_component31_fa17_xor1;
  wire [0:0] csa_component31_fa17_or0;
  wire [0:0] csa_component31_fa18_xor1;
  wire [0:0] csa_component31_fa18_or0;
  wire [0:0] csa_component31_fa19_xor1;
  wire [0:0] csa_component31_fa19_or0;
  wire [0:0] csa_component31_fa20_xor1;
  wire [0:0] csa_component31_fa20_or0;
  wire [0:0] csa_component31_fa21_xor1;
  wire [0:0] csa_component31_fa21_or0;
  wire [0:0] csa_component31_fa22_xor1;
  wire [0:0] csa_component31_fa22_or0;
  wire [0:0] csa_component31_fa23_xor1;
  wire [0:0] csa_component31_fa23_or0;
  wire [0:0] csa_component31_fa24_xor1;
  wire [0:0] csa_component31_fa24_or0;
  wire [0:0] csa_component31_fa25_xor1;
  wire [0:0] csa_component31_fa25_or0;
  wire [0:0] csa_component31_fa26_xor1;
  wire [0:0] csa_component31_fa26_or0;
  wire [0:0] csa_component31_fa27_xor1;
  wire [0:0] csa_component31_fa27_or0;
  wire [0:0] csa_component31_fa28_xor1;
  wire [0:0] csa_component31_fa28_or0;
  wire [0:0] csa_component31_fa29_xor1;
  wire [0:0] csa_component31_fa29_or0;
  wire [0:0] csa_component31_fa30_xor1;
  wire [0:0] csa_component31_fa30_or0;

  fa fa_csa_component31_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component31_fa0_xor1), .fa_or0(csa_component31_fa0_or0));
  fa fa_csa_component31_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component31_fa1_xor1), .fa_or0(csa_component31_fa1_or0));
  fa fa_csa_component31_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component31_fa2_xor1), .fa_or0(csa_component31_fa2_or0));
  fa fa_csa_component31_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component31_fa3_xor1), .fa_or0(csa_component31_fa3_or0));
  fa fa_csa_component31_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component31_fa4_xor1), .fa_or0(csa_component31_fa4_or0));
  fa fa_csa_component31_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component31_fa5_xor1), .fa_or0(csa_component31_fa5_or0));
  fa fa_csa_component31_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component31_fa6_xor1), .fa_or0(csa_component31_fa6_or0));
  fa fa_csa_component31_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component31_fa7_xor1), .fa_or0(csa_component31_fa7_or0));
  fa fa_csa_component31_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component31_fa8_xor1), .fa_or0(csa_component31_fa8_or0));
  fa fa_csa_component31_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component31_fa9_xor1), .fa_or0(csa_component31_fa9_or0));
  fa fa_csa_component31_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component31_fa10_xor1), .fa_or0(csa_component31_fa10_or0));
  fa fa_csa_component31_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component31_fa11_xor1), .fa_or0(csa_component31_fa11_or0));
  fa fa_csa_component31_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component31_fa12_xor1), .fa_or0(csa_component31_fa12_or0));
  fa fa_csa_component31_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component31_fa13_xor1), .fa_or0(csa_component31_fa13_or0));
  fa fa_csa_component31_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component31_fa14_xor1), .fa_or0(csa_component31_fa14_or0));
  fa fa_csa_component31_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component31_fa15_xor1), .fa_or0(csa_component31_fa15_or0));
  fa fa_csa_component31_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component31_fa16_xor1), .fa_or0(csa_component31_fa16_or0));
  fa fa_csa_component31_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component31_fa17_xor1), .fa_or0(csa_component31_fa17_or0));
  fa fa_csa_component31_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component31_fa18_xor1), .fa_or0(csa_component31_fa18_or0));
  fa fa_csa_component31_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component31_fa19_xor1), .fa_or0(csa_component31_fa19_or0));
  fa fa_csa_component31_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component31_fa20_xor1), .fa_or0(csa_component31_fa20_or0));
  fa fa_csa_component31_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component31_fa21_xor1), .fa_or0(csa_component31_fa21_or0));
  fa fa_csa_component31_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component31_fa22_xor1), .fa_or0(csa_component31_fa22_or0));
  fa fa_csa_component31_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component31_fa23_xor1), .fa_or0(csa_component31_fa23_or0));
  fa fa_csa_component31_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component31_fa24_xor1), .fa_or0(csa_component31_fa24_or0));
  fa fa_csa_component31_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component31_fa25_xor1), .fa_or0(csa_component31_fa25_or0));
  fa fa_csa_component31_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component31_fa26_xor1), .fa_or0(csa_component31_fa26_or0));
  fa fa_csa_component31_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component31_fa27_xor1), .fa_or0(csa_component31_fa27_or0));
  fa fa_csa_component31_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component31_fa28_xor1), .fa_or0(csa_component31_fa28_or0));
  fa fa_csa_component31_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component31_fa29_xor1), .fa_or0(csa_component31_fa29_or0));
  fa fa_csa_component31_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component31_fa30_xor1), .fa_or0(csa_component31_fa30_or0));

  assign csa_component31_out[0] = csa_component31_fa0_xor1[0];
  assign csa_component31_out[1] = csa_component31_fa1_xor1[0];
  assign csa_component31_out[2] = csa_component31_fa2_xor1[0];
  assign csa_component31_out[3] = csa_component31_fa3_xor1[0];
  assign csa_component31_out[4] = csa_component31_fa4_xor1[0];
  assign csa_component31_out[5] = csa_component31_fa5_xor1[0];
  assign csa_component31_out[6] = csa_component31_fa6_xor1[0];
  assign csa_component31_out[7] = csa_component31_fa7_xor1[0];
  assign csa_component31_out[8] = csa_component31_fa8_xor1[0];
  assign csa_component31_out[9] = csa_component31_fa9_xor1[0];
  assign csa_component31_out[10] = csa_component31_fa10_xor1[0];
  assign csa_component31_out[11] = csa_component31_fa11_xor1[0];
  assign csa_component31_out[12] = csa_component31_fa12_xor1[0];
  assign csa_component31_out[13] = csa_component31_fa13_xor1[0];
  assign csa_component31_out[14] = csa_component31_fa14_xor1[0];
  assign csa_component31_out[15] = csa_component31_fa15_xor1[0];
  assign csa_component31_out[16] = csa_component31_fa16_xor1[0];
  assign csa_component31_out[17] = csa_component31_fa17_xor1[0];
  assign csa_component31_out[18] = csa_component31_fa18_xor1[0];
  assign csa_component31_out[19] = csa_component31_fa19_xor1[0];
  assign csa_component31_out[20] = csa_component31_fa20_xor1[0];
  assign csa_component31_out[21] = csa_component31_fa21_xor1[0];
  assign csa_component31_out[22] = csa_component31_fa22_xor1[0];
  assign csa_component31_out[23] = csa_component31_fa23_xor1[0];
  assign csa_component31_out[24] = csa_component31_fa24_xor1[0];
  assign csa_component31_out[25] = csa_component31_fa25_xor1[0];
  assign csa_component31_out[26] = csa_component31_fa26_xor1[0];
  assign csa_component31_out[27] = csa_component31_fa27_xor1[0];
  assign csa_component31_out[28] = csa_component31_fa28_xor1[0];
  assign csa_component31_out[29] = csa_component31_fa29_xor1[0];
  assign csa_component31_out[30] = csa_component31_fa30_xor1[0];
  assign csa_component31_out[31] = 1'b0;
  assign csa_component31_out[32] = 1'b0;
  assign csa_component31_out[33] = csa_component31_fa0_or0[0];
  assign csa_component31_out[34] = csa_component31_fa1_or0[0];
  assign csa_component31_out[35] = csa_component31_fa2_or0[0];
  assign csa_component31_out[36] = csa_component31_fa3_or0[0];
  assign csa_component31_out[37] = csa_component31_fa4_or0[0];
  assign csa_component31_out[38] = csa_component31_fa5_or0[0];
  assign csa_component31_out[39] = csa_component31_fa6_or0[0];
  assign csa_component31_out[40] = csa_component31_fa7_or0[0];
  assign csa_component31_out[41] = csa_component31_fa8_or0[0];
  assign csa_component31_out[42] = csa_component31_fa9_or0[0];
  assign csa_component31_out[43] = csa_component31_fa10_or0[0];
  assign csa_component31_out[44] = csa_component31_fa11_or0[0];
  assign csa_component31_out[45] = csa_component31_fa12_or0[0];
  assign csa_component31_out[46] = csa_component31_fa13_or0[0];
  assign csa_component31_out[47] = csa_component31_fa14_or0[0];
  assign csa_component31_out[48] = csa_component31_fa15_or0[0];
  assign csa_component31_out[49] = csa_component31_fa16_or0[0];
  assign csa_component31_out[50] = csa_component31_fa17_or0[0];
  assign csa_component31_out[51] = csa_component31_fa18_or0[0];
  assign csa_component31_out[52] = csa_component31_fa19_or0[0];
  assign csa_component31_out[53] = csa_component31_fa20_or0[0];
  assign csa_component31_out[54] = csa_component31_fa21_or0[0];
  assign csa_component31_out[55] = csa_component31_fa22_or0[0];
  assign csa_component31_out[56] = csa_component31_fa23_or0[0];
  assign csa_component31_out[57] = csa_component31_fa24_or0[0];
  assign csa_component31_out[58] = csa_component31_fa25_or0[0];
  assign csa_component31_out[59] = csa_component31_fa26_or0[0];
  assign csa_component31_out[60] = csa_component31_fa27_or0[0];
  assign csa_component31_out[61] = csa_component31_fa28_or0[0];
  assign csa_component31_out[62] = csa_component31_fa29_or0[0];
  assign csa_component31_out[63] = csa_component31_fa30_or0[0];
endmodule

module csa_component26(input [25:0] a, input [25:0] b, input [25:0] c, output [53:0] csa_component26_out);
  wire [0:0] csa_component26_fa0_xor1;
  wire [0:0] csa_component26_fa0_or0;
  wire [0:0] csa_component26_fa1_xor1;
  wire [0:0] csa_component26_fa1_or0;
  wire [0:0] csa_component26_fa2_xor1;
  wire [0:0] csa_component26_fa2_or0;
  wire [0:0] csa_component26_fa3_xor1;
  wire [0:0] csa_component26_fa3_or0;
  wire [0:0] csa_component26_fa4_xor1;
  wire [0:0] csa_component26_fa4_or0;
  wire [0:0] csa_component26_fa5_xor1;
  wire [0:0] csa_component26_fa5_or0;
  wire [0:0] csa_component26_fa6_xor1;
  wire [0:0] csa_component26_fa6_or0;
  wire [0:0] csa_component26_fa7_xor1;
  wire [0:0] csa_component26_fa7_or0;
  wire [0:0] csa_component26_fa8_xor1;
  wire [0:0] csa_component26_fa8_or0;
  wire [0:0] csa_component26_fa9_xor1;
  wire [0:0] csa_component26_fa9_or0;
  wire [0:0] csa_component26_fa10_xor1;
  wire [0:0] csa_component26_fa10_or0;
  wire [0:0] csa_component26_fa11_xor1;
  wire [0:0] csa_component26_fa11_or0;
  wire [0:0] csa_component26_fa12_xor1;
  wire [0:0] csa_component26_fa12_or0;
  wire [0:0] csa_component26_fa13_xor1;
  wire [0:0] csa_component26_fa13_or0;
  wire [0:0] csa_component26_fa14_xor1;
  wire [0:0] csa_component26_fa14_or0;
  wire [0:0] csa_component26_fa15_xor1;
  wire [0:0] csa_component26_fa15_or0;
  wire [0:0] csa_component26_fa16_xor1;
  wire [0:0] csa_component26_fa16_or0;
  wire [0:0] csa_component26_fa17_xor1;
  wire [0:0] csa_component26_fa17_or0;
  wire [0:0] csa_component26_fa18_xor1;
  wire [0:0] csa_component26_fa18_or0;
  wire [0:0] csa_component26_fa19_xor1;
  wire [0:0] csa_component26_fa19_or0;
  wire [0:0] csa_component26_fa20_xor1;
  wire [0:0] csa_component26_fa20_or0;
  wire [0:0] csa_component26_fa21_xor1;
  wire [0:0] csa_component26_fa21_or0;
  wire [0:0] csa_component26_fa22_xor1;
  wire [0:0] csa_component26_fa22_or0;
  wire [0:0] csa_component26_fa23_xor1;
  wire [0:0] csa_component26_fa23_or0;
  wire [0:0] csa_component26_fa24_xor1;
  wire [0:0] csa_component26_fa24_or0;
  wire [0:0] csa_component26_fa25_xor1;
  wire [0:0] csa_component26_fa25_or0;

  fa fa_csa_component26_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component26_fa0_xor1), .fa_or0(csa_component26_fa0_or0));
  fa fa_csa_component26_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component26_fa1_xor1), .fa_or0(csa_component26_fa1_or0));
  fa fa_csa_component26_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component26_fa2_xor1), .fa_or0(csa_component26_fa2_or0));
  fa fa_csa_component26_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component26_fa3_xor1), .fa_or0(csa_component26_fa3_or0));
  fa fa_csa_component26_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component26_fa4_xor1), .fa_or0(csa_component26_fa4_or0));
  fa fa_csa_component26_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component26_fa5_xor1), .fa_or0(csa_component26_fa5_or0));
  fa fa_csa_component26_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component26_fa6_xor1), .fa_or0(csa_component26_fa6_or0));
  fa fa_csa_component26_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component26_fa7_xor1), .fa_or0(csa_component26_fa7_or0));
  fa fa_csa_component26_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component26_fa8_xor1), .fa_or0(csa_component26_fa8_or0));
  fa fa_csa_component26_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component26_fa9_xor1), .fa_or0(csa_component26_fa9_or0));
  fa fa_csa_component26_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component26_fa10_xor1), .fa_or0(csa_component26_fa10_or0));
  fa fa_csa_component26_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component26_fa11_xor1), .fa_or0(csa_component26_fa11_or0));
  fa fa_csa_component26_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component26_fa12_xor1), .fa_or0(csa_component26_fa12_or0));
  fa fa_csa_component26_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component26_fa13_xor1), .fa_or0(csa_component26_fa13_or0));
  fa fa_csa_component26_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component26_fa14_xor1), .fa_or0(csa_component26_fa14_or0));
  fa fa_csa_component26_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component26_fa15_xor1), .fa_or0(csa_component26_fa15_or0));
  fa fa_csa_component26_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component26_fa16_xor1), .fa_or0(csa_component26_fa16_or0));
  fa fa_csa_component26_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component26_fa17_xor1), .fa_or0(csa_component26_fa17_or0));
  fa fa_csa_component26_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component26_fa18_xor1), .fa_or0(csa_component26_fa18_or0));
  fa fa_csa_component26_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component26_fa19_xor1), .fa_or0(csa_component26_fa19_or0));
  fa fa_csa_component26_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component26_fa20_xor1), .fa_or0(csa_component26_fa20_or0));
  fa fa_csa_component26_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component26_fa21_xor1), .fa_or0(csa_component26_fa21_or0));
  fa fa_csa_component26_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component26_fa22_xor1), .fa_or0(csa_component26_fa22_or0));
  fa fa_csa_component26_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component26_fa23_xor1), .fa_or0(csa_component26_fa23_or0));
  fa fa_csa_component26_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component26_fa24_xor1), .fa_or0(csa_component26_fa24_or0));
  fa fa_csa_component26_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component26_fa25_xor1), .fa_or0(csa_component26_fa25_or0));

  assign csa_component26_out[0] = csa_component26_fa0_xor1[0];
  assign csa_component26_out[1] = csa_component26_fa1_xor1[0];
  assign csa_component26_out[2] = csa_component26_fa2_xor1[0];
  assign csa_component26_out[3] = csa_component26_fa3_xor1[0];
  assign csa_component26_out[4] = csa_component26_fa4_xor1[0];
  assign csa_component26_out[5] = csa_component26_fa5_xor1[0];
  assign csa_component26_out[6] = csa_component26_fa6_xor1[0];
  assign csa_component26_out[7] = csa_component26_fa7_xor1[0];
  assign csa_component26_out[8] = csa_component26_fa8_xor1[0];
  assign csa_component26_out[9] = csa_component26_fa9_xor1[0];
  assign csa_component26_out[10] = csa_component26_fa10_xor1[0];
  assign csa_component26_out[11] = csa_component26_fa11_xor1[0];
  assign csa_component26_out[12] = csa_component26_fa12_xor1[0];
  assign csa_component26_out[13] = csa_component26_fa13_xor1[0];
  assign csa_component26_out[14] = csa_component26_fa14_xor1[0];
  assign csa_component26_out[15] = csa_component26_fa15_xor1[0];
  assign csa_component26_out[16] = csa_component26_fa16_xor1[0];
  assign csa_component26_out[17] = csa_component26_fa17_xor1[0];
  assign csa_component26_out[18] = csa_component26_fa18_xor1[0];
  assign csa_component26_out[19] = csa_component26_fa19_xor1[0];
  assign csa_component26_out[20] = csa_component26_fa20_xor1[0];
  assign csa_component26_out[21] = csa_component26_fa21_xor1[0];
  assign csa_component26_out[22] = csa_component26_fa22_xor1[0];
  assign csa_component26_out[23] = csa_component26_fa23_xor1[0];
  assign csa_component26_out[24] = csa_component26_fa24_xor1[0];
  assign csa_component26_out[25] = csa_component26_fa25_xor1[0];
  assign csa_component26_out[26] = 1'b0;
  assign csa_component26_out[27] = 1'b0;
  assign csa_component26_out[28] = csa_component26_fa0_or0[0];
  assign csa_component26_out[29] = csa_component26_fa1_or0[0];
  assign csa_component26_out[30] = csa_component26_fa2_or0[0];
  assign csa_component26_out[31] = csa_component26_fa3_or0[0];
  assign csa_component26_out[32] = csa_component26_fa4_or0[0];
  assign csa_component26_out[33] = csa_component26_fa5_or0[0];
  assign csa_component26_out[34] = csa_component26_fa6_or0[0];
  assign csa_component26_out[35] = csa_component26_fa7_or0[0];
  assign csa_component26_out[36] = csa_component26_fa8_or0[0];
  assign csa_component26_out[37] = csa_component26_fa9_or0[0];
  assign csa_component26_out[38] = csa_component26_fa10_or0[0];
  assign csa_component26_out[39] = csa_component26_fa11_or0[0];
  assign csa_component26_out[40] = csa_component26_fa12_or0[0];
  assign csa_component26_out[41] = csa_component26_fa13_or0[0];
  assign csa_component26_out[42] = csa_component26_fa14_or0[0];
  assign csa_component26_out[43] = csa_component26_fa15_or0[0];
  assign csa_component26_out[44] = csa_component26_fa16_or0[0];
  assign csa_component26_out[45] = csa_component26_fa17_or0[0];
  assign csa_component26_out[46] = csa_component26_fa18_or0[0];
  assign csa_component26_out[47] = csa_component26_fa19_or0[0];
  assign csa_component26_out[48] = csa_component26_fa20_or0[0];
  assign csa_component26_out[49] = csa_component26_fa21_or0[0];
  assign csa_component26_out[50] = csa_component26_fa22_or0[0];
  assign csa_component26_out[51] = csa_component26_fa23_or0[0];
  assign csa_component26_out[52] = csa_component26_fa24_or0[0];
  assign csa_component26_out[53] = csa_component26_fa25_or0[0];
endmodule

module csa_component32(input [31:0] a, input [31:0] b, input [31:0] c, output [65:0] csa_component32_out);
  wire [0:0] csa_component32_fa0_xor1;
  wire [0:0] csa_component32_fa0_or0;
  wire [0:0] csa_component32_fa1_xor1;
  wire [0:0] csa_component32_fa1_or0;
  wire [0:0] csa_component32_fa2_xor1;
  wire [0:0] csa_component32_fa2_or0;
  wire [0:0] csa_component32_fa3_xor1;
  wire [0:0] csa_component32_fa3_or0;
  wire [0:0] csa_component32_fa4_xor1;
  wire [0:0] csa_component32_fa4_or0;
  wire [0:0] csa_component32_fa5_xor1;
  wire [0:0] csa_component32_fa5_or0;
  wire [0:0] csa_component32_fa6_xor1;
  wire [0:0] csa_component32_fa6_or0;
  wire [0:0] csa_component32_fa7_xor1;
  wire [0:0] csa_component32_fa7_or0;
  wire [0:0] csa_component32_fa8_xor1;
  wire [0:0] csa_component32_fa8_or0;
  wire [0:0] csa_component32_fa9_xor1;
  wire [0:0] csa_component32_fa9_or0;
  wire [0:0] csa_component32_fa10_xor1;
  wire [0:0] csa_component32_fa10_or0;
  wire [0:0] csa_component32_fa11_xor1;
  wire [0:0] csa_component32_fa11_or0;
  wire [0:0] csa_component32_fa12_xor1;
  wire [0:0] csa_component32_fa12_or0;
  wire [0:0] csa_component32_fa13_xor1;
  wire [0:0] csa_component32_fa13_or0;
  wire [0:0] csa_component32_fa14_xor1;
  wire [0:0] csa_component32_fa14_or0;
  wire [0:0] csa_component32_fa15_xor1;
  wire [0:0] csa_component32_fa15_or0;
  wire [0:0] csa_component32_fa16_xor1;
  wire [0:0] csa_component32_fa16_or0;
  wire [0:0] csa_component32_fa17_xor1;
  wire [0:0] csa_component32_fa17_or0;
  wire [0:0] csa_component32_fa18_xor1;
  wire [0:0] csa_component32_fa18_or0;
  wire [0:0] csa_component32_fa19_xor1;
  wire [0:0] csa_component32_fa19_or0;
  wire [0:0] csa_component32_fa20_xor1;
  wire [0:0] csa_component32_fa20_or0;
  wire [0:0] csa_component32_fa21_xor1;
  wire [0:0] csa_component32_fa21_or0;
  wire [0:0] csa_component32_fa22_xor1;
  wire [0:0] csa_component32_fa22_or0;
  wire [0:0] csa_component32_fa23_xor1;
  wire [0:0] csa_component32_fa23_or0;
  wire [0:0] csa_component32_fa24_xor1;
  wire [0:0] csa_component32_fa24_or0;
  wire [0:0] csa_component32_fa25_xor1;
  wire [0:0] csa_component32_fa25_or0;
  wire [0:0] csa_component32_fa26_xor1;
  wire [0:0] csa_component32_fa26_or0;
  wire [0:0] csa_component32_fa27_xor1;
  wire [0:0] csa_component32_fa27_or0;
  wire [0:0] csa_component32_fa28_xor1;
  wire [0:0] csa_component32_fa28_or0;
  wire [0:0] csa_component32_fa29_xor1;
  wire [0:0] csa_component32_fa29_or0;
  wire [0:0] csa_component32_fa30_xor1;
  wire [0:0] csa_component32_fa30_or0;
  wire [0:0] csa_component32_fa31_xor1;
  wire [0:0] csa_component32_fa31_or0;

  fa fa_csa_component32_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component32_fa0_xor1), .fa_or0(csa_component32_fa0_or0));
  fa fa_csa_component32_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component32_fa1_xor1), .fa_or0(csa_component32_fa1_or0));
  fa fa_csa_component32_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component32_fa2_xor1), .fa_or0(csa_component32_fa2_or0));
  fa fa_csa_component32_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component32_fa3_xor1), .fa_or0(csa_component32_fa3_or0));
  fa fa_csa_component32_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component32_fa4_xor1), .fa_or0(csa_component32_fa4_or0));
  fa fa_csa_component32_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component32_fa5_xor1), .fa_or0(csa_component32_fa5_or0));
  fa fa_csa_component32_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component32_fa6_xor1), .fa_or0(csa_component32_fa6_or0));
  fa fa_csa_component32_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component32_fa7_xor1), .fa_or0(csa_component32_fa7_or0));
  fa fa_csa_component32_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component32_fa8_xor1), .fa_or0(csa_component32_fa8_or0));
  fa fa_csa_component32_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component32_fa9_xor1), .fa_or0(csa_component32_fa9_or0));
  fa fa_csa_component32_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component32_fa10_xor1), .fa_or0(csa_component32_fa10_or0));
  fa fa_csa_component32_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component32_fa11_xor1), .fa_or0(csa_component32_fa11_or0));
  fa fa_csa_component32_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component32_fa12_xor1), .fa_or0(csa_component32_fa12_or0));
  fa fa_csa_component32_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component32_fa13_xor1), .fa_or0(csa_component32_fa13_or0));
  fa fa_csa_component32_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component32_fa14_xor1), .fa_or0(csa_component32_fa14_or0));
  fa fa_csa_component32_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component32_fa15_xor1), .fa_or0(csa_component32_fa15_or0));
  fa fa_csa_component32_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component32_fa16_xor1), .fa_or0(csa_component32_fa16_or0));
  fa fa_csa_component32_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component32_fa17_xor1), .fa_or0(csa_component32_fa17_or0));
  fa fa_csa_component32_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component32_fa18_xor1), .fa_or0(csa_component32_fa18_or0));
  fa fa_csa_component32_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component32_fa19_xor1), .fa_or0(csa_component32_fa19_or0));
  fa fa_csa_component32_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component32_fa20_xor1), .fa_or0(csa_component32_fa20_or0));
  fa fa_csa_component32_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component32_fa21_xor1), .fa_or0(csa_component32_fa21_or0));
  fa fa_csa_component32_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component32_fa22_xor1), .fa_or0(csa_component32_fa22_or0));
  fa fa_csa_component32_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component32_fa23_xor1), .fa_or0(csa_component32_fa23_or0));
  fa fa_csa_component32_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component32_fa24_xor1), .fa_or0(csa_component32_fa24_or0));
  fa fa_csa_component32_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component32_fa25_xor1), .fa_or0(csa_component32_fa25_or0));
  fa fa_csa_component32_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component32_fa26_xor1), .fa_or0(csa_component32_fa26_or0));
  fa fa_csa_component32_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component32_fa27_xor1), .fa_or0(csa_component32_fa27_or0));
  fa fa_csa_component32_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component32_fa28_xor1), .fa_or0(csa_component32_fa28_or0));
  fa fa_csa_component32_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component32_fa29_xor1), .fa_or0(csa_component32_fa29_or0));
  fa fa_csa_component32_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component32_fa30_xor1), .fa_or0(csa_component32_fa30_or0));
  fa fa_csa_component32_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component32_fa31_xor1), .fa_or0(csa_component32_fa31_or0));

  assign csa_component32_out[0] = csa_component32_fa0_xor1[0];
  assign csa_component32_out[1] = csa_component32_fa1_xor1[0];
  assign csa_component32_out[2] = csa_component32_fa2_xor1[0];
  assign csa_component32_out[3] = csa_component32_fa3_xor1[0];
  assign csa_component32_out[4] = csa_component32_fa4_xor1[0];
  assign csa_component32_out[5] = csa_component32_fa5_xor1[0];
  assign csa_component32_out[6] = csa_component32_fa6_xor1[0];
  assign csa_component32_out[7] = csa_component32_fa7_xor1[0];
  assign csa_component32_out[8] = csa_component32_fa8_xor1[0];
  assign csa_component32_out[9] = csa_component32_fa9_xor1[0];
  assign csa_component32_out[10] = csa_component32_fa10_xor1[0];
  assign csa_component32_out[11] = csa_component32_fa11_xor1[0];
  assign csa_component32_out[12] = csa_component32_fa12_xor1[0];
  assign csa_component32_out[13] = csa_component32_fa13_xor1[0];
  assign csa_component32_out[14] = csa_component32_fa14_xor1[0];
  assign csa_component32_out[15] = csa_component32_fa15_xor1[0];
  assign csa_component32_out[16] = csa_component32_fa16_xor1[0];
  assign csa_component32_out[17] = csa_component32_fa17_xor1[0];
  assign csa_component32_out[18] = csa_component32_fa18_xor1[0];
  assign csa_component32_out[19] = csa_component32_fa19_xor1[0];
  assign csa_component32_out[20] = csa_component32_fa20_xor1[0];
  assign csa_component32_out[21] = csa_component32_fa21_xor1[0];
  assign csa_component32_out[22] = csa_component32_fa22_xor1[0];
  assign csa_component32_out[23] = csa_component32_fa23_xor1[0];
  assign csa_component32_out[24] = csa_component32_fa24_xor1[0];
  assign csa_component32_out[25] = csa_component32_fa25_xor1[0];
  assign csa_component32_out[26] = csa_component32_fa26_xor1[0];
  assign csa_component32_out[27] = csa_component32_fa27_xor1[0];
  assign csa_component32_out[28] = csa_component32_fa28_xor1[0];
  assign csa_component32_out[29] = csa_component32_fa29_xor1[0];
  assign csa_component32_out[30] = csa_component32_fa30_xor1[0];
  assign csa_component32_out[31] = csa_component32_fa31_xor1[0];
  assign csa_component32_out[32] = 1'b0;
  assign csa_component32_out[33] = 1'b0;
  assign csa_component32_out[34] = csa_component32_fa0_or0[0];
  assign csa_component32_out[35] = csa_component32_fa1_or0[0];
  assign csa_component32_out[36] = csa_component32_fa2_or0[0];
  assign csa_component32_out[37] = csa_component32_fa3_or0[0];
  assign csa_component32_out[38] = csa_component32_fa4_or0[0];
  assign csa_component32_out[39] = csa_component32_fa5_or0[0];
  assign csa_component32_out[40] = csa_component32_fa6_or0[0];
  assign csa_component32_out[41] = csa_component32_fa7_or0[0];
  assign csa_component32_out[42] = csa_component32_fa8_or0[0];
  assign csa_component32_out[43] = csa_component32_fa9_or0[0];
  assign csa_component32_out[44] = csa_component32_fa10_or0[0];
  assign csa_component32_out[45] = csa_component32_fa11_or0[0];
  assign csa_component32_out[46] = csa_component32_fa12_or0[0];
  assign csa_component32_out[47] = csa_component32_fa13_or0[0];
  assign csa_component32_out[48] = csa_component32_fa14_or0[0];
  assign csa_component32_out[49] = csa_component32_fa15_or0[0];
  assign csa_component32_out[50] = csa_component32_fa16_or0[0];
  assign csa_component32_out[51] = csa_component32_fa17_or0[0];
  assign csa_component32_out[52] = csa_component32_fa18_or0[0];
  assign csa_component32_out[53] = csa_component32_fa19_or0[0];
  assign csa_component32_out[54] = csa_component32_fa20_or0[0];
  assign csa_component32_out[55] = csa_component32_fa21_or0[0];
  assign csa_component32_out[56] = csa_component32_fa22_or0[0];
  assign csa_component32_out[57] = csa_component32_fa23_or0[0];
  assign csa_component32_out[58] = csa_component32_fa24_or0[0];
  assign csa_component32_out[59] = csa_component32_fa25_or0[0];
  assign csa_component32_out[60] = csa_component32_fa26_or0[0];
  assign csa_component32_out[61] = csa_component32_fa27_or0[0];
  assign csa_component32_out[62] = csa_component32_fa28_or0[0];
  assign csa_component32_out[63] = csa_component32_fa29_or0[0];
  assign csa_component32_out[64] = csa_component32_fa30_or0[0];
  assign csa_component32_out[65] = csa_component32_fa31_or0[0];
endmodule

module u_pg_rca32(input [31:0] a, input [31:0] b, output [32:0] u_pg_rca32_out);
  wire [0:0] u_pg_rca32_pg_fa0_xor0;
  wire [0:0] u_pg_rca32_pg_fa0_and0;
  wire [0:0] u_pg_rca32_pg_fa1_xor0;
  wire [0:0] u_pg_rca32_pg_fa1_and0;
  wire [0:0] u_pg_rca32_pg_fa1_xor1;
  wire [0:0] u_pg_rca32_and1;
  wire [0:0] u_pg_rca32_or1;
  wire [0:0] u_pg_rca32_pg_fa2_xor0;
  wire [0:0] u_pg_rca32_pg_fa2_and0;
  wire [0:0] u_pg_rca32_pg_fa2_xor1;
  wire [0:0] u_pg_rca32_and2;
  wire [0:0] u_pg_rca32_or2;
  wire [0:0] u_pg_rca32_pg_fa3_xor0;
  wire [0:0] u_pg_rca32_pg_fa3_and0;
  wire [0:0] u_pg_rca32_pg_fa3_xor1;
  wire [0:0] u_pg_rca32_and3;
  wire [0:0] u_pg_rca32_or3;
  wire [0:0] u_pg_rca32_pg_fa4_xor0;
  wire [0:0] u_pg_rca32_pg_fa4_and0;
  wire [0:0] u_pg_rca32_pg_fa4_xor1;
  wire [0:0] u_pg_rca32_and4;
  wire [0:0] u_pg_rca32_or4;
  wire [0:0] u_pg_rca32_pg_fa5_xor0;
  wire [0:0] u_pg_rca32_pg_fa5_and0;
  wire [0:0] u_pg_rca32_pg_fa5_xor1;
  wire [0:0] u_pg_rca32_and5;
  wire [0:0] u_pg_rca32_or5;
  wire [0:0] u_pg_rca32_pg_fa6_xor0;
  wire [0:0] u_pg_rca32_pg_fa6_and0;
  wire [0:0] u_pg_rca32_pg_fa6_xor1;
  wire [0:0] u_pg_rca32_and6;
  wire [0:0] u_pg_rca32_or6;
  wire [0:0] u_pg_rca32_pg_fa7_xor0;
  wire [0:0] u_pg_rca32_pg_fa7_and0;
  wire [0:0] u_pg_rca32_pg_fa7_xor1;
  wire [0:0] u_pg_rca32_and7;
  wire [0:0] u_pg_rca32_or7;
  wire [0:0] u_pg_rca32_pg_fa8_xor0;
  wire [0:0] u_pg_rca32_pg_fa8_and0;
  wire [0:0] u_pg_rca32_pg_fa8_xor1;
  wire [0:0] u_pg_rca32_and8;
  wire [0:0] u_pg_rca32_or8;
  wire [0:0] u_pg_rca32_pg_fa9_xor0;
  wire [0:0] u_pg_rca32_pg_fa9_and0;
  wire [0:0] u_pg_rca32_pg_fa9_xor1;
  wire [0:0] u_pg_rca32_and9;
  wire [0:0] u_pg_rca32_or9;
  wire [0:0] u_pg_rca32_pg_fa10_xor0;
  wire [0:0] u_pg_rca32_pg_fa10_and0;
  wire [0:0] u_pg_rca32_pg_fa10_xor1;
  wire [0:0] u_pg_rca32_and10;
  wire [0:0] u_pg_rca32_or10;
  wire [0:0] u_pg_rca32_pg_fa11_xor0;
  wire [0:0] u_pg_rca32_pg_fa11_and0;
  wire [0:0] u_pg_rca32_pg_fa11_xor1;
  wire [0:0] u_pg_rca32_and11;
  wire [0:0] u_pg_rca32_or11;
  wire [0:0] u_pg_rca32_pg_fa12_xor0;
  wire [0:0] u_pg_rca32_pg_fa12_and0;
  wire [0:0] u_pg_rca32_pg_fa12_xor1;
  wire [0:0] u_pg_rca32_and12;
  wire [0:0] u_pg_rca32_or12;
  wire [0:0] u_pg_rca32_pg_fa13_xor0;
  wire [0:0] u_pg_rca32_pg_fa13_and0;
  wire [0:0] u_pg_rca32_pg_fa13_xor1;
  wire [0:0] u_pg_rca32_and13;
  wire [0:0] u_pg_rca32_or13;
  wire [0:0] u_pg_rca32_pg_fa14_xor0;
  wire [0:0] u_pg_rca32_pg_fa14_and0;
  wire [0:0] u_pg_rca32_pg_fa14_xor1;
  wire [0:0] u_pg_rca32_and14;
  wire [0:0] u_pg_rca32_or14;
  wire [0:0] u_pg_rca32_pg_fa15_xor0;
  wire [0:0] u_pg_rca32_pg_fa15_and0;
  wire [0:0] u_pg_rca32_pg_fa15_xor1;
  wire [0:0] u_pg_rca32_and15;
  wire [0:0] u_pg_rca32_or15;
  wire [0:0] u_pg_rca32_pg_fa16_xor0;
  wire [0:0] u_pg_rca32_pg_fa16_and0;
  wire [0:0] u_pg_rca32_pg_fa16_xor1;
  wire [0:0] u_pg_rca32_and16;
  wire [0:0] u_pg_rca32_or16;
  wire [0:0] u_pg_rca32_pg_fa17_xor0;
  wire [0:0] u_pg_rca32_pg_fa17_and0;
  wire [0:0] u_pg_rca32_pg_fa17_xor1;
  wire [0:0] u_pg_rca32_and17;
  wire [0:0] u_pg_rca32_or17;
  wire [0:0] u_pg_rca32_pg_fa18_xor0;
  wire [0:0] u_pg_rca32_pg_fa18_and0;
  wire [0:0] u_pg_rca32_pg_fa18_xor1;
  wire [0:0] u_pg_rca32_and18;
  wire [0:0] u_pg_rca32_or18;
  wire [0:0] u_pg_rca32_pg_fa19_xor0;
  wire [0:0] u_pg_rca32_pg_fa19_and0;
  wire [0:0] u_pg_rca32_pg_fa19_xor1;
  wire [0:0] u_pg_rca32_and19;
  wire [0:0] u_pg_rca32_or19;
  wire [0:0] u_pg_rca32_pg_fa20_xor0;
  wire [0:0] u_pg_rca32_pg_fa20_and0;
  wire [0:0] u_pg_rca32_pg_fa20_xor1;
  wire [0:0] u_pg_rca32_and20;
  wire [0:0] u_pg_rca32_or20;
  wire [0:0] u_pg_rca32_pg_fa21_xor0;
  wire [0:0] u_pg_rca32_pg_fa21_and0;
  wire [0:0] u_pg_rca32_pg_fa21_xor1;
  wire [0:0] u_pg_rca32_and21;
  wire [0:0] u_pg_rca32_or21;
  wire [0:0] u_pg_rca32_pg_fa22_xor0;
  wire [0:0] u_pg_rca32_pg_fa22_and0;
  wire [0:0] u_pg_rca32_pg_fa22_xor1;
  wire [0:0] u_pg_rca32_and22;
  wire [0:0] u_pg_rca32_or22;
  wire [0:0] u_pg_rca32_pg_fa23_xor0;
  wire [0:0] u_pg_rca32_pg_fa23_and0;
  wire [0:0] u_pg_rca32_pg_fa23_xor1;
  wire [0:0] u_pg_rca32_and23;
  wire [0:0] u_pg_rca32_or23;
  wire [0:0] u_pg_rca32_pg_fa24_xor0;
  wire [0:0] u_pg_rca32_pg_fa24_and0;
  wire [0:0] u_pg_rca32_pg_fa24_xor1;
  wire [0:0] u_pg_rca32_and24;
  wire [0:0] u_pg_rca32_or24;
  wire [0:0] u_pg_rca32_pg_fa25_xor0;
  wire [0:0] u_pg_rca32_pg_fa25_and0;
  wire [0:0] u_pg_rca32_pg_fa25_xor1;
  wire [0:0] u_pg_rca32_and25;
  wire [0:0] u_pg_rca32_or25;
  wire [0:0] u_pg_rca32_pg_fa26_xor0;
  wire [0:0] u_pg_rca32_pg_fa26_and0;
  wire [0:0] u_pg_rca32_pg_fa26_xor1;
  wire [0:0] u_pg_rca32_and26;
  wire [0:0] u_pg_rca32_or26;
  wire [0:0] u_pg_rca32_pg_fa27_xor0;
  wire [0:0] u_pg_rca32_pg_fa27_and0;
  wire [0:0] u_pg_rca32_pg_fa27_xor1;
  wire [0:0] u_pg_rca32_and27;
  wire [0:0] u_pg_rca32_or27;
  wire [0:0] u_pg_rca32_pg_fa28_xor0;
  wire [0:0] u_pg_rca32_pg_fa28_and0;
  wire [0:0] u_pg_rca32_pg_fa28_xor1;
  wire [0:0] u_pg_rca32_and28;
  wire [0:0] u_pg_rca32_or28;
  wire [0:0] u_pg_rca32_pg_fa29_xor0;
  wire [0:0] u_pg_rca32_pg_fa29_and0;
  wire [0:0] u_pg_rca32_pg_fa29_xor1;
  wire [0:0] u_pg_rca32_and29;
  wire [0:0] u_pg_rca32_or29;
  wire [0:0] u_pg_rca32_pg_fa30_xor0;
  wire [0:0] u_pg_rca32_pg_fa30_and0;
  wire [0:0] u_pg_rca32_pg_fa30_xor1;
  wire [0:0] u_pg_rca32_and30;
  wire [0:0] u_pg_rca32_or30;
  wire [0:0] u_pg_rca32_pg_fa31_xor0;
  wire [0:0] u_pg_rca32_pg_fa31_and0;
  wire [0:0] u_pg_rca32_pg_fa31_xor1;
  wire [0:0] u_pg_rca32_and31;
  wire [0:0] u_pg_rca32_or31;

  pg_fa pg_fa_u_pg_rca32_pg_fa0_out(.a(a[0]), .b(b[0]), .cin(1'b0), .pg_fa_xor0(u_pg_rca32_pg_fa0_xor0), .pg_fa_and0(u_pg_rca32_pg_fa0_and0), .pg_fa_xor1());
  pg_fa pg_fa_u_pg_rca32_pg_fa1_out(.a(a[1]), .b(b[1]), .cin(u_pg_rca32_pg_fa0_and0[0]), .pg_fa_xor0(u_pg_rca32_pg_fa1_xor0), .pg_fa_and0(u_pg_rca32_pg_fa1_and0), .pg_fa_xor1(u_pg_rca32_pg_fa1_xor1));
  and_gate and_gate_u_pg_rca32_and1(.a(u_pg_rca32_pg_fa0_and0[0]), .b(u_pg_rca32_pg_fa1_xor0[0]), .out(u_pg_rca32_and1));
  or_gate or_gate_u_pg_rca32_or1(.a(u_pg_rca32_and1[0]), .b(u_pg_rca32_pg_fa1_and0[0]), .out(u_pg_rca32_or1));
  pg_fa pg_fa_u_pg_rca32_pg_fa2_out(.a(a[2]), .b(b[2]), .cin(u_pg_rca32_or1[0]), .pg_fa_xor0(u_pg_rca32_pg_fa2_xor0), .pg_fa_and0(u_pg_rca32_pg_fa2_and0), .pg_fa_xor1(u_pg_rca32_pg_fa2_xor1));
  and_gate and_gate_u_pg_rca32_and2(.a(u_pg_rca32_or1[0]), .b(u_pg_rca32_pg_fa2_xor0[0]), .out(u_pg_rca32_and2));
  or_gate or_gate_u_pg_rca32_or2(.a(u_pg_rca32_and2[0]), .b(u_pg_rca32_pg_fa2_and0[0]), .out(u_pg_rca32_or2));
  pg_fa pg_fa_u_pg_rca32_pg_fa3_out(.a(a[3]), .b(b[3]), .cin(u_pg_rca32_or2[0]), .pg_fa_xor0(u_pg_rca32_pg_fa3_xor0), .pg_fa_and0(u_pg_rca32_pg_fa3_and0), .pg_fa_xor1(u_pg_rca32_pg_fa3_xor1));
  and_gate and_gate_u_pg_rca32_and3(.a(u_pg_rca32_or2[0]), .b(u_pg_rca32_pg_fa3_xor0[0]), .out(u_pg_rca32_and3));
  or_gate or_gate_u_pg_rca32_or3(.a(u_pg_rca32_and3[0]), .b(u_pg_rca32_pg_fa3_and0[0]), .out(u_pg_rca32_or3));
  pg_fa pg_fa_u_pg_rca32_pg_fa4_out(.a(a[4]), .b(b[4]), .cin(u_pg_rca32_or3[0]), .pg_fa_xor0(u_pg_rca32_pg_fa4_xor0), .pg_fa_and0(u_pg_rca32_pg_fa4_and0), .pg_fa_xor1(u_pg_rca32_pg_fa4_xor1));
  and_gate and_gate_u_pg_rca32_and4(.a(u_pg_rca32_or3[0]), .b(u_pg_rca32_pg_fa4_xor0[0]), .out(u_pg_rca32_and4));
  or_gate or_gate_u_pg_rca32_or4(.a(u_pg_rca32_and4[0]), .b(u_pg_rca32_pg_fa4_and0[0]), .out(u_pg_rca32_or4));
  pg_fa pg_fa_u_pg_rca32_pg_fa5_out(.a(a[5]), .b(b[5]), .cin(u_pg_rca32_or4[0]), .pg_fa_xor0(u_pg_rca32_pg_fa5_xor0), .pg_fa_and0(u_pg_rca32_pg_fa5_and0), .pg_fa_xor1(u_pg_rca32_pg_fa5_xor1));
  and_gate and_gate_u_pg_rca32_and5(.a(u_pg_rca32_or4[0]), .b(u_pg_rca32_pg_fa5_xor0[0]), .out(u_pg_rca32_and5));
  or_gate or_gate_u_pg_rca32_or5(.a(u_pg_rca32_and5[0]), .b(u_pg_rca32_pg_fa5_and0[0]), .out(u_pg_rca32_or5));
  pg_fa pg_fa_u_pg_rca32_pg_fa6_out(.a(a[6]), .b(b[6]), .cin(u_pg_rca32_or5[0]), .pg_fa_xor0(u_pg_rca32_pg_fa6_xor0), .pg_fa_and0(u_pg_rca32_pg_fa6_and0), .pg_fa_xor1(u_pg_rca32_pg_fa6_xor1));
  and_gate and_gate_u_pg_rca32_and6(.a(u_pg_rca32_or5[0]), .b(u_pg_rca32_pg_fa6_xor0[0]), .out(u_pg_rca32_and6));
  or_gate or_gate_u_pg_rca32_or6(.a(u_pg_rca32_and6[0]), .b(u_pg_rca32_pg_fa6_and0[0]), .out(u_pg_rca32_or6));
  pg_fa pg_fa_u_pg_rca32_pg_fa7_out(.a(a[7]), .b(b[7]), .cin(u_pg_rca32_or6[0]), .pg_fa_xor0(u_pg_rca32_pg_fa7_xor0), .pg_fa_and0(u_pg_rca32_pg_fa7_and0), .pg_fa_xor1(u_pg_rca32_pg_fa7_xor1));
  and_gate and_gate_u_pg_rca32_and7(.a(u_pg_rca32_or6[0]), .b(u_pg_rca32_pg_fa7_xor0[0]), .out(u_pg_rca32_and7));
  or_gate or_gate_u_pg_rca32_or7(.a(u_pg_rca32_and7[0]), .b(u_pg_rca32_pg_fa7_and0[0]), .out(u_pg_rca32_or7));
  pg_fa pg_fa_u_pg_rca32_pg_fa8_out(.a(a[8]), .b(b[8]), .cin(u_pg_rca32_or7[0]), .pg_fa_xor0(u_pg_rca32_pg_fa8_xor0), .pg_fa_and0(u_pg_rca32_pg_fa8_and0), .pg_fa_xor1(u_pg_rca32_pg_fa8_xor1));
  and_gate and_gate_u_pg_rca32_and8(.a(u_pg_rca32_or7[0]), .b(u_pg_rca32_pg_fa8_xor0[0]), .out(u_pg_rca32_and8));
  or_gate or_gate_u_pg_rca32_or8(.a(u_pg_rca32_and8[0]), .b(u_pg_rca32_pg_fa8_and0[0]), .out(u_pg_rca32_or8));
  pg_fa pg_fa_u_pg_rca32_pg_fa9_out(.a(a[9]), .b(b[9]), .cin(u_pg_rca32_or8[0]), .pg_fa_xor0(u_pg_rca32_pg_fa9_xor0), .pg_fa_and0(u_pg_rca32_pg_fa9_and0), .pg_fa_xor1(u_pg_rca32_pg_fa9_xor1));
  and_gate and_gate_u_pg_rca32_and9(.a(u_pg_rca32_or8[0]), .b(u_pg_rca32_pg_fa9_xor0[0]), .out(u_pg_rca32_and9));
  or_gate or_gate_u_pg_rca32_or9(.a(u_pg_rca32_and9[0]), .b(u_pg_rca32_pg_fa9_and0[0]), .out(u_pg_rca32_or9));
  pg_fa pg_fa_u_pg_rca32_pg_fa10_out(.a(a[10]), .b(b[10]), .cin(u_pg_rca32_or9[0]), .pg_fa_xor0(u_pg_rca32_pg_fa10_xor0), .pg_fa_and0(u_pg_rca32_pg_fa10_and0), .pg_fa_xor1(u_pg_rca32_pg_fa10_xor1));
  and_gate and_gate_u_pg_rca32_and10(.a(u_pg_rca32_or9[0]), .b(u_pg_rca32_pg_fa10_xor0[0]), .out(u_pg_rca32_and10));
  or_gate or_gate_u_pg_rca32_or10(.a(u_pg_rca32_and10[0]), .b(u_pg_rca32_pg_fa10_and0[0]), .out(u_pg_rca32_or10));
  pg_fa pg_fa_u_pg_rca32_pg_fa11_out(.a(a[11]), .b(b[11]), .cin(u_pg_rca32_or10[0]), .pg_fa_xor0(u_pg_rca32_pg_fa11_xor0), .pg_fa_and0(u_pg_rca32_pg_fa11_and0), .pg_fa_xor1(u_pg_rca32_pg_fa11_xor1));
  and_gate and_gate_u_pg_rca32_and11(.a(u_pg_rca32_or10[0]), .b(u_pg_rca32_pg_fa11_xor0[0]), .out(u_pg_rca32_and11));
  or_gate or_gate_u_pg_rca32_or11(.a(u_pg_rca32_and11[0]), .b(u_pg_rca32_pg_fa11_and0[0]), .out(u_pg_rca32_or11));
  pg_fa pg_fa_u_pg_rca32_pg_fa12_out(.a(a[12]), .b(b[12]), .cin(u_pg_rca32_or11[0]), .pg_fa_xor0(u_pg_rca32_pg_fa12_xor0), .pg_fa_and0(u_pg_rca32_pg_fa12_and0), .pg_fa_xor1(u_pg_rca32_pg_fa12_xor1));
  and_gate and_gate_u_pg_rca32_and12(.a(u_pg_rca32_or11[0]), .b(u_pg_rca32_pg_fa12_xor0[0]), .out(u_pg_rca32_and12));
  or_gate or_gate_u_pg_rca32_or12(.a(u_pg_rca32_and12[0]), .b(u_pg_rca32_pg_fa12_and0[0]), .out(u_pg_rca32_or12));
  pg_fa pg_fa_u_pg_rca32_pg_fa13_out(.a(a[13]), .b(b[13]), .cin(u_pg_rca32_or12[0]), .pg_fa_xor0(u_pg_rca32_pg_fa13_xor0), .pg_fa_and0(u_pg_rca32_pg_fa13_and0), .pg_fa_xor1(u_pg_rca32_pg_fa13_xor1));
  and_gate and_gate_u_pg_rca32_and13(.a(u_pg_rca32_or12[0]), .b(u_pg_rca32_pg_fa13_xor0[0]), .out(u_pg_rca32_and13));
  or_gate or_gate_u_pg_rca32_or13(.a(u_pg_rca32_and13[0]), .b(u_pg_rca32_pg_fa13_and0[0]), .out(u_pg_rca32_or13));
  pg_fa pg_fa_u_pg_rca32_pg_fa14_out(.a(a[14]), .b(b[14]), .cin(u_pg_rca32_or13[0]), .pg_fa_xor0(u_pg_rca32_pg_fa14_xor0), .pg_fa_and0(u_pg_rca32_pg_fa14_and0), .pg_fa_xor1(u_pg_rca32_pg_fa14_xor1));
  and_gate and_gate_u_pg_rca32_and14(.a(u_pg_rca32_or13[0]), .b(u_pg_rca32_pg_fa14_xor0[0]), .out(u_pg_rca32_and14));
  or_gate or_gate_u_pg_rca32_or14(.a(u_pg_rca32_and14[0]), .b(u_pg_rca32_pg_fa14_and0[0]), .out(u_pg_rca32_or14));
  pg_fa pg_fa_u_pg_rca32_pg_fa15_out(.a(a[15]), .b(b[15]), .cin(u_pg_rca32_or14[0]), .pg_fa_xor0(u_pg_rca32_pg_fa15_xor0), .pg_fa_and0(u_pg_rca32_pg_fa15_and0), .pg_fa_xor1(u_pg_rca32_pg_fa15_xor1));
  and_gate and_gate_u_pg_rca32_and15(.a(u_pg_rca32_or14[0]), .b(u_pg_rca32_pg_fa15_xor0[0]), .out(u_pg_rca32_and15));
  or_gate or_gate_u_pg_rca32_or15(.a(u_pg_rca32_and15[0]), .b(u_pg_rca32_pg_fa15_and0[0]), .out(u_pg_rca32_or15));
  pg_fa pg_fa_u_pg_rca32_pg_fa16_out(.a(a[16]), .b(b[16]), .cin(u_pg_rca32_or15[0]), .pg_fa_xor0(u_pg_rca32_pg_fa16_xor0), .pg_fa_and0(u_pg_rca32_pg_fa16_and0), .pg_fa_xor1(u_pg_rca32_pg_fa16_xor1));
  and_gate and_gate_u_pg_rca32_and16(.a(u_pg_rca32_or15[0]), .b(u_pg_rca32_pg_fa16_xor0[0]), .out(u_pg_rca32_and16));
  or_gate or_gate_u_pg_rca32_or16(.a(u_pg_rca32_and16[0]), .b(u_pg_rca32_pg_fa16_and0[0]), .out(u_pg_rca32_or16));
  pg_fa pg_fa_u_pg_rca32_pg_fa17_out(.a(a[17]), .b(b[17]), .cin(u_pg_rca32_or16[0]), .pg_fa_xor0(u_pg_rca32_pg_fa17_xor0), .pg_fa_and0(u_pg_rca32_pg_fa17_and0), .pg_fa_xor1(u_pg_rca32_pg_fa17_xor1));
  and_gate and_gate_u_pg_rca32_and17(.a(u_pg_rca32_or16[0]), .b(u_pg_rca32_pg_fa17_xor0[0]), .out(u_pg_rca32_and17));
  or_gate or_gate_u_pg_rca32_or17(.a(u_pg_rca32_and17[0]), .b(u_pg_rca32_pg_fa17_and0[0]), .out(u_pg_rca32_or17));
  pg_fa pg_fa_u_pg_rca32_pg_fa18_out(.a(a[18]), .b(b[18]), .cin(u_pg_rca32_or17[0]), .pg_fa_xor0(u_pg_rca32_pg_fa18_xor0), .pg_fa_and0(u_pg_rca32_pg_fa18_and0), .pg_fa_xor1(u_pg_rca32_pg_fa18_xor1));
  and_gate and_gate_u_pg_rca32_and18(.a(u_pg_rca32_or17[0]), .b(u_pg_rca32_pg_fa18_xor0[0]), .out(u_pg_rca32_and18));
  or_gate or_gate_u_pg_rca32_or18(.a(u_pg_rca32_and18[0]), .b(u_pg_rca32_pg_fa18_and0[0]), .out(u_pg_rca32_or18));
  pg_fa pg_fa_u_pg_rca32_pg_fa19_out(.a(a[19]), .b(b[19]), .cin(u_pg_rca32_or18[0]), .pg_fa_xor0(u_pg_rca32_pg_fa19_xor0), .pg_fa_and0(u_pg_rca32_pg_fa19_and0), .pg_fa_xor1(u_pg_rca32_pg_fa19_xor1));
  and_gate and_gate_u_pg_rca32_and19(.a(u_pg_rca32_or18[0]), .b(u_pg_rca32_pg_fa19_xor0[0]), .out(u_pg_rca32_and19));
  or_gate or_gate_u_pg_rca32_or19(.a(u_pg_rca32_and19[0]), .b(u_pg_rca32_pg_fa19_and0[0]), .out(u_pg_rca32_or19));
  pg_fa pg_fa_u_pg_rca32_pg_fa20_out(.a(a[20]), .b(b[20]), .cin(u_pg_rca32_or19[0]), .pg_fa_xor0(u_pg_rca32_pg_fa20_xor0), .pg_fa_and0(u_pg_rca32_pg_fa20_and0), .pg_fa_xor1(u_pg_rca32_pg_fa20_xor1));
  and_gate and_gate_u_pg_rca32_and20(.a(u_pg_rca32_or19[0]), .b(u_pg_rca32_pg_fa20_xor0[0]), .out(u_pg_rca32_and20));
  or_gate or_gate_u_pg_rca32_or20(.a(u_pg_rca32_and20[0]), .b(u_pg_rca32_pg_fa20_and0[0]), .out(u_pg_rca32_or20));
  pg_fa pg_fa_u_pg_rca32_pg_fa21_out(.a(a[21]), .b(b[21]), .cin(u_pg_rca32_or20[0]), .pg_fa_xor0(u_pg_rca32_pg_fa21_xor0), .pg_fa_and0(u_pg_rca32_pg_fa21_and0), .pg_fa_xor1(u_pg_rca32_pg_fa21_xor1));
  and_gate and_gate_u_pg_rca32_and21(.a(u_pg_rca32_or20[0]), .b(u_pg_rca32_pg_fa21_xor0[0]), .out(u_pg_rca32_and21));
  or_gate or_gate_u_pg_rca32_or21(.a(u_pg_rca32_and21[0]), .b(u_pg_rca32_pg_fa21_and0[0]), .out(u_pg_rca32_or21));
  pg_fa pg_fa_u_pg_rca32_pg_fa22_out(.a(a[22]), .b(b[22]), .cin(u_pg_rca32_or21[0]), .pg_fa_xor0(u_pg_rca32_pg_fa22_xor0), .pg_fa_and0(u_pg_rca32_pg_fa22_and0), .pg_fa_xor1(u_pg_rca32_pg_fa22_xor1));
  and_gate and_gate_u_pg_rca32_and22(.a(u_pg_rca32_or21[0]), .b(u_pg_rca32_pg_fa22_xor0[0]), .out(u_pg_rca32_and22));
  or_gate or_gate_u_pg_rca32_or22(.a(u_pg_rca32_and22[0]), .b(u_pg_rca32_pg_fa22_and0[0]), .out(u_pg_rca32_or22));
  pg_fa pg_fa_u_pg_rca32_pg_fa23_out(.a(a[23]), .b(b[23]), .cin(u_pg_rca32_or22[0]), .pg_fa_xor0(u_pg_rca32_pg_fa23_xor0), .pg_fa_and0(u_pg_rca32_pg_fa23_and0), .pg_fa_xor1(u_pg_rca32_pg_fa23_xor1));
  and_gate and_gate_u_pg_rca32_and23(.a(u_pg_rca32_or22[0]), .b(u_pg_rca32_pg_fa23_xor0[0]), .out(u_pg_rca32_and23));
  or_gate or_gate_u_pg_rca32_or23(.a(u_pg_rca32_and23[0]), .b(u_pg_rca32_pg_fa23_and0[0]), .out(u_pg_rca32_or23));
  pg_fa pg_fa_u_pg_rca32_pg_fa24_out(.a(a[24]), .b(b[24]), .cin(u_pg_rca32_or23[0]), .pg_fa_xor0(u_pg_rca32_pg_fa24_xor0), .pg_fa_and0(u_pg_rca32_pg_fa24_and0), .pg_fa_xor1(u_pg_rca32_pg_fa24_xor1));
  and_gate and_gate_u_pg_rca32_and24(.a(u_pg_rca32_or23[0]), .b(u_pg_rca32_pg_fa24_xor0[0]), .out(u_pg_rca32_and24));
  or_gate or_gate_u_pg_rca32_or24(.a(u_pg_rca32_and24[0]), .b(u_pg_rca32_pg_fa24_and0[0]), .out(u_pg_rca32_or24));
  pg_fa pg_fa_u_pg_rca32_pg_fa25_out(.a(a[25]), .b(b[25]), .cin(u_pg_rca32_or24[0]), .pg_fa_xor0(u_pg_rca32_pg_fa25_xor0), .pg_fa_and0(u_pg_rca32_pg_fa25_and0), .pg_fa_xor1(u_pg_rca32_pg_fa25_xor1));
  and_gate and_gate_u_pg_rca32_and25(.a(u_pg_rca32_or24[0]), .b(u_pg_rca32_pg_fa25_xor0[0]), .out(u_pg_rca32_and25));
  or_gate or_gate_u_pg_rca32_or25(.a(u_pg_rca32_and25[0]), .b(u_pg_rca32_pg_fa25_and0[0]), .out(u_pg_rca32_or25));
  pg_fa pg_fa_u_pg_rca32_pg_fa26_out(.a(a[26]), .b(b[26]), .cin(u_pg_rca32_or25[0]), .pg_fa_xor0(u_pg_rca32_pg_fa26_xor0), .pg_fa_and0(u_pg_rca32_pg_fa26_and0), .pg_fa_xor1(u_pg_rca32_pg_fa26_xor1));
  and_gate and_gate_u_pg_rca32_and26(.a(u_pg_rca32_or25[0]), .b(u_pg_rca32_pg_fa26_xor0[0]), .out(u_pg_rca32_and26));
  or_gate or_gate_u_pg_rca32_or26(.a(u_pg_rca32_and26[0]), .b(u_pg_rca32_pg_fa26_and0[0]), .out(u_pg_rca32_or26));
  pg_fa pg_fa_u_pg_rca32_pg_fa27_out(.a(a[27]), .b(b[27]), .cin(u_pg_rca32_or26[0]), .pg_fa_xor0(u_pg_rca32_pg_fa27_xor0), .pg_fa_and0(u_pg_rca32_pg_fa27_and0), .pg_fa_xor1(u_pg_rca32_pg_fa27_xor1));
  and_gate and_gate_u_pg_rca32_and27(.a(u_pg_rca32_or26[0]), .b(u_pg_rca32_pg_fa27_xor0[0]), .out(u_pg_rca32_and27));
  or_gate or_gate_u_pg_rca32_or27(.a(u_pg_rca32_and27[0]), .b(u_pg_rca32_pg_fa27_and0[0]), .out(u_pg_rca32_or27));
  pg_fa pg_fa_u_pg_rca32_pg_fa28_out(.a(a[28]), .b(b[28]), .cin(u_pg_rca32_or27[0]), .pg_fa_xor0(u_pg_rca32_pg_fa28_xor0), .pg_fa_and0(u_pg_rca32_pg_fa28_and0), .pg_fa_xor1(u_pg_rca32_pg_fa28_xor1));
  and_gate and_gate_u_pg_rca32_and28(.a(u_pg_rca32_or27[0]), .b(u_pg_rca32_pg_fa28_xor0[0]), .out(u_pg_rca32_and28));
  or_gate or_gate_u_pg_rca32_or28(.a(u_pg_rca32_and28[0]), .b(u_pg_rca32_pg_fa28_and0[0]), .out(u_pg_rca32_or28));
  pg_fa pg_fa_u_pg_rca32_pg_fa29_out(.a(a[29]), .b(b[29]), .cin(u_pg_rca32_or28[0]), .pg_fa_xor0(u_pg_rca32_pg_fa29_xor0), .pg_fa_and0(u_pg_rca32_pg_fa29_and0), .pg_fa_xor1(u_pg_rca32_pg_fa29_xor1));
  and_gate and_gate_u_pg_rca32_and29(.a(u_pg_rca32_or28[0]), .b(u_pg_rca32_pg_fa29_xor0[0]), .out(u_pg_rca32_and29));
  or_gate or_gate_u_pg_rca32_or29(.a(u_pg_rca32_and29[0]), .b(u_pg_rca32_pg_fa29_and0[0]), .out(u_pg_rca32_or29));
  pg_fa pg_fa_u_pg_rca32_pg_fa30_out(.a(a[30]), .b(b[30]), .cin(u_pg_rca32_or29[0]), .pg_fa_xor0(u_pg_rca32_pg_fa30_xor0), .pg_fa_and0(u_pg_rca32_pg_fa30_and0), .pg_fa_xor1(u_pg_rca32_pg_fa30_xor1));
  and_gate and_gate_u_pg_rca32_and30(.a(u_pg_rca32_or29[0]), .b(u_pg_rca32_pg_fa30_xor0[0]), .out(u_pg_rca32_and30));
  or_gate or_gate_u_pg_rca32_or30(.a(u_pg_rca32_and30[0]), .b(u_pg_rca32_pg_fa30_and0[0]), .out(u_pg_rca32_or30));
  pg_fa pg_fa_u_pg_rca32_pg_fa31_out(.a(a[31]), .b(b[31]), .cin(u_pg_rca32_or30[0]), .pg_fa_xor0(u_pg_rca32_pg_fa31_xor0), .pg_fa_and0(u_pg_rca32_pg_fa31_and0), .pg_fa_xor1(u_pg_rca32_pg_fa31_xor1));
  and_gate and_gate_u_pg_rca32_and31(.a(u_pg_rca32_or30[0]), .b(u_pg_rca32_pg_fa31_xor0[0]), .out(u_pg_rca32_and31));
  or_gate or_gate_u_pg_rca32_or31(.a(u_pg_rca32_and31[0]), .b(u_pg_rca32_pg_fa31_and0[0]), .out(u_pg_rca32_or31));

  assign u_pg_rca32_out[0] = u_pg_rca32_pg_fa0_xor0[0];
  assign u_pg_rca32_out[1] = u_pg_rca32_pg_fa1_xor1[0];
  assign u_pg_rca32_out[2] = u_pg_rca32_pg_fa2_xor1[0];
  assign u_pg_rca32_out[3] = u_pg_rca32_pg_fa3_xor1[0];
  assign u_pg_rca32_out[4] = u_pg_rca32_pg_fa4_xor1[0];
  assign u_pg_rca32_out[5] = u_pg_rca32_pg_fa5_xor1[0];
  assign u_pg_rca32_out[6] = u_pg_rca32_pg_fa6_xor1[0];
  assign u_pg_rca32_out[7] = u_pg_rca32_pg_fa7_xor1[0];
  assign u_pg_rca32_out[8] = u_pg_rca32_pg_fa8_xor1[0];
  assign u_pg_rca32_out[9] = u_pg_rca32_pg_fa9_xor1[0];
  assign u_pg_rca32_out[10] = u_pg_rca32_pg_fa10_xor1[0];
  assign u_pg_rca32_out[11] = u_pg_rca32_pg_fa11_xor1[0];
  assign u_pg_rca32_out[12] = u_pg_rca32_pg_fa12_xor1[0];
  assign u_pg_rca32_out[13] = u_pg_rca32_pg_fa13_xor1[0];
  assign u_pg_rca32_out[14] = u_pg_rca32_pg_fa14_xor1[0];
  assign u_pg_rca32_out[15] = u_pg_rca32_pg_fa15_xor1[0];
  assign u_pg_rca32_out[16] = u_pg_rca32_pg_fa16_xor1[0];
  assign u_pg_rca32_out[17] = u_pg_rca32_pg_fa17_xor1[0];
  assign u_pg_rca32_out[18] = u_pg_rca32_pg_fa18_xor1[0];
  assign u_pg_rca32_out[19] = u_pg_rca32_pg_fa19_xor1[0];
  assign u_pg_rca32_out[20] = u_pg_rca32_pg_fa20_xor1[0];
  assign u_pg_rca32_out[21] = u_pg_rca32_pg_fa21_xor1[0];
  assign u_pg_rca32_out[22] = u_pg_rca32_pg_fa22_xor1[0];
  assign u_pg_rca32_out[23] = u_pg_rca32_pg_fa23_xor1[0];
  assign u_pg_rca32_out[24] = u_pg_rca32_pg_fa24_xor1[0];
  assign u_pg_rca32_out[25] = u_pg_rca32_pg_fa25_xor1[0];
  assign u_pg_rca32_out[26] = u_pg_rca32_pg_fa26_xor1[0];
  assign u_pg_rca32_out[27] = u_pg_rca32_pg_fa27_xor1[0];
  assign u_pg_rca32_out[28] = u_pg_rca32_pg_fa28_xor1[0];
  assign u_pg_rca32_out[29] = u_pg_rca32_pg_fa29_xor1[0];
  assign u_pg_rca32_out[30] = u_pg_rca32_pg_fa30_xor1[0];
  assign u_pg_rca32_out[31] = u_pg_rca32_pg_fa31_xor1[0];
  assign u_pg_rca32_out[32] = u_pg_rca32_or31[0];
endmodule

module u_CSAwallace_pg_rca16(input [15:0] a, input [15:0] b, output [31:0] u_CSAwallace_pg_rca16_out);
  wire [0:0] u_CSAwallace_pg_rca16_and_0_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_0;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_1;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_2;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_3;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_4;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_5;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_6;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_7;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_8;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_9;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_10;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_11;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_12;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_13;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_14;
  wire [0:0] u_CSAwallace_pg_rca16_and_0_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_1_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_2_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_3_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_4_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_5_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_6_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_7_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_8_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_9_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_10_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_11_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_12_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_13_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_14_15;
  wire [0:0] u_CSAwallace_pg_rca16_and_15_15;
  wire [17:0] u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0;
  wire [17:0] u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1;
  wire [17:0] u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2;
  wire [37:0] u_CSAwallace_pg_rca16_csa0_csa_component_out;
  wire [20:0] u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3;
  wire [20:0] u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4;
  wire [20:0] u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5;
  wire [43:0] u_CSAwallace_pg_rca16_csa1_csa_component_out;
  wire [23:0] u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6;
  wire [23:0] u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7;
  wire [23:0] u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8;
  wire [49:0] u_CSAwallace_pg_rca16_csa2_csa_component_out;
  wire [26:0] u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9;
  wire [26:0] u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10;
  wire [26:0] u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11;
  wire [55:0] u_CSAwallace_pg_rca16_csa3_csa_component_out;
  wire [29:0] u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12;
  wire [29:0] u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13;
  wire [29:0] u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14;
  wire [61:0] u_CSAwallace_pg_rca16_csa4_csa_component_out;
  wire [21:0] u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1;
  wire [21:0] u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1;
  wire [21:0] u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2;
  wire [45:0] u_CSAwallace_pg_rca16_csa5_csa_component_out;
  wire [24:0] u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2;
  wire [24:0] u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3;
  wire [24:0] u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3;
  wire [51:0] u_CSAwallace_pg_rca16_csa6_csa_component_out;
  wire [30:0] u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4;
  wire [30:0] u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4;
  wire [30:0] u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5;
  wire [63:0] u_CSAwallace_pg_rca16_csa7_csa_component_out;
  wire [25:0] u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6;
  wire [25:0] u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6;
  wire [25:0] u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7;
  wire [53:0] u_CSAwallace_pg_rca16_csa8_csa_component_out;
  wire [31:0] u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7;
  wire [31:0] u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8;
  wire [31:0] u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8;
  wire [65:0] u_CSAwallace_pg_rca16_csa9_csa_component_out;
  wire [31:0] u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9;
  wire [31:0] u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9;
  wire [31:0] u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10;
  wire [65:0] u_CSAwallace_pg_rca16_csa10_csa_component_out;
  wire [31:0] u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10;
  wire [31:0] u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5;
  wire [31:0] u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15;
  wire [65:0] u_CSAwallace_pg_rca16_csa11_csa_component_out;
  wire [31:0] u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11;
  wire [31:0] u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11;
  wire [31:0] u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12;
  wire [65:0] u_CSAwallace_pg_rca16_csa12_csa_component_out;
  wire [31:0] u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13;
  wire [31:0] u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13;
  wire [31:0] u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12;
  wire [65:0] u_CSAwallace_pg_rca16_csa13_csa_component_out;
  wire [31:0] u_CSAwallace_pg_rca16_u_pg_rca32_a;
  wire [31:0] u_CSAwallace_pg_rca16_u_pg_rca32_b;
  wire [32:0] u_CSAwallace_pg_rca16_u_pg_rca32_out;

  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_0(.a(a[0]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_0_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_0(.a(a[1]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_1_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_0(.a(a[2]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_2_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_0(.a(a[3]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_3_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_0(.a(a[4]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_4_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_0(.a(a[5]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_5_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_0(.a(a[6]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_6_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_0(.a(a[7]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_7_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_0(.a(a[8]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_8_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_0(.a(a[9]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_9_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_0(.a(a[10]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_10_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_0(.a(a[11]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_11_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_0(.a(a[12]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_12_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_0(.a(a[13]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_13_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_0(.a(a[14]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_14_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_0(.a(a[15]), .b(b[0]), .out(u_CSAwallace_pg_rca16_and_15_0));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_1(.a(a[0]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_0_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_1(.a(a[1]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_1_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_1(.a(a[2]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_2_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_1(.a(a[3]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_3_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_1(.a(a[4]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_4_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_1(.a(a[5]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_5_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_1(.a(a[6]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_6_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_1(.a(a[7]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_7_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_1(.a(a[8]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_8_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_1(.a(a[9]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_9_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_1(.a(a[10]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_10_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_1(.a(a[11]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_11_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_1(.a(a[12]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_12_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_1(.a(a[13]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_13_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_1(.a(a[14]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_14_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_1(.a(a[15]), .b(b[1]), .out(u_CSAwallace_pg_rca16_and_15_1));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_2(.a(a[0]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_0_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_2(.a(a[1]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_1_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_2(.a(a[2]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_2_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_2(.a(a[3]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_3_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_2(.a(a[4]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_4_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_2(.a(a[5]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_5_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_2(.a(a[6]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_6_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_2(.a(a[7]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_7_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_2(.a(a[8]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_8_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_2(.a(a[9]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_9_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_2(.a(a[10]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_10_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_2(.a(a[11]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_11_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_2(.a(a[12]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_12_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_2(.a(a[13]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_13_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_2(.a(a[14]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_14_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_2(.a(a[15]), .b(b[2]), .out(u_CSAwallace_pg_rca16_and_15_2));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_3(.a(a[0]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_0_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_3(.a(a[1]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_1_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_3(.a(a[2]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_2_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_3(.a(a[3]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_3_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_3(.a(a[4]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_4_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_3(.a(a[5]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_5_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_3(.a(a[6]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_6_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_3(.a(a[7]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_7_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_3(.a(a[8]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_8_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_3(.a(a[9]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_9_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_3(.a(a[10]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_10_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_3(.a(a[11]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_11_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_3(.a(a[12]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_12_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_3(.a(a[13]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_13_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_3(.a(a[14]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_14_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_3(.a(a[15]), .b(b[3]), .out(u_CSAwallace_pg_rca16_and_15_3));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_4(.a(a[0]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_0_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_4(.a(a[1]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_1_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_4(.a(a[2]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_2_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_4(.a(a[3]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_3_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_4(.a(a[4]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_4_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_4(.a(a[5]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_5_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_4(.a(a[6]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_6_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_4(.a(a[7]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_7_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_4(.a(a[8]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_8_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_4(.a(a[9]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_9_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_4(.a(a[10]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_10_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_4(.a(a[11]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_11_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_4(.a(a[12]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_12_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_4(.a(a[13]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_13_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_4(.a(a[14]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_14_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_4(.a(a[15]), .b(b[4]), .out(u_CSAwallace_pg_rca16_and_15_4));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_5(.a(a[0]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_0_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_5(.a(a[1]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_1_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_5(.a(a[2]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_2_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_5(.a(a[3]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_3_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_5(.a(a[4]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_4_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_5(.a(a[5]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_5_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_5(.a(a[6]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_6_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_5(.a(a[7]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_7_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_5(.a(a[8]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_8_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_5(.a(a[9]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_9_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_5(.a(a[10]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_10_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_5(.a(a[11]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_11_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_5(.a(a[12]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_12_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_5(.a(a[13]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_13_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_5(.a(a[14]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_14_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_5(.a(a[15]), .b(b[5]), .out(u_CSAwallace_pg_rca16_and_15_5));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_6(.a(a[0]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_0_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_6(.a(a[1]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_1_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_6(.a(a[2]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_2_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_6(.a(a[3]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_3_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_6(.a(a[4]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_4_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_6(.a(a[5]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_5_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_6(.a(a[6]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_6_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_6(.a(a[7]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_7_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_6(.a(a[8]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_8_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_6(.a(a[9]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_9_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_6(.a(a[10]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_10_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_6(.a(a[11]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_11_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_6(.a(a[12]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_12_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_6(.a(a[13]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_13_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_6(.a(a[14]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_14_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_6(.a(a[15]), .b(b[6]), .out(u_CSAwallace_pg_rca16_and_15_6));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_7(.a(a[0]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_0_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_7(.a(a[1]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_1_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_7(.a(a[2]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_2_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_7(.a(a[3]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_3_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_7(.a(a[4]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_4_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_7(.a(a[5]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_5_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_7(.a(a[6]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_6_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_7(.a(a[7]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_7_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_7(.a(a[8]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_8_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_7(.a(a[9]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_9_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_7(.a(a[10]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_10_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_7(.a(a[11]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_11_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_7(.a(a[12]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_12_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_7(.a(a[13]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_13_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_7(.a(a[14]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_14_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_7(.a(a[15]), .b(b[7]), .out(u_CSAwallace_pg_rca16_and_15_7));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_8(.a(a[0]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_0_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_8(.a(a[1]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_1_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_8(.a(a[2]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_2_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_8(.a(a[3]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_3_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_8(.a(a[4]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_4_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_8(.a(a[5]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_5_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_8(.a(a[6]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_6_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_8(.a(a[7]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_7_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_8(.a(a[8]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_8_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_8(.a(a[9]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_9_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_8(.a(a[10]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_10_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_8(.a(a[11]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_11_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_8(.a(a[12]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_12_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_8(.a(a[13]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_13_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_8(.a(a[14]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_14_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_8(.a(a[15]), .b(b[8]), .out(u_CSAwallace_pg_rca16_and_15_8));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_9(.a(a[0]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_0_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_9(.a(a[1]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_1_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_9(.a(a[2]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_2_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_9(.a(a[3]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_3_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_9(.a(a[4]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_4_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_9(.a(a[5]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_5_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_9(.a(a[6]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_6_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_9(.a(a[7]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_7_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_9(.a(a[8]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_8_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_9(.a(a[9]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_9_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_9(.a(a[10]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_10_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_9(.a(a[11]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_11_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_9(.a(a[12]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_12_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_9(.a(a[13]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_13_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_9(.a(a[14]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_14_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_9(.a(a[15]), .b(b[9]), .out(u_CSAwallace_pg_rca16_and_15_9));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_10(.a(a[0]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_0_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_10(.a(a[1]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_1_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_10(.a(a[2]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_2_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_10(.a(a[3]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_3_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_10(.a(a[4]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_4_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_10(.a(a[5]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_5_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_10(.a(a[6]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_6_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_10(.a(a[7]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_7_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_10(.a(a[8]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_8_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_10(.a(a[9]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_9_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_10(.a(a[10]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_10_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_10(.a(a[11]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_11_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_10(.a(a[12]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_12_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_10(.a(a[13]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_13_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_10(.a(a[14]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_14_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_10(.a(a[15]), .b(b[10]), .out(u_CSAwallace_pg_rca16_and_15_10));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_11(.a(a[0]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_0_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_11(.a(a[1]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_1_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_11(.a(a[2]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_2_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_11(.a(a[3]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_3_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_11(.a(a[4]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_4_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_11(.a(a[5]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_5_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_11(.a(a[6]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_6_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_11(.a(a[7]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_7_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_11(.a(a[8]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_8_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_11(.a(a[9]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_9_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_11(.a(a[10]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_10_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_11(.a(a[11]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_11_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_11(.a(a[12]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_12_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_11(.a(a[13]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_13_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_11(.a(a[14]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_14_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_11(.a(a[15]), .b(b[11]), .out(u_CSAwallace_pg_rca16_and_15_11));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_12(.a(a[0]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_0_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_12(.a(a[1]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_1_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_12(.a(a[2]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_2_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_12(.a(a[3]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_3_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_12(.a(a[4]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_4_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_12(.a(a[5]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_5_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_12(.a(a[6]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_6_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_12(.a(a[7]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_7_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_12(.a(a[8]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_8_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_12(.a(a[9]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_9_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_12(.a(a[10]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_10_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_12(.a(a[11]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_11_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_12(.a(a[12]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_12_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_12(.a(a[13]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_13_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_12(.a(a[14]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_14_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_12(.a(a[15]), .b(b[12]), .out(u_CSAwallace_pg_rca16_and_15_12));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_13(.a(a[0]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_0_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_13(.a(a[1]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_1_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_13(.a(a[2]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_2_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_13(.a(a[3]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_3_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_13(.a(a[4]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_4_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_13(.a(a[5]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_5_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_13(.a(a[6]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_6_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_13(.a(a[7]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_7_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_13(.a(a[8]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_8_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_13(.a(a[9]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_9_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_13(.a(a[10]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_10_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_13(.a(a[11]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_11_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_13(.a(a[12]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_12_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_13(.a(a[13]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_13_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_13(.a(a[14]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_14_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_13(.a(a[15]), .b(b[13]), .out(u_CSAwallace_pg_rca16_and_15_13));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_14(.a(a[0]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_0_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_14(.a(a[1]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_1_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_14(.a(a[2]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_2_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_14(.a(a[3]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_3_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_14(.a(a[4]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_4_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_14(.a(a[5]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_5_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_14(.a(a[6]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_6_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_14(.a(a[7]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_7_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_14(.a(a[8]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_8_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_14(.a(a[9]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_9_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_14(.a(a[10]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_10_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_14(.a(a[11]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_11_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_14(.a(a[12]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_12_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_14(.a(a[13]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_13_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_14(.a(a[14]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_14_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_14(.a(a[15]), .b(b[14]), .out(u_CSAwallace_pg_rca16_and_15_14));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_0_15(.a(a[0]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_0_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_1_15(.a(a[1]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_1_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_2_15(.a(a[2]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_2_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_3_15(.a(a[3]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_3_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_4_15(.a(a[4]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_4_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_5_15(.a(a[5]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_5_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_6_15(.a(a[6]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_6_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_7_15(.a(a[7]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_7_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_8_15(.a(a[8]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_8_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_9_15(.a(a[9]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_9_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_10_15(.a(a[10]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_10_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_11_15(.a(a[11]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_11_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_12_15(.a(a[12]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_12_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_13_15(.a(a[13]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_13_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_14_15(.a(a[14]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_14_15));
  and_gate and_gate_u_CSAwallace_pg_rca16_and_15_15(.a(a[15]), .b(b[15]), .out(u_CSAwallace_pg_rca16_and_15_15));
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[0] = u_CSAwallace_pg_rca16_and_0_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[1] = u_CSAwallace_pg_rca16_and_1_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[2] = u_CSAwallace_pg_rca16_and_2_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[3] = u_CSAwallace_pg_rca16_and_3_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[4] = u_CSAwallace_pg_rca16_and_4_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[5] = u_CSAwallace_pg_rca16_and_5_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[6] = u_CSAwallace_pg_rca16_and_6_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[7] = u_CSAwallace_pg_rca16_and_7_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[8] = u_CSAwallace_pg_rca16_and_8_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[9] = u_CSAwallace_pg_rca16_and_9_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[10] = u_CSAwallace_pg_rca16_and_10_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[11] = u_CSAwallace_pg_rca16_and_11_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[12] = u_CSAwallace_pg_rca16_and_12_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[13] = u_CSAwallace_pg_rca16_and_13_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[14] = u_CSAwallace_pg_rca16_and_14_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[15] = u_CSAwallace_pg_rca16_and_15_0[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[16] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0[17] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[1] = u_CSAwallace_pg_rca16_and_0_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[2] = u_CSAwallace_pg_rca16_and_1_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[3] = u_CSAwallace_pg_rca16_and_2_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[4] = u_CSAwallace_pg_rca16_and_3_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[5] = u_CSAwallace_pg_rca16_and_4_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[6] = u_CSAwallace_pg_rca16_and_5_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[7] = u_CSAwallace_pg_rca16_and_6_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[8] = u_CSAwallace_pg_rca16_and_7_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[9] = u_CSAwallace_pg_rca16_and_8_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[10] = u_CSAwallace_pg_rca16_and_9_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[11] = u_CSAwallace_pg_rca16_and_10_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[12] = u_CSAwallace_pg_rca16_and_11_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[13] = u_CSAwallace_pg_rca16_and_12_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[14] = u_CSAwallace_pg_rca16_and_13_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[15] = u_CSAwallace_pg_rca16_and_14_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[16] = u_CSAwallace_pg_rca16_and_15_1[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1[17] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[2] = u_CSAwallace_pg_rca16_and_0_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[3] = u_CSAwallace_pg_rca16_and_1_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[4] = u_CSAwallace_pg_rca16_and_2_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[5] = u_CSAwallace_pg_rca16_and_3_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[6] = u_CSAwallace_pg_rca16_and_4_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[7] = u_CSAwallace_pg_rca16_and_5_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[8] = u_CSAwallace_pg_rca16_and_6_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[9] = u_CSAwallace_pg_rca16_and_7_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[10] = u_CSAwallace_pg_rca16_and_8_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[11] = u_CSAwallace_pg_rca16_and_9_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[12] = u_CSAwallace_pg_rca16_and_10_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[13] = u_CSAwallace_pg_rca16_and_11_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[14] = u_CSAwallace_pg_rca16_and_12_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[15] = u_CSAwallace_pg_rca16_and_13_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[16] = u_CSAwallace_pg_rca16_and_14_2[0];
  assign u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2[17] = u_CSAwallace_pg_rca16_and_15_2[0];
  csa_component18 csa_component18_u_CSAwallace_pg_rca16_csa0_csa_component_out(.a(u_CSAwallace_pg_rca16_csa0_csa_component_pp_row0), .b(u_CSAwallace_pg_rca16_csa0_csa_component_pp_row1), .c(u_CSAwallace_pg_rca16_csa0_csa_component_pp_row2), .csa_component18_out(u_CSAwallace_pg_rca16_csa0_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[3] = u_CSAwallace_pg_rca16_and_0_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[4] = u_CSAwallace_pg_rca16_and_1_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[5] = u_CSAwallace_pg_rca16_and_2_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[6] = u_CSAwallace_pg_rca16_and_3_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[7] = u_CSAwallace_pg_rca16_and_4_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[8] = u_CSAwallace_pg_rca16_and_5_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[9] = u_CSAwallace_pg_rca16_and_6_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[10] = u_CSAwallace_pg_rca16_and_7_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[11] = u_CSAwallace_pg_rca16_and_8_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[12] = u_CSAwallace_pg_rca16_and_9_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[13] = u_CSAwallace_pg_rca16_and_10_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[14] = u_CSAwallace_pg_rca16_and_11_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[15] = u_CSAwallace_pg_rca16_and_12_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[16] = u_CSAwallace_pg_rca16_and_13_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[17] = u_CSAwallace_pg_rca16_and_14_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[18] = u_CSAwallace_pg_rca16_and_15_3[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[19] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3[20] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[4] = u_CSAwallace_pg_rca16_and_0_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[5] = u_CSAwallace_pg_rca16_and_1_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[6] = u_CSAwallace_pg_rca16_and_2_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[7] = u_CSAwallace_pg_rca16_and_3_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[8] = u_CSAwallace_pg_rca16_and_4_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[9] = u_CSAwallace_pg_rca16_and_5_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[10] = u_CSAwallace_pg_rca16_and_6_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[11] = u_CSAwallace_pg_rca16_and_7_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[12] = u_CSAwallace_pg_rca16_and_8_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[13] = u_CSAwallace_pg_rca16_and_9_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[14] = u_CSAwallace_pg_rca16_and_10_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[15] = u_CSAwallace_pg_rca16_and_11_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[16] = u_CSAwallace_pg_rca16_and_12_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[17] = u_CSAwallace_pg_rca16_and_13_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[18] = u_CSAwallace_pg_rca16_and_14_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[19] = u_CSAwallace_pg_rca16_and_15_4[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4[20] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[5] = u_CSAwallace_pg_rca16_and_0_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[6] = u_CSAwallace_pg_rca16_and_1_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[7] = u_CSAwallace_pg_rca16_and_2_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[8] = u_CSAwallace_pg_rca16_and_3_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[9] = u_CSAwallace_pg_rca16_and_4_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[10] = u_CSAwallace_pg_rca16_and_5_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[11] = u_CSAwallace_pg_rca16_and_6_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[12] = u_CSAwallace_pg_rca16_and_7_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[13] = u_CSAwallace_pg_rca16_and_8_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[14] = u_CSAwallace_pg_rca16_and_9_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[15] = u_CSAwallace_pg_rca16_and_10_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[16] = u_CSAwallace_pg_rca16_and_11_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[17] = u_CSAwallace_pg_rca16_and_12_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[18] = u_CSAwallace_pg_rca16_and_13_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[19] = u_CSAwallace_pg_rca16_and_14_5[0];
  assign u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5[20] = u_CSAwallace_pg_rca16_and_15_5[0];
  csa_component21 csa_component21_u_CSAwallace_pg_rca16_csa1_csa_component_out(.a(u_CSAwallace_pg_rca16_csa1_csa_component_pp_row3), .b(u_CSAwallace_pg_rca16_csa1_csa_component_pp_row4), .c(u_CSAwallace_pg_rca16_csa1_csa_component_pp_row5), .csa_component21_out(u_CSAwallace_pg_rca16_csa1_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[6] = u_CSAwallace_pg_rca16_and_0_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[7] = u_CSAwallace_pg_rca16_and_1_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[8] = u_CSAwallace_pg_rca16_and_2_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[9] = u_CSAwallace_pg_rca16_and_3_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[10] = u_CSAwallace_pg_rca16_and_4_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[11] = u_CSAwallace_pg_rca16_and_5_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[12] = u_CSAwallace_pg_rca16_and_6_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[13] = u_CSAwallace_pg_rca16_and_7_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[14] = u_CSAwallace_pg_rca16_and_8_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[15] = u_CSAwallace_pg_rca16_and_9_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[16] = u_CSAwallace_pg_rca16_and_10_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[17] = u_CSAwallace_pg_rca16_and_11_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[18] = u_CSAwallace_pg_rca16_and_12_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[19] = u_CSAwallace_pg_rca16_and_13_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[20] = u_CSAwallace_pg_rca16_and_14_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[21] = u_CSAwallace_pg_rca16_and_15_6[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[22] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6[23] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[7] = u_CSAwallace_pg_rca16_and_0_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[8] = u_CSAwallace_pg_rca16_and_1_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[9] = u_CSAwallace_pg_rca16_and_2_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[10] = u_CSAwallace_pg_rca16_and_3_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[11] = u_CSAwallace_pg_rca16_and_4_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[12] = u_CSAwallace_pg_rca16_and_5_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[13] = u_CSAwallace_pg_rca16_and_6_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[14] = u_CSAwallace_pg_rca16_and_7_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[15] = u_CSAwallace_pg_rca16_and_8_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[16] = u_CSAwallace_pg_rca16_and_9_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[17] = u_CSAwallace_pg_rca16_and_10_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[18] = u_CSAwallace_pg_rca16_and_11_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[19] = u_CSAwallace_pg_rca16_and_12_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[20] = u_CSAwallace_pg_rca16_and_13_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[21] = u_CSAwallace_pg_rca16_and_14_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[22] = u_CSAwallace_pg_rca16_and_15_7[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7[23] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[8] = u_CSAwallace_pg_rca16_and_0_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[9] = u_CSAwallace_pg_rca16_and_1_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[10] = u_CSAwallace_pg_rca16_and_2_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[11] = u_CSAwallace_pg_rca16_and_3_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[12] = u_CSAwallace_pg_rca16_and_4_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[13] = u_CSAwallace_pg_rca16_and_5_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[14] = u_CSAwallace_pg_rca16_and_6_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[15] = u_CSAwallace_pg_rca16_and_7_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[16] = u_CSAwallace_pg_rca16_and_8_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[17] = u_CSAwallace_pg_rca16_and_9_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[18] = u_CSAwallace_pg_rca16_and_10_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[19] = u_CSAwallace_pg_rca16_and_11_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[20] = u_CSAwallace_pg_rca16_and_12_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[21] = u_CSAwallace_pg_rca16_and_13_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[22] = u_CSAwallace_pg_rca16_and_14_8[0];
  assign u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8[23] = u_CSAwallace_pg_rca16_and_15_8[0];
  csa_component24 csa_component24_u_CSAwallace_pg_rca16_csa2_csa_component_out(.a(u_CSAwallace_pg_rca16_csa2_csa_component_pp_row6), .b(u_CSAwallace_pg_rca16_csa2_csa_component_pp_row7), .c(u_CSAwallace_pg_rca16_csa2_csa_component_pp_row8), .csa_component24_out(u_CSAwallace_pg_rca16_csa2_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[9] = u_CSAwallace_pg_rca16_and_0_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[10] = u_CSAwallace_pg_rca16_and_1_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[11] = u_CSAwallace_pg_rca16_and_2_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[12] = u_CSAwallace_pg_rca16_and_3_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[13] = u_CSAwallace_pg_rca16_and_4_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[14] = u_CSAwallace_pg_rca16_and_5_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[15] = u_CSAwallace_pg_rca16_and_6_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[16] = u_CSAwallace_pg_rca16_and_7_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[17] = u_CSAwallace_pg_rca16_and_8_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[18] = u_CSAwallace_pg_rca16_and_9_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[19] = u_CSAwallace_pg_rca16_and_10_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[20] = u_CSAwallace_pg_rca16_and_11_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[21] = u_CSAwallace_pg_rca16_and_12_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[22] = u_CSAwallace_pg_rca16_and_13_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[23] = u_CSAwallace_pg_rca16_and_14_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[24] = u_CSAwallace_pg_rca16_and_15_9[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9[26] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[10] = u_CSAwallace_pg_rca16_and_0_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[11] = u_CSAwallace_pg_rca16_and_1_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[12] = u_CSAwallace_pg_rca16_and_2_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[13] = u_CSAwallace_pg_rca16_and_3_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[14] = u_CSAwallace_pg_rca16_and_4_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[15] = u_CSAwallace_pg_rca16_and_5_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[16] = u_CSAwallace_pg_rca16_and_6_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[17] = u_CSAwallace_pg_rca16_and_7_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[18] = u_CSAwallace_pg_rca16_and_8_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[19] = u_CSAwallace_pg_rca16_and_9_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[20] = u_CSAwallace_pg_rca16_and_10_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[21] = u_CSAwallace_pg_rca16_and_11_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[22] = u_CSAwallace_pg_rca16_and_12_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[23] = u_CSAwallace_pg_rca16_and_13_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[24] = u_CSAwallace_pg_rca16_and_14_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[25] = u_CSAwallace_pg_rca16_and_15_10[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10[26] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[11] = u_CSAwallace_pg_rca16_and_0_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[12] = u_CSAwallace_pg_rca16_and_1_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[13] = u_CSAwallace_pg_rca16_and_2_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[14] = u_CSAwallace_pg_rca16_and_3_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[15] = u_CSAwallace_pg_rca16_and_4_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[16] = u_CSAwallace_pg_rca16_and_5_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[17] = u_CSAwallace_pg_rca16_and_6_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[18] = u_CSAwallace_pg_rca16_and_7_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[19] = u_CSAwallace_pg_rca16_and_8_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[20] = u_CSAwallace_pg_rca16_and_9_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[21] = u_CSAwallace_pg_rca16_and_10_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[22] = u_CSAwallace_pg_rca16_and_11_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[23] = u_CSAwallace_pg_rca16_and_12_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[24] = u_CSAwallace_pg_rca16_and_13_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[25] = u_CSAwallace_pg_rca16_and_14_11[0];
  assign u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11[26] = u_CSAwallace_pg_rca16_and_15_11[0];
  csa_component27 csa_component27_u_CSAwallace_pg_rca16_csa3_csa_component_out(.a(u_CSAwallace_pg_rca16_csa3_csa_component_pp_row9), .b(u_CSAwallace_pg_rca16_csa3_csa_component_pp_row10), .c(u_CSAwallace_pg_rca16_csa3_csa_component_pp_row11), .csa_component27_out(u_CSAwallace_pg_rca16_csa3_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[12] = u_CSAwallace_pg_rca16_and_0_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[13] = u_CSAwallace_pg_rca16_and_1_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[14] = u_CSAwallace_pg_rca16_and_2_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[15] = u_CSAwallace_pg_rca16_and_3_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[16] = u_CSAwallace_pg_rca16_and_4_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[17] = u_CSAwallace_pg_rca16_and_5_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[18] = u_CSAwallace_pg_rca16_and_6_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[19] = u_CSAwallace_pg_rca16_and_7_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[20] = u_CSAwallace_pg_rca16_and_8_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[21] = u_CSAwallace_pg_rca16_and_9_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[22] = u_CSAwallace_pg_rca16_and_10_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[23] = u_CSAwallace_pg_rca16_and_11_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[24] = u_CSAwallace_pg_rca16_and_12_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[25] = u_CSAwallace_pg_rca16_and_13_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[26] = u_CSAwallace_pg_rca16_and_14_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[27] = u_CSAwallace_pg_rca16_and_15_12[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[12] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[13] = u_CSAwallace_pg_rca16_and_0_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[14] = u_CSAwallace_pg_rca16_and_1_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[15] = u_CSAwallace_pg_rca16_and_2_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[16] = u_CSAwallace_pg_rca16_and_3_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[17] = u_CSAwallace_pg_rca16_and_4_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[18] = u_CSAwallace_pg_rca16_and_5_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[19] = u_CSAwallace_pg_rca16_and_6_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[20] = u_CSAwallace_pg_rca16_and_7_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[21] = u_CSAwallace_pg_rca16_and_8_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[22] = u_CSAwallace_pg_rca16_and_9_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[23] = u_CSAwallace_pg_rca16_and_10_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[24] = u_CSAwallace_pg_rca16_and_11_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[25] = u_CSAwallace_pg_rca16_and_12_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[26] = u_CSAwallace_pg_rca16_and_13_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[27] = u_CSAwallace_pg_rca16_and_14_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[28] = u_CSAwallace_pg_rca16_and_15_13[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[12] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[13] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[14] = u_CSAwallace_pg_rca16_and_0_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[15] = u_CSAwallace_pg_rca16_and_1_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[16] = u_CSAwallace_pg_rca16_and_2_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[17] = u_CSAwallace_pg_rca16_and_3_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[18] = u_CSAwallace_pg_rca16_and_4_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[19] = u_CSAwallace_pg_rca16_and_5_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[20] = u_CSAwallace_pg_rca16_and_6_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[21] = u_CSAwallace_pg_rca16_and_7_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[22] = u_CSAwallace_pg_rca16_and_8_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[23] = u_CSAwallace_pg_rca16_and_9_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[24] = u_CSAwallace_pg_rca16_and_10_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[25] = u_CSAwallace_pg_rca16_and_11_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[26] = u_CSAwallace_pg_rca16_and_12_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[27] = u_CSAwallace_pg_rca16_and_13_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[28] = u_CSAwallace_pg_rca16_and_14_14[0];
  assign u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14[29] = u_CSAwallace_pg_rca16_and_15_14[0];
  csa_component30 csa_component30_u_CSAwallace_pg_rca16_csa4_csa_component_out(.a(u_CSAwallace_pg_rca16_csa4_csa_component_pp_row12), .b(u_CSAwallace_pg_rca16_csa4_csa_component_pp_row13), .c(u_CSAwallace_pg_rca16_csa4_csa_component_pp_row14), .csa_component30_out(u_CSAwallace_pg_rca16_csa4_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[0] = u_CSAwallace_pg_rca16_csa0_csa_component_out[0];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[1] = u_CSAwallace_pg_rca16_csa0_csa_component_out[1];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[2] = u_CSAwallace_pg_rca16_csa0_csa_component_out[2];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[3] = u_CSAwallace_pg_rca16_csa0_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[4] = u_CSAwallace_pg_rca16_csa0_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[5] = u_CSAwallace_pg_rca16_csa0_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[6] = u_CSAwallace_pg_rca16_csa0_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[7] = u_CSAwallace_pg_rca16_csa0_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[8] = u_CSAwallace_pg_rca16_csa0_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[9] = u_CSAwallace_pg_rca16_csa0_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[10] = u_CSAwallace_pg_rca16_csa0_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[11] = u_CSAwallace_pg_rca16_csa0_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[12] = u_CSAwallace_pg_rca16_csa0_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[13] = u_CSAwallace_pg_rca16_csa0_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[14] = u_CSAwallace_pg_rca16_csa0_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[15] = u_CSAwallace_pg_rca16_csa0_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[16] = u_CSAwallace_pg_rca16_csa0_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[17] = u_CSAwallace_pg_rca16_csa0_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[18] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[19] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[20] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1[21] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[2] = u_CSAwallace_pg_rca16_csa0_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[3] = u_CSAwallace_pg_rca16_csa0_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[4] = u_CSAwallace_pg_rca16_csa0_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[5] = u_CSAwallace_pg_rca16_csa0_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[6] = u_CSAwallace_pg_rca16_csa0_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[7] = u_CSAwallace_pg_rca16_csa0_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[8] = u_CSAwallace_pg_rca16_csa0_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[9] = u_CSAwallace_pg_rca16_csa0_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[10] = u_CSAwallace_pg_rca16_csa0_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[11] = u_CSAwallace_pg_rca16_csa0_csa_component_out[30];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[12] = u_CSAwallace_pg_rca16_csa0_csa_component_out[31];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[13] = u_CSAwallace_pg_rca16_csa0_csa_component_out[32];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[14] = u_CSAwallace_pg_rca16_csa0_csa_component_out[33];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[15] = u_CSAwallace_pg_rca16_csa0_csa_component_out[34];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[16] = u_CSAwallace_pg_rca16_csa0_csa_component_out[35];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[17] = u_CSAwallace_pg_rca16_csa0_csa_component_out[36];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[18] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[19] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[20] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1[21] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[3] = u_CSAwallace_pg_rca16_csa1_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[4] = u_CSAwallace_pg_rca16_csa1_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[5] = u_CSAwallace_pg_rca16_csa1_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[6] = u_CSAwallace_pg_rca16_csa1_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[7] = u_CSAwallace_pg_rca16_csa1_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[8] = u_CSAwallace_pg_rca16_csa1_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[9] = u_CSAwallace_pg_rca16_csa1_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[10] = u_CSAwallace_pg_rca16_csa1_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[11] = u_CSAwallace_pg_rca16_csa1_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[12] = u_CSAwallace_pg_rca16_csa1_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[13] = u_CSAwallace_pg_rca16_csa1_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[14] = u_CSAwallace_pg_rca16_csa1_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[15] = u_CSAwallace_pg_rca16_csa1_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[16] = u_CSAwallace_pg_rca16_csa1_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[17] = u_CSAwallace_pg_rca16_csa1_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[18] = u_CSAwallace_pg_rca16_csa1_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[19] = u_CSAwallace_pg_rca16_csa1_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[20] = u_CSAwallace_pg_rca16_csa1_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2[21] = 1'b0;
  csa_component22 csa_component22_u_CSAwallace_pg_rca16_csa5_csa_component_out(.a(u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s1), .b(u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_c1), .c(u_CSAwallace_pg_rca16_csa5_csa_component_u_CSAwallace_pg_rca16_csa_s2), .csa_component22_out(u_CSAwallace_pg_rca16_csa5_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[5] = u_CSAwallace_pg_rca16_csa1_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[6] = u_CSAwallace_pg_rca16_csa1_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[7] = u_CSAwallace_pg_rca16_csa1_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[8] = u_CSAwallace_pg_rca16_csa1_csa_component_out[30];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[9] = u_CSAwallace_pg_rca16_csa1_csa_component_out[31];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[10] = u_CSAwallace_pg_rca16_csa1_csa_component_out[32];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[11] = u_CSAwallace_pg_rca16_csa1_csa_component_out[33];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[12] = u_CSAwallace_pg_rca16_csa1_csa_component_out[34];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[13] = u_CSAwallace_pg_rca16_csa1_csa_component_out[35];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[14] = u_CSAwallace_pg_rca16_csa1_csa_component_out[36];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[15] = u_CSAwallace_pg_rca16_csa1_csa_component_out[37];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[16] = u_CSAwallace_pg_rca16_csa1_csa_component_out[38];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[17] = u_CSAwallace_pg_rca16_csa1_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[18] = u_CSAwallace_pg_rca16_csa1_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[19] = u_CSAwallace_pg_rca16_csa1_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[20] = u_CSAwallace_pg_rca16_csa1_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[21] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[22] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[23] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[6] = u_CSAwallace_pg_rca16_csa2_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[7] = u_CSAwallace_pg_rca16_csa2_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[8] = u_CSAwallace_pg_rca16_csa2_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[9] = u_CSAwallace_pg_rca16_csa2_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[10] = u_CSAwallace_pg_rca16_csa2_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[11] = u_CSAwallace_pg_rca16_csa2_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[12] = u_CSAwallace_pg_rca16_csa2_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[13] = u_CSAwallace_pg_rca16_csa2_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[14] = u_CSAwallace_pg_rca16_csa2_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[15] = u_CSAwallace_pg_rca16_csa2_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[16] = u_CSAwallace_pg_rca16_csa2_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[17] = u_CSAwallace_pg_rca16_csa2_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[18] = u_CSAwallace_pg_rca16_csa2_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[19] = u_CSAwallace_pg_rca16_csa2_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[20] = u_CSAwallace_pg_rca16_csa2_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[21] = u_CSAwallace_pg_rca16_csa2_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[22] = u_CSAwallace_pg_rca16_csa2_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[23] = u_CSAwallace_pg_rca16_csa2_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[8] = u_CSAwallace_pg_rca16_csa2_csa_component_out[33];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[9] = u_CSAwallace_pg_rca16_csa2_csa_component_out[34];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[10] = u_CSAwallace_pg_rca16_csa2_csa_component_out[35];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[11] = u_CSAwallace_pg_rca16_csa2_csa_component_out[36];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[12] = u_CSAwallace_pg_rca16_csa2_csa_component_out[37];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[13] = u_CSAwallace_pg_rca16_csa2_csa_component_out[38];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[14] = u_CSAwallace_pg_rca16_csa2_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[15] = u_CSAwallace_pg_rca16_csa2_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[16] = u_CSAwallace_pg_rca16_csa2_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[17] = u_CSAwallace_pg_rca16_csa2_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[18] = u_CSAwallace_pg_rca16_csa2_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[19] = u_CSAwallace_pg_rca16_csa2_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[20] = u_CSAwallace_pg_rca16_csa2_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[21] = u_CSAwallace_pg_rca16_csa2_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[22] = u_CSAwallace_pg_rca16_csa2_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[23] = u_CSAwallace_pg_rca16_csa2_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3[24] = 1'b0;
  csa_component25 csa_component25_u_CSAwallace_pg_rca16_csa6_csa_component_out(.a(u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c2), .b(u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_s3), .c(u_CSAwallace_pg_rca16_csa6_csa_component_u_CSAwallace_pg_rca16_csa_c3), .csa_component25_out(u_CSAwallace_pg_rca16_csa6_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[9] = u_CSAwallace_pg_rca16_csa3_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[10] = u_CSAwallace_pg_rca16_csa3_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[11] = u_CSAwallace_pg_rca16_csa3_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[12] = u_CSAwallace_pg_rca16_csa3_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[13] = u_CSAwallace_pg_rca16_csa3_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[14] = u_CSAwallace_pg_rca16_csa3_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[15] = u_CSAwallace_pg_rca16_csa3_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[16] = u_CSAwallace_pg_rca16_csa3_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[17] = u_CSAwallace_pg_rca16_csa3_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[18] = u_CSAwallace_pg_rca16_csa3_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[19] = u_CSAwallace_pg_rca16_csa3_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[20] = u_CSAwallace_pg_rca16_csa3_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[21] = u_CSAwallace_pg_rca16_csa3_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[22] = u_CSAwallace_pg_rca16_csa3_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[23] = u_CSAwallace_pg_rca16_csa3_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[24] = u_CSAwallace_pg_rca16_csa3_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[25] = u_CSAwallace_pg_rca16_csa3_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[26] = u_CSAwallace_pg_rca16_csa3_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[27] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[11] = u_CSAwallace_pg_rca16_csa3_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[12] = u_CSAwallace_pg_rca16_csa3_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[13] = u_CSAwallace_pg_rca16_csa3_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[14] = u_CSAwallace_pg_rca16_csa3_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[15] = u_CSAwallace_pg_rca16_csa3_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[16] = u_CSAwallace_pg_rca16_csa3_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[17] = u_CSAwallace_pg_rca16_csa3_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[18] = u_CSAwallace_pg_rca16_csa3_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[19] = u_CSAwallace_pg_rca16_csa3_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[20] = u_CSAwallace_pg_rca16_csa3_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[21] = u_CSAwallace_pg_rca16_csa3_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[22] = u_CSAwallace_pg_rca16_csa3_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[23] = u_CSAwallace_pg_rca16_csa3_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[24] = u_CSAwallace_pg_rca16_csa3_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[25] = u_CSAwallace_pg_rca16_csa3_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[26] = u_CSAwallace_pg_rca16_csa3_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[27] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[12] = u_CSAwallace_pg_rca16_csa4_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[13] = u_CSAwallace_pg_rca16_csa4_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[14] = u_CSAwallace_pg_rca16_csa4_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[15] = u_CSAwallace_pg_rca16_csa4_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[16] = u_CSAwallace_pg_rca16_csa4_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[17] = u_CSAwallace_pg_rca16_csa4_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[18] = u_CSAwallace_pg_rca16_csa4_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[19] = u_CSAwallace_pg_rca16_csa4_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[20] = u_CSAwallace_pg_rca16_csa4_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[21] = u_CSAwallace_pg_rca16_csa4_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[22] = u_CSAwallace_pg_rca16_csa4_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[23] = u_CSAwallace_pg_rca16_csa4_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[24] = u_CSAwallace_pg_rca16_csa4_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[25] = u_CSAwallace_pg_rca16_csa4_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[26] = u_CSAwallace_pg_rca16_csa4_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[27] = u_CSAwallace_pg_rca16_csa4_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[28] = u_CSAwallace_pg_rca16_csa4_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[29] = u_CSAwallace_pg_rca16_csa4_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5[30] = 1'b0;
  csa_component31 csa_component31_u_CSAwallace_pg_rca16_csa7_csa_component_out(.a(u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s4), .b(u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_c4), .c(u_CSAwallace_pg_rca16_csa7_csa_component_u_CSAwallace_pg_rca16_csa_s5), .csa_component31_out(u_CSAwallace_pg_rca16_csa7_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[0] = u_CSAwallace_pg_rca16_csa5_csa_component_out[0];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[1] = u_CSAwallace_pg_rca16_csa5_csa_component_out[1];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[2] = u_CSAwallace_pg_rca16_csa5_csa_component_out[2];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[3] = u_CSAwallace_pg_rca16_csa5_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[4] = u_CSAwallace_pg_rca16_csa5_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[5] = u_CSAwallace_pg_rca16_csa5_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[6] = u_CSAwallace_pg_rca16_csa5_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[7] = u_CSAwallace_pg_rca16_csa5_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[8] = u_CSAwallace_pg_rca16_csa5_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[9] = u_CSAwallace_pg_rca16_csa5_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[10] = u_CSAwallace_pg_rca16_csa5_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[11] = u_CSAwallace_pg_rca16_csa5_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[12] = u_CSAwallace_pg_rca16_csa5_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[13] = u_CSAwallace_pg_rca16_csa5_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[14] = u_CSAwallace_pg_rca16_csa5_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[15] = u_CSAwallace_pg_rca16_csa5_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[16] = u_CSAwallace_pg_rca16_csa5_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[17] = u_CSAwallace_pg_rca16_csa5_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[18] = u_CSAwallace_pg_rca16_csa5_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[19] = u_CSAwallace_pg_rca16_csa5_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[20] = u_CSAwallace_pg_rca16_csa5_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[21] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[22] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[23] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[3] = u_CSAwallace_pg_rca16_csa5_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[4] = u_CSAwallace_pg_rca16_csa5_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[5] = u_CSAwallace_pg_rca16_csa5_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[6] = u_CSAwallace_pg_rca16_csa5_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[7] = u_CSAwallace_pg_rca16_csa5_csa_component_out[30];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[8] = u_CSAwallace_pg_rca16_csa5_csa_component_out[31];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[9] = u_CSAwallace_pg_rca16_csa5_csa_component_out[32];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[10] = u_CSAwallace_pg_rca16_csa5_csa_component_out[33];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[11] = u_CSAwallace_pg_rca16_csa5_csa_component_out[34];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[12] = u_CSAwallace_pg_rca16_csa5_csa_component_out[35];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[13] = u_CSAwallace_pg_rca16_csa5_csa_component_out[36];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[14] = u_CSAwallace_pg_rca16_csa5_csa_component_out[37];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[15] = u_CSAwallace_pg_rca16_csa5_csa_component_out[38];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[16] = u_CSAwallace_pg_rca16_csa5_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[17] = u_CSAwallace_pg_rca16_csa5_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[18] = u_CSAwallace_pg_rca16_csa5_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[19] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[20] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[21] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[22] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[23] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[5] = u_CSAwallace_pg_rca16_csa6_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[6] = u_CSAwallace_pg_rca16_csa6_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[7] = u_CSAwallace_pg_rca16_csa6_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[8] = u_CSAwallace_pg_rca16_csa6_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[9] = u_CSAwallace_pg_rca16_csa6_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[10] = u_CSAwallace_pg_rca16_csa6_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[11] = u_CSAwallace_pg_rca16_csa6_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[12] = u_CSAwallace_pg_rca16_csa6_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[13] = u_CSAwallace_pg_rca16_csa6_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[14] = u_CSAwallace_pg_rca16_csa6_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[15] = u_CSAwallace_pg_rca16_csa6_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[16] = u_CSAwallace_pg_rca16_csa6_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[17] = u_CSAwallace_pg_rca16_csa6_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[18] = u_CSAwallace_pg_rca16_csa6_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[19] = u_CSAwallace_pg_rca16_csa6_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[20] = u_CSAwallace_pg_rca16_csa6_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[21] = u_CSAwallace_pg_rca16_csa6_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[22] = u_CSAwallace_pg_rca16_csa6_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[23] = u_CSAwallace_pg_rca16_csa6_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7[25] = 1'b0;
  csa_component26 csa_component26_u_CSAwallace_pg_rca16_csa8_csa_component_out(.a(u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s6), .b(u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_c6), .c(u_CSAwallace_pg_rca16_csa8_csa_component_u_CSAwallace_pg_rca16_csa_s7), .csa_component26_out(u_CSAwallace_pg_rca16_csa8_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[7] = u_CSAwallace_pg_rca16_csa6_csa_component_out[33];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[8] = u_CSAwallace_pg_rca16_csa6_csa_component_out[34];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[9] = u_CSAwallace_pg_rca16_csa6_csa_component_out[35];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[10] = u_CSAwallace_pg_rca16_csa6_csa_component_out[36];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[11] = u_CSAwallace_pg_rca16_csa6_csa_component_out[37];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[12] = u_CSAwallace_pg_rca16_csa6_csa_component_out[38];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[13] = u_CSAwallace_pg_rca16_csa6_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[14] = u_CSAwallace_pg_rca16_csa6_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[15] = u_CSAwallace_pg_rca16_csa6_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[16] = u_CSAwallace_pg_rca16_csa6_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[17] = u_CSAwallace_pg_rca16_csa6_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[18] = u_CSAwallace_pg_rca16_csa6_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[19] = u_CSAwallace_pg_rca16_csa6_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[20] = u_CSAwallace_pg_rca16_csa6_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[21] = u_CSAwallace_pg_rca16_csa6_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[22] = u_CSAwallace_pg_rca16_csa6_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[23] = u_CSAwallace_pg_rca16_csa6_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[24] = u_CSAwallace_pg_rca16_csa6_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[26] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[27] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[9] = u_CSAwallace_pg_rca16_csa7_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[10] = u_CSAwallace_pg_rca16_csa7_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[11] = u_CSAwallace_pg_rca16_csa7_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[12] = u_CSAwallace_pg_rca16_csa7_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[13] = u_CSAwallace_pg_rca16_csa7_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[14] = u_CSAwallace_pg_rca16_csa7_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[15] = u_CSAwallace_pg_rca16_csa7_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[16] = u_CSAwallace_pg_rca16_csa7_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[17] = u_CSAwallace_pg_rca16_csa7_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[18] = u_CSAwallace_pg_rca16_csa7_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[19] = u_CSAwallace_pg_rca16_csa7_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[20] = u_CSAwallace_pg_rca16_csa7_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[21] = u_CSAwallace_pg_rca16_csa7_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[22] = u_CSAwallace_pg_rca16_csa7_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[23] = u_CSAwallace_pg_rca16_csa7_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[24] = u_CSAwallace_pg_rca16_csa7_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[25] = u_CSAwallace_pg_rca16_csa7_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[26] = u_CSAwallace_pg_rca16_csa7_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[27] = u_CSAwallace_pg_rca16_csa7_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[28] = u_CSAwallace_pg_rca16_csa7_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[29] = u_CSAwallace_pg_rca16_csa7_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[12] = u_CSAwallace_pg_rca16_csa7_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[13] = u_CSAwallace_pg_rca16_csa7_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[14] = u_CSAwallace_pg_rca16_csa7_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[15] = u_CSAwallace_pg_rca16_csa7_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[16] = u_CSAwallace_pg_rca16_csa7_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[17] = u_CSAwallace_pg_rca16_csa7_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[18] = u_CSAwallace_pg_rca16_csa7_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[19] = u_CSAwallace_pg_rca16_csa7_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[20] = u_CSAwallace_pg_rca16_csa7_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[21] = u_CSAwallace_pg_rca16_csa7_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[22] = u_CSAwallace_pg_rca16_csa7_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[23] = u_CSAwallace_pg_rca16_csa7_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[24] = u_CSAwallace_pg_rca16_csa7_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[25] = u_CSAwallace_pg_rca16_csa7_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[26] = u_CSAwallace_pg_rca16_csa7_csa_component_out[58];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[27] = u_CSAwallace_pg_rca16_csa7_csa_component_out[59];
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8[31] = 1'b0;
  csa_component32 csa_component32_u_CSAwallace_pg_rca16_csa9_csa_component_out(.a(u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c7), .b(u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_s8), .c(u_CSAwallace_pg_rca16_csa9_csa_component_u_CSAwallace_pg_rca16_csa_c8), .csa_component32_out(u_CSAwallace_pg_rca16_csa9_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[0] = u_CSAwallace_pg_rca16_csa8_csa_component_out[0];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[1] = u_CSAwallace_pg_rca16_csa8_csa_component_out[1];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[2] = u_CSAwallace_pg_rca16_csa8_csa_component_out[2];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[3] = u_CSAwallace_pg_rca16_csa8_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[4] = u_CSAwallace_pg_rca16_csa8_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[5] = u_CSAwallace_pg_rca16_csa8_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[6] = u_CSAwallace_pg_rca16_csa8_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[7] = u_CSAwallace_pg_rca16_csa8_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[8] = u_CSAwallace_pg_rca16_csa8_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[9] = u_CSAwallace_pg_rca16_csa8_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[10] = u_CSAwallace_pg_rca16_csa8_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[11] = u_CSAwallace_pg_rca16_csa8_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[12] = u_CSAwallace_pg_rca16_csa8_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[13] = u_CSAwallace_pg_rca16_csa8_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[14] = u_CSAwallace_pg_rca16_csa8_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[15] = u_CSAwallace_pg_rca16_csa8_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[16] = u_CSAwallace_pg_rca16_csa8_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[17] = u_CSAwallace_pg_rca16_csa8_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[18] = u_CSAwallace_pg_rca16_csa8_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[19] = u_CSAwallace_pg_rca16_csa8_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[20] = u_CSAwallace_pg_rca16_csa8_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[21] = u_CSAwallace_pg_rca16_csa8_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[22] = u_CSAwallace_pg_rca16_csa8_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[23] = u_CSAwallace_pg_rca16_csa8_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[26] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[27] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[4] = u_CSAwallace_pg_rca16_csa8_csa_component_out[31];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[5] = u_CSAwallace_pg_rca16_csa8_csa_component_out[32];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[6] = u_CSAwallace_pg_rca16_csa8_csa_component_out[33];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[7] = u_CSAwallace_pg_rca16_csa8_csa_component_out[34];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[8] = u_CSAwallace_pg_rca16_csa8_csa_component_out[35];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[9] = u_CSAwallace_pg_rca16_csa8_csa_component_out[36];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[10] = u_CSAwallace_pg_rca16_csa8_csa_component_out[37];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[11] = u_CSAwallace_pg_rca16_csa8_csa_component_out[38];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[12] = u_CSAwallace_pg_rca16_csa8_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[13] = u_CSAwallace_pg_rca16_csa8_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[14] = u_CSAwallace_pg_rca16_csa8_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[15] = u_CSAwallace_pg_rca16_csa8_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[16] = u_CSAwallace_pg_rca16_csa8_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[17] = u_CSAwallace_pg_rca16_csa8_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[18] = u_CSAwallace_pg_rca16_csa8_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[19] = u_CSAwallace_pg_rca16_csa8_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[20] = u_CSAwallace_pg_rca16_csa8_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[21] = u_CSAwallace_pg_rca16_csa8_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[22] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[23] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[24] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[26] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[27] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[7] = u_CSAwallace_pg_rca16_csa9_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[8] = u_CSAwallace_pg_rca16_csa9_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[9] = u_CSAwallace_pg_rca16_csa9_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[10] = u_CSAwallace_pg_rca16_csa9_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[11] = u_CSAwallace_pg_rca16_csa9_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[12] = u_CSAwallace_pg_rca16_csa9_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[13] = u_CSAwallace_pg_rca16_csa9_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[14] = u_CSAwallace_pg_rca16_csa9_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[15] = u_CSAwallace_pg_rca16_csa9_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[16] = u_CSAwallace_pg_rca16_csa9_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[17] = u_CSAwallace_pg_rca16_csa9_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[18] = u_CSAwallace_pg_rca16_csa9_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[19] = u_CSAwallace_pg_rca16_csa9_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[20] = u_CSAwallace_pg_rca16_csa9_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[21] = u_CSAwallace_pg_rca16_csa9_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[22] = u_CSAwallace_pg_rca16_csa9_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[23] = u_CSAwallace_pg_rca16_csa9_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[24] = u_CSAwallace_pg_rca16_csa9_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[25] = u_CSAwallace_pg_rca16_csa9_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[26] = u_CSAwallace_pg_rca16_csa9_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[27] = u_CSAwallace_pg_rca16_csa9_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[28] = u_CSAwallace_pg_rca16_csa9_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[29] = u_CSAwallace_pg_rca16_csa9_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10[31] = 1'b0;
  csa_component32 csa_component32_u_CSAwallace_pg_rca16_csa10_csa_component_out(.a(u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s9), .b(u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_c9), .c(u_CSAwallace_pg_rca16_csa10_csa_component_u_CSAwallace_pg_rca16_csa_s10), .csa_component32_out(u_CSAwallace_pg_rca16_csa10_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[10] = u_CSAwallace_pg_rca16_csa9_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[11] = u_CSAwallace_pg_rca16_csa9_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[12] = u_CSAwallace_pg_rca16_csa9_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[13] = u_CSAwallace_pg_rca16_csa9_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[14] = u_CSAwallace_pg_rca16_csa9_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[15] = u_CSAwallace_pg_rca16_csa9_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[16] = u_CSAwallace_pg_rca16_csa9_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[17] = u_CSAwallace_pg_rca16_csa9_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[18] = u_CSAwallace_pg_rca16_csa9_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[19] = u_CSAwallace_pg_rca16_csa9_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[20] = u_CSAwallace_pg_rca16_csa9_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[21] = u_CSAwallace_pg_rca16_csa9_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[22] = u_CSAwallace_pg_rca16_csa9_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[23] = u_CSAwallace_pg_rca16_csa9_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[24] = u_CSAwallace_pg_rca16_csa9_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[25] = u_CSAwallace_pg_rca16_csa9_csa_component_out[58];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[26] = u_CSAwallace_pg_rca16_csa9_csa_component_out[59];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[27] = u_CSAwallace_pg_rca16_csa9_csa_component_out[60];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[28] = u_CSAwallace_pg_rca16_csa9_csa_component_out[61];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[12] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[13] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[14] = u_CSAwallace_pg_rca16_csa4_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[15] = u_CSAwallace_pg_rca16_csa4_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[16] = u_CSAwallace_pg_rca16_csa4_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[17] = u_CSAwallace_pg_rca16_csa4_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[18] = u_CSAwallace_pg_rca16_csa4_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[19] = u_CSAwallace_pg_rca16_csa4_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[20] = u_CSAwallace_pg_rca16_csa4_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[21] = u_CSAwallace_pg_rca16_csa4_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[22] = u_CSAwallace_pg_rca16_csa4_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[23] = u_CSAwallace_pg_rca16_csa4_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[24] = u_CSAwallace_pg_rca16_csa4_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[25] = u_CSAwallace_pg_rca16_csa4_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[26] = u_CSAwallace_pg_rca16_csa4_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[27] = u_CSAwallace_pg_rca16_csa4_csa_component_out[58];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[28] = u_CSAwallace_pg_rca16_csa4_csa_component_out[59];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[29] = u_CSAwallace_pg_rca16_csa4_csa_component_out[60];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[12] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[13] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[14] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[15] = u_CSAwallace_pg_rca16_and_0_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[16] = u_CSAwallace_pg_rca16_and_1_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[17] = u_CSAwallace_pg_rca16_and_2_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[18] = u_CSAwallace_pg_rca16_and_3_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[19] = u_CSAwallace_pg_rca16_and_4_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[20] = u_CSAwallace_pg_rca16_and_5_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[21] = u_CSAwallace_pg_rca16_and_6_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[22] = u_CSAwallace_pg_rca16_and_7_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[23] = u_CSAwallace_pg_rca16_and_8_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[24] = u_CSAwallace_pg_rca16_and_9_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[25] = u_CSAwallace_pg_rca16_and_10_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[26] = u_CSAwallace_pg_rca16_and_11_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[27] = u_CSAwallace_pg_rca16_and_12_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[28] = u_CSAwallace_pg_rca16_and_13_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[29] = u_CSAwallace_pg_rca16_and_14_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[30] = u_CSAwallace_pg_rca16_and_15_15[0];
  assign u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15[31] = 1'b0;
  csa_component32 csa_component32_u_CSAwallace_pg_rca16_csa11_csa_component_out(.a(u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c10), .b(u_CSAwallace_pg_rca16_csa11_csa_component_u_CSAwallace_pg_rca16_csa_c5), .c(u_CSAwallace_pg_rca16_csa11_csa_component_pp_row15), .csa_component32_out(u_CSAwallace_pg_rca16_csa11_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[0] = u_CSAwallace_pg_rca16_csa10_csa_component_out[0];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[1] = u_CSAwallace_pg_rca16_csa10_csa_component_out[1];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[2] = u_CSAwallace_pg_rca16_csa10_csa_component_out[2];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[3] = u_CSAwallace_pg_rca16_csa10_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[4] = u_CSAwallace_pg_rca16_csa10_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[5] = u_CSAwallace_pg_rca16_csa10_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[6] = u_CSAwallace_pg_rca16_csa10_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[7] = u_CSAwallace_pg_rca16_csa10_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[8] = u_CSAwallace_pg_rca16_csa10_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[9] = u_CSAwallace_pg_rca16_csa10_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[10] = u_CSAwallace_pg_rca16_csa10_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[11] = u_CSAwallace_pg_rca16_csa10_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[12] = u_CSAwallace_pg_rca16_csa10_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[13] = u_CSAwallace_pg_rca16_csa10_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[14] = u_CSAwallace_pg_rca16_csa10_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[15] = u_CSAwallace_pg_rca16_csa10_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[16] = u_CSAwallace_pg_rca16_csa10_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[17] = u_CSAwallace_pg_rca16_csa10_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[18] = u_CSAwallace_pg_rca16_csa10_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[19] = u_CSAwallace_pg_rca16_csa10_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[20] = u_CSAwallace_pg_rca16_csa10_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[21] = u_CSAwallace_pg_rca16_csa10_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[22] = u_CSAwallace_pg_rca16_csa10_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[23] = u_CSAwallace_pg_rca16_csa10_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[24] = u_CSAwallace_pg_rca16_csa10_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[25] = u_CSAwallace_pg_rca16_csa10_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[26] = u_CSAwallace_pg_rca16_csa10_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[27] = u_CSAwallace_pg_rca16_csa10_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[28] = u_CSAwallace_pg_rca16_csa10_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[29] = u_CSAwallace_pg_rca16_csa10_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[5] = u_CSAwallace_pg_rca16_csa10_csa_component_out[38];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[6] = u_CSAwallace_pg_rca16_csa10_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[7] = u_CSAwallace_pg_rca16_csa10_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[8] = u_CSAwallace_pg_rca16_csa10_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[9] = u_CSAwallace_pg_rca16_csa10_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[10] = u_CSAwallace_pg_rca16_csa10_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[11] = u_CSAwallace_pg_rca16_csa10_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[12] = u_CSAwallace_pg_rca16_csa10_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[13] = u_CSAwallace_pg_rca16_csa10_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[14] = u_CSAwallace_pg_rca16_csa10_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[15] = u_CSAwallace_pg_rca16_csa10_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[16] = u_CSAwallace_pg_rca16_csa10_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[17] = u_CSAwallace_pg_rca16_csa10_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[18] = u_CSAwallace_pg_rca16_csa10_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[19] = u_CSAwallace_pg_rca16_csa10_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[20] = u_CSAwallace_pg_rca16_csa10_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[21] = u_CSAwallace_pg_rca16_csa10_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[22] = u_CSAwallace_pg_rca16_csa10_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[23] = u_CSAwallace_pg_rca16_csa10_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[24] = u_CSAwallace_pg_rca16_csa10_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[25] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[26] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[27] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[28] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[29] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[30] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[10] = u_CSAwallace_pg_rca16_csa11_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[11] = u_CSAwallace_pg_rca16_csa11_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[12] = u_CSAwallace_pg_rca16_csa11_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[13] = u_CSAwallace_pg_rca16_csa11_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[14] = u_CSAwallace_pg_rca16_csa11_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[15] = u_CSAwallace_pg_rca16_csa11_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[16] = u_CSAwallace_pg_rca16_csa11_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[17] = u_CSAwallace_pg_rca16_csa11_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[18] = u_CSAwallace_pg_rca16_csa11_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[19] = u_CSAwallace_pg_rca16_csa11_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[20] = u_CSAwallace_pg_rca16_csa11_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[21] = u_CSAwallace_pg_rca16_csa11_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[22] = u_CSAwallace_pg_rca16_csa11_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[23] = u_CSAwallace_pg_rca16_csa11_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[24] = u_CSAwallace_pg_rca16_csa11_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[25] = u_CSAwallace_pg_rca16_csa11_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[26] = u_CSAwallace_pg_rca16_csa11_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[27] = u_CSAwallace_pg_rca16_csa11_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[28] = u_CSAwallace_pg_rca16_csa11_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[29] = u_CSAwallace_pg_rca16_csa11_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[30] = u_CSAwallace_pg_rca16_csa11_csa_component_out[30];
  assign u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12[31] = 1'b0;
  csa_component32 csa_component32_u_CSAwallace_pg_rca16_csa12_csa_component_out(.a(u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s11), .b(u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_c11), .c(u_CSAwallace_pg_rca16_csa12_csa_component_u_CSAwallace_pg_rca16_csa_s12), .csa_component32_out(u_CSAwallace_pg_rca16_csa12_csa_component_out));
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[0] = u_CSAwallace_pg_rca16_csa12_csa_component_out[0];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[1] = u_CSAwallace_pg_rca16_csa12_csa_component_out[1];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[2] = u_CSAwallace_pg_rca16_csa12_csa_component_out[2];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[3] = u_CSAwallace_pg_rca16_csa12_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[4] = u_CSAwallace_pg_rca16_csa12_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[5] = u_CSAwallace_pg_rca16_csa12_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[6] = u_CSAwallace_pg_rca16_csa12_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[7] = u_CSAwallace_pg_rca16_csa12_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[8] = u_CSAwallace_pg_rca16_csa12_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[9] = u_CSAwallace_pg_rca16_csa12_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[10] = u_CSAwallace_pg_rca16_csa12_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[11] = u_CSAwallace_pg_rca16_csa12_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[12] = u_CSAwallace_pg_rca16_csa12_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[13] = u_CSAwallace_pg_rca16_csa12_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[14] = u_CSAwallace_pg_rca16_csa12_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[15] = u_CSAwallace_pg_rca16_csa12_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[16] = u_CSAwallace_pg_rca16_csa12_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[17] = u_CSAwallace_pg_rca16_csa12_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[18] = u_CSAwallace_pg_rca16_csa12_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[19] = u_CSAwallace_pg_rca16_csa12_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[20] = u_CSAwallace_pg_rca16_csa12_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[21] = u_CSAwallace_pg_rca16_csa12_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[22] = u_CSAwallace_pg_rca16_csa12_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[23] = u_CSAwallace_pg_rca16_csa12_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[24] = u_CSAwallace_pg_rca16_csa12_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[25] = u_CSAwallace_pg_rca16_csa12_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[26] = u_CSAwallace_pg_rca16_csa12_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[27] = u_CSAwallace_pg_rca16_csa12_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[28] = u_CSAwallace_pg_rca16_csa12_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[29] = u_CSAwallace_pg_rca16_csa12_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[30] = u_CSAwallace_pg_rca16_csa12_csa_component_out[30];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[6] = u_CSAwallace_pg_rca16_csa12_csa_component_out[39];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[7] = u_CSAwallace_pg_rca16_csa12_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[8] = u_CSAwallace_pg_rca16_csa12_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[9] = u_CSAwallace_pg_rca16_csa12_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[10] = u_CSAwallace_pg_rca16_csa12_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[11] = u_CSAwallace_pg_rca16_csa12_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[12] = u_CSAwallace_pg_rca16_csa12_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[13] = u_CSAwallace_pg_rca16_csa12_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[14] = u_CSAwallace_pg_rca16_csa12_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[15] = u_CSAwallace_pg_rca16_csa12_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[16] = u_CSAwallace_pg_rca16_csa12_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[17] = u_CSAwallace_pg_rca16_csa12_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[18] = u_CSAwallace_pg_rca16_csa12_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[19] = u_CSAwallace_pg_rca16_csa12_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[20] = u_CSAwallace_pg_rca16_csa12_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[21] = u_CSAwallace_pg_rca16_csa12_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[22] = u_CSAwallace_pg_rca16_csa12_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[23] = u_CSAwallace_pg_rca16_csa12_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[24] = u_CSAwallace_pg_rca16_csa12_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[25] = u_CSAwallace_pg_rca16_csa12_csa_component_out[58];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[26] = u_CSAwallace_pg_rca16_csa12_csa_component_out[59];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[27] = u_CSAwallace_pg_rca16_csa12_csa_component_out[60];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[28] = u_CSAwallace_pg_rca16_csa12_csa_component_out[61];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[29] = u_CSAwallace_pg_rca16_csa12_csa_component_out[62];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[30] = u_CSAwallace_pg_rca16_csa12_csa_component_out[63];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[7] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[8] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[9] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[10] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[11] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[12] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[13] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[14] = 1'b0;
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[15] = u_CSAwallace_pg_rca16_csa11_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[16] = u_CSAwallace_pg_rca16_csa11_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[17] = u_CSAwallace_pg_rca16_csa11_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[18] = u_CSAwallace_pg_rca16_csa11_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[19] = u_CSAwallace_pg_rca16_csa11_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[20] = u_CSAwallace_pg_rca16_csa11_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[21] = u_CSAwallace_pg_rca16_csa11_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[22] = u_CSAwallace_pg_rca16_csa11_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[23] = u_CSAwallace_pg_rca16_csa11_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[24] = u_CSAwallace_pg_rca16_csa11_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[25] = u_CSAwallace_pg_rca16_csa11_csa_component_out[58];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[26] = u_CSAwallace_pg_rca16_csa11_csa_component_out[59];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[27] = u_CSAwallace_pg_rca16_csa11_csa_component_out[60];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[28] = u_CSAwallace_pg_rca16_csa11_csa_component_out[61];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[29] = u_CSAwallace_pg_rca16_csa11_csa_component_out[62];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[30] = u_CSAwallace_pg_rca16_csa11_csa_component_out[63];
  assign u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12[31] = 1'b0;
  csa_component32 csa_component32_u_CSAwallace_pg_rca16_csa13_csa_component_out(.a(u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_s13), .b(u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c13), .c(u_CSAwallace_pg_rca16_csa13_csa_component_u_CSAwallace_pg_rca16_csa_c12), .csa_component32_out(u_CSAwallace_pg_rca16_csa13_csa_component_out));
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[0] = u_CSAwallace_pg_rca16_csa13_csa_component_out[0];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[1] = u_CSAwallace_pg_rca16_csa13_csa_component_out[1];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[2] = u_CSAwallace_pg_rca16_csa13_csa_component_out[2];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[3] = u_CSAwallace_pg_rca16_csa13_csa_component_out[3];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[4] = u_CSAwallace_pg_rca16_csa13_csa_component_out[4];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[5] = u_CSAwallace_pg_rca16_csa13_csa_component_out[5];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[6] = u_CSAwallace_pg_rca16_csa13_csa_component_out[6];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[7] = u_CSAwallace_pg_rca16_csa13_csa_component_out[7];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[8] = u_CSAwallace_pg_rca16_csa13_csa_component_out[8];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[9] = u_CSAwallace_pg_rca16_csa13_csa_component_out[9];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[10] = u_CSAwallace_pg_rca16_csa13_csa_component_out[10];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[11] = u_CSAwallace_pg_rca16_csa13_csa_component_out[11];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[12] = u_CSAwallace_pg_rca16_csa13_csa_component_out[12];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[13] = u_CSAwallace_pg_rca16_csa13_csa_component_out[13];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[14] = u_CSAwallace_pg_rca16_csa13_csa_component_out[14];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[15] = u_CSAwallace_pg_rca16_csa13_csa_component_out[15];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[16] = u_CSAwallace_pg_rca16_csa13_csa_component_out[16];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[17] = u_CSAwallace_pg_rca16_csa13_csa_component_out[17];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[18] = u_CSAwallace_pg_rca16_csa13_csa_component_out[18];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[19] = u_CSAwallace_pg_rca16_csa13_csa_component_out[19];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[20] = u_CSAwallace_pg_rca16_csa13_csa_component_out[20];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[21] = u_CSAwallace_pg_rca16_csa13_csa_component_out[21];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[22] = u_CSAwallace_pg_rca16_csa13_csa_component_out[22];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[23] = u_CSAwallace_pg_rca16_csa13_csa_component_out[23];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[24] = u_CSAwallace_pg_rca16_csa13_csa_component_out[24];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[25] = u_CSAwallace_pg_rca16_csa13_csa_component_out[25];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[26] = u_CSAwallace_pg_rca16_csa13_csa_component_out[26];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[27] = u_CSAwallace_pg_rca16_csa13_csa_component_out[27];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[28] = u_CSAwallace_pg_rca16_csa13_csa_component_out[28];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[29] = u_CSAwallace_pg_rca16_csa13_csa_component_out[29];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[30] = u_CSAwallace_pg_rca16_csa13_csa_component_out[30];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_a[31] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[0] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[1] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[2] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[3] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[4] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[5] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[6] = 1'b0;
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[7] = u_CSAwallace_pg_rca16_csa13_csa_component_out[40];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[8] = u_CSAwallace_pg_rca16_csa13_csa_component_out[41];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[9] = u_CSAwallace_pg_rca16_csa13_csa_component_out[42];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[10] = u_CSAwallace_pg_rca16_csa13_csa_component_out[43];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[11] = u_CSAwallace_pg_rca16_csa13_csa_component_out[44];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[12] = u_CSAwallace_pg_rca16_csa13_csa_component_out[45];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[13] = u_CSAwallace_pg_rca16_csa13_csa_component_out[46];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[14] = u_CSAwallace_pg_rca16_csa13_csa_component_out[47];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[15] = u_CSAwallace_pg_rca16_csa13_csa_component_out[48];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[16] = u_CSAwallace_pg_rca16_csa13_csa_component_out[49];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[17] = u_CSAwallace_pg_rca16_csa13_csa_component_out[50];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[18] = u_CSAwallace_pg_rca16_csa13_csa_component_out[51];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[19] = u_CSAwallace_pg_rca16_csa13_csa_component_out[52];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[20] = u_CSAwallace_pg_rca16_csa13_csa_component_out[53];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[21] = u_CSAwallace_pg_rca16_csa13_csa_component_out[54];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[22] = u_CSAwallace_pg_rca16_csa13_csa_component_out[55];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[23] = u_CSAwallace_pg_rca16_csa13_csa_component_out[56];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[24] = u_CSAwallace_pg_rca16_csa13_csa_component_out[57];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[25] = u_CSAwallace_pg_rca16_csa13_csa_component_out[58];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[26] = u_CSAwallace_pg_rca16_csa13_csa_component_out[59];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[27] = u_CSAwallace_pg_rca16_csa13_csa_component_out[60];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[28] = u_CSAwallace_pg_rca16_csa13_csa_component_out[61];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[29] = u_CSAwallace_pg_rca16_csa13_csa_component_out[62];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[30] = u_CSAwallace_pg_rca16_csa13_csa_component_out[63];
  assign u_CSAwallace_pg_rca16_u_pg_rca32_b[31] = u_CSAwallace_pg_rca16_csa13_csa_component_out[64];
  u_pg_rca32 u_pg_rca32_u_CSAwallace_pg_rca16_u_pg_rca32_out(.a(u_CSAwallace_pg_rca16_u_pg_rca32_a), .b(u_CSAwallace_pg_rca16_u_pg_rca32_b), .u_pg_rca32_out(u_CSAwallace_pg_rca16_u_pg_rca32_out));

  assign u_CSAwallace_pg_rca16_out[0] = u_CSAwallace_pg_rca16_u_pg_rca32_out[0];
  assign u_CSAwallace_pg_rca16_out[1] = u_CSAwallace_pg_rca16_u_pg_rca32_out[1];
  assign u_CSAwallace_pg_rca16_out[2] = u_CSAwallace_pg_rca16_u_pg_rca32_out[2];
  assign u_CSAwallace_pg_rca16_out[3] = u_CSAwallace_pg_rca16_u_pg_rca32_out[3];
  assign u_CSAwallace_pg_rca16_out[4] = u_CSAwallace_pg_rca16_u_pg_rca32_out[4];
  assign u_CSAwallace_pg_rca16_out[5] = u_CSAwallace_pg_rca16_u_pg_rca32_out[5];
  assign u_CSAwallace_pg_rca16_out[6] = u_CSAwallace_pg_rca16_u_pg_rca32_out[6];
  assign u_CSAwallace_pg_rca16_out[7] = u_CSAwallace_pg_rca16_u_pg_rca32_out[7];
  assign u_CSAwallace_pg_rca16_out[8] = u_CSAwallace_pg_rca16_u_pg_rca32_out[8];
  assign u_CSAwallace_pg_rca16_out[9] = u_CSAwallace_pg_rca16_u_pg_rca32_out[9];
  assign u_CSAwallace_pg_rca16_out[10] = u_CSAwallace_pg_rca16_u_pg_rca32_out[10];
  assign u_CSAwallace_pg_rca16_out[11] = u_CSAwallace_pg_rca16_u_pg_rca32_out[11];
  assign u_CSAwallace_pg_rca16_out[12] = u_CSAwallace_pg_rca16_u_pg_rca32_out[12];
  assign u_CSAwallace_pg_rca16_out[13] = u_CSAwallace_pg_rca16_u_pg_rca32_out[13];
  assign u_CSAwallace_pg_rca16_out[14] = u_CSAwallace_pg_rca16_u_pg_rca32_out[14];
  assign u_CSAwallace_pg_rca16_out[15] = u_CSAwallace_pg_rca16_u_pg_rca32_out[15];
  assign u_CSAwallace_pg_rca16_out[16] = u_CSAwallace_pg_rca16_u_pg_rca32_out[16];
  assign u_CSAwallace_pg_rca16_out[17] = u_CSAwallace_pg_rca16_u_pg_rca32_out[17];
  assign u_CSAwallace_pg_rca16_out[18] = u_CSAwallace_pg_rca16_u_pg_rca32_out[18];
  assign u_CSAwallace_pg_rca16_out[19] = u_CSAwallace_pg_rca16_u_pg_rca32_out[19];
  assign u_CSAwallace_pg_rca16_out[20] = u_CSAwallace_pg_rca16_u_pg_rca32_out[20];
  assign u_CSAwallace_pg_rca16_out[21] = u_CSAwallace_pg_rca16_u_pg_rca32_out[21];
  assign u_CSAwallace_pg_rca16_out[22] = u_CSAwallace_pg_rca16_u_pg_rca32_out[22];
  assign u_CSAwallace_pg_rca16_out[23] = u_CSAwallace_pg_rca16_u_pg_rca32_out[23];
  assign u_CSAwallace_pg_rca16_out[24] = u_CSAwallace_pg_rca16_u_pg_rca32_out[24];
  assign u_CSAwallace_pg_rca16_out[25] = u_CSAwallace_pg_rca16_u_pg_rca32_out[25];
  assign u_CSAwallace_pg_rca16_out[26] = u_CSAwallace_pg_rca16_u_pg_rca32_out[26];
  assign u_CSAwallace_pg_rca16_out[27] = u_CSAwallace_pg_rca16_u_pg_rca32_out[27];
  assign u_CSAwallace_pg_rca16_out[28] = u_CSAwallace_pg_rca16_u_pg_rca32_out[28];
  assign u_CSAwallace_pg_rca16_out[29] = u_CSAwallace_pg_rca16_u_pg_rca32_out[29];
  assign u_CSAwallace_pg_rca16_out[30] = u_CSAwallace_pg_rca16_u_pg_rca32_out[30];
  assign u_CSAwallace_pg_rca16_out[31] = u_CSAwallace_pg_rca16_u_pg_rca32_out[31];
endmodule