module f_u_arr_mul8(input [7:0] a, input [7:0] b, output [15:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire f_u_arr_mul8_and_0_0_a_0;
  wire f_u_arr_mul8_and_0_0_b_0;
  wire f_u_arr_mul8_and_0_0_y0;
  wire f_u_arr_mul8_and_1_0_a_1;
  wire f_u_arr_mul8_and_1_0_b_0;
  wire f_u_arr_mul8_and_1_0_y0;
  wire f_u_arr_mul8_and_2_0_a_2;
  wire f_u_arr_mul8_and_2_0_b_0;
  wire f_u_arr_mul8_and_2_0_y0;
  wire f_u_arr_mul8_and_3_0_a_3;
  wire f_u_arr_mul8_and_3_0_b_0;
  wire f_u_arr_mul8_and_3_0_y0;
  wire f_u_arr_mul8_and_4_0_a_4;
  wire f_u_arr_mul8_and_4_0_b_0;
  wire f_u_arr_mul8_and_4_0_y0;
  wire f_u_arr_mul8_and_5_0_a_5;
  wire f_u_arr_mul8_and_5_0_b_0;
  wire f_u_arr_mul8_and_5_0_y0;
  wire f_u_arr_mul8_and_6_0_a_6;
  wire f_u_arr_mul8_and_6_0_b_0;
  wire f_u_arr_mul8_and_6_0_y0;
  wire f_u_arr_mul8_and_7_0_a_7;
  wire f_u_arr_mul8_and_7_0_b_0;
  wire f_u_arr_mul8_and_7_0_y0;
  wire f_u_arr_mul8_and_0_1_a_0;
  wire f_u_arr_mul8_and_0_1_b_1;
  wire f_u_arr_mul8_and_0_1_y0;
  wire f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_0_1_y0;
  wire f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_1_0_y0;
  wire f_u_arr_mul8_ha_0_1_y0;
  wire f_u_arr_mul8_ha_0_1_y1;
  wire f_u_arr_mul8_and_1_1_a_1;
  wire f_u_arr_mul8_and_1_1_b_1;
  wire f_u_arr_mul8_and_1_1_y0;
  wire f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_1_1_y0;
  wire f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_2_0_y0;
  wire f_u_arr_mul8_fa_1_1_y0;
  wire f_u_arr_mul8_fa_1_1_y1;
  wire f_u_arr_mul8_fa_1_1_f_u_arr_mul8_ha_0_1_y1;
  wire f_u_arr_mul8_fa_1_1_y2;
  wire f_u_arr_mul8_fa_1_1_y3;
  wire f_u_arr_mul8_fa_1_1_y4;
  wire f_u_arr_mul8_and_2_1_a_2;
  wire f_u_arr_mul8_and_2_1_b_1;
  wire f_u_arr_mul8_and_2_1_y0;
  wire f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_2_1_y0;
  wire f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_3_0_y0;
  wire f_u_arr_mul8_fa_2_1_y0;
  wire f_u_arr_mul8_fa_2_1_y1;
  wire f_u_arr_mul8_fa_2_1_f_u_arr_mul8_fa_1_1_y4;
  wire f_u_arr_mul8_fa_2_1_y2;
  wire f_u_arr_mul8_fa_2_1_y3;
  wire f_u_arr_mul8_fa_2_1_y4;
  wire f_u_arr_mul8_and_3_1_a_3;
  wire f_u_arr_mul8_and_3_1_b_1;
  wire f_u_arr_mul8_and_3_1_y0;
  wire f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_3_1_y0;
  wire f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_4_0_y0;
  wire f_u_arr_mul8_fa_3_1_y0;
  wire f_u_arr_mul8_fa_3_1_y1;
  wire f_u_arr_mul8_fa_3_1_f_u_arr_mul8_fa_2_1_y4;
  wire f_u_arr_mul8_fa_3_1_y2;
  wire f_u_arr_mul8_fa_3_1_y3;
  wire f_u_arr_mul8_fa_3_1_y4;
  wire f_u_arr_mul8_and_4_1_a_4;
  wire f_u_arr_mul8_and_4_1_b_1;
  wire f_u_arr_mul8_and_4_1_y0;
  wire f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_4_1_y0;
  wire f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_5_0_y0;
  wire f_u_arr_mul8_fa_4_1_y0;
  wire f_u_arr_mul8_fa_4_1_y1;
  wire f_u_arr_mul8_fa_4_1_f_u_arr_mul8_fa_3_1_y4;
  wire f_u_arr_mul8_fa_4_1_y2;
  wire f_u_arr_mul8_fa_4_1_y3;
  wire f_u_arr_mul8_fa_4_1_y4;
  wire f_u_arr_mul8_and_5_1_a_5;
  wire f_u_arr_mul8_and_5_1_b_1;
  wire f_u_arr_mul8_and_5_1_y0;
  wire f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_5_1_y0;
  wire f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_6_0_y0;
  wire f_u_arr_mul8_fa_5_1_y0;
  wire f_u_arr_mul8_fa_5_1_y1;
  wire f_u_arr_mul8_fa_5_1_f_u_arr_mul8_fa_4_1_y4;
  wire f_u_arr_mul8_fa_5_1_y2;
  wire f_u_arr_mul8_fa_5_1_y3;
  wire f_u_arr_mul8_fa_5_1_y4;
  wire f_u_arr_mul8_and_6_1_a_6;
  wire f_u_arr_mul8_and_6_1_b_1;
  wire f_u_arr_mul8_and_6_1_y0;
  wire f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_6_1_y0;
  wire f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_7_0_y0;
  wire f_u_arr_mul8_fa_6_1_y0;
  wire f_u_arr_mul8_fa_6_1_y1;
  wire f_u_arr_mul8_fa_6_1_f_u_arr_mul8_fa_5_1_y4;
  wire f_u_arr_mul8_fa_6_1_y2;
  wire f_u_arr_mul8_fa_6_1_y3;
  wire f_u_arr_mul8_fa_6_1_y4;
  wire f_u_arr_mul8_and_7_1_a_7;
  wire f_u_arr_mul8_and_7_1_b_1;
  wire f_u_arr_mul8_and_7_1_y0;
  wire f_u_arr_mul8_ha_7_1_f_u_arr_mul8_and_7_1_y0;
  wire f_u_arr_mul8_ha_7_1_f_u_arr_mul8_fa_6_1_y4;
  wire f_u_arr_mul8_ha_7_1_y0;
  wire f_u_arr_mul8_ha_7_1_y1;
  wire f_u_arr_mul8_and_0_2_a_0;
  wire f_u_arr_mul8_and_0_2_b_2;
  wire f_u_arr_mul8_and_0_2_y0;
  wire f_u_arr_mul8_ha_0_2_f_u_arr_mul8_and_0_2_y0;
  wire f_u_arr_mul8_ha_0_2_f_u_arr_mul8_fa_1_1_y2;
  wire f_u_arr_mul8_ha_0_2_y0;
  wire f_u_arr_mul8_ha_0_2_y1;
  wire f_u_arr_mul8_and_1_2_a_1;
  wire f_u_arr_mul8_and_1_2_b_2;
  wire f_u_arr_mul8_and_1_2_y0;
  wire f_u_arr_mul8_fa_1_2_f_u_arr_mul8_and_1_2_y0;
  wire f_u_arr_mul8_fa_1_2_f_u_arr_mul8_fa_2_1_y2;
  wire f_u_arr_mul8_fa_1_2_y0;
  wire f_u_arr_mul8_fa_1_2_y1;
  wire f_u_arr_mul8_fa_1_2_f_u_arr_mul8_ha_0_2_y1;
  wire f_u_arr_mul8_fa_1_2_y2;
  wire f_u_arr_mul8_fa_1_2_y3;
  wire f_u_arr_mul8_fa_1_2_y4;
  wire f_u_arr_mul8_and_2_2_a_2;
  wire f_u_arr_mul8_and_2_2_b_2;
  wire f_u_arr_mul8_and_2_2_y0;
  wire f_u_arr_mul8_fa_2_2_f_u_arr_mul8_and_2_2_y0;
  wire f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_3_1_y2;
  wire f_u_arr_mul8_fa_2_2_y0;
  wire f_u_arr_mul8_fa_2_2_y1;
  wire f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_1_2_y4;
  wire f_u_arr_mul8_fa_2_2_y2;
  wire f_u_arr_mul8_fa_2_2_y3;
  wire f_u_arr_mul8_fa_2_2_y4;
  wire f_u_arr_mul8_and_3_2_a_3;
  wire f_u_arr_mul8_and_3_2_b_2;
  wire f_u_arr_mul8_and_3_2_y0;
  wire f_u_arr_mul8_fa_3_2_f_u_arr_mul8_and_3_2_y0;
  wire f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_4_1_y2;
  wire f_u_arr_mul8_fa_3_2_y0;
  wire f_u_arr_mul8_fa_3_2_y1;
  wire f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_2_2_y4;
  wire f_u_arr_mul8_fa_3_2_y2;
  wire f_u_arr_mul8_fa_3_2_y3;
  wire f_u_arr_mul8_fa_3_2_y4;
  wire f_u_arr_mul8_and_4_2_a_4;
  wire f_u_arr_mul8_and_4_2_b_2;
  wire f_u_arr_mul8_and_4_2_y0;
  wire f_u_arr_mul8_fa_4_2_f_u_arr_mul8_and_4_2_y0;
  wire f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_5_1_y2;
  wire f_u_arr_mul8_fa_4_2_y0;
  wire f_u_arr_mul8_fa_4_2_y1;
  wire f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_3_2_y4;
  wire f_u_arr_mul8_fa_4_2_y2;
  wire f_u_arr_mul8_fa_4_2_y3;
  wire f_u_arr_mul8_fa_4_2_y4;
  wire f_u_arr_mul8_and_5_2_a_5;
  wire f_u_arr_mul8_and_5_2_b_2;
  wire f_u_arr_mul8_and_5_2_y0;
  wire f_u_arr_mul8_fa_5_2_f_u_arr_mul8_and_5_2_y0;
  wire f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_6_1_y2;
  wire f_u_arr_mul8_fa_5_2_y0;
  wire f_u_arr_mul8_fa_5_2_y1;
  wire f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_4_2_y4;
  wire f_u_arr_mul8_fa_5_2_y2;
  wire f_u_arr_mul8_fa_5_2_y3;
  wire f_u_arr_mul8_fa_5_2_y4;
  wire f_u_arr_mul8_and_6_2_a_6;
  wire f_u_arr_mul8_and_6_2_b_2;
  wire f_u_arr_mul8_and_6_2_y0;
  wire f_u_arr_mul8_fa_6_2_f_u_arr_mul8_and_6_2_y0;
  wire f_u_arr_mul8_fa_6_2_f_u_arr_mul8_ha_7_1_y0;
  wire f_u_arr_mul8_fa_6_2_y0;
  wire f_u_arr_mul8_fa_6_2_y1;
  wire f_u_arr_mul8_fa_6_2_f_u_arr_mul8_fa_5_2_y4;
  wire f_u_arr_mul8_fa_6_2_y2;
  wire f_u_arr_mul8_fa_6_2_y3;
  wire f_u_arr_mul8_fa_6_2_y4;
  wire f_u_arr_mul8_and_7_2_a_7;
  wire f_u_arr_mul8_and_7_2_b_2;
  wire f_u_arr_mul8_and_7_2_y0;
  wire f_u_arr_mul8_fa_7_2_f_u_arr_mul8_and_7_2_y0;
  wire f_u_arr_mul8_fa_7_2_f_u_arr_mul8_ha_7_1_y1;
  wire f_u_arr_mul8_fa_7_2_y0;
  wire f_u_arr_mul8_fa_7_2_y1;
  wire f_u_arr_mul8_fa_7_2_f_u_arr_mul8_fa_6_2_y4;
  wire f_u_arr_mul8_fa_7_2_y2;
  wire f_u_arr_mul8_fa_7_2_y3;
  wire f_u_arr_mul8_fa_7_2_y4;
  wire f_u_arr_mul8_and_0_3_a_0;
  wire f_u_arr_mul8_and_0_3_b_3;
  wire f_u_arr_mul8_and_0_3_y0;
  wire f_u_arr_mul8_ha_0_3_f_u_arr_mul8_and_0_3_y0;
  wire f_u_arr_mul8_ha_0_3_f_u_arr_mul8_fa_1_2_y2;
  wire f_u_arr_mul8_ha_0_3_y0;
  wire f_u_arr_mul8_ha_0_3_y1;
  wire f_u_arr_mul8_and_1_3_a_1;
  wire f_u_arr_mul8_and_1_3_b_3;
  wire f_u_arr_mul8_and_1_3_y0;
  wire f_u_arr_mul8_fa_1_3_f_u_arr_mul8_and_1_3_y0;
  wire f_u_arr_mul8_fa_1_3_f_u_arr_mul8_fa_2_2_y2;
  wire f_u_arr_mul8_fa_1_3_y0;
  wire f_u_arr_mul8_fa_1_3_y1;
  wire f_u_arr_mul8_fa_1_3_f_u_arr_mul8_ha_0_3_y1;
  wire f_u_arr_mul8_fa_1_3_y2;
  wire f_u_arr_mul8_fa_1_3_y3;
  wire f_u_arr_mul8_fa_1_3_y4;
  wire f_u_arr_mul8_and_2_3_a_2;
  wire f_u_arr_mul8_and_2_3_b_3;
  wire f_u_arr_mul8_and_2_3_y0;
  wire f_u_arr_mul8_fa_2_3_f_u_arr_mul8_and_2_3_y0;
  wire f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_3_2_y2;
  wire f_u_arr_mul8_fa_2_3_y0;
  wire f_u_arr_mul8_fa_2_3_y1;
  wire f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_1_3_y4;
  wire f_u_arr_mul8_fa_2_3_y2;
  wire f_u_arr_mul8_fa_2_3_y3;
  wire f_u_arr_mul8_fa_2_3_y4;
  wire f_u_arr_mul8_and_3_3_a_3;
  wire f_u_arr_mul8_and_3_3_b_3;
  wire f_u_arr_mul8_and_3_3_y0;
  wire f_u_arr_mul8_fa_3_3_f_u_arr_mul8_and_3_3_y0;
  wire f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_4_2_y2;
  wire f_u_arr_mul8_fa_3_3_y0;
  wire f_u_arr_mul8_fa_3_3_y1;
  wire f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_2_3_y4;
  wire f_u_arr_mul8_fa_3_3_y2;
  wire f_u_arr_mul8_fa_3_3_y3;
  wire f_u_arr_mul8_fa_3_3_y4;
  wire f_u_arr_mul8_and_4_3_a_4;
  wire f_u_arr_mul8_and_4_3_b_3;
  wire f_u_arr_mul8_and_4_3_y0;
  wire f_u_arr_mul8_fa_4_3_f_u_arr_mul8_and_4_3_y0;
  wire f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_5_2_y2;
  wire f_u_arr_mul8_fa_4_3_y0;
  wire f_u_arr_mul8_fa_4_3_y1;
  wire f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_3_3_y4;
  wire f_u_arr_mul8_fa_4_3_y2;
  wire f_u_arr_mul8_fa_4_3_y3;
  wire f_u_arr_mul8_fa_4_3_y4;
  wire f_u_arr_mul8_and_5_3_a_5;
  wire f_u_arr_mul8_and_5_3_b_3;
  wire f_u_arr_mul8_and_5_3_y0;
  wire f_u_arr_mul8_fa_5_3_f_u_arr_mul8_and_5_3_y0;
  wire f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_6_2_y2;
  wire f_u_arr_mul8_fa_5_3_y0;
  wire f_u_arr_mul8_fa_5_3_y1;
  wire f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_4_3_y4;
  wire f_u_arr_mul8_fa_5_3_y2;
  wire f_u_arr_mul8_fa_5_3_y3;
  wire f_u_arr_mul8_fa_5_3_y4;
  wire f_u_arr_mul8_and_6_3_a_6;
  wire f_u_arr_mul8_and_6_3_b_3;
  wire f_u_arr_mul8_and_6_3_y0;
  wire f_u_arr_mul8_fa_6_3_f_u_arr_mul8_and_6_3_y0;
  wire f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_7_2_y2;
  wire f_u_arr_mul8_fa_6_3_y0;
  wire f_u_arr_mul8_fa_6_3_y1;
  wire f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_5_3_y4;
  wire f_u_arr_mul8_fa_6_3_y2;
  wire f_u_arr_mul8_fa_6_3_y3;
  wire f_u_arr_mul8_fa_6_3_y4;
  wire f_u_arr_mul8_and_7_3_a_7;
  wire f_u_arr_mul8_and_7_3_b_3;
  wire f_u_arr_mul8_and_7_3_y0;
  wire f_u_arr_mul8_fa_7_3_f_u_arr_mul8_and_7_3_y0;
  wire f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_7_2_y4;
  wire f_u_arr_mul8_fa_7_3_y0;
  wire f_u_arr_mul8_fa_7_3_y1;
  wire f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_6_3_y4;
  wire f_u_arr_mul8_fa_7_3_y2;
  wire f_u_arr_mul8_fa_7_3_y3;
  wire f_u_arr_mul8_fa_7_3_y4;
  wire f_u_arr_mul8_and_0_4_a_0;
  wire f_u_arr_mul8_and_0_4_b_4;
  wire f_u_arr_mul8_and_0_4_y0;
  wire f_u_arr_mul8_ha_0_4_f_u_arr_mul8_and_0_4_y0;
  wire f_u_arr_mul8_ha_0_4_f_u_arr_mul8_fa_1_3_y2;
  wire f_u_arr_mul8_ha_0_4_y0;
  wire f_u_arr_mul8_ha_0_4_y1;
  wire f_u_arr_mul8_and_1_4_a_1;
  wire f_u_arr_mul8_and_1_4_b_4;
  wire f_u_arr_mul8_and_1_4_y0;
  wire f_u_arr_mul8_fa_1_4_f_u_arr_mul8_and_1_4_y0;
  wire f_u_arr_mul8_fa_1_4_f_u_arr_mul8_fa_2_3_y2;
  wire f_u_arr_mul8_fa_1_4_y0;
  wire f_u_arr_mul8_fa_1_4_y1;
  wire f_u_arr_mul8_fa_1_4_f_u_arr_mul8_ha_0_4_y1;
  wire f_u_arr_mul8_fa_1_4_y2;
  wire f_u_arr_mul8_fa_1_4_y3;
  wire f_u_arr_mul8_fa_1_4_y4;
  wire f_u_arr_mul8_and_2_4_a_2;
  wire f_u_arr_mul8_and_2_4_b_4;
  wire f_u_arr_mul8_and_2_4_y0;
  wire f_u_arr_mul8_fa_2_4_f_u_arr_mul8_and_2_4_y0;
  wire f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_3_3_y2;
  wire f_u_arr_mul8_fa_2_4_y0;
  wire f_u_arr_mul8_fa_2_4_y1;
  wire f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_1_4_y4;
  wire f_u_arr_mul8_fa_2_4_y2;
  wire f_u_arr_mul8_fa_2_4_y3;
  wire f_u_arr_mul8_fa_2_4_y4;
  wire f_u_arr_mul8_and_3_4_a_3;
  wire f_u_arr_mul8_and_3_4_b_4;
  wire f_u_arr_mul8_and_3_4_y0;
  wire f_u_arr_mul8_fa_3_4_f_u_arr_mul8_and_3_4_y0;
  wire f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_4_3_y2;
  wire f_u_arr_mul8_fa_3_4_y0;
  wire f_u_arr_mul8_fa_3_4_y1;
  wire f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_2_4_y4;
  wire f_u_arr_mul8_fa_3_4_y2;
  wire f_u_arr_mul8_fa_3_4_y3;
  wire f_u_arr_mul8_fa_3_4_y4;
  wire f_u_arr_mul8_and_4_4_a_4;
  wire f_u_arr_mul8_and_4_4_b_4;
  wire f_u_arr_mul8_and_4_4_y0;
  wire f_u_arr_mul8_fa_4_4_f_u_arr_mul8_and_4_4_y0;
  wire f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_5_3_y2;
  wire f_u_arr_mul8_fa_4_4_y0;
  wire f_u_arr_mul8_fa_4_4_y1;
  wire f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_3_4_y4;
  wire f_u_arr_mul8_fa_4_4_y2;
  wire f_u_arr_mul8_fa_4_4_y3;
  wire f_u_arr_mul8_fa_4_4_y4;
  wire f_u_arr_mul8_and_5_4_a_5;
  wire f_u_arr_mul8_and_5_4_b_4;
  wire f_u_arr_mul8_and_5_4_y0;
  wire f_u_arr_mul8_fa_5_4_f_u_arr_mul8_and_5_4_y0;
  wire f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_6_3_y2;
  wire f_u_arr_mul8_fa_5_4_y0;
  wire f_u_arr_mul8_fa_5_4_y1;
  wire f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_4_4_y4;
  wire f_u_arr_mul8_fa_5_4_y2;
  wire f_u_arr_mul8_fa_5_4_y3;
  wire f_u_arr_mul8_fa_5_4_y4;
  wire f_u_arr_mul8_and_6_4_a_6;
  wire f_u_arr_mul8_and_6_4_b_4;
  wire f_u_arr_mul8_and_6_4_y0;
  wire f_u_arr_mul8_fa_6_4_f_u_arr_mul8_and_6_4_y0;
  wire f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_7_3_y2;
  wire f_u_arr_mul8_fa_6_4_y0;
  wire f_u_arr_mul8_fa_6_4_y1;
  wire f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_5_4_y4;
  wire f_u_arr_mul8_fa_6_4_y2;
  wire f_u_arr_mul8_fa_6_4_y3;
  wire f_u_arr_mul8_fa_6_4_y4;
  wire f_u_arr_mul8_and_7_4_a_7;
  wire f_u_arr_mul8_and_7_4_b_4;
  wire f_u_arr_mul8_and_7_4_y0;
  wire f_u_arr_mul8_fa_7_4_f_u_arr_mul8_and_7_4_y0;
  wire f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_7_3_y4;
  wire f_u_arr_mul8_fa_7_4_y0;
  wire f_u_arr_mul8_fa_7_4_y1;
  wire f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_6_4_y4;
  wire f_u_arr_mul8_fa_7_4_y2;
  wire f_u_arr_mul8_fa_7_4_y3;
  wire f_u_arr_mul8_fa_7_4_y4;
  wire f_u_arr_mul8_and_0_5_a_0;
  wire f_u_arr_mul8_and_0_5_b_5;
  wire f_u_arr_mul8_and_0_5_y0;
  wire f_u_arr_mul8_ha_0_5_f_u_arr_mul8_and_0_5_y0;
  wire f_u_arr_mul8_ha_0_5_f_u_arr_mul8_fa_1_4_y2;
  wire f_u_arr_mul8_ha_0_5_y0;
  wire f_u_arr_mul8_ha_0_5_y1;
  wire f_u_arr_mul8_and_1_5_a_1;
  wire f_u_arr_mul8_and_1_5_b_5;
  wire f_u_arr_mul8_and_1_5_y0;
  wire f_u_arr_mul8_fa_1_5_f_u_arr_mul8_and_1_5_y0;
  wire f_u_arr_mul8_fa_1_5_f_u_arr_mul8_fa_2_4_y2;
  wire f_u_arr_mul8_fa_1_5_y0;
  wire f_u_arr_mul8_fa_1_5_y1;
  wire f_u_arr_mul8_fa_1_5_f_u_arr_mul8_ha_0_5_y1;
  wire f_u_arr_mul8_fa_1_5_y2;
  wire f_u_arr_mul8_fa_1_5_y3;
  wire f_u_arr_mul8_fa_1_5_y4;
  wire f_u_arr_mul8_and_2_5_a_2;
  wire f_u_arr_mul8_and_2_5_b_5;
  wire f_u_arr_mul8_and_2_5_y0;
  wire f_u_arr_mul8_fa_2_5_f_u_arr_mul8_and_2_5_y0;
  wire f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_3_4_y2;
  wire f_u_arr_mul8_fa_2_5_y0;
  wire f_u_arr_mul8_fa_2_5_y1;
  wire f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_1_5_y4;
  wire f_u_arr_mul8_fa_2_5_y2;
  wire f_u_arr_mul8_fa_2_5_y3;
  wire f_u_arr_mul8_fa_2_5_y4;
  wire f_u_arr_mul8_and_3_5_a_3;
  wire f_u_arr_mul8_and_3_5_b_5;
  wire f_u_arr_mul8_and_3_5_y0;
  wire f_u_arr_mul8_fa_3_5_f_u_arr_mul8_and_3_5_y0;
  wire f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_4_4_y2;
  wire f_u_arr_mul8_fa_3_5_y0;
  wire f_u_arr_mul8_fa_3_5_y1;
  wire f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_2_5_y4;
  wire f_u_arr_mul8_fa_3_5_y2;
  wire f_u_arr_mul8_fa_3_5_y3;
  wire f_u_arr_mul8_fa_3_5_y4;
  wire f_u_arr_mul8_and_4_5_a_4;
  wire f_u_arr_mul8_and_4_5_b_5;
  wire f_u_arr_mul8_and_4_5_y0;
  wire f_u_arr_mul8_fa_4_5_f_u_arr_mul8_and_4_5_y0;
  wire f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_5_4_y2;
  wire f_u_arr_mul8_fa_4_5_y0;
  wire f_u_arr_mul8_fa_4_5_y1;
  wire f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_3_5_y4;
  wire f_u_arr_mul8_fa_4_5_y2;
  wire f_u_arr_mul8_fa_4_5_y3;
  wire f_u_arr_mul8_fa_4_5_y4;
  wire f_u_arr_mul8_and_5_5_a_5;
  wire f_u_arr_mul8_and_5_5_b_5;
  wire f_u_arr_mul8_and_5_5_y0;
  wire f_u_arr_mul8_fa_5_5_f_u_arr_mul8_and_5_5_y0;
  wire f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_6_4_y2;
  wire f_u_arr_mul8_fa_5_5_y0;
  wire f_u_arr_mul8_fa_5_5_y1;
  wire f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_4_5_y4;
  wire f_u_arr_mul8_fa_5_5_y2;
  wire f_u_arr_mul8_fa_5_5_y3;
  wire f_u_arr_mul8_fa_5_5_y4;
  wire f_u_arr_mul8_and_6_5_a_6;
  wire f_u_arr_mul8_and_6_5_b_5;
  wire f_u_arr_mul8_and_6_5_y0;
  wire f_u_arr_mul8_fa_6_5_f_u_arr_mul8_and_6_5_y0;
  wire f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_7_4_y2;
  wire f_u_arr_mul8_fa_6_5_y0;
  wire f_u_arr_mul8_fa_6_5_y1;
  wire f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_5_5_y4;
  wire f_u_arr_mul8_fa_6_5_y2;
  wire f_u_arr_mul8_fa_6_5_y3;
  wire f_u_arr_mul8_fa_6_5_y4;
  wire f_u_arr_mul8_and_7_5_a_7;
  wire f_u_arr_mul8_and_7_5_b_5;
  wire f_u_arr_mul8_and_7_5_y0;
  wire f_u_arr_mul8_fa_7_5_f_u_arr_mul8_and_7_5_y0;
  wire f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_7_4_y4;
  wire f_u_arr_mul8_fa_7_5_y0;
  wire f_u_arr_mul8_fa_7_5_y1;
  wire f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_6_5_y4;
  wire f_u_arr_mul8_fa_7_5_y2;
  wire f_u_arr_mul8_fa_7_5_y3;
  wire f_u_arr_mul8_fa_7_5_y4;
  wire f_u_arr_mul8_and_0_6_a_0;
  wire f_u_arr_mul8_and_0_6_b_6;
  wire f_u_arr_mul8_and_0_6_y0;
  wire f_u_arr_mul8_ha_0_6_f_u_arr_mul8_and_0_6_y0;
  wire f_u_arr_mul8_ha_0_6_f_u_arr_mul8_fa_1_5_y2;
  wire f_u_arr_mul8_ha_0_6_y0;
  wire f_u_arr_mul8_ha_0_6_y1;
  wire f_u_arr_mul8_and_1_6_a_1;
  wire f_u_arr_mul8_and_1_6_b_6;
  wire f_u_arr_mul8_and_1_6_y0;
  wire f_u_arr_mul8_fa_1_6_f_u_arr_mul8_and_1_6_y0;
  wire f_u_arr_mul8_fa_1_6_f_u_arr_mul8_fa_2_5_y2;
  wire f_u_arr_mul8_fa_1_6_y0;
  wire f_u_arr_mul8_fa_1_6_y1;
  wire f_u_arr_mul8_fa_1_6_f_u_arr_mul8_ha_0_6_y1;
  wire f_u_arr_mul8_fa_1_6_y2;
  wire f_u_arr_mul8_fa_1_6_y3;
  wire f_u_arr_mul8_fa_1_6_y4;
  wire f_u_arr_mul8_and_2_6_a_2;
  wire f_u_arr_mul8_and_2_6_b_6;
  wire f_u_arr_mul8_and_2_6_y0;
  wire f_u_arr_mul8_fa_2_6_f_u_arr_mul8_and_2_6_y0;
  wire f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_3_5_y2;
  wire f_u_arr_mul8_fa_2_6_y0;
  wire f_u_arr_mul8_fa_2_6_y1;
  wire f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_1_6_y4;
  wire f_u_arr_mul8_fa_2_6_y2;
  wire f_u_arr_mul8_fa_2_6_y3;
  wire f_u_arr_mul8_fa_2_6_y4;
  wire f_u_arr_mul8_and_3_6_a_3;
  wire f_u_arr_mul8_and_3_6_b_6;
  wire f_u_arr_mul8_and_3_6_y0;
  wire f_u_arr_mul8_fa_3_6_f_u_arr_mul8_and_3_6_y0;
  wire f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_4_5_y2;
  wire f_u_arr_mul8_fa_3_6_y0;
  wire f_u_arr_mul8_fa_3_6_y1;
  wire f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_2_6_y4;
  wire f_u_arr_mul8_fa_3_6_y2;
  wire f_u_arr_mul8_fa_3_6_y3;
  wire f_u_arr_mul8_fa_3_6_y4;
  wire f_u_arr_mul8_and_4_6_a_4;
  wire f_u_arr_mul8_and_4_6_b_6;
  wire f_u_arr_mul8_and_4_6_y0;
  wire f_u_arr_mul8_fa_4_6_f_u_arr_mul8_and_4_6_y0;
  wire f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_5_5_y2;
  wire f_u_arr_mul8_fa_4_6_y0;
  wire f_u_arr_mul8_fa_4_6_y1;
  wire f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_3_6_y4;
  wire f_u_arr_mul8_fa_4_6_y2;
  wire f_u_arr_mul8_fa_4_6_y3;
  wire f_u_arr_mul8_fa_4_6_y4;
  wire f_u_arr_mul8_and_5_6_a_5;
  wire f_u_arr_mul8_and_5_6_b_6;
  wire f_u_arr_mul8_and_5_6_y0;
  wire f_u_arr_mul8_fa_5_6_f_u_arr_mul8_and_5_6_y0;
  wire f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_6_5_y2;
  wire f_u_arr_mul8_fa_5_6_y0;
  wire f_u_arr_mul8_fa_5_6_y1;
  wire f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_4_6_y4;
  wire f_u_arr_mul8_fa_5_6_y2;
  wire f_u_arr_mul8_fa_5_6_y3;
  wire f_u_arr_mul8_fa_5_6_y4;
  wire f_u_arr_mul8_and_6_6_a_6;
  wire f_u_arr_mul8_and_6_6_b_6;
  wire f_u_arr_mul8_and_6_6_y0;
  wire f_u_arr_mul8_fa_6_6_f_u_arr_mul8_and_6_6_y0;
  wire f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_7_5_y2;
  wire f_u_arr_mul8_fa_6_6_y0;
  wire f_u_arr_mul8_fa_6_6_y1;
  wire f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_5_6_y4;
  wire f_u_arr_mul8_fa_6_6_y2;
  wire f_u_arr_mul8_fa_6_6_y3;
  wire f_u_arr_mul8_fa_6_6_y4;
  wire f_u_arr_mul8_and_7_6_a_7;
  wire f_u_arr_mul8_and_7_6_b_6;
  wire f_u_arr_mul8_and_7_6_y0;
  wire f_u_arr_mul8_fa_7_6_f_u_arr_mul8_and_7_6_y0;
  wire f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_7_5_y4;
  wire f_u_arr_mul8_fa_7_6_y0;
  wire f_u_arr_mul8_fa_7_6_y1;
  wire f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_6_6_y4;
  wire f_u_arr_mul8_fa_7_6_y2;
  wire f_u_arr_mul8_fa_7_6_y3;
  wire f_u_arr_mul8_fa_7_6_y4;
  wire f_u_arr_mul8_and_0_7_a_0;
  wire f_u_arr_mul8_and_0_7_b_7;
  wire f_u_arr_mul8_and_0_7_y0;
  wire f_u_arr_mul8_ha_0_7_f_u_arr_mul8_and_0_7_y0;
  wire f_u_arr_mul8_ha_0_7_f_u_arr_mul8_fa_1_6_y2;
  wire f_u_arr_mul8_ha_0_7_y0;
  wire f_u_arr_mul8_ha_0_7_y1;
  wire f_u_arr_mul8_and_1_7_a_1;
  wire f_u_arr_mul8_and_1_7_b_7;
  wire f_u_arr_mul8_and_1_7_y0;
  wire f_u_arr_mul8_fa_1_7_f_u_arr_mul8_and_1_7_y0;
  wire f_u_arr_mul8_fa_1_7_f_u_arr_mul8_fa_2_6_y2;
  wire f_u_arr_mul8_fa_1_7_y0;
  wire f_u_arr_mul8_fa_1_7_y1;
  wire f_u_arr_mul8_fa_1_7_f_u_arr_mul8_ha_0_7_y1;
  wire f_u_arr_mul8_fa_1_7_y2;
  wire f_u_arr_mul8_fa_1_7_y3;
  wire f_u_arr_mul8_fa_1_7_y4;
  wire f_u_arr_mul8_and_2_7_a_2;
  wire f_u_arr_mul8_and_2_7_b_7;
  wire f_u_arr_mul8_and_2_7_y0;
  wire f_u_arr_mul8_fa_2_7_f_u_arr_mul8_and_2_7_y0;
  wire f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_3_6_y2;
  wire f_u_arr_mul8_fa_2_7_y0;
  wire f_u_arr_mul8_fa_2_7_y1;
  wire f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_1_7_y4;
  wire f_u_arr_mul8_fa_2_7_y2;
  wire f_u_arr_mul8_fa_2_7_y3;
  wire f_u_arr_mul8_fa_2_7_y4;
  wire f_u_arr_mul8_and_3_7_a_3;
  wire f_u_arr_mul8_and_3_7_b_7;
  wire f_u_arr_mul8_and_3_7_y0;
  wire f_u_arr_mul8_fa_3_7_f_u_arr_mul8_and_3_7_y0;
  wire f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_4_6_y2;
  wire f_u_arr_mul8_fa_3_7_y0;
  wire f_u_arr_mul8_fa_3_7_y1;
  wire f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_2_7_y4;
  wire f_u_arr_mul8_fa_3_7_y2;
  wire f_u_arr_mul8_fa_3_7_y3;
  wire f_u_arr_mul8_fa_3_7_y4;
  wire f_u_arr_mul8_and_4_7_a_4;
  wire f_u_arr_mul8_and_4_7_b_7;
  wire f_u_arr_mul8_and_4_7_y0;
  wire f_u_arr_mul8_fa_4_7_f_u_arr_mul8_and_4_7_y0;
  wire f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_5_6_y2;
  wire f_u_arr_mul8_fa_4_7_y0;
  wire f_u_arr_mul8_fa_4_7_y1;
  wire f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_3_7_y4;
  wire f_u_arr_mul8_fa_4_7_y2;
  wire f_u_arr_mul8_fa_4_7_y3;
  wire f_u_arr_mul8_fa_4_7_y4;
  wire f_u_arr_mul8_and_5_7_a_5;
  wire f_u_arr_mul8_and_5_7_b_7;
  wire f_u_arr_mul8_and_5_7_y0;
  wire f_u_arr_mul8_fa_5_7_f_u_arr_mul8_and_5_7_y0;
  wire f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_6_6_y2;
  wire f_u_arr_mul8_fa_5_7_y0;
  wire f_u_arr_mul8_fa_5_7_y1;
  wire f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_4_7_y4;
  wire f_u_arr_mul8_fa_5_7_y2;
  wire f_u_arr_mul8_fa_5_7_y3;
  wire f_u_arr_mul8_fa_5_7_y4;
  wire f_u_arr_mul8_and_6_7_a_6;
  wire f_u_arr_mul8_and_6_7_b_7;
  wire f_u_arr_mul8_and_6_7_y0;
  wire f_u_arr_mul8_fa_6_7_f_u_arr_mul8_and_6_7_y0;
  wire f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_7_6_y2;
  wire f_u_arr_mul8_fa_6_7_y0;
  wire f_u_arr_mul8_fa_6_7_y1;
  wire f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_5_7_y4;
  wire f_u_arr_mul8_fa_6_7_y2;
  wire f_u_arr_mul8_fa_6_7_y3;
  wire f_u_arr_mul8_fa_6_7_y4;
  wire f_u_arr_mul8_and_7_7_a_7;
  wire f_u_arr_mul8_and_7_7_b_7;
  wire f_u_arr_mul8_and_7_7_y0;
  wire f_u_arr_mul8_fa_7_7_f_u_arr_mul8_and_7_7_y0;
  wire f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_7_6_y4;
  wire f_u_arr_mul8_fa_7_7_y0;
  wire f_u_arr_mul8_fa_7_7_y1;
  wire f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_6_7_y4;
  wire f_u_arr_mul8_fa_7_7_y2;
  wire f_u_arr_mul8_fa_7_7_y3;
  wire f_u_arr_mul8_fa_7_7_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign f_u_arr_mul8_and_0_0_a_0 = a_0;
  assign f_u_arr_mul8_and_0_0_b_0 = b_0;
  assign f_u_arr_mul8_and_0_0_y0 = f_u_arr_mul8_and_0_0_a_0 & f_u_arr_mul8_and_0_0_b_0;
  assign f_u_arr_mul8_and_1_0_a_1 = a_1;
  assign f_u_arr_mul8_and_1_0_b_0 = b_0;
  assign f_u_arr_mul8_and_1_0_y0 = f_u_arr_mul8_and_1_0_a_1 & f_u_arr_mul8_and_1_0_b_0;
  assign f_u_arr_mul8_and_2_0_a_2 = a_2;
  assign f_u_arr_mul8_and_2_0_b_0 = b_0;
  assign f_u_arr_mul8_and_2_0_y0 = f_u_arr_mul8_and_2_0_a_2 & f_u_arr_mul8_and_2_0_b_0;
  assign f_u_arr_mul8_and_3_0_a_3 = a_3;
  assign f_u_arr_mul8_and_3_0_b_0 = b_0;
  assign f_u_arr_mul8_and_3_0_y0 = f_u_arr_mul8_and_3_0_a_3 & f_u_arr_mul8_and_3_0_b_0;
  assign f_u_arr_mul8_and_4_0_a_4 = a_4;
  assign f_u_arr_mul8_and_4_0_b_0 = b_0;
  assign f_u_arr_mul8_and_4_0_y0 = f_u_arr_mul8_and_4_0_a_4 & f_u_arr_mul8_and_4_0_b_0;
  assign f_u_arr_mul8_and_5_0_a_5 = a_5;
  assign f_u_arr_mul8_and_5_0_b_0 = b_0;
  assign f_u_arr_mul8_and_5_0_y0 = f_u_arr_mul8_and_5_0_a_5 & f_u_arr_mul8_and_5_0_b_0;
  assign f_u_arr_mul8_and_6_0_a_6 = a_6;
  assign f_u_arr_mul8_and_6_0_b_0 = b_0;
  assign f_u_arr_mul8_and_6_0_y0 = f_u_arr_mul8_and_6_0_a_6 & f_u_arr_mul8_and_6_0_b_0;
  assign f_u_arr_mul8_and_7_0_a_7 = a_7;
  assign f_u_arr_mul8_and_7_0_b_0 = b_0;
  assign f_u_arr_mul8_and_7_0_y0 = f_u_arr_mul8_and_7_0_a_7 & f_u_arr_mul8_and_7_0_b_0;
  assign f_u_arr_mul8_and_0_1_a_0 = a_0;
  assign f_u_arr_mul8_and_0_1_b_1 = b_1;
  assign f_u_arr_mul8_and_0_1_y0 = f_u_arr_mul8_and_0_1_a_0 & f_u_arr_mul8_and_0_1_b_1;
  assign f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_0_1_y0 = f_u_arr_mul8_and_0_1_y0;
  assign f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_1_0_y0 = f_u_arr_mul8_and_1_0_y0;
  assign f_u_arr_mul8_ha_0_1_y0 = f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_0_1_y0 ^ f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_1_0_y0;
  assign f_u_arr_mul8_ha_0_1_y1 = f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_0_1_y0 & f_u_arr_mul8_ha_0_1_f_u_arr_mul8_and_1_0_y0;
  assign f_u_arr_mul8_and_1_1_a_1 = a_1;
  assign f_u_arr_mul8_and_1_1_b_1 = b_1;
  assign f_u_arr_mul8_and_1_1_y0 = f_u_arr_mul8_and_1_1_a_1 & f_u_arr_mul8_and_1_1_b_1;
  assign f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_1_1_y0 = f_u_arr_mul8_and_1_1_y0;
  assign f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_2_0_y0 = f_u_arr_mul8_and_2_0_y0;
  assign f_u_arr_mul8_fa_1_1_f_u_arr_mul8_ha_0_1_y1 = f_u_arr_mul8_ha_0_1_y1;
  assign f_u_arr_mul8_fa_1_1_y0 = f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_1_1_y0 ^ f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_2_0_y0;
  assign f_u_arr_mul8_fa_1_1_y1 = f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_1_1_y0 & f_u_arr_mul8_fa_1_1_f_u_arr_mul8_and_2_0_y0;
  assign f_u_arr_mul8_fa_1_1_y2 = f_u_arr_mul8_fa_1_1_y0 ^ f_u_arr_mul8_fa_1_1_f_u_arr_mul8_ha_0_1_y1;
  assign f_u_arr_mul8_fa_1_1_y3 = f_u_arr_mul8_fa_1_1_y0 & f_u_arr_mul8_fa_1_1_f_u_arr_mul8_ha_0_1_y1;
  assign f_u_arr_mul8_fa_1_1_y4 = f_u_arr_mul8_fa_1_1_y1 | f_u_arr_mul8_fa_1_1_y3;
  assign f_u_arr_mul8_and_2_1_a_2 = a_2;
  assign f_u_arr_mul8_and_2_1_b_1 = b_1;
  assign f_u_arr_mul8_and_2_1_y0 = f_u_arr_mul8_and_2_1_a_2 & f_u_arr_mul8_and_2_1_b_1;
  assign f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_2_1_y0 = f_u_arr_mul8_and_2_1_y0;
  assign f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_3_0_y0 = f_u_arr_mul8_and_3_0_y0;
  assign f_u_arr_mul8_fa_2_1_f_u_arr_mul8_fa_1_1_y4 = f_u_arr_mul8_fa_1_1_y4;
  assign f_u_arr_mul8_fa_2_1_y0 = f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_2_1_y0 ^ f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_3_0_y0;
  assign f_u_arr_mul8_fa_2_1_y1 = f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_2_1_y0 & f_u_arr_mul8_fa_2_1_f_u_arr_mul8_and_3_0_y0;
  assign f_u_arr_mul8_fa_2_1_y2 = f_u_arr_mul8_fa_2_1_y0 ^ f_u_arr_mul8_fa_2_1_f_u_arr_mul8_fa_1_1_y4;
  assign f_u_arr_mul8_fa_2_1_y3 = f_u_arr_mul8_fa_2_1_y0 & f_u_arr_mul8_fa_2_1_f_u_arr_mul8_fa_1_1_y4;
  assign f_u_arr_mul8_fa_2_1_y4 = f_u_arr_mul8_fa_2_1_y1 | f_u_arr_mul8_fa_2_1_y3;
  assign f_u_arr_mul8_and_3_1_a_3 = a_3;
  assign f_u_arr_mul8_and_3_1_b_1 = b_1;
  assign f_u_arr_mul8_and_3_1_y0 = f_u_arr_mul8_and_3_1_a_3 & f_u_arr_mul8_and_3_1_b_1;
  assign f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_3_1_y0 = f_u_arr_mul8_and_3_1_y0;
  assign f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_4_0_y0 = f_u_arr_mul8_and_4_0_y0;
  assign f_u_arr_mul8_fa_3_1_f_u_arr_mul8_fa_2_1_y4 = f_u_arr_mul8_fa_2_1_y4;
  assign f_u_arr_mul8_fa_3_1_y0 = f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_3_1_y0 ^ f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_4_0_y0;
  assign f_u_arr_mul8_fa_3_1_y1 = f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_3_1_y0 & f_u_arr_mul8_fa_3_1_f_u_arr_mul8_and_4_0_y0;
  assign f_u_arr_mul8_fa_3_1_y2 = f_u_arr_mul8_fa_3_1_y0 ^ f_u_arr_mul8_fa_3_1_f_u_arr_mul8_fa_2_1_y4;
  assign f_u_arr_mul8_fa_3_1_y3 = f_u_arr_mul8_fa_3_1_y0 & f_u_arr_mul8_fa_3_1_f_u_arr_mul8_fa_2_1_y4;
  assign f_u_arr_mul8_fa_3_1_y4 = f_u_arr_mul8_fa_3_1_y1 | f_u_arr_mul8_fa_3_1_y3;
  assign f_u_arr_mul8_and_4_1_a_4 = a_4;
  assign f_u_arr_mul8_and_4_1_b_1 = b_1;
  assign f_u_arr_mul8_and_4_1_y0 = f_u_arr_mul8_and_4_1_a_4 & f_u_arr_mul8_and_4_1_b_1;
  assign f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_4_1_y0 = f_u_arr_mul8_and_4_1_y0;
  assign f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_5_0_y0 = f_u_arr_mul8_and_5_0_y0;
  assign f_u_arr_mul8_fa_4_1_f_u_arr_mul8_fa_3_1_y4 = f_u_arr_mul8_fa_3_1_y4;
  assign f_u_arr_mul8_fa_4_1_y0 = f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_4_1_y0 ^ f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_5_0_y0;
  assign f_u_arr_mul8_fa_4_1_y1 = f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_4_1_y0 & f_u_arr_mul8_fa_4_1_f_u_arr_mul8_and_5_0_y0;
  assign f_u_arr_mul8_fa_4_1_y2 = f_u_arr_mul8_fa_4_1_y0 ^ f_u_arr_mul8_fa_4_1_f_u_arr_mul8_fa_3_1_y4;
  assign f_u_arr_mul8_fa_4_1_y3 = f_u_arr_mul8_fa_4_1_y0 & f_u_arr_mul8_fa_4_1_f_u_arr_mul8_fa_3_1_y4;
  assign f_u_arr_mul8_fa_4_1_y4 = f_u_arr_mul8_fa_4_1_y1 | f_u_arr_mul8_fa_4_1_y3;
  assign f_u_arr_mul8_and_5_1_a_5 = a_5;
  assign f_u_arr_mul8_and_5_1_b_1 = b_1;
  assign f_u_arr_mul8_and_5_1_y0 = f_u_arr_mul8_and_5_1_a_5 & f_u_arr_mul8_and_5_1_b_1;
  assign f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_5_1_y0 = f_u_arr_mul8_and_5_1_y0;
  assign f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_6_0_y0 = f_u_arr_mul8_and_6_0_y0;
  assign f_u_arr_mul8_fa_5_1_f_u_arr_mul8_fa_4_1_y4 = f_u_arr_mul8_fa_4_1_y4;
  assign f_u_arr_mul8_fa_5_1_y0 = f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_5_1_y0 ^ f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_6_0_y0;
  assign f_u_arr_mul8_fa_5_1_y1 = f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_5_1_y0 & f_u_arr_mul8_fa_5_1_f_u_arr_mul8_and_6_0_y0;
  assign f_u_arr_mul8_fa_5_1_y2 = f_u_arr_mul8_fa_5_1_y0 ^ f_u_arr_mul8_fa_5_1_f_u_arr_mul8_fa_4_1_y4;
  assign f_u_arr_mul8_fa_5_1_y3 = f_u_arr_mul8_fa_5_1_y0 & f_u_arr_mul8_fa_5_1_f_u_arr_mul8_fa_4_1_y4;
  assign f_u_arr_mul8_fa_5_1_y4 = f_u_arr_mul8_fa_5_1_y1 | f_u_arr_mul8_fa_5_1_y3;
  assign f_u_arr_mul8_and_6_1_a_6 = a_6;
  assign f_u_arr_mul8_and_6_1_b_1 = b_1;
  assign f_u_arr_mul8_and_6_1_y0 = f_u_arr_mul8_and_6_1_a_6 & f_u_arr_mul8_and_6_1_b_1;
  assign f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_6_1_y0 = f_u_arr_mul8_and_6_1_y0;
  assign f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_7_0_y0 = f_u_arr_mul8_and_7_0_y0;
  assign f_u_arr_mul8_fa_6_1_f_u_arr_mul8_fa_5_1_y4 = f_u_arr_mul8_fa_5_1_y4;
  assign f_u_arr_mul8_fa_6_1_y0 = f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_6_1_y0 ^ f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_7_0_y0;
  assign f_u_arr_mul8_fa_6_1_y1 = f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_6_1_y0 & f_u_arr_mul8_fa_6_1_f_u_arr_mul8_and_7_0_y0;
  assign f_u_arr_mul8_fa_6_1_y2 = f_u_arr_mul8_fa_6_1_y0 ^ f_u_arr_mul8_fa_6_1_f_u_arr_mul8_fa_5_1_y4;
  assign f_u_arr_mul8_fa_6_1_y3 = f_u_arr_mul8_fa_6_1_y0 & f_u_arr_mul8_fa_6_1_f_u_arr_mul8_fa_5_1_y4;
  assign f_u_arr_mul8_fa_6_1_y4 = f_u_arr_mul8_fa_6_1_y1 | f_u_arr_mul8_fa_6_1_y3;
  assign f_u_arr_mul8_and_7_1_a_7 = a_7;
  assign f_u_arr_mul8_and_7_1_b_1 = b_1;
  assign f_u_arr_mul8_and_7_1_y0 = f_u_arr_mul8_and_7_1_a_7 & f_u_arr_mul8_and_7_1_b_1;
  assign f_u_arr_mul8_ha_7_1_f_u_arr_mul8_and_7_1_y0 = f_u_arr_mul8_and_7_1_y0;
  assign f_u_arr_mul8_ha_7_1_f_u_arr_mul8_fa_6_1_y4 = f_u_arr_mul8_fa_6_1_y4;
  assign f_u_arr_mul8_ha_7_1_y0 = f_u_arr_mul8_ha_7_1_f_u_arr_mul8_and_7_1_y0 ^ f_u_arr_mul8_ha_7_1_f_u_arr_mul8_fa_6_1_y4;
  assign f_u_arr_mul8_ha_7_1_y1 = f_u_arr_mul8_ha_7_1_f_u_arr_mul8_and_7_1_y0 & f_u_arr_mul8_ha_7_1_f_u_arr_mul8_fa_6_1_y4;
  assign f_u_arr_mul8_and_0_2_a_0 = a_0;
  assign f_u_arr_mul8_and_0_2_b_2 = b_2;
  assign f_u_arr_mul8_and_0_2_y0 = f_u_arr_mul8_and_0_2_a_0 & f_u_arr_mul8_and_0_2_b_2;
  assign f_u_arr_mul8_ha_0_2_f_u_arr_mul8_and_0_2_y0 = f_u_arr_mul8_and_0_2_y0;
  assign f_u_arr_mul8_ha_0_2_f_u_arr_mul8_fa_1_1_y2 = f_u_arr_mul8_fa_1_1_y2;
  assign f_u_arr_mul8_ha_0_2_y0 = f_u_arr_mul8_ha_0_2_f_u_arr_mul8_and_0_2_y0 ^ f_u_arr_mul8_ha_0_2_f_u_arr_mul8_fa_1_1_y2;
  assign f_u_arr_mul8_ha_0_2_y1 = f_u_arr_mul8_ha_0_2_f_u_arr_mul8_and_0_2_y0 & f_u_arr_mul8_ha_0_2_f_u_arr_mul8_fa_1_1_y2;
  assign f_u_arr_mul8_and_1_2_a_1 = a_1;
  assign f_u_arr_mul8_and_1_2_b_2 = b_2;
  assign f_u_arr_mul8_and_1_2_y0 = f_u_arr_mul8_and_1_2_a_1 & f_u_arr_mul8_and_1_2_b_2;
  assign f_u_arr_mul8_fa_1_2_f_u_arr_mul8_and_1_2_y0 = f_u_arr_mul8_and_1_2_y0;
  assign f_u_arr_mul8_fa_1_2_f_u_arr_mul8_fa_2_1_y2 = f_u_arr_mul8_fa_2_1_y2;
  assign f_u_arr_mul8_fa_1_2_f_u_arr_mul8_ha_0_2_y1 = f_u_arr_mul8_ha_0_2_y1;
  assign f_u_arr_mul8_fa_1_2_y0 = f_u_arr_mul8_fa_1_2_f_u_arr_mul8_and_1_2_y0 ^ f_u_arr_mul8_fa_1_2_f_u_arr_mul8_fa_2_1_y2;
  assign f_u_arr_mul8_fa_1_2_y1 = f_u_arr_mul8_fa_1_2_f_u_arr_mul8_and_1_2_y0 & f_u_arr_mul8_fa_1_2_f_u_arr_mul8_fa_2_1_y2;
  assign f_u_arr_mul8_fa_1_2_y2 = f_u_arr_mul8_fa_1_2_y0 ^ f_u_arr_mul8_fa_1_2_f_u_arr_mul8_ha_0_2_y1;
  assign f_u_arr_mul8_fa_1_2_y3 = f_u_arr_mul8_fa_1_2_y0 & f_u_arr_mul8_fa_1_2_f_u_arr_mul8_ha_0_2_y1;
  assign f_u_arr_mul8_fa_1_2_y4 = f_u_arr_mul8_fa_1_2_y1 | f_u_arr_mul8_fa_1_2_y3;
  assign f_u_arr_mul8_and_2_2_a_2 = a_2;
  assign f_u_arr_mul8_and_2_2_b_2 = b_2;
  assign f_u_arr_mul8_and_2_2_y0 = f_u_arr_mul8_and_2_2_a_2 & f_u_arr_mul8_and_2_2_b_2;
  assign f_u_arr_mul8_fa_2_2_f_u_arr_mul8_and_2_2_y0 = f_u_arr_mul8_and_2_2_y0;
  assign f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_3_1_y2 = f_u_arr_mul8_fa_3_1_y2;
  assign f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_1_2_y4 = f_u_arr_mul8_fa_1_2_y4;
  assign f_u_arr_mul8_fa_2_2_y0 = f_u_arr_mul8_fa_2_2_f_u_arr_mul8_and_2_2_y0 ^ f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_3_1_y2;
  assign f_u_arr_mul8_fa_2_2_y1 = f_u_arr_mul8_fa_2_2_f_u_arr_mul8_and_2_2_y0 & f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_3_1_y2;
  assign f_u_arr_mul8_fa_2_2_y2 = f_u_arr_mul8_fa_2_2_y0 ^ f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_1_2_y4;
  assign f_u_arr_mul8_fa_2_2_y3 = f_u_arr_mul8_fa_2_2_y0 & f_u_arr_mul8_fa_2_2_f_u_arr_mul8_fa_1_2_y4;
  assign f_u_arr_mul8_fa_2_2_y4 = f_u_arr_mul8_fa_2_2_y1 | f_u_arr_mul8_fa_2_2_y3;
  assign f_u_arr_mul8_and_3_2_a_3 = a_3;
  assign f_u_arr_mul8_and_3_2_b_2 = b_2;
  assign f_u_arr_mul8_and_3_2_y0 = f_u_arr_mul8_and_3_2_a_3 & f_u_arr_mul8_and_3_2_b_2;
  assign f_u_arr_mul8_fa_3_2_f_u_arr_mul8_and_3_2_y0 = f_u_arr_mul8_and_3_2_y0;
  assign f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_4_1_y2 = f_u_arr_mul8_fa_4_1_y2;
  assign f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_2_2_y4 = f_u_arr_mul8_fa_2_2_y4;
  assign f_u_arr_mul8_fa_3_2_y0 = f_u_arr_mul8_fa_3_2_f_u_arr_mul8_and_3_2_y0 ^ f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_4_1_y2;
  assign f_u_arr_mul8_fa_3_2_y1 = f_u_arr_mul8_fa_3_2_f_u_arr_mul8_and_3_2_y0 & f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_4_1_y2;
  assign f_u_arr_mul8_fa_3_2_y2 = f_u_arr_mul8_fa_3_2_y0 ^ f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_2_2_y4;
  assign f_u_arr_mul8_fa_3_2_y3 = f_u_arr_mul8_fa_3_2_y0 & f_u_arr_mul8_fa_3_2_f_u_arr_mul8_fa_2_2_y4;
  assign f_u_arr_mul8_fa_3_2_y4 = f_u_arr_mul8_fa_3_2_y1 | f_u_arr_mul8_fa_3_2_y3;
  assign f_u_arr_mul8_and_4_2_a_4 = a_4;
  assign f_u_arr_mul8_and_4_2_b_2 = b_2;
  assign f_u_arr_mul8_and_4_2_y0 = f_u_arr_mul8_and_4_2_a_4 & f_u_arr_mul8_and_4_2_b_2;
  assign f_u_arr_mul8_fa_4_2_f_u_arr_mul8_and_4_2_y0 = f_u_arr_mul8_and_4_2_y0;
  assign f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_5_1_y2 = f_u_arr_mul8_fa_5_1_y2;
  assign f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_3_2_y4 = f_u_arr_mul8_fa_3_2_y4;
  assign f_u_arr_mul8_fa_4_2_y0 = f_u_arr_mul8_fa_4_2_f_u_arr_mul8_and_4_2_y0 ^ f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_5_1_y2;
  assign f_u_arr_mul8_fa_4_2_y1 = f_u_arr_mul8_fa_4_2_f_u_arr_mul8_and_4_2_y0 & f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_5_1_y2;
  assign f_u_arr_mul8_fa_4_2_y2 = f_u_arr_mul8_fa_4_2_y0 ^ f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_3_2_y4;
  assign f_u_arr_mul8_fa_4_2_y3 = f_u_arr_mul8_fa_4_2_y0 & f_u_arr_mul8_fa_4_2_f_u_arr_mul8_fa_3_2_y4;
  assign f_u_arr_mul8_fa_4_2_y4 = f_u_arr_mul8_fa_4_2_y1 | f_u_arr_mul8_fa_4_2_y3;
  assign f_u_arr_mul8_and_5_2_a_5 = a_5;
  assign f_u_arr_mul8_and_5_2_b_2 = b_2;
  assign f_u_arr_mul8_and_5_2_y0 = f_u_arr_mul8_and_5_2_a_5 & f_u_arr_mul8_and_5_2_b_2;
  assign f_u_arr_mul8_fa_5_2_f_u_arr_mul8_and_5_2_y0 = f_u_arr_mul8_and_5_2_y0;
  assign f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_6_1_y2 = f_u_arr_mul8_fa_6_1_y2;
  assign f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_4_2_y4 = f_u_arr_mul8_fa_4_2_y4;
  assign f_u_arr_mul8_fa_5_2_y0 = f_u_arr_mul8_fa_5_2_f_u_arr_mul8_and_5_2_y0 ^ f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_6_1_y2;
  assign f_u_arr_mul8_fa_5_2_y1 = f_u_arr_mul8_fa_5_2_f_u_arr_mul8_and_5_2_y0 & f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_6_1_y2;
  assign f_u_arr_mul8_fa_5_2_y2 = f_u_arr_mul8_fa_5_2_y0 ^ f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_4_2_y4;
  assign f_u_arr_mul8_fa_5_2_y3 = f_u_arr_mul8_fa_5_2_y0 & f_u_arr_mul8_fa_5_2_f_u_arr_mul8_fa_4_2_y4;
  assign f_u_arr_mul8_fa_5_2_y4 = f_u_arr_mul8_fa_5_2_y1 | f_u_arr_mul8_fa_5_2_y3;
  assign f_u_arr_mul8_and_6_2_a_6 = a_6;
  assign f_u_arr_mul8_and_6_2_b_2 = b_2;
  assign f_u_arr_mul8_and_6_2_y0 = f_u_arr_mul8_and_6_2_a_6 & f_u_arr_mul8_and_6_2_b_2;
  assign f_u_arr_mul8_fa_6_2_f_u_arr_mul8_and_6_2_y0 = f_u_arr_mul8_and_6_2_y0;
  assign f_u_arr_mul8_fa_6_2_f_u_arr_mul8_ha_7_1_y0 = f_u_arr_mul8_ha_7_1_y0;
  assign f_u_arr_mul8_fa_6_2_f_u_arr_mul8_fa_5_2_y4 = f_u_arr_mul8_fa_5_2_y4;
  assign f_u_arr_mul8_fa_6_2_y0 = f_u_arr_mul8_fa_6_2_f_u_arr_mul8_and_6_2_y0 ^ f_u_arr_mul8_fa_6_2_f_u_arr_mul8_ha_7_1_y0;
  assign f_u_arr_mul8_fa_6_2_y1 = f_u_arr_mul8_fa_6_2_f_u_arr_mul8_and_6_2_y0 & f_u_arr_mul8_fa_6_2_f_u_arr_mul8_ha_7_1_y0;
  assign f_u_arr_mul8_fa_6_2_y2 = f_u_arr_mul8_fa_6_2_y0 ^ f_u_arr_mul8_fa_6_2_f_u_arr_mul8_fa_5_2_y4;
  assign f_u_arr_mul8_fa_6_2_y3 = f_u_arr_mul8_fa_6_2_y0 & f_u_arr_mul8_fa_6_2_f_u_arr_mul8_fa_5_2_y4;
  assign f_u_arr_mul8_fa_6_2_y4 = f_u_arr_mul8_fa_6_2_y1 | f_u_arr_mul8_fa_6_2_y3;
  assign f_u_arr_mul8_and_7_2_a_7 = a_7;
  assign f_u_arr_mul8_and_7_2_b_2 = b_2;
  assign f_u_arr_mul8_and_7_2_y0 = f_u_arr_mul8_and_7_2_a_7 & f_u_arr_mul8_and_7_2_b_2;
  assign f_u_arr_mul8_fa_7_2_f_u_arr_mul8_and_7_2_y0 = f_u_arr_mul8_and_7_2_y0;
  assign f_u_arr_mul8_fa_7_2_f_u_arr_mul8_ha_7_1_y1 = f_u_arr_mul8_ha_7_1_y1;
  assign f_u_arr_mul8_fa_7_2_f_u_arr_mul8_fa_6_2_y4 = f_u_arr_mul8_fa_6_2_y4;
  assign f_u_arr_mul8_fa_7_2_y0 = f_u_arr_mul8_fa_7_2_f_u_arr_mul8_and_7_2_y0 ^ f_u_arr_mul8_fa_7_2_f_u_arr_mul8_ha_7_1_y1;
  assign f_u_arr_mul8_fa_7_2_y1 = f_u_arr_mul8_fa_7_2_f_u_arr_mul8_and_7_2_y0 & f_u_arr_mul8_fa_7_2_f_u_arr_mul8_ha_7_1_y1;
  assign f_u_arr_mul8_fa_7_2_y2 = f_u_arr_mul8_fa_7_2_y0 ^ f_u_arr_mul8_fa_7_2_f_u_arr_mul8_fa_6_2_y4;
  assign f_u_arr_mul8_fa_7_2_y3 = f_u_arr_mul8_fa_7_2_y0 & f_u_arr_mul8_fa_7_2_f_u_arr_mul8_fa_6_2_y4;
  assign f_u_arr_mul8_fa_7_2_y4 = f_u_arr_mul8_fa_7_2_y1 | f_u_arr_mul8_fa_7_2_y3;
  assign f_u_arr_mul8_and_0_3_a_0 = a_0;
  assign f_u_arr_mul8_and_0_3_b_3 = b_3;
  assign f_u_arr_mul8_and_0_3_y0 = f_u_arr_mul8_and_0_3_a_0 & f_u_arr_mul8_and_0_3_b_3;
  assign f_u_arr_mul8_ha_0_3_f_u_arr_mul8_and_0_3_y0 = f_u_arr_mul8_and_0_3_y0;
  assign f_u_arr_mul8_ha_0_3_f_u_arr_mul8_fa_1_2_y2 = f_u_arr_mul8_fa_1_2_y2;
  assign f_u_arr_mul8_ha_0_3_y0 = f_u_arr_mul8_ha_0_3_f_u_arr_mul8_and_0_3_y0 ^ f_u_arr_mul8_ha_0_3_f_u_arr_mul8_fa_1_2_y2;
  assign f_u_arr_mul8_ha_0_3_y1 = f_u_arr_mul8_ha_0_3_f_u_arr_mul8_and_0_3_y0 & f_u_arr_mul8_ha_0_3_f_u_arr_mul8_fa_1_2_y2;
  assign f_u_arr_mul8_and_1_3_a_1 = a_1;
  assign f_u_arr_mul8_and_1_3_b_3 = b_3;
  assign f_u_arr_mul8_and_1_3_y0 = f_u_arr_mul8_and_1_3_a_1 & f_u_arr_mul8_and_1_3_b_3;
  assign f_u_arr_mul8_fa_1_3_f_u_arr_mul8_and_1_3_y0 = f_u_arr_mul8_and_1_3_y0;
  assign f_u_arr_mul8_fa_1_3_f_u_arr_mul8_fa_2_2_y2 = f_u_arr_mul8_fa_2_2_y2;
  assign f_u_arr_mul8_fa_1_3_f_u_arr_mul8_ha_0_3_y1 = f_u_arr_mul8_ha_0_3_y1;
  assign f_u_arr_mul8_fa_1_3_y0 = f_u_arr_mul8_fa_1_3_f_u_arr_mul8_and_1_3_y0 ^ f_u_arr_mul8_fa_1_3_f_u_arr_mul8_fa_2_2_y2;
  assign f_u_arr_mul8_fa_1_3_y1 = f_u_arr_mul8_fa_1_3_f_u_arr_mul8_and_1_3_y0 & f_u_arr_mul8_fa_1_3_f_u_arr_mul8_fa_2_2_y2;
  assign f_u_arr_mul8_fa_1_3_y2 = f_u_arr_mul8_fa_1_3_y0 ^ f_u_arr_mul8_fa_1_3_f_u_arr_mul8_ha_0_3_y1;
  assign f_u_arr_mul8_fa_1_3_y3 = f_u_arr_mul8_fa_1_3_y0 & f_u_arr_mul8_fa_1_3_f_u_arr_mul8_ha_0_3_y1;
  assign f_u_arr_mul8_fa_1_3_y4 = f_u_arr_mul8_fa_1_3_y1 | f_u_arr_mul8_fa_1_3_y3;
  assign f_u_arr_mul8_and_2_3_a_2 = a_2;
  assign f_u_arr_mul8_and_2_3_b_3 = b_3;
  assign f_u_arr_mul8_and_2_3_y0 = f_u_arr_mul8_and_2_3_a_2 & f_u_arr_mul8_and_2_3_b_3;
  assign f_u_arr_mul8_fa_2_3_f_u_arr_mul8_and_2_3_y0 = f_u_arr_mul8_and_2_3_y0;
  assign f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_3_2_y2 = f_u_arr_mul8_fa_3_2_y2;
  assign f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_1_3_y4 = f_u_arr_mul8_fa_1_3_y4;
  assign f_u_arr_mul8_fa_2_3_y0 = f_u_arr_mul8_fa_2_3_f_u_arr_mul8_and_2_3_y0 ^ f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_3_2_y2;
  assign f_u_arr_mul8_fa_2_3_y1 = f_u_arr_mul8_fa_2_3_f_u_arr_mul8_and_2_3_y0 & f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_3_2_y2;
  assign f_u_arr_mul8_fa_2_3_y2 = f_u_arr_mul8_fa_2_3_y0 ^ f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_1_3_y4;
  assign f_u_arr_mul8_fa_2_3_y3 = f_u_arr_mul8_fa_2_3_y0 & f_u_arr_mul8_fa_2_3_f_u_arr_mul8_fa_1_3_y4;
  assign f_u_arr_mul8_fa_2_3_y4 = f_u_arr_mul8_fa_2_3_y1 | f_u_arr_mul8_fa_2_3_y3;
  assign f_u_arr_mul8_and_3_3_a_3 = a_3;
  assign f_u_arr_mul8_and_3_3_b_3 = b_3;
  assign f_u_arr_mul8_and_3_3_y0 = f_u_arr_mul8_and_3_3_a_3 & f_u_arr_mul8_and_3_3_b_3;
  assign f_u_arr_mul8_fa_3_3_f_u_arr_mul8_and_3_3_y0 = f_u_arr_mul8_and_3_3_y0;
  assign f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_4_2_y2 = f_u_arr_mul8_fa_4_2_y2;
  assign f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_2_3_y4 = f_u_arr_mul8_fa_2_3_y4;
  assign f_u_arr_mul8_fa_3_3_y0 = f_u_arr_mul8_fa_3_3_f_u_arr_mul8_and_3_3_y0 ^ f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_4_2_y2;
  assign f_u_arr_mul8_fa_3_3_y1 = f_u_arr_mul8_fa_3_3_f_u_arr_mul8_and_3_3_y0 & f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_4_2_y2;
  assign f_u_arr_mul8_fa_3_3_y2 = f_u_arr_mul8_fa_3_3_y0 ^ f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_2_3_y4;
  assign f_u_arr_mul8_fa_3_3_y3 = f_u_arr_mul8_fa_3_3_y0 & f_u_arr_mul8_fa_3_3_f_u_arr_mul8_fa_2_3_y4;
  assign f_u_arr_mul8_fa_3_3_y4 = f_u_arr_mul8_fa_3_3_y1 | f_u_arr_mul8_fa_3_3_y3;
  assign f_u_arr_mul8_and_4_3_a_4 = a_4;
  assign f_u_arr_mul8_and_4_3_b_3 = b_3;
  assign f_u_arr_mul8_and_4_3_y0 = f_u_arr_mul8_and_4_3_a_4 & f_u_arr_mul8_and_4_3_b_3;
  assign f_u_arr_mul8_fa_4_3_f_u_arr_mul8_and_4_3_y0 = f_u_arr_mul8_and_4_3_y0;
  assign f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_5_2_y2 = f_u_arr_mul8_fa_5_2_y2;
  assign f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_3_3_y4 = f_u_arr_mul8_fa_3_3_y4;
  assign f_u_arr_mul8_fa_4_3_y0 = f_u_arr_mul8_fa_4_3_f_u_arr_mul8_and_4_3_y0 ^ f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_5_2_y2;
  assign f_u_arr_mul8_fa_4_3_y1 = f_u_arr_mul8_fa_4_3_f_u_arr_mul8_and_4_3_y0 & f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_5_2_y2;
  assign f_u_arr_mul8_fa_4_3_y2 = f_u_arr_mul8_fa_4_3_y0 ^ f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_3_3_y4;
  assign f_u_arr_mul8_fa_4_3_y3 = f_u_arr_mul8_fa_4_3_y0 & f_u_arr_mul8_fa_4_3_f_u_arr_mul8_fa_3_3_y4;
  assign f_u_arr_mul8_fa_4_3_y4 = f_u_arr_mul8_fa_4_3_y1 | f_u_arr_mul8_fa_4_3_y3;
  assign f_u_arr_mul8_and_5_3_a_5 = a_5;
  assign f_u_arr_mul8_and_5_3_b_3 = b_3;
  assign f_u_arr_mul8_and_5_3_y0 = f_u_arr_mul8_and_5_3_a_5 & f_u_arr_mul8_and_5_3_b_3;
  assign f_u_arr_mul8_fa_5_3_f_u_arr_mul8_and_5_3_y0 = f_u_arr_mul8_and_5_3_y0;
  assign f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_6_2_y2 = f_u_arr_mul8_fa_6_2_y2;
  assign f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_4_3_y4 = f_u_arr_mul8_fa_4_3_y4;
  assign f_u_arr_mul8_fa_5_3_y0 = f_u_arr_mul8_fa_5_3_f_u_arr_mul8_and_5_3_y0 ^ f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_6_2_y2;
  assign f_u_arr_mul8_fa_5_3_y1 = f_u_arr_mul8_fa_5_3_f_u_arr_mul8_and_5_3_y0 & f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_6_2_y2;
  assign f_u_arr_mul8_fa_5_3_y2 = f_u_arr_mul8_fa_5_3_y0 ^ f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_4_3_y4;
  assign f_u_arr_mul8_fa_5_3_y3 = f_u_arr_mul8_fa_5_3_y0 & f_u_arr_mul8_fa_5_3_f_u_arr_mul8_fa_4_3_y4;
  assign f_u_arr_mul8_fa_5_3_y4 = f_u_arr_mul8_fa_5_3_y1 | f_u_arr_mul8_fa_5_3_y3;
  assign f_u_arr_mul8_and_6_3_a_6 = a_6;
  assign f_u_arr_mul8_and_6_3_b_3 = b_3;
  assign f_u_arr_mul8_and_6_3_y0 = f_u_arr_mul8_and_6_3_a_6 & f_u_arr_mul8_and_6_3_b_3;
  assign f_u_arr_mul8_fa_6_3_f_u_arr_mul8_and_6_3_y0 = f_u_arr_mul8_and_6_3_y0;
  assign f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_7_2_y2 = f_u_arr_mul8_fa_7_2_y2;
  assign f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_5_3_y4 = f_u_arr_mul8_fa_5_3_y4;
  assign f_u_arr_mul8_fa_6_3_y0 = f_u_arr_mul8_fa_6_3_f_u_arr_mul8_and_6_3_y0 ^ f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_7_2_y2;
  assign f_u_arr_mul8_fa_6_3_y1 = f_u_arr_mul8_fa_6_3_f_u_arr_mul8_and_6_3_y0 & f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_7_2_y2;
  assign f_u_arr_mul8_fa_6_3_y2 = f_u_arr_mul8_fa_6_3_y0 ^ f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_5_3_y4;
  assign f_u_arr_mul8_fa_6_3_y3 = f_u_arr_mul8_fa_6_3_y0 & f_u_arr_mul8_fa_6_3_f_u_arr_mul8_fa_5_3_y4;
  assign f_u_arr_mul8_fa_6_3_y4 = f_u_arr_mul8_fa_6_3_y1 | f_u_arr_mul8_fa_6_3_y3;
  assign f_u_arr_mul8_and_7_3_a_7 = a_7;
  assign f_u_arr_mul8_and_7_3_b_3 = b_3;
  assign f_u_arr_mul8_and_7_3_y0 = f_u_arr_mul8_and_7_3_a_7 & f_u_arr_mul8_and_7_3_b_3;
  assign f_u_arr_mul8_fa_7_3_f_u_arr_mul8_and_7_3_y0 = f_u_arr_mul8_and_7_3_y0;
  assign f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_7_2_y4 = f_u_arr_mul8_fa_7_2_y4;
  assign f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_6_3_y4 = f_u_arr_mul8_fa_6_3_y4;
  assign f_u_arr_mul8_fa_7_3_y0 = f_u_arr_mul8_fa_7_3_f_u_arr_mul8_and_7_3_y0 ^ f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_7_2_y4;
  assign f_u_arr_mul8_fa_7_3_y1 = f_u_arr_mul8_fa_7_3_f_u_arr_mul8_and_7_3_y0 & f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_7_2_y4;
  assign f_u_arr_mul8_fa_7_3_y2 = f_u_arr_mul8_fa_7_3_y0 ^ f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_6_3_y4;
  assign f_u_arr_mul8_fa_7_3_y3 = f_u_arr_mul8_fa_7_3_y0 & f_u_arr_mul8_fa_7_3_f_u_arr_mul8_fa_6_3_y4;
  assign f_u_arr_mul8_fa_7_3_y4 = f_u_arr_mul8_fa_7_3_y1 | f_u_arr_mul8_fa_7_3_y3;
  assign f_u_arr_mul8_and_0_4_a_0 = a_0;
  assign f_u_arr_mul8_and_0_4_b_4 = b_4;
  assign f_u_arr_mul8_and_0_4_y0 = f_u_arr_mul8_and_0_4_a_0 & f_u_arr_mul8_and_0_4_b_4;
  assign f_u_arr_mul8_ha_0_4_f_u_arr_mul8_and_0_4_y0 = f_u_arr_mul8_and_0_4_y0;
  assign f_u_arr_mul8_ha_0_4_f_u_arr_mul8_fa_1_3_y2 = f_u_arr_mul8_fa_1_3_y2;
  assign f_u_arr_mul8_ha_0_4_y0 = f_u_arr_mul8_ha_0_4_f_u_arr_mul8_and_0_4_y0 ^ f_u_arr_mul8_ha_0_4_f_u_arr_mul8_fa_1_3_y2;
  assign f_u_arr_mul8_ha_0_4_y1 = f_u_arr_mul8_ha_0_4_f_u_arr_mul8_and_0_4_y0 & f_u_arr_mul8_ha_0_4_f_u_arr_mul8_fa_1_3_y2;
  assign f_u_arr_mul8_and_1_4_a_1 = a_1;
  assign f_u_arr_mul8_and_1_4_b_4 = b_4;
  assign f_u_arr_mul8_and_1_4_y0 = f_u_arr_mul8_and_1_4_a_1 & f_u_arr_mul8_and_1_4_b_4;
  assign f_u_arr_mul8_fa_1_4_f_u_arr_mul8_and_1_4_y0 = f_u_arr_mul8_and_1_4_y0;
  assign f_u_arr_mul8_fa_1_4_f_u_arr_mul8_fa_2_3_y2 = f_u_arr_mul8_fa_2_3_y2;
  assign f_u_arr_mul8_fa_1_4_f_u_arr_mul8_ha_0_4_y1 = f_u_arr_mul8_ha_0_4_y1;
  assign f_u_arr_mul8_fa_1_4_y0 = f_u_arr_mul8_fa_1_4_f_u_arr_mul8_and_1_4_y0 ^ f_u_arr_mul8_fa_1_4_f_u_arr_mul8_fa_2_3_y2;
  assign f_u_arr_mul8_fa_1_4_y1 = f_u_arr_mul8_fa_1_4_f_u_arr_mul8_and_1_4_y0 & f_u_arr_mul8_fa_1_4_f_u_arr_mul8_fa_2_3_y2;
  assign f_u_arr_mul8_fa_1_4_y2 = f_u_arr_mul8_fa_1_4_y0 ^ f_u_arr_mul8_fa_1_4_f_u_arr_mul8_ha_0_4_y1;
  assign f_u_arr_mul8_fa_1_4_y3 = f_u_arr_mul8_fa_1_4_y0 & f_u_arr_mul8_fa_1_4_f_u_arr_mul8_ha_0_4_y1;
  assign f_u_arr_mul8_fa_1_4_y4 = f_u_arr_mul8_fa_1_4_y1 | f_u_arr_mul8_fa_1_4_y3;
  assign f_u_arr_mul8_and_2_4_a_2 = a_2;
  assign f_u_arr_mul8_and_2_4_b_4 = b_4;
  assign f_u_arr_mul8_and_2_4_y0 = f_u_arr_mul8_and_2_4_a_2 & f_u_arr_mul8_and_2_4_b_4;
  assign f_u_arr_mul8_fa_2_4_f_u_arr_mul8_and_2_4_y0 = f_u_arr_mul8_and_2_4_y0;
  assign f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_3_3_y2 = f_u_arr_mul8_fa_3_3_y2;
  assign f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_1_4_y4 = f_u_arr_mul8_fa_1_4_y4;
  assign f_u_arr_mul8_fa_2_4_y0 = f_u_arr_mul8_fa_2_4_f_u_arr_mul8_and_2_4_y0 ^ f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_3_3_y2;
  assign f_u_arr_mul8_fa_2_4_y1 = f_u_arr_mul8_fa_2_4_f_u_arr_mul8_and_2_4_y0 & f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_3_3_y2;
  assign f_u_arr_mul8_fa_2_4_y2 = f_u_arr_mul8_fa_2_4_y0 ^ f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_1_4_y4;
  assign f_u_arr_mul8_fa_2_4_y3 = f_u_arr_mul8_fa_2_4_y0 & f_u_arr_mul8_fa_2_4_f_u_arr_mul8_fa_1_4_y4;
  assign f_u_arr_mul8_fa_2_4_y4 = f_u_arr_mul8_fa_2_4_y1 | f_u_arr_mul8_fa_2_4_y3;
  assign f_u_arr_mul8_and_3_4_a_3 = a_3;
  assign f_u_arr_mul8_and_3_4_b_4 = b_4;
  assign f_u_arr_mul8_and_3_4_y0 = f_u_arr_mul8_and_3_4_a_3 & f_u_arr_mul8_and_3_4_b_4;
  assign f_u_arr_mul8_fa_3_4_f_u_arr_mul8_and_3_4_y0 = f_u_arr_mul8_and_3_4_y0;
  assign f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_4_3_y2 = f_u_arr_mul8_fa_4_3_y2;
  assign f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_2_4_y4 = f_u_arr_mul8_fa_2_4_y4;
  assign f_u_arr_mul8_fa_3_4_y0 = f_u_arr_mul8_fa_3_4_f_u_arr_mul8_and_3_4_y0 ^ f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_4_3_y2;
  assign f_u_arr_mul8_fa_3_4_y1 = f_u_arr_mul8_fa_3_4_f_u_arr_mul8_and_3_4_y0 & f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_4_3_y2;
  assign f_u_arr_mul8_fa_3_4_y2 = f_u_arr_mul8_fa_3_4_y0 ^ f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_2_4_y4;
  assign f_u_arr_mul8_fa_3_4_y3 = f_u_arr_mul8_fa_3_4_y0 & f_u_arr_mul8_fa_3_4_f_u_arr_mul8_fa_2_4_y4;
  assign f_u_arr_mul8_fa_3_4_y4 = f_u_arr_mul8_fa_3_4_y1 | f_u_arr_mul8_fa_3_4_y3;
  assign f_u_arr_mul8_and_4_4_a_4 = a_4;
  assign f_u_arr_mul8_and_4_4_b_4 = b_4;
  assign f_u_arr_mul8_and_4_4_y0 = f_u_arr_mul8_and_4_4_a_4 & f_u_arr_mul8_and_4_4_b_4;
  assign f_u_arr_mul8_fa_4_4_f_u_arr_mul8_and_4_4_y0 = f_u_arr_mul8_and_4_4_y0;
  assign f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_5_3_y2 = f_u_arr_mul8_fa_5_3_y2;
  assign f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_3_4_y4 = f_u_arr_mul8_fa_3_4_y4;
  assign f_u_arr_mul8_fa_4_4_y0 = f_u_arr_mul8_fa_4_4_f_u_arr_mul8_and_4_4_y0 ^ f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_5_3_y2;
  assign f_u_arr_mul8_fa_4_4_y1 = f_u_arr_mul8_fa_4_4_f_u_arr_mul8_and_4_4_y0 & f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_5_3_y2;
  assign f_u_arr_mul8_fa_4_4_y2 = f_u_arr_mul8_fa_4_4_y0 ^ f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_3_4_y4;
  assign f_u_arr_mul8_fa_4_4_y3 = f_u_arr_mul8_fa_4_4_y0 & f_u_arr_mul8_fa_4_4_f_u_arr_mul8_fa_3_4_y4;
  assign f_u_arr_mul8_fa_4_4_y4 = f_u_arr_mul8_fa_4_4_y1 | f_u_arr_mul8_fa_4_4_y3;
  assign f_u_arr_mul8_and_5_4_a_5 = a_5;
  assign f_u_arr_mul8_and_5_4_b_4 = b_4;
  assign f_u_arr_mul8_and_5_4_y0 = f_u_arr_mul8_and_5_4_a_5 & f_u_arr_mul8_and_5_4_b_4;
  assign f_u_arr_mul8_fa_5_4_f_u_arr_mul8_and_5_4_y0 = f_u_arr_mul8_and_5_4_y0;
  assign f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_6_3_y2 = f_u_arr_mul8_fa_6_3_y2;
  assign f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_4_4_y4 = f_u_arr_mul8_fa_4_4_y4;
  assign f_u_arr_mul8_fa_5_4_y0 = f_u_arr_mul8_fa_5_4_f_u_arr_mul8_and_5_4_y0 ^ f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_6_3_y2;
  assign f_u_arr_mul8_fa_5_4_y1 = f_u_arr_mul8_fa_5_4_f_u_arr_mul8_and_5_4_y0 & f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_6_3_y2;
  assign f_u_arr_mul8_fa_5_4_y2 = f_u_arr_mul8_fa_5_4_y0 ^ f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_4_4_y4;
  assign f_u_arr_mul8_fa_5_4_y3 = f_u_arr_mul8_fa_5_4_y0 & f_u_arr_mul8_fa_5_4_f_u_arr_mul8_fa_4_4_y4;
  assign f_u_arr_mul8_fa_5_4_y4 = f_u_arr_mul8_fa_5_4_y1 | f_u_arr_mul8_fa_5_4_y3;
  assign f_u_arr_mul8_and_6_4_a_6 = a_6;
  assign f_u_arr_mul8_and_6_4_b_4 = b_4;
  assign f_u_arr_mul8_and_6_4_y0 = f_u_arr_mul8_and_6_4_a_6 & f_u_arr_mul8_and_6_4_b_4;
  assign f_u_arr_mul8_fa_6_4_f_u_arr_mul8_and_6_4_y0 = f_u_arr_mul8_and_6_4_y0;
  assign f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_7_3_y2 = f_u_arr_mul8_fa_7_3_y2;
  assign f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_5_4_y4 = f_u_arr_mul8_fa_5_4_y4;
  assign f_u_arr_mul8_fa_6_4_y0 = f_u_arr_mul8_fa_6_4_f_u_arr_mul8_and_6_4_y0 ^ f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_7_3_y2;
  assign f_u_arr_mul8_fa_6_4_y1 = f_u_arr_mul8_fa_6_4_f_u_arr_mul8_and_6_4_y0 & f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_7_3_y2;
  assign f_u_arr_mul8_fa_6_4_y2 = f_u_arr_mul8_fa_6_4_y0 ^ f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_5_4_y4;
  assign f_u_arr_mul8_fa_6_4_y3 = f_u_arr_mul8_fa_6_4_y0 & f_u_arr_mul8_fa_6_4_f_u_arr_mul8_fa_5_4_y4;
  assign f_u_arr_mul8_fa_6_4_y4 = f_u_arr_mul8_fa_6_4_y1 | f_u_arr_mul8_fa_6_4_y3;
  assign f_u_arr_mul8_and_7_4_a_7 = a_7;
  assign f_u_arr_mul8_and_7_4_b_4 = b_4;
  assign f_u_arr_mul8_and_7_4_y0 = f_u_arr_mul8_and_7_4_a_7 & f_u_arr_mul8_and_7_4_b_4;
  assign f_u_arr_mul8_fa_7_4_f_u_arr_mul8_and_7_4_y0 = f_u_arr_mul8_and_7_4_y0;
  assign f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_7_3_y4 = f_u_arr_mul8_fa_7_3_y4;
  assign f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_6_4_y4 = f_u_arr_mul8_fa_6_4_y4;
  assign f_u_arr_mul8_fa_7_4_y0 = f_u_arr_mul8_fa_7_4_f_u_arr_mul8_and_7_4_y0 ^ f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_7_3_y4;
  assign f_u_arr_mul8_fa_7_4_y1 = f_u_arr_mul8_fa_7_4_f_u_arr_mul8_and_7_4_y0 & f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_7_3_y4;
  assign f_u_arr_mul8_fa_7_4_y2 = f_u_arr_mul8_fa_7_4_y0 ^ f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_6_4_y4;
  assign f_u_arr_mul8_fa_7_4_y3 = f_u_arr_mul8_fa_7_4_y0 & f_u_arr_mul8_fa_7_4_f_u_arr_mul8_fa_6_4_y4;
  assign f_u_arr_mul8_fa_7_4_y4 = f_u_arr_mul8_fa_7_4_y1 | f_u_arr_mul8_fa_7_4_y3;
  assign f_u_arr_mul8_and_0_5_a_0 = a_0;
  assign f_u_arr_mul8_and_0_5_b_5 = b_5;
  assign f_u_arr_mul8_and_0_5_y0 = f_u_arr_mul8_and_0_5_a_0 & f_u_arr_mul8_and_0_5_b_5;
  assign f_u_arr_mul8_ha_0_5_f_u_arr_mul8_and_0_5_y0 = f_u_arr_mul8_and_0_5_y0;
  assign f_u_arr_mul8_ha_0_5_f_u_arr_mul8_fa_1_4_y2 = f_u_arr_mul8_fa_1_4_y2;
  assign f_u_arr_mul8_ha_0_5_y0 = f_u_arr_mul8_ha_0_5_f_u_arr_mul8_and_0_5_y0 ^ f_u_arr_mul8_ha_0_5_f_u_arr_mul8_fa_1_4_y2;
  assign f_u_arr_mul8_ha_0_5_y1 = f_u_arr_mul8_ha_0_5_f_u_arr_mul8_and_0_5_y0 & f_u_arr_mul8_ha_0_5_f_u_arr_mul8_fa_1_4_y2;
  assign f_u_arr_mul8_and_1_5_a_1 = a_1;
  assign f_u_arr_mul8_and_1_5_b_5 = b_5;
  assign f_u_arr_mul8_and_1_5_y0 = f_u_arr_mul8_and_1_5_a_1 & f_u_arr_mul8_and_1_5_b_5;
  assign f_u_arr_mul8_fa_1_5_f_u_arr_mul8_and_1_5_y0 = f_u_arr_mul8_and_1_5_y0;
  assign f_u_arr_mul8_fa_1_5_f_u_arr_mul8_fa_2_4_y2 = f_u_arr_mul8_fa_2_4_y2;
  assign f_u_arr_mul8_fa_1_5_f_u_arr_mul8_ha_0_5_y1 = f_u_arr_mul8_ha_0_5_y1;
  assign f_u_arr_mul8_fa_1_5_y0 = f_u_arr_mul8_fa_1_5_f_u_arr_mul8_and_1_5_y0 ^ f_u_arr_mul8_fa_1_5_f_u_arr_mul8_fa_2_4_y2;
  assign f_u_arr_mul8_fa_1_5_y1 = f_u_arr_mul8_fa_1_5_f_u_arr_mul8_and_1_5_y0 & f_u_arr_mul8_fa_1_5_f_u_arr_mul8_fa_2_4_y2;
  assign f_u_arr_mul8_fa_1_5_y2 = f_u_arr_mul8_fa_1_5_y0 ^ f_u_arr_mul8_fa_1_5_f_u_arr_mul8_ha_0_5_y1;
  assign f_u_arr_mul8_fa_1_5_y3 = f_u_arr_mul8_fa_1_5_y0 & f_u_arr_mul8_fa_1_5_f_u_arr_mul8_ha_0_5_y1;
  assign f_u_arr_mul8_fa_1_5_y4 = f_u_arr_mul8_fa_1_5_y1 | f_u_arr_mul8_fa_1_5_y3;
  assign f_u_arr_mul8_and_2_5_a_2 = a_2;
  assign f_u_arr_mul8_and_2_5_b_5 = b_5;
  assign f_u_arr_mul8_and_2_5_y0 = f_u_arr_mul8_and_2_5_a_2 & f_u_arr_mul8_and_2_5_b_5;
  assign f_u_arr_mul8_fa_2_5_f_u_arr_mul8_and_2_5_y0 = f_u_arr_mul8_and_2_5_y0;
  assign f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_3_4_y2 = f_u_arr_mul8_fa_3_4_y2;
  assign f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_1_5_y4 = f_u_arr_mul8_fa_1_5_y4;
  assign f_u_arr_mul8_fa_2_5_y0 = f_u_arr_mul8_fa_2_5_f_u_arr_mul8_and_2_5_y0 ^ f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_3_4_y2;
  assign f_u_arr_mul8_fa_2_5_y1 = f_u_arr_mul8_fa_2_5_f_u_arr_mul8_and_2_5_y0 & f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_3_4_y2;
  assign f_u_arr_mul8_fa_2_5_y2 = f_u_arr_mul8_fa_2_5_y0 ^ f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_1_5_y4;
  assign f_u_arr_mul8_fa_2_5_y3 = f_u_arr_mul8_fa_2_5_y0 & f_u_arr_mul8_fa_2_5_f_u_arr_mul8_fa_1_5_y4;
  assign f_u_arr_mul8_fa_2_5_y4 = f_u_arr_mul8_fa_2_5_y1 | f_u_arr_mul8_fa_2_5_y3;
  assign f_u_arr_mul8_and_3_5_a_3 = a_3;
  assign f_u_arr_mul8_and_3_5_b_5 = b_5;
  assign f_u_arr_mul8_and_3_5_y0 = f_u_arr_mul8_and_3_5_a_3 & f_u_arr_mul8_and_3_5_b_5;
  assign f_u_arr_mul8_fa_3_5_f_u_arr_mul8_and_3_5_y0 = f_u_arr_mul8_and_3_5_y0;
  assign f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_4_4_y2 = f_u_arr_mul8_fa_4_4_y2;
  assign f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_2_5_y4 = f_u_arr_mul8_fa_2_5_y4;
  assign f_u_arr_mul8_fa_3_5_y0 = f_u_arr_mul8_fa_3_5_f_u_arr_mul8_and_3_5_y0 ^ f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_4_4_y2;
  assign f_u_arr_mul8_fa_3_5_y1 = f_u_arr_mul8_fa_3_5_f_u_arr_mul8_and_3_5_y0 & f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_4_4_y2;
  assign f_u_arr_mul8_fa_3_5_y2 = f_u_arr_mul8_fa_3_5_y0 ^ f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_2_5_y4;
  assign f_u_arr_mul8_fa_3_5_y3 = f_u_arr_mul8_fa_3_5_y0 & f_u_arr_mul8_fa_3_5_f_u_arr_mul8_fa_2_5_y4;
  assign f_u_arr_mul8_fa_3_5_y4 = f_u_arr_mul8_fa_3_5_y1 | f_u_arr_mul8_fa_3_5_y3;
  assign f_u_arr_mul8_and_4_5_a_4 = a_4;
  assign f_u_arr_mul8_and_4_5_b_5 = b_5;
  assign f_u_arr_mul8_and_4_5_y0 = f_u_arr_mul8_and_4_5_a_4 & f_u_arr_mul8_and_4_5_b_5;
  assign f_u_arr_mul8_fa_4_5_f_u_arr_mul8_and_4_5_y0 = f_u_arr_mul8_and_4_5_y0;
  assign f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_5_4_y2 = f_u_arr_mul8_fa_5_4_y2;
  assign f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_3_5_y4 = f_u_arr_mul8_fa_3_5_y4;
  assign f_u_arr_mul8_fa_4_5_y0 = f_u_arr_mul8_fa_4_5_f_u_arr_mul8_and_4_5_y0 ^ f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_5_4_y2;
  assign f_u_arr_mul8_fa_4_5_y1 = f_u_arr_mul8_fa_4_5_f_u_arr_mul8_and_4_5_y0 & f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_5_4_y2;
  assign f_u_arr_mul8_fa_4_5_y2 = f_u_arr_mul8_fa_4_5_y0 ^ f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_3_5_y4;
  assign f_u_arr_mul8_fa_4_5_y3 = f_u_arr_mul8_fa_4_5_y0 & f_u_arr_mul8_fa_4_5_f_u_arr_mul8_fa_3_5_y4;
  assign f_u_arr_mul8_fa_4_5_y4 = f_u_arr_mul8_fa_4_5_y1 | f_u_arr_mul8_fa_4_5_y3;
  assign f_u_arr_mul8_and_5_5_a_5 = a_5;
  assign f_u_arr_mul8_and_5_5_b_5 = b_5;
  assign f_u_arr_mul8_and_5_5_y0 = f_u_arr_mul8_and_5_5_a_5 & f_u_arr_mul8_and_5_5_b_5;
  assign f_u_arr_mul8_fa_5_5_f_u_arr_mul8_and_5_5_y0 = f_u_arr_mul8_and_5_5_y0;
  assign f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_6_4_y2 = f_u_arr_mul8_fa_6_4_y2;
  assign f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_4_5_y4 = f_u_arr_mul8_fa_4_5_y4;
  assign f_u_arr_mul8_fa_5_5_y0 = f_u_arr_mul8_fa_5_5_f_u_arr_mul8_and_5_5_y0 ^ f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_6_4_y2;
  assign f_u_arr_mul8_fa_5_5_y1 = f_u_arr_mul8_fa_5_5_f_u_arr_mul8_and_5_5_y0 & f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_6_4_y2;
  assign f_u_arr_mul8_fa_5_5_y2 = f_u_arr_mul8_fa_5_5_y0 ^ f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_4_5_y4;
  assign f_u_arr_mul8_fa_5_5_y3 = f_u_arr_mul8_fa_5_5_y0 & f_u_arr_mul8_fa_5_5_f_u_arr_mul8_fa_4_5_y4;
  assign f_u_arr_mul8_fa_5_5_y4 = f_u_arr_mul8_fa_5_5_y1 | f_u_arr_mul8_fa_5_5_y3;
  assign f_u_arr_mul8_and_6_5_a_6 = a_6;
  assign f_u_arr_mul8_and_6_5_b_5 = b_5;
  assign f_u_arr_mul8_and_6_5_y0 = f_u_arr_mul8_and_6_5_a_6 & f_u_arr_mul8_and_6_5_b_5;
  assign f_u_arr_mul8_fa_6_5_f_u_arr_mul8_and_6_5_y0 = f_u_arr_mul8_and_6_5_y0;
  assign f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_7_4_y2 = f_u_arr_mul8_fa_7_4_y2;
  assign f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_5_5_y4 = f_u_arr_mul8_fa_5_5_y4;
  assign f_u_arr_mul8_fa_6_5_y0 = f_u_arr_mul8_fa_6_5_f_u_arr_mul8_and_6_5_y0 ^ f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_7_4_y2;
  assign f_u_arr_mul8_fa_6_5_y1 = f_u_arr_mul8_fa_6_5_f_u_arr_mul8_and_6_5_y0 & f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_7_4_y2;
  assign f_u_arr_mul8_fa_6_5_y2 = f_u_arr_mul8_fa_6_5_y0 ^ f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_5_5_y4;
  assign f_u_arr_mul8_fa_6_5_y3 = f_u_arr_mul8_fa_6_5_y0 & f_u_arr_mul8_fa_6_5_f_u_arr_mul8_fa_5_5_y4;
  assign f_u_arr_mul8_fa_6_5_y4 = f_u_arr_mul8_fa_6_5_y1 | f_u_arr_mul8_fa_6_5_y3;
  assign f_u_arr_mul8_and_7_5_a_7 = a_7;
  assign f_u_arr_mul8_and_7_5_b_5 = b_5;
  assign f_u_arr_mul8_and_7_5_y0 = f_u_arr_mul8_and_7_5_a_7 & f_u_arr_mul8_and_7_5_b_5;
  assign f_u_arr_mul8_fa_7_5_f_u_arr_mul8_and_7_5_y0 = f_u_arr_mul8_and_7_5_y0;
  assign f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_7_4_y4 = f_u_arr_mul8_fa_7_4_y4;
  assign f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_6_5_y4 = f_u_arr_mul8_fa_6_5_y4;
  assign f_u_arr_mul8_fa_7_5_y0 = f_u_arr_mul8_fa_7_5_f_u_arr_mul8_and_7_5_y0 ^ f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_7_4_y4;
  assign f_u_arr_mul8_fa_7_5_y1 = f_u_arr_mul8_fa_7_5_f_u_arr_mul8_and_7_5_y0 & f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_7_4_y4;
  assign f_u_arr_mul8_fa_7_5_y2 = f_u_arr_mul8_fa_7_5_y0 ^ f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_6_5_y4;
  assign f_u_arr_mul8_fa_7_5_y3 = f_u_arr_mul8_fa_7_5_y0 & f_u_arr_mul8_fa_7_5_f_u_arr_mul8_fa_6_5_y4;
  assign f_u_arr_mul8_fa_7_5_y4 = f_u_arr_mul8_fa_7_5_y1 | f_u_arr_mul8_fa_7_5_y3;
  assign f_u_arr_mul8_and_0_6_a_0 = a_0;
  assign f_u_arr_mul8_and_0_6_b_6 = b_6;
  assign f_u_arr_mul8_and_0_6_y0 = f_u_arr_mul8_and_0_6_a_0 & f_u_arr_mul8_and_0_6_b_6;
  assign f_u_arr_mul8_ha_0_6_f_u_arr_mul8_and_0_6_y0 = f_u_arr_mul8_and_0_6_y0;
  assign f_u_arr_mul8_ha_0_6_f_u_arr_mul8_fa_1_5_y2 = f_u_arr_mul8_fa_1_5_y2;
  assign f_u_arr_mul8_ha_0_6_y0 = f_u_arr_mul8_ha_0_6_f_u_arr_mul8_and_0_6_y0 ^ f_u_arr_mul8_ha_0_6_f_u_arr_mul8_fa_1_5_y2;
  assign f_u_arr_mul8_ha_0_6_y1 = f_u_arr_mul8_ha_0_6_f_u_arr_mul8_and_0_6_y0 & f_u_arr_mul8_ha_0_6_f_u_arr_mul8_fa_1_5_y2;
  assign f_u_arr_mul8_and_1_6_a_1 = a_1;
  assign f_u_arr_mul8_and_1_6_b_6 = b_6;
  assign f_u_arr_mul8_and_1_6_y0 = f_u_arr_mul8_and_1_6_a_1 & f_u_arr_mul8_and_1_6_b_6;
  assign f_u_arr_mul8_fa_1_6_f_u_arr_mul8_and_1_6_y0 = f_u_arr_mul8_and_1_6_y0;
  assign f_u_arr_mul8_fa_1_6_f_u_arr_mul8_fa_2_5_y2 = f_u_arr_mul8_fa_2_5_y2;
  assign f_u_arr_mul8_fa_1_6_f_u_arr_mul8_ha_0_6_y1 = f_u_arr_mul8_ha_0_6_y1;
  assign f_u_arr_mul8_fa_1_6_y0 = f_u_arr_mul8_fa_1_6_f_u_arr_mul8_and_1_6_y0 ^ f_u_arr_mul8_fa_1_6_f_u_arr_mul8_fa_2_5_y2;
  assign f_u_arr_mul8_fa_1_6_y1 = f_u_arr_mul8_fa_1_6_f_u_arr_mul8_and_1_6_y0 & f_u_arr_mul8_fa_1_6_f_u_arr_mul8_fa_2_5_y2;
  assign f_u_arr_mul8_fa_1_6_y2 = f_u_arr_mul8_fa_1_6_y0 ^ f_u_arr_mul8_fa_1_6_f_u_arr_mul8_ha_0_6_y1;
  assign f_u_arr_mul8_fa_1_6_y3 = f_u_arr_mul8_fa_1_6_y0 & f_u_arr_mul8_fa_1_6_f_u_arr_mul8_ha_0_6_y1;
  assign f_u_arr_mul8_fa_1_6_y4 = f_u_arr_mul8_fa_1_6_y1 | f_u_arr_mul8_fa_1_6_y3;
  assign f_u_arr_mul8_and_2_6_a_2 = a_2;
  assign f_u_arr_mul8_and_2_6_b_6 = b_6;
  assign f_u_arr_mul8_and_2_6_y0 = f_u_arr_mul8_and_2_6_a_2 & f_u_arr_mul8_and_2_6_b_6;
  assign f_u_arr_mul8_fa_2_6_f_u_arr_mul8_and_2_6_y0 = f_u_arr_mul8_and_2_6_y0;
  assign f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_3_5_y2 = f_u_arr_mul8_fa_3_5_y2;
  assign f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_1_6_y4 = f_u_arr_mul8_fa_1_6_y4;
  assign f_u_arr_mul8_fa_2_6_y0 = f_u_arr_mul8_fa_2_6_f_u_arr_mul8_and_2_6_y0 ^ f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_3_5_y2;
  assign f_u_arr_mul8_fa_2_6_y1 = f_u_arr_mul8_fa_2_6_f_u_arr_mul8_and_2_6_y0 & f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_3_5_y2;
  assign f_u_arr_mul8_fa_2_6_y2 = f_u_arr_mul8_fa_2_6_y0 ^ f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_1_6_y4;
  assign f_u_arr_mul8_fa_2_6_y3 = f_u_arr_mul8_fa_2_6_y0 & f_u_arr_mul8_fa_2_6_f_u_arr_mul8_fa_1_6_y4;
  assign f_u_arr_mul8_fa_2_6_y4 = f_u_arr_mul8_fa_2_6_y1 | f_u_arr_mul8_fa_2_6_y3;
  assign f_u_arr_mul8_and_3_6_a_3 = a_3;
  assign f_u_arr_mul8_and_3_6_b_6 = b_6;
  assign f_u_arr_mul8_and_3_6_y0 = f_u_arr_mul8_and_3_6_a_3 & f_u_arr_mul8_and_3_6_b_6;
  assign f_u_arr_mul8_fa_3_6_f_u_arr_mul8_and_3_6_y0 = f_u_arr_mul8_and_3_6_y0;
  assign f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_4_5_y2 = f_u_arr_mul8_fa_4_5_y2;
  assign f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_2_6_y4 = f_u_arr_mul8_fa_2_6_y4;
  assign f_u_arr_mul8_fa_3_6_y0 = f_u_arr_mul8_fa_3_6_f_u_arr_mul8_and_3_6_y0 ^ f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_4_5_y2;
  assign f_u_arr_mul8_fa_3_6_y1 = f_u_arr_mul8_fa_3_6_f_u_arr_mul8_and_3_6_y0 & f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_4_5_y2;
  assign f_u_arr_mul8_fa_3_6_y2 = f_u_arr_mul8_fa_3_6_y0 ^ f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_2_6_y4;
  assign f_u_arr_mul8_fa_3_6_y3 = f_u_arr_mul8_fa_3_6_y0 & f_u_arr_mul8_fa_3_6_f_u_arr_mul8_fa_2_6_y4;
  assign f_u_arr_mul8_fa_3_6_y4 = f_u_arr_mul8_fa_3_6_y1 | f_u_arr_mul8_fa_3_6_y3;
  assign f_u_arr_mul8_and_4_6_a_4 = a_4;
  assign f_u_arr_mul8_and_4_6_b_6 = b_6;
  assign f_u_arr_mul8_and_4_6_y0 = f_u_arr_mul8_and_4_6_a_4 & f_u_arr_mul8_and_4_6_b_6;
  assign f_u_arr_mul8_fa_4_6_f_u_arr_mul8_and_4_6_y0 = f_u_arr_mul8_and_4_6_y0;
  assign f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_5_5_y2 = f_u_arr_mul8_fa_5_5_y2;
  assign f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_3_6_y4 = f_u_arr_mul8_fa_3_6_y4;
  assign f_u_arr_mul8_fa_4_6_y0 = f_u_arr_mul8_fa_4_6_f_u_arr_mul8_and_4_6_y0 ^ f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_5_5_y2;
  assign f_u_arr_mul8_fa_4_6_y1 = f_u_arr_mul8_fa_4_6_f_u_arr_mul8_and_4_6_y0 & f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_5_5_y2;
  assign f_u_arr_mul8_fa_4_6_y2 = f_u_arr_mul8_fa_4_6_y0 ^ f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_3_6_y4;
  assign f_u_arr_mul8_fa_4_6_y3 = f_u_arr_mul8_fa_4_6_y0 & f_u_arr_mul8_fa_4_6_f_u_arr_mul8_fa_3_6_y4;
  assign f_u_arr_mul8_fa_4_6_y4 = f_u_arr_mul8_fa_4_6_y1 | f_u_arr_mul8_fa_4_6_y3;
  assign f_u_arr_mul8_and_5_6_a_5 = a_5;
  assign f_u_arr_mul8_and_5_6_b_6 = b_6;
  assign f_u_arr_mul8_and_5_6_y0 = f_u_arr_mul8_and_5_6_a_5 & f_u_arr_mul8_and_5_6_b_6;
  assign f_u_arr_mul8_fa_5_6_f_u_arr_mul8_and_5_6_y0 = f_u_arr_mul8_and_5_6_y0;
  assign f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_6_5_y2 = f_u_arr_mul8_fa_6_5_y2;
  assign f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_4_6_y4 = f_u_arr_mul8_fa_4_6_y4;
  assign f_u_arr_mul8_fa_5_6_y0 = f_u_arr_mul8_fa_5_6_f_u_arr_mul8_and_5_6_y0 ^ f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_6_5_y2;
  assign f_u_arr_mul8_fa_5_6_y1 = f_u_arr_mul8_fa_5_6_f_u_arr_mul8_and_5_6_y0 & f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_6_5_y2;
  assign f_u_arr_mul8_fa_5_6_y2 = f_u_arr_mul8_fa_5_6_y0 ^ f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_4_6_y4;
  assign f_u_arr_mul8_fa_5_6_y3 = f_u_arr_mul8_fa_5_6_y0 & f_u_arr_mul8_fa_5_6_f_u_arr_mul8_fa_4_6_y4;
  assign f_u_arr_mul8_fa_5_6_y4 = f_u_arr_mul8_fa_5_6_y1 | f_u_arr_mul8_fa_5_6_y3;
  assign f_u_arr_mul8_and_6_6_a_6 = a_6;
  assign f_u_arr_mul8_and_6_6_b_6 = b_6;
  assign f_u_arr_mul8_and_6_6_y0 = f_u_arr_mul8_and_6_6_a_6 & f_u_arr_mul8_and_6_6_b_6;
  assign f_u_arr_mul8_fa_6_6_f_u_arr_mul8_and_6_6_y0 = f_u_arr_mul8_and_6_6_y0;
  assign f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_7_5_y2 = f_u_arr_mul8_fa_7_5_y2;
  assign f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_5_6_y4 = f_u_arr_mul8_fa_5_6_y4;
  assign f_u_arr_mul8_fa_6_6_y0 = f_u_arr_mul8_fa_6_6_f_u_arr_mul8_and_6_6_y0 ^ f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_7_5_y2;
  assign f_u_arr_mul8_fa_6_6_y1 = f_u_arr_mul8_fa_6_6_f_u_arr_mul8_and_6_6_y0 & f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_7_5_y2;
  assign f_u_arr_mul8_fa_6_6_y2 = f_u_arr_mul8_fa_6_6_y0 ^ f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_5_6_y4;
  assign f_u_arr_mul8_fa_6_6_y3 = f_u_arr_mul8_fa_6_6_y0 & f_u_arr_mul8_fa_6_6_f_u_arr_mul8_fa_5_6_y4;
  assign f_u_arr_mul8_fa_6_6_y4 = f_u_arr_mul8_fa_6_6_y1 | f_u_arr_mul8_fa_6_6_y3;
  assign f_u_arr_mul8_and_7_6_a_7 = a_7;
  assign f_u_arr_mul8_and_7_6_b_6 = b_6;
  assign f_u_arr_mul8_and_7_6_y0 = f_u_arr_mul8_and_7_6_a_7 & f_u_arr_mul8_and_7_6_b_6;
  assign f_u_arr_mul8_fa_7_6_f_u_arr_mul8_and_7_6_y0 = f_u_arr_mul8_and_7_6_y0;
  assign f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_7_5_y4 = f_u_arr_mul8_fa_7_5_y4;
  assign f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_6_6_y4 = f_u_arr_mul8_fa_6_6_y4;
  assign f_u_arr_mul8_fa_7_6_y0 = f_u_arr_mul8_fa_7_6_f_u_arr_mul8_and_7_6_y0 ^ f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_7_5_y4;
  assign f_u_arr_mul8_fa_7_6_y1 = f_u_arr_mul8_fa_7_6_f_u_arr_mul8_and_7_6_y0 & f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_7_5_y4;
  assign f_u_arr_mul8_fa_7_6_y2 = f_u_arr_mul8_fa_7_6_y0 ^ f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_6_6_y4;
  assign f_u_arr_mul8_fa_7_6_y3 = f_u_arr_mul8_fa_7_6_y0 & f_u_arr_mul8_fa_7_6_f_u_arr_mul8_fa_6_6_y4;
  assign f_u_arr_mul8_fa_7_6_y4 = f_u_arr_mul8_fa_7_6_y1 | f_u_arr_mul8_fa_7_6_y3;
  assign f_u_arr_mul8_and_0_7_a_0 = a_0;
  assign f_u_arr_mul8_and_0_7_b_7 = b_7;
  assign f_u_arr_mul8_and_0_7_y0 = f_u_arr_mul8_and_0_7_a_0 & f_u_arr_mul8_and_0_7_b_7;
  assign f_u_arr_mul8_ha_0_7_f_u_arr_mul8_and_0_7_y0 = f_u_arr_mul8_and_0_7_y0;
  assign f_u_arr_mul8_ha_0_7_f_u_arr_mul8_fa_1_6_y2 = f_u_arr_mul8_fa_1_6_y2;
  assign f_u_arr_mul8_ha_0_7_y0 = f_u_arr_mul8_ha_0_7_f_u_arr_mul8_and_0_7_y0 ^ f_u_arr_mul8_ha_0_7_f_u_arr_mul8_fa_1_6_y2;
  assign f_u_arr_mul8_ha_0_7_y1 = f_u_arr_mul8_ha_0_7_f_u_arr_mul8_and_0_7_y0 & f_u_arr_mul8_ha_0_7_f_u_arr_mul8_fa_1_6_y2;
  assign f_u_arr_mul8_and_1_7_a_1 = a_1;
  assign f_u_arr_mul8_and_1_7_b_7 = b_7;
  assign f_u_arr_mul8_and_1_7_y0 = f_u_arr_mul8_and_1_7_a_1 & f_u_arr_mul8_and_1_7_b_7;
  assign f_u_arr_mul8_fa_1_7_f_u_arr_mul8_and_1_7_y0 = f_u_arr_mul8_and_1_7_y0;
  assign f_u_arr_mul8_fa_1_7_f_u_arr_mul8_fa_2_6_y2 = f_u_arr_mul8_fa_2_6_y2;
  assign f_u_arr_mul8_fa_1_7_f_u_arr_mul8_ha_0_7_y1 = f_u_arr_mul8_ha_0_7_y1;
  assign f_u_arr_mul8_fa_1_7_y0 = f_u_arr_mul8_fa_1_7_f_u_arr_mul8_and_1_7_y0 ^ f_u_arr_mul8_fa_1_7_f_u_arr_mul8_fa_2_6_y2;
  assign f_u_arr_mul8_fa_1_7_y1 = f_u_arr_mul8_fa_1_7_f_u_arr_mul8_and_1_7_y0 & f_u_arr_mul8_fa_1_7_f_u_arr_mul8_fa_2_6_y2;
  assign f_u_arr_mul8_fa_1_7_y2 = f_u_arr_mul8_fa_1_7_y0 ^ f_u_arr_mul8_fa_1_7_f_u_arr_mul8_ha_0_7_y1;
  assign f_u_arr_mul8_fa_1_7_y3 = f_u_arr_mul8_fa_1_7_y0 & f_u_arr_mul8_fa_1_7_f_u_arr_mul8_ha_0_7_y1;
  assign f_u_arr_mul8_fa_1_7_y4 = f_u_arr_mul8_fa_1_7_y1 | f_u_arr_mul8_fa_1_7_y3;
  assign f_u_arr_mul8_and_2_7_a_2 = a_2;
  assign f_u_arr_mul8_and_2_7_b_7 = b_7;
  assign f_u_arr_mul8_and_2_7_y0 = f_u_arr_mul8_and_2_7_a_2 & f_u_arr_mul8_and_2_7_b_7;
  assign f_u_arr_mul8_fa_2_7_f_u_arr_mul8_and_2_7_y0 = f_u_arr_mul8_and_2_7_y0;
  assign f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_3_6_y2 = f_u_arr_mul8_fa_3_6_y2;
  assign f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_1_7_y4 = f_u_arr_mul8_fa_1_7_y4;
  assign f_u_arr_mul8_fa_2_7_y0 = f_u_arr_mul8_fa_2_7_f_u_arr_mul8_and_2_7_y0 ^ f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_3_6_y2;
  assign f_u_arr_mul8_fa_2_7_y1 = f_u_arr_mul8_fa_2_7_f_u_arr_mul8_and_2_7_y0 & f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_3_6_y2;
  assign f_u_arr_mul8_fa_2_7_y2 = f_u_arr_mul8_fa_2_7_y0 ^ f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_1_7_y4;
  assign f_u_arr_mul8_fa_2_7_y3 = f_u_arr_mul8_fa_2_7_y0 & f_u_arr_mul8_fa_2_7_f_u_arr_mul8_fa_1_7_y4;
  assign f_u_arr_mul8_fa_2_7_y4 = f_u_arr_mul8_fa_2_7_y1 | f_u_arr_mul8_fa_2_7_y3;
  assign f_u_arr_mul8_and_3_7_a_3 = a_3;
  assign f_u_arr_mul8_and_3_7_b_7 = b_7;
  assign f_u_arr_mul8_and_3_7_y0 = f_u_arr_mul8_and_3_7_a_3 & f_u_arr_mul8_and_3_7_b_7;
  assign f_u_arr_mul8_fa_3_7_f_u_arr_mul8_and_3_7_y0 = f_u_arr_mul8_and_3_7_y0;
  assign f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_4_6_y2 = f_u_arr_mul8_fa_4_6_y2;
  assign f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_2_7_y4 = f_u_arr_mul8_fa_2_7_y4;
  assign f_u_arr_mul8_fa_3_7_y0 = f_u_arr_mul8_fa_3_7_f_u_arr_mul8_and_3_7_y0 ^ f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_4_6_y2;
  assign f_u_arr_mul8_fa_3_7_y1 = f_u_arr_mul8_fa_3_7_f_u_arr_mul8_and_3_7_y0 & f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_4_6_y2;
  assign f_u_arr_mul8_fa_3_7_y2 = f_u_arr_mul8_fa_3_7_y0 ^ f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_2_7_y4;
  assign f_u_arr_mul8_fa_3_7_y3 = f_u_arr_mul8_fa_3_7_y0 & f_u_arr_mul8_fa_3_7_f_u_arr_mul8_fa_2_7_y4;
  assign f_u_arr_mul8_fa_3_7_y4 = f_u_arr_mul8_fa_3_7_y1 | f_u_arr_mul8_fa_3_7_y3;
  assign f_u_arr_mul8_and_4_7_a_4 = a_4;
  assign f_u_arr_mul8_and_4_7_b_7 = b_7;
  assign f_u_arr_mul8_and_4_7_y0 = f_u_arr_mul8_and_4_7_a_4 & f_u_arr_mul8_and_4_7_b_7;
  assign f_u_arr_mul8_fa_4_7_f_u_arr_mul8_and_4_7_y0 = f_u_arr_mul8_and_4_7_y0;
  assign f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_5_6_y2 = f_u_arr_mul8_fa_5_6_y2;
  assign f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_3_7_y4 = f_u_arr_mul8_fa_3_7_y4;
  assign f_u_arr_mul8_fa_4_7_y0 = f_u_arr_mul8_fa_4_7_f_u_arr_mul8_and_4_7_y0 ^ f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_5_6_y2;
  assign f_u_arr_mul8_fa_4_7_y1 = f_u_arr_mul8_fa_4_7_f_u_arr_mul8_and_4_7_y0 & f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_5_6_y2;
  assign f_u_arr_mul8_fa_4_7_y2 = f_u_arr_mul8_fa_4_7_y0 ^ f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_3_7_y4;
  assign f_u_arr_mul8_fa_4_7_y3 = f_u_arr_mul8_fa_4_7_y0 & f_u_arr_mul8_fa_4_7_f_u_arr_mul8_fa_3_7_y4;
  assign f_u_arr_mul8_fa_4_7_y4 = f_u_arr_mul8_fa_4_7_y1 | f_u_arr_mul8_fa_4_7_y3;
  assign f_u_arr_mul8_and_5_7_a_5 = a_5;
  assign f_u_arr_mul8_and_5_7_b_7 = b_7;
  assign f_u_arr_mul8_and_5_7_y0 = f_u_arr_mul8_and_5_7_a_5 & f_u_arr_mul8_and_5_7_b_7;
  assign f_u_arr_mul8_fa_5_7_f_u_arr_mul8_and_5_7_y0 = f_u_arr_mul8_and_5_7_y0;
  assign f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_6_6_y2 = f_u_arr_mul8_fa_6_6_y2;
  assign f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_4_7_y4 = f_u_arr_mul8_fa_4_7_y4;
  assign f_u_arr_mul8_fa_5_7_y0 = f_u_arr_mul8_fa_5_7_f_u_arr_mul8_and_5_7_y0 ^ f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_6_6_y2;
  assign f_u_arr_mul8_fa_5_7_y1 = f_u_arr_mul8_fa_5_7_f_u_arr_mul8_and_5_7_y0 & f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_6_6_y2;
  assign f_u_arr_mul8_fa_5_7_y2 = f_u_arr_mul8_fa_5_7_y0 ^ f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_4_7_y4;
  assign f_u_arr_mul8_fa_5_7_y3 = f_u_arr_mul8_fa_5_7_y0 & f_u_arr_mul8_fa_5_7_f_u_arr_mul8_fa_4_7_y4;
  assign f_u_arr_mul8_fa_5_7_y4 = f_u_arr_mul8_fa_5_7_y1 | f_u_arr_mul8_fa_5_7_y3;
  assign f_u_arr_mul8_and_6_7_a_6 = a_6;
  assign f_u_arr_mul8_and_6_7_b_7 = b_7;
  assign f_u_arr_mul8_and_6_7_y0 = f_u_arr_mul8_and_6_7_a_6 & f_u_arr_mul8_and_6_7_b_7;
  assign f_u_arr_mul8_fa_6_7_f_u_arr_mul8_and_6_7_y0 = f_u_arr_mul8_and_6_7_y0;
  assign f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_7_6_y2 = f_u_arr_mul8_fa_7_6_y2;
  assign f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_5_7_y4 = f_u_arr_mul8_fa_5_7_y4;
  assign f_u_arr_mul8_fa_6_7_y0 = f_u_arr_mul8_fa_6_7_f_u_arr_mul8_and_6_7_y0 ^ f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_7_6_y2;
  assign f_u_arr_mul8_fa_6_7_y1 = f_u_arr_mul8_fa_6_7_f_u_arr_mul8_and_6_7_y0 & f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_7_6_y2;
  assign f_u_arr_mul8_fa_6_7_y2 = f_u_arr_mul8_fa_6_7_y0 ^ f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_5_7_y4;
  assign f_u_arr_mul8_fa_6_7_y3 = f_u_arr_mul8_fa_6_7_y0 & f_u_arr_mul8_fa_6_7_f_u_arr_mul8_fa_5_7_y4;
  assign f_u_arr_mul8_fa_6_7_y4 = f_u_arr_mul8_fa_6_7_y1 | f_u_arr_mul8_fa_6_7_y3;
  assign f_u_arr_mul8_and_7_7_a_7 = a_7;
  assign f_u_arr_mul8_and_7_7_b_7 = b_7;
  assign f_u_arr_mul8_and_7_7_y0 = f_u_arr_mul8_and_7_7_a_7 & f_u_arr_mul8_and_7_7_b_7;
  assign f_u_arr_mul8_fa_7_7_f_u_arr_mul8_and_7_7_y0 = f_u_arr_mul8_and_7_7_y0;
  assign f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_7_6_y4 = f_u_arr_mul8_fa_7_6_y4;
  assign f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_6_7_y4 = f_u_arr_mul8_fa_6_7_y4;
  assign f_u_arr_mul8_fa_7_7_y0 = f_u_arr_mul8_fa_7_7_f_u_arr_mul8_and_7_7_y0 ^ f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_7_6_y4;
  assign f_u_arr_mul8_fa_7_7_y1 = f_u_arr_mul8_fa_7_7_f_u_arr_mul8_and_7_7_y0 & f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_7_6_y4;
  assign f_u_arr_mul8_fa_7_7_y2 = f_u_arr_mul8_fa_7_7_y0 ^ f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_6_7_y4;
  assign f_u_arr_mul8_fa_7_7_y3 = f_u_arr_mul8_fa_7_7_y0 & f_u_arr_mul8_fa_7_7_f_u_arr_mul8_fa_6_7_y4;
  assign f_u_arr_mul8_fa_7_7_y4 = f_u_arr_mul8_fa_7_7_y1 | f_u_arr_mul8_fa_7_7_y3;

  assign out[0] = f_u_arr_mul8_and_0_0_y0;
  assign out[1] = f_u_arr_mul8_ha_0_1_y0;
  assign out[2] = f_u_arr_mul8_ha_0_2_y0;
  assign out[3] = f_u_arr_mul8_ha_0_3_y0;
  assign out[4] = f_u_arr_mul8_ha_0_4_y0;
  assign out[5] = f_u_arr_mul8_ha_0_5_y0;
  assign out[6] = f_u_arr_mul8_ha_0_6_y0;
  assign out[7] = f_u_arr_mul8_ha_0_7_y0;
  assign out[8] = f_u_arr_mul8_fa_1_7_y2;
  assign out[9] = f_u_arr_mul8_fa_2_7_y2;
  assign out[10] = f_u_arr_mul8_fa_3_7_y2;
  assign out[11] = f_u_arr_mul8_fa_4_7_y2;
  assign out[12] = f_u_arr_mul8_fa_5_7_y2;
  assign out[13] = f_u_arr_mul8_fa_6_7_y2;
  assign out[14] = f_u_arr_mul8_fa_7_7_y2;
  assign out[15] = f_u_arr_mul8_fa_7_7_y4;
endmodule