module s_cska8(input [7:0] a, input [7:0] b, output [8:0] s_cska8_out);
  wire s_cska8_xor0;
  wire s_cska8_ha0_xor0;
  wire s_cska8_ha0_and0;
  wire s_cska8_xor1;
  wire s_cska8_fa0_xor0;
  wire s_cska8_fa0_and0;
  wire s_cska8_fa0_xor1;
  wire s_cska8_fa0_and1;
  wire s_cska8_fa0_or0;
  wire s_cska8_xor2;
  wire s_cska8_fa1_xor0;
  wire s_cska8_fa1_and0;
  wire s_cska8_fa1_xor1;
  wire s_cska8_fa1_and1;
  wire s_cska8_fa1_or0;
  wire s_cska8_xor3;
  wire s_cska8_fa2_xor0;
  wire s_cska8_fa2_and0;
  wire s_cska8_fa2_xor1;
  wire s_cska8_fa2_and1;
  wire s_cska8_fa2_or0;
  wire s_cska8_and_propagate00;
  wire s_cska8_and_propagate01;
  wire s_cska8_and_propagate02;
  wire s_cska8_mux2to10_not0;
  wire s_cska8_mux2to10_and1;
  wire s_cska8_xor4;
  wire s_cska8_fa3_xor0;
  wire s_cska8_fa3_and0;
  wire s_cska8_fa3_xor1;
  wire s_cska8_fa3_and1;
  wire s_cska8_fa3_or0;
  wire s_cska8_xor5;
  wire s_cska8_fa4_xor0;
  wire s_cska8_fa4_and0;
  wire s_cska8_fa4_xor1;
  wire s_cska8_fa4_and1;
  wire s_cska8_fa4_or0;
  wire s_cska8_xor6;
  wire s_cska8_fa5_xor0;
  wire s_cska8_fa5_and0;
  wire s_cska8_fa5_xor1;
  wire s_cska8_fa5_and1;
  wire s_cska8_fa5_or0;
  wire s_cska8_xor7;
  wire s_cska8_fa6_xor0;
  wire s_cska8_fa6_and0;
  wire s_cska8_fa6_xor1;
  wire s_cska8_fa6_and1;
  wire s_cska8_fa6_or0;
  wire s_cska8_and_propagate13;
  wire s_cska8_and_propagate14;
  wire s_cska8_and_propagate15;
  wire s_cska8_mux2to11_and0;
  wire s_cska8_mux2to11_not0;
  wire s_cska8_mux2to11_and1;
  wire s_cska8_mux2to11_xor0;
  wire s_cska8_xor8;
  wire s_cska8_xor9;

  assign s_cska8_xor0 = a[0] ^ b[0];
  assign s_cska8_ha0_xor0 = a[0] ^ b[0];
  assign s_cska8_ha0_and0 = a[0] & b[0];
  assign s_cska8_xor1 = a[1] ^ b[1];
  assign s_cska8_fa0_xor0 = a[1] ^ b[1];
  assign s_cska8_fa0_and0 = a[1] & b[1];
  assign s_cska8_fa0_xor1 = s_cska8_fa0_xor0 ^ s_cska8_ha0_and0;
  assign s_cska8_fa0_and1 = s_cska8_fa0_xor0 & s_cska8_ha0_and0;
  assign s_cska8_fa0_or0 = s_cska8_fa0_and0 | s_cska8_fa0_and1;
  assign s_cska8_xor2 = a[2] ^ b[2];
  assign s_cska8_fa1_xor0 = a[2] ^ b[2];
  assign s_cska8_fa1_and0 = a[2] & b[2];
  assign s_cska8_fa1_xor1 = s_cska8_fa1_xor0 ^ s_cska8_fa0_or0;
  assign s_cska8_fa1_and1 = s_cska8_fa1_xor0 & s_cska8_fa0_or0;
  assign s_cska8_fa1_or0 = s_cska8_fa1_and0 | s_cska8_fa1_and1;
  assign s_cska8_xor3 = a[3] ^ b[3];
  assign s_cska8_fa2_xor0 = a[3] ^ b[3];
  assign s_cska8_fa2_and0 = a[3] & b[3];
  assign s_cska8_fa2_xor1 = s_cska8_fa2_xor0 ^ s_cska8_fa1_or0;
  assign s_cska8_fa2_and1 = s_cska8_fa2_xor0 & s_cska8_fa1_or0;
  assign s_cska8_fa2_or0 = s_cska8_fa2_and0 | s_cska8_fa2_and1;
  assign s_cska8_and_propagate00 = s_cska8_xor0 & s_cska8_xor2;
  assign s_cska8_and_propagate01 = s_cska8_xor1 & s_cska8_xor3;
  assign s_cska8_and_propagate02 = s_cska8_and_propagate00 & s_cska8_and_propagate01;
  assign s_cska8_mux2to10_not0 = ~s_cska8_and_propagate02;
  assign s_cska8_mux2to10_and1 = s_cska8_fa2_or0 & s_cska8_mux2to10_not0;
  assign s_cska8_xor4 = a[4] ^ b[4];
  assign s_cska8_fa3_xor0 = a[4] ^ b[4];
  assign s_cska8_fa3_and0 = a[4] & b[4];
  assign s_cska8_fa3_xor1 = s_cska8_fa3_xor0 ^ s_cska8_mux2to10_and1;
  assign s_cska8_fa3_and1 = s_cska8_fa3_xor0 & s_cska8_mux2to10_and1;
  assign s_cska8_fa3_or0 = s_cska8_fa3_and0 | s_cska8_fa3_and1;
  assign s_cska8_xor5 = a[5] ^ b[5];
  assign s_cska8_fa4_xor0 = a[5] ^ b[5];
  assign s_cska8_fa4_and0 = a[5] & b[5];
  assign s_cska8_fa4_xor1 = s_cska8_fa4_xor0 ^ s_cska8_fa3_or0;
  assign s_cska8_fa4_and1 = s_cska8_fa4_xor0 & s_cska8_fa3_or0;
  assign s_cska8_fa4_or0 = s_cska8_fa4_and0 | s_cska8_fa4_and1;
  assign s_cska8_xor6 = a[6] ^ b[6];
  assign s_cska8_fa5_xor0 = a[6] ^ b[6];
  assign s_cska8_fa5_and0 = a[6] & b[6];
  assign s_cska8_fa5_xor1 = s_cska8_fa5_xor0 ^ s_cska8_fa4_or0;
  assign s_cska8_fa5_and1 = s_cska8_fa5_xor0 & s_cska8_fa4_or0;
  assign s_cska8_fa5_or0 = s_cska8_fa5_and0 | s_cska8_fa5_and1;
  assign s_cska8_xor7 = a[7] ^ b[7];
  assign s_cska8_fa6_xor0 = a[7] ^ b[7];
  assign s_cska8_fa6_and0 = a[7] & b[7];
  assign s_cska8_fa6_xor1 = s_cska8_fa6_xor0 ^ s_cska8_fa5_or0;
  assign s_cska8_fa6_and1 = s_cska8_fa6_xor0 & s_cska8_fa5_or0;
  assign s_cska8_fa6_or0 = s_cska8_fa6_and0 | s_cska8_fa6_and1;
  assign s_cska8_and_propagate13 = s_cska8_xor4 & s_cska8_xor6;
  assign s_cska8_and_propagate14 = s_cska8_xor5 & s_cska8_xor7;
  assign s_cska8_and_propagate15 = s_cska8_and_propagate13 & s_cska8_and_propagate14;
  assign s_cska8_mux2to11_and0 = s_cska8_mux2to10_and1 & s_cska8_and_propagate15;
  assign s_cska8_mux2to11_not0 = ~s_cska8_and_propagate15;
  assign s_cska8_mux2to11_and1 = s_cska8_fa6_or0 & s_cska8_mux2to11_not0;
  assign s_cska8_mux2to11_xor0 = s_cska8_mux2to11_and0 ^ s_cska8_mux2to11_and1;
  assign s_cska8_xor8 = a[7] ^ b[7];
  assign s_cska8_xor9 = s_cska8_xor8 ^ s_cska8_mux2to11_xor0;

  assign s_cska8_out[0] = s_cska8_ha0_xor0;
  assign s_cska8_out[1] = s_cska8_fa0_xor1;
  assign s_cska8_out[2] = s_cska8_fa1_xor1;
  assign s_cska8_out[3] = s_cska8_fa2_xor1;
  assign s_cska8_out[4] = s_cska8_fa3_xor1;
  assign s_cska8_out[5] = s_cska8_fa4_xor1;
  assign s_cska8_out[6] = s_cska8_fa5_xor1;
  assign s_cska8_out[7] = s_cska8_fa6_xor1;
  assign s_cska8_out[8] = s_cska8_xor9;
endmodule