module f_arrdiv24(input [23:0] a, input [23:0] b, output [23:0] f_arrdiv24_out);
  wire f_arrdiv24_fs0_xor0;
  wire f_arrdiv24_fs0_not0;
  wire f_arrdiv24_fs0_and0;
  wire f_arrdiv24_fs0_not1;
  wire f_arrdiv24_fs1_xor1;
  wire f_arrdiv24_fs1_not1;
  wire f_arrdiv24_fs1_and1;
  wire f_arrdiv24_fs1_or0;
  wire f_arrdiv24_fs2_xor1;
  wire f_arrdiv24_fs2_not1;
  wire f_arrdiv24_fs2_and1;
  wire f_arrdiv24_fs2_or0;
  wire f_arrdiv24_fs3_xor1;
  wire f_arrdiv24_fs3_not1;
  wire f_arrdiv24_fs3_and1;
  wire f_arrdiv24_fs3_or0;
  wire f_arrdiv24_fs4_xor1;
  wire f_arrdiv24_fs4_not1;
  wire f_arrdiv24_fs4_and1;
  wire f_arrdiv24_fs4_or0;
  wire f_arrdiv24_fs5_xor1;
  wire f_arrdiv24_fs5_not1;
  wire f_arrdiv24_fs5_and1;
  wire f_arrdiv24_fs5_or0;
  wire f_arrdiv24_fs6_xor1;
  wire f_arrdiv24_fs6_not1;
  wire f_arrdiv24_fs6_and1;
  wire f_arrdiv24_fs6_or0;
  wire f_arrdiv24_fs7_xor1;
  wire f_arrdiv24_fs7_not1;
  wire f_arrdiv24_fs7_and1;
  wire f_arrdiv24_fs7_or0;
  wire f_arrdiv24_fs8_xor1;
  wire f_arrdiv24_fs8_not1;
  wire f_arrdiv24_fs8_and1;
  wire f_arrdiv24_fs8_or0;
  wire f_arrdiv24_fs9_xor1;
  wire f_arrdiv24_fs9_not1;
  wire f_arrdiv24_fs9_and1;
  wire f_arrdiv24_fs9_or0;
  wire f_arrdiv24_fs10_xor1;
  wire f_arrdiv24_fs10_not1;
  wire f_arrdiv24_fs10_and1;
  wire f_arrdiv24_fs10_or0;
  wire f_arrdiv24_fs11_xor1;
  wire f_arrdiv24_fs11_not1;
  wire f_arrdiv24_fs11_and1;
  wire f_arrdiv24_fs11_or0;
  wire f_arrdiv24_fs12_xor1;
  wire f_arrdiv24_fs12_not1;
  wire f_arrdiv24_fs12_and1;
  wire f_arrdiv24_fs12_or0;
  wire f_arrdiv24_fs13_xor1;
  wire f_arrdiv24_fs13_not1;
  wire f_arrdiv24_fs13_and1;
  wire f_arrdiv24_fs13_or0;
  wire f_arrdiv24_fs14_xor1;
  wire f_arrdiv24_fs14_not1;
  wire f_arrdiv24_fs14_and1;
  wire f_arrdiv24_fs14_or0;
  wire f_arrdiv24_fs15_xor1;
  wire f_arrdiv24_fs15_not1;
  wire f_arrdiv24_fs15_and1;
  wire f_arrdiv24_fs15_or0;
  wire f_arrdiv24_fs16_xor1;
  wire f_arrdiv24_fs16_not1;
  wire f_arrdiv24_fs16_and1;
  wire f_arrdiv24_fs16_or0;
  wire f_arrdiv24_fs17_xor1;
  wire f_arrdiv24_fs17_not1;
  wire f_arrdiv24_fs17_and1;
  wire f_arrdiv24_fs17_or0;
  wire f_arrdiv24_fs18_xor1;
  wire f_arrdiv24_fs18_not1;
  wire f_arrdiv24_fs18_and1;
  wire f_arrdiv24_fs18_or0;
  wire f_arrdiv24_fs19_xor1;
  wire f_arrdiv24_fs19_not1;
  wire f_arrdiv24_fs19_and1;
  wire f_arrdiv24_fs19_or0;
  wire f_arrdiv24_fs20_xor1;
  wire f_arrdiv24_fs20_not1;
  wire f_arrdiv24_fs20_and1;
  wire f_arrdiv24_fs20_or0;
  wire f_arrdiv24_fs21_xor1;
  wire f_arrdiv24_fs21_not1;
  wire f_arrdiv24_fs21_and1;
  wire f_arrdiv24_fs21_or0;
  wire f_arrdiv24_fs22_xor1;
  wire f_arrdiv24_fs22_not1;
  wire f_arrdiv24_fs22_and1;
  wire f_arrdiv24_fs22_or0;
  wire f_arrdiv24_fs23_xor1;
  wire f_arrdiv24_fs23_not1;
  wire f_arrdiv24_fs23_and1;
  wire f_arrdiv24_fs23_or0;
  wire f_arrdiv24_mux2to10_and0;
  wire f_arrdiv24_mux2to10_not0;
  wire f_arrdiv24_mux2to10_and1;
  wire f_arrdiv24_mux2to10_xor0;
  wire f_arrdiv24_mux2to11_not0;
  wire f_arrdiv24_mux2to11_and1;
  wire f_arrdiv24_mux2to12_not0;
  wire f_arrdiv24_mux2to12_and1;
  wire f_arrdiv24_mux2to13_not0;
  wire f_arrdiv24_mux2to13_and1;
  wire f_arrdiv24_mux2to14_not0;
  wire f_arrdiv24_mux2to14_and1;
  wire f_arrdiv24_mux2to15_not0;
  wire f_arrdiv24_mux2to15_and1;
  wire f_arrdiv24_mux2to16_not0;
  wire f_arrdiv24_mux2to16_and1;
  wire f_arrdiv24_mux2to17_not0;
  wire f_arrdiv24_mux2to17_and1;
  wire f_arrdiv24_mux2to18_not0;
  wire f_arrdiv24_mux2to18_and1;
  wire f_arrdiv24_mux2to19_not0;
  wire f_arrdiv24_mux2to19_and1;
  wire f_arrdiv24_mux2to110_not0;
  wire f_arrdiv24_mux2to110_and1;
  wire f_arrdiv24_mux2to111_not0;
  wire f_arrdiv24_mux2to111_and1;
  wire f_arrdiv24_mux2to112_not0;
  wire f_arrdiv24_mux2to112_and1;
  wire f_arrdiv24_mux2to113_not0;
  wire f_arrdiv24_mux2to113_and1;
  wire f_arrdiv24_mux2to114_not0;
  wire f_arrdiv24_mux2to114_and1;
  wire f_arrdiv24_mux2to115_not0;
  wire f_arrdiv24_mux2to115_and1;
  wire f_arrdiv24_mux2to116_not0;
  wire f_arrdiv24_mux2to116_and1;
  wire f_arrdiv24_mux2to117_not0;
  wire f_arrdiv24_mux2to117_and1;
  wire f_arrdiv24_mux2to118_not0;
  wire f_arrdiv24_mux2to118_and1;
  wire f_arrdiv24_mux2to119_not0;
  wire f_arrdiv24_mux2to119_and1;
  wire f_arrdiv24_mux2to120_not0;
  wire f_arrdiv24_mux2to120_and1;
  wire f_arrdiv24_mux2to121_not0;
  wire f_arrdiv24_mux2to121_and1;
  wire f_arrdiv24_mux2to122_not0;
  wire f_arrdiv24_mux2to122_and1;
  wire f_arrdiv24_not0;
  wire f_arrdiv24_fs24_xor0;
  wire f_arrdiv24_fs24_not0;
  wire f_arrdiv24_fs24_and0;
  wire f_arrdiv24_fs24_not1;
  wire f_arrdiv24_fs25_xor0;
  wire f_arrdiv24_fs25_not0;
  wire f_arrdiv24_fs25_and0;
  wire f_arrdiv24_fs25_xor1;
  wire f_arrdiv24_fs25_not1;
  wire f_arrdiv24_fs25_and1;
  wire f_arrdiv24_fs25_or0;
  wire f_arrdiv24_fs26_xor0;
  wire f_arrdiv24_fs26_not0;
  wire f_arrdiv24_fs26_and0;
  wire f_arrdiv24_fs26_xor1;
  wire f_arrdiv24_fs26_not1;
  wire f_arrdiv24_fs26_and1;
  wire f_arrdiv24_fs26_or0;
  wire f_arrdiv24_fs27_xor0;
  wire f_arrdiv24_fs27_not0;
  wire f_arrdiv24_fs27_and0;
  wire f_arrdiv24_fs27_xor1;
  wire f_arrdiv24_fs27_not1;
  wire f_arrdiv24_fs27_and1;
  wire f_arrdiv24_fs27_or0;
  wire f_arrdiv24_fs28_xor0;
  wire f_arrdiv24_fs28_not0;
  wire f_arrdiv24_fs28_and0;
  wire f_arrdiv24_fs28_xor1;
  wire f_arrdiv24_fs28_not1;
  wire f_arrdiv24_fs28_and1;
  wire f_arrdiv24_fs28_or0;
  wire f_arrdiv24_fs29_xor0;
  wire f_arrdiv24_fs29_not0;
  wire f_arrdiv24_fs29_and0;
  wire f_arrdiv24_fs29_xor1;
  wire f_arrdiv24_fs29_not1;
  wire f_arrdiv24_fs29_and1;
  wire f_arrdiv24_fs29_or0;
  wire f_arrdiv24_fs30_xor0;
  wire f_arrdiv24_fs30_not0;
  wire f_arrdiv24_fs30_and0;
  wire f_arrdiv24_fs30_xor1;
  wire f_arrdiv24_fs30_not1;
  wire f_arrdiv24_fs30_and1;
  wire f_arrdiv24_fs30_or0;
  wire f_arrdiv24_fs31_xor0;
  wire f_arrdiv24_fs31_not0;
  wire f_arrdiv24_fs31_and0;
  wire f_arrdiv24_fs31_xor1;
  wire f_arrdiv24_fs31_not1;
  wire f_arrdiv24_fs31_and1;
  wire f_arrdiv24_fs31_or0;
  wire f_arrdiv24_fs32_xor0;
  wire f_arrdiv24_fs32_not0;
  wire f_arrdiv24_fs32_and0;
  wire f_arrdiv24_fs32_xor1;
  wire f_arrdiv24_fs32_not1;
  wire f_arrdiv24_fs32_and1;
  wire f_arrdiv24_fs32_or0;
  wire f_arrdiv24_fs33_xor0;
  wire f_arrdiv24_fs33_not0;
  wire f_arrdiv24_fs33_and0;
  wire f_arrdiv24_fs33_xor1;
  wire f_arrdiv24_fs33_not1;
  wire f_arrdiv24_fs33_and1;
  wire f_arrdiv24_fs33_or0;
  wire f_arrdiv24_fs34_xor0;
  wire f_arrdiv24_fs34_not0;
  wire f_arrdiv24_fs34_and0;
  wire f_arrdiv24_fs34_xor1;
  wire f_arrdiv24_fs34_not1;
  wire f_arrdiv24_fs34_and1;
  wire f_arrdiv24_fs34_or0;
  wire f_arrdiv24_fs35_xor0;
  wire f_arrdiv24_fs35_not0;
  wire f_arrdiv24_fs35_and0;
  wire f_arrdiv24_fs35_xor1;
  wire f_arrdiv24_fs35_not1;
  wire f_arrdiv24_fs35_and1;
  wire f_arrdiv24_fs35_or0;
  wire f_arrdiv24_fs36_xor0;
  wire f_arrdiv24_fs36_not0;
  wire f_arrdiv24_fs36_and0;
  wire f_arrdiv24_fs36_xor1;
  wire f_arrdiv24_fs36_not1;
  wire f_arrdiv24_fs36_and1;
  wire f_arrdiv24_fs36_or0;
  wire f_arrdiv24_fs37_xor0;
  wire f_arrdiv24_fs37_not0;
  wire f_arrdiv24_fs37_and0;
  wire f_arrdiv24_fs37_xor1;
  wire f_arrdiv24_fs37_not1;
  wire f_arrdiv24_fs37_and1;
  wire f_arrdiv24_fs37_or0;
  wire f_arrdiv24_fs38_xor0;
  wire f_arrdiv24_fs38_not0;
  wire f_arrdiv24_fs38_and0;
  wire f_arrdiv24_fs38_xor1;
  wire f_arrdiv24_fs38_not1;
  wire f_arrdiv24_fs38_and1;
  wire f_arrdiv24_fs38_or0;
  wire f_arrdiv24_fs39_xor0;
  wire f_arrdiv24_fs39_not0;
  wire f_arrdiv24_fs39_and0;
  wire f_arrdiv24_fs39_xor1;
  wire f_arrdiv24_fs39_not1;
  wire f_arrdiv24_fs39_and1;
  wire f_arrdiv24_fs39_or0;
  wire f_arrdiv24_fs40_xor0;
  wire f_arrdiv24_fs40_not0;
  wire f_arrdiv24_fs40_and0;
  wire f_arrdiv24_fs40_xor1;
  wire f_arrdiv24_fs40_not1;
  wire f_arrdiv24_fs40_and1;
  wire f_arrdiv24_fs40_or0;
  wire f_arrdiv24_fs41_xor0;
  wire f_arrdiv24_fs41_not0;
  wire f_arrdiv24_fs41_and0;
  wire f_arrdiv24_fs41_xor1;
  wire f_arrdiv24_fs41_not1;
  wire f_arrdiv24_fs41_and1;
  wire f_arrdiv24_fs41_or0;
  wire f_arrdiv24_fs42_xor0;
  wire f_arrdiv24_fs42_not0;
  wire f_arrdiv24_fs42_and0;
  wire f_arrdiv24_fs42_xor1;
  wire f_arrdiv24_fs42_not1;
  wire f_arrdiv24_fs42_and1;
  wire f_arrdiv24_fs42_or0;
  wire f_arrdiv24_fs43_xor0;
  wire f_arrdiv24_fs43_not0;
  wire f_arrdiv24_fs43_and0;
  wire f_arrdiv24_fs43_xor1;
  wire f_arrdiv24_fs43_not1;
  wire f_arrdiv24_fs43_and1;
  wire f_arrdiv24_fs43_or0;
  wire f_arrdiv24_fs44_xor0;
  wire f_arrdiv24_fs44_not0;
  wire f_arrdiv24_fs44_and0;
  wire f_arrdiv24_fs44_xor1;
  wire f_arrdiv24_fs44_not1;
  wire f_arrdiv24_fs44_and1;
  wire f_arrdiv24_fs44_or0;
  wire f_arrdiv24_fs45_xor0;
  wire f_arrdiv24_fs45_not0;
  wire f_arrdiv24_fs45_and0;
  wire f_arrdiv24_fs45_xor1;
  wire f_arrdiv24_fs45_not1;
  wire f_arrdiv24_fs45_and1;
  wire f_arrdiv24_fs45_or0;
  wire f_arrdiv24_fs46_xor0;
  wire f_arrdiv24_fs46_not0;
  wire f_arrdiv24_fs46_and0;
  wire f_arrdiv24_fs46_xor1;
  wire f_arrdiv24_fs46_not1;
  wire f_arrdiv24_fs46_and1;
  wire f_arrdiv24_fs46_or0;
  wire f_arrdiv24_fs47_xor0;
  wire f_arrdiv24_fs47_not0;
  wire f_arrdiv24_fs47_and0;
  wire f_arrdiv24_fs47_xor1;
  wire f_arrdiv24_fs47_not1;
  wire f_arrdiv24_fs47_and1;
  wire f_arrdiv24_fs47_or0;
  wire f_arrdiv24_mux2to123_and0;
  wire f_arrdiv24_mux2to123_not0;
  wire f_arrdiv24_mux2to123_and1;
  wire f_arrdiv24_mux2to123_xor0;
  wire f_arrdiv24_mux2to124_and0;
  wire f_arrdiv24_mux2to124_not0;
  wire f_arrdiv24_mux2to124_and1;
  wire f_arrdiv24_mux2to124_xor0;
  wire f_arrdiv24_mux2to125_and0;
  wire f_arrdiv24_mux2to125_not0;
  wire f_arrdiv24_mux2to125_and1;
  wire f_arrdiv24_mux2to125_xor0;
  wire f_arrdiv24_mux2to126_and0;
  wire f_arrdiv24_mux2to126_not0;
  wire f_arrdiv24_mux2to126_and1;
  wire f_arrdiv24_mux2to126_xor0;
  wire f_arrdiv24_mux2to127_and0;
  wire f_arrdiv24_mux2to127_not0;
  wire f_arrdiv24_mux2to127_and1;
  wire f_arrdiv24_mux2to127_xor0;
  wire f_arrdiv24_mux2to128_and0;
  wire f_arrdiv24_mux2to128_not0;
  wire f_arrdiv24_mux2to128_and1;
  wire f_arrdiv24_mux2to128_xor0;
  wire f_arrdiv24_mux2to129_and0;
  wire f_arrdiv24_mux2to129_not0;
  wire f_arrdiv24_mux2to129_and1;
  wire f_arrdiv24_mux2to129_xor0;
  wire f_arrdiv24_mux2to130_and0;
  wire f_arrdiv24_mux2to130_not0;
  wire f_arrdiv24_mux2to130_and1;
  wire f_arrdiv24_mux2to130_xor0;
  wire f_arrdiv24_mux2to131_and0;
  wire f_arrdiv24_mux2to131_not0;
  wire f_arrdiv24_mux2to131_and1;
  wire f_arrdiv24_mux2to131_xor0;
  wire f_arrdiv24_mux2to132_and0;
  wire f_arrdiv24_mux2to132_not0;
  wire f_arrdiv24_mux2to132_and1;
  wire f_arrdiv24_mux2to132_xor0;
  wire f_arrdiv24_mux2to133_and0;
  wire f_arrdiv24_mux2to133_not0;
  wire f_arrdiv24_mux2to133_and1;
  wire f_arrdiv24_mux2to133_xor0;
  wire f_arrdiv24_mux2to134_and0;
  wire f_arrdiv24_mux2to134_not0;
  wire f_arrdiv24_mux2to134_and1;
  wire f_arrdiv24_mux2to134_xor0;
  wire f_arrdiv24_mux2to135_and0;
  wire f_arrdiv24_mux2to135_not0;
  wire f_arrdiv24_mux2to135_and1;
  wire f_arrdiv24_mux2to135_xor0;
  wire f_arrdiv24_mux2to136_and0;
  wire f_arrdiv24_mux2to136_not0;
  wire f_arrdiv24_mux2to136_and1;
  wire f_arrdiv24_mux2to136_xor0;
  wire f_arrdiv24_mux2to137_and0;
  wire f_arrdiv24_mux2to137_not0;
  wire f_arrdiv24_mux2to137_and1;
  wire f_arrdiv24_mux2to137_xor0;
  wire f_arrdiv24_mux2to138_and0;
  wire f_arrdiv24_mux2to138_not0;
  wire f_arrdiv24_mux2to138_and1;
  wire f_arrdiv24_mux2to138_xor0;
  wire f_arrdiv24_mux2to139_and0;
  wire f_arrdiv24_mux2to139_not0;
  wire f_arrdiv24_mux2to139_and1;
  wire f_arrdiv24_mux2to139_xor0;
  wire f_arrdiv24_mux2to140_and0;
  wire f_arrdiv24_mux2to140_not0;
  wire f_arrdiv24_mux2to140_and1;
  wire f_arrdiv24_mux2to140_xor0;
  wire f_arrdiv24_mux2to141_and0;
  wire f_arrdiv24_mux2to141_not0;
  wire f_arrdiv24_mux2to141_and1;
  wire f_arrdiv24_mux2to141_xor0;
  wire f_arrdiv24_mux2to142_and0;
  wire f_arrdiv24_mux2to142_not0;
  wire f_arrdiv24_mux2to142_and1;
  wire f_arrdiv24_mux2to142_xor0;
  wire f_arrdiv24_mux2to143_and0;
  wire f_arrdiv24_mux2to143_not0;
  wire f_arrdiv24_mux2to143_and1;
  wire f_arrdiv24_mux2to143_xor0;
  wire f_arrdiv24_mux2to144_and0;
  wire f_arrdiv24_mux2to144_not0;
  wire f_arrdiv24_mux2to144_and1;
  wire f_arrdiv24_mux2to144_xor0;
  wire f_arrdiv24_mux2to145_and0;
  wire f_arrdiv24_mux2to145_not0;
  wire f_arrdiv24_mux2to145_and1;
  wire f_arrdiv24_mux2to145_xor0;
  wire f_arrdiv24_not1;
  wire f_arrdiv24_fs48_xor0;
  wire f_arrdiv24_fs48_not0;
  wire f_arrdiv24_fs48_and0;
  wire f_arrdiv24_fs48_not1;
  wire f_arrdiv24_fs49_xor0;
  wire f_arrdiv24_fs49_not0;
  wire f_arrdiv24_fs49_and0;
  wire f_arrdiv24_fs49_xor1;
  wire f_arrdiv24_fs49_not1;
  wire f_arrdiv24_fs49_and1;
  wire f_arrdiv24_fs49_or0;
  wire f_arrdiv24_fs50_xor0;
  wire f_arrdiv24_fs50_not0;
  wire f_arrdiv24_fs50_and0;
  wire f_arrdiv24_fs50_xor1;
  wire f_arrdiv24_fs50_not1;
  wire f_arrdiv24_fs50_and1;
  wire f_arrdiv24_fs50_or0;
  wire f_arrdiv24_fs51_xor0;
  wire f_arrdiv24_fs51_not0;
  wire f_arrdiv24_fs51_and0;
  wire f_arrdiv24_fs51_xor1;
  wire f_arrdiv24_fs51_not1;
  wire f_arrdiv24_fs51_and1;
  wire f_arrdiv24_fs51_or0;
  wire f_arrdiv24_fs52_xor0;
  wire f_arrdiv24_fs52_not0;
  wire f_arrdiv24_fs52_and0;
  wire f_arrdiv24_fs52_xor1;
  wire f_arrdiv24_fs52_not1;
  wire f_arrdiv24_fs52_and1;
  wire f_arrdiv24_fs52_or0;
  wire f_arrdiv24_fs53_xor0;
  wire f_arrdiv24_fs53_not0;
  wire f_arrdiv24_fs53_and0;
  wire f_arrdiv24_fs53_xor1;
  wire f_arrdiv24_fs53_not1;
  wire f_arrdiv24_fs53_and1;
  wire f_arrdiv24_fs53_or0;
  wire f_arrdiv24_fs54_xor0;
  wire f_arrdiv24_fs54_not0;
  wire f_arrdiv24_fs54_and0;
  wire f_arrdiv24_fs54_xor1;
  wire f_arrdiv24_fs54_not1;
  wire f_arrdiv24_fs54_and1;
  wire f_arrdiv24_fs54_or0;
  wire f_arrdiv24_fs55_xor0;
  wire f_arrdiv24_fs55_not0;
  wire f_arrdiv24_fs55_and0;
  wire f_arrdiv24_fs55_xor1;
  wire f_arrdiv24_fs55_not1;
  wire f_arrdiv24_fs55_and1;
  wire f_arrdiv24_fs55_or0;
  wire f_arrdiv24_fs56_xor0;
  wire f_arrdiv24_fs56_not0;
  wire f_arrdiv24_fs56_and0;
  wire f_arrdiv24_fs56_xor1;
  wire f_arrdiv24_fs56_not1;
  wire f_arrdiv24_fs56_and1;
  wire f_arrdiv24_fs56_or0;
  wire f_arrdiv24_fs57_xor0;
  wire f_arrdiv24_fs57_not0;
  wire f_arrdiv24_fs57_and0;
  wire f_arrdiv24_fs57_xor1;
  wire f_arrdiv24_fs57_not1;
  wire f_arrdiv24_fs57_and1;
  wire f_arrdiv24_fs57_or0;
  wire f_arrdiv24_fs58_xor0;
  wire f_arrdiv24_fs58_not0;
  wire f_arrdiv24_fs58_and0;
  wire f_arrdiv24_fs58_xor1;
  wire f_arrdiv24_fs58_not1;
  wire f_arrdiv24_fs58_and1;
  wire f_arrdiv24_fs58_or0;
  wire f_arrdiv24_fs59_xor0;
  wire f_arrdiv24_fs59_not0;
  wire f_arrdiv24_fs59_and0;
  wire f_arrdiv24_fs59_xor1;
  wire f_arrdiv24_fs59_not1;
  wire f_arrdiv24_fs59_and1;
  wire f_arrdiv24_fs59_or0;
  wire f_arrdiv24_fs60_xor0;
  wire f_arrdiv24_fs60_not0;
  wire f_arrdiv24_fs60_and0;
  wire f_arrdiv24_fs60_xor1;
  wire f_arrdiv24_fs60_not1;
  wire f_arrdiv24_fs60_and1;
  wire f_arrdiv24_fs60_or0;
  wire f_arrdiv24_fs61_xor0;
  wire f_arrdiv24_fs61_not0;
  wire f_arrdiv24_fs61_and0;
  wire f_arrdiv24_fs61_xor1;
  wire f_arrdiv24_fs61_not1;
  wire f_arrdiv24_fs61_and1;
  wire f_arrdiv24_fs61_or0;
  wire f_arrdiv24_fs62_xor0;
  wire f_arrdiv24_fs62_not0;
  wire f_arrdiv24_fs62_and0;
  wire f_arrdiv24_fs62_xor1;
  wire f_arrdiv24_fs62_not1;
  wire f_arrdiv24_fs62_and1;
  wire f_arrdiv24_fs62_or0;
  wire f_arrdiv24_fs63_xor0;
  wire f_arrdiv24_fs63_not0;
  wire f_arrdiv24_fs63_and0;
  wire f_arrdiv24_fs63_xor1;
  wire f_arrdiv24_fs63_not1;
  wire f_arrdiv24_fs63_and1;
  wire f_arrdiv24_fs63_or0;
  wire f_arrdiv24_fs64_xor0;
  wire f_arrdiv24_fs64_not0;
  wire f_arrdiv24_fs64_and0;
  wire f_arrdiv24_fs64_xor1;
  wire f_arrdiv24_fs64_not1;
  wire f_arrdiv24_fs64_and1;
  wire f_arrdiv24_fs64_or0;
  wire f_arrdiv24_fs65_xor0;
  wire f_arrdiv24_fs65_not0;
  wire f_arrdiv24_fs65_and0;
  wire f_arrdiv24_fs65_xor1;
  wire f_arrdiv24_fs65_not1;
  wire f_arrdiv24_fs65_and1;
  wire f_arrdiv24_fs65_or0;
  wire f_arrdiv24_fs66_xor0;
  wire f_arrdiv24_fs66_not0;
  wire f_arrdiv24_fs66_and0;
  wire f_arrdiv24_fs66_xor1;
  wire f_arrdiv24_fs66_not1;
  wire f_arrdiv24_fs66_and1;
  wire f_arrdiv24_fs66_or0;
  wire f_arrdiv24_fs67_xor0;
  wire f_arrdiv24_fs67_not0;
  wire f_arrdiv24_fs67_and0;
  wire f_arrdiv24_fs67_xor1;
  wire f_arrdiv24_fs67_not1;
  wire f_arrdiv24_fs67_and1;
  wire f_arrdiv24_fs67_or0;
  wire f_arrdiv24_fs68_xor0;
  wire f_arrdiv24_fs68_not0;
  wire f_arrdiv24_fs68_and0;
  wire f_arrdiv24_fs68_xor1;
  wire f_arrdiv24_fs68_not1;
  wire f_arrdiv24_fs68_and1;
  wire f_arrdiv24_fs68_or0;
  wire f_arrdiv24_fs69_xor0;
  wire f_arrdiv24_fs69_not0;
  wire f_arrdiv24_fs69_and0;
  wire f_arrdiv24_fs69_xor1;
  wire f_arrdiv24_fs69_not1;
  wire f_arrdiv24_fs69_and1;
  wire f_arrdiv24_fs69_or0;
  wire f_arrdiv24_fs70_xor0;
  wire f_arrdiv24_fs70_not0;
  wire f_arrdiv24_fs70_and0;
  wire f_arrdiv24_fs70_xor1;
  wire f_arrdiv24_fs70_not1;
  wire f_arrdiv24_fs70_and1;
  wire f_arrdiv24_fs70_or0;
  wire f_arrdiv24_fs71_xor0;
  wire f_arrdiv24_fs71_not0;
  wire f_arrdiv24_fs71_and0;
  wire f_arrdiv24_fs71_xor1;
  wire f_arrdiv24_fs71_not1;
  wire f_arrdiv24_fs71_and1;
  wire f_arrdiv24_fs71_or0;
  wire f_arrdiv24_mux2to146_and0;
  wire f_arrdiv24_mux2to146_not0;
  wire f_arrdiv24_mux2to146_and1;
  wire f_arrdiv24_mux2to146_xor0;
  wire f_arrdiv24_mux2to147_and0;
  wire f_arrdiv24_mux2to147_not0;
  wire f_arrdiv24_mux2to147_and1;
  wire f_arrdiv24_mux2to147_xor0;
  wire f_arrdiv24_mux2to148_and0;
  wire f_arrdiv24_mux2to148_not0;
  wire f_arrdiv24_mux2to148_and1;
  wire f_arrdiv24_mux2to148_xor0;
  wire f_arrdiv24_mux2to149_and0;
  wire f_arrdiv24_mux2to149_not0;
  wire f_arrdiv24_mux2to149_and1;
  wire f_arrdiv24_mux2to149_xor0;
  wire f_arrdiv24_mux2to150_and0;
  wire f_arrdiv24_mux2to150_not0;
  wire f_arrdiv24_mux2to150_and1;
  wire f_arrdiv24_mux2to150_xor0;
  wire f_arrdiv24_mux2to151_and0;
  wire f_arrdiv24_mux2to151_not0;
  wire f_arrdiv24_mux2to151_and1;
  wire f_arrdiv24_mux2to151_xor0;
  wire f_arrdiv24_mux2to152_and0;
  wire f_arrdiv24_mux2to152_not0;
  wire f_arrdiv24_mux2to152_and1;
  wire f_arrdiv24_mux2to152_xor0;
  wire f_arrdiv24_mux2to153_and0;
  wire f_arrdiv24_mux2to153_not0;
  wire f_arrdiv24_mux2to153_and1;
  wire f_arrdiv24_mux2to153_xor0;
  wire f_arrdiv24_mux2to154_and0;
  wire f_arrdiv24_mux2to154_not0;
  wire f_arrdiv24_mux2to154_and1;
  wire f_arrdiv24_mux2to154_xor0;
  wire f_arrdiv24_mux2to155_and0;
  wire f_arrdiv24_mux2to155_not0;
  wire f_arrdiv24_mux2to155_and1;
  wire f_arrdiv24_mux2to155_xor0;
  wire f_arrdiv24_mux2to156_and0;
  wire f_arrdiv24_mux2to156_not0;
  wire f_arrdiv24_mux2to156_and1;
  wire f_arrdiv24_mux2to156_xor0;
  wire f_arrdiv24_mux2to157_and0;
  wire f_arrdiv24_mux2to157_not0;
  wire f_arrdiv24_mux2to157_and1;
  wire f_arrdiv24_mux2to157_xor0;
  wire f_arrdiv24_mux2to158_and0;
  wire f_arrdiv24_mux2to158_not0;
  wire f_arrdiv24_mux2to158_and1;
  wire f_arrdiv24_mux2to158_xor0;
  wire f_arrdiv24_mux2to159_and0;
  wire f_arrdiv24_mux2to159_not0;
  wire f_arrdiv24_mux2to159_and1;
  wire f_arrdiv24_mux2to159_xor0;
  wire f_arrdiv24_mux2to160_and0;
  wire f_arrdiv24_mux2to160_not0;
  wire f_arrdiv24_mux2to160_and1;
  wire f_arrdiv24_mux2to160_xor0;
  wire f_arrdiv24_mux2to161_and0;
  wire f_arrdiv24_mux2to161_not0;
  wire f_arrdiv24_mux2to161_and1;
  wire f_arrdiv24_mux2to161_xor0;
  wire f_arrdiv24_mux2to162_and0;
  wire f_arrdiv24_mux2to162_not0;
  wire f_arrdiv24_mux2to162_and1;
  wire f_arrdiv24_mux2to162_xor0;
  wire f_arrdiv24_mux2to163_and0;
  wire f_arrdiv24_mux2to163_not0;
  wire f_arrdiv24_mux2to163_and1;
  wire f_arrdiv24_mux2to163_xor0;
  wire f_arrdiv24_mux2to164_and0;
  wire f_arrdiv24_mux2to164_not0;
  wire f_arrdiv24_mux2to164_and1;
  wire f_arrdiv24_mux2to164_xor0;
  wire f_arrdiv24_mux2to165_and0;
  wire f_arrdiv24_mux2to165_not0;
  wire f_arrdiv24_mux2to165_and1;
  wire f_arrdiv24_mux2to165_xor0;
  wire f_arrdiv24_mux2to166_and0;
  wire f_arrdiv24_mux2to166_not0;
  wire f_arrdiv24_mux2to166_and1;
  wire f_arrdiv24_mux2to166_xor0;
  wire f_arrdiv24_mux2to167_and0;
  wire f_arrdiv24_mux2to167_not0;
  wire f_arrdiv24_mux2to167_and1;
  wire f_arrdiv24_mux2to167_xor0;
  wire f_arrdiv24_mux2to168_and0;
  wire f_arrdiv24_mux2to168_not0;
  wire f_arrdiv24_mux2to168_and1;
  wire f_arrdiv24_mux2to168_xor0;
  wire f_arrdiv24_not2;
  wire f_arrdiv24_fs72_xor0;
  wire f_arrdiv24_fs72_not0;
  wire f_arrdiv24_fs72_and0;
  wire f_arrdiv24_fs72_not1;
  wire f_arrdiv24_fs73_xor0;
  wire f_arrdiv24_fs73_not0;
  wire f_arrdiv24_fs73_and0;
  wire f_arrdiv24_fs73_xor1;
  wire f_arrdiv24_fs73_not1;
  wire f_arrdiv24_fs73_and1;
  wire f_arrdiv24_fs73_or0;
  wire f_arrdiv24_fs74_xor0;
  wire f_arrdiv24_fs74_not0;
  wire f_arrdiv24_fs74_and0;
  wire f_arrdiv24_fs74_xor1;
  wire f_arrdiv24_fs74_not1;
  wire f_arrdiv24_fs74_and1;
  wire f_arrdiv24_fs74_or0;
  wire f_arrdiv24_fs75_xor0;
  wire f_arrdiv24_fs75_not0;
  wire f_arrdiv24_fs75_and0;
  wire f_arrdiv24_fs75_xor1;
  wire f_arrdiv24_fs75_not1;
  wire f_arrdiv24_fs75_and1;
  wire f_arrdiv24_fs75_or0;
  wire f_arrdiv24_fs76_xor0;
  wire f_arrdiv24_fs76_not0;
  wire f_arrdiv24_fs76_and0;
  wire f_arrdiv24_fs76_xor1;
  wire f_arrdiv24_fs76_not1;
  wire f_arrdiv24_fs76_and1;
  wire f_arrdiv24_fs76_or0;
  wire f_arrdiv24_fs77_xor0;
  wire f_arrdiv24_fs77_not0;
  wire f_arrdiv24_fs77_and0;
  wire f_arrdiv24_fs77_xor1;
  wire f_arrdiv24_fs77_not1;
  wire f_arrdiv24_fs77_and1;
  wire f_arrdiv24_fs77_or0;
  wire f_arrdiv24_fs78_xor0;
  wire f_arrdiv24_fs78_not0;
  wire f_arrdiv24_fs78_and0;
  wire f_arrdiv24_fs78_xor1;
  wire f_arrdiv24_fs78_not1;
  wire f_arrdiv24_fs78_and1;
  wire f_arrdiv24_fs78_or0;
  wire f_arrdiv24_fs79_xor0;
  wire f_arrdiv24_fs79_not0;
  wire f_arrdiv24_fs79_and0;
  wire f_arrdiv24_fs79_xor1;
  wire f_arrdiv24_fs79_not1;
  wire f_arrdiv24_fs79_and1;
  wire f_arrdiv24_fs79_or0;
  wire f_arrdiv24_fs80_xor0;
  wire f_arrdiv24_fs80_not0;
  wire f_arrdiv24_fs80_and0;
  wire f_arrdiv24_fs80_xor1;
  wire f_arrdiv24_fs80_not1;
  wire f_arrdiv24_fs80_and1;
  wire f_arrdiv24_fs80_or0;
  wire f_arrdiv24_fs81_xor0;
  wire f_arrdiv24_fs81_not0;
  wire f_arrdiv24_fs81_and0;
  wire f_arrdiv24_fs81_xor1;
  wire f_arrdiv24_fs81_not1;
  wire f_arrdiv24_fs81_and1;
  wire f_arrdiv24_fs81_or0;
  wire f_arrdiv24_fs82_xor0;
  wire f_arrdiv24_fs82_not0;
  wire f_arrdiv24_fs82_and0;
  wire f_arrdiv24_fs82_xor1;
  wire f_arrdiv24_fs82_not1;
  wire f_arrdiv24_fs82_and1;
  wire f_arrdiv24_fs82_or0;
  wire f_arrdiv24_fs83_xor0;
  wire f_arrdiv24_fs83_not0;
  wire f_arrdiv24_fs83_and0;
  wire f_arrdiv24_fs83_xor1;
  wire f_arrdiv24_fs83_not1;
  wire f_arrdiv24_fs83_and1;
  wire f_arrdiv24_fs83_or0;
  wire f_arrdiv24_fs84_xor0;
  wire f_arrdiv24_fs84_not0;
  wire f_arrdiv24_fs84_and0;
  wire f_arrdiv24_fs84_xor1;
  wire f_arrdiv24_fs84_not1;
  wire f_arrdiv24_fs84_and1;
  wire f_arrdiv24_fs84_or0;
  wire f_arrdiv24_fs85_xor0;
  wire f_arrdiv24_fs85_not0;
  wire f_arrdiv24_fs85_and0;
  wire f_arrdiv24_fs85_xor1;
  wire f_arrdiv24_fs85_not1;
  wire f_arrdiv24_fs85_and1;
  wire f_arrdiv24_fs85_or0;
  wire f_arrdiv24_fs86_xor0;
  wire f_arrdiv24_fs86_not0;
  wire f_arrdiv24_fs86_and0;
  wire f_arrdiv24_fs86_xor1;
  wire f_arrdiv24_fs86_not1;
  wire f_arrdiv24_fs86_and1;
  wire f_arrdiv24_fs86_or0;
  wire f_arrdiv24_fs87_xor0;
  wire f_arrdiv24_fs87_not0;
  wire f_arrdiv24_fs87_and0;
  wire f_arrdiv24_fs87_xor1;
  wire f_arrdiv24_fs87_not1;
  wire f_arrdiv24_fs87_and1;
  wire f_arrdiv24_fs87_or0;
  wire f_arrdiv24_fs88_xor0;
  wire f_arrdiv24_fs88_not0;
  wire f_arrdiv24_fs88_and0;
  wire f_arrdiv24_fs88_xor1;
  wire f_arrdiv24_fs88_not1;
  wire f_arrdiv24_fs88_and1;
  wire f_arrdiv24_fs88_or0;
  wire f_arrdiv24_fs89_xor0;
  wire f_arrdiv24_fs89_not0;
  wire f_arrdiv24_fs89_and0;
  wire f_arrdiv24_fs89_xor1;
  wire f_arrdiv24_fs89_not1;
  wire f_arrdiv24_fs89_and1;
  wire f_arrdiv24_fs89_or0;
  wire f_arrdiv24_fs90_xor0;
  wire f_arrdiv24_fs90_not0;
  wire f_arrdiv24_fs90_and0;
  wire f_arrdiv24_fs90_xor1;
  wire f_arrdiv24_fs90_not1;
  wire f_arrdiv24_fs90_and1;
  wire f_arrdiv24_fs90_or0;
  wire f_arrdiv24_fs91_xor0;
  wire f_arrdiv24_fs91_not0;
  wire f_arrdiv24_fs91_and0;
  wire f_arrdiv24_fs91_xor1;
  wire f_arrdiv24_fs91_not1;
  wire f_arrdiv24_fs91_and1;
  wire f_arrdiv24_fs91_or0;
  wire f_arrdiv24_fs92_xor0;
  wire f_arrdiv24_fs92_not0;
  wire f_arrdiv24_fs92_and0;
  wire f_arrdiv24_fs92_xor1;
  wire f_arrdiv24_fs92_not1;
  wire f_arrdiv24_fs92_and1;
  wire f_arrdiv24_fs92_or0;
  wire f_arrdiv24_fs93_xor0;
  wire f_arrdiv24_fs93_not0;
  wire f_arrdiv24_fs93_and0;
  wire f_arrdiv24_fs93_xor1;
  wire f_arrdiv24_fs93_not1;
  wire f_arrdiv24_fs93_and1;
  wire f_arrdiv24_fs93_or0;
  wire f_arrdiv24_fs94_xor0;
  wire f_arrdiv24_fs94_not0;
  wire f_arrdiv24_fs94_and0;
  wire f_arrdiv24_fs94_xor1;
  wire f_arrdiv24_fs94_not1;
  wire f_arrdiv24_fs94_and1;
  wire f_arrdiv24_fs94_or0;
  wire f_arrdiv24_fs95_xor0;
  wire f_arrdiv24_fs95_not0;
  wire f_arrdiv24_fs95_and0;
  wire f_arrdiv24_fs95_xor1;
  wire f_arrdiv24_fs95_not1;
  wire f_arrdiv24_fs95_and1;
  wire f_arrdiv24_fs95_or0;
  wire f_arrdiv24_mux2to169_and0;
  wire f_arrdiv24_mux2to169_not0;
  wire f_arrdiv24_mux2to169_and1;
  wire f_arrdiv24_mux2to169_xor0;
  wire f_arrdiv24_mux2to170_and0;
  wire f_arrdiv24_mux2to170_not0;
  wire f_arrdiv24_mux2to170_and1;
  wire f_arrdiv24_mux2to170_xor0;
  wire f_arrdiv24_mux2to171_and0;
  wire f_arrdiv24_mux2to171_not0;
  wire f_arrdiv24_mux2to171_and1;
  wire f_arrdiv24_mux2to171_xor0;
  wire f_arrdiv24_mux2to172_and0;
  wire f_arrdiv24_mux2to172_not0;
  wire f_arrdiv24_mux2to172_and1;
  wire f_arrdiv24_mux2to172_xor0;
  wire f_arrdiv24_mux2to173_and0;
  wire f_arrdiv24_mux2to173_not0;
  wire f_arrdiv24_mux2to173_and1;
  wire f_arrdiv24_mux2to173_xor0;
  wire f_arrdiv24_mux2to174_and0;
  wire f_arrdiv24_mux2to174_not0;
  wire f_arrdiv24_mux2to174_and1;
  wire f_arrdiv24_mux2to174_xor0;
  wire f_arrdiv24_mux2to175_and0;
  wire f_arrdiv24_mux2to175_not0;
  wire f_arrdiv24_mux2to175_and1;
  wire f_arrdiv24_mux2to175_xor0;
  wire f_arrdiv24_mux2to176_and0;
  wire f_arrdiv24_mux2to176_not0;
  wire f_arrdiv24_mux2to176_and1;
  wire f_arrdiv24_mux2to176_xor0;
  wire f_arrdiv24_mux2to177_and0;
  wire f_arrdiv24_mux2to177_not0;
  wire f_arrdiv24_mux2to177_and1;
  wire f_arrdiv24_mux2to177_xor0;
  wire f_arrdiv24_mux2to178_and0;
  wire f_arrdiv24_mux2to178_not0;
  wire f_arrdiv24_mux2to178_and1;
  wire f_arrdiv24_mux2to178_xor0;
  wire f_arrdiv24_mux2to179_and0;
  wire f_arrdiv24_mux2to179_not0;
  wire f_arrdiv24_mux2to179_and1;
  wire f_arrdiv24_mux2to179_xor0;
  wire f_arrdiv24_mux2to180_and0;
  wire f_arrdiv24_mux2to180_not0;
  wire f_arrdiv24_mux2to180_and1;
  wire f_arrdiv24_mux2to180_xor0;
  wire f_arrdiv24_mux2to181_and0;
  wire f_arrdiv24_mux2to181_not0;
  wire f_arrdiv24_mux2to181_and1;
  wire f_arrdiv24_mux2to181_xor0;
  wire f_arrdiv24_mux2to182_and0;
  wire f_arrdiv24_mux2to182_not0;
  wire f_arrdiv24_mux2to182_and1;
  wire f_arrdiv24_mux2to182_xor0;
  wire f_arrdiv24_mux2to183_and0;
  wire f_arrdiv24_mux2to183_not0;
  wire f_arrdiv24_mux2to183_and1;
  wire f_arrdiv24_mux2to183_xor0;
  wire f_arrdiv24_mux2to184_and0;
  wire f_arrdiv24_mux2to184_not0;
  wire f_arrdiv24_mux2to184_and1;
  wire f_arrdiv24_mux2to184_xor0;
  wire f_arrdiv24_mux2to185_and0;
  wire f_arrdiv24_mux2to185_not0;
  wire f_arrdiv24_mux2to185_and1;
  wire f_arrdiv24_mux2to185_xor0;
  wire f_arrdiv24_mux2to186_and0;
  wire f_arrdiv24_mux2to186_not0;
  wire f_arrdiv24_mux2to186_and1;
  wire f_arrdiv24_mux2to186_xor0;
  wire f_arrdiv24_mux2to187_and0;
  wire f_arrdiv24_mux2to187_not0;
  wire f_arrdiv24_mux2to187_and1;
  wire f_arrdiv24_mux2to187_xor0;
  wire f_arrdiv24_mux2to188_and0;
  wire f_arrdiv24_mux2to188_not0;
  wire f_arrdiv24_mux2to188_and1;
  wire f_arrdiv24_mux2to188_xor0;
  wire f_arrdiv24_mux2to189_and0;
  wire f_arrdiv24_mux2to189_not0;
  wire f_arrdiv24_mux2to189_and1;
  wire f_arrdiv24_mux2to189_xor0;
  wire f_arrdiv24_mux2to190_and0;
  wire f_arrdiv24_mux2to190_not0;
  wire f_arrdiv24_mux2to190_and1;
  wire f_arrdiv24_mux2to190_xor0;
  wire f_arrdiv24_mux2to191_and0;
  wire f_arrdiv24_mux2to191_not0;
  wire f_arrdiv24_mux2to191_and1;
  wire f_arrdiv24_mux2to191_xor0;
  wire f_arrdiv24_not3;
  wire f_arrdiv24_fs96_xor0;
  wire f_arrdiv24_fs96_not0;
  wire f_arrdiv24_fs96_and0;
  wire f_arrdiv24_fs96_not1;
  wire f_arrdiv24_fs97_xor0;
  wire f_arrdiv24_fs97_not0;
  wire f_arrdiv24_fs97_and0;
  wire f_arrdiv24_fs97_xor1;
  wire f_arrdiv24_fs97_not1;
  wire f_arrdiv24_fs97_and1;
  wire f_arrdiv24_fs97_or0;
  wire f_arrdiv24_fs98_xor0;
  wire f_arrdiv24_fs98_not0;
  wire f_arrdiv24_fs98_and0;
  wire f_arrdiv24_fs98_xor1;
  wire f_arrdiv24_fs98_not1;
  wire f_arrdiv24_fs98_and1;
  wire f_arrdiv24_fs98_or0;
  wire f_arrdiv24_fs99_xor0;
  wire f_arrdiv24_fs99_not0;
  wire f_arrdiv24_fs99_and0;
  wire f_arrdiv24_fs99_xor1;
  wire f_arrdiv24_fs99_not1;
  wire f_arrdiv24_fs99_and1;
  wire f_arrdiv24_fs99_or0;
  wire f_arrdiv24_fs100_xor0;
  wire f_arrdiv24_fs100_not0;
  wire f_arrdiv24_fs100_and0;
  wire f_arrdiv24_fs100_xor1;
  wire f_arrdiv24_fs100_not1;
  wire f_arrdiv24_fs100_and1;
  wire f_arrdiv24_fs100_or0;
  wire f_arrdiv24_fs101_xor0;
  wire f_arrdiv24_fs101_not0;
  wire f_arrdiv24_fs101_and0;
  wire f_arrdiv24_fs101_xor1;
  wire f_arrdiv24_fs101_not1;
  wire f_arrdiv24_fs101_and1;
  wire f_arrdiv24_fs101_or0;
  wire f_arrdiv24_fs102_xor0;
  wire f_arrdiv24_fs102_not0;
  wire f_arrdiv24_fs102_and0;
  wire f_arrdiv24_fs102_xor1;
  wire f_arrdiv24_fs102_not1;
  wire f_arrdiv24_fs102_and1;
  wire f_arrdiv24_fs102_or0;
  wire f_arrdiv24_fs103_xor0;
  wire f_arrdiv24_fs103_not0;
  wire f_arrdiv24_fs103_and0;
  wire f_arrdiv24_fs103_xor1;
  wire f_arrdiv24_fs103_not1;
  wire f_arrdiv24_fs103_and1;
  wire f_arrdiv24_fs103_or0;
  wire f_arrdiv24_fs104_xor0;
  wire f_arrdiv24_fs104_not0;
  wire f_arrdiv24_fs104_and0;
  wire f_arrdiv24_fs104_xor1;
  wire f_arrdiv24_fs104_not1;
  wire f_arrdiv24_fs104_and1;
  wire f_arrdiv24_fs104_or0;
  wire f_arrdiv24_fs105_xor0;
  wire f_arrdiv24_fs105_not0;
  wire f_arrdiv24_fs105_and0;
  wire f_arrdiv24_fs105_xor1;
  wire f_arrdiv24_fs105_not1;
  wire f_arrdiv24_fs105_and1;
  wire f_arrdiv24_fs105_or0;
  wire f_arrdiv24_fs106_xor0;
  wire f_arrdiv24_fs106_not0;
  wire f_arrdiv24_fs106_and0;
  wire f_arrdiv24_fs106_xor1;
  wire f_arrdiv24_fs106_not1;
  wire f_arrdiv24_fs106_and1;
  wire f_arrdiv24_fs106_or0;
  wire f_arrdiv24_fs107_xor0;
  wire f_arrdiv24_fs107_not0;
  wire f_arrdiv24_fs107_and0;
  wire f_arrdiv24_fs107_xor1;
  wire f_arrdiv24_fs107_not1;
  wire f_arrdiv24_fs107_and1;
  wire f_arrdiv24_fs107_or0;
  wire f_arrdiv24_fs108_xor0;
  wire f_arrdiv24_fs108_not0;
  wire f_arrdiv24_fs108_and0;
  wire f_arrdiv24_fs108_xor1;
  wire f_arrdiv24_fs108_not1;
  wire f_arrdiv24_fs108_and1;
  wire f_arrdiv24_fs108_or0;
  wire f_arrdiv24_fs109_xor0;
  wire f_arrdiv24_fs109_not0;
  wire f_arrdiv24_fs109_and0;
  wire f_arrdiv24_fs109_xor1;
  wire f_arrdiv24_fs109_not1;
  wire f_arrdiv24_fs109_and1;
  wire f_arrdiv24_fs109_or0;
  wire f_arrdiv24_fs110_xor0;
  wire f_arrdiv24_fs110_not0;
  wire f_arrdiv24_fs110_and0;
  wire f_arrdiv24_fs110_xor1;
  wire f_arrdiv24_fs110_not1;
  wire f_arrdiv24_fs110_and1;
  wire f_arrdiv24_fs110_or0;
  wire f_arrdiv24_fs111_xor0;
  wire f_arrdiv24_fs111_not0;
  wire f_arrdiv24_fs111_and0;
  wire f_arrdiv24_fs111_xor1;
  wire f_arrdiv24_fs111_not1;
  wire f_arrdiv24_fs111_and1;
  wire f_arrdiv24_fs111_or0;
  wire f_arrdiv24_fs112_xor0;
  wire f_arrdiv24_fs112_not0;
  wire f_arrdiv24_fs112_and0;
  wire f_arrdiv24_fs112_xor1;
  wire f_arrdiv24_fs112_not1;
  wire f_arrdiv24_fs112_and1;
  wire f_arrdiv24_fs112_or0;
  wire f_arrdiv24_fs113_xor0;
  wire f_arrdiv24_fs113_not0;
  wire f_arrdiv24_fs113_and0;
  wire f_arrdiv24_fs113_xor1;
  wire f_arrdiv24_fs113_not1;
  wire f_arrdiv24_fs113_and1;
  wire f_arrdiv24_fs113_or0;
  wire f_arrdiv24_fs114_xor0;
  wire f_arrdiv24_fs114_not0;
  wire f_arrdiv24_fs114_and0;
  wire f_arrdiv24_fs114_xor1;
  wire f_arrdiv24_fs114_not1;
  wire f_arrdiv24_fs114_and1;
  wire f_arrdiv24_fs114_or0;
  wire f_arrdiv24_fs115_xor0;
  wire f_arrdiv24_fs115_not0;
  wire f_arrdiv24_fs115_and0;
  wire f_arrdiv24_fs115_xor1;
  wire f_arrdiv24_fs115_not1;
  wire f_arrdiv24_fs115_and1;
  wire f_arrdiv24_fs115_or0;
  wire f_arrdiv24_fs116_xor0;
  wire f_arrdiv24_fs116_not0;
  wire f_arrdiv24_fs116_and0;
  wire f_arrdiv24_fs116_xor1;
  wire f_arrdiv24_fs116_not1;
  wire f_arrdiv24_fs116_and1;
  wire f_arrdiv24_fs116_or0;
  wire f_arrdiv24_fs117_xor0;
  wire f_arrdiv24_fs117_not0;
  wire f_arrdiv24_fs117_and0;
  wire f_arrdiv24_fs117_xor1;
  wire f_arrdiv24_fs117_not1;
  wire f_arrdiv24_fs117_and1;
  wire f_arrdiv24_fs117_or0;
  wire f_arrdiv24_fs118_xor0;
  wire f_arrdiv24_fs118_not0;
  wire f_arrdiv24_fs118_and0;
  wire f_arrdiv24_fs118_xor1;
  wire f_arrdiv24_fs118_not1;
  wire f_arrdiv24_fs118_and1;
  wire f_arrdiv24_fs118_or0;
  wire f_arrdiv24_fs119_xor0;
  wire f_arrdiv24_fs119_not0;
  wire f_arrdiv24_fs119_and0;
  wire f_arrdiv24_fs119_xor1;
  wire f_arrdiv24_fs119_not1;
  wire f_arrdiv24_fs119_and1;
  wire f_arrdiv24_fs119_or0;
  wire f_arrdiv24_mux2to192_and0;
  wire f_arrdiv24_mux2to192_not0;
  wire f_arrdiv24_mux2to192_and1;
  wire f_arrdiv24_mux2to192_xor0;
  wire f_arrdiv24_mux2to193_and0;
  wire f_arrdiv24_mux2to193_not0;
  wire f_arrdiv24_mux2to193_and1;
  wire f_arrdiv24_mux2to193_xor0;
  wire f_arrdiv24_mux2to194_and0;
  wire f_arrdiv24_mux2to194_not0;
  wire f_arrdiv24_mux2to194_and1;
  wire f_arrdiv24_mux2to194_xor0;
  wire f_arrdiv24_mux2to195_and0;
  wire f_arrdiv24_mux2to195_not0;
  wire f_arrdiv24_mux2to195_and1;
  wire f_arrdiv24_mux2to195_xor0;
  wire f_arrdiv24_mux2to196_and0;
  wire f_arrdiv24_mux2to196_not0;
  wire f_arrdiv24_mux2to196_and1;
  wire f_arrdiv24_mux2to196_xor0;
  wire f_arrdiv24_mux2to197_and0;
  wire f_arrdiv24_mux2to197_not0;
  wire f_arrdiv24_mux2to197_and1;
  wire f_arrdiv24_mux2to197_xor0;
  wire f_arrdiv24_mux2to198_and0;
  wire f_arrdiv24_mux2to198_not0;
  wire f_arrdiv24_mux2to198_and1;
  wire f_arrdiv24_mux2to198_xor0;
  wire f_arrdiv24_mux2to199_and0;
  wire f_arrdiv24_mux2to199_not0;
  wire f_arrdiv24_mux2to199_and1;
  wire f_arrdiv24_mux2to199_xor0;
  wire f_arrdiv24_mux2to1100_and0;
  wire f_arrdiv24_mux2to1100_not0;
  wire f_arrdiv24_mux2to1100_and1;
  wire f_arrdiv24_mux2to1100_xor0;
  wire f_arrdiv24_mux2to1101_and0;
  wire f_arrdiv24_mux2to1101_not0;
  wire f_arrdiv24_mux2to1101_and1;
  wire f_arrdiv24_mux2to1101_xor0;
  wire f_arrdiv24_mux2to1102_and0;
  wire f_arrdiv24_mux2to1102_not0;
  wire f_arrdiv24_mux2to1102_and1;
  wire f_arrdiv24_mux2to1102_xor0;
  wire f_arrdiv24_mux2to1103_and0;
  wire f_arrdiv24_mux2to1103_not0;
  wire f_arrdiv24_mux2to1103_and1;
  wire f_arrdiv24_mux2to1103_xor0;
  wire f_arrdiv24_mux2to1104_and0;
  wire f_arrdiv24_mux2to1104_not0;
  wire f_arrdiv24_mux2to1104_and1;
  wire f_arrdiv24_mux2to1104_xor0;
  wire f_arrdiv24_mux2to1105_and0;
  wire f_arrdiv24_mux2to1105_not0;
  wire f_arrdiv24_mux2to1105_and1;
  wire f_arrdiv24_mux2to1105_xor0;
  wire f_arrdiv24_mux2to1106_and0;
  wire f_arrdiv24_mux2to1106_not0;
  wire f_arrdiv24_mux2to1106_and1;
  wire f_arrdiv24_mux2to1106_xor0;
  wire f_arrdiv24_mux2to1107_and0;
  wire f_arrdiv24_mux2to1107_not0;
  wire f_arrdiv24_mux2to1107_and1;
  wire f_arrdiv24_mux2to1107_xor0;
  wire f_arrdiv24_mux2to1108_and0;
  wire f_arrdiv24_mux2to1108_not0;
  wire f_arrdiv24_mux2to1108_and1;
  wire f_arrdiv24_mux2to1108_xor0;
  wire f_arrdiv24_mux2to1109_and0;
  wire f_arrdiv24_mux2to1109_not0;
  wire f_arrdiv24_mux2to1109_and1;
  wire f_arrdiv24_mux2to1109_xor0;
  wire f_arrdiv24_mux2to1110_and0;
  wire f_arrdiv24_mux2to1110_not0;
  wire f_arrdiv24_mux2to1110_and1;
  wire f_arrdiv24_mux2to1110_xor0;
  wire f_arrdiv24_mux2to1111_and0;
  wire f_arrdiv24_mux2to1111_not0;
  wire f_arrdiv24_mux2to1111_and1;
  wire f_arrdiv24_mux2to1111_xor0;
  wire f_arrdiv24_mux2to1112_and0;
  wire f_arrdiv24_mux2to1112_not0;
  wire f_arrdiv24_mux2to1112_and1;
  wire f_arrdiv24_mux2to1112_xor0;
  wire f_arrdiv24_mux2to1113_and0;
  wire f_arrdiv24_mux2to1113_not0;
  wire f_arrdiv24_mux2to1113_and1;
  wire f_arrdiv24_mux2to1113_xor0;
  wire f_arrdiv24_mux2to1114_and0;
  wire f_arrdiv24_mux2to1114_not0;
  wire f_arrdiv24_mux2to1114_and1;
  wire f_arrdiv24_mux2to1114_xor0;
  wire f_arrdiv24_not4;
  wire f_arrdiv24_fs120_xor0;
  wire f_arrdiv24_fs120_not0;
  wire f_arrdiv24_fs120_and0;
  wire f_arrdiv24_fs120_not1;
  wire f_arrdiv24_fs121_xor0;
  wire f_arrdiv24_fs121_not0;
  wire f_arrdiv24_fs121_and0;
  wire f_arrdiv24_fs121_xor1;
  wire f_arrdiv24_fs121_not1;
  wire f_arrdiv24_fs121_and1;
  wire f_arrdiv24_fs121_or0;
  wire f_arrdiv24_fs122_xor0;
  wire f_arrdiv24_fs122_not0;
  wire f_arrdiv24_fs122_and0;
  wire f_arrdiv24_fs122_xor1;
  wire f_arrdiv24_fs122_not1;
  wire f_arrdiv24_fs122_and1;
  wire f_arrdiv24_fs122_or0;
  wire f_arrdiv24_fs123_xor0;
  wire f_arrdiv24_fs123_not0;
  wire f_arrdiv24_fs123_and0;
  wire f_arrdiv24_fs123_xor1;
  wire f_arrdiv24_fs123_not1;
  wire f_arrdiv24_fs123_and1;
  wire f_arrdiv24_fs123_or0;
  wire f_arrdiv24_fs124_xor0;
  wire f_arrdiv24_fs124_not0;
  wire f_arrdiv24_fs124_and0;
  wire f_arrdiv24_fs124_xor1;
  wire f_arrdiv24_fs124_not1;
  wire f_arrdiv24_fs124_and1;
  wire f_arrdiv24_fs124_or0;
  wire f_arrdiv24_fs125_xor0;
  wire f_arrdiv24_fs125_not0;
  wire f_arrdiv24_fs125_and0;
  wire f_arrdiv24_fs125_xor1;
  wire f_arrdiv24_fs125_not1;
  wire f_arrdiv24_fs125_and1;
  wire f_arrdiv24_fs125_or0;
  wire f_arrdiv24_fs126_xor0;
  wire f_arrdiv24_fs126_not0;
  wire f_arrdiv24_fs126_and0;
  wire f_arrdiv24_fs126_xor1;
  wire f_arrdiv24_fs126_not1;
  wire f_arrdiv24_fs126_and1;
  wire f_arrdiv24_fs126_or0;
  wire f_arrdiv24_fs127_xor0;
  wire f_arrdiv24_fs127_not0;
  wire f_arrdiv24_fs127_and0;
  wire f_arrdiv24_fs127_xor1;
  wire f_arrdiv24_fs127_not1;
  wire f_arrdiv24_fs127_and1;
  wire f_arrdiv24_fs127_or0;
  wire f_arrdiv24_fs128_xor0;
  wire f_arrdiv24_fs128_not0;
  wire f_arrdiv24_fs128_and0;
  wire f_arrdiv24_fs128_xor1;
  wire f_arrdiv24_fs128_not1;
  wire f_arrdiv24_fs128_and1;
  wire f_arrdiv24_fs128_or0;
  wire f_arrdiv24_fs129_xor0;
  wire f_arrdiv24_fs129_not0;
  wire f_arrdiv24_fs129_and0;
  wire f_arrdiv24_fs129_xor1;
  wire f_arrdiv24_fs129_not1;
  wire f_arrdiv24_fs129_and1;
  wire f_arrdiv24_fs129_or0;
  wire f_arrdiv24_fs130_xor0;
  wire f_arrdiv24_fs130_not0;
  wire f_arrdiv24_fs130_and0;
  wire f_arrdiv24_fs130_xor1;
  wire f_arrdiv24_fs130_not1;
  wire f_arrdiv24_fs130_and1;
  wire f_arrdiv24_fs130_or0;
  wire f_arrdiv24_fs131_xor0;
  wire f_arrdiv24_fs131_not0;
  wire f_arrdiv24_fs131_and0;
  wire f_arrdiv24_fs131_xor1;
  wire f_arrdiv24_fs131_not1;
  wire f_arrdiv24_fs131_and1;
  wire f_arrdiv24_fs131_or0;
  wire f_arrdiv24_fs132_xor0;
  wire f_arrdiv24_fs132_not0;
  wire f_arrdiv24_fs132_and0;
  wire f_arrdiv24_fs132_xor1;
  wire f_arrdiv24_fs132_not1;
  wire f_arrdiv24_fs132_and1;
  wire f_arrdiv24_fs132_or0;
  wire f_arrdiv24_fs133_xor0;
  wire f_arrdiv24_fs133_not0;
  wire f_arrdiv24_fs133_and0;
  wire f_arrdiv24_fs133_xor1;
  wire f_arrdiv24_fs133_not1;
  wire f_arrdiv24_fs133_and1;
  wire f_arrdiv24_fs133_or0;
  wire f_arrdiv24_fs134_xor0;
  wire f_arrdiv24_fs134_not0;
  wire f_arrdiv24_fs134_and0;
  wire f_arrdiv24_fs134_xor1;
  wire f_arrdiv24_fs134_not1;
  wire f_arrdiv24_fs134_and1;
  wire f_arrdiv24_fs134_or0;
  wire f_arrdiv24_fs135_xor0;
  wire f_arrdiv24_fs135_not0;
  wire f_arrdiv24_fs135_and0;
  wire f_arrdiv24_fs135_xor1;
  wire f_arrdiv24_fs135_not1;
  wire f_arrdiv24_fs135_and1;
  wire f_arrdiv24_fs135_or0;
  wire f_arrdiv24_fs136_xor0;
  wire f_arrdiv24_fs136_not0;
  wire f_arrdiv24_fs136_and0;
  wire f_arrdiv24_fs136_xor1;
  wire f_arrdiv24_fs136_not1;
  wire f_arrdiv24_fs136_and1;
  wire f_arrdiv24_fs136_or0;
  wire f_arrdiv24_fs137_xor0;
  wire f_arrdiv24_fs137_not0;
  wire f_arrdiv24_fs137_and0;
  wire f_arrdiv24_fs137_xor1;
  wire f_arrdiv24_fs137_not1;
  wire f_arrdiv24_fs137_and1;
  wire f_arrdiv24_fs137_or0;
  wire f_arrdiv24_fs138_xor0;
  wire f_arrdiv24_fs138_not0;
  wire f_arrdiv24_fs138_and0;
  wire f_arrdiv24_fs138_xor1;
  wire f_arrdiv24_fs138_not1;
  wire f_arrdiv24_fs138_and1;
  wire f_arrdiv24_fs138_or0;
  wire f_arrdiv24_fs139_xor0;
  wire f_arrdiv24_fs139_not0;
  wire f_arrdiv24_fs139_and0;
  wire f_arrdiv24_fs139_xor1;
  wire f_arrdiv24_fs139_not1;
  wire f_arrdiv24_fs139_and1;
  wire f_arrdiv24_fs139_or0;
  wire f_arrdiv24_fs140_xor0;
  wire f_arrdiv24_fs140_not0;
  wire f_arrdiv24_fs140_and0;
  wire f_arrdiv24_fs140_xor1;
  wire f_arrdiv24_fs140_not1;
  wire f_arrdiv24_fs140_and1;
  wire f_arrdiv24_fs140_or0;
  wire f_arrdiv24_fs141_xor0;
  wire f_arrdiv24_fs141_not0;
  wire f_arrdiv24_fs141_and0;
  wire f_arrdiv24_fs141_xor1;
  wire f_arrdiv24_fs141_not1;
  wire f_arrdiv24_fs141_and1;
  wire f_arrdiv24_fs141_or0;
  wire f_arrdiv24_fs142_xor0;
  wire f_arrdiv24_fs142_not0;
  wire f_arrdiv24_fs142_and0;
  wire f_arrdiv24_fs142_xor1;
  wire f_arrdiv24_fs142_not1;
  wire f_arrdiv24_fs142_and1;
  wire f_arrdiv24_fs142_or0;
  wire f_arrdiv24_fs143_xor0;
  wire f_arrdiv24_fs143_not0;
  wire f_arrdiv24_fs143_and0;
  wire f_arrdiv24_fs143_xor1;
  wire f_arrdiv24_fs143_not1;
  wire f_arrdiv24_fs143_and1;
  wire f_arrdiv24_fs143_or0;
  wire f_arrdiv24_mux2to1115_and0;
  wire f_arrdiv24_mux2to1115_not0;
  wire f_arrdiv24_mux2to1115_and1;
  wire f_arrdiv24_mux2to1115_xor0;
  wire f_arrdiv24_mux2to1116_and0;
  wire f_arrdiv24_mux2to1116_not0;
  wire f_arrdiv24_mux2to1116_and1;
  wire f_arrdiv24_mux2to1116_xor0;
  wire f_arrdiv24_mux2to1117_and0;
  wire f_arrdiv24_mux2to1117_not0;
  wire f_arrdiv24_mux2to1117_and1;
  wire f_arrdiv24_mux2to1117_xor0;
  wire f_arrdiv24_mux2to1118_and0;
  wire f_arrdiv24_mux2to1118_not0;
  wire f_arrdiv24_mux2to1118_and1;
  wire f_arrdiv24_mux2to1118_xor0;
  wire f_arrdiv24_mux2to1119_and0;
  wire f_arrdiv24_mux2to1119_not0;
  wire f_arrdiv24_mux2to1119_and1;
  wire f_arrdiv24_mux2to1119_xor0;
  wire f_arrdiv24_mux2to1120_and0;
  wire f_arrdiv24_mux2to1120_not0;
  wire f_arrdiv24_mux2to1120_and1;
  wire f_arrdiv24_mux2to1120_xor0;
  wire f_arrdiv24_mux2to1121_and0;
  wire f_arrdiv24_mux2to1121_not0;
  wire f_arrdiv24_mux2to1121_and1;
  wire f_arrdiv24_mux2to1121_xor0;
  wire f_arrdiv24_mux2to1122_and0;
  wire f_arrdiv24_mux2to1122_not0;
  wire f_arrdiv24_mux2to1122_and1;
  wire f_arrdiv24_mux2to1122_xor0;
  wire f_arrdiv24_mux2to1123_and0;
  wire f_arrdiv24_mux2to1123_not0;
  wire f_arrdiv24_mux2to1123_and1;
  wire f_arrdiv24_mux2to1123_xor0;
  wire f_arrdiv24_mux2to1124_and0;
  wire f_arrdiv24_mux2to1124_not0;
  wire f_arrdiv24_mux2to1124_and1;
  wire f_arrdiv24_mux2to1124_xor0;
  wire f_arrdiv24_mux2to1125_and0;
  wire f_arrdiv24_mux2to1125_not0;
  wire f_arrdiv24_mux2to1125_and1;
  wire f_arrdiv24_mux2to1125_xor0;
  wire f_arrdiv24_mux2to1126_and0;
  wire f_arrdiv24_mux2to1126_not0;
  wire f_arrdiv24_mux2to1126_and1;
  wire f_arrdiv24_mux2to1126_xor0;
  wire f_arrdiv24_mux2to1127_and0;
  wire f_arrdiv24_mux2to1127_not0;
  wire f_arrdiv24_mux2to1127_and1;
  wire f_arrdiv24_mux2to1127_xor0;
  wire f_arrdiv24_mux2to1128_and0;
  wire f_arrdiv24_mux2to1128_not0;
  wire f_arrdiv24_mux2to1128_and1;
  wire f_arrdiv24_mux2to1128_xor0;
  wire f_arrdiv24_mux2to1129_and0;
  wire f_arrdiv24_mux2to1129_not0;
  wire f_arrdiv24_mux2to1129_and1;
  wire f_arrdiv24_mux2to1129_xor0;
  wire f_arrdiv24_mux2to1130_and0;
  wire f_arrdiv24_mux2to1130_not0;
  wire f_arrdiv24_mux2to1130_and1;
  wire f_arrdiv24_mux2to1130_xor0;
  wire f_arrdiv24_mux2to1131_and0;
  wire f_arrdiv24_mux2to1131_not0;
  wire f_arrdiv24_mux2to1131_and1;
  wire f_arrdiv24_mux2to1131_xor0;
  wire f_arrdiv24_mux2to1132_and0;
  wire f_arrdiv24_mux2to1132_not0;
  wire f_arrdiv24_mux2to1132_and1;
  wire f_arrdiv24_mux2to1132_xor0;
  wire f_arrdiv24_mux2to1133_and0;
  wire f_arrdiv24_mux2to1133_not0;
  wire f_arrdiv24_mux2to1133_and1;
  wire f_arrdiv24_mux2to1133_xor0;
  wire f_arrdiv24_mux2to1134_and0;
  wire f_arrdiv24_mux2to1134_not0;
  wire f_arrdiv24_mux2to1134_and1;
  wire f_arrdiv24_mux2to1134_xor0;
  wire f_arrdiv24_mux2to1135_and0;
  wire f_arrdiv24_mux2to1135_not0;
  wire f_arrdiv24_mux2to1135_and1;
  wire f_arrdiv24_mux2to1135_xor0;
  wire f_arrdiv24_mux2to1136_and0;
  wire f_arrdiv24_mux2to1136_not0;
  wire f_arrdiv24_mux2to1136_and1;
  wire f_arrdiv24_mux2to1136_xor0;
  wire f_arrdiv24_mux2to1137_and0;
  wire f_arrdiv24_mux2to1137_not0;
  wire f_arrdiv24_mux2to1137_and1;
  wire f_arrdiv24_mux2to1137_xor0;
  wire f_arrdiv24_not5;
  wire f_arrdiv24_fs144_xor0;
  wire f_arrdiv24_fs144_not0;
  wire f_arrdiv24_fs144_and0;
  wire f_arrdiv24_fs144_not1;
  wire f_arrdiv24_fs145_xor0;
  wire f_arrdiv24_fs145_not0;
  wire f_arrdiv24_fs145_and0;
  wire f_arrdiv24_fs145_xor1;
  wire f_arrdiv24_fs145_not1;
  wire f_arrdiv24_fs145_and1;
  wire f_arrdiv24_fs145_or0;
  wire f_arrdiv24_fs146_xor0;
  wire f_arrdiv24_fs146_not0;
  wire f_arrdiv24_fs146_and0;
  wire f_arrdiv24_fs146_xor1;
  wire f_arrdiv24_fs146_not1;
  wire f_arrdiv24_fs146_and1;
  wire f_arrdiv24_fs146_or0;
  wire f_arrdiv24_fs147_xor0;
  wire f_arrdiv24_fs147_not0;
  wire f_arrdiv24_fs147_and0;
  wire f_arrdiv24_fs147_xor1;
  wire f_arrdiv24_fs147_not1;
  wire f_arrdiv24_fs147_and1;
  wire f_arrdiv24_fs147_or0;
  wire f_arrdiv24_fs148_xor0;
  wire f_arrdiv24_fs148_not0;
  wire f_arrdiv24_fs148_and0;
  wire f_arrdiv24_fs148_xor1;
  wire f_arrdiv24_fs148_not1;
  wire f_arrdiv24_fs148_and1;
  wire f_arrdiv24_fs148_or0;
  wire f_arrdiv24_fs149_xor0;
  wire f_arrdiv24_fs149_not0;
  wire f_arrdiv24_fs149_and0;
  wire f_arrdiv24_fs149_xor1;
  wire f_arrdiv24_fs149_not1;
  wire f_arrdiv24_fs149_and1;
  wire f_arrdiv24_fs149_or0;
  wire f_arrdiv24_fs150_xor0;
  wire f_arrdiv24_fs150_not0;
  wire f_arrdiv24_fs150_and0;
  wire f_arrdiv24_fs150_xor1;
  wire f_arrdiv24_fs150_not1;
  wire f_arrdiv24_fs150_and1;
  wire f_arrdiv24_fs150_or0;
  wire f_arrdiv24_fs151_xor0;
  wire f_arrdiv24_fs151_not0;
  wire f_arrdiv24_fs151_and0;
  wire f_arrdiv24_fs151_xor1;
  wire f_arrdiv24_fs151_not1;
  wire f_arrdiv24_fs151_and1;
  wire f_arrdiv24_fs151_or0;
  wire f_arrdiv24_fs152_xor0;
  wire f_arrdiv24_fs152_not0;
  wire f_arrdiv24_fs152_and0;
  wire f_arrdiv24_fs152_xor1;
  wire f_arrdiv24_fs152_not1;
  wire f_arrdiv24_fs152_and1;
  wire f_arrdiv24_fs152_or0;
  wire f_arrdiv24_fs153_xor0;
  wire f_arrdiv24_fs153_not0;
  wire f_arrdiv24_fs153_and0;
  wire f_arrdiv24_fs153_xor1;
  wire f_arrdiv24_fs153_not1;
  wire f_arrdiv24_fs153_and1;
  wire f_arrdiv24_fs153_or0;
  wire f_arrdiv24_fs154_xor0;
  wire f_arrdiv24_fs154_not0;
  wire f_arrdiv24_fs154_and0;
  wire f_arrdiv24_fs154_xor1;
  wire f_arrdiv24_fs154_not1;
  wire f_arrdiv24_fs154_and1;
  wire f_arrdiv24_fs154_or0;
  wire f_arrdiv24_fs155_xor0;
  wire f_arrdiv24_fs155_not0;
  wire f_arrdiv24_fs155_and0;
  wire f_arrdiv24_fs155_xor1;
  wire f_arrdiv24_fs155_not1;
  wire f_arrdiv24_fs155_and1;
  wire f_arrdiv24_fs155_or0;
  wire f_arrdiv24_fs156_xor0;
  wire f_arrdiv24_fs156_not0;
  wire f_arrdiv24_fs156_and0;
  wire f_arrdiv24_fs156_xor1;
  wire f_arrdiv24_fs156_not1;
  wire f_arrdiv24_fs156_and1;
  wire f_arrdiv24_fs156_or0;
  wire f_arrdiv24_fs157_xor0;
  wire f_arrdiv24_fs157_not0;
  wire f_arrdiv24_fs157_and0;
  wire f_arrdiv24_fs157_xor1;
  wire f_arrdiv24_fs157_not1;
  wire f_arrdiv24_fs157_and1;
  wire f_arrdiv24_fs157_or0;
  wire f_arrdiv24_fs158_xor0;
  wire f_arrdiv24_fs158_not0;
  wire f_arrdiv24_fs158_and0;
  wire f_arrdiv24_fs158_xor1;
  wire f_arrdiv24_fs158_not1;
  wire f_arrdiv24_fs158_and1;
  wire f_arrdiv24_fs158_or0;
  wire f_arrdiv24_fs159_xor0;
  wire f_arrdiv24_fs159_not0;
  wire f_arrdiv24_fs159_and0;
  wire f_arrdiv24_fs159_xor1;
  wire f_arrdiv24_fs159_not1;
  wire f_arrdiv24_fs159_and1;
  wire f_arrdiv24_fs159_or0;
  wire f_arrdiv24_fs160_xor0;
  wire f_arrdiv24_fs160_not0;
  wire f_arrdiv24_fs160_and0;
  wire f_arrdiv24_fs160_xor1;
  wire f_arrdiv24_fs160_not1;
  wire f_arrdiv24_fs160_and1;
  wire f_arrdiv24_fs160_or0;
  wire f_arrdiv24_fs161_xor0;
  wire f_arrdiv24_fs161_not0;
  wire f_arrdiv24_fs161_and0;
  wire f_arrdiv24_fs161_xor1;
  wire f_arrdiv24_fs161_not1;
  wire f_arrdiv24_fs161_and1;
  wire f_arrdiv24_fs161_or0;
  wire f_arrdiv24_fs162_xor0;
  wire f_arrdiv24_fs162_not0;
  wire f_arrdiv24_fs162_and0;
  wire f_arrdiv24_fs162_xor1;
  wire f_arrdiv24_fs162_not1;
  wire f_arrdiv24_fs162_and1;
  wire f_arrdiv24_fs162_or0;
  wire f_arrdiv24_fs163_xor0;
  wire f_arrdiv24_fs163_not0;
  wire f_arrdiv24_fs163_and0;
  wire f_arrdiv24_fs163_xor1;
  wire f_arrdiv24_fs163_not1;
  wire f_arrdiv24_fs163_and1;
  wire f_arrdiv24_fs163_or0;
  wire f_arrdiv24_fs164_xor0;
  wire f_arrdiv24_fs164_not0;
  wire f_arrdiv24_fs164_and0;
  wire f_arrdiv24_fs164_xor1;
  wire f_arrdiv24_fs164_not1;
  wire f_arrdiv24_fs164_and1;
  wire f_arrdiv24_fs164_or0;
  wire f_arrdiv24_fs165_xor0;
  wire f_arrdiv24_fs165_not0;
  wire f_arrdiv24_fs165_and0;
  wire f_arrdiv24_fs165_xor1;
  wire f_arrdiv24_fs165_not1;
  wire f_arrdiv24_fs165_and1;
  wire f_arrdiv24_fs165_or0;
  wire f_arrdiv24_fs166_xor0;
  wire f_arrdiv24_fs166_not0;
  wire f_arrdiv24_fs166_and0;
  wire f_arrdiv24_fs166_xor1;
  wire f_arrdiv24_fs166_not1;
  wire f_arrdiv24_fs166_and1;
  wire f_arrdiv24_fs166_or0;
  wire f_arrdiv24_fs167_xor0;
  wire f_arrdiv24_fs167_not0;
  wire f_arrdiv24_fs167_and0;
  wire f_arrdiv24_fs167_xor1;
  wire f_arrdiv24_fs167_not1;
  wire f_arrdiv24_fs167_and1;
  wire f_arrdiv24_fs167_or0;
  wire f_arrdiv24_mux2to1138_and0;
  wire f_arrdiv24_mux2to1138_not0;
  wire f_arrdiv24_mux2to1138_and1;
  wire f_arrdiv24_mux2to1138_xor0;
  wire f_arrdiv24_mux2to1139_and0;
  wire f_arrdiv24_mux2to1139_not0;
  wire f_arrdiv24_mux2to1139_and1;
  wire f_arrdiv24_mux2to1139_xor0;
  wire f_arrdiv24_mux2to1140_and0;
  wire f_arrdiv24_mux2to1140_not0;
  wire f_arrdiv24_mux2to1140_and1;
  wire f_arrdiv24_mux2to1140_xor0;
  wire f_arrdiv24_mux2to1141_and0;
  wire f_arrdiv24_mux2to1141_not0;
  wire f_arrdiv24_mux2to1141_and1;
  wire f_arrdiv24_mux2to1141_xor0;
  wire f_arrdiv24_mux2to1142_and0;
  wire f_arrdiv24_mux2to1142_not0;
  wire f_arrdiv24_mux2to1142_and1;
  wire f_arrdiv24_mux2to1142_xor0;
  wire f_arrdiv24_mux2to1143_and0;
  wire f_arrdiv24_mux2to1143_not0;
  wire f_arrdiv24_mux2to1143_and1;
  wire f_arrdiv24_mux2to1143_xor0;
  wire f_arrdiv24_mux2to1144_and0;
  wire f_arrdiv24_mux2to1144_not0;
  wire f_arrdiv24_mux2to1144_and1;
  wire f_arrdiv24_mux2to1144_xor0;
  wire f_arrdiv24_mux2to1145_and0;
  wire f_arrdiv24_mux2to1145_not0;
  wire f_arrdiv24_mux2to1145_and1;
  wire f_arrdiv24_mux2to1145_xor0;
  wire f_arrdiv24_mux2to1146_and0;
  wire f_arrdiv24_mux2to1146_not0;
  wire f_arrdiv24_mux2to1146_and1;
  wire f_arrdiv24_mux2to1146_xor0;
  wire f_arrdiv24_mux2to1147_and0;
  wire f_arrdiv24_mux2to1147_not0;
  wire f_arrdiv24_mux2to1147_and1;
  wire f_arrdiv24_mux2to1147_xor0;
  wire f_arrdiv24_mux2to1148_and0;
  wire f_arrdiv24_mux2to1148_not0;
  wire f_arrdiv24_mux2to1148_and1;
  wire f_arrdiv24_mux2to1148_xor0;
  wire f_arrdiv24_mux2to1149_and0;
  wire f_arrdiv24_mux2to1149_not0;
  wire f_arrdiv24_mux2to1149_and1;
  wire f_arrdiv24_mux2to1149_xor0;
  wire f_arrdiv24_mux2to1150_and0;
  wire f_arrdiv24_mux2to1150_not0;
  wire f_arrdiv24_mux2to1150_and1;
  wire f_arrdiv24_mux2to1150_xor0;
  wire f_arrdiv24_mux2to1151_and0;
  wire f_arrdiv24_mux2to1151_not0;
  wire f_arrdiv24_mux2to1151_and1;
  wire f_arrdiv24_mux2to1151_xor0;
  wire f_arrdiv24_mux2to1152_and0;
  wire f_arrdiv24_mux2to1152_not0;
  wire f_arrdiv24_mux2to1152_and1;
  wire f_arrdiv24_mux2to1152_xor0;
  wire f_arrdiv24_mux2to1153_and0;
  wire f_arrdiv24_mux2to1153_not0;
  wire f_arrdiv24_mux2to1153_and1;
  wire f_arrdiv24_mux2to1153_xor0;
  wire f_arrdiv24_mux2to1154_and0;
  wire f_arrdiv24_mux2to1154_not0;
  wire f_arrdiv24_mux2to1154_and1;
  wire f_arrdiv24_mux2to1154_xor0;
  wire f_arrdiv24_mux2to1155_and0;
  wire f_arrdiv24_mux2to1155_not0;
  wire f_arrdiv24_mux2to1155_and1;
  wire f_arrdiv24_mux2to1155_xor0;
  wire f_arrdiv24_mux2to1156_and0;
  wire f_arrdiv24_mux2to1156_not0;
  wire f_arrdiv24_mux2to1156_and1;
  wire f_arrdiv24_mux2to1156_xor0;
  wire f_arrdiv24_mux2to1157_and0;
  wire f_arrdiv24_mux2to1157_not0;
  wire f_arrdiv24_mux2to1157_and1;
  wire f_arrdiv24_mux2to1157_xor0;
  wire f_arrdiv24_mux2to1158_and0;
  wire f_arrdiv24_mux2to1158_not0;
  wire f_arrdiv24_mux2to1158_and1;
  wire f_arrdiv24_mux2to1158_xor0;
  wire f_arrdiv24_mux2to1159_and0;
  wire f_arrdiv24_mux2to1159_not0;
  wire f_arrdiv24_mux2to1159_and1;
  wire f_arrdiv24_mux2to1159_xor0;
  wire f_arrdiv24_mux2to1160_and0;
  wire f_arrdiv24_mux2to1160_not0;
  wire f_arrdiv24_mux2to1160_and1;
  wire f_arrdiv24_mux2to1160_xor0;
  wire f_arrdiv24_not6;
  wire f_arrdiv24_fs168_xor0;
  wire f_arrdiv24_fs168_not0;
  wire f_arrdiv24_fs168_and0;
  wire f_arrdiv24_fs168_not1;
  wire f_arrdiv24_fs169_xor0;
  wire f_arrdiv24_fs169_not0;
  wire f_arrdiv24_fs169_and0;
  wire f_arrdiv24_fs169_xor1;
  wire f_arrdiv24_fs169_not1;
  wire f_arrdiv24_fs169_and1;
  wire f_arrdiv24_fs169_or0;
  wire f_arrdiv24_fs170_xor0;
  wire f_arrdiv24_fs170_not0;
  wire f_arrdiv24_fs170_and0;
  wire f_arrdiv24_fs170_xor1;
  wire f_arrdiv24_fs170_not1;
  wire f_arrdiv24_fs170_and1;
  wire f_arrdiv24_fs170_or0;
  wire f_arrdiv24_fs171_xor0;
  wire f_arrdiv24_fs171_not0;
  wire f_arrdiv24_fs171_and0;
  wire f_arrdiv24_fs171_xor1;
  wire f_arrdiv24_fs171_not1;
  wire f_arrdiv24_fs171_and1;
  wire f_arrdiv24_fs171_or0;
  wire f_arrdiv24_fs172_xor0;
  wire f_arrdiv24_fs172_not0;
  wire f_arrdiv24_fs172_and0;
  wire f_arrdiv24_fs172_xor1;
  wire f_arrdiv24_fs172_not1;
  wire f_arrdiv24_fs172_and1;
  wire f_arrdiv24_fs172_or0;
  wire f_arrdiv24_fs173_xor0;
  wire f_arrdiv24_fs173_not0;
  wire f_arrdiv24_fs173_and0;
  wire f_arrdiv24_fs173_xor1;
  wire f_arrdiv24_fs173_not1;
  wire f_arrdiv24_fs173_and1;
  wire f_arrdiv24_fs173_or0;
  wire f_arrdiv24_fs174_xor0;
  wire f_arrdiv24_fs174_not0;
  wire f_arrdiv24_fs174_and0;
  wire f_arrdiv24_fs174_xor1;
  wire f_arrdiv24_fs174_not1;
  wire f_arrdiv24_fs174_and1;
  wire f_arrdiv24_fs174_or0;
  wire f_arrdiv24_fs175_xor0;
  wire f_arrdiv24_fs175_not0;
  wire f_arrdiv24_fs175_and0;
  wire f_arrdiv24_fs175_xor1;
  wire f_arrdiv24_fs175_not1;
  wire f_arrdiv24_fs175_and1;
  wire f_arrdiv24_fs175_or0;
  wire f_arrdiv24_fs176_xor0;
  wire f_arrdiv24_fs176_not0;
  wire f_arrdiv24_fs176_and0;
  wire f_arrdiv24_fs176_xor1;
  wire f_arrdiv24_fs176_not1;
  wire f_arrdiv24_fs176_and1;
  wire f_arrdiv24_fs176_or0;
  wire f_arrdiv24_fs177_xor0;
  wire f_arrdiv24_fs177_not0;
  wire f_arrdiv24_fs177_and0;
  wire f_arrdiv24_fs177_xor1;
  wire f_arrdiv24_fs177_not1;
  wire f_arrdiv24_fs177_and1;
  wire f_arrdiv24_fs177_or0;
  wire f_arrdiv24_fs178_xor0;
  wire f_arrdiv24_fs178_not0;
  wire f_arrdiv24_fs178_and0;
  wire f_arrdiv24_fs178_xor1;
  wire f_arrdiv24_fs178_not1;
  wire f_arrdiv24_fs178_and1;
  wire f_arrdiv24_fs178_or0;
  wire f_arrdiv24_fs179_xor0;
  wire f_arrdiv24_fs179_not0;
  wire f_arrdiv24_fs179_and0;
  wire f_arrdiv24_fs179_xor1;
  wire f_arrdiv24_fs179_not1;
  wire f_arrdiv24_fs179_and1;
  wire f_arrdiv24_fs179_or0;
  wire f_arrdiv24_fs180_xor0;
  wire f_arrdiv24_fs180_not0;
  wire f_arrdiv24_fs180_and0;
  wire f_arrdiv24_fs180_xor1;
  wire f_arrdiv24_fs180_not1;
  wire f_arrdiv24_fs180_and1;
  wire f_arrdiv24_fs180_or0;
  wire f_arrdiv24_fs181_xor0;
  wire f_arrdiv24_fs181_not0;
  wire f_arrdiv24_fs181_and0;
  wire f_arrdiv24_fs181_xor1;
  wire f_arrdiv24_fs181_not1;
  wire f_arrdiv24_fs181_and1;
  wire f_arrdiv24_fs181_or0;
  wire f_arrdiv24_fs182_xor0;
  wire f_arrdiv24_fs182_not0;
  wire f_arrdiv24_fs182_and0;
  wire f_arrdiv24_fs182_xor1;
  wire f_arrdiv24_fs182_not1;
  wire f_arrdiv24_fs182_and1;
  wire f_arrdiv24_fs182_or0;
  wire f_arrdiv24_fs183_xor0;
  wire f_arrdiv24_fs183_not0;
  wire f_arrdiv24_fs183_and0;
  wire f_arrdiv24_fs183_xor1;
  wire f_arrdiv24_fs183_not1;
  wire f_arrdiv24_fs183_and1;
  wire f_arrdiv24_fs183_or0;
  wire f_arrdiv24_fs184_xor0;
  wire f_arrdiv24_fs184_not0;
  wire f_arrdiv24_fs184_and0;
  wire f_arrdiv24_fs184_xor1;
  wire f_arrdiv24_fs184_not1;
  wire f_arrdiv24_fs184_and1;
  wire f_arrdiv24_fs184_or0;
  wire f_arrdiv24_fs185_xor0;
  wire f_arrdiv24_fs185_not0;
  wire f_arrdiv24_fs185_and0;
  wire f_arrdiv24_fs185_xor1;
  wire f_arrdiv24_fs185_not1;
  wire f_arrdiv24_fs185_and1;
  wire f_arrdiv24_fs185_or0;
  wire f_arrdiv24_fs186_xor0;
  wire f_arrdiv24_fs186_not0;
  wire f_arrdiv24_fs186_and0;
  wire f_arrdiv24_fs186_xor1;
  wire f_arrdiv24_fs186_not1;
  wire f_arrdiv24_fs186_and1;
  wire f_arrdiv24_fs186_or0;
  wire f_arrdiv24_fs187_xor0;
  wire f_arrdiv24_fs187_not0;
  wire f_arrdiv24_fs187_and0;
  wire f_arrdiv24_fs187_xor1;
  wire f_arrdiv24_fs187_not1;
  wire f_arrdiv24_fs187_and1;
  wire f_arrdiv24_fs187_or0;
  wire f_arrdiv24_fs188_xor0;
  wire f_arrdiv24_fs188_not0;
  wire f_arrdiv24_fs188_and0;
  wire f_arrdiv24_fs188_xor1;
  wire f_arrdiv24_fs188_not1;
  wire f_arrdiv24_fs188_and1;
  wire f_arrdiv24_fs188_or0;
  wire f_arrdiv24_fs189_xor0;
  wire f_arrdiv24_fs189_not0;
  wire f_arrdiv24_fs189_and0;
  wire f_arrdiv24_fs189_xor1;
  wire f_arrdiv24_fs189_not1;
  wire f_arrdiv24_fs189_and1;
  wire f_arrdiv24_fs189_or0;
  wire f_arrdiv24_fs190_xor0;
  wire f_arrdiv24_fs190_not0;
  wire f_arrdiv24_fs190_and0;
  wire f_arrdiv24_fs190_xor1;
  wire f_arrdiv24_fs190_not1;
  wire f_arrdiv24_fs190_and1;
  wire f_arrdiv24_fs190_or0;
  wire f_arrdiv24_fs191_xor0;
  wire f_arrdiv24_fs191_not0;
  wire f_arrdiv24_fs191_and0;
  wire f_arrdiv24_fs191_xor1;
  wire f_arrdiv24_fs191_not1;
  wire f_arrdiv24_fs191_and1;
  wire f_arrdiv24_fs191_or0;
  wire f_arrdiv24_mux2to1161_and0;
  wire f_arrdiv24_mux2to1161_not0;
  wire f_arrdiv24_mux2to1161_and1;
  wire f_arrdiv24_mux2to1161_xor0;
  wire f_arrdiv24_mux2to1162_and0;
  wire f_arrdiv24_mux2to1162_not0;
  wire f_arrdiv24_mux2to1162_and1;
  wire f_arrdiv24_mux2to1162_xor0;
  wire f_arrdiv24_mux2to1163_and0;
  wire f_arrdiv24_mux2to1163_not0;
  wire f_arrdiv24_mux2to1163_and1;
  wire f_arrdiv24_mux2to1163_xor0;
  wire f_arrdiv24_mux2to1164_and0;
  wire f_arrdiv24_mux2to1164_not0;
  wire f_arrdiv24_mux2to1164_and1;
  wire f_arrdiv24_mux2to1164_xor0;
  wire f_arrdiv24_mux2to1165_and0;
  wire f_arrdiv24_mux2to1165_not0;
  wire f_arrdiv24_mux2to1165_and1;
  wire f_arrdiv24_mux2to1165_xor0;
  wire f_arrdiv24_mux2to1166_and0;
  wire f_arrdiv24_mux2to1166_not0;
  wire f_arrdiv24_mux2to1166_and1;
  wire f_arrdiv24_mux2to1166_xor0;
  wire f_arrdiv24_mux2to1167_and0;
  wire f_arrdiv24_mux2to1167_not0;
  wire f_arrdiv24_mux2to1167_and1;
  wire f_arrdiv24_mux2to1167_xor0;
  wire f_arrdiv24_mux2to1168_and0;
  wire f_arrdiv24_mux2to1168_not0;
  wire f_arrdiv24_mux2to1168_and1;
  wire f_arrdiv24_mux2to1168_xor0;
  wire f_arrdiv24_mux2to1169_and0;
  wire f_arrdiv24_mux2to1169_not0;
  wire f_arrdiv24_mux2to1169_and1;
  wire f_arrdiv24_mux2to1169_xor0;
  wire f_arrdiv24_mux2to1170_and0;
  wire f_arrdiv24_mux2to1170_not0;
  wire f_arrdiv24_mux2to1170_and1;
  wire f_arrdiv24_mux2to1170_xor0;
  wire f_arrdiv24_mux2to1171_and0;
  wire f_arrdiv24_mux2to1171_not0;
  wire f_arrdiv24_mux2to1171_and1;
  wire f_arrdiv24_mux2to1171_xor0;
  wire f_arrdiv24_mux2to1172_and0;
  wire f_arrdiv24_mux2to1172_not0;
  wire f_arrdiv24_mux2to1172_and1;
  wire f_arrdiv24_mux2to1172_xor0;
  wire f_arrdiv24_mux2to1173_and0;
  wire f_arrdiv24_mux2to1173_not0;
  wire f_arrdiv24_mux2to1173_and1;
  wire f_arrdiv24_mux2to1173_xor0;
  wire f_arrdiv24_mux2to1174_and0;
  wire f_arrdiv24_mux2to1174_not0;
  wire f_arrdiv24_mux2to1174_and1;
  wire f_arrdiv24_mux2to1174_xor0;
  wire f_arrdiv24_mux2to1175_and0;
  wire f_arrdiv24_mux2to1175_not0;
  wire f_arrdiv24_mux2to1175_and1;
  wire f_arrdiv24_mux2to1175_xor0;
  wire f_arrdiv24_mux2to1176_and0;
  wire f_arrdiv24_mux2to1176_not0;
  wire f_arrdiv24_mux2to1176_and1;
  wire f_arrdiv24_mux2to1176_xor0;
  wire f_arrdiv24_mux2to1177_and0;
  wire f_arrdiv24_mux2to1177_not0;
  wire f_arrdiv24_mux2to1177_and1;
  wire f_arrdiv24_mux2to1177_xor0;
  wire f_arrdiv24_mux2to1178_and0;
  wire f_arrdiv24_mux2to1178_not0;
  wire f_arrdiv24_mux2to1178_and1;
  wire f_arrdiv24_mux2to1178_xor0;
  wire f_arrdiv24_mux2to1179_and0;
  wire f_arrdiv24_mux2to1179_not0;
  wire f_arrdiv24_mux2to1179_and1;
  wire f_arrdiv24_mux2to1179_xor0;
  wire f_arrdiv24_mux2to1180_and0;
  wire f_arrdiv24_mux2to1180_not0;
  wire f_arrdiv24_mux2to1180_and1;
  wire f_arrdiv24_mux2to1180_xor0;
  wire f_arrdiv24_mux2to1181_and0;
  wire f_arrdiv24_mux2to1181_not0;
  wire f_arrdiv24_mux2to1181_and1;
  wire f_arrdiv24_mux2to1181_xor0;
  wire f_arrdiv24_mux2to1182_and0;
  wire f_arrdiv24_mux2to1182_not0;
  wire f_arrdiv24_mux2to1182_and1;
  wire f_arrdiv24_mux2to1182_xor0;
  wire f_arrdiv24_mux2to1183_and0;
  wire f_arrdiv24_mux2to1183_not0;
  wire f_arrdiv24_mux2to1183_and1;
  wire f_arrdiv24_mux2to1183_xor0;
  wire f_arrdiv24_not7;
  wire f_arrdiv24_fs192_xor0;
  wire f_arrdiv24_fs192_not0;
  wire f_arrdiv24_fs192_and0;
  wire f_arrdiv24_fs192_not1;
  wire f_arrdiv24_fs193_xor0;
  wire f_arrdiv24_fs193_not0;
  wire f_arrdiv24_fs193_and0;
  wire f_arrdiv24_fs193_xor1;
  wire f_arrdiv24_fs193_not1;
  wire f_arrdiv24_fs193_and1;
  wire f_arrdiv24_fs193_or0;
  wire f_arrdiv24_fs194_xor0;
  wire f_arrdiv24_fs194_not0;
  wire f_arrdiv24_fs194_and0;
  wire f_arrdiv24_fs194_xor1;
  wire f_arrdiv24_fs194_not1;
  wire f_arrdiv24_fs194_and1;
  wire f_arrdiv24_fs194_or0;
  wire f_arrdiv24_fs195_xor0;
  wire f_arrdiv24_fs195_not0;
  wire f_arrdiv24_fs195_and0;
  wire f_arrdiv24_fs195_xor1;
  wire f_arrdiv24_fs195_not1;
  wire f_arrdiv24_fs195_and1;
  wire f_arrdiv24_fs195_or0;
  wire f_arrdiv24_fs196_xor0;
  wire f_arrdiv24_fs196_not0;
  wire f_arrdiv24_fs196_and0;
  wire f_arrdiv24_fs196_xor1;
  wire f_arrdiv24_fs196_not1;
  wire f_arrdiv24_fs196_and1;
  wire f_arrdiv24_fs196_or0;
  wire f_arrdiv24_fs197_xor0;
  wire f_arrdiv24_fs197_not0;
  wire f_arrdiv24_fs197_and0;
  wire f_arrdiv24_fs197_xor1;
  wire f_arrdiv24_fs197_not1;
  wire f_arrdiv24_fs197_and1;
  wire f_arrdiv24_fs197_or0;
  wire f_arrdiv24_fs198_xor0;
  wire f_arrdiv24_fs198_not0;
  wire f_arrdiv24_fs198_and0;
  wire f_arrdiv24_fs198_xor1;
  wire f_arrdiv24_fs198_not1;
  wire f_arrdiv24_fs198_and1;
  wire f_arrdiv24_fs198_or0;
  wire f_arrdiv24_fs199_xor0;
  wire f_arrdiv24_fs199_not0;
  wire f_arrdiv24_fs199_and0;
  wire f_arrdiv24_fs199_xor1;
  wire f_arrdiv24_fs199_not1;
  wire f_arrdiv24_fs199_and1;
  wire f_arrdiv24_fs199_or0;
  wire f_arrdiv24_fs200_xor0;
  wire f_arrdiv24_fs200_not0;
  wire f_arrdiv24_fs200_and0;
  wire f_arrdiv24_fs200_xor1;
  wire f_arrdiv24_fs200_not1;
  wire f_arrdiv24_fs200_and1;
  wire f_arrdiv24_fs200_or0;
  wire f_arrdiv24_fs201_xor0;
  wire f_arrdiv24_fs201_not0;
  wire f_arrdiv24_fs201_and0;
  wire f_arrdiv24_fs201_xor1;
  wire f_arrdiv24_fs201_not1;
  wire f_arrdiv24_fs201_and1;
  wire f_arrdiv24_fs201_or0;
  wire f_arrdiv24_fs202_xor0;
  wire f_arrdiv24_fs202_not0;
  wire f_arrdiv24_fs202_and0;
  wire f_arrdiv24_fs202_xor1;
  wire f_arrdiv24_fs202_not1;
  wire f_arrdiv24_fs202_and1;
  wire f_arrdiv24_fs202_or0;
  wire f_arrdiv24_fs203_xor0;
  wire f_arrdiv24_fs203_not0;
  wire f_arrdiv24_fs203_and0;
  wire f_arrdiv24_fs203_xor1;
  wire f_arrdiv24_fs203_not1;
  wire f_arrdiv24_fs203_and1;
  wire f_arrdiv24_fs203_or0;
  wire f_arrdiv24_fs204_xor0;
  wire f_arrdiv24_fs204_not0;
  wire f_arrdiv24_fs204_and0;
  wire f_arrdiv24_fs204_xor1;
  wire f_arrdiv24_fs204_not1;
  wire f_arrdiv24_fs204_and1;
  wire f_arrdiv24_fs204_or0;
  wire f_arrdiv24_fs205_xor0;
  wire f_arrdiv24_fs205_not0;
  wire f_arrdiv24_fs205_and0;
  wire f_arrdiv24_fs205_xor1;
  wire f_arrdiv24_fs205_not1;
  wire f_arrdiv24_fs205_and1;
  wire f_arrdiv24_fs205_or0;
  wire f_arrdiv24_fs206_xor0;
  wire f_arrdiv24_fs206_not0;
  wire f_arrdiv24_fs206_and0;
  wire f_arrdiv24_fs206_xor1;
  wire f_arrdiv24_fs206_not1;
  wire f_arrdiv24_fs206_and1;
  wire f_arrdiv24_fs206_or0;
  wire f_arrdiv24_fs207_xor0;
  wire f_arrdiv24_fs207_not0;
  wire f_arrdiv24_fs207_and0;
  wire f_arrdiv24_fs207_xor1;
  wire f_arrdiv24_fs207_not1;
  wire f_arrdiv24_fs207_and1;
  wire f_arrdiv24_fs207_or0;
  wire f_arrdiv24_fs208_xor0;
  wire f_arrdiv24_fs208_not0;
  wire f_arrdiv24_fs208_and0;
  wire f_arrdiv24_fs208_xor1;
  wire f_arrdiv24_fs208_not1;
  wire f_arrdiv24_fs208_and1;
  wire f_arrdiv24_fs208_or0;
  wire f_arrdiv24_fs209_xor0;
  wire f_arrdiv24_fs209_not0;
  wire f_arrdiv24_fs209_and0;
  wire f_arrdiv24_fs209_xor1;
  wire f_arrdiv24_fs209_not1;
  wire f_arrdiv24_fs209_and1;
  wire f_arrdiv24_fs209_or0;
  wire f_arrdiv24_fs210_xor0;
  wire f_arrdiv24_fs210_not0;
  wire f_arrdiv24_fs210_and0;
  wire f_arrdiv24_fs210_xor1;
  wire f_arrdiv24_fs210_not1;
  wire f_arrdiv24_fs210_and1;
  wire f_arrdiv24_fs210_or0;
  wire f_arrdiv24_fs211_xor0;
  wire f_arrdiv24_fs211_not0;
  wire f_arrdiv24_fs211_and0;
  wire f_arrdiv24_fs211_xor1;
  wire f_arrdiv24_fs211_not1;
  wire f_arrdiv24_fs211_and1;
  wire f_arrdiv24_fs211_or0;
  wire f_arrdiv24_fs212_xor0;
  wire f_arrdiv24_fs212_not0;
  wire f_arrdiv24_fs212_and0;
  wire f_arrdiv24_fs212_xor1;
  wire f_arrdiv24_fs212_not1;
  wire f_arrdiv24_fs212_and1;
  wire f_arrdiv24_fs212_or0;
  wire f_arrdiv24_fs213_xor0;
  wire f_arrdiv24_fs213_not0;
  wire f_arrdiv24_fs213_and0;
  wire f_arrdiv24_fs213_xor1;
  wire f_arrdiv24_fs213_not1;
  wire f_arrdiv24_fs213_and1;
  wire f_arrdiv24_fs213_or0;
  wire f_arrdiv24_fs214_xor0;
  wire f_arrdiv24_fs214_not0;
  wire f_arrdiv24_fs214_and0;
  wire f_arrdiv24_fs214_xor1;
  wire f_arrdiv24_fs214_not1;
  wire f_arrdiv24_fs214_and1;
  wire f_arrdiv24_fs214_or0;
  wire f_arrdiv24_fs215_xor0;
  wire f_arrdiv24_fs215_not0;
  wire f_arrdiv24_fs215_and0;
  wire f_arrdiv24_fs215_xor1;
  wire f_arrdiv24_fs215_not1;
  wire f_arrdiv24_fs215_and1;
  wire f_arrdiv24_fs215_or0;
  wire f_arrdiv24_mux2to1184_and0;
  wire f_arrdiv24_mux2to1184_not0;
  wire f_arrdiv24_mux2to1184_and1;
  wire f_arrdiv24_mux2to1184_xor0;
  wire f_arrdiv24_mux2to1185_and0;
  wire f_arrdiv24_mux2to1185_not0;
  wire f_arrdiv24_mux2to1185_and1;
  wire f_arrdiv24_mux2to1185_xor0;
  wire f_arrdiv24_mux2to1186_and0;
  wire f_arrdiv24_mux2to1186_not0;
  wire f_arrdiv24_mux2to1186_and1;
  wire f_arrdiv24_mux2to1186_xor0;
  wire f_arrdiv24_mux2to1187_and0;
  wire f_arrdiv24_mux2to1187_not0;
  wire f_arrdiv24_mux2to1187_and1;
  wire f_arrdiv24_mux2to1187_xor0;
  wire f_arrdiv24_mux2to1188_and0;
  wire f_arrdiv24_mux2to1188_not0;
  wire f_arrdiv24_mux2to1188_and1;
  wire f_arrdiv24_mux2to1188_xor0;
  wire f_arrdiv24_mux2to1189_and0;
  wire f_arrdiv24_mux2to1189_not0;
  wire f_arrdiv24_mux2to1189_and1;
  wire f_arrdiv24_mux2to1189_xor0;
  wire f_arrdiv24_mux2to1190_and0;
  wire f_arrdiv24_mux2to1190_not0;
  wire f_arrdiv24_mux2to1190_and1;
  wire f_arrdiv24_mux2to1190_xor0;
  wire f_arrdiv24_mux2to1191_and0;
  wire f_arrdiv24_mux2to1191_not0;
  wire f_arrdiv24_mux2to1191_and1;
  wire f_arrdiv24_mux2to1191_xor0;
  wire f_arrdiv24_mux2to1192_and0;
  wire f_arrdiv24_mux2to1192_not0;
  wire f_arrdiv24_mux2to1192_and1;
  wire f_arrdiv24_mux2to1192_xor0;
  wire f_arrdiv24_mux2to1193_and0;
  wire f_arrdiv24_mux2to1193_not0;
  wire f_arrdiv24_mux2to1193_and1;
  wire f_arrdiv24_mux2to1193_xor0;
  wire f_arrdiv24_mux2to1194_and0;
  wire f_arrdiv24_mux2to1194_not0;
  wire f_arrdiv24_mux2to1194_and1;
  wire f_arrdiv24_mux2to1194_xor0;
  wire f_arrdiv24_mux2to1195_and0;
  wire f_arrdiv24_mux2to1195_not0;
  wire f_arrdiv24_mux2to1195_and1;
  wire f_arrdiv24_mux2to1195_xor0;
  wire f_arrdiv24_mux2to1196_and0;
  wire f_arrdiv24_mux2to1196_not0;
  wire f_arrdiv24_mux2to1196_and1;
  wire f_arrdiv24_mux2to1196_xor0;
  wire f_arrdiv24_mux2to1197_and0;
  wire f_arrdiv24_mux2to1197_not0;
  wire f_arrdiv24_mux2to1197_and1;
  wire f_arrdiv24_mux2to1197_xor0;
  wire f_arrdiv24_mux2to1198_and0;
  wire f_arrdiv24_mux2to1198_not0;
  wire f_arrdiv24_mux2to1198_and1;
  wire f_arrdiv24_mux2to1198_xor0;
  wire f_arrdiv24_mux2to1199_and0;
  wire f_arrdiv24_mux2to1199_not0;
  wire f_arrdiv24_mux2to1199_and1;
  wire f_arrdiv24_mux2to1199_xor0;
  wire f_arrdiv24_mux2to1200_and0;
  wire f_arrdiv24_mux2to1200_not0;
  wire f_arrdiv24_mux2to1200_and1;
  wire f_arrdiv24_mux2to1200_xor0;
  wire f_arrdiv24_mux2to1201_and0;
  wire f_arrdiv24_mux2to1201_not0;
  wire f_arrdiv24_mux2to1201_and1;
  wire f_arrdiv24_mux2to1201_xor0;
  wire f_arrdiv24_mux2to1202_and0;
  wire f_arrdiv24_mux2to1202_not0;
  wire f_arrdiv24_mux2to1202_and1;
  wire f_arrdiv24_mux2to1202_xor0;
  wire f_arrdiv24_mux2to1203_and0;
  wire f_arrdiv24_mux2to1203_not0;
  wire f_arrdiv24_mux2to1203_and1;
  wire f_arrdiv24_mux2to1203_xor0;
  wire f_arrdiv24_mux2to1204_and0;
  wire f_arrdiv24_mux2to1204_not0;
  wire f_arrdiv24_mux2to1204_and1;
  wire f_arrdiv24_mux2to1204_xor0;
  wire f_arrdiv24_mux2to1205_and0;
  wire f_arrdiv24_mux2to1205_not0;
  wire f_arrdiv24_mux2to1205_and1;
  wire f_arrdiv24_mux2to1205_xor0;
  wire f_arrdiv24_mux2to1206_and0;
  wire f_arrdiv24_mux2to1206_not0;
  wire f_arrdiv24_mux2to1206_and1;
  wire f_arrdiv24_mux2to1206_xor0;
  wire f_arrdiv24_not8;
  wire f_arrdiv24_fs216_xor0;
  wire f_arrdiv24_fs216_not0;
  wire f_arrdiv24_fs216_and0;
  wire f_arrdiv24_fs216_not1;
  wire f_arrdiv24_fs217_xor0;
  wire f_arrdiv24_fs217_not0;
  wire f_arrdiv24_fs217_and0;
  wire f_arrdiv24_fs217_xor1;
  wire f_arrdiv24_fs217_not1;
  wire f_arrdiv24_fs217_and1;
  wire f_arrdiv24_fs217_or0;
  wire f_arrdiv24_fs218_xor0;
  wire f_arrdiv24_fs218_not0;
  wire f_arrdiv24_fs218_and0;
  wire f_arrdiv24_fs218_xor1;
  wire f_arrdiv24_fs218_not1;
  wire f_arrdiv24_fs218_and1;
  wire f_arrdiv24_fs218_or0;
  wire f_arrdiv24_fs219_xor0;
  wire f_arrdiv24_fs219_not0;
  wire f_arrdiv24_fs219_and0;
  wire f_arrdiv24_fs219_xor1;
  wire f_arrdiv24_fs219_not1;
  wire f_arrdiv24_fs219_and1;
  wire f_arrdiv24_fs219_or0;
  wire f_arrdiv24_fs220_xor0;
  wire f_arrdiv24_fs220_not0;
  wire f_arrdiv24_fs220_and0;
  wire f_arrdiv24_fs220_xor1;
  wire f_arrdiv24_fs220_not1;
  wire f_arrdiv24_fs220_and1;
  wire f_arrdiv24_fs220_or0;
  wire f_arrdiv24_fs221_xor0;
  wire f_arrdiv24_fs221_not0;
  wire f_arrdiv24_fs221_and0;
  wire f_arrdiv24_fs221_xor1;
  wire f_arrdiv24_fs221_not1;
  wire f_arrdiv24_fs221_and1;
  wire f_arrdiv24_fs221_or0;
  wire f_arrdiv24_fs222_xor0;
  wire f_arrdiv24_fs222_not0;
  wire f_arrdiv24_fs222_and0;
  wire f_arrdiv24_fs222_xor1;
  wire f_arrdiv24_fs222_not1;
  wire f_arrdiv24_fs222_and1;
  wire f_arrdiv24_fs222_or0;
  wire f_arrdiv24_fs223_xor0;
  wire f_arrdiv24_fs223_not0;
  wire f_arrdiv24_fs223_and0;
  wire f_arrdiv24_fs223_xor1;
  wire f_arrdiv24_fs223_not1;
  wire f_arrdiv24_fs223_and1;
  wire f_arrdiv24_fs223_or0;
  wire f_arrdiv24_fs224_xor0;
  wire f_arrdiv24_fs224_not0;
  wire f_arrdiv24_fs224_and0;
  wire f_arrdiv24_fs224_xor1;
  wire f_arrdiv24_fs224_not1;
  wire f_arrdiv24_fs224_and1;
  wire f_arrdiv24_fs224_or0;
  wire f_arrdiv24_fs225_xor0;
  wire f_arrdiv24_fs225_not0;
  wire f_arrdiv24_fs225_and0;
  wire f_arrdiv24_fs225_xor1;
  wire f_arrdiv24_fs225_not1;
  wire f_arrdiv24_fs225_and1;
  wire f_arrdiv24_fs225_or0;
  wire f_arrdiv24_fs226_xor0;
  wire f_arrdiv24_fs226_not0;
  wire f_arrdiv24_fs226_and0;
  wire f_arrdiv24_fs226_xor1;
  wire f_arrdiv24_fs226_not1;
  wire f_arrdiv24_fs226_and1;
  wire f_arrdiv24_fs226_or0;
  wire f_arrdiv24_fs227_xor0;
  wire f_arrdiv24_fs227_not0;
  wire f_arrdiv24_fs227_and0;
  wire f_arrdiv24_fs227_xor1;
  wire f_arrdiv24_fs227_not1;
  wire f_arrdiv24_fs227_and1;
  wire f_arrdiv24_fs227_or0;
  wire f_arrdiv24_fs228_xor0;
  wire f_arrdiv24_fs228_not0;
  wire f_arrdiv24_fs228_and0;
  wire f_arrdiv24_fs228_xor1;
  wire f_arrdiv24_fs228_not1;
  wire f_arrdiv24_fs228_and1;
  wire f_arrdiv24_fs228_or0;
  wire f_arrdiv24_fs229_xor0;
  wire f_arrdiv24_fs229_not0;
  wire f_arrdiv24_fs229_and0;
  wire f_arrdiv24_fs229_xor1;
  wire f_arrdiv24_fs229_not1;
  wire f_arrdiv24_fs229_and1;
  wire f_arrdiv24_fs229_or0;
  wire f_arrdiv24_fs230_xor0;
  wire f_arrdiv24_fs230_not0;
  wire f_arrdiv24_fs230_and0;
  wire f_arrdiv24_fs230_xor1;
  wire f_arrdiv24_fs230_not1;
  wire f_arrdiv24_fs230_and1;
  wire f_arrdiv24_fs230_or0;
  wire f_arrdiv24_fs231_xor0;
  wire f_arrdiv24_fs231_not0;
  wire f_arrdiv24_fs231_and0;
  wire f_arrdiv24_fs231_xor1;
  wire f_arrdiv24_fs231_not1;
  wire f_arrdiv24_fs231_and1;
  wire f_arrdiv24_fs231_or0;
  wire f_arrdiv24_fs232_xor0;
  wire f_arrdiv24_fs232_not0;
  wire f_arrdiv24_fs232_and0;
  wire f_arrdiv24_fs232_xor1;
  wire f_arrdiv24_fs232_not1;
  wire f_arrdiv24_fs232_and1;
  wire f_arrdiv24_fs232_or0;
  wire f_arrdiv24_fs233_xor0;
  wire f_arrdiv24_fs233_not0;
  wire f_arrdiv24_fs233_and0;
  wire f_arrdiv24_fs233_xor1;
  wire f_arrdiv24_fs233_not1;
  wire f_arrdiv24_fs233_and1;
  wire f_arrdiv24_fs233_or0;
  wire f_arrdiv24_fs234_xor0;
  wire f_arrdiv24_fs234_not0;
  wire f_arrdiv24_fs234_and0;
  wire f_arrdiv24_fs234_xor1;
  wire f_arrdiv24_fs234_not1;
  wire f_arrdiv24_fs234_and1;
  wire f_arrdiv24_fs234_or0;
  wire f_arrdiv24_fs235_xor0;
  wire f_arrdiv24_fs235_not0;
  wire f_arrdiv24_fs235_and0;
  wire f_arrdiv24_fs235_xor1;
  wire f_arrdiv24_fs235_not1;
  wire f_arrdiv24_fs235_and1;
  wire f_arrdiv24_fs235_or0;
  wire f_arrdiv24_fs236_xor0;
  wire f_arrdiv24_fs236_not0;
  wire f_arrdiv24_fs236_and0;
  wire f_arrdiv24_fs236_xor1;
  wire f_arrdiv24_fs236_not1;
  wire f_arrdiv24_fs236_and1;
  wire f_arrdiv24_fs236_or0;
  wire f_arrdiv24_fs237_xor0;
  wire f_arrdiv24_fs237_not0;
  wire f_arrdiv24_fs237_and0;
  wire f_arrdiv24_fs237_xor1;
  wire f_arrdiv24_fs237_not1;
  wire f_arrdiv24_fs237_and1;
  wire f_arrdiv24_fs237_or0;
  wire f_arrdiv24_fs238_xor0;
  wire f_arrdiv24_fs238_not0;
  wire f_arrdiv24_fs238_and0;
  wire f_arrdiv24_fs238_xor1;
  wire f_arrdiv24_fs238_not1;
  wire f_arrdiv24_fs238_and1;
  wire f_arrdiv24_fs238_or0;
  wire f_arrdiv24_fs239_xor0;
  wire f_arrdiv24_fs239_not0;
  wire f_arrdiv24_fs239_and0;
  wire f_arrdiv24_fs239_xor1;
  wire f_arrdiv24_fs239_not1;
  wire f_arrdiv24_fs239_and1;
  wire f_arrdiv24_fs239_or0;
  wire f_arrdiv24_mux2to1207_and0;
  wire f_arrdiv24_mux2to1207_not0;
  wire f_arrdiv24_mux2to1207_and1;
  wire f_arrdiv24_mux2to1207_xor0;
  wire f_arrdiv24_mux2to1208_and0;
  wire f_arrdiv24_mux2to1208_not0;
  wire f_arrdiv24_mux2to1208_and1;
  wire f_arrdiv24_mux2to1208_xor0;
  wire f_arrdiv24_mux2to1209_and0;
  wire f_arrdiv24_mux2to1209_not0;
  wire f_arrdiv24_mux2to1209_and1;
  wire f_arrdiv24_mux2to1209_xor0;
  wire f_arrdiv24_mux2to1210_and0;
  wire f_arrdiv24_mux2to1210_not0;
  wire f_arrdiv24_mux2to1210_and1;
  wire f_arrdiv24_mux2to1210_xor0;
  wire f_arrdiv24_mux2to1211_and0;
  wire f_arrdiv24_mux2to1211_not0;
  wire f_arrdiv24_mux2to1211_and1;
  wire f_arrdiv24_mux2to1211_xor0;
  wire f_arrdiv24_mux2to1212_and0;
  wire f_arrdiv24_mux2to1212_not0;
  wire f_arrdiv24_mux2to1212_and1;
  wire f_arrdiv24_mux2to1212_xor0;
  wire f_arrdiv24_mux2to1213_and0;
  wire f_arrdiv24_mux2to1213_not0;
  wire f_arrdiv24_mux2to1213_and1;
  wire f_arrdiv24_mux2to1213_xor0;
  wire f_arrdiv24_mux2to1214_and0;
  wire f_arrdiv24_mux2to1214_not0;
  wire f_arrdiv24_mux2to1214_and1;
  wire f_arrdiv24_mux2to1214_xor0;
  wire f_arrdiv24_mux2to1215_and0;
  wire f_arrdiv24_mux2to1215_not0;
  wire f_arrdiv24_mux2to1215_and1;
  wire f_arrdiv24_mux2to1215_xor0;
  wire f_arrdiv24_mux2to1216_and0;
  wire f_arrdiv24_mux2to1216_not0;
  wire f_arrdiv24_mux2to1216_and1;
  wire f_arrdiv24_mux2to1216_xor0;
  wire f_arrdiv24_mux2to1217_and0;
  wire f_arrdiv24_mux2to1217_not0;
  wire f_arrdiv24_mux2to1217_and1;
  wire f_arrdiv24_mux2to1217_xor0;
  wire f_arrdiv24_mux2to1218_and0;
  wire f_arrdiv24_mux2to1218_not0;
  wire f_arrdiv24_mux2to1218_and1;
  wire f_arrdiv24_mux2to1218_xor0;
  wire f_arrdiv24_mux2to1219_and0;
  wire f_arrdiv24_mux2to1219_not0;
  wire f_arrdiv24_mux2to1219_and1;
  wire f_arrdiv24_mux2to1219_xor0;
  wire f_arrdiv24_mux2to1220_and0;
  wire f_arrdiv24_mux2to1220_not0;
  wire f_arrdiv24_mux2to1220_and1;
  wire f_arrdiv24_mux2to1220_xor0;
  wire f_arrdiv24_mux2to1221_and0;
  wire f_arrdiv24_mux2to1221_not0;
  wire f_arrdiv24_mux2to1221_and1;
  wire f_arrdiv24_mux2to1221_xor0;
  wire f_arrdiv24_mux2to1222_and0;
  wire f_arrdiv24_mux2to1222_not0;
  wire f_arrdiv24_mux2to1222_and1;
  wire f_arrdiv24_mux2to1222_xor0;
  wire f_arrdiv24_mux2to1223_and0;
  wire f_arrdiv24_mux2to1223_not0;
  wire f_arrdiv24_mux2to1223_and1;
  wire f_arrdiv24_mux2to1223_xor0;
  wire f_arrdiv24_mux2to1224_and0;
  wire f_arrdiv24_mux2to1224_not0;
  wire f_arrdiv24_mux2to1224_and1;
  wire f_arrdiv24_mux2to1224_xor0;
  wire f_arrdiv24_mux2to1225_and0;
  wire f_arrdiv24_mux2to1225_not0;
  wire f_arrdiv24_mux2to1225_and1;
  wire f_arrdiv24_mux2to1225_xor0;
  wire f_arrdiv24_mux2to1226_and0;
  wire f_arrdiv24_mux2to1226_not0;
  wire f_arrdiv24_mux2to1226_and1;
  wire f_arrdiv24_mux2to1226_xor0;
  wire f_arrdiv24_mux2to1227_and0;
  wire f_arrdiv24_mux2to1227_not0;
  wire f_arrdiv24_mux2to1227_and1;
  wire f_arrdiv24_mux2to1227_xor0;
  wire f_arrdiv24_mux2to1228_and0;
  wire f_arrdiv24_mux2to1228_not0;
  wire f_arrdiv24_mux2to1228_and1;
  wire f_arrdiv24_mux2to1228_xor0;
  wire f_arrdiv24_mux2to1229_and0;
  wire f_arrdiv24_mux2to1229_not0;
  wire f_arrdiv24_mux2to1229_and1;
  wire f_arrdiv24_mux2to1229_xor0;
  wire f_arrdiv24_not9;
  wire f_arrdiv24_fs240_xor0;
  wire f_arrdiv24_fs240_not0;
  wire f_arrdiv24_fs240_and0;
  wire f_arrdiv24_fs240_not1;
  wire f_arrdiv24_fs241_xor0;
  wire f_arrdiv24_fs241_not0;
  wire f_arrdiv24_fs241_and0;
  wire f_arrdiv24_fs241_xor1;
  wire f_arrdiv24_fs241_not1;
  wire f_arrdiv24_fs241_and1;
  wire f_arrdiv24_fs241_or0;
  wire f_arrdiv24_fs242_xor0;
  wire f_arrdiv24_fs242_not0;
  wire f_arrdiv24_fs242_and0;
  wire f_arrdiv24_fs242_xor1;
  wire f_arrdiv24_fs242_not1;
  wire f_arrdiv24_fs242_and1;
  wire f_arrdiv24_fs242_or0;
  wire f_arrdiv24_fs243_xor0;
  wire f_arrdiv24_fs243_not0;
  wire f_arrdiv24_fs243_and0;
  wire f_arrdiv24_fs243_xor1;
  wire f_arrdiv24_fs243_not1;
  wire f_arrdiv24_fs243_and1;
  wire f_arrdiv24_fs243_or0;
  wire f_arrdiv24_fs244_xor0;
  wire f_arrdiv24_fs244_not0;
  wire f_arrdiv24_fs244_and0;
  wire f_arrdiv24_fs244_xor1;
  wire f_arrdiv24_fs244_not1;
  wire f_arrdiv24_fs244_and1;
  wire f_arrdiv24_fs244_or0;
  wire f_arrdiv24_fs245_xor0;
  wire f_arrdiv24_fs245_not0;
  wire f_arrdiv24_fs245_and0;
  wire f_arrdiv24_fs245_xor1;
  wire f_arrdiv24_fs245_not1;
  wire f_arrdiv24_fs245_and1;
  wire f_arrdiv24_fs245_or0;
  wire f_arrdiv24_fs246_xor0;
  wire f_arrdiv24_fs246_not0;
  wire f_arrdiv24_fs246_and0;
  wire f_arrdiv24_fs246_xor1;
  wire f_arrdiv24_fs246_not1;
  wire f_arrdiv24_fs246_and1;
  wire f_arrdiv24_fs246_or0;
  wire f_arrdiv24_fs247_xor0;
  wire f_arrdiv24_fs247_not0;
  wire f_arrdiv24_fs247_and0;
  wire f_arrdiv24_fs247_xor1;
  wire f_arrdiv24_fs247_not1;
  wire f_arrdiv24_fs247_and1;
  wire f_arrdiv24_fs247_or0;
  wire f_arrdiv24_fs248_xor0;
  wire f_arrdiv24_fs248_not0;
  wire f_arrdiv24_fs248_and0;
  wire f_arrdiv24_fs248_xor1;
  wire f_arrdiv24_fs248_not1;
  wire f_arrdiv24_fs248_and1;
  wire f_arrdiv24_fs248_or0;
  wire f_arrdiv24_fs249_xor0;
  wire f_arrdiv24_fs249_not0;
  wire f_arrdiv24_fs249_and0;
  wire f_arrdiv24_fs249_xor1;
  wire f_arrdiv24_fs249_not1;
  wire f_arrdiv24_fs249_and1;
  wire f_arrdiv24_fs249_or0;
  wire f_arrdiv24_fs250_xor0;
  wire f_arrdiv24_fs250_not0;
  wire f_arrdiv24_fs250_and0;
  wire f_arrdiv24_fs250_xor1;
  wire f_arrdiv24_fs250_not1;
  wire f_arrdiv24_fs250_and1;
  wire f_arrdiv24_fs250_or0;
  wire f_arrdiv24_fs251_xor0;
  wire f_arrdiv24_fs251_not0;
  wire f_arrdiv24_fs251_and0;
  wire f_arrdiv24_fs251_xor1;
  wire f_arrdiv24_fs251_not1;
  wire f_arrdiv24_fs251_and1;
  wire f_arrdiv24_fs251_or0;
  wire f_arrdiv24_fs252_xor0;
  wire f_arrdiv24_fs252_not0;
  wire f_arrdiv24_fs252_and0;
  wire f_arrdiv24_fs252_xor1;
  wire f_arrdiv24_fs252_not1;
  wire f_arrdiv24_fs252_and1;
  wire f_arrdiv24_fs252_or0;
  wire f_arrdiv24_fs253_xor0;
  wire f_arrdiv24_fs253_not0;
  wire f_arrdiv24_fs253_and0;
  wire f_arrdiv24_fs253_xor1;
  wire f_arrdiv24_fs253_not1;
  wire f_arrdiv24_fs253_and1;
  wire f_arrdiv24_fs253_or0;
  wire f_arrdiv24_fs254_xor0;
  wire f_arrdiv24_fs254_not0;
  wire f_arrdiv24_fs254_and0;
  wire f_arrdiv24_fs254_xor1;
  wire f_arrdiv24_fs254_not1;
  wire f_arrdiv24_fs254_and1;
  wire f_arrdiv24_fs254_or0;
  wire f_arrdiv24_fs255_xor0;
  wire f_arrdiv24_fs255_not0;
  wire f_arrdiv24_fs255_and0;
  wire f_arrdiv24_fs255_xor1;
  wire f_arrdiv24_fs255_not1;
  wire f_arrdiv24_fs255_and1;
  wire f_arrdiv24_fs255_or0;
  wire f_arrdiv24_fs256_xor0;
  wire f_arrdiv24_fs256_not0;
  wire f_arrdiv24_fs256_and0;
  wire f_arrdiv24_fs256_xor1;
  wire f_arrdiv24_fs256_not1;
  wire f_arrdiv24_fs256_and1;
  wire f_arrdiv24_fs256_or0;
  wire f_arrdiv24_fs257_xor0;
  wire f_arrdiv24_fs257_not0;
  wire f_arrdiv24_fs257_and0;
  wire f_arrdiv24_fs257_xor1;
  wire f_arrdiv24_fs257_not1;
  wire f_arrdiv24_fs257_and1;
  wire f_arrdiv24_fs257_or0;
  wire f_arrdiv24_fs258_xor0;
  wire f_arrdiv24_fs258_not0;
  wire f_arrdiv24_fs258_and0;
  wire f_arrdiv24_fs258_xor1;
  wire f_arrdiv24_fs258_not1;
  wire f_arrdiv24_fs258_and1;
  wire f_arrdiv24_fs258_or0;
  wire f_arrdiv24_fs259_xor0;
  wire f_arrdiv24_fs259_not0;
  wire f_arrdiv24_fs259_and0;
  wire f_arrdiv24_fs259_xor1;
  wire f_arrdiv24_fs259_not1;
  wire f_arrdiv24_fs259_and1;
  wire f_arrdiv24_fs259_or0;
  wire f_arrdiv24_fs260_xor0;
  wire f_arrdiv24_fs260_not0;
  wire f_arrdiv24_fs260_and0;
  wire f_arrdiv24_fs260_xor1;
  wire f_arrdiv24_fs260_not1;
  wire f_arrdiv24_fs260_and1;
  wire f_arrdiv24_fs260_or0;
  wire f_arrdiv24_fs261_xor0;
  wire f_arrdiv24_fs261_not0;
  wire f_arrdiv24_fs261_and0;
  wire f_arrdiv24_fs261_xor1;
  wire f_arrdiv24_fs261_not1;
  wire f_arrdiv24_fs261_and1;
  wire f_arrdiv24_fs261_or0;
  wire f_arrdiv24_fs262_xor0;
  wire f_arrdiv24_fs262_not0;
  wire f_arrdiv24_fs262_and0;
  wire f_arrdiv24_fs262_xor1;
  wire f_arrdiv24_fs262_not1;
  wire f_arrdiv24_fs262_and1;
  wire f_arrdiv24_fs262_or0;
  wire f_arrdiv24_fs263_xor0;
  wire f_arrdiv24_fs263_not0;
  wire f_arrdiv24_fs263_and0;
  wire f_arrdiv24_fs263_xor1;
  wire f_arrdiv24_fs263_not1;
  wire f_arrdiv24_fs263_and1;
  wire f_arrdiv24_fs263_or0;
  wire f_arrdiv24_mux2to1230_and0;
  wire f_arrdiv24_mux2to1230_not0;
  wire f_arrdiv24_mux2to1230_and1;
  wire f_arrdiv24_mux2to1230_xor0;
  wire f_arrdiv24_mux2to1231_and0;
  wire f_arrdiv24_mux2to1231_not0;
  wire f_arrdiv24_mux2to1231_and1;
  wire f_arrdiv24_mux2to1231_xor0;
  wire f_arrdiv24_mux2to1232_and0;
  wire f_arrdiv24_mux2to1232_not0;
  wire f_arrdiv24_mux2to1232_and1;
  wire f_arrdiv24_mux2to1232_xor0;
  wire f_arrdiv24_mux2to1233_and0;
  wire f_arrdiv24_mux2to1233_not0;
  wire f_arrdiv24_mux2to1233_and1;
  wire f_arrdiv24_mux2to1233_xor0;
  wire f_arrdiv24_mux2to1234_and0;
  wire f_arrdiv24_mux2to1234_not0;
  wire f_arrdiv24_mux2to1234_and1;
  wire f_arrdiv24_mux2to1234_xor0;
  wire f_arrdiv24_mux2to1235_and0;
  wire f_arrdiv24_mux2to1235_not0;
  wire f_arrdiv24_mux2to1235_and1;
  wire f_arrdiv24_mux2to1235_xor0;
  wire f_arrdiv24_mux2to1236_and0;
  wire f_arrdiv24_mux2to1236_not0;
  wire f_arrdiv24_mux2to1236_and1;
  wire f_arrdiv24_mux2to1236_xor0;
  wire f_arrdiv24_mux2to1237_and0;
  wire f_arrdiv24_mux2to1237_not0;
  wire f_arrdiv24_mux2to1237_and1;
  wire f_arrdiv24_mux2to1237_xor0;
  wire f_arrdiv24_mux2to1238_and0;
  wire f_arrdiv24_mux2to1238_not0;
  wire f_arrdiv24_mux2to1238_and1;
  wire f_arrdiv24_mux2to1238_xor0;
  wire f_arrdiv24_mux2to1239_and0;
  wire f_arrdiv24_mux2to1239_not0;
  wire f_arrdiv24_mux2to1239_and1;
  wire f_arrdiv24_mux2to1239_xor0;
  wire f_arrdiv24_mux2to1240_and0;
  wire f_arrdiv24_mux2to1240_not0;
  wire f_arrdiv24_mux2to1240_and1;
  wire f_arrdiv24_mux2to1240_xor0;
  wire f_arrdiv24_mux2to1241_and0;
  wire f_arrdiv24_mux2to1241_not0;
  wire f_arrdiv24_mux2to1241_and1;
  wire f_arrdiv24_mux2to1241_xor0;
  wire f_arrdiv24_mux2to1242_and0;
  wire f_arrdiv24_mux2to1242_not0;
  wire f_arrdiv24_mux2to1242_and1;
  wire f_arrdiv24_mux2to1242_xor0;
  wire f_arrdiv24_mux2to1243_and0;
  wire f_arrdiv24_mux2to1243_not0;
  wire f_arrdiv24_mux2to1243_and1;
  wire f_arrdiv24_mux2to1243_xor0;
  wire f_arrdiv24_mux2to1244_and0;
  wire f_arrdiv24_mux2to1244_not0;
  wire f_arrdiv24_mux2to1244_and1;
  wire f_arrdiv24_mux2to1244_xor0;
  wire f_arrdiv24_mux2to1245_and0;
  wire f_arrdiv24_mux2to1245_not0;
  wire f_arrdiv24_mux2to1245_and1;
  wire f_arrdiv24_mux2to1245_xor0;
  wire f_arrdiv24_mux2to1246_and0;
  wire f_arrdiv24_mux2to1246_not0;
  wire f_arrdiv24_mux2to1246_and1;
  wire f_arrdiv24_mux2to1246_xor0;
  wire f_arrdiv24_mux2to1247_and0;
  wire f_arrdiv24_mux2to1247_not0;
  wire f_arrdiv24_mux2to1247_and1;
  wire f_arrdiv24_mux2to1247_xor0;
  wire f_arrdiv24_mux2to1248_and0;
  wire f_arrdiv24_mux2to1248_not0;
  wire f_arrdiv24_mux2to1248_and1;
  wire f_arrdiv24_mux2to1248_xor0;
  wire f_arrdiv24_mux2to1249_and0;
  wire f_arrdiv24_mux2to1249_not0;
  wire f_arrdiv24_mux2to1249_and1;
  wire f_arrdiv24_mux2to1249_xor0;
  wire f_arrdiv24_mux2to1250_and0;
  wire f_arrdiv24_mux2to1250_not0;
  wire f_arrdiv24_mux2to1250_and1;
  wire f_arrdiv24_mux2to1250_xor0;
  wire f_arrdiv24_mux2to1251_and0;
  wire f_arrdiv24_mux2to1251_not0;
  wire f_arrdiv24_mux2to1251_and1;
  wire f_arrdiv24_mux2to1251_xor0;
  wire f_arrdiv24_mux2to1252_and0;
  wire f_arrdiv24_mux2to1252_not0;
  wire f_arrdiv24_mux2to1252_and1;
  wire f_arrdiv24_mux2to1252_xor0;
  wire f_arrdiv24_not10;
  wire f_arrdiv24_fs264_xor0;
  wire f_arrdiv24_fs264_not0;
  wire f_arrdiv24_fs264_and0;
  wire f_arrdiv24_fs264_not1;
  wire f_arrdiv24_fs265_xor0;
  wire f_arrdiv24_fs265_not0;
  wire f_arrdiv24_fs265_and0;
  wire f_arrdiv24_fs265_xor1;
  wire f_arrdiv24_fs265_not1;
  wire f_arrdiv24_fs265_and1;
  wire f_arrdiv24_fs265_or0;
  wire f_arrdiv24_fs266_xor0;
  wire f_arrdiv24_fs266_not0;
  wire f_arrdiv24_fs266_and0;
  wire f_arrdiv24_fs266_xor1;
  wire f_arrdiv24_fs266_not1;
  wire f_arrdiv24_fs266_and1;
  wire f_arrdiv24_fs266_or0;
  wire f_arrdiv24_fs267_xor0;
  wire f_arrdiv24_fs267_not0;
  wire f_arrdiv24_fs267_and0;
  wire f_arrdiv24_fs267_xor1;
  wire f_arrdiv24_fs267_not1;
  wire f_arrdiv24_fs267_and1;
  wire f_arrdiv24_fs267_or0;
  wire f_arrdiv24_fs268_xor0;
  wire f_arrdiv24_fs268_not0;
  wire f_arrdiv24_fs268_and0;
  wire f_arrdiv24_fs268_xor1;
  wire f_arrdiv24_fs268_not1;
  wire f_arrdiv24_fs268_and1;
  wire f_arrdiv24_fs268_or0;
  wire f_arrdiv24_fs269_xor0;
  wire f_arrdiv24_fs269_not0;
  wire f_arrdiv24_fs269_and0;
  wire f_arrdiv24_fs269_xor1;
  wire f_arrdiv24_fs269_not1;
  wire f_arrdiv24_fs269_and1;
  wire f_arrdiv24_fs269_or0;
  wire f_arrdiv24_fs270_xor0;
  wire f_arrdiv24_fs270_not0;
  wire f_arrdiv24_fs270_and0;
  wire f_arrdiv24_fs270_xor1;
  wire f_arrdiv24_fs270_not1;
  wire f_arrdiv24_fs270_and1;
  wire f_arrdiv24_fs270_or0;
  wire f_arrdiv24_fs271_xor0;
  wire f_arrdiv24_fs271_not0;
  wire f_arrdiv24_fs271_and0;
  wire f_arrdiv24_fs271_xor1;
  wire f_arrdiv24_fs271_not1;
  wire f_arrdiv24_fs271_and1;
  wire f_arrdiv24_fs271_or0;
  wire f_arrdiv24_fs272_xor0;
  wire f_arrdiv24_fs272_not0;
  wire f_arrdiv24_fs272_and0;
  wire f_arrdiv24_fs272_xor1;
  wire f_arrdiv24_fs272_not1;
  wire f_arrdiv24_fs272_and1;
  wire f_arrdiv24_fs272_or0;
  wire f_arrdiv24_fs273_xor0;
  wire f_arrdiv24_fs273_not0;
  wire f_arrdiv24_fs273_and0;
  wire f_arrdiv24_fs273_xor1;
  wire f_arrdiv24_fs273_not1;
  wire f_arrdiv24_fs273_and1;
  wire f_arrdiv24_fs273_or0;
  wire f_arrdiv24_fs274_xor0;
  wire f_arrdiv24_fs274_not0;
  wire f_arrdiv24_fs274_and0;
  wire f_arrdiv24_fs274_xor1;
  wire f_arrdiv24_fs274_not1;
  wire f_arrdiv24_fs274_and1;
  wire f_arrdiv24_fs274_or0;
  wire f_arrdiv24_fs275_xor0;
  wire f_arrdiv24_fs275_not0;
  wire f_arrdiv24_fs275_and0;
  wire f_arrdiv24_fs275_xor1;
  wire f_arrdiv24_fs275_not1;
  wire f_arrdiv24_fs275_and1;
  wire f_arrdiv24_fs275_or0;
  wire f_arrdiv24_fs276_xor0;
  wire f_arrdiv24_fs276_not0;
  wire f_arrdiv24_fs276_and0;
  wire f_arrdiv24_fs276_xor1;
  wire f_arrdiv24_fs276_not1;
  wire f_arrdiv24_fs276_and1;
  wire f_arrdiv24_fs276_or0;
  wire f_arrdiv24_fs277_xor0;
  wire f_arrdiv24_fs277_not0;
  wire f_arrdiv24_fs277_and0;
  wire f_arrdiv24_fs277_xor1;
  wire f_arrdiv24_fs277_not1;
  wire f_arrdiv24_fs277_and1;
  wire f_arrdiv24_fs277_or0;
  wire f_arrdiv24_fs278_xor0;
  wire f_arrdiv24_fs278_not0;
  wire f_arrdiv24_fs278_and0;
  wire f_arrdiv24_fs278_xor1;
  wire f_arrdiv24_fs278_not1;
  wire f_arrdiv24_fs278_and1;
  wire f_arrdiv24_fs278_or0;
  wire f_arrdiv24_fs279_xor0;
  wire f_arrdiv24_fs279_not0;
  wire f_arrdiv24_fs279_and0;
  wire f_arrdiv24_fs279_xor1;
  wire f_arrdiv24_fs279_not1;
  wire f_arrdiv24_fs279_and1;
  wire f_arrdiv24_fs279_or0;
  wire f_arrdiv24_fs280_xor0;
  wire f_arrdiv24_fs280_not0;
  wire f_arrdiv24_fs280_and0;
  wire f_arrdiv24_fs280_xor1;
  wire f_arrdiv24_fs280_not1;
  wire f_arrdiv24_fs280_and1;
  wire f_arrdiv24_fs280_or0;
  wire f_arrdiv24_fs281_xor0;
  wire f_arrdiv24_fs281_not0;
  wire f_arrdiv24_fs281_and0;
  wire f_arrdiv24_fs281_xor1;
  wire f_arrdiv24_fs281_not1;
  wire f_arrdiv24_fs281_and1;
  wire f_arrdiv24_fs281_or0;
  wire f_arrdiv24_fs282_xor0;
  wire f_arrdiv24_fs282_not0;
  wire f_arrdiv24_fs282_and0;
  wire f_arrdiv24_fs282_xor1;
  wire f_arrdiv24_fs282_not1;
  wire f_arrdiv24_fs282_and1;
  wire f_arrdiv24_fs282_or0;
  wire f_arrdiv24_fs283_xor0;
  wire f_arrdiv24_fs283_not0;
  wire f_arrdiv24_fs283_and0;
  wire f_arrdiv24_fs283_xor1;
  wire f_arrdiv24_fs283_not1;
  wire f_arrdiv24_fs283_and1;
  wire f_arrdiv24_fs283_or0;
  wire f_arrdiv24_fs284_xor0;
  wire f_arrdiv24_fs284_not0;
  wire f_arrdiv24_fs284_and0;
  wire f_arrdiv24_fs284_xor1;
  wire f_arrdiv24_fs284_not1;
  wire f_arrdiv24_fs284_and1;
  wire f_arrdiv24_fs284_or0;
  wire f_arrdiv24_fs285_xor0;
  wire f_arrdiv24_fs285_not0;
  wire f_arrdiv24_fs285_and0;
  wire f_arrdiv24_fs285_xor1;
  wire f_arrdiv24_fs285_not1;
  wire f_arrdiv24_fs285_and1;
  wire f_arrdiv24_fs285_or0;
  wire f_arrdiv24_fs286_xor0;
  wire f_arrdiv24_fs286_not0;
  wire f_arrdiv24_fs286_and0;
  wire f_arrdiv24_fs286_xor1;
  wire f_arrdiv24_fs286_not1;
  wire f_arrdiv24_fs286_and1;
  wire f_arrdiv24_fs286_or0;
  wire f_arrdiv24_fs287_xor0;
  wire f_arrdiv24_fs287_not0;
  wire f_arrdiv24_fs287_and0;
  wire f_arrdiv24_fs287_xor1;
  wire f_arrdiv24_fs287_not1;
  wire f_arrdiv24_fs287_and1;
  wire f_arrdiv24_fs287_or0;
  wire f_arrdiv24_mux2to1253_and0;
  wire f_arrdiv24_mux2to1253_not0;
  wire f_arrdiv24_mux2to1253_and1;
  wire f_arrdiv24_mux2to1253_xor0;
  wire f_arrdiv24_mux2to1254_and0;
  wire f_arrdiv24_mux2to1254_not0;
  wire f_arrdiv24_mux2to1254_and1;
  wire f_arrdiv24_mux2to1254_xor0;
  wire f_arrdiv24_mux2to1255_and0;
  wire f_arrdiv24_mux2to1255_not0;
  wire f_arrdiv24_mux2to1255_and1;
  wire f_arrdiv24_mux2to1255_xor0;
  wire f_arrdiv24_mux2to1256_and0;
  wire f_arrdiv24_mux2to1256_not0;
  wire f_arrdiv24_mux2to1256_and1;
  wire f_arrdiv24_mux2to1256_xor0;
  wire f_arrdiv24_mux2to1257_and0;
  wire f_arrdiv24_mux2to1257_not0;
  wire f_arrdiv24_mux2to1257_and1;
  wire f_arrdiv24_mux2to1257_xor0;
  wire f_arrdiv24_mux2to1258_and0;
  wire f_arrdiv24_mux2to1258_not0;
  wire f_arrdiv24_mux2to1258_and1;
  wire f_arrdiv24_mux2to1258_xor0;
  wire f_arrdiv24_mux2to1259_and0;
  wire f_arrdiv24_mux2to1259_not0;
  wire f_arrdiv24_mux2to1259_and1;
  wire f_arrdiv24_mux2to1259_xor0;
  wire f_arrdiv24_mux2to1260_and0;
  wire f_arrdiv24_mux2to1260_not0;
  wire f_arrdiv24_mux2to1260_and1;
  wire f_arrdiv24_mux2to1260_xor0;
  wire f_arrdiv24_mux2to1261_and0;
  wire f_arrdiv24_mux2to1261_not0;
  wire f_arrdiv24_mux2to1261_and1;
  wire f_arrdiv24_mux2to1261_xor0;
  wire f_arrdiv24_mux2to1262_and0;
  wire f_arrdiv24_mux2to1262_not0;
  wire f_arrdiv24_mux2to1262_and1;
  wire f_arrdiv24_mux2to1262_xor0;
  wire f_arrdiv24_mux2to1263_and0;
  wire f_arrdiv24_mux2to1263_not0;
  wire f_arrdiv24_mux2to1263_and1;
  wire f_arrdiv24_mux2to1263_xor0;
  wire f_arrdiv24_mux2to1264_and0;
  wire f_arrdiv24_mux2to1264_not0;
  wire f_arrdiv24_mux2to1264_and1;
  wire f_arrdiv24_mux2to1264_xor0;
  wire f_arrdiv24_mux2to1265_and0;
  wire f_arrdiv24_mux2to1265_not0;
  wire f_arrdiv24_mux2to1265_and1;
  wire f_arrdiv24_mux2to1265_xor0;
  wire f_arrdiv24_mux2to1266_and0;
  wire f_arrdiv24_mux2to1266_not0;
  wire f_arrdiv24_mux2to1266_and1;
  wire f_arrdiv24_mux2to1266_xor0;
  wire f_arrdiv24_mux2to1267_and0;
  wire f_arrdiv24_mux2to1267_not0;
  wire f_arrdiv24_mux2to1267_and1;
  wire f_arrdiv24_mux2to1267_xor0;
  wire f_arrdiv24_mux2to1268_and0;
  wire f_arrdiv24_mux2to1268_not0;
  wire f_arrdiv24_mux2to1268_and1;
  wire f_arrdiv24_mux2to1268_xor0;
  wire f_arrdiv24_mux2to1269_and0;
  wire f_arrdiv24_mux2to1269_not0;
  wire f_arrdiv24_mux2to1269_and1;
  wire f_arrdiv24_mux2to1269_xor0;
  wire f_arrdiv24_mux2to1270_and0;
  wire f_arrdiv24_mux2to1270_not0;
  wire f_arrdiv24_mux2to1270_and1;
  wire f_arrdiv24_mux2to1270_xor0;
  wire f_arrdiv24_mux2to1271_and0;
  wire f_arrdiv24_mux2to1271_not0;
  wire f_arrdiv24_mux2to1271_and1;
  wire f_arrdiv24_mux2to1271_xor0;
  wire f_arrdiv24_mux2to1272_and0;
  wire f_arrdiv24_mux2to1272_not0;
  wire f_arrdiv24_mux2to1272_and1;
  wire f_arrdiv24_mux2to1272_xor0;
  wire f_arrdiv24_mux2to1273_and0;
  wire f_arrdiv24_mux2to1273_not0;
  wire f_arrdiv24_mux2to1273_and1;
  wire f_arrdiv24_mux2to1273_xor0;
  wire f_arrdiv24_mux2to1274_and0;
  wire f_arrdiv24_mux2to1274_not0;
  wire f_arrdiv24_mux2to1274_and1;
  wire f_arrdiv24_mux2to1274_xor0;
  wire f_arrdiv24_mux2to1275_and0;
  wire f_arrdiv24_mux2to1275_not0;
  wire f_arrdiv24_mux2to1275_and1;
  wire f_arrdiv24_mux2to1275_xor0;
  wire f_arrdiv24_not11;
  wire f_arrdiv24_fs288_xor0;
  wire f_arrdiv24_fs288_not0;
  wire f_arrdiv24_fs288_and0;
  wire f_arrdiv24_fs288_not1;
  wire f_arrdiv24_fs289_xor0;
  wire f_arrdiv24_fs289_not0;
  wire f_arrdiv24_fs289_and0;
  wire f_arrdiv24_fs289_xor1;
  wire f_arrdiv24_fs289_not1;
  wire f_arrdiv24_fs289_and1;
  wire f_arrdiv24_fs289_or0;
  wire f_arrdiv24_fs290_xor0;
  wire f_arrdiv24_fs290_not0;
  wire f_arrdiv24_fs290_and0;
  wire f_arrdiv24_fs290_xor1;
  wire f_arrdiv24_fs290_not1;
  wire f_arrdiv24_fs290_and1;
  wire f_arrdiv24_fs290_or0;
  wire f_arrdiv24_fs291_xor0;
  wire f_arrdiv24_fs291_not0;
  wire f_arrdiv24_fs291_and0;
  wire f_arrdiv24_fs291_xor1;
  wire f_arrdiv24_fs291_not1;
  wire f_arrdiv24_fs291_and1;
  wire f_arrdiv24_fs291_or0;
  wire f_arrdiv24_fs292_xor0;
  wire f_arrdiv24_fs292_not0;
  wire f_arrdiv24_fs292_and0;
  wire f_arrdiv24_fs292_xor1;
  wire f_arrdiv24_fs292_not1;
  wire f_arrdiv24_fs292_and1;
  wire f_arrdiv24_fs292_or0;
  wire f_arrdiv24_fs293_xor0;
  wire f_arrdiv24_fs293_not0;
  wire f_arrdiv24_fs293_and0;
  wire f_arrdiv24_fs293_xor1;
  wire f_arrdiv24_fs293_not1;
  wire f_arrdiv24_fs293_and1;
  wire f_arrdiv24_fs293_or0;
  wire f_arrdiv24_fs294_xor0;
  wire f_arrdiv24_fs294_not0;
  wire f_arrdiv24_fs294_and0;
  wire f_arrdiv24_fs294_xor1;
  wire f_arrdiv24_fs294_not1;
  wire f_arrdiv24_fs294_and1;
  wire f_arrdiv24_fs294_or0;
  wire f_arrdiv24_fs295_xor0;
  wire f_arrdiv24_fs295_not0;
  wire f_arrdiv24_fs295_and0;
  wire f_arrdiv24_fs295_xor1;
  wire f_arrdiv24_fs295_not1;
  wire f_arrdiv24_fs295_and1;
  wire f_arrdiv24_fs295_or0;
  wire f_arrdiv24_fs296_xor0;
  wire f_arrdiv24_fs296_not0;
  wire f_arrdiv24_fs296_and0;
  wire f_arrdiv24_fs296_xor1;
  wire f_arrdiv24_fs296_not1;
  wire f_arrdiv24_fs296_and1;
  wire f_arrdiv24_fs296_or0;
  wire f_arrdiv24_fs297_xor0;
  wire f_arrdiv24_fs297_not0;
  wire f_arrdiv24_fs297_and0;
  wire f_arrdiv24_fs297_xor1;
  wire f_arrdiv24_fs297_not1;
  wire f_arrdiv24_fs297_and1;
  wire f_arrdiv24_fs297_or0;
  wire f_arrdiv24_fs298_xor0;
  wire f_arrdiv24_fs298_not0;
  wire f_arrdiv24_fs298_and0;
  wire f_arrdiv24_fs298_xor1;
  wire f_arrdiv24_fs298_not1;
  wire f_arrdiv24_fs298_and1;
  wire f_arrdiv24_fs298_or0;
  wire f_arrdiv24_fs299_xor0;
  wire f_arrdiv24_fs299_not0;
  wire f_arrdiv24_fs299_and0;
  wire f_arrdiv24_fs299_xor1;
  wire f_arrdiv24_fs299_not1;
  wire f_arrdiv24_fs299_and1;
  wire f_arrdiv24_fs299_or0;
  wire f_arrdiv24_fs300_xor0;
  wire f_arrdiv24_fs300_not0;
  wire f_arrdiv24_fs300_and0;
  wire f_arrdiv24_fs300_xor1;
  wire f_arrdiv24_fs300_not1;
  wire f_arrdiv24_fs300_and1;
  wire f_arrdiv24_fs300_or0;
  wire f_arrdiv24_fs301_xor0;
  wire f_arrdiv24_fs301_not0;
  wire f_arrdiv24_fs301_and0;
  wire f_arrdiv24_fs301_xor1;
  wire f_arrdiv24_fs301_not1;
  wire f_arrdiv24_fs301_and1;
  wire f_arrdiv24_fs301_or0;
  wire f_arrdiv24_fs302_xor0;
  wire f_arrdiv24_fs302_not0;
  wire f_arrdiv24_fs302_and0;
  wire f_arrdiv24_fs302_xor1;
  wire f_arrdiv24_fs302_not1;
  wire f_arrdiv24_fs302_and1;
  wire f_arrdiv24_fs302_or0;
  wire f_arrdiv24_fs303_xor0;
  wire f_arrdiv24_fs303_not0;
  wire f_arrdiv24_fs303_and0;
  wire f_arrdiv24_fs303_xor1;
  wire f_arrdiv24_fs303_not1;
  wire f_arrdiv24_fs303_and1;
  wire f_arrdiv24_fs303_or0;
  wire f_arrdiv24_fs304_xor0;
  wire f_arrdiv24_fs304_not0;
  wire f_arrdiv24_fs304_and0;
  wire f_arrdiv24_fs304_xor1;
  wire f_arrdiv24_fs304_not1;
  wire f_arrdiv24_fs304_and1;
  wire f_arrdiv24_fs304_or0;
  wire f_arrdiv24_fs305_xor0;
  wire f_arrdiv24_fs305_not0;
  wire f_arrdiv24_fs305_and0;
  wire f_arrdiv24_fs305_xor1;
  wire f_arrdiv24_fs305_not1;
  wire f_arrdiv24_fs305_and1;
  wire f_arrdiv24_fs305_or0;
  wire f_arrdiv24_fs306_xor0;
  wire f_arrdiv24_fs306_not0;
  wire f_arrdiv24_fs306_and0;
  wire f_arrdiv24_fs306_xor1;
  wire f_arrdiv24_fs306_not1;
  wire f_arrdiv24_fs306_and1;
  wire f_arrdiv24_fs306_or0;
  wire f_arrdiv24_fs307_xor0;
  wire f_arrdiv24_fs307_not0;
  wire f_arrdiv24_fs307_and0;
  wire f_arrdiv24_fs307_xor1;
  wire f_arrdiv24_fs307_not1;
  wire f_arrdiv24_fs307_and1;
  wire f_arrdiv24_fs307_or0;
  wire f_arrdiv24_fs308_xor0;
  wire f_arrdiv24_fs308_not0;
  wire f_arrdiv24_fs308_and0;
  wire f_arrdiv24_fs308_xor1;
  wire f_arrdiv24_fs308_not1;
  wire f_arrdiv24_fs308_and1;
  wire f_arrdiv24_fs308_or0;
  wire f_arrdiv24_fs309_xor0;
  wire f_arrdiv24_fs309_not0;
  wire f_arrdiv24_fs309_and0;
  wire f_arrdiv24_fs309_xor1;
  wire f_arrdiv24_fs309_not1;
  wire f_arrdiv24_fs309_and1;
  wire f_arrdiv24_fs309_or0;
  wire f_arrdiv24_fs310_xor0;
  wire f_arrdiv24_fs310_not0;
  wire f_arrdiv24_fs310_and0;
  wire f_arrdiv24_fs310_xor1;
  wire f_arrdiv24_fs310_not1;
  wire f_arrdiv24_fs310_and1;
  wire f_arrdiv24_fs310_or0;
  wire f_arrdiv24_fs311_xor0;
  wire f_arrdiv24_fs311_not0;
  wire f_arrdiv24_fs311_and0;
  wire f_arrdiv24_fs311_xor1;
  wire f_arrdiv24_fs311_not1;
  wire f_arrdiv24_fs311_and1;
  wire f_arrdiv24_fs311_or0;
  wire f_arrdiv24_mux2to1276_and0;
  wire f_arrdiv24_mux2to1276_not0;
  wire f_arrdiv24_mux2to1276_and1;
  wire f_arrdiv24_mux2to1276_xor0;
  wire f_arrdiv24_mux2to1277_and0;
  wire f_arrdiv24_mux2to1277_not0;
  wire f_arrdiv24_mux2to1277_and1;
  wire f_arrdiv24_mux2to1277_xor0;
  wire f_arrdiv24_mux2to1278_and0;
  wire f_arrdiv24_mux2to1278_not0;
  wire f_arrdiv24_mux2to1278_and1;
  wire f_arrdiv24_mux2to1278_xor0;
  wire f_arrdiv24_mux2to1279_and0;
  wire f_arrdiv24_mux2to1279_not0;
  wire f_arrdiv24_mux2to1279_and1;
  wire f_arrdiv24_mux2to1279_xor0;
  wire f_arrdiv24_mux2to1280_and0;
  wire f_arrdiv24_mux2to1280_not0;
  wire f_arrdiv24_mux2to1280_and1;
  wire f_arrdiv24_mux2to1280_xor0;
  wire f_arrdiv24_mux2to1281_and0;
  wire f_arrdiv24_mux2to1281_not0;
  wire f_arrdiv24_mux2to1281_and1;
  wire f_arrdiv24_mux2to1281_xor0;
  wire f_arrdiv24_mux2to1282_and0;
  wire f_arrdiv24_mux2to1282_not0;
  wire f_arrdiv24_mux2to1282_and1;
  wire f_arrdiv24_mux2to1282_xor0;
  wire f_arrdiv24_mux2to1283_and0;
  wire f_arrdiv24_mux2to1283_not0;
  wire f_arrdiv24_mux2to1283_and1;
  wire f_arrdiv24_mux2to1283_xor0;
  wire f_arrdiv24_mux2to1284_and0;
  wire f_arrdiv24_mux2to1284_not0;
  wire f_arrdiv24_mux2to1284_and1;
  wire f_arrdiv24_mux2to1284_xor0;
  wire f_arrdiv24_mux2to1285_and0;
  wire f_arrdiv24_mux2to1285_not0;
  wire f_arrdiv24_mux2to1285_and1;
  wire f_arrdiv24_mux2to1285_xor0;
  wire f_arrdiv24_mux2to1286_and0;
  wire f_arrdiv24_mux2to1286_not0;
  wire f_arrdiv24_mux2to1286_and1;
  wire f_arrdiv24_mux2to1286_xor0;
  wire f_arrdiv24_mux2to1287_and0;
  wire f_arrdiv24_mux2to1287_not0;
  wire f_arrdiv24_mux2to1287_and1;
  wire f_arrdiv24_mux2to1287_xor0;
  wire f_arrdiv24_mux2to1288_and0;
  wire f_arrdiv24_mux2to1288_not0;
  wire f_arrdiv24_mux2to1288_and1;
  wire f_arrdiv24_mux2to1288_xor0;
  wire f_arrdiv24_mux2to1289_and0;
  wire f_arrdiv24_mux2to1289_not0;
  wire f_arrdiv24_mux2to1289_and1;
  wire f_arrdiv24_mux2to1289_xor0;
  wire f_arrdiv24_mux2to1290_and0;
  wire f_arrdiv24_mux2to1290_not0;
  wire f_arrdiv24_mux2to1290_and1;
  wire f_arrdiv24_mux2to1290_xor0;
  wire f_arrdiv24_mux2to1291_and0;
  wire f_arrdiv24_mux2to1291_not0;
  wire f_arrdiv24_mux2to1291_and1;
  wire f_arrdiv24_mux2to1291_xor0;
  wire f_arrdiv24_mux2to1292_and0;
  wire f_arrdiv24_mux2to1292_not0;
  wire f_arrdiv24_mux2to1292_and1;
  wire f_arrdiv24_mux2to1292_xor0;
  wire f_arrdiv24_mux2to1293_and0;
  wire f_arrdiv24_mux2to1293_not0;
  wire f_arrdiv24_mux2to1293_and1;
  wire f_arrdiv24_mux2to1293_xor0;
  wire f_arrdiv24_mux2to1294_and0;
  wire f_arrdiv24_mux2to1294_not0;
  wire f_arrdiv24_mux2to1294_and1;
  wire f_arrdiv24_mux2to1294_xor0;
  wire f_arrdiv24_mux2to1295_and0;
  wire f_arrdiv24_mux2to1295_not0;
  wire f_arrdiv24_mux2to1295_and1;
  wire f_arrdiv24_mux2to1295_xor0;
  wire f_arrdiv24_mux2to1296_and0;
  wire f_arrdiv24_mux2to1296_not0;
  wire f_arrdiv24_mux2to1296_and1;
  wire f_arrdiv24_mux2to1296_xor0;
  wire f_arrdiv24_mux2to1297_and0;
  wire f_arrdiv24_mux2to1297_not0;
  wire f_arrdiv24_mux2to1297_and1;
  wire f_arrdiv24_mux2to1297_xor0;
  wire f_arrdiv24_mux2to1298_and0;
  wire f_arrdiv24_mux2to1298_not0;
  wire f_arrdiv24_mux2to1298_and1;
  wire f_arrdiv24_mux2to1298_xor0;
  wire f_arrdiv24_not12;
  wire f_arrdiv24_fs312_xor0;
  wire f_arrdiv24_fs312_not0;
  wire f_arrdiv24_fs312_and0;
  wire f_arrdiv24_fs312_not1;
  wire f_arrdiv24_fs313_xor0;
  wire f_arrdiv24_fs313_not0;
  wire f_arrdiv24_fs313_and0;
  wire f_arrdiv24_fs313_xor1;
  wire f_arrdiv24_fs313_not1;
  wire f_arrdiv24_fs313_and1;
  wire f_arrdiv24_fs313_or0;
  wire f_arrdiv24_fs314_xor0;
  wire f_arrdiv24_fs314_not0;
  wire f_arrdiv24_fs314_and0;
  wire f_arrdiv24_fs314_xor1;
  wire f_arrdiv24_fs314_not1;
  wire f_arrdiv24_fs314_and1;
  wire f_arrdiv24_fs314_or0;
  wire f_arrdiv24_fs315_xor0;
  wire f_arrdiv24_fs315_not0;
  wire f_arrdiv24_fs315_and0;
  wire f_arrdiv24_fs315_xor1;
  wire f_arrdiv24_fs315_not1;
  wire f_arrdiv24_fs315_and1;
  wire f_arrdiv24_fs315_or0;
  wire f_arrdiv24_fs316_xor0;
  wire f_arrdiv24_fs316_not0;
  wire f_arrdiv24_fs316_and0;
  wire f_arrdiv24_fs316_xor1;
  wire f_arrdiv24_fs316_not1;
  wire f_arrdiv24_fs316_and1;
  wire f_arrdiv24_fs316_or0;
  wire f_arrdiv24_fs317_xor0;
  wire f_arrdiv24_fs317_not0;
  wire f_arrdiv24_fs317_and0;
  wire f_arrdiv24_fs317_xor1;
  wire f_arrdiv24_fs317_not1;
  wire f_arrdiv24_fs317_and1;
  wire f_arrdiv24_fs317_or0;
  wire f_arrdiv24_fs318_xor0;
  wire f_arrdiv24_fs318_not0;
  wire f_arrdiv24_fs318_and0;
  wire f_arrdiv24_fs318_xor1;
  wire f_arrdiv24_fs318_not1;
  wire f_arrdiv24_fs318_and1;
  wire f_arrdiv24_fs318_or0;
  wire f_arrdiv24_fs319_xor0;
  wire f_arrdiv24_fs319_not0;
  wire f_arrdiv24_fs319_and0;
  wire f_arrdiv24_fs319_xor1;
  wire f_arrdiv24_fs319_not1;
  wire f_arrdiv24_fs319_and1;
  wire f_arrdiv24_fs319_or0;
  wire f_arrdiv24_fs320_xor0;
  wire f_arrdiv24_fs320_not0;
  wire f_arrdiv24_fs320_and0;
  wire f_arrdiv24_fs320_xor1;
  wire f_arrdiv24_fs320_not1;
  wire f_arrdiv24_fs320_and1;
  wire f_arrdiv24_fs320_or0;
  wire f_arrdiv24_fs321_xor0;
  wire f_arrdiv24_fs321_not0;
  wire f_arrdiv24_fs321_and0;
  wire f_arrdiv24_fs321_xor1;
  wire f_arrdiv24_fs321_not1;
  wire f_arrdiv24_fs321_and1;
  wire f_arrdiv24_fs321_or0;
  wire f_arrdiv24_fs322_xor0;
  wire f_arrdiv24_fs322_not0;
  wire f_arrdiv24_fs322_and0;
  wire f_arrdiv24_fs322_xor1;
  wire f_arrdiv24_fs322_not1;
  wire f_arrdiv24_fs322_and1;
  wire f_arrdiv24_fs322_or0;
  wire f_arrdiv24_fs323_xor0;
  wire f_arrdiv24_fs323_not0;
  wire f_arrdiv24_fs323_and0;
  wire f_arrdiv24_fs323_xor1;
  wire f_arrdiv24_fs323_not1;
  wire f_arrdiv24_fs323_and1;
  wire f_arrdiv24_fs323_or0;
  wire f_arrdiv24_fs324_xor0;
  wire f_arrdiv24_fs324_not0;
  wire f_arrdiv24_fs324_and0;
  wire f_arrdiv24_fs324_xor1;
  wire f_arrdiv24_fs324_not1;
  wire f_arrdiv24_fs324_and1;
  wire f_arrdiv24_fs324_or0;
  wire f_arrdiv24_fs325_xor0;
  wire f_arrdiv24_fs325_not0;
  wire f_arrdiv24_fs325_and0;
  wire f_arrdiv24_fs325_xor1;
  wire f_arrdiv24_fs325_not1;
  wire f_arrdiv24_fs325_and1;
  wire f_arrdiv24_fs325_or0;
  wire f_arrdiv24_fs326_xor0;
  wire f_arrdiv24_fs326_not0;
  wire f_arrdiv24_fs326_and0;
  wire f_arrdiv24_fs326_xor1;
  wire f_arrdiv24_fs326_not1;
  wire f_arrdiv24_fs326_and1;
  wire f_arrdiv24_fs326_or0;
  wire f_arrdiv24_fs327_xor0;
  wire f_arrdiv24_fs327_not0;
  wire f_arrdiv24_fs327_and0;
  wire f_arrdiv24_fs327_xor1;
  wire f_arrdiv24_fs327_not1;
  wire f_arrdiv24_fs327_and1;
  wire f_arrdiv24_fs327_or0;
  wire f_arrdiv24_fs328_xor0;
  wire f_arrdiv24_fs328_not0;
  wire f_arrdiv24_fs328_and0;
  wire f_arrdiv24_fs328_xor1;
  wire f_arrdiv24_fs328_not1;
  wire f_arrdiv24_fs328_and1;
  wire f_arrdiv24_fs328_or0;
  wire f_arrdiv24_fs329_xor0;
  wire f_arrdiv24_fs329_not0;
  wire f_arrdiv24_fs329_and0;
  wire f_arrdiv24_fs329_xor1;
  wire f_arrdiv24_fs329_not1;
  wire f_arrdiv24_fs329_and1;
  wire f_arrdiv24_fs329_or0;
  wire f_arrdiv24_fs330_xor0;
  wire f_arrdiv24_fs330_not0;
  wire f_arrdiv24_fs330_and0;
  wire f_arrdiv24_fs330_xor1;
  wire f_arrdiv24_fs330_not1;
  wire f_arrdiv24_fs330_and1;
  wire f_arrdiv24_fs330_or0;
  wire f_arrdiv24_fs331_xor0;
  wire f_arrdiv24_fs331_not0;
  wire f_arrdiv24_fs331_and0;
  wire f_arrdiv24_fs331_xor1;
  wire f_arrdiv24_fs331_not1;
  wire f_arrdiv24_fs331_and1;
  wire f_arrdiv24_fs331_or0;
  wire f_arrdiv24_fs332_xor0;
  wire f_arrdiv24_fs332_not0;
  wire f_arrdiv24_fs332_and0;
  wire f_arrdiv24_fs332_xor1;
  wire f_arrdiv24_fs332_not1;
  wire f_arrdiv24_fs332_and1;
  wire f_arrdiv24_fs332_or0;
  wire f_arrdiv24_fs333_xor0;
  wire f_arrdiv24_fs333_not0;
  wire f_arrdiv24_fs333_and0;
  wire f_arrdiv24_fs333_xor1;
  wire f_arrdiv24_fs333_not1;
  wire f_arrdiv24_fs333_and1;
  wire f_arrdiv24_fs333_or0;
  wire f_arrdiv24_fs334_xor0;
  wire f_arrdiv24_fs334_not0;
  wire f_arrdiv24_fs334_and0;
  wire f_arrdiv24_fs334_xor1;
  wire f_arrdiv24_fs334_not1;
  wire f_arrdiv24_fs334_and1;
  wire f_arrdiv24_fs334_or0;
  wire f_arrdiv24_fs335_xor0;
  wire f_arrdiv24_fs335_not0;
  wire f_arrdiv24_fs335_and0;
  wire f_arrdiv24_fs335_xor1;
  wire f_arrdiv24_fs335_not1;
  wire f_arrdiv24_fs335_and1;
  wire f_arrdiv24_fs335_or0;
  wire f_arrdiv24_mux2to1299_and0;
  wire f_arrdiv24_mux2to1299_not0;
  wire f_arrdiv24_mux2to1299_and1;
  wire f_arrdiv24_mux2to1299_xor0;
  wire f_arrdiv24_mux2to1300_and0;
  wire f_arrdiv24_mux2to1300_not0;
  wire f_arrdiv24_mux2to1300_and1;
  wire f_arrdiv24_mux2to1300_xor0;
  wire f_arrdiv24_mux2to1301_and0;
  wire f_arrdiv24_mux2to1301_not0;
  wire f_arrdiv24_mux2to1301_and1;
  wire f_arrdiv24_mux2to1301_xor0;
  wire f_arrdiv24_mux2to1302_and0;
  wire f_arrdiv24_mux2to1302_not0;
  wire f_arrdiv24_mux2to1302_and1;
  wire f_arrdiv24_mux2to1302_xor0;
  wire f_arrdiv24_mux2to1303_and0;
  wire f_arrdiv24_mux2to1303_not0;
  wire f_arrdiv24_mux2to1303_and1;
  wire f_arrdiv24_mux2to1303_xor0;
  wire f_arrdiv24_mux2to1304_and0;
  wire f_arrdiv24_mux2to1304_not0;
  wire f_arrdiv24_mux2to1304_and1;
  wire f_arrdiv24_mux2to1304_xor0;
  wire f_arrdiv24_mux2to1305_and0;
  wire f_arrdiv24_mux2to1305_not0;
  wire f_arrdiv24_mux2to1305_and1;
  wire f_arrdiv24_mux2to1305_xor0;
  wire f_arrdiv24_mux2to1306_and0;
  wire f_arrdiv24_mux2to1306_not0;
  wire f_arrdiv24_mux2to1306_and1;
  wire f_arrdiv24_mux2to1306_xor0;
  wire f_arrdiv24_mux2to1307_and0;
  wire f_arrdiv24_mux2to1307_not0;
  wire f_arrdiv24_mux2to1307_and1;
  wire f_arrdiv24_mux2to1307_xor0;
  wire f_arrdiv24_mux2to1308_and0;
  wire f_arrdiv24_mux2to1308_not0;
  wire f_arrdiv24_mux2to1308_and1;
  wire f_arrdiv24_mux2to1308_xor0;
  wire f_arrdiv24_mux2to1309_and0;
  wire f_arrdiv24_mux2to1309_not0;
  wire f_arrdiv24_mux2to1309_and1;
  wire f_arrdiv24_mux2to1309_xor0;
  wire f_arrdiv24_mux2to1310_and0;
  wire f_arrdiv24_mux2to1310_not0;
  wire f_arrdiv24_mux2to1310_and1;
  wire f_arrdiv24_mux2to1310_xor0;
  wire f_arrdiv24_mux2to1311_and0;
  wire f_arrdiv24_mux2to1311_not0;
  wire f_arrdiv24_mux2to1311_and1;
  wire f_arrdiv24_mux2to1311_xor0;
  wire f_arrdiv24_mux2to1312_and0;
  wire f_arrdiv24_mux2to1312_not0;
  wire f_arrdiv24_mux2to1312_and1;
  wire f_arrdiv24_mux2to1312_xor0;
  wire f_arrdiv24_mux2to1313_and0;
  wire f_arrdiv24_mux2to1313_not0;
  wire f_arrdiv24_mux2to1313_and1;
  wire f_arrdiv24_mux2to1313_xor0;
  wire f_arrdiv24_mux2to1314_and0;
  wire f_arrdiv24_mux2to1314_not0;
  wire f_arrdiv24_mux2to1314_and1;
  wire f_arrdiv24_mux2to1314_xor0;
  wire f_arrdiv24_mux2to1315_and0;
  wire f_arrdiv24_mux2to1315_not0;
  wire f_arrdiv24_mux2to1315_and1;
  wire f_arrdiv24_mux2to1315_xor0;
  wire f_arrdiv24_mux2to1316_and0;
  wire f_arrdiv24_mux2to1316_not0;
  wire f_arrdiv24_mux2to1316_and1;
  wire f_arrdiv24_mux2to1316_xor0;
  wire f_arrdiv24_mux2to1317_and0;
  wire f_arrdiv24_mux2to1317_not0;
  wire f_arrdiv24_mux2to1317_and1;
  wire f_arrdiv24_mux2to1317_xor0;
  wire f_arrdiv24_mux2to1318_and0;
  wire f_arrdiv24_mux2to1318_not0;
  wire f_arrdiv24_mux2to1318_and1;
  wire f_arrdiv24_mux2to1318_xor0;
  wire f_arrdiv24_mux2to1319_and0;
  wire f_arrdiv24_mux2to1319_not0;
  wire f_arrdiv24_mux2to1319_and1;
  wire f_arrdiv24_mux2to1319_xor0;
  wire f_arrdiv24_mux2to1320_and0;
  wire f_arrdiv24_mux2to1320_not0;
  wire f_arrdiv24_mux2to1320_and1;
  wire f_arrdiv24_mux2to1320_xor0;
  wire f_arrdiv24_mux2to1321_and0;
  wire f_arrdiv24_mux2to1321_not0;
  wire f_arrdiv24_mux2to1321_and1;
  wire f_arrdiv24_mux2to1321_xor0;
  wire f_arrdiv24_not13;
  wire f_arrdiv24_fs336_xor0;
  wire f_arrdiv24_fs336_not0;
  wire f_arrdiv24_fs336_and0;
  wire f_arrdiv24_fs336_not1;
  wire f_arrdiv24_fs337_xor0;
  wire f_arrdiv24_fs337_not0;
  wire f_arrdiv24_fs337_and0;
  wire f_arrdiv24_fs337_xor1;
  wire f_arrdiv24_fs337_not1;
  wire f_arrdiv24_fs337_and1;
  wire f_arrdiv24_fs337_or0;
  wire f_arrdiv24_fs338_xor0;
  wire f_arrdiv24_fs338_not0;
  wire f_arrdiv24_fs338_and0;
  wire f_arrdiv24_fs338_xor1;
  wire f_arrdiv24_fs338_not1;
  wire f_arrdiv24_fs338_and1;
  wire f_arrdiv24_fs338_or0;
  wire f_arrdiv24_fs339_xor0;
  wire f_arrdiv24_fs339_not0;
  wire f_arrdiv24_fs339_and0;
  wire f_arrdiv24_fs339_xor1;
  wire f_arrdiv24_fs339_not1;
  wire f_arrdiv24_fs339_and1;
  wire f_arrdiv24_fs339_or0;
  wire f_arrdiv24_fs340_xor0;
  wire f_arrdiv24_fs340_not0;
  wire f_arrdiv24_fs340_and0;
  wire f_arrdiv24_fs340_xor1;
  wire f_arrdiv24_fs340_not1;
  wire f_arrdiv24_fs340_and1;
  wire f_arrdiv24_fs340_or0;
  wire f_arrdiv24_fs341_xor0;
  wire f_arrdiv24_fs341_not0;
  wire f_arrdiv24_fs341_and0;
  wire f_arrdiv24_fs341_xor1;
  wire f_arrdiv24_fs341_not1;
  wire f_arrdiv24_fs341_and1;
  wire f_arrdiv24_fs341_or0;
  wire f_arrdiv24_fs342_xor0;
  wire f_arrdiv24_fs342_not0;
  wire f_arrdiv24_fs342_and0;
  wire f_arrdiv24_fs342_xor1;
  wire f_arrdiv24_fs342_not1;
  wire f_arrdiv24_fs342_and1;
  wire f_arrdiv24_fs342_or0;
  wire f_arrdiv24_fs343_xor0;
  wire f_arrdiv24_fs343_not0;
  wire f_arrdiv24_fs343_and0;
  wire f_arrdiv24_fs343_xor1;
  wire f_arrdiv24_fs343_not1;
  wire f_arrdiv24_fs343_and1;
  wire f_arrdiv24_fs343_or0;
  wire f_arrdiv24_fs344_xor0;
  wire f_arrdiv24_fs344_not0;
  wire f_arrdiv24_fs344_and0;
  wire f_arrdiv24_fs344_xor1;
  wire f_arrdiv24_fs344_not1;
  wire f_arrdiv24_fs344_and1;
  wire f_arrdiv24_fs344_or0;
  wire f_arrdiv24_fs345_xor0;
  wire f_arrdiv24_fs345_not0;
  wire f_arrdiv24_fs345_and0;
  wire f_arrdiv24_fs345_xor1;
  wire f_arrdiv24_fs345_not1;
  wire f_arrdiv24_fs345_and1;
  wire f_arrdiv24_fs345_or0;
  wire f_arrdiv24_fs346_xor0;
  wire f_arrdiv24_fs346_not0;
  wire f_arrdiv24_fs346_and0;
  wire f_arrdiv24_fs346_xor1;
  wire f_arrdiv24_fs346_not1;
  wire f_arrdiv24_fs346_and1;
  wire f_arrdiv24_fs346_or0;
  wire f_arrdiv24_fs347_xor0;
  wire f_arrdiv24_fs347_not0;
  wire f_arrdiv24_fs347_and0;
  wire f_arrdiv24_fs347_xor1;
  wire f_arrdiv24_fs347_not1;
  wire f_arrdiv24_fs347_and1;
  wire f_arrdiv24_fs347_or0;
  wire f_arrdiv24_fs348_xor0;
  wire f_arrdiv24_fs348_not0;
  wire f_arrdiv24_fs348_and0;
  wire f_arrdiv24_fs348_xor1;
  wire f_arrdiv24_fs348_not1;
  wire f_arrdiv24_fs348_and1;
  wire f_arrdiv24_fs348_or0;
  wire f_arrdiv24_fs349_xor0;
  wire f_arrdiv24_fs349_not0;
  wire f_arrdiv24_fs349_and0;
  wire f_arrdiv24_fs349_xor1;
  wire f_arrdiv24_fs349_not1;
  wire f_arrdiv24_fs349_and1;
  wire f_arrdiv24_fs349_or0;
  wire f_arrdiv24_fs350_xor0;
  wire f_arrdiv24_fs350_not0;
  wire f_arrdiv24_fs350_and0;
  wire f_arrdiv24_fs350_xor1;
  wire f_arrdiv24_fs350_not1;
  wire f_arrdiv24_fs350_and1;
  wire f_arrdiv24_fs350_or0;
  wire f_arrdiv24_fs351_xor0;
  wire f_arrdiv24_fs351_not0;
  wire f_arrdiv24_fs351_and0;
  wire f_arrdiv24_fs351_xor1;
  wire f_arrdiv24_fs351_not1;
  wire f_arrdiv24_fs351_and1;
  wire f_arrdiv24_fs351_or0;
  wire f_arrdiv24_fs352_xor0;
  wire f_arrdiv24_fs352_not0;
  wire f_arrdiv24_fs352_and0;
  wire f_arrdiv24_fs352_xor1;
  wire f_arrdiv24_fs352_not1;
  wire f_arrdiv24_fs352_and1;
  wire f_arrdiv24_fs352_or0;
  wire f_arrdiv24_fs353_xor0;
  wire f_arrdiv24_fs353_not0;
  wire f_arrdiv24_fs353_and0;
  wire f_arrdiv24_fs353_xor1;
  wire f_arrdiv24_fs353_not1;
  wire f_arrdiv24_fs353_and1;
  wire f_arrdiv24_fs353_or0;
  wire f_arrdiv24_fs354_xor0;
  wire f_arrdiv24_fs354_not0;
  wire f_arrdiv24_fs354_and0;
  wire f_arrdiv24_fs354_xor1;
  wire f_arrdiv24_fs354_not1;
  wire f_arrdiv24_fs354_and1;
  wire f_arrdiv24_fs354_or0;
  wire f_arrdiv24_fs355_xor0;
  wire f_arrdiv24_fs355_not0;
  wire f_arrdiv24_fs355_and0;
  wire f_arrdiv24_fs355_xor1;
  wire f_arrdiv24_fs355_not1;
  wire f_arrdiv24_fs355_and1;
  wire f_arrdiv24_fs355_or0;
  wire f_arrdiv24_fs356_xor0;
  wire f_arrdiv24_fs356_not0;
  wire f_arrdiv24_fs356_and0;
  wire f_arrdiv24_fs356_xor1;
  wire f_arrdiv24_fs356_not1;
  wire f_arrdiv24_fs356_and1;
  wire f_arrdiv24_fs356_or0;
  wire f_arrdiv24_fs357_xor0;
  wire f_arrdiv24_fs357_not0;
  wire f_arrdiv24_fs357_and0;
  wire f_arrdiv24_fs357_xor1;
  wire f_arrdiv24_fs357_not1;
  wire f_arrdiv24_fs357_and1;
  wire f_arrdiv24_fs357_or0;
  wire f_arrdiv24_fs358_xor0;
  wire f_arrdiv24_fs358_not0;
  wire f_arrdiv24_fs358_and0;
  wire f_arrdiv24_fs358_xor1;
  wire f_arrdiv24_fs358_not1;
  wire f_arrdiv24_fs358_and1;
  wire f_arrdiv24_fs358_or0;
  wire f_arrdiv24_fs359_xor0;
  wire f_arrdiv24_fs359_not0;
  wire f_arrdiv24_fs359_and0;
  wire f_arrdiv24_fs359_xor1;
  wire f_arrdiv24_fs359_not1;
  wire f_arrdiv24_fs359_and1;
  wire f_arrdiv24_fs359_or0;
  wire f_arrdiv24_mux2to1322_and0;
  wire f_arrdiv24_mux2to1322_not0;
  wire f_arrdiv24_mux2to1322_and1;
  wire f_arrdiv24_mux2to1322_xor0;
  wire f_arrdiv24_mux2to1323_and0;
  wire f_arrdiv24_mux2to1323_not0;
  wire f_arrdiv24_mux2to1323_and1;
  wire f_arrdiv24_mux2to1323_xor0;
  wire f_arrdiv24_mux2to1324_and0;
  wire f_arrdiv24_mux2to1324_not0;
  wire f_arrdiv24_mux2to1324_and1;
  wire f_arrdiv24_mux2to1324_xor0;
  wire f_arrdiv24_mux2to1325_and0;
  wire f_arrdiv24_mux2to1325_not0;
  wire f_arrdiv24_mux2to1325_and1;
  wire f_arrdiv24_mux2to1325_xor0;
  wire f_arrdiv24_mux2to1326_and0;
  wire f_arrdiv24_mux2to1326_not0;
  wire f_arrdiv24_mux2to1326_and1;
  wire f_arrdiv24_mux2to1326_xor0;
  wire f_arrdiv24_mux2to1327_and0;
  wire f_arrdiv24_mux2to1327_not0;
  wire f_arrdiv24_mux2to1327_and1;
  wire f_arrdiv24_mux2to1327_xor0;
  wire f_arrdiv24_mux2to1328_and0;
  wire f_arrdiv24_mux2to1328_not0;
  wire f_arrdiv24_mux2to1328_and1;
  wire f_arrdiv24_mux2to1328_xor0;
  wire f_arrdiv24_mux2to1329_and0;
  wire f_arrdiv24_mux2to1329_not0;
  wire f_arrdiv24_mux2to1329_and1;
  wire f_arrdiv24_mux2to1329_xor0;
  wire f_arrdiv24_mux2to1330_and0;
  wire f_arrdiv24_mux2to1330_not0;
  wire f_arrdiv24_mux2to1330_and1;
  wire f_arrdiv24_mux2to1330_xor0;
  wire f_arrdiv24_mux2to1331_and0;
  wire f_arrdiv24_mux2to1331_not0;
  wire f_arrdiv24_mux2to1331_and1;
  wire f_arrdiv24_mux2to1331_xor0;
  wire f_arrdiv24_mux2to1332_and0;
  wire f_arrdiv24_mux2to1332_not0;
  wire f_arrdiv24_mux2to1332_and1;
  wire f_arrdiv24_mux2to1332_xor0;
  wire f_arrdiv24_mux2to1333_and0;
  wire f_arrdiv24_mux2to1333_not0;
  wire f_arrdiv24_mux2to1333_and1;
  wire f_arrdiv24_mux2to1333_xor0;
  wire f_arrdiv24_mux2to1334_and0;
  wire f_arrdiv24_mux2to1334_not0;
  wire f_arrdiv24_mux2to1334_and1;
  wire f_arrdiv24_mux2to1334_xor0;
  wire f_arrdiv24_mux2to1335_and0;
  wire f_arrdiv24_mux2to1335_not0;
  wire f_arrdiv24_mux2to1335_and1;
  wire f_arrdiv24_mux2to1335_xor0;
  wire f_arrdiv24_mux2to1336_and0;
  wire f_arrdiv24_mux2to1336_not0;
  wire f_arrdiv24_mux2to1336_and1;
  wire f_arrdiv24_mux2to1336_xor0;
  wire f_arrdiv24_mux2to1337_and0;
  wire f_arrdiv24_mux2to1337_not0;
  wire f_arrdiv24_mux2to1337_and1;
  wire f_arrdiv24_mux2to1337_xor0;
  wire f_arrdiv24_mux2to1338_and0;
  wire f_arrdiv24_mux2to1338_not0;
  wire f_arrdiv24_mux2to1338_and1;
  wire f_arrdiv24_mux2to1338_xor0;
  wire f_arrdiv24_mux2to1339_and0;
  wire f_arrdiv24_mux2to1339_not0;
  wire f_arrdiv24_mux2to1339_and1;
  wire f_arrdiv24_mux2to1339_xor0;
  wire f_arrdiv24_mux2to1340_and0;
  wire f_arrdiv24_mux2to1340_not0;
  wire f_arrdiv24_mux2to1340_and1;
  wire f_arrdiv24_mux2to1340_xor0;
  wire f_arrdiv24_mux2to1341_and0;
  wire f_arrdiv24_mux2to1341_not0;
  wire f_arrdiv24_mux2to1341_and1;
  wire f_arrdiv24_mux2to1341_xor0;
  wire f_arrdiv24_mux2to1342_and0;
  wire f_arrdiv24_mux2to1342_not0;
  wire f_arrdiv24_mux2to1342_and1;
  wire f_arrdiv24_mux2to1342_xor0;
  wire f_arrdiv24_mux2to1343_and0;
  wire f_arrdiv24_mux2to1343_not0;
  wire f_arrdiv24_mux2to1343_and1;
  wire f_arrdiv24_mux2to1343_xor0;
  wire f_arrdiv24_mux2to1344_and0;
  wire f_arrdiv24_mux2to1344_not0;
  wire f_arrdiv24_mux2to1344_and1;
  wire f_arrdiv24_mux2to1344_xor0;
  wire f_arrdiv24_not14;
  wire f_arrdiv24_fs360_xor0;
  wire f_arrdiv24_fs360_not0;
  wire f_arrdiv24_fs360_and0;
  wire f_arrdiv24_fs360_not1;
  wire f_arrdiv24_fs361_xor0;
  wire f_arrdiv24_fs361_not0;
  wire f_arrdiv24_fs361_and0;
  wire f_arrdiv24_fs361_xor1;
  wire f_arrdiv24_fs361_not1;
  wire f_arrdiv24_fs361_and1;
  wire f_arrdiv24_fs361_or0;
  wire f_arrdiv24_fs362_xor0;
  wire f_arrdiv24_fs362_not0;
  wire f_arrdiv24_fs362_and0;
  wire f_arrdiv24_fs362_xor1;
  wire f_arrdiv24_fs362_not1;
  wire f_arrdiv24_fs362_and1;
  wire f_arrdiv24_fs362_or0;
  wire f_arrdiv24_fs363_xor0;
  wire f_arrdiv24_fs363_not0;
  wire f_arrdiv24_fs363_and0;
  wire f_arrdiv24_fs363_xor1;
  wire f_arrdiv24_fs363_not1;
  wire f_arrdiv24_fs363_and1;
  wire f_arrdiv24_fs363_or0;
  wire f_arrdiv24_fs364_xor0;
  wire f_arrdiv24_fs364_not0;
  wire f_arrdiv24_fs364_and0;
  wire f_arrdiv24_fs364_xor1;
  wire f_arrdiv24_fs364_not1;
  wire f_arrdiv24_fs364_and1;
  wire f_arrdiv24_fs364_or0;
  wire f_arrdiv24_fs365_xor0;
  wire f_arrdiv24_fs365_not0;
  wire f_arrdiv24_fs365_and0;
  wire f_arrdiv24_fs365_xor1;
  wire f_arrdiv24_fs365_not1;
  wire f_arrdiv24_fs365_and1;
  wire f_arrdiv24_fs365_or0;
  wire f_arrdiv24_fs366_xor0;
  wire f_arrdiv24_fs366_not0;
  wire f_arrdiv24_fs366_and0;
  wire f_arrdiv24_fs366_xor1;
  wire f_arrdiv24_fs366_not1;
  wire f_arrdiv24_fs366_and1;
  wire f_arrdiv24_fs366_or0;
  wire f_arrdiv24_fs367_xor0;
  wire f_arrdiv24_fs367_not0;
  wire f_arrdiv24_fs367_and0;
  wire f_arrdiv24_fs367_xor1;
  wire f_arrdiv24_fs367_not1;
  wire f_arrdiv24_fs367_and1;
  wire f_arrdiv24_fs367_or0;
  wire f_arrdiv24_fs368_xor0;
  wire f_arrdiv24_fs368_not0;
  wire f_arrdiv24_fs368_and0;
  wire f_arrdiv24_fs368_xor1;
  wire f_arrdiv24_fs368_not1;
  wire f_arrdiv24_fs368_and1;
  wire f_arrdiv24_fs368_or0;
  wire f_arrdiv24_fs369_xor0;
  wire f_arrdiv24_fs369_not0;
  wire f_arrdiv24_fs369_and0;
  wire f_arrdiv24_fs369_xor1;
  wire f_arrdiv24_fs369_not1;
  wire f_arrdiv24_fs369_and1;
  wire f_arrdiv24_fs369_or0;
  wire f_arrdiv24_fs370_xor0;
  wire f_arrdiv24_fs370_not0;
  wire f_arrdiv24_fs370_and0;
  wire f_arrdiv24_fs370_xor1;
  wire f_arrdiv24_fs370_not1;
  wire f_arrdiv24_fs370_and1;
  wire f_arrdiv24_fs370_or0;
  wire f_arrdiv24_fs371_xor0;
  wire f_arrdiv24_fs371_not0;
  wire f_arrdiv24_fs371_and0;
  wire f_arrdiv24_fs371_xor1;
  wire f_arrdiv24_fs371_not1;
  wire f_arrdiv24_fs371_and1;
  wire f_arrdiv24_fs371_or0;
  wire f_arrdiv24_fs372_xor0;
  wire f_arrdiv24_fs372_not0;
  wire f_arrdiv24_fs372_and0;
  wire f_arrdiv24_fs372_xor1;
  wire f_arrdiv24_fs372_not1;
  wire f_arrdiv24_fs372_and1;
  wire f_arrdiv24_fs372_or0;
  wire f_arrdiv24_fs373_xor0;
  wire f_arrdiv24_fs373_not0;
  wire f_arrdiv24_fs373_and0;
  wire f_arrdiv24_fs373_xor1;
  wire f_arrdiv24_fs373_not1;
  wire f_arrdiv24_fs373_and1;
  wire f_arrdiv24_fs373_or0;
  wire f_arrdiv24_fs374_xor0;
  wire f_arrdiv24_fs374_not0;
  wire f_arrdiv24_fs374_and0;
  wire f_arrdiv24_fs374_xor1;
  wire f_arrdiv24_fs374_not1;
  wire f_arrdiv24_fs374_and1;
  wire f_arrdiv24_fs374_or0;
  wire f_arrdiv24_fs375_xor0;
  wire f_arrdiv24_fs375_not0;
  wire f_arrdiv24_fs375_and0;
  wire f_arrdiv24_fs375_xor1;
  wire f_arrdiv24_fs375_not1;
  wire f_arrdiv24_fs375_and1;
  wire f_arrdiv24_fs375_or0;
  wire f_arrdiv24_fs376_xor0;
  wire f_arrdiv24_fs376_not0;
  wire f_arrdiv24_fs376_and0;
  wire f_arrdiv24_fs376_xor1;
  wire f_arrdiv24_fs376_not1;
  wire f_arrdiv24_fs376_and1;
  wire f_arrdiv24_fs376_or0;
  wire f_arrdiv24_fs377_xor0;
  wire f_arrdiv24_fs377_not0;
  wire f_arrdiv24_fs377_and0;
  wire f_arrdiv24_fs377_xor1;
  wire f_arrdiv24_fs377_not1;
  wire f_arrdiv24_fs377_and1;
  wire f_arrdiv24_fs377_or0;
  wire f_arrdiv24_fs378_xor0;
  wire f_arrdiv24_fs378_not0;
  wire f_arrdiv24_fs378_and0;
  wire f_arrdiv24_fs378_xor1;
  wire f_arrdiv24_fs378_not1;
  wire f_arrdiv24_fs378_and1;
  wire f_arrdiv24_fs378_or0;
  wire f_arrdiv24_fs379_xor0;
  wire f_arrdiv24_fs379_not0;
  wire f_arrdiv24_fs379_and0;
  wire f_arrdiv24_fs379_xor1;
  wire f_arrdiv24_fs379_not1;
  wire f_arrdiv24_fs379_and1;
  wire f_arrdiv24_fs379_or0;
  wire f_arrdiv24_fs380_xor0;
  wire f_arrdiv24_fs380_not0;
  wire f_arrdiv24_fs380_and0;
  wire f_arrdiv24_fs380_xor1;
  wire f_arrdiv24_fs380_not1;
  wire f_arrdiv24_fs380_and1;
  wire f_arrdiv24_fs380_or0;
  wire f_arrdiv24_fs381_xor0;
  wire f_arrdiv24_fs381_not0;
  wire f_arrdiv24_fs381_and0;
  wire f_arrdiv24_fs381_xor1;
  wire f_arrdiv24_fs381_not1;
  wire f_arrdiv24_fs381_and1;
  wire f_arrdiv24_fs381_or0;
  wire f_arrdiv24_fs382_xor0;
  wire f_arrdiv24_fs382_not0;
  wire f_arrdiv24_fs382_and0;
  wire f_arrdiv24_fs382_xor1;
  wire f_arrdiv24_fs382_not1;
  wire f_arrdiv24_fs382_and1;
  wire f_arrdiv24_fs382_or0;
  wire f_arrdiv24_fs383_xor0;
  wire f_arrdiv24_fs383_not0;
  wire f_arrdiv24_fs383_and0;
  wire f_arrdiv24_fs383_xor1;
  wire f_arrdiv24_fs383_not1;
  wire f_arrdiv24_fs383_and1;
  wire f_arrdiv24_fs383_or0;
  wire f_arrdiv24_mux2to1345_and0;
  wire f_arrdiv24_mux2to1345_not0;
  wire f_arrdiv24_mux2to1345_and1;
  wire f_arrdiv24_mux2to1345_xor0;
  wire f_arrdiv24_mux2to1346_and0;
  wire f_arrdiv24_mux2to1346_not0;
  wire f_arrdiv24_mux2to1346_and1;
  wire f_arrdiv24_mux2to1346_xor0;
  wire f_arrdiv24_mux2to1347_and0;
  wire f_arrdiv24_mux2to1347_not0;
  wire f_arrdiv24_mux2to1347_and1;
  wire f_arrdiv24_mux2to1347_xor0;
  wire f_arrdiv24_mux2to1348_and0;
  wire f_arrdiv24_mux2to1348_not0;
  wire f_arrdiv24_mux2to1348_and1;
  wire f_arrdiv24_mux2to1348_xor0;
  wire f_arrdiv24_mux2to1349_and0;
  wire f_arrdiv24_mux2to1349_not0;
  wire f_arrdiv24_mux2to1349_and1;
  wire f_arrdiv24_mux2to1349_xor0;
  wire f_arrdiv24_mux2to1350_and0;
  wire f_arrdiv24_mux2to1350_not0;
  wire f_arrdiv24_mux2to1350_and1;
  wire f_arrdiv24_mux2to1350_xor0;
  wire f_arrdiv24_mux2to1351_and0;
  wire f_arrdiv24_mux2to1351_not0;
  wire f_arrdiv24_mux2to1351_and1;
  wire f_arrdiv24_mux2to1351_xor0;
  wire f_arrdiv24_mux2to1352_and0;
  wire f_arrdiv24_mux2to1352_not0;
  wire f_arrdiv24_mux2to1352_and1;
  wire f_arrdiv24_mux2to1352_xor0;
  wire f_arrdiv24_mux2to1353_and0;
  wire f_arrdiv24_mux2to1353_not0;
  wire f_arrdiv24_mux2to1353_and1;
  wire f_arrdiv24_mux2to1353_xor0;
  wire f_arrdiv24_mux2to1354_and0;
  wire f_arrdiv24_mux2to1354_not0;
  wire f_arrdiv24_mux2to1354_and1;
  wire f_arrdiv24_mux2to1354_xor0;
  wire f_arrdiv24_mux2to1355_and0;
  wire f_arrdiv24_mux2to1355_not0;
  wire f_arrdiv24_mux2to1355_and1;
  wire f_arrdiv24_mux2to1355_xor0;
  wire f_arrdiv24_mux2to1356_and0;
  wire f_arrdiv24_mux2to1356_not0;
  wire f_arrdiv24_mux2to1356_and1;
  wire f_arrdiv24_mux2to1356_xor0;
  wire f_arrdiv24_mux2to1357_and0;
  wire f_arrdiv24_mux2to1357_not0;
  wire f_arrdiv24_mux2to1357_and1;
  wire f_arrdiv24_mux2to1357_xor0;
  wire f_arrdiv24_mux2to1358_and0;
  wire f_arrdiv24_mux2to1358_not0;
  wire f_arrdiv24_mux2to1358_and1;
  wire f_arrdiv24_mux2to1358_xor0;
  wire f_arrdiv24_mux2to1359_and0;
  wire f_arrdiv24_mux2to1359_not0;
  wire f_arrdiv24_mux2to1359_and1;
  wire f_arrdiv24_mux2to1359_xor0;
  wire f_arrdiv24_mux2to1360_and0;
  wire f_arrdiv24_mux2to1360_not0;
  wire f_arrdiv24_mux2to1360_and1;
  wire f_arrdiv24_mux2to1360_xor0;
  wire f_arrdiv24_mux2to1361_and0;
  wire f_arrdiv24_mux2to1361_not0;
  wire f_arrdiv24_mux2to1361_and1;
  wire f_arrdiv24_mux2to1361_xor0;
  wire f_arrdiv24_mux2to1362_and0;
  wire f_arrdiv24_mux2to1362_not0;
  wire f_arrdiv24_mux2to1362_and1;
  wire f_arrdiv24_mux2to1362_xor0;
  wire f_arrdiv24_mux2to1363_and0;
  wire f_arrdiv24_mux2to1363_not0;
  wire f_arrdiv24_mux2to1363_and1;
  wire f_arrdiv24_mux2to1363_xor0;
  wire f_arrdiv24_mux2to1364_and0;
  wire f_arrdiv24_mux2to1364_not0;
  wire f_arrdiv24_mux2to1364_and1;
  wire f_arrdiv24_mux2to1364_xor0;
  wire f_arrdiv24_mux2to1365_and0;
  wire f_arrdiv24_mux2to1365_not0;
  wire f_arrdiv24_mux2to1365_and1;
  wire f_arrdiv24_mux2to1365_xor0;
  wire f_arrdiv24_mux2to1366_and0;
  wire f_arrdiv24_mux2to1366_not0;
  wire f_arrdiv24_mux2to1366_and1;
  wire f_arrdiv24_mux2to1366_xor0;
  wire f_arrdiv24_mux2to1367_and0;
  wire f_arrdiv24_mux2to1367_not0;
  wire f_arrdiv24_mux2to1367_and1;
  wire f_arrdiv24_mux2to1367_xor0;
  wire f_arrdiv24_not15;
  wire f_arrdiv24_fs384_xor0;
  wire f_arrdiv24_fs384_not0;
  wire f_arrdiv24_fs384_and0;
  wire f_arrdiv24_fs384_not1;
  wire f_arrdiv24_fs385_xor0;
  wire f_arrdiv24_fs385_not0;
  wire f_arrdiv24_fs385_and0;
  wire f_arrdiv24_fs385_xor1;
  wire f_arrdiv24_fs385_not1;
  wire f_arrdiv24_fs385_and1;
  wire f_arrdiv24_fs385_or0;
  wire f_arrdiv24_fs386_xor0;
  wire f_arrdiv24_fs386_not0;
  wire f_arrdiv24_fs386_and0;
  wire f_arrdiv24_fs386_xor1;
  wire f_arrdiv24_fs386_not1;
  wire f_arrdiv24_fs386_and1;
  wire f_arrdiv24_fs386_or0;
  wire f_arrdiv24_fs387_xor0;
  wire f_arrdiv24_fs387_not0;
  wire f_arrdiv24_fs387_and0;
  wire f_arrdiv24_fs387_xor1;
  wire f_arrdiv24_fs387_not1;
  wire f_arrdiv24_fs387_and1;
  wire f_arrdiv24_fs387_or0;
  wire f_arrdiv24_fs388_xor0;
  wire f_arrdiv24_fs388_not0;
  wire f_arrdiv24_fs388_and0;
  wire f_arrdiv24_fs388_xor1;
  wire f_arrdiv24_fs388_not1;
  wire f_arrdiv24_fs388_and1;
  wire f_arrdiv24_fs388_or0;
  wire f_arrdiv24_fs389_xor0;
  wire f_arrdiv24_fs389_not0;
  wire f_arrdiv24_fs389_and0;
  wire f_arrdiv24_fs389_xor1;
  wire f_arrdiv24_fs389_not1;
  wire f_arrdiv24_fs389_and1;
  wire f_arrdiv24_fs389_or0;
  wire f_arrdiv24_fs390_xor0;
  wire f_arrdiv24_fs390_not0;
  wire f_arrdiv24_fs390_and0;
  wire f_arrdiv24_fs390_xor1;
  wire f_arrdiv24_fs390_not1;
  wire f_arrdiv24_fs390_and1;
  wire f_arrdiv24_fs390_or0;
  wire f_arrdiv24_fs391_xor0;
  wire f_arrdiv24_fs391_not0;
  wire f_arrdiv24_fs391_and0;
  wire f_arrdiv24_fs391_xor1;
  wire f_arrdiv24_fs391_not1;
  wire f_arrdiv24_fs391_and1;
  wire f_arrdiv24_fs391_or0;
  wire f_arrdiv24_fs392_xor0;
  wire f_arrdiv24_fs392_not0;
  wire f_arrdiv24_fs392_and0;
  wire f_arrdiv24_fs392_xor1;
  wire f_arrdiv24_fs392_not1;
  wire f_arrdiv24_fs392_and1;
  wire f_arrdiv24_fs392_or0;
  wire f_arrdiv24_fs393_xor0;
  wire f_arrdiv24_fs393_not0;
  wire f_arrdiv24_fs393_and0;
  wire f_arrdiv24_fs393_xor1;
  wire f_arrdiv24_fs393_not1;
  wire f_arrdiv24_fs393_and1;
  wire f_arrdiv24_fs393_or0;
  wire f_arrdiv24_fs394_xor0;
  wire f_arrdiv24_fs394_not0;
  wire f_arrdiv24_fs394_and0;
  wire f_arrdiv24_fs394_xor1;
  wire f_arrdiv24_fs394_not1;
  wire f_arrdiv24_fs394_and1;
  wire f_arrdiv24_fs394_or0;
  wire f_arrdiv24_fs395_xor0;
  wire f_arrdiv24_fs395_not0;
  wire f_arrdiv24_fs395_and0;
  wire f_arrdiv24_fs395_xor1;
  wire f_arrdiv24_fs395_not1;
  wire f_arrdiv24_fs395_and1;
  wire f_arrdiv24_fs395_or0;
  wire f_arrdiv24_fs396_xor0;
  wire f_arrdiv24_fs396_not0;
  wire f_arrdiv24_fs396_and0;
  wire f_arrdiv24_fs396_xor1;
  wire f_arrdiv24_fs396_not1;
  wire f_arrdiv24_fs396_and1;
  wire f_arrdiv24_fs396_or0;
  wire f_arrdiv24_fs397_xor0;
  wire f_arrdiv24_fs397_not0;
  wire f_arrdiv24_fs397_and0;
  wire f_arrdiv24_fs397_xor1;
  wire f_arrdiv24_fs397_not1;
  wire f_arrdiv24_fs397_and1;
  wire f_arrdiv24_fs397_or0;
  wire f_arrdiv24_fs398_xor0;
  wire f_arrdiv24_fs398_not0;
  wire f_arrdiv24_fs398_and0;
  wire f_arrdiv24_fs398_xor1;
  wire f_arrdiv24_fs398_not1;
  wire f_arrdiv24_fs398_and1;
  wire f_arrdiv24_fs398_or0;
  wire f_arrdiv24_fs399_xor0;
  wire f_arrdiv24_fs399_not0;
  wire f_arrdiv24_fs399_and0;
  wire f_arrdiv24_fs399_xor1;
  wire f_arrdiv24_fs399_not1;
  wire f_arrdiv24_fs399_and1;
  wire f_arrdiv24_fs399_or0;
  wire f_arrdiv24_fs400_xor0;
  wire f_arrdiv24_fs400_not0;
  wire f_arrdiv24_fs400_and0;
  wire f_arrdiv24_fs400_xor1;
  wire f_arrdiv24_fs400_not1;
  wire f_arrdiv24_fs400_and1;
  wire f_arrdiv24_fs400_or0;
  wire f_arrdiv24_fs401_xor0;
  wire f_arrdiv24_fs401_not0;
  wire f_arrdiv24_fs401_and0;
  wire f_arrdiv24_fs401_xor1;
  wire f_arrdiv24_fs401_not1;
  wire f_arrdiv24_fs401_and1;
  wire f_arrdiv24_fs401_or0;
  wire f_arrdiv24_fs402_xor0;
  wire f_arrdiv24_fs402_not0;
  wire f_arrdiv24_fs402_and0;
  wire f_arrdiv24_fs402_xor1;
  wire f_arrdiv24_fs402_not1;
  wire f_arrdiv24_fs402_and1;
  wire f_arrdiv24_fs402_or0;
  wire f_arrdiv24_fs403_xor0;
  wire f_arrdiv24_fs403_not0;
  wire f_arrdiv24_fs403_and0;
  wire f_arrdiv24_fs403_xor1;
  wire f_arrdiv24_fs403_not1;
  wire f_arrdiv24_fs403_and1;
  wire f_arrdiv24_fs403_or0;
  wire f_arrdiv24_fs404_xor0;
  wire f_arrdiv24_fs404_not0;
  wire f_arrdiv24_fs404_and0;
  wire f_arrdiv24_fs404_xor1;
  wire f_arrdiv24_fs404_not1;
  wire f_arrdiv24_fs404_and1;
  wire f_arrdiv24_fs404_or0;
  wire f_arrdiv24_fs405_xor0;
  wire f_arrdiv24_fs405_not0;
  wire f_arrdiv24_fs405_and0;
  wire f_arrdiv24_fs405_xor1;
  wire f_arrdiv24_fs405_not1;
  wire f_arrdiv24_fs405_and1;
  wire f_arrdiv24_fs405_or0;
  wire f_arrdiv24_fs406_xor0;
  wire f_arrdiv24_fs406_not0;
  wire f_arrdiv24_fs406_and0;
  wire f_arrdiv24_fs406_xor1;
  wire f_arrdiv24_fs406_not1;
  wire f_arrdiv24_fs406_and1;
  wire f_arrdiv24_fs406_or0;
  wire f_arrdiv24_fs407_xor0;
  wire f_arrdiv24_fs407_not0;
  wire f_arrdiv24_fs407_and0;
  wire f_arrdiv24_fs407_xor1;
  wire f_arrdiv24_fs407_not1;
  wire f_arrdiv24_fs407_and1;
  wire f_arrdiv24_fs407_or0;
  wire f_arrdiv24_mux2to1368_and0;
  wire f_arrdiv24_mux2to1368_not0;
  wire f_arrdiv24_mux2to1368_and1;
  wire f_arrdiv24_mux2to1368_xor0;
  wire f_arrdiv24_mux2to1369_and0;
  wire f_arrdiv24_mux2to1369_not0;
  wire f_arrdiv24_mux2to1369_and1;
  wire f_arrdiv24_mux2to1369_xor0;
  wire f_arrdiv24_mux2to1370_and0;
  wire f_arrdiv24_mux2to1370_not0;
  wire f_arrdiv24_mux2to1370_and1;
  wire f_arrdiv24_mux2to1370_xor0;
  wire f_arrdiv24_mux2to1371_and0;
  wire f_arrdiv24_mux2to1371_not0;
  wire f_arrdiv24_mux2to1371_and1;
  wire f_arrdiv24_mux2to1371_xor0;
  wire f_arrdiv24_mux2to1372_and0;
  wire f_arrdiv24_mux2to1372_not0;
  wire f_arrdiv24_mux2to1372_and1;
  wire f_arrdiv24_mux2to1372_xor0;
  wire f_arrdiv24_mux2to1373_and0;
  wire f_arrdiv24_mux2to1373_not0;
  wire f_arrdiv24_mux2to1373_and1;
  wire f_arrdiv24_mux2to1373_xor0;
  wire f_arrdiv24_mux2to1374_and0;
  wire f_arrdiv24_mux2to1374_not0;
  wire f_arrdiv24_mux2to1374_and1;
  wire f_arrdiv24_mux2to1374_xor0;
  wire f_arrdiv24_mux2to1375_and0;
  wire f_arrdiv24_mux2to1375_not0;
  wire f_arrdiv24_mux2to1375_and1;
  wire f_arrdiv24_mux2to1375_xor0;
  wire f_arrdiv24_mux2to1376_and0;
  wire f_arrdiv24_mux2to1376_not0;
  wire f_arrdiv24_mux2to1376_and1;
  wire f_arrdiv24_mux2to1376_xor0;
  wire f_arrdiv24_mux2to1377_and0;
  wire f_arrdiv24_mux2to1377_not0;
  wire f_arrdiv24_mux2to1377_and1;
  wire f_arrdiv24_mux2to1377_xor0;
  wire f_arrdiv24_mux2to1378_and0;
  wire f_arrdiv24_mux2to1378_not0;
  wire f_arrdiv24_mux2to1378_and1;
  wire f_arrdiv24_mux2to1378_xor0;
  wire f_arrdiv24_mux2to1379_and0;
  wire f_arrdiv24_mux2to1379_not0;
  wire f_arrdiv24_mux2to1379_and1;
  wire f_arrdiv24_mux2to1379_xor0;
  wire f_arrdiv24_mux2to1380_and0;
  wire f_arrdiv24_mux2to1380_not0;
  wire f_arrdiv24_mux2to1380_and1;
  wire f_arrdiv24_mux2to1380_xor0;
  wire f_arrdiv24_mux2to1381_and0;
  wire f_arrdiv24_mux2to1381_not0;
  wire f_arrdiv24_mux2to1381_and1;
  wire f_arrdiv24_mux2to1381_xor0;
  wire f_arrdiv24_mux2to1382_and0;
  wire f_arrdiv24_mux2to1382_not0;
  wire f_arrdiv24_mux2to1382_and1;
  wire f_arrdiv24_mux2to1382_xor0;
  wire f_arrdiv24_mux2to1383_and0;
  wire f_arrdiv24_mux2to1383_not0;
  wire f_arrdiv24_mux2to1383_and1;
  wire f_arrdiv24_mux2to1383_xor0;
  wire f_arrdiv24_mux2to1384_and0;
  wire f_arrdiv24_mux2to1384_not0;
  wire f_arrdiv24_mux2to1384_and1;
  wire f_arrdiv24_mux2to1384_xor0;
  wire f_arrdiv24_mux2to1385_and0;
  wire f_arrdiv24_mux2to1385_not0;
  wire f_arrdiv24_mux2to1385_and1;
  wire f_arrdiv24_mux2to1385_xor0;
  wire f_arrdiv24_mux2to1386_and0;
  wire f_arrdiv24_mux2to1386_not0;
  wire f_arrdiv24_mux2to1386_and1;
  wire f_arrdiv24_mux2to1386_xor0;
  wire f_arrdiv24_mux2to1387_and0;
  wire f_arrdiv24_mux2to1387_not0;
  wire f_arrdiv24_mux2to1387_and1;
  wire f_arrdiv24_mux2to1387_xor0;
  wire f_arrdiv24_mux2to1388_and0;
  wire f_arrdiv24_mux2to1388_not0;
  wire f_arrdiv24_mux2to1388_and1;
  wire f_arrdiv24_mux2to1388_xor0;
  wire f_arrdiv24_mux2to1389_and0;
  wire f_arrdiv24_mux2to1389_not0;
  wire f_arrdiv24_mux2to1389_and1;
  wire f_arrdiv24_mux2to1389_xor0;
  wire f_arrdiv24_mux2to1390_and0;
  wire f_arrdiv24_mux2to1390_not0;
  wire f_arrdiv24_mux2to1390_and1;
  wire f_arrdiv24_mux2to1390_xor0;
  wire f_arrdiv24_not16;
  wire f_arrdiv24_fs408_xor0;
  wire f_arrdiv24_fs408_not0;
  wire f_arrdiv24_fs408_and0;
  wire f_arrdiv24_fs408_not1;
  wire f_arrdiv24_fs409_xor0;
  wire f_arrdiv24_fs409_not0;
  wire f_arrdiv24_fs409_and0;
  wire f_arrdiv24_fs409_xor1;
  wire f_arrdiv24_fs409_not1;
  wire f_arrdiv24_fs409_and1;
  wire f_arrdiv24_fs409_or0;
  wire f_arrdiv24_fs410_xor0;
  wire f_arrdiv24_fs410_not0;
  wire f_arrdiv24_fs410_and0;
  wire f_arrdiv24_fs410_xor1;
  wire f_arrdiv24_fs410_not1;
  wire f_arrdiv24_fs410_and1;
  wire f_arrdiv24_fs410_or0;
  wire f_arrdiv24_fs411_xor0;
  wire f_arrdiv24_fs411_not0;
  wire f_arrdiv24_fs411_and0;
  wire f_arrdiv24_fs411_xor1;
  wire f_arrdiv24_fs411_not1;
  wire f_arrdiv24_fs411_and1;
  wire f_arrdiv24_fs411_or0;
  wire f_arrdiv24_fs412_xor0;
  wire f_arrdiv24_fs412_not0;
  wire f_arrdiv24_fs412_and0;
  wire f_arrdiv24_fs412_xor1;
  wire f_arrdiv24_fs412_not1;
  wire f_arrdiv24_fs412_and1;
  wire f_arrdiv24_fs412_or0;
  wire f_arrdiv24_fs413_xor0;
  wire f_arrdiv24_fs413_not0;
  wire f_arrdiv24_fs413_and0;
  wire f_arrdiv24_fs413_xor1;
  wire f_arrdiv24_fs413_not1;
  wire f_arrdiv24_fs413_and1;
  wire f_arrdiv24_fs413_or0;
  wire f_arrdiv24_fs414_xor0;
  wire f_arrdiv24_fs414_not0;
  wire f_arrdiv24_fs414_and0;
  wire f_arrdiv24_fs414_xor1;
  wire f_arrdiv24_fs414_not1;
  wire f_arrdiv24_fs414_and1;
  wire f_arrdiv24_fs414_or0;
  wire f_arrdiv24_fs415_xor0;
  wire f_arrdiv24_fs415_not0;
  wire f_arrdiv24_fs415_and0;
  wire f_arrdiv24_fs415_xor1;
  wire f_arrdiv24_fs415_not1;
  wire f_arrdiv24_fs415_and1;
  wire f_arrdiv24_fs415_or0;
  wire f_arrdiv24_fs416_xor0;
  wire f_arrdiv24_fs416_not0;
  wire f_arrdiv24_fs416_and0;
  wire f_arrdiv24_fs416_xor1;
  wire f_arrdiv24_fs416_not1;
  wire f_arrdiv24_fs416_and1;
  wire f_arrdiv24_fs416_or0;
  wire f_arrdiv24_fs417_xor0;
  wire f_arrdiv24_fs417_not0;
  wire f_arrdiv24_fs417_and0;
  wire f_arrdiv24_fs417_xor1;
  wire f_arrdiv24_fs417_not1;
  wire f_arrdiv24_fs417_and1;
  wire f_arrdiv24_fs417_or0;
  wire f_arrdiv24_fs418_xor0;
  wire f_arrdiv24_fs418_not0;
  wire f_arrdiv24_fs418_and0;
  wire f_arrdiv24_fs418_xor1;
  wire f_arrdiv24_fs418_not1;
  wire f_arrdiv24_fs418_and1;
  wire f_arrdiv24_fs418_or0;
  wire f_arrdiv24_fs419_xor0;
  wire f_arrdiv24_fs419_not0;
  wire f_arrdiv24_fs419_and0;
  wire f_arrdiv24_fs419_xor1;
  wire f_arrdiv24_fs419_not1;
  wire f_arrdiv24_fs419_and1;
  wire f_arrdiv24_fs419_or0;
  wire f_arrdiv24_fs420_xor0;
  wire f_arrdiv24_fs420_not0;
  wire f_arrdiv24_fs420_and0;
  wire f_arrdiv24_fs420_xor1;
  wire f_arrdiv24_fs420_not1;
  wire f_arrdiv24_fs420_and1;
  wire f_arrdiv24_fs420_or0;
  wire f_arrdiv24_fs421_xor0;
  wire f_arrdiv24_fs421_not0;
  wire f_arrdiv24_fs421_and0;
  wire f_arrdiv24_fs421_xor1;
  wire f_arrdiv24_fs421_not1;
  wire f_arrdiv24_fs421_and1;
  wire f_arrdiv24_fs421_or0;
  wire f_arrdiv24_fs422_xor0;
  wire f_arrdiv24_fs422_not0;
  wire f_arrdiv24_fs422_and0;
  wire f_arrdiv24_fs422_xor1;
  wire f_arrdiv24_fs422_not1;
  wire f_arrdiv24_fs422_and1;
  wire f_arrdiv24_fs422_or0;
  wire f_arrdiv24_fs423_xor0;
  wire f_arrdiv24_fs423_not0;
  wire f_arrdiv24_fs423_and0;
  wire f_arrdiv24_fs423_xor1;
  wire f_arrdiv24_fs423_not1;
  wire f_arrdiv24_fs423_and1;
  wire f_arrdiv24_fs423_or0;
  wire f_arrdiv24_fs424_xor0;
  wire f_arrdiv24_fs424_not0;
  wire f_arrdiv24_fs424_and0;
  wire f_arrdiv24_fs424_xor1;
  wire f_arrdiv24_fs424_not1;
  wire f_arrdiv24_fs424_and1;
  wire f_arrdiv24_fs424_or0;
  wire f_arrdiv24_fs425_xor0;
  wire f_arrdiv24_fs425_not0;
  wire f_arrdiv24_fs425_and0;
  wire f_arrdiv24_fs425_xor1;
  wire f_arrdiv24_fs425_not1;
  wire f_arrdiv24_fs425_and1;
  wire f_arrdiv24_fs425_or0;
  wire f_arrdiv24_fs426_xor0;
  wire f_arrdiv24_fs426_not0;
  wire f_arrdiv24_fs426_and0;
  wire f_arrdiv24_fs426_xor1;
  wire f_arrdiv24_fs426_not1;
  wire f_arrdiv24_fs426_and1;
  wire f_arrdiv24_fs426_or0;
  wire f_arrdiv24_fs427_xor0;
  wire f_arrdiv24_fs427_not0;
  wire f_arrdiv24_fs427_and0;
  wire f_arrdiv24_fs427_xor1;
  wire f_arrdiv24_fs427_not1;
  wire f_arrdiv24_fs427_and1;
  wire f_arrdiv24_fs427_or0;
  wire f_arrdiv24_fs428_xor0;
  wire f_arrdiv24_fs428_not0;
  wire f_arrdiv24_fs428_and0;
  wire f_arrdiv24_fs428_xor1;
  wire f_arrdiv24_fs428_not1;
  wire f_arrdiv24_fs428_and1;
  wire f_arrdiv24_fs428_or0;
  wire f_arrdiv24_fs429_xor0;
  wire f_arrdiv24_fs429_not0;
  wire f_arrdiv24_fs429_and0;
  wire f_arrdiv24_fs429_xor1;
  wire f_arrdiv24_fs429_not1;
  wire f_arrdiv24_fs429_and1;
  wire f_arrdiv24_fs429_or0;
  wire f_arrdiv24_fs430_xor0;
  wire f_arrdiv24_fs430_not0;
  wire f_arrdiv24_fs430_and0;
  wire f_arrdiv24_fs430_xor1;
  wire f_arrdiv24_fs430_not1;
  wire f_arrdiv24_fs430_and1;
  wire f_arrdiv24_fs430_or0;
  wire f_arrdiv24_fs431_xor0;
  wire f_arrdiv24_fs431_not0;
  wire f_arrdiv24_fs431_and0;
  wire f_arrdiv24_fs431_xor1;
  wire f_arrdiv24_fs431_not1;
  wire f_arrdiv24_fs431_and1;
  wire f_arrdiv24_fs431_or0;
  wire f_arrdiv24_mux2to1391_and0;
  wire f_arrdiv24_mux2to1391_not0;
  wire f_arrdiv24_mux2to1391_and1;
  wire f_arrdiv24_mux2to1391_xor0;
  wire f_arrdiv24_mux2to1392_and0;
  wire f_arrdiv24_mux2to1392_not0;
  wire f_arrdiv24_mux2to1392_and1;
  wire f_arrdiv24_mux2to1392_xor0;
  wire f_arrdiv24_mux2to1393_and0;
  wire f_arrdiv24_mux2to1393_not0;
  wire f_arrdiv24_mux2to1393_and1;
  wire f_arrdiv24_mux2to1393_xor0;
  wire f_arrdiv24_mux2to1394_and0;
  wire f_arrdiv24_mux2to1394_not0;
  wire f_arrdiv24_mux2to1394_and1;
  wire f_arrdiv24_mux2to1394_xor0;
  wire f_arrdiv24_mux2to1395_and0;
  wire f_arrdiv24_mux2to1395_not0;
  wire f_arrdiv24_mux2to1395_and1;
  wire f_arrdiv24_mux2to1395_xor0;
  wire f_arrdiv24_mux2to1396_and0;
  wire f_arrdiv24_mux2to1396_not0;
  wire f_arrdiv24_mux2to1396_and1;
  wire f_arrdiv24_mux2to1396_xor0;
  wire f_arrdiv24_mux2to1397_and0;
  wire f_arrdiv24_mux2to1397_not0;
  wire f_arrdiv24_mux2to1397_and1;
  wire f_arrdiv24_mux2to1397_xor0;
  wire f_arrdiv24_mux2to1398_and0;
  wire f_arrdiv24_mux2to1398_not0;
  wire f_arrdiv24_mux2to1398_and1;
  wire f_arrdiv24_mux2to1398_xor0;
  wire f_arrdiv24_mux2to1399_and0;
  wire f_arrdiv24_mux2to1399_not0;
  wire f_arrdiv24_mux2to1399_and1;
  wire f_arrdiv24_mux2to1399_xor0;
  wire f_arrdiv24_mux2to1400_and0;
  wire f_arrdiv24_mux2to1400_not0;
  wire f_arrdiv24_mux2to1400_and1;
  wire f_arrdiv24_mux2to1400_xor0;
  wire f_arrdiv24_mux2to1401_and0;
  wire f_arrdiv24_mux2to1401_not0;
  wire f_arrdiv24_mux2to1401_and1;
  wire f_arrdiv24_mux2to1401_xor0;
  wire f_arrdiv24_mux2to1402_and0;
  wire f_arrdiv24_mux2to1402_not0;
  wire f_arrdiv24_mux2to1402_and1;
  wire f_arrdiv24_mux2to1402_xor0;
  wire f_arrdiv24_mux2to1403_and0;
  wire f_arrdiv24_mux2to1403_not0;
  wire f_arrdiv24_mux2to1403_and1;
  wire f_arrdiv24_mux2to1403_xor0;
  wire f_arrdiv24_mux2to1404_and0;
  wire f_arrdiv24_mux2to1404_not0;
  wire f_arrdiv24_mux2to1404_and1;
  wire f_arrdiv24_mux2to1404_xor0;
  wire f_arrdiv24_mux2to1405_and0;
  wire f_arrdiv24_mux2to1405_not0;
  wire f_arrdiv24_mux2to1405_and1;
  wire f_arrdiv24_mux2to1405_xor0;
  wire f_arrdiv24_mux2to1406_and0;
  wire f_arrdiv24_mux2to1406_not0;
  wire f_arrdiv24_mux2to1406_and1;
  wire f_arrdiv24_mux2to1406_xor0;
  wire f_arrdiv24_mux2to1407_and0;
  wire f_arrdiv24_mux2to1407_not0;
  wire f_arrdiv24_mux2to1407_and1;
  wire f_arrdiv24_mux2to1407_xor0;
  wire f_arrdiv24_mux2to1408_and0;
  wire f_arrdiv24_mux2to1408_not0;
  wire f_arrdiv24_mux2to1408_and1;
  wire f_arrdiv24_mux2to1408_xor0;
  wire f_arrdiv24_mux2to1409_and0;
  wire f_arrdiv24_mux2to1409_not0;
  wire f_arrdiv24_mux2to1409_and1;
  wire f_arrdiv24_mux2to1409_xor0;
  wire f_arrdiv24_mux2to1410_and0;
  wire f_arrdiv24_mux2to1410_not0;
  wire f_arrdiv24_mux2to1410_and1;
  wire f_arrdiv24_mux2to1410_xor0;
  wire f_arrdiv24_mux2to1411_and0;
  wire f_arrdiv24_mux2to1411_not0;
  wire f_arrdiv24_mux2to1411_and1;
  wire f_arrdiv24_mux2to1411_xor0;
  wire f_arrdiv24_mux2to1412_and0;
  wire f_arrdiv24_mux2to1412_not0;
  wire f_arrdiv24_mux2to1412_and1;
  wire f_arrdiv24_mux2to1412_xor0;
  wire f_arrdiv24_mux2to1413_and0;
  wire f_arrdiv24_mux2to1413_not0;
  wire f_arrdiv24_mux2to1413_and1;
  wire f_arrdiv24_mux2to1413_xor0;
  wire f_arrdiv24_not17;
  wire f_arrdiv24_fs432_xor0;
  wire f_arrdiv24_fs432_not0;
  wire f_arrdiv24_fs432_and0;
  wire f_arrdiv24_fs432_not1;
  wire f_arrdiv24_fs433_xor0;
  wire f_arrdiv24_fs433_not0;
  wire f_arrdiv24_fs433_and0;
  wire f_arrdiv24_fs433_xor1;
  wire f_arrdiv24_fs433_not1;
  wire f_arrdiv24_fs433_and1;
  wire f_arrdiv24_fs433_or0;
  wire f_arrdiv24_fs434_xor0;
  wire f_arrdiv24_fs434_not0;
  wire f_arrdiv24_fs434_and0;
  wire f_arrdiv24_fs434_xor1;
  wire f_arrdiv24_fs434_not1;
  wire f_arrdiv24_fs434_and1;
  wire f_arrdiv24_fs434_or0;
  wire f_arrdiv24_fs435_xor0;
  wire f_arrdiv24_fs435_not0;
  wire f_arrdiv24_fs435_and0;
  wire f_arrdiv24_fs435_xor1;
  wire f_arrdiv24_fs435_not1;
  wire f_arrdiv24_fs435_and1;
  wire f_arrdiv24_fs435_or0;
  wire f_arrdiv24_fs436_xor0;
  wire f_arrdiv24_fs436_not0;
  wire f_arrdiv24_fs436_and0;
  wire f_arrdiv24_fs436_xor1;
  wire f_arrdiv24_fs436_not1;
  wire f_arrdiv24_fs436_and1;
  wire f_arrdiv24_fs436_or0;
  wire f_arrdiv24_fs437_xor0;
  wire f_arrdiv24_fs437_not0;
  wire f_arrdiv24_fs437_and0;
  wire f_arrdiv24_fs437_xor1;
  wire f_arrdiv24_fs437_not1;
  wire f_arrdiv24_fs437_and1;
  wire f_arrdiv24_fs437_or0;
  wire f_arrdiv24_fs438_xor0;
  wire f_arrdiv24_fs438_not0;
  wire f_arrdiv24_fs438_and0;
  wire f_arrdiv24_fs438_xor1;
  wire f_arrdiv24_fs438_not1;
  wire f_arrdiv24_fs438_and1;
  wire f_arrdiv24_fs438_or0;
  wire f_arrdiv24_fs439_xor0;
  wire f_arrdiv24_fs439_not0;
  wire f_arrdiv24_fs439_and0;
  wire f_arrdiv24_fs439_xor1;
  wire f_arrdiv24_fs439_not1;
  wire f_arrdiv24_fs439_and1;
  wire f_arrdiv24_fs439_or0;
  wire f_arrdiv24_fs440_xor0;
  wire f_arrdiv24_fs440_not0;
  wire f_arrdiv24_fs440_and0;
  wire f_arrdiv24_fs440_xor1;
  wire f_arrdiv24_fs440_not1;
  wire f_arrdiv24_fs440_and1;
  wire f_arrdiv24_fs440_or0;
  wire f_arrdiv24_fs441_xor0;
  wire f_arrdiv24_fs441_not0;
  wire f_arrdiv24_fs441_and0;
  wire f_arrdiv24_fs441_xor1;
  wire f_arrdiv24_fs441_not1;
  wire f_arrdiv24_fs441_and1;
  wire f_arrdiv24_fs441_or0;
  wire f_arrdiv24_fs442_xor0;
  wire f_arrdiv24_fs442_not0;
  wire f_arrdiv24_fs442_and0;
  wire f_arrdiv24_fs442_xor1;
  wire f_arrdiv24_fs442_not1;
  wire f_arrdiv24_fs442_and1;
  wire f_arrdiv24_fs442_or0;
  wire f_arrdiv24_fs443_xor0;
  wire f_arrdiv24_fs443_not0;
  wire f_arrdiv24_fs443_and0;
  wire f_arrdiv24_fs443_xor1;
  wire f_arrdiv24_fs443_not1;
  wire f_arrdiv24_fs443_and1;
  wire f_arrdiv24_fs443_or0;
  wire f_arrdiv24_fs444_xor0;
  wire f_arrdiv24_fs444_not0;
  wire f_arrdiv24_fs444_and0;
  wire f_arrdiv24_fs444_xor1;
  wire f_arrdiv24_fs444_not1;
  wire f_arrdiv24_fs444_and1;
  wire f_arrdiv24_fs444_or0;
  wire f_arrdiv24_fs445_xor0;
  wire f_arrdiv24_fs445_not0;
  wire f_arrdiv24_fs445_and0;
  wire f_arrdiv24_fs445_xor1;
  wire f_arrdiv24_fs445_not1;
  wire f_arrdiv24_fs445_and1;
  wire f_arrdiv24_fs445_or0;
  wire f_arrdiv24_fs446_xor0;
  wire f_arrdiv24_fs446_not0;
  wire f_arrdiv24_fs446_and0;
  wire f_arrdiv24_fs446_xor1;
  wire f_arrdiv24_fs446_not1;
  wire f_arrdiv24_fs446_and1;
  wire f_arrdiv24_fs446_or0;
  wire f_arrdiv24_fs447_xor0;
  wire f_arrdiv24_fs447_not0;
  wire f_arrdiv24_fs447_and0;
  wire f_arrdiv24_fs447_xor1;
  wire f_arrdiv24_fs447_not1;
  wire f_arrdiv24_fs447_and1;
  wire f_arrdiv24_fs447_or0;
  wire f_arrdiv24_fs448_xor0;
  wire f_arrdiv24_fs448_not0;
  wire f_arrdiv24_fs448_and0;
  wire f_arrdiv24_fs448_xor1;
  wire f_arrdiv24_fs448_not1;
  wire f_arrdiv24_fs448_and1;
  wire f_arrdiv24_fs448_or0;
  wire f_arrdiv24_fs449_xor0;
  wire f_arrdiv24_fs449_not0;
  wire f_arrdiv24_fs449_and0;
  wire f_arrdiv24_fs449_xor1;
  wire f_arrdiv24_fs449_not1;
  wire f_arrdiv24_fs449_and1;
  wire f_arrdiv24_fs449_or0;
  wire f_arrdiv24_fs450_xor0;
  wire f_arrdiv24_fs450_not0;
  wire f_arrdiv24_fs450_and0;
  wire f_arrdiv24_fs450_xor1;
  wire f_arrdiv24_fs450_not1;
  wire f_arrdiv24_fs450_and1;
  wire f_arrdiv24_fs450_or0;
  wire f_arrdiv24_fs451_xor0;
  wire f_arrdiv24_fs451_not0;
  wire f_arrdiv24_fs451_and0;
  wire f_arrdiv24_fs451_xor1;
  wire f_arrdiv24_fs451_not1;
  wire f_arrdiv24_fs451_and1;
  wire f_arrdiv24_fs451_or0;
  wire f_arrdiv24_fs452_xor0;
  wire f_arrdiv24_fs452_not0;
  wire f_arrdiv24_fs452_and0;
  wire f_arrdiv24_fs452_xor1;
  wire f_arrdiv24_fs452_not1;
  wire f_arrdiv24_fs452_and1;
  wire f_arrdiv24_fs452_or0;
  wire f_arrdiv24_fs453_xor0;
  wire f_arrdiv24_fs453_not0;
  wire f_arrdiv24_fs453_and0;
  wire f_arrdiv24_fs453_xor1;
  wire f_arrdiv24_fs453_not1;
  wire f_arrdiv24_fs453_and1;
  wire f_arrdiv24_fs453_or0;
  wire f_arrdiv24_fs454_xor0;
  wire f_arrdiv24_fs454_not0;
  wire f_arrdiv24_fs454_and0;
  wire f_arrdiv24_fs454_xor1;
  wire f_arrdiv24_fs454_not1;
  wire f_arrdiv24_fs454_and1;
  wire f_arrdiv24_fs454_or0;
  wire f_arrdiv24_fs455_xor0;
  wire f_arrdiv24_fs455_not0;
  wire f_arrdiv24_fs455_and0;
  wire f_arrdiv24_fs455_xor1;
  wire f_arrdiv24_fs455_not1;
  wire f_arrdiv24_fs455_and1;
  wire f_arrdiv24_fs455_or0;
  wire f_arrdiv24_mux2to1414_and0;
  wire f_arrdiv24_mux2to1414_not0;
  wire f_arrdiv24_mux2to1414_and1;
  wire f_arrdiv24_mux2to1414_xor0;
  wire f_arrdiv24_mux2to1415_and0;
  wire f_arrdiv24_mux2to1415_not0;
  wire f_arrdiv24_mux2to1415_and1;
  wire f_arrdiv24_mux2to1415_xor0;
  wire f_arrdiv24_mux2to1416_and0;
  wire f_arrdiv24_mux2to1416_not0;
  wire f_arrdiv24_mux2to1416_and1;
  wire f_arrdiv24_mux2to1416_xor0;
  wire f_arrdiv24_mux2to1417_and0;
  wire f_arrdiv24_mux2to1417_not0;
  wire f_arrdiv24_mux2to1417_and1;
  wire f_arrdiv24_mux2to1417_xor0;
  wire f_arrdiv24_mux2to1418_and0;
  wire f_arrdiv24_mux2to1418_not0;
  wire f_arrdiv24_mux2to1418_and1;
  wire f_arrdiv24_mux2to1418_xor0;
  wire f_arrdiv24_mux2to1419_and0;
  wire f_arrdiv24_mux2to1419_not0;
  wire f_arrdiv24_mux2to1419_and1;
  wire f_arrdiv24_mux2to1419_xor0;
  wire f_arrdiv24_mux2to1420_and0;
  wire f_arrdiv24_mux2to1420_not0;
  wire f_arrdiv24_mux2to1420_and1;
  wire f_arrdiv24_mux2to1420_xor0;
  wire f_arrdiv24_mux2to1421_and0;
  wire f_arrdiv24_mux2to1421_not0;
  wire f_arrdiv24_mux2to1421_and1;
  wire f_arrdiv24_mux2to1421_xor0;
  wire f_arrdiv24_mux2to1422_and0;
  wire f_arrdiv24_mux2to1422_not0;
  wire f_arrdiv24_mux2to1422_and1;
  wire f_arrdiv24_mux2to1422_xor0;
  wire f_arrdiv24_mux2to1423_and0;
  wire f_arrdiv24_mux2to1423_not0;
  wire f_arrdiv24_mux2to1423_and1;
  wire f_arrdiv24_mux2to1423_xor0;
  wire f_arrdiv24_mux2to1424_and0;
  wire f_arrdiv24_mux2to1424_not0;
  wire f_arrdiv24_mux2to1424_and1;
  wire f_arrdiv24_mux2to1424_xor0;
  wire f_arrdiv24_mux2to1425_and0;
  wire f_arrdiv24_mux2to1425_not0;
  wire f_arrdiv24_mux2to1425_and1;
  wire f_arrdiv24_mux2to1425_xor0;
  wire f_arrdiv24_mux2to1426_and0;
  wire f_arrdiv24_mux2to1426_not0;
  wire f_arrdiv24_mux2to1426_and1;
  wire f_arrdiv24_mux2to1426_xor0;
  wire f_arrdiv24_mux2to1427_and0;
  wire f_arrdiv24_mux2to1427_not0;
  wire f_arrdiv24_mux2to1427_and1;
  wire f_arrdiv24_mux2to1427_xor0;
  wire f_arrdiv24_mux2to1428_and0;
  wire f_arrdiv24_mux2to1428_not0;
  wire f_arrdiv24_mux2to1428_and1;
  wire f_arrdiv24_mux2to1428_xor0;
  wire f_arrdiv24_mux2to1429_and0;
  wire f_arrdiv24_mux2to1429_not0;
  wire f_arrdiv24_mux2to1429_and1;
  wire f_arrdiv24_mux2to1429_xor0;
  wire f_arrdiv24_mux2to1430_and0;
  wire f_arrdiv24_mux2to1430_not0;
  wire f_arrdiv24_mux2to1430_and1;
  wire f_arrdiv24_mux2to1430_xor0;
  wire f_arrdiv24_mux2to1431_and0;
  wire f_arrdiv24_mux2to1431_not0;
  wire f_arrdiv24_mux2to1431_and1;
  wire f_arrdiv24_mux2to1431_xor0;
  wire f_arrdiv24_mux2to1432_and0;
  wire f_arrdiv24_mux2to1432_not0;
  wire f_arrdiv24_mux2to1432_and1;
  wire f_arrdiv24_mux2to1432_xor0;
  wire f_arrdiv24_mux2to1433_and0;
  wire f_arrdiv24_mux2to1433_not0;
  wire f_arrdiv24_mux2to1433_and1;
  wire f_arrdiv24_mux2to1433_xor0;
  wire f_arrdiv24_mux2to1434_and0;
  wire f_arrdiv24_mux2to1434_not0;
  wire f_arrdiv24_mux2to1434_and1;
  wire f_arrdiv24_mux2to1434_xor0;
  wire f_arrdiv24_mux2to1435_and0;
  wire f_arrdiv24_mux2to1435_not0;
  wire f_arrdiv24_mux2to1435_and1;
  wire f_arrdiv24_mux2to1435_xor0;
  wire f_arrdiv24_mux2to1436_and0;
  wire f_arrdiv24_mux2to1436_not0;
  wire f_arrdiv24_mux2to1436_and1;
  wire f_arrdiv24_mux2to1436_xor0;
  wire f_arrdiv24_not18;
  wire f_arrdiv24_fs456_xor0;
  wire f_arrdiv24_fs456_not0;
  wire f_arrdiv24_fs456_and0;
  wire f_arrdiv24_fs456_not1;
  wire f_arrdiv24_fs457_xor0;
  wire f_arrdiv24_fs457_not0;
  wire f_arrdiv24_fs457_and0;
  wire f_arrdiv24_fs457_xor1;
  wire f_arrdiv24_fs457_not1;
  wire f_arrdiv24_fs457_and1;
  wire f_arrdiv24_fs457_or0;
  wire f_arrdiv24_fs458_xor0;
  wire f_arrdiv24_fs458_not0;
  wire f_arrdiv24_fs458_and0;
  wire f_arrdiv24_fs458_xor1;
  wire f_arrdiv24_fs458_not1;
  wire f_arrdiv24_fs458_and1;
  wire f_arrdiv24_fs458_or0;
  wire f_arrdiv24_fs459_xor0;
  wire f_arrdiv24_fs459_not0;
  wire f_arrdiv24_fs459_and0;
  wire f_arrdiv24_fs459_xor1;
  wire f_arrdiv24_fs459_not1;
  wire f_arrdiv24_fs459_and1;
  wire f_arrdiv24_fs459_or0;
  wire f_arrdiv24_fs460_xor0;
  wire f_arrdiv24_fs460_not0;
  wire f_arrdiv24_fs460_and0;
  wire f_arrdiv24_fs460_xor1;
  wire f_arrdiv24_fs460_not1;
  wire f_arrdiv24_fs460_and1;
  wire f_arrdiv24_fs460_or0;
  wire f_arrdiv24_fs461_xor0;
  wire f_arrdiv24_fs461_not0;
  wire f_arrdiv24_fs461_and0;
  wire f_arrdiv24_fs461_xor1;
  wire f_arrdiv24_fs461_not1;
  wire f_arrdiv24_fs461_and1;
  wire f_arrdiv24_fs461_or0;
  wire f_arrdiv24_fs462_xor0;
  wire f_arrdiv24_fs462_not0;
  wire f_arrdiv24_fs462_and0;
  wire f_arrdiv24_fs462_xor1;
  wire f_arrdiv24_fs462_not1;
  wire f_arrdiv24_fs462_and1;
  wire f_arrdiv24_fs462_or0;
  wire f_arrdiv24_fs463_xor0;
  wire f_arrdiv24_fs463_not0;
  wire f_arrdiv24_fs463_and0;
  wire f_arrdiv24_fs463_xor1;
  wire f_arrdiv24_fs463_not1;
  wire f_arrdiv24_fs463_and1;
  wire f_arrdiv24_fs463_or0;
  wire f_arrdiv24_fs464_xor0;
  wire f_arrdiv24_fs464_not0;
  wire f_arrdiv24_fs464_and0;
  wire f_arrdiv24_fs464_xor1;
  wire f_arrdiv24_fs464_not1;
  wire f_arrdiv24_fs464_and1;
  wire f_arrdiv24_fs464_or0;
  wire f_arrdiv24_fs465_xor0;
  wire f_arrdiv24_fs465_not0;
  wire f_arrdiv24_fs465_and0;
  wire f_arrdiv24_fs465_xor1;
  wire f_arrdiv24_fs465_not1;
  wire f_arrdiv24_fs465_and1;
  wire f_arrdiv24_fs465_or0;
  wire f_arrdiv24_fs466_xor0;
  wire f_arrdiv24_fs466_not0;
  wire f_arrdiv24_fs466_and0;
  wire f_arrdiv24_fs466_xor1;
  wire f_arrdiv24_fs466_not1;
  wire f_arrdiv24_fs466_and1;
  wire f_arrdiv24_fs466_or0;
  wire f_arrdiv24_fs467_xor0;
  wire f_arrdiv24_fs467_not0;
  wire f_arrdiv24_fs467_and0;
  wire f_arrdiv24_fs467_xor1;
  wire f_arrdiv24_fs467_not1;
  wire f_arrdiv24_fs467_and1;
  wire f_arrdiv24_fs467_or0;
  wire f_arrdiv24_fs468_xor0;
  wire f_arrdiv24_fs468_not0;
  wire f_arrdiv24_fs468_and0;
  wire f_arrdiv24_fs468_xor1;
  wire f_arrdiv24_fs468_not1;
  wire f_arrdiv24_fs468_and1;
  wire f_arrdiv24_fs468_or0;
  wire f_arrdiv24_fs469_xor0;
  wire f_arrdiv24_fs469_not0;
  wire f_arrdiv24_fs469_and0;
  wire f_arrdiv24_fs469_xor1;
  wire f_arrdiv24_fs469_not1;
  wire f_arrdiv24_fs469_and1;
  wire f_arrdiv24_fs469_or0;
  wire f_arrdiv24_fs470_xor0;
  wire f_arrdiv24_fs470_not0;
  wire f_arrdiv24_fs470_and0;
  wire f_arrdiv24_fs470_xor1;
  wire f_arrdiv24_fs470_not1;
  wire f_arrdiv24_fs470_and1;
  wire f_arrdiv24_fs470_or0;
  wire f_arrdiv24_fs471_xor0;
  wire f_arrdiv24_fs471_not0;
  wire f_arrdiv24_fs471_and0;
  wire f_arrdiv24_fs471_xor1;
  wire f_arrdiv24_fs471_not1;
  wire f_arrdiv24_fs471_and1;
  wire f_arrdiv24_fs471_or0;
  wire f_arrdiv24_fs472_xor0;
  wire f_arrdiv24_fs472_not0;
  wire f_arrdiv24_fs472_and0;
  wire f_arrdiv24_fs472_xor1;
  wire f_arrdiv24_fs472_not1;
  wire f_arrdiv24_fs472_and1;
  wire f_arrdiv24_fs472_or0;
  wire f_arrdiv24_fs473_xor0;
  wire f_arrdiv24_fs473_not0;
  wire f_arrdiv24_fs473_and0;
  wire f_arrdiv24_fs473_xor1;
  wire f_arrdiv24_fs473_not1;
  wire f_arrdiv24_fs473_and1;
  wire f_arrdiv24_fs473_or0;
  wire f_arrdiv24_fs474_xor0;
  wire f_arrdiv24_fs474_not0;
  wire f_arrdiv24_fs474_and0;
  wire f_arrdiv24_fs474_xor1;
  wire f_arrdiv24_fs474_not1;
  wire f_arrdiv24_fs474_and1;
  wire f_arrdiv24_fs474_or0;
  wire f_arrdiv24_fs475_xor0;
  wire f_arrdiv24_fs475_not0;
  wire f_arrdiv24_fs475_and0;
  wire f_arrdiv24_fs475_xor1;
  wire f_arrdiv24_fs475_not1;
  wire f_arrdiv24_fs475_and1;
  wire f_arrdiv24_fs475_or0;
  wire f_arrdiv24_fs476_xor0;
  wire f_arrdiv24_fs476_not0;
  wire f_arrdiv24_fs476_and0;
  wire f_arrdiv24_fs476_xor1;
  wire f_arrdiv24_fs476_not1;
  wire f_arrdiv24_fs476_and1;
  wire f_arrdiv24_fs476_or0;
  wire f_arrdiv24_fs477_xor0;
  wire f_arrdiv24_fs477_not0;
  wire f_arrdiv24_fs477_and0;
  wire f_arrdiv24_fs477_xor1;
  wire f_arrdiv24_fs477_not1;
  wire f_arrdiv24_fs477_and1;
  wire f_arrdiv24_fs477_or0;
  wire f_arrdiv24_fs478_xor0;
  wire f_arrdiv24_fs478_not0;
  wire f_arrdiv24_fs478_and0;
  wire f_arrdiv24_fs478_xor1;
  wire f_arrdiv24_fs478_not1;
  wire f_arrdiv24_fs478_and1;
  wire f_arrdiv24_fs478_or0;
  wire f_arrdiv24_fs479_xor0;
  wire f_arrdiv24_fs479_not0;
  wire f_arrdiv24_fs479_and0;
  wire f_arrdiv24_fs479_xor1;
  wire f_arrdiv24_fs479_not1;
  wire f_arrdiv24_fs479_and1;
  wire f_arrdiv24_fs479_or0;
  wire f_arrdiv24_mux2to1437_and0;
  wire f_arrdiv24_mux2to1437_not0;
  wire f_arrdiv24_mux2to1437_and1;
  wire f_arrdiv24_mux2to1437_xor0;
  wire f_arrdiv24_mux2to1438_and0;
  wire f_arrdiv24_mux2to1438_not0;
  wire f_arrdiv24_mux2to1438_and1;
  wire f_arrdiv24_mux2to1438_xor0;
  wire f_arrdiv24_mux2to1439_and0;
  wire f_arrdiv24_mux2to1439_not0;
  wire f_arrdiv24_mux2to1439_and1;
  wire f_arrdiv24_mux2to1439_xor0;
  wire f_arrdiv24_mux2to1440_and0;
  wire f_arrdiv24_mux2to1440_not0;
  wire f_arrdiv24_mux2to1440_and1;
  wire f_arrdiv24_mux2to1440_xor0;
  wire f_arrdiv24_mux2to1441_and0;
  wire f_arrdiv24_mux2to1441_not0;
  wire f_arrdiv24_mux2to1441_and1;
  wire f_arrdiv24_mux2to1441_xor0;
  wire f_arrdiv24_mux2to1442_and0;
  wire f_arrdiv24_mux2to1442_not0;
  wire f_arrdiv24_mux2to1442_and1;
  wire f_arrdiv24_mux2to1442_xor0;
  wire f_arrdiv24_mux2to1443_and0;
  wire f_arrdiv24_mux2to1443_not0;
  wire f_arrdiv24_mux2to1443_and1;
  wire f_arrdiv24_mux2to1443_xor0;
  wire f_arrdiv24_mux2to1444_and0;
  wire f_arrdiv24_mux2to1444_not0;
  wire f_arrdiv24_mux2to1444_and1;
  wire f_arrdiv24_mux2to1444_xor0;
  wire f_arrdiv24_mux2to1445_and0;
  wire f_arrdiv24_mux2to1445_not0;
  wire f_arrdiv24_mux2to1445_and1;
  wire f_arrdiv24_mux2to1445_xor0;
  wire f_arrdiv24_mux2to1446_and0;
  wire f_arrdiv24_mux2to1446_not0;
  wire f_arrdiv24_mux2to1446_and1;
  wire f_arrdiv24_mux2to1446_xor0;
  wire f_arrdiv24_mux2to1447_and0;
  wire f_arrdiv24_mux2to1447_not0;
  wire f_arrdiv24_mux2to1447_and1;
  wire f_arrdiv24_mux2to1447_xor0;
  wire f_arrdiv24_mux2to1448_and0;
  wire f_arrdiv24_mux2to1448_not0;
  wire f_arrdiv24_mux2to1448_and1;
  wire f_arrdiv24_mux2to1448_xor0;
  wire f_arrdiv24_mux2to1449_and0;
  wire f_arrdiv24_mux2to1449_not0;
  wire f_arrdiv24_mux2to1449_and1;
  wire f_arrdiv24_mux2to1449_xor0;
  wire f_arrdiv24_mux2to1450_and0;
  wire f_arrdiv24_mux2to1450_not0;
  wire f_arrdiv24_mux2to1450_and1;
  wire f_arrdiv24_mux2to1450_xor0;
  wire f_arrdiv24_mux2to1451_and0;
  wire f_arrdiv24_mux2to1451_not0;
  wire f_arrdiv24_mux2to1451_and1;
  wire f_arrdiv24_mux2to1451_xor0;
  wire f_arrdiv24_mux2to1452_and0;
  wire f_arrdiv24_mux2to1452_not0;
  wire f_arrdiv24_mux2to1452_and1;
  wire f_arrdiv24_mux2to1452_xor0;
  wire f_arrdiv24_mux2to1453_and0;
  wire f_arrdiv24_mux2to1453_not0;
  wire f_arrdiv24_mux2to1453_and1;
  wire f_arrdiv24_mux2to1453_xor0;
  wire f_arrdiv24_mux2to1454_and0;
  wire f_arrdiv24_mux2to1454_not0;
  wire f_arrdiv24_mux2to1454_and1;
  wire f_arrdiv24_mux2to1454_xor0;
  wire f_arrdiv24_mux2to1455_and0;
  wire f_arrdiv24_mux2to1455_not0;
  wire f_arrdiv24_mux2to1455_and1;
  wire f_arrdiv24_mux2to1455_xor0;
  wire f_arrdiv24_mux2to1456_and0;
  wire f_arrdiv24_mux2to1456_not0;
  wire f_arrdiv24_mux2to1456_and1;
  wire f_arrdiv24_mux2to1456_xor0;
  wire f_arrdiv24_mux2to1457_and0;
  wire f_arrdiv24_mux2to1457_not0;
  wire f_arrdiv24_mux2to1457_and1;
  wire f_arrdiv24_mux2to1457_xor0;
  wire f_arrdiv24_mux2to1458_and0;
  wire f_arrdiv24_mux2to1458_not0;
  wire f_arrdiv24_mux2to1458_and1;
  wire f_arrdiv24_mux2to1458_xor0;
  wire f_arrdiv24_mux2to1459_and0;
  wire f_arrdiv24_mux2to1459_not0;
  wire f_arrdiv24_mux2to1459_and1;
  wire f_arrdiv24_mux2to1459_xor0;
  wire f_arrdiv24_not19;
  wire f_arrdiv24_fs480_xor0;
  wire f_arrdiv24_fs480_not0;
  wire f_arrdiv24_fs480_and0;
  wire f_arrdiv24_fs480_not1;
  wire f_arrdiv24_fs481_xor0;
  wire f_arrdiv24_fs481_not0;
  wire f_arrdiv24_fs481_and0;
  wire f_arrdiv24_fs481_xor1;
  wire f_arrdiv24_fs481_not1;
  wire f_arrdiv24_fs481_and1;
  wire f_arrdiv24_fs481_or0;
  wire f_arrdiv24_fs482_xor0;
  wire f_arrdiv24_fs482_not0;
  wire f_arrdiv24_fs482_and0;
  wire f_arrdiv24_fs482_xor1;
  wire f_arrdiv24_fs482_not1;
  wire f_arrdiv24_fs482_and1;
  wire f_arrdiv24_fs482_or0;
  wire f_arrdiv24_fs483_xor0;
  wire f_arrdiv24_fs483_not0;
  wire f_arrdiv24_fs483_and0;
  wire f_arrdiv24_fs483_xor1;
  wire f_arrdiv24_fs483_not1;
  wire f_arrdiv24_fs483_and1;
  wire f_arrdiv24_fs483_or0;
  wire f_arrdiv24_fs484_xor0;
  wire f_arrdiv24_fs484_not0;
  wire f_arrdiv24_fs484_and0;
  wire f_arrdiv24_fs484_xor1;
  wire f_arrdiv24_fs484_not1;
  wire f_arrdiv24_fs484_and1;
  wire f_arrdiv24_fs484_or0;
  wire f_arrdiv24_fs485_xor0;
  wire f_arrdiv24_fs485_not0;
  wire f_arrdiv24_fs485_and0;
  wire f_arrdiv24_fs485_xor1;
  wire f_arrdiv24_fs485_not1;
  wire f_arrdiv24_fs485_and1;
  wire f_arrdiv24_fs485_or0;
  wire f_arrdiv24_fs486_xor0;
  wire f_arrdiv24_fs486_not0;
  wire f_arrdiv24_fs486_and0;
  wire f_arrdiv24_fs486_xor1;
  wire f_arrdiv24_fs486_not1;
  wire f_arrdiv24_fs486_and1;
  wire f_arrdiv24_fs486_or0;
  wire f_arrdiv24_fs487_xor0;
  wire f_arrdiv24_fs487_not0;
  wire f_arrdiv24_fs487_and0;
  wire f_arrdiv24_fs487_xor1;
  wire f_arrdiv24_fs487_not1;
  wire f_arrdiv24_fs487_and1;
  wire f_arrdiv24_fs487_or0;
  wire f_arrdiv24_fs488_xor0;
  wire f_arrdiv24_fs488_not0;
  wire f_arrdiv24_fs488_and0;
  wire f_arrdiv24_fs488_xor1;
  wire f_arrdiv24_fs488_not1;
  wire f_arrdiv24_fs488_and1;
  wire f_arrdiv24_fs488_or0;
  wire f_arrdiv24_fs489_xor0;
  wire f_arrdiv24_fs489_not0;
  wire f_arrdiv24_fs489_and0;
  wire f_arrdiv24_fs489_xor1;
  wire f_arrdiv24_fs489_not1;
  wire f_arrdiv24_fs489_and1;
  wire f_arrdiv24_fs489_or0;
  wire f_arrdiv24_fs490_xor0;
  wire f_arrdiv24_fs490_not0;
  wire f_arrdiv24_fs490_and0;
  wire f_arrdiv24_fs490_xor1;
  wire f_arrdiv24_fs490_not1;
  wire f_arrdiv24_fs490_and1;
  wire f_arrdiv24_fs490_or0;
  wire f_arrdiv24_fs491_xor0;
  wire f_arrdiv24_fs491_not0;
  wire f_arrdiv24_fs491_and0;
  wire f_arrdiv24_fs491_xor1;
  wire f_arrdiv24_fs491_not1;
  wire f_arrdiv24_fs491_and1;
  wire f_arrdiv24_fs491_or0;
  wire f_arrdiv24_fs492_xor0;
  wire f_arrdiv24_fs492_not0;
  wire f_arrdiv24_fs492_and0;
  wire f_arrdiv24_fs492_xor1;
  wire f_arrdiv24_fs492_not1;
  wire f_arrdiv24_fs492_and1;
  wire f_arrdiv24_fs492_or0;
  wire f_arrdiv24_fs493_xor0;
  wire f_arrdiv24_fs493_not0;
  wire f_arrdiv24_fs493_and0;
  wire f_arrdiv24_fs493_xor1;
  wire f_arrdiv24_fs493_not1;
  wire f_arrdiv24_fs493_and1;
  wire f_arrdiv24_fs493_or0;
  wire f_arrdiv24_fs494_xor0;
  wire f_arrdiv24_fs494_not0;
  wire f_arrdiv24_fs494_and0;
  wire f_arrdiv24_fs494_xor1;
  wire f_arrdiv24_fs494_not1;
  wire f_arrdiv24_fs494_and1;
  wire f_arrdiv24_fs494_or0;
  wire f_arrdiv24_fs495_xor0;
  wire f_arrdiv24_fs495_not0;
  wire f_arrdiv24_fs495_and0;
  wire f_arrdiv24_fs495_xor1;
  wire f_arrdiv24_fs495_not1;
  wire f_arrdiv24_fs495_and1;
  wire f_arrdiv24_fs495_or0;
  wire f_arrdiv24_fs496_xor0;
  wire f_arrdiv24_fs496_not0;
  wire f_arrdiv24_fs496_and0;
  wire f_arrdiv24_fs496_xor1;
  wire f_arrdiv24_fs496_not1;
  wire f_arrdiv24_fs496_and1;
  wire f_arrdiv24_fs496_or0;
  wire f_arrdiv24_fs497_xor0;
  wire f_arrdiv24_fs497_not0;
  wire f_arrdiv24_fs497_and0;
  wire f_arrdiv24_fs497_xor1;
  wire f_arrdiv24_fs497_not1;
  wire f_arrdiv24_fs497_and1;
  wire f_arrdiv24_fs497_or0;
  wire f_arrdiv24_fs498_xor0;
  wire f_arrdiv24_fs498_not0;
  wire f_arrdiv24_fs498_and0;
  wire f_arrdiv24_fs498_xor1;
  wire f_arrdiv24_fs498_not1;
  wire f_arrdiv24_fs498_and1;
  wire f_arrdiv24_fs498_or0;
  wire f_arrdiv24_fs499_xor0;
  wire f_arrdiv24_fs499_not0;
  wire f_arrdiv24_fs499_and0;
  wire f_arrdiv24_fs499_xor1;
  wire f_arrdiv24_fs499_not1;
  wire f_arrdiv24_fs499_and1;
  wire f_arrdiv24_fs499_or0;
  wire f_arrdiv24_fs500_xor0;
  wire f_arrdiv24_fs500_not0;
  wire f_arrdiv24_fs500_and0;
  wire f_arrdiv24_fs500_xor1;
  wire f_arrdiv24_fs500_not1;
  wire f_arrdiv24_fs500_and1;
  wire f_arrdiv24_fs500_or0;
  wire f_arrdiv24_fs501_xor0;
  wire f_arrdiv24_fs501_not0;
  wire f_arrdiv24_fs501_and0;
  wire f_arrdiv24_fs501_xor1;
  wire f_arrdiv24_fs501_not1;
  wire f_arrdiv24_fs501_and1;
  wire f_arrdiv24_fs501_or0;
  wire f_arrdiv24_fs502_xor0;
  wire f_arrdiv24_fs502_not0;
  wire f_arrdiv24_fs502_and0;
  wire f_arrdiv24_fs502_xor1;
  wire f_arrdiv24_fs502_not1;
  wire f_arrdiv24_fs502_and1;
  wire f_arrdiv24_fs502_or0;
  wire f_arrdiv24_fs503_xor0;
  wire f_arrdiv24_fs503_not0;
  wire f_arrdiv24_fs503_and0;
  wire f_arrdiv24_fs503_xor1;
  wire f_arrdiv24_fs503_not1;
  wire f_arrdiv24_fs503_and1;
  wire f_arrdiv24_fs503_or0;
  wire f_arrdiv24_mux2to1460_and0;
  wire f_arrdiv24_mux2to1460_not0;
  wire f_arrdiv24_mux2to1460_and1;
  wire f_arrdiv24_mux2to1460_xor0;
  wire f_arrdiv24_mux2to1461_and0;
  wire f_arrdiv24_mux2to1461_not0;
  wire f_arrdiv24_mux2to1461_and1;
  wire f_arrdiv24_mux2to1461_xor0;
  wire f_arrdiv24_mux2to1462_and0;
  wire f_arrdiv24_mux2to1462_not0;
  wire f_arrdiv24_mux2to1462_and1;
  wire f_arrdiv24_mux2to1462_xor0;
  wire f_arrdiv24_mux2to1463_and0;
  wire f_arrdiv24_mux2to1463_not0;
  wire f_arrdiv24_mux2to1463_and1;
  wire f_arrdiv24_mux2to1463_xor0;
  wire f_arrdiv24_mux2to1464_and0;
  wire f_arrdiv24_mux2to1464_not0;
  wire f_arrdiv24_mux2to1464_and1;
  wire f_arrdiv24_mux2to1464_xor0;
  wire f_arrdiv24_mux2to1465_and0;
  wire f_arrdiv24_mux2to1465_not0;
  wire f_arrdiv24_mux2to1465_and1;
  wire f_arrdiv24_mux2to1465_xor0;
  wire f_arrdiv24_mux2to1466_and0;
  wire f_arrdiv24_mux2to1466_not0;
  wire f_arrdiv24_mux2to1466_and1;
  wire f_arrdiv24_mux2to1466_xor0;
  wire f_arrdiv24_mux2to1467_and0;
  wire f_arrdiv24_mux2to1467_not0;
  wire f_arrdiv24_mux2to1467_and1;
  wire f_arrdiv24_mux2to1467_xor0;
  wire f_arrdiv24_mux2to1468_and0;
  wire f_arrdiv24_mux2to1468_not0;
  wire f_arrdiv24_mux2to1468_and1;
  wire f_arrdiv24_mux2to1468_xor0;
  wire f_arrdiv24_mux2to1469_and0;
  wire f_arrdiv24_mux2to1469_not0;
  wire f_arrdiv24_mux2to1469_and1;
  wire f_arrdiv24_mux2to1469_xor0;
  wire f_arrdiv24_mux2to1470_and0;
  wire f_arrdiv24_mux2to1470_not0;
  wire f_arrdiv24_mux2to1470_and1;
  wire f_arrdiv24_mux2to1470_xor0;
  wire f_arrdiv24_mux2to1471_and0;
  wire f_arrdiv24_mux2to1471_not0;
  wire f_arrdiv24_mux2to1471_and1;
  wire f_arrdiv24_mux2to1471_xor0;
  wire f_arrdiv24_mux2to1472_and0;
  wire f_arrdiv24_mux2to1472_not0;
  wire f_arrdiv24_mux2to1472_and1;
  wire f_arrdiv24_mux2to1472_xor0;
  wire f_arrdiv24_mux2to1473_and0;
  wire f_arrdiv24_mux2to1473_not0;
  wire f_arrdiv24_mux2to1473_and1;
  wire f_arrdiv24_mux2to1473_xor0;
  wire f_arrdiv24_mux2to1474_and0;
  wire f_arrdiv24_mux2to1474_not0;
  wire f_arrdiv24_mux2to1474_and1;
  wire f_arrdiv24_mux2to1474_xor0;
  wire f_arrdiv24_mux2to1475_and0;
  wire f_arrdiv24_mux2to1475_not0;
  wire f_arrdiv24_mux2to1475_and1;
  wire f_arrdiv24_mux2to1475_xor0;
  wire f_arrdiv24_mux2to1476_and0;
  wire f_arrdiv24_mux2to1476_not0;
  wire f_arrdiv24_mux2to1476_and1;
  wire f_arrdiv24_mux2to1476_xor0;
  wire f_arrdiv24_mux2to1477_and0;
  wire f_arrdiv24_mux2to1477_not0;
  wire f_arrdiv24_mux2to1477_and1;
  wire f_arrdiv24_mux2to1477_xor0;
  wire f_arrdiv24_mux2to1478_and0;
  wire f_arrdiv24_mux2to1478_not0;
  wire f_arrdiv24_mux2to1478_and1;
  wire f_arrdiv24_mux2to1478_xor0;
  wire f_arrdiv24_mux2to1479_and0;
  wire f_arrdiv24_mux2to1479_not0;
  wire f_arrdiv24_mux2to1479_and1;
  wire f_arrdiv24_mux2to1479_xor0;
  wire f_arrdiv24_mux2to1480_and0;
  wire f_arrdiv24_mux2to1480_not0;
  wire f_arrdiv24_mux2to1480_and1;
  wire f_arrdiv24_mux2to1480_xor0;
  wire f_arrdiv24_mux2to1481_and0;
  wire f_arrdiv24_mux2to1481_not0;
  wire f_arrdiv24_mux2to1481_and1;
  wire f_arrdiv24_mux2to1481_xor0;
  wire f_arrdiv24_mux2to1482_and0;
  wire f_arrdiv24_mux2to1482_not0;
  wire f_arrdiv24_mux2to1482_and1;
  wire f_arrdiv24_mux2to1482_xor0;
  wire f_arrdiv24_not20;
  wire f_arrdiv24_fs504_xor0;
  wire f_arrdiv24_fs504_not0;
  wire f_arrdiv24_fs504_and0;
  wire f_arrdiv24_fs504_not1;
  wire f_arrdiv24_fs505_xor0;
  wire f_arrdiv24_fs505_not0;
  wire f_arrdiv24_fs505_and0;
  wire f_arrdiv24_fs505_xor1;
  wire f_arrdiv24_fs505_not1;
  wire f_arrdiv24_fs505_and1;
  wire f_arrdiv24_fs505_or0;
  wire f_arrdiv24_fs506_xor0;
  wire f_arrdiv24_fs506_not0;
  wire f_arrdiv24_fs506_and0;
  wire f_arrdiv24_fs506_xor1;
  wire f_arrdiv24_fs506_not1;
  wire f_arrdiv24_fs506_and1;
  wire f_arrdiv24_fs506_or0;
  wire f_arrdiv24_fs507_xor0;
  wire f_arrdiv24_fs507_not0;
  wire f_arrdiv24_fs507_and0;
  wire f_arrdiv24_fs507_xor1;
  wire f_arrdiv24_fs507_not1;
  wire f_arrdiv24_fs507_and1;
  wire f_arrdiv24_fs507_or0;
  wire f_arrdiv24_fs508_xor0;
  wire f_arrdiv24_fs508_not0;
  wire f_arrdiv24_fs508_and0;
  wire f_arrdiv24_fs508_xor1;
  wire f_arrdiv24_fs508_not1;
  wire f_arrdiv24_fs508_and1;
  wire f_arrdiv24_fs508_or0;
  wire f_arrdiv24_fs509_xor0;
  wire f_arrdiv24_fs509_not0;
  wire f_arrdiv24_fs509_and0;
  wire f_arrdiv24_fs509_xor1;
  wire f_arrdiv24_fs509_not1;
  wire f_arrdiv24_fs509_and1;
  wire f_arrdiv24_fs509_or0;
  wire f_arrdiv24_fs510_xor0;
  wire f_arrdiv24_fs510_not0;
  wire f_arrdiv24_fs510_and0;
  wire f_arrdiv24_fs510_xor1;
  wire f_arrdiv24_fs510_not1;
  wire f_arrdiv24_fs510_and1;
  wire f_arrdiv24_fs510_or0;
  wire f_arrdiv24_fs511_xor0;
  wire f_arrdiv24_fs511_not0;
  wire f_arrdiv24_fs511_and0;
  wire f_arrdiv24_fs511_xor1;
  wire f_arrdiv24_fs511_not1;
  wire f_arrdiv24_fs511_and1;
  wire f_arrdiv24_fs511_or0;
  wire f_arrdiv24_fs512_xor0;
  wire f_arrdiv24_fs512_not0;
  wire f_arrdiv24_fs512_and0;
  wire f_arrdiv24_fs512_xor1;
  wire f_arrdiv24_fs512_not1;
  wire f_arrdiv24_fs512_and1;
  wire f_arrdiv24_fs512_or0;
  wire f_arrdiv24_fs513_xor0;
  wire f_arrdiv24_fs513_not0;
  wire f_arrdiv24_fs513_and0;
  wire f_arrdiv24_fs513_xor1;
  wire f_arrdiv24_fs513_not1;
  wire f_arrdiv24_fs513_and1;
  wire f_arrdiv24_fs513_or0;
  wire f_arrdiv24_fs514_xor0;
  wire f_arrdiv24_fs514_not0;
  wire f_arrdiv24_fs514_and0;
  wire f_arrdiv24_fs514_xor1;
  wire f_arrdiv24_fs514_not1;
  wire f_arrdiv24_fs514_and1;
  wire f_arrdiv24_fs514_or0;
  wire f_arrdiv24_fs515_xor0;
  wire f_arrdiv24_fs515_not0;
  wire f_arrdiv24_fs515_and0;
  wire f_arrdiv24_fs515_xor1;
  wire f_arrdiv24_fs515_not1;
  wire f_arrdiv24_fs515_and1;
  wire f_arrdiv24_fs515_or0;
  wire f_arrdiv24_fs516_xor0;
  wire f_arrdiv24_fs516_not0;
  wire f_arrdiv24_fs516_and0;
  wire f_arrdiv24_fs516_xor1;
  wire f_arrdiv24_fs516_not1;
  wire f_arrdiv24_fs516_and1;
  wire f_arrdiv24_fs516_or0;
  wire f_arrdiv24_fs517_xor0;
  wire f_arrdiv24_fs517_not0;
  wire f_arrdiv24_fs517_and0;
  wire f_arrdiv24_fs517_xor1;
  wire f_arrdiv24_fs517_not1;
  wire f_arrdiv24_fs517_and1;
  wire f_arrdiv24_fs517_or0;
  wire f_arrdiv24_fs518_xor0;
  wire f_arrdiv24_fs518_not0;
  wire f_arrdiv24_fs518_and0;
  wire f_arrdiv24_fs518_xor1;
  wire f_arrdiv24_fs518_not1;
  wire f_arrdiv24_fs518_and1;
  wire f_arrdiv24_fs518_or0;
  wire f_arrdiv24_fs519_xor0;
  wire f_arrdiv24_fs519_not0;
  wire f_arrdiv24_fs519_and0;
  wire f_arrdiv24_fs519_xor1;
  wire f_arrdiv24_fs519_not1;
  wire f_arrdiv24_fs519_and1;
  wire f_arrdiv24_fs519_or0;
  wire f_arrdiv24_fs520_xor0;
  wire f_arrdiv24_fs520_not0;
  wire f_arrdiv24_fs520_and0;
  wire f_arrdiv24_fs520_xor1;
  wire f_arrdiv24_fs520_not1;
  wire f_arrdiv24_fs520_and1;
  wire f_arrdiv24_fs520_or0;
  wire f_arrdiv24_fs521_xor0;
  wire f_arrdiv24_fs521_not0;
  wire f_arrdiv24_fs521_and0;
  wire f_arrdiv24_fs521_xor1;
  wire f_arrdiv24_fs521_not1;
  wire f_arrdiv24_fs521_and1;
  wire f_arrdiv24_fs521_or0;
  wire f_arrdiv24_fs522_xor0;
  wire f_arrdiv24_fs522_not0;
  wire f_arrdiv24_fs522_and0;
  wire f_arrdiv24_fs522_xor1;
  wire f_arrdiv24_fs522_not1;
  wire f_arrdiv24_fs522_and1;
  wire f_arrdiv24_fs522_or0;
  wire f_arrdiv24_fs523_xor0;
  wire f_arrdiv24_fs523_not0;
  wire f_arrdiv24_fs523_and0;
  wire f_arrdiv24_fs523_xor1;
  wire f_arrdiv24_fs523_not1;
  wire f_arrdiv24_fs523_and1;
  wire f_arrdiv24_fs523_or0;
  wire f_arrdiv24_fs524_xor0;
  wire f_arrdiv24_fs524_not0;
  wire f_arrdiv24_fs524_and0;
  wire f_arrdiv24_fs524_xor1;
  wire f_arrdiv24_fs524_not1;
  wire f_arrdiv24_fs524_and1;
  wire f_arrdiv24_fs524_or0;
  wire f_arrdiv24_fs525_xor0;
  wire f_arrdiv24_fs525_not0;
  wire f_arrdiv24_fs525_and0;
  wire f_arrdiv24_fs525_xor1;
  wire f_arrdiv24_fs525_not1;
  wire f_arrdiv24_fs525_and1;
  wire f_arrdiv24_fs525_or0;
  wire f_arrdiv24_fs526_xor0;
  wire f_arrdiv24_fs526_not0;
  wire f_arrdiv24_fs526_and0;
  wire f_arrdiv24_fs526_xor1;
  wire f_arrdiv24_fs526_not1;
  wire f_arrdiv24_fs526_and1;
  wire f_arrdiv24_fs526_or0;
  wire f_arrdiv24_fs527_xor0;
  wire f_arrdiv24_fs527_not0;
  wire f_arrdiv24_fs527_and0;
  wire f_arrdiv24_fs527_xor1;
  wire f_arrdiv24_fs527_not1;
  wire f_arrdiv24_fs527_and1;
  wire f_arrdiv24_fs527_or0;
  wire f_arrdiv24_mux2to1483_and0;
  wire f_arrdiv24_mux2to1483_not0;
  wire f_arrdiv24_mux2to1483_and1;
  wire f_arrdiv24_mux2to1483_xor0;
  wire f_arrdiv24_mux2to1484_and0;
  wire f_arrdiv24_mux2to1484_not0;
  wire f_arrdiv24_mux2to1484_and1;
  wire f_arrdiv24_mux2to1484_xor0;
  wire f_arrdiv24_mux2to1485_and0;
  wire f_arrdiv24_mux2to1485_not0;
  wire f_arrdiv24_mux2to1485_and1;
  wire f_arrdiv24_mux2to1485_xor0;
  wire f_arrdiv24_mux2to1486_and0;
  wire f_arrdiv24_mux2to1486_not0;
  wire f_arrdiv24_mux2to1486_and1;
  wire f_arrdiv24_mux2to1486_xor0;
  wire f_arrdiv24_mux2to1487_and0;
  wire f_arrdiv24_mux2to1487_not0;
  wire f_arrdiv24_mux2to1487_and1;
  wire f_arrdiv24_mux2to1487_xor0;
  wire f_arrdiv24_mux2to1488_and0;
  wire f_arrdiv24_mux2to1488_not0;
  wire f_arrdiv24_mux2to1488_and1;
  wire f_arrdiv24_mux2to1488_xor0;
  wire f_arrdiv24_mux2to1489_and0;
  wire f_arrdiv24_mux2to1489_not0;
  wire f_arrdiv24_mux2to1489_and1;
  wire f_arrdiv24_mux2to1489_xor0;
  wire f_arrdiv24_mux2to1490_and0;
  wire f_arrdiv24_mux2to1490_not0;
  wire f_arrdiv24_mux2to1490_and1;
  wire f_arrdiv24_mux2to1490_xor0;
  wire f_arrdiv24_mux2to1491_and0;
  wire f_arrdiv24_mux2to1491_not0;
  wire f_arrdiv24_mux2to1491_and1;
  wire f_arrdiv24_mux2to1491_xor0;
  wire f_arrdiv24_mux2to1492_and0;
  wire f_arrdiv24_mux2to1492_not0;
  wire f_arrdiv24_mux2to1492_and1;
  wire f_arrdiv24_mux2to1492_xor0;
  wire f_arrdiv24_mux2to1493_and0;
  wire f_arrdiv24_mux2to1493_not0;
  wire f_arrdiv24_mux2to1493_and1;
  wire f_arrdiv24_mux2to1493_xor0;
  wire f_arrdiv24_mux2to1494_and0;
  wire f_arrdiv24_mux2to1494_not0;
  wire f_arrdiv24_mux2to1494_and1;
  wire f_arrdiv24_mux2to1494_xor0;
  wire f_arrdiv24_mux2to1495_and0;
  wire f_arrdiv24_mux2to1495_not0;
  wire f_arrdiv24_mux2to1495_and1;
  wire f_arrdiv24_mux2to1495_xor0;
  wire f_arrdiv24_mux2to1496_and0;
  wire f_arrdiv24_mux2to1496_not0;
  wire f_arrdiv24_mux2to1496_and1;
  wire f_arrdiv24_mux2to1496_xor0;
  wire f_arrdiv24_mux2to1497_and0;
  wire f_arrdiv24_mux2to1497_not0;
  wire f_arrdiv24_mux2to1497_and1;
  wire f_arrdiv24_mux2to1497_xor0;
  wire f_arrdiv24_mux2to1498_and0;
  wire f_arrdiv24_mux2to1498_not0;
  wire f_arrdiv24_mux2to1498_and1;
  wire f_arrdiv24_mux2to1498_xor0;
  wire f_arrdiv24_mux2to1499_and0;
  wire f_arrdiv24_mux2to1499_not0;
  wire f_arrdiv24_mux2to1499_and1;
  wire f_arrdiv24_mux2to1499_xor0;
  wire f_arrdiv24_mux2to1500_and0;
  wire f_arrdiv24_mux2to1500_not0;
  wire f_arrdiv24_mux2to1500_and1;
  wire f_arrdiv24_mux2to1500_xor0;
  wire f_arrdiv24_mux2to1501_and0;
  wire f_arrdiv24_mux2to1501_not0;
  wire f_arrdiv24_mux2to1501_and1;
  wire f_arrdiv24_mux2to1501_xor0;
  wire f_arrdiv24_mux2to1502_and0;
  wire f_arrdiv24_mux2to1502_not0;
  wire f_arrdiv24_mux2to1502_and1;
  wire f_arrdiv24_mux2to1502_xor0;
  wire f_arrdiv24_mux2to1503_and0;
  wire f_arrdiv24_mux2to1503_not0;
  wire f_arrdiv24_mux2to1503_and1;
  wire f_arrdiv24_mux2to1503_xor0;
  wire f_arrdiv24_mux2to1504_and0;
  wire f_arrdiv24_mux2to1504_not0;
  wire f_arrdiv24_mux2to1504_and1;
  wire f_arrdiv24_mux2to1504_xor0;
  wire f_arrdiv24_mux2to1505_and0;
  wire f_arrdiv24_mux2to1505_not0;
  wire f_arrdiv24_mux2to1505_and1;
  wire f_arrdiv24_mux2to1505_xor0;
  wire f_arrdiv24_not21;
  wire f_arrdiv24_fs528_xor0;
  wire f_arrdiv24_fs528_not0;
  wire f_arrdiv24_fs528_and0;
  wire f_arrdiv24_fs528_not1;
  wire f_arrdiv24_fs529_xor0;
  wire f_arrdiv24_fs529_not0;
  wire f_arrdiv24_fs529_and0;
  wire f_arrdiv24_fs529_xor1;
  wire f_arrdiv24_fs529_not1;
  wire f_arrdiv24_fs529_and1;
  wire f_arrdiv24_fs529_or0;
  wire f_arrdiv24_fs530_xor0;
  wire f_arrdiv24_fs530_not0;
  wire f_arrdiv24_fs530_and0;
  wire f_arrdiv24_fs530_xor1;
  wire f_arrdiv24_fs530_not1;
  wire f_arrdiv24_fs530_and1;
  wire f_arrdiv24_fs530_or0;
  wire f_arrdiv24_fs531_xor0;
  wire f_arrdiv24_fs531_not0;
  wire f_arrdiv24_fs531_and0;
  wire f_arrdiv24_fs531_xor1;
  wire f_arrdiv24_fs531_not1;
  wire f_arrdiv24_fs531_and1;
  wire f_arrdiv24_fs531_or0;
  wire f_arrdiv24_fs532_xor0;
  wire f_arrdiv24_fs532_not0;
  wire f_arrdiv24_fs532_and0;
  wire f_arrdiv24_fs532_xor1;
  wire f_arrdiv24_fs532_not1;
  wire f_arrdiv24_fs532_and1;
  wire f_arrdiv24_fs532_or0;
  wire f_arrdiv24_fs533_xor0;
  wire f_arrdiv24_fs533_not0;
  wire f_arrdiv24_fs533_and0;
  wire f_arrdiv24_fs533_xor1;
  wire f_arrdiv24_fs533_not1;
  wire f_arrdiv24_fs533_and1;
  wire f_arrdiv24_fs533_or0;
  wire f_arrdiv24_fs534_xor0;
  wire f_arrdiv24_fs534_not0;
  wire f_arrdiv24_fs534_and0;
  wire f_arrdiv24_fs534_xor1;
  wire f_arrdiv24_fs534_not1;
  wire f_arrdiv24_fs534_and1;
  wire f_arrdiv24_fs534_or0;
  wire f_arrdiv24_fs535_xor0;
  wire f_arrdiv24_fs535_not0;
  wire f_arrdiv24_fs535_and0;
  wire f_arrdiv24_fs535_xor1;
  wire f_arrdiv24_fs535_not1;
  wire f_arrdiv24_fs535_and1;
  wire f_arrdiv24_fs535_or0;
  wire f_arrdiv24_fs536_xor0;
  wire f_arrdiv24_fs536_not0;
  wire f_arrdiv24_fs536_and0;
  wire f_arrdiv24_fs536_xor1;
  wire f_arrdiv24_fs536_not1;
  wire f_arrdiv24_fs536_and1;
  wire f_arrdiv24_fs536_or0;
  wire f_arrdiv24_fs537_xor0;
  wire f_arrdiv24_fs537_not0;
  wire f_arrdiv24_fs537_and0;
  wire f_arrdiv24_fs537_xor1;
  wire f_arrdiv24_fs537_not1;
  wire f_arrdiv24_fs537_and1;
  wire f_arrdiv24_fs537_or0;
  wire f_arrdiv24_fs538_xor0;
  wire f_arrdiv24_fs538_not0;
  wire f_arrdiv24_fs538_and0;
  wire f_arrdiv24_fs538_xor1;
  wire f_arrdiv24_fs538_not1;
  wire f_arrdiv24_fs538_and1;
  wire f_arrdiv24_fs538_or0;
  wire f_arrdiv24_fs539_xor0;
  wire f_arrdiv24_fs539_not0;
  wire f_arrdiv24_fs539_and0;
  wire f_arrdiv24_fs539_xor1;
  wire f_arrdiv24_fs539_not1;
  wire f_arrdiv24_fs539_and1;
  wire f_arrdiv24_fs539_or0;
  wire f_arrdiv24_fs540_xor0;
  wire f_arrdiv24_fs540_not0;
  wire f_arrdiv24_fs540_and0;
  wire f_arrdiv24_fs540_xor1;
  wire f_arrdiv24_fs540_not1;
  wire f_arrdiv24_fs540_and1;
  wire f_arrdiv24_fs540_or0;
  wire f_arrdiv24_fs541_xor0;
  wire f_arrdiv24_fs541_not0;
  wire f_arrdiv24_fs541_and0;
  wire f_arrdiv24_fs541_xor1;
  wire f_arrdiv24_fs541_not1;
  wire f_arrdiv24_fs541_and1;
  wire f_arrdiv24_fs541_or0;
  wire f_arrdiv24_fs542_xor0;
  wire f_arrdiv24_fs542_not0;
  wire f_arrdiv24_fs542_and0;
  wire f_arrdiv24_fs542_xor1;
  wire f_arrdiv24_fs542_not1;
  wire f_arrdiv24_fs542_and1;
  wire f_arrdiv24_fs542_or0;
  wire f_arrdiv24_fs543_xor0;
  wire f_arrdiv24_fs543_not0;
  wire f_arrdiv24_fs543_and0;
  wire f_arrdiv24_fs543_xor1;
  wire f_arrdiv24_fs543_not1;
  wire f_arrdiv24_fs543_and1;
  wire f_arrdiv24_fs543_or0;
  wire f_arrdiv24_fs544_xor0;
  wire f_arrdiv24_fs544_not0;
  wire f_arrdiv24_fs544_and0;
  wire f_arrdiv24_fs544_xor1;
  wire f_arrdiv24_fs544_not1;
  wire f_arrdiv24_fs544_and1;
  wire f_arrdiv24_fs544_or0;
  wire f_arrdiv24_fs545_xor0;
  wire f_arrdiv24_fs545_not0;
  wire f_arrdiv24_fs545_and0;
  wire f_arrdiv24_fs545_xor1;
  wire f_arrdiv24_fs545_not1;
  wire f_arrdiv24_fs545_and1;
  wire f_arrdiv24_fs545_or0;
  wire f_arrdiv24_fs546_xor0;
  wire f_arrdiv24_fs546_not0;
  wire f_arrdiv24_fs546_and0;
  wire f_arrdiv24_fs546_xor1;
  wire f_arrdiv24_fs546_not1;
  wire f_arrdiv24_fs546_and1;
  wire f_arrdiv24_fs546_or0;
  wire f_arrdiv24_fs547_xor0;
  wire f_arrdiv24_fs547_not0;
  wire f_arrdiv24_fs547_and0;
  wire f_arrdiv24_fs547_xor1;
  wire f_arrdiv24_fs547_not1;
  wire f_arrdiv24_fs547_and1;
  wire f_arrdiv24_fs547_or0;
  wire f_arrdiv24_fs548_xor0;
  wire f_arrdiv24_fs548_not0;
  wire f_arrdiv24_fs548_and0;
  wire f_arrdiv24_fs548_xor1;
  wire f_arrdiv24_fs548_not1;
  wire f_arrdiv24_fs548_and1;
  wire f_arrdiv24_fs548_or0;
  wire f_arrdiv24_fs549_xor0;
  wire f_arrdiv24_fs549_not0;
  wire f_arrdiv24_fs549_and0;
  wire f_arrdiv24_fs549_xor1;
  wire f_arrdiv24_fs549_not1;
  wire f_arrdiv24_fs549_and1;
  wire f_arrdiv24_fs549_or0;
  wire f_arrdiv24_fs550_xor0;
  wire f_arrdiv24_fs550_not0;
  wire f_arrdiv24_fs550_and0;
  wire f_arrdiv24_fs550_xor1;
  wire f_arrdiv24_fs550_not1;
  wire f_arrdiv24_fs550_and1;
  wire f_arrdiv24_fs550_or0;
  wire f_arrdiv24_fs551_xor0;
  wire f_arrdiv24_fs551_not0;
  wire f_arrdiv24_fs551_and0;
  wire f_arrdiv24_fs551_xor1;
  wire f_arrdiv24_fs551_not1;
  wire f_arrdiv24_fs551_and1;
  wire f_arrdiv24_fs551_or0;
  wire f_arrdiv24_mux2to1506_and0;
  wire f_arrdiv24_mux2to1506_not0;
  wire f_arrdiv24_mux2to1506_and1;
  wire f_arrdiv24_mux2to1506_xor0;
  wire f_arrdiv24_mux2to1507_and0;
  wire f_arrdiv24_mux2to1507_not0;
  wire f_arrdiv24_mux2to1507_and1;
  wire f_arrdiv24_mux2to1507_xor0;
  wire f_arrdiv24_mux2to1508_and0;
  wire f_arrdiv24_mux2to1508_not0;
  wire f_arrdiv24_mux2to1508_and1;
  wire f_arrdiv24_mux2to1508_xor0;
  wire f_arrdiv24_mux2to1509_and0;
  wire f_arrdiv24_mux2to1509_not0;
  wire f_arrdiv24_mux2to1509_and1;
  wire f_arrdiv24_mux2to1509_xor0;
  wire f_arrdiv24_mux2to1510_and0;
  wire f_arrdiv24_mux2to1510_not0;
  wire f_arrdiv24_mux2to1510_and1;
  wire f_arrdiv24_mux2to1510_xor0;
  wire f_arrdiv24_mux2to1511_and0;
  wire f_arrdiv24_mux2to1511_not0;
  wire f_arrdiv24_mux2to1511_and1;
  wire f_arrdiv24_mux2to1511_xor0;
  wire f_arrdiv24_mux2to1512_and0;
  wire f_arrdiv24_mux2to1512_not0;
  wire f_arrdiv24_mux2to1512_and1;
  wire f_arrdiv24_mux2to1512_xor0;
  wire f_arrdiv24_mux2to1513_and0;
  wire f_arrdiv24_mux2to1513_not0;
  wire f_arrdiv24_mux2to1513_and1;
  wire f_arrdiv24_mux2to1513_xor0;
  wire f_arrdiv24_mux2to1514_and0;
  wire f_arrdiv24_mux2to1514_not0;
  wire f_arrdiv24_mux2to1514_and1;
  wire f_arrdiv24_mux2to1514_xor0;
  wire f_arrdiv24_mux2to1515_and0;
  wire f_arrdiv24_mux2to1515_not0;
  wire f_arrdiv24_mux2to1515_and1;
  wire f_arrdiv24_mux2to1515_xor0;
  wire f_arrdiv24_mux2to1516_and0;
  wire f_arrdiv24_mux2to1516_not0;
  wire f_arrdiv24_mux2to1516_and1;
  wire f_arrdiv24_mux2to1516_xor0;
  wire f_arrdiv24_mux2to1517_and0;
  wire f_arrdiv24_mux2to1517_not0;
  wire f_arrdiv24_mux2to1517_and1;
  wire f_arrdiv24_mux2to1517_xor0;
  wire f_arrdiv24_mux2to1518_and0;
  wire f_arrdiv24_mux2to1518_not0;
  wire f_arrdiv24_mux2to1518_and1;
  wire f_arrdiv24_mux2to1518_xor0;
  wire f_arrdiv24_mux2to1519_and0;
  wire f_arrdiv24_mux2to1519_not0;
  wire f_arrdiv24_mux2to1519_and1;
  wire f_arrdiv24_mux2to1519_xor0;
  wire f_arrdiv24_mux2to1520_and0;
  wire f_arrdiv24_mux2to1520_not0;
  wire f_arrdiv24_mux2to1520_and1;
  wire f_arrdiv24_mux2to1520_xor0;
  wire f_arrdiv24_mux2to1521_and0;
  wire f_arrdiv24_mux2to1521_not0;
  wire f_arrdiv24_mux2to1521_and1;
  wire f_arrdiv24_mux2to1521_xor0;
  wire f_arrdiv24_mux2to1522_and0;
  wire f_arrdiv24_mux2to1522_not0;
  wire f_arrdiv24_mux2to1522_and1;
  wire f_arrdiv24_mux2to1522_xor0;
  wire f_arrdiv24_mux2to1523_and0;
  wire f_arrdiv24_mux2to1523_not0;
  wire f_arrdiv24_mux2to1523_and1;
  wire f_arrdiv24_mux2to1523_xor0;
  wire f_arrdiv24_mux2to1524_and0;
  wire f_arrdiv24_mux2to1524_not0;
  wire f_arrdiv24_mux2to1524_and1;
  wire f_arrdiv24_mux2to1524_xor0;
  wire f_arrdiv24_mux2to1525_and0;
  wire f_arrdiv24_mux2to1525_not0;
  wire f_arrdiv24_mux2to1525_and1;
  wire f_arrdiv24_mux2to1525_xor0;
  wire f_arrdiv24_mux2to1526_and0;
  wire f_arrdiv24_mux2to1526_not0;
  wire f_arrdiv24_mux2to1526_and1;
  wire f_arrdiv24_mux2to1526_xor0;
  wire f_arrdiv24_mux2to1527_and0;
  wire f_arrdiv24_mux2to1527_not0;
  wire f_arrdiv24_mux2to1527_and1;
  wire f_arrdiv24_mux2to1527_xor0;
  wire f_arrdiv24_mux2to1528_and0;
  wire f_arrdiv24_mux2to1528_not0;
  wire f_arrdiv24_mux2to1528_and1;
  wire f_arrdiv24_mux2to1528_xor0;
  wire f_arrdiv24_not22;
  wire f_arrdiv24_fs552_xor0;
  wire f_arrdiv24_fs552_not0;
  wire f_arrdiv24_fs552_and0;
  wire f_arrdiv24_fs552_not1;
  wire f_arrdiv24_fs553_xor0;
  wire f_arrdiv24_fs553_not0;
  wire f_arrdiv24_fs553_and0;
  wire f_arrdiv24_fs553_xor1;
  wire f_arrdiv24_fs553_not1;
  wire f_arrdiv24_fs553_and1;
  wire f_arrdiv24_fs553_or0;
  wire f_arrdiv24_fs554_xor0;
  wire f_arrdiv24_fs554_not0;
  wire f_arrdiv24_fs554_and0;
  wire f_arrdiv24_fs554_xor1;
  wire f_arrdiv24_fs554_not1;
  wire f_arrdiv24_fs554_and1;
  wire f_arrdiv24_fs554_or0;
  wire f_arrdiv24_fs555_xor0;
  wire f_arrdiv24_fs555_not0;
  wire f_arrdiv24_fs555_and0;
  wire f_arrdiv24_fs555_xor1;
  wire f_arrdiv24_fs555_not1;
  wire f_arrdiv24_fs555_and1;
  wire f_arrdiv24_fs555_or0;
  wire f_arrdiv24_fs556_xor0;
  wire f_arrdiv24_fs556_not0;
  wire f_arrdiv24_fs556_and0;
  wire f_arrdiv24_fs556_xor1;
  wire f_arrdiv24_fs556_not1;
  wire f_arrdiv24_fs556_and1;
  wire f_arrdiv24_fs556_or0;
  wire f_arrdiv24_fs557_xor0;
  wire f_arrdiv24_fs557_not0;
  wire f_arrdiv24_fs557_and0;
  wire f_arrdiv24_fs557_xor1;
  wire f_arrdiv24_fs557_not1;
  wire f_arrdiv24_fs557_and1;
  wire f_arrdiv24_fs557_or0;
  wire f_arrdiv24_fs558_xor0;
  wire f_arrdiv24_fs558_not0;
  wire f_arrdiv24_fs558_and0;
  wire f_arrdiv24_fs558_xor1;
  wire f_arrdiv24_fs558_not1;
  wire f_arrdiv24_fs558_and1;
  wire f_arrdiv24_fs558_or0;
  wire f_arrdiv24_fs559_xor0;
  wire f_arrdiv24_fs559_not0;
  wire f_arrdiv24_fs559_and0;
  wire f_arrdiv24_fs559_xor1;
  wire f_arrdiv24_fs559_not1;
  wire f_arrdiv24_fs559_and1;
  wire f_arrdiv24_fs559_or0;
  wire f_arrdiv24_fs560_xor0;
  wire f_arrdiv24_fs560_not0;
  wire f_arrdiv24_fs560_and0;
  wire f_arrdiv24_fs560_xor1;
  wire f_arrdiv24_fs560_not1;
  wire f_arrdiv24_fs560_and1;
  wire f_arrdiv24_fs560_or0;
  wire f_arrdiv24_fs561_xor0;
  wire f_arrdiv24_fs561_not0;
  wire f_arrdiv24_fs561_and0;
  wire f_arrdiv24_fs561_xor1;
  wire f_arrdiv24_fs561_not1;
  wire f_arrdiv24_fs561_and1;
  wire f_arrdiv24_fs561_or0;
  wire f_arrdiv24_fs562_xor0;
  wire f_arrdiv24_fs562_not0;
  wire f_arrdiv24_fs562_and0;
  wire f_arrdiv24_fs562_xor1;
  wire f_arrdiv24_fs562_not1;
  wire f_arrdiv24_fs562_and1;
  wire f_arrdiv24_fs562_or0;
  wire f_arrdiv24_fs563_xor0;
  wire f_arrdiv24_fs563_not0;
  wire f_arrdiv24_fs563_and0;
  wire f_arrdiv24_fs563_xor1;
  wire f_arrdiv24_fs563_not1;
  wire f_arrdiv24_fs563_and1;
  wire f_arrdiv24_fs563_or0;
  wire f_arrdiv24_fs564_xor0;
  wire f_arrdiv24_fs564_not0;
  wire f_arrdiv24_fs564_and0;
  wire f_arrdiv24_fs564_xor1;
  wire f_arrdiv24_fs564_not1;
  wire f_arrdiv24_fs564_and1;
  wire f_arrdiv24_fs564_or0;
  wire f_arrdiv24_fs565_xor0;
  wire f_arrdiv24_fs565_not0;
  wire f_arrdiv24_fs565_and0;
  wire f_arrdiv24_fs565_xor1;
  wire f_arrdiv24_fs565_not1;
  wire f_arrdiv24_fs565_and1;
  wire f_arrdiv24_fs565_or0;
  wire f_arrdiv24_fs566_xor0;
  wire f_arrdiv24_fs566_not0;
  wire f_arrdiv24_fs566_and0;
  wire f_arrdiv24_fs566_xor1;
  wire f_arrdiv24_fs566_not1;
  wire f_arrdiv24_fs566_and1;
  wire f_arrdiv24_fs566_or0;
  wire f_arrdiv24_fs567_xor0;
  wire f_arrdiv24_fs567_not0;
  wire f_arrdiv24_fs567_and0;
  wire f_arrdiv24_fs567_xor1;
  wire f_arrdiv24_fs567_not1;
  wire f_arrdiv24_fs567_and1;
  wire f_arrdiv24_fs567_or0;
  wire f_arrdiv24_fs568_xor0;
  wire f_arrdiv24_fs568_not0;
  wire f_arrdiv24_fs568_and0;
  wire f_arrdiv24_fs568_xor1;
  wire f_arrdiv24_fs568_not1;
  wire f_arrdiv24_fs568_and1;
  wire f_arrdiv24_fs568_or0;
  wire f_arrdiv24_fs569_xor0;
  wire f_arrdiv24_fs569_not0;
  wire f_arrdiv24_fs569_and0;
  wire f_arrdiv24_fs569_xor1;
  wire f_arrdiv24_fs569_not1;
  wire f_arrdiv24_fs569_and1;
  wire f_arrdiv24_fs569_or0;
  wire f_arrdiv24_fs570_xor0;
  wire f_arrdiv24_fs570_not0;
  wire f_arrdiv24_fs570_and0;
  wire f_arrdiv24_fs570_xor1;
  wire f_arrdiv24_fs570_not1;
  wire f_arrdiv24_fs570_and1;
  wire f_arrdiv24_fs570_or0;
  wire f_arrdiv24_fs571_xor0;
  wire f_arrdiv24_fs571_not0;
  wire f_arrdiv24_fs571_and0;
  wire f_arrdiv24_fs571_xor1;
  wire f_arrdiv24_fs571_not1;
  wire f_arrdiv24_fs571_and1;
  wire f_arrdiv24_fs571_or0;
  wire f_arrdiv24_fs572_xor0;
  wire f_arrdiv24_fs572_not0;
  wire f_arrdiv24_fs572_and0;
  wire f_arrdiv24_fs572_xor1;
  wire f_arrdiv24_fs572_not1;
  wire f_arrdiv24_fs572_and1;
  wire f_arrdiv24_fs572_or0;
  wire f_arrdiv24_fs573_xor0;
  wire f_arrdiv24_fs573_not0;
  wire f_arrdiv24_fs573_and0;
  wire f_arrdiv24_fs573_xor1;
  wire f_arrdiv24_fs573_not1;
  wire f_arrdiv24_fs573_and1;
  wire f_arrdiv24_fs573_or0;
  wire f_arrdiv24_fs574_xor0;
  wire f_arrdiv24_fs574_not0;
  wire f_arrdiv24_fs574_and0;
  wire f_arrdiv24_fs574_xor1;
  wire f_arrdiv24_fs574_not1;
  wire f_arrdiv24_fs574_and1;
  wire f_arrdiv24_fs574_or0;
  wire f_arrdiv24_fs575_xor0;
  wire f_arrdiv24_fs575_not0;
  wire f_arrdiv24_fs575_and0;
  wire f_arrdiv24_fs575_xor1;
  wire f_arrdiv24_fs575_not1;
  wire f_arrdiv24_fs575_and1;
  wire f_arrdiv24_fs575_or0;
  wire f_arrdiv24_not23;

  assign f_arrdiv24_fs0_xor0 = a[23] ^ b[0];
  assign f_arrdiv24_fs0_not0 = ~a[23];
  assign f_arrdiv24_fs0_and0 = f_arrdiv24_fs0_not0 & b[0];
  assign f_arrdiv24_fs0_not1 = ~f_arrdiv24_fs0_xor0;
  assign f_arrdiv24_fs1_xor1 = f_arrdiv24_fs0_and0 ^ b[1];
  assign f_arrdiv24_fs1_not1 = ~b[1];
  assign f_arrdiv24_fs1_and1 = f_arrdiv24_fs1_not1 & f_arrdiv24_fs0_and0;
  assign f_arrdiv24_fs1_or0 = f_arrdiv24_fs1_and1 | b[1];
  assign f_arrdiv24_fs2_xor1 = f_arrdiv24_fs1_or0 ^ b[2];
  assign f_arrdiv24_fs2_not1 = ~b[2];
  assign f_arrdiv24_fs2_and1 = f_arrdiv24_fs2_not1 & f_arrdiv24_fs1_or0;
  assign f_arrdiv24_fs2_or0 = f_arrdiv24_fs2_and1 | b[2];
  assign f_arrdiv24_fs3_xor1 = f_arrdiv24_fs2_or0 ^ b[3];
  assign f_arrdiv24_fs3_not1 = ~b[3];
  assign f_arrdiv24_fs3_and1 = f_arrdiv24_fs3_not1 & f_arrdiv24_fs2_or0;
  assign f_arrdiv24_fs3_or0 = f_arrdiv24_fs3_and1 | b[3];
  assign f_arrdiv24_fs4_xor1 = f_arrdiv24_fs3_or0 ^ b[4];
  assign f_arrdiv24_fs4_not1 = ~b[4];
  assign f_arrdiv24_fs4_and1 = f_arrdiv24_fs4_not1 & f_arrdiv24_fs3_or0;
  assign f_arrdiv24_fs4_or0 = f_arrdiv24_fs4_and1 | b[4];
  assign f_arrdiv24_fs5_xor1 = f_arrdiv24_fs4_or0 ^ b[5];
  assign f_arrdiv24_fs5_not1 = ~b[5];
  assign f_arrdiv24_fs5_and1 = f_arrdiv24_fs5_not1 & f_arrdiv24_fs4_or0;
  assign f_arrdiv24_fs5_or0 = f_arrdiv24_fs5_and1 | b[5];
  assign f_arrdiv24_fs6_xor1 = f_arrdiv24_fs5_or0 ^ b[6];
  assign f_arrdiv24_fs6_not1 = ~b[6];
  assign f_arrdiv24_fs6_and1 = f_arrdiv24_fs6_not1 & f_arrdiv24_fs5_or0;
  assign f_arrdiv24_fs6_or0 = f_arrdiv24_fs6_and1 | b[6];
  assign f_arrdiv24_fs7_xor1 = f_arrdiv24_fs6_or0 ^ b[7];
  assign f_arrdiv24_fs7_not1 = ~b[7];
  assign f_arrdiv24_fs7_and1 = f_arrdiv24_fs7_not1 & f_arrdiv24_fs6_or0;
  assign f_arrdiv24_fs7_or0 = f_arrdiv24_fs7_and1 | b[7];
  assign f_arrdiv24_fs8_xor1 = f_arrdiv24_fs7_or0 ^ b[8];
  assign f_arrdiv24_fs8_not1 = ~b[8];
  assign f_arrdiv24_fs8_and1 = f_arrdiv24_fs8_not1 & f_arrdiv24_fs7_or0;
  assign f_arrdiv24_fs8_or0 = f_arrdiv24_fs8_and1 | b[8];
  assign f_arrdiv24_fs9_xor1 = f_arrdiv24_fs8_or0 ^ b[9];
  assign f_arrdiv24_fs9_not1 = ~b[9];
  assign f_arrdiv24_fs9_and1 = f_arrdiv24_fs9_not1 & f_arrdiv24_fs8_or0;
  assign f_arrdiv24_fs9_or0 = f_arrdiv24_fs9_and1 | b[9];
  assign f_arrdiv24_fs10_xor1 = f_arrdiv24_fs9_or0 ^ b[10];
  assign f_arrdiv24_fs10_not1 = ~b[10];
  assign f_arrdiv24_fs10_and1 = f_arrdiv24_fs10_not1 & f_arrdiv24_fs9_or0;
  assign f_arrdiv24_fs10_or0 = f_arrdiv24_fs10_and1 | b[10];
  assign f_arrdiv24_fs11_xor1 = f_arrdiv24_fs10_or0 ^ b[11];
  assign f_arrdiv24_fs11_not1 = ~b[11];
  assign f_arrdiv24_fs11_and1 = f_arrdiv24_fs11_not1 & f_arrdiv24_fs10_or0;
  assign f_arrdiv24_fs11_or0 = f_arrdiv24_fs11_and1 | b[11];
  assign f_arrdiv24_fs12_xor1 = f_arrdiv24_fs11_or0 ^ b[12];
  assign f_arrdiv24_fs12_not1 = ~b[12];
  assign f_arrdiv24_fs12_and1 = f_arrdiv24_fs12_not1 & f_arrdiv24_fs11_or0;
  assign f_arrdiv24_fs12_or0 = f_arrdiv24_fs12_and1 | b[12];
  assign f_arrdiv24_fs13_xor1 = f_arrdiv24_fs12_or0 ^ b[13];
  assign f_arrdiv24_fs13_not1 = ~b[13];
  assign f_arrdiv24_fs13_and1 = f_arrdiv24_fs13_not1 & f_arrdiv24_fs12_or0;
  assign f_arrdiv24_fs13_or0 = f_arrdiv24_fs13_and1 | b[13];
  assign f_arrdiv24_fs14_xor1 = f_arrdiv24_fs13_or0 ^ b[14];
  assign f_arrdiv24_fs14_not1 = ~b[14];
  assign f_arrdiv24_fs14_and1 = f_arrdiv24_fs14_not1 & f_arrdiv24_fs13_or0;
  assign f_arrdiv24_fs14_or0 = f_arrdiv24_fs14_and1 | b[14];
  assign f_arrdiv24_fs15_xor1 = f_arrdiv24_fs14_or0 ^ b[15];
  assign f_arrdiv24_fs15_not1 = ~b[15];
  assign f_arrdiv24_fs15_and1 = f_arrdiv24_fs15_not1 & f_arrdiv24_fs14_or0;
  assign f_arrdiv24_fs15_or0 = f_arrdiv24_fs15_and1 | b[15];
  assign f_arrdiv24_fs16_xor1 = f_arrdiv24_fs15_or0 ^ b[16];
  assign f_arrdiv24_fs16_not1 = ~b[16];
  assign f_arrdiv24_fs16_and1 = f_arrdiv24_fs16_not1 & f_arrdiv24_fs15_or0;
  assign f_arrdiv24_fs16_or0 = f_arrdiv24_fs16_and1 | b[16];
  assign f_arrdiv24_fs17_xor1 = f_arrdiv24_fs16_or0 ^ b[17];
  assign f_arrdiv24_fs17_not1 = ~b[17];
  assign f_arrdiv24_fs17_and1 = f_arrdiv24_fs17_not1 & f_arrdiv24_fs16_or0;
  assign f_arrdiv24_fs17_or0 = f_arrdiv24_fs17_and1 | b[17];
  assign f_arrdiv24_fs18_xor1 = f_arrdiv24_fs17_or0 ^ b[18];
  assign f_arrdiv24_fs18_not1 = ~b[18];
  assign f_arrdiv24_fs18_and1 = f_arrdiv24_fs18_not1 & f_arrdiv24_fs17_or0;
  assign f_arrdiv24_fs18_or0 = f_arrdiv24_fs18_and1 | b[18];
  assign f_arrdiv24_fs19_xor1 = f_arrdiv24_fs18_or0 ^ b[19];
  assign f_arrdiv24_fs19_not1 = ~b[19];
  assign f_arrdiv24_fs19_and1 = f_arrdiv24_fs19_not1 & f_arrdiv24_fs18_or0;
  assign f_arrdiv24_fs19_or0 = f_arrdiv24_fs19_and1 | b[19];
  assign f_arrdiv24_fs20_xor1 = f_arrdiv24_fs19_or0 ^ b[20];
  assign f_arrdiv24_fs20_not1 = ~b[20];
  assign f_arrdiv24_fs20_and1 = f_arrdiv24_fs20_not1 & f_arrdiv24_fs19_or0;
  assign f_arrdiv24_fs20_or0 = f_arrdiv24_fs20_and1 | b[20];
  assign f_arrdiv24_fs21_xor1 = f_arrdiv24_fs20_or0 ^ b[21];
  assign f_arrdiv24_fs21_not1 = ~b[21];
  assign f_arrdiv24_fs21_and1 = f_arrdiv24_fs21_not1 & f_arrdiv24_fs20_or0;
  assign f_arrdiv24_fs21_or0 = f_arrdiv24_fs21_and1 | b[21];
  assign f_arrdiv24_fs22_xor1 = f_arrdiv24_fs21_or0 ^ b[22];
  assign f_arrdiv24_fs22_not1 = ~b[22];
  assign f_arrdiv24_fs22_and1 = f_arrdiv24_fs22_not1 & f_arrdiv24_fs21_or0;
  assign f_arrdiv24_fs22_or0 = f_arrdiv24_fs22_and1 | b[22];
  assign f_arrdiv24_fs23_xor1 = f_arrdiv24_fs22_or0 ^ b[23];
  assign f_arrdiv24_fs23_not1 = ~b[23];
  assign f_arrdiv24_fs23_and1 = f_arrdiv24_fs23_not1 & f_arrdiv24_fs22_or0;
  assign f_arrdiv24_fs23_or0 = f_arrdiv24_fs23_and1 | b[23];
  assign f_arrdiv24_mux2to10_and0 = a[23] & f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to10_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to10_and1 = f_arrdiv24_fs0_xor0 & f_arrdiv24_mux2to10_not0;
  assign f_arrdiv24_mux2to10_xor0 = f_arrdiv24_mux2to10_and0 ^ f_arrdiv24_mux2to10_and1;
  assign f_arrdiv24_mux2to11_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to11_and1 = f_arrdiv24_fs1_xor1 & f_arrdiv24_mux2to11_not0;
  assign f_arrdiv24_mux2to12_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to12_and1 = f_arrdiv24_fs2_xor1 & f_arrdiv24_mux2to12_not0;
  assign f_arrdiv24_mux2to13_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to13_and1 = f_arrdiv24_fs3_xor1 & f_arrdiv24_mux2to13_not0;
  assign f_arrdiv24_mux2to14_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to14_and1 = f_arrdiv24_fs4_xor1 & f_arrdiv24_mux2to14_not0;
  assign f_arrdiv24_mux2to15_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to15_and1 = f_arrdiv24_fs5_xor1 & f_arrdiv24_mux2to15_not0;
  assign f_arrdiv24_mux2to16_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to16_and1 = f_arrdiv24_fs6_xor1 & f_arrdiv24_mux2to16_not0;
  assign f_arrdiv24_mux2to17_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to17_and1 = f_arrdiv24_fs7_xor1 & f_arrdiv24_mux2to17_not0;
  assign f_arrdiv24_mux2to18_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to18_and1 = f_arrdiv24_fs8_xor1 & f_arrdiv24_mux2to18_not0;
  assign f_arrdiv24_mux2to19_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to19_and1 = f_arrdiv24_fs9_xor1 & f_arrdiv24_mux2to19_not0;
  assign f_arrdiv24_mux2to110_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to110_and1 = f_arrdiv24_fs10_xor1 & f_arrdiv24_mux2to110_not0;
  assign f_arrdiv24_mux2to111_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to111_and1 = f_arrdiv24_fs11_xor1 & f_arrdiv24_mux2to111_not0;
  assign f_arrdiv24_mux2to112_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to112_and1 = f_arrdiv24_fs12_xor1 & f_arrdiv24_mux2to112_not0;
  assign f_arrdiv24_mux2to113_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to113_and1 = f_arrdiv24_fs13_xor1 & f_arrdiv24_mux2to113_not0;
  assign f_arrdiv24_mux2to114_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to114_and1 = f_arrdiv24_fs14_xor1 & f_arrdiv24_mux2to114_not0;
  assign f_arrdiv24_mux2to115_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to115_and1 = f_arrdiv24_fs15_xor1 & f_arrdiv24_mux2to115_not0;
  assign f_arrdiv24_mux2to116_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to116_and1 = f_arrdiv24_fs16_xor1 & f_arrdiv24_mux2to116_not0;
  assign f_arrdiv24_mux2to117_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to117_and1 = f_arrdiv24_fs17_xor1 & f_arrdiv24_mux2to117_not0;
  assign f_arrdiv24_mux2to118_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to118_and1 = f_arrdiv24_fs18_xor1 & f_arrdiv24_mux2to118_not0;
  assign f_arrdiv24_mux2to119_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to119_and1 = f_arrdiv24_fs19_xor1 & f_arrdiv24_mux2to119_not0;
  assign f_arrdiv24_mux2to120_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to120_and1 = f_arrdiv24_fs20_xor1 & f_arrdiv24_mux2to120_not0;
  assign f_arrdiv24_mux2to121_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to121_and1 = f_arrdiv24_fs21_xor1 & f_arrdiv24_mux2to121_not0;
  assign f_arrdiv24_mux2to122_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_mux2to122_and1 = f_arrdiv24_fs22_xor1 & f_arrdiv24_mux2to122_not0;
  assign f_arrdiv24_not0 = ~f_arrdiv24_fs23_or0;
  assign f_arrdiv24_fs24_xor0 = a[22] ^ b[0];
  assign f_arrdiv24_fs24_not0 = ~a[22];
  assign f_arrdiv24_fs24_and0 = f_arrdiv24_fs24_not0 & b[0];
  assign f_arrdiv24_fs24_not1 = ~f_arrdiv24_fs24_xor0;
  assign f_arrdiv24_fs25_xor0 = f_arrdiv24_mux2to10_xor0 ^ b[1];
  assign f_arrdiv24_fs25_not0 = ~f_arrdiv24_mux2to10_xor0;
  assign f_arrdiv24_fs25_and0 = f_arrdiv24_fs25_not0 & b[1];
  assign f_arrdiv24_fs25_xor1 = f_arrdiv24_fs24_and0 ^ f_arrdiv24_fs25_xor0;
  assign f_arrdiv24_fs25_not1 = ~f_arrdiv24_fs25_xor0;
  assign f_arrdiv24_fs25_and1 = f_arrdiv24_fs25_not1 & f_arrdiv24_fs24_and0;
  assign f_arrdiv24_fs25_or0 = f_arrdiv24_fs25_and1 | f_arrdiv24_fs25_and0;
  assign f_arrdiv24_fs26_xor0 = f_arrdiv24_mux2to11_and1 ^ b[2];
  assign f_arrdiv24_fs26_not0 = ~f_arrdiv24_mux2to11_and1;
  assign f_arrdiv24_fs26_and0 = f_arrdiv24_fs26_not0 & b[2];
  assign f_arrdiv24_fs26_xor1 = f_arrdiv24_fs25_or0 ^ f_arrdiv24_fs26_xor0;
  assign f_arrdiv24_fs26_not1 = ~f_arrdiv24_fs26_xor0;
  assign f_arrdiv24_fs26_and1 = f_arrdiv24_fs26_not1 & f_arrdiv24_fs25_or0;
  assign f_arrdiv24_fs26_or0 = f_arrdiv24_fs26_and1 | f_arrdiv24_fs26_and0;
  assign f_arrdiv24_fs27_xor0 = f_arrdiv24_mux2to12_and1 ^ b[3];
  assign f_arrdiv24_fs27_not0 = ~f_arrdiv24_mux2to12_and1;
  assign f_arrdiv24_fs27_and0 = f_arrdiv24_fs27_not0 & b[3];
  assign f_arrdiv24_fs27_xor1 = f_arrdiv24_fs26_or0 ^ f_arrdiv24_fs27_xor0;
  assign f_arrdiv24_fs27_not1 = ~f_arrdiv24_fs27_xor0;
  assign f_arrdiv24_fs27_and1 = f_arrdiv24_fs27_not1 & f_arrdiv24_fs26_or0;
  assign f_arrdiv24_fs27_or0 = f_arrdiv24_fs27_and1 | f_arrdiv24_fs27_and0;
  assign f_arrdiv24_fs28_xor0 = f_arrdiv24_mux2to13_and1 ^ b[4];
  assign f_arrdiv24_fs28_not0 = ~f_arrdiv24_mux2to13_and1;
  assign f_arrdiv24_fs28_and0 = f_arrdiv24_fs28_not0 & b[4];
  assign f_arrdiv24_fs28_xor1 = f_arrdiv24_fs27_or0 ^ f_arrdiv24_fs28_xor0;
  assign f_arrdiv24_fs28_not1 = ~f_arrdiv24_fs28_xor0;
  assign f_arrdiv24_fs28_and1 = f_arrdiv24_fs28_not1 & f_arrdiv24_fs27_or0;
  assign f_arrdiv24_fs28_or0 = f_arrdiv24_fs28_and1 | f_arrdiv24_fs28_and0;
  assign f_arrdiv24_fs29_xor0 = f_arrdiv24_mux2to14_and1 ^ b[5];
  assign f_arrdiv24_fs29_not0 = ~f_arrdiv24_mux2to14_and1;
  assign f_arrdiv24_fs29_and0 = f_arrdiv24_fs29_not0 & b[5];
  assign f_arrdiv24_fs29_xor1 = f_arrdiv24_fs28_or0 ^ f_arrdiv24_fs29_xor0;
  assign f_arrdiv24_fs29_not1 = ~f_arrdiv24_fs29_xor0;
  assign f_arrdiv24_fs29_and1 = f_arrdiv24_fs29_not1 & f_arrdiv24_fs28_or0;
  assign f_arrdiv24_fs29_or0 = f_arrdiv24_fs29_and1 | f_arrdiv24_fs29_and0;
  assign f_arrdiv24_fs30_xor0 = f_arrdiv24_mux2to15_and1 ^ b[6];
  assign f_arrdiv24_fs30_not0 = ~f_arrdiv24_mux2to15_and1;
  assign f_arrdiv24_fs30_and0 = f_arrdiv24_fs30_not0 & b[6];
  assign f_arrdiv24_fs30_xor1 = f_arrdiv24_fs29_or0 ^ f_arrdiv24_fs30_xor0;
  assign f_arrdiv24_fs30_not1 = ~f_arrdiv24_fs30_xor0;
  assign f_arrdiv24_fs30_and1 = f_arrdiv24_fs30_not1 & f_arrdiv24_fs29_or0;
  assign f_arrdiv24_fs30_or0 = f_arrdiv24_fs30_and1 | f_arrdiv24_fs30_and0;
  assign f_arrdiv24_fs31_xor0 = f_arrdiv24_mux2to16_and1 ^ b[7];
  assign f_arrdiv24_fs31_not0 = ~f_arrdiv24_mux2to16_and1;
  assign f_arrdiv24_fs31_and0 = f_arrdiv24_fs31_not0 & b[7];
  assign f_arrdiv24_fs31_xor1 = f_arrdiv24_fs30_or0 ^ f_arrdiv24_fs31_xor0;
  assign f_arrdiv24_fs31_not1 = ~f_arrdiv24_fs31_xor0;
  assign f_arrdiv24_fs31_and1 = f_arrdiv24_fs31_not1 & f_arrdiv24_fs30_or0;
  assign f_arrdiv24_fs31_or0 = f_arrdiv24_fs31_and1 | f_arrdiv24_fs31_and0;
  assign f_arrdiv24_fs32_xor0 = f_arrdiv24_mux2to17_and1 ^ b[8];
  assign f_arrdiv24_fs32_not0 = ~f_arrdiv24_mux2to17_and1;
  assign f_arrdiv24_fs32_and0 = f_arrdiv24_fs32_not0 & b[8];
  assign f_arrdiv24_fs32_xor1 = f_arrdiv24_fs31_or0 ^ f_arrdiv24_fs32_xor0;
  assign f_arrdiv24_fs32_not1 = ~f_arrdiv24_fs32_xor0;
  assign f_arrdiv24_fs32_and1 = f_arrdiv24_fs32_not1 & f_arrdiv24_fs31_or0;
  assign f_arrdiv24_fs32_or0 = f_arrdiv24_fs32_and1 | f_arrdiv24_fs32_and0;
  assign f_arrdiv24_fs33_xor0 = f_arrdiv24_mux2to18_and1 ^ b[9];
  assign f_arrdiv24_fs33_not0 = ~f_arrdiv24_mux2to18_and1;
  assign f_arrdiv24_fs33_and0 = f_arrdiv24_fs33_not0 & b[9];
  assign f_arrdiv24_fs33_xor1 = f_arrdiv24_fs32_or0 ^ f_arrdiv24_fs33_xor0;
  assign f_arrdiv24_fs33_not1 = ~f_arrdiv24_fs33_xor0;
  assign f_arrdiv24_fs33_and1 = f_arrdiv24_fs33_not1 & f_arrdiv24_fs32_or0;
  assign f_arrdiv24_fs33_or0 = f_arrdiv24_fs33_and1 | f_arrdiv24_fs33_and0;
  assign f_arrdiv24_fs34_xor0 = f_arrdiv24_mux2to19_and1 ^ b[10];
  assign f_arrdiv24_fs34_not0 = ~f_arrdiv24_mux2to19_and1;
  assign f_arrdiv24_fs34_and0 = f_arrdiv24_fs34_not0 & b[10];
  assign f_arrdiv24_fs34_xor1 = f_arrdiv24_fs33_or0 ^ f_arrdiv24_fs34_xor0;
  assign f_arrdiv24_fs34_not1 = ~f_arrdiv24_fs34_xor0;
  assign f_arrdiv24_fs34_and1 = f_arrdiv24_fs34_not1 & f_arrdiv24_fs33_or0;
  assign f_arrdiv24_fs34_or0 = f_arrdiv24_fs34_and1 | f_arrdiv24_fs34_and0;
  assign f_arrdiv24_fs35_xor0 = f_arrdiv24_mux2to110_and1 ^ b[11];
  assign f_arrdiv24_fs35_not0 = ~f_arrdiv24_mux2to110_and1;
  assign f_arrdiv24_fs35_and0 = f_arrdiv24_fs35_not0 & b[11];
  assign f_arrdiv24_fs35_xor1 = f_arrdiv24_fs34_or0 ^ f_arrdiv24_fs35_xor0;
  assign f_arrdiv24_fs35_not1 = ~f_arrdiv24_fs35_xor0;
  assign f_arrdiv24_fs35_and1 = f_arrdiv24_fs35_not1 & f_arrdiv24_fs34_or0;
  assign f_arrdiv24_fs35_or0 = f_arrdiv24_fs35_and1 | f_arrdiv24_fs35_and0;
  assign f_arrdiv24_fs36_xor0 = f_arrdiv24_mux2to111_and1 ^ b[12];
  assign f_arrdiv24_fs36_not0 = ~f_arrdiv24_mux2to111_and1;
  assign f_arrdiv24_fs36_and0 = f_arrdiv24_fs36_not0 & b[12];
  assign f_arrdiv24_fs36_xor1 = f_arrdiv24_fs35_or0 ^ f_arrdiv24_fs36_xor0;
  assign f_arrdiv24_fs36_not1 = ~f_arrdiv24_fs36_xor0;
  assign f_arrdiv24_fs36_and1 = f_arrdiv24_fs36_not1 & f_arrdiv24_fs35_or0;
  assign f_arrdiv24_fs36_or0 = f_arrdiv24_fs36_and1 | f_arrdiv24_fs36_and0;
  assign f_arrdiv24_fs37_xor0 = f_arrdiv24_mux2to112_and1 ^ b[13];
  assign f_arrdiv24_fs37_not0 = ~f_arrdiv24_mux2to112_and1;
  assign f_arrdiv24_fs37_and0 = f_arrdiv24_fs37_not0 & b[13];
  assign f_arrdiv24_fs37_xor1 = f_arrdiv24_fs36_or0 ^ f_arrdiv24_fs37_xor0;
  assign f_arrdiv24_fs37_not1 = ~f_arrdiv24_fs37_xor0;
  assign f_arrdiv24_fs37_and1 = f_arrdiv24_fs37_not1 & f_arrdiv24_fs36_or0;
  assign f_arrdiv24_fs37_or0 = f_arrdiv24_fs37_and1 | f_arrdiv24_fs37_and0;
  assign f_arrdiv24_fs38_xor0 = f_arrdiv24_mux2to113_and1 ^ b[14];
  assign f_arrdiv24_fs38_not0 = ~f_arrdiv24_mux2to113_and1;
  assign f_arrdiv24_fs38_and0 = f_arrdiv24_fs38_not0 & b[14];
  assign f_arrdiv24_fs38_xor1 = f_arrdiv24_fs37_or0 ^ f_arrdiv24_fs38_xor0;
  assign f_arrdiv24_fs38_not1 = ~f_arrdiv24_fs38_xor0;
  assign f_arrdiv24_fs38_and1 = f_arrdiv24_fs38_not1 & f_arrdiv24_fs37_or0;
  assign f_arrdiv24_fs38_or0 = f_arrdiv24_fs38_and1 | f_arrdiv24_fs38_and0;
  assign f_arrdiv24_fs39_xor0 = f_arrdiv24_mux2to114_and1 ^ b[15];
  assign f_arrdiv24_fs39_not0 = ~f_arrdiv24_mux2to114_and1;
  assign f_arrdiv24_fs39_and0 = f_arrdiv24_fs39_not0 & b[15];
  assign f_arrdiv24_fs39_xor1 = f_arrdiv24_fs38_or0 ^ f_arrdiv24_fs39_xor0;
  assign f_arrdiv24_fs39_not1 = ~f_arrdiv24_fs39_xor0;
  assign f_arrdiv24_fs39_and1 = f_arrdiv24_fs39_not1 & f_arrdiv24_fs38_or0;
  assign f_arrdiv24_fs39_or0 = f_arrdiv24_fs39_and1 | f_arrdiv24_fs39_and0;
  assign f_arrdiv24_fs40_xor0 = f_arrdiv24_mux2to115_and1 ^ b[16];
  assign f_arrdiv24_fs40_not0 = ~f_arrdiv24_mux2to115_and1;
  assign f_arrdiv24_fs40_and0 = f_arrdiv24_fs40_not0 & b[16];
  assign f_arrdiv24_fs40_xor1 = f_arrdiv24_fs39_or0 ^ f_arrdiv24_fs40_xor0;
  assign f_arrdiv24_fs40_not1 = ~f_arrdiv24_fs40_xor0;
  assign f_arrdiv24_fs40_and1 = f_arrdiv24_fs40_not1 & f_arrdiv24_fs39_or0;
  assign f_arrdiv24_fs40_or0 = f_arrdiv24_fs40_and1 | f_arrdiv24_fs40_and0;
  assign f_arrdiv24_fs41_xor0 = f_arrdiv24_mux2to116_and1 ^ b[17];
  assign f_arrdiv24_fs41_not0 = ~f_arrdiv24_mux2to116_and1;
  assign f_arrdiv24_fs41_and0 = f_arrdiv24_fs41_not0 & b[17];
  assign f_arrdiv24_fs41_xor1 = f_arrdiv24_fs40_or0 ^ f_arrdiv24_fs41_xor0;
  assign f_arrdiv24_fs41_not1 = ~f_arrdiv24_fs41_xor0;
  assign f_arrdiv24_fs41_and1 = f_arrdiv24_fs41_not1 & f_arrdiv24_fs40_or0;
  assign f_arrdiv24_fs41_or0 = f_arrdiv24_fs41_and1 | f_arrdiv24_fs41_and0;
  assign f_arrdiv24_fs42_xor0 = f_arrdiv24_mux2to117_and1 ^ b[18];
  assign f_arrdiv24_fs42_not0 = ~f_arrdiv24_mux2to117_and1;
  assign f_arrdiv24_fs42_and0 = f_arrdiv24_fs42_not0 & b[18];
  assign f_arrdiv24_fs42_xor1 = f_arrdiv24_fs41_or0 ^ f_arrdiv24_fs42_xor0;
  assign f_arrdiv24_fs42_not1 = ~f_arrdiv24_fs42_xor0;
  assign f_arrdiv24_fs42_and1 = f_arrdiv24_fs42_not1 & f_arrdiv24_fs41_or0;
  assign f_arrdiv24_fs42_or0 = f_arrdiv24_fs42_and1 | f_arrdiv24_fs42_and0;
  assign f_arrdiv24_fs43_xor0 = f_arrdiv24_mux2to118_and1 ^ b[19];
  assign f_arrdiv24_fs43_not0 = ~f_arrdiv24_mux2to118_and1;
  assign f_arrdiv24_fs43_and0 = f_arrdiv24_fs43_not0 & b[19];
  assign f_arrdiv24_fs43_xor1 = f_arrdiv24_fs42_or0 ^ f_arrdiv24_fs43_xor0;
  assign f_arrdiv24_fs43_not1 = ~f_arrdiv24_fs43_xor0;
  assign f_arrdiv24_fs43_and1 = f_arrdiv24_fs43_not1 & f_arrdiv24_fs42_or0;
  assign f_arrdiv24_fs43_or0 = f_arrdiv24_fs43_and1 | f_arrdiv24_fs43_and0;
  assign f_arrdiv24_fs44_xor0 = f_arrdiv24_mux2to119_and1 ^ b[20];
  assign f_arrdiv24_fs44_not0 = ~f_arrdiv24_mux2to119_and1;
  assign f_arrdiv24_fs44_and0 = f_arrdiv24_fs44_not0 & b[20];
  assign f_arrdiv24_fs44_xor1 = f_arrdiv24_fs43_or0 ^ f_arrdiv24_fs44_xor0;
  assign f_arrdiv24_fs44_not1 = ~f_arrdiv24_fs44_xor0;
  assign f_arrdiv24_fs44_and1 = f_arrdiv24_fs44_not1 & f_arrdiv24_fs43_or0;
  assign f_arrdiv24_fs44_or0 = f_arrdiv24_fs44_and1 | f_arrdiv24_fs44_and0;
  assign f_arrdiv24_fs45_xor0 = f_arrdiv24_mux2to120_and1 ^ b[21];
  assign f_arrdiv24_fs45_not0 = ~f_arrdiv24_mux2to120_and1;
  assign f_arrdiv24_fs45_and0 = f_arrdiv24_fs45_not0 & b[21];
  assign f_arrdiv24_fs45_xor1 = f_arrdiv24_fs44_or0 ^ f_arrdiv24_fs45_xor0;
  assign f_arrdiv24_fs45_not1 = ~f_arrdiv24_fs45_xor0;
  assign f_arrdiv24_fs45_and1 = f_arrdiv24_fs45_not1 & f_arrdiv24_fs44_or0;
  assign f_arrdiv24_fs45_or0 = f_arrdiv24_fs45_and1 | f_arrdiv24_fs45_and0;
  assign f_arrdiv24_fs46_xor0 = f_arrdiv24_mux2to121_and1 ^ b[22];
  assign f_arrdiv24_fs46_not0 = ~f_arrdiv24_mux2to121_and1;
  assign f_arrdiv24_fs46_and0 = f_arrdiv24_fs46_not0 & b[22];
  assign f_arrdiv24_fs46_xor1 = f_arrdiv24_fs45_or0 ^ f_arrdiv24_fs46_xor0;
  assign f_arrdiv24_fs46_not1 = ~f_arrdiv24_fs46_xor0;
  assign f_arrdiv24_fs46_and1 = f_arrdiv24_fs46_not1 & f_arrdiv24_fs45_or0;
  assign f_arrdiv24_fs46_or0 = f_arrdiv24_fs46_and1 | f_arrdiv24_fs46_and0;
  assign f_arrdiv24_fs47_xor0 = f_arrdiv24_mux2to122_and1 ^ b[23];
  assign f_arrdiv24_fs47_not0 = ~f_arrdiv24_mux2to122_and1;
  assign f_arrdiv24_fs47_and0 = f_arrdiv24_fs47_not0 & b[23];
  assign f_arrdiv24_fs47_xor1 = f_arrdiv24_fs46_or0 ^ f_arrdiv24_fs47_xor0;
  assign f_arrdiv24_fs47_not1 = ~f_arrdiv24_fs47_xor0;
  assign f_arrdiv24_fs47_and1 = f_arrdiv24_fs47_not1 & f_arrdiv24_fs46_or0;
  assign f_arrdiv24_fs47_or0 = f_arrdiv24_fs47_and1 | f_arrdiv24_fs47_and0;
  assign f_arrdiv24_mux2to123_and0 = a[22] & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to123_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to123_and1 = f_arrdiv24_fs24_xor0 & f_arrdiv24_mux2to123_not0;
  assign f_arrdiv24_mux2to123_xor0 = f_arrdiv24_mux2to123_and0 ^ f_arrdiv24_mux2to123_and1;
  assign f_arrdiv24_mux2to124_and0 = f_arrdiv24_mux2to10_xor0 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to124_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to124_and1 = f_arrdiv24_fs25_xor1 & f_arrdiv24_mux2to124_not0;
  assign f_arrdiv24_mux2to124_xor0 = f_arrdiv24_mux2to124_and0 ^ f_arrdiv24_mux2to124_and1;
  assign f_arrdiv24_mux2to125_and0 = f_arrdiv24_mux2to11_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to125_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to125_and1 = f_arrdiv24_fs26_xor1 & f_arrdiv24_mux2to125_not0;
  assign f_arrdiv24_mux2to125_xor0 = f_arrdiv24_mux2to125_and0 ^ f_arrdiv24_mux2to125_and1;
  assign f_arrdiv24_mux2to126_and0 = f_arrdiv24_mux2to12_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to126_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to126_and1 = f_arrdiv24_fs27_xor1 & f_arrdiv24_mux2to126_not0;
  assign f_arrdiv24_mux2to126_xor0 = f_arrdiv24_mux2to126_and0 ^ f_arrdiv24_mux2to126_and1;
  assign f_arrdiv24_mux2to127_and0 = f_arrdiv24_mux2to13_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to127_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to127_and1 = f_arrdiv24_fs28_xor1 & f_arrdiv24_mux2to127_not0;
  assign f_arrdiv24_mux2to127_xor0 = f_arrdiv24_mux2to127_and0 ^ f_arrdiv24_mux2to127_and1;
  assign f_arrdiv24_mux2to128_and0 = f_arrdiv24_mux2to14_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to128_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to128_and1 = f_arrdiv24_fs29_xor1 & f_arrdiv24_mux2to128_not0;
  assign f_arrdiv24_mux2to128_xor0 = f_arrdiv24_mux2to128_and0 ^ f_arrdiv24_mux2to128_and1;
  assign f_arrdiv24_mux2to129_and0 = f_arrdiv24_mux2to15_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to129_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to129_and1 = f_arrdiv24_fs30_xor1 & f_arrdiv24_mux2to129_not0;
  assign f_arrdiv24_mux2to129_xor0 = f_arrdiv24_mux2to129_and0 ^ f_arrdiv24_mux2to129_and1;
  assign f_arrdiv24_mux2to130_and0 = f_arrdiv24_mux2to16_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to130_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to130_and1 = f_arrdiv24_fs31_xor1 & f_arrdiv24_mux2to130_not0;
  assign f_arrdiv24_mux2to130_xor0 = f_arrdiv24_mux2to130_and0 ^ f_arrdiv24_mux2to130_and1;
  assign f_arrdiv24_mux2to131_and0 = f_arrdiv24_mux2to17_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to131_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to131_and1 = f_arrdiv24_fs32_xor1 & f_arrdiv24_mux2to131_not0;
  assign f_arrdiv24_mux2to131_xor0 = f_arrdiv24_mux2to131_and0 ^ f_arrdiv24_mux2to131_and1;
  assign f_arrdiv24_mux2to132_and0 = f_arrdiv24_mux2to18_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to132_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to132_and1 = f_arrdiv24_fs33_xor1 & f_arrdiv24_mux2to132_not0;
  assign f_arrdiv24_mux2to132_xor0 = f_arrdiv24_mux2to132_and0 ^ f_arrdiv24_mux2to132_and1;
  assign f_arrdiv24_mux2to133_and0 = f_arrdiv24_mux2to19_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to133_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to133_and1 = f_arrdiv24_fs34_xor1 & f_arrdiv24_mux2to133_not0;
  assign f_arrdiv24_mux2to133_xor0 = f_arrdiv24_mux2to133_and0 ^ f_arrdiv24_mux2to133_and1;
  assign f_arrdiv24_mux2to134_and0 = f_arrdiv24_mux2to110_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to134_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to134_and1 = f_arrdiv24_fs35_xor1 & f_arrdiv24_mux2to134_not0;
  assign f_arrdiv24_mux2to134_xor0 = f_arrdiv24_mux2to134_and0 ^ f_arrdiv24_mux2to134_and1;
  assign f_arrdiv24_mux2to135_and0 = f_arrdiv24_mux2to111_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to135_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to135_and1 = f_arrdiv24_fs36_xor1 & f_arrdiv24_mux2to135_not0;
  assign f_arrdiv24_mux2to135_xor0 = f_arrdiv24_mux2to135_and0 ^ f_arrdiv24_mux2to135_and1;
  assign f_arrdiv24_mux2to136_and0 = f_arrdiv24_mux2to112_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to136_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to136_and1 = f_arrdiv24_fs37_xor1 & f_arrdiv24_mux2to136_not0;
  assign f_arrdiv24_mux2to136_xor0 = f_arrdiv24_mux2to136_and0 ^ f_arrdiv24_mux2to136_and1;
  assign f_arrdiv24_mux2to137_and0 = f_arrdiv24_mux2to113_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to137_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to137_and1 = f_arrdiv24_fs38_xor1 & f_arrdiv24_mux2to137_not0;
  assign f_arrdiv24_mux2to137_xor0 = f_arrdiv24_mux2to137_and0 ^ f_arrdiv24_mux2to137_and1;
  assign f_arrdiv24_mux2to138_and0 = f_arrdiv24_mux2to114_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to138_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to138_and1 = f_arrdiv24_fs39_xor1 & f_arrdiv24_mux2to138_not0;
  assign f_arrdiv24_mux2to138_xor0 = f_arrdiv24_mux2to138_and0 ^ f_arrdiv24_mux2to138_and1;
  assign f_arrdiv24_mux2to139_and0 = f_arrdiv24_mux2to115_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to139_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to139_and1 = f_arrdiv24_fs40_xor1 & f_arrdiv24_mux2to139_not0;
  assign f_arrdiv24_mux2to139_xor0 = f_arrdiv24_mux2to139_and0 ^ f_arrdiv24_mux2to139_and1;
  assign f_arrdiv24_mux2to140_and0 = f_arrdiv24_mux2to116_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to140_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to140_and1 = f_arrdiv24_fs41_xor1 & f_arrdiv24_mux2to140_not0;
  assign f_arrdiv24_mux2to140_xor0 = f_arrdiv24_mux2to140_and0 ^ f_arrdiv24_mux2to140_and1;
  assign f_arrdiv24_mux2to141_and0 = f_arrdiv24_mux2to117_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to141_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to141_and1 = f_arrdiv24_fs42_xor1 & f_arrdiv24_mux2to141_not0;
  assign f_arrdiv24_mux2to141_xor0 = f_arrdiv24_mux2to141_and0 ^ f_arrdiv24_mux2to141_and1;
  assign f_arrdiv24_mux2to142_and0 = f_arrdiv24_mux2to118_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to142_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to142_and1 = f_arrdiv24_fs43_xor1 & f_arrdiv24_mux2to142_not0;
  assign f_arrdiv24_mux2to142_xor0 = f_arrdiv24_mux2to142_and0 ^ f_arrdiv24_mux2to142_and1;
  assign f_arrdiv24_mux2to143_and0 = f_arrdiv24_mux2to119_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to143_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to143_and1 = f_arrdiv24_fs44_xor1 & f_arrdiv24_mux2to143_not0;
  assign f_arrdiv24_mux2to143_xor0 = f_arrdiv24_mux2to143_and0 ^ f_arrdiv24_mux2to143_and1;
  assign f_arrdiv24_mux2to144_and0 = f_arrdiv24_mux2to120_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to144_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to144_and1 = f_arrdiv24_fs45_xor1 & f_arrdiv24_mux2to144_not0;
  assign f_arrdiv24_mux2to144_xor0 = f_arrdiv24_mux2to144_and0 ^ f_arrdiv24_mux2to144_and1;
  assign f_arrdiv24_mux2to145_and0 = f_arrdiv24_mux2to121_and1 & f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to145_not0 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_mux2to145_and1 = f_arrdiv24_fs46_xor1 & f_arrdiv24_mux2to145_not0;
  assign f_arrdiv24_mux2to145_xor0 = f_arrdiv24_mux2to145_and0 ^ f_arrdiv24_mux2to145_and1;
  assign f_arrdiv24_not1 = ~f_arrdiv24_fs47_or0;
  assign f_arrdiv24_fs48_xor0 = a[21] ^ b[0];
  assign f_arrdiv24_fs48_not0 = ~a[21];
  assign f_arrdiv24_fs48_and0 = f_arrdiv24_fs48_not0 & b[0];
  assign f_arrdiv24_fs48_not1 = ~f_arrdiv24_fs48_xor0;
  assign f_arrdiv24_fs49_xor0 = f_arrdiv24_mux2to123_xor0 ^ b[1];
  assign f_arrdiv24_fs49_not0 = ~f_arrdiv24_mux2to123_xor0;
  assign f_arrdiv24_fs49_and0 = f_arrdiv24_fs49_not0 & b[1];
  assign f_arrdiv24_fs49_xor1 = f_arrdiv24_fs48_and0 ^ f_arrdiv24_fs49_xor0;
  assign f_arrdiv24_fs49_not1 = ~f_arrdiv24_fs49_xor0;
  assign f_arrdiv24_fs49_and1 = f_arrdiv24_fs49_not1 & f_arrdiv24_fs48_and0;
  assign f_arrdiv24_fs49_or0 = f_arrdiv24_fs49_and1 | f_arrdiv24_fs49_and0;
  assign f_arrdiv24_fs50_xor0 = f_arrdiv24_mux2to124_xor0 ^ b[2];
  assign f_arrdiv24_fs50_not0 = ~f_arrdiv24_mux2to124_xor0;
  assign f_arrdiv24_fs50_and0 = f_arrdiv24_fs50_not0 & b[2];
  assign f_arrdiv24_fs50_xor1 = f_arrdiv24_fs49_or0 ^ f_arrdiv24_fs50_xor0;
  assign f_arrdiv24_fs50_not1 = ~f_arrdiv24_fs50_xor0;
  assign f_arrdiv24_fs50_and1 = f_arrdiv24_fs50_not1 & f_arrdiv24_fs49_or0;
  assign f_arrdiv24_fs50_or0 = f_arrdiv24_fs50_and1 | f_arrdiv24_fs50_and0;
  assign f_arrdiv24_fs51_xor0 = f_arrdiv24_mux2to125_xor0 ^ b[3];
  assign f_arrdiv24_fs51_not0 = ~f_arrdiv24_mux2to125_xor0;
  assign f_arrdiv24_fs51_and0 = f_arrdiv24_fs51_not0 & b[3];
  assign f_arrdiv24_fs51_xor1 = f_arrdiv24_fs50_or0 ^ f_arrdiv24_fs51_xor0;
  assign f_arrdiv24_fs51_not1 = ~f_arrdiv24_fs51_xor0;
  assign f_arrdiv24_fs51_and1 = f_arrdiv24_fs51_not1 & f_arrdiv24_fs50_or0;
  assign f_arrdiv24_fs51_or0 = f_arrdiv24_fs51_and1 | f_arrdiv24_fs51_and0;
  assign f_arrdiv24_fs52_xor0 = f_arrdiv24_mux2to126_xor0 ^ b[4];
  assign f_arrdiv24_fs52_not0 = ~f_arrdiv24_mux2to126_xor0;
  assign f_arrdiv24_fs52_and0 = f_arrdiv24_fs52_not0 & b[4];
  assign f_arrdiv24_fs52_xor1 = f_arrdiv24_fs51_or0 ^ f_arrdiv24_fs52_xor0;
  assign f_arrdiv24_fs52_not1 = ~f_arrdiv24_fs52_xor0;
  assign f_arrdiv24_fs52_and1 = f_arrdiv24_fs52_not1 & f_arrdiv24_fs51_or0;
  assign f_arrdiv24_fs52_or0 = f_arrdiv24_fs52_and1 | f_arrdiv24_fs52_and0;
  assign f_arrdiv24_fs53_xor0 = f_arrdiv24_mux2to127_xor0 ^ b[5];
  assign f_arrdiv24_fs53_not0 = ~f_arrdiv24_mux2to127_xor0;
  assign f_arrdiv24_fs53_and0 = f_arrdiv24_fs53_not0 & b[5];
  assign f_arrdiv24_fs53_xor1 = f_arrdiv24_fs52_or0 ^ f_arrdiv24_fs53_xor0;
  assign f_arrdiv24_fs53_not1 = ~f_arrdiv24_fs53_xor0;
  assign f_arrdiv24_fs53_and1 = f_arrdiv24_fs53_not1 & f_arrdiv24_fs52_or0;
  assign f_arrdiv24_fs53_or0 = f_arrdiv24_fs53_and1 | f_arrdiv24_fs53_and0;
  assign f_arrdiv24_fs54_xor0 = f_arrdiv24_mux2to128_xor0 ^ b[6];
  assign f_arrdiv24_fs54_not0 = ~f_arrdiv24_mux2to128_xor0;
  assign f_arrdiv24_fs54_and0 = f_arrdiv24_fs54_not0 & b[6];
  assign f_arrdiv24_fs54_xor1 = f_arrdiv24_fs53_or0 ^ f_arrdiv24_fs54_xor0;
  assign f_arrdiv24_fs54_not1 = ~f_arrdiv24_fs54_xor0;
  assign f_arrdiv24_fs54_and1 = f_arrdiv24_fs54_not1 & f_arrdiv24_fs53_or0;
  assign f_arrdiv24_fs54_or0 = f_arrdiv24_fs54_and1 | f_arrdiv24_fs54_and0;
  assign f_arrdiv24_fs55_xor0 = f_arrdiv24_mux2to129_xor0 ^ b[7];
  assign f_arrdiv24_fs55_not0 = ~f_arrdiv24_mux2to129_xor0;
  assign f_arrdiv24_fs55_and0 = f_arrdiv24_fs55_not0 & b[7];
  assign f_arrdiv24_fs55_xor1 = f_arrdiv24_fs54_or0 ^ f_arrdiv24_fs55_xor0;
  assign f_arrdiv24_fs55_not1 = ~f_arrdiv24_fs55_xor0;
  assign f_arrdiv24_fs55_and1 = f_arrdiv24_fs55_not1 & f_arrdiv24_fs54_or0;
  assign f_arrdiv24_fs55_or0 = f_arrdiv24_fs55_and1 | f_arrdiv24_fs55_and0;
  assign f_arrdiv24_fs56_xor0 = f_arrdiv24_mux2to130_xor0 ^ b[8];
  assign f_arrdiv24_fs56_not0 = ~f_arrdiv24_mux2to130_xor0;
  assign f_arrdiv24_fs56_and0 = f_arrdiv24_fs56_not0 & b[8];
  assign f_arrdiv24_fs56_xor1 = f_arrdiv24_fs55_or0 ^ f_arrdiv24_fs56_xor0;
  assign f_arrdiv24_fs56_not1 = ~f_arrdiv24_fs56_xor0;
  assign f_arrdiv24_fs56_and1 = f_arrdiv24_fs56_not1 & f_arrdiv24_fs55_or0;
  assign f_arrdiv24_fs56_or0 = f_arrdiv24_fs56_and1 | f_arrdiv24_fs56_and0;
  assign f_arrdiv24_fs57_xor0 = f_arrdiv24_mux2to131_xor0 ^ b[9];
  assign f_arrdiv24_fs57_not0 = ~f_arrdiv24_mux2to131_xor0;
  assign f_arrdiv24_fs57_and0 = f_arrdiv24_fs57_not0 & b[9];
  assign f_arrdiv24_fs57_xor1 = f_arrdiv24_fs56_or0 ^ f_arrdiv24_fs57_xor0;
  assign f_arrdiv24_fs57_not1 = ~f_arrdiv24_fs57_xor0;
  assign f_arrdiv24_fs57_and1 = f_arrdiv24_fs57_not1 & f_arrdiv24_fs56_or0;
  assign f_arrdiv24_fs57_or0 = f_arrdiv24_fs57_and1 | f_arrdiv24_fs57_and0;
  assign f_arrdiv24_fs58_xor0 = f_arrdiv24_mux2to132_xor0 ^ b[10];
  assign f_arrdiv24_fs58_not0 = ~f_arrdiv24_mux2to132_xor0;
  assign f_arrdiv24_fs58_and0 = f_arrdiv24_fs58_not0 & b[10];
  assign f_arrdiv24_fs58_xor1 = f_arrdiv24_fs57_or0 ^ f_arrdiv24_fs58_xor0;
  assign f_arrdiv24_fs58_not1 = ~f_arrdiv24_fs58_xor0;
  assign f_arrdiv24_fs58_and1 = f_arrdiv24_fs58_not1 & f_arrdiv24_fs57_or0;
  assign f_arrdiv24_fs58_or0 = f_arrdiv24_fs58_and1 | f_arrdiv24_fs58_and0;
  assign f_arrdiv24_fs59_xor0 = f_arrdiv24_mux2to133_xor0 ^ b[11];
  assign f_arrdiv24_fs59_not0 = ~f_arrdiv24_mux2to133_xor0;
  assign f_arrdiv24_fs59_and0 = f_arrdiv24_fs59_not0 & b[11];
  assign f_arrdiv24_fs59_xor1 = f_arrdiv24_fs58_or0 ^ f_arrdiv24_fs59_xor0;
  assign f_arrdiv24_fs59_not1 = ~f_arrdiv24_fs59_xor0;
  assign f_arrdiv24_fs59_and1 = f_arrdiv24_fs59_not1 & f_arrdiv24_fs58_or0;
  assign f_arrdiv24_fs59_or0 = f_arrdiv24_fs59_and1 | f_arrdiv24_fs59_and0;
  assign f_arrdiv24_fs60_xor0 = f_arrdiv24_mux2to134_xor0 ^ b[12];
  assign f_arrdiv24_fs60_not0 = ~f_arrdiv24_mux2to134_xor0;
  assign f_arrdiv24_fs60_and0 = f_arrdiv24_fs60_not0 & b[12];
  assign f_arrdiv24_fs60_xor1 = f_arrdiv24_fs59_or0 ^ f_arrdiv24_fs60_xor0;
  assign f_arrdiv24_fs60_not1 = ~f_arrdiv24_fs60_xor0;
  assign f_arrdiv24_fs60_and1 = f_arrdiv24_fs60_not1 & f_arrdiv24_fs59_or0;
  assign f_arrdiv24_fs60_or0 = f_arrdiv24_fs60_and1 | f_arrdiv24_fs60_and0;
  assign f_arrdiv24_fs61_xor0 = f_arrdiv24_mux2to135_xor0 ^ b[13];
  assign f_arrdiv24_fs61_not0 = ~f_arrdiv24_mux2to135_xor0;
  assign f_arrdiv24_fs61_and0 = f_arrdiv24_fs61_not0 & b[13];
  assign f_arrdiv24_fs61_xor1 = f_arrdiv24_fs60_or0 ^ f_arrdiv24_fs61_xor0;
  assign f_arrdiv24_fs61_not1 = ~f_arrdiv24_fs61_xor0;
  assign f_arrdiv24_fs61_and1 = f_arrdiv24_fs61_not1 & f_arrdiv24_fs60_or0;
  assign f_arrdiv24_fs61_or0 = f_arrdiv24_fs61_and1 | f_arrdiv24_fs61_and0;
  assign f_arrdiv24_fs62_xor0 = f_arrdiv24_mux2to136_xor0 ^ b[14];
  assign f_arrdiv24_fs62_not0 = ~f_arrdiv24_mux2to136_xor0;
  assign f_arrdiv24_fs62_and0 = f_arrdiv24_fs62_not0 & b[14];
  assign f_arrdiv24_fs62_xor1 = f_arrdiv24_fs61_or0 ^ f_arrdiv24_fs62_xor0;
  assign f_arrdiv24_fs62_not1 = ~f_arrdiv24_fs62_xor0;
  assign f_arrdiv24_fs62_and1 = f_arrdiv24_fs62_not1 & f_arrdiv24_fs61_or0;
  assign f_arrdiv24_fs62_or0 = f_arrdiv24_fs62_and1 | f_arrdiv24_fs62_and0;
  assign f_arrdiv24_fs63_xor0 = f_arrdiv24_mux2to137_xor0 ^ b[15];
  assign f_arrdiv24_fs63_not0 = ~f_arrdiv24_mux2to137_xor0;
  assign f_arrdiv24_fs63_and0 = f_arrdiv24_fs63_not0 & b[15];
  assign f_arrdiv24_fs63_xor1 = f_arrdiv24_fs62_or0 ^ f_arrdiv24_fs63_xor0;
  assign f_arrdiv24_fs63_not1 = ~f_arrdiv24_fs63_xor0;
  assign f_arrdiv24_fs63_and1 = f_arrdiv24_fs63_not1 & f_arrdiv24_fs62_or0;
  assign f_arrdiv24_fs63_or0 = f_arrdiv24_fs63_and1 | f_arrdiv24_fs63_and0;
  assign f_arrdiv24_fs64_xor0 = f_arrdiv24_mux2to138_xor0 ^ b[16];
  assign f_arrdiv24_fs64_not0 = ~f_arrdiv24_mux2to138_xor0;
  assign f_arrdiv24_fs64_and0 = f_arrdiv24_fs64_not0 & b[16];
  assign f_arrdiv24_fs64_xor1 = f_arrdiv24_fs63_or0 ^ f_arrdiv24_fs64_xor0;
  assign f_arrdiv24_fs64_not1 = ~f_arrdiv24_fs64_xor0;
  assign f_arrdiv24_fs64_and1 = f_arrdiv24_fs64_not1 & f_arrdiv24_fs63_or0;
  assign f_arrdiv24_fs64_or0 = f_arrdiv24_fs64_and1 | f_arrdiv24_fs64_and0;
  assign f_arrdiv24_fs65_xor0 = f_arrdiv24_mux2to139_xor0 ^ b[17];
  assign f_arrdiv24_fs65_not0 = ~f_arrdiv24_mux2to139_xor0;
  assign f_arrdiv24_fs65_and0 = f_arrdiv24_fs65_not0 & b[17];
  assign f_arrdiv24_fs65_xor1 = f_arrdiv24_fs64_or0 ^ f_arrdiv24_fs65_xor0;
  assign f_arrdiv24_fs65_not1 = ~f_arrdiv24_fs65_xor0;
  assign f_arrdiv24_fs65_and1 = f_arrdiv24_fs65_not1 & f_arrdiv24_fs64_or0;
  assign f_arrdiv24_fs65_or0 = f_arrdiv24_fs65_and1 | f_arrdiv24_fs65_and0;
  assign f_arrdiv24_fs66_xor0 = f_arrdiv24_mux2to140_xor0 ^ b[18];
  assign f_arrdiv24_fs66_not0 = ~f_arrdiv24_mux2to140_xor0;
  assign f_arrdiv24_fs66_and0 = f_arrdiv24_fs66_not0 & b[18];
  assign f_arrdiv24_fs66_xor1 = f_arrdiv24_fs65_or0 ^ f_arrdiv24_fs66_xor0;
  assign f_arrdiv24_fs66_not1 = ~f_arrdiv24_fs66_xor0;
  assign f_arrdiv24_fs66_and1 = f_arrdiv24_fs66_not1 & f_arrdiv24_fs65_or0;
  assign f_arrdiv24_fs66_or0 = f_arrdiv24_fs66_and1 | f_arrdiv24_fs66_and0;
  assign f_arrdiv24_fs67_xor0 = f_arrdiv24_mux2to141_xor0 ^ b[19];
  assign f_arrdiv24_fs67_not0 = ~f_arrdiv24_mux2to141_xor0;
  assign f_arrdiv24_fs67_and0 = f_arrdiv24_fs67_not0 & b[19];
  assign f_arrdiv24_fs67_xor1 = f_arrdiv24_fs66_or0 ^ f_arrdiv24_fs67_xor0;
  assign f_arrdiv24_fs67_not1 = ~f_arrdiv24_fs67_xor0;
  assign f_arrdiv24_fs67_and1 = f_arrdiv24_fs67_not1 & f_arrdiv24_fs66_or0;
  assign f_arrdiv24_fs67_or0 = f_arrdiv24_fs67_and1 | f_arrdiv24_fs67_and0;
  assign f_arrdiv24_fs68_xor0 = f_arrdiv24_mux2to142_xor0 ^ b[20];
  assign f_arrdiv24_fs68_not0 = ~f_arrdiv24_mux2to142_xor0;
  assign f_arrdiv24_fs68_and0 = f_arrdiv24_fs68_not0 & b[20];
  assign f_arrdiv24_fs68_xor1 = f_arrdiv24_fs67_or0 ^ f_arrdiv24_fs68_xor0;
  assign f_arrdiv24_fs68_not1 = ~f_arrdiv24_fs68_xor0;
  assign f_arrdiv24_fs68_and1 = f_arrdiv24_fs68_not1 & f_arrdiv24_fs67_or0;
  assign f_arrdiv24_fs68_or0 = f_arrdiv24_fs68_and1 | f_arrdiv24_fs68_and0;
  assign f_arrdiv24_fs69_xor0 = f_arrdiv24_mux2to143_xor0 ^ b[21];
  assign f_arrdiv24_fs69_not0 = ~f_arrdiv24_mux2to143_xor0;
  assign f_arrdiv24_fs69_and0 = f_arrdiv24_fs69_not0 & b[21];
  assign f_arrdiv24_fs69_xor1 = f_arrdiv24_fs68_or0 ^ f_arrdiv24_fs69_xor0;
  assign f_arrdiv24_fs69_not1 = ~f_arrdiv24_fs69_xor0;
  assign f_arrdiv24_fs69_and1 = f_arrdiv24_fs69_not1 & f_arrdiv24_fs68_or0;
  assign f_arrdiv24_fs69_or0 = f_arrdiv24_fs69_and1 | f_arrdiv24_fs69_and0;
  assign f_arrdiv24_fs70_xor0 = f_arrdiv24_mux2to144_xor0 ^ b[22];
  assign f_arrdiv24_fs70_not0 = ~f_arrdiv24_mux2to144_xor0;
  assign f_arrdiv24_fs70_and0 = f_arrdiv24_fs70_not0 & b[22];
  assign f_arrdiv24_fs70_xor1 = f_arrdiv24_fs69_or0 ^ f_arrdiv24_fs70_xor0;
  assign f_arrdiv24_fs70_not1 = ~f_arrdiv24_fs70_xor0;
  assign f_arrdiv24_fs70_and1 = f_arrdiv24_fs70_not1 & f_arrdiv24_fs69_or0;
  assign f_arrdiv24_fs70_or0 = f_arrdiv24_fs70_and1 | f_arrdiv24_fs70_and0;
  assign f_arrdiv24_fs71_xor0 = f_arrdiv24_mux2to145_xor0 ^ b[23];
  assign f_arrdiv24_fs71_not0 = ~f_arrdiv24_mux2to145_xor0;
  assign f_arrdiv24_fs71_and0 = f_arrdiv24_fs71_not0 & b[23];
  assign f_arrdiv24_fs71_xor1 = f_arrdiv24_fs70_or0 ^ f_arrdiv24_fs71_xor0;
  assign f_arrdiv24_fs71_not1 = ~f_arrdiv24_fs71_xor0;
  assign f_arrdiv24_fs71_and1 = f_arrdiv24_fs71_not1 & f_arrdiv24_fs70_or0;
  assign f_arrdiv24_fs71_or0 = f_arrdiv24_fs71_and1 | f_arrdiv24_fs71_and0;
  assign f_arrdiv24_mux2to146_and0 = a[21] & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to146_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to146_and1 = f_arrdiv24_fs48_xor0 & f_arrdiv24_mux2to146_not0;
  assign f_arrdiv24_mux2to146_xor0 = f_arrdiv24_mux2to146_and0 ^ f_arrdiv24_mux2to146_and1;
  assign f_arrdiv24_mux2to147_and0 = f_arrdiv24_mux2to123_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to147_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to147_and1 = f_arrdiv24_fs49_xor1 & f_arrdiv24_mux2to147_not0;
  assign f_arrdiv24_mux2to147_xor0 = f_arrdiv24_mux2to147_and0 ^ f_arrdiv24_mux2to147_and1;
  assign f_arrdiv24_mux2to148_and0 = f_arrdiv24_mux2to124_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to148_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to148_and1 = f_arrdiv24_fs50_xor1 & f_arrdiv24_mux2to148_not0;
  assign f_arrdiv24_mux2to148_xor0 = f_arrdiv24_mux2to148_and0 ^ f_arrdiv24_mux2to148_and1;
  assign f_arrdiv24_mux2to149_and0 = f_arrdiv24_mux2to125_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to149_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to149_and1 = f_arrdiv24_fs51_xor1 & f_arrdiv24_mux2to149_not0;
  assign f_arrdiv24_mux2to149_xor0 = f_arrdiv24_mux2to149_and0 ^ f_arrdiv24_mux2to149_and1;
  assign f_arrdiv24_mux2to150_and0 = f_arrdiv24_mux2to126_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to150_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to150_and1 = f_arrdiv24_fs52_xor1 & f_arrdiv24_mux2to150_not0;
  assign f_arrdiv24_mux2to150_xor0 = f_arrdiv24_mux2to150_and0 ^ f_arrdiv24_mux2to150_and1;
  assign f_arrdiv24_mux2to151_and0 = f_arrdiv24_mux2to127_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to151_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to151_and1 = f_arrdiv24_fs53_xor1 & f_arrdiv24_mux2to151_not0;
  assign f_arrdiv24_mux2to151_xor0 = f_arrdiv24_mux2to151_and0 ^ f_arrdiv24_mux2to151_and1;
  assign f_arrdiv24_mux2to152_and0 = f_arrdiv24_mux2to128_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to152_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to152_and1 = f_arrdiv24_fs54_xor1 & f_arrdiv24_mux2to152_not0;
  assign f_arrdiv24_mux2to152_xor0 = f_arrdiv24_mux2to152_and0 ^ f_arrdiv24_mux2to152_and1;
  assign f_arrdiv24_mux2to153_and0 = f_arrdiv24_mux2to129_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to153_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to153_and1 = f_arrdiv24_fs55_xor1 & f_arrdiv24_mux2to153_not0;
  assign f_arrdiv24_mux2to153_xor0 = f_arrdiv24_mux2to153_and0 ^ f_arrdiv24_mux2to153_and1;
  assign f_arrdiv24_mux2to154_and0 = f_arrdiv24_mux2to130_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to154_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to154_and1 = f_arrdiv24_fs56_xor1 & f_arrdiv24_mux2to154_not0;
  assign f_arrdiv24_mux2to154_xor0 = f_arrdiv24_mux2to154_and0 ^ f_arrdiv24_mux2to154_and1;
  assign f_arrdiv24_mux2to155_and0 = f_arrdiv24_mux2to131_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to155_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to155_and1 = f_arrdiv24_fs57_xor1 & f_arrdiv24_mux2to155_not0;
  assign f_arrdiv24_mux2to155_xor0 = f_arrdiv24_mux2to155_and0 ^ f_arrdiv24_mux2to155_and1;
  assign f_arrdiv24_mux2to156_and0 = f_arrdiv24_mux2to132_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to156_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to156_and1 = f_arrdiv24_fs58_xor1 & f_arrdiv24_mux2to156_not0;
  assign f_arrdiv24_mux2to156_xor0 = f_arrdiv24_mux2to156_and0 ^ f_arrdiv24_mux2to156_and1;
  assign f_arrdiv24_mux2to157_and0 = f_arrdiv24_mux2to133_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to157_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to157_and1 = f_arrdiv24_fs59_xor1 & f_arrdiv24_mux2to157_not0;
  assign f_arrdiv24_mux2to157_xor0 = f_arrdiv24_mux2to157_and0 ^ f_arrdiv24_mux2to157_and1;
  assign f_arrdiv24_mux2to158_and0 = f_arrdiv24_mux2to134_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to158_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to158_and1 = f_arrdiv24_fs60_xor1 & f_arrdiv24_mux2to158_not0;
  assign f_arrdiv24_mux2to158_xor0 = f_arrdiv24_mux2to158_and0 ^ f_arrdiv24_mux2to158_and1;
  assign f_arrdiv24_mux2to159_and0 = f_arrdiv24_mux2to135_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to159_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to159_and1 = f_arrdiv24_fs61_xor1 & f_arrdiv24_mux2to159_not0;
  assign f_arrdiv24_mux2to159_xor0 = f_arrdiv24_mux2to159_and0 ^ f_arrdiv24_mux2to159_and1;
  assign f_arrdiv24_mux2to160_and0 = f_arrdiv24_mux2to136_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to160_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to160_and1 = f_arrdiv24_fs62_xor1 & f_arrdiv24_mux2to160_not0;
  assign f_arrdiv24_mux2to160_xor0 = f_arrdiv24_mux2to160_and0 ^ f_arrdiv24_mux2to160_and1;
  assign f_arrdiv24_mux2to161_and0 = f_arrdiv24_mux2to137_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to161_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to161_and1 = f_arrdiv24_fs63_xor1 & f_arrdiv24_mux2to161_not0;
  assign f_arrdiv24_mux2to161_xor0 = f_arrdiv24_mux2to161_and0 ^ f_arrdiv24_mux2to161_and1;
  assign f_arrdiv24_mux2to162_and0 = f_arrdiv24_mux2to138_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to162_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to162_and1 = f_arrdiv24_fs64_xor1 & f_arrdiv24_mux2to162_not0;
  assign f_arrdiv24_mux2to162_xor0 = f_arrdiv24_mux2to162_and0 ^ f_arrdiv24_mux2to162_and1;
  assign f_arrdiv24_mux2to163_and0 = f_arrdiv24_mux2to139_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to163_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to163_and1 = f_arrdiv24_fs65_xor1 & f_arrdiv24_mux2to163_not0;
  assign f_arrdiv24_mux2to163_xor0 = f_arrdiv24_mux2to163_and0 ^ f_arrdiv24_mux2to163_and1;
  assign f_arrdiv24_mux2to164_and0 = f_arrdiv24_mux2to140_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to164_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to164_and1 = f_arrdiv24_fs66_xor1 & f_arrdiv24_mux2to164_not0;
  assign f_arrdiv24_mux2to164_xor0 = f_arrdiv24_mux2to164_and0 ^ f_arrdiv24_mux2to164_and1;
  assign f_arrdiv24_mux2to165_and0 = f_arrdiv24_mux2to141_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to165_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to165_and1 = f_arrdiv24_fs67_xor1 & f_arrdiv24_mux2to165_not0;
  assign f_arrdiv24_mux2to165_xor0 = f_arrdiv24_mux2to165_and0 ^ f_arrdiv24_mux2to165_and1;
  assign f_arrdiv24_mux2to166_and0 = f_arrdiv24_mux2to142_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to166_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to166_and1 = f_arrdiv24_fs68_xor1 & f_arrdiv24_mux2to166_not0;
  assign f_arrdiv24_mux2to166_xor0 = f_arrdiv24_mux2to166_and0 ^ f_arrdiv24_mux2to166_and1;
  assign f_arrdiv24_mux2to167_and0 = f_arrdiv24_mux2to143_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to167_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to167_and1 = f_arrdiv24_fs69_xor1 & f_arrdiv24_mux2to167_not0;
  assign f_arrdiv24_mux2to167_xor0 = f_arrdiv24_mux2to167_and0 ^ f_arrdiv24_mux2to167_and1;
  assign f_arrdiv24_mux2to168_and0 = f_arrdiv24_mux2to144_xor0 & f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to168_not0 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_mux2to168_and1 = f_arrdiv24_fs70_xor1 & f_arrdiv24_mux2to168_not0;
  assign f_arrdiv24_mux2to168_xor0 = f_arrdiv24_mux2to168_and0 ^ f_arrdiv24_mux2to168_and1;
  assign f_arrdiv24_not2 = ~f_arrdiv24_fs71_or0;
  assign f_arrdiv24_fs72_xor0 = a[20] ^ b[0];
  assign f_arrdiv24_fs72_not0 = ~a[20];
  assign f_arrdiv24_fs72_and0 = f_arrdiv24_fs72_not0 & b[0];
  assign f_arrdiv24_fs72_not1 = ~f_arrdiv24_fs72_xor0;
  assign f_arrdiv24_fs73_xor0 = f_arrdiv24_mux2to146_xor0 ^ b[1];
  assign f_arrdiv24_fs73_not0 = ~f_arrdiv24_mux2to146_xor0;
  assign f_arrdiv24_fs73_and0 = f_arrdiv24_fs73_not0 & b[1];
  assign f_arrdiv24_fs73_xor1 = f_arrdiv24_fs72_and0 ^ f_arrdiv24_fs73_xor0;
  assign f_arrdiv24_fs73_not1 = ~f_arrdiv24_fs73_xor0;
  assign f_arrdiv24_fs73_and1 = f_arrdiv24_fs73_not1 & f_arrdiv24_fs72_and0;
  assign f_arrdiv24_fs73_or0 = f_arrdiv24_fs73_and1 | f_arrdiv24_fs73_and0;
  assign f_arrdiv24_fs74_xor0 = f_arrdiv24_mux2to147_xor0 ^ b[2];
  assign f_arrdiv24_fs74_not0 = ~f_arrdiv24_mux2to147_xor0;
  assign f_arrdiv24_fs74_and0 = f_arrdiv24_fs74_not0 & b[2];
  assign f_arrdiv24_fs74_xor1 = f_arrdiv24_fs73_or0 ^ f_arrdiv24_fs74_xor0;
  assign f_arrdiv24_fs74_not1 = ~f_arrdiv24_fs74_xor0;
  assign f_arrdiv24_fs74_and1 = f_arrdiv24_fs74_not1 & f_arrdiv24_fs73_or0;
  assign f_arrdiv24_fs74_or0 = f_arrdiv24_fs74_and1 | f_arrdiv24_fs74_and0;
  assign f_arrdiv24_fs75_xor0 = f_arrdiv24_mux2to148_xor0 ^ b[3];
  assign f_arrdiv24_fs75_not0 = ~f_arrdiv24_mux2to148_xor0;
  assign f_arrdiv24_fs75_and0 = f_arrdiv24_fs75_not0 & b[3];
  assign f_arrdiv24_fs75_xor1 = f_arrdiv24_fs74_or0 ^ f_arrdiv24_fs75_xor0;
  assign f_arrdiv24_fs75_not1 = ~f_arrdiv24_fs75_xor0;
  assign f_arrdiv24_fs75_and1 = f_arrdiv24_fs75_not1 & f_arrdiv24_fs74_or0;
  assign f_arrdiv24_fs75_or0 = f_arrdiv24_fs75_and1 | f_arrdiv24_fs75_and0;
  assign f_arrdiv24_fs76_xor0 = f_arrdiv24_mux2to149_xor0 ^ b[4];
  assign f_arrdiv24_fs76_not0 = ~f_arrdiv24_mux2to149_xor0;
  assign f_arrdiv24_fs76_and0 = f_arrdiv24_fs76_not0 & b[4];
  assign f_arrdiv24_fs76_xor1 = f_arrdiv24_fs75_or0 ^ f_arrdiv24_fs76_xor0;
  assign f_arrdiv24_fs76_not1 = ~f_arrdiv24_fs76_xor0;
  assign f_arrdiv24_fs76_and1 = f_arrdiv24_fs76_not1 & f_arrdiv24_fs75_or0;
  assign f_arrdiv24_fs76_or0 = f_arrdiv24_fs76_and1 | f_arrdiv24_fs76_and0;
  assign f_arrdiv24_fs77_xor0 = f_arrdiv24_mux2to150_xor0 ^ b[5];
  assign f_arrdiv24_fs77_not0 = ~f_arrdiv24_mux2to150_xor0;
  assign f_arrdiv24_fs77_and0 = f_arrdiv24_fs77_not0 & b[5];
  assign f_arrdiv24_fs77_xor1 = f_arrdiv24_fs76_or0 ^ f_arrdiv24_fs77_xor0;
  assign f_arrdiv24_fs77_not1 = ~f_arrdiv24_fs77_xor0;
  assign f_arrdiv24_fs77_and1 = f_arrdiv24_fs77_not1 & f_arrdiv24_fs76_or0;
  assign f_arrdiv24_fs77_or0 = f_arrdiv24_fs77_and1 | f_arrdiv24_fs77_and0;
  assign f_arrdiv24_fs78_xor0 = f_arrdiv24_mux2to151_xor0 ^ b[6];
  assign f_arrdiv24_fs78_not0 = ~f_arrdiv24_mux2to151_xor0;
  assign f_arrdiv24_fs78_and0 = f_arrdiv24_fs78_not0 & b[6];
  assign f_arrdiv24_fs78_xor1 = f_arrdiv24_fs77_or0 ^ f_arrdiv24_fs78_xor0;
  assign f_arrdiv24_fs78_not1 = ~f_arrdiv24_fs78_xor0;
  assign f_arrdiv24_fs78_and1 = f_arrdiv24_fs78_not1 & f_arrdiv24_fs77_or0;
  assign f_arrdiv24_fs78_or0 = f_arrdiv24_fs78_and1 | f_arrdiv24_fs78_and0;
  assign f_arrdiv24_fs79_xor0 = f_arrdiv24_mux2to152_xor0 ^ b[7];
  assign f_arrdiv24_fs79_not0 = ~f_arrdiv24_mux2to152_xor0;
  assign f_arrdiv24_fs79_and0 = f_arrdiv24_fs79_not0 & b[7];
  assign f_arrdiv24_fs79_xor1 = f_arrdiv24_fs78_or0 ^ f_arrdiv24_fs79_xor0;
  assign f_arrdiv24_fs79_not1 = ~f_arrdiv24_fs79_xor0;
  assign f_arrdiv24_fs79_and1 = f_arrdiv24_fs79_not1 & f_arrdiv24_fs78_or0;
  assign f_arrdiv24_fs79_or0 = f_arrdiv24_fs79_and1 | f_arrdiv24_fs79_and0;
  assign f_arrdiv24_fs80_xor0 = f_arrdiv24_mux2to153_xor0 ^ b[8];
  assign f_arrdiv24_fs80_not0 = ~f_arrdiv24_mux2to153_xor0;
  assign f_arrdiv24_fs80_and0 = f_arrdiv24_fs80_not0 & b[8];
  assign f_arrdiv24_fs80_xor1 = f_arrdiv24_fs79_or0 ^ f_arrdiv24_fs80_xor0;
  assign f_arrdiv24_fs80_not1 = ~f_arrdiv24_fs80_xor0;
  assign f_arrdiv24_fs80_and1 = f_arrdiv24_fs80_not1 & f_arrdiv24_fs79_or0;
  assign f_arrdiv24_fs80_or0 = f_arrdiv24_fs80_and1 | f_arrdiv24_fs80_and0;
  assign f_arrdiv24_fs81_xor0 = f_arrdiv24_mux2to154_xor0 ^ b[9];
  assign f_arrdiv24_fs81_not0 = ~f_arrdiv24_mux2to154_xor0;
  assign f_arrdiv24_fs81_and0 = f_arrdiv24_fs81_not0 & b[9];
  assign f_arrdiv24_fs81_xor1 = f_arrdiv24_fs80_or0 ^ f_arrdiv24_fs81_xor0;
  assign f_arrdiv24_fs81_not1 = ~f_arrdiv24_fs81_xor0;
  assign f_arrdiv24_fs81_and1 = f_arrdiv24_fs81_not1 & f_arrdiv24_fs80_or0;
  assign f_arrdiv24_fs81_or0 = f_arrdiv24_fs81_and1 | f_arrdiv24_fs81_and0;
  assign f_arrdiv24_fs82_xor0 = f_arrdiv24_mux2to155_xor0 ^ b[10];
  assign f_arrdiv24_fs82_not0 = ~f_arrdiv24_mux2to155_xor0;
  assign f_arrdiv24_fs82_and0 = f_arrdiv24_fs82_not0 & b[10];
  assign f_arrdiv24_fs82_xor1 = f_arrdiv24_fs81_or0 ^ f_arrdiv24_fs82_xor0;
  assign f_arrdiv24_fs82_not1 = ~f_arrdiv24_fs82_xor0;
  assign f_arrdiv24_fs82_and1 = f_arrdiv24_fs82_not1 & f_arrdiv24_fs81_or0;
  assign f_arrdiv24_fs82_or0 = f_arrdiv24_fs82_and1 | f_arrdiv24_fs82_and0;
  assign f_arrdiv24_fs83_xor0 = f_arrdiv24_mux2to156_xor0 ^ b[11];
  assign f_arrdiv24_fs83_not0 = ~f_arrdiv24_mux2to156_xor0;
  assign f_arrdiv24_fs83_and0 = f_arrdiv24_fs83_not0 & b[11];
  assign f_arrdiv24_fs83_xor1 = f_arrdiv24_fs82_or0 ^ f_arrdiv24_fs83_xor0;
  assign f_arrdiv24_fs83_not1 = ~f_arrdiv24_fs83_xor0;
  assign f_arrdiv24_fs83_and1 = f_arrdiv24_fs83_not1 & f_arrdiv24_fs82_or0;
  assign f_arrdiv24_fs83_or0 = f_arrdiv24_fs83_and1 | f_arrdiv24_fs83_and0;
  assign f_arrdiv24_fs84_xor0 = f_arrdiv24_mux2to157_xor0 ^ b[12];
  assign f_arrdiv24_fs84_not0 = ~f_arrdiv24_mux2to157_xor0;
  assign f_arrdiv24_fs84_and0 = f_arrdiv24_fs84_not0 & b[12];
  assign f_arrdiv24_fs84_xor1 = f_arrdiv24_fs83_or0 ^ f_arrdiv24_fs84_xor0;
  assign f_arrdiv24_fs84_not1 = ~f_arrdiv24_fs84_xor0;
  assign f_arrdiv24_fs84_and1 = f_arrdiv24_fs84_not1 & f_arrdiv24_fs83_or0;
  assign f_arrdiv24_fs84_or0 = f_arrdiv24_fs84_and1 | f_arrdiv24_fs84_and0;
  assign f_arrdiv24_fs85_xor0 = f_arrdiv24_mux2to158_xor0 ^ b[13];
  assign f_arrdiv24_fs85_not0 = ~f_arrdiv24_mux2to158_xor0;
  assign f_arrdiv24_fs85_and0 = f_arrdiv24_fs85_not0 & b[13];
  assign f_arrdiv24_fs85_xor1 = f_arrdiv24_fs84_or0 ^ f_arrdiv24_fs85_xor0;
  assign f_arrdiv24_fs85_not1 = ~f_arrdiv24_fs85_xor0;
  assign f_arrdiv24_fs85_and1 = f_arrdiv24_fs85_not1 & f_arrdiv24_fs84_or0;
  assign f_arrdiv24_fs85_or0 = f_arrdiv24_fs85_and1 | f_arrdiv24_fs85_and0;
  assign f_arrdiv24_fs86_xor0 = f_arrdiv24_mux2to159_xor0 ^ b[14];
  assign f_arrdiv24_fs86_not0 = ~f_arrdiv24_mux2to159_xor0;
  assign f_arrdiv24_fs86_and0 = f_arrdiv24_fs86_not0 & b[14];
  assign f_arrdiv24_fs86_xor1 = f_arrdiv24_fs85_or0 ^ f_arrdiv24_fs86_xor0;
  assign f_arrdiv24_fs86_not1 = ~f_arrdiv24_fs86_xor0;
  assign f_arrdiv24_fs86_and1 = f_arrdiv24_fs86_not1 & f_arrdiv24_fs85_or0;
  assign f_arrdiv24_fs86_or0 = f_arrdiv24_fs86_and1 | f_arrdiv24_fs86_and0;
  assign f_arrdiv24_fs87_xor0 = f_arrdiv24_mux2to160_xor0 ^ b[15];
  assign f_arrdiv24_fs87_not0 = ~f_arrdiv24_mux2to160_xor0;
  assign f_arrdiv24_fs87_and0 = f_arrdiv24_fs87_not0 & b[15];
  assign f_arrdiv24_fs87_xor1 = f_arrdiv24_fs86_or0 ^ f_arrdiv24_fs87_xor0;
  assign f_arrdiv24_fs87_not1 = ~f_arrdiv24_fs87_xor0;
  assign f_arrdiv24_fs87_and1 = f_arrdiv24_fs87_not1 & f_arrdiv24_fs86_or0;
  assign f_arrdiv24_fs87_or0 = f_arrdiv24_fs87_and1 | f_arrdiv24_fs87_and0;
  assign f_arrdiv24_fs88_xor0 = f_arrdiv24_mux2to161_xor0 ^ b[16];
  assign f_arrdiv24_fs88_not0 = ~f_arrdiv24_mux2to161_xor0;
  assign f_arrdiv24_fs88_and0 = f_arrdiv24_fs88_not0 & b[16];
  assign f_arrdiv24_fs88_xor1 = f_arrdiv24_fs87_or0 ^ f_arrdiv24_fs88_xor0;
  assign f_arrdiv24_fs88_not1 = ~f_arrdiv24_fs88_xor0;
  assign f_arrdiv24_fs88_and1 = f_arrdiv24_fs88_not1 & f_arrdiv24_fs87_or0;
  assign f_arrdiv24_fs88_or0 = f_arrdiv24_fs88_and1 | f_arrdiv24_fs88_and0;
  assign f_arrdiv24_fs89_xor0 = f_arrdiv24_mux2to162_xor0 ^ b[17];
  assign f_arrdiv24_fs89_not0 = ~f_arrdiv24_mux2to162_xor0;
  assign f_arrdiv24_fs89_and0 = f_arrdiv24_fs89_not0 & b[17];
  assign f_arrdiv24_fs89_xor1 = f_arrdiv24_fs88_or0 ^ f_arrdiv24_fs89_xor0;
  assign f_arrdiv24_fs89_not1 = ~f_arrdiv24_fs89_xor0;
  assign f_arrdiv24_fs89_and1 = f_arrdiv24_fs89_not1 & f_arrdiv24_fs88_or0;
  assign f_arrdiv24_fs89_or0 = f_arrdiv24_fs89_and1 | f_arrdiv24_fs89_and0;
  assign f_arrdiv24_fs90_xor0 = f_arrdiv24_mux2to163_xor0 ^ b[18];
  assign f_arrdiv24_fs90_not0 = ~f_arrdiv24_mux2to163_xor0;
  assign f_arrdiv24_fs90_and0 = f_arrdiv24_fs90_not0 & b[18];
  assign f_arrdiv24_fs90_xor1 = f_arrdiv24_fs89_or0 ^ f_arrdiv24_fs90_xor0;
  assign f_arrdiv24_fs90_not1 = ~f_arrdiv24_fs90_xor0;
  assign f_arrdiv24_fs90_and1 = f_arrdiv24_fs90_not1 & f_arrdiv24_fs89_or0;
  assign f_arrdiv24_fs90_or0 = f_arrdiv24_fs90_and1 | f_arrdiv24_fs90_and0;
  assign f_arrdiv24_fs91_xor0 = f_arrdiv24_mux2to164_xor0 ^ b[19];
  assign f_arrdiv24_fs91_not0 = ~f_arrdiv24_mux2to164_xor0;
  assign f_arrdiv24_fs91_and0 = f_arrdiv24_fs91_not0 & b[19];
  assign f_arrdiv24_fs91_xor1 = f_arrdiv24_fs90_or0 ^ f_arrdiv24_fs91_xor0;
  assign f_arrdiv24_fs91_not1 = ~f_arrdiv24_fs91_xor0;
  assign f_arrdiv24_fs91_and1 = f_arrdiv24_fs91_not1 & f_arrdiv24_fs90_or0;
  assign f_arrdiv24_fs91_or0 = f_arrdiv24_fs91_and1 | f_arrdiv24_fs91_and0;
  assign f_arrdiv24_fs92_xor0 = f_arrdiv24_mux2to165_xor0 ^ b[20];
  assign f_arrdiv24_fs92_not0 = ~f_arrdiv24_mux2to165_xor0;
  assign f_arrdiv24_fs92_and0 = f_arrdiv24_fs92_not0 & b[20];
  assign f_arrdiv24_fs92_xor1 = f_arrdiv24_fs91_or0 ^ f_arrdiv24_fs92_xor0;
  assign f_arrdiv24_fs92_not1 = ~f_arrdiv24_fs92_xor0;
  assign f_arrdiv24_fs92_and1 = f_arrdiv24_fs92_not1 & f_arrdiv24_fs91_or0;
  assign f_arrdiv24_fs92_or0 = f_arrdiv24_fs92_and1 | f_arrdiv24_fs92_and0;
  assign f_arrdiv24_fs93_xor0 = f_arrdiv24_mux2to166_xor0 ^ b[21];
  assign f_arrdiv24_fs93_not0 = ~f_arrdiv24_mux2to166_xor0;
  assign f_arrdiv24_fs93_and0 = f_arrdiv24_fs93_not0 & b[21];
  assign f_arrdiv24_fs93_xor1 = f_arrdiv24_fs92_or0 ^ f_arrdiv24_fs93_xor0;
  assign f_arrdiv24_fs93_not1 = ~f_arrdiv24_fs93_xor0;
  assign f_arrdiv24_fs93_and1 = f_arrdiv24_fs93_not1 & f_arrdiv24_fs92_or0;
  assign f_arrdiv24_fs93_or0 = f_arrdiv24_fs93_and1 | f_arrdiv24_fs93_and0;
  assign f_arrdiv24_fs94_xor0 = f_arrdiv24_mux2to167_xor0 ^ b[22];
  assign f_arrdiv24_fs94_not0 = ~f_arrdiv24_mux2to167_xor0;
  assign f_arrdiv24_fs94_and0 = f_arrdiv24_fs94_not0 & b[22];
  assign f_arrdiv24_fs94_xor1 = f_arrdiv24_fs93_or0 ^ f_arrdiv24_fs94_xor0;
  assign f_arrdiv24_fs94_not1 = ~f_arrdiv24_fs94_xor0;
  assign f_arrdiv24_fs94_and1 = f_arrdiv24_fs94_not1 & f_arrdiv24_fs93_or0;
  assign f_arrdiv24_fs94_or0 = f_arrdiv24_fs94_and1 | f_arrdiv24_fs94_and0;
  assign f_arrdiv24_fs95_xor0 = f_arrdiv24_mux2to168_xor0 ^ b[23];
  assign f_arrdiv24_fs95_not0 = ~f_arrdiv24_mux2to168_xor0;
  assign f_arrdiv24_fs95_and0 = f_arrdiv24_fs95_not0 & b[23];
  assign f_arrdiv24_fs95_xor1 = f_arrdiv24_fs94_or0 ^ f_arrdiv24_fs95_xor0;
  assign f_arrdiv24_fs95_not1 = ~f_arrdiv24_fs95_xor0;
  assign f_arrdiv24_fs95_and1 = f_arrdiv24_fs95_not1 & f_arrdiv24_fs94_or0;
  assign f_arrdiv24_fs95_or0 = f_arrdiv24_fs95_and1 | f_arrdiv24_fs95_and0;
  assign f_arrdiv24_mux2to169_and0 = a[20] & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to169_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to169_and1 = f_arrdiv24_fs72_xor0 & f_arrdiv24_mux2to169_not0;
  assign f_arrdiv24_mux2to169_xor0 = f_arrdiv24_mux2to169_and0 ^ f_arrdiv24_mux2to169_and1;
  assign f_arrdiv24_mux2to170_and0 = f_arrdiv24_mux2to146_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to170_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to170_and1 = f_arrdiv24_fs73_xor1 & f_arrdiv24_mux2to170_not0;
  assign f_arrdiv24_mux2to170_xor0 = f_arrdiv24_mux2to170_and0 ^ f_arrdiv24_mux2to170_and1;
  assign f_arrdiv24_mux2to171_and0 = f_arrdiv24_mux2to147_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to171_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to171_and1 = f_arrdiv24_fs74_xor1 & f_arrdiv24_mux2to171_not0;
  assign f_arrdiv24_mux2to171_xor0 = f_arrdiv24_mux2to171_and0 ^ f_arrdiv24_mux2to171_and1;
  assign f_arrdiv24_mux2to172_and0 = f_arrdiv24_mux2to148_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to172_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to172_and1 = f_arrdiv24_fs75_xor1 & f_arrdiv24_mux2to172_not0;
  assign f_arrdiv24_mux2to172_xor0 = f_arrdiv24_mux2to172_and0 ^ f_arrdiv24_mux2to172_and1;
  assign f_arrdiv24_mux2to173_and0 = f_arrdiv24_mux2to149_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to173_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to173_and1 = f_arrdiv24_fs76_xor1 & f_arrdiv24_mux2to173_not0;
  assign f_arrdiv24_mux2to173_xor0 = f_arrdiv24_mux2to173_and0 ^ f_arrdiv24_mux2to173_and1;
  assign f_arrdiv24_mux2to174_and0 = f_arrdiv24_mux2to150_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to174_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to174_and1 = f_arrdiv24_fs77_xor1 & f_arrdiv24_mux2to174_not0;
  assign f_arrdiv24_mux2to174_xor0 = f_arrdiv24_mux2to174_and0 ^ f_arrdiv24_mux2to174_and1;
  assign f_arrdiv24_mux2to175_and0 = f_arrdiv24_mux2to151_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to175_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to175_and1 = f_arrdiv24_fs78_xor1 & f_arrdiv24_mux2to175_not0;
  assign f_arrdiv24_mux2to175_xor0 = f_arrdiv24_mux2to175_and0 ^ f_arrdiv24_mux2to175_and1;
  assign f_arrdiv24_mux2to176_and0 = f_arrdiv24_mux2to152_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to176_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to176_and1 = f_arrdiv24_fs79_xor1 & f_arrdiv24_mux2to176_not0;
  assign f_arrdiv24_mux2to176_xor0 = f_arrdiv24_mux2to176_and0 ^ f_arrdiv24_mux2to176_and1;
  assign f_arrdiv24_mux2to177_and0 = f_arrdiv24_mux2to153_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to177_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to177_and1 = f_arrdiv24_fs80_xor1 & f_arrdiv24_mux2to177_not0;
  assign f_arrdiv24_mux2to177_xor0 = f_arrdiv24_mux2to177_and0 ^ f_arrdiv24_mux2to177_and1;
  assign f_arrdiv24_mux2to178_and0 = f_arrdiv24_mux2to154_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to178_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to178_and1 = f_arrdiv24_fs81_xor1 & f_arrdiv24_mux2to178_not0;
  assign f_arrdiv24_mux2to178_xor0 = f_arrdiv24_mux2to178_and0 ^ f_arrdiv24_mux2to178_and1;
  assign f_arrdiv24_mux2to179_and0 = f_arrdiv24_mux2to155_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to179_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to179_and1 = f_arrdiv24_fs82_xor1 & f_arrdiv24_mux2to179_not0;
  assign f_arrdiv24_mux2to179_xor0 = f_arrdiv24_mux2to179_and0 ^ f_arrdiv24_mux2to179_and1;
  assign f_arrdiv24_mux2to180_and0 = f_arrdiv24_mux2to156_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to180_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to180_and1 = f_arrdiv24_fs83_xor1 & f_arrdiv24_mux2to180_not0;
  assign f_arrdiv24_mux2to180_xor0 = f_arrdiv24_mux2to180_and0 ^ f_arrdiv24_mux2to180_and1;
  assign f_arrdiv24_mux2to181_and0 = f_arrdiv24_mux2to157_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to181_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to181_and1 = f_arrdiv24_fs84_xor1 & f_arrdiv24_mux2to181_not0;
  assign f_arrdiv24_mux2to181_xor0 = f_arrdiv24_mux2to181_and0 ^ f_arrdiv24_mux2to181_and1;
  assign f_arrdiv24_mux2to182_and0 = f_arrdiv24_mux2to158_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to182_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to182_and1 = f_arrdiv24_fs85_xor1 & f_arrdiv24_mux2to182_not0;
  assign f_arrdiv24_mux2to182_xor0 = f_arrdiv24_mux2to182_and0 ^ f_arrdiv24_mux2to182_and1;
  assign f_arrdiv24_mux2to183_and0 = f_arrdiv24_mux2to159_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to183_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to183_and1 = f_arrdiv24_fs86_xor1 & f_arrdiv24_mux2to183_not0;
  assign f_arrdiv24_mux2to183_xor0 = f_arrdiv24_mux2to183_and0 ^ f_arrdiv24_mux2to183_and1;
  assign f_arrdiv24_mux2to184_and0 = f_arrdiv24_mux2to160_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to184_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to184_and1 = f_arrdiv24_fs87_xor1 & f_arrdiv24_mux2to184_not0;
  assign f_arrdiv24_mux2to184_xor0 = f_arrdiv24_mux2to184_and0 ^ f_arrdiv24_mux2to184_and1;
  assign f_arrdiv24_mux2to185_and0 = f_arrdiv24_mux2to161_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to185_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to185_and1 = f_arrdiv24_fs88_xor1 & f_arrdiv24_mux2to185_not0;
  assign f_arrdiv24_mux2to185_xor0 = f_arrdiv24_mux2to185_and0 ^ f_arrdiv24_mux2to185_and1;
  assign f_arrdiv24_mux2to186_and0 = f_arrdiv24_mux2to162_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to186_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to186_and1 = f_arrdiv24_fs89_xor1 & f_arrdiv24_mux2to186_not0;
  assign f_arrdiv24_mux2to186_xor0 = f_arrdiv24_mux2to186_and0 ^ f_arrdiv24_mux2to186_and1;
  assign f_arrdiv24_mux2to187_and0 = f_arrdiv24_mux2to163_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to187_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to187_and1 = f_arrdiv24_fs90_xor1 & f_arrdiv24_mux2to187_not0;
  assign f_arrdiv24_mux2to187_xor0 = f_arrdiv24_mux2to187_and0 ^ f_arrdiv24_mux2to187_and1;
  assign f_arrdiv24_mux2to188_and0 = f_arrdiv24_mux2to164_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to188_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to188_and1 = f_arrdiv24_fs91_xor1 & f_arrdiv24_mux2to188_not0;
  assign f_arrdiv24_mux2to188_xor0 = f_arrdiv24_mux2to188_and0 ^ f_arrdiv24_mux2to188_and1;
  assign f_arrdiv24_mux2to189_and0 = f_arrdiv24_mux2to165_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to189_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to189_and1 = f_arrdiv24_fs92_xor1 & f_arrdiv24_mux2to189_not0;
  assign f_arrdiv24_mux2to189_xor0 = f_arrdiv24_mux2to189_and0 ^ f_arrdiv24_mux2to189_and1;
  assign f_arrdiv24_mux2to190_and0 = f_arrdiv24_mux2to166_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to190_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to190_and1 = f_arrdiv24_fs93_xor1 & f_arrdiv24_mux2to190_not0;
  assign f_arrdiv24_mux2to190_xor0 = f_arrdiv24_mux2to190_and0 ^ f_arrdiv24_mux2to190_and1;
  assign f_arrdiv24_mux2to191_and0 = f_arrdiv24_mux2to167_xor0 & f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to191_not0 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_mux2to191_and1 = f_arrdiv24_fs94_xor1 & f_arrdiv24_mux2to191_not0;
  assign f_arrdiv24_mux2to191_xor0 = f_arrdiv24_mux2to191_and0 ^ f_arrdiv24_mux2to191_and1;
  assign f_arrdiv24_not3 = ~f_arrdiv24_fs95_or0;
  assign f_arrdiv24_fs96_xor0 = a[19] ^ b[0];
  assign f_arrdiv24_fs96_not0 = ~a[19];
  assign f_arrdiv24_fs96_and0 = f_arrdiv24_fs96_not0 & b[0];
  assign f_arrdiv24_fs96_not1 = ~f_arrdiv24_fs96_xor0;
  assign f_arrdiv24_fs97_xor0 = f_arrdiv24_mux2to169_xor0 ^ b[1];
  assign f_arrdiv24_fs97_not0 = ~f_arrdiv24_mux2to169_xor0;
  assign f_arrdiv24_fs97_and0 = f_arrdiv24_fs97_not0 & b[1];
  assign f_arrdiv24_fs97_xor1 = f_arrdiv24_fs96_and0 ^ f_arrdiv24_fs97_xor0;
  assign f_arrdiv24_fs97_not1 = ~f_arrdiv24_fs97_xor0;
  assign f_arrdiv24_fs97_and1 = f_arrdiv24_fs97_not1 & f_arrdiv24_fs96_and0;
  assign f_arrdiv24_fs97_or0 = f_arrdiv24_fs97_and1 | f_arrdiv24_fs97_and0;
  assign f_arrdiv24_fs98_xor0 = f_arrdiv24_mux2to170_xor0 ^ b[2];
  assign f_arrdiv24_fs98_not0 = ~f_arrdiv24_mux2to170_xor0;
  assign f_arrdiv24_fs98_and0 = f_arrdiv24_fs98_not0 & b[2];
  assign f_arrdiv24_fs98_xor1 = f_arrdiv24_fs97_or0 ^ f_arrdiv24_fs98_xor0;
  assign f_arrdiv24_fs98_not1 = ~f_arrdiv24_fs98_xor0;
  assign f_arrdiv24_fs98_and1 = f_arrdiv24_fs98_not1 & f_arrdiv24_fs97_or0;
  assign f_arrdiv24_fs98_or0 = f_arrdiv24_fs98_and1 | f_arrdiv24_fs98_and0;
  assign f_arrdiv24_fs99_xor0 = f_arrdiv24_mux2to171_xor0 ^ b[3];
  assign f_arrdiv24_fs99_not0 = ~f_arrdiv24_mux2to171_xor0;
  assign f_arrdiv24_fs99_and0 = f_arrdiv24_fs99_not0 & b[3];
  assign f_arrdiv24_fs99_xor1 = f_arrdiv24_fs98_or0 ^ f_arrdiv24_fs99_xor0;
  assign f_arrdiv24_fs99_not1 = ~f_arrdiv24_fs99_xor0;
  assign f_arrdiv24_fs99_and1 = f_arrdiv24_fs99_not1 & f_arrdiv24_fs98_or0;
  assign f_arrdiv24_fs99_or0 = f_arrdiv24_fs99_and1 | f_arrdiv24_fs99_and0;
  assign f_arrdiv24_fs100_xor0 = f_arrdiv24_mux2to172_xor0 ^ b[4];
  assign f_arrdiv24_fs100_not0 = ~f_arrdiv24_mux2to172_xor0;
  assign f_arrdiv24_fs100_and0 = f_arrdiv24_fs100_not0 & b[4];
  assign f_arrdiv24_fs100_xor1 = f_arrdiv24_fs99_or0 ^ f_arrdiv24_fs100_xor0;
  assign f_arrdiv24_fs100_not1 = ~f_arrdiv24_fs100_xor0;
  assign f_arrdiv24_fs100_and1 = f_arrdiv24_fs100_not1 & f_arrdiv24_fs99_or0;
  assign f_arrdiv24_fs100_or0 = f_arrdiv24_fs100_and1 | f_arrdiv24_fs100_and0;
  assign f_arrdiv24_fs101_xor0 = f_arrdiv24_mux2to173_xor0 ^ b[5];
  assign f_arrdiv24_fs101_not0 = ~f_arrdiv24_mux2to173_xor0;
  assign f_arrdiv24_fs101_and0 = f_arrdiv24_fs101_not0 & b[5];
  assign f_arrdiv24_fs101_xor1 = f_arrdiv24_fs100_or0 ^ f_arrdiv24_fs101_xor0;
  assign f_arrdiv24_fs101_not1 = ~f_arrdiv24_fs101_xor0;
  assign f_arrdiv24_fs101_and1 = f_arrdiv24_fs101_not1 & f_arrdiv24_fs100_or0;
  assign f_arrdiv24_fs101_or0 = f_arrdiv24_fs101_and1 | f_arrdiv24_fs101_and0;
  assign f_arrdiv24_fs102_xor0 = f_arrdiv24_mux2to174_xor0 ^ b[6];
  assign f_arrdiv24_fs102_not0 = ~f_arrdiv24_mux2to174_xor0;
  assign f_arrdiv24_fs102_and0 = f_arrdiv24_fs102_not0 & b[6];
  assign f_arrdiv24_fs102_xor1 = f_arrdiv24_fs101_or0 ^ f_arrdiv24_fs102_xor0;
  assign f_arrdiv24_fs102_not1 = ~f_arrdiv24_fs102_xor0;
  assign f_arrdiv24_fs102_and1 = f_arrdiv24_fs102_not1 & f_arrdiv24_fs101_or0;
  assign f_arrdiv24_fs102_or0 = f_arrdiv24_fs102_and1 | f_arrdiv24_fs102_and0;
  assign f_arrdiv24_fs103_xor0 = f_arrdiv24_mux2to175_xor0 ^ b[7];
  assign f_arrdiv24_fs103_not0 = ~f_arrdiv24_mux2to175_xor0;
  assign f_arrdiv24_fs103_and0 = f_arrdiv24_fs103_not0 & b[7];
  assign f_arrdiv24_fs103_xor1 = f_arrdiv24_fs102_or0 ^ f_arrdiv24_fs103_xor0;
  assign f_arrdiv24_fs103_not1 = ~f_arrdiv24_fs103_xor0;
  assign f_arrdiv24_fs103_and1 = f_arrdiv24_fs103_not1 & f_arrdiv24_fs102_or0;
  assign f_arrdiv24_fs103_or0 = f_arrdiv24_fs103_and1 | f_arrdiv24_fs103_and0;
  assign f_arrdiv24_fs104_xor0 = f_arrdiv24_mux2to176_xor0 ^ b[8];
  assign f_arrdiv24_fs104_not0 = ~f_arrdiv24_mux2to176_xor0;
  assign f_arrdiv24_fs104_and0 = f_arrdiv24_fs104_not0 & b[8];
  assign f_arrdiv24_fs104_xor1 = f_arrdiv24_fs103_or0 ^ f_arrdiv24_fs104_xor0;
  assign f_arrdiv24_fs104_not1 = ~f_arrdiv24_fs104_xor0;
  assign f_arrdiv24_fs104_and1 = f_arrdiv24_fs104_not1 & f_arrdiv24_fs103_or0;
  assign f_arrdiv24_fs104_or0 = f_arrdiv24_fs104_and1 | f_arrdiv24_fs104_and0;
  assign f_arrdiv24_fs105_xor0 = f_arrdiv24_mux2to177_xor0 ^ b[9];
  assign f_arrdiv24_fs105_not0 = ~f_arrdiv24_mux2to177_xor0;
  assign f_arrdiv24_fs105_and0 = f_arrdiv24_fs105_not0 & b[9];
  assign f_arrdiv24_fs105_xor1 = f_arrdiv24_fs104_or0 ^ f_arrdiv24_fs105_xor0;
  assign f_arrdiv24_fs105_not1 = ~f_arrdiv24_fs105_xor0;
  assign f_arrdiv24_fs105_and1 = f_arrdiv24_fs105_not1 & f_arrdiv24_fs104_or0;
  assign f_arrdiv24_fs105_or0 = f_arrdiv24_fs105_and1 | f_arrdiv24_fs105_and0;
  assign f_arrdiv24_fs106_xor0 = f_arrdiv24_mux2to178_xor0 ^ b[10];
  assign f_arrdiv24_fs106_not0 = ~f_arrdiv24_mux2to178_xor0;
  assign f_arrdiv24_fs106_and0 = f_arrdiv24_fs106_not0 & b[10];
  assign f_arrdiv24_fs106_xor1 = f_arrdiv24_fs105_or0 ^ f_arrdiv24_fs106_xor0;
  assign f_arrdiv24_fs106_not1 = ~f_arrdiv24_fs106_xor0;
  assign f_arrdiv24_fs106_and1 = f_arrdiv24_fs106_not1 & f_arrdiv24_fs105_or0;
  assign f_arrdiv24_fs106_or0 = f_arrdiv24_fs106_and1 | f_arrdiv24_fs106_and0;
  assign f_arrdiv24_fs107_xor0 = f_arrdiv24_mux2to179_xor0 ^ b[11];
  assign f_arrdiv24_fs107_not0 = ~f_arrdiv24_mux2to179_xor0;
  assign f_arrdiv24_fs107_and0 = f_arrdiv24_fs107_not0 & b[11];
  assign f_arrdiv24_fs107_xor1 = f_arrdiv24_fs106_or0 ^ f_arrdiv24_fs107_xor0;
  assign f_arrdiv24_fs107_not1 = ~f_arrdiv24_fs107_xor0;
  assign f_arrdiv24_fs107_and1 = f_arrdiv24_fs107_not1 & f_arrdiv24_fs106_or0;
  assign f_arrdiv24_fs107_or0 = f_arrdiv24_fs107_and1 | f_arrdiv24_fs107_and0;
  assign f_arrdiv24_fs108_xor0 = f_arrdiv24_mux2to180_xor0 ^ b[12];
  assign f_arrdiv24_fs108_not0 = ~f_arrdiv24_mux2to180_xor0;
  assign f_arrdiv24_fs108_and0 = f_arrdiv24_fs108_not0 & b[12];
  assign f_arrdiv24_fs108_xor1 = f_arrdiv24_fs107_or0 ^ f_arrdiv24_fs108_xor0;
  assign f_arrdiv24_fs108_not1 = ~f_arrdiv24_fs108_xor0;
  assign f_arrdiv24_fs108_and1 = f_arrdiv24_fs108_not1 & f_arrdiv24_fs107_or0;
  assign f_arrdiv24_fs108_or0 = f_arrdiv24_fs108_and1 | f_arrdiv24_fs108_and0;
  assign f_arrdiv24_fs109_xor0 = f_arrdiv24_mux2to181_xor0 ^ b[13];
  assign f_arrdiv24_fs109_not0 = ~f_arrdiv24_mux2to181_xor0;
  assign f_arrdiv24_fs109_and0 = f_arrdiv24_fs109_not0 & b[13];
  assign f_arrdiv24_fs109_xor1 = f_arrdiv24_fs108_or0 ^ f_arrdiv24_fs109_xor0;
  assign f_arrdiv24_fs109_not1 = ~f_arrdiv24_fs109_xor0;
  assign f_arrdiv24_fs109_and1 = f_arrdiv24_fs109_not1 & f_arrdiv24_fs108_or0;
  assign f_arrdiv24_fs109_or0 = f_arrdiv24_fs109_and1 | f_arrdiv24_fs109_and0;
  assign f_arrdiv24_fs110_xor0 = f_arrdiv24_mux2to182_xor0 ^ b[14];
  assign f_arrdiv24_fs110_not0 = ~f_arrdiv24_mux2to182_xor0;
  assign f_arrdiv24_fs110_and0 = f_arrdiv24_fs110_not0 & b[14];
  assign f_arrdiv24_fs110_xor1 = f_arrdiv24_fs109_or0 ^ f_arrdiv24_fs110_xor0;
  assign f_arrdiv24_fs110_not1 = ~f_arrdiv24_fs110_xor0;
  assign f_arrdiv24_fs110_and1 = f_arrdiv24_fs110_not1 & f_arrdiv24_fs109_or0;
  assign f_arrdiv24_fs110_or0 = f_arrdiv24_fs110_and1 | f_arrdiv24_fs110_and0;
  assign f_arrdiv24_fs111_xor0 = f_arrdiv24_mux2to183_xor0 ^ b[15];
  assign f_arrdiv24_fs111_not0 = ~f_arrdiv24_mux2to183_xor0;
  assign f_arrdiv24_fs111_and0 = f_arrdiv24_fs111_not0 & b[15];
  assign f_arrdiv24_fs111_xor1 = f_arrdiv24_fs110_or0 ^ f_arrdiv24_fs111_xor0;
  assign f_arrdiv24_fs111_not1 = ~f_arrdiv24_fs111_xor0;
  assign f_arrdiv24_fs111_and1 = f_arrdiv24_fs111_not1 & f_arrdiv24_fs110_or0;
  assign f_arrdiv24_fs111_or0 = f_arrdiv24_fs111_and1 | f_arrdiv24_fs111_and0;
  assign f_arrdiv24_fs112_xor0 = f_arrdiv24_mux2to184_xor0 ^ b[16];
  assign f_arrdiv24_fs112_not0 = ~f_arrdiv24_mux2to184_xor0;
  assign f_arrdiv24_fs112_and0 = f_arrdiv24_fs112_not0 & b[16];
  assign f_arrdiv24_fs112_xor1 = f_arrdiv24_fs111_or0 ^ f_arrdiv24_fs112_xor0;
  assign f_arrdiv24_fs112_not1 = ~f_arrdiv24_fs112_xor0;
  assign f_arrdiv24_fs112_and1 = f_arrdiv24_fs112_not1 & f_arrdiv24_fs111_or0;
  assign f_arrdiv24_fs112_or0 = f_arrdiv24_fs112_and1 | f_arrdiv24_fs112_and0;
  assign f_arrdiv24_fs113_xor0 = f_arrdiv24_mux2to185_xor0 ^ b[17];
  assign f_arrdiv24_fs113_not0 = ~f_arrdiv24_mux2to185_xor0;
  assign f_arrdiv24_fs113_and0 = f_arrdiv24_fs113_not0 & b[17];
  assign f_arrdiv24_fs113_xor1 = f_arrdiv24_fs112_or0 ^ f_arrdiv24_fs113_xor0;
  assign f_arrdiv24_fs113_not1 = ~f_arrdiv24_fs113_xor0;
  assign f_arrdiv24_fs113_and1 = f_arrdiv24_fs113_not1 & f_arrdiv24_fs112_or0;
  assign f_arrdiv24_fs113_or0 = f_arrdiv24_fs113_and1 | f_arrdiv24_fs113_and0;
  assign f_arrdiv24_fs114_xor0 = f_arrdiv24_mux2to186_xor0 ^ b[18];
  assign f_arrdiv24_fs114_not0 = ~f_arrdiv24_mux2to186_xor0;
  assign f_arrdiv24_fs114_and0 = f_arrdiv24_fs114_not0 & b[18];
  assign f_arrdiv24_fs114_xor1 = f_arrdiv24_fs113_or0 ^ f_arrdiv24_fs114_xor0;
  assign f_arrdiv24_fs114_not1 = ~f_arrdiv24_fs114_xor0;
  assign f_arrdiv24_fs114_and1 = f_arrdiv24_fs114_not1 & f_arrdiv24_fs113_or0;
  assign f_arrdiv24_fs114_or0 = f_arrdiv24_fs114_and1 | f_arrdiv24_fs114_and0;
  assign f_arrdiv24_fs115_xor0 = f_arrdiv24_mux2to187_xor0 ^ b[19];
  assign f_arrdiv24_fs115_not0 = ~f_arrdiv24_mux2to187_xor0;
  assign f_arrdiv24_fs115_and0 = f_arrdiv24_fs115_not0 & b[19];
  assign f_arrdiv24_fs115_xor1 = f_arrdiv24_fs114_or0 ^ f_arrdiv24_fs115_xor0;
  assign f_arrdiv24_fs115_not1 = ~f_arrdiv24_fs115_xor0;
  assign f_arrdiv24_fs115_and1 = f_arrdiv24_fs115_not1 & f_arrdiv24_fs114_or0;
  assign f_arrdiv24_fs115_or0 = f_arrdiv24_fs115_and1 | f_arrdiv24_fs115_and0;
  assign f_arrdiv24_fs116_xor0 = f_arrdiv24_mux2to188_xor0 ^ b[20];
  assign f_arrdiv24_fs116_not0 = ~f_arrdiv24_mux2to188_xor0;
  assign f_arrdiv24_fs116_and0 = f_arrdiv24_fs116_not0 & b[20];
  assign f_arrdiv24_fs116_xor1 = f_arrdiv24_fs115_or0 ^ f_arrdiv24_fs116_xor0;
  assign f_arrdiv24_fs116_not1 = ~f_arrdiv24_fs116_xor0;
  assign f_arrdiv24_fs116_and1 = f_arrdiv24_fs116_not1 & f_arrdiv24_fs115_or0;
  assign f_arrdiv24_fs116_or0 = f_arrdiv24_fs116_and1 | f_arrdiv24_fs116_and0;
  assign f_arrdiv24_fs117_xor0 = f_arrdiv24_mux2to189_xor0 ^ b[21];
  assign f_arrdiv24_fs117_not0 = ~f_arrdiv24_mux2to189_xor0;
  assign f_arrdiv24_fs117_and0 = f_arrdiv24_fs117_not0 & b[21];
  assign f_arrdiv24_fs117_xor1 = f_arrdiv24_fs116_or0 ^ f_arrdiv24_fs117_xor0;
  assign f_arrdiv24_fs117_not1 = ~f_arrdiv24_fs117_xor0;
  assign f_arrdiv24_fs117_and1 = f_arrdiv24_fs117_not1 & f_arrdiv24_fs116_or0;
  assign f_arrdiv24_fs117_or0 = f_arrdiv24_fs117_and1 | f_arrdiv24_fs117_and0;
  assign f_arrdiv24_fs118_xor0 = f_arrdiv24_mux2to190_xor0 ^ b[22];
  assign f_arrdiv24_fs118_not0 = ~f_arrdiv24_mux2to190_xor0;
  assign f_arrdiv24_fs118_and0 = f_arrdiv24_fs118_not0 & b[22];
  assign f_arrdiv24_fs118_xor1 = f_arrdiv24_fs117_or0 ^ f_arrdiv24_fs118_xor0;
  assign f_arrdiv24_fs118_not1 = ~f_arrdiv24_fs118_xor0;
  assign f_arrdiv24_fs118_and1 = f_arrdiv24_fs118_not1 & f_arrdiv24_fs117_or0;
  assign f_arrdiv24_fs118_or0 = f_arrdiv24_fs118_and1 | f_arrdiv24_fs118_and0;
  assign f_arrdiv24_fs119_xor0 = f_arrdiv24_mux2to191_xor0 ^ b[23];
  assign f_arrdiv24_fs119_not0 = ~f_arrdiv24_mux2to191_xor0;
  assign f_arrdiv24_fs119_and0 = f_arrdiv24_fs119_not0 & b[23];
  assign f_arrdiv24_fs119_xor1 = f_arrdiv24_fs118_or0 ^ f_arrdiv24_fs119_xor0;
  assign f_arrdiv24_fs119_not1 = ~f_arrdiv24_fs119_xor0;
  assign f_arrdiv24_fs119_and1 = f_arrdiv24_fs119_not1 & f_arrdiv24_fs118_or0;
  assign f_arrdiv24_fs119_or0 = f_arrdiv24_fs119_and1 | f_arrdiv24_fs119_and0;
  assign f_arrdiv24_mux2to192_and0 = a[19] & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to192_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to192_and1 = f_arrdiv24_fs96_xor0 & f_arrdiv24_mux2to192_not0;
  assign f_arrdiv24_mux2to192_xor0 = f_arrdiv24_mux2to192_and0 ^ f_arrdiv24_mux2to192_and1;
  assign f_arrdiv24_mux2to193_and0 = f_arrdiv24_mux2to169_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to193_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to193_and1 = f_arrdiv24_fs97_xor1 & f_arrdiv24_mux2to193_not0;
  assign f_arrdiv24_mux2to193_xor0 = f_arrdiv24_mux2to193_and0 ^ f_arrdiv24_mux2to193_and1;
  assign f_arrdiv24_mux2to194_and0 = f_arrdiv24_mux2to170_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to194_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to194_and1 = f_arrdiv24_fs98_xor1 & f_arrdiv24_mux2to194_not0;
  assign f_arrdiv24_mux2to194_xor0 = f_arrdiv24_mux2to194_and0 ^ f_arrdiv24_mux2to194_and1;
  assign f_arrdiv24_mux2to195_and0 = f_arrdiv24_mux2to171_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to195_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to195_and1 = f_arrdiv24_fs99_xor1 & f_arrdiv24_mux2to195_not0;
  assign f_arrdiv24_mux2to195_xor0 = f_arrdiv24_mux2to195_and0 ^ f_arrdiv24_mux2to195_and1;
  assign f_arrdiv24_mux2to196_and0 = f_arrdiv24_mux2to172_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to196_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to196_and1 = f_arrdiv24_fs100_xor1 & f_arrdiv24_mux2to196_not0;
  assign f_arrdiv24_mux2to196_xor0 = f_arrdiv24_mux2to196_and0 ^ f_arrdiv24_mux2to196_and1;
  assign f_arrdiv24_mux2to197_and0 = f_arrdiv24_mux2to173_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to197_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to197_and1 = f_arrdiv24_fs101_xor1 & f_arrdiv24_mux2to197_not0;
  assign f_arrdiv24_mux2to197_xor0 = f_arrdiv24_mux2to197_and0 ^ f_arrdiv24_mux2to197_and1;
  assign f_arrdiv24_mux2to198_and0 = f_arrdiv24_mux2to174_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to198_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to198_and1 = f_arrdiv24_fs102_xor1 & f_arrdiv24_mux2to198_not0;
  assign f_arrdiv24_mux2to198_xor0 = f_arrdiv24_mux2to198_and0 ^ f_arrdiv24_mux2to198_and1;
  assign f_arrdiv24_mux2to199_and0 = f_arrdiv24_mux2to175_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to199_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to199_and1 = f_arrdiv24_fs103_xor1 & f_arrdiv24_mux2to199_not0;
  assign f_arrdiv24_mux2to199_xor0 = f_arrdiv24_mux2to199_and0 ^ f_arrdiv24_mux2to199_and1;
  assign f_arrdiv24_mux2to1100_and0 = f_arrdiv24_mux2to176_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1100_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1100_and1 = f_arrdiv24_fs104_xor1 & f_arrdiv24_mux2to1100_not0;
  assign f_arrdiv24_mux2to1100_xor0 = f_arrdiv24_mux2to1100_and0 ^ f_arrdiv24_mux2to1100_and1;
  assign f_arrdiv24_mux2to1101_and0 = f_arrdiv24_mux2to177_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1101_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1101_and1 = f_arrdiv24_fs105_xor1 & f_arrdiv24_mux2to1101_not0;
  assign f_arrdiv24_mux2to1101_xor0 = f_arrdiv24_mux2to1101_and0 ^ f_arrdiv24_mux2to1101_and1;
  assign f_arrdiv24_mux2to1102_and0 = f_arrdiv24_mux2to178_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1102_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1102_and1 = f_arrdiv24_fs106_xor1 & f_arrdiv24_mux2to1102_not0;
  assign f_arrdiv24_mux2to1102_xor0 = f_arrdiv24_mux2to1102_and0 ^ f_arrdiv24_mux2to1102_and1;
  assign f_arrdiv24_mux2to1103_and0 = f_arrdiv24_mux2to179_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1103_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1103_and1 = f_arrdiv24_fs107_xor1 & f_arrdiv24_mux2to1103_not0;
  assign f_arrdiv24_mux2to1103_xor0 = f_arrdiv24_mux2to1103_and0 ^ f_arrdiv24_mux2to1103_and1;
  assign f_arrdiv24_mux2to1104_and0 = f_arrdiv24_mux2to180_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1104_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1104_and1 = f_arrdiv24_fs108_xor1 & f_arrdiv24_mux2to1104_not0;
  assign f_arrdiv24_mux2to1104_xor0 = f_arrdiv24_mux2to1104_and0 ^ f_arrdiv24_mux2to1104_and1;
  assign f_arrdiv24_mux2to1105_and0 = f_arrdiv24_mux2to181_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1105_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1105_and1 = f_arrdiv24_fs109_xor1 & f_arrdiv24_mux2to1105_not0;
  assign f_arrdiv24_mux2to1105_xor0 = f_arrdiv24_mux2to1105_and0 ^ f_arrdiv24_mux2to1105_and1;
  assign f_arrdiv24_mux2to1106_and0 = f_arrdiv24_mux2to182_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1106_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1106_and1 = f_arrdiv24_fs110_xor1 & f_arrdiv24_mux2to1106_not0;
  assign f_arrdiv24_mux2to1106_xor0 = f_arrdiv24_mux2to1106_and0 ^ f_arrdiv24_mux2to1106_and1;
  assign f_arrdiv24_mux2to1107_and0 = f_arrdiv24_mux2to183_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1107_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1107_and1 = f_arrdiv24_fs111_xor1 & f_arrdiv24_mux2to1107_not0;
  assign f_arrdiv24_mux2to1107_xor0 = f_arrdiv24_mux2to1107_and0 ^ f_arrdiv24_mux2to1107_and1;
  assign f_arrdiv24_mux2to1108_and0 = f_arrdiv24_mux2to184_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1108_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1108_and1 = f_arrdiv24_fs112_xor1 & f_arrdiv24_mux2to1108_not0;
  assign f_arrdiv24_mux2to1108_xor0 = f_arrdiv24_mux2to1108_and0 ^ f_arrdiv24_mux2to1108_and1;
  assign f_arrdiv24_mux2to1109_and0 = f_arrdiv24_mux2to185_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1109_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1109_and1 = f_arrdiv24_fs113_xor1 & f_arrdiv24_mux2to1109_not0;
  assign f_arrdiv24_mux2to1109_xor0 = f_arrdiv24_mux2to1109_and0 ^ f_arrdiv24_mux2to1109_and1;
  assign f_arrdiv24_mux2to1110_and0 = f_arrdiv24_mux2to186_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1110_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1110_and1 = f_arrdiv24_fs114_xor1 & f_arrdiv24_mux2to1110_not0;
  assign f_arrdiv24_mux2to1110_xor0 = f_arrdiv24_mux2to1110_and0 ^ f_arrdiv24_mux2to1110_and1;
  assign f_arrdiv24_mux2to1111_and0 = f_arrdiv24_mux2to187_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1111_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1111_and1 = f_arrdiv24_fs115_xor1 & f_arrdiv24_mux2to1111_not0;
  assign f_arrdiv24_mux2to1111_xor0 = f_arrdiv24_mux2to1111_and0 ^ f_arrdiv24_mux2to1111_and1;
  assign f_arrdiv24_mux2to1112_and0 = f_arrdiv24_mux2to188_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1112_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1112_and1 = f_arrdiv24_fs116_xor1 & f_arrdiv24_mux2to1112_not0;
  assign f_arrdiv24_mux2to1112_xor0 = f_arrdiv24_mux2to1112_and0 ^ f_arrdiv24_mux2to1112_and1;
  assign f_arrdiv24_mux2to1113_and0 = f_arrdiv24_mux2to189_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1113_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1113_and1 = f_arrdiv24_fs117_xor1 & f_arrdiv24_mux2to1113_not0;
  assign f_arrdiv24_mux2to1113_xor0 = f_arrdiv24_mux2to1113_and0 ^ f_arrdiv24_mux2to1113_and1;
  assign f_arrdiv24_mux2to1114_and0 = f_arrdiv24_mux2to190_xor0 & f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1114_not0 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_mux2to1114_and1 = f_arrdiv24_fs118_xor1 & f_arrdiv24_mux2to1114_not0;
  assign f_arrdiv24_mux2to1114_xor0 = f_arrdiv24_mux2to1114_and0 ^ f_arrdiv24_mux2to1114_and1;
  assign f_arrdiv24_not4 = ~f_arrdiv24_fs119_or0;
  assign f_arrdiv24_fs120_xor0 = a[18] ^ b[0];
  assign f_arrdiv24_fs120_not0 = ~a[18];
  assign f_arrdiv24_fs120_and0 = f_arrdiv24_fs120_not0 & b[0];
  assign f_arrdiv24_fs120_not1 = ~f_arrdiv24_fs120_xor0;
  assign f_arrdiv24_fs121_xor0 = f_arrdiv24_mux2to192_xor0 ^ b[1];
  assign f_arrdiv24_fs121_not0 = ~f_arrdiv24_mux2to192_xor0;
  assign f_arrdiv24_fs121_and0 = f_arrdiv24_fs121_not0 & b[1];
  assign f_arrdiv24_fs121_xor1 = f_arrdiv24_fs120_and0 ^ f_arrdiv24_fs121_xor0;
  assign f_arrdiv24_fs121_not1 = ~f_arrdiv24_fs121_xor0;
  assign f_arrdiv24_fs121_and1 = f_arrdiv24_fs121_not1 & f_arrdiv24_fs120_and0;
  assign f_arrdiv24_fs121_or0 = f_arrdiv24_fs121_and1 | f_arrdiv24_fs121_and0;
  assign f_arrdiv24_fs122_xor0 = f_arrdiv24_mux2to193_xor0 ^ b[2];
  assign f_arrdiv24_fs122_not0 = ~f_arrdiv24_mux2to193_xor0;
  assign f_arrdiv24_fs122_and0 = f_arrdiv24_fs122_not0 & b[2];
  assign f_arrdiv24_fs122_xor1 = f_arrdiv24_fs121_or0 ^ f_arrdiv24_fs122_xor0;
  assign f_arrdiv24_fs122_not1 = ~f_arrdiv24_fs122_xor0;
  assign f_arrdiv24_fs122_and1 = f_arrdiv24_fs122_not1 & f_arrdiv24_fs121_or0;
  assign f_arrdiv24_fs122_or0 = f_arrdiv24_fs122_and1 | f_arrdiv24_fs122_and0;
  assign f_arrdiv24_fs123_xor0 = f_arrdiv24_mux2to194_xor0 ^ b[3];
  assign f_arrdiv24_fs123_not0 = ~f_arrdiv24_mux2to194_xor0;
  assign f_arrdiv24_fs123_and0 = f_arrdiv24_fs123_not0 & b[3];
  assign f_arrdiv24_fs123_xor1 = f_arrdiv24_fs122_or0 ^ f_arrdiv24_fs123_xor0;
  assign f_arrdiv24_fs123_not1 = ~f_arrdiv24_fs123_xor0;
  assign f_arrdiv24_fs123_and1 = f_arrdiv24_fs123_not1 & f_arrdiv24_fs122_or0;
  assign f_arrdiv24_fs123_or0 = f_arrdiv24_fs123_and1 | f_arrdiv24_fs123_and0;
  assign f_arrdiv24_fs124_xor0 = f_arrdiv24_mux2to195_xor0 ^ b[4];
  assign f_arrdiv24_fs124_not0 = ~f_arrdiv24_mux2to195_xor0;
  assign f_arrdiv24_fs124_and0 = f_arrdiv24_fs124_not0 & b[4];
  assign f_arrdiv24_fs124_xor1 = f_arrdiv24_fs123_or0 ^ f_arrdiv24_fs124_xor0;
  assign f_arrdiv24_fs124_not1 = ~f_arrdiv24_fs124_xor0;
  assign f_arrdiv24_fs124_and1 = f_arrdiv24_fs124_not1 & f_arrdiv24_fs123_or0;
  assign f_arrdiv24_fs124_or0 = f_arrdiv24_fs124_and1 | f_arrdiv24_fs124_and0;
  assign f_arrdiv24_fs125_xor0 = f_arrdiv24_mux2to196_xor0 ^ b[5];
  assign f_arrdiv24_fs125_not0 = ~f_arrdiv24_mux2to196_xor0;
  assign f_arrdiv24_fs125_and0 = f_arrdiv24_fs125_not0 & b[5];
  assign f_arrdiv24_fs125_xor1 = f_arrdiv24_fs124_or0 ^ f_arrdiv24_fs125_xor0;
  assign f_arrdiv24_fs125_not1 = ~f_arrdiv24_fs125_xor0;
  assign f_arrdiv24_fs125_and1 = f_arrdiv24_fs125_not1 & f_arrdiv24_fs124_or0;
  assign f_arrdiv24_fs125_or0 = f_arrdiv24_fs125_and1 | f_arrdiv24_fs125_and0;
  assign f_arrdiv24_fs126_xor0 = f_arrdiv24_mux2to197_xor0 ^ b[6];
  assign f_arrdiv24_fs126_not0 = ~f_arrdiv24_mux2to197_xor0;
  assign f_arrdiv24_fs126_and0 = f_arrdiv24_fs126_not0 & b[6];
  assign f_arrdiv24_fs126_xor1 = f_arrdiv24_fs125_or0 ^ f_arrdiv24_fs126_xor0;
  assign f_arrdiv24_fs126_not1 = ~f_arrdiv24_fs126_xor0;
  assign f_arrdiv24_fs126_and1 = f_arrdiv24_fs126_not1 & f_arrdiv24_fs125_or0;
  assign f_arrdiv24_fs126_or0 = f_arrdiv24_fs126_and1 | f_arrdiv24_fs126_and0;
  assign f_arrdiv24_fs127_xor0 = f_arrdiv24_mux2to198_xor0 ^ b[7];
  assign f_arrdiv24_fs127_not0 = ~f_arrdiv24_mux2to198_xor0;
  assign f_arrdiv24_fs127_and0 = f_arrdiv24_fs127_not0 & b[7];
  assign f_arrdiv24_fs127_xor1 = f_arrdiv24_fs126_or0 ^ f_arrdiv24_fs127_xor0;
  assign f_arrdiv24_fs127_not1 = ~f_arrdiv24_fs127_xor0;
  assign f_arrdiv24_fs127_and1 = f_arrdiv24_fs127_not1 & f_arrdiv24_fs126_or0;
  assign f_arrdiv24_fs127_or0 = f_arrdiv24_fs127_and1 | f_arrdiv24_fs127_and0;
  assign f_arrdiv24_fs128_xor0 = f_arrdiv24_mux2to199_xor0 ^ b[8];
  assign f_arrdiv24_fs128_not0 = ~f_arrdiv24_mux2to199_xor0;
  assign f_arrdiv24_fs128_and0 = f_arrdiv24_fs128_not0 & b[8];
  assign f_arrdiv24_fs128_xor1 = f_arrdiv24_fs127_or0 ^ f_arrdiv24_fs128_xor0;
  assign f_arrdiv24_fs128_not1 = ~f_arrdiv24_fs128_xor0;
  assign f_arrdiv24_fs128_and1 = f_arrdiv24_fs128_not1 & f_arrdiv24_fs127_or0;
  assign f_arrdiv24_fs128_or0 = f_arrdiv24_fs128_and1 | f_arrdiv24_fs128_and0;
  assign f_arrdiv24_fs129_xor0 = f_arrdiv24_mux2to1100_xor0 ^ b[9];
  assign f_arrdiv24_fs129_not0 = ~f_arrdiv24_mux2to1100_xor0;
  assign f_arrdiv24_fs129_and0 = f_arrdiv24_fs129_not0 & b[9];
  assign f_arrdiv24_fs129_xor1 = f_arrdiv24_fs128_or0 ^ f_arrdiv24_fs129_xor0;
  assign f_arrdiv24_fs129_not1 = ~f_arrdiv24_fs129_xor0;
  assign f_arrdiv24_fs129_and1 = f_arrdiv24_fs129_not1 & f_arrdiv24_fs128_or0;
  assign f_arrdiv24_fs129_or0 = f_arrdiv24_fs129_and1 | f_arrdiv24_fs129_and0;
  assign f_arrdiv24_fs130_xor0 = f_arrdiv24_mux2to1101_xor0 ^ b[10];
  assign f_arrdiv24_fs130_not0 = ~f_arrdiv24_mux2to1101_xor0;
  assign f_arrdiv24_fs130_and0 = f_arrdiv24_fs130_not0 & b[10];
  assign f_arrdiv24_fs130_xor1 = f_arrdiv24_fs129_or0 ^ f_arrdiv24_fs130_xor0;
  assign f_arrdiv24_fs130_not1 = ~f_arrdiv24_fs130_xor0;
  assign f_arrdiv24_fs130_and1 = f_arrdiv24_fs130_not1 & f_arrdiv24_fs129_or0;
  assign f_arrdiv24_fs130_or0 = f_arrdiv24_fs130_and1 | f_arrdiv24_fs130_and0;
  assign f_arrdiv24_fs131_xor0 = f_arrdiv24_mux2to1102_xor0 ^ b[11];
  assign f_arrdiv24_fs131_not0 = ~f_arrdiv24_mux2to1102_xor0;
  assign f_arrdiv24_fs131_and0 = f_arrdiv24_fs131_not0 & b[11];
  assign f_arrdiv24_fs131_xor1 = f_arrdiv24_fs130_or0 ^ f_arrdiv24_fs131_xor0;
  assign f_arrdiv24_fs131_not1 = ~f_arrdiv24_fs131_xor0;
  assign f_arrdiv24_fs131_and1 = f_arrdiv24_fs131_not1 & f_arrdiv24_fs130_or0;
  assign f_arrdiv24_fs131_or0 = f_arrdiv24_fs131_and1 | f_arrdiv24_fs131_and0;
  assign f_arrdiv24_fs132_xor0 = f_arrdiv24_mux2to1103_xor0 ^ b[12];
  assign f_arrdiv24_fs132_not0 = ~f_arrdiv24_mux2to1103_xor0;
  assign f_arrdiv24_fs132_and0 = f_arrdiv24_fs132_not0 & b[12];
  assign f_arrdiv24_fs132_xor1 = f_arrdiv24_fs131_or0 ^ f_arrdiv24_fs132_xor0;
  assign f_arrdiv24_fs132_not1 = ~f_arrdiv24_fs132_xor0;
  assign f_arrdiv24_fs132_and1 = f_arrdiv24_fs132_not1 & f_arrdiv24_fs131_or0;
  assign f_arrdiv24_fs132_or0 = f_arrdiv24_fs132_and1 | f_arrdiv24_fs132_and0;
  assign f_arrdiv24_fs133_xor0 = f_arrdiv24_mux2to1104_xor0 ^ b[13];
  assign f_arrdiv24_fs133_not0 = ~f_arrdiv24_mux2to1104_xor0;
  assign f_arrdiv24_fs133_and0 = f_arrdiv24_fs133_not0 & b[13];
  assign f_arrdiv24_fs133_xor1 = f_arrdiv24_fs132_or0 ^ f_arrdiv24_fs133_xor0;
  assign f_arrdiv24_fs133_not1 = ~f_arrdiv24_fs133_xor0;
  assign f_arrdiv24_fs133_and1 = f_arrdiv24_fs133_not1 & f_arrdiv24_fs132_or0;
  assign f_arrdiv24_fs133_or0 = f_arrdiv24_fs133_and1 | f_arrdiv24_fs133_and0;
  assign f_arrdiv24_fs134_xor0 = f_arrdiv24_mux2to1105_xor0 ^ b[14];
  assign f_arrdiv24_fs134_not0 = ~f_arrdiv24_mux2to1105_xor0;
  assign f_arrdiv24_fs134_and0 = f_arrdiv24_fs134_not0 & b[14];
  assign f_arrdiv24_fs134_xor1 = f_arrdiv24_fs133_or0 ^ f_arrdiv24_fs134_xor0;
  assign f_arrdiv24_fs134_not1 = ~f_arrdiv24_fs134_xor0;
  assign f_arrdiv24_fs134_and1 = f_arrdiv24_fs134_not1 & f_arrdiv24_fs133_or0;
  assign f_arrdiv24_fs134_or0 = f_arrdiv24_fs134_and1 | f_arrdiv24_fs134_and0;
  assign f_arrdiv24_fs135_xor0 = f_arrdiv24_mux2to1106_xor0 ^ b[15];
  assign f_arrdiv24_fs135_not0 = ~f_arrdiv24_mux2to1106_xor0;
  assign f_arrdiv24_fs135_and0 = f_arrdiv24_fs135_not0 & b[15];
  assign f_arrdiv24_fs135_xor1 = f_arrdiv24_fs134_or0 ^ f_arrdiv24_fs135_xor0;
  assign f_arrdiv24_fs135_not1 = ~f_arrdiv24_fs135_xor0;
  assign f_arrdiv24_fs135_and1 = f_arrdiv24_fs135_not1 & f_arrdiv24_fs134_or0;
  assign f_arrdiv24_fs135_or0 = f_arrdiv24_fs135_and1 | f_arrdiv24_fs135_and0;
  assign f_arrdiv24_fs136_xor0 = f_arrdiv24_mux2to1107_xor0 ^ b[16];
  assign f_arrdiv24_fs136_not0 = ~f_arrdiv24_mux2to1107_xor0;
  assign f_arrdiv24_fs136_and0 = f_arrdiv24_fs136_not0 & b[16];
  assign f_arrdiv24_fs136_xor1 = f_arrdiv24_fs135_or0 ^ f_arrdiv24_fs136_xor0;
  assign f_arrdiv24_fs136_not1 = ~f_arrdiv24_fs136_xor0;
  assign f_arrdiv24_fs136_and1 = f_arrdiv24_fs136_not1 & f_arrdiv24_fs135_or0;
  assign f_arrdiv24_fs136_or0 = f_arrdiv24_fs136_and1 | f_arrdiv24_fs136_and0;
  assign f_arrdiv24_fs137_xor0 = f_arrdiv24_mux2to1108_xor0 ^ b[17];
  assign f_arrdiv24_fs137_not0 = ~f_arrdiv24_mux2to1108_xor0;
  assign f_arrdiv24_fs137_and0 = f_arrdiv24_fs137_not0 & b[17];
  assign f_arrdiv24_fs137_xor1 = f_arrdiv24_fs136_or0 ^ f_arrdiv24_fs137_xor0;
  assign f_arrdiv24_fs137_not1 = ~f_arrdiv24_fs137_xor0;
  assign f_arrdiv24_fs137_and1 = f_arrdiv24_fs137_not1 & f_arrdiv24_fs136_or0;
  assign f_arrdiv24_fs137_or0 = f_arrdiv24_fs137_and1 | f_arrdiv24_fs137_and0;
  assign f_arrdiv24_fs138_xor0 = f_arrdiv24_mux2to1109_xor0 ^ b[18];
  assign f_arrdiv24_fs138_not0 = ~f_arrdiv24_mux2to1109_xor0;
  assign f_arrdiv24_fs138_and0 = f_arrdiv24_fs138_not0 & b[18];
  assign f_arrdiv24_fs138_xor1 = f_arrdiv24_fs137_or0 ^ f_arrdiv24_fs138_xor0;
  assign f_arrdiv24_fs138_not1 = ~f_arrdiv24_fs138_xor0;
  assign f_arrdiv24_fs138_and1 = f_arrdiv24_fs138_not1 & f_arrdiv24_fs137_or0;
  assign f_arrdiv24_fs138_or0 = f_arrdiv24_fs138_and1 | f_arrdiv24_fs138_and0;
  assign f_arrdiv24_fs139_xor0 = f_arrdiv24_mux2to1110_xor0 ^ b[19];
  assign f_arrdiv24_fs139_not0 = ~f_arrdiv24_mux2to1110_xor0;
  assign f_arrdiv24_fs139_and0 = f_arrdiv24_fs139_not0 & b[19];
  assign f_arrdiv24_fs139_xor1 = f_arrdiv24_fs138_or0 ^ f_arrdiv24_fs139_xor0;
  assign f_arrdiv24_fs139_not1 = ~f_arrdiv24_fs139_xor0;
  assign f_arrdiv24_fs139_and1 = f_arrdiv24_fs139_not1 & f_arrdiv24_fs138_or0;
  assign f_arrdiv24_fs139_or0 = f_arrdiv24_fs139_and1 | f_arrdiv24_fs139_and0;
  assign f_arrdiv24_fs140_xor0 = f_arrdiv24_mux2to1111_xor0 ^ b[20];
  assign f_arrdiv24_fs140_not0 = ~f_arrdiv24_mux2to1111_xor0;
  assign f_arrdiv24_fs140_and0 = f_arrdiv24_fs140_not0 & b[20];
  assign f_arrdiv24_fs140_xor1 = f_arrdiv24_fs139_or0 ^ f_arrdiv24_fs140_xor0;
  assign f_arrdiv24_fs140_not1 = ~f_arrdiv24_fs140_xor0;
  assign f_arrdiv24_fs140_and1 = f_arrdiv24_fs140_not1 & f_arrdiv24_fs139_or0;
  assign f_arrdiv24_fs140_or0 = f_arrdiv24_fs140_and1 | f_arrdiv24_fs140_and0;
  assign f_arrdiv24_fs141_xor0 = f_arrdiv24_mux2to1112_xor0 ^ b[21];
  assign f_arrdiv24_fs141_not0 = ~f_arrdiv24_mux2to1112_xor0;
  assign f_arrdiv24_fs141_and0 = f_arrdiv24_fs141_not0 & b[21];
  assign f_arrdiv24_fs141_xor1 = f_arrdiv24_fs140_or0 ^ f_arrdiv24_fs141_xor0;
  assign f_arrdiv24_fs141_not1 = ~f_arrdiv24_fs141_xor0;
  assign f_arrdiv24_fs141_and1 = f_arrdiv24_fs141_not1 & f_arrdiv24_fs140_or0;
  assign f_arrdiv24_fs141_or0 = f_arrdiv24_fs141_and1 | f_arrdiv24_fs141_and0;
  assign f_arrdiv24_fs142_xor0 = f_arrdiv24_mux2to1113_xor0 ^ b[22];
  assign f_arrdiv24_fs142_not0 = ~f_arrdiv24_mux2to1113_xor0;
  assign f_arrdiv24_fs142_and0 = f_arrdiv24_fs142_not0 & b[22];
  assign f_arrdiv24_fs142_xor1 = f_arrdiv24_fs141_or0 ^ f_arrdiv24_fs142_xor0;
  assign f_arrdiv24_fs142_not1 = ~f_arrdiv24_fs142_xor0;
  assign f_arrdiv24_fs142_and1 = f_arrdiv24_fs142_not1 & f_arrdiv24_fs141_or0;
  assign f_arrdiv24_fs142_or0 = f_arrdiv24_fs142_and1 | f_arrdiv24_fs142_and0;
  assign f_arrdiv24_fs143_xor0 = f_arrdiv24_mux2to1114_xor0 ^ b[23];
  assign f_arrdiv24_fs143_not0 = ~f_arrdiv24_mux2to1114_xor0;
  assign f_arrdiv24_fs143_and0 = f_arrdiv24_fs143_not0 & b[23];
  assign f_arrdiv24_fs143_xor1 = f_arrdiv24_fs142_or0 ^ f_arrdiv24_fs143_xor0;
  assign f_arrdiv24_fs143_not1 = ~f_arrdiv24_fs143_xor0;
  assign f_arrdiv24_fs143_and1 = f_arrdiv24_fs143_not1 & f_arrdiv24_fs142_or0;
  assign f_arrdiv24_fs143_or0 = f_arrdiv24_fs143_and1 | f_arrdiv24_fs143_and0;
  assign f_arrdiv24_mux2to1115_and0 = a[18] & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1115_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1115_and1 = f_arrdiv24_fs120_xor0 & f_arrdiv24_mux2to1115_not0;
  assign f_arrdiv24_mux2to1115_xor0 = f_arrdiv24_mux2to1115_and0 ^ f_arrdiv24_mux2to1115_and1;
  assign f_arrdiv24_mux2to1116_and0 = f_arrdiv24_mux2to192_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1116_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1116_and1 = f_arrdiv24_fs121_xor1 & f_arrdiv24_mux2to1116_not0;
  assign f_arrdiv24_mux2to1116_xor0 = f_arrdiv24_mux2to1116_and0 ^ f_arrdiv24_mux2to1116_and1;
  assign f_arrdiv24_mux2to1117_and0 = f_arrdiv24_mux2to193_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1117_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1117_and1 = f_arrdiv24_fs122_xor1 & f_arrdiv24_mux2to1117_not0;
  assign f_arrdiv24_mux2to1117_xor0 = f_arrdiv24_mux2to1117_and0 ^ f_arrdiv24_mux2to1117_and1;
  assign f_arrdiv24_mux2to1118_and0 = f_arrdiv24_mux2to194_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1118_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1118_and1 = f_arrdiv24_fs123_xor1 & f_arrdiv24_mux2to1118_not0;
  assign f_arrdiv24_mux2to1118_xor0 = f_arrdiv24_mux2to1118_and0 ^ f_arrdiv24_mux2to1118_and1;
  assign f_arrdiv24_mux2to1119_and0 = f_arrdiv24_mux2to195_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1119_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1119_and1 = f_arrdiv24_fs124_xor1 & f_arrdiv24_mux2to1119_not0;
  assign f_arrdiv24_mux2to1119_xor0 = f_arrdiv24_mux2to1119_and0 ^ f_arrdiv24_mux2to1119_and1;
  assign f_arrdiv24_mux2to1120_and0 = f_arrdiv24_mux2to196_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1120_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1120_and1 = f_arrdiv24_fs125_xor1 & f_arrdiv24_mux2to1120_not0;
  assign f_arrdiv24_mux2to1120_xor0 = f_arrdiv24_mux2to1120_and0 ^ f_arrdiv24_mux2to1120_and1;
  assign f_arrdiv24_mux2to1121_and0 = f_arrdiv24_mux2to197_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1121_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1121_and1 = f_arrdiv24_fs126_xor1 & f_arrdiv24_mux2to1121_not0;
  assign f_arrdiv24_mux2to1121_xor0 = f_arrdiv24_mux2to1121_and0 ^ f_arrdiv24_mux2to1121_and1;
  assign f_arrdiv24_mux2to1122_and0 = f_arrdiv24_mux2to198_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1122_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1122_and1 = f_arrdiv24_fs127_xor1 & f_arrdiv24_mux2to1122_not0;
  assign f_arrdiv24_mux2to1122_xor0 = f_arrdiv24_mux2to1122_and0 ^ f_arrdiv24_mux2to1122_and1;
  assign f_arrdiv24_mux2to1123_and0 = f_arrdiv24_mux2to199_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1123_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1123_and1 = f_arrdiv24_fs128_xor1 & f_arrdiv24_mux2to1123_not0;
  assign f_arrdiv24_mux2to1123_xor0 = f_arrdiv24_mux2to1123_and0 ^ f_arrdiv24_mux2to1123_and1;
  assign f_arrdiv24_mux2to1124_and0 = f_arrdiv24_mux2to1100_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1124_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1124_and1 = f_arrdiv24_fs129_xor1 & f_arrdiv24_mux2to1124_not0;
  assign f_arrdiv24_mux2to1124_xor0 = f_arrdiv24_mux2to1124_and0 ^ f_arrdiv24_mux2to1124_and1;
  assign f_arrdiv24_mux2to1125_and0 = f_arrdiv24_mux2to1101_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1125_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1125_and1 = f_arrdiv24_fs130_xor1 & f_arrdiv24_mux2to1125_not0;
  assign f_arrdiv24_mux2to1125_xor0 = f_arrdiv24_mux2to1125_and0 ^ f_arrdiv24_mux2to1125_and1;
  assign f_arrdiv24_mux2to1126_and0 = f_arrdiv24_mux2to1102_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1126_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1126_and1 = f_arrdiv24_fs131_xor1 & f_arrdiv24_mux2to1126_not0;
  assign f_arrdiv24_mux2to1126_xor0 = f_arrdiv24_mux2to1126_and0 ^ f_arrdiv24_mux2to1126_and1;
  assign f_arrdiv24_mux2to1127_and0 = f_arrdiv24_mux2to1103_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1127_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1127_and1 = f_arrdiv24_fs132_xor1 & f_arrdiv24_mux2to1127_not0;
  assign f_arrdiv24_mux2to1127_xor0 = f_arrdiv24_mux2to1127_and0 ^ f_arrdiv24_mux2to1127_and1;
  assign f_arrdiv24_mux2to1128_and0 = f_arrdiv24_mux2to1104_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1128_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1128_and1 = f_arrdiv24_fs133_xor1 & f_arrdiv24_mux2to1128_not0;
  assign f_arrdiv24_mux2to1128_xor0 = f_arrdiv24_mux2to1128_and0 ^ f_arrdiv24_mux2to1128_and1;
  assign f_arrdiv24_mux2to1129_and0 = f_arrdiv24_mux2to1105_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1129_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1129_and1 = f_arrdiv24_fs134_xor1 & f_arrdiv24_mux2to1129_not0;
  assign f_arrdiv24_mux2to1129_xor0 = f_arrdiv24_mux2to1129_and0 ^ f_arrdiv24_mux2to1129_and1;
  assign f_arrdiv24_mux2to1130_and0 = f_arrdiv24_mux2to1106_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1130_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1130_and1 = f_arrdiv24_fs135_xor1 & f_arrdiv24_mux2to1130_not0;
  assign f_arrdiv24_mux2to1130_xor0 = f_arrdiv24_mux2to1130_and0 ^ f_arrdiv24_mux2to1130_and1;
  assign f_arrdiv24_mux2to1131_and0 = f_arrdiv24_mux2to1107_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1131_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1131_and1 = f_arrdiv24_fs136_xor1 & f_arrdiv24_mux2to1131_not0;
  assign f_arrdiv24_mux2to1131_xor0 = f_arrdiv24_mux2to1131_and0 ^ f_arrdiv24_mux2to1131_and1;
  assign f_arrdiv24_mux2to1132_and0 = f_arrdiv24_mux2to1108_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1132_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1132_and1 = f_arrdiv24_fs137_xor1 & f_arrdiv24_mux2to1132_not0;
  assign f_arrdiv24_mux2to1132_xor0 = f_arrdiv24_mux2to1132_and0 ^ f_arrdiv24_mux2to1132_and1;
  assign f_arrdiv24_mux2to1133_and0 = f_arrdiv24_mux2to1109_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1133_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1133_and1 = f_arrdiv24_fs138_xor1 & f_arrdiv24_mux2to1133_not0;
  assign f_arrdiv24_mux2to1133_xor0 = f_arrdiv24_mux2to1133_and0 ^ f_arrdiv24_mux2to1133_and1;
  assign f_arrdiv24_mux2to1134_and0 = f_arrdiv24_mux2to1110_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1134_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1134_and1 = f_arrdiv24_fs139_xor1 & f_arrdiv24_mux2to1134_not0;
  assign f_arrdiv24_mux2to1134_xor0 = f_arrdiv24_mux2to1134_and0 ^ f_arrdiv24_mux2to1134_and1;
  assign f_arrdiv24_mux2to1135_and0 = f_arrdiv24_mux2to1111_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1135_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1135_and1 = f_arrdiv24_fs140_xor1 & f_arrdiv24_mux2to1135_not0;
  assign f_arrdiv24_mux2to1135_xor0 = f_arrdiv24_mux2to1135_and0 ^ f_arrdiv24_mux2to1135_and1;
  assign f_arrdiv24_mux2to1136_and0 = f_arrdiv24_mux2to1112_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1136_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1136_and1 = f_arrdiv24_fs141_xor1 & f_arrdiv24_mux2to1136_not0;
  assign f_arrdiv24_mux2to1136_xor0 = f_arrdiv24_mux2to1136_and0 ^ f_arrdiv24_mux2to1136_and1;
  assign f_arrdiv24_mux2to1137_and0 = f_arrdiv24_mux2to1113_xor0 & f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1137_not0 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_mux2to1137_and1 = f_arrdiv24_fs142_xor1 & f_arrdiv24_mux2to1137_not0;
  assign f_arrdiv24_mux2to1137_xor0 = f_arrdiv24_mux2to1137_and0 ^ f_arrdiv24_mux2to1137_and1;
  assign f_arrdiv24_not5 = ~f_arrdiv24_fs143_or0;
  assign f_arrdiv24_fs144_xor0 = a[17] ^ b[0];
  assign f_arrdiv24_fs144_not0 = ~a[17];
  assign f_arrdiv24_fs144_and0 = f_arrdiv24_fs144_not0 & b[0];
  assign f_arrdiv24_fs144_not1 = ~f_arrdiv24_fs144_xor0;
  assign f_arrdiv24_fs145_xor0 = f_arrdiv24_mux2to1115_xor0 ^ b[1];
  assign f_arrdiv24_fs145_not0 = ~f_arrdiv24_mux2to1115_xor0;
  assign f_arrdiv24_fs145_and0 = f_arrdiv24_fs145_not0 & b[1];
  assign f_arrdiv24_fs145_xor1 = f_arrdiv24_fs144_and0 ^ f_arrdiv24_fs145_xor0;
  assign f_arrdiv24_fs145_not1 = ~f_arrdiv24_fs145_xor0;
  assign f_arrdiv24_fs145_and1 = f_arrdiv24_fs145_not1 & f_arrdiv24_fs144_and0;
  assign f_arrdiv24_fs145_or0 = f_arrdiv24_fs145_and1 | f_arrdiv24_fs145_and0;
  assign f_arrdiv24_fs146_xor0 = f_arrdiv24_mux2to1116_xor0 ^ b[2];
  assign f_arrdiv24_fs146_not0 = ~f_arrdiv24_mux2to1116_xor0;
  assign f_arrdiv24_fs146_and0 = f_arrdiv24_fs146_not0 & b[2];
  assign f_arrdiv24_fs146_xor1 = f_arrdiv24_fs145_or0 ^ f_arrdiv24_fs146_xor0;
  assign f_arrdiv24_fs146_not1 = ~f_arrdiv24_fs146_xor0;
  assign f_arrdiv24_fs146_and1 = f_arrdiv24_fs146_not1 & f_arrdiv24_fs145_or0;
  assign f_arrdiv24_fs146_or0 = f_arrdiv24_fs146_and1 | f_arrdiv24_fs146_and0;
  assign f_arrdiv24_fs147_xor0 = f_arrdiv24_mux2to1117_xor0 ^ b[3];
  assign f_arrdiv24_fs147_not0 = ~f_arrdiv24_mux2to1117_xor0;
  assign f_arrdiv24_fs147_and0 = f_arrdiv24_fs147_not0 & b[3];
  assign f_arrdiv24_fs147_xor1 = f_arrdiv24_fs146_or0 ^ f_arrdiv24_fs147_xor0;
  assign f_arrdiv24_fs147_not1 = ~f_arrdiv24_fs147_xor0;
  assign f_arrdiv24_fs147_and1 = f_arrdiv24_fs147_not1 & f_arrdiv24_fs146_or0;
  assign f_arrdiv24_fs147_or0 = f_arrdiv24_fs147_and1 | f_arrdiv24_fs147_and0;
  assign f_arrdiv24_fs148_xor0 = f_arrdiv24_mux2to1118_xor0 ^ b[4];
  assign f_arrdiv24_fs148_not0 = ~f_arrdiv24_mux2to1118_xor0;
  assign f_arrdiv24_fs148_and0 = f_arrdiv24_fs148_not0 & b[4];
  assign f_arrdiv24_fs148_xor1 = f_arrdiv24_fs147_or0 ^ f_arrdiv24_fs148_xor0;
  assign f_arrdiv24_fs148_not1 = ~f_arrdiv24_fs148_xor0;
  assign f_arrdiv24_fs148_and1 = f_arrdiv24_fs148_not1 & f_arrdiv24_fs147_or0;
  assign f_arrdiv24_fs148_or0 = f_arrdiv24_fs148_and1 | f_arrdiv24_fs148_and0;
  assign f_arrdiv24_fs149_xor0 = f_arrdiv24_mux2to1119_xor0 ^ b[5];
  assign f_arrdiv24_fs149_not0 = ~f_arrdiv24_mux2to1119_xor0;
  assign f_arrdiv24_fs149_and0 = f_arrdiv24_fs149_not0 & b[5];
  assign f_arrdiv24_fs149_xor1 = f_arrdiv24_fs148_or0 ^ f_arrdiv24_fs149_xor0;
  assign f_arrdiv24_fs149_not1 = ~f_arrdiv24_fs149_xor0;
  assign f_arrdiv24_fs149_and1 = f_arrdiv24_fs149_not1 & f_arrdiv24_fs148_or0;
  assign f_arrdiv24_fs149_or0 = f_arrdiv24_fs149_and1 | f_arrdiv24_fs149_and0;
  assign f_arrdiv24_fs150_xor0 = f_arrdiv24_mux2to1120_xor0 ^ b[6];
  assign f_arrdiv24_fs150_not0 = ~f_arrdiv24_mux2to1120_xor0;
  assign f_arrdiv24_fs150_and0 = f_arrdiv24_fs150_not0 & b[6];
  assign f_arrdiv24_fs150_xor1 = f_arrdiv24_fs149_or0 ^ f_arrdiv24_fs150_xor0;
  assign f_arrdiv24_fs150_not1 = ~f_arrdiv24_fs150_xor0;
  assign f_arrdiv24_fs150_and1 = f_arrdiv24_fs150_not1 & f_arrdiv24_fs149_or0;
  assign f_arrdiv24_fs150_or0 = f_arrdiv24_fs150_and1 | f_arrdiv24_fs150_and0;
  assign f_arrdiv24_fs151_xor0 = f_arrdiv24_mux2to1121_xor0 ^ b[7];
  assign f_arrdiv24_fs151_not0 = ~f_arrdiv24_mux2to1121_xor0;
  assign f_arrdiv24_fs151_and0 = f_arrdiv24_fs151_not0 & b[7];
  assign f_arrdiv24_fs151_xor1 = f_arrdiv24_fs150_or0 ^ f_arrdiv24_fs151_xor0;
  assign f_arrdiv24_fs151_not1 = ~f_arrdiv24_fs151_xor0;
  assign f_arrdiv24_fs151_and1 = f_arrdiv24_fs151_not1 & f_arrdiv24_fs150_or0;
  assign f_arrdiv24_fs151_or0 = f_arrdiv24_fs151_and1 | f_arrdiv24_fs151_and0;
  assign f_arrdiv24_fs152_xor0 = f_arrdiv24_mux2to1122_xor0 ^ b[8];
  assign f_arrdiv24_fs152_not0 = ~f_arrdiv24_mux2to1122_xor0;
  assign f_arrdiv24_fs152_and0 = f_arrdiv24_fs152_not0 & b[8];
  assign f_arrdiv24_fs152_xor1 = f_arrdiv24_fs151_or0 ^ f_arrdiv24_fs152_xor0;
  assign f_arrdiv24_fs152_not1 = ~f_arrdiv24_fs152_xor0;
  assign f_arrdiv24_fs152_and1 = f_arrdiv24_fs152_not1 & f_arrdiv24_fs151_or0;
  assign f_arrdiv24_fs152_or0 = f_arrdiv24_fs152_and1 | f_arrdiv24_fs152_and0;
  assign f_arrdiv24_fs153_xor0 = f_arrdiv24_mux2to1123_xor0 ^ b[9];
  assign f_arrdiv24_fs153_not0 = ~f_arrdiv24_mux2to1123_xor0;
  assign f_arrdiv24_fs153_and0 = f_arrdiv24_fs153_not0 & b[9];
  assign f_arrdiv24_fs153_xor1 = f_arrdiv24_fs152_or0 ^ f_arrdiv24_fs153_xor0;
  assign f_arrdiv24_fs153_not1 = ~f_arrdiv24_fs153_xor0;
  assign f_arrdiv24_fs153_and1 = f_arrdiv24_fs153_not1 & f_arrdiv24_fs152_or0;
  assign f_arrdiv24_fs153_or0 = f_arrdiv24_fs153_and1 | f_arrdiv24_fs153_and0;
  assign f_arrdiv24_fs154_xor0 = f_arrdiv24_mux2to1124_xor0 ^ b[10];
  assign f_arrdiv24_fs154_not0 = ~f_arrdiv24_mux2to1124_xor0;
  assign f_arrdiv24_fs154_and0 = f_arrdiv24_fs154_not0 & b[10];
  assign f_arrdiv24_fs154_xor1 = f_arrdiv24_fs153_or0 ^ f_arrdiv24_fs154_xor0;
  assign f_arrdiv24_fs154_not1 = ~f_arrdiv24_fs154_xor0;
  assign f_arrdiv24_fs154_and1 = f_arrdiv24_fs154_not1 & f_arrdiv24_fs153_or0;
  assign f_arrdiv24_fs154_or0 = f_arrdiv24_fs154_and1 | f_arrdiv24_fs154_and0;
  assign f_arrdiv24_fs155_xor0 = f_arrdiv24_mux2to1125_xor0 ^ b[11];
  assign f_arrdiv24_fs155_not0 = ~f_arrdiv24_mux2to1125_xor0;
  assign f_arrdiv24_fs155_and0 = f_arrdiv24_fs155_not0 & b[11];
  assign f_arrdiv24_fs155_xor1 = f_arrdiv24_fs154_or0 ^ f_arrdiv24_fs155_xor0;
  assign f_arrdiv24_fs155_not1 = ~f_arrdiv24_fs155_xor0;
  assign f_arrdiv24_fs155_and1 = f_arrdiv24_fs155_not1 & f_arrdiv24_fs154_or0;
  assign f_arrdiv24_fs155_or0 = f_arrdiv24_fs155_and1 | f_arrdiv24_fs155_and0;
  assign f_arrdiv24_fs156_xor0 = f_arrdiv24_mux2to1126_xor0 ^ b[12];
  assign f_arrdiv24_fs156_not0 = ~f_arrdiv24_mux2to1126_xor0;
  assign f_arrdiv24_fs156_and0 = f_arrdiv24_fs156_not0 & b[12];
  assign f_arrdiv24_fs156_xor1 = f_arrdiv24_fs155_or0 ^ f_arrdiv24_fs156_xor0;
  assign f_arrdiv24_fs156_not1 = ~f_arrdiv24_fs156_xor0;
  assign f_arrdiv24_fs156_and1 = f_arrdiv24_fs156_not1 & f_arrdiv24_fs155_or0;
  assign f_arrdiv24_fs156_or0 = f_arrdiv24_fs156_and1 | f_arrdiv24_fs156_and0;
  assign f_arrdiv24_fs157_xor0 = f_arrdiv24_mux2to1127_xor0 ^ b[13];
  assign f_arrdiv24_fs157_not0 = ~f_arrdiv24_mux2to1127_xor0;
  assign f_arrdiv24_fs157_and0 = f_arrdiv24_fs157_not0 & b[13];
  assign f_arrdiv24_fs157_xor1 = f_arrdiv24_fs156_or0 ^ f_arrdiv24_fs157_xor0;
  assign f_arrdiv24_fs157_not1 = ~f_arrdiv24_fs157_xor0;
  assign f_arrdiv24_fs157_and1 = f_arrdiv24_fs157_not1 & f_arrdiv24_fs156_or0;
  assign f_arrdiv24_fs157_or0 = f_arrdiv24_fs157_and1 | f_arrdiv24_fs157_and0;
  assign f_arrdiv24_fs158_xor0 = f_arrdiv24_mux2to1128_xor0 ^ b[14];
  assign f_arrdiv24_fs158_not0 = ~f_arrdiv24_mux2to1128_xor0;
  assign f_arrdiv24_fs158_and0 = f_arrdiv24_fs158_not0 & b[14];
  assign f_arrdiv24_fs158_xor1 = f_arrdiv24_fs157_or0 ^ f_arrdiv24_fs158_xor0;
  assign f_arrdiv24_fs158_not1 = ~f_arrdiv24_fs158_xor0;
  assign f_arrdiv24_fs158_and1 = f_arrdiv24_fs158_not1 & f_arrdiv24_fs157_or0;
  assign f_arrdiv24_fs158_or0 = f_arrdiv24_fs158_and1 | f_arrdiv24_fs158_and0;
  assign f_arrdiv24_fs159_xor0 = f_arrdiv24_mux2to1129_xor0 ^ b[15];
  assign f_arrdiv24_fs159_not0 = ~f_arrdiv24_mux2to1129_xor0;
  assign f_arrdiv24_fs159_and0 = f_arrdiv24_fs159_not0 & b[15];
  assign f_arrdiv24_fs159_xor1 = f_arrdiv24_fs158_or0 ^ f_arrdiv24_fs159_xor0;
  assign f_arrdiv24_fs159_not1 = ~f_arrdiv24_fs159_xor0;
  assign f_arrdiv24_fs159_and1 = f_arrdiv24_fs159_not1 & f_arrdiv24_fs158_or0;
  assign f_arrdiv24_fs159_or0 = f_arrdiv24_fs159_and1 | f_arrdiv24_fs159_and0;
  assign f_arrdiv24_fs160_xor0 = f_arrdiv24_mux2to1130_xor0 ^ b[16];
  assign f_arrdiv24_fs160_not0 = ~f_arrdiv24_mux2to1130_xor0;
  assign f_arrdiv24_fs160_and0 = f_arrdiv24_fs160_not0 & b[16];
  assign f_arrdiv24_fs160_xor1 = f_arrdiv24_fs159_or0 ^ f_arrdiv24_fs160_xor0;
  assign f_arrdiv24_fs160_not1 = ~f_arrdiv24_fs160_xor0;
  assign f_arrdiv24_fs160_and1 = f_arrdiv24_fs160_not1 & f_arrdiv24_fs159_or0;
  assign f_arrdiv24_fs160_or0 = f_arrdiv24_fs160_and1 | f_arrdiv24_fs160_and0;
  assign f_arrdiv24_fs161_xor0 = f_arrdiv24_mux2to1131_xor0 ^ b[17];
  assign f_arrdiv24_fs161_not0 = ~f_arrdiv24_mux2to1131_xor0;
  assign f_arrdiv24_fs161_and0 = f_arrdiv24_fs161_not0 & b[17];
  assign f_arrdiv24_fs161_xor1 = f_arrdiv24_fs160_or0 ^ f_arrdiv24_fs161_xor0;
  assign f_arrdiv24_fs161_not1 = ~f_arrdiv24_fs161_xor0;
  assign f_arrdiv24_fs161_and1 = f_arrdiv24_fs161_not1 & f_arrdiv24_fs160_or0;
  assign f_arrdiv24_fs161_or0 = f_arrdiv24_fs161_and1 | f_arrdiv24_fs161_and0;
  assign f_arrdiv24_fs162_xor0 = f_arrdiv24_mux2to1132_xor0 ^ b[18];
  assign f_arrdiv24_fs162_not0 = ~f_arrdiv24_mux2to1132_xor0;
  assign f_arrdiv24_fs162_and0 = f_arrdiv24_fs162_not0 & b[18];
  assign f_arrdiv24_fs162_xor1 = f_arrdiv24_fs161_or0 ^ f_arrdiv24_fs162_xor0;
  assign f_arrdiv24_fs162_not1 = ~f_arrdiv24_fs162_xor0;
  assign f_arrdiv24_fs162_and1 = f_arrdiv24_fs162_not1 & f_arrdiv24_fs161_or0;
  assign f_arrdiv24_fs162_or0 = f_arrdiv24_fs162_and1 | f_arrdiv24_fs162_and0;
  assign f_arrdiv24_fs163_xor0 = f_arrdiv24_mux2to1133_xor0 ^ b[19];
  assign f_arrdiv24_fs163_not0 = ~f_arrdiv24_mux2to1133_xor0;
  assign f_arrdiv24_fs163_and0 = f_arrdiv24_fs163_not0 & b[19];
  assign f_arrdiv24_fs163_xor1 = f_arrdiv24_fs162_or0 ^ f_arrdiv24_fs163_xor0;
  assign f_arrdiv24_fs163_not1 = ~f_arrdiv24_fs163_xor0;
  assign f_arrdiv24_fs163_and1 = f_arrdiv24_fs163_not1 & f_arrdiv24_fs162_or0;
  assign f_arrdiv24_fs163_or0 = f_arrdiv24_fs163_and1 | f_arrdiv24_fs163_and0;
  assign f_arrdiv24_fs164_xor0 = f_arrdiv24_mux2to1134_xor0 ^ b[20];
  assign f_arrdiv24_fs164_not0 = ~f_arrdiv24_mux2to1134_xor0;
  assign f_arrdiv24_fs164_and0 = f_arrdiv24_fs164_not0 & b[20];
  assign f_arrdiv24_fs164_xor1 = f_arrdiv24_fs163_or0 ^ f_arrdiv24_fs164_xor0;
  assign f_arrdiv24_fs164_not1 = ~f_arrdiv24_fs164_xor0;
  assign f_arrdiv24_fs164_and1 = f_arrdiv24_fs164_not1 & f_arrdiv24_fs163_or0;
  assign f_arrdiv24_fs164_or0 = f_arrdiv24_fs164_and1 | f_arrdiv24_fs164_and0;
  assign f_arrdiv24_fs165_xor0 = f_arrdiv24_mux2to1135_xor0 ^ b[21];
  assign f_arrdiv24_fs165_not0 = ~f_arrdiv24_mux2to1135_xor0;
  assign f_arrdiv24_fs165_and0 = f_arrdiv24_fs165_not0 & b[21];
  assign f_arrdiv24_fs165_xor1 = f_arrdiv24_fs164_or0 ^ f_arrdiv24_fs165_xor0;
  assign f_arrdiv24_fs165_not1 = ~f_arrdiv24_fs165_xor0;
  assign f_arrdiv24_fs165_and1 = f_arrdiv24_fs165_not1 & f_arrdiv24_fs164_or0;
  assign f_arrdiv24_fs165_or0 = f_arrdiv24_fs165_and1 | f_arrdiv24_fs165_and0;
  assign f_arrdiv24_fs166_xor0 = f_arrdiv24_mux2to1136_xor0 ^ b[22];
  assign f_arrdiv24_fs166_not0 = ~f_arrdiv24_mux2to1136_xor0;
  assign f_arrdiv24_fs166_and0 = f_arrdiv24_fs166_not0 & b[22];
  assign f_arrdiv24_fs166_xor1 = f_arrdiv24_fs165_or0 ^ f_arrdiv24_fs166_xor0;
  assign f_arrdiv24_fs166_not1 = ~f_arrdiv24_fs166_xor0;
  assign f_arrdiv24_fs166_and1 = f_arrdiv24_fs166_not1 & f_arrdiv24_fs165_or0;
  assign f_arrdiv24_fs166_or0 = f_arrdiv24_fs166_and1 | f_arrdiv24_fs166_and0;
  assign f_arrdiv24_fs167_xor0 = f_arrdiv24_mux2to1137_xor0 ^ b[23];
  assign f_arrdiv24_fs167_not0 = ~f_arrdiv24_mux2to1137_xor0;
  assign f_arrdiv24_fs167_and0 = f_arrdiv24_fs167_not0 & b[23];
  assign f_arrdiv24_fs167_xor1 = f_arrdiv24_fs166_or0 ^ f_arrdiv24_fs167_xor0;
  assign f_arrdiv24_fs167_not1 = ~f_arrdiv24_fs167_xor0;
  assign f_arrdiv24_fs167_and1 = f_arrdiv24_fs167_not1 & f_arrdiv24_fs166_or0;
  assign f_arrdiv24_fs167_or0 = f_arrdiv24_fs167_and1 | f_arrdiv24_fs167_and0;
  assign f_arrdiv24_mux2to1138_and0 = a[17] & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1138_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1138_and1 = f_arrdiv24_fs144_xor0 & f_arrdiv24_mux2to1138_not0;
  assign f_arrdiv24_mux2to1138_xor0 = f_arrdiv24_mux2to1138_and0 ^ f_arrdiv24_mux2to1138_and1;
  assign f_arrdiv24_mux2to1139_and0 = f_arrdiv24_mux2to1115_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1139_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1139_and1 = f_arrdiv24_fs145_xor1 & f_arrdiv24_mux2to1139_not0;
  assign f_arrdiv24_mux2to1139_xor0 = f_arrdiv24_mux2to1139_and0 ^ f_arrdiv24_mux2to1139_and1;
  assign f_arrdiv24_mux2to1140_and0 = f_arrdiv24_mux2to1116_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1140_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1140_and1 = f_arrdiv24_fs146_xor1 & f_arrdiv24_mux2to1140_not0;
  assign f_arrdiv24_mux2to1140_xor0 = f_arrdiv24_mux2to1140_and0 ^ f_arrdiv24_mux2to1140_and1;
  assign f_arrdiv24_mux2to1141_and0 = f_arrdiv24_mux2to1117_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1141_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1141_and1 = f_arrdiv24_fs147_xor1 & f_arrdiv24_mux2to1141_not0;
  assign f_arrdiv24_mux2to1141_xor0 = f_arrdiv24_mux2to1141_and0 ^ f_arrdiv24_mux2to1141_and1;
  assign f_arrdiv24_mux2to1142_and0 = f_arrdiv24_mux2to1118_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1142_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1142_and1 = f_arrdiv24_fs148_xor1 & f_arrdiv24_mux2to1142_not0;
  assign f_arrdiv24_mux2to1142_xor0 = f_arrdiv24_mux2to1142_and0 ^ f_arrdiv24_mux2to1142_and1;
  assign f_arrdiv24_mux2to1143_and0 = f_arrdiv24_mux2to1119_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1143_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1143_and1 = f_arrdiv24_fs149_xor1 & f_arrdiv24_mux2to1143_not0;
  assign f_arrdiv24_mux2to1143_xor0 = f_arrdiv24_mux2to1143_and0 ^ f_arrdiv24_mux2to1143_and1;
  assign f_arrdiv24_mux2to1144_and0 = f_arrdiv24_mux2to1120_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1144_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1144_and1 = f_arrdiv24_fs150_xor1 & f_arrdiv24_mux2to1144_not0;
  assign f_arrdiv24_mux2to1144_xor0 = f_arrdiv24_mux2to1144_and0 ^ f_arrdiv24_mux2to1144_and1;
  assign f_arrdiv24_mux2to1145_and0 = f_arrdiv24_mux2to1121_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1145_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1145_and1 = f_arrdiv24_fs151_xor1 & f_arrdiv24_mux2to1145_not0;
  assign f_arrdiv24_mux2to1145_xor0 = f_arrdiv24_mux2to1145_and0 ^ f_arrdiv24_mux2to1145_and1;
  assign f_arrdiv24_mux2to1146_and0 = f_arrdiv24_mux2to1122_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1146_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1146_and1 = f_arrdiv24_fs152_xor1 & f_arrdiv24_mux2to1146_not0;
  assign f_arrdiv24_mux2to1146_xor0 = f_arrdiv24_mux2to1146_and0 ^ f_arrdiv24_mux2to1146_and1;
  assign f_arrdiv24_mux2to1147_and0 = f_arrdiv24_mux2to1123_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1147_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1147_and1 = f_arrdiv24_fs153_xor1 & f_arrdiv24_mux2to1147_not0;
  assign f_arrdiv24_mux2to1147_xor0 = f_arrdiv24_mux2to1147_and0 ^ f_arrdiv24_mux2to1147_and1;
  assign f_arrdiv24_mux2to1148_and0 = f_arrdiv24_mux2to1124_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1148_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1148_and1 = f_arrdiv24_fs154_xor1 & f_arrdiv24_mux2to1148_not0;
  assign f_arrdiv24_mux2to1148_xor0 = f_arrdiv24_mux2to1148_and0 ^ f_arrdiv24_mux2to1148_and1;
  assign f_arrdiv24_mux2to1149_and0 = f_arrdiv24_mux2to1125_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1149_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1149_and1 = f_arrdiv24_fs155_xor1 & f_arrdiv24_mux2to1149_not0;
  assign f_arrdiv24_mux2to1149_xor0 = f_arrdiv24_mux2to1149_and0 ^ f_arrdiv24_mux2to1149_and1;
  assign f_arrdiv24_mux2to1150_and0 = f_arrdiv24_mux2to1126_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1150_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1150_and1 = f_arrdiv24_fs156_xor1 & f_arrdiv24_mux2to1150_not0;
  assign f_arrdiv24_mux2to1150_xor0 = f_arrdiv24_mux2to1150_and0 ^ f_arrdiv24_mux2to1150_and1;
  assign f_arrdiv24_mux2to1151_and0 = f_arrdiv24_mux2to1127_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1151_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1151_and1 = f_arrdiv24_fs157_xor1 & f_arrdiv24_mux2to1151_not0;
  assign f_arrdiv24_mux2to1151_xor0 = f_arrdiv24_mux2to1151_and0 ^ f_arrdiv24_mux2to1151_and1;
  assign f_arrdiv24_mux2to1152_and0 = f_arrdiv24_mux2to1128_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1152_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1152_and1 = f_arrdiv24_fs158_xor1 & f_arrdiv24_mux2to1152_not0;
  assign f_arrdiv24_mux2to1152_xor0 = f_arrdiv24_mux2to1152_and0 ^ f_arrdiv24_mux2to1152_and1;
  assign f_arrdiv24_mux2to1153_and0 = f_arrdiv24_mux2to1129_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1153_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1153_and1 = f_arrdiv24_fs159_xor1 & f_arrdiv24_mux2to1153_not0;
  assign f_arrdiv24_mux2to1153_xor0 = f_arrdiv24_mux2to1153_and0 ^ f_arrdiv24_mux2to1153_and1;
  assign f_arrdiv24_mux2to1154_and0 = f_arrdiv24_mux2to1130_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1154_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1154_and1 = f_arrdiv24_fs160_xor1 & f_arrdiv24_mux2to1154_not0;
  assign f_arrdiv24_mux2to1154_xor0 = f_arrdiv24_mux2to1154_and0 ^ f_arrdiv24_mux2to1154_and1;
  assign f_arrdiv24_mux2to1155_and0 = f_arrdiv24_mux2to1131_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1155_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1155_and1 = f_arrdiv24_fs161_xor1 & f_arrdiv24_mux2to1155_not0;
  assign f_arrdiv24_mux2to1155_xor0 = f_arrdiv24_mux2to1155_and0 ^ f_arrdiv24_mux2to1155_and1;
  assign f_arrdiv24_mux2to1156_and0 = f_arrdiv24_mux2to1132_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1156_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1156_and1 = f_arrdiv24_fs162_xor1 & f_arrdiv24_mux2to1156_not0;
  assign f_arrdiv24_mux2to1156_xor0 = f_arrdiv24_mux2to1156_and0 ^ f_arrdiv24_mux2to1156_and1;
  assign f_arrdiv24_mux2to1157_and0 = f_arrdiv24_mux2to1133_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1157_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1157_and1 = f_arrdiv24_fs163_xor1 & f_arrdiv24_mux2to1157_not0;
  assign f_arrdiv24_mux2to1157_xor0 = f_arrdiv24_mux2to1157_and0 ^ f_arrdiv24_mux2to1157_and1;
  assign f_arrdiv24_mux2to1158_and0 = f_arrdiv24_mux2to1134_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1158_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1158_and1 = f_arrdiv24_fs164_xor1 & f_arrdiv24_mux2to1158_not0;
  assign f_arrdiv24_mux2to1158_xor0 = f_arrdiv24_mux2to1158_and0 ^ f_arrdiv24_mux2to1158_and1;
  assign f_arrdiv24_mux2to1159_and0 = f_arrdiv24_mux2to1135_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1159_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1159_and1 = f_arrdiv24_fs165_xor1 & f_arrdiv24_mux2to1159_not0;
  assign f_arrdiv24_mux2to1159_xor0 = f_arrdiv24_mux2to1159_and0 ^ f_arrdiv24_mux2to1159_and1;
  assign f_arrdiv24_mux2to1160_and0 = f_arrdiv24_mux2to1136_xor0 & f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1160_not0 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_mux2to1160_and1 = f_arrdiv24_fs166_xor1 & f_arrdiv24_mux2to1160_not0;
  assign f_arrdiv24_mux2to1160_xor0 = f_arrdiv24_mux2to1160_and0 ^ f_arrdiv24_mux2to1160_and1;
  assign f_arrdiv24_not6 = ~f_arrdiv24_fs167_or0;
  assign f_arrdiv24_fs168_xor0 = a[16] ^ b[0];
  assign f_arrdiv24_fs168_not0 = ~a[16];
  assign f_arrdiv24_fs168_and0 = f_arrdiv24_fs168_not0 & b[0];
  assign f_arrdiv24_fs168_not1 = ~f_arrdiv24_fs168_xor0;
  assign f_arrdiv24_fs169_xor0 = f_arrdiv24_mux2to1138_xor0 ^ b[1];
  assign f_arrdiv24_fs169_not0 = ~f_arrdiv24_mux2to1138_xor0;
  assign f_arrdiv24_fs169_and0 = f_arrdiv24_fs169_not0 & b[1];
  assign f_arrdiv24_fs169_xor1 = f_arrdiv24_fs168_and0 ^ f_arrdiv24_fs169_xor0;
  assign f_arrdiv24_fs169_not1 = ~f_arrdiv24_fs169_xor0;
  assign f_arrdiv24_fs169_and1 = f_arrdiv24_fs169_not1 & f_arrdiv24_fs168_and0;
  assign f_arrdiv24_fs169_or0 = f_arrdiv24_fs169_and1 | f_arrdiv24_fs169_and0;
  assign f_arrdiv24_fs170_xor0 = f_arrdiv24_mux2to1139_xor0 ^ b[2];
  assign f_arrdiv24_fs170_not0 = ~f_arrdiv24_mux2to1139_xor0;
  assign f_arrdiv24_fs170_and0 = f_arrdiv24_fs170_not0 & b[2];
  assign f_arrdiv24_fs170_xor1 = f_arrdiv24_fs169_or0 ^ f_arrdiv24_fs170_xor0;
  assign f_arrdiv24_fs170_not1 = ~f_arrdiv24_fs170_xor0;
  assign f_arrdiv24_fs170_and1 = f_arrdiv24_fs170_not1 & f_arrdiv24_fs169_or0;
  assign f_arrdiv24_fs170_or0 = f_arrdiv24_fs170_and1 | f_arrdiv24_fs170_and0;
  assign f_arrdiv24_fs171_xor0 = f_arrdiv24_mux2to1140_xor0 ^ b[3];
  assign f_arrdiv24_fs171_not0 = ~f_arrdiv24_mux2to1140_xor0;
  assign f_arrdiv24_fs171_and0 = f_arrdiv24_fs171_not0 & b[3];
  assign f_arrdiv24_fs171_xor1 = f_arrdiv24_fs170_or0 ^ f_arrdiv24_fs171_xor0;
  assign f_arrdiv24_fs171_not1 = ~f_arrdiv24_fs171_xor0;
  assign f_arrdiv24_fs171_and1 = f_arrdiv24_fs171_not1 & f_arrdiv24_fs170_or0;
  assign f_arrdiv24_fs171_or0 = f_arrdiv24_fs171_and1 | f_arrdiv24_fs171_and0;
  assign f_arrdiv24_fs172_xor0 = f_arrdiv24_mux2to1141_xor0 ^ b[4];
  assign f_arrdiv24_fs172_not0 = ~f_arrdiv24_mux2to1141_xor0;
  assign f_arrdiv24_fs172_and0 = f_arrdiv24_fs172_not0 & b[4];
  assign f_arrdiv24_fs172_xor1 = f_arrdiv24_fs171_or0 ^ f_arrdiv24_fs172_xor0;
  assign f_arrdiv24_fs172_not1 = ~f_arrdiv24_fs172_xor0;
  assign f_arrdiv24_fs172_and1 = f_arrdiv24_fs172_not1 & f_arrdiv24_fs171_or0;
  assign f_arrdiv24_fs172_or0 = f_arrdiv24_fs172_and1 | f_arrdiv24_fs172_and0;
  assign f_arrdiv24_fs173_xor0 = f_arrdiv24_mux2to1142_xor0 ^ b[5];
  assign f_arrdiv24_fs173_not0 = ~f_arrdiv24_mux2to1142_xor0;
  assign f_arrdiv24_fs173_and0 = f_arrdiv24_fs173_not0 & b[5];
  assign f_arrdiv24_fs173_xor1 = f_arrdiv24_fs172_or0 ^ f_arrdiv24_fs173_xor0;
  assign f_arrdiv24_fs173_not1 = ~f_arrdiv24_fs173_xor0;
  assign f_arrdiv24_fs173_and1 = f_arrdiv24_fs173_not1 & f_arrdiv24_fs172_or0;
  assign f_arrdiv24_fs173_or0 = f_arrdiv24_fs173_and1 | f_arrdiv24_fs173_and0;
  assign f_arrdiv24_fs174_xor0 = f_arrdiv24_mux2to1143_xor0 ^ b[6];
  assign f_arrdiv24_fs174_not0 = ~f_arrdiv24_mux2to1143_xor0;
  assign f_arrdiv24_fs174_and0 = f_arrdiv24_fs174_not0 & b[6];
  assign f_arrdiv24_fs174_xor1 = f_arrdiv24_fs173_or0 ^ f_arrdiv24_fs174_xor0;
  assign f_arrdiv24_fs174_not1 = ~f_arrdiv24_fs174_xor0;
  assign f_arrdiv24_fs174_and1 = f_arrdiv24_fs174_not1 & f_arrdiv24_fs173_or0;
  assign f_arrdiv24_fs174_or0 = f_arrdiv24_fs174_and1 | f_arrdiv24_fs174_and0;
  assign f_arrdiv24_fs175_xor0 = f_arrdiv24_mux2to1144_xor0 ^ b[7];
  assign f_arrdiv24_fs175_not0 = ~f_arrdiv24_mux2to1144_xor0;
  assign f_arrdiv24_fs175_and0 = f_arrdiv24_fs175_not0 & b[7];
  assign f_arrdiv24_fs175_xor1 = f_arrdiv24_fs174_or0 ^ f_arrdiv24_fs175_xor0;
  assign f_arrdiv24_fs175_not1 = ~f_arrdiv24_fs175_xor0;
  assign f_arrdiv24_fs175_and1 = f_arrdiv24_fs175_not1 & f_arrdiv24_fs174_or0;
  assign f_arrdiv24_fs175_or0 = f_arrdiv24_fs175_and1 | f_arrdiv24_fs175_and0;
  assign f_arrdiv24_fs176_xor0 = f_arrdiv24_mux2to1145_xor0 ^ b[8];
  assign f_arrdiv24_fs176_not0 = ~f_arrdiv24_mux2to1145_xor0;
  assign f_arrdiv24_fs176_and0 = f_arrdiv24_fs176_not0 & b[8];
  assign f_arrdiv24_fs176_xor1 = f_arrdiv24_fs175_or0 ^ f_arrdiv24_fs176_xor0;
  assign f_arrdiv24_fs176_not1 = ~f_arrdiv24_fs176_xor0;
  assign f_arrdiv24_fs176_and1 = f_arrdiv24_fs176_not1 & f_arrdiv24_fs175_or0;
  assign f_arrdiv24_fs176_or0 = f_arrdiv24_fs176_and1 | f_arrdiv24_fs176_and0;
  assign f_arrdiv24_fs177_xor0 = f_arrdiv24_mux2to1146_xor0 ^ b[9];
  assign f_arrdiv24_fs177_not0 = ~f_arrdiv24_mux2to1146_xor0;
  assign f_arrdiv24_fs177_and0 = f_arrdiv24_fs177_not0 & b[9];
  assign f_arrdiv24_fs177_xor1 = f_arrdiv24_fs176_or0 ^ f_arrdiv24_fs177_xor0;
  assign f_arrdiv24_fs177_not1 = ~f_arrdiv24_fs177_xor0;
  assign f_arrdiv24_fs177_and1 = f_arrdiv24_fs177_not1 & f_arrdiv24_fs176_or0;
  assign f_arrdiv24_fs177_or0 = f_arrdiv24_fs177_and1 | f_arrdiv24_fs177_and0;
  assign f_arrdiv24_fs178_xor0 = f_arrdiv24_mux2to1147_xor0 ^ b[10];
  assign f_arrdiv24_fs178_not0 = ~f_arrdiv24_mux2to1147_xor0;
  assign f_arrdiv24_fs178_and0 = f_arrdiv24_fs178_not0 & b[10];
  assign f_arrdiv24_fs178_xor1 = f_arrdiv24_fs177_or0 ^ f_arrdiv24_fs178_xor0;
  assign f_arrdiv24_fs178_not1 = ~f_arrdiv24_fs178_xor0;
  assign f_arrdiv24_fs178_and1 = f_arrdiv24_fs178_not1 & f_arrdiv24_fs177_or0;
  assign f_arrdiv24_fs178_or0 = f_arrdiv24_fs178_and1 | f_arrdiv24_fs178_and0;
  assign f_arrdiv24_fs179_xor0 = f_arrdiv24_mux2to1148_xor0 ^ b[11];
  assign f_arrdiv24_fs179_not0 = ~f_arrdiv24_mux2to1148_xor0;
  assign f_arrdiv24_fs179_and0 = f_arrdiv24_fs179_not0 & b[11];
  assign f_arrdiv24_fs179_xor1 = f_arrdiv24_fs178_or0 ^ f_arrdiv24_fs179_xor0;
  assign f_arrdiv24_fs179_not1 = ~f_arrdiv24_fs179_xor0;
  assign f_arrdiv24_fs179_and1 = f_arrdiv24_fs179_not1 & f_arrdiv24_fs178_or0;
  assign f_arrdiv24_fs179_or0 = f_arrdiv24_fs179_and1 | f_arrdiv24_fs179_and0;
  assign f_arrdiv24_fs180_xor0 = f_arrdiv24_mux2to1149_xor0 ^ b[12];
  assign f_arrdiv24_fs180_not0 = ~f_arrdiv24_mux2to1149_xor0;
  assign f_arrdiv24_fs180_and0 = f_arrdiv24_fs180_not0 & b[12];
  assign f_arrdiv24_fs180_xor1 = f_arrdiv24_fs179_or0 ^ f_arrdiv24_fs180_xor0;
  assign f_arrdiv24_fs180_not1 = ~f_arrdiv24_fs180_xor0;
  assign f_arrdiv24_fs180_and1 = f_arrdiv24_fs180_not1 & f_arrdiv24_fs179_or0;
  assign f_arrdiv24_fs180_or0 = f_arrdiv24_fs180_and1 | f_arrdiv24_fs180_and0;
  assign f_arrdiv24_fs181_xor0 = f_arrdiv24_mux2to1150_xor0 ^ b[13];
  assign f_arrdiv24_fs181_not0 = ~f_arrdiv24_mux2to1150_xor0;
  assign f_arrdiv24_fs181_and0 = f_arrdiv24_fs181_not0 & b[13];
  assign f_arrdiv24_fs181_xor1 = f_arrdiv24_fs180_or0 ^ f_arrdiv24_fs181_xor0;
  assign f_arrdiv24_fs181_not1 = ~f_arrdiv24_fs181_xor0;
  assign f_arrdiv24_fs181_and1 = f_arrdiv24_fs181_not1 & f_arrdiv24_fs180_or0;
  assign f_arrdiv24_fs181_or0 = f_arrdiv24_fs181_and1 | f_arrdiv24_fs181_and0;
  assign f_arrdiv24_fs182_xor0 = f_arrdiv24_mux2to1151_xor0 ^ b[14];
  assign f_arrdiv24_fs182_not0 = ~f_arrdiv24_mux2to1151_xor0;
  assign f_arrdiv24_fs182_and0 = f_arrdiv24_fs182_not0 & b[14];
  assign f_arrdiv24_fs182_xor1 = f_arrdiv24_fs181_or0 ^ f_arrdiv24_fs182_xor0;
  assign f_arrdiv24_fs182_not1 = ~f_arrdiv24_fs182_xor0;
  assign f_arrdiv24_fs182_and1 = f_arrdiv24_fs182_not1 & f_arrdiv24_fs181_or0;
  assign f_arrdiv24_fs182_or0 = f_arrdiv24_fs182_and1 | f_arrdiv24_fs182_and0;
  assign f_arrdiv24_fs183_xor0 = f_arrdiv24_mux2to1152_xor0 ^ b[15];
  assign f_arrdiv24_fs183_not0 = ~f_arrdiv24_mux2to1152_xor0;
  assign f_arrdiv24_fs183_and0 = f_arrdiv24_fs183_not0 & b[15];
  assign f_arrdiv24_fs183_xor1 = f_arrdiv24_fs182_or0 ^ f_arrdiv24_fs183_xor0;
  assign f_arrdiv24_fs183_not1 = ~f_arrdiv24_fs183_xor0;
  assign f_arrdiv24_fs183_and1 = f_arrdiv24_fs183_not1 & f_arrdiv24_fs182_or0;
  assign f_arrdiv24_fs183_or0 = f_arrdiv24_fs183_and1 | f_arrdiv24_fs183_and0;
  assign f_arrdiv24_fs184_xor0 = f_arrdiv24_mux2to1153_xor0 ^ b[16];
  assign f_arrdiv24_fs184_not0 = ~f_arrdiv24_mux2to1153_xor0;
  assign f_arrdiv24_fs184_and0 = f_arrdiv24_fs184_not0 & b[16];
  assign f_arrdiv24_fs184_xor1 = f_arrdiv24_fs183_or0 ^ f_arrdiv24_fs184_xor0;
  assign f_arrdiv24_fs184_not1 = ~f_arrdiv24_fs184_xor0;
  assign f_arrdiv24_fs184_and1 = f_arrdiv24_fs184_not1 & f_arrdiv24_fs183_or0;
  assign f_arrdiv24_fs184_or0 = f_arrdiv24_fs184_and1 | f_arrdiv24_fs184_and0;
  assign f_arrdiv24_fs185_xor0 = f_arrdiv24_mux2to1154_xor0 ^ b[17];
  assign f_arrdiv24_fs185_not0 = ~f_arrdiv24_mux2to1154_xor0;
  assign f_arrdiv24_fs185_and0 = f_arrdiv24_fs185_not0 & b[17];
  assign f_arrdiv24_fs185_xor1 = f_arrdiv24_fs184_or0 ^ f_arrdiv24_fs185_xor0;
  assign f_arrdiv24_fs185_not1 = ~f_arrdiv24_fs185_xor0;
  assign f_arrdiv24_fs185_and1 = f_arrdiv24_fs185_not1 & f_arrdiv24_fs184_or0;
  assign f_arrdiv24_fs185_or0 = f_arrdiv24_fs185_and1 | f_arrdiv24_fs185_and0;
  assign f_arrdiv24_fs186_xor0 = f_arrdiv24_mux2to1155_xor0 ^ b[18];
  assign f_arrdiv24_fs186_not0 = ~f_arrdiv24_mux2to1155_xor0;
  assign f_arrdiv24_fs186_and0 = f_arrdiv24_fs186_not0 & b[18];
  assign f_arrdiv24_fs186_xor1 = f_arrdiv24_fs185_or0 ^ f_arrdiv24_fs186_xor0;
  assign f_arrdiv24_fs186_not1 = ~f_arrdiv24_fs186_xor0;
  assign f_arrdiv24_fs186_and1 = f_arrdiv24_fs186_not1 & f_arrdiv24_fs185_or0;
  assign f_arrdiv24_fs186_or0 = f_arrdiv24_fs186_and1 | f_arrdiv24_fs186_and0;
  assign f_arrdiv24_fs187_xor0 = f_arrdiv24_mux2to1156_xor0 ^ b[19];
  assign f_arrdiv24_fs187_not0 = ~f_arrdiv24_mux2to1156_xor0;
  assign f_arrdiv24_fs187_and0 = f_arrdiv24_fs187_not0 & b[19];
  assign f_arrdiv24_fs187_xor1 = f_arrdiv24_fs186_or0 ^ f_arrdiv24_fs187_xor0;
  assign f_arrdiv24_fs187_not1 = ~f_arrdiv24_fs187_xor0;
  assign f_arrdiv24_fs187_and1 = f_arrdiv24_fs187_not1 & f_arrdiv24_fs186_or0;
  assign f_arrdiv24_fs187_or0 = f_arrdiv24_fs187_and1 | f_arrdiv24_fs187_and0;
  assign f_arrdiv24_fs188_xor0 = f_arrdiv24_mux2to1157_xor0 ^ b[20];
  assign f_arrdiv24_fs188_not0 = ~f_arrdiv24_mux2to1157_xor0;
  assign f_arrdiv24_fs188_and0 = f_arrdiv24_fs188_not0 & b[20];
  assign f_arrdiv24_fs188_xor1 = f_arrdiv24_fs187_or0 ^ f_arrdiv24_fs188_xor0;
  assign f_arrdiv24_fs188_not1 = ~f_arrdiv24_fs188_xor0;
  assign f_arrdiv24_fs188_and1 = f_arrdiv24_fs188_not1 & f_arrdiv24_fs187_or0;
  assign f_arrdiv24_fs188_or0 = f_arrdiv24_fs188_and1 | f_arrdiv24_fs188_and0;
  assign f_arrdiv24_fs189_xor0 = f_arrdiv24_mux2to1158_xor0 ^ b[21];
  assign f_arrdiv24_fs189_not0 = ~f_arrdiv24_mux2to1158_xor0;
  assign f_arrdiv24_fs189_and0 = f_arrdiv24_fs189_not0 & b[21];
  assign f_arrdiv24_fs189_xor1 = f_arrdiv24_fs188_or0 ^ f_arrdiv24_fs189_xor0;
  assign f_arrdiv24_fs189_not1 = ~f_arrdiv24_fs189_xor0;
  assign f_arrdiv24_fs189_and1 = f_arrdiv24_fs189_not1 & f_arrdiv24_fs188_or0;
  assign f_arrdiv24_fs189_or0 = f_arrdiv24_fs189_and1 | f_arrdiv24_fs189_and0;
  assign f_arrdiv24_fs190_xor0 = f_arrdiv24_mux2to1159_xor0 ^ b[22];
  assign f_arrdiv24_fs190_not0 = ~f_arrdiv24_mux2to1159_xor0;
  assign f_arrdiv24_fs190_and0 = f_arrdiv24_fs190_not0 & b[22];
  assign f_arrdiv24_fs190_xor1 = f_arrdiv24_fs189_or0 ^ f_arrdiv24_fs190_xor0;
  assign f_arrdiv24_fs190_not1 = ~f_arrdiv24_fs190_xor0;
  assign f_arrdiv24_fs190_and1 = f_arrdiv24_fs190_not1 & f_arrdiv24_fs189_or0;
  assign f_arrdiv24_fs190_or0 = f_arrdiv24_fs190_and1 | f_arrdiv24_fs190_and0;
  assign f_arrdiv24_fs191_xor0 = f_arrdiv24_mux2to1160_xor0 ^ b[23];
  assign f_arrdiv24_fs191_not0 = ~f_arrdiv24_mux2to1160_xor0;
  assign f_arrdiv24_fs191_and0 = f_arrdiv24_fs191_not0 & b[23];
  assign f_arrdiv24_fs191_xor1 = f_arrdiv24_fs190_or0 ^ f_arrdiv24_fs191_xor0;
  assign f_arrdiv24_fs191_not1 = ~f_arrdiv24_fs191_xor0;
  assign f_arrdiv24_fs191_and1 = f_arrdiv24_fs191_not1 & f_arrdiv24_fs190_or0;
  assign f_arrdiv24_fs191_or0 = f_arrdiv24_fs191_and1 | f_arrdiv24_fs191_and0;
  assign f_arrdiv24_mux2to1161_and0 = a[16] & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1161_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1161_and1 = f_arrdiv24_fs168_xor0 & f_arrdiv24_mux2to1161_not0;
  assign f_arrdiv24_mux2to1161_xor0 = f_arrdiv24_mux2to1161_and0 ^ f_arrdiv24_mux2to1161_and1;
  assign f_arrdiv24_mux2to1162_and0 = f_arrdiv24_mux2to1138_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1162_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1162_and1 = f_arrdiv24_fs169_xor1 & f_arrdiv24_mux2to1162_not0;
  assign f_arrdiv24_mux2to1162_xor0 = f_arrdiv24_mux2to1162_and0 ^ f_arrdiv24_mux2to1162_and1;
  assign f_arrdiv24_mux2to1163_and0 = f_arrdiv24_mux2to1139_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1163_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1163_and1 = f_arrdiv24_fs170_xor1 & f_arrdiv24_mux2to1163_not0;
  assign f_arrdiv24_mux2to1163_xor0 = f_arrdiv24_mux2to1163_and0 ^ f_arrdiv24_mux2to1163_and1;
  assign f_arrdiv24_mux2to1164_and0 = f_arrdiv24_mux2to1140_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1164_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1164_and1 = f_arrdiv24_fs171_xor1 & f_arrdiv24_mux2to1164_not0;
  assign f_arrdiv24_mux2to1164_xor0 = f_arrdiv24_mux2to1164_and0 ^ f_arrdiv24_mux2to1164_and1;
  assign f_arrdiv24_mux2to1165_and0 = f_arrdiv24_mux2to1141_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1165_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1165_and1 = f_arrdiv24_fs172_xor1 & f_arrdiv24_mux2to1165_not0;
  assign f_arrdiv24_mux2to1165_xor0 = f_arrdiv24_mux2to1165_and0 ^ f_arrdiv24_mux2to1165_and1;
  assign f_arrdiv24_mux2to1166_and0 = f_arrdiv24_mux2to1142_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1166_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1166_and1 = f_arrdiv24_fs173_xor1 & f_arrdiv24_mux2to1166_not0;
  assign f_arrdiv24_mux2to1166_xor0 = f_arrdiv24_mux2to1166_and0 ^ f_arrdiv24_mux2to1166_and1;
  assign f_arrdiv24_mux2to1167_and0 = f_arrdiv24_mux2to1143_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1167_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1167_and1 = f_arrdiv24_fs174_xor1 & f_arrdiv24_mux2to1167_not0;
  assign f_arrdiv24_mux2to1167_xor0 = f_arrdiv24_mux2to1167_and0 ^ f_arrdiv24_mux2to1167_and1;
  assign f_arrdiv24_mux2to1168_and0 = f_arrdiv24_mux2to1144_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1168_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1168_and1 = f_arrdiv24_fs175_xor1 & f_arrdiv24_mux2to1168_not0;
  assign f_arrdiv24_mux2to1168_xor0 = f_arrdiv24_mux2to1168_and0 ^ f_arrdiv24_mux2to1168_and1;
  assign f_arrdiv24_mux2to1169_and0 = f_arrdiv24_mux2to1145_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1169_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1169_and1 = f_arrdiv24_fs176_xor1 & f_arrdiv24_mux2to1169_not0;
  assign f_arrdiv24_mux2to1169_xor0 = f_arrdiv24_mux2to1169_and0 ^ f_arrdiv24_mux2to1169_and1;
  assign f_arrdiv24_mux2to1170_and0 = f_arrdiv24_mux2to1146_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1170_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1170_and1 = f_arrdiv24_fs177_xor1 & f_arrdiv24_mux2to1170_not0;
  assign f_arrdiv24_mux2to1170_xor0 = f_arrdiv24_mux2to1170_and0 ^ f_arrdiv24_mux2to1170_and1;
  assign f_arrdiv24_mux2to1171_and0 = f_arrdiv24_mux2to1147_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1171_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1171_and1 = f_arrdiv24_fs178_xor1 & f_arrdiv24_mux2to1171_not0;
  assign f_arrdiv24_mux2to1171_xor0 = f_arrdiv24_mux2to1171_and0 ^ f_arrdiv24_mux2to1171_and1;
  assign f_arrdiv24_mux2to1172_and0 = f_arrdiv24_mux2to1148_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1172_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1172_and1 = f_arrdiv24_fs179_xor1 & f_arrdiv24_mux2to1172_not0;
  assign f_arrdiv24_mux2to1172_xor0 = f_arrdiv24_mux2to1172_and0 ^ f_arrdiv24_mux2to1172_and1;
  assign f_arrdiv24_mux2to1173_and0 = f_arrdiv24_mux2to1149_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1173_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1173_and1 = f_arrdiv24_fs180_xor1 & f_arrdiv24_mux2to1173_not0;
  assign f_arrdiv24_mux2to1173_xor0 = f_arrdiv24_mux2to1173_and0 ^ f_arrdiv24_mux2to1173_and1;
  assign f_arrdiv24_mux2to1174_and0 = f_arrdiv24_mux2to1150_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1174_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1174_and1 = f_arrdiv24_fs181_xor1 & f_arrdiv24_mux2to1174_not0;
  assign f_arrdiv24_mux2to1174_xor0 = f_arrdiv24_mux2to1174_and0 ^ f_arrdiv24_mux2to1174_and1;
  assign f_arrdiv24_mux2to1175_and0 = f_arrdiv24_mux2to1151_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1175_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1175_and1 = f_arrdiv24_fs182_xor1 & f_arrdiv24_mux2to1175_not0;
  assign f_arrdiv24_mux2to1175_xor0 = f_arrdiv24_mux2to1175_and0 ^ f_arrdiv24_mux2to1175_and1;
  assign f_arrdiv24_mux2to1176_and0 = f_arrdiv24_mux2to1152_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1176_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1176_and1 = f_arrdiv24_fs183_xor1 & f_arrdiv24_mux2to1176_not0;
  assign f_arrdiv24_mux2to1176_xor0 = f_arrdiv24_mux2to1176_and0 ^ f_arrdiv24_mux2to1176_and1;
  assign f_arrdiv24_mux2to1177_and0 = f_arrdiv24_mux2to1153_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1177_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1177_and1 = f_arrdiv24_fs184_xor1 & f_arrdiv24_mux2to1177_not0;
  assign f_arrdiv24_mux2to1177_xor0 = f_arrdiv24_mux2to1177_and0 ^ f_arrdiv24_mux2to1177_and1;
  assign f_arrdiv24_mux2to1178_and0 = f_arrdiv24_mux2to1154_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1178_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1178_and1 = f_arrdiv24_fs185_xor1 & f_arrdiv24_mux2to1178_not0;
  assign f_arrdiv24_mux2to1178_xor0 = f_arrdiv24_mux2to1178_and0 ^ f_arrdiv24_mux2to1178_and1;
  assign f_arrdiv24_mux2to1179_and0 = f_arrdiv24_mux2to1155_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1179_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1179_and1 = f_arrdiv24_fs186_xor1 & f_arrdiv24_mux2to1179_not0;
  assign f_arrdiv24_mux2to1179_xor0 = f_arrdiv24_mux2to1179_and0 ^ f_arrdiv24_mux2to1179_and1;
  assign f_arrdiv24_mux2to1180_and0 = f_arrdiv24_mux2to1156_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1180_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1180_and1 = f_arrdiv24_fs187_xor1 & f_arrdiv24_mux2to1180_not0;
  assign f_arrdiv24_mux2to1180_xor0 = f_arrdiv24_mux2to1180_and0 ^ f_arrdiv24_mux2to1180_and1;
  assign f_arrdiv24_mux2to1181_and0 = f_arrdiv24_mux2to1157_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1181_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1181_and1 = f_arrdiv24_fs188_xor1 & f_arrdiv24_mux2to1181_not0;
  assign f_arrdiv24_mux2to1181_xor0 = f_arrdiv24_mux2to1181_and0 ^ f_arrdiv24_mux2to1181_and1;
  assign f_arrdiv24_mux2to1182_and0 = f_arrdiv24_mux2to1158_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1182_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1182_and1 = f_arrdiv24_fs189_xor1 & f_arrdiv24_mux2to1182_not0;
  assign f_arrdiv24_mux2to1182_xor0 = f_arrdiv24_mux2to1182_and0 ^ f_arrdiv24_mux2to1182_and1;
  assign f_arrdiv24_mux2to1183_and0 = f_arrdiv24_mux2to1159_xor0 & f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1183_not0 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_mux2to1183_and1 = f_arrdiv24_fs190_xor1 & f_arrdiv24_mux2to1183_not0;
  assign f_arrdiv24_mux2to1183_xor0 = f_arrdiv24_mux2to1183_and0 ^ f_arrdiv24_mux2to1183_and1;
  assign f_arrdiv24_not7 = ~f_arrdiv24_fs191_or0;
  assign f_arrdiv24_fs192_xor0 = a[15] ^ b[0];
  assign f_arrdiv24_fs192_not0 = ~a[15];
  assign f_arrdiv24_fs192_and0 = f_arrdiv24_fs192_not0 & b[0];
  assign f_arrdiv24_fs192_not1 = ~f_arrdiv24_fs192_xor0;
  assign f_arrdiv24_fs193_xor0 = f_arrdiv24_mux2to1161_xor0 ^ b[1];
  assign f_arrdiv24_fs193_not0 = ~f_arrdiv24_mux2to1161_xor0;
  assign f_arrdiv24_fs193_and0 = f_arrdiv24_fs193_not0 & b[1];
  assign f_arrdiv24_fs193_xor1 = f_arrdiv24_fs192_and0 ^ f_arrdiv24_fs193_xor0;
  assign f_arrdiv24_fs193_not1 = ~f_arrdiv24_fs193_xor0;
  assign f_arrdiv24_fs193_and1 = f_arrdiv24_fs193_not1 & f_arrdiv24_fs192_and0;
  assign f_arrdiv24_fs193_or0 = f_arrdiv24_fs193_and1 | f_arrdiv24_fs193_and0;
  assign f_arrdiv24_fs194_xor0 = f_arrdiv24_mux2to1162_xor0 ^ b[2];
  assign f_arrdiv24_fs194_not0 = ~f_arrdiv24_mux2to1162_xor0;
  assign f_arrdiv24_fs194_and0 = f_arrdiv24_fs194_not0 & b[2];
  assign f_arrdiv24_fs194_xor1 = f_arrdiv24_fs193_or0 ^ f_arrdiv24_fs194_xor0;
  assign f_arrdiv24_fs194_not1 = ~f_arrdiv24_fs194_xor0;
  assign f_arrdiv24_fs194_and1 = f_arrdiv24_fs194_not1 & f_arrdiv24_fs193_or0;
  assign f_arrdiv24_fs194_or0 = f_arrdiv24_fs194_and1 | f_arrdiv24_fs194_and0;
  assign f_arrdiv24_fs195_xor0 = f_arrdiv24_mux2to1163_xor0 ^ b[3];
  assign f_arrdiv24_fs195_not0 = ~f_arrdiv24_mux2to1163_xor0;
  assign f_arrdiv24_fs195_and0 = f_arrdiv24_fs195_not0 & b[3];
  assign f_arrdiv24_fs195_xor1 = f_arrdiv24_fs194_or0 ^ f_arrdiv24_fs195_xor0;
  assign f_arrdiv24_fs195_not1 = ~f_arrdiv24_fs195_xor0;
  assign f_arrdiv24_fs195_and1 = f_arrdiv24_fs195_not1 & f_arrdiv24_fs194_or0;
  assign f_arrdiv24_fs195_or0 = f_arrdiv24_fs195_and1 | f_arrdiv24_fs195_and0;
  assign f_arrdiv24_fs196_xor0 = f_arrdiv24_mux2to1164_xor0 ^ b[4];
  assign f_arrdiv24_fs196_not0 = ~f_arrdiv24_mux2to1164_xor0;
  assign f_arrdiv24_fs196_and0 = f_arrdiv24_fs196_not0 & b[4];
  assign f_arrdiv24_fs196_xor1 = f_arrdiv24_fs195_or0 ^ f_arrdiv24_fs196_xor0;
  assign f_arrdiv24_fs196_not1 = ~f_arrdiv24_fs196_xor0;
  assign f_arrdiv24_fs196_and1 = f_arrdiv24_fs196_not1 & f_arrdiv24_fs195_or0;
  assign f_arrdiv24_fs196_or0 = f_arrdiv24_fs196_and1 | f_arrdiv24_fs196_and0;
  assign f_arrdiv24_fs197_xor0 = f_arrdiv24_mux2to1165_xor0 ^ b[5];
  assign f_arrdiv24_fs197_not0 = ~f_arrdiv24_mux2to1165_xor0;
  assign f_arrdiv24_fs197_and0 = f_arrdiv24_fs197_not0 & b[5];
  assign f_arrdiv24_fs197_xor1 = f_arrdiv24_fs196_or0 ^ f_arrdiv24_fs197_xor0;
  assign f_arrdiv24_fs197_not1 = ~f_arrdiv24_fs197_xor0;
  assign f_arrdiv24_fs197_and1 = f_arrdiv24_fs197_not1 & f_arrdiv24_fs196_or0;
  assign f_arrdiv24_fs197_or0 = f_arrdiv24_fs197_and1 | f_arrdiv24_fs197_and0;
  assign f_arrdiv24_fs198_xor0 = f_arrdiv24_mux2to1166_xor0 ^ b[6];
  assign f_arrdiv24_fs198_not0 = ~f_arrdiv24_mux2to1166_xor0;
  assign f_arrdiv24_fs198_and0 = f_arrdiv24_fs198_not0 & b[6];
  assign f_arrdiv24_fs198_xor1 = f_arrdiv24_fs197_or0 ^ f_arrdiv24_fs198_xor0;
  assign f_arrdiv24_fs198_not1 = ~f_arrdiv24_fs198_xor0;
  assign f_arrdiv24_fs198_and1 = f_arrdiv24_fs198_not1 & f_arrdiv24_fs197_or0;
  assign f_arrdiv24_fs198_or0 = f_arrdiv24_fs198_and1 | f_arrdiv24_fs198_and0;
  assign f_arrdiv24_fs199_xor0 = f_arrdiv24_mux2to1167_xor0 ^ b[7];
  assign f_arrdiv24_fs199_not0 = ~f_arrdiv24_mux2to1167_xor0;
  assign f_arrdiv24_fs199_and0 = f_arrdiv24_fs199_not0 & b[7];
  assign f_arrdiv24_fs199_xor1 = f_arrdiv24_fs198_or0 ^ f_arrdiv24_fs199_xor0;
  assign f_arrdiv24_fs199_not1 = ~f_arrdiv24_fs199_xor0;
  assign f_arrdiv24_fs199_and1 = f_arrdiv24_fs199_not1 & f_arrdiv24_fs198_or0;
  assign f_arrdiv24_fs199_or0 = f_arrdiv24_fs199_and1 | f_arrdiv24_fs199_and0;
  assign f_arrdiv24_fs200_xor0 = f_arrdiv24_mux2to1168_xor0 ^ b[8];
  assign f_arrdiv24_fs200_not0 = ~f_arrdiv24_mux2to1168_xor0;
  assign f_arrdiv24_fs200_and0 = f_arrdiv24_fs200_not0 & b[8];
  assign f_arrdiv24_fs200_xor1 = f_arrdiv24_fs199_or0 ^ f_arrdiv24_fs200_xor0;
  assign f_arrdiv24_fs200_not1 = ~f_arrdiv24_fs200_xor0;
  assign f_arrdiv24_fs200_and1 = f_arrdiv24_fs200_not1 & f_arrdiv24_fs199_or0;
  assign f_arrdiv24_fs200_or0 = f_arrdiv24_fs200_and1 | f_arrdiv24_fs200_and0;
  assign f_arrdiv24_fs201_xor0 = f_arrdiv24_mux2to1169_xor0 ^ b[9];
  assign f_arrdiv24_fs201_not0 = ~f_arrdiv24_mux2to1169_xor0;
  assign f_arrdiv24_fs201_and0 = f_arrdiv24_fs201_not0 & b[9];
  assign f_arrdiv24_fs201_xor1 = f_arrdiv24_fs200_or0 ^ f_arrdiv24_fs201_xor0;
  assign f_arrdiv24_fs201_not1 = ~f_arrdiv24_fs201_xor0;
  assign f_arrdiv24_fs201_and1 = f_arrdiv24_fs201_not1 & f_arrdiv24_fs200_or0;
  assign f_arrdiv24_fs201_or0 = f_arrdiv24_fs201_and1 | f_arrdiv24_fs201_and0;
  assign f_arrdiv24_fs202_xor0 = f_arrdiv24_mux2to1170_xor0 ^ b[10];
  assign f_arrdiv24_fs202_not0 = ~f_arrdiv24_mux2to1170_xor0;
  assign f_arrdiv24_fs202_and0 = f_arrdiv24_fs202_not0 & b[10];
  assign f_arrdiv24_fs202_xor1 = f_arrdiv24_fs201_or0 ^ f_arrdiv24_fs202_xor0;
  assign f_arrdiv24_fs202_not1 = ~f_arrdiv24_fs202_xor0;
  assign f_arrdiv24_fs202_and1 = f_arrdiv24_fs202_not1 & f_arrdiv24_fs201_or0;
  assign f_arrdiv24_fs202_or0 = f_arrdiv24_fs202_and1 | f_arrdiv24_fs202_and0;
  assign f_arrdiv24_fs203_xor0 = f_arrdiv24_mux2to1171_xor0 ^ b[11];
  assign f_arrdiv24_fs203_not0 = ~f_arrdiv24_mux2to1171_xor0;
  assign f_arrdiv24_fs203_and0 = f_arrdiv24_fs203_not0 & b[11];
  assign f_arrdiv24_fs203_xor1 = f_arrdiv24_fs202_or0 ^ f_arrdiv24_fs203_xor0;
  assign f_arrdiv24_fs203_not1 = ~f_arrdiv24_fs203_xor0;
  assign f_arrdiv24_fs203_and1 = f_arrdiv24_fs203_not1 & f_arrdiv24_fs202_or0;
  assign f_arrdiv24_fs203_or0 = f_arrdiv24_fs203_and1 | f_arrdiv24_fs203_and0;
  assign f_arrdiv24_fs204_xor0 = f_arrdiv24_mux2to1172_xor0 ^ b[12];
  assign f_arrdiv24_fs204_not0 = ~f_arrdiv24_mux2to1172_xor0;
  assign f_arrdiv24_fs204_and0 = f_arrdiv24_fs204_not0 & b[12];
  assign f_arrdiv24_fs204_xor1 = f_arrdiv24_fs203_or0 ^ f_arrdiv24_fs204_xor0;
  assign f_arrdiv24_fs204_not1 = ~f_arrdiv24_fs204_xor0;
  assign f_arrdiv24_fs204_and1 = f_arrdiv24_fs204_not1 & f_arrdiv24_fs203_or0;
  assign f_arrdiv24_fs204_or0 = f_arrdiv24_fs204_and1 | f_arrdiv24_fs204_and0;
  assign f_arrdiv24_fs205_xor0 = f_arrdiv24_mux2to1173_xor0 ^ b[13];
  assign f_arrdiv24_fs205_not0 = ~f_arrdiv24_mux2to1173_xor0;
  assign f_arrdiv24_fs205_and0 = f_arrdiv24_fs205_not0 & b[13];
  assign f_arrdiv24_fs205_xor1 = f_arrdiv24_fs204_or0 ^ f_arrdiv24_fs205_xor0;
  assign f_arrdiv24_fs205_not1 = ~f_arrdiv24_fs205_xor0;
  assign f_arrdiv24_fs205_and1 = f_arrdiv24_fs205_not1 & f_arrdiv24_fs204_or0;
  assign f_arrdiv24_fs205_or0 = f_arrdiv24_fs205_and1 | f_arrdiv24_fs205_and0;
  assign f_arrdiv24_fs206_xor0 = f_arrdiv24_mux2to1174_xor0 ^ b[14];
  assign f_arrdiv24_fs206_not0 = ~f_arrdiv24_mux2to1174_xor0;
  assign f_arrdiv24_fs206_and0 = f_arrdiv24_fs206_not0 & b[14];
  assign f_arrdiv24_fs206_xor1 = f_arrdiv24_fs205_or0 ^ f_arrdiv24_fs206_xor0;
  assign f_arrdiv24_fs206_not1 = ~f_arrdiv24_fs206_xor0;
  assign f_arrdiv24_fs206_and1 = f_arrdiv24_fs206_not1 & f_arrdiv24_fs205_or0;
  assign f_arrdiv24_fs206_or0 = f_arrdiv24_fs206_and1 | f_arrdiv24_fs206_and0;
  assign f_arrdiv24_fs207_xor0 = f_arrdiv24_mux2to1175_xor0 ^ b[15];
  assign f_arrdiv24_fs207_not0 = ~f_arrdiv24_mux2to1175_xor0;
  assign f_arrdiv24_fs207_and0 = f_arrdiv24_fs207_not0 & b[15];
  assign f_arrdiv24_fs207_xor1 = f_arrdiv24_fs206_or0 ^ f_arrdiv24_fs207_xor0;
  assign f_arrdiv24_fs207_not1 = ~f_arrdiv24_fs207_xor0;
  assign f_arrdiv24_fs207_and1 = f_arrdiv24_fs207_not1 & f_arrdiv24_fs206_or0;
  assign f_arrdiv24_fs207_or0 = f_arrdiv24_fs207_and1 | f_arrdiv24_fs207_and0;
  assign f_arrdiv24_fs208_xor0 = f_arrdiv24_mux2to1176_xor0 ^ b[16];
  assign f_arrdiv24_fs208_not0 = ~f_arrdiv24_mux2to1176_xor0;
  assign f_arrdiv24_fs208_and0 = f_arrdiv24_fs208_not0 & b[16];
  assign f_arrdiv24_fs208_xor1 = f_arrdiv24_fs207_or0 ^ f_arrdiv24_fs208_xor0;
  assign f_arrdiv24_fs208_not1 = ~f_arrdiv24_fs208_xor0;
  assign f_arrdiv24_fs208_and1 = f_arrdiv24_fs208_not1 & f_arrdiv24_fs207_or0;
  assign f_arrdiv24_fs208_or0 = f_arrdiv24_fs208_and1 | f_arrdiv24_fs208_and0;
  assign f_arrdiv24_fs209_xor0 = f_arrdiv24_mux2to1177_xor0 ^ b[17];
  assign f_arrdiv24_fs209_not0 = ~f_arrdiv24_mux2to1177_xor0;
  assign f_arrdiv24_fs209_and0 = f_arrdiv24_fs209_not0 & b[17];
  assign f_arrdiv24_fs209_xor1 = f_arrdiv24_fs208_or0 ^ f_arrdiv24_fs209_xor0;
  assign f_arrdiv24_fs209_not1 = ~f_arrdiv24_fs209_xor0;
  assign f_arrdiv24_fs209_and1 = f_arrdiv24_fs209_not1 & f_arrdiv24_fs208_or0;
  assign f_arrdiv24_fs209_or0 = f_arrdiv24_fs209_and1 | f_arrdiv24_fs209_and0;
  assign f_arrdiv24_fs210_xor0 = f_arrdiv24_mux2to1178_xor0 ^ b[18];
  assign f_arrdiv24_fs210_not0 = ~f_arrdiv24_mux2to1178_xor0;
  assign f_arrdiv24_fs210_and0 = f_arrdiv24_fs210_not0 & b[18];
  assign f_arrdiv24_fs210_xor1 = f_arrdiv24_fs209_or0 ^ f_arrdiv24_fs210_xor0;
  assign f_arrdiv24_fs210_not1 = ~f_arrdiv24_fs210_xor0;
  assign f_arrdiv24_fs210_and1 = f_arrdiv24_fs210_not1 & f_arrdiv24_fs209_or0;
  assign f_arrdiv24_fs210_or0 = f_arrdiv24_fs210_and1 | f_arrdiv24_fs210_and0;
  assign f_arrdiv24_fs211_xor0 = f_arrdiv24_mux2to1179_xor0 ^ b[19];
  assign f_arrdiv24_fs211_not0 = ~f_arrdiv24_mux2to1179_xor0;
  assign f_arrdiv24_fs211_and0 = f_arrdiv24_fs211_not0 & b[19];
  assign f_arrdiv24_fs211_xor1 = f_arrdiv24_fs210_or0 ^ f_arrdiv24_fs211_xor0;
  assign f_arrdiv24_fs211_not1 = ~f_arrdiv24_fs211_xor0;
  assign f_arrdiv24_fs211_and1 = f_arrdiv24_fs211_not1 & f_arrdiv24_fs210_or0;
  assign f_arrdiv24_fs211_or0 = f_arrdiv24_fs211_and1 | f_arrdiv24_fs211_and0;
  assign f_arrdiv24_fs212_xor0 = f_arrdiv24_mux2to1180_xor0 ^ b[20];
  assign f_arrdiv24_fs212_not0 = ~f_arrdiv24_mux2to1180_xor0;
  assign f_arrdiv24_fs212_and0 = f_arrdiv24_fs212_not0 & b[20];
  assign f_arrdiv24_fs212_xor1 = f_arrdiv24_fs211_or0 ^ f_arrdiv24_fs212_xor0;
  assign f_arrdiv24_fs212_not1 = ~f_arrdiv24_fs212_xor0;
  assign f_arrdiv24_fs212_and1 = f_arrdiv24_fs212_not1 & f_arrdiv24_fs211_or0;
  assign f_arrdiv24_fs212_or0 = f_arrdiv24_fs212_and1 | f_arrdiv24_fs212_and0;
  assign f_arrdiv24_fs213_xor0 = f_arrdiv24_mux2to1181_xor0 ^ b[21];
  assign f_arrdiv24_fs213_not0 = ~f_arrdiv24_mux2to1181_xor0;
  assign f_arrdiv24_fs213_and0 = f_arrdiv24_fs213_not0 & b[21];
  assign f_arrdiv24_fs213_xor1 = f_arrdiv24_fs212_or0 ^ f_arrdiv24_fs213_xor0;
  assign f_arrdiv24_fs213_not1 = ~f_arrdiv24_fs213_xor0;
  assign f_arrdiv24_fs213_and1 = f_arrdiv24_fs213_not1 & f_arrdiv24_fs212_or0;
  assign f_arrdiv24_fs213_or0 = f_arrdiv24_fs213_and1 | f_arrdiv24_fs213_and0;
  assign f_arrdiv24_fs214_xor0 = f_arrdiv24_mux2to1182_xor0 ^ b[22];
  assign f_arrdiv24_fs214_not0 = ~f_arrdiv24_mux2to1182_xor0;
  assign f_arrdiv24_fs214_and0 = f_arrdiv24_fs214_not0 & b[22];
  assign f_arrdiv24_fs214_xor1 = f_arrdiv24_fs213_or0 ^ f_arrdiv24_fs214_xor0;
  assign f_arrdiv24_fs214_not1 = ~f_arrdiv24_fs214_xor0;
  assign f_arrdiv24_fs214_and1 = f_arrdiv24_fs214_not1 & f_arrdiv24_fs213_or0;
  assign f_arrdiv24_fs214_or0 = f_arrdiv24_fs214_and1 | f_arrdiv24_fs214_and0;
  assign f_arrdiv24_fs215_xor0 = f_arrdiv24_mux2to1183_xor0 ^ b[23];
  assign f_arrdiv24_fs215_not0 = ~f_arrdiv24_mux2to1183_xor0;
  assign f_arrdiv24_fs215_and0 = f_arrdiv24_fs215_not0 & b[23];
  assign f_arrdiv24_fs215_xor1 = f_arrdiv24_fs214_or0 ^ f_arrdiv24_fs215_xor0;
  assign f_arrdiv24_fs215_not1 = ~f_arrdiv24_fs215_xor0;
  assign f_arrdiv24_fs215_and1 = f_arrdiv24_fs215_not1 & f_arrdiv24_fs214_or0;
  assign f_arrdiv24_fs215_or0 = f_arrdiv24_fs215_and1 | f_arrdiv24_fs215_and0;
  assign f_arrdiv24_mux2to1184_and0 = a[15] & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1184_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1184_and1 = f_arrdiv24_fs192_xor0 & f_arrdiv24_mux2to1184_not0;
  assign f_arrdiv24_mux2to1184_xor0 = f_arrdiv24_mux2to1184_and0 ^ f_arrdiv24_mux2to1184_and1;
  assign f_arrdiv24_mux2to1185_and0 = f_arrdiv24_mux2to1161_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1185_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1185_and1 = f_arrdiv24_fs193_xor1 & f_arrdiv24_mux2to1185_not0;
  assign f_arrdiv24_mux2to1185_xor0 = f_arrdiv24_mux2to1185_and0 ^ f_arrdiv24_mux2to1185_and1;
  assign f_arrdiv24_mux2to1186_and0 = f_arrdiv24_mux2to1162_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1186_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1186_and1 = f_arrdiv24_fs194_xor1 & f_arrdiv24_mux2to1186_not0;
  assign f_arrdiv24_mux2to1186_xor0 = f_arrdiv24_mux2to1186_and0 ^ f_arrdiv24_mux2to1186_and1;
  assign f_arrdiv24_mux2to1187_and0 = f_arrdiv24_mux2to1163_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1187_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1187_and1 = f_arrdiv24_fs195_xor1 & f_arrdiv24_mux2to1187_not0;
  assign f_arrdiv24_mux2to1187_xor0 = f_arrdiv24_mux2to1187_and0 ^ f_arrdiv24_mux2to1187_and1;
  assign f_arrdiv24_mux2to1188_and0 = f_arrdiv24_mux2to1164_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1188_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1188_and1 = f_arrdiv24_fs196_xor1 & f_arrdiv24_mux2to1188_not0;
  assign f_arrdiv24_mux2to1188_xor0 = f_arrdiv24_mux2to1188_and0 ^ f_arrdiv24_mux2to1188_and1;
  assign f_arrdiv24_mux2to1189_and0 = f_arrdiv24_mux2to1165_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1189_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1189_and1 = f_arrdiv24_fs197_xor1 & f_arrdiv24_mux2to1189_not0;
  assign f_arrdiv24_mux2to1189_xor0 = f_arrdiv24_mux2to1189_and0 ^ f_arrdiv24_mux2to1189_and1;
  assign f_arrdiv24_mux2to1190_and0 = f_arrdiv24_mux2to1166_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1190_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1190_and1 = f_arrdiv24_fs198_xor1 & f_arrdiv24_mux2to1190_not0;
  assign f_arrdiv24_mux2to1190_xor0 = f_arrdiv24_mux2to1190_and0 ^ f_arrdiv24_mux2to1190_and1;
  assign f_arrdiv24_mux2to1191_and0 = f_arrdiv24_mux2to1167_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1191_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1191_and1 = f_arrdiv24_fs199_xor1 & f_arrdiv24_mux2to1191_not0;
  assign f_arrdiv24_mux2to1191_xor0 = f_arrdiv24_mux2to1191_and0 ^ f_arrdiv24_mux2to1191_and1;
  assign f_arrdiv24_mux2to1192_and0 = f_arrdiv24_mux2to1168_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1192_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1192_and1 = f_arrdiv24_fs200_xor1 & f_arrdiv24_mux2to1192_not0;
  assign f_arrdiv24_mux2to1192_xor0 = f_arrdiv24_mux2to1192_and0 ^ f_arrdiv24_mux2to1192_and1;
  assign f_arrdiv24_mux2to1193_and0 = f_arrdiv24_mux2to1169_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1193_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1193_and1 = f_arrdiv24_fs201_xor1 & f_arrdiv24_mux2to1193_not0;
  assign f_arrdiv24_mux2to1193_xor0 = f_arrdiv24_mux2to1193_and0 ^ f_arrdiv24_mux2to1193_and1;
  assign f_arrdiv24_mux2to1194_and0 = f_arrdiv24_mux2to1170_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1194_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1194_and1 = f_arrdiv24_fs202_xor1 & f_arrdiv24_mux2to1194_not0;
  assign f_arrdiv24_mux2to1194_xor0 = f_arrdiv24_mux2to1194_and0 ^ f_arrdiv24_mux2to1194_and1;
  assign f_arrdiv24_mux2to1195_and0 = f_arrdiv24_mux2to1171_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1195_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1195_and1 = f_arrdiv24_fs203_xor1 & f_arrdiv24_mux2to1195_not0;
  assign f_arrdiv24_mux2to1195_xor0 = f_arrdiv24_mux2to1195_and0 ^ f_arrdiv24_mux2to1195_and1;
  assign f_arrdiv24_mux2to1196_and0 = f_arrdiv24_mux2to1172_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1196_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1196_and1 = f_arrdiv24_fs204_xor1 & f_arrdiv24_mux2to1196_not0;
  assign f_arrdiv24_mux2to1196_xor0 = f_arrdiv24_mux2to1196_and0 ^ f_arrdiv24_mux2to1196_and1;
  assign f_arrdiv24_mux2to1197_and0 = f_arrdiv24_mux2to1173_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1197_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1197_and1 = f_arrdiv24_fs205_xor1 & f_arrdiv24_mux2to1197_not0;
  assign f_arrdiv24_mux2to1197_xor0 = f_arrdiv24_mux2to1197_and0 ^ f_arrdiv24_mux2to1197_and1;
  assign f_arrdiv24_mux2to1198_and0 = f_arrdiv24_mux2to1174_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1198_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1198_and1 = f_arrdiv24_fs206_xor1 & f_arrdiv24_mux2to1198_not0;
  assign f_arrdiv24_mux2to1198_xor0 = f_arrdiv24_mux2to1198_and0 ^ f_arrdiv24_mux2to1198_and1;
  assign f_arrdiv24_mux2to1199_and0 = f_arrdiv24_mux2to1175_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1199_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1199_and1 = f_arrdiv24_fs207_xor1 & f_arrdiv24_mux2to1199_not0;
  assign f_arrdiv24_mux2to1199_xor0 = f_arrdiv24_mux2to1199_and0 ^ f_arrdiv24_mux2to1199_and1;
  assign f_arrdiv24_mux2to1200_and0 = f_arrdiv24_mux2to1176_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1200_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1200_and1 = f_arrdiv24_fs208_xor1 & f_arrdiv24_mux2to1200_not0;
  assign f_arrdiv24_mux2to1200_xor0 = f_arrdiv24_mux2to1200_and0 ^ f_arrdiv24_mux2to1200_and1;
  assign f_arrdiv24_mux2to1201_and0 = f_arrdiv24_mux2to1177_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1201_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1201_and1 = f_arrdiv24_fs209_xor1 & f_arrdiv24_mux2to1201_not0;
  assign f_arrdiv24_mux2to1201_xor0 = f_arrdiv24_mux2to1201_and0 ^ f_arrdiv24_mux2to1201_and1;
  assign f_arrdiv24_mux2to1202_and0 = f_arrdiv24_mux2to1178_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1202_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1202_and1 = f_arrdiv24_fs210_xor1 & f_arrdiv24_mux2to1202_not0;
  assign f_arrdiv24_mux2to1202_xor0 = f_arrdiv24_mux2to1202_and0 ^ f_arrdiv24_mux2to1202_and1;
  assign f_arrdiv24_mux2to1203_and0 = f_arrdiv24_mux2to1179_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1203_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1203_and1 = f_arrdiv24_fs211_xor1 & f_arrdiv24_mux2to1203_not0;
  assign f_arrdiv24_mux2to1203_xor0 = f_arrdiv24_mux2to1203_and0 ^ f_arrdiv24_mux2to1203_and1;
  assign f_arrdiv24_mux2to1204_and0 = f_arrdiv24_mux2to1180_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1204_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1204_and1 = f_arrdiv24_fs212_xor1 & f_arrdiv24_mux2to1204_not0;
  assign f_arrdiv24_mux2to1204_xor0 = f_arrdiv24_mux2to1204_and0 ^ f_arrdiv24_mux2to1204_and1;
  assign f_arrdiv24_mux2to1205_and0 = f_arrdiv24_mux2to1181_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1205_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1205_and1 = f_arrdiv24_fs213_xor1 & f_arrdiv24_mux2to1205_not0;
  assign f_arrdiv24_mux2to1205_xor0 = f_arrdiv24_mux2to1205_and0 ^ f_arrdiv24_mux2to1205_and1;
  assign f_arrdiv24_mux2to1206_and0 = f_arrdiv24_mux2to1182_xor0 & f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1206_not0 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_mux2to1206_and1 = f_arrdiv24_fs214_xor1 & f_arrdiv24_mux2to1206_not0;
  assign f_arrdiv24_mux2to1206_xor0 = f_arrdiv24_mux2to1206_and0 ^ f_arrdiv24_mux2to1206_and1;
  assign f_arrdiv24_not8 = ~f_arrdiv24_fs215_or0;
  assign f_arrdiv24_fs216_xor0 = a[14] ^ b[0];
  assign f_arrdiv24_fs216_not0 = ~a[14];
  assign f_arrdiv24_fs216_and0 = f_arrdiv24_fs216_not0 & b[0];
  assign f_arrdiv24_fs216_not1 = ~f_arrdiv24_fs216_xor0;
  assign f_arrdiv24_fs217_xor0 = f_arrdiv24_mux2to1184_xor0 ^ b[1];
  assign f_arrdiv24_fs217_not0 = ~f_arrdiv24_mux2to1184_xor0;
  assign f_arrdiv24_fs217_and0 = f_arrdiv24_fs217_not0 & b[1];
  assign f_arrdiv24_fs217_xor1 = f_arrdiv24_fs216_and0 ^ f_arrdiv24_fs217_xor0;
  assign f_arrdiv24_fs217_not1 = ~f_arrdiv24_fs217_xor0;
  assign f_arrdiv24_fs217_and1 = f_arrdiv24_fs217_not1 & f_arrdiv24_fs216_and0;
  assign f_arrdiv24_fs217_or0 = f_arrdiv24_fs217_and1 | f_arrdiv24_fs217_and0;
  assign f_arrdiv24_fs218_xor0 = f_arrdiv24_mux2to1185_xor0 ^ b[2];
  assign f_arrdiv24_fs218_not0 = ~f_arrdiv24_mux2to1185_xor0;
  assign f_arrdiv24_fs218_and0 = f_arrdiv24_fs218_not0 & b[2];
  assign f_arrdiv24_fs218_xor1 = f_arrdiv24_fs217_or0 ^ f_arrdiv24_fs218_xor0;
  assign f_arrdiv24_fs218_not1 = ~f_arrdiv24_fs218_xor0;
  assign f_arrdiv24_fs218_and1 = f_arrdiv24_fs218_not1 & f_arrdiv24_fs217_or0;
  assign f_arrdiv24_fs218_or0 = f_arrdiv24_fs218_and1 | f_arrdiv24_fs218_and0;
  assign f_arrdiv24_fs219_xor0 = f_arrdiv24_mux2to1186_xor0 ^ b[3];
  assign f_arrdiv24_fs219_not0 = ~f_arrdiv24_mux2to1186_xor0;
  assign f_arrdiv24_fs219_and0 = f_arrdiv24_fs219_not0 & b[3];
  assign f_arrdiv24_fs219_xor1 = f_arrdiv24_fs218_or0 ^ f_arrdiv24_fs219_xor0;
  assign f_arrdiv24_fs219_not1 = ~f_arrdiv24_fs219_xor0;
  assign f_arrdiv24_fs219_and1 = f_arrdiv24_fs219_not1 & f_arrdiv24_fs218_or0;
  assign f_arrdiv24_fs219_or0 = f_arrdiv24_fs219_and1 | f_arrdiv24_fs219_and0;
  assign f_arrdiv24_fs220_xor0 = f_arrdiv24_mux2to1187_xor0 ^ b[4];
  assign f_arrdiv24_fs220_not0 = ~f_arrdiv24_mux2to1187_xor0;
  assign f_arrdiv24_fs220_and0 = f_arrdiv24_fs220_not0 & b[4];
  assign f_arrdiv24_fs220_xor1 = f_arrdiv24_fs219_or0 ^ f_arrdiv24_fs220_xor0;
  assign f_arrdiv24_fs220_not1 = ~f_arrdiv24_fs220_xor0;
  assign f_arrdiv24_fs220_and1 = f_arrdiv24_fs220_not1 & f_arrdiv24_fs219_or0;
  assign f_arrdiv24_fs220_or0 = f_arrdiv24_fs220_and1 | f_arrdiv24_fs220_and0;
  assign f_arrdiv24_fs221_xor0 = f_arrdiv24_mux2to1188_xor0 ^ b[5];
  assign f_arrdiv24_fs221_not0 = ~f_arrdiv24_mux2to1188_xor0;
  assign f_arrdiv24_fs221_and0 = f_arrdiv24_fs221_not0 & b[5];
  assign f_arrdiv24_fs221_xor1 = f_arrdiv24_fs220_or0 ^ f_arrdiv24_fs221_xor0;
  assign f_arrdiv24_fs221_not1 = ~f_arrdiv24_fs221_xor0;
  assign f_arrdiv24_fs221_and1 = f_arrdiv24_fs221_not1 & f_arrdiv24_fs220_or0;
  assign f_arrdiv24_fs221_or0 = f_arrdiv24_fs221_and1 | f_arrdiv24_fs221_and0;
  assign f_arrdiv24_fs222_xor0 = f_arrdiv24_mux2to1189_xor0 ^ b[6];
  assign f_arrdiv24_fs222_not0 = ~f_arrdiv24_mux2to1189_xor0;
  assign f_arrdiv24_fs222_and0 = f_arrdiv24_fs222_not0 & b[6];
  assign f_arrdiv24_fs222_xor1 = f_arrdiv24_fs221_or0 ^ f_arrdiv24_fs222_xor0;
  assign f_arrdiv24_fs222_not1 = ~f_arrdiv24_fs222_xor0;
  assign f_arrdiv24_fs222_and1 = f_arrdiv24_fs222_not1 & f_arrdiv24_fs221_or0;
  assign f_arrdiv24_fs222_or0 = f_arrdiv24_fs222_and1 | f_arrdiv24_fs222_and0;
  assign f_arrdiv24_fs223_xor0 = f_arrdiv24_mux2to1190_xor0 ^ b[7];
  assign f_arrdiv24_fs223_not0 = ~f_arrdiv24_mux2to1190_xor0;
  assign f_arrdiv24_fs223_and0 = f_arrdiv24_fs223_not0 & b[7];
  assign f_arrdiv24_fs223_xor1 = f_arrdiv24_fs222_or0 ^ f_arrdiv24_fs223_xor0;
  assign f_arrdiv24_fs223_not1 = ~f_arrdiv24_fs223_xor0;
  assign f_arrdiv24_fs223_and1 = f_arrdiv24_fs223_not1 & f_arrdiv24_fs222_or0;
  assign f_arrdiv24_fs223_or0 = f_arrdiv24_fs223_and1 | f_arrdiv24_fs223_and0;
  assign f_arrdiv24_fs224_xor0 = f_arrdiv24_mux2to1191_xor0 ^ b[8];
  assign f_arrdiv24_fs224_not0 = ~f_arrdiv24_mux2to1191_xor0;
  assign f_arrdiv24_fs224_and0 = f_arrdiv24_fs224_not0 & b[8];
  assign f_arrdiv24_fs224_xor1 = f_arrdiv24_fs223_or0 ^ f_arrdiv24_fs224_xor0;
  assign f_arrdiv24_fs224_not1 = ~f_arrdiv24_fs224_xor0;
  assign f_arrdiv24_fs224_and1 = f_arrdiv24_fs224_not1 & f_arrdiv24_fs223_or0;
  assign f_arrdiv24_fs224_or0 = f_arrdiv24_fs224_and1 | f_arrdiv24_fs224_and0;
  assign f_arrdiv24_fs225_xor0 = f_arrdiv24_mux2to1192_xor0 ^ b[9];
  assign f_arrdiv24_fs225_not0 = ~f_arrdiv24_mux2to1192_xor0;
  assign f_arrdiv24_fs225_and0 = f_arrdiv24_fs225_not0 & b[9];
  assign f_arrdiv24_fs225_xor1 = f_arrdiv24_fs224_or0 ^ f_arrdiv24_fs225_xor0;
  assign f_arrdiv24_fs225_not1 = ~f_arrdiv24_fs225_xor0;
  assign f_arrdiv24_fs225_and1 = f_arrdiv24_fs225_not1 & f_arrdiv24_fs224_or0;
  assign f_arrdiv24_fs225_or0 = f_arrdiv24_fs225_and1 | f_arrdiv24_fs225_and0;
  assign f_arrdiv24_fs226_xor0 = f_arrdiv24_mux2to1193_xor0 ^ b[10];
  assign f_arrdiv24_fs226_not0 = ~f_arrdiv24_mux2to1193_xor0;
  assign f_arrdiv24_fs226_and0 = f_arrdiv24_fs226_not0 & b[10];
  assign f_arrdiv24_fs226_xor1 = f_arrdiv24_fs225_or0 ^ f_arrdiv24_fs226_xor0;
  assign f_arrdiv24_fs226_not1 = ~f_arrdiv24_fs226_xor0;
  assign f_arrdiv24_fs226_and1 = f_arrdiv24_fs226_not1 & f_arrdiv24_fs225_or0;
  assign f_arrdiv24_fs226_or0 = f_arrdiv24_fs226_and1 | f_arrdiv24_fs226_and0;
  assign f_arrdiv24_fs227_xor0 = f_arrdiv24_mux2to1194_xor0 ^ b[11];
  assign f_arrdiv24_fs227_not0 = ~f_arrdiv24_mux2to1194_xor0;
  assign f_arrdiv24_fs227_and0 = f_arrdiv24_fs227_not0 & b[11];
  assign f_arrdiv24_fs227_xor1 = f_arrdiv24_fs226_or0 ^ f_arrdiv24_fs227_xor0;
  assign f_arrdiv24_fs227_not1 = ~f_arrdiv24_fs227_xor0;
  assign f_arrdiv24_fs227_and1 = f_arrdiv24_fs227_not1 & f_arrdiv24_fs226_or0;
  assign f_arrdiv24_fs227_or0 = f_arrdiv24_fs227_and1 | f_arrdiv24_fs227_and0;
  assign f_arrdiv24_fs228_xor0 = f_arrdiv24_mux2to1195_xor0 ^ b[12];
  assign f_arrdiv24_fs228_not0 = ~f_arrdiv24_mux2to1195_xor0;
  assign f_arrdiv24_fs228_and0 = f_arrdiv24_fs228_not0 & b[12];
  assign f_arrdiv24_fs228_xor1 = f_arrdiv24_fs227_or0 ^ f_arrdiv24_fs228_xor0;
  assign f_arrdiv24_fs228_not1 = ~f_arrdiv24_fs228_xor0;
  assign f_arrdiv24_fs228_and1 = f_arrdiv24_fs228_not1 & f_arrdiv24_fs227_or0;
  assign f_arrdiv24_fs228_or0 = f_arrdiv24_fs228_and1 | f_arrdiv24_fs228_and0;
  assign f_arrdiv24_fs229_xor0 = f_arrdiv24_mux2to1196_xor0 ^ b[13];
  assign f_arrdiv24_fs229_not0 = ~f_arrdiv24_mux2to1196_xor0;
  assign f_arrdiv24_fs229_and0 = f_arrdiv24_fs229_not0 & b[13];
  assign f_arrdiv24_fs229_xor1 = f_arrdiv24_fs228_or0 ^ f_arrdiv24_fs229_xor0;
  assign f_arrdiv24_fs229_not1 = ~f_arrdiv24_fs229_xor0;
  assign f_arrdiv24_fs229_and1 = f_arrdiv24_fs229_not1 & f_arrdiv24_fs228_or0;
  assign f_arrdiv24_fs229_or0 = f_arrdiv24_fs229_and1 | f_arrdiv24_fs229_and0;
  assign f_arrdiv24_fs230_xor0 = f_arrdiv24_mux2to1197_xor0 ^ b[14];
  assign f_arrdiv24_fs230_not0 = ~f_arrdiv24_mux2to1197_xor0;
  assign f_arrdiv24_fs230_and0 = f_arrdiv24_fs230_not0 & b[14];
  assign f_arrdiv24_fs230_xor1 = f_arrdiv24_fs229_or0 ^ f_arrdiv24_fs230_xor0;
  assign f_arrdiv24_fs230_not1 = ~f_arrdiv24_fs230_xor0;
  assign f_arrdiv24_fs230_and1 = f_arrdiv24_fs230_not1 & f_arrdiv24_fs229_or0;
  assign f_arrdiv24_fs230_or0 = f_arrdiv24_fs230_and1 | f_arrdiv24_fs230_and0;
  assign f_arrdiv24_fs231_xor0 = f_arrdiv24_mux2to1198_xor0 ^ b[15];
  assign f_arrdiv24_fs231_not0 = ~f_arrdiv24_mux2to1198_xor0;
  assign f_arrdiv24_fs231_and0 = f_arrdiv24_fs231_not0 & b[15];
  assign f_arrdiv24_fs231_xor1 = f_arrdiv24_fs230_or0 ^ f_arrdiv24_fs231_xor0;
  assign f_arrdiv24_fs231_not1 = ~f_arrdiv24_fs231_xor0;
  assign f_arrdiv24_fs231_and1 = f_arrdiv24_fs231_not1 & f_arrdiv24_fs230_or0;
  assign f_arrdiv24_fs231_or0 = f_arrdiv24_fs231_and1 | f_arrdiv24_fs231_and0;
  assign f_arrdiv24_fs232_xor0 = f_arrdiv24_mux2to1199_xor0 ^ b[16];
  assign f_arrdiv24_fs232_not0 = ~f_arrdiv24_mux2to1199_xor0;
  assign f_arrdiv24_fs232_and0 = f_arrdiv24_fs232_not0 & b[16];
  assign f_arrdiv24_fs232_xor1 = f_arrdiv24_fs231_or0 ^ f_arrdiv24_fs232_xor0;
  assign f_arrdiv24_fs232_not1 = ~f_arrdiv24_fs232_xor0;
  assign f_arrdiv24_fs232_and1 = f_arrdiv24_fs232_not1 & f_arrdiv24_fs231_or0;
  assign f_arrdiv24_fs232_or0 = f_arrdiv24_fs232_and1 | f_arrdiv24_fs232_and0;
  assign f_arrdiv24_fs233_xor0 = f_arrdiv24_mux2to1200_xor0 ^ b[17];
  assign f_arrdiv24_fs233_not0 = ~f_arrdiv24_mux2to1200_xor0;
  assign f_arrdiv24_fs233_and0 = f_arrdiv24_fs233_not0 & b[17];
  assign f_arrdiv24_fs233_xor1 = f_arrdiv24_fs232_or0 ^ f_arrdiv24_fs233_xor0;
  assign f_arrdiv24_fs233_not1 = ~f_arrdiv24_fs233_xor0;
  assign f_arrdiv24_fs233_and1 = f_arrdiv24_fs233_not1 & f_arrdiv24_fs232_or0;
  assign f_arrdiv24_fs233_or0 = f_arrdiv24_fs233_and1 | f_arrdiv24_fs233_and0;
  assign f_arrdiv24_fs234_xor0 = f_arrdiv24_mux2to1201_xor0 ^ b[18];
  assign f_arrdiv24_fs234_not0 = ~f_arrdiv24_mux2to1201_xor0;
  assign f_arrdiv24_fs234_and0 = f_arrdiv24_fs234_not0 & b[18];
  assign f_arrdiv24_fs234_xor1 = f_arrdiv24_fs233_or0 ^ f_arrdiv24_fs234_xor0;
  assign f_arrdiv24_fs234_not1 = ~f_arrdiv24_fs234_xor0;
  assign f_arrdiv24_fs234_and1 = f_arrdiv24_fs234_not1 & f_arrdiv24_fs233_or0;
  assign f_arrdiv24_fs234_or0 = f_arrdiv24_fs234_and1 | f_arrdiv24_fs234_and0;
  assign f_arrdiv24_fs235_xor0 = f_arrdiv24_mux2to1202_xor0 ^ b[19];
  assign f_arrdiv24_fs235_not0 = ~f_arrdiv24_mux2to1202_xor0;
  assign f_arrdiv24_fs235_and0 = f_arrdiv24_fs235_not0 & b[19];
  assign f_arrdiv24_fs235_xor1 = f_arrdiv24_fs234_or0 ^ f_arrdiv24_fs235_xor0;
  assign f_arrdiv24_fs235_not1 = ~f_arrdiv24_fs235_xor0;
  assign f_arrdiv24_fs235_and1 = f_arrdiv24_fs235_not1 & f_arrdiv24_fs234_or0;
  assign f_arrdiv24_fs235_or0 = f_arrdiv24_fs235_and1 | f_arrdiv24_fs235_and0;
  assign f_arrdiv24_fs236_xor0 = f_arrdiv24_mux2to1203_xor0 ^ b[20];
  assign f_arrdiv24_fs236_not0 = ~f_arrdiv24_mux2to1203_xor0;
  assign f_arrdiv24_fs236_and0 = f_arrdiv24_fs236_not0 & b[20];
  assign f_arrdiv24_fs236_xor1 = f_arrdiv24_fs235_or0 ^ f_arrdiv24_fs236_xor0;
  assign f_arrdiv24_fs236_not1 = ~f_arrdiv24_fs236_xor0;
  assign f_arrdiv24_fs236_and1 = f_arrdiv24_fs236_not1 & f_arrdiv24_fs235_or0;
  assign f_arrdiv24_fs236_or0 = f_arrdiv24_fs236_and1 | f_arrdiv24_fs236_and0;
  assign f_arrdiv24_fs237_xor0 = f_arrdiv24_mux2to1204_xor0 ^ b[21];
  assign f_arrdiv24_fs237_not0 = ~f_arrdiv24_mux2to1204_xor0;
  assign f_arrdiv24_fs237_and0 = f_arrdiv24_fs237_not0 & b[21];
  assign f_arrdiv24_fs237_xor1 = f_arrdiv24_fs236_or0 ^ f_arrdiv24_fs237_xor0;
  assign f_arrdiv24_fs237_not1 = ~f_arrdiv24_fs237_xor0;
  assign f_arrdiv24_fs237_and1 = f_arrdiv24_fs237_not1 & f_arrdiv24_fs236_or0;
  assign f_arrdiv24_fs237_or0 = f_arrdiv24_fs237_and1 | f_arrdiv24_fs237_and0;
  assign f_arrdiv24_fs238_xor0 = f_arrdiv24_mux2to1205_xor0 ^ b[22];
  assign f_arrdiv24_fs238_not0 = ~f_arrdiv24_mux2to1205_xor0;
  assign f_arrdiv24_fs238_and0 = f_arrdiv24_fs238_not0 & b[22];
  assign f_arrdiv24_fs238_xor1 = f_arrdiv24_fs237_or0 ^ f_arrdiv24_fs238_xor0;
  assign f_arrdiv24_fs238_not1 = ~f_arrdiv24_fs238_xor0;
  assign f_arrdiv24_fs238_and1 = f_arrdiv24_fs238_not1 & f_arrdiv24_fs237_or0;
  assign f_arrdiv24_fs238_or0 = f_arrdiv24_fs238_and1 | f_arrdiv24_fs238_and0;
  assign f_arrdiv24_fs239_xor0 = f_arrdiv24_mux2to1206_xor0 ^ b[23];
  assign f_arrdiv24_fs239_not0 = ~f_arrdiv24_mux2to1206_xor0;
  assign f_arrdiv24_fs239_and0 = f_arrdiv24_fs239_not0 & b[23];
  assign f_arrdiv24_fs239_xor1 = f_arrdiv24_fs238_or0 ^ f_arrdiv24_fs239_xor0;
  assign f_arrdiv24_fs239_not1 = ~f_arrdiv24_fs239_xor0;
  assign f_arrdiv24_fs239_and1 = f_arrdiv24_fs239_not1 & f_arrdiv24_fs238_or0;
  assign f_arrdiv24_fs239_or0 = f_arrdiv24_fs239_and1 | f_arrdiv24_fs239_and0;
  assign f_arrdiv24_mux2to1207_and0 = a[14] & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1207_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1207_and1 = f_arrdiv24_fs216_xor0 & f_arrdiv24_mux2to1207_not0;
  assign f_arrdiv24_mux2to1207_xor0 = f_arrdiv24_mux2to1207_and0 ^ f_arrdiv24_mux2to1207_and1;
  assign f_arrdiv24_mux2to1208_and0 = f_arrdiv24_mux2to1184_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1208_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1208_and1 = f_arrdiv24_fs217_xor1 & f_arrdiv24_mux2to1208_not0;
  assign f_arrdiv24_mux2to1208_xor0 = f_arrdiv24_mux2to1208_and0 ^ f_arrdiv24_mux2to1208_and1;
  assign f_arrdiv24_mux2to1209_and0 = f_arrdiv24_mux2to1185_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1209_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1209_and1 = f_arrdiv24_fs218_xor1 & f_arrdiv24_mux2to1209_not0;
  assign f_arrdiv24_mux2to1209_xor0 = f_arrdiv24_mux2to1209_and0 ^ f_arrdiv24_mux2to1209_and1;
  assign f_arrdiv24_mux2to1210_and0 = f_arrdiv24_mux2to1186_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1210_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1210_and1 = f_arrdiv24_fs219_xor1 & f_arrdiv24_mux2to1210_not0;
  assign f_arrdiv24_mux2to1210_xor0 = f_arrdiv24_mux2to1210_and0 ^ f_arrdiv24_mux2to1210_and1;
  assign f_arrdiv24_mux2to1211_and0 = f_arrdiv24_mux2to1187_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1211_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1211_and1 = f_arrdiv24_fs220_xor1 & f_arrdiv24_mux2to1211_not0;
  assign f_arrdiv24_mux2to1211_xor0 = f_arrdiv24_mux2to1211_and0 ^ f_arrdiv24_mux2to1211_and1;
  assign f_arrdiv24_mux2to1212_and0 = f_arrdiv24_mux2to1188_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1212_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1212_and1 = f_arrdiv24_fs221_xor1 & f_arrdiv24_mux2to1212_not0;
  assign f_arrdiv24_mux2to1212_xor0 = f_arrdiv24_mux2to1212_and0 ^ f_arrdiv24_mux2to1212_and1;
  assign f_arrdiv24_mux2to1213_and0 = f_arrdiv24_mux2to1189_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1213_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1213_and1 = f_arrdiv24_fs222_xor1 & f_arrdiv24_mux2to1213_not0;
  assign f_arrdiv24_mux2to1213_xor0 = f_arrdiv24_mux2to1213_and0 ^ f_arrdiv24_mux2to1213_and1;
  assign f_arrdiv24_mux2to1214_and0 = f_arrdiv24_mux2to1190_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1214_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1214_and1 = f_arrdiv24_fs223_xor1 & f_arrdiv24_mux2to1214_not0;
  assign f_arrdiv24_mux2to1214_xor0 = f_arrdiv24_mux2to1214_and0 ^ f_arrdiv24_mux2to1214_and1;
  assign f_arrdiv24_mux2to1215_and0 = f_arrdiv24_mux2to1191_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1215_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1215_and1 = f_arrdiv24_fs224_xor1 & f_arrdiv24_mux2to1215_not0;
  assign f_arrdiv24_mux2to1215_xor0 = f_arrdiv24_mux2to1215_and0 ^ f_arrdiv24_mux2to1215_and1;
  assign f_arrdiv24_mux2to1216_and0 = f_arrdiv24_mux2to1192_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1216_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1216_and1 = f_arrdiv24_fs225_xor1 & f_arrdiv24_mux2to1216_not0;
  assign f_arrdiv24_mux2to1216_xor0 = f_arrdiv24_mux2to1216_and0 ^ f_arrdiv24_mux2to1216_and1;
  assign f_arrdiv24_mux2to1217_and0 = f_arrdiv24_mux2to1193_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1217_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1217_and1 = f_arrdiv24_fs226_xor1 & f_arrdiv24_mux2to1217_not0;
  assign f_arrdiv24_mux2to1217_xor0 = f_arrdiv24_mux2to1217_and0 ^ f_arrdiv24_mux2to1217_and1;
  assign f_arrdiv24_mux2to1218_and0 = f_arrdiv24_mux2to1194_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1218_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1218_and1 = f_arrdiv24_fs227_xor1 & f_arrdiv24_mux2to1218_not0;
  assign f_arrdiv24_mux2to1218_xor0 = f_arrdiv24_mux2to1218_and0 ^ f_arrdiv24_mux2to1218_and1;
  assign f_arrdiv24_mux2to1219_and0 = f_arrdiv24_mux2to1195_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1219_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1219_and1 = f_arrdiv24_fs228_xor1 & f_arrdiv24_mux2to1219_not0;
  assign f_arrdiv24_mux2to1219_xor0 = f_arrdiv24_mux2to1219_and0 ^ f_arrdiv24_mux2to1219_and1;
  assign f_arrdiv24_mux2to1220_and0 = f_arrdiv24_mux2to1196_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1220_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1220_and1 = f_arrdiv24_fs229_xor1 & f_arrdiv24_mux2to1220_not0;
  assign f_arrdiv24_mux2to1220_xor0 = f_arrdiv24_mux2to1220_and0 ^ f_arrdiv24_mux2to1220_and1;
  assign f_arrdiv24_mux2to1221_and0 = f_arrdiv24_mux2to1197_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1221_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1221_and1 = f_arrdiv24_fs230_xor1 & f_arrdiv24_mux2to1221_not0;
  assign f_arrdiv24_mux2to1221_xor0 = f_arrdiv24_mux2to1221_and0 ^ f_arrdiv24_mux2to1221_and1;
  assign f_arrdiv24_mux2to1222_and0 = f_arrdiv24_mux2to1198_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1222_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1222_and1 = f_arrdiv24_fs231_xor1 & f_arrdiv24_mux2to1222_not0;
  assign f_arrdiv24_mux2to1222_xor0 = f_arrdiv24_mux2to1222_and0 ^ f_arrdiv24_mux2to1222_and1;
  assign f_arrdiv24_mux2to1223_and0 = f_arrdiv24_mux2to1199_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1223_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1223_and1 = f_arrdiv24_fs232_xor1 & f_arrdiv24_mux2to1223_not0;
  assign f_arrdiv24_mux2to1223_xor0 = f_arrdiv24_mux2to1223_and0 ^ f_arrdiv24_mux2to1223_and1;
  assign f_arrdiv24_mux2to1224_and0 = f_arrdiv24_mux2to1200_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1224_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1224_and1 = f_arrdiv24_fs233_xor1 & f_arrdiv24_mux2to1224_not0;
  assign f_arrdiv24_mux2to1224_xor0 = f_arrdiv24_mux2to1224_and0 ^ f_arrdiv24_mux2to1224_and1;
  assign f_arrdiv24_mux2to1225_and0 = f_arrdiv24_mux2to1201_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1225_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1225_and1 = f_arrdiv24_fs234_xor1 & f_arrdiv24_mux2to1225_not0;
  assign f_arrdiv24_mux2to1225_xor0 = f_arrdiv24_mux2to1225_and0 ^ f_arrdiv24_mux2to1225_and1;
  assign f_arrdiv24_mux2to1226_and0 = f_arrdiv24_mux2to1202_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1226_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1226_and1 = f_arrdiv24_fs235_xor1 & f_arrdiv24_mux2to1226_not0;
  assign f_arrdiv24_mux2to1226_xor0 = f_arrdiv24_mux2to1226_and0 ^ f_arrdiv24_mux2to1226_and1;
  assign f_arrdiv24_mux2to1227_and0 = f_arrdiv24_mux2to1203_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1227_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1227_and1 = f_arrdiv24_fs236_xor1 & f_arrdiv24_mux2to1227_not0;
  assign f_arrdiv24_mux2to1227_xor0 = f_arrdiv24_mux2to1227_and0 ^ f_arrdiv24_mux2to1227_and1;
  assign f_arrdiv24_mux2to1228_and0 = f_arrdiv24_mux2to1204_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1228_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1228_and1 = f_arrdiv24_fs237_xor1 & f_arrdiv24_mux2to1228_not0;
  assign f_arrdiv24_mux2to1228_xor0 = f_arrdiv24_mux2to1228_and0 ^ f_arrdiv24_mux2to1228_and1;
  assign f_arrdiv24_mux2to1229_and0 = f_arrdiv24_mux2to1205_xor0 & f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1229_not0 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_mux2to1229_and1 = f_arrdiv24_fs238_xor1 & f_arrdiv24_mux2to1229_not0;
  assign f_arrdiv24_mux2to1229_xor0 = f_arrdiv24_mux2to1229_and0 ^ f_arrdiv24_mux2to1229_and1;
  assign f_arrdiv24_not9 = ~f_arrdiv24_fs239_or0;
  assign f_arrdiv24_fs240_xor0 = a[13] ^ b[0];
  assign f_arrdiv24_fs240_not0 = ~a[13];
  assign f_arrdiv24_fs240_and0 = f_arrdiv24_fs240_not0 & b[0];
  assign f_arrdiv24_fs240_not1 = ~f_arrdiv24_fs240_xor0;
  assign f_arrdiv24_fs241_xor0 = f_arrdiv24_mux2to1207_xor0 ^ b[1];
  assign f_arrdiv24_fs241_not0 = ~f_arrdiv24_mux2to1207_xor0;
  assign f_arrdiv24_fs241_and0 = f_arrdiv24_fs241_not0 & b[1];
  assign f_arrdiv24_fs241_xor1 = f_arrdiv24_fs240_and0 ^ f_arrdiv24_fs241_xor0;
  assign f_arrdiv24_fs241_not1 = ~f_arrdiv24_fs241_xor0;
  assign f_arrdiv24_fs241_and1 = f_arrdiv24_fs241_not1 & f_arrdiv24_fs240_and0;
  assign f_arrdiv24_fs241_or0 = f_arrdiv24_fs241_and1 | f_arrdiv24_fs241_and0;
  assign f_arrdiv24_fs242_xor0 = f_arrdiv24_mux2to1208_xor0 ^ b[2];
  assign f_arrdiv24_fs242_not0 = ~f_arrdiv24_mux2to1208_xor0;
  assign f_arrdiv24_fs242_and0 = f_arrdiv24_fs242_not0 & b[2];
  assign f_arrdiv24_fs242_xor1 = f_arrdiv24_fs241_or0 ^ f_arrdiv24_fs242_xor0;
  assign f_arrdiv24_fs242_not1 = ~f_arrdiv24_fs242_xor0;
  assign f_arrdiv24_fs242_and1 = f_arrdiv24_fs242_not1 & f_arrdiv24_fs241_or0;
  assign f_arrdiv24_fs242_or0 = f_arrdiv24_fs242_and1 | f_arrdiv24_fs242_and0;
  assign f_arrdiv24_fs243_xor0 = f_arrdiv24_mux2to1209_xor0 ^ b[3];
  assign f_arrdiv24_fs243_not0 = ~f_arrdiv24_mux2to1209_xor0;
  assign f_arrdiv24_fs243_and0 = f_arrdiv24_fs243_not0 & b[3];
  assign f_arrdiv24_fs243_xor1 = f_arrdiv24_fs242_or0 ^ f_arrdiv24_fs243_xor0;
  assign f_arrdiv24_fs243_not1 = ~f_arrdiv24_fs243_xor0;
  assign f_arrdiv24_fs243_and1 = f_arrdiv24_fs243_not1 & f_arrdiv24_fs242_or0;
  assign f_arrdiv24_fs243_or0 = f_arrdiv24_fs243_and1 | f_arrdiv24_fs243_and0;
  assign f_arrdiv24_fs244_xor0 = f_arrdiv24_mux2to1210_xor0 ^ b[4];
  assign f_arrdiv24_fs244_not0 = ~f_arrdiv24_mux2to1210_xor0;
  assign f_arrdiv24_fs244_and0 = f_arrdiv24_fs244_not0 & b[4];
  assign f_arrdiv24_fs244_xor1 = f_arrdiv24_fs243_or0 ^ f_arrdiv24_fs244_xor0;
  assign f_arrdiv24_fs244_not1 = ~f_arrdiv24_fs244_xor0;
  assign f_arrdiv24_fs244_and1 = f_arrdiv24_fs244_not1 & f_arrdiv24_fs243_or0;
  assign f_arrdiv24_fs244_or0 = f_arrdiv24_fs244_and1 | f_arrdiv24_fs244_and0;
  assign f_arrdiv24_fs245_xor0 = f_arrdiv24_mux2to1211_xor0 ^ b[5];
  assign f_arrdiv24_fs245_not0 = ~f_arrdiv24_mux2to1211_xor0;
  assign f_arrdiv24_fs245_and0 = f_arrdiv24_fs245_not0 & b[5];
  assign f_arrdiv24_fs245_xor1 = f_arrdiv24_fs244_or0 ^ f_arrdiv24_fs245_xor0;
  assign f_arrdiv24_fs245_not1 = ~f_arrdiv24_fs245_xor0;
  assign f_arrdiv24_fs245_and1 = f_arrdiv24_fs245_not1 & f_arrdiv24_fs244_or0;
  assign f_arrdiv24_fs245_or0 = f_arrdiv24_fs245_and1 | f_arrdiv24_fs245_and0;
  assign f_arrdiv24_fs246_xor0 = f_arrdiv24_mux2to1212_xor0 ^ b[6];
  assign f_arrdiv24_fs246_not0 = ~f_arrdiv24_mux2to1212_xor0;
  assign f_arrdiv24_fs246_and0 = f_arrdiv24_fs246_not0 & b[6];
  assign f_arrdiv24_fs246_xor1 = f_arrdiv24_fs245_or0 ^ f_arrdiv24_fs246_xor0;
  assign f_arrdiv24_fs246_not1 = ~f_arrdiv24_fs246_xor0;
  assign f_arrdiv24_fs246_and1 = f_arrdiv24_fs246_not1 & f_arrdiv24_fs245_or0;
  assign f_arrdiv24_fs246_or0 = f_arrdiv24_fs246_and1 | f_arrdiv24_fs246_and0;
  assign f_arrdiv24_fs247_xor0 = f_arrdiv24_mux2to1213_xor0 ^ b[7];
  assign f_arrdiv24_fs247_not0 = ~f_arrdiv24_mux2to1213_xor0;
  assign f_arrdiv24_fs247_and0 = f_arrdiv24_fs247_not0 & b[7];
  assign f_arrdiv24_fs247_xor1 = f_arrdiv24_fs246_or0 ^ f_arrdiv24_fs247_xor0;
  assign f_arrdiv24_fs247_not1 = ~f_arrdiv24_fs247_xor0;
  assign f_arrdiv24_fs247_and1 = f_arrdiv24_fs247_not1 & f_arrdiv24_fs246_or0;
  assign f_arrdiv24_fs247_or0 = f_arrdiv24_fs247_and1 | f_arrdiv24_fs247_and0;
  assign f_arrdiv24_fs248_xor0 = f_arrdiv24_mux2to1214_xor0 ^ b[8];
  assign f_arrdiv24_fs248_not0 = ~f_arrdiv24_mux2to1214_xor0;
  assign f_arrdiv24_fs248_and0 = f_arrdiv24_fs248_not0 & b[8];
  assign f_arrdiv24_fs248_xor1 = f_arrdiv24_fs247_or0 ^ f_arrdiv24_fs248_xor0;
  assign f_arrdiv24_fs248_not1 = ~f_arrdiv24_fs248_xor0;
  assign f_arrdiv24_fs248_and1 = f_arrdiv24_fs248_not1 & f_arrdiv24_fs247_or0;
  assign f_arrdiv24_fs248_or0 = f_arrdiv24_fs248_and1 | f_arrdiv24_fs248_and0;
  assign f_arrdiv24_fs249_xor0 = f_arrdiv24_mux2to1215_xor0 ^ b[9];
  assign f_arrdiv24_fs249_not0 = ~f_arrdiv24_mux2to1215_xor0;
  assign f_arrdiv24_fs249_and0 = f_arrdiv24_fs249_not0 & b[9];
  assign f_arrdiv24_fs249_xor1 = f_arrdiv24_fs248_or0 ^ f_arrdiv24_fs249_xor0;
  assign f_arrdiv24_fs249_not1 = ~f_arrdiv24_fs249_xor0;
  assign f_arrdiv24_fs249_and1 = f_arrdiv24_fs249_not1 & f_arrdiv24_fs248_or0;
  assign f_arrdiv24_fs249_or0 = f_arrdiv24_fs249_and1 | f_arrdiv24_fs249_and0;
  assign f_arrdiv24_fs250_xor0 = f_arrdiv24_mux2to1216_xor0 ^ b[10];
  assign f_arrdiv24_fs250_not0 = ~f_arrdiv24_mux2to1216_xor0;
  assign f_arrdiv24_fs250_and0 = f_arrdiv24_fs250_not0 & b[10];
  assign f_arrdiv24_fs250_xor1 = f_arrdiv24_fs249_or0 ^ f_arrdiv24_fs250_xor0;
  assign f_arrdiv24_fs250_not1 = ~f_arrdiv24_fs250_xor0;
  assign f_arrdiv24_fs250_and1 = f_arrdiv24_fs250_not1 & f_arrdiv24_fs249_or0;
  assign f_arrdiv24_fs250_or0 = f_arrdiv24_fs250_and1 | f_arrdiv24_fs250_and0;
  assign f_arrdiv24_fs251_xor0 = f_arrdiv24_mux2to1217_xor0 ^ b[11];
  assign f_arrdiv24_fs251_not0 = ~f_arrdiv24_mux2to1217_xor0;
  assign f_arrdiv24_fs251_and0 = f_arrdiv24_fs251_not0 & b[11];
  assign f_arrdiv24_fs251_xor1 = f_arrdiv24_fs250_or0 ^ f_arrdiv24_fs251_xor0;
  assign f_arrdiv24_fs251_not1 = ~f_arrdiv24_fs251_xor0;
  assign f_arrdiv24_fs251_and1 = f_arrdiv24_fs251_not1 & f_arrdiv24_fs250_or0;
  assign f_arrdiv24_fs251_or0 = f_arrdiv24_fs251_and1 | f_arrdiv24_fs251_and0;
  assign f_arrdiv24_fs252_xor0 = f_arrdiv24_mux2to1218_xor0 ^ b[12];
  assign f_arrdiv24_fs252_not0 = ~f_arrdiv24_mux2to1218_xor0;
  assign f_arrdiv24_fs252_and0 = f_arrdiv24_fs252_not0 & b[12];
  assign f_arrdiv24_fs252_xor1 = f_arrdiv24_fs251_or0 ^ f_arrdiv24_fs252_xor0;
  assign f_arrdiv24_fs252_not1 = ~f_arrdiv24_fs252_xor0;
  assign f_arrdiv24_fs252_and1 = f_arrdiv24_fs252_not1 & f_arrdiv24_fs251_or0;
  assign f_arrdiv24_fs252_or0 = f_arrdiv24_fs252_and1 | f_arrdiv24_fs252_and0;
  assign f_arrdiv24_fs253_xor0 = f_arrdiv24_mux2to1219_xor0 ^ b[13];
  assign f_arrdiv24_fs253_not0 = ~f_arrdiv24_mux2to1219_xor0;
  assign f_arrdiv24_fs253_and0 = f_arrdiv24_fs253_not0 & b[13];
  assign f_arrdiv24_fs253_xor1 = f_arrdiv24_fs252_or0 ^ f_arrdiv24_fs253_xor0;
  assign f_arrdiv24_fs253_not1 = ~f_arrdiv24_fs253_xor0;
  assign f_arrdiv24_fs253_and1 = f_arrdiv24_fs253_not1 & f_arrdiv24_fs252_or0;
  assign f_arrdiv24_fs253_or0 = f_arrdiv24_fs253_and1 | f_arrdiv24_fs253_and0;
  assign f_arrdiv24_fs254_xor0 = f_arrdiv24_mux2to1220_xor0 ^ b[14];
  assign f_arrdiv24_fs254_not0 = ~f_arrdiv24_mux2to1220_xor0;
  assign f_arrdiv24_fs254_and0 = f_arrdiv24_fs254_not0 & b[14];
  assign f_arrdiv24_fs254_xor1 = f_arrdiv24_fs253_or0 ^ f_arrdiv24_fs254_xor0;
  assign f_arrdiv24_fs254_not1 = ~f_arrdiv24_fs254_xor0;
  assign f_arrdiv24_fs254_and1 = f_arrdiv24_fs254_not1 & f_arrdiv24_fs253_or0;
  assign f_arrdiv24_fs254_or0 = f_arrdiv24_fs254_and1 | f_arrdiv24_fs254_and0;
  assign f_arrdiv24_fs255_xor0 = f_arrdiv24_mux2to1221_xor0 ^ b[15];
  assign f_arrdiv24_fs255_not0 = ~f_arrdiv24_mux2to1221_xor0;
  assign f_arrdiv24_fs255_and0 = f_arrdiv24_fs255_not0 & b[15];
  assign f_arrdiv24_fs255_xor1 = f_arrdiv24_fs254_or0 ^ f_arrdiv24_fs255_xor0;
  assign f_arrdiv24_fs255_not1 = ~f_arrdiv24_fs255_xor0;
  assign f_arrdiv24_fs255_and1 = f_arrdiv24_fs255_not1 & f_arrdiv24_fs254_or0;
  assign f_arrdiv24_fs255_or0 = f_arrdiv24_fs255_and1 | f_arrdiv24_fs255_and0;
  assign f_arrdiv24_fs256_xor0 = f_arrdiv24_mux2to1222_xor0 ^ b[16];
  assign f_arrdiv24_fs256_not0 = ~f_arrdiv24_mux2to1222_xor0;
  assign f_arrdiv24_fs256_and0 = f_arrdiv24_fs256_not0 & b[16];
  assign f_arrdiv24_fs256_xor1 = f_arrdiv24_fs255_or0 ^ f_arrdiv24_fs256_xor0;
  assign f_arrdiv24_fs256_not1 = ~f_arrdiv24_fs256_xor0;
  assign f_arrdiv24_fs256_and1 = f_arrdiv24_fs256_not1 & f_arrdiv24_fs255_or0;
  assign f_arrdiv24_fs256_or0 = f_arrdiv24_fs256_and1 | f_arrdiv24_fs256_and0;
  assign f_arrdiv24_fs257_xor0 = f_arrdiv24_mux2to1223_xor0 ^ b[17];
  assign f_arrdiv24_fs257_not0 = ~f_arrdiv24_mux2to1223_xor0;
  assign f_arrdiv24_fs257_and0 = f_arrdiv24_fs257_not0 & b[17];
  assign f_arrdiv24_fs257_xor1 = f_arrdiv24_fs256_or0 ^ f_arrdiv24_fs257_xor0;
  assign f_arrdiv24_fs257_not1 = ~f_arrdiv24_fs257_xor0;
  assign f_arrdiv24_fs257_and1 = f_arrdiv24_fs257_not1 & f_arrdiv24_fs256_or0;
  assign f_arrdiv24_fs257_or0 = f_arrdiv24_fs257_and1 | f_arrdiv24_fs257_and0;
  assign f_arrdiv24_fs258_xor0 = f_arrdiv24_mux2to1224_xor0 ^ b[18];
  assign f_arrdiv24_fs258_not0 = ~f_arrdiv24_mux2to1224_xor0;
  assign f_arrdiv24_fs258_and0 = f_arrdiv24_fs258_not0 & b[18];
  assign f_arrdiv24_fs258_xor1 = f_arrdiv24_fs257_or0 ^ f_arrdiv24_fs258_xor0;
  assign f_arrdiv24_fs258_not1 = ~f_arrdiv24_fs258_xor0;
  assign f_arrdiv24_fs258_and1 = f_arrdiv24_fs258_not1 & f_arrdiv24_fs257_or0;
  assign f_arrdiv24_fs258_or0 = f_arrdiv24_fs258_and1 | f_arrdiv24_fs258_and0;
  assign f_arrdiv24_fs259_xor0 = f_arrdiv24_mux2to1225_xor0 ^ b[19];
  assign f_arrdiv24_fs259_not0 = ~f_arrdiv24_mux2to1225_xor0;
  assign f_arrdiv24_fs259_and0 = f_arrdiv24_fs259_not0 & b[19];
  assign f_arrdiv24_fs259_xor1 = f_arrdiv24_fs258_or0 ^ f_arrdiv24_fs259_xor0;
  assign f_arrdiv24_fs259_not1 = ~f_arrdiv24_fs259_xor0;
  assign f_arrdiv24_fs259_and1 = f_arrdiv24_fs259_not1 & f_arrdiv24_fs258_or0;
  assign f_arrdiv24_fs259_or0 = f_arrdiv24_fs259_and1 | f_arrdiv24_fs259_and0;
  assign f_arrdiv24_fs260_xor0 = f_arrdiv24_mux2to1226_xor0 ^ b[20];
  assign f_arrdiv24_fs260_not0 = ~f_arrdiv24_mux2to1226_xor0;
  assign f_arrdiv24_fs260_and0 = f_arrdiv24_fs260_not0 & b[20];
  assign f_arrdiv24_fs260_xor1 = f_arrdiv24_fs259_or0 ^ f_arrdiv24_fs260_xor0;
  assign f_arrdiv24_fs260_not1 = ~f_arrdiv24_fs260_xor0;
  assign f_arrdiv24_fs260_and1 = f_arrdiv24_fs260_not1 & f_arrdiv24_fs259_or0;
  assign f_arrdiv24_fs260_or0 = f_arrdiv24_fs260_and1 | f_arrdiv24_fs260_and0;
  assign f_arrdiv24_fs261_xor0 = f_arrdiv24_mux2to1227_xor0 ^ b[21];
  assign f_arrdiv24_fs261_not0 = ~f_arrdiv24_mux2to1227_xor0;
  assign f_arrdiv24_fs261_and0 = f_arrdiv24_fs261_not0 & b[21];
  assign f_arrdiv24_fs261_xor1 = f_arrdiv24_fs260_or0 ^ f_arrdiv24_fs261_xor0;
  assign f_arrdiv24_fs261_not1 = ~f_arrdiv24_fs261_xor0;
  assign f_arrdiv24_fs261_and1 = f_arrdiv24_fs261_not1 & f_arrdiv24_fs260_or0;
  assign f_arrdiv24_fs261_or0 = f_arrdiv24_fs261_and1 | f_arrdiv24_fs261_and0;
  assign f_arrdiv24_fs262_xor0 = f_arrdiv24_mux2to1228_xor0 ^ b[22];
  assign f_arrdiv24_fs262_not0 = ~f_arrdiv24_mux2to1228_xor0;
  assign f_arrdiv24_fs262_and0 = f_arrdiv24_fs262_not0 & b[22];
  assign f_arrdiv24_fs262_xor1 = f_arrdiv24_fs261_or0 ^ f_arrdiv24_fs262_xor0;
  assign f_arrdiv24_fs262_not1 = ~f_arrdiv24_fs262_xor0;
  assign f_arrdiv24_fs262_and1 = f_arrdiv24_fs262_not1 & f_arrdiv24_fs261_or0;
  assign f_arrdiv24_fs262_or0 = f_arrdiv24_fs262_and1 | f_arrdiv24_fs262_and0;
  assign f_arrdiv24_fs263_xor0 = f_arrdiv24_mux2to1229_xor0 ^ b[23];
  assign f_arrdiv24_fs263_not0 = ~f_arrdiv24_mux2to1229_xor0;
  assign f_arrdiv24_fs263_and0 = f_arrdiv24_fs263_not0 & b[23];
  assign f_arrdiv24_fs263_xor1 = f_arrdiv24_fs262_or0 ^ f_arrdiv24_fs263_xor0;
  assign f_arrdiv24_fs263_not1 = ~f_arrdiv24_fs263_xor0;
  assign f_arrdiv24_fs263_and1 = f_arrdiv24_fs263_not1 & f_arrdiv24_fs262_or0;
  assign f_arrdiv24_fs263_or0 = f_arrdiv24_fs263_and1 | f_arrdiv24_fs263_and0;
  assign f_arrdiv24_mux2to1230_and0 = a[13] & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1230_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1230_and1 = f_arrdiv24_fs240_xor0 & f_arrdiv24_mux2to1230_not0;
  assign f_arrdiv24_mux2to1230_xor0 = f_arrdiv24_mux2to1230_and0 ^ f_arrdiv24_mux2to1230_and1;
  assign f_arrdiv24_mux2to1231_and0 = f_arrdiv24_mux2to1207_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1231_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1231_and1 = f_arrdiv24_fs241_xor1 & f_arrdiv24_mux2to1231_not0;
  assign f_arrdiv24_mux2to1231_xor0 = f_arrdiv24_mux2to1231_and0 ^ f_arrdiv24_mux2to1231_and1;
  assign f_arrdiv24_mux2to1232_and0 = f_arrdiv24_mux2to1208_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1232_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1232_and1 = f_arrdiv24_fs242_xor1 & f_arrdiv24_mux2to1232_not0;
  assign f_arrdiv24_mux2to1232_xor0 = f_arrdiv24_mux2to1232_and0 ^ f_arrdiv24_mux2to1232_and1;
  assign f_arrdiv24_mux2to1233_and0 = f_arrdiv24_mux2to1209_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1233_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1233_and1 = f_arrdiv24_fs243_xor1 & f_arrdiv24_mux2to1233_not0;
  assign f_arrdiv24_mux2to1233_xor0 = f_arrdiv24_mux2to1233_and0 ^ f_arrdiv24_mux2to1233_and1;
  assign f_arrdiv24_mux2to1234_and0 = f_arrdiv24_mux2to1210_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1234_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1234_and1 = f_arrdiv24_fs244_xor1 & f_arrdiv24_mux2to1234_not0;
  assign f_arrdiv24_mux2to1234_xor0 = f_arrdiv24_mux2to1234_and0 ^ f_arrdiv24_mux2to1234_and1;
  assign f_arrdiv24_mux2to1235_and0 = f_arrdiv24_mux2to1211_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1235_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1235_and1 = f_arrdiv24_fs245_xor1 & f_arrdiv24_mux2to1235_not0;
  assign f_arrdiv24_mux2to1235_xor0 = f_arrdiv24_mux2to1235_and0 ^ f_arrdiv24_mux2to1235_and1;
  assign f_arrdiv24_mux2to1236_and0 = f_arrdiv24_mux2to1212_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1236_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1236_and1 = f_arrdiv24_fs246_xor1 & f_arrdiv24_mux2to1236_not0;
  assign f_arrdiv24_mux2to1236_xor0 = f_arrdiv24_mux2to1236_and0 ^ f_arrdiv24_mux2to1236_and1;
  assign f_arrdiv24_mux2to1237_and0 = f_arrdiv24_mux2to1213_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1237_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1237_and1 = f_arrdiv24_fs247_xor1 & f_arrdiv24_mux2to1237_not0;
  assign f_arrdiv24_mux2to1237_xor0 = f_arrdiv24_mux2to1237_and0 ^ f_arrdiv24_mux2to1237_and1;
  assign f_arrdiv24_mux2to1238_and0 = f_arrdiv24_mux2to1214_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1238_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1238_and1 = f_arrdiv24_fs248_xor1 & f_arrdiv24_mux2to1238_not0;
  assign f_arrdiv24_mux2to1238_xor0 = f_arrdiv24_mux2to1238_and0 ^ f_arrdiv24_mux2to1238_and1;
  assign f_arrdiv24_mux2to1239_and0 = f_arrdiv24_mux2to1215_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1239_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1239_and1 = f_arrdiv24_fs249_xor1 & f_arrdiv24_mux2to1239_not0;
  assign f_arrdiv24_mux2to1239_xor0 = f_arrdiv24_mux2to1239_and0 ^ f_arrdiv24_mux2to1239_and1;
  assign f_arrdiv24_mux2to1240_and0 = f_arrdiv24_mux2to1216_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1240_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1240_and1 = f_arrdiv24_fs250_xor1 & f_arrdiv24_mux2to1240_not0;
  assign f_arrdiv24_mux2to1240_xor0 = f_arrdiv24_mux2to1240_and0 ^ f_arrdiv24_mux2to1240_and1;
  assign f_arrdiv24_mux2to1241_and0 = f_arrdiv24_mux2to1217_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1241_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1241_and1 = f_arrdiv24_fs251_xor1 & f_arrdiv24_mux2to1241_not0;
  assign f_arrdiv24_mux2to1241_xor0 = f_arrdiv24_mux2to1241_and0 ^ f_arrdiv24_mux2to1241_and1;
  assign f_arrdiv24_mux2to1242_and0 = f_arrdiv24_mux2to1218_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1242_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1242_and1 = f_arrdiv24_fs252_xor1 & f_arrdiv24_mux2to1242_not0;
  assign f_arrdiv24_mux2to1242_xor0 = f_arrdiv24_mux2to1242_and0 ^ f_arrdiv24_mux2to1242_and1;
  assign f_arrdiv24_mux2to1243_and0 = f_arrdiv24_mux2to1219_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1243_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1243_and1 = f_arrdiv24_fs253_xor1 & f_arrdiv24_mux2to1243_not0;
  assign f_arrdiv24_mux2to1243_xor0 = f_arrdiv24_mux2to1243_and0 ^ f_arrdiv24_mux2to1243_and1;
  assign f_arrdiv24_mux2to1244_and0 = f_arrdiv24_mux2to1220_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1244_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1244_and1 = f_arrdiv24_fs254_xor1 & f_arrdiv24_mux2to1244_not0;
  assign f_arrdiv24_mux2to1244_xor0 = f_arrdiv24_mux2to1244_and0 ^ f_arrdiv24_mux2to1244_and1;
  assign f_arrdiv24_mux2to1245_and0 = f_arrdiv24_mux2to1221_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1245_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1245_and1 = f_arrdiv24_fs255_xor1 & f_arrdiv24_mux2to1245_not0;
  assign f_arrdiv24_mux2to1245_xor0 = f_arrdiv24_mux2to1245_and0 ^ f_arrdiv24_mux2to1245_and1;
  assign f_arrdiv24_mux2to1246_and0 = f_arrdiv24_mux2to1222_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1246_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1246_and1 = f_arrdiv24_fs256_xor1 & f_arrdiv24_mux2to1246_not0;
  assign f_arrdiv24_mux2to1246_xor0 = f_arrdiv24_mux2to1246_and0 ^ f_arrdiv24_mux2to1246_and1;
  assign f_arrdiv24_mux2to1247_and0 = f_arrdiv24_mux2to1223_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1247_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1247_and1 = f_arrdiv24_fs257_xor1 & f_arrdiv24_mux2to1247_not0;
  assign f_arrdiv24_mux2to1247_xor0 = f_arrdiv24_mux2to1247_and0 ^ f_arrdiv24_mux2to1247_and1;
  assign f_arrdiv24_mux2to1248_and0 = f_arrdiv24_mux2to1224_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1248_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1248_and1 = f_arrdiv24_fs258_xor1 & f_arrdiv24_mux2to1248_not0;
  assign f_arrdiv24_mux2to1248_xor0 = f_arrdiv24_mux2to1248_and0 ^ f_arrdiv24_mux2to1248_and1;
  assign f_arrdiv24_mux2to1249_and0 = f_arrdiv24_mux2to1225_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1249_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1249_and1 = f_arrdiv24_fs259_xor1 & f_arrdiv24_mux2to1249_not0;
  assign f_arrdiv24_mux2to1249_xor0 = f_arrdiv24_mux2to1249_and0 ^ f_arrdiv24_mux2to1249_and1;
  assign f_arrdiv24_mux2to1250_and0 = f_arrdiv24_mux2to1226_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1250_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1250_and1 = f_arrdiv24_fs260_xor1 & f_arrdiv24_mux2to1250_not0;
  assign f_arrdiv24_mux2to1250_xor0 = f_arrdiv24_mux2to1250_and0 ^ f_arrdiv24_mux2to1250_and1;
  assign f_arrdiv24_mux2to1251_and0 = f_arrdiv24_mux2to1227_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1251_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1251_and1 = f_arrdiv24_fs261_xor1 & f_arrdiv24_mux2to1251_not0;
  assign f_arrdiv24_mux2to1251_xor0 = f_arrdiv24_mux2to1251_and0 ^ f_arrdiv24_mux2to1251_and1;
  assign f_arrdiv24_mux2to1252_and0 = f_arrdiv24_mux2to1228_xor0 & f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1252_not0 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_mux2to1252_and1 = f_arrdiv24_fs262_xor1 & f_arrdiv24_mux2to1252_not0;
  assign f_arrdiv24_mux2to1252_xor0 = f_arrdiv24_mux2to1252_and0 ^ f_arrdiv24_mux2to1252_and1;
  assign f_arrdiv24_not10 = ~f_arrdiv24_fs263_or0;
  assign f_arrdiv24_fs264_xor0 = a[12] ^ b[0];
  assign f_arrdiv24_fs264_not0 = ~a[12];
  assign f_arrdiv24_fs264_and0 = f_arrdiv24_fs264_not0 & b[0];
  assign f_arrdiv24_fs264_not1 = ~f_arrdiv24_fs264_xor0;
  assign f_arrdiv24_fs265_xor0 = f_arrdiv24_mux2to1230_xor0 ^ b[1];
  assign f_arrdiv24_fs265_not0 = ~f_arrdiv24_mux2to1230_xor0;
  assign f_arrdiv24_fs265_and0 = f_arrdiv24_fs265_not0 & b[1];
  assign f_arrdiv24_fs265_xor1 = f_arrdiv24_fs264_and0 ^ f_arrdiv24_fs265_xor0;
  assign f_arrdiv24_fs265_not1 = ~f_arrdiv24_fs265_xor0;
  assign f_arrdiv24_fs265_and1 = f_arrdiv24_fs265_not1 & f_arrdiv24_fs264_and0;
  assign f_arrdiv24_fs265_or0 = f_arrdiv24_fs265_and1 | f_arrdiv24_fs265_and0;
  assign f_arrdiv24_fs266_xor0 = f_arrdiv24_mux2to1231_xor0 ^ b[2];
  assign f_arrdiv24_fs266_not0 = ~f_arrdiv24_mux2to1231_xor0;
  assign f_arrdiv24_fs266_and0 = f_arrdiv24_fs266_not0 & b[2];
  assign f_arrdiv24_fs266_xor1 = f_arrdiv24_fs265_or0 ^ f_arrdiv24_fs266_xor0;
  assign f_arrdiv24_fs266_not1 = ~f_arrdiv24_fs266_xor0;
  assign f_arrdiv24_fs266_and1 = f_arrdiv24_fs266_not1 & f_arrdiv24_fs265_or0;
  assign f_arrdiv24_fs266_or0 = f_arrdiv24_fs266_and1 | f_arrdiv24_fs266_and0;
  assign f_arrdiv24_fs267_xor0 = f_arrdiv24_mux2to1232_xor0 ^ b[3];
  assign f_arrdiv24_fs267_not0 = ~f_arrdiv24_mux2to1232_xor0;
  assign f_arrdiv24_fs267_and0 = f_arrdiv24_fs267_not0 & b[3];
  assign f_arrdiv24_fs267_xor1 = f_arrdiv24_fs266_or0 ^ f_arrdiv24_fs267_xor0;
  assign f_arrdiv24_fs267_not1 = ~f_arrdiv24_fs267_xor0;
  assign f_arrdiv24_fs267_and1 = f_arrdiv24_fs267_not1 & f_arrdiv24_fs266_or0;
  assign f_arrdiv24_fs267_or0 = f_arrdiv24_fs267_and1 | f_arrdiv24_fs267_and0;
  assign f_arrdiv24_fs268_xor0 = f_arrdiv24_mux2to1233_xor0 ^ b[4];
  assign f_arrdiv24_fs268_not0 = ~f_arrdiv24_mux2to1233_xor0;
  assign f_arrdiv24_fs268_and0 = f_arrdiv24_fs268_not0 & b[4];
  assign f_arrdiv24_fs268_xor1 = f_arrdiv24_fs267_or0 ^ f_arrdiv24_fs268_xor0;
  assign f_arrdiv24_fs268_not1 = ~f_arrdiv24_fs268_xor0;
  assign f_arrdiv24_fs268_and1 = f_arrdiv24_fs268_not1 & f_arrdiv24_fs267_or0;
  assign f_arrdiv24_fs268_or0 = f_arrdiv24_fs268_and1 | f_arrdiv24_fs268_and0;
  assign f_arrdiv24_fs269_xor0 = f_arrdiv24_mux2to1234_xor0 ^ b[5];
  assign f_arrdiv24_fs269_not0 = ~f_arrdiv24_mux2to1234_xor0;
  assign f_arrdiv24_fs269_and0 = f_arrdiv24_fs269_not0 & b[5];
  assign f_arrdiv24_fs269_xor1 = f_arrdiv24_fs268_or0 ^ f_arrdiv24_fs269_xor0;
  assign f_arrdiv24_fs269_not1 = ~f_arrdiv24_fs269_xor0;
  assign f_arrdiv24_fs269_and1 = f_arrdiv24_fs269_not1 & f_arrdiv24_fs268_or0;
  assign f_arrdiv24_fs269_or0 = f_arrdiv24_fs269_and1 | f_arrdiv24_fs269_and0;
  assign f_arrdiv24_fs270_xor0 = f_arrdiv24_mux2to1235_xor0 ^ b[6];
  assign f_arrdiv24_fs270_not0 = ~f_arrdiv24_mux2to1235_xor0;
  assign f_arrdiv24_fs270_and0 = f_arrdiv24_fs270_not0 & b[6];
  assign f_arrdiv24_fs270_xor1 = f_arrdiv24_fs269_or0 ^ f_arrdiv24_fs270_xor0;
  assign f_arrdiv24_fs270_not1 = ~f_arrdiv24_fs270_xor0;
  assign f_arrdiv24_fs270_and1 = f_arrdiv24_fs270_not1 & f_arrdiv24_fs269_or0;
  assign f_arrdiv24_fs270_or0 = f_arrdiv24_fs270_and1 | f_arrdiv24_fs270_and0;
  assign f_arrdiv24_fs271_xor0 = f_arrdiv24_mux2to1236_xor0 ^ b[7];
  assign f_arrdiv24_fs271_not0 = ~f_arrdiv24_mux2to1236_xor0;
  assign f_arrdiv24_fs271_and0 = f_arrdiv24_fs271_not0 & b[7];
  assign f_arrdiv24_fs271_xor1 = f_arrdiv24_fs270_or0 ^ f_arrdiv24_fs271_xor0;
  assign f_arrdiv24_fs271_not1 = ~f_arrdiv24_fs271_xor0;
  assign f_arrdiv24_fs271_and1 = f_arrdiv24_fs271_not1 & f_arrdiv24_fs270_or0;
  assign f_arrdiv24_fs271_or0 = f_arrdiv24_fs271_and1 | f_arrdiv24_fs271_and0;
  assign f_arrdiv24_fs272_xor0 = f_arrdiv24_mux2to1237_xor0 ^ b[8];
  assign f_arrdiv24_fs272_not0 = ~f_arrdiv24_mux2to1237_xor0;
  assign f_arrdiv24_fs272_and0 = f_arrdiv24_fs272_not0 & b[8];
  assign f_arrdiv24_fs272_xor1 = f_arrdiv24_fs271_or0 ^ f_arrdiv24_fs272_xor0;
  assign f_arrdiv24_fs272_not1 = ~f_arrdiv24_fs272_xor0;
  assign f_arrdiv24_fs272_and1 = f_arrdiv24_fs272_not1 & f_arrdiv24_fs271_or0;
  assign f_arrdiv24_fs272_or0 = f_arrdiv24_fs272_and1 | f_arrdiv24_fs272_and0;
  assign f_arrdiv24_fs273_xor0 = f_arrdiv24_mux2to1238_xor0 ^ b[9];
  assign f_arrdiv24_fs273_not0 = ~f_arrdiv24_mux2to1238_xor0;
  assign f_arrdiv24_fs273_and0 = f_arrdiv24_fs273_not0 & b[9];
  assign f_arrdiv24_fs273_xor1 = f_arrdiv24_fs272_or0 ^ f_arrdiv24_fs273_xor0;
  assign f_arrdiv24_fs273_not1 = ~f_arrdiv24_fs273_xor0;
  assign f_arrdiv24_fs273_and1 = f_arrdiv24_fs273_not1 & f_arrdiv24_fs272_or0;
  assign f_arrdiv24_fs273_or0 = f_arrdiv24_fs273_and1 | f_arrdiv24_fs273_and0;
  assign f_arrdiv24_fs274_xor0 = f_arrdiv24_mux2to1239_xor0 ^ b[10];
  assign f_arrdiv24_fs274_not0 = ~f_arrdiv24_mux2to1239_xor0;
  assign f_arrdiv24_fs274_and0 = f_arrdiv24_fs274_not0 & b[10];
  assign f_arrdiv24_fs274_xor1 = f_arrdiv24_fs273_or0 ^ f_arrdiv24_fs274_xor0;
  assign f_arrdiv24_fs274_not1 = ~f_arrdiv24_fs274_xor0;
  assign f_arrdiv24_fs274_and1 = f_arrdiv24_fs274_not1 & f_arrdiv24_fs273_or0;
  assign f_arrdiv24_fs274_or0 = f_arrdiv24_fs274_and1 | f_arrdiv24_fs274_and0;
  assign f_arrdiv24_fs275_xor0 = f_arrdiv24_mux2to1240_xor0 ^ b[11];
  assign f_arrdiv24_fs275_not0 = ~f_arrdiv24_mux2to1240_xor0;
  assign f_arrdiv24_fs275_and0 = f_arrdiv24_fs275_not0 & b[11];
  assign f_arrdiv24_fs275_xor1 = f_arrdiv24_fs274_or0 ^ f_arrdiv24_fs275_xor0;
  assign f_arrdiv24_fs275_not1 = ~f_arrdiv24_fs275_xor0;
  assign f_arrdiv24_fs275_and1 = f_arrdiv24_fs275_not1 & f_arrdiv24_fs274_or0;
  assign f_arrdiv24_fs275_or0 = f_arrdiv24_fs275_and1 | f_arrdiv24_fs275_and0;
  assign f_arrdiv24_fs276_xor0 = f_arrdiv24_mux2to1241_xor0 ^ b[12];
  assign f_arrdiv24_fs276_not0 = ~f_arrdiv24_mux2to1241_xor0;
  assign f_arrdiv24_fs276_and0 = f_arrdiv24_fs276_not0 & b[12];
  assign f_arrdiv24_fs276_xor1 = f_arrdiv24_fs275_or0 ^ f_arrdiv24_fs276_xor0;
  assign f_arrdiv24_fs276_not1 = ~f_arrdiv24_fs276_xor0;
  assign f_arrdiv24_fs276_and1 = f_arrdiv24_fs276_not1 & f_arrdiv24_fs275_or0;
  assign f_arrdiv24_fs276_or0 = f_arrdiv24_fs276_and1 | f_arrdiv24_fs276_and0;
  assign f_arrdiv24_fs277_xor0 = f_arrdiv24_mux2to1242_xor0 ^ b[13];
  assign f_arrdiv24_fs277_not0 = ~f_arrdiv24_mux2to1242_xor0;
  assign f_arrdiv24_fs277_and0 = f_arrdiv24_fs277_not0 & b[13];
  assign f_arrdiv24_fs277_xor1 = f_arrdiv24_fs276_or0 ^ f_arrdiv24_fs277_xor0;
  assign f_arrdiv24_fs277_not1 = ~f_arrdiv24_fs277_xor0;
  assign f_arrdiv24_fs277_and1 = f_arrdiv24_fs277_not1 & f_arrdiv24_fs276_or0;
  assign f_arrdiv24_fs277_or0 = f_arrdiv24_fs277_and1 | f_arrdiv24_fs277_and0;
  assign f_arrdiv24_fs278_xor0 = f_arrdiv24_mux2to1243_xor0 ^ b[14];
  assign f_arrdiv24_fs278_not0 = ~f_arrdiv24_mux2to1243_xor0;
  assign f_arrdiv24_fs278_and0 = f_arrdiv24_fs278_not0 & b[14];
  assign f_arrdiv24_fs278_xor1 = f_arrdiv24_fs277_or0 ^ f_arrdiv24_fs278_xor0;
  assign f_arrdiv24_fs278_not1 = ~f_arrdiv24_fs278_xor0;
  assign f_arrdiv24_fs278_and1 = f_arrdiv24_fs278_not1 & f_arrdiv24_fs277_or0;
  assign f_arrdiv24_fs278_or0 = f_arrdiv24_fs278_and1 | f_arrdiv24_fs278_and0;
  assign f_arrdiv24_fs279_xor0 = f_arrdiv24_mux2to1244_xor0 ^ b[15];
  assign f_arrdiv24_fs279_not0 = ~f_arrdiv24_mux2to1244_xor0;
  assign f_arrdiv24_fs279_and0 = f_arrdiv24_fs279_not0 & b[15];
  assign f_arrdiv24_fs279_xor1 = f_arrdiv24_fs278_or0 ^ f_arrdiv24_fs279_xor0;
  assign f_arrdiv24_fs279_not1 = ~f_arrdiv24_fs279_xor0;
  assign f_arrdiv24_fs279_and1 = f_arrdiv24_fs279_not1 & f_arrdiv24_fs278_or0;
  assign f_arrdiv24_fs279_or0 = f_arrdiv24_fs279_and1 | f_arrdiv24_fs279_and0;
  assign f_arrdiv24_fs280_xor0 = f_arrdiv24_mux2to1245_xor0 ^ b[16];
  assign f_arrdiv24_fs280_not0 = ~f_arrdiv24_mux2to1245_xor0;
  assign f_arrdiv24_fs280_and0 = f_arrdiv24_fs280_not0 & b[16];
  assign f_arrdiv24_fs280_xor1 = f_arrdiv24_fs279_or0 ^ f_arrdiv24_fs280_xor0;
  assign f_arrdiv24_fs280_not1 = ~f_arrdiv24_fs280_xor0;
  assign f_arrdiv24_fs280_and1 = f_arrdiv24_fs280_not1 & f_arrdiv24_fs279_or0;
  assign f_arrdiv24_fs280_or0 = f_arrdiv24_fs280_and1 | f_arrdiv24_fs280_and0;
  assign f_arrdiv24_fs281_xor0 = f_arrdiv24_mux2to1246_xor0 ^ b[17];
  assign f_arrdiv24_fs281_not0 = ~f_arrdiv24_mux2to1246_xor0;
  assign f_arrdiv24_fs281_and0 = f_arrdiv24_fs281_not0 & b[17];
  assign f_arrdiv24_fs281_xor1 = f_arrdiv24_fs280_or0 ^ f_arrdiv24_fs281_xor0;
  assign f_arrdiv24_fs281_not1 = ~f_arrdiv24_fs281_xor0;
  assign f_arrdiv24_fs281_and1 = f_arrdiv24_fs281_not1 & f_arrdiv24_fs280_or0;
  assign f_arrdiv24_fs281_or0 = f_arrdiv24_fs281_and1 | f_arrdiv24_fs281_and0;
  assign f_arrdiv24_fs282_xor0 = f_arrdiv24_mux2to1247_xor0 ^ b[18];
  assign f_arrdiv24_fs282_not0 = ~f_arrdiv24_mux2to1247_xor0;
  assign f_arrdiv24_fs282_and0 = f_arrdiv24_fs282_not0 & b[18];
  assign f_arrdiv24_fs282_xor1 = f_arrdiv24_fs281_or0 ^ f_arrdiv24_fs282_xor0;
  assign f_arrdiv24_fs282_not1 = ~f_arrdiv24_fs282_xor0;
  assign f_arrdiv24_fs282_and1 = f_arrdiv24_fs282_not1 & f_arrdiv24_fs281_or0;
  assign f_arrdiv24_fs282_or0 = f_arrdiv24_fs282_and1 | f_arrdiv24_fs282_and0;
  assign f_arrdiv24_fs283_xor0 = f_arrdiv24_mux2to1248_xor0 ^ b[19];
  assign f_arrdiv24_fs283_not0 = ~f_arrdiv24_mux2to1248_xor0;
  assign f_arrdiv24_fs283_and0 = f_arrdiv24_fs283_not0 & b[19];
  assign f_arrdiv24_fs283_xor1 = f_arrdiv24_fs282_or0 ^ f_arrdiv24_fs283_xor0;
  assign f_arrdiv24_fs283_not1 = ~f_arrdiv24_fs283_xor0;
  assign f_arrdiv24_fs283_and1 = f_arrdiv24_fs283_not1 & f_arrdiv24_fs282_or0;
  assign f_arrdiv24_fs283_or0 = f_arrdiv24_fs283_and1 | f_arrdiv24_fs283_and0;
  assign f_arrdiv24_fs284_xor0 = f_arrdiv24_mux2to1249_xor0 ^ b[20];
  assign f_arrdiv24_fs284_not0 = ~f_arrdiv24_mux2to1249_xor0;
  assign f_arrdiv24_fs284_and0 = f_arrdiv24_fs284_not0 & b[20];
  assign f_arrdiv24_fs284_xor1 = f_arrdiv24_fs283_or0 ^ f_arrdiv24_fs284_xor0;
  assign f_arrdiv24_fs284_not1 = ~f_arrdiv24_fs284_xor0;
  assign f_arrdiv24_fs284_and1 = f_arrdiv24_fs284_not1 & f_arrdiv24_fs283_or0;
  assign f_arrdiv24_fs284_or0 = f_arrdiv24_fs284_and1 | f_arrdiv24_fs284_and0;
  assign f_arrdiv24_fs285_xor0 = f_arrdiv24_mux2to1250_xor0 ^ b[21];
  assign f_arrdiv24_fs285_not0 = ~f_arrdiv24_mux2to1250_xor0;
  assign f_arrdiv24_fs285_and0 = f_arrdiv24_fs285_not0 & b[21];
  assign f_arrdiv24_fs285_xor1 = f_arrdiv24_fs284_or0 ^ f_arrdiv24_fs285_xor0;
  assign f_arrdiv24_fs285_not1 = ~f_arrdiv24_fs285_xor0;
  assign f_arrdiv24_fs285_and1 = f_arrdiv24_fs285_not1 & f_arrdiv24_fs284_or0;
  assign f_arrdiv24_fs285_or0 = f_arrdiv24_fs285_and1 | f_arrdiv24_fs285_and0;
  assign f_arrdiv24_fs286_xor0 = f_arrdiv24_mux2to1251_xor0 ^ b[22];
  assign f_arrdiv24_fs286_not0 = ~f_arrdiv24_mux2to1251_xor0;
  assign f_arrdiv24_fs286_and0 = f_arrdiv24_fs286_not0 & b[22];
  assign f_arrdiv24_fs286_xor1 = f_arrdiv24_fs285_or0 ^ f_arrdiv24_fs286_xor0;
  assign f_arrdiv24_fs286_not1 = ~f_arrdiv24_fs286_xor0;
  assign f_arrdiv24_fs286_and1 = f_arrdiv24_fs286_not1 & f_arrdiv24_fs285_or0;
  assign f_arrdiv24_fs286_or0 = f_arrdiv24_fs286_and1 | f_arrdiv24_fs286_and0;
  assign f_arrdiv24_fs287_xor0 = f_arrdiv24_mux2to1252_xor0 ^ b[23];
  assign f_arrdiv24_fs287_not0 = ~f_arrdiv24_mux2to1252_xor0;
  assign f_arrdiv24_fs287_and0 = f_arrdiv24_fs287_not0 & b[23];
  assign f_arrdiv24_fs287_xor1 = f_arrdiv24_fs286_or0 ^ f_arrdiv24_fs287_xor0;
  assign f_arrdiv24_fs287_not1 = ~f_arrdiv24_fs287_xor0;
  assign f_arrdiv24_fs287_and1 = f_arrdiv24_fs287_not1 & f_arrdiv24_fs286_or0;
  assign f_arrdiv24_fs287_or0 = f_arrdiv24_fs287_and1 | f_arrdiv24_fs287_and0;
  assign f_arrdiv24_mux2to1253_and0 = a[12] & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1253_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1253_and1 = f_arrdiv24_fs264_xor0 & f_arrdiv24_mux2to1253_not0;
  assign f_arrdiv24_mux2to1253_xor0 = f_arrdiv24_mux2to1253_and0 ^ f_arrdiv24_mux2to1253_and1;
  assign f_arrdiv24_mux2to1254_and0 = f_arrdiv24_mux2to1230_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1254_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1254_and1 = f_arrdiv24_fs265_xor1 & f_arrdiv24_mux2to1254_not0;
  assign f_arrdiv24_mux2to1254_xor0 = f_arrdiv24_mux2to1254_and0 ^ f_arrdiv24_mux2to1254_and1;
  assign f_arrdiv24_mux2to1255_and0 = f_arrdiv24_mux2to1231_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1255_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1255_and1 = f_arrdiv24_fs266_xor1 & f_arrdiv24_mux2to1255_not0;
  assign f_arrdiv24_mux2to1255_xor0 = f_arrdiv24_mux2to1255_and0 ^ f_arrdiv24_mux2to1255_and1;
  assign f_arrdiv24_mux2to1256_and0 = f_arrdiv24_mux2to1232_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1256_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1256_and1 = f_arrdiv24_fs267_xor1 & f_arrdiv24_mux2to1256_not0;
  assign f_arrdiv24_mux2to1256_xor0 = f_arrdiv24_mux2to1256_and0 ^ f_arrdiv24_mux2to1256_and1;
  assign f_arrdiv24_mux2to1257_and0 = f_arrdiv24_mux2to1233_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1257_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1257_and1 = f_arrdiv24_fs268_xor1 & f_arrdiv24_mux2to1257_not0;
  assign f_arrdiv24_mux2to1257_xor0 = f_arrdiv24_mux2to1257_and0 ^ f_arrdiv24_mux2to1257_and1;
  assign f_arrdiv24_mux2to1258_and0 = f_arrdiv24_mux2to1234_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1258_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1258_and1 = f_arrdiv24_fs269_xor1 & f_arrdiv24_mux2to1258_not0;
  assign f_arrdiv24_mux2to1258_xor0 = f_arrdiv24_mux2to1258_and0 ^ f_arrdiv24_mux2to1258_and1;
  assign f_arrdiv24_mux2to1259_and0 = f_arrdiv24_mux2to1235_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1259_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1259_and1 = f_arrdiv24_fs270_xor1 & f_arrdiv24_mux2to1259_not0;
  assign f_arrdiv24_mux2to1259_xor0 = f_arrdiv24_mux2to1259_and0 ^ f_arrdiv24_mux2to1259_and1;
  assign f_arrdiv24_mux2to1260_and0 = f_arrdiv24_mux2to1236_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1260_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1260_and1 = f_arrdiv24_fs271_xor1 & f_arrdiv24_mux2to1260_not0;
  assign f_arrdiv24_mux2to1260_xor0 = f_arrdiv24_mux2to1260_and0 ^ f_arrdiv24_mux2to1260_and1;
  assign f_arrdiv24_mux2to1261_and0 = f_arrdiv24_mux2to1237_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1261_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1261_and1 = f_arrdiv24_fs272_xor1 & f_arrdiv24_mux2to1261_not0;
  assign f_arrdiv24_mux2to1261_xor0 = f_arrdiv24_mux2to1261_and0 ^ f_arrdiv24_mux2to1261_and1;
  assign f_arrdiv24_mux2to1262_and0 = f_arrdiv24_mux2to1238_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1262_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1262_and1 = f_arrdiv24_fs273_xor1 & f_arrdiv24_mux2to1262_not0;
  assign f_arrdiv24_mux2to1262_xor0 = f_arrdiv24_mux2to1262_and0 ^ f_arrdiv24_mux2to1262_and1;
  assign f_arrdiv24_mux2to1263_and0 = f_arrdiv24_mux2to1239_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1263_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1263_and1 = f_arrdiv24_fs274_xor1 & f_arrdiv24_mux2to1263_not0;
  assign f_arrdiv24_mux2to1263_xor0 = f_arrdiv24_mux2to1263_and0 ^ f_arrdiv24_mux2to1263_and1;
  assign f_arrdiv24_mux2to1264_and0 = f_arrdiv24_mux2to1240_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1264_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1264_and1 = f_arrdiv24_fs275_xor1 & f_arrdiv24_mux2to1264_not0;
  assign f_arrdiv24_mux2to1264_xor0 = f_arrdiv24_mux2to1264_and0 ^ f_arrdiv24_mux2to1264_and1;
  assign f_arrdiv24_mux2to1265_and0 = f_arrdiv24_mux2to1241_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1265_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1265_and1 = f_arrdiv24_fs276_xor1 & f_arrdiv24_mux2to1265_not0;
  assign f_arrdiv24_mux2to1265_xor0 = f_arrdiv24_mux2to1265_and0 ^ f_arrdiv24_mux2to1265_and1;
  assign f_arrdiv24_mux2to1266_and0 = f_arrdiv24_mux2to1242_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1266_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1266_and1 = f_arrdiv24_fs277_xor1 & f_arrdiv24_mux2to1266_not0;
  assign f_arrdiv24_mux2to1266_xor0 = f_arrdiv24_mux2to1266_and0 ^ f_arrdiv24_mux2to1266_and1;
  assign f_arrdiv24_mux2to1267_and0 = f_arrdiv24_mux2to1243_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1267_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1267_and1 = f_arrdiv24_fs278_xor1 & f_arrdiv24_mux2to1267_not0;
  assign f_arrdiv24_mux2to1267_xor0 = f_arrdiv24_mux2to1267_and0 ^ f_arrdiv24_mux2to1267_and1;
  assign f_arrdiv24_mux2to1268_and0 = f_arrdiv24_mux2to1244_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1268_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1268_and1 = f_arrdiv24_fs279_xor1 & f_arrdiv24_mux2to1268_not0;
  assign f_arrdiv24_mux2to1268_xor0 = f_arrdiv24_mux2to1268_and0 ^ f_arrdiv24_mux2to1268_and1;
  assign f_arrdiv24_mux2to1269_and0 = f_arrdiv24_mux2to1245_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1269_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1269_and1 = f_arrdiv24_fs280_xor1 & f_arrdiv24_mux2to1269_not0;
  assign f_arrdiv24_mux2to1269_xor0 = f_arrdiv24_mux2to1269_and0 ^ f_arrdiv24_mux2to1269_and1;
  assign f_arrdiv24_mux2to1270_and0 = f_arrdiv24_mux2to1246_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1270_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1270_and1 = f_arrdiv24_fs281_xor1 & f_arrdiv24_mux2to1270_not0;
  assign f_arrdiv24_mux2to1270_xor0 = f_arrdiv24_mux2to1270_and0 ^ f_arrdiv24_mux2to1270_and1;
  assign f_arrdiv24_mux2to1271_and0 = f_arrdiv24_mux2to1247_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1271_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1271_and1 = f_arrdiv24_fs282_xor1 & f_arrdiv24_mux2to1271_not0;
  assign f_arrdiv24_mux2to1271_xor0 = f_arrdiv24_mux2to1271_and0 ^ f_arrdiv24_mux2to1271_and1;
  assign f_arrdiv24_mux2to1272_and0 = f_arrdiv24_mux2to1248_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1272_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1272_and1 = f_arrdiv24_fs283_xor1 & f_arrdiv24_mux2to1272_not0;
  assign f_arrdiv24_mux2to1272_xor0 = f_arrdiv24_mux2to1272_and0 ^ f_arrdiv24_mux2to1272_and1;
  assign f_arrdiv24_mux2to1273_and0 = f_arrdiv24_mux2to1249_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1273_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1273_and1 = f_arrdiv24_fs284_xor1 & f_arrdiv24_mux2to1273_not0;
  assign f_arrdiv24_mux2to1273_xor0 = f_arrdiv24_mux2to1273_and0 ^ f_arrdiv24_mux2to1273_and1;
  assign f_arrdiv24_mux2to1274_and0 = f_arrdiv24_mux2to1250_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1274_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1274_and1 = f_arrdiv24_fs285_xor1 & f_arrdiv24_mux2to1274_not0;
  assign f_arrdiv24_mux2to1274_xor0 = f_arrdiv24_mux2to1274_and0 ^ f_arrdiv24_mux2to1274_and1;
  assign f_arrdiv24_mux2to1275_and0 = f_arrdiv24_mux2to1251_xor0 & f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1275_not0 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_mux2to1275_and1 = f_arrdiv24_fs286_xor1 & f_arrdiv24_mux2to1275_not0;
  assign f_arrdiv24_mux2to1275_xor0 = f_arrdiv24_mux2to1275_and0 ^ f_arrdiv24_mux2to1275_and1;
  assign f_arrdiv24_not11 = ~f_arrdiv24_fs287_or0;
  assign f_arrdiv24_fs288_xor0 = a[11] ^ b[0];
  assign f_arrdiv24_fs288_not0 = ~a[11];
  assign f_arrdiv24_fs288_and0 = f_arrdiv24_fs288_not0 & b[0];
  assign f_arrdiv24_fs288_not1 = ~f_arrdiv24_fs288_xor0;
  assign f_arrdiv24_fs289_xor0 = f_arrdiv24_mux2to1253_xor0 ^ b[1];
  assign f_arrdiv24_fs289_not0 = ~f_arrdiv24_mux2to1253_xor0;
  assign f_arrdiv24_fs289_and0 = f_arrdiv24_fs289_not0 & b[1];
  assign f_arrdiv24_fs289_xor1 = f_arrdiv24_fs288_and0 ^ f_arrdiv24_fs289_xor0;
  assign f_arrdiv24_fs289_not1 = ~f_arrdiv24_fs289_xor0;
  assign f_arrdiv24_fs289_and1 = f_arrdiv24_fs289_not1 & f_arrdiv24_fs288_and0;
  assign f_arrdiv24_fs289_or0 = f_arrdiv24_fs289_and1 | f_arrdiv24_fs289_and0;
  assign f_arrdiv24_fs290_xor0 = f_arrdiv24_mux2to1254_xor0 ^ b[2];
  assign f_arrdiv24_fs290_not0 = ~f_arrdiv24_mux2to1254_xor0;
  assign f_arrdiv24_fs290_and0 = f_arrdiv24_fs290_not0 & b[2];
  assign f_arrdiv24_fs290_xor1 = f_arrdiv24_fs289_or0 ^ f_arrdiv24_fs290_xor0;
  assign f_arrdiv24_fs290_not1 = ~f_arrdiv24_fs290_xor0;
  assign f_arrdiv24_fs290_and1 = f_arrdiv24_fs290_not1 & f_arrdiv24_fs289_or0;
  assign f_arrdiv24_fs290_or0 = f_arrdiv24_fs290_and1 | f_arrdiv24_fs290_and0;
  assign f_arrdiv24_fs291_xor0 = f_arrdiv24_mux2to1255_xor0 ^ b[3];
  assign f_arrdiv24_fs291_not0 = ~f_arrdiv24_mux2to1255_xor0;
  assign f_arrdiv24_fs291_and0 = f_arrdiv24_fs291_not0 & b[3];
  assign f_arrdiv24_fs291_xor1 = f_arrdiv24_fs290_or0 ^ f_arrdiv24_fs291_xor0;
  assign f_arrdiv24_fs291_not1 = ~f_arrdiv24_fs291_xor0;
  assign f_arrdiv24_fs291_and1 = f_arrdiv24_fs291_not1 & f_arrdiv24_fs290_or0;
  assign f_arrdiv24_fs291_or0 = f_arrdiv24_fs291_and1 | f_arrdiv24_fs291_and0;
  assign f_arrdiv24_fs292_xor0 = f_arrdiv24_mux2to1256_xor0 ^ b[4];
  assign f_arrdiv24_fs292_not0 = ~f_arrdiv24_mux2to1256_xor0;
  assign f_arrdiv24_fs292_and0 = f_arrdiv24_fs292_not0 & b[4];
  assign f_arrdiv24_fs292_xor1 = f_arrdiv24_fs291_or0 ^ f_arrdiv24_fs292_xor0;
  assign f_arrdiv24_fs292_not1 = ~f_arrdiv24_fs292_xor0;
  assign f_arrdiv24_fs292_and1 = f_arrdiv24_fs292_not1 & f_arrdiv24_fs291_or0;
  assign f_arrdiv24_fs292_or0 = f_arrdiv24_fs292_and1 | f_arrdiv24_fs292_and0;
  assign f_arrdiv24_fs293_xor0 = f_arrdiv24_mux2to1257_xor0 ^ b[5];
  assign f_arrdiv24_fs293_not0 = ~f_arrdiv24_mux2to1257_xor0;
  assign f_arrdiv24_fs293_and0 = f_arrdiv24_fs293_not0 & b[5];
  assign f_arrdiv24_fs293_xor1 = f_arrdiv24_fs292_or0 ^ f_arrdiv24_fs293_xor0;
  assign f_arrdiv24_fs293_not1 = ~f_arrdiv24_fs293_xor0;
  assign f_arrdiv24_fs293_and1 = f_arrdiv24_fs293_not1 & f_arrdiv24_fs292_or0;
  assign f_arrdiv24_fs293_or0 = f_arrdiv24_fs293_and1 | f_arrdiv24_fs293_and0;
  assign f_arrdiv24_fs294_xor0 = f_arrdiv24_mux2to1258_xor0 ^ b[6];
  assign f_arrdiv24_fs294_not0 = ~f_arrdiv24_mux2to1258_xor0;
  assign f_arrdiv24_fs294_and0 = f_arrdiv24_fs294_not0 & b[6];
  assign f_arrdiv24_fs294_xor1 = f_arrdiv24_fs293_or0 ^ f_arrdiv24_fs294_xor0;
  assign f_arrdiv24_fs294_not1 = ~f_arrdiv24_fs294_xor0;
  assign f_arrdiv24_fs294_and1 = f_arrdiv24_fs294_not1 & f_arrdiv24_fs293_or0;
  assign f_arrdiv24_fs294_or0 = f_arrdiv24_fs294_and1 | f_arrdiv24_fs294_and0;
  assign f_arrdiv24_fs295_xor0 = f_arrdiv24_mux2to1259_xor0 ^ b[7];
  assign f_arrdiv24_fs295_not0 = ~f_arrdiv24_mux2to1259_xor0;
  assign f_arrdiv24_fs295_and0 = f_arrdiv24_fs295_not0 & b[7];
  assign f_arrdiv24_fs295_xor1 = f_arrdiv24_fs294_or0 ^ f_arrdiv24_fs295_xor0;
  assign f_arrdiv24_fs295_not1 = ~f_arrdiv24_fs295_xor0;
  assign f_arrdiv24_fs295_and1 = f_arrdiv24_fs295_not1 & f_arrdiv24_fs294_or0;
  assign f_arrdiv24_fs295_or0 = f_arrdiv24_fs295_and1 | f_arrdiv24_fs295_and0;
  assign f_arrdiv24_fs296_xor0 = f_arrdiv24_mux2to1260_xor0 ^ b[8];
  assign f_arrdiv24_fs296_not0 = ~f_arrdiv24_mux2to1260_xor0;
  assign f_arrdiv24_fs296_and0 = f_arrdiv24_fs296_not0 & b[8];
  assign f_arrdiv24_fs296_xor1 = f_arrdiv24_fs295_or0 ^ f_arrdiv24_fs296_xor0;
  assign f_arrdiv24_fs296_not1 = ~f_arrdiv24_fs296_xor0;
  assign f_arrdiv24_fs296_and1 = f_arrdiv24_fs296_not1 & f_arrdiv24_fs295_or0;
  assign f_arrdiv24_fs296_or0 = f_arrdiv24_fs296_and1 | f_arrdiv24_fs296_and0;
  assign f_arrdiv24_fs297_xor0 = f_arrdiv24_mux2to1261_xor0 ^ b[9];
  assign f_arrdiv24_fs297_not0 = ~f_arrdiv24_mux2to1261_xor0;
  assign f_arrdiv24_fs297_and0 = f_arrdiv24_fs297_not0 & b[9];
  assign f_arrdiv24_fs297_xor1 = f_arrdiv24_fs296_or0 ^ f_arrdiv24_fs297_xor0;
  assign f_arrdiv24_fs297_not1 = ~f_arrdiv24_fs297_xor0;
  assign f_arrdiv24_fs297_and1 = f_arrdiv24_fs297_not1 & f_arrdiv24_fs296_or0;
  assign f_arrdiv24_fs297_or0 = f_arrdiv24_fs297_and1 | f_arrdiv24_fs297_and0;
  assign f_arrdiv24_fs298_xor0 = f_arrdiv24_mux2to1262_xor0 ^ b[10];
  assign f_arrdiv24_fs298_not0 = ~f_arrdiv24_mux2to1262_xor0;
  assign f_arrdiv24_fs298_and0 = f_arrdiv24_fs298_not0 & b[10];
  assign f_arrdiv24_fs298_xor1 = f_arrdiv24_fs297_or0 ^ f_arrdiv24_fs298_xor0;
  assign f_arrdiv24_fs298_not1 = ~f_arrdiv24_fs298_xor0;
  assign f_arrdiv24_fs298_and1 = f_arrdiv24_fs298_not1 & f_arrdiv24_fs297_or0;
  assign f_arrdiv24_fs298_or0 = f_arrdiv24_fs298_and1 | f_arrdiv24_fs298_and0;
  assign f_arrdiv24_fs299_xor0 = f_arrdiv24_mux2to1263_xor0 ^ b[11];
  assign f_arrdiv24_fs299_not0 = ~f_arrdiv24_mux2to1263_xor0;
  assign f_arrdiv24_fs299_and0 = f_arrdiv24_fs299_not0 & b[11];
  assign f_arrdiv24_fs299_xor1 = f_arrdiv24_fs298_or0 ^ f_arrdiv24_fs299_xor0;
  assign f_arrdiv24_fs299_not1 = ~f_arrdiv24_fs299_xor0;
  assign f_arrdiv24_fs299_and1 = f_arrdiv24_fs299_not1 & f_arrdiv24_fs298_or0;
  assign f_arrdiv24_fs299_or0 = f_arrdiv24_fs299_and1 | f_arrdiv24_fs299_and0;
  assign f_arrdiv24_fs300_xor0 = f_arrdiv24_mux2to1264_xor0 ^ b[12];
  assign f_arrdiv24_fs300_not0 = ~f_arrdiv24_mux2to1264_xor0;
  assign f_arrdiv24_fs300_and0 = f_arrdiv24_fs300_not0 & b[12];
  assign f_arrdiv24_fs300_xor1 = f_arrdiv24_fs299_or0 ^ f_arrdiv24_fs300_xor0;
  assign f_arrdiv24_fs300_not1 = ~f_arrdiv24_fs300_xor0;
  assign f_arrdiv24_fs300_and1 = f_arrdiv24_fs300_not1 & f_arrdiv24_fs299_or0;
  assign f_arrdiv24_fs300_or0 = f_arrdiv24_fs300_and1 | f_arrdiv24_fs300_and0;
  assign f_arrdiv24_fs301_xor0 = f_arrdiv24_mux2to1265_xor0 ^ b[13];
  assign f_arrdiv24_fs301_not0 = ~f_arrdiv24_mux2to1265_xor0;
  assign f_arrdiv24_fs301_and0 = f_arrdiv24_fs301_not0 & b[13];
  assign f_arrdiv24_fs301_xor1 = f_arrdiv24_fs300_or0 ^ f_arrdiv24_fs301_xor0;
  assign f_arrdiv24_fs301_not1 = ~f_arrdiv24_fs301_xor0;
  assign f_arrdiv24_fs301_and1 = f_arrdiv24_fs301_not1 & f_arrdiv24_fs300_or0;
  assign f_arrdiv24_fs301_or0 = f_arrdiv24_fs301_and1 | f_arrdiv24_fs301_and0;
  assign f_arrdiv24_fs302_xor0 = f_arrdiv24_mux2to1266_xor0 ^ b[14];
  assign f_arrdiv24_fs302_not0 = ~f_arrdiv24_mux2to1266_xor0;
  assign f_arrdiv24_fs302_and0 = f_arrdiv24_fs302_not0 & b[14];
  assign f_arrdiv24_fs302_xor1 = f_arrdiv24_fs301_or0 ^ f_arrdiv24_fs302_xor0;
  assign f_arrdiv24_fs302_not1 = ~f_arrdiv24_fs302_xor0;
  assign f_arrdiv24_fs302_and1 = f_arrdiv24_fs302_not1 & f_arrdiv24_fs301_or0;
  assign f_arrdiv24_fs302_or0 = f_arrdiv24_fs302_and1 | f_arrdiv24_fs302_and0;
  assign f_arrdiv24_fs303_xor0 = f_arrdiv24_mux2to1267_xor0 ^ b[15];
  assign f_arrdiv24_fs303_not0 = ~f_arrdiv24_mux2to1267_xor0;
  assign f_arrdiv24_fs303_and0 = f_arrdiv24_fs303_not0 & b[15];
  assign f_arrdiv24_fs303_xor1 = f_arrdiv24_fs302_or0 ^ f_arrdiv24_fs303_xor0;
  assign f_arrdiv24_fs303_not1 = ~f_arrdiv24_fs303_xor0;
  assign f_arrdiv24_fs303_and1 = f_arrdiv24_fs303_not1 & f_arrdiv24_fs302_or0;
  assign f_arrdiv24_fs303_or0 = f_arrdiv24_fs303_and1 | f_arrdiv24_fs303_and0;
  assign f_arrdiv24_fs304_xor0 = f_arrdiv24_mux2to1268_xor0 ^ b[16];
  assign f_arrdiv24_fs304_not0 = ~f_arrdiv24_mux2to1268_xor0;
  assign f_arrdiv24_fs304_and0 = f_arrdiv24_fs304_not0 & b[16];
  assign f_arrdiv24_fs304_xor1 = f_arrdiv24_fs303_or0 ^ f_arrdiv24_fs304_xor0;
  assign f_arrdiv24_fs304_not1 = ~f_arrdiv24_fs304_xor0;
  assign f_arrdiv24_fs304_and1 = f_arrdiv24_fs304_not1 & f_arrdiv24_fs303_or0;
  assign f_arrdiv24_fs304_or0 = f_arrdiv24_fs304_and1 | f_arrdiv24_fs304_and0;
  assign f_arrdiv24_fs305_xor0 = f_arrdiv24_mux2to1269_xor0 ^ b[17];
  assign f_arrdiv24_fs305_not0 = ~f_arrdiv24_mux2to1269_xor0;
  assign f_arrdiv24_fs305_and0 = f_arrdiv24_fs305_not0 & b[17];
  assign f_arrdiv24_fs305_xor1 = f_arrdiv24_fs304_or0 ^ f_arrdiv24_fs305_xor0;
  assign f_arrdiv24_fs305_not1 = ~f_arrdiv24_fs305_xor0;
  assign f_arrdiv24_fs305_and1 = f_arrdiv24_fs305_not1 & f_arrdiv24_fs304_or0;
  assign f_arrdiv24_fs305_or0 = f_arrdiv24_fs305_and1 | f_arrdiv24_fs305_and0;
  assign f_arrdiv24_fs306_xor0 = f_arrdiv24_mux2to1270_xor0 ^ b[18];
  assign f_arrdiv24_fs306_not0 = ~f_arrdiv24_mux2to1270_xor0;
  assign f_arrdiv24_fs306_and0 = f_arrdiv24_fs306_not0 & b[18];
  assign f_arrdiv24_fs306_xor1 = f_arrdiv24_fs305_or0 ^ f_arrdiv24_fs306_xor0;
  assign f_arrdiv24_fs306_not1 = ~f_arrdiv24_fs306_xor0;
  assign f_arrdiv24_fs306_and1 = f_arrdiv24_fs306_not1 & f_arrdiv24_fs305_or0;
  assign f_arrdiv24_fs306_or0 = f_arrdiv24_fs306_and1 | f_arrdiv24_fs306_and0;
  assign f_arrdiv24_fs307_xor0 = f_arrdiv24_mux2to1271_xor0 ^ b[19];
  assign f_arrdiv24_fs307_not0 = ~f_arrdiv24_mux2to1271_xor0;
  assign f_arrdiv24_fs307_and0 = f_arrdiv24_fs307_not0 & b[19];
  assign f_arrdiv24_fs307_xor1 = f_arrdiv24_fs306_or0 ^ f_arrdiv24_fs307_xor0;
  assign f_arrdiv24_fs307_not1 = ~f_arrdiv24_fs307_xor0;
  assign f_arrdiv24_fs307_and1 = f_arrdiv24_fs307_not1 & f_arrdiv24_fs306_or0;
  assign f_arrdiv24_fs307_or0 = f_arrdiv24_fs307_and1 | f_arrdiv24_fs307_and0;
  assign f_arrdiv24_fs308_xor0 = f_arrdiv24_mux2to1272_xor0 ^ b[20];
  assign f_arrdiv24_fs308_not0 = ~f_arrdiv24_mux2to1272_xor0;
  assign f_arrdiv24_fs308_and0 = f_arrdiv24_fs308_not0 & b[20];
  assign f_arrdiv24_fs308_xor1 = f_arrdiv24_fs307_or0 ^ f_arrdiv24_fs308_xor0;
  assign f_arrdiv24_fs308_not1 = ~f_arrdiv24_fs308_xor0;
  assign f_arrdiv24_fs308_and1 = f_arrdiv24_fs308_not1 & f_arrdiv24_fs307_or0;
  assign f_arrdiv24_fs308_or0 = f_arrdiv24_fs308_and1 | f_arrdiv24_fs308_and0;
  assign f_arrdiv24_fs309_xor0 = f_arrdiv24_mux2to1273_xor0 ^ b[21];
  assign f_arrdiv24_fs309_not0 = ~f_arrdiv24_mux2to1273_xor0;
  assign f_arrdiv24_fs309_and0 = f_arrdiv24_fs309_not0 & b[21];
  assign f_arrdiv24_fs309_xor1 = f_arrdiv24_fs308_or0 ^ f_arrdiv24_fs309_xor0;
  assign f_arrdiv24_fs309_not1 = ~f_arrdiv24_fs309_xor0;
  assign f_arrdiv24_fs309_and1 = f_arrdiv24_fs309_not1 & f_arrdiv24_fs308_or0;
  assign f_arrdiv24_fs309_or0 = f_arrdiv24_fs309_and1 | f_arrdiv24_fs309_and0;
  assign f_arrdiv24_fs310_xor0 = f_arrdiv24_mux2to1274_xor0 ^ b[22];
  assign f_arrdiv24_fs310_not0 = ~f_arrdiv24_mux2to1274_xor0;
  assign f_arrdiv24_fs310_and0 = f_arrdiv24_fs310_not0 & b[22];
  assign f_arrdiv24_fs310_xor1 = f_arrdiv24_fs309_or0 ^ f_arrdiv24_fs310_xor0;
  assign f_arrdiv24_fs310_not1 = ~f_arrdiv24_fs310_xor0;
  assign f_arrdiv24_fs310_and1 = f_arrdiv24_fs310_not1 & f_arrdiv24_fs309_or0;
  assign f_arrdiv24_fs310_or0 = f_arrdiv24_fs310_and1 | f_arrdiv24_fs310_and0;
  assign f_arrdiv24_fs311_xor0 = f_arrdiv24_mux2to1275_xor0 ^ b[23];
  assign f_arrdiv24_fs311_not0 = ~f_arrdiv24_mux2to1275_xor0;
  assign f_arrdiv24_fs311_and0 = f_arrdiv24_fs311_not0 & b[23];
  assign f_arrdiv24_fs311_xor1 = f_arrdiv24_fs310_or0 ^ f_arrdiv24_fs311_xor0;
  assign f_arrdiv24_fs311_not1 = ~f_arrdiv24_fs311_xor0;
  assign f_arrdiv24_fs311_and1 = f_arrdiv24_fs311_not1 & f_arrdiv24_fs310_or0;
  assign f_arrdiv24_fs311_or0 = f_arrdiv24_fs311_and1 | f_arrdiv24_fs311_and0;
  assign f_arrdiv24_mux2to1276_and0 = a[11] & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1276_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1276_and1 = f_arrdiv24_fs288_xor0 & f_arrdiv24_mux2to1276_not0;
  assign f_arrdiv24_mux2to1276_xor0 = f_arrdiv24_mux2to1276_and0 ^ f_arrdiv24_mux2to1276_and1;
  assign f_arrdiv24_mux2to1277_and0 = f_arrdiv24_mux2to1253_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1277_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1277_and1 = f_arrdiv24_fs289_xor1 & f_arrdiv24_mux2to1277_not0;
  assign f_arrdiv24_mux2to1277_xor0 = f_arrdiv24_mux2to1277_and0 ^ f_arrdiv24_mux2to1277_and1;
  assign f_arrdiv24_mux2to1278_and0 = f_arrdiv24_mux2to1254_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1278_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1278_and1 = f_arrdiv24_fs290_xor1 & f_arrdiv24_mux2to1278_not0;
  assign f_arrdiv24_mux2to1278_xor0 = f_arrdiv24_mux2to1278_and0 ^ f_arrdiv24_mux2to1278_and1;
  assign f_arrdiv24_mux2to1279_and0 = f_arrdiv24_mux2to1255_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1279_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1279_and1 = f_arrdiv24_fs291_xor1 & f_arrdiv24_mux2to1279_not0;
  assign f_arrdiv24_mux2to1279_xor0 = f_arrdiv24_mux2to1279_and0 ^ f_arrdiv24_mux2to1279_and1;
  assign f_arrdiv24_mux2to1280_and0 = f_arrdiv24_mux2to1256_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1280_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1280_and1 = f_arrdiv24_fs292_xor1 & f_arrdiv24_mux2to1280_not0;
  assign f_arrdiv24_mux2to1280_xor0 = f_arrdiv24_mux2to1280_and0 ^ f_arrdiv24_mux2to1280_and1;
  assign f_arrdiv24_mux2to1281_and0 = f_arrdiv24_mux2to1257_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1281_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1281_and1 = f_arrdiv24_fs293_xor1 & f_arrdiv24_mux2to1281_not0;
  assign f_arrdiv24_mux2to1281_xor0 = f_arrdiv24_mux2to1281_and0 ^ f_arrdiv24_mux2to1281_and1;
  assign f_arrdiv24_mux2to1282_and0 = f_arrdiv24_mux2to1258_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1282_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1282_and1 = f_arrdiv24_fs294_xor1 & f_arrdiv24_mux2to1282_not0;
  assign f_arrdiv24_mux2to1282_xor0 = f_arrdiv24_mux2to1282_and0 ^ f_arrdiv24_mux2to1282_and1;
  assign f_arrdiv24_mux2to1283_and0 = f_arrdiv24_mux2to1259_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1283_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1283_and1 = f_arrdiv24_fs295_xor1 & f_arrdiv24_mux2to1283_not0;
  assign f_arrdiv24_mux2to1283_xor0 = f_arrdiv24_mux2to1283_and0 ^ f_arrdiv24_mux2to1283_and1;
  assign f_arrdiv24_mux2to1284_and0 = f_arrdiv24_mux2to1260_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1284_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1284_and1 = f_arrdiv24_fs296_xor1 & f_arrdiv24_mux2to1284_not0;
  assign f_arrdiv24_mux2to1284_xor0 = f_arrdiv24_mux2to1284_and0 ^ f_arrdiv24_mux2to1284_and1;
  assign f_arrdiv24_mux2to1285_and0 = f_arrdiv24_mux2to1261_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1285_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1285_and1 = f_arrdiv24_fs297_xor1 & f_arrdiv24_mux2to1285_not0;
  assign f_arrdiv24_mux2to1285_xor0 = f_arrdiv24_mux2to1285_and0 ^ f_arrdiv24_mux2to1285_and1;
  assign f_arrdiv24_mux2to1286_and0 = f_arrdiv24_mux2to1262_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1286_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1286_and1 = f_arrdiv24_fs298_xor1 & f_arrdiv24_mux2to1286_not0;
  assign f_arrdiv24_mux2to1286_xor0 = f_arrdiv24_mux2to1286_and0 ^ f_arrdiv24_mux2to1286_and1;
  assign f_arrdiv24_mux2to1287_and0 = f_arrdiv24_mux2to1263_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1287_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1287_and1 = f_arrdiv24_fs299_xor1 & f_arrdiv24_mux2to1287_not0;
  assign f_arrdiv24_mux2to1287_xor0 = f_arrdiv24_mux2to1287_and0 ^ f_arrdiv24_mux2to1287_and1;
  assign f_arrdiv24_mux2to1288_and0 = f_arrdiv24_mux2to1264_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1288_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1288_and1 = f_arrdiv24_fs300_xor1 & f_arrdiv24_mux2to1288_not0;
  assign f_arrdiv24_mux2to1288_xor0 = f_arrdiv24_mux2to1288_and0 ^ f_arrdiv24_mux2to1288_and1;
  assign f_arrdiv24_mux2to1289_and0 = f_arrdiv24_mux2to1265_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1289_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1289_and1 = f_arrdiv24_fs301_xor1 & f_arrdiv24_mux2to1289_not0;
  assign f_arrdiv24_mux2to1289_xor0 = f_arrdiv24_mux2to1289_and0 ^ f_arrdiv24_mux2to1289_and1;
  assign f_arrdiv24_mux2to1290_and0 = f_arrdiv24_mux2to1266_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1290_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1290_and1 = f_arrdiv24_fs302_xor1 & f_arrdiv24_mux2to1290_not0;
  assign f_arrdiv24_mux2to1290_xor0 = f_arrdiv24_mux2to1290_and0 ^ f_arrdiv24_mux2to1290_and1;
  assign f_arrdiv24_mux2to1291_and0 = f_arrdiv24_mux2to1267_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1291_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1291_and1 = f_arrdiv24_fs303_xor1 & f_arrdiv24_mux2to1291_not0;
  assign f_arrdiv24_mux2to1291_xor0 = f_arrdiv24_mux2to1291_and0 ^ f_arrdiv24_mux2to1291_and1;
  assign f_arrdiv24_mux2to1292_and0 = f_arrdiv24_mux2to1268_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1292_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1292_and1 = f_arrdiv24_fs304_xor1 & f_arrdiv24_mux2to1292_not0;
  assign f_arrdiv24_mux2to1292_xor0 = f_arrdiv24_mux2to1292_and0 ^ f_arrdiv24_mux2to1292_and1;
  assign f_arrdiv24_mux2to1293_and0 = f_arrdiv24_mux2to1269_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1293_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1293_and1 = f_arrdiv24_fs305_xor1 & f_arrdiv24_mux2to1293_not0;
  assign f_arrdiv24_mux2to1293_xor0 = f_arrdiv24_mux2to1293_and0 ^ f_arrdiv24_mux2to1293_and1;
  assign f_arrdiv24_mux2to1294_and0 = f_arrdiv24_mux2to1270_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1294_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1294_and1 = f_arrdiv24_fs306_xor1 & f_arrdiv24_mux2to1294_not0;
  assign f_arrdiv24_mux2to1294_xor0 = f_arrdiv24_mux2to1294_and0 ^ f_arrdiv24_mux2to1294_and1;
  assign f_arrdiv24_mux2to1295_and0 = f_arrdiv24_mux2to1271_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1295_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1295_and1 = f_arrdiv24_fs307_xor1 & f_arrdiv24_mux2to1295_not0;
  assign f_arrdiv24_mux2to1295_xor0 = f_arrdiv24_mux2to1295_and0 ^ f_arrdiv24_mux2to1295_and1;
  assign f_arrdiv24_mux2to1296_and0 = f_arrdiv24_mux2to1272_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1296_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1296_and1 = f_arrdiv24_fs308_xor1 & f_arrdiv24_mux2to1296_not0;
  assign f_arrdiv24_mux2to1296_xor0 = f_arrdiv24_mux2to1296_and0 ^ f_arrdiv24_mux2to1296_and1;
  assign f_arrdiv24_mux2to1297_and0 = f_arrdiv24_mux2to1273_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1297_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1297_and1 = f_arrdiv24_fs309_xor1 & f_arrdiv24_mux2to1297_not0;
  assign f_arrdiv24_mux2to1297_xor0 = f_arrdiv24_mux2to1297_and0 ^ f_arrdiv24_mux2to1297_and1;
  assign f_arrdiv24_mux2to1298_and0 = f_arrdiv24_mux2to1274_xor0 & f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1298_not0 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_mux2to1298_and1 = f_arrdiv24_fs310_xor1 & f_arrdiv24_mux2to1298_not0;
  assign f_arrdiv24_mux2to1298_xor0 = f_arrdiv24_mux2to1298_and0 ^ f_arrdiv24_mux2to1298_and1;
  assign f_arrdiv24_not12 = ~f_arrdiv24_fs311_or0;
  assign f_arrdiv24_fs312_xor0 = a[10] ^ b[0];
  assign f_arrdiv24_fs312_not0 = ~a[10];
  assign f_arrdiv24_fs312_and0 = f_arrdiv24_fs312_not0 & b[0];
  assign f_arrdiv24_fs312_not1 = ~f_arrdiv24_fs312_xor0;
  assign f_arrdiv24_fs313_xor0 = f_arrdiv24_mux2to1276_xor0 ^ b[1];
  assign f_arrdiv24_fs313_not0 = ~f_arrdiv24_mux2to1276_xor0;
  assign f_arrdiv24_fs313_and0 = f_arrdiv24_fs313_not0 & b[1];
  assign f_arrdiv24_fs313_xor1 = f_arrdiv24_fs312_and0 ^ f_arrdiv24_fs313_xor0;
  assign f_arrdiv24_fs313_not1 = ~f_arrdiv24_fs313_xor0;
  assign f_arrdiv24_fs313_and1 = f_arrdiv24_fs313_not1 & f_arrdiv24_fs312_and0;
  assign f_arrdiv24_fs313_or0 = f_arrdiv24_fs313_and1 | f_arrdiv24_fs313_and0;
  assign f_arrdiv24_fs314_xor0 = f_arrdiv24_mux2to1277_xor0 ^ b[2];
  assign f_arrdiv24_fs314_not0 = ~f_arrdiv24_mux2to1277_xor0;
  assign f_arrdiv24_fs314_and0 = f_arrdiv24_fs314_not0 & b[2];
  assign f_arrdiv24_fs314_xor1 = f_arrdiv24_fs313_or0 ^ f_arrdiv24_fs314_xor0;
  assign f_arrdiv24_fs314_not1 = ~f_arrdiv24_fs314_xor0;
  assign f_arrdiv24_fs314_and1 = f_arrdiv24_fs314_not1 & f_arrdiv24_fs313_or0;
  assign f_arrdiv24_fs314_or0 = f_arrdiv24_fs314_and1 | f_arrdiv24_fs314_and0;
  assign f_arrdiv24_fs315_xor0 = f_arrdiv24_mux2to1278_xor0 ^ b[3];
  assign f_arrdiv24_fs315_not0 = ~f_arrdiv24_mux2to1278_xor0;
  assign f_arrdiv24_fs315_and0 = f_arrdiv24_fs315_not0 & b[3];
  assign f_arrdiv24_fs315_xor1 = f_arrdiv24_fs314_or0 ^ f_arrdiv24_fs315_xor0;
  assign f_arrdiv24_fs315_not1 = ~f_arrdiv24_fs315_xor0;
  assign f_arrdiv24_fs315_and1 = f_arrdiv24_fs315_not1 & f_arrdiv24_fs314_or0;
  assign f_arrdiv24_fs315_or0 = f_arrdiv24_fs315_and1 | f_arrdiv24_fs315_and0;
  assign f_arrdiv24_fs316_xor0 = f_arrdiv24_mux2to1279_xor0 ^ b[4];
  assign f_arrdiv24_fs316_not0 = ~f_arrdiv24_mux2to1279_xor0;
  assign f_arrdiv24_fs316_and0 = f_arrdiv24_fs316_not0 & b[4];
  assign f_arrdiv24_fs316_xor1 = f_arrdiv24_fs315_or0 ^ f_arrdiv24_fs316_xor0;
  assign f_arrdiv24_fs316_not1 = ~f_arrdiv24_fs316_xor0;
  assign f_arrdiv24_fs316_and1 = f_arrdiv24_fs316_not1 & f_arrdiv24_fs315_or0;
  assign f_arrdiv24_fs316_or0 = f_arrdiv24_fs316_and1 | f_arrdiv24_fs316_and0;
  assign f_arrdiv24_fs317_xor0 = f_arrdiv24_mux2to1280_xor0 ^ b[5];
  assign f_arrdiv24_fs317_not0 = ~f_arrdiv24_mux2to1280_xor0;
  assign f_arrdiv24_fs317_and0 = f_arrdiv24_fs317_not0 & b[5];
  assign f_arrdiv24_fs317_xor1 = f_arrdiv24_fs316_or0 ^ f_arrdiv24_fs317_xor0;
  assign f_arrdiv24_fs317_not1 = ~f_arrdiv24_fs317_xor0;
  assign f_arrdiv24_fs317_and1 = f_arrdiv24_fs317_not1 & f_arrdiv24_fs316_or0;
  assign f_arrdiv24_fs317_or0 = f_arrdiv24_fs317_and1 | f_arrdiv24_fs317_and0;
  assign f_arrdiv24_fs318_xor0 = f_arrdiv24_mux2to1281_xor0 ^ b[6];
  assign f_arrdiv24_fs318_not0 = ~f_arrdiv24_mux2to1281_xor0;
  assign f_arrdiv24_fs318_and0 = f_arrdiv24_fs318_not0 & b[6];
  assign f_arrdiv24_fs318_xor1 = f_arrdiv24_fs317_or0 ^ f_arrdiv24_fs318_xor0;
  assign f_arrdiv24_fs318_not1 = ~f_arrdiv24_fs318_xor0;
  assign f_arrdiv24_fs318_and1 = f_arrdiv24_fs318_not1 & f_arrdiv24_fs317_or0;
  assign f_arrdiv24_fs318_or0 = f_arrdiv24_fs318_and1 | f_arrdiv24_fs318_and0;
  assign f_arrdiv24_fs319_xor0 = f_arrdiv24_mux2to1282_xor0 ^ b[7];
  assign f_arrdiv24_fs319_not0 = ~f_arrdiv24_mux2to1282_xor0;
  assign f_arrdiv24_fs319_and0 = f_arrdiv24_fs319_not0 & b[7];
  assign f_arrdiv24_fs319_xor1 = f_arrdiv24_fs318_or0 ^ f_arrdiv24_fs319_xor0;
  assign f_arrdiv24_fs319_not1 = ~f_arrdiv24_fs319_xor0;
  assign f_arrdiv24_fs319_and1 = f_arrdiv24_fs319_not1 & f_arrdiv24_fs318_or0;
  assign f_arrdiv24_fs319_or0 = f_arrdiv24_fs319_and1 | f_arrdiv24_fs319_and0;
  assign f_arrdiv24_fs320_xor0 = f_arrdiv24_mux2to1283_xor0 ^ b[8];
  assign f_arrdiv24_fs320_not0 = ~f_arrdiv24_mux2to1283_xor0;
  assign f_arrdiv24_fs320_and0 = f_arrdiv24_fs320_not0 & b[8];
  assign f_arrdiv24_fs320_xor1 = f_arrdiv24_fs319_or0 ^ f_arrdiv24_fs320_xor0;
  assign f_arrdiv24_fs320_not1 = ~f_arrdiv24_fs320_xor0;
  assign f_arrdiv24_fs320_and1 = f_arrdiv24_fs320_not1 & f_arrdiv24_fs319_or0;
  assign f_arrdiv24_fs320_or0 = f_arrdiv24_fs320_and1 | f_arrdiv24_fs320_and0;
  assign f_arrdiv24_fs321_xor0 = f_arrdiv24_mux2to1284_xor0 ^ b[9];
  assign f_arrdiv24_fs321_not0 = ~f_arrdiv24_mux2to1284_xor0;
  assign f_arrdiv24_fs321_and0 = f_arrdiv24_fs321_not0 & b[9];
  assign f_arrdiv24_fs321_xor1 = f_arrdiv24_fs320_or0 ^ f_arrdiv24_fs321_xor0;
  assign f_arrdiv24_fs321_not1 = ~f_arrdiv24_fs321_xor0;
  assign f_arrdiv24_fs321_and1 = f_arrdiv24_fs321_not1 & f_arrdiv24_fs320_or0;
  assign f_arrdiv24_fs321_or0 = f_arrdiv24_fs321_and1 | f_arrdiv24_fs321_and0;
  assign f_arrdiv24_fs322_xor0 = f_arrdiv24_mux2to1285_xor0 ^ b[10];
  assign f_arrdiv24_fs322_not0 = ~f_arrdiv24_mux2to1285_xor0;
  assign f_arrdiv24_fs322_and0 = f_arrdiv24_fs322_not0 & b[10];
  assign f_arrdiv24_fs322_xor1 = f_arrdiv24_fs321_or0 ^ f_arrdiv24_fs322_xor0;
  assign f_arrdiv24_fs322_not1 = ~f_arrdiv24_fs322_xor0;
  assign f_arrdiv24_fs322_and1 = f_arrdiv24_fs322_not1 & f_arrdiv24_fs321_or0;
  assign f_arrdiv24_fs322_or0 = f_arrdiv24_fs322_and1 | f_arrdiv24_fs322_and0;
  assign f_arrdiv24_fs323_xor0 = f_arrdiv24_mux2to1286_xor0 ^ b[11];
  assign f_arrdiv24_fs323_not0 = ~f_arrdiv24_mux2to1286_xor0;
  assign f_arrdiv24_fs323_and0 = f_arrdiv24_fs323_not0 & b[11];
  assign f_arrdiv24_fs323_xor1 = f_arrdiv24_fs322_or0 ^ f_arrdiv24_fs323_xor0;
  assign f_arrdiv24_fs323_not1 = ~f_arrdiv24_fs323_xor0;
  assign f_arrdiv24_fs323_and1 = f_arrdiv24_fs323_not1 & f_arrdiv24_fs322_or0;
  assign f_arrdiv24_fs323_or0 = f_arrdiv24_fs323_and1 | f_arrdiv24_fs323_and0;
  assign f_arrdiv24_fs324_xor0 = f_arrdiv24_mux2to1287_xor0 ^ b[12];
  assign f_arrdiv24_fs324_not0 = ~f_arrdiv24_mux2to1287_xor0;
  assign f_arrdiv24_fs324_and0 = f_arrdiv24_fs324_not0 & b[12];
  assign f_arrdiv24_fs324_xor1 = f_arrdiv24_fs323_or0 ^ f_arrdiv24_fs324_xor0;
  assign f_arrdiv24_fs324_not1 = ~f_arrdiv24_fs324_xor0;
  assign f_arrdiv24_fs324_and1 = f_arrdiv24_fs324_not1 & f_arrdiv24_fs323_or0;
  assign f_arrdiv24_fs324_or0 = f_arrdiv24_fs324_and1 | f_arrdiv24_fs324_and0;
  assign f_arrdiv24_fs325_xor0 = f_arrdiv24_mux2to1288_xor0 ^ b[13];
  assign f_arrdiv24_fs325_not0 = ~f_arrdiv24_mux2to1288_xor0;
  assign f_arrdiv24_fs325_and0 = f_arrdiv24_fs325_not0 & b[13];
  assign f_arrdiv24_fs325_xor1 = f_arrdiv24_fs324_or0 ^ f_arrdiv24_fs325_xor0;
  assign f_arrdiv24_fs325_not1 = ~f_arrdiv24_fs325_xor0;
  assign f_arrdiv24_fs325_and1 = f_arrdiv24_fs325_not1 & f_arrdiv24_fs324_or0;
  assign f_arrdiv24_fs325_or0 = f_arrdiv24_fs325_and1 | f_arrdiv24_fs325_and0;
  assign f_arrdiv24_fs326_xor0 = f_arrdiv24_mux2to1289_xor0 ^ b[14];
  assign f_arrdiv24_fs326_not0 = ~f_arrdiv24_mux2to1289_xor0;
  assign f_arrdiv24_fs326_and0 = f_arrdiv24_fs326_not0 & b[14];
  assign f_arrdiv24_fs326_xor1 = f_arrdiv24_fs325_or0 ^ f_arrdiv24_fs326_xor0;
  assign f_arrdiv24_fs326_not1 = ~f_arrdiv24_fs326_xor0;
  assign f_arrdiv24_fs326_and1 = f_arrdiv24_fs326_not1 & f_arrdiv24_fs325_or0;
  assign f_arrdiv24_fs326_or0 = f_arrdiv24_fs326_and1 | f_arrdiv24_fs326_and0;
  assign f_arrdiv24_fs327_xor0 = f_arrdiv24_mux2to1290_xor0 ^ b[15];
  assign f_arrdiv24_fs327_not0 = ~f_arrdiv24_mux2to1290_xor0;
  assign f_arrdiv24_fs327_and0 = f_arrdiv24_fs327_not0 & b[15];
  assign f_arrdiv24_fs327_xor1 = f_arrdiv24_fs326_or0 ^ f_arrdiv24_fs327_xor0;
  assign f_arrdiv24_fs327_not1 = ~f_arrdiv24_fs327_xor0;
  assign f_arrdiv24_fs327_and1 = f_arrdiv24_fs327_not1 & f_arrdiv24_fs326_or0;
  assign f_arrdiv24_fs327_or0 = f_arrdiv24_fs327_and1 | f_arrdiv24_fs327_and0;
  assign f_arrdiv24_fs328_xor0 = f_arrdiv24_mux2to1291_xor0 ^ b[16];
  assign f_arrdiv24_fs328_not0 = ~f_arrdiv24_mux2to1291_xor0;
  assign f_arrdiv24_fs328_and0 = f_arrdiv24_fs328_not0 & b[16];
  assign f_arrdiv24_fs328_xor1 = f_arrdiv24_fs327_or0 ^ f_arrdiv24_fs328_xor0;
  assign f_arrdiv24_fs328_not1 = ~f_arrdiv24_fs328_xor0;
  assign f_arrdiv24_fs328_and1 = f_arrdiv24_fs328_not1 & f_arrdiv24_fs327_or0;
  assign f_arrdiv24_fs328_or0 = f_arrdiv24_fs328_and1 | f_arrdiv24_fs328_and0;
  assign f_arrdiv24_fs329_xor0 = f_arrdiv24_mux2to1292_xor0 ^ b[17];
  assign f_arrdiv24_fs329_not0 = ~f_arrdiv24_mux2to1292_xor0;
  assign f_arrdiv24_fs329_and0 = f_arrdiv24_fs329_not0 & b[17];
  assign f_arrdiv24_fs329_xor1 = f_arrdiv24_fs328_or0 ^ f_arrdiv24_fs329_xor0;
  assign f_arrdiv24_fs329_not1 = ~f_arrdiv24_fs329_xor0;
  assign f_arrdiv24_fs329_and1 = f_arrdiv24_fs329_not1 & f_arrdiv24_fs328_or0;
  assign f_arrdiv24_fs329_or0 = f_arrdiv24_fs329_and1 | f_arrdiv24_fs329_and0;
  assign f_arrdiv24_fs330_xor0 = f_arrdiv24_mux2to1293_xor0 ^ b[18];
  assign f_arrdiv24_fs330_not0 = ~f_arrdiv24_mux2to1293_xor0;
  assign f_arrdiv24_fs330_and0 = f_arrdiv24_fs330_not0 & b[18];
  assign f_arrdiv24_fs330_xor1 = f_arrdiv24_fs329_or0 ^ f_arrdiv24_fs330_xor0;
  assign f_arrdiv24_fs330_not1 = ~f_arrdiv24_fs330_xor0;
  assign f_arrdiv24_fs330_and1 = f_arrdiv24_fs330_not1 & f_arrdiv24_fs329_or0;
  assign f_arrdiv24_fs330_or0 = f_arrdiv24_fs330_and1 | f_arrdiv24_fs330_and0;
  assign f_arrdiv24_fs331_xor0 = f_arrdiv24_mux2to1294_xor0 ^ b[19];
  assign f_arrdiv24_fs331_not0 = ~f_arrdiv24_mux2to1294_xor0;
  assign f_arrdiv24_fs331_and0 = f_arrdiv24_fs331_not0 & b[19];
  assign f_arrdiv24_fs331_xor1 = f_arrdiv24_fs330_or0 ^ f_arrdiv24_fs331_xor0;
  assign f_arrdiv24_fs331_not1 = ~f_arrdiv24_fs331_xor0;
  assign f_arrdiv24_fs331_and1 = f_arrdiv24_fs331_not1 & f_arrdiv24_fs330_or0;
  assign f_arrdiv24_fs331_or0 = f_arrdiv24_fs331_and1 | f_arrdiv24_fs331_and0;
  assign f_arrdiv24_fs332_xor0 = f_arrdiv24_mux2to1295_xor0 ^ b[20];
  assign f_arrdiv24_fs332_not0 = ~f_arrdiv24_mux2to1295_xor0;
  assign f_arrdiv24_fs332_and0 = f_arrdiv24_fs332_not0 & b[20];
  assign f_arrdiv24_fs332_xor1 = f_arrdiv24_fs331_or0 ^ f_arrdiv24_fs332_xor0;
  assign f_arrdiv24_fs332_not1 = ~f_arrdiv24_fs332_xor0;
  assign f_arrdiv24_fs332_and1 = f_arrdiv24_fs332_not1 & f_arrdiv24_fs331_or0;
  assign f_arrdiv24_fs332_or0 = f_arrdiv24_fs332_and1 | f_arrdiv24_fs332_and0;
  assign f_arrdiv24_fs333_xor0 = f_arrdiv24_mux2to1296_xor0 ^ b[21];
  assign f_arrdiv24_fs333_not0 = ~f_arrdiv24_mux2to1296_xor0;
  assign f_arrdiv24_fs333_and0 = f_arrdiv24_fs333_not0 & b[21];
  assign f_arrdiv24_fs333_xor1 = f_arrdiv24_fs332_or0 ^ f_arrdiv24_fs333_xor0;
  assign f_arrdiv24_fs333_not1 = ~f_arrdiv24_fs333_xor0;
  assign f_arrdiv24_fs333_and1 = f_arrdiv24_fs333_not1 & f_arrdiv24_fs332_or0;
  assign f_arrdiv24_fs333_or0 = f_arrdiv24_fs333_and1 | f_arrdiv24_fs333_and0;
  assign f_arrdiv24_fs334_xor0 = f_arrdiv24_mux2to1297_xor0 ^ b[22];
  assign f_arrdiv24_fs334_not0 = ~f_arrdiv24_mux2to1297_xor0;
  assign f_arrdiv24_fs334_and0 = f_arrdiv24_fs334_not0 & b[22];
  assign f_arrdiv24_fs334_xor1 = f_arrdiv24_fs333_or0 ^ f_arrdiv24_fs334_xor0;
  assign f_arrdiv24_fs334_not1 = ~f_arrdiv24_fs334_xor0;
  assign f_arrdiv24_fs334_and1 = f_arrdiv24_fs334_not1 & f_arrdiv24_fs333_or0;
  assign f_arrdiv24_fs334_or0 = f_arrdiv24_fs334_and1 | f_arrdiv24_fs334_and0;
  assign f_arrdiv24_fs335_xor0 = f_arrdiv24_mux2to1298_xor0 ^ b[23];
  assign f_arrdiv24_fs335_not0 = ~f_arrdiv24_mux2to1298_xor0;
  assign f_arrdiv24_fs335_and0 = f_arrdiv24_fs335_not0 & b[23];
  assign f_arrdiv24_fs335_xor1 = f_arrdiv24_fs334_or0 ^ f_arrdiv24_fs335_xor0;
  assign f_arrdiv24_fs335_not1 = ~f_arrdiv24_fs335_xor0;
  assign f_arrdiv24_fs335_and1 = f_arrdiv24_fs335_not1 & f_arrdiv24_fs334_or0;
  assign f_arrdiv24_fs335_or0 = f_arrdiv24_fs335_and1 | f_arrdiv24_fs335_and0;
  assign f_arrdiv24_mux2to1299_and0 = a[10] & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1299_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1299_and1 = f_arrdiv24_fs312_xor0 & f_arrdiv24_mux2to1299_not0;
  assign f_arrdiv24_mux2to1299_xor0 = f_arrdiv24_mux2to1299_and0 ^ f_arrdiv24_mux2to1299_and1;
  assign f_arrdiv24_mux2to1300_and0 = f_arrdiv24_mux2to1276_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1300_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1300_and1 = f_arrdiv24_fs313_xor1 & f_arrdiv24_mux2to1300_not0;
  assign f_arrdiv24_mux2to1300_xor0 = f_arrdiv24_mux2to1300_and0 ^ f_arrdiv24_mux2to1300_and1;
  assign f_arrdiv24_mux2to1301_and0 = f_arrdiv24_mux2to1277_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1301_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1301_and1 = f_arrdiv24_fs314_xor1 & f_arrdiv24_mux2to1301_not0;
  assign f_arrdiv24_mux2to1301_xor0 = f_arrdiv24_mux2to1301_and0 ^ f_arrdiv24_mux2to1301_and1;
  assign f_arrdiv24_mux2to1302_and0 = f_arrdiv24_mux2to1278_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1302_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1302_and1 = f_arrdiv24_fs315_xor1 & f_arrdiv24_mux2to1302_not0;
  assign f_arrdiv24_mux2to1302_xor0 = f_arrdiv24_mux2to1302_and0 ^ f_arrdiv24_mux2to1302_and1;
  assign f_arrdiv24_mux2to1303_and0 = f_arrdiv24_mux2to1279_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1303_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1303_and1 = f_arrdiv24_fs316_xor1 & f_arrdiv24_mux2to1303_not0;
  assign f_arrdiv24_mux2to1303_xor0 = f_arrdiv24_mux2to1303_and0 ^ f_arrdiv24_mux2to1303_and1;
  assign f_arrdiv24_mux2to1304_and0 = f_arrdiv24_mux2to1280_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1304_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1304_and1 = f_arrdiv24_fs317_xor1 & f_arrdiv24_mux2to1304_not0;
  assign f_arrdiv24_mux2to1304_xor0 = f_arrdiv24_mux2to1304_and0 ^ f_arrdiv24_mux2to1304_and1;
  assign f_arrdiv24_mux2to1305_and0 = f_arrdiv24_mux2to1281_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1305_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1305_and1 = f_arrdiv24_fs318_xor1 & f_arrdiv24_mux2to1305_not0;
  assign f_arrdiv24_mux2to1305_xor0 = f_arrdiv24_mux2to1305_and0 ^ f_arrdiv24_mux2to1305_and1;
  assign f_arrdiv24_mux2to1306_and0 = f_arrdiv24_mux2to1282_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1306_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1306_and1 = f_arrdiv24_fs319_xor1 & f_arrdiv24_mux2to1306_not0;
  assign f_arrdiv24_mux2to1306_xor0 = f_arrdiv24_mux2to1306_and0 ^ f_arrdiv24_mux2to1306_and1;
  assign f_arrdiv24_mux2to1307_and0 = f_arrdiv24_mux2to1283_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1307_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1307_and1 = f_arrdiv24_fs320_xor1 & f_arrdiv24_mux2to1307_not0;
  assign f_arrdiv24_mux2to1307_xor0 = f_arrdiv24_mux2to1307_and0 ^ f_arrdiv24_mux2to1307_and1;
  assign f_arrdiv24_mux2to1308_and0 = f_arrdiv24_mux2to1284_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1308_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1308_and1 = f_arrdiv24_fs321_xor1 & f_arrdiv24_mux2to1308_not0;
  assign f_arrdiv24_mux2to1308_xor0 = f_arrdiv24_mux2to1308_and0 ^ f_arrdiv24_mux2to1308_and1;
  assign f_arrdiv24_mux2to1309_and0 = f_arrdiv24_mux2to1285_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1309_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1309_and1 = f_arrdiv24_fs322_xor1 & f_arrdiv24_mux2to1309_not0;
  assign f_arrdiv24_mux2to1309_xor0 = f_arrdiv24_mux2to1309_and0 ^ f_arrdiv24_mux2to1309_and1;
  assign f_arrdiv24_mux2to1310_and0 = f_arrdiv24_mux2to1286_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1310_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1310_and1 = f_arrdiv24_fs323_xor1 & f_arrdiv24_mux2to1310_not0;
  assign f_arrdiv24_mux2to1310_xor0 = f_arrdiv24_mux2to1310_and0 ^ f_arrdiv24_mux2to1310_and1;
  assign f_arrdiv24_mux2to1311_and0 = f_arrdiv24_mux2to1287_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1311_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1311_and1 = f_arrdiv24_fs324_xor1 & f_arrdiv24_mux2to1311_not0;
  assign f_arrdiv24_mux2to1311_xor0 = f_arrdiv24_mux2to1311_and0 ^ f_arrdiv24_mux2to1311_and1;
  assign f_arrdiv24_mux2to1312_and0 = f_arrdiv24_mux2to1288_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1312_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1312_and1 = f_arrdiv24_fs325_xor1 & f_arrdiv24_mux2to1312_not0;
  assign f_arrdiv24_mux2to1312_xor0 = f_arrdiv24_mux2to1312_and0 ^ f_arrdiv24_mux2to1312_and1;
  assign f_arrdiv24_mux2to1313_and0 = f_arrdiv24_mux2to1289_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1313_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1313_and1 = f_arrdiv24_fs326_xor1 & f_arrdiv24_mux2to1313_not0;
  assign f_arrdiv24_mux2to1313_xor0 = f_arrdiv24_mux2to1313_and0 ^ f_arrdiv24_mux2to1313_and1;
  assign f_arrdiv24_mux2to1314_and0 = f_arrdiv24_mux2to1290_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1314_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1314_and1 = f_arrdiv24_fs327_xor1 & f_arrdiv24_mux2to1314_not0;
  assign f_arrdiv24_mux2to1314_xor0 = f_arrdiv24_mux2to1314_and0 ^ f_arrdiv24_mux2to1314_and1;
  assign f_arrdiv24_mux2to1315_and0 = f_arrdiv24_mux2to1291_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1315_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1315_and1 = f_arrdiv24_fs328_xor1 & f_arrdiv24_mux2to1315_not0;
  assign f_arrdiv24_mux2to1315_xor0 = f_arrdiv24_mux2to1315_and0 ^ f_arrdiv24_mux2to1315_and1;
  assign f_arrdiv24_mux2to1316_and0 = f_arrdiv24_mux2to1292_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1316_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1316_and1 = f_arrdiv24_fs329_xor1 & f_arrdiv24_mux2to1316_not0;
  assign f_arrdiv24_mux2to1316_xor0 = f_arrdiv24_mux2to1316_and0 ^ f_arrdiv24_mux2to1316_and1;
  assign f_arrdiv24_mux2to1317_and0 = f_arrdiv24_mux2to1293_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1317_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1317_and1 = f_arrdiv24_fs330_xor1 & f_arrdiv24_mux2to1317_not0;
  assign f_arrdiv24_mux2to1317_xor0 = f_arrdiv24_mux2to1317_and0 ^ f_arrdiv24_mux2to1317_and1;
  assign f_arrdiv24_mux2to1318_and0 = f_arrdiv24_mux2to1294_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1318_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1318_and1 = f_arrdiv24_fs331_xor1 & f_arrdiv24_mux2to1318_not0;
  assign f_arrdiv24_mux2to1318_xor0 = f_arrdiv24_mux2to1318_and0 ^ f_arrdiv24_mux2to1318_and1;
  assign f_arrdiv24_mux2to1319_and0 = f_arrdiv24_mux2to1295_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1319_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1319_and1 = f_arrdiv24_fs332_xor1 & f_arrdiv24_mux2to1319_not0;
  assign f_arrdiv24_mux2to1319_xor0 = f_arrdiv24_mux2to1319_and0 ^ f_arrdiv24_mux2to1319_and1;
  assign f_arrdiv24_mux2to1320_and0 = f_arrdiv24_mux2to1296_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1320_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1320_and1 = f_arrdiv24_fs333_xor1 & f_arrdiv24_mux2to1320_not0;
  assign f_arrdiv24_mux2to1320_xor0 = f_arrdiv24_mux2to1320_and0 ^ f_arrdiv24_mux2to1320_and1;
  assign f_arrdiv24_mux2to1321_and0 = f_arrdiv24_mux2to1297_xor0 & f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1321_not0 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_mux2to1321_and1 = f_arrdiv24_fs334_xor1 & f_arrdiv24_mux2to1321_not0;
  assign f_arrdiv24_mux2to1321_xor0 = f_arrdiv24_mux2to1321_and0 ^ f_arrdiv24_mux2to1321_and1;
  assign f_arrdiv24_not13 = ~f_arrdiv24_fs335_or0;
  assign f_arrdiv24_fs336_xor0 = a[9] ^ b[0];
  assign f_arrdiv24_fs336_not0 = ~a[9];
  assign f_arrdiv24_fs336_and0 = f_arrdiv24_fs336_not0 & b[0];
  assign f_arrdiv24_fs336_not1 = ~f_arrdiv24_fs336_xor0;
  assign f_arrdiv24_fs337_xor0 = f_arrdiv24_mux2to1299_xor0 ^ b[1];
  assign f_arrdiv24_fs337_not0 = ~f_arrdiv24_mux2to1299_xor0;
  assign f_arrdiv24_fs337_and0 = f_arrdiv24_fs337_not0 & b[1];
  assign f_arrdiv24_fs337_xor1 = f_arrdiv24_fs336_and0 ^ f_arrdiv24_fs337_xor0;
  assign f_arrdiv24_fs337_not1 = ~f_arrdiv24_fs337_xor0;
  assign f_arrdiv24_fs337_and1 = f_arrdiv24_fs337_not1 & f_arrdiv24_fs336_and0;
  assign f_arrdiv24_fs337_or0 = f_arrdiv24_fs337_and1 | f_arrdiv24_fs337_and0;
  assign f_arrdiv24_fs338_xor0 = f_arrdiv24_mux2to1300_xor0 ^ b[2];
  assign f_arrdiv24_fs338_not0 = ~f_arrdiv24_mux2to1300_xor0;
  assign f_arrdiv24_fs338_and0 = f_arrdiv24_fs338_not0 & b[2];
  assign f_arrdiv24_fs338_xor1 = f_arrdiv24_fs337_or0 ^ f_arrdiv24_fs338_xor0;
  assign f_arrdiv24_fs338_not1 = ~f_arrdiv24_fs338_xor0;
  assign f_arrdiv24_fs338_and1 = f_arrdiv24_fs338_not1 & f_arrdiv24_fs337_or0;
  assign f_arrdiv24_fs338_or0 = f_arrdiv24_fs338_and1 | f_arrdiv24_fs338_and0;
  assign f_arrdiv24_fs339_xor0 = f_arrdiv24_mux2to1301_xor0 ^ b[3];
  assign f_arrdiv24_fs339_not0 = ~f_arrdiv24_mux2to1301_xor0;
  assign f_arrdiv24_fs339_and0 = f_arrdiv24_fs339_not0 & b[3];
  assign f_arrdiv24_fs339_xor1 = f_arrdiv24_fs338_or0 ^ f_arrdiv24_fs339_xor0;
  assign f_arrdiv24_fs339_not1 = ~f_arrdiv24_fs339_xor0;
  assign f_arrdiv24_fs339_and1 = f_arrdiv24_fs339_not1 & f_arrdiv24_fs338_or0;
  assign f_arrdiv24_fs339_or0 = f_arrdiv24_fs339_and1 | f_arrdiv24_fs339_and0;
  assign f_arrdiv24_fs340_xor0 = f_arrdiv24_mux2to1302_xor0 ^ b[4];
  assign f_arrdiv24_fs340_not0 = ~f_arrdiv24_mux2to1302_xor0;
  assign f_arrdiv24_fs340_and0 = f_arrdiv24_fs340_not0 & b[4];
  assign f_arrdiv24_fs340_xor1 = f_arrdiv24_fs339_or0 ^ f_arrdiv24_fs340_xor0;
  assign f_arrdiv24_fs340_not1 = ~f_arrdiv24_fs340_xor0;
  assign f_arrdiv24_fs340_and1 = f_arrdiv24_fs340_not1 & f_arrdiv24_fs339_or0;
  assign f_arrdiv24_fs340_or0 = f_arrdiv24_fs340_and1 | f_arrdiv24_fs340_and0;
  assign f_arrdiv24_fs341_xor0 = f_arrdiv24_mux2to1303_xor0 ^ b[5];
  assign f_arrdiv24_fs341_not0 = ~f_arrdiv24_mux2to1303_xor0;
  assign f_arrdiv24_fs341_and0 = f_arrdiv24_fs341_not0 & b[5];
  assign f_arrdiv24_fs341_xor1 = f_arrdiv24_fs340_or0 ^ f_arrdiv24_fs341_xor0;
  assign f_arrdiv24_fs341_not1 = ~f_arrdiv24_fs341_xor0;
  assign f_arrdiv24_fs341_and1 = f_arrdiv24_fs341_not1 & f_arrdiv24_fs340_or0;
  assign f_arrdiv24_fs341_or0 = f_arrdiv24_fs341_and1 | f_arrdiv24_fs341_and0;
  assign f_arrdiv24_fs342_xor0 = f_arrdiv24_mux2to1304_xor0 ^ b[6];
  assign f_arrdiv24_fs342_not0 = ~f_arrdiv24_mux2to1304_xor0;
  assign f_arrdiv24_fs342_and0 = f_arrdiv24_fs342_not0 & b[6];
  assign f_arrdiv24_fs342_xor1 = f_arrdiv24_fs341_or0 ^ f_arrdiv24_fs342_xor0;
  assign f_arrdiv24_fs342_not1 = ~f_arrdiv24_fs342_xor0;
  assign f_arrdiv24_fs342_and1 = f_arrdiv24_fs342_not1 & f_arrdiv24_fs341_or0;
  assign f_arrdiv24_fs342_or0 = f_arrdiv24_fs342_and1 | f_arrdiv24_fs342_and0;
  assign f_arrdiv24_fs343_xor0 = f_arrdiv24_mux2to1305_xor0 ^ b[7];
  assign f_arrdiv24_fs343_not0 = ~f_arrdiv24_mux2to1305_xor0;
  assign f_arrdiv24_fs343_and0 = f_arrdiv24_fs343_not0 & b[7];
  assign f_arrdiv24_fs343_xor1 = f_arrdiv24_fs342_or0 ^ f_arrdiv24_fs343_xor0;
  assign f_arrdiv24_fs343_not1 = ~f_arrdiv24_fs343_xor0;
  assign f_arrdiv24_fs343_and1 = f_arrdiv24_fs343_not1 & f_arrdiv24_fs342_or0;
  assign f_arrdiv24_fs343_or0 = f_arrdiv24_fs343_and1 | f_arrdiv24_fs343_and0;
  assign f_arrdiv24_fs344_xor0 = f_arrdiv24_mux2to1306_xor0 ^ b[8];
  assign f_arrdiv24_fs344_not0 = ~f_arrdiv24_mux2to1306_xor0;
  assign f_arrdiv24_fs344_and0 = f_arrdiv24_fs344_not0 & b[8];
  assign f_arrdiv24_fs344_xor1 = f_arrdiv24_fs343_or0 ^ f_arrdiv24_fs344_xor0;
  assign f_arrdiv24_fs344_not1 = ~f_arrdiv24_fs344_xor0;
  assign f_arrdiv24_fs344_and1 = f_arrdiv24_fs344_not1 & f_arrdiv24_fs343_or0;
  assign f_arrdiv24_fs344_or0 = f_arrdiv24_fs344_and1 | f_arrdiv24_fs344_and0;
  assign f_arrdiv24_fs345_xor0 = f_arrdiv24_mux2to1307_xor0 ^ b[9];
  assign f_arrdiv24_fs345_not0 = ~f_arrdiv24_mux2to1307_xor0;
  assign f_arrdiv24_fs345_and0 = f_arrdiv24_fs345_not0 & b[9];
  assign f_arrdiv24_fs345_xor1 = f_arrdiv24_fs344_or0 ^ f_arrdiv24_fs345_xor0;
  assign f_arrdiv24_fs345_not1 = ~f_arrdiv24_fs345_xor0;
  assign f_arrdiv24_fs345_and1 = f_arrdiv24_fs345_not1 & f_arrdiv24_fs344_or0;
  assign f_arrdiv24_fs345_or0 = f_arrdiv24_fs345_and1 | f_arrdiv24_fs345_and0;
  assign f_arrdiv24_fs346_xor0 = f_arrdiv24_mux2to1308_xor0 ^ b[10];
  assign f_arrdiv24_fs346_not0 = ~f_arrdiv24_mux2to1308_xor0;
  assign f_arrdiv24_fs346_and0 = f_arrdiv24_fs346_not0 & b[10];
  assign f_arrdiv24_fs346_xor1 = f_arrdiv24_fs345_or0 ^ f_arrdiv24_fs346_xor0;
  assign f_arrdiv24_fs346_not1 = ~f_arrdiv24_fs346_xor0;
  assign f_arrdiv24_fs346_and1 = f_arrdiv24_fs346_not1 & f_arrdiv24_fs345_or0;
  assign f_arrdiv24_fs346_or0 = f_arrdiv24_fs346_and1 | f_arrdiv24_fs346_and0;
  assign f_arrdiv24_fs347_xor0 = f_arrdiv24_mux2to1309_xor0 ^ b[11];
  assign f_arrdiv24_fs347_not0 = ~f_arrdiv24_mux2to1309_xor0;
  assign f_arrdiv24_fs347_and0 = f_arrdiv24_fs347_not0 & b[11];
  assign f_arrdiv24_fs347_xor1 = f_arrdiv24_fs346_or0 ^ f_arrdiv24_fs347_xor0;
  assign f_arrdiv24_fs347_not1 = ~f_arrdiv24_fs347_xor0;
  assign f_arrdiv24_fs347_and1 = f_arrdiv24_fs347_not1 & f_arrdiv24_fs346_or0;
  assign f_arrdiv24_fs347_or0 = f_arrdiv24_fs347_and1 | f_arrdiv24_fs347_and0;
  assign f_arrdiv24_fs348_xor0 = f_arrdiv24_mux2to1310_xor0 ^ b[12];
  assign f_arrdiv24_fs348_not0 = ~f_arrdiv24_mux2to1310_xor0;
  assign f_arrdiv24_fs348_and0 = f_arrdiv24_fs348_not0 & b[12];
  assign f_arrdiv24_fs348_xor1 = f_arrdiv24_fs347_or0 ^ f_arrdiv24_fs348_xor0;
  assign f_arrdiv24_fs348_not1 = ~f_arrdiv24_fs348_xor0;
  assign f_arrdiv24_fs348_and1 = f_arrdiv24_fs348_not1 & f_arrdiv24_fs347_or0;
  assign f_arrdiv24_fs348_or0 = f_arrdiv24_fs348_and1 | f_arrdiv24_fs348_and0;
  assign f_arrdiv24_fs349_xor0 = f_arrdiv24_mux2to1311_xor0 ^ b[13];
  assign f_arrdiv24_fs349_not0 = ~f_arrdiv24_mux2to1311_xor0;
  assign f_arrdiv24_fs349_and0 = f_arrdiv24_fs349_not0 & b[13];
  assign f_arrdiv24_fs349_xor1 = f_arrdiv24_fs348_or0 ^ f_arrdiv24_fs349_xor0;
  assign f_arrdiv24_fs349_not1 = ~f_arrdiv24_fs349_xor0;
  assign f_arrdiv24_fs349_and1 = f_arrdiv24_fs349_not1 & f_arrdiv24_fs348_or0;
  assign f_arrdiv24_fs349_or0 = f_arrdiv24_fs349_and1 | f_arrdiv24_fs349_and0;
  assign f_arrdiv24_fs350_xor0 = f_arrdiv24_mux2to1312_xor0 ^ b[14];
  assign f_arrdiv24_fs350_not0 = ~f_arrdiv24_mux2to1312_xor0;
  assign f_arrdiv24_fs350_and0 = f_arrdiv24_fs350_not0 & b[14];
  assign f_arrdiv24_fs350_xor1 = f_arrdiv24_fs349_or0 ^ f_arrdiv24_fs350_xor0;
  assign f_arrdiv24_fs350_not1 = ~f_arrdiv24_fs350_xor0;
  assign f_arrdiv24_fs350_and1 = f_arrdiv24_fs350_not1 & f_arrdiv24_fs349_or0;
  assign f_arrdiv24_fs350_or0 = f_arrdiv24_fs350_and1 | f_arrdiv24_fs350_and0;
  assign f_arrdiv24_fs351_xor0 = f_arrdiv24_mux2to1313_xor0 ^ b[15];
  assign f_arrdiv24_fs351_not0 = ~f_arrdiv24_mux2to1313_xor0;
  assign f_arrdiv24_fs351_and0 = f_arrdiv24_fs351_not0 & b[15];
  assign f_arrdiv24_fs351_xor1 = f_arrdiv24_fs350_or0 ^ f_arrdiv24_fs351_xor0;
  assign f_arrdiv24_fs351_not1 = ~f_arrdiv24_fs351_xor0;
  assign f_arrdiv24_fs351_and1 = f_arrdiv24_fs351_not1 & f_arrdiv24_fs350_or0;
  assign f_arrdiv24_fs351_or0 = f_arrdiv24_fs351_and1 | f_arrdiv24_fs351_and0;
  assign f_arrdiv24_fs352_xor0 = f_arrdiv24_mux2to1314_xor0 ^ b[16];
  assign f_arrdiv24_fs352_not0 = ~f_arrdiv24_mux2to1314_xor0;
  assign f_arrdiv24_fs352_and0 = f_arrdiv24_fs352_not0 & b[16];
  assign f_arrdiv24_fs352_xor1 = f_arrdiv24_fs351_or0 ^ f_arrdiv24_fs352_xor0;
  assign f_arrdiv24_fs352_not1 = ~f_arrdiv24_fs352_xor0;
  assign f_arrdiv24_fs352_and1 = f_arrdiv24_fs352_not1 & f_arrdiv24_fs351_or0;
  assign f_arrdiv24_fs352_or0 = f_arrdiv24_fs352_and1 | f_arrdiv24_fs352_and0;
  assign f_arrdiv24_fs353_xor0 = f_arrdiv24_mux2to1315_xor0 ^ b[17];
  assign f_arrdiv24_fs353_not0 = ~f_arrdiv24_mux2to1315_xor0;
  assign f_arrdiv24_fs353_and0 = f_arrdiv24_fs353_not0 & b[17];
  assign f_arrdiv24_fs353_xor1 = f_arrdiv24_fs352_or0 ^ f_arrdiv24_fs353_xor0;
  assign f_arrdiv24_fs353_not1 = ~f_arrdiv24_fs353_xor0;
  assign f_arrdiv24_fs353_and1 = f_arrdiv24_fs353_not1 & f_arrdiv24_fs352_or0;
  assign f_arrdiv24_fs353_or0 = f_arrdiv24_fs353_and1 | f_arrdiv24_fs353_and0;
  assign f_arrdiv24_fs354_xor0 = f_arrdiv24_mux2to1316_xor0 ^ b[18];
  assign f_arrdiv24_fs354_not0 = ~f_arrdiv24_mux2to1316_xor0;
  assign f_arrdiv24_fs354_and0 = f_arrdiv24_fs354_not0 & b[18];
  assign f_arrdiv24_fs354_xor1 = f_arrdiv24_fs353_or0 ^ f_arrdiv24_fs354_xor0;
  assign f_arrdiv24_fs354_not1 = ~f_arrdiv24_fs354_xor0;
  assign f_arrdiv24_fs354_and1 = f_arrdiv24_fs354_not1 & f_arrdiv24_fs353_or0;
  assign f_arrdiv24_fs354_or0 = f_arrdiv24_fs354_and1 | f_arrdiv24_fs354_and0;
  assign f_arrdiv24_fs355_xor0 = f_arrdiv24_mux2to1317_xor0 ^ b[19];
  assign f_arrdiv24_fs355_not0 = ~f_arrdiv24_mux2to1317_xor0;
  assign f_arrdiv24_fs355_and0 = f_arrdiv24_fs355_not0 & b[19];
  assign f_arrdiv24_fs355_xor1 = f_arrdiv24_fs354_or0 ^ f_arrdiv24_fs355_xor0;
  assign f_arrdiv24_fs355_not1 = ~f_arrdiv24_fs355_xor0;
  assign f_arrdiv24_fs355_and1 = f_arrdiv24_fs355_not1 & f_arrdiv24_fs354_or0;
  assign f_arrdiv24_fs355_or0 = f_arrdiv24_fs355_and1 | f_arrdiv24_fs355_and0;
  assign f_arrdiv24_fs356_xor0 = f_arrdiv24_mux2to1318_xor0 ^ b[20];
  assign f_arrdiv24_fs356_not0 = ~f_arrdiv24_mux2to1318_xor0;
  assign f_arrdiv24_fs356_and0 = f_arrdiv24_fs356_not0 & b[20];
  assign f_arrdiv24_fs356_xor1 = f_arrdiv24_fs355_or0 ^ f_arrdiv24_fs356_xor0;
  assign f_arrdiv24_fs356_not1 = ~f_arrdiv24_fs356_xor0;
  assign f_arrdiv24_fs356_and1 = f_arrdiv24_fs356_not1 & f_arrdiv24_fs355_or0;
  assign f_arrdiv24_fs356_or0 = f_arrdiv24_fs356_and1 | f_arrdiv24_fs356_and0;
  assign f_arrdiv24_fs357_xor0 = f_arrdiv24_mux2to1319_xor0 ^ b[21];
  assign f_arrdiv24_fs357_not0 = ~f_arrdiv24_mux2to1319_xor0;
  assign f_arrdiv24_fs357_and0 = f_arrdiv24_fs357_not0 & b[21];
  assign f_arrdiv24_fs357_xor1 = f_arrdiv24_fs356_or0 ^ f_arrdiv24_fs357_xor0;
  assign f_arrdiv24_fs357_not1 = ~f_arrdiv24_fs357_xor0;
  assign f_arrdiv24_fs357_and1 = f_arrdiv24_fs357_not1 & f_arrdiv24_fs356_or0;
  assign f_arrdiv24_fs357_or0 = f_arrdiv24_fs357_and1 | f_arrdiv24_fs357_and0;
  assign f_arrdiv24_fs358_xor0 = f_arrdiv24_mux2to1320_xor0 ^ b[22];
  assign f_arrdiv24_fs358_not0 = ~f_arrdiv24_mux2to1320_xor0;
  assign f_arrdiv24_fs358_and0 = f_arrdiv24_fs358_not0 & b[22];
  assign f_arrdiv24_fs358_xor1 = f_arrdiv24_fs357_or0 ^ f_arrdiv24_fs358_xor0;
  assign f_arrdiv24_fs358_not1 = ~f_arrdiv24_fs358_xor0;
  assign f_arrdiv24_fs358_and1 = f_arrdiv24_fs358_not1 & f_arrdiv24_fs357_or0;
  assign f_arrdiv24_fs358_or0 = f_arrdiv24_fs358_and1 | f_arrdiv24_fs358_and0;
  assign f_arrdiv24_fs359_xor0 = f_arrdiv24_mux2to1321_xor0 ^ b[23];
  assign f_arrdiv24_fs359_not0 = ~f_arrdiv24_mux2to1321_xor0;
  assign f_arrdiv24_fs359_and0 = f_arrdiv24_fs359_not0 & b[23];
  assign f_arrdiv24_fs359_xor1 = f_arrdiv24_fs358_or0 ^ f_arrdiv24_fs359_xor0;
  assign f_arrdiv24_fs359_not1 = ~f_arrdiv24_fs359_xor0;
  assign f_arrdiv24_fs359_and1 = f_arrdiv24_fs359_not1 & f_arrdiv24_fs358_or0;
  assign f_arrdiv24_fs359_or0 = f_arrdiv24_fs359_and1 | f_arrdiv24_fs359_and0;
  assign f_arrdiv24_mux2to1322_and0 = a[9] & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1322_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1322_and1 = f_arrdiv24_fs336_xor0 & f_arrdiv24_mux2to1322_not0;
  assign f_arrdiv24_mux2to1322_xor0 = f_arrdiv24_mux2to1322_and0 ^ f_arrdiv24_mux2to1322_and1;
  assign f_arrdiv24_mux2to1323_and0 = f_arrdiv24_mux2to1299_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1323_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1323_and1 = f_arrdiv24_fs337_xor1 & f_arrdiv24_mux2to1323_not0;
  assign f_arrdiv24_mux2to1323_xor0 = f_arrdiv24_mux2to1323_and0 ^ f_arrdiv24_mux2to1323_and1;
  assign f_arrdiv24_mux2to1324_and0 = f_arrdiv24_mux2to1300_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1324_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1324_and1 = f_arrdiv24_fs338_xor1 & f_arrdiv24_mux2to1324_not0;
  assign f_arrdiv24_mux2to1324_xor0 = f_arrdiv24_mux2to1324_and0 ^ f_arrdiv24_mux2to1324_and1;
  assign f_arrdiv24_mux2to1325_and0 = f_arrdiv24_mux2to1301_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1325_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1325_and1 = f_arrdiv24_fs339_xor1 & f_arrdiv24_mux2to1325_not0;
  assign f_arrdiv24_mux2to1325_xor0 = f_arrdiv24_mux2to1325_and0 ^ f_arrdiv24_mux2to1325_and1;
  assign f_arrdiv24_mux2to1326_and0 = f_arrdiv24_mux2to1302_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1326_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1326_and1 = f_arrdiv24_fs340_xor1 & f_arrdiv24_mux2to1326_not0;
  assign f_arrdiv24_mux2to1326_xor0 = f_arrdiv24_mux2to1326_and0 ^ f_arrdiv24_mux2to1326_and1;
  assign f_arrdiv24_mux2to1327_and0 = f_arrdiv24_mux2to1303_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1327_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1327_and1 = f_arrdiv24_fs341_xor1 & f_arrdiv24_mux2to1327_not0;
  assign f_arrdiv24_mux2to1327_xor0 = f_arrdiv24_mux2to1327_and0 ^ f_arrdiv24_mux2to1327_and1;
  assign f_arrdiv24_mux2to1328_and0 = f_arrdiv24_mux2to1304_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1328_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1328_and1 = f_arrdiv24_fs342_xor1 & f_arrdiv24_mux2to1328_not0;
  assign f_arrdiv24_mux2to1328_xor0 = f_arrdiv24_mux2to1328_and0 ^ f_arrdiv24_mux2to1328_and1;
  assign f_arrdiv24_mux2to1329_and0 = f_arrdiv24_mux2to1305_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1329_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1329_and1 = f_arrdiv24_fs343_xor1 & f_arrdiv24_mux2to1329_not0;
  assign f_arrdiv24_mux2to1329_xor0 = f_arrdiv24_mux2to1329_and0 ^ f_arrdiv24_mux2to1329_and1;
  assign f_arrdiv24_mux2to1330_and0 = f_arrdiv24_mux2to1306_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1330_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1330_and1 = f_arrdiv24_fs344_xor1 & f_arrdiv24_mux2to1330_not0;
  assign f_arrdiv24_mux2to1330_xor0 = f_arrdiv24_mux2to1330_and0 ^ f_arrdiv24_mux2to1330_and1;
  assign f_arrdiv24_mux2to1331_and0 = f_arrdiv24_mux2to1307_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1331_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1331_and1 = f_arrdiv24_fs345_xor1 & f_arrdiv24_mux2to1331_not0;
  assign f_arrdiv24_mux2to1331_xor0 = f_arrdiv24_mux2to1331_and0 ^ f_arrdiv24_mux2to1331_and1;
  assign f_arrdiv24_mux2to1332_and0 = f_arrdiv24_mux2to1308_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1332_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1332_and1 = f_arrdiv24_fs346_xor1 & f_arrdiv24_mux2to1332_not0;
  assign f_arrdiv24_mux2to1332_xor0 = f_arrdiv24_mux2to1332_and0 ^ f_arrdiv24_mux2to1332_and1;
  assign f_arrdiv24_mux2to1333_and0 = f_arrdiv24_mux2to1309_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1333_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1333_and1 = f_arrdiv24_fs347_xor1 & f_arrdiv24_mux2to1333_not0;
  assign f_arrdiv24_mux2to1333_xor0 = f_arrdiv24_mux2to1333_and0 ^ f_arrdiv24_mux2to1333_and1;
  assign f_arrdiv24_mux2to1334_and0 = f_arrdiv24_mux2to1310_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1334_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1334_and1 = f_arrdiv24_fs348_xor1 & f_arrdiv24_mux2to1334_not0;
  assign f_arrdiv24_mux2to1334_xor0 = f_arrdiv24_mux2to1334_and0 ^ f_arrdiv24_mux2to1334_and1;
  assign f_arrdiv24_mux2to1335_and0 = f_arrdiv24_mux2to1311_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1335_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1335_and1 = f_arrdiv24_fs349_xor1 & f_arrdiv24_mux2to1335_not0;
  assign f_arrdiv24_mux2to1335_xor0 = f_arrdiv24_mux2to1335_and0 ^ f_arrdiv24_mux2to1335_and1;
  assign f_arrdiv24_mux2to1336_and0 = f_arrdiv24_mux2to1312_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1336_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1336_and1 = f_arrdiv24_fs350_xor1 & f_arrdiv24_mux2to1336_not0;
  assign f_arrdiv24_mux2to1336_xor0 = f_arrdiv24_mux2to1336_and0 ^ f_arrdiv24_mux2to1336_and1;
  assign f_arrdiv24_mux2to1337_and0 = f_arrdiv24_mux2to1313_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1337_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1337_and1 = f_arrdiv24_fs351_xor1 & f_arrdiv24_mux2to1337_not0;
  assign f_arrdiv24_mux2to1337_xor0 = f_arrdiv24_mux2to1337_and0 ^ f_arrdiv24_mux2to1337_and1;
  assign f_arrdiv24_mux2to1338_and0 = f_arrdiv24_mux2to1314_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1338_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1338_and1 = f_arrdiv24_fs352_xor1 & f_arrdiv24_mux2to1338_not0;
  assign f_arrdiv24_mux2to1338_xor0 = f_arrdiv24_mux2to1338_and0 ^ f_arrdiv24_mux2to1338_and1;
  assign f_arrdiv24_mux2to1339_and0 = f_arrdiv24_mux2to1315_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1339_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1339_and1 = f_arrdiv24_fs353_xor1 & f_arrdiv24_mux2to1339_not0;
  assign f_arrdiv24_mux2to1339_xor0 = f_arrdiv24_mux2to1339_and0 ^ f_arrdiv24_mux2to1339_and1;
  assign f_arrdiv24_mux2to1340_and0 = f_arrdiv24_mux2to1316_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1340_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1340_and1 = f_arrdiv24_fs354_xor1 & f_arrdiv24_mux2to1340_not0;
  assign f_arrdiv24_mux2to1340_xor0 = f_arrdiv24_mux2to1340_and0 ^ f_arrdiv24_mux2to1340_and1;
  assign f_arrdiv24_mux2to1341_and0 = f_arrdiv24_mux2to1317_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1341_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1341_and1 = f_arrdiv24_fs355_xor1 & f_arrdiv24_mux2to1341_not0;
  assign f_arrdiv24_mux2to1341_xor0 = f_arrdiv24_mux2to1341_and0 ^ f_arrdiv24_mux2to1341_and1;
  assign f_arrdiv24_mux2to1342_and0 = f_arrdiv24_mux2to1318_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1342_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1342_and1 = f_arrdiv24_fs356_xor1 & f_arrdiv24_mux2to1342_not0;
  assign f_arrdiv24_mux2to1342_xor0 = f_arrdiv24_mux2to1342_and0 ^ f_arrdiv24_mux2to1342_and1;
  assign f_arrdiv24_mux2to1343_and0 = f_arrdiv24_mux2to1319_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1343_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1343_and1 = f_arrdiv24_fs357_xor1 & f_arrdiv24_mux2to1343_not0;
  assign f_arrdiv24_mux2to1343_xor0 = f_arrdiv24_mux2to1343_and0 ^ f_arrdiv24_mux2to1343_and1;
  assign f_arrdiv24_mux2to1344_and0 = f_arrdiv24_mux2to1320_xor0 & f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1344_not0 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_mux2to1344_and1 = f_arrdiv24_fs358_xor1 & f_arrdiv24_mux2to1344_not0;
  assign f_arrdiv24_mux2to1344_xor0 = f_arrdiv24_mux2to1344_and0 ^ f_arrdiv24_mux2to1344_and1;
  assign f_arrdiv24_not14 = ~f_arrdiv24_fs359_or0;
  assign f_arrdiv24_fs360_xor0 = a[8] ^ b[0];
  assign f_arrdiv24_fs360_not0 = ~a[8];
  assign f_arrdiv24_fs360_and0 = f_arrdiv24_fs360_not0 & b[0];
  assign f_arrdiv24_fs360_not1 = ~f_arrdiv24_fs360_xor0;
  assign f_arrdiv24_fs361_xor0 = f_arrdiv24_mux2to1322_xor0 ^ b[1];
  assign f_arrdiv24_fs361_not0 = ~f_arrdiv24_mux2to1322_xor0;
  assign f_arrdiv24_fs361_and0 = f_arrdiv24_fs361_not0 & b[1];
  assign f_arrdiv24_fs361_xor1 = f_arrdiv24_fs360_and0 ^ f_arrdiv24_fs361_xor0;
  assign f_arrdiv24_fs361_not1 = ~f_arrdiv24_fs361_xor0;
  assign f_arrdiv24_fs361_and1 = f_arrdiv24_fs361_not1 & f_arrdiv24_fs360_and0;
  assign f_arrdiv24_fs361_or0 = f_arrdiv24_fs361_and1 | f_arrdiv24_fs361_and0;
  assign f_arrdiv24_fs362_xor0 = f_arrdiv24_mux2to1323_xor0 ^ b[2];
  assign f_arrdiv24_fs362_not0 = ~f_arrdiv24_mux2to1323_xor0;
  assign f_arrdiv24_fs362_and0 = f_arrdiv24_fs362_not0 & b[2];
  assign f_arrdiv24_fs362_xor1 = f_arrdiv24_fs361_or0 ^ f_arrdiv24_fs362_xor0;
  assign f_arrdiv24_fs362_not1 = ~f_arrdiv24_fs362_xor0;
  assign f_arrdiv24_fs362_and1 = f_arrdiv24_fs362_not1 & f_arrdiv24_fs361_or0;
  assign f_arrdiv24_fs362_or0 = f_arrdiv24_fs362_and1 | f_arrdiv24_fs362_and0;
  assign f_arrdiv24_fs363_xor0 = f_arrdiv24_mux2to1324_xor0 ^ b[3];
  assign f_arrdiv24_fs363_not0 = ~f_arrdiv24_mux2to1324_xor0;
  assign f_arrdiv24_fs363_and0 = f_arrdiv24_fs363_not0 & b[3];
  assign f_arrdiv24_fs363_xor1 = f_arrdiv24_fs362_or0 ^ f_arrdiv24_fs363_xor0;
  assign f_arrdiv24_fs363_not1 = ~f_arrdiv24_fs363_xor0;
  assign f_arrdiv24_fs363_and1 = f_arrdiv24_fs363_not1 & f_arrdiv24_fs362_or0;
  assign f_arrdiv24_fs363_or0 = f_arrdiv24_fs363_and1 | f_arrdiv24_fs363_and0;
  assign f_arrdiv24_fs364_xor0 = f_arrdiv24_mux2to1325_xor0 ^ b[4];
  assign f_arrdiv24_fs364_not0 = ~f_arrdiv24_mux2to1325_xor0;
  assign f_arrdiv24_fs364_and0 = f_arrdiv24_fs364_not0 & b[4];
  assign f_arrdiv24_fs364_xor1 = f_arrdiv24_fs363_or0 ^ f_arrdiv24_fs364_xor0;
  assign f_arrdiv24_fs364_not1 = ~f_arrdiv24_fs364_xor0;
  assign f_arrdiv24_fs364_and1 = f_arrdiv24_fs364_not1 & f_arrdiv24_fs363_or0;
  assign f_arrdiv24_fs364_or0 = f_arrdiv24_fs364_and1 | f_arrdiv24_fs364_and0;
  assign f_arrdiv24_fs365_xor0 = f_arrdiv24_mux2to1326_xor0 ^ b[5];
  assign f_arrdiv24_fs365_not0 = ~f_arrdiv24_mux2to1326_xor0;
  assign f_arrdiv24_fs365_and0 = f_arrdiv24_fs365_not0 & b[5];
  assign f_arrdiv24_fs365_xor1 = f_arrdiv24_fs364_or0 ^ f_arrdiv24_fs365_xor0;
  assign f_arrdiv24_fs365_not1 = ~f_arrdiv24_fs365_xor0;
  assign f_arrdiv24_fs365_and1 = f_arrdiv24_fs365_not1 & f_arrdiv24_fs364_or0;
  assign f_arrdiv24_fs365_or0 = f_arrdiv24_fs365_and1 | f_arrdiv24_fs365_and0;
  assign f_arrdiv24_fs366_xor0 = f_arrdiv24_mux2to1327_xor0 ^ b[6];
  assign f_arrdiv24_fs366_not0 = ~f_arrdiv24_mux2to1327_xor0;
  assign f_arrdiv24_fs366_and0 = f_arrdiv24_fs366_not0 & b[6];
  assign f_arrdiv24_fs366_xor1 = f_arrdiv24_fs365_or0 ^ f_arrdiv24_fs366_xor0;
  assign f_arrdiv24_fs366_not1 = ~f_arrdiv24_fs366_xor0;
  assign f_arrdiv24_fs366_and1 = f_arrdiv24_fs366_not1 & f_arrdiv24_fs365_or0;
  assign f_arrdiv24_fs366_or0 = f_arrdiv24_fs366_and1 | f_arrdiv24_fs366_and0;
  assign f_arrdiv24_fs367_xor0 = f_arrdiv24_mux2to1328_xor0 ^ b[7];
  assign f_arrdiv24_fs367_not0 = ~f_arrdiv24_mux2to1328_xor0;
  assign f_arrdiv24_fs367_and0 = f_arrdiv24_fs367_not0 & b[7];
  assign f_arrdiv24_fs367_xor1 = f_arrdiv24_fs366_or0 ^ f_arrdiv24_fs367_xor0;
  assign f_arrdiv24_fs367_not1 = ~f_arrdiv24_fs367_xor0;
  assign f_arrdiv24_fs367_and1 = f_arrdiv24_fs367_not1 & f_arrdiv24_fs366_or0;
  assign f_arrdiv24_fs367_or0 = f_arrdiv24_fs367_and1 | f_arrdiv24_fs367_and0;
  assign f_arrdiv24_fs368_xor0 = f_arrdiv24_mux2to1329_xor0 ^ b[8];
  assign f_arrdiv24_fs368_not0 = ~f_arrdiv24_mux2to1329_xor0;
  assign f_arrdiv24_fs368_and0 = f_arrdiv24_fs368_not0 & b[8];
  assign f_arrdiv24_fs368_xor1 = f_arrdiv24_fs367_or0 ^ f_arrdiv24_fs368_xor0;
  assign f_arrdiv24_fs368_not1 = ~f_arrdiv24_fs368_xor0;
  assign f_arrdiv24_fs368_and1 = f_arrdiv24_fs368_not1 & f_arrdiv24_fs367_or0;
  assign f_arrdiv24_fs368_or0 = f_arrdiv24_fs368_and1 | f_arrdiv24_fs368_and0;
  assign f_arrdiv24_fs369_xor0 = f_arrdiv24_mux2to1330_xor0 ^ b[9];
  assign f_arrdiv24_fs369_not0 = ~f_arrdiv24_mux2to1330_xor0;
  assign f_arrdiv24_fs369_and0 = f_arrdiv24_fs369_not0 & b[9];
  assign f_arrdiv24_fs369_xor1 = f_arrdiv24_fs368_or0 ^ f_arrdiv24_fs369_xor0;
  assign f_arrdiv24_fs369_not1 = ~f_arrdiv24_fs369_xor0;
  assign f_arrdiv24_fs369_and1 = f_arrdiv24_fs369_not1 & f_arrdiv24_fs368_or0;
  assign f_arrdiv24_fs369_or0 = f_arrdiv24_fs369_and1 | f_arrdiv24_fs369_and0;
  assign f_arrdiv24_fs370_xor0 = f_arrdiv24_mux2to1331_xor0 ^ b[10];
  assign f_arrdiv24_fs370_not0 = ~f_arrdiv24_mux2to1331_xor0;
  assign f_arrdiv24_fs370_and0 = f_arrdiv24_fs370_not0 & b[10];
  assign f_arrdiv24_fs370_xor1 = f_arrdiv24_fs369_or0 ^ f_arrdiv24_fs370_xor0;
  assign f_arrdiv24_fs370_not1 = ~f_arrdiv24_fs370_xor0;
  assign f_arrdiv24_fs370_and1 = f_arrdiv24_fs370_not1 & f_arrdiv24_fs369_or0;
  assign f_arrdiv24_fs370_or0 = f_arrdiv24_fs370_and1 | f_arrdiv24_fs370_and0;
  assign f_arrdiv24_fs371_xor0 = f_arrdiv24_mux2to1332_xor0 ^ b[11];
  assign f_arrdiv24_fs371_not0 = ~f_arrdiv24_mux2to1332_xor0;
  assign f_arrdiv24_fs371_and0 = f_arrdiv24_fs371_not0 & b[11];
  assign f_arrdiv24_fs371_xor1 = f_arrdiv24_fs370_or0 ^ f_arrdiv24_fs371_xor0;
  assign f_arrdiv24_fs371_not1 = ~f_arrdiv24_fs371_xor0;
  assign f_arrdiv24_fs371_and1 = f_arrdiv24_fs371_not1 & f_arrdiv24_fs370_or0;
  assign f_arrdiv24_fs371_or0 = f_arrdiv24_fs371_and1 | f_arrdiv24_fs371_and0;
  assign f_arrdiv24_fs372_xor0 = f_arrdiv24_mux2to1333_xor0 ^ b[12];
  assign f_arrdiv24_fs372_not0 = ~f_arrdiv24_mux2to1333_xor0;
  assign f_arrdiv24_fs372_and0 = f_arrdiv24_fs372_not0 & b[12];
  assign f_arrdiv24_fs372_xor1 = f_arrdiv24_fs371_or0 ^ f_arrdiv24_fs372_xor0;
  assign f_arrdiv24_fs372_not1 = ~f_arrdiv24_fs372_xor0;
  assign f_arrdiv24_fs372_and1 = f_arrdiv24_fs372_not1 & f_arrdiv24_fs371_or0;
  assign f_arrdiv24_fs372_or0 = f_arrdiv24_fs372_and1 | f_arrdiv24_fs372_and0;
  assign f_arrdiv24_fs373_xor0 = f_arrdiv24_mux2to1334_xor0 ^ b[13];
  assign f_arrdiv24_fs373_not0 = ~f_arrdiv24_mux2to1334_xor0;
  assign f_arrdiv24_fs373_and0 = f_arrdiv24_fs373_not0 & b[13];
  assign f_arrdiv24_fs373_xor1 = f_arrdiv24_fs372_or0 ^ f_arrdiv24_fs373_xor0;
  assign f_arrdiv24_fs373_not1 = ~f_arrdiv24_fs373_xor0;
  assign f_arrdiv24_fs373_and1 = f_arrdiv24_fs373_not1 & f_arrdiv24_fs372_or0;
  assign f_arrdiv24_fs373_or0 = f_arrdiv24_fs373_and1 | f_arrdiv24_fs373_and0;
  assign f_arrdiv24_fs374_xor0 = f_arrdiv24_mux2to1335_xor0 ^ b[14];
  assign f_arrdiv24_fs374_not0 = ~f_arrdiv24_mux2to1335_xor0;
  assign f_arrdiv24_fs374_and0 = f_arrdiv24_fs374_not0 & b[14];
  assign f_arrdiv24_fs374_xor1 = f_arrdiv24_fs373_or0 ^ f_arrdiv24_fs374_xor0;
  assign f_arrdiv24_fs374_not1 = ~f_arrdiv24_fs374_xor0;
  assign f_arrdiv24_fs374_and1 = f_arrdiv24_fs374_not1 & f_arrdiv24_fs373_or0;
  assign f_arrdiv24_fs374_or0 = f_arrdiv24_fs374_and1 | f_arrdiv24_fs374_and0;
  assign f_arrdiv24_fs375_xor0 = f_arrdiv24_mux2to1336_xor0 ^ b[15];
  assign f_arrdiv24_fs375_not0 = ~f_arrdiv24_mux2to1336_xor0;
  assign f_arrdiv24_fs375_and0 = f_arrdiv24_fs375_not0 & b[15];
  assign f_arrdiv24_fs375_xor1 = f_arrdiv24_fs374_or0 ^ f_arrdiv24_fs375_xor0;
  assign f_arrdiv24_fs375_not1 = ~f_arrdiv24_fs375_xor0;
  assign f_arrdiv24_fs375_and1 = f_arrdiv24_fs375_not1 & f_arrdiv24_fs374_or0;
  assign f_arrdiv24_fs375_or0 = f_arrdiv24_fs375_and1 | f_arrdiv24_fs375_and0;
  assign f_arrdiv24_fs376_xor0 = f_arrdiv24_mux2to1337_xor0 ^ b[16];
  assign f_arrdiv24_fs376_not0 = ~f_arrdiv24_mux2to1337_xor0;
  assign f_arrdiv24_fs376_and0 = f_arrdiv24_fs376_not0 & b[16];
  assign f_arrdiv24_fs376_xor1 = f_arrdiv24_fs375_or0 ^ f_arrdiv24_fs376_xor0;
  assign f_arrdiv24_fs376_not1 = ~f_arrdiv24_fs376_xor0;
  assign f_arrdiv24_fs376_and1 = f_arrdiv24_fs376_not1 & f_arrdiv24_fs375_or0;
  assign f_arrdiv24_fs376_or0 = f_arrdiv24_fs376_and1 | f_arrdiv24_fs376_and0;
  assign f_arrdiv24_fs377_xor0 = f_arrdiv24_mux2to1338_xor0 ^ b[17];
  assign f_arrdiv24_fs377_not0 = ~f_arrdiv24_mux2to1338_xor0;
  assign f_arrdiv24_fs377_and0 = f_arrdiv24_fs377_not0 & b[17];
  assign f_arrdiv24_fs377_xor1 = f_arrdiv24_fs376_or0 ^ f_arrdiv24_fs377_xor0;
  assign f_arrdiv24_fs377_not1 = ~f_arrdiv24_fs377_xor0;
  assign f_arrdiv24_fs377_and1 = f_arrdiv24_fs377_not1 & f_arrdiv24_fs376_or0;
  assign f_arrdiv24_fs377_or0 = f_arrdiv24_fs377_and1 | f_arrdiv24_fs377_and0;
  assign f_arrdiv24_fs378_xor0 = f_arrdiv24_mux2to1339_xor0 ^ b[18];
  assign f_arrdiv24_fs378_not0 = ~f_arrdiv24_mux2to1339_xor0;
  assign f_arrdiv24_fs378_and0 = f_arrdiv24_fs378_not0 & b[18];
  assign f_arrdiv24_fs378_xor1 = f_arrdiv24_fs377_or0 ^ f_arrdiv24_fs378_xor0;
  assign f_arrdiv24_fs378_not1 = ~f_arrdiv24_fs378_xor0;
  assign f_arrdiv24_fs378_and1 = f_arrdiv24_fs378_not1 & f_arrdiv24_fs377_or0;
  assign f_arrdiv24_fs378_or0 = f_arrdiv24_fs378_and1 | f_arrdiv24_fs378_and0;
  assign f_arrdiv24_fs379_xor0 = f_arrdiv24_mux2to1340_xor0 ^ b[19];
  assign f_arrdiv24_fs379_not0 = ~f_arrdiv24_mux2to1340_xor0;
  assign f_arrdiv24_fs379_and0 = f_arrdiv24_fs379_not0 & b[19];
  assign f_arrdiv24_fs379_xor1 = f_arrdiv24_fs378_or0 ^ f_arrdiv24_fs379_xor0;
  assign f_arrdiv24_fs379_not1 = ~f_arrdiv24_fs379_xor0;
  assign f_arrdiv24_fs379_and1 = f_arrdiv24_fs379_not1 & f_arrdiv24_fs378_or0;
  assign f_arrdiv24_fs379_or0 = f_arrdiv24_fs379_and1 | f_arrdiv24_fs379_and0;
  assign f_arrdiv24_fs380_xor0 = f_arrdiv24_mux2to1341_xor0 ^ b[20];
  assign f_arrdiv24_fs380_not0 = ~f_arrdiv24_mux2to1341_xor0;
  assign f_arrdiv24_fs380_and0 = f_arrdiv24_fs380_not0 & b[20];
  assign f_arrdiv24_fs380_xor1 = f_arrdiv24_fs379_or0 ^ f_arrdiv24_fs380_xor0;
  assign f_arrdiv24_fs380_not1 = ~f_arrdiv24_fs380_xor0;
  assign f_arrdiv24_fs380_and1 = f_arrdiv24_fs380_not1 & f_arrdiv24_fs379_or0;
  assign f_arrdiv24_fs380_or0 = f_arrdiv24_fs380_and1 | f_arrdiv24_fs380_and0;
  assign f_arrdiv24_fs381_xor0 = f_arrdiv24_mux2to1342_xor0 ^ b[21];
  assign f_arrdiv24_fs381_not0 = ~f_arrdiv24_mux2to1342_xor0;
  assign f_arrdiv24_fs381_and0 = f_arrdiv24_fs381_not0 & b[21];
  assign f_arrdiv24_fs381_xor1 = f_arrdiv24_fs380_or0 ^ f_arrdiv24_fs381_xor0;
  assign f_arrdiv24_fs381_not1 = ~f_arrdiv24_fs381_xor0;
  assign f_arrdiv24_fs381_and1 = f_arrdiv24_fs381_not1 & f_arrdiv24_fs380_or0;
  assign f_arrdiv24_fs381_or0 = f_arrdiv24_fs381_and1 | f_arrdiv24_fs381_and0;
  assign f_arrdiv24_fs382_xor0 = f_arrdiv24_mux2to1343_xor0 ^ b[22];
  assign f_arrdiv24_fs382_not0 = ~f_arrdiv24_mux2to1343_xor0;
  assign f_arrdiv24_fs382_and0 = f_arrdiv24_fs382_not0 & b[22];
  assign f_arrdiv24_fs382_xor1 = f_arrdiv24_fs381_or0 ^ f_arrdiv24_fs382_xor0;
  assign f_arrdiv24_fs382_not1 = ~f_arrdiv24_fs382_xor0;
  assign f_arrdiv24_fs382_and1 = f_arrdiv24_fs382_not1 & f_arrdiv24_fs381_or0;
  assign f_arrdiv24_fs382_or0 = f_arrdiv24_fs382_and1 | f_arrdiv24_fs382_and0;
  assign f_arrdiv24_fs383_xor0 = f_arrdiv24_mux2to1344_xor0 ^ b[23];
  assign f_arrdiv24_fs383_not0 = ~f_arrdiv24_mux2to1344_xor0;
  assign f_arrdiv24_fs383_and0 = f_arrdiv24_fs383_not0 & b[23];
  assign f_arrdiv24_fs383_xor1 = f_arrdiv24_fs382_or0 ^ f_arrdiv24_fs383_xor0;
  assign f_arrdiv24_fs383_not1 = ~f_arrdiv24_fs383_xor0;
  assign f_arrdiv24_fs383_and1 = f_arrdiv24_fs383_not1 & f_arrdiv24_fs382_or0;
  assign f_arrdiv24_fs383_or0 = f_arrdiv24_fs383_and1 | f_arrdiv24_fs383_and0;
  assign f_arrdiv24_mux2to1345_and0 = a[8] & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1345_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1345_and1 = f_arrdiv24_fs360_xor0 & f_arrdiv24_mux2to1345_not0;
  assign f_arrdiv24_mux2to1345_xor0 = f_arrdiv24_mux2to1345_and0 ^ f_arrdiv24_mux2to1345_and1;
  assign f_arrdiv24_mux2to1346_and0 = f_arrdiv24_mux2to1322_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1346_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1346_and1 = f_arrdiv24_fs361_xor1 & f_arrdiv24_mux2to1346_not0;
  assign f_arrdiv24_mux2to1346_xor0 = f_arrdiv24_mux2to1346_and0 ^ f_arrdiv24_mux2to1346_and1;
  assign f_arrdiv24_mux2to1347_and0 = f_arrdiv24_mux2to1323_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1347_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1347_and1 = f_arrdiv24_fs362_xor1 & f_arrdiv24_mux2to1347_not0;
  assign f_arrdiv24_mux2to1347_xor0 = f_arrdiv24_mux2to1347_and0 ^ f_arrdiv24_mux2to1347_and1;
  assign f_arrdiv24_mux2to1348_and0 = f_arrdiv24_mux2to1324_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1348_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1348_and1 = f_arrdiv24_fs363_xor1 & f_arrdiv24_mux2to1348_not0;
  assign f_arrdiv24_mux2to1348_xor0 = f_arrdiv24_mux2to1348_and0 ^ f_arrdiv24_mux2to1348_and1;
  assign f_arrdiv24_mux2to1349_and0 = f_arrdiv24_mux2to1325_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1349_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1349_and1 = f_arrdiv24_fs364_xor1 & f_arrdiv24_mux2to1349_not0;
  assign f_arrdiv24_mux2to1349_xor0 = f_arrdiv24_mux2to1349_and0 ^ f_arrdiv24_mux2to1349_and1;
  assign f_arrdiv24_mux2to1350_and0 = f_arrdiv24_mux2to1326_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1350_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1350_and1 = f_arrdiv24_fs365_xor1 & f_arrdiv24_mux2to1350_not0;
  assign f_arrdiv24_mux2to1350_xor0 = f_arrdiv24_mux2to1350_and0 ^ f_arrdiv24_mux2to1350_and1;
  assign f_arrdiv24_mux2to1351_and0 = f_arrdiv24_mux2to1327_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1351_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1351_and1 = f_arrdiv24_fs366_xor1 & f_arrdiv24_mux2to1351_not0;
  assign f_arrdiv24_mux2to1351_xor0 = f_arrdiv24_mux2to1351_and0 ^ f_arrdiv24_mux2to1351_and1;
  assign f_arrdiv24_mux2to1352_and0 = f_arrdiv24_mux2to1328_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1352_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1352_and1 = f_arrdiv24_fs367_xor1 & f_arrdiv24_mux2to1352_not0;
  assign f_arrdiv24_mux2to1352_xor0 = f_arrdiv24_mux2to1352_and0 ^ f_arrdiv24_mux2to1352_and1;
  assign f_arrdiv24_mux2to1353_and0 = f_arrdiv24_mux2to1329_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1353_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1353_and1 = f_arrdiv24_fs368_xor1 & f_arrdiv24_mux2to1353_not0;
  assign f_arrdiv24_mux2to1353_xor0 = f_arrdiv24_mux2to1353_and0 ^ f_arrdiv24_mux2to1353_and1;
  assign f_arrdiv24_mux2to1354_and0 = f_arrdiv24_mux2to1330_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1354_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1354_and1 = f_arrdiv24_fs369_xor1 & f_arrdiv24_mux2to1354_not0;
  assign f_arrdiv24_mux2to1354_xor0 = f_arrdiv24_mux2to1354_and0 ^ f_arrdiv24_mux2to1354_and1;
  assign f_arrdiv24_mux2to1355_and0 = f_arrdiv24_mux2to1331_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1355_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1355_and1 = f_arrdiv24_fs370_xor1 & f_arrdiv24_mux2to1355_not0;
  assign f_arrdiv24_mux2to1355_xor0 = f_arrdiv24_mux2to1355_and0 ^ f_arrdiv24_mux2to1355_and1;
  assign f_arrdiv24_mux2to1356_and0 = f_arrdiv24_mux2to1332_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1356_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1356_and1 = f_arrdiv24_fs371_xor1 & f_arrdiv24_mux2to1356_not0;
  assign f_arrdiv24_mux2to1356_xor0 = f_arrdiv24_mux2to1356_and0 ^ f_arrdiv24_mux2to1356_and1;
  assign f_arrdiv24_mux2to1357_and0 = f_arrdiv24_mux2to1333_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1357_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1357_and1 = f_arrdiv24_fs372_xor1 & f_arrdiv24_mux2to1357_not0;
  assign f_arrdiv24_mux2to1357_xor0 = f_arrdiv24_mux2to1357_and0 ^ f_arrdiv24_mux2to1357_and1;
  assign f_arrdiv24_mux2to1358_and0 = f_arrdiv24_mux2to1334_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1358_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1358_and1 = f_arrdiv24_fs373_xor1 & f_arrdiv24_mux2to1358_not0;
  assign f_arrdiv24_mux2to1358_xor0 = f_arrdiv24_mux2to1358_and0 ^ f_arrdiv24_mux2to1358_and1;
  assign f_arrdiv24_mux2to1359_and0 = f_arrdiv24_mux2to1335_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1359_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1359_and1 = f_arrdiv24_fs374_xor1 & f_arrdiv24_mux2to1359_not0;
  assign f_arrdiv24_mux2to1359_xor0 = f_arrdiv24_mux2to1359_and0 ^ f_arrdiv24_mux2to1359_and1;
  assign f_arrdiv24_mux2to1360_and0 = f_arrdiv24_mux2to1336_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1360_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1360_and1 = f_arrdiv24_fs375_xor1 & f_arrdiv24_mux2to1360_not0;
  assign f_arrdiv24_mux2to1360_xor0 = f_arrdiv24_mux2to1360_and0 ^ f_arrdiv24_mux2to1360_and1;
  assign f_arrdiv24_mux2to1361_and0 = f_arrdiv24_mux2to1337_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1361_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1361_and1 = f_arrdiv24_fs376_xor1 & f_arrdiv24_mux2to1361_not0;
  assign f_arrdiv24_mux2to1361_xor0 = f_arrdiv24_mux2to1361_and0 ^ f_arrdiv24_mux2to1361_and1;
  assign f_arrdiv24_mux2to1362_and0 = f_arrdiv24_mux2to1338_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1362_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1362_and1 = f_arrdiv24_fs377_xor1 & f_arrdiv24_mux2to1362_not0;
  assign f_arrdiv24_mux2to1362_xor0 = f_arrdiv24_mux2to1362_and0 ^ f_arrdiv24_mux2to1362_and1;
  assign f_arrdiv24_mux2to1363_and0 = f_arrdiv24_mux2to1339_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1363_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1363_and1 = f_arrdiv24_fs378_xor1 & f_arrdiv24_mux2to1363_not0;
  assign f_arrdiv24_mux2to1363_xor0 = f_arrdiv24_mux2to1363_and0 ^ f_arrdiv24_mux2to1363_and1;
  assign f_arrdiv24_mux2to1364_and0 = f_arrdiv24_mux2to1340_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1364_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1364_and1 = f_arrdiv24_fs379_xor1 & f_arrdiv24_mux2to1364_not0;
  assign f_arrdiv24_mux2to1364_xor0 = f_arrdiv24_mux2to1364_and0 ^ f_arrdiv24_mux2to1364_and1;
  assign f_arrdiv24_mux2to1365_and0 = f_arrdiv24_mux2to1341_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1365_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1365_and1 = f_arrdiv24_fs380_xor1 & f_arrdiv24_mux2to1365_not0;
  assign f_arrdiv24_mux2to1365_xor0 = f_arrdiv24_mux2to1365_and0 ^ f_arrdiv24_mux2to1365_and1;
  assign f_arrdiv24_mux2to1366_and0 = f_arrdiv24_mux2to1342_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1366_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1366_and1 = f_arrdiv24_fs381_xor1 & f_arrdiv24_mux2to1366_not0;
  assign f_arrdiv24_mux2to1366_xor0 = f_arrdiv24_mux2to1366_and0 ^ f_arrdiv24_mux2to1366_and1;
  assign f_arrdiv24_mux2to1367_and0 = f_arrdiv24_mux2to1343_xor0 & f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1367_not0 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_mux2to1367_and1 = f_arrdiv24_fs382_xor1 & f_arrdiv24_mux2to1367_not0;
  assign f_arrdiv24_mux2to1367_xor0 = f_arrdiv24_mux2to1367_and0 ^ f_arrdiv24_mux2to1367_and1;
  assign f_arrdiv24_not15 = ~f_arrdiv24_fs383_or0;
  assign f_arrdiv24_fs384_xor0 = a[7] ^ b[0];
  assign f_arrdiv24_fs384_not0 = ~a[7];
  assign f_arrdiv24_fs384_and0 = f_arrdiv24_fs384_not0 & b[0];
  assign f_arrdiv24_fs384_not1 = ~f_arrdiv24_fs384_xor0;
  assign f_arrdiv24_fs385_xor0 = f_arrdiv24_mux2to1345_xor0 ^ b[1];
  assign f_arrdiv24_fs385_not0 = ~f_arrdiv24_mux2to1345_xor0;
  assign f_arrdiv24_fs385_and0 = f_arrdiv24_fs385_not0 & b[1];
  assign f_arrdiv24_fs385_xor1 = f_arrdiv24_fs384_and0 ^ f_arrdiv24_fs385_xor0;
  assign f_arrdiv24_fs385_not1 = ~f_arrdiv24_fs385_xor0;
  assign f_arrdiv24_fs385_and1 = f_arrdiv24_fs385_not1 & f_arrdiv24_fs384_and0;
  assign f_arrdiv24_fs385_or0 = f_arrdiv24_fs385_and1 | f_arrdiv24_fs385_and0;
  assign f_arrdiv24_fs386_xor0 = f_arrdiv24_mux2to1346_xor0 ^ b[2];
  assign f_arrdiv24_fs386_not0 = ~f_arrdiv24_mux2to1346_xor0;
  assign f_arrdiv24_fs386_and0 = f_arrdiv24_fs386_not0 & b[2];
  assign f_arrdiv24_fs386_xor1 = f_arrdiv24_fs385_or0 ^ f_arrdiv24_fs386_xor0;
  assign f_arrdiv24_fs386_not1 = ~f_arrdiv24_fs386_xor0;
  assign f_arrdiv24_fs386_and1 = f_arrdiv24_fs386_not1 & f_arrdiv24_fs385_or0;
  assign f_arrdiv24_fs386_or0 = f_arrdiv24_fs386_and1 | f_arrdiv24_fs386_and0;
  assign f_arrdiv24_fs387_xor0 = f_arrdiv24_mux2to1347_xor0 ^ b[3];
  assign f_arrdiv24_fs387_not0 = ~f_arrdiv24_mux2to1347_xor0;
  assign f_arrdiv24_fs387_and0 = f_arrdiv24_fs387_not0 & b[3];
  assign f_arrdiv24_fs387_xor1 = f_arrdiv24_fs386_or0 ^ f_arrdiv24_fs387_xor0;
  assign f_arrdiv24_fs387_not1 = ~f_arrdiv24_fs387_xor0;
  assign f_arrdiv24_fs387_and1 = f_arrdiv24_fs387_not1 & f_arrdiv24_fs386_or0;
  assign f_arrdiv24_fs387_or0 = f_arrdiv24_fs387_and1 | f_arrdiv24_fs387_and0;
  assign f_arrdiv24_fs388_xor0 = f_arrdiv24_mux2to1348_xor0 ^ b[4];
  assign f_arrdiv24_fs388_not0 = ~f_arrdiv24_mux2to1348_xor0;
  assign f_arrdiv24_fs388_and0 = f_arrdiv24_fs388_not0 & b[4];
  assign f_arrdiv24_fs388_xor1 = f_arrdiv24_fs387_or0 ^ f_arrdiv24_fs388_xor0;
  assign f_arrdiv24_fs388_not1 = ~f_arrdiv24_fs388_xor0;
  assign f_arrdiv24_fs388_and1 = f_arrdiv24_fs388_not1 & f_arrdiv24_fs387_or0;
  assign f_arrdiv24_fs388_or0 = f_arrdiv24_fs388_and1 | f_arrdiv24_fs388_and0;
  assign f_arrdiv24_fs389_xor0 = f_arrdiv24_mux2to1349_xor0 ^ b[5];
  assign f_arrdiv24_fs389_not0 = ~f_arrdiv24_mux2to1349_xor0;
  assign f_arrdiv24_fs389_and0 = f_arrdiv24_fs389_not0 & b[5];
  assign f_arrdiv24_fs389_xor1 = f_arrdiv24_fs388_or0 ^ f_arrdiv24_fs389_xor0;
  assign f_arrdiv24_fs389_not1 = ~f_arrdiv24_fs389_xor0;
  assign f_arrdiv24_fs389_and1 = f_arrdiv24_fs389_not1 & f_arrdiv24_fs388_or0;
  assign f_arrdiv24_fs389_or0 = f_arrdiv24_fs389_and1 | f_arrdiv24_fs389_and0;
  assign f_arrdiv24_fs390_xor0 = f_arrdiv24_mux2to1350_xor0 ^ b[6];
  assign f_arrdiv24_fs390_not0 = ~f_arrdiv24_mux2to1350_xor0;
  assign f_arrdiv24_fs390_and0 = f_arrdiv24_fs390_not0 & b[6];
  assign f_arrdiv24_fs390_xor1 = f_arrdiv24_fs389_or0 ^ f_arrdiv24_fs390_xor0;
  assign f_arrdiv24_fs390_not1 = ~f_arrdiv24_fs390_xor0;
  assign f_arrdiv24_fs390_and1 = f_arrdiv24_fs390_not1 & f_arrdiv24_fs389_or0;
  assign f_arrdiv24_fs390_or0 = f_arrdiv24_fs390_and1 | f_arrdiv24_fs390_and0;
  assign f_arrdiv24_fs391_xor0 = f_arrdiv24_mux2to1351_xor0 ^ b[7];
  assign f_arrdiv24_fs391_not0 = ~f_arrdiv24_mux2to1351_xor0;
  assign f_arrdiv24_fs391_and0 = f_arrdiv24_fs391_not0 & b[7];
  assign f_arrdiv24_fs391_xor1 = f_arrdiv24_fs390_or0 ^ f_arrdiv24_fs391_xor0;
  assign f_arrdiv24_fs391_not1 = ~f_arrdiv24_fs391_xor0;
  assign f_arrdiv24_fs391_and1 = f_arrdiv24_fs391_not1 & f_arrdiv24_fs390_or0;
  assign f_arrdiv24_fs391_or0 = f_arrdiv24_fs391_and1 | f_arrdiv24_fs391_and0;
  assign f_arrdiv24_fs392_xor0 = f_arrdiv24_mux2to1352_xor0 ^ b[8];
  assign f_arrdiv24_fs392_not0 = ~f_arrdiv24_mux2to1352_xor0;
  assign f_arrdiv24_fs392_and0 = f_arrdiv24_fs392_not0 & b[8];
  assign f_arrdiv24_fs392_xor1 = f_arrdiv24_fs391_or0 ^ f_arrdiv24_fs392_xor0;
  assign f_arrdiv24_fs392_not1 = ~f_arrdiv24_fs392_xor0;
  assign f_arrdiv24_fs392_and1 = f_arrdiv24_fs392_not1 & f_arrdiv24_fs391_or0;
  assign f_arrdiv24_fs392_or0 = f_arrdiv24_fs392_and1 | f_arrdiv24_fs392_and0;
  assign f_arrdiv24_fs393_xor0 = f_arrdiv24_mux2to1353_xor0 ^ b[9];
  assign f_arrdiv24_fs393_not0 = ~f_arrdiv24_mux2to1353_xor0;
  assign f_arrdiv24_fs393_and0 = f_arrdiv24_fs393_not0 & b[9];
  assign f_arrdiv24_fs393_xor1 = f_arrdiv24_fs392_or0 ^ f_arrdiv24_fs393_xor0;
  assign f_arrdiv24_fs393_not1 = ~f_arrdiv24_fs393_xor0;
  assign f_arrdiv24_fs393_and1 = f_arrdiv24_fs393_not1 & f_arrdiv24_fs392_or0;
  assign f_arrdiv24_fs393_or0 = f_arrdiv24_fs393_and1 | f_arrdiv24_fs393_and0;
  assign f_arrdiv24_fs394_xor0 = f_arrdiv24_mux2to1354_xor0 ^ b[10];
  assign f_arrdiv24_fs394_not0 = ~f_arrdiv24_mux2to1354_xor0;
  assign f_arrdiv24_fs394_and0 = f_arrdiv24_fs394_not0 & b[10];
  assign f_arrdiv24_fs394_xor1 = f_arrdiv24_fs393_or0 ^ f_arrdiv24_fs394_xor0;
  assign f_arrdiv24_fs394_not1 = ~f_arrdiv24_fs394_xor0;
  assign f_arrdiv24_fs394_and1 = f_arrdiv24_fs394_not1 & f_arrdiv24_fs393_or0;
  assign f_arrdiv24_fs394_or0 = f_arrdiv24_fs394_and1 | f_arrdiv24_fs394_and0;
  assign f_arrdiv24_fs395_xor0 = f_arrdiv24_mux2to1355_xor0 ^ b[11];
  assign f_arrdiv24_fs395_not0 = ~f_arrdiv24_mux2to1355_xor0;
  assign f_arrdiv24_fs395_and0 = f_arrdiv24_fs395_not0 & b[11];
  assign f_arrdiv24_fs395_xor1 = f_arrdiv24_fs394_or0 ^ f_arrdiv24_fs395_xor0;
  assign f_arrdiv24_fs395_not1 = ~f_arrdiv24_fs395_xor0;
  assign f_arrdiv24_fs395_and1 = f_arrdiv24_fs395_not1 & f_arrdiv24_fs394_or0;
  assign f_arrdiv24_fs395_or0 = f_arrdiv24_fs395_and1 | f_arrdiv24_fs395_and0;
  assign f_arrdiv24_fs396_xor0 = f_arrdiv24_mux2to1356_xor0 ^ b[12];
  assign f_arrdiv24_fs396_not0 = ~f_arrdiv24_mux2to1356_xor0;
  assign f_arrdiv24_fs396_and0 = f_arrdiv24_fs396_not0 & b[12];
  assign f_arrdiv24_fs396_xor1 = f_arrdiv24_fs395_or0 ^ f_arrdiv24_fs396_xor0;
  assign f_arrdiv24_fs396_not1 = ~f_arrdiv24_fs396_xor0;
  assign f_arrdiv24_fs396_and1 = f_arrdiv24_fs396_not1 & f_arrdiv24_fs395_or0;
  assign f_arrdiv24_fs396_or0 = f_arrdiv24_fs396_and1 | f_arrdiv24_fs396_and0;
  assign f_arrdiv24_fs397_xor0 = f_arrdiv24_mux2to1357_xor0 ^ b[13];
  assign f_arrdiv24_fs397_not0 = ~f_arrdiv24_mux2to1357_xor0;
  assign f_arrdiv24_fs397_and0 = f_arrdiv24_fs397_not0 & b[13];
  assign f_arrdiv24_fs397_xor1 = f_arrdiv24_fs396_or0 ^ f_arrdiv24_fs397_xor0;
  assign f_arrdiv24_fs397_not1 = ~f_arrdiv24_fs397_xor0;
  assign f_arrdiv24_fs397_and1 = f_arrdiv24_fs397_not1 & f_arrdiv24_fs396_or0;
  assign f_arrdiv24_fs397_or0 = f_arrdiv24_fs397_and1 | f_arrdiv24_fs397_and0;
  assign f_arrdiv24_fs398_xor0 = f_arrdiv24_mux2to1358_xor0 ^ b[14];
  assign f_arrdiv24_fs398_not0 = ~f_arrdiv24_mux2to1358_xor0;
  assign f_arrdiv24_fs398_and0 = f_arrdiv24_fs398_not0 & b[14];
  assign f_arrdiv24_fs398_xor1 = f_arrdiv24_fs397_or0 ^ f_arrdiv24_fs398_xor0;
  assign f_arrdiv24_fs398_not1 = ~f_arrdiv24_fs398_xor0;
  assign f_arrdiv24_fs398_and1 = f_arrdiv24_fs398_not1 & f_arrdiv24_fs397_or0;
  assign f_arrdiv24_fs398_or0 = f_arrdiv24_fs398_and1 | f_arrdiv24_fs398_and0;
  assign f_arrdiv24_fs399_xor0 = f_arrdiv24_mux2to1359_xor0 ^ b[15];
  assign f_arrdiv24_fs399_not0 = ~f_arrdiv24_mux2to1359_xor0;
  assign f_arrdiv24_fs399_and0 = f_arrdiv24_fs399_not0 & b[15];
  assign f_arrdiv24_fs399_xor1 = f_arrdiv24_fs398_or0 ^ f_arrdiv24_fs399_xor0;
  assign f_arrdiv24_fs399_not1 = ~f_arrdiv24_fs399_xor0;
  assign f_arrdiv24_fs399_and1 = f_arrdiv24_fs399_not1 & f_arrdiv24_fs398_or0;
  assign f_arrdiv24_fs399_or0 = f_arrdiv24_fs399_and1 | f_arrdiv24_fs399_and0;
  assign f_arrdiv24_fs400_xor0 = f_arrdiv24_mux2to1360_xor0 ^ b[16];
  assign f_arrdiv24_fs400_not0 = ~f_arrdiv24_mux2to1360_xor0;
  assign f_arrdiv24_fs400_and0 = f_arrdiv24_fs400_not0 & b[16];
  assign f_arrdiv24_fs400_xor1 = f_arrdiv24_fs399_or0 ^ f_arrdiv24_fs400_xor0;
  assign f_arrdiv24_fs400_not1 = ~f_arrdiv24_fs400_xor0;
  assign f_arrdiv24_fs400_and1 = f_arrdiv24_fs400_not1 & f_arrdiv24_fs399_or0;
  assign f_arrdiv24_fs400_or0 = f_arrdiv24_fs400_and1 | f_arrdiv24_fs400_and0;
  assign f_arrdiv24_fs401_xor0 = f_arrdiv24_mux2to1361_xor0 ^ b[17];
  assign f_arrdiv24_fs401_not0 = ~f_arrdiv24_mux2to1361_xor0;
  assign f_arrdiv24_fs401_and0 = f_arrdiv24_fs401_not0 & b[17];
  assign f_arrdiv24_fs401_xor1 = f_arrdiv24_fs400_or0 ^ f_arrdiv24_fs401_xor0;
  assign f_arrdiv24_fs401_not1 = ~f_arrdiv24_fs401_xor0;
  assign f_arrdiv24_fs401_and1 = f_arrdiv24_fs401_not1 & f_arrdiv24_fs400_or0;
  assign f_arrdiv24_fs401_or0 = f_arrdiv24_fs401_and1 | f_arrdiv24_fs401_and0;
  assign f_arrdiv24_fs402_xor0 = f_arrdiv24_mux2to1362_xor0 ^ b[18];
  assign f_arrdiv24_fs402_not0 = ~f_arrdiv24_mux2to1362_xor0;
  assign f_arrdiv24_fs402_and0 = f_arrdiv24_fs402_not0 & b[18];
  assign f_arrdiv24_fs402_xor1 = f_arrdiv24_fs401_or0 ^ f_arrdiv24_fs402_xor0;
  assign f_arrdiv24_fs402_not1 = ~f_arrdiv24_fs402_xor0;
  assign f_arrdiv24_fs402_and1 = f_arrdiv24_fs402_not1 & f_arrdiv24_fs401_or0;
  assign f_arrdiv24_fs402_or0 = f_arrdiv24_fs402_and1 | f_arrdiv24_fs402_and0;
  assign f_arrdiv24_fs403_xor0 = f_arrdiv24_mux2to1363_xor0 ^ b[19];
  assign f_arrdiv24_fs403_not0 = ~f_arrdiv24_mux2to1363_xor0;
  assign f_arrdiv24_fs403_and0 = f_arrdiv24_fs403_not0 & b[19];
  assign f_arrdiv24_fs403_xor1 = f_arrdiv24_fs402_or0 ^ f_arrdiv24_fs403_xor0;
  assign f_arrdiv24_fs403_not1 = ~f_arrdiv24_fs403_xor0;
  assign f_arrdiv24_fs403_and1 = f_arrdiv24_fs403_not1 & f_arrdiv24_fs402_or0;
  assign f_arrdiv24_fs403_or0 = f_arrdiv24_fs403_and1 | f_arrdiv24_fs403_and0;
  assign f_arrdiv24_fs404_xor0 = f_arrdiv24_mux2to1364_xor0 ^ b[20];
  assign f_arrdiv24_fs404_not0 = ~f_arrdiv24_mux2to1364_xor0;
  assign f_arrdiv24_fs404_and0 = f_arrdiv24_fs404_not0 & b[20];
  assign f_arrdiv24_fs404_xor1 = f_arrdiv24_fs403_or0 ^ f_arrdiv24_fs404_xor0;
  assign f_arrdiv24_fs404_not1 = ~f_arrdiv24_fs404_xor0;
  assign f_arrdiv24_fs404_and1 = f_arrdiv24_fs404_not1 & f_arrdiv24_fs403_or0;
  assign f_arrdiv24_fs404_or0 = f_arrdiv24_fs404_and1 | f_arrdiv24_fs404_and0;
  assign f_arrdiv24_fs405_xor0 = f_arrdiv24_mux2to1365_xor0 ^ b[21];
  assign f_arrdiv24_fs405_not0 = ~f_arrdiv24_mux2to1365_xor0;
  assign f_arrdiv24_fs405_and0 = f_arrdiv24_fs405_not0 & b[21];
  assign f_arrdiv24_fs405_xor1 = f_arrdiv24_fs404_or0 ^ f_arrdiv24_fs405_xor0;
  assign f_arrdiv24_fs405_not1 = ~f_arrdiv24_fs405_xor0;
  assign f_arrdiv24_fs405_and1 = f_arrdiv24_fs405_not1 & f_arrdiv24_fs404_or0;
  assign f_arrdiv24_fs405_or0 = f_arrdiv24_fs405_and1 | f_arrdiv24_fs405_and0;
  assign f_arrdiv24_fs406_xor0 = f_arrdiv24_mux2to1366_xor0 ^ b[22];
  assign f_arrdiv24_fs406_not0 = ~f_arrdiv24_mux2to1366_xor0;
  assign f_arrdiv24_fs406_and0 = f_arrdiv24_fs406_not0 & b[22];
  assign f_arrdiv24_fs406_xor1 = f_arrdiv24_fs405_or0 ^ f_arrdiv24_fs406_xor0;
  assign f_arrdiv24_fs406_not1 = ~f_arrdiv24_fs406_xor0;
  assign f_arrdiv24_fs406_and1 = f_arrdiv24_fs406_not1 & f_arrdiv24_fs405_or0;
  assign f_arrdiv24_fs406_or0 = f_arrdiv24_fs406_and1 | f_arrdiv24_fs406_and0;
  assign f_arrdiv24_fs407_xor0 = f_arrdiv24_mux2to1367_xor0 ^ b[23];
  assign f_arrdiv24_fs407_not0 = ~f_arrdiv24_mux2to1367_xor0;
  assign f_arrdiv24_fs407_and0 = f_arrdiv24_fs407_not0 & b[23];
  assign f_arrdiv24_fs407_xor1 = f_arrdiv24_fs406_or0 ^ f_arrdiv24_fs407_xor0;
  assign f_arrdiv24_fs407_not1 = ~f_arrdiv24_fs407_xor0;
  assign f_arrdiv24_fs407_and1 = f_arrdiv24_fs407_not1 & f_arrdiv24_fs406_or0;
  assign f_arrdiv24_fs407_or0 = f_arrdiv24_fs407_and1 | f_arrdiv24_fs407_and0;
  assign f_arrdiv24_mux2to1368_and0 = a[7] & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1368_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1368_and1 = f_arrdiv24_fs384_xor0 & f_arrdiv24_mux2to1368_not0;
  assign f_arrdiv24_mux2to1368_xor0 = f_arrdiv24_mux2to1368_and0 ^ f_arrdiv24_mux2to1368_and1;
  assign f_arrdiv24_mux2to1369_and0 = f_arrdiv24_mux2to1345_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1369_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1369_and1 = f_arrdiv24_fs385_xor1 & f_arrdiv24_mux2to1369_not0;
  assign f_arrdiv24_mux2to1369_xor0 = f_arrdiv24_mux2to1369_and0 ^ f_arrdiv24_mux2to1369_and1;
  assign f_arrdiv24_mux2to1370_and0 = f_arrdiv24_mux2to1346_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1370_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1370_and1 = f_arrdiv24_fs386_xor1 & f_arrdiv24_mux2to1370_not0;
  assign f_arrdiv24_mux2to1370_xor0 = f_arrdiv24_mux2to1370_and0 ^ f_arrdiv24_mux2to1370_and1;
  assign f_arrdiv24_mux2to1371_and0 = f_arrdiv24_mux2to1347_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1371_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1371_and1 = f_arrdiv24_fs387_xor1 & f_arrdiv24_mux2to1371_not0;
  assign f_arrdiv24_mux2to1371_xor0 = f_arrdiv24_mux2to1371_and0 ^ f_arrdiv24_mux2to1371_and1;
  assign f_arrdiv24_mux2to1372_and0 = f_arrdiv24_mux2to1348_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1372_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1372_and1 = f_arrdiv24_fs388_xor1 & f_arrdiv24_mux2to1372_not0;
  assign f_arrdiv24_mux2to1372_xor0 = f_arrdiv24_mux2to1372_and0 ^ f_arrdiv24_mux2to1372_and1;
  assign f_arrdiv24_mux2to1373_and0 = f_arrdiv24_mux2to1349_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1373_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1373_and1 = f_arrdiv24_fs389_xor1 & f_arrdiv24_mux2to1373_not0;
  assign f_arrdiv24_mux2to1373_xor0 = f_arrdiv24_mux2to1373_and0 ^ f_arrdiv24_mux2to1373_and1;
  assign f_arrdiv24_mux2to1374_and0 = f_arrdiv24_mux2to1350_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1374_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1374_and1 = f_arrdiv24_fs390_xor1 & f_arrdiv24_mux2to1374_not0;
  assign f_arrdiv24_mux2to1374_xor0 = f_arrdiv24_mux2to1374_and0 ^ f_arrdiv24_mux2to1374_and1;
  assign f_arrdiv24_mux2to1375_and0 = f_arrdiv24_mux2to1351_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1375_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1375_and1 = f_arrdiv24_fs391_xor1 & f_arrdiv24_mux2to1375_not0;
  assign f_arrdiv24_mux2to1375_xor0 = f_arrdiv24_mux2to1375_and0 ^ f_arrdiv24_mux2to1375_and1;
  assign f_arrdiv24_mux2to1376_and0 = f_arrdiv24_mux2to1352_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1376_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1376_and1 = f_arrdiv24_fs392_xor1 & f_arrdiv24_mux2to1376_not0;
  assign f_arrdiv24_mux2to1376_xor0 = f_arrdiv24_mux2to1376_and0 ^ f_arrdiv24_mux2to1376_and1;
  assign f_arrdiv24_mux2to1377_and0 = f_arrdiv24_mux2to1353_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1377_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1377_and1 = f_arrdiv24_fs393_xor1 & f_arrdiv24_mux2to1377_not0;
  assign f_arrdiv24_mux2to1377_xor0 = f_arrdiv24_mux2to1377_and0 ^ f_arrdiv24_mux2to1377_and1;
  assign f_arrdiv24_mux2to1378_and0 = f_arrdiv24_mux2to1354_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1378_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1378_and1 = f_arrdiv24_fs394_xor1 & f_arrdiv24_mux2to1378_not0;
  assign f_arrdiv24_mux2to1378_xor0 = f_arrdiv24_mux2to1378_and0 ^ f_arrdiv24_mux2to1378_and1;
  assign f_arrdiv24_mux2to1379_and0 = f_arrdiv24_mux2to1355_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1379_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1379_and1 = f_arrdiv24_fs395_xor1 & f_arrdiv24_mux2to1379_not0;
  assign f_arrdiv24_mux2to1379_xor0 = f_arrdiv24_mux2to1379_and0 ^ f_arrdiv24_mux2to1379_and1;
  assign f_arrdiv24_mux2to1380_and0 = f_arrdiv24_mux2to1356_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1380_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1380_and1 = f_arrdiv24_fs396_xor1 & f_arrdiv24_mux2to1380_not0;
  assign f_arrdiv24_mux2to1380_xor0 = f_arrdiv24_mux2to1380_and0 ^ f_arrdiv24_mux2to1380_and1;
  assign f_arrdiv24_mux2to1381_and0 = f_arrdiv24_mux2to1357_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1381_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1381_and1 = f_arrdiv24_fs397_xor1 & f_arrdiv24_mux2to1381_not0;
  assign f_arrdiv24_mux2to1381_xor0 = f_arrdiv24_mux2to1381_and0 ^ f_arrdiv24_mux2to1381_and1;
  assign f_arrdiv24_mux2to1382_and0 = f_arrdiv24_mux2to1358_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1382_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1382_and1 = f_arrdiv24_fs398_xor1 & f_arrdiv24_mux2to1382_not0;
  assign f_arrdiv24_mux2to1382_xor0 = f_arrdiv24_mux2to1382_and0 ^ f_arrdiv24_mux2to1382_and1;
  assign f_arrdiv24_mux2to1383_and0 = f_arrdiv24_mux2to1359_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1383_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1383_and1 = f_arrdiv24_fs399_xor1 & f_arrdiv24_mux2to1383_not0;
  assign f_arrdiv24_mux2to1383_xor0 = f_arrdiv24_mux2to1383_and0 ^ f_arrdiv24_mux2to1383_and1;
  assign f_arrdiv24_mux2to1384_and0 = f_arrdiv24_mux2to1360_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1384_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1384_and1 = f_arrdiv24_fs400_xor1 & f_arrdiv24_mux2to1384_not0;
  assign f_arrdiv24_mux2to1384_xor0 = f_arrdiv24_mux2to1384_and0 ^ f_arrdiv24_mux2to1384_and1;
  assign f_arrdiv24_mux2to1385_and0 = f_arrdiv24_mux2to1361_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1385_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1385_and1 = f_arrdiv24_fs401_xor1 & f_arrdiv24_mux2to1385_not0;
  assign f_arrdiv24_mux2to1385_xor0 = f_arrdiv24_mux2to1385_and0 ^ f_arrdiv24_mux2to1385_and1;
  assign f_arrdiv24_mux2to1386_and0 = f_arrdiv24_mux2to1362_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1386_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1386_and1 = f_arrdiv24_fs402_xor1 & f_arrdiv24_mux2to1386_not0;
  assign f_arrdiv24_mux2to1386_xor0 = f_arrdiv24_mux2to1386_and0 ^ f_arrdiv24_mux2to1386_and1;
  assign f_arrdiv24_mux2to1387_and0 = f_arrdiv24_mux2to1363_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1387_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1387_and1 = f_arrdiv24_fs403_xor1 & f_arrdiv24_mux2to1387_not0;
  assign f_arrdiv24_mux2to1387_xor0 = f_arrdiv24_mux2to1387_and0 ^ f_arrdiv24_mux2to1387_and1;
  assign f_arrdiv24_mux2to1388_and0 = f_arrdiv24_mux2to1364_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1388_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1388_and1 = f_arrdiv24_fs404_xor1 & f_arrdiv24_mux2to1388_not0;
  assign f_arrdiv24_mux2to1388_xor0 = f_arrdiv24_mux2to1388_and0 ^ f_arrdiv24_mux2to1388_and1;
  assign f_arrdiv24_mux2to1389_and0 = f_arrdiv24_mux2to1365_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1389_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1389_and1 = f_arrdiv24_fs405_xor1 & f_arrdiv24_mux2to1389_not0;
  assign f_arrdiv24_mux2to1389_xor0 = f_arrdiv24_mux2to1389_and0 ^ f_arrdiv24_mux2to1389_and1;
  assign f_arrdiv24_mux2to1390_and0 = f_arrdiv24_mux2to1366_xor0 & f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1390_not0 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_mux2to1390_and1 = f_arrdiv24_fs406_xor1 & f_arrdiv24_mux2to1390_not0;
  assign f_arrdiv24_mux2to1390_xor0 = f_arrdiv24_mux2to1390_and0 ^ f_arrdiv24_mux2to1390_and1;
  assign f_arrdiv24_not16 = ~f_arrdiv24_fs407_or0;
  assign f_arrdiv24_fs408_xor0 = a[6] ^ b[0];
  assign f_arrdiv24_fs408_not0 = ~a[6];
  assign f_arrdiv24_fs408_and0 = f_arrdiv24_fs408_not0 & b[0];
  assign f_arrdiv24_fs408_not1 = ~f_arrdiv24_fs408_xor0;
  assign f_arrdiv24_fs409_xor0 = f_arrdiv24_mux2to1368_xor0 ^ b[1];
  assign f_arrdiv24_fs409_not0 = ~f_arrdiv24_mux2to1368_xor0;
  assign f_arrdiv24_fs409_and0 = f_arrdiv24_fs409_not0 & b[1];
  assign f_arrdiv24_fs409_xor1 = f_arrdiv24_fs408_and0 ^ f_arrdiv24_fs409_xor0;
  assign f_arrdiv24_fs409_not1 = ~f_arrdiv24_fs409_xor0;
  assign f_arrdiv24_fs409_and1 = f_arrdiv24_fs409_not1 & f_arrdiv24_fs408_and0;
  assign f_arrdiv24_fs409_or0 = f_arrdiv24_fs409_and1 | f_arrdiv24_fs409_and0;
  assign f_arrdiv24_fs410_xor0 = f_arrdiv24_mux2to1369_xor0 ^ b[2];
  assign f_arrdiv24_fs410_not0 = ~f_arrdiv24_mux2to1369_xor0;
  assign f_arrdiv24_fs410_and0 = f_arrdiv24_fs410_not0 & b[2];
  assign f_arrdiv24_fs410_xor1 = f_arrdiv24_fs409_or0 ^ f_arrdiv24_fs410_xor0;
  assign f_arrdiv24_fs410_not1 = ~f_arrdiv24_fs410_xor0;
  assign f_arrdiv24_fs410_and1 = f_arrdiv24_fs410_not1 & f_arrdiv24_fs409_or0;
  assign f_arrdiv24_fs410_or0 = f_arrdiv24_fs410_and1 | f_arrdiv24_fs410_and0;
  assign f_arrdiv24_fs411_xor0 = f_arrdiv24_mux2to1370_xor0 ^ b[3];
  assign f_arrdiv24_fs411_not0 = ~f_arrdiv24_mux2to1370_xor0;
  assign f_arrdiv24_fs411_and0 = f_arrdiv24_fs411_not0 & b[3];
  assign f_arrdiv24_fs411_xor1 = f_arrdiv24_fs410_or0 ^ f_arrdiv24_fs411_xor0;
  assign f_arrdiv24_fs411_not1 = ~f_arrdiv24_fs411_xor0;
  assign f_arrdiv24_fs411_and1 = f_arrdiv24_fs411_not1 & f_arrdiv24_fs410_or0;
  assign f_arrdiv24_fs411_or0 = f_arrdiv24_fs411_and1 | f_arrdiv24_fs411_and0;
  assign f_arrdiv24_fs412_xor0 = f_arrdiv24_mux2to1371_xor0 ^ b[4];
  assign f_arrdiv24_fs412_not0 = ~f_arrdiv24_mux2to1371_xor0;
  assign f_arrdiv24_fs412_and0 = f_arrdiv24_fs412_not0 & b[4];
  assign f_arrdiv24_fs412_xor1 = f_arrdiv24_fs411_or0 ^ f_arrdiv24_fs412_xor0;
  assign f_arrdiv24_fs412_not1 = ~f_arrdiv24_fs412_xor0;
  assign f_arrdiv24_fs412_and1 = f_arrdiv24_fs412_not1 & f_arrdiv24_fs411_or0;
  assign f_arrdiv24_fs412_or0 = f_arrdiv24_fs412_and1 | f_arrdiv24_fs412_and0;
  assign f_arrdiv24_fs413_xor0 = f_arrdiv24_mux2to1372_xor0 ^ b[5];
  assign f_arrdiv24_fs413_not0 = ~f_arrdiv24_mux2to1372_xor0;
  assign f_arrdiv24_fs413_and0 = f_arrdiv24_fs413_not0 & b[5];
  assign f_arrdiv24_fs413_xor1 = f_arrdiv24_fs412_or0 ^ f_arrdiv24_fs413_xor0;
  assign f_arrdiv24_fs413_not1 = ~f_arrdiv24_fs413_xor0;
  assign f_arrdiv24_fs413_and1 = f_arrdiv24_fs413_not1 & f_arrdiv24_fs412_or0;
  assign f_arrdiv24_fs413_or0 = f_arrdiv24_fs413_and1 | f_arrdiv24_fs413_and0;
  assign f_arrdiv24_fs414_xor0 = f_arrdiv24_mux2to1373_xor0 ^ b[6];
  assign f_arrdiv24_fs414_not0 = ~f_arrdiv24_mux2to1373_xor0;
  assign f_arrdiv24_fs414_and0 = f_arrdiv24_fs414_not0 & b[6];
  assign f_arrdiv24_fs414_xor1 = f_arrdiv24_fs413_or0 ^ f_arrdiv24_fs414_xor0;
  assign f_arrdiv24_fs414_not1 = ~f_arrdiv24_fs414_xor0;
  assign f_arrdiv24_fs414_and1 = f_arrdiv24_fs414_not1 & f_arrdiv24_fs413_or0;
  assign f_arrdiv24_fs414_or0 = f_arrdiv24_fs414_and1 | f_arrdiv24_fs414_and0;
  assign f_arrdiv24_fs415_xor0 = f_arrdiv24_mux2to1374_xor0 ^ b[7];
  assign f_arrdiv24_fs415_not0 = ~f_arrdiv24_mux2to1374_xor0;
  assign f_arrdiv24_fs415_and0 = f_arrdiv24_fs415_not0 & b[7];
  assign f_arrdiv24_fs415_xor1 = f_arrdiv24_fs414_or0 ^ f_arrdiv24_fs415_xor0;
  assign f_arrdiv24_fs415_not1 = ~f_arrdiv24_fs415_xor0;
  assign f_arrdiv24_fs415_and1 = f_arrdiv24_fs415_not1 & f_arrdiv24_fs414_or0;
  assign f_arrdiv24_fs415_or0 = f_arrdiv24_fs415_and1 | f_arrdiv24_fs415_and0;
  assign f_arrdiv24_fs416_xor0 = f_arrdiv24_mux2to1375_xor0 ^ b[8];
  assign f_arrdiv24_fs416_not0 = ~f_arrdiv24_mux2to1375_xor0;
  assign f_arrdiv24_fs416_and0 = f_arrdiv24_fs416_not0 & b[8];
  assign f_arrdiv24_fs416_xor1 = f_arrdiv24_fs415_or0 ^ f_arrdiv24_fs416_xor0;
  assign f_arrdiv24_fs416_not1 = ~f_arrdiv24_fs416_xor0;
  assign f_arrdiv24_fs416_and1 = f_arrdiv24_fs416_not1 & f_arrdiv24_fs415_or0;
  assign f_arrdiv24_fs416_or0 = f_arrdiv24_fs416_and1 | f_arrdiv24_fs416_and0;
  assign f_arrdiv24_fs417_xor0 = f_arrdiv24_mux2to1376_xor0 ^ b[9];
  assign f_arrdiv24_fs417_not0 = ~f_arrdiv24_mux2to1376_xor0;
  assign f_arrdiv24_fs417_and0 = f_arrdiv24_fs417_not0 & b[9];
  assign f_arrdiv24_fs417_xor1 = f_arrdiv24_fs416_or0 ^ f_arrdiv24_fs417_xor0;
  assign f_arrdiv24_fs417_not1 = ~f_arrdiv24_fs417_xor0;
  assign f_arrdiv24_fs417_and1 = f_arrdiv24_fs417_not1 & f_arrdiv24_fs416_or0;
  assign f_arrdiv24_fs417_or0 = f_arrdiv24_fs417_and1 | f_arrdiv24_fs417_and0;
  assign f_arrdiv24_fs418_xor0 = f_arrdiv24_mux2to1377_xor0 ^ b[10];
  assign f_arrdiv24_fs418_not0 = ~f_arrdiv24_mux2to1377_xor0;
  assign f_arrdiv24_fs418_and0 = f_arrdiv24_fs418_not0 & b[10];
  assign f_arrdiv24_fs418_xor1 = f_arrdiv24_fs417_or0 ^ f_arrdiv24_fs418_xor0;
  assign f_arrdiv24_fs418_not1 = ~f_arrdiv24_fs418_xor0;
  assign f_arrdiv24_fs418_and1 = f_arrdiv24_fs418_not1 & f_arrdiv24_fs417_or0;
  assign f_arrdiv24_fs418_or0 = f_arrdiv24_fs418_and1 | f_arrdiv24_fs418_and0;
  assign f_arrdiv24_fs419_xor0 = f_arrdiv24_mux2to1378_xor0 ^ b[11];
  assign f_arrdiv24_fs419_not0 = ~f_arrdiv24_mux2to1378_xor0;
  assign f_arrdiv24_fs419_and0 = f_arrdiv24_fs419_not0 & b[11];
  assign f_arrdiv24_fs419_xor1 = f_arrdiv24_fs418_or0 ^ f_arrdiv24_fs419_xor0;
  assign f_arrdiv24_fs419_not1 = ~f_arrdiv24_fs419_xor0;
  assign f_arrdiv24_fs419_and1 = f_arrdiv24_fs419_not1 & f_arrdiv24_fs418_or0;
  assign f_arrdiv24_fs419_or0 = f_arrdiv24_fs419_and1 | f_arrdiv24_fs419_and0;
  assign f_arrdiv24_fs420_xor0 = f_arrdiv24_mux2to1379_xor0 ^ b[12];
  assign f_arrdiv24_fs420_not0 = ~f_arrdiv24_mux2to1379_xor0;
  assign f_arrdiv24_fs420_and0 = f_arrdiv24_fs420_not0 & b[12];
  assign f_arrdiv24_fs420_xor1 = f_arrdiv24_fs419_or0 ^ f_arrdiv24_fs420_xor0;
  assign f_arrdiv24_fs420_not1 = ~f_arrdiv24_fs420_xor0;
  assign f_arrdiv24_fs420_and1 = f_arrdiv24_fs420_not1 & f_arrdiv24_fs419_or0;
  assign f_arrdiv24_fs420_or0 = f_arrdiv24_fs420_and1 | f_arrdiv24_fs420_and0;
  assign f_arrdiv24_fs421_xor0 = f_arrdiv24_mux2to1380_xor0 ^ b[13];
  assign f_arrdiv24_fs421_not0 = ~f_arrdiv24_mux2to1380_xor0;
  assign f_arrdiv24_fs421_and0 = f_arrdiv24_fs421_not0 & b[13];
  assign f_arrdiv24_fs421_xor1 = f_arrdiv24_fs420_or0 ^ f_arrdiv24_fs421_xor0;
  assign f_arrdiv24_fs421_not1 = ~f_arrdiv24_fs421_xor0;
  assign f_arrdiv24_fs421_and1 = f_arrdiv24_fs421_not1 & f_arrdiv24_fs420_or0;
  assign f_arrdiv24_fs421_or0 = f_arrdiv24_fs421_and1 | f_arrdiv24_fs421_and0;
  assign f_arrdiv24_fs422_xor0 = f_arrdiv24_mux2to1381_xor0 ^ b[14];
  assign f_arrdiv24_fs422_not0 = ~f_arrdiv24_mux2to1381_xor0;
  assign f_arrdiv24_fs422_and0 = f_arrdiv24_fs422_not0 & b[14];
  assign f_arrdiv24_fs422_xor1 = f_arrdiv24_fs421_or0 ^ f_arrdiv24_fs422_xor0;
  assign f_arrdiv24_fs422_not1 = ~f_arrdiv24_fs422_xor0;
  assign f_arrdiv24_fs422_and1 = f_arrdiv24_fs422_not1 & f_arrdiv24_fs421_or0;
  assign f_arrdiv24_fs422_or0 = f_arrdiv24_fs422_and1 | f_arrdiv24_fs422_and0;
  assign f_arrdiv24_fs423_xor0 = f_arrdiv24_mux2to1382_xor0 ^ b[15];
  assign f_arrdiv24_fs423_not0 = ~f_arrdiv24_mux2to1382_xor0;
  assign f_arrdiv24_fs423_and0 = f_arrdiv24_fs423_not0 & b[15];
  assign f_arrdiv24_fs423_xor1 = f_arrdiv24_fs422_or0 ^ f_arrdiv24_fs423_xor0;
  assign f_arrdiv24_fs423_not1 = ~f_arrdiv24_fs423_xor0;
  assign f_arrdiv24_fs423_and1 = f_arrdiv24_fs423_not1 & f_arrdiv24_fs422_or0;
  assign f_arrdiv24_fs423_or0 = f_arrdiv24_fs423_and1 | f_arrdiv24_fs423_and0;
  assign f_arrdiv24_fs424_xor0 = f_arrdiv24_mux2to1383_xor0 ^ b[16];
  assign f_arrdiv24_fs424_not0 = ~f_arrdiv24_mux2to1383_xor0;
  assign f_arrdiv24_fs424_and0 = f_arrdiv24_fs424_not0 & b[16];
  assign f_arrdiv24_fs424_xor1 = f_arrdiv24_fs423_or0 ^ f_arrdiv24_fs424_xor0;
  assign f_arrdiv24_fs424_not1 = ~f_arrdiv24_fs424_xor0;
  assign f_arrdiv24_fs424_and1 = f_arrdiv24_fs424_not1 & f_arrdiv24_fs423_or0;
  assign f_arrdiv24_fs424_or0 = f_arrdiv24_fs424_and1 | f_arrdiv24_fs424_and0;
  assign f_arrdiv24_fs425_xor0 = f_arrdiv24_mux2to1384_xor0 ^ b[17];
  assign f_arrdiv24_fs425_not0 = ~f_arrdiv24_mux2to1384_xor0;
  assign f_arrdiv24_fs425_and0 = f_arrdiv24_fs425_not0 & b[17];
  assign f_arrdiv24_fs425_xor1 = f_arrdiv24_fs424_or0 ^ f_arrdiv24_fs425_xor0;
  assign f_arrdiv24_fs425_not1 = ~f_arrdiv24_fs425_xor0;
  assign f_arrdiv24_fs425_and1 = f_arrdiv24_fs425_not1 & f_arrdiv24_fs424_or0;
  assign f_arrdiv24_fs425_or0 = f_arrdiv24_fs425_and1 | f_arrdiv24_fs425_and0;
  assign f_arrdiv24_fs426_xor0 = f_arrdiv24_mux2to1385_xor0 ^ b[18];
  assign f_arrdiv24_fs426_not0 = ~f_arrdiv24_mux2to1385_xor0;
  assign f_arrdiv24_fs426_and0 = f_arrdiv24_fs426_not0 & b[18];
  assign f_arrdiv24_fs426_xor1 = f_arrdiv24_fs425_or0 ^ f_arrdiv24_fs426_xor0;
  assign f_arrdiv24_fs426_not1 = ~f_arrdiv24_fs426_xor0;
  assign f_arrdiv24_fs426_and1 = f_arrdiv24_fs426_not1 & f_arrdiv24_fs425_or0;
  assign f_arrdiv24_fs426_or0 = f_arrdiv24_fs426_and1 | f_arrdiv24_fs426_and0;
  assign f_arrdiv24_fs427_xor0 = f_arrdiv24_mux2to1386_xor0 ^ b[19];
  assign f_arrdiv24_fs427_not0 = ~f_arrdiv24_mux2to1386_xor0;
  assign f_arrdiv24_fs427_and0 = f_arrdiv24_fs427_not0 & b[19];
  assign f_arrdiv24_fs427_xor1 = f_arrdiv24_fs426_or0 ^ f_arrdiv24_fs427_xor0;
  assign f_arrdiv24_fs427_not1 = ~f_arrdiv24_fs427_xor0;
  assign f_arrdiv24_fs427_and1 = f_arrdiv24_fs427_not1 & f_arrdiv24_fs426_or0;
  assign f_arrdiv24_fs427_or0 = f_arrdiv24_fs427_and1 | f_arrdiv24_fs427_and0;
  assign f_arrdiv24_fs428_xor0 = f_arrdiv24_mux2to1387_xor0 ^ b[20];
  assign f_arrdiv24_fs428_not0 = ~f_arrdiv24_mux2to1387_xor0;
  assign f_arrdiv24_fs428_and0 = f_arrdiv24_fs428_not0 & b[20];
  assign f_arrdiv24_fs428_xor1 = f_arrdiv24_fs427_or0 ^ f_arrdiv24_fs428_xor0;
  assign f_arrdiv24_fs428_not1 = ~f_arrdiv24_fs428_xor0;
  assign f_arrdiv24_fs428_and1 = f_arrdiv24_fs428_not1 & f_arrdiv24_fs427_or0;
  assign f_arrdiv24_fs428_or0 = f_arrdiv24_fs428_and1 | f_arrdiv24_fs428_and0;
  assign f_arrdiv24_fs429_xor0 = f_arrdiv24_mux2to1388_xor0 ^ b[21];
  assign f_arrdiv24_fs429_not0 = ~f_arrdiv24_mux2to1388_xor0;
  assign f_arrdiv24_fs429_and0 = f_arrdiv24_fs429_not0 & b[21];
  assign f_arrdiv24_fs429_xor1 = f_arrdiv24_fs428_or0 ^ f_arrdiv24_fs429_xor0;
  assign f_arrdiv24_fs429_not1 = ~f_arrdiv24_fs429_xor0;
  assign f_arrdiv24_fs429_and1 = f_arrdiv24_fs429_not1 & f_arrdiv24_fs428_or0;
  assign f_arrdiv24_fs429_or0 = f_arrdiv24_fs429_and1 | f_arrdiv24_fs429_and0;
  assign f_arrdiv24_fs430_xor0 = f_arrdiv24_mux2to1389_xor0 ^ b[22];
  assign f_arrdiv24_fs430_not0 = ~f_arrdiv24_mux2to1389_xor0;
  assign f_arrdiv24_fs430_and0 = f_arrdiv24_fs430_not0 & b[22];
  assign f_arrdiv24_fs430_xor1 = f_arrdiv24_fs429_or0 ^ f_arrdiv24_fs430_xor0;
  assign f_arrdiv24_fs430_not1 = ~f_arrdiv24_fs430_xor0;
  assign f_arrdiv24_fs430_and1 = f_arrdiv24_fs430_not1 & f_arrdiv24_fs429_or0;
  assign f_arrdiv24_fs430_or0 = f_arrdiv24_fs430_and1 | f_arrdiv24_fs430_and0;
  assign f_arrdiv24_fs431_xor0 = f_arrdiv24_mux2to1390_xor0 ^ b[23];
  assign f_arrdiv24_fs431_not0 = ~f_arrdiv24_mux2to1390_xor0;
  assign f_arrdiv24_fs431_and0 = f_arrdiv24_fs431_not0 & b[23];
  assign f_arrdiv24_fs431_xor1 = f_arrdiv24_fs430_or0 ^ f_arrdiv24_fs431_xor0;
  assign f_arrdiv24_fs431_not1 = ~f_arrdiv24_fs431_xor0;
  assign f_arrdiv24_fs431_and1 = f_arrdiv24_fs431_not1 & f_arrdiv24_fs430_or0;
  assign f_arrdiv24_fs431_or0 = f_arrdiv24_fs431_and1 | f_arrdiv24_fs431_and0;
  assign f_arrdiv24_mux2to1391_and0 = a[6] & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1391_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1391_and1 = f_arrdiv24_fs408_xor0 & f_arrdiv24_mux2to1391_not0;
  assign f_arrdiv24_mux2to1391_xor0 = f_arrdiv24_mux2to1391_and0 ^ f_arrdiv24_mux2to1391_and1;
  assign f_arrdiv24_mux2to1392_and0 = f_arrdiv24_mux2to1368_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1392_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1392_and1 = f_arrdiv24_fs409_xor1 & f_arrdiv24_mux2to1392_not0;
  assign f_arrdiv24_mux2to1392_xor0 = f_arrdiv24_mux2to1392_and0 ^ f_arrdiv24_mux2to1392_and1;
  assign f_arrdiv24_mux2to1393_and0 = f_arrdiv24_mux2to1369_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1393_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1393_and1 = f_arrdiv24_fs410_xor1 & f_arrdiv24_mux2to1393_not0;
  assign f_arrdiv24_mux2to1393_xor0 = f_arrdiv24_mux2to1393_and0 ^ f_arrdiv24_mux2to1393_and1;
  assign f_arrdiv24_mux2to1394_and0 = f_arrdiv24_mux2to1370_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1394_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1394_and1 = f_arrdiv24_fs411_xor1 & f_arrdiv24_mux2to1394_not0;
  assign f_arrdiv24_mux2to1394_xor0 = f_arrdiv24_mux2to1394_and0 ^ f_arrdiv24_mux2to1394_and1;
  assign f_arrdiv24_mux2to1395_and0 = f_arrdiv24_mux2to1371_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1395_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1395_and1 = f_arrdiv24_fs412_xor1 & f_arrdiv24_mux2to1395_not0;
  assign f_arrdiv24_mux2to1395_xor0 = f_arrdiv24_mux2to1395_and0 ^ f_arrdiv24_mux2to1395_and1;
  assign f_arrdiv24_mux2to1396_and0 = f_arrdiv24_mux2to1372_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1396_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1396_and1 = f_arrdiv24_fs413_xor1 & f_arrdiv24_mux2to1396_not0;
  assign f_arrdiv24_mux2to1396_xor0 = f_arrdiv24_mux2to1396_and0 ^ f_arrdiv24_mux2to1396_and1;
  assign f_arrdiv24_mux2to1397_and0 = f_arrdiv24_mux2to1373_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1397_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1397_and1 = f_arrdiv24_fs414_xor1 & f_arrdiv24_mux2to1397_not0;
  assign f_arrdiv24_mux2to1397_xor0 = f_arrdiv24_mux2to1397_and0 ^ f_arrdiv24_mux2to1397_and1;
  assign f_arrdiv24_mux2to1398_and0 = f_arrdiv24_mux2to1374_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1398_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1398_and1 = f_arrdiv24_fs415_xor1 & f_arrdiv24_mux2to1398_not0;
  assign f_arrdiv24_mux2to1398_xor0 = f_arrdiv24_mux2to1398_and0 ^ f_arrdiv24_mux2to1398_and1;
  assign f_arrdiv24_mux2to1399_and0 = f_arrdiv24_mux2to1375_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1399_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1399_and1 = f_arrdiv24_fs416_xor1 & f_arrdiv24_mux2to1399_not0;
  assign f_arrdiv24_mux2to1399_xor0 = f_arrdiv24_mux2to1399_and0 ^ f_arrdiv24_mux2to1399_and1;
  assign f_arrdiv24_mux2to1400_and0 = f_arrdiv24_mux2to1376_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1400_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1400_and1 = f_arrdiv24_fs417_xor1 & f_arrdiv24_mux2to1400_not0;
  assign f_arrdiv24_mux2to1400_xor0 = f_arrdiv24_mux2to1400_and0 ^ f_arrdiv24_mux2to1400_and1;
  assign f_arrdiv24_mux2to1401_and0 = f_arrdiv24_mux2to1377_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1401_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1401_and1 = f_arrdiv24_fs418_xor1 & f_arrdiv24_mux2to1401_not0;
  assign f_arrdiv24_mux2to1401_xor0 = f_arrdiv24_mux2to1401_and0 ^ f_arrdiv24_mux2to1401_and1;
  assign f_arrdiv24_mux2to1402_and0 = f_arrdiv24_mux2to1378_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1402_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1402_and1 = f_arrdiv24_fs419_xor1 & f_arrdiv24_mux2to1402_not0;
  assign f_arrdiv24_mux2to1402_xor0 = f_arrdiv24_mux2to1402_and0 ^ f_arrdiv24_mux2to1402_and1;
  assign f_arrdiv24_mux2to1403_and0 = f_arrdiv24_mux2to1379_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1403_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1403_and1 = f_arrdiv24_fs420_xor1 & f_arrdiv24_mux2to1403_not0;
  assign f_arrdiv24_mux2to1403_xor0 = f_arrdiv24_mux2to1403_and0 ^ f_arrdiv24_mux2to1403_and1;
  assign f_arrdiv24_mux2to1404_and0 = f_arrdiv24_mux2to1380_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1404_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1404_and1 = f_arrdiv24_fs421_xor1 & f_arrdiv24_mux2to1404_not0;
  assign f_arrdiv24_mux2to1404_xor0 = f_arrdiv24_mux2to1404_and0 ^ f_arrdiv24_mux2to1404_and1;
  assign f_arrdiv24_mux2to1405_and0 = f_arrdiv24_mux2to1381_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1405_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1405_and1 = f_arrdiv24_fs422_xor1 & f_arrdiv24_mux2to1405_not0;
  assign f_arrdiv24_mux2to1405_xor0 = f_arrdiv24_mux2to1405_and0 ^ f_arrdiv24_mux2to1405_and1;
  assign f_arrdiv24_mux2to1406_and0 = f_arrdiv24_mux2to1382_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1406_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1406_and1 = f_arrdiv24_fs423_xor1 & f_arrdiv24_mux2to1406_not0;
  assign f_arrdiv24_mux2to1406_xor0 = f_arrdiv24_mux2to1406_and0 ^ f_arrdiv24_mux2to1406_and1;
  assign f_arrdiv24_mux2to1407_and0 = f_arrdiv24_mux2to1383_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1407_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1407_and1 = f_arrdiv24_fs424_xor1 & f_arrdiv24_mux2to1407_not0;
  assign f_arrdiv24_mux2to1407_xor0 = f_arrdiv24_mux2to1407_and0 ^ f_arrdiv24_mux2to1407_and1;
  assign f_arrdiv24_mux2to1408_and0 = f_arrdiv24_mux2to1384_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1408_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1408_and1 = f_arrdiv24_fs425_xor1 & f_arrdiv24_mux2to1408_not0;
  assign f_arrdiv24_mux2to1408_xor0 = f_arrdiv24_mux2to1408_and0 ^ f_arrdiv24_mux2to1408_and1;
  assign f_arrdiv24_mux2to1409_and0 = f_arrdiv24_mux2to1385_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1409_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1409_and1 = f_arrdiv24_fs426_xor1 & f_arrdiv24_mux2to1409_not0;
  assign f_arrdiv24_mux2to1409_xor0 = f_arrdiv24_mux2to1409_and0 ^ f_arrdiv24_mux2to1409_and1;
  assign f_arrdiv24_mux2to1410_and0 = f_arrdiv24_mux2to1386_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1410_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1410_and1 = f_arrdiv24_fs427_xor1 & f_arrdiv24_mux2to1410_not0;
  assign f_arrdiv24_mux2to1410_xor0 = f_arrdiv24_mux2to1410_and0 ^ f_arrdiv24_mux2to1410_and1;
  assign f_arrdiv24_mux2to1411_and0 = f_arrdiv24_mux2to1387_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1411_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1411_and1 = f_arrdiv24_fs428_xor1 & f_arrdiv24_mux2to1411_not0;
  assign f_arrdiv24_mux2to1411_xor0 = f_arrdiv24_mux2to1411_and0 ^ f_arrdiv24_mux2to1411_and1;
  assign f_arrdiv24_mux2to1412_and0 = f_arrdiv24_mux2to1388_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1412_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1412_and1 = f_arrdiv24_fs429_xor1 & f_arrdiv24_mux2to1412_not0;
  assign f_arrdiv24_mux2to1412_xor0 = f_arrdiv24_mux2to1412_and0 ^ f_arrdiv24_mux2to1412_and1;
  assign f_arrdiv24_mux2to1413_and0 = f_arrdiv24_mux2to1389_xor0 & f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1413_not0 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_mux2to1413_and1 = f_arrdiv24_fs430_xor1 & f_arrdiv24_mux2to1413_not0;
  assign f_arrdiv24_mux2to1413_xor0 = f_arrdiv24_mux2to1413_and0 ^ f_arrdiv24_mux2to1413_and1;
  assign f_arrdiv24_not17 = ~f_arrdiv24_fs431_or0;
  assign f_arrdiv24_fs432_xor0 = a[5] ^ b[0];
  assign f_arrdiv24_fs432_not0 = ~a[5];
  assign f_arrdiv24_fs432_and0 = f_arrdiv24_fs432_not0 & b[0];
  assign f_arrdiv24_fs432_not1 = ~f_arrdiv24_fs432_xor0;
  assign f_arrdiv24_fs433_xor0 = f_arrdiv24_mux2to1391_xor0 ^ b[1];
  assign f_arrdiv24_fs433_not0 = ~f_arrdiv24_mux2to1391_xor0;
  assign f_arrdiv24_fs433_and0 = f_arrdiv24_fs433_not0 & b[1];
  assign f_arrdiv24_fs433_xor1 = f_arrdiv24_fs432_and0 ^ f_arrdiv24_fs433_xor0;
  assign f_arrdiv24_fs433_not1 = ~f_arrdiv24_fs433_xor0;
  assign f_arrdiv24_fs433_and1 = f_arrdiv24_fs433_not1 & f_arrdiv24_fs432_and0;
  assign f_arrdiv24_fs433_or0 = f_arrdiv24_fs433_and1 | f_arrdiv24_fs433_and0;
  assign f_arrdiv24_fs434_xor0 = f_arrdiv24_mux2to1392_xor0 ^ b[2];
  assign f_arrdiv24_fs434_not0 = ~f_arrdiv24_mux2to1392_xor0;
  assign f_arrdiv24_fs434_and0 = f_arrdiv24_fs434_not0 & b[2];
  assign f_arrdiv24_fs434_xor1 = f_arrdiv24_fs433_or0 ^ f_arrdiv24_fs434_xor0;
  assign f_arrdiv24_fs434_not1 = ~f_arrdiv24_fs434_xor0;
  assign f_arrdiv24_fs434_and1 = f_arrdiv24_fs434_not1 & f_arrdiv24_fs433_or0;
  assign f_arrdiv24_fs434_or0 = f_arrdiv24_fs434_and1 | f_arrdiv24_fs434_and0;
  assign f_arrdiv24_fs435_xor0 = f_arrdiv24_mux2to1393_xor0 ^ b[3];
  assign f_arrdiv24_fs435_not0 = ~f_arrdiv24_mux2to1393_xor0;
  assign f_arrdiv24_fs435_and0 = f_arrdiv24_fs435_not0 & b[3];
  assign f_arrdiv24_fs435_xor1 = f_arrdiv24_fs434_or0 ^ f_arrdiv24_fs435_xor0;
  assign f_arrdiv24_fs435_not1 = ~f_arrdiv24_fs435_xor0;
  assign f_arrdiv24_fs435_and1 = f_arrdiv24_fs435_not1 & f_arrdiv24_fs434_or0;
  assign f_arrdiv24_fs435_or0 = f_arrdiv24_fs435_and1 | f_arrdiv24_fs435_and0;
  assign f_arrdiv24_fs436_xor0 = f_arrdiv24_mux2to1394_xor0 ^ b[4];
  assign f_arrdiv24_fs436_not0 = ~f_arrdiv24_mux2to1394_xor0;
  assign f_arrdiv24_fs436_and0 = f_arrdiv24_fs436_not0 & b[4];
  assign f_arrdiv24_fs436_xor1 = f_arrdiv24_fs435_or0 ^ f_arrdiv24_fs436_xor0;
  assign f_arrdiv24_fs436_not1 = ~f_arrdiv24_fs436_xor0;
  assign f_arrdiv24_fs436_and1 = f_arrdiv24_fs436_not1 & f_arrdiv24_fs435_or0;
  assign f_arrdiv24_fs436_or0 = f_arrdiv24_fs436_and1 | f_arrdiv24_fs436_and0;
  assign f_arrdiv24_fs437_xor0 = f_arrdiv24_mux2to1395_xor0 ^ b[5];
  assign f_arrdiv24_fs437_not0 = ~f_arrdiv24_mux2to1395_xor0;
  assign f_arrdiv24_fs437_and0 = f_arrdiv24_fs437_not0 & b[5];
  assign f_arrdiv24_fs437_xor1 = f_arrdiv24_fs436_or0 ^ f_arrdiv24_fs437_xor0;
  assign f_arrdiv24_fs437_not1 = ~f_arrdiv24_fs437_xor0;
  assign f_arrdiv24_fs437_and1 = f_arrdiv24_fs437_not1 & f_arrdiv24_fs436_or0;
  assign f_arrdiv24_fs437_or0 = f_arrdiv24_fs437_and1 | f_arrdiv24_fs437_and0;
  assign f_arrdiv24_fs438_xor0 = f_arrdiv24_mux2to1396_xor0 ^ b[6];
  assign f_arrdiv24_fs438_not0 = ~f_arrdiv24_mux2to1396_xor0;
  assign f_arrdiv24_fs438_and0 = f_arrdiv24_fs438_not0 & b[6];
  assign f_arrdiv24_fs438_xor1 = f_arrdiv24_fs437_or0 ^ f_arrdiv24_fs438_xor0;
  assign f_arrdiv24_fs438_not1 = ~f_arrdiv24_fs438_xor0;
  assign f_arrdiv24_fs438_and1 = f_arrdiv24_fs438_not1 & f_arrdiv24_fs437_or0;
  assign f_arrdiv24_fs438_or0 = f_arrdiv24_fs438_and1 | f_arrdiv24_fs438_and0;
  assign f_arrdiv24_fs439_xor0 = f_arrdiv24_mux2to1397_xor0 ^ b[7];
  assign f_arrdiv24_fs439_not0 = ~f_arrdiv24_mux2to1397_xor0;
  assign f_arrdiv24_fs439_and0 = f_arrdiv24_fs439_not0 & b[7];
  assign f_arrdiv24_fs439_xor1 = f_arrdiv24_fs438_or0 ^ f_arrdiv24_fs439_xor0;
  assign f_arrdiv24_fs439_not1 = ~f_arrdiv24_fs439_xor0;
  assign f_arrdiv24_fs439_and1 = f_arrdiv24_fs439_not1 & f_arrdiv24_fs438_or0;
  assign f_arrdiv24_fs439_or0 = f_arrdiv24_fs439_and1 | f_arrdiv24_fs439_and0;
  assign f_arrdiv24_fs440_xor0 = f_arrdiv24_mux2to1398_xor0 ^ b[8];
  assign f_arrdiv24_fs440_not0 = ~f_arrdiv24_mux2to1398_xor0;
  assign f_arrdiv24_fs440_and0 = f_arrdiv24_fs440_not0 & b[8];
  assign f_arrdiv24_fs440_xor1 = f_arrdiv24_fs439_or0 ^ f_arrdiv24_fs440_xor0;
  assign f_arrdiv24_fs440_not1 = ~f_arrdiv24_fs440_xor0;
  assign f_arrdiv24_fs440_and1 = f_arrdiv24_fs440_not1 & f_arrdiv24_fs439_or0;
  assign f_arrdiv24_fs440_or0 = f_arrdiv24_fs440_and1 | f_arrdiv24_fs440_and0;
  assign f_arrdiv24_fs441_xor0 = f_arrdiv24_mux2to1399_xor0 ^ b[9];
  assign f_arrdiv24_fs441_not0 = ~f_arrdiv24_mux2to1399_xor0;
  assign f_arrdiv24_fs441_and0 = f_arrdiv24_fs441_not0 & b[9];
  assign f_arrdiv24_fs441_xor1 = f_arrdiv24_fs440_or0 ^ f_arrdiv24_fs441_xor0;
  assign f_arrdiv24_fs441_not1 = ~f_arrdiv24_fs441_xor0;
  assign f_arrdiv24_fs441_and1 = f_arrdiv24_fs441_not1 & f_arrdiv24_fs440_or0;
  assign f_arrdiv24_fs441_or0 = f_arrdiv24_fs441_and1 | f_arrdiv24_fs441_and0;
  assign f_arrdiv24_fs442_xor0 = f_arrdiv24_mux2to1400_xor0 ^ b[10];
  assign f_arrdiv24_fs442_not0 = ~f_arrdiv24_mux2to1400_xor0;
  assign f_arrdiv24_fs442_and0 = f_arrdiv24_fs442_not0 & b[10];
  assign f_arrdiv24_fs442_xor1 = f_arrdiv24_fs441_or0 ^ f_arrdiv24_fs442_xor0;
  assign f_arrdiv24_fs442_not1 = ~f_arrdiv24_fs442_xor0;
  assign f_arrdiv24_fs442_and1 = f_arrdiv24_fs442_not1 & f_arrdiv24_fs441_or0;
  assign f_arrdiv24_fs442_or0 = f_arrdiv24_fs442_and1 | f_arrdiv24_fs442_and0;
  assign f_arrdiv24_fs443_xor0 = f_arrdiv24_mux2to1401_xor0 ^ b[11];
  assign f_arrdiv24_fs443_not0 = ~f_arrdiv24_mux2to1401_xor0;
  assign f_arrdiv24_fs443_and0 = f_arrdiv24_fs443_not0 & b[11];
  assign f_arrdiv24_fs443_xor1 = f_arrdiv24_fs442_or0 ^ f_arrdiv24_fs443_xor0;
  assign f_arrdiv24_fs443_not1 = ~f_arrdiv24_fs443_xor0;
  assign f_arrdiv24_fs443_and1 = f_arrdiv24_fs443_not1 & f_arrdiv24_fs442_or0;
  assign f_arrdiv24_fs443_or0 = f_arrdiv24_fs443_and1 | f_arrdiv24_fs443_and0;
  assign f_arrdiv24_fs444_xor0 = f_arrdiv24_mux2to1402_xor0 ^ b[12];
  assign f_arrdiv24_fs444_not0 = ~f_arrdiv24_mux2to1402_xor0;
  assign f_arrdiv24_fs444_and0 = f_arrdiv24_fs444_not0 & b[12];
  assign f_arrdiv24_fs444_xor1 = f_arrdiv24_fs443_or0 ^ f_arrdiv24_fs444_xor0;
  assign f_arrdiv24_fs444_not1 = ~f_arrdiv24_fs444_xor0;
  assign f_arrdiv24_fs444_and1 = f_arrdiv24_fs444_not1 & f_arrdiv24_fs443_or0;
  assign f_arrdiv24_fs444_or0 = f_arrdiv24_fs444_and1 | f_arrdiv24_fs444_and0;
  assign f_arrdiv24_fs445_xor0 = f_arrdiv24_mux2to1403_xor0 ^ b[13];
  assign f_arrdiv24_fs445_not0 = ~f_arrdiv24_mux2to1403_xor0;
  assign f_arrdiv24_fs445_and0 = f_arrdiv24_fs445_not0 & b[13];
  assign f_arrdiv24_fs445_xor1 = f_arrdiv24_fs444_or0 ^ f_arrdiv24_fs445_xor0;
  assign f_arrdiv24_fs445_not1 = ~f_arrdiv24_fs445_xor0;
  assign f_arrdiv24_fs445_and1 = f_arrdiv24_fs445_not1 & f_arrdiv24_fs444_or0;
  assign f_arrdiv24_fs445_or0 = f_arrdiv24_fs445_and1 | f_arrdiv24_fs445_and0;
  assign f_arrdiv24_fs446_xor0 = f_arrdiv24_mux2to1404_xor0 ^ b[14];
  assign f_arrdiv24_fs446_not0 = ~f_arrdiv24_mux2to1404_xor0;
  assign f_arrdiv24_fs446_and0 = f_arrdiv24_fs446_not0 & b[14];
  assign f_arrdiv24_fs446_xor1 = f_arrdiv24_fs445_or0 ^ f_arrdiv24_fs446_xor0;
  assign f_arrdiv24_fs446_not1 = ~f_arrdiv24_fs446_xor0;
  assign f_arrdiv24_fs446_and1 = f_arrdiv24_fs446_not1 & f_arrdiv24_fs445_or0;
  assign f_arrdiv24_fs446_or0 = f_arrdiv24_fs446_and1 | f_arrdiv24_fs446_and0;
  assign f_arrdiv24_fs447_xor0 = f_arrdiv24_mux2to1405_xor0 ^ b[15];
  assign f_arrdiv24_fs447_not0 = ~f_arrdiv24_mux2to1405_xor0;
  assign f_arrdiv24_fs447_and0 = f_arrdiv24_fs447_not0 & b[15];
  assign f_arrdiv24_fs447_xor1 = f_arrdiv24_fs446_or0 ^ f_arrdiv24_fs447_xor0;
  assign f_arrdiv24_fs447_not1 = ~f_arrdiv24_fs447_xor0;
  assign f_arrdiv24_fs447_and1 = f_arrdiv24_fs447_not1 & f_arrdiv24_fs446_or0;
  assign f_arrdiv24_fs447_or0 = f_arrdiv24_fs447_and1 | f_arrdiv24_fs447_and0;
  assign f_arrdiv24_fs448_xor0 = f_arrdiv24_mux2to1406_xor0 ^ b[16];
  assign f_arrdiv24_fs448_not0 = ~f_arrdiv24_mux2to1406_xor0;
  assign f_arrdiv24_fs448_and0 = f_arrdiv24_fs448_not0 & b[16];
  assign f_arrdiv24_fs448_xor1 = f_arrdiv24_fs447_or0 ^ f_arrdiv24_fs448_xor0;
  assign f_arrdiv24_fs448_not1 = ~f_arrdiv24_fs448_xor0;
  assign f_arrdiv24_fs448_and1 = f_arrdiv24_fs448_not1 & f_arrdiv24_fs447_or0;
  assign f_arrdiv24_fs448_or0 = f_arrdiv24_fs448_and1 | f_arrdiv24_fs448_and0;
  assign f_arrdiv24_fs449_xor0 = f_arrdiv24_mux2to1407_xor0 ^ b[17];
  assign f_arrdiv24_fs449_not0 = ~f_arrdiv24_mux2to1407_xor0;
  assign f_arrdiv24_fs449_and0 = f_arrdiv24_fs449_not0 & b[17];
  assign f_arrdiv24_fs449_xor1 = f_arrdiv24_fs448_or0 ^ f_arrdiv24_fs449_xor0;
  assign f_arrdiv24_fs449_not1 = ~f_arrdiv24_fs449_xor0;
  assign f_arrdiv24_fs449_and1 = f_arrdiv24_fs449_not1 & f_arrdiv24_fs448_or0;
  assign f_arrdiv24_fs449_or0 = f_arrdiv24_fs449_and1 | f_arrdiv24_fs449_and0;
  assign f_arrdiv24_fs450_xor0 = f_arrdiv24_mux2to1408_xor0 ^ b[18];
  assign f_arrdiv24_fs450_not0 = ~f_arrdiv24_mux2to1408_xor0;
  assign f_arrdiv24_fs450_and0 = f_arrdiv24_fs450_not0 & b[18];
  assign f_arrdiv24_fs450_xor1 = f_arrdiv24_fs449_or0 ^ f_arrdiv24_fs450_xor0;
  assign f_arrdiv24_fs450_not1 = ~f_arrdiv24_fs450_xor0;
  assign f_arrdiv24_fs450_and1 = f_arrdiv24_fs450_not1 & f_arrdiv24_fs449_or0;
  assign f_arrdiv24_fs450_or0 = f_arrdiv24_fs450_and1 | f_arrdiv24_fs450_and0;
  assign f_arrdiv24_fs451_xor0 = f_arrdiv24_mux2to1409_xor0 ^ b[19];
  assign f_arrdiv24_fs451_not0 = ~f_arrdiv24_mux2to1409_xor0;
  assign f_arrdiv24_fs451_and0 = f_arrdiv24_fs451_not0 & b[19];
  assign f_arrdiv24_fs451_xor1 = f_arrdiv24_fs450_or0 ^ f_arrdiv24_fs451_xor0;
  assign f_arrdiv24_fs451_not1 = ~f_arrdiv24_fs451_xor0;
  assign f_arrdiv24_fs451_and1 = f_arrdiv24_fs451_not1 & f_arrdiv24_fs450_or0;
  assign f_arrdiv24_fs451_or0 = f_arrdiv24_fs451_and1 | f_arrdiv24_fs451_and0;
  assign f_arrdiv24_fs452_xor0 = f_arrdiv24_mux2to1410_xor0 ^ b[20];
  assign f_arrdiv24_fs452_not0 = ~f_arrdiv24_mux2to1410_xor0;
  assign f_arrdiv24_fs452_and0 = f_arrdiv24_fs452_not0 & b[20];
  assign f_arrdiv24_fs452_xor1 = f_arrdiv24_fs451_or0 ^ f_arrdiv24_fs452_xor0;
  assign f_arrdiv24_fs452_not1 = ~f_arrdiv24_fs452_xor0;
  assign f_arrdiv24_fs452_and1 = f_arrdiv24_fs452_not1 & f_arrdiv24_fs451_or0;
  assign f_arrdiv24_fs452_or0 = f_arrdiv24_fs452_and1 | f_arrdiv24_fs452_and0;
  assign f_arrdiv24_fs453_xor0 = f_arrdiv24_mux2to1411_xor0 ^ b[21];
  assign f_arrdiv24_fs453_not0 = ~f_arrdiv24_mux2to1411_xor0;
  assign f_arrdiv24_fs453_and0 = f_arrdiv24_fs453_not0 & b[21];
  assign f_arrdiv24_fs453_xor1 = f_arrdiv24_fs452_or0 ^ f_arrdiv24_fs453_xor0;
  assign f_arrdiv24_fs453_not1 = ~f_arrdiv24_fs453_xor0;
  assign f_arrdiv24_fs453_and1 = f_arrdiv24_fs453_not1 & f_arrdiv24_fs452_or0;
  assign f_arrdiv24_fs453_or0 = f_arrdiv24_fs453_and1 | f_arrdiv24_fs453_and0;
  assign f_arrdiv24_fs454_xor0 = f_arrdiv24_mux2to1412_xor0 ^ b[22];
  assign f_arrdiv24_fs454_not0 = ~f_arrdiv24_mux2to1412_xor0;
  assign f_arrdiv24_fs454_and0 = f_arrdiv24_fs454_not0 & b[22];
  assign f_arrdiv24_fs454_xor1 = f_arrdiv24_fs453_or0 ^ f_arrdiv24_fs454_xor0;
  assign f_arrdiv24_fs454_not1 = ~f_arrdiv24_fs454_xor0;
  assign f_arrdiv24_fs454_and1 = f_arrdiv24_fs454_not1 & f_arrdiv24_fs453_or0;
  assign f_arrdiv24_fs454_or0 = f_arrdiv24_fs454_and1 | f_arrdiv24_fs454_and0;
  assign f_arrdiv24_fs455_xor0 = f_arrdiv24_mux2to1413_xor0 ^ b[23];
  assign f_arrdiv24_fs455_not0 = ~f_arrdiv24_mux2to1413_xor0;
  assign f_arrdiv24_fs455_and0 = f_arrdiv24_fs455_not0 & b[23];
  assign f_arrdiv24_fs455_xor1 = f_arrdiv24_fs454_or0 ^ f_arrdiv24_fs455_xor0;
  assign f_arrdiv24_fs455_not1 = ~f_arrdiv24_fs455_xor0;
  assign f_arrdiv24_fs455_and1 = f_arrdiv24_fs455_not1 & f_arrdiv24_fs454_or0;
  assign f_arrdiv24_fs455_or0 = f_arrdiv24_fs455_and1 | f_arrdiv24_fs455_and0;
  assign f_arrdiv24_mux2to1414_and0 = a[5] & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1414_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1414_and1 = f_arrdiv24_fs432_xor0 & f_arrdiv24_mux2to1414_not0;
  assign f_arrdiv24_mux2to1414_xor0 = f_arrdiv24_mux2to1414_and0 ^ f_arrdiv24_mux2to1414_and1;
  assign f_arrdiv24_mux2to1415_and0 = f_arrdiv24_mux2to1391_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1415_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1415_and1 = f_arrdiv24_fs433_xor1 & f_arrdiv24_mux2to1415_not0;
  assign f_arrdiv24_mux2to1415_xor0 = f_arrdiv24_mux2to1415_and0 ^ f_arrdiv24_mux2to1415_and1;
  assign f_arrdiv24_mux2to1416_and0 = f_arrdiv24_mux2to1392_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1416_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1416_and1 = f_arrdiv24_fs434_xor1 & f_arrdiv24_mux2to1416_not0;
  assign f_arrdiv24_mux2to1416_xor0 = f_arrdiv24_mux2to1416_and0 ^ f_arrdiv24_mux2to1416_and1;
  assign f_arrdiv24_mux2to1417_and0 = f_arrdiv24_mux2to1393_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1417_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1417_and1 = f_arrdiv24_fs435_xor1 & f_arrdiv24_mux2to1417_not0;
  assign f_arrdiv24_mux2to1417_xor0 = f_arrdiv24_mux2to1417_and0 ^ f_arrdiv24_mux2to1417_and1;
  assign f_arrdiv24_mux2to1418_and0 = f_arrdiv24_mux2to1394_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1418_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1418_and1 = f_arrdiv24_fs436_xor1 & f_arrdiv24_mux2to1418_not0;
  assign f_arrdiv24_mux2to1418_xor0 = f_arrdiv24_mux2to1418_and0 ^ f_arrdiv24_mux2to1418_and1;
  assign f_arrdiv24_mux2to1419_and0 = f_arrdiv24_mux2to1395_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1419_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1419_and1 = f_arrdiv24_fs437_xor1 & f_arrdiv24_mux2to1419_not0;
  assign f_arrdiv24_mux2to1419_xor0 = f_arrdiv24_mux2to1419_and0 ^ f_arrdiv24_mux2to1419_and1;
  assign f_arrdiv24_mux2to1420_and0 = f_arrdiv24_mux2to1396_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1420_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1420_and1 = f_arrdiv24_fs438_xor1 & f_arrdiv24_mux2to1420_not0;
  assign f_arrdiv24_mux2to1420_xor0 = f_arrdiv24_mux2to1420_and0 ^ f_arrdiv24_mux2to1420_and1;
  assign f_arrdiv24_mux2to1421_and0 = f_arrdiv24_mux2to1397_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1421_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1421_and1 = f_arrdiv24_fs439_xor1 & f_arrdiv24_mux2to1421_not0;
  assign f_arrdiv24_mux2to1421_xor0 = f_arrdiv24_mux2to1421_and0 ^ f_arrdiv24_mux2to1421_and1;
  assign f_arrdiv24_mux2to1422_and0 = f_arrdiv24_mux2to1398_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1422_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1422_and1 = f_arrdiv24_fs440_xor1 & f_arrdiv24_mux2to1422_not0;
  assign f_arrdiv24_mux2to1422_xor0 = f_arrdiv24_mux2to1422_and0 ^ f_arrdiv24_mux2to1422_and1;
  assign f_arrdiv24_mux2to1423_and0 = f_arrdiv24_mux2to1399_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1423_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1423_and1 = f_arrdiv24_fs441_xor1 & f_arrdiv24_mux2to1423_not0;
  assign f_arrdiv24_mux2to1423_xor0 = f_arrdiv24_mux2to1423_and0 ^ f_arrdiv24_mux2to1423_and1;
  assign f_arrdiv24_mux2to1424_and0 = f_arrdiv24_mux2to1400_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1424_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1424_and1 = f_arrdiv24_fs442_xor1 & f_arrdiv24_mux2to1424_not0;
  assign f_arrdiv24_mux2to1424_xor0 = f_arrdiv24_mux2to1424_and0 ^ f_arrdiv24_mux2to1424_and1;
  assign f_arrdiv24_mux2to1425_and0 = f_arrdiv24_mux2to1401_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1425_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1425_and1 = f_arrdiv24_fs443_xor1 & f_arrdiv24_mux2to1425_not0;
  assign f_arrdiv24_mux2to1425_xor0 = f_arrdiv24_mux2to1425_and0 ^ f_arrdiv24_mux2to1425_and1;
  assign f_arrdiv24_mux2to1426_and0 = f_arrdiv24_mux2to1402_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1426_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1426_and1 = f_arrdiv24_fs444_xor1 & f_arrdiv24_mux2to1426_not0;
  assign f_arrdiv24_mux2to1426_xor0 = f_arrdiv24_mux2to1426_and0 ^ f_arrdiv24_mux2to1426_and1;
  assign f_arrdiv24_mux2to1427_and0 = f_arrdiv24_mux2to1403_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1427_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1427_and1 = f_arrdiv24_fs445_xor1 & f_arrdiv24_mux2to1427_not0;
  assign f_arrdiv24_mux2to1427_xor0 = f_arrdiv24_mux2to1427_and0 ^ f_arrdiv24_mux2to1427_and1;
  assign f_arrdiv24_mux2to1428_and0 = f_arrdiv24_mux2to1404_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1428_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1428_and1 = f_arrdiv24_fs446_xor1 & f_arrdiv24_mux2to1428_not0;
  assign f_arrdiv24_mux2to1428_xor0 = f_arrdiv24_mux2to1428_and0 ^ f_arrdiv24_mux2to1428_and1;
  assign f_arrdiv24_mux2to1429_and0 = f_arrdiv24_mux2to1405_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1429_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1429_and1 = f_arrdiv24_fs447_xor1 & f_arrdiv24_mux2to1429_not0;
  assign f_arrdiv24_mux2to1429_xor0 = f_arrdiv24_mux2to1429_and0 ^ f_arrdiv24_mux2to1429_and1;
  assign f_arrdiv24_mux2to1430_and0 = f_arrdiv24_mux2to1406_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1430_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1430_and1 = f_arrdiv24_fs448_xor1 & f_arrdiv24_mux2to1430_not0;
  assign f_arrdiv24_mux2to1430_xor0 = f_arrdiv24_mux2to1430_and0 ^ f_arrdiv24_mux2to1430_and1;
  assign f_arrdiv24_mux2to1431_and0 = f_arrdiv24_mux2to1407_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1431_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1431_and1 = f_arrdiv24_fs449_xor1 & f_arrdiv24_mux2to1431_not0;
  assign f_arrdiv24_mux2to1431_xor0 = f_arrdiv24_mux2to1431_and0 ^ f_arrdiv24_mux2to1431_and1;
  assign f_arrdiv24_mux2to1432_and0 = f_arrdiv24_mux2to1408_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1432_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1432_and1 = f_arrdiv24_fs450_xor1 & f_arrdiv24_mux2to1432_not0;
  assign f_arrdiv24_mux2to1432_xor0 = f_arrdiv24_mux2to1432_and0 ^ f_arrdiv24_mux2to1432_and1;
  assign f_arrdiv24_mux2to1433_and0 = f_arrdiv24_mux2to1409_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1433_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1433_and1 = f_arrdiv24_fs451_xor1 & f_arrdiv24_mux2to1433_not0;
  assign f_arrdiv24_mux2to1433_xor0 = f_arrdiv24_mux2to1433_and0 ^ f_arrdiv24_mux2to1433_and1;
  assign f_arrdiv24_mux2to1434_and0 = f_arrdiv24_mux2to1410_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1434_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1434_and1 = f_arrdiv24_fs452_xor1 & f_arrdiv24_mux2to1434_not0;
  assign f_arrdiv24_mux2to1434_xor0 = f_arrdiv24_mux2to1434_and0 ^ f_arrdiv24_mux2to1434_and1;
  assign f_arrdiv24_mux2to1435_and0 = f_arrdiv24_mux2to1411_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1435_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1435_and1 = f_arrdiv24_fs453_xor1 & f_arrdiv24_mux2to1435_not0;
  assign f_arrdiv24_mux2to1435_xor0 = f_arrdiv24_mux2to1435_and0 ^ f_arrdiv24_mux2to1435_and1;
  assign f_arrdiv24_mux2to1436_and0 = f_arrdiv24_mux2to1412_xor0 & f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1436_not0 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_mux2to1436_and1 = f_arrdiv24_fs454_xor1 & f_arrdiv24_mux2to1436_not0;
  assign f_arrdiv24_mux2to1436_xor0 = f_arrdiv24_mux2to1436_and0 ^ f_arrdiv24_mux2to1436_and1;
  assign f_arrdiv24_not18 = ~f_arrdiv24_fs455_or0;
  assign f_arrdiv24_fs456_xor0 = a[4] ^ b[0];
  assign f_arrdiv24_fs456_not0 = ~a[4];
  assign f_arrdiv24_fs456_and0 = f_arrdiv24_fs456_not0 & b[0];
  assign f_arrdiv24_fs456_not1 = ~f_arrdiv24_fs456_xor0;
  assign f_arrdiv24_fs457_xor0 = f_arrdiv24_mux2to1414_xor0 ^ b[1];
  assign f_arrdiv24_fs457_not0 = ~f_arrdiv24_mux2to1414_xor0;
  assign f_arrdiv24_fs457_and0 = f_arrdiv24_fs457_not0 & b[1];
  assign f_arrdiv24_fs457_xor1 = f_arrdiv24_fs456_and0 ^ f_arrdiv24_fs457_xor0;
  assign f_arrdiv24_fs457_not1 = ~f_arrdiv24_fs457_xor0;
  assign f_arrdiv24_fs457_and1 = f_arrdiv24_fs457_not1 & f_arrdiv24_fs456_and0;
  assign f_arrdiv24_fs457_or0 = f_arrdiv24_fs457_and1 | f_arrdiv24_fs457_and0;
  assign f_arrdiv24_fs458_xor0 = f_arrdiv24_mux2to1415_xor0 ^ b[2];
  assign f_arrdiv24_fs458_not0 = ~f_arrdiv24_mux2to1415_xor0;
  assign f_arrdiv24_fs458_and0 = f_arrdiv24_fs458_not0 & b[2];
  assign f_arrdiv24_fs458_xor1 = f_arrdiv24_fs457_or0 ^ f_arrdiv24_fs458_xor0;
  assign f_arrdiv24_fs458_not1 = ~f_arrdiv24_fs458_xor0;
  assign f_arrdiv24_fs458_and1 = f_arrdiv24_fs458_not1 & f_arrdiv24_fs457_or0;
  assign f_arrdiv24_fs458_or0 = f_arrdiv24_fs458_and1 | f_arrdiv24_fs458_and0;
  assign f_arrdiv24_fs459_xor0 = f_arrdiv24_mux2to1416_xor0 ^ b[3];
  assign f_arrdiv24_fs459_not0 = ~f_arrdiv24_mux2to1416_xor0;
  assign f_arrdiv24_fs459_and0 = f_arrdiv24_fs459_not0 & b[3];
  assign f_arrdiv24_fs459_xor1 = f_arrdiv24_fs458_or0 ^ f_arrdiv24_fs459_xor0;
  assign f_arrdiv24_fs459_not1 = ~f_arrdiv24_fs459_xor0;
  assign f_arrdiv24_fs459_and1 = f_arrdiv24_fs459_not1 & f_arrdiv24_fs458_or0;
  assign f_arrdiv24_fs459_or0 = f_arrdiv24_fs459_and1 | f_arrdiv24_fs459_and0;
  assign f_arrdiv24_fs460_xor0 = f_arrdiv24_mux2to1417_xor0 ^ b[4];
  assign f_arrdiv24_fs460_not0 = ~f_arrdiv24_mux2to1417_xor0;
  assign f_arrdiv24_fs460_and0 = f_arrdiv24_fs460_not0 & b[4];
  assign f_arrdiv24_fs460_xor1 = f_arrdiv24_fs459_or0 ^ f_arrdiv24_fs460_xor0;
  assign f_arrdiv24_fs460_not1 = ~f_arrdiv24_fs460_xor0;
  assign f_arrdiv24_fs460_and1 = f_arrdiv24_fs460_not1 & f_arrdiv24_fs459_or0;
  assign f_arrdiv24_fs460_or0 = f_arrdiv24_fs460_and1 | f_arrdiv24_fs460_and0;
  assign f_arrdiv24_fs461_xor0 = f_arrdiv24_mux2to1418_xor0 ^ b[5];
  assign f_arrdiv24_fs461_not0 = ~f_arrdiv24_mux2to1418_xor0;
  assign f_arrdiv24_fs461_and0 = f_arrdiv24_fs461_not0 & b[5];
  assign f_arrdiv24_fs461_xor1 = f_arrdiv24_fs460_or0 ^ f_arrdiv24_fs461_xor0;
  assign f_arrdiv24_fs461_not1 = ~f_arrdiv24_fs461_xor0;
  assign f_arrdiv24_fs461_and1 = f_arrdiv24_fs461_not1 & f_arrdiv24_fs460_or0;
  assign f_arrdiv24_fs461_or0 = f_arrdiv24_fs461_and1 | f_arrdiv24_fs461_and0;
  assign f_arrdiv24_fs462_xor0 = f_arrdiv24_mux2to1419_xor0 ^ b[6];
  assign f_arrdiv24_fs462_not0 = ~f_arrdiv24_mux2to1419_xor0;
  assign f_arrdiv24_fs462_and0 = f_arrdiv24_fs462_not0 & b[6];
  assign f_arrdiv24_fs462_xor1 = f_arrdiv24_fs461_or0 ^ f_arrdiv24_fs462_xor0;
  assign f_arrdiv24_fs462_not1 = ~f_arrdiv24_fs462_xor0;
  assign f_arrdiv24_fs462_and1 = f_arrdiv24_fs462_not1 & f_arrdiv24_fs461_or0;
  assign f_arrdiv24_fs462_or0 = f_arrdiv24_fs462_and1 | f_arrdiv24_fs462_and0;
  assign f_arrdiv24_fs463_xor0 = f_arrdiv24_mux2to1420_xor0 ^ b[7];
  assign f_arrdiv24_fs463_not0 = ~f_arrdiv24_mux2to1420_xor0;
  assign f_arrdiv24_fs463_and0 = f_arrdiv24_fs463_not0 & b[7];
  assign f_arrdiv24_fs463_xor1 = f_arrdiv24_fs462_or0 ^ f_arrdiv24_fs463_xor0;
  assign f_arrdiv24_fs463_not1 = ~f_arrdiv24_fs463_xor0;
  assign f_arrdiv24_fs463_and1 = f_arrdiv24_fs463_not1 & f_arrdiv24_fs462_or0;
  assign f_arrdiv24_fs463_or0 = f_arrdiv24_fs463_and1 | f_arrdiv24_fs463_and0;
  assign f_arrdiv24_fs464_xor0 = f_arrdiv24_mux2to1421_xor0 ^ b[8];
  assign f_arrdiv24_fs464_not0 = ~f_arrdiv24_mux2to1421_xor0;
  assign f_arrdiv24_fs464_and0 = f_arrdiv24_fs464_not0 & b[8];
  assign f_arrdiv24_fs464_xor1 = f_arrdiv24_fs463_or0 ^ f_arrdiv24_fs464_xor0;
  assign f_arrdiv24_fs464_not1 = ~f_arrdiv24_fs464_xor0;
  assign f_arrdiv24_fs464_and1 = f_arrdiv24_fs464_not1 & f_arrdiv24_fs463_or0;
  assign f_arrdiv24_fs464_or0 = f_arrdiv24_fs464_and1 | f_arrdiv24_fs464_and0;
  assign f_arrdiv24_fs465_xor0 = f_arrdiv24_mux2to1422_xor0 ^ b[9];
  assign f_arrdiv24_fs465_not0 = ~f_arrdiv24_mux2to1422_xor0;
  assign f_arrdiv24_fs465_and0 = f_arrdiv24_fs465_not0 & b[9];
  assign f_arrdiv24_fs465_xor1 = f_arrdiv24_fs464_or0 ^ f_arrdiv24_fs465_xor0;
  assign f_arrdiv24_fs465_not1 = ~f_arrdiv24_fs465_xor0;
  assign f_arrdiv24_fs465_and1 = f_arrdiv24_fs465_not1 & f_arrdiv24_fs464_or0;
  assign f_arrdiv24_fs465_or0 = f_arrdiv24_fs465_and1 | f_arrdiv24_fs465_and0;
  assign f_arrdiv24_fs466_xor0 = f_arrdiv24_mux2to1423_xor0 ^ b[10];
  assign f_arrdiv24_fs466_not0 = ~f_arrdiv24_mux2to1423_xor0;
  assign f_arrdiv24_fs466_and0 = f_arrdiv24_fs466_not0 & b[10];
  assign f_arrdiv24_fs466_xor1 = f_arrdiv24_fs465_or0 ^ f_arrdiv24_fs466_xor0;
  assign f_arrdiv24_fs466_not1 = ~f_arrdiv24_fs466_xor0;
  assign f_arrdiv24_fs466_and1 = f_arrdiv24_fs466_not1 & f_arrdiv24_fs465_or0;
  assign f_arrdiv24_fs466_or0 = f_arrdiv24_fs466_and1 | f_arrdiv24_fs466_and0;
  assign f_arrdiv24_fs467_xor0 = f_arrdiv24_mux2to1424_xor0 ^ b[11];
  assign f_arrdiv24_fs467_not0 = ~f_arrdiv24_mux2to1424_xor0;
  assign f_arrdiv24_fs467_and0 = f_arrdiv24_fs467_not0 & b[11];
  assign f_arrdiv24_fs467_xor1 = f_arrdiv24_fs466_or0 ^ f_arrdiv24_fs467_xor0;
  assign f_arrdiv24_fs467_not1 = ~f_arrdiv24_fs467_xor0;
  assign f_arrdiv24_fs467_and1 = f_arrdiv24_fs467_not1 & f_arrdiv24_fs466_or0;
  assign f_arrdiv24_fs467_or0 = f_arrdiv24_fs467_and1 | f_arrdiv24_fs467_and0;
  assign f_arrdiv24_fs468_xor0 = f_arrdiv24_mux2to1425_xor0 ^ b[12];
  assign f_arrdiv24_fs468_not0 = ~f_arrdiv24_mux2to1425_xor0;
  assign f_arrdiv24_fs468_and0 = f_arrdiv24_fs468_not0 & b[12];
  assign f_arrdiv24_fs468_xor1 = f_arrdiv24_fs467_or0 ^ f_arrdiv24_fs468_xor0;
  assign f_arrdiv24_fs468_not1 = ~f_arrdiv24_fs468_xor0;
  assign f_arrdiv24_fs468_and1 = f_arrdiv24_fs468_not1 & f_arrdiv24_fs467_or0;
  assign f_arrdiv24_fs468_or0 = f_arrdiv24_fs468_and1 | f_arrdiv24_fs468_and0;
  assign f_arrdiv24_fs469_xor0 = f_arrdiv24_mux2to1426_xor0 ^ b[13];
  assign f_arrdiv24_fs469_not0 = ~f_arrdiv24_mux2to1426_xor0;
  assign f_arrdiv24_fs469_and0 = f_arrdiv24_fs469_not0 & b[13];
  assign f_arrdiv24_fs469_xor1 = f_arrdiv24_fs468_or0 ^ f_arrdiv24_fs469_xor0;
  assign f_arrdiv24_fs469_not1 = ~f_arrdiv24_fs469_xor0;
  assign f_arrdiv24_fs469_and1 = f_arrdiv24_fs469_not1 & f_arrdiv24_fs468_or0;
  assign f_arrdiv24_fs469_or0 = f_arrdiv24_fs469_and1 | f_arrdiv24_fs469_and0;
  assign f_arrdiv24_fs470_xor0 = f_arrdiv24_mux2to1427_xor0 ^ b[14];
  assign f_arrdiv24_fs470_not0 = ~f_arrdiv24_mux2to1427_xor0;
  assign f_arrdiv24_fs470_and0 = f_arrdiv24_fs470_not0 & b[14];
  assign f_arrdiv24_fs470_xor1 = f_arrdiv24_fs469_or0 ^ f_arrdiv24_fs470_xor0;
  assign f_arrdiv24_fs470_not1 = ~f_arrdiv24_fs470_xor0;
  assign f_arrdiv24_fs470_and1 = f_arrdiv24_fs470_not1 & f_arrdiv24_fs469_or0;
  assign f_arrdiv24_fs470_or0 = f_arrdiv24_fs470_and1 | f_arrdiv24_fs470_and0;
  assign f_arrdiv24_fs471_xor0 = f_arrdiv24_mux2to1428_xor0 ^ b[15];
  assign f_arrdiv24_fs471_not0 = ~f_arrdiv24_mux2to1428_xor0;
  assign f_arrdiv24_fs471_and0 = f_arrdiv24_fs471_not0 & b[15];
  assign f_arrdiv24_fs471_xor1 = f_arrdiv24_fs470_or0 ^ f_arrdiv24_fs471_xor0;
  assign f_arrdiv24_fs471_not1 = ~f_arrdiv24_fs471_xor0;
  assign f_arrdiv24_fs471_and1 = f_arrdiv24_fs471_not1 & f_arrdiv24_fs470_or0;
  assign f_arrdiv24_fs471_or0 = f_arrdiv24_fs471_and1 | f_arrdiv24_fs471_and0;
  assign f_arrdiv24_fs472_xor0 = f_arrdiv24_mux2to1429_xor0 ^ b[16];
  assign f_arrdiv24_fs472_not0 = ~f_arrdiv24_mux2to1429_xor0;
  assign f_arrdiv24_fs472_and0 = f_arrdiv24_fs472_not0 & b[16];
  assign f_arrdiv24_fs472_xor1 = f_arrdiv24_fs471_or0 ^ f_arrdiv24_fs472_xor0;
  assign f_arrdiv24_fs472_not1 = ~f_arrdiv24_fs472_xor0;
  assign f_arrdiv24_fs472_and1 = f_arrdiv24_fs472_not1 & f_arrdiv24_fs471_or0;
  assign f_arrdiv24_fs472_or0 = f_arrdiv24_fs472_and1 | f_arrdiv24_fs472_and0;
  assign f_arrdiv24_fs473_xor0 = f_arrdiv24_mux2to1430_xor0 ^ b[17];
  assign f_arrdiv24_fs473_not0 = ~f_arrdiv24_mux2to1430_xor0;
  assign f_arrdiv24_fs473_and0 = f_arrdiv24_fs473_not0 & b[17];
  assign f_arrdiv24_fs473_xor1 = f_arrdiv24_fs472_or0 ^ f_arrdiv24_fs473_xor0;
  assign f_arrdiv24_fs473_not1 = ~f_arrdiv24_fs473_xor0;
  assign f_arrdiv24_fs473_and1 = f_arrdiv24_fs473_not1 & f_arrdiv24_fs472_or0;
  assign f_arrdiv24_fs473_or0 = f_arrdiv24_fs473_and1 | f_arrdiv24_fs473_and0;
  assign f_arrdiv24_fs474_xor0 = f_arrdiv24_mux2to1431_xor0 ^ b[18];
  assign f_arrdiv24_fs474_not0 = ~f_arrdiv24_mux2to1431_xor0;
  assign f_arrdiv24_fs474_and0 = f_arrdiv24_fs474_not0 & b[18];
  assign f_arrdiv24_fs474_xor1 = f_arrdiv24_fs473_or0 ^ f_arrdiv24_fs474_xor0;
  assign f_arrdiv24_fs474_not1 = ~f_arrdiv24_fs474_xor0;
  assign f_arrdiv24_fs474_and1 = f_arrdiv24_fs474_not1 & f_arrdiv24_fs473_or0;
  assign f_arrdiv24_fs474_or0 = f_arrdiv24_fs474_and1 | f_arrdiv24_fs474_and0;
  assign f_arrdiv24_fs475_xor0 = f_arrdiv24_mux2to1432_xor0 ^ b[19];
  assign f_arrdiv24_fs475_not0 = ~f_arrdiv24_mux2to1432_xor0;
  assign f_arrdiv24_fs475_and0 = f_arrdiv24_fs475_not0 & b[19];
  assign f_arrdiv24_fs475_xor1 = f_arrdiv24_fs474_or0 ^ f_arrdiv24_fs475_xor0;
  assign f_arrdiv24_fs475_not1 = ~f_arrdiv24_fs475_xor0;
  assign f_arrdiv24_fs475_and1 = f_arrdiv24_fs475_not1 & f_arrdiv24_fs474_or0;
  assign f_arrdiv24_fs475_or0 = f_arrdiv24_fs475_and1 | f_arrdiv24_fs475_and0;
  assign f_arrdiv24_fs476_xor0 = f_arrdiv24_mux2to1433_xor0 ^ b[20];
  assign f_arrdiv24_fs476_not0 = ~f_arrdiv24_mux2to1433_xor0;
  assign f_arrdiv24_fs476_and0 = f_arrdiv24_fs476_not0 & b[20];
  assign f_arrdiv24_fs476_xor1 = f_arrdiv24_fs475_or0 ^ f_arrdiv24_fs476_xor0;
  assign f_arrdiv24_fs476_not1 = ~f_arrdiv24_fs476_xor0;
  assign f_arrdiv24_fs476_and1 = f_arrdiv24_fs476_not1 & f_arrdiv24_fs475_or0;
  assign f_arrdiv24_fs476_or0 = f_arrdiv24_fs476_and1 | f_arrdiv24_fs476_and0;
  assign f_arrdiv24_fs477_xor0 = f_arrdiv24_mux2to1434_xor0 ^ b[21];
  assign f_arrdiv24_fs477_not0 = ~f_arrdiv24_mux2to1434_xor0;
  assign f_arrdiv24_fs477_and0 = f_arrdiv24_fs477_not0 & b[21];
  assign f_arrdiv24_fs477_xor1 = f_arrdiv24_fs476_or0 ^ f_arrdiv24_fs477_xor0;
  assign f_arrdiv24_fs477_not1 = ~f_arrdiv24_fs477_xor0;
  assign f_arrdiv24_fs477_and1 = f_arrdiv24_fs477_not1 & f_arrdiv24_fs476_or0;
  assign f_arrdiv24_fs477_or0 = f_arrdiv24_fs477_and1 | f_arrdiv24_fs477_and0;
  assign f_arrdiv24_fs478_xor0 = f_arrdiv24_mux2to1435_xor0 ^ b[22];
  assign f_arrdiv24_fs478_not0 = ~f_arrdiv24_mux2to1435_xor0;
  assign f_arrdiv24_fs478_and0 = f_arrdiv24_fs478_not0 & b[22];
  assign f_arrdiv24_fs478_xor1 = f_arrdiv24_fs477_or0 ^ f_arrdiv24_fs478_xor0;
  assign f_arrdiv24_fs478_not1 = ~f_arrdiv24_fs478_xor0;
  assign f_arrdiv24_fs478_and1 = f_arrdiv24_fs478_not1 & f_arrdiv24_fs477_or0;
  assign f_arrdiv24_fs478_or0 = f_arrdiv24_fs478_and1 | f_arrdiv24_fs478_and0;
  assign f_arrdiv24_fs479_xor0 = f_arrdiv24_mux2to1436_xor0 ^ b[23];
  assign f_arrdiv24_fs479_not0 = ~f_arrdiv24_mux2to1436_xor0;
  assign f_arrdiv24_fs479_and0 = f_arrdiv24_fs479_not0 & b[23];
  assign f_arrdiv24_fs479_xor1 = f_arrdiv24_fs478_or0 ^ f_arrdiv24_fs479_xor0;
  assign f_arrdiv24_fs479_not1 = ~f_arrdiv24_fs479_xor0;
  assign f_arrdiv24_fs479_and1 = f_arrdiv24_fs479_not1 & f_arrdiv24_fs478_or0;
  assign f_arrdiv24_fs479_or0 = f_arrdiv24_fs479_and1 | f_arrdiv24_fs479_and0;
  assign f_arrdiv24_mux2to1437_and0 = a[4] & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1437_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1437_and1 = f_arrdiv24_fs456_xor0 & f_arrdiv24_mux2to1437_not0;
  assign f_arrdiv24_mux2to1437_xor0 = f_arrdiv24_mux2to1437_and0 ^ f_arrdiv24_mux2to1437_and1;
  assign f_arrdiv24_mux2to1438_and0 = f_arrdiv24_mux2to1414_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1438_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1438_and1 = f_arrdiv24_fs457_xor1 & f_arrdiv24_mux2to1438_not0;
  assign f_arrdiv24_mux2to1438_xor0 = f_arrdiv24_mux2to1438_and0 ^ f_arrdiv24_mux2to1438_and1;
  assign f_arrdiv24_mux2to1439_and0 = f_arrdiv24_mux2to1415_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1439_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1439_and1 = f_arrdiv24_fs458_xor1 & f_arrdiv24_mux2to1439_not0;
  assign f_arrdiv24_mux2to1439_xor0 = f_arrdiv24_mux2to1439_and0 ^ f_arrdiv24_mux2to1439_and1;
  assign f_arrdiv24_mux2to1440_and0 = f_arrdiv24_mux2to1416_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1440_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1440_and1 = f_arrdiv24_fs459_xor1 & f_arrdiv24_mux2to1440_not0;
  assign f_arrdiv24_mux2to1440_xor0 = f_arrdiv24_mux2to1440_and0 ^ f_arrdiv24_mux2to1440_and1;
  assign f_arrdiv24_mux2to1441_and0 = f_arrdiv24_mux2to1417_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1441_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1441_and1 = f_arrdiv24_fs460_xor1 & f_arrdiv24_mux2to1441_not0;
  assign f_arrdiv24_mux2to1441_xor0 = f_arrdiv24_mux2to1441_and0 ^ f_arrdiv24_mux2to1441_and1;
  assign f_arrdiv24_mux2to1442_and0 = f_arrdiv24_mux2to1418_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1442_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1442_and1 = f_arrdiv24_fs461_xor1 & f_arrdiv24_mux2to1442_not0;
  assign f_arrdiv24_mux2to1442_xor0 = f_arrdiv24_mux2to1442_and0 ^ f_arrdiv24_mux2to1442_and1;
  assign f_arrdiv24_mux2to1443_and0 = f_arrdiv24_mux2to1419_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1443_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1443_and1 = f_arrdiv24_fs462_xor1 & f_arrdiv24_mux2to1443_not0;
  assign f_arrdiv24_mux2to1443_xor0 = f_arrdiv24_mux2to1443_and0 ^ f_arrdiv24_mux2to1443_and1;
  assign f_arrdiv24_mux2to1444_and0 = f_arrdiv24_mux2to1420_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1444_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1444_and1 = f_arrdiv24_fs463_xor1 & f_arrdiv24_mux2to1444_not0;
  assign f_arrdiv24_mux2to1444_xor0 = f_arrdiv24_mux2to1444_and0 ^ f_arrdiv24_mux2to1444_and1;
  assign f_arrdiv24_mux2to1445_and0 = f_arrdiv24_mux2to1421_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1445_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1445_and1 = f_arrdiv24_fs464_xor1 & f_arrdiv24_mux2to1445_not0;
  assign f_arrdiv24_mux2to1445_xor0 = f_arrdiv24_mux2to1445_and0 ^ f_arrdiv24_mux2to1445_and1;
  assign f_arrdiv24_mux2to1446_and0 = f_arrdiv24_mux2to1422_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1446_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1446_and1 = f_arrdiv24_fs465_xor1 & f_arrdiv24_mux2to1446_not0;
  assign f_arrdiv24_mux2to1446_xor0 = f_arrdiv24_mux2to1446_and0 ^ f_arrdiv24_mux2to1446_and1;
  assign f_arrdiv24_mux2to1447_and0 = f_arrdiv24_mux2to1423_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1447_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1447_and1 = f_arrdiv24_fs466_xor1 & f_arrdiv24_mux2to1447_not0;
  assign f_arrdiv24_mux2to1447_xor0 = f_arrdiv24_mux2to1447_and0 ^ f_arrdiv24_mux2to1447_and1;
  assign f_arrdiv24_mux2to1448_and0 = f_arrdiv24_mux2to1424_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1448_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1448_and1 = f_arrdiv24_fs467_xor1 & f_arrdiv24_mux2to1448_not0;
  assign f_arrdiv24_mux2to1448_xor0 = f_arrdiv24_mux2to1448_and0 ^ f_arrdiv24_mux2to1448_and1;
  assign f_arrdiv24_mux2to1449_and0 = f_arrdiv24_mux2to1425_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1449_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1449_and1 = f_arrdiv24_fs468_xor1 & f_arrdiv24_mux2to1449_not0;
  assign f_arrdiv24_mux2to1449_xor0 = f_arrdiv24_mux2to1449_and0 ^ f_arrdiv24_mux2to1449_and1;
  assign f_arrdiv24_mux2to1450_and0 = f_arrdiv24_mux2to1426_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1450_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1450_and1 = f_arrdiv24_fs469_xor1 & f_arrdiv24_mux2to1450_not0;
  assign f_arrdiv24_mux2to1450_xor0 = f_arrdiv24_mux2to1450_and0 ^ f_arrdiv24_mux2to1450_and1;
  assign f_arrdiv24_mux2to1451_and0 = f_arrdiv24_mux2to1427_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1451_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1451_and1 = f_arrdiv24_fs470_xor1 & f_arrdiv24_mux2to1451_not0;
  assign f_arrdiv24_mux2to1451_xor0 = f_arrdiv24_mux2to1451_and0 ^ f_arrdiv24_mux2to1451_and1;
  assign f_arrdiv24_mux2to1452_and0 = f_arrdiv24_mux2to1428_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1452_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1452_and1 = f_arrdiv24_fs471_xor1 & f_arrdiv24_mux2to1452_not0;
  assign f_arrdiv24_mux2to1452_xor0 = f_arrdiv24_mux2to1452_and0 ^ f_arrdiv24_mux2to1452_and1;
  assign f_arrdiv24_mux2to1453_and0 = f_arrdiv24_mux2to1429_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1453_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1453_and1 = f_arrdiv24_fs472_xor1 & f_arrdiv24_mux2to1453_not0;
  assign f_arrdiv24_mux2to1453_xor0 = f_arrdiv24_mux2to1453_and0 ^ f_arrdiv24_mux2to1453_and1;
  assign f_arrdiv24_mux2to1454_and0 = f_arrdiv24_mux2to1430_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1454_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1454_and1 = f_arrdiv24_fs473_xor1 & f_arrdiv24_mux2to1454_not0;
  assign f_arrdiv24_mux2to1454_xor0 = f_arrdiv24_mux2to1454_and0 ^ f_arrdiv24_mux2to1454_and1;
  assign f_arrdiv24_mux2to1455_and0 = f_arrdiv24_mux2to1431_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1455_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1455_and1 = f_arrdiv24_fs474_xor1 & f_arrdiv24_mux2to1455_not0;
  assign f_arrdiv24_mux2to1455_xor0 = f_arrdiv24_mux2to1455_and0 ^ f_arrdiv24_mux2to1455_and1;
  assign f_arrdiv24_mux2to1456_and0 = f_arrdiv24_mux2to1432_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1456_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1456_and1 = f_arrdiv24_fs475_xor1 & f_arrdiv24_mux2to1456_not0;
  assign f_arrdiv24_mux2to1456_xor0 = f_arrdiv24_mux2to1456_and0 ^ f_arrdiv24_mux2to1456_and1;
  assign f_arrdiv24_mux2to1457_and0 = f_arrdiv24_mux2to1433_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1457_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1457_and1 = f_arrdiv24_fs476_xor1 & f_arrdiv24_mux2to1457_not0;
  assign f_arrdiv24_mux2to1457_xor0 = f_arrdiv24_mux2to1457_and0 ^ f_arrdiv24_mux2to1457_and1;
  assign f_arrdiv24_mux2to1458_and0 = f_arrdiv24_mux2to1434_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1458_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1458_and1 = f_arrdiv24_fs477_xor1 & f_arrdiv24_mux2to1458_not0;
  assign f_arrdiv24_mux2to1458_xor0 = f_arrdiv24_mux2to1458_and0 ^ f_arrdiv24_mux2to1458_and1;
  assign f_arrdiv24_mux2to1459_and0 = f_arrdiv24_mux2to1435_xor0 & f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1459_not0 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_mux2to1459_and1 = f_arrdiv24_fs478_xor1 & f_arrdiv24_mux2to1459_not0;
  assign f_arrdiv24_mux2to1459_xor0 = f_arrdiv24_mux2to1459_and0 ^ f_arrdiv24_mux2to1459_and1;
  assign f_arrdiv24_not19 = ~f_arrdiv24_fs479_or0;
  assign f_arrdiv24_fs480_xor0 = a[3] ^ b[0];
  assign f_arrdiv24_fs480_not0 = ~a[3];
  assign f_arrdiv24_fs480_and0 = f_arrdiv24_fs480_not0 & b[0];
  assign f_arrdiv24_fs480_not1 = ~f_arrdiv24_fs480_xor0;
  assign f_arrdiv24_fs481_xor0 = f_arrdiv24_mux2to1437_xor0 ^ b[1];
  assign f_arrdiv24_fs481_not0 = ~f_arrdiv24_mux2to1437_xor0;
  assign f_arrdiv24_fs481_and0 = f_arrdiv24_fs481_not0 & b[1];
  assign f_arrdiv24_fs481_xor1 = f_arrdiv24_fs480_and0 ^ f_arrdiv24_fs481_xor0;
  assign f_arrdiv24_fs481_not1 = ~f_arrdiv24_fs481_xor0;
  assign f_arrdiv24_fs481_and1 = f_arrdiv24_fs481_not1 & f_arrdiv24_fs480_and0;
  assign f_arrdiv24_fs481_or0 = f_arrdiv24_fs481_and1 | f_arrdiv24_fs481_and0;
  assign f_arrdiv24_fs482_xor0 = f_arrdiv24_mux2to1438_xor0 ^ b[2];
  assign f_arrdiv24_fs482_not0 = ~f_arrdiv24_mux2to1438_xor0;
  assign f_arrdiv24_fs482_and0 = f_arrdiv24_fs482_not0 & b[2];
  assign f_arrdiv24_fs482_xor1 = f_arrdiv24_fs481_or0 ^ f_arrdiv24_fs482_xor0;
  assign f_arrdiv24_fs482_not1 = ~f_arrdiv24_fs482_xor0;
  assign f_arrdiv24_fs482_and1 = f_arrdiv24_fs482_not1 & f_arrdiv24_fs481_or0;
  assign f_arrdiv24_fs482_or0 = f_arrdiv24_fs482_and1 | f_arrdiv24_fs482_and0;
  assign f_arrdiv24_fs483_xor0 = f_arrdiv24_mux2to1439_xor0 ^ b[3];
  assign f_arrdiv24_fs483_not0 = ~f_arrdiv24_mux2to1439_xor0;
  assign f_arrdiv24_fs483_and0 = f_arrdiv24_fs483_not0 & b[3];
  assign f_arrdiv24_fs483_xor1 = f_arrdiv24_fs482_or0 ^ f_arrdiv24_fs483_xor0;
  assign f_arrdiv24_fs483_not1 = ~f_arrdiv24_fs483_xor0;
  assign f_arrdiv24_fs483_and1 = f_arrdiv24_fs483_not1 & f_arrdiv24_fs482_or0;
  assign f_arrdiv24_fs483_or0 = f_arrdiv24_fs483_and1 | f_arrdiv24_fs483_and0;
  assign f_arrdiv24_fs484_xor0 = f_arrdiv24_mux2to1440_xor0 ^ b[4];
  assign f_arrdiv24_fs484_not0 = ~f_arrdiv24_mux2to1440_xor0;
  assign f_arrdiv24_fs484_and0 = f_arrdiv24_fs484_not0 & b[4];
  assign f_arrdiv24_fs484_xor1 = f_arrdiv24_fs483_or0 ^ f_arrdiv24_fs484_xor0;
  assign f_arrdiv24_fs484_not1 = ~f_arrdiv24_fs484_xor0;
  assign f_arrdiv24_fs484_and1 = f_arrdiv24_fs484_not1 & f_arrdiv24_fs483_or0;
  assign f_arrdiv24_fs484_or0 = f_arrdiv24_fs484_and1 | f_arrdiv24_fs484_and0;
  assign f_arrdiv24_fs485_xor0 = f_arrdiv24_mux2to1441_xor0 ^ b[5];
  assign f_arrdiv24_fs485_not0 = ~f_arrdiv24_mux2to1441_xor0;
  assign f_arrdiv24_fs485_and0 = f_arrdiv24_fs485_not0 & b[5];
  assign f_arrdiv24_fs485_xor1 = f_arrdiv24_fs484_or0 ^ f_arrdiv24_fs485_xor0;
  assign f_arrdiv24_fs485_not1 = ~f_arrdiv24_fs485_xor0;
  assign f_arrdiv24_fs485_and1 = f_arrdiv24_fs485_not1 & f_arrdiv24_fs484_or0;
  assign f_arrdiv24_fs485_or0 = f_arrdiv24_fs485_and1 | f_arrdiv24_fs485_and0;
  assign f_arrdiv24_fs486_xor0 = f_arrdiv24_mux2to1442_xor0 ^ b[6];
  assign f_arrdiv24_fs486_not0 = ~f_arrdiv24_mux2to1442_xor0;
  assign f_arrdiv24_fs486_and0 = f_arrdiv24_fs486_not0 & b[6];
  assign f_arrdiv24_fs486_xor1 = f_arrdiv24_fs485_or0 ^ f_arrdiv24_fs486_xor0;
  assign f_arrdiv24_fs486_not1 = ~f_arrdiv24_fs486_xor0;
  assign f_arrdiv24_fs486_and1 = f_arrdiv24_fs486_not1 & f_arrdiv24_fs485_or0;
  assign f_arrdiv24_fs486_or0 = f_arrdiv24_fs486_and1 | f_arrdiv24_fs486_and0;
  assign f_arrdiv24_fs487_xor0 = f_arrdiv24_mux2to1443_xor0 ^ b[7];
  assign f_arrdiv24_fs487_not0 = ~f_arrdiv24_mux2to1443_xor0;
  assign f_arrdiv24_fs487_and0 = f_arrdiv24_fs487_not0 & b[7];
  assign f_arrdiv24_fs487_xor1 = f_arrdiv24_fs486_or0 ^ f_arrdiv24_fs487_xor0;
  assign f_arrdiv24_fs487_not1 = ~f_arrdiv24_fs487_xor0;
  assign f_arrdiv24_fs487_and1 = f_arrdiv24_fs487_not1 & f_arrdiv24_fs486_or0;
  assign f_arrdiv24_fs487_or0 = f_arrdiv24_fs487_and1 | f_arrdiv24_fs487_and0;
  assign f_arrdiv24_fs488_xor0 = f_arrdiv24_mux2to1444_xor0 ^ b[8];
  assign f_arrdiv24_fs488_not0 = ~f_arrdiv24_mux2to1444_xor0;
  assign f_arrdiv24_fs488_and0 = f_arrdiv24_fs488_not0 & b[8];
  assign f_arrdiv24_fs488_xor1 = f_arrdiv24_fs487_or0 ^ f_arrdiv24_fs488_xor0;
  assign f_arrdiv24_fs488_not1 = ~f_arrdiv24_fs488_xor0;
  assign f_arrdiv24_fs488_and1 = f_arrdiv24_fs488_not1 & f_arrdiv24_fs487_or0;
  assign f_arrdiv24_fs488_or0 = f_arrdiv24_fs488_and1 | f_arrdiv24_fs488_and0;
  assign f_arrdiv24_fs489_xor0 = f_arrdiv24_mux2to1445_xor0 ^ b[9];
  assign f_arrdiv24_fs489_not0 = ~f_arrdiv24_mux2to1445_xor0;
  assign f_arrdiv24_fs489_and0 = f_arrdiv24_fs489_not0 & b[9];
  assign f_arrdiv24_fs489_xor1 = f_arrdiv24_fs488_or0 ^ f_arrdiv24_fs489_xor0;
  assign f_arrdiv24_fs489_not1 = ~f_arrdiv24_fs489_xor0;
  assign f_arrdiv24_fs489_and1 = f_arrdiv24_fs489_not1 & f_arrdiv24_fs488_or0;
  assign f_arrdiv24_fs489_or0 = f_arrdiv24_fs489_and1 | f_arrdiv24_fs489_and0;
  assign f_arrdiv24_fs490_xor0 = f_arrdiv24_mux2to1446_xor0 ^ b[10];
  assign f_arrdiv24_fs490_not0 = ~f_arrdiv24_mux2to1446_xor0;
  assign f_arrdiv24_fs490_and0 = f_arrdiv24_fs490_not0 & b[10];
  assign f_arrdiv24_fs490_xor1 = f_arrdiv24_fs489_or0 ^ f_arrdiv24_fs490_xor0;
  assign f_arrdiv24_fs490_not1 = ~f_arrdiv24_fs490_xor0;
  assign f_arrdiv24_fs490_and1 = f_arrdiv24_fs490_not1 & f_arrdiv24_fs489_or0;
  assign f_arrdiv24_fs490_or0 = f_arrdiv24_fs490_and1 | f_arrdiv24_fs490_and0;
  assign f_arrdiv24_fs491_xor0 = f_arrdiv24_mux2to1447_xor0 ^ b[11];
  assign f_arrdiv24_fs491_not0 = ~f_arrdiv24_mux2to1447_xor0;
  assign f_arrdiv24_fs491_and0 = f_arrdiv24_fs491_not0 & b[11];
  assign f_arrdiv24_fs491_xor1 = f_arrdiv24_fs490_or0 ^ f_arrdiv24_fs491_xor0;
  assign f_arrdiv24_fs491_not1 = ~f_arrdiv24_fs491_xor0;
  assign f_arrdiv24_fs491_and1 = f_arrdiv24_fs491_not1 & f_arrdiv24_fs490_or0;
  assign f_arrdiv24_fs491_or0 = f_arrdiv24_fs491_and1 | f_arrdiv24_fs491_and0;
  assign f_arrdiv24_fs492_xor0 = f_arrdiv24_mux2to1448_xor0 ^ b[12];
  assign f_arrdiv24_fs492_not0 = ~f_arrdiv24_mux2to1448_xor0;
  assign f_arrdiv24_fs492_and0 = f_arrdiv24_fs492_not0 & b[12];
  assign f_arrdiv24_fs492_xor1 = f_arrdiv24_fs491_or0 ^ f_arrdiv24_fs492_xor0;
  assign f_arrdiv24_fs492_not1 = ~f_arrdiv24_fs492_xor0;
  assign f_arrdiv24_fs492_and1 = f_arrdiv24_fs492_not1 & f_arrdiv24_fs491_or0;
  assign f_arrdiv24_fs492_or0 = f_arrdiv24_fs492_and1 | f_arrdiv24_fs492_and0;
  assign f_arrdiv24_fs493_xor0 = f_arrdiv24_mux2to1449_xor0 ^ b[13];
  assign f_arrdiv24_fs493_not0 = ~f_arrdiv24_mux2to1449_xor0;
  assign f_arrdiv24_fs493_and0 = f_arrdiv24_fs493_not0 & b[13];
  assign f_arrdiv24_fs493_xor1 = f_arrdiv24_fs492_or0 ^ f_arrdiv24_fs493_xor0;
  assign f_arrdiv24_fs493_not1 = ~f_arrdiv24_fs493_xor0;
  assign f_arrdiv24_fs493_and1 = f_arrdiv24_fs493_not1 & f_arrdiv24_fs492_or0;
  assign f_arrdiv24_fs493_or0 = f_arrdiv24_fs493_and1 | f_arrdiv24_fs493_and0;
  assign f_arrdiv24_fs494_xor0 = f_arrdiv24_mux2to1450_xor0 ^ b[14];
  assign f_arrdiv24_fs494_not0 = ~f_arrdiv24_mux2to1450_xor0;
  assign f_arrdiv24_fs494_and0 = f_arrdiv24_fs494_not0 & b[14];
  assign f_arrdiv24_fs494_xor1 = f_arrdiv24_fs493_or0 ^ f_arrdiv24_fs494_xor0;
  assign f_arrdiv24_fs494_not1 = ~f_arrdiv24_fs494_xor0;
  assign f_arrdiv24_fs494_and1 = f_arrdiv24_fs494_not1 & f_arrdiv24_fs493_or0;
  assign f_arrdiv24_fs494_or0 = f_arrdiv24_fs494_and1 | f_arrdiv24_fs494_and0;
  assign f_arrdiv24_fs495_xor0 = f_arrdiv24_mux2to1451_xor0 ^ b[15];
  assign f_arrdiv24_fs495_not0 = ~f_arrdiv24_mux2to1451_xor0;
  assign f_arrdiv24_fs495_and0 = f_arrdiv24_fs495_not0 & b[15];
  assign f_arrdiv24_fs495_xor1 = f_arrdiv24_fs494_or0 ^ f_arrdiv24_fs495_xor0;
  assign f_arrdiv24_fs495_not1 = ~f_arrdiv24_fs495_xor0;
  assign f_arrdiv24_fs495_and1 = f_arrdiv24_fs495_not1 & f_arrdiv24_fs494_or0;
  assign f_arrdiv24_fs495_or0 = f_arrdiv24_fs495_and1 | f_arrdiv24_fs495_and0;
  assign f_arrdiv24_fs496_xor0 = f_arrdiv24_mux2to1452_xor0 ^ b[16];
  assign f_arrdiv24_fs496_not0 = ~f_arrdiv24_mux2to1452_xor0;
  assign f_arrdiv24_fs496_and0 = f_arrdiv24_fs496_not0 & b[16];
  assign f_arrdiv24_fs496_xor1 = f_arrdiv24_fs495_or0 ^ f_arrdiv24_fs496_xor0;
  assign f_arrdiv24_fs496_not1 = ~f_arrdiv24_fs496_xor0;
  assign f_arrdiv24_fs496_and1 = f_arrdiv24_fs496_not1 & f_arrdiv24_fs495_or0;
  assign f_arrdiv24_fs496_or0 = f_arrdiv24_fs496_and1 | f_arrdiv24_fs496_and0;
  assign f_arrdiv24_fs497_xor0 = f_arrdiv24_mux2to1453_xor0 ^ b[17];
  assign f_arrdiv24_fs497_not0 = ~f_arrdiv24_mux2to1453_xor0;
  assign f_arrdiv24_fs497_and0 = f_arrdiv24_fs497_not0 & b[17];
  assign f_arrdiv24_fs497_xor1 = f_arrdiv24_fs496_or0 ^ f_arrdiv24_fs497_xor0;
  assign f_arrdiv24_fs497_not1 = ~f_arrdiv24_fs497_xor0;
  assign f_arrdiv24_fs497_and1 = f_arrdiv24_fs497_not1 & f_arrdiv24_fs496_or0;
  assign f_arrdiv24_fs497_or0 = f_arrdiv24_fs497_and1 | f_arrdiv24_fs497_and0;
  assign f_arrdiv24_fs498_xor0 = f_arrdiv24_mux2to1454_xor0 ^ b[18];
  assign f_arrdiv24_fs498_not0 = ~f_arrdiv24_mux2to1454_xor0;
  assign f_arrdiv24_fs498_and0 = f_arrdiv24_fs498_not0 & b[18];
  assign f_arrdiv24_fs498_xor1 = f_arrdiv24_fs497_or0 ^ f_arrdiv24_fs498_xor0;
  assign f_arrdiv24_fs498_not1 = ~f_arrdiv24_fs498_xor0;
  assign f_arrdiv24_fs498_and1 = f_arrdiv24_fs498_not1 & f_arrdiv24_fs497_or0;
  assign f_arrdiv24_fs498_or0 = f_arrdiv24_fs498_and1 | f_arrdiv24_fs498_and0;
  assign f_arrdiv24_fs499_xor0 = f_arrdiv24_mux2to1455_xor0 ^ b[19];
  assign f_arrdiv24_fs499_not0 = ~f_arrdiv24_mux2to1455_xor0;
  assign f_arrdiv24_fs499_and0 = f_arrdiv24_fs499_not0 & b[19];
  assign f_arrdiv24_fs499_xor1 = f_arrdiv24_fs498_or0 ^ f_arrdiv24_fs499_xor0;
  assign f_arrdiv24_fs499_not1 = ~f_arrdiv24_fs499_xor0;
  assign f_arrdiv24_fs499_and1 = f_arrdiv24_fs499_not1 & f_arrdiv24_fs498_or0;
  assign f_arrdiv24_fs499_or0 = f_arrdiv24_fs499_and1 | f_arrdiv24_fs499_and0;
  assign f_arrdiv24_fs500_xor0 = f_arrdiv24_mux2to1456_xor0 ^ b[20];
  assign f_arrdiv24_fs500_not0 = ~f_arrdiv24_mux2to1456_xor0;
  assign f_arrdiv24_fs500_and0 = f_arrdiv24_fs500_not0 & b[20];
  assign f_arrdiv24_fs500_xor1 = f_arrdiv24_fs499_or0 ^ f_arrdiv24_fs500_xor0;
  assign f_arrdiv24_fs500_not1 = ~f_arrdiv24_fs500_xor0;
  assign f_arrdiv24_fs500_and1 = f_arrdiv24_fs500_not1 & f_arrdiv24_fs499_or0;
  assign f_arrdiv24_fs500_or0 = f_arrdiv24_fs500_and1 | f_arrdiv24_fs500_and0;
  assign f_arrdiv24_fs501_xor0 = f_arrdiv24_mux2to1457_xor0 ^ b[21];
  assign f_arrdiv24_fs501_not0 = ~f_arrdiv24_mux2to1457_xor0;
  assign f_arrdiv24_fs501_and0 = f_arrdiv24_fs501_not0 & b[21];
  assign f_arrdiv24_fs501_xor1 = f_arrdiv24_fs500_or0 ^ f_arrdiv24_fs501_xor0;
  assign f_arrdiv24_fs501_not1 = ~f_arrdiv24_fs501_xor0;
  assign f_arrdiv24_fs501_and1 = f_arrdiv24_fs501_not1 & f_arrdiv24_fs500_or0;
  assign f_arrdiv24_fs501_or0 = f_arrdiv24_fs501_and1 | f_arrdiv24_fs501_and0;
  assign f_arrdiv24_fs502_xor0 = f_arrdiv24_mux2to1458_xor0 ^ b[22];
  assign f_arrdiv24_fs502_not0 = ~f_arrdiv24_mux2to1458_xor0;
  assign f_arrdiv24_fs502_and0 = f_arrdiv24_fs502_not0 & b[22];
  assign f_arrdiv24_fs502_xor1 = f_arrdiv24_fs501_or0 ^ f_arrdiv24_fs502_xor0;
  assign f_arrdiv24_fs502_not1 = ~f_arrdiv24_fs502_xor0;
  assign f_arrdiv24_fs502_and1 = f_arrdiv24_fs502_not1 & f_arrdiv24_fs501_or0;
  assign f_arrdiv24_fs502_or0 = f_arrdiv24_fs502_and1 | f_arrdiv24_fs502_and0;
  assign f_arrdiv24_fs503_xor0 = f_arrdiv24_mux2to1459_xor0 ^ b[23];
  assign f_arrdiv24_fs503_not0 = ~f_arrdiv24_mux2to1459_xor0;
  assign f_arrdiv24_fs503_and0 = f_arrdiv24_fs503_not0 & b[23];
  assign f_arrdiv24_fs503_xor1 = f_arrdiv24_fs502_or0 ^ f_arrdiv24_fs503_xor0;
  assign f_arrdiv24_fs503_not1 = ~f_arrdiv24_fs503_xor0;
  assign f_arrdiv24_fs503_and1 = f_arrdiv24_fs503_not1 & f_arrdiv24_fs502_or0;
  assign f_arrdiv24_fs503_or0 = f_arrdiv24_fs503_and1 | f_arrdiv24_fs503_and0;
  assign f_arrdiv24_mux2to1460_and0 = a[3] & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1460_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1460_and1 = f_arrdiv24_fs480_xor0 & f_arrdiv24_mux2to1460_not0;
  assign f_arrdiv24_mux2to1460_xor0 = f_arrdiv24_mux2to1460_and0 ^ f_arrdiv24_mux2to1460_and1;
  assign f_arrdiv24_mux2to1461_and0 = f_arrdiv24_mux2to1437_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1461_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1461_and1 = f_arrdiv24_fs481_xor1 & f_arrdiv24_mux2to1461_not0;
  assign f_arrdiv24_mux2to1461_xor0 = f_arrdiv24_mux2to1461_and0 ^ f_arrdiv24_mux2to1461_and1;
  assign f_arrdiv24_mux2to1462_and0 = f_arrdiv24_mux2to1438_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1462_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1462_and1 = f_arrdiv24_fs482_xor1 & f_arrdiv24_mux2to1462_not0;
  assign f_arrdiv24_mux2to1462_xor0 = f_arrdiv24_mux2to1462_and0 ^ f_arrdiv24_mux2to1462_and1;
  assign f_arrdiv24_mux2to1463_and0 = f_arrdiv24_mux2to1439_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1463_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1463_and1 = f_arrdiv24_fs483_xor1 & f_arrdiv24_mux2to1463_not0;
  assign f_arrdiv24_mux2to1463_xor0 = f_arrdiv24_mux2to1463_and0 ^ f_arrdiv24_mux2to1463_and1;
  assign f_arrdiv24_mux2to1464_and0 = f_arrdiv24_mux2to1440_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1464_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1464_and1 = f_arrdiv24_fs484_xor1 & f_arrdiv24_mux2to1464_not0;
  assign f_arrdiv24_mux2to1464_xor0 = f_arrdiv24_mux2to1464_and0 ^ f_arrdiv24_mux2to1464_and1;
  assign f_arrdiv24_mux2to1465_and0 = f_arrdiv24_mux2to1441_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1465_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1465_and1 = f_arrdiv24_fs485_xor1 & f_arrdiv24_mux2to1465_not0;
  assign f_arrdiv24_mux2to1465_xor0 = f_arrdiv24_mux2to1465_and0 ^ f_arrdiv24_mux2to1465_and1;
  assign f_arrdiv24_mux2to1466_and0 = f_arrdiv24_mux2to1442_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1466_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1466_and1 = f_arrdiv24_fs486_xor1 & f_arrdiv24_mux2to1466_not0;
  assign f_arrdiv24_mux2to1466_xor0 = f_arrdiv24_mux2to1466_and0 ^ f_arrdiv24_mux2to1466_and1;
  assign f_arrdiv24_mux2to1467_and0 = f_arrdiv24_mux2to1443_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1467_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1467_and1 = f_arrdiv24_fs487_xor1 & f_arrdiv24_mux2to1467_not0;
  assign f_arrdiv24_mux2to1467_xor0 = f_arrdiv24_mux2to1467_and0 ^ f_arrdiv24_mux2to1467_and1;
  assign f_arrdiv24_mux2to1468_and0 = f_arrdiv24_mux2to1444_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1468_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1468_and1 = f_arrdiv24_fs488_xor1 & f_arrdiv24_mux2to1468_not0;
  assign f_arrdiv24_mux2to1468_xor0 = f_arrdiv24_mux2to1468_and0 ^ f_arrdiv24_mux2to1468_and1;
  assign f_arrdiv24_mux2to1469_and0 = f_arrdiv24_mux2to1445_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1469_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1469_and1 = f_arrdiv24_fs489_xor1 & f_arrdiv24_mux2to1469_not0;
  assign f_arrdiv24_mux2to1469_xor0 = f_arrdiv24_mux2to1469_and0 ^ f_arrdiv24_mux2to1469_and1;
  assign f_arrdiv24_mux2to1470_and0 = f_arrdiv24_mux2to1446_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1470_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1470_and1 = f_arrdiv24_fs490_xor1 & f_arrdiv24_mux2to1470_not0;
  assign f_arrdiv24_mux2to1470_xor0 = f_arrdiv24_mux2to1470_and0 ^ f_arrdiv24_mux2to1470_and1;
  assign f_arrdiv24_mux2to1471_and0 = f_arrdiv24_mux2to1447_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1471_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1471_and1 = f_arrdiv24_fs491_xor1 & f_arrdiv24_mux2to1471_not0;
  assign f_arrdiv24_mux2to1471_xor0 = f_arrdiv24_mux2to1471_and0 ^ f_arrdiv24_mux2to1471_and1;
  assign f_arrdiv24_mux2to1472_and0 = f_arrdiv24_mux2to1448_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1472_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1472_and1 = f_arrdiv24_fs492_xor1 & f_arrdiv24_mux2to1472_not0;
  assign f_arrdiv24_mux2to1472_xor0 = f_arrdiv24_mux2to1472_and0 ^ f_arrdiv24_mux2to1472_and1;
  assign f_arrdiv24_mux2to1473_and0 = f_arrdiv24_mux2to1449_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1473_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1473_and1 = f_arrdiv24_fs493_xor1 & f_arrdiv24_mux2to1473_not0;
  assign f_arrdiv24_mux2to1473_xor0 = f_arrdiv24_mux2to1473_and0 ^ f_arrdiv24_mux2to1473_and1;
  assign f_arrdiv24_mux2to1474_and0 = f_arrdiv24_mux2to1450_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1474_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1474_and1 = f_arrdiv24_fs494_xor1 & f_arrdiv24_mux2to1474_not0;
  assign f_arrdiv24_mux2to1474_xor0 = f_arrdiv24_mux2to1474_and0 ^ f_arrdiv24_mux2to1474_and1;
  assign f_arrdiv24_mux2to1475_and0 = f_arrdiv24_mux2to1451_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1475_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1475_and1 = f_arrdiv24_fs495_xor1 & f_arrdiv24_mux2to1475_not0;
  assign f_arrdiv24_mux2to1475_xor0 = f_arrdiv24_mux2to1475_and0 ^ f_arrdiv24_mux2to1475_and1;
  assign f_arrdiv24_mux2to1476_and0 = f_arrdiv24_mux2to1452_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1476_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1476_and1 = f_arrdiv24_fs496_xor1 & f_arrdiv24_mux2to1476_not0;
  assign f_arrdiv24_mux2to1476_xor0 = f_arrdiv24_mux2to1476_and0 ^ f_arrdiv24_mux2to1476_and1;
  assign f_arrdiv24_mux2to1477_and0 = f_arrdiv24_mux2to1453_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1477_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1477_and1 = f_arrdiv24_fs497_xor1 & f_arrdiv24_mux2to1477_not0;
  assign f_arrdiv24_mux2to1477_xor0 = f_arrdiv24_mux2to1477_and0 ^ f_arrdiv24_mux2to1477_and1;
  assign f_arrdiv24_mux2to1478_and0 = f_arrdiv24_mux2to1454_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1478_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1478_and1 = f_arrdiv24_fs498_xor1 & f_arrdiv24_mux2to1478_not0;
  assign f_arrdiv24_mux2to1478_xor0 = f_arrdiv24_mux2to1478_and0 ^ f_arrdiv24_mux2to1478_and1;
  assign f_arrdiv24_mux2to1479_and0 = f_arrdiv24_mux2to1455_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1479_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1479_and1 = f_arrdiv24_fs499_xor1 & f_arrdiv24_mux2to1479_not0;
  assign f_arrdiv24_mux2to1479_xor0 = f_arrdiv24_mux2to1479_and0 ^ f_arrdiv24_mux2to1479_and1;
  assign f_arrdiv24_mux2to1480_and0 = f_arrdiv24_mux2to1456_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1480_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1480_and1 = f_arrdiv24_fs500_xor1 & f_arrdiv24_mux2to1480_not0;
  assign f_arrdiv24_mux2to1480_xor0 = f_arrdiv24_mux2to1480_and0 ^ f_arrdiv24_mux2to1480_and1;
  assign f_arrdiv24_mux2to1481_and0 = f_arrdiv24_mux2to1457_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1481_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1481_and1 = f_arrdiv24_fs501_xor1 & f_arrdiv24_mux2to1481_not0;
  assign f_arrdiv24_mux2to1481_xor0 = f_arrdiv24_mux2to1481_and0 ^ f_arrdiv24_mux2to1481_and1;
  assign f_arrdiv24_mux2to1482_and0 = f_arrdiv24_mux2to1458_xor0 & f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1482_not0 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_mux2to1482_and1 = f_arrdiv24_fs502_xor1 & f_arrdiv24_mux2to1482_not0;
  assign f_arrdiv24_mux2to1482_xor0 = f_arrdiv24_mux2to1482_and0 ^ f_arrdiv24_mux2to1482_and1;
  assign f_arrdiv24_not20 = ~f_arrdiv24_fs503_or0;
  assign f_arrdiv24_fs504_xor0 = a[2] ^ b[0];
  assign f_arrdiv24_fs504_not0 = ~a[2];
  assign f_arrdiv24_fs504_and0 = f_arrdiv24_fs504_not0 & b[0];
  assign f_arrdiv24_fs504_not1 = ~f_arrdiv24_fs504_xor0;
  assign f_arrdiv24_fs505_xor0 = f_arrdiv24_mux2to1460_xor0 ^ b[1];
  assign f_arrdiv24_fs505_not0 = ~f_arrdiv24_mux2to1460_xor0;
  assign f_arrdiv24_fs505_and0 = f_arrdiv24_fs505_not0 & b[1];
  assign f_arrdiv24_fs505_xor1 = f_arrdiv24_fs504_and0 ^ f_arrdiv24_fs505_xor0;
  assign f_arrdiv24_fs505_not1 = ~f_arrdiv24_fs505_xor0;
  assign f_arrdiv24_fs505_and1 = f_arrdiv24_fs505_not1 & f_arrdiv24_fs504_and0;
  assign f_arrdiv24_fs505_or0 = f_arrdiv24_fs505_and1 | f_arrdiv24_fs505_and0;
  assign f_arrdiv24_fs506_xor0 = f_arrdiv24_mux2to1461_xor0 ^ b[2];
  assign f_arrdiv24_fs506_not0 = ~f_arrdiv24_mux2to1461_xor0;
  assign f_arrdiv24_fs506_and0 = f_arrdiv24_fs506_not0 & b[2];
  assign f_arrdiv24_fs506_xor1 = f_arrdiv24_fs505_or0 ^ f_arrdiv24_fs506_xor0;
  assign f_arrdiv24_fs506_not1 = ~f_arrdiv24_fs506_xor0;
  assign f_arrdiv24_fs506_and1 = f_arrdiv24_fs506_not1 & f_arrdiv24_fs505_or0;
  assign f_arrdiv24_fs506_or0 = f_arrdiv24_fs506_and1 | f_arrdiv24_fs506_and0;
  assign f_arrdiv24_fs507_xor0 = f_arrdiv24_mux2to1462_xor0 ^ b[3];
  assign f_arrdiv24_fs507_not0 = ~f_arrdiv24_mux2to1462_xor0;
  assign f_arrdiv24_fs507_and0 = f_arrdiv24_fs507_not0 & b[3];
  assign f_arrdiv24_fs507_xor1 = f_arrdiv24_fs506_or0 ^ f_arrdiv24_fs507_xor0;
  assign f_arrdiv24_fs507_not1 = ~f_arrdiv24_fs507_xor0;
  assign f_arrdiv24_fs507_and1 = f_arrdiv24_fs507_not1 & f_arrdiv24_fs506_or0;
  assign f_arrdiv24_fs507_or0 = f_arrdiv24_fs507_and1 | f_arrdiv24_fs507_and0;
  assign f_arrdiv24_fs508_xor0 = f_arrdiv24_mux2to1463_xor0 ^ b[4];
  assign f_arrdiv24_fs508_not0 = ~f_arrdiv24_mux2to1463_xor0;
  assign f_arrdiv24_fs508_and0 = f_arrdiv24_fs508_not0 & b[4];
  assign f_arrdiv24_fs508_xor1 = f_arrdiv24_fs507_or0 ^ f_arrdiv24_fs508_xor0;
  assign f_arrdiv24_fs508_not1 = ~f_arrdiv24_fs508_xor0;
  assign f_arrdiv24_fs508_and1 = f_arrdiv24_fs508_not1 & f_arrdiv24_fs507_or0;
  assign f_arrdiv24_fs508_or0 = f_arrdiv24_fs508_and1 | f_arrdiv24_fs508_and0;
  assign f_arrdiv24_fs509_xor0 = f_arrdiv24_mux2to1464_xor0 ^ b[5];
  assign f_arrdiv24_fs509_not0 = ~f_arrdiv24_mux2to1464_xor0;
  assign f_arrdiv24_fs509_and0 = f_arrdiv24_fs509_not0 & b[5];
  assign f_arrdiv24_fs509_xor1 = f_arrdiv24_fs508_or0 ^ f_arrdiv24_fs509_xor0;
  assign f_arrdiv24_fs509_not1 = ~f_arrdiv24_fs509_xor0;
  assign f_arrdiv24_fs509_and1 = f_arrdiv24_fs509_not1 & f_arrdiv24_fs508_or0;
  assign f_arrdiv24_fs509_or0 = f_arrdiv24_fs509_and1 | f_arrdiv24_fs509_and0;
  assign f_arrdiv24_fs510_xor0 = f_arrdiv24_mux2to1465_xor0 ^ b[6];
  assign f_arrdiv24_fs510_not0 = ~f_arrdiv24_mux2to1465_xor0;
  assign f_arrdiv24_fs510_and0 = f_arrdiv24_fs510_not0 & b[6];
  assign f_arrdiv24_fs510_xor1 = f_arrdiv24_fs509_or0 ^ f_arrdiv24_fs510_xor0;
  assign f_arrdiv24_fs510_not1 = ~f_arrdiv24_fs510_xor0;
  assign f_arrdiv24_fs510_and1 = f_arrdiv24_fs510_not1 & f_arrdiv24_fs509_or0;
  assign f_arrdiv24_fs510_or0 = f_arrdiv24_fs510_and1 | f_arrdiv24_fs510_and0;
  assign f_arrdiv24_fs511_xor0 = f_arrdiv24_mux2to1466_xor0 ^ b[7];
  assign f_arrdiv24_fs511_not0 = ~f_arrdiv24_mux2to1466_xor0;
  assign f_arrdiv24_fs511_and0 = f_arrdiv24_fs511_not0 & b[7];
  assign f_arrdiv24_fs511_xor1 = f_arrdiv24_fs510_or0 ^ f_arrdiv24_fs511_xor0;
  assign f_arrdiv24_fs511_not1 = ~f_arrdiv24_fs511_xor0;
  assign f_arrdiv24_fs511_and1 = f_arrdiv24_fs511_not1 & f_arrdiv24_fs510_or0;
  assign f_arrdiv24_fs511_or0 = f_arrdiv24_fs511_and1 | f_arrdiv24_fs511_and0;
  assign f_arrdiv24_fs512_xor0 = f_arrdiv24_mux2to1467_xor0 ^ b[8];
  assign f_arrdiv24_fs512_not0 = ~f_arrdiv24_mux2to1467_xor0;
  assign f_arrdiv24_fs512_and0 = f_arrdiv24_fs512_not0 & b[8];
  assign f_arrdiv24_fs512_xor1 = f_arrdiv24_fs511_or0 ^ f_arrdiv24_fs512_xor0;
  assign f_arrdiv24_fs512_not1 = ~f_arrdiv24_fs512_xor0;
  assign f_arrdiv24_fs512_and1 = f_arrdiv24_fs512_not1 & f_arrdiv24_fs511_or0;
  assign f_arrdiv24_fs512_or0 = f_arrdiv24_fs512_and1 | f_arrdiv24_fs512_and0;
  assign f_arrdiv24_fs513_xor0 = f_arrdiv24_mux2to1468_xor0 ^ b[9];
  assign f_arrdiv24_fs513_not0 = ~f_arrdiv24_mux2to1468_xor0;
  assign f_arrdiv24_fs513_and0 = f_arrdiv24_fs513_not0 & b[9];
  assign f_arrdiv24_fs513_xor1 = f_arrdiv24_fs512_or0 ^ f_arrdiv24_fs513_xor0;
  assign f_arrdiv24_fs513_not1 = ~f_arrdiv24_fs513_xor0;
  assign f_arrdiv24_fs513_and1 = f_arrdiv24_fs513_not1 & f_arrdiv24_fs512_or0;
  assign f_arrdiv24_fs513_or0 = f_arrdiv24_fs513_and1 | f_arrdiv24_fs513_and0;
  assign f_arrdiv24_fs514_xor0 = f_arrdiv24_mux2to1469_xor0 ^ b[10];
  assign f_arrdiv24_fs514_not0 = ~f_arrdiv24_mux2to1469_xor0;
  assign f_arrdiv24_fs514_and0 = f_arrdiv24_fs514_not0 & b[10];
  assign f_arrdiv24_fs514_xor1 = f_arrdiv24_fs513_or0 ^ f_arrdiv24_fs514_xor0;
  assign f_arrdiv24_fs514_not1 = ~f_arrdiv24_fs514_xor0;
  assign f_arrdiv24_fs514_and1 = f_arrdiv24_fs514_not1 & f_arrdiv24_fs513_or0;
  assign f_arrdiv24_fs514_or0 = f_arrdiv24_fs514_and1 | f_arrdiv24_fs514_and0;
  assign f_arrdiv24_fs515_xor0 = f_arrdiv24_mux2to1470_xor0 ^ b[11];
  assign f_arrdiv24_fs515_not0 = ~f_arrdiv24_mux2to1470_xor0;
  assign f_arrdiv24_fs515_and0 = f_arrdiv24_fs515_not0 & b[11];
  assign f_arrdiv24_fs515_xor1 = f_arrdiv24_fs514_or0 ^ f_arrdiv24_fs515_xor0;
  assign f_arrdiv24_fs515_not1 = ~f_arrdiv24_fs515_xor0;
  assign f_arrdiv24_fs515_and1 = f_arrdiv24_fs515_not1 & f_arrdiv24_fs514_or0;
  assign f_arrdiv24_fs515_or0 = f_arrdiv24_fs515_and1 | f_arrdiv24_fs515_and0;
  assign f_arrdiv24_fs516_xor0 = f_arrdiv24_mux2to1471_xor0 ^ b[12];
  assign f_arrdiv24_fs516_not0 = ~f_arrdiv24_mux2to1471_xor0;
  assign f_arrdiv24_fs516_and0 = f_arrdiv24_fs516_not0 & b[12];
  assign f_arrdiv24_fs516_xor1 = f_arrdiv24_fs515_or0 ^ f_arrdiv24_fs516_xor0;
  assign f_arrdiv24_fs516_not1 = ~f_arrdiv24_fs516_xor0;
  assign f_arrdiv24_fs516_and1 = f_arrdiv24_fs516_not1 & f_arrdiv24_fs515_or0;
  assign f_arrdiv24_fs516_or0 = f_arrdiv24_fs516_and1 | f_arrdiv24_fs516_and0;
  assign f_arrdiv24_fs517_xor0 = f_arrdiv24_mux2to1472_xor0 ^ b[13];
  assign f_arrdiv24_fs517_not0 = ~f_arrdiv24_mux2to1472_xor0;
  assign f_arrdiv24_fs517_and0 = f_arrdiv24_fs517_not0 & b[13];
  assign f_arrdiv24_fs517_xor1 = f_arrdiv24_fs516_or0 ^ f_arrdiv24_fs517_xor0;
  assign f_arrdiv24_fs517_not1 = ~f_arrdiv24_fs517_xor0;
  assign f_arrdiv24_fs517_and1 = f_arrdiv24_fs517_not1 & f_arrdiv24_fs516_or0;
  assign f_arrdiv24_fs517_or0 = f_arrdiv24_fs517_and1 | f_arrdiv24_fs517_and0;
  assign f_arrdiv24_fs518_xor0 = f_arrdiv24_mux2to1473_xor0 ^ b[14];
  assign f_arrdiv24_fs518_not0 = ~f_arrdiv24_mux2to1473_xor0;
  assign f_arrdiv24_fs518_and0 = f_arrdiv24_fs518_not0 & b[14];
  assign f_arrdiv24_fs518_xor1 = f_arrdiv24_fs517_or0 ^ f_arrdiv24_fs518_xor0;
  assign f_arrdiv24_fs518_not1 = ~f_arrdiv24_fs518_xor0;
  assign f_arrdiv24_fs518_and1 = f_arrdiv24_fs518_not1 & f_arrdiv24_fs517_or0;
  assign f_arrdiv24_fs518_or0 = f_arrdiv24_fs518_and1 | f_arrdiv24_fs518_and0;
  assign f_arrdiv24_fs519_xor0 = f_arrdiv24_mux2to1474_xor0 ^ b[15];
  assign f_arrdiv24_fs519_not0 = ~f_arrdiv24_mux2to1474_xor0;
  assign f_arrdiv24_fs519_and0 = f_arrdiv24_fs519_not0 & b[15];
  assign f_arrdiv24_fs519_xor1 = f_arrdiv24_fs518_or0 ^ f_arrdiv24_fs519_xor0;
  assign f_arrdiv24_fs519_not1 = ~f_arrdiv24_fs519_xor0;
  assign f_arrdiv24_fs519_and1 = f_arrdiv24_fs519_not1 & f_arrdiv24_fs518_or0;
  assign f_arrdiv24_fs519_or0 = f_arrdiv24_fs519_and1 | f_arrdiv24_fs519_and0;
  assign f_arrdiv24_fs520_xor0 = f_arrdiv24_mux2to1475_xor0 ^ b[16];
  assign f_arrdiv24_fs520_not0 = ~f_arrdiv24_mux2to1475_xor0;
  assign f_arrdiv24_fs520_and0 = f_arrdiv24_fs520_not0 & b[16];
  assign f_arrdiv24_fs520_xor1 = f_arrdiv24_fs519_or0 ^ f_arrdiv24_fs520_xor0;
  assign f_arrdiv24_fs520_not1 = ~f_arrdiv24_fs520_xor0;
  assign f_arrdiv24_fs520_and1 = f_arrdiv24_fs520_not1 & f_arrdiv24_fs519_or0;
  assign f_arrdiv24_fs520_or0 = f_arrdiv24_fs520_and1 | f_arrdiv24_fs520_and0;
  assign f_arrdiv24_fs521_xor0 = f_arrdiv24_mux2to1476_xor0 ^ b[17];
  assign f_arrdiv24_fs521_not0 = ~f_arrdiv24_mux2to1476_xor0;
  assign f_arrdiv24_fs521_and0 = f_arrdiv24_fs521_not0 & b[17];
  assign f_arrdiv24_fs521_xor1 = f_arrdiv24_fs520_or0 ^ f_arrdiv24_fs521_xor0;
  assign f_arrdiv24_fs521_not1 = ~f_arrdiv24_fs521_xor0;
  assign f_arrdiv24_fs521_and1 = f_arrdiv24_fs521_not1 & f_arrdiv24_fs520_or0;
  assign f_arrdiv24_fs521_or0 = f_arrdiv24_fs521_and1 | f_arrdiv24_fs521_and0;
  assign f_arrdiv24_fs522_xor0 = f_arrdiv24_mux2to1477_xor0 ^ b[18];
  assign f_arrdiv24_fs522_not0 = ~f_arrdiv24_mux2to1477_xor0;
  assign f_arrdiv24_fs522_and0 = f_arrdiv24_fs522_not0 & b[18];
  assign f_arrdiv24_fs522_xor1 = f_arrdiv24_fs521_or0 ^ f_arrdiv24_fs522_xor0;
  assign f_arrdiv24_fs522_not1 = ~f_arrdiv24_fs522_xor0;
  assign f_arrdiv24_fs522_and1 = f_arrdiv24_fs522_not1 & f_arrdiv24_fs521_or0;
  assign f_arrdiv24_fs522_or0 = f_arrdiv24_fs522_and1 | f_arrdiv24_fs522_and0;
  assign f_arrdiv24_fs523_xor0 = f_arrdiv24_mux2to1478_xor0 ^ b[19];
  assign f_arrdiv24_fs523_not0 = ~f_arrdiv24_mux2to1478_xor0;
  assign f_arrdiv24_fs523_and0 = f_arrdiv24_fs523_not0 & b[19];
  assign f_arrdiv24_fs523_xor1 = f_arrdiv24_fs522_or0 ^ f_arrdiv24_fs523_xor0;
  assign f_arrdiv24_fs523_not1 = ~f_arrdiv24_fs523_xor0;
  assign f_arrdiv24_fs523_and1 = f_arrdiv24_fs523_not1 & f_arrdiv24_fs522_or0;
  assign f_arrdiv24_fs523_or0 = f_arrdiv24_fs523_and1 | f_arrdiv24_fs523_and0;
  assign f_arrdiv24_fs524_xor0 = f_arrdiv24_mux2to1479_xor0 ^ b[20];
  assign f_arrdiv24_fs524_not0 = ~f_arrdiv24_mux2to1479_xor0;
  assign f_arrdiv24_fs524_and0 = f_arrdiv24_fs524_not0 & b[20];
  assign f_arrdiv24_fs524_xor1 = f_arrdiv24_fs523_or0 ^ f_arrdiv24_fs524_xor0;
  assign f_arrdiv24_fs524_not1 = ~f_arrdiv24_fs524_xor0;
  assign f_arrdiv24_fs524_and1 = f_arrdiv24_fs524_not1 & f_arrdiv24_fs523_or0;
  assign f_arrdiv24_fs524_or0 = f_arrdiv24_fs524_and1 | f_arrdiv24_fs524_and0;
  assign f_arrdiv24_fs525_xor0 = f_arrdiv24_mux2to1480_xor0 ^ b[21];
  assign f_arrdiv24_fs525_not0 = ~f_arrdiv24_mux2to1480_xor0;
  assign f_arrdiv24_fs525_and0 = f_arrdiv24_fs525_not0 & b[21];
  assign f_arrdiv24_fs525_xor1 = f_arrdiv24_fs524_or0 ^ f_arrdiv24_fs525_xor0;
  assign f_arrdiv24_fs525_not1 = ~f_arrdiv24_fs525_xor0;
  assign f_arrdiv24_fs525_and1 = f_arrdiv24_fs525_not1 & f_arrdiv24_fs524_or0;
  assign f_arrdiv24_fs525_or0 = f_arrdiv24_fs525_and1 | f_arrdiv24_fs525_and0;
  assign f_arrdiv24_fs526_xor0 = f_arrdiv24_mux2to1481_xor0 ^ b[22];
  assign f_arrdiv24_fs526_not0 = ~f_arrdiv24_mux2to1481_xor0;
  assign f_arrdiv24_fs526_and0 = f_arrdiv24_fs526_not0 & b[22];
  assign f_arrdiv24_fs526_xor1 = f_arrdiv24_fs525_or0 ^ f_arrdiv24_fs526_xor0;
  assign f_arrdiv24_fs526_not1 = ~f_arrdiv24_fs526_xor0;
  assign f_arrdiv24_fs526_and1 = f_arrdiv24_fs526_not1 & f_arrdiv24_fs525_or0;
  assign f_arrdiv24_fs526_or0 = f_arrdiv24_fs526_and1 | f_arrdiv24_fs526_and0;
  assign f_arrdiv24_fs527_xor0 = f_arrdiv24_mux2to1482_xor0 ^ b[23];
  assign f_arrdiv24_fs527_not0 = ~f_arrdiv24_mux2to1482_xor0;
  assign f_arrdiv24_fs527_and0 = f_arrdiv24_fs527_not0 & b[23];
  assign f_arrdiv24_fs527_xor1 = f_arrdiv24_fs526_or0 ^ f_arrdiv24_fs527_xor0;
  assign f_arrdiv24_fs527_not1 = ~f_arrdiv24_fs527_xor0;
  assign f_arrdiv24_fs527_and1 = f_arrdiv24_fs527_not1 & f_arrdiv24_fs526_or0;
  assign f_arrdiv24_fs527_or0 = f_arrdiv24_fs527_and1 | f_arrdiv24_fs527_and0;
  assign f_arrdiv24_mux2to1483_and0 = a[2] & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1483_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1483_and1 = f_arrdiv24_fs504_xor0 & f_arrdiv24_mux2to1483_not0;
  assign f_arrdiv24_mux2to1483_xor0 = f_arrdiv24_mux2to1483_and0 ^ f_arrdiv24_mux2to1483_and1;
  assign f_arrdiv24_mux2to1484_and0 = f_arrdiv24_mux2to1460_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1484_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1484_and1 = f_arrdiv24_fs505_xor1 & f_arrdiv24_mux2to1484_not0;
  assign f_arrdiv24_mux2to1484_xor0 = f_arrdiv24_mux2to1484_and0 ^ f_arrdiv24_mux2to1484_and1;
  assign f_arrdiv24_mux2to1485_and0 = f_arrdiv24_mux2to1461_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1485_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1485_and1 = f_arrdiv24_fs506_xor1 & f_arrdiv24_mux2to1485_not0;
  assign f_arrdiv24_mux2to1485_xor0 = f_arrdiv24_mux2to1485_and0 ^ f_arrdiv24_mux2to1485_and1;
  assign f_arrdiv24_mux2to1486_and0 = f_arrdiv24_mux2to1462_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1486_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1486_and1 = f_arrdiv24_fs507_xor1 & f_arrdiv24_mux2to1486_not0;
  assign f_arrdiv24_mux2to1486_xor0 = f_arrdiv24_mux2to1486_and0 ^ f_arrdiv24_mux2to1486_and1;
  assign f_arrdiv24_mux2to1487_and0 = f_arrdiv24_mux2to1463_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1487_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1487_and1 = f_arrdiv24_fs508_xor1 & f_arrdiv24_mux2to1487_not0;
  assign f_arrdiv24_mux2to1487_xor0 = f_arrdiv24_mux2to1487_and0 ^ f_arrdiv24_mux2to1487_and1;
  assign f_arrdiv24_mux2to1488_and0 = f_arrdiv24_mux2to1464_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1488_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1488_and1 = f_arrdiv24_fs509_xor1 & f_arrdiv24_mux2to1488_not0;
  assign f_arrdiv24_mux2to1488_xor0 = f_arrdiv24_mux2to1488_and0 ^ f_arrdiv24_mux2to1488_and1;
  assign f_arrdiv24_mux2to1489_and0 = f_arrdiv24_mux2to1465_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1489_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1489_and1 = f_arrdiv24_fs510_xor1 & f_arrdiv24_mux2to1489_not0;
  assign f_arrdiv24_mux2to1489_xor0 = f_arrdiv24_mux2to1489_and0 ^ f_arrdiv24_mux2to1489_and1;
  assign f_arrdiv24_mux2to1490_and0 = f_arrdiv24_mux2to1466_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1490_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1490_and1 = f_arrdiv24_fs511_xor1 & f_arrdiv24_mux2to1490_not0;
  assign f_arrdiv24_mux2to1490_xor0 = f_arrdiv24_mux2to1490_and0 ^ f_arrdiv24_mux2to1490_and1;
  assign f_arrdiv24_mux2to1491_and0 = f_arrdiv24_mux2to1467_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1491_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1491_and1 = f_arrdiv24_fs512_xor1 & f_arrdiv24_mux2to1491_not0;
  assign f_arrdiv24_mux2to1491_xor0 = f_arrdiv24_mux2to1491_and0 ^ f_arrdiv24_mux2to1491_and1;
  assign f_arrdiv24_mux2to1492_and0 = f_arrdiv24_mux2to1468_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1492_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1492_and1 = f_arrdiv24_fs513_xor1 & f_arrdiv24_mux2to1492_not0;
  assign f_arrdiv24_mux2to1492_xor0 = f_arrdiv24_mux2to1492_and0 ^ f_arrdiv24_mux2to1492_and1;
  assign f_arrdiv24_mux2to1493_and0 = f_arrdiv24_mux2to1469_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1493_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1493_and1 = f_arrdiv24_fs514_xor1 & f_arrdiv24_mux2to1493_not0;
  assign f_arrdiv24_mux2to1493_xor0 = f_arrdiv24_mux2to1493_and0 ^ f_arrdiv24_mux2to1493_and1;
  assign f_arrdiv24_mux2to1494_and0 = f_arrdiv24_mux2to1470_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1494_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1494_and1 = f_arrdiv24_fs515_xor1 & f_arrdiv24_mux2to1494_not0;
  assign f_arrdiv24_mux2to1494_xor0 = f_arrdiv24_mux2to1494_and0 ^ f_arrdiv24_mux2to1494_and1;
  assign f_arrdiv24_mux2to1495_and0 = f_arrdiv24_mux2to1471_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1495_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1495_and1 = f_arrdiv24_fs516_xor1 & f_arrdiv24_mux2to1495_not0;
  assign f_arrdiv24_mux2to1495_xor0 = f_arrdiv24_mux2to1495_and0 ^ f_arrdiv24_mux2to1495_and1;
  assign f_arrdiv24_mux2to1496_and0 = f_arrdiv24_mux2to1472_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1496_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1496_and1 = f_arrdiv24_fs517_xor1 & f_arrdiv24_mux2to1496_not0;
  assign f_arrdiv24_mux2to1496_xor0 = f_arrdiv24_mux2to1496_and0 ^ f_arrdiv24_mux2to1496_and1;
  assign f_arrdiv24_mux2to1497_and0 = f_arrdiv24_mux2to1473_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1497_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1497_and1 = f_arrdiv24_fs518_xor1 & f_arrdiv24_mux2to1497_not0;
  assign f_arrdiv24_mux2to1497_xor0 = f_arrdiv24_mux2to1497_and0 ^ f_arrdiv24_mux2to1497_and1;
  assign f_arrdiv24_mux2to1498_and0 = f_arrdiv24_mux2to1474_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1498_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1498_and1 = f_arrdiv24_fs519_xor1 & f_arrdiv24_mux2to1498_not0;
  assign f_arrdiv24_mux2to1498_xor0 = f_arrdiv24_mux2to1498_and0 ^ f_arrdiv24_mux2to1498_and1;
  assign f_arrdiv24_mux2to1499_and0 = f_arrdiv24_mux2to1475_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1499_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1499_and1 = f_arrdiv24_fs520_xor1 & f_arrdiv24_mux2to1499_not0;
  assign f_arrdiv24_mux2to1499_xor0 = f_arrdiv24_mux2to1499_and0 ^ f_arrdiv24_mux2to1499_and1;
  assign f_arrdiv24_mux2to1500_and0 = f_arrdiv24_mux2to1476_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1500_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1500_and1 = f_arrdiv24_fs521_xor1 & f_arrdiv24_mux2to1500_not0;
  assign f_arrdiv24_mux2to1500_xor0 = f_arrdiv24_mux2to1500_and0 ^ f_arrdiv24_mux2to1500_and1;
  assign f_arrdiv24_mux2to1501_and0 = f_arrdiv24_mux2to1477_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1501_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1501_and1 = f_arrdiv24_fs522_xor1 & f_arrdiv24_mux2to1501_not0;
  assign f_arrdiv24_mux2to1501_xor0 = f_arrdiv24_mux2to1501_and0 ^ f_arrdiv24_mux2to1501_and1;
  assign f_arrdiv24_mux2to1502_and0 = f_arrdiv24_mux2to1478_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1502_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1502_and1 = f_arrdiv24_fs523_xor1 & f_arrdiv24_mux2to1502_not0;
  assign f_arrdiv24_mux2to1502_xor0 = f_arrdiv24_mux2to1502_and0 ^ f_arrdiv24_mux2to1502_and1;
  assign f_arrdiv24_mux2to1503_and0 = f_arrdiv24_mux2to1479_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1503_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1503_and1 = f_arrdiv24_fs524_xor1 & f_arrdiv24_mux2to1503_not0;
  assign f_arrdiv24_mux2to1503_xor0 = f_arrdiv24_mux2to1503_and0 ^ f_arrdiv24_mux2to1503_and1;
  assign f_arrdiv24_mux2to1504_and0 = f_arrdiv24_mux2to1480_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1504_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1504_and1 = f_arrdiv24_fs525_xor1 & f_arrdiv24_mux2to1504_not0;
  assign f_arrdiv24_mux2to1504_xor0 = f_arrdiv24_mux2to1504_and0 ^ f_arrdiv24_mux2to1504_and1;
  assign f_arrdiv24_mux2to1505_and0 = f_arrdiv24_mux2to1481_xor0 & f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1505_not0 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_mux2to1505_and1 = f_arrdiv24_fs526_xor1 & f_arrdiv24_mux2to1505_not0;
  assign f_arrdiv24_mux2to1505_xor0 = f_arrdiv24_mux2to1505_and0 ^ f_arrdiv24_mux2to1505_and1;
  assign f_arrdiv24_not21 = ~f_arrdiv24_fs527_or0;
  assign f_arrdiv24_fs528_xor0 = a[1] ^ b[0];
  assign f_arrdiv24_fs528_not0 = ~a[1];
  assign f_arrdiv24_fs528_and0 = f_arrdiv24_fs528_not0 & b[0];
  assign f_arrdiv24_fs528_not1 = ~f_arrdiv24_fs528_xor0;
  assign f_arrdiv24_fs529_xor0 = f_arrdiv24_mux2to1483_xor0 ^ b[1];
  assign f_arrdiv24_fs529_not0 = ~f_arrdiv24_mux2to1483_xor0;
  assign f_arrdiv24_fs529_and0 = f_arrdiv24_fs529_not0 & b[1];
  assign f_arrdiv24_fs529_xor1 = f_arrdiv24_fs528_and0 ^ f_arrdiv24_fs529_xor0;
  assign f_arrdiv24_fs529_not1 = ~f_arrdiv24_fs529_xor0;
  assign f_arrdiv24_fs529_and1 = f_arrdiv24_fs529_not1 & f_arrdiv24_fs528_and0;
  assign f_arrdiv24_fs529_or0 = f_arrdiv24_fs529_and1 | f_arrdiv24_fs529_and0;
  assign f_arrdiv24_fs530_xor0 = f_arrdiv24_mux2to1484_xor0 ^ b[2];
  assign f_arrdiv24_fs530_not0 = ~f_arrdiv24_mux2to1484_xor0;
  assign f_arrdiv24_fs530_and0 = f_arrdiv24_fs530_not0 & b[2];
  assign f_arrdiv24_fs530_xor1 = f_arrdiv24_fs529_or0 ^ f_arrdiv24_fs530_xor0;
  assign f_arrdiv24_fs530_not1 = ~f_arrdiv24_fs530_xor0;
  assign f_arrdiv24_fs530_and1 = f_arrdiv24_fs530_not1 & f_arrdiv24_fs529_or0;
  assign f_arrdiv24_fs530_or0 = f_arrdiv24_fs530_and1 | f_arrdiv24_fs530_and0;
  assign f_arrdiv24_fs531_xor0 = f_arrdiv24_mux2to1485_xor0 ^ b[3];
  assign f_arrdiv24_fs531_not0 = ~f_arrdiv24_mux2to1485_xor0;
  assign f_arrdiv24_fs531_and0 = f_arrdiv24_fs531_not0 & b[3];
  assign f_arrdiv24_fs531_xor1 = f_arrdiv24_fs530_or0 ^ f_arrdiv24_fs531_xor0;
  assign f_arrdiv24_fs531_not1 = ~f_arrdiv24_fs531_xor0;
  assign f_arrdiv24_fs531_and1 = f_arrdiv24_fs531_not1 & f_arrdiv24_fs530_or0;
  assign f_arrdiv24_fs531_or0 = f_arrdiv24_fs531_and1 | f_arrdiv24_fs531_and0;
  assign f_arrdiv24_fs532_xor0 = f_arrdiv24_mux2to1486_xor0 ^ b[4];
  assign f_arrdiv24_fs532_not0 = ~f_arrdiv24_mux2to1486_xor0;
  assign f_arrdiv24_fs532_and0 = f_arrdiv24_fs532_not0 & b[4];
  assign f_arrdiv24_fs532_xor1 = f_arrdiv24_fs531_or0 ^ f_arrdiv24_fs532_xor0;
  assign f_arrdiv24_fs532_not1 = ~f_arrdiv24_fs532_xor0;
  assign f_arrdiv24_fs532_and1 = f_arrdiv24_fs532_not1 & f_arrdiv24_fs531_or0;
  assign f_arrdiv24_fs532_or0 = f_arrdiv24_fs532_and1 | f_arrdiv24_fs532_and0;
  assign f_arrdiv24_fs533_xor0 = f_arrdiv24_mux2to1487_xor0 ^ b[5];
  assign f_arrdiv24_fs533_not0 = ~f_arrdiv24_mux2to1487_xor0;
  assign f_arrdiv24_fs533_and0 = f_arrdiv24_fs533_not0 & b[5];
  assign f_arrdiv24_fs533_xor1 = f_arrdiv24_fs532_or0 ^ f_arrdiv24_fs533_xor0;
  assign f_arrdiv24_fs533_not1 = ~f_arrdiv24_fs533_xor0;
  assign f_arrdiv24_fs533_and1 = f_arrdiv24_fs533_not1 & f_arrdiv24_fs532_or0;
  assign f_arrdiv24_fs533_or0 = f_arrdiv24_fs533_and1 | f_arrdiv24_fs533_and0;
  assign f_arrdiv24_fs534_xor0 = f_arrdiv24_mux2to1488_xor0 ^ b[6];
  assign f_arrdiv24_fs534_not0 = ~f_arrdiv24_mux2to1488_xor0;
  assign f_arrdiv24_fs534_and0 = f_arrdiv24_fs534_not0 & b[6];
  assign f_arrdiv24_fs534_xor1 = f_arrdiv24_fs533_or0 ^ f_arrdiv24_fs534_xor0;
  assign f_arrdiv24_fs534_not1 = ~f_arrdiv24_fs534_xor0;
  assign f_arrdiv24_fs534_and1 = f_arrdiv24_fs534_not1 & f_arrdiv24_fs533_or0;
  assign f_arrdiv24_fs534_or0 = f_arrdiv24_fs534_and1 | f_arrdiv24_fs534_and0;
  assign f_arrdiv24_fs535_xor0 = f_arrdiv24_mux2to1489_xor0 ^ b[7];
  assign f_arrdiv24_fs535_not0 = ~f_arrdiv24_mux2to1489_xor0;
  assign f_arrdiv24_fs535_and0 = f_arrdiv24_fs535_not0 & b[7];
  assign f_arrdiv24_fs535_xor1 = f_arrdiv24_fs534_or0 ^ f_arrdiv24_fs535_xor0;
  assign f_arrdiv24_fs535_not1 = ~f_arrdiv24_fs535_xor0;
  assign f_arrdiv24_fs535_and1 = f_arrdiv24_fs535_not1 & f_arrdiv24_fs534_or0;
  assign f_arrdiv24_fs535_or0 = f_arrdiv24_fs535_and1 | f_arrdiv24_fs535_and0;
  assign f_arrdiv24_fs536_xor0 = f_arrdiv24_mux2to1490_xor0 ^ b[8];
  assign f_arrdiv24_fs536_not0 = ~f_arrdiv24_mux2to1490_xor0;
  assign f_arrdiv24_fs536_and0 = f_arrdiv24_fs536_not0 & b[8];
  assign f_arrdiv24_fs536_xor1 = f_arrdiv24_fs535_or0 ^ f_arrdiv24_fs536_xor0;
  assign f_arrdiv24_fs536_not1 = ~f_arrdiv24_fs536_xor0;
  assign f_arrdiv24_fs536_and1 = f_arrdiv24_fs536_not1 & f_arrdiv24_fs535_or0;
  assign f_arrdiv24_fs536_or0 = f_arrdiv24_fs536_and1 | f_arrdiv24_fs536_and0;
  assign f_arrdiv24_fs537_xor0 = f_arrdiv24_mux2to1491_xor0 ^ b[9];
  assign f_arrdiv24_fs537_not0 = ~f_arrdiv24_mux2to1491_xor0;
  assign f_arrdiv24_fs537_and0 = f_arrdiv24_fs537_not0 & b[9];
  assign f_arrdiv24_fs537_xor1 = f_arrdiv24_fs536_or0 ^ f_arrdiv24_fs537_xor0;
  assign f_arrdiv24_fs537_not1 = ~f_arrdiv24_fs537_xor0;
  assign f_arrdiv24_fs537_and1 = f_arrdiv24_fs537_not1 & f_arrdiv24_fs536_or0;
  assign f_arrdiv24_fs537_or0 = f_arrdiv24_fs537_and1 | f_arrdiv24_fs537_and0;
  assign f_arrdiv24_fs538_xor0 = f_arrdiv24_mux2to1492_xor0 ^ b[10];
  assign f_arrdiv24_fs538_not0 = ~f_arrdiv24_mux2to1492_xor0;
  assign f_arrdiv24_fs538_and0 = f_arrdiv24_fs538_not0 & b[10];
  assign f_arrdiv24_fs538_xor1 = f_arrdiv24_fs537_or0 ^ f_arrdiv24_fs538_xor0;
  assign f_arrdiv24_fs538_not1 = ~f_arrdiv24_fs538_xor0;
  assign f_arrdiv24_fs538_and1 = f_arrdiv24_fs538_not1 & f_arrdiv24_fs537_or0;
  assign f_arrdiv24_fs538_or0 = f_arrdiv24_fs538_and1 | f_arrdiv24_fs538_and0;
  assign f_arrdiv24_fs539_xor0 = f_arrdiv24_mux2to1493_xor0 ^ b[11];
  assign f_arrdiv24_fs539_not0 = ~f_arrdiv24_mux2to1493_xor0;
  assign f_arrdiv24_fs539_and0 = f_arrdiv24_fs539_not0 & b[11];
  assign f_arrdiv24_fs539_xor1 = f_arrdiv24_fs538_or0 ^ f_arrdiv24_fs539_xor0;
  assign f_arrdiv24_fs539_not1 = ~f_arrdiv24_fs539_xor0;
  assign f_arrdiv24_fs539_and1 = f_arrdiv24_fs539_not1 & f_arrdiv24_fs538_or0;
  assign f_arrdiv24_fs539_or0 = f_arrdiv24_fs539_and1 | f_arrdiv24_fs539_and0;
  assign f_arrdiv24_fs540_xor0 = f_arrdiv24_mux2to1494_xor0 ^ b[12];
  assign f_arrdiv24_fs540_not0 = ~f_arrdiv24_mux2to1494_xor0;
  assign f_arrdiv24_fs540_and0 = f_arrdiv24_fs540_not0 & b[12];
  assign f_arrdiv24_fs540_xor1 = f_arrdiv24_fs539_or0 ^ f_arrdiv24_fs540_xor0;
  assign f_arrdiv24_fs540_not1 = ~f_arrdiv24_fs540_xor0;
  assign f_arrdiv24_fs540_and1 = f_arrdiv24_fs540_not1 & f_arrdiv24_fs539_or0;
  assign f_arrdiv24_fs540_or0 = f_arrdiv24_fs540_and1 | f_arrdiv24_fs540_and0;
  assign f_arrdiv24_fs541_xor0 = f_arrdiv24_mux2to1495_xor0 ^ b[13];
  assign f_arrdiv24_fs541_not0 = ~f_arrdiv24_mux2to1495_xor0;
  assign f_arrdiv24_fs541_and0 = f_arrdiv24_fs541_not0 & b[13];
  assign f_arrdiv24_fs541_xor1 = f_arrdiv24_fs540_or0 ^ f_arrdiv24_fs541_xor0;
  assign f_arrdiv24_fs541_not1 = ~f_arrdiv24_fs541_xor0;
  assign f_arrdiv24_fs541_and1 = f_arrdiv24_fs541_not1 & f_arrdiv24_fs540_or0;
  assign f_arrdiv24_fs541_or0 = f_arrdiv24_fs541_and1 | f_arrdiv24_fs541_and0;
  assign f_arrdiv24_fs542_xor0 = f_arrdiv24_mux2to1496_xor0 ^ b[14];
  assign f_arrdiv24_fs542_not0 = ~f_arrdiv24_mux2to1496_xor0;
  assign f_arrdiv24_fs542_and0 = f_arrdiv24_fs542_not0 & b[14];
  assign f_arrdiv24_fs542_xor1 = f_arrdiv24_fs541_or0 ^ f_arrdiv24_fs542_xor0;
  assign f_arrdiv24_fs542_not1 = ~f_arrdiv24_fs542_xor0;
  assign f_arrdiv24_fs542_and1 = f_arrdiv24_fs542_not1 & f_arrdiv24_fs541_or0;
  assign f_arrdiv24_fs542_or0 = f_arrdiv24_fs542_and1 | f_arrdiv24_fs542_and0;
  assign f_arrdiv24_fs543_xor0 = f_arrdiv24_mux2to1497_xor0 ^ b[15];
  assign f_arrdiv24_fs543_not0 = ~f_arrdiv24_mux2to1497_xor0;
  assign f_arrdiv24_fs543_and0 = f_arrdiv24_fs543_not0 & b[15];
  assign f_arrdiv24_fs543_xor1 = f_arrdiv24_fs542_or0 ^ f_arrdiv24_fs543_xor0;
  assign f_arrdiv24_fs543_not1 = ~f_arrdiv24_fs543_xor0;
  assign f_arrdiv24_fs543_and1 = f_arrdiv24_fs543_not1 & f_arrdiv24_fs542_or0;
  assign f_arrdiv24_fs543_or0 = f_arrdiv24_fs543_and1 | f_arrdiv24_fs543_and0;
  assign f_arrdiv24_fs544_xor0 = f_arrdiv24_mux2to1498_xor0 ^ b[16];
  assign f_arrdiv24_fs544_not0 = ~f_arrdiv24_mux2to1498_xor0;
  assign f_arrdiv24_fs544_and0 = f_arrdiv24_fs544_not0 & b[16];
  assign f_arrdiv24_fs544_xor1 = f_arrdiv24_fs543_or0 ^ f_arrdiv24_fs544_xor0;
  assign f_arrdiv24_fs544_not1 = ~f_arrdiv24_fs544_xor0;
  assign f_arrdiv24_fs544_and1 = f_arrdiv24_fs544_not1 & f_arrdiv24_fs543_or0;
  assign f_arrdiv24_fs544_or0 = f_arrdiv24_fs544_and1 | f_arrdiv24_fs544_and0;
  assign f_arrdiv24_fs545_xor0 = f_arrdiv24_mux2to1499_xor0 ^ b[17];
  assign f_arrdiv24_fs545_not0 = ~f_arrdiv24_mux2to1499_xor0;
  assign f_arrdiv24_fs545_and0 = f_arrdiv24_fs545_not0 & b[17];
  assign f_arrdiv24_fs545_xor1 = f_arrdiv24_fs544_or0 ^ f_arrdiv24_fs545_xor0;
  assign f_arrdiv24_fs545_not1 = ~f_arrdiv24_fs545_xor0;
  assign f_arrdiv24_fs545_and1 = f_arrdiv24_fs545_not1 & f_arrdiv24_fs544_or0;
  assign f_arrdiv24_fs545_or0 = f_arrdiv24_fs545_and1 | f_arrdiv24_fs545_and0;
  assign f_arrdiv24_fs546_xor0 = f_arrdiv24_mux2to1500_xor0 ^ b[18];
  assign f_arrdiv24_fs546_not0 = ~f_arrdiv24_mux2to1500_xor0;
  assign f_arrdiv24_fs546_and0 = f_arrdiv24_fs546_not0 & b[18];
  assign f_arrdiv24_fs546_xor1 = f_arrdiv24_fs545_or0 ^ f_arrdiv24_fs546_xor0;
  assign f_arrdiv24_fs546_not1 = ~f_arrdiv24_fs546_xor0;
  assign f_arrdiv24_fs546_and1 = f_arrdiv24_fs546_not1 & f_arrdiv24_fs545_or0;
  assign f_arrdiv24_fs546_or0 = f_arrdiv24_fs546_and1 | f_arrdiv24_fs546_and0;
  assign f_arrdiv24_fs547_xor0 = f_arrdiv24_mux2to1501_xor0 ^ b[19];
  assign f_arrdiv24_fs547_not0 = ~f_arrdiv24_mux2to1501_xor0;
  assign f_arrdiv24_fs547_and0 = f_arrdiv24_fs547_not0 & b[19];
  assign f_arrdiv24_fs547_xor1 = f_arrdiv24_fs546_or0 ^ f_arrdiv24_fs547_xor0;
  assign f_arrdiv24_fs547_not1 = ~f_arrdiv24_fs547_xor0;
  assign f_arrdiv24_fs547_and1 = f_arrdiv24_fs547_not1 & f_arrdiv24_fs546_or0;
  assign f_arrdiv24_fs547_or0 = f_arrdiv24_fs547_and1 | f_arrdiv24_fs547_and0;
  assign f_arrdiv24_fs548_xor0 = f_arrdiv24_mux2to1502_xor0 ^ b[20];
  assign f_arrdiv24_fs548_not0 = ~f_arrdiv24_mux2to1502_xor0;
  assign f_arrdiv24_fs548_and0 = f_arrdiv24_fs548_not0 & b[20];
  assign f_arrdiv24_fs548_xor1 = f_arrdiv24_fs547_or0 ^ f_arrdiv24_fs548_xor0;
  assign f_arrdiv24_fs548_not1 = ~f_arrdiv24_fs548_xor0;
  assign f_arrdiv24_fs548_and1 = f_arrdiv24_fs548_not1 & f_arrdiv24_fs547_or0;
  assign f_arrdiv24_fs548_or0 = f_arrdiv24_fs548_and1 | f_arrdiv24_fs548_and0;
  assign f_arrdiv24_fs549_xor0 = f_arrdiv24_mux2to1503_xor0 ^ b[21];
  assign f_arrdiv24_fs549_not0 = ~f_arrdiv24_mux2to1503_xor0;
  assign f_arrdiv24_fs549_and0 = f_arrdiv24_fs549_not0 & b[21];
  assign f_arrdiv24_fs549_xor1 = f_arrdiv24_fs548_or0 ^ f_arrdiv24_fs549_xor0;
  assign f_arrdiv24_fs549_not1 = ~f_arrdiv24_fs549_xor0;
  assign f_arrdiv24_fs549_and1 = f_arrdiv24_fs549_not1 & f_arrdiv24_fs548_or0;
  assign f_arrdiv24_fs549_or0 = f_arrdiv24_fs549_and1 | f_arrdiv24_fs549_and0;
  assign f_arrdiv24_fs550_xor0 = f_arrdiv24_mux2to1504_xor0 ^ b[22];
  assign f_arrdiv24_fs550_not0 = ~f_arrdiv24_mux2to1504_xor0;
  assign f_arrdiv24_fs550_and0 = f_arrdiv24_fs550_not0 & b[22];
  assign f_arrdiv24_fs550_xor1 = f_arrdiv24_fs549_or0 ^ f_arrdiv24_fs550_xor0;
  assign f_arrdiv24_fs550_not1 = ~f_arrdiv24_fs550_xor0;
  assign f_arrdiv24_fs550_and1 = f_arrdiv24_fs550_not1 & f_arrdiv24_fs549_or0;
  assign f_arrdiv24_fs550_or0 = f_arrdiv24_fs550_and1 | f_arrdiv24_fs550_and0;
  assign f_arrdiv24_fs551_xor0 = f_arrdiv24_mux2to1505_xor0 ^ b[23];
  assign f_arrdiv24_fs551_not0 = ~f_arrdiv24_mux2to1505_xor0;
  assign f_arrdiv24_fs551_and0 = f_arrdiv24_fs551_not0 & b[23];
  assign f_arrdiv24_fs551_xor1 = f_arrdiv24_fs550_or0 ^ f_arrdiv24_fs551_xor0;
  assign f_arrdiv24_fs551_not1 = ~f_arrdiv24_fs551_xor0;
  assign f_arrdiv24_fs551_and1 = f_arrdiv24_fs551_not1 & f_arrdiv24_fs550_or0;
  assign f_arrdiv24_fs551_or0 = f_arrdiv24_fs551_and1 | f_arrdiv24_fs551_and0;
  assign f_arrdiv24_mux2to1506_and0 = a[1] & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1506_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1506_and1 = f_arrdiv24_fs528_xor0 & f_arrdiv24_mux2to1506_not0;
  assign f_arrdiv24_mux2to1506_xor0 = f_arrdiv24_mux2to1506_and0 ^ f_arrdiv24_mux2to1506_and1;
  assign f_arrdiv24_mux2to1507_and0 = f_arrdiv24_mux2to1483_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1507_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1507_and1 = f_arrdiv24_fs529_xor1 & f_arrdiv24_mux2to1507_not0;
  assign f_arrdiv24_mux2to1507_xor0 = f_arrdiv24_mux2to1507_and0 ^ f_arrdiv24_mux2to1507_and1;
  assign f_arrdiv24_mux2to1508_and0 = f_arrdiv24_mux2to1484_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1508_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1508_and1 = f_arrdiv24_fs530_xor1 & f_arrdiv24_mux2to1508_not0;
  assign f_arrdiv24_mux2to1508_xor0 = f_arrdiv24_mux2to1508_and0 ^ f_arrdiv24_mux2to1508_and1;
  assign f_arrdiv24_mux2to1509_and0 = f_arrdiv24_mux2to1485_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1509_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1509_and1 = f_arrdiv24_fs531_xor1 & f_arrdiv24_mux2to1509_not0;
  assign f_arrdiv24_mux2to1509_xor0 = f_arrdiv24_mux2to1509_and0 ^ f_arrdiv24_mux2to1509_and1;
  assign f_arrdiv24_mux2to1510_and0 = f_arrdiv24_mux2to1486_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1510_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1510_and1 = f_arrdiv24_fs532_xor1 & f_arrdiv24_mux2to1510_not0;
  assign f_arrdiv24_mux2to1510_xor0 = f_arrdiv24_mux2to1510_and0 ^ f_arrdiv24_mux2to1510_and1;
  assign f_arrdiv24_mux2to1511_and0 = f_arrdiv24_mux2to1487_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1511_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1511_and1 = f_arrdiv24_fs533_xor1 & f_arrdiv24_mux2to1511_not0;
  assign f_arrdiv24_mux2to1511_xor0 = f_arrdiv24_mux2to1511_and0 ^ f_arrdiv24_mux2to1511_and1;
  assign f_arrdiv24_mux2to1512_and0 = f_arrdiv24_mux2to1488_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1512_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1512_and1 = f_arrdiv24_fs534_xor1 & f_arrdiv24_mux2to1512_not0;
  assign f_arrdiv24_mux2to1512_xor0 = f_arrdiv24_mux2to1512_and0 ^ f_arrdiv24_mux2to1512_and1;
  assign f_arrdiv24_mux2to1513_and0 = f_arrdiv24_mux2to1489_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1513_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1513_and1 = f_arrdiv24_fs535_xor1 & f_arrdiv24_mux2to1513_not0;
  assign f_arrdiv24_mux2to1513_xor0 = f_arrdiv24_mux2to1513_and0 ^ f_arrdiv24_mux2to1513_and1;
  assign f_arrdiv24_mux2to1514_and0 = f_arrdiv24_mux2to1490_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1514_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1514_and1 = f_arrdiv24_fs536_xor1 & f_arrdiv24_mux2to1514_not0;
  assign f_arrdiv24_mux2to1514_xor0 = f_arrdiv24_mux2to1514_and0 ^ f_arrdiv24_mux2to1514_and1;
  assign f_arrdiv24_mux2to1515_and0 = f_arrdiv24_mux2to1491_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1515_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1515_and1 = f_arrdiv24_fs537_xor1 & f_arrdiv24_mux2to1515_not0;
  assign f_arrdiv24_mux2to1515_xor0 = f_arrdiv24_mux2to1515_and0 ^ f_arrdiv24_mux2to1515_and1;
  assign f_arrdiv24_mux2to1516_and0 = f_arrdiv24_mux2to1492_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1516_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1516_and1 = f_arrdiv24_fs538_xor1 & f_arrdiv24_mux2to1516_not0;
  assign f_arrdiv24_mux2to1516_xor0 = f_arrdiv24_mux2to1516_and0 ^ f_arrdiv24_mux2to1516_and1;
  assign f_arrdiv24_mux2to1517_and0 = f_arrdiv24_mux2to1493_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1517_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1517_and1 = f_arrdiv24_fs539_xor1 & f_arrdiv24_mux2to1517_not0;
  assign f_arrdiv24_mux2to1517_xor0 = f_arrdiv24_mux2to1517_and0 ^ f_arrdiv24_mux2to1517_and1;
  assign f_arrdiv24_mux2to1518_and0 = f_arrdiv24_mux2to1494_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1518_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1518_and1 = f_arrdiv24_fs540_xor1 & f_arrdiv24_mux2to1518_not0;
  assign f_arrdiv24_mux2to1518_xor0 = f_arrdiv24_mux2to1518_and0 ^ f_arrdiv24_mux2to1518_and1;
  assign f_arrdiv24_mux2to1519_and0 = f_arrdiv24_mux2to1495_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1519_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1519_and1 = f_arrdiv24_fs541_xor1 & f_arrdiv24_mux2to1519_not0;
  assign f_arrdiv24_mux2to1519_xor0 = f_arrdiv24_mux2to1519_and0 ^ f_arrdiv24_mux2to1519_and1;
  assign f_arrdiv24_mux2to1520_and0 = f_arrdiv24_mux2to1496_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1520_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1520_and1 = f_arrdiv24_fs542_xor1 & f_arrdiv24_mux2to1520_not0;
  assign f_arrdiv24_mux2to1520_xor0 = f_arrdiv24_mux2to1520_and0 ^ f_arrdiv24_mux2to1520_and1;
  assign f_arrdiv24_mux2to1521_and0 = f_arrdiv24_mux2to1497_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1521_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1521_and1 = f_arrdiv24_fs543_xor1 & f_arrdiv24_mux2to1521_not0;
  assign f_arrdiv24_mux2to1521_xor0 = f_arrdiv24_mux2to1521_and0 ^ f_arrdiv24_mux2to1521_and1;
  assign f_arrdiv24_mux2to1522_and0 = f_arrdiv24_mux2to1498_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1522_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1522_and1 = f_arrdiv24_fs544_xor1 & f_arrdiv24_mux2to1522_not0;
  assign f_arrdiv24_mux2to1522_xor0 = f_arrdiv24_mux2to1522_and0 ^ f_arrdiv24_mux2to1522_and1;
  assign f_arrdiv24_mux2to1523_and0 = f_arrdiv24_mux2to1499_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1523_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1523_and1 = f_arrdiv24_fs545_xor1 & f_arrdiv24_mux2to1523_not0;
  assign f_arrdiv24_mux2to1523_xor0 = f_arrdiv24_mux2to1523_and0 ^ f_arrdiv24_mux2to1523_and1;
  assign f_arrdiv24_mux2to1524_and0 = f_arrdiv24_mux2to1500_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1524_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1524_and1 = f_arrdiv24_fs546_xor1 & f_arrdiv24_mux2to1524_not0;
  assign f_arrdiv24_mux2to1524_xor0 = f_arrdiv24_mux2to1524_and0 ^ f_arrdiv24_mux2to1524_and1;
  assign f_arrdiv24_mux2to1525_and0 = f_arrdiv24_mux2to1501_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1525_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1525_and1 = f_arrdiv24_fs547_xor1 & f_arrdiv24_mux2to1525_not0;
  assign f_arrdiv24_mux2to1525_xor0 = f_arrdiv24_mux2to1525_and0 ^ f_arrdiv24_mux2to1525_and1;
  assign f_arrdiv24_mux2to1526_and0 = f_arrdiv24_mux2to1502_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1526_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1526_and1 = f_arrdiv24_fs548_xor1 & f_arrdiv24_mux2to1526_not0;
  assign f_arrdiv24_mux2to1526_xor0 = f_arrdiv24_mux2to1526_and0 ^ f_arrdiv24_mux2to1526_and1;
  assign f_arrdiv24_mux2to1527_and0 = f_arrdiv24_mux2to1503_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1527_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1527_and1 = f_arrdiv24_fs549_xor1 & f_arrdiv24_mux2to1527_not0;
  assign f_arrdiv24_mux2to1527_xor0 = f_arrdiv24_mux2to1527_and0 ^ f_arrdiv24_mux2to1527_and1;
  assign f_arrdiv24_mux2to1528_and0 = f_arrdiv24_mux2to1504_xor0 & f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1528_not0 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_mux2to1528_and1 = f_arrdiv24_fs550_xor1 & f_arrdiv24_mux2to1528_not0;
  assign f_arrdiv24_mux2to1528_xor0 = f_arrdiv24_mux2to1528_and0 ^ f_arrdiv24_mux2to1528_and1;
  assign f_arrdiv24_not22 = ~f_arrdiv24_fs551_or0;
  assign f_arrdiv24_fs552_xor0 = a[0] ^ b[0];
  assign f_arrdiv24_fs552_not0 = ~a[0];
  assign f_arrdiv24_fs552_and0 = f_arrdiv24_fs552_not0 & b[0];
  assign f_arrdiv24_fs552_not1 = ~f_arrdiv24_fs552_xor0;
  assign f_arrdiv24_fs553_xor0 = f_arrdiv24_mux2to1506_xor0 ^ b[1];
  assign f_arrdiv24_fs553_not0 = ~f_arrdiv24_mux2to1506_xor0;
  assign f_arrdiv24_fs553_and0 = f_arrdiv24_fs553_not0 & b[1];
  assign f_arrdiv24_fs553_xor1 = f_arrdiv24_fs552_and0 ^ f_arrdiv24_fs553_xor0;
  assign f_arrdiv24_fs553_not1 = ~f_arrdiv24_fs553_xor0;
  assign f_arrdiv24_fs553_and1 = f_arrdiv24_fs553_not1 & f_arrdiv24_fs552_and0;
  assign f_arrdiv24_fs553_or0 = f_arrdiv24_fs553_and1 | f_arrdiv24_fs553_and0;
  assign f_arrdiv24_fs554_xor0 = f_arrdiv24_mux2to1507_xor0 ^ b[2];
  assign f_arrdiv24_fs554_not0 = ~f_arrdiv24_mux2to1507_xor0;
  assign f_arrdiv24_fs554_and0 = f_arrdiv24_fs554_not0 & b[2];
  assign f_arrdiv24_fs554_xor1 = f_arrdiv24_fs553_or0 ^ f_arrdiv24_fs554_xor0;
  assign f_arrdiv24_fs554_not1 = ~f_arrdiv24_fs554_xor0;
  assign f_arrdiv24_fs554_and1 = f_arrdiv24_fs554_not1 & f_arrdiv24_fs553_or0;
  assign f_arrdiv24_fs554_or0 = f_arrdiv24_fs554_and1 | f_arrdiv24_fs554_and0;
  assign f_arrdiv24_fs555_xor0 = f_arrdiv24_mux2to1508_xor0 ^ b[3];
  assign f_arrdiv24_fs555_not0 = ~f_arrdiv24_mux2to1508_xor0;
  assign f_arrdiv24_fs555_and0 = f_arrdiv24_fs555_not0 & b[3];
  assign f_arrdiv24_fs555_xor1 = f_arrdiv24_fs554_or0 ^ f_arrdiv24_fs555_xor0;
  assign f_arrdiv24_fs555_not1 = ~f_arrdiv24_fs555_xor0;
  assign f_arrdiv24_fs555_and1 = f_arrdiv24_fs555_not1 & f_arrdiv24_fs554_or0;
  assign f_arrdiv24_fs555_or0 = f_arrdiv24_fs555_and1 | f_arrdiv24_fs555_and0;
  assign f_arrdiv24_fs556_xor0 = f_arrdiv24_mux2to1509_xor0 ^ b[4];
  assign f_arrdiv24_fs556_not0 = ~f_arrdiv24_mux2to1509_xor0;
  assign f_arrdiv24_fs556_and0 = f_arrdiv24_fs556_not0 & b[4];
  assign f_arrdiv24_fs556_xor1 = f_arrdiv24_fs555_or0 ^ f_arrdiv24_fs556_xor0;
  assign f_arrdiv24_fs556_not1 = ~f_arrdiv24_fs556_xor0;
  assign f_arrdiv24_fs556_and1 = f_arrdiv24_fs556_not1 & f_arrdiv24_fs555_or0;
  assign f_arrdiv24_fs556_or0 = f_arrdiv24_fs556_and1 | f_arrdiv24_fs556_and0;
  assign f_arrdiv24_fs557_xor0 = f_arrdiv24_mux2to1510_xor0 ^ b[5];
  assign f_arrdiv24_fs557_not0 = ~f_arrdiv24_mux2to1510_xor0;
  assign f_arrdiv24_fs557_and0 = f_arrdiv24_fs557_not0 & b[5];
  assign f_arrdiv24_fs557_xor1 = f_arrdiv24_fs556_or0 ^ f_arrdiv24_fs557_xor0;
  assign f_arrdiv24_fs557_not1 = ~f_arrdiv24_fs557_xor0;
  assign f_arrdiv24_fs557_and1 = f_arrdiv24_fs557_not1 & f_arrdiv24_fs556_or0;
  assign f_arrdiv24_fs557_or0 = f_arrdiv24_fs557_and1 | f_arrdiv24_fs557_and0;
  assign f_arrdiv24_fs558_xor0 = f_arrdiv24_mux2to1511_xor0 ^ b[6];
  assign f_arrdiv24_fs558_not0 = ~f_arrdiv24_mux2to1511_xor0;
  assign f_arrdiv24_fs558_and0 = f_arrdiv24_fs558_not0 & b[6];
  assign f_arrdiv24_fs558_xor1 = f_arrdiv24_fs557_or0 ^ f_arrdiv24_fs558_xor0;
  assign f_arrdiv24_fs558_not1 = ~f_arrdiv24_fs558_xor0;
  assign f_arrdiv24_fs558_and1 = f_arrdiv24_fs558_not1 & f_arrdiv24_fs557_or0;
  assign f_arrdiv24_fs558_or0 = f_arrdiv24_fs558_and1 | f_arrdiv24_fs558_and0;
  assign f_arrdiv24_fs559_xor0 = f_arrdiv24_mux2to1512_xor0 ^ b[7];
  assign f_arrdiv24_fs559_not0 = ~f_arrdiv24_mux2to1512_xor0;
  assign f_arrdiv24_fs559_and0 = f_arrdiv24_fs559_not0 & b[7];
  assign f_arrdiv24_fs559_xor1 = f_arrdiv24_fs558_or0 ^ f_arrdiv24_fs559_xor0;
  assign f_arrdiv24_fs559_not1 = ~f_arrdiv24_fs559_xor0;
  assign f_arrdiv24_fs559_and1 = f_arrdiv24_fs559_not1 & f_arrdiv24_fs558_or0;
  assign f_arrdiv24_fs559_or0 = f_arrdiv24_fs559_and1 | f_arrdiv24_fs559_and0;
  assign f_arrdiv24_fs560_xor0 = f_arrdiv24_mux2to1513_xor0 ^ b[8];
  assign f_arrdiv24_fs560_not0 = ~f_arrdiv24_mux2to1513_xor0;
  assign f_arrdiv24_fs560_and0 = f_arrdiv24_fs560_not0 & b[8];
  assign f_arrdiv24_fs560_xor1 = f_arrdiv24_fs559_or0 ^ f_arrdiv24_fs560_xor0;
  assign f_arrdiv24_fs560_not1 = ~f_arrdiv24_fs560_xor0;
  assign f_arrdiv24_fs560_and1 = f_arrdiv24_fs560_not1 & f_arrdiv24_fs559_or0;
  assign f_arrdiv24_fs560_or0 = f_arrdiv24_fs560_and1 | f_arrdiv24_fs560_and0;
  assign f_arrdiv24_fs561_xor0 = f_arrdiv24_mux2to1514_xor0 ^ b[9];
  assign f_arrdiv24_fs561_not0 = ~f_arrdiv24_mux2to1514_xor0;
  assign f_arrdiv24_fs561_and0 = f_arrdiv24_fs561_not0 & b[9];
  assign f_arrdiv24_fs561_xor1 = f_arrdiv24_fs560_or0 ^ f_arrdiv24_fs561_xor0;
  assign f_arrdiv24_fs561_not1 = ~f_arrdiv24_fs561_xor0;
  assign f_arrdiv24_fs561_and1 = f_arrdiv24_fs561_not1 & f_arrdiv24_fs560_or0;
  assign f_arrdiv24_fs561_or0 = f_arrdiv24_fs561_and1 | f_arrdiv24_fs561_and0;
  assign f_arrdiv24_fs562_xor0 = f_arrdiv24_mux2to1515_xor0 ^ b[10];
  assign f_arrdiv24_fs562_not0 = ~f_arrdiv24_mux2to1515_xor0;
  assign f_arrdiv24_fs562_and0 = f_arrdiv24_fs562_not0 & b[10];
  assign f_arrdiv24_fs562_xor1 = f_arrdiv24_fs561_or0 ^ f_arrdiv24_fs562_xor0;
  assign f_arrdiv24_fs562_not1 = ~f_arrdiv24_fs562_xor0;
  assign f_arrdiv24_fs562_and1 = f_arrdiv24_fs562_not1 & f_arrdiv24_fs561_or0;
  assign f_arrdiv24_fs562_or0 = f_arrdiv24_fs562_and1 | f_arrdiv24_fs562_and0;
  assign f_arrdiv24_fs563_xor0 = f_arrdiv24_mux2to1516_xor0 ^ b[11];
  assign f_arrdiv24_fs563_not0 = ~f_arrdiv24_mux2to1516_xor0;
  assign f_arrdiv24_fs563_and0 = f_arrdiv24_fs563_not0 & b[11];
  assign f_arrdiv24_fs563_xor1 = f_arrdiv24_fs562_or0 ^ f_arrdiv24_fs563_xor0;
  assign f_arrdiv24_fs563_not1 = ~f_arrdiv24_fs563_xor0;
  assign f_arrdiv24_fs563_and1 = f_arrdiv24_fs563_not1 & f_arrdiv24_fs562_or0;
  assign f_arrdiv24_fs563_or0 = f_arrdiv24_fs563_and1 | f_arrdiv24_fs563_and0;
  assign f_arrdiv24_fs564_xor0 = f_arrdiv24_mux2to1517_xor0 ^ b[12];
  assign f_arrdiv24_fs564_not0 = ~f_arrdiv24_mux2to1517_xor0;
  assign f_arrdiv24_fs564_and0 = f_arrdiv24_fs564_not0 & b[12];
  assign f_arrdiv24_fs564_xor1 = f_arrdiv24_fs563_or0 ^ f_arrdiv24_fs564_xor0;
  assign f_arrdiv24_fs564_not1 = ~f_arrdiv24_fs564_xor0;
  assign f_arrdiv24_fs564_and1 = f_arrdiv24_fs564_not1 & f_arrdiv24_fs563_or0;
  assign f_arrdiv24_fs564_or0 = f_arrdiv24_fs564_and1 | f_arrdiv24_fs564_and0;
  assign f_arrdiv24_fs565_xor0 = f_arrdiv24_mux2to1518_xor0 ^ b[13];
  assign f_arrdiv24_fs565_not0 = ~f_arrdiv24_mux2to1518_xor0;
  assign f_arrdiv24_fs565_and0 = f_arrdiv24_fs565_not0 & b[13];
  assign f_arrdiv24_fs565_xor1 = f_arrdiv24_fs564_or0 ^ f_arrdiv24_fs565_xor0;
  assign f_arrdiv24_fs565_not1 = ~f_arrdiv24_fs565_xor0;
  assign f_arrdiv24_fs565_and1 = f_arrdiv24_fs565_not1 & f_arrdiv24_fs564_or0;
  assign f_arrdiv24_fs565_or0 = f_arrdiv24_fs565_and1 | f_arrdiv24_fs565_and0;
  assign f_arrdiv24_fs566_xor0 = f_arrdiv24_mux2to1519_xor0 ^ b[14];
  assign f_arrdiv24_fs566_not0 = ~f_arrdiv24_mux2to1519_xor0;
  assign f_arrdiv24_fs566_and0 = f_arrdiv24_fs566_not0 & b[14];
  assign f_arrdiv24_fs566_xor1 = f_arrdiv24_fs565_or0 ^ f_arrdiv24_fs566_xor0;
  assign f_arrdiv24_fs566_not1 = ~f_arrdiv24_fs566_xor0;
  assign f_arrdiv24_fs566_and1 = f_arrdiv24_fs566_not1 & f_arrdiv24_fs565_or0;
  assign f_arrdiv24_fs566_or0 = f_arrdiv24_fs566_and1 | f_arrdiv24_fs566_and0;
  assign f_arrdiv24_fs567_xor0 = f_arrdiv24_mux2to1520_xor0 ^ b[15];
  assign f_arrdiv24_fs567_not0 = ~f_arrdiv24_mux2to1520_xor0;
  assign f_arrdiv24_fs567_and0 = f_arrdiv24_fs567_not0 & b[15];
  assign f_arrdiv24_fs567_xor1 = f_arrdiv24_fs566_or0 ^ f_arrdiv24_fs567_xor0;
  assign f_arrdiv24_fs567_not1 = ~f_arrdiv24_fs567_xor0;
  assign f_arrdiv24_fs567_and1 = f_arrdiv24_fs567_not1 & f_arrdiv24_fs566_or0;
  assign f_arrdiv24_fs567_or0 = f_arrdiv24_fs567_and1 | f_arrdiv24_fs567_and0;
  assign f_arrdiv24_fs568_xor0 = f_arrdiv24_mux2to1521_xor0 ^ b[16];
  assign f_arrdiv24_fs568_not0 = ~f_arrdiv24_mux2to1521_xor0;
  assign f_arrdiv24_fs568_and0 = f_arrdiv24_fs568_not0 & b[16];
  assign f_arrdiv24_fs568_xor1 = f_arrdiv24_fs567_or0 ^ f_arrdiv24_fs568_xor0;
  assign f_arrdiv24_fs568_not1 = ~f_arrdiv24_fs568_xor0;
  assign f_arrdiv24_fs568_and1 = f_arrdiv24_fs568_not1 & f_arrdiv24_fs567_or0;
  assign f_arrdiv24_fs568_or0 = f_arrdiv24_fs568_and1 | f_arrdiv24_fs568_and0;
  assign f_arrdiv24_fs569_xor0 = f_arrdiv24_mux2to1522_xor0 ^ b[17];
  assign f_arrdiv24_fs569_not0 = ~f_arrdiv24_mux2to1522_xor0;
  assign f_arrdiv24_fs569_and0 = f_arrdiv24_fs569_not0 & b[17];
  assign f_arrdiv24_fs569_xor1 = f_arrdiv24_fs568_or0 ^ f_arrdiv24_fs569_xor0;
  assign f_arrdiv24_fs569_not1 = ~f_arrdiv24_fs569_xor0;
  assign f_arrdiv24_fs569_and1 = f_arrdiv24_fs569_not1 & f_arrdiv24_fs568_or0;
  assign f_arrdiv24_fs569_or0 = f_arrdiv24_fs569_and1 | f_arrdiv24_fs569_and0;
  assign f_arrdiv24_fs570_xor0 = f_arrdiv24_mux2to1523_xor0 ^ b[18];
  assign f_arrdiv24_fs570_not0 = ~f_arrdiv24_mux2to1523_xor0;
  assign f_arrdiv24_fs570_and0 = f_arrdiv24_fs570_not0 & b[18];
  assign f_arrdiv24_fs570_xor1 = f_arrdiv24_fs569_or0 ^ f_arrdiv24_fs570_xor0;
  assign f_arrdiv24_fs570_not1 = ~f_arrdiv24_fs570_xor0;
  assign f_arrdiv24_fs570_and1 = f_arrdiv24_fs570_not1 & f_arrdiv24_fs569_or0;
  assign f_arrdiv24_fs570_or0 = f_arrdiv24_fs570_and1 | f_arrdiv24_fs570_and0;
  assign f_arrdiv24_fs571_xor0 = f_arrdiv24_mux2to1524_xor0 ^ b[19];
  assign f_arrdiv24_fs571_not0 = ~f_arrdiv24_mux2to1524_xor0;
  assign f_arrdiv24_fs571_and0 = f_arrdiv24_fs571_not0 & b[19];
  assign f_arrdiv24_fs571_xor1 = f_arrdiv24_fs570_or0 ^ f_arrdiv24_fs571_xor0;
  assign f_arrdiv24_fs571_not1 = ~f_arrdiv24_fs571_xor0;
  assign f_arrdiv24_fs571_and1 = f_arrdiv24_fs571_not1 & f_arrdiv24_fs570_or0;
  assign f_arrdiv24_fs571_or0 = f_arrdiv24_fs571_and1 | f_arrdiv24_fs571_and0;
  assign f_arrdiv24_fs572_xor0 = f_arrdiv24_mux2to1525_xor0 ^ b[20];
  assign f_arrdiv24_fs572_not0 = ~f_arrdiv24_mux2to1525_xor0;
  assign f_arrdiv24_fs572_and0 = f_arrdiv24_fs572_not0 & b[20];
  assign f_arrdiv24_fs572_xor1 = f_arrdiv24_fs571_or0 ^ f_arrdiv24_fs572_xor0;
  assign f_arrdiv24_fs572_not1 = ~f_arrdiv24_fs572_xor0;
  assign f_arrdiv24_fs572_and1 = f_arrdiv24_fs572_not1 & f_arrdiv24_fs571_or0;
  assign f_arrdiv24_fs572_or0 = f_arrdiv24_fs572_and1 | f_arrdiv24_fs572_and0;
  assign f_arrdiv24_fs573_xor0 = f_arrdiv24_mux2to1526_xor0 ^ b[21];
  assign f_arrdiv24_fs573_not0 = ~f_arrdiv24_mux2to1526_xor0;
  assign f_arrdiv24_fs573_and0 = f_arrdiv24_fs573_not0 & b[21];
  assign f_arrdiv24_fs573_xor1 = f_arrdiv24_fs572_or0 ^ f_arrdiv24_fs573_xor0;
  assign f_arrdiv24_fs573_not1 = ~f_arrdiv24_fs573_xor0;
  assign f_arrdiv24_fs573_and1 = f_arrdiv24_fs573_not1 & f_arrdiv24_fs572_or0;
  assign f_arrdiv24_fs573_or0 = f_arrdiv24_fs573_and1 | f_arrdiv24_fs573_and0;
  assign f_arrdiv24_fs574_xor0 = f_arrdiv24_mux2to1527_xor0 ^ b[22];
  assign f_arrdiv24_fs574_not0 = ~f_arrdiv24_mux2to1527_xor0;
  assign f_arrdiv24_fs574_and0 = f_arrdiv24_fs574_not0 & b[22];
  assign f_arrdiv24_fs574_xor1 = f_arrdiv24_fs573_or0 ^ f_arrdiv24_fs574_xor0;
  assign f_arrdiv24_fs574_not1 = ~f_arrdiv24_fs574_xor0;
  assign f_arrdiv24_fs574_and1 = f_arrdiv24_fs574_not1 & f_arrdiv24_fs573_or0;
  assign f_arrdiv24_fs574_or0 = f_arrdiv24_fs574_and1 | f_arrdiv24_fs574_and0;
  assign f_arrdiv24_fs575_xor0 = f_arrdiv24_mux2to1528_xor0 ^ b[23];
  assign f_arrdiv24_fs575_not0 = ~f_arrdiv24_mux2to1528_xor0;
  assign f_arrdiv24_fs575_and0 = f_arrdiv24_fs575_not0 & b[23];
  assign f_arrdiv24_fs575_xor1 = f_arrdiv24_fs574_or0 ^ f_arrdiv24_fs575_xor0;
  assign f_arrdiv24_fs575_not1 = ~f_arrdiv24_fs575_xor0;
  assign f_arrdiv24_fs575_and1 = f_arrdiv24_fs575_not1 & f_arrdiv24_fs574_or0;
  assign f_arrdiv24_fs575_or0 = f_arrdiv24_fs575_and1 | f_arrdiv24_fs575_and0;
  assign f_arrdiv24_not23 = ~f_arrdiv24_fs575_or0;

  assign f_arrdiv24_out[0] = f_arrdiv24_not23;
  assign f_arrdiv24_out[1] = f_arrdiv24_not22;
  assign f_arrdiv24_out[2] = f_arrdiv24_not21;
  assign f_arrdiv24_out[3] = f_arrdiv24_not20;
  assign f_arrdiv24_out[4] = f_arrdiv24_not19;
  assign f_arrdiv24_out[5] = f_arrdiv24_not18;
  assign f_arrdiv24_out[6] = f_arrdiv24_not17;
  assign f_arrdiv24_out[7] = f_arrdiv24_not16;
  assign f_arrdiv24_out[8] = f_arrdiv24_not15;
  assign f_arrdiv24_out[9] = f_arrdiv24_not14;
  assign f_arrdiv24_out[10] = f_arrdiv24_not13;
  assign f_arrdiv24_out[11] = f_arrdiv24_not12;
  assign f_arrdiv24_out[12] = f_arrdiv24_not11;
  assign f_arrdiv24_out[13] = f_arrdiv24_not10;
  assign f_arrdiv24_out[14] = f_arrdiv24_not9;
  assign f_arrdiv24_out[15] = f_arrdiv24_not8;
  assign f_arrdiv24_out[16] = f_arrdiv24_not7;
  assign f_arrdiv24_out[17] = f_arrdiv24_not6;
  assign f_arrdiv24_out[18] = f_arrdiv24_not5;
  assign f_arrdiv24_out[19] = f_arrdiv24_not4;
  assign f_arrdiv24_out[20] = f_arrdiv24_not3;
  assign f_arrdiv24_out[21] = f_arrdiv24_not2;
  assign f_arrdiv24_out[22] = f_arrdiv24_not1;
  assign f_arrdiv24_out[23] = f_arrdiv24_not0;
endmodule