module f_u_csabam8_cla_h0_v6(input [7:0] a, input [7:0] b, output [15:0] f_u_csabam8_cla_h0_v6_out);
  wire f_u_csabam8_cla_h0_v6_and6_0;
  wire f_u_csabam8_cla_h0_v6_and7_0;
  wire f_u_csabam8_cla_h0_v6_and5_1;
  wire f_u_csabam8_cla_h0_v6_ha5_1_xor0;
  wire f_u_csabam8_cla_h0_v6_ha5_1_and0;
  wire f_u_csabam8_cla_h0_v6_and6_1;
  wire f_u_csabam8_cla_h0_v6_ha6_1_xor0;
  wire f_u_csabam8_cla_h0_v6_ha6_1_and0;
  wire f_u_csabam8_cla_h0_v6_and7_1;
  wire f_u_csabam8_cla_h0_v6_and4_2;
  wire f_u_csabam8_cla_h0_v6_ha4_2_xor0;
  wire f_u_csabam8_cla_h0_v6_ha4_2_and0;
  wire f_u_csabam8_cla_h0_v6_and5_2;
  wire f_u_csabam8_cla_h0_v6_fa5_2_xor0;
  wire f_u_csabam8_cla_h0_v6_fa5_2_and0;
  wire f_u_csabam8_cla_h0_v6_fa5_2_xor1;
  wire f_u_csabam8_cla_h0_v6_fa5_2_and1;
  wire f_u_csabam8_cla_h0_v6_fa5_2_or0;
  wire f_u_csabam8_cla_h0_v6_and6_2;
  wire f_u_csabam8_cla_h0_v6_fa6_2_xor0;
  wire f_u_csabam8_cla_h0_v6_fa6_2_and0;
  wire f_u_csabam8_cla_h0_v6_fa6_2_xor1;
  wire f_u_csabam8_cla_h0_v6_fa6_2_and1;
  wire f_u_csabam8_cla_h0_v6_fa6_2_or0;
  wire f_u_csabam8_cla_h0_v6_and7_2;
  wire f_u_csabam8_cla_h0_v6_and3_3;
  wire f_u_csabam8_cla_h0_v6_ha3_3_xor0;
  wire f_u_csabam8_cla_h0_v6_ha3_3_and0;
  wire f_u_csabam8_cla_h0_v6_and4_3;
  wire f_u_csabam8_cla_h0_v6_fa4_3_xor0;
  wire f_u_csabam8_cla_h0_v6_fa4_3_and0;
  wire f_u_csabam8_cla_h0_v6_fa4_3_xor1;
  wire f_u_csabam8_cla_h0_v6_fa4_3_and1;
  wire f_u_csabam8_cla_h0_v6_fa4_3_or0;
  wire f_u_csabam8_cla_h0_v6_and5_3;
  wire f_u_csabam8_cla_h0_v6_fa5_3_xor0;
  wire f_u_csabam8_cla_h0_v6_fa5_3_and0;
  wire f_u_csabam8_cla_h0_v6_fa5_3_xor1;
  wire f_u_csabam8_cla_h0_v6_fa5_3_and1;
  wire f_u_csabam8_cla_h0_v6_fa5_3_or0;
  wire f_u_csabam8_cla_h0_v6_and6_3;
  wire f_u_csabam8_cla_h0_v6_fa6_3_xor0;
  wire f_u_csabam8_cla_h0_v6_fa6_3_and0;
  wire f_u_csabam8_cla_h0_v6_fa6_3_xor1;
  wire f_u_csabam8_cla_h0_v6_fa6_3_and1;
  wire f_u_csabam8_cla_h0_v6_fa6_3_or0;
  wire f_u_csabam8_cla_h0_v6_and7_3;
  wire f_u_csabam8_cla_h0_v6_and2_4;
  wire f_u_csabam8_cla_h0_v6_ha2_4_xor0;
  wire f_u_csabam8_cla_h0_v6_ha2_4_and0;
  wire f_u_csabam8_cla_h0_v6_and3_4;
  wire f_u_csabam8_cla_h0_v6_fa3_4_xor0;
  wire f_u_csabam8_cla_h0_v6_fa3_4_and0;
  wire f_u_csabam8_cla_h0_v6_fa3_4_xor1;
  wire f_u_csabam8_cla_h0_v6_fa3_4_and1;
  wire f_u_csabam8_cla_h0_v6_fa3_4_or0;
  wire f_u_csabam8_cla_h0_v6_and4_4;
  wire f_u_csabam8_cla_h0_v6_fa4_4_xor0;
  wire f_u_csabam8_cla_h0_v6_fa4_4_and0;
  wire f_u_csabam8_cla_h0_v6_fa4_4_xor1;
  wire f_u_csabam8_cla_h0_v6_fa4_4_and1;
  wire f_u_csabam8_cla_h0_v6_fa4_4_or0;
  wire f_u_csabam8_cla_h0_v6_and5_4;
  wire f_u_csabam8_cla_h0_v6_fa5_4_xor0;
  wire f_u_csabam8_cla_h0_v6_fa5_4_and0;
  wire f_u_csabam8_cla_h0_v6_fa5_4_xor1;
  wire f_u_csabam8_cla_h0_v6_fa5_4_and1;
  wire f_u_csabam8_cla_h0_v6_fa5_4_or0;
  wire f_u_csabam8_cla_h0_v6_and6_4;
  wire f_u_csabam8_cla_h0_v6_fa6_4_xor0;
  wire f_u_csabam8_cla_h0_v6_fa6_4_and0;
  wire f_u_csabam8_cla_h0_v6_fa6_4_xor1;
  wire f_u_csabam8_cla_h0_v6_fa6_4_and1;
  wire f_u_csabam8_cla_h0_v6_fa6_4_or0;
  wire f_u_csabam8_cla_h0_v6_and7_4;
  wire f_u_csabam8_cla_h0_v6_and1_5;
  wire f_u_csabam8_cla_h0_v6_ha1_5_xor0;
  wire f_u_csabam8_cla_h0_v6_ha1_5_and0;
  wire f_u_csabam8_cla_h0_v6_and2_5;
  wire f_u_csabam8_cla_h0_v6_fa2_5_xor0;
  wire f_u_csabam8_cla_h0_v6_fa2_5_and0;
  wire f_u_csabam8_cla_h0_v6_fa2_5_xor1;
  wire f_u_csabam8_cla_h0_v6_fa2_5_and1;
  wire f_u_csabam8_cla_h0_v6_fa2_5_or0;
  wire f_u_csabam8_cla_h0_v6_and3_5;
  wire f_u_csabam8_cla_h0_v6_fa3_5_xor0;
  wire f_u_csabam8_cla_h0_v6_fa3_5_and0;
  wire f_u_csabam8_cla_h0_v6_fa3_5_xor1;
  wire f_u_csabam8_cla_h0_v6_fa3_5_and1;
  wire f_u_csabam8_cla_h0_v6_fa3_5_or0;
  wire f_u_csabam8_cla_h0_v6_and4_5;
  wire f_u_csabam8_cla_h0_v6_fa4_5_xor0;
  wire f_u_csabam8_cla_h0_v6_fa4_5_and0;
  wire f_u_csabam8_cla_h0_v6_fa4_5_xor1;
  wire f_u_csabam8_cla_h0_v6_fa4_5_and1;
  wire f_u_csabam8_cla_h0_v6_fa4_5_or0;
  wire f_u_csabam8_cla_h0_v6_and5_5;
  wire f_u_csabam8_cla_h0_v6_fa5_5_xor0;
  wire f_u_csabam8_cla_h0_v6_fa5_5_and0;
  wire f_u_csabam8_cla_h0_v6_fa5_5_xor1;
  wire f_u_csabam8_cla_h0_v6_fa5_5_and1;
  wire f_u_csabam8_cla_h0_v6_fa5_5_or0;
  wire f_u_csabam8_cla_h0_v6_and6_5;
  wire f_u_csabam8_cla_h0_v6_fa6_5_xor0;
  wire f_u_csabam8_cla_h0_v6_fa6_5_and0;
  wire f_u_csabam8_cla_h0_v6_fa6_5_xor1;
  wire f_u_csabam8_cla_h0_v6_fa6_5_and1;
  wire f_u_csabam8_cla_h0_v6_fa6_5_or0;
  wire f_u_csabam8_cla_h0_v6_and7_5;
  wire f_u_csabam8_cla_h0_v6_and0_6;
  wire f_u_csabam8_cla_h0_v6_ha0_6_xor0;
  wire f_u_csabam8_cla_h0_v6_ha0_6_and0;
  wire f_u_csabam8_cla_h0_v6_and1_6;
  wire f_u_csabam8_cla_h0_v6_fa1_6_xor0;
  wire f_u_csabam8_cla_h0_v6_fa1_6_and0;
  wire f_u_csabam8_cla_h0_v6_fa1_6_xor1;
  wire f_u_csabam8_cla_h0_v6_fa1_6_and1;
  wire f_u_csabam8_cla_h0_v6_fa1_6_or0;
  wire f_u_csabam8_cla_h0_v6_and2_6;
  wire f_u_csabam8_cla_h0_v6_fa2_6_xor0;
  wire f_u_csabam8_cla_h0_v6_fa2_6_and0;
  wire f_u_csabam8_cla_h0_v6_fa2_6_xor1;
  wire f_u_csabam8_cla_h0_v6_fa2_6_and1;
  wire f_u_csabam8_cla_h0_v6_fa2_6_or0;
  wire f_u_csabam8_cla_h0_v6_and3_6;
  wire f_u_csabam8_cla_h0_v6_fa3_6_xor0;
  wire f_u_csabam8_cla_h0_v6_fa3_6_and0;
  wire f_u_csabam8_cla_h0_v6_fa3_6_xor1;
  wire f_u_csabam8_cla_h0_v6_fa3_6_and1;
  wire f_u_csabam8_cla_h0_v6_fa3_6_or0;
  wire f_u_csabam8_cla_h0_v6_and4_6;
  wire f_u_csabam8_cla_h0_v6_fa4_6_xor0;
  wire f_u_csabam8_cla_h0_v6_fa4_6_and0;
  wire f_u_csabam8_cla_h0_v6_fa4_6_xor1;
  wire f_u_csabam8_cla_h0_v6_fa4_6_and1;
  wire f_u_csabam8_cla_h0_v6_fa4_6_or0;
  wire f_u_csabam8_cla_h0_v6_and5_6;
  wire f_u_csabam8_cla_h0_v6_fa5_6_xor0;
  wire f_u_csabam8_cla_h0_v6_fa5_6_and0;
  wire f_u_csabam8_cla_h0_v6_fa5_6_xor1;
  wire f_u_csabam8_cla_h0_v6_fa5_6_and1;
  wire f_u_csabam8_cla_h0_v6_fa5_6_or0;
  wire f_u_csabam8_cla_h0_v6_and6_6;
  wire f_u_csabam8_cla_h0_v6_fa6_6_xor0;
  wire f_u_csabam8_cla_h0_v6_fa6_6_and0;
  wire f_u_csabam8_cla_h0_v6_fa6_6_xor1;
  wire f_u_csabam8_cla_h0_v6_fa6_6_and1;
  wire f_u_csabam8_cla_h0_v6_fa6_6_or0;
  wire f_u_csabam8_cla_h0_v6_and7_6;
  wire f_u_csabam8_cla_h0_v6_and0_7;
  wire f_u_csabam8_cla_h0_v6_fa0_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa0_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa0_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa0_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa0_7_or0;
  wire f_u_csabam8_cla_h0_v6_and1_7;
  wire f_u_csabam8_cla_h0_v6_fa1_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa1_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa1_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa1_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa1_7_or0;
  wire f_u_csabam8_cla_h0_v6_and2_7;
  wire f_u_csabam8_cla_h0_v6_fa2_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa2_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa2_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa2_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa2_7_or0;
  wire f_u_csabam8_cla_h0_v6_and3_7;
  wire f_u_csabam8_cla_h0_v6_fa3_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa3_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa3_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa3_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa3_7_or0;
  wire f_u_csabam8_cla_h0_v6_and4_7;
  wire f_u_csabam8_cla_h0_v6_fa4_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa4_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa4_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa4_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa4_7_or0;
  wire f_u_csabam8_cla_h0_v6_and5_7;
  wire f_u_csabam8_cla_h0_v6_fa5_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa5_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa5_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa5_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa5_7_or0;
  wire f_u_csabam8_cla_h0_v6_and6_7;
  wire f_u_csabam8_cla_h0_v6_fa6_7_xor0;
  wire f_u_csabam8_cla_h0_v6_fa6_7_and0;
  wire f_u_csabam8_cla_h0_v6_fa6_7_xor1;
  wire f_u_csabam8_cla_h0_v6_fa6_7_and1;
  wire f_u_csabam8_cla_h0_v6_fa6_7_or0;
  wire f_u_csabam8_cla_h0_v6_and7_7;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_xor1;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_xor2;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and1;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and2;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and3;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and4;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or1;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or2;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_xor3;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and5;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and6;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and7;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and8;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and9;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and10;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and11;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or3;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or4;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or5;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_xor4;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and12;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or6;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_xor5;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and13;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and14;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and15;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or7;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or8;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_and0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_xor0;
  wire f_u_csabam8_cla_h0_v6_u_cla8_xor6;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and16;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and17;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and18;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and19;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and20;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and21;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or9;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or10;
  wire f_u_csabam8_cla_h0_v6_u_cla8_or11;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and22;
  wire f_u_csabam8_cla_h0_v6_u_cla8_and23;

  assign f_u_csabam8_cla_h0_v6_and6_0 = a[6] & b[0];
  assign f_u_csabam8_cla_h0_v6_and7_0 = a[7] & b[0];
  assign f_u_csabam8_cla_h0_v6_and5_1 = a[5] & b[1];
  assign f_u_csabam8_cla_h0_v6_ha5_1_xor0 = f_u_csabam8_cla_h0_v6_and5_1 ^ f_u_csabam8_cla_h0_v6_and6_0;
  assign f_u_csabam8_cla_h0_v6_ha5_1_and0 = f_u_csabam8_cla_h0_v6_and5_1 & f_u_csabam8_cla_h0_v6_and6_0;
  assign f_u_csabam8_cla_h0_v6_and6_1 = a[6] & b[1];
  assign f_u_csabam8_cla_h0_v6_ha6_1_xor0 = f_u_csabam8_cla_h0_v6_and6_1 ^ f_u_csabam8_cla_h0_v6_and7_0;
  assign f_u_csabam8_cla_h0_v6_ha6_1_and0 = f_u_csabam8_cla_h0_v6_and6_1 & f_u_csabam8_cla_h0_v6_and7_0;
  assign f_u_csabam8_cla_h0_v6_and7_1 = a[7] & b[1];
  assign f_u_csabam8_cla_h0_v6_and4_2 = a[4] & b[2];
  assign f_u_csabam8_cla_h0_v6_ha4_2_xor0 = f_u_csabam8_cla_h0_v6_and4_2 ^ f_u_csabam8_cla_h0_v6_ha5_1_xor0;
  assign f_u_csabam8_cla_h0_v6_ha4_2_and0 = f_u_csabam8_cla_h0_v6_and4_2 & f_u_csabam8_cla_h0_v6_ha5_1_xor0;
  assign f_u_csabam8_cla_h0_v6_and5_2 = a[5] & b[2];
  assign f_u_csabam8_cla_h0_v6_fa5_2_xor0 = f_u_csabam8_cla_h0_v6_and5_2 ^ f_u_csabam8_cla_h0_v6_ha6_1_xor0;
  assign f_u_csabam8_cla_h0_v6_fa5_2_and0 = f_u_csabam8_cla_h0_v6_and5_2 & f_u_csabam8_cla_h0_v6_ha6_1_xor0;
  assign f_u_csabam8_cla_h0_v6_fa5_2_xor1 = f_u_csabam8_cla_h0_v6_fa5_2_xor0 ^ f_u_csabam8_cla_h0_v6_ha5_1_and0;
  assign f_u_csabam8_cla_h0_v6_fa5_2_and1 = f_u_csabam8_cla_h0_v6_fa5_2_xor0 & f_u_csabam8_cla_h0_v6_ha5_1_and0;
  assign f_u_csabam8_cla_h0_v6_fa5_2_or0 = f_u_csabam8_cla_h0_v6_fa5_2_and0 | f_u_csabam8_cla_h0_v6_fa5_2_and1;
  assign f_u_csabam8_cla_h0_v6_and6_2 = a[6] & b[2];
  assign f_u_csabam8_cla_h0_v6_fa6_2_xor0 = f_u_csabam8_cla_h0_v6_and6_2 ^ f_u_csabam8_cla_h0_v6_and7_1;
  assign f_u_csabam8_cla_h0_v6_fa6_2_and0 = f_u_csabam8_cla_h0_v6_and6_2 & f_u_csabam8_cla_h0_v6_and7_1;
  assign f_u_csabam8_cla_h0_v6_fa6_2_xor1 = f_u_csabam8_cla_h0_v6_fa6_2_xor0 ^ f_u_csabam8_cla_h0_v6_ha6_1_and0;
  assign f_u_csabam8_cla_h0_v6_fa6_2_and1 = f_u_csabam8_cla_h0_v6_fa6_2_xor0 & f_u_csabam8_cla_h0_v6_ha6_1_and0;
  assign f_u_csabam8_cla_h0_v6_fa6_2_or0 = f_u_csabam8_cla_h0_v6_fa6_2_and0 | f_u_csabam8_cla_h0_v6_fa6_2_and1;
  assign f_u_csabam8_cla_h0_v6_and7_2 = a[7] & b[2];
  assign f_u_csabam8_cla_h0_v6_and3_3 = a[3] & b[3];
  assign f_u_csabam8_cla_h0_v6_ha3_3_xor0 = f_u_csabam8_cla_h0_v6_and3_3 ^ f_u_csabam8_cla_h0_v6_ha4_2_xor0;
  assign f_u_csabam8_cla_h0_v6_ha3_3_and0 = f_u_csabam8_cla_h0_v6_and3_3 & f_u_csabam8_cla_h0_v6_ha4_2_xor0;
  assign f_u_csabam8_cla_h0_v6_and4_3 = a[4] & b[3];
  assign f_u_csabam8_cla_h0_v6_fa4_3_xor0 = f_u_csabam8_cla_h0_v6_and4_3 ^ f_u_csabam8_cla_h0_v6_fa5_2_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_3_and0 = f_u_csabam8_cla_h0_v6_and4_3 & f_u_csabam8_cla_h0_v6_fa5_2_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_3_xor1 = f_u_csabam8_cla_h0_v6_fa4_3_xor0 ^ f_u_csabam8_cla_h0_v6_ha4_2_and0;
  assign f_u_csabam8_cla_h0_v6_fa4_3_and1 = f_u_csabam8_cla_h0_v6_fa4_3_xor0 & f_u_csabam8_cla_h0_v6_ha4_2_and0;
  assign f_u_csabam8_cla_h0_v6_fa4_3_or0 = f_u_csabam8_cla_h0_v6_fa4_3_and0 | f_u_csabam8_cla_h0_v6_fa4_3_and1;
  assign f_u_csabam8_cla_h0_v6_and5_3 = a[5] & b[3];
  assign f_u_csabam8_cla_h0_v6_fa5_3_xor0 = f_u_csabam8_cla_h0_v6_and5_3 ^ f_u_csabam8_cla_h0_v6_fa6_2_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_3_and0 = f_u_csabam8_cla_h0_v6_and5_3 & f_u_csabam8_cla_h0_v6_fa6_2_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_3_xor1 = f_u_csabam8_cla_h0_v6_fa5_3_xor0 ^ f_u_csabam8_cla_h0_v6_fa5_2_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_3_and1 = f_u_csabam8_cla_h0_v6_fa5_3_xor0 & f_u_csabam8_cla_h0_v6_fa5_2_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_3_or0 = f_u_csabam8_cla_h0_v6_fa5_3_and0 | f_u_csabam8_cla_h0_v6_fa5_3_and1;
  assign f_u_csabam8_cla_h0_v6_and6_3 = a[6] & b[3];
  assign f_u_csabam8_cla_h0_v6_fa6_3_xor0 = f_u_csabam8_cla_h0_v6_and6_3 ^ f_u_csabam8_cla_h0_v6_and7_2;
  assign f_u_csabam8_cla_h0_v6_fa6_3_and0 = f_u_csabam8_cla_h0_v6_and6_3 & f_u_csabam8_cla_h0_v6_and7_2;
  assign f_u_csabam8_cla_h0_v6_fa6_3_xor1 = f_u_csabam8_cla_h0_v6_fa6_3_xor0 ^ f_u_csabam8_cla_h0_v6_fa6_2_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_3_and1 = f_u_csabam8_cla_h0_v6_fa6_3_xor0 & f_u_csabam8_cla_h0_v6_fa6_2_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_3_or0 = f_u_csabam8_cla_h0_v6_fa6_3_and0 | f_u_csabam8_cla_h0_v6_fa6_3_and1;
  assign f_u_csabam8_cla_h0_v6_and7_3 = a[7] & b[3];
  assign f_u_csabam8_cla_h0_v6_and2_4 = a[2] & b[4];
  assign f_u_csabam8_cla_h0_v6_ha2_4_xor0 = f_u_csabam8_cla_h0_v6_and2_4 ^ f_u_csabam8_cla_h0_v6_ha3_3_xor0;
  assign f_u_csabam8_cla_h0_v6_ha2_4_and0 = f_u_csabam8_cla_h0_v6_and2_4 & f_u_csabam8_cla_h0_v6_ha3_3_xor0;
  assign f_u_csabam8_cla_h0_v6_and3_4 = a[3] & b[4];
  assign f_u_csabam8_cla_h0_v6_fa3_4_xor0 = f_u_csabam8_cla_h0_v6_and3_4 ^ f_u_csabam8_cla_h0_v6_fa4_3_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_4_and0 = f_u_csabam8_cla_h0_v6_and3_4 & f_u_csabam8_cla_h0_v6_fa4_3_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_4_xor1 = f_u_csabam8_cla_h0_v6_fa3_4_xor0 ^ f_u_csabam8_cla_h0_v6_ha3_3_and0;
  assign f_u_csabam8_cla_h0_v6_fa3_4_and1 = f_u_csabam8_cla_h0_v6_fa3_4_xor0 & f_u_csabam8_cla_h0_v6_ha3_3_and0;
  assign f_u_csabam8_cla_h0_v6_fa3_4_or0 = f_u_csabam8_cla_h0_v6_fa3_4_and0 | f_u_csabam8_cla_h0_v6_fa3_4_and1;
  assign f_u_csabam8_cla_h0_v6_and4_4 = a[4] & b[4];
  assign f_u_csabam8_cla_h0_v6_fa4_4_xor0 = f_u_csabam8_cla_h0_v6_and4_4 ^ f_u_csabam8_cla_h0_v6_fa5_3_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_4_and0 = f_u_csabam8_cla_h0_v6_and4_4 & f_u_csabam8_cla_h0_v6_fa5_3_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_4_xor1 = f_u_csabam8_cla_h0_v6_fa4_4_xor0 ^ f_u_csabam8_cla_h0_v6_fa4_3_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_4_and1 = f_u_csabam8_cla_h0_v6_fa4_4_xor0 & f_u_csabam8_cla_h0_v6_fa4_3_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_4_or0 = f_u_csabam8_cla_h0_v6_fa4_4_and0 | f_u_csabam8_cla_h0_v6_fa4_4_and1;
  assign f_u_csabam8_cla_h0_v6_and5_4 = a[5] & b[4];
  assign f_u_csabam8_cla_h0_v6_fa5_4_xor0 = f_u_csabam8_cla_h0_v6_and5_4 ^ f_u_csabam8_cla_h0_v6_fa6_3_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_4_and0 = f_u_csabam8_cla_h0_v6_and5_4 & f_u_csabam8_cla_h0_v6_fa6_3_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_4_xor1 = f_u_csabam8_cla_h0_v6_fa5_4_xor0 ^ f_u_csabam8_cla_h0_v6_fa5_3_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_4_and1 = f_u_csabam8_cla_h0_v6_fa5_4_xor0 & f_u_csabam8_cla_h0_v6_fa5_3_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_4_or0 = f_u_csabam8_cla_h0_v6_fa5_4_and0 | f_u_csabam8_cla_h0_v6_fa5_4_and1;
  assign f_u_csabam8_cla_h0_v6_and6_4 = a[6] & b[4];
  assign f_u_csabam8_cla_h0_v6_fa6_4_xor0 = f_u_csabam8_cla_h0_v6_and6_4 ^ f_u_csabam8_cla_h0_v6_and7_3;
  assign f_u_csabam8_cla_h0_v6_fa6_4_and0 = f_u_csabam8_cla_h0_v6_and6_4 & f_u_csabam8_cla_h0_v6_and7_3;
  assign f_u_csabam8_cla_h0_v6_fa6_4_xor1 = f_u_csabam8_cla_h0_v6_fa6_4_xor0 ^ f_u_csabam8_cla_h0_v6_fa6_3_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_4_and1 = f_u_csabam8_cla_h0_v6_fa6_4_xor0 & f_u_csabam8_cla_h0_v6_fa6_3_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_4_or0 = f_u_csabam8_cla_h0_v6_fa6_4_and0 | f_u_csabam8_cla_h0_v6_fa6_4_and1;
  assign f_u_csabam8_cla_h0_v6_and7_4 = a[7] & b[4];
  assign f_u_csabam8_cla_h0_v6_and1_5 = a[1] & b[5];
  assign f_u_csabam8_cla_h0_v6_ha1_5_xor0 = f_u_csabam8_cla_h0_v6_and1_5 ^ f_u_csabam8_cla_h0_v6_ha2_4_xor0;
  assign f_u_csabam8_cla_h0_v6_ha1_5_and0 = f_u_csabam8_cla_h0_v6_and1_5 & f_u_csabam8_cla_h0_v6_ha2_4_xor0;
  assign f_u_csabam8_cla_h0_v6_and2_5 = a[2] & b[5];
  assign f_u_csabam8_cla_h0_v6_fa2_5_xor0 = f_u_csabam8_cla_h0_v6_and2_5 ^ f_u_csabam8_cla_h0_v6_fa3_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa2_5_and0 = f_u_csabam8_cla_h0_v6_and2_5 & f_u_csabam8_cla_h0_v6_fa3_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa2_5_xor1 = f_u_csabam8_cla_h0_v6_fa2_5_xor0 ^ f_u_csabam8_cla_h0_v6_ha2_4_and0;
  assign f_u_csabam8_cla_h0_v6_fa2_5_and1 = f_u_csabam8_cla_h0_v6_fa2_5_xor0 & f_u_csabam8_cla_h0_v6_ha2_4_and0;
  assign f_u_csabam8_cla_h0_v6_fa2_5_or0 = f_u_csabam8_cla_h0_v6_fa2_5_and0 | f_u_csabam8_cla_h0_v6_fa2_5_and1;
  assign f_u_csabam8_cla_h0_v6_and3_5 = a[3] & b[5];
  assign f_u_csabam8_cla_h0_v6_fa3_5_xor0 = f_u_csabam8_cla_h0_v6_and3_5 ^ f_u_csabam8_cla_h0_v6_fa4_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_5_and0 = f_u_csabam8_cla_h0_v6_and3_5 & f_u_csabam8_cla_h0_v6_fa4_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_5_xor1 = f_u_csabam8_cla_h0_v6_fa3_5_xor0 ^ f_u_csabam8_cla_h0_v6_fa3_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa3_5_and1 = f_u_csabam8_cla_h0_v6_fa3_5_xor0 & f_u_csabam8_cla_h0_v6_fa3_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa3_5_or0 = f_u_csabam8_cla_h0_v6_fa3_5_and0 | f_u_csabam8_cla_h0_v6_fa3_5_and1;
  assign f_u_csabam8_cla_h0_v6_and4_5 = a[4] & b[5];
  assign f_u_csabam8_cla_h0_v6_fa4_5_xor0 = f_u_csabam8_cla_h0_v6_and4_5 ^ f_u_csabam8_cla_h0_v6_fa5_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_5_and0 = f_u_csabam8_cla_h0_v6_and4_5 & f_u_csabam8_cla_h0_v6_fa5_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_5_xor1 = f_u_csabam8_cla_h0_v6_fa4_5_xor0 ^ f_u_csabam8_cla_h0_v6_fa4_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_5_and1 = f_u_csabam8_cla_h0_v6_fa4_5_xor0 & f_u_csabam8_cla_h0_v6_fa4_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_5_or0 = f_u_csabam8_cla_h0_v6_fa4_5_and0 | f_u_csabam8_cla_h0_v6_fa4_5_and1;
  assign f_u_csabam8_cla_h0_v6_and5_5 = a[5] & b[5];
  assign f_u_csabam8_cla_h0_v6_fa5_5_xor0 = f_u_csabam8_cla_h0_v6_and5_5 ^ f_u_csabam8_cla_h0_v6_fa6_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_5_and0 = f_u_csabam8_cla_h0_v6_and5_5 & f_u_csabam8_cla_h0_v6_fa6_4_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_5_xor1 = f_u_csabam8_cla_h0_v6_fa5_5_xor0 ^ f_u_csabam8_cla_h0_v6_fa5_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_5_and1 = f_u_csabam8_cla_h0_v6_fa5_5_xor0 & f_u_csabam8_cla_h0_v6_fa5_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_5_or0 = f_u_csabam8_cla_h0_v6_fa5_5_and0 | f_u_csabam8_cla_h0_v6_fa5_5_and1;
  assign f_u_csabam8_cla_h0_v6_and6_5 = a[6] & b[5];
  assign f_u_csabam8_cla_h0_v6_fa6_5_xor0 = f_u_csabam8_cla_h0_v6_and6_5 ^ f_u_csabam8_cla_h0_v6_and7_4;
  assign f_u_csabam8_cla_h0_v6_fa6_5_and0 = f_u_csabam8_cla_h0_v6_and6_5 & f_u_csabam8_cla_h0_v6_and7_4;
  assign f_u_csabam8_cla_h0_v6_fa6_5_xor1 = f_u_csabam8_cla_h0_v6_fa6_5_xor0 ^ f_u_csabam8_cla_h0_v6_fa6_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_5_and1 = f_u_csabam8_cla_h0_v6_fa6_5_xor0 & f_u_csabam8_cla_h0_v6_fa6_4_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_5_or0 = f_u_csabam8_cla_h0_v6_fa6_5_and0 | f_u_csabam8_cla_h0_v6_fa6_5_and1;
  assign f_u_csabam8_cla_h0_v6_and7_5 = a[7] & b[5];
  assign f_u_csabam8_cla_h0_v6_and0_6 = a[0] & b[6];
  assign f_u_csabam8_cla_h0_v6_ha0_6_xor0 = f_u_csabam8_cla_h0_v6_and0_6 ^ f_u_csabam8_cla_h0_v6_ha1_5_xor0;
  assign f_u_csabam8_cla_h0_v6_ha0_6_and0 = f_u_csabam8_cla_h0_v6_and0_6 & f_u_csabam8_cla_h0_v6_ha1_5_xor0;
  assign f_u_csabam8_cla_h0_v6_and1_6 = a[1] & b[6];
  assign f_u_csabam8_cla_h0_v6_fa1_6_xor0 = f_u_csabam8_cla_h0_v6_and1_6 ^ f_u_csabam8_cla_h0_v6_fa2_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa1_6_and0 = f_u_csabam8_cla_h0_v6_and1_6 & f_u_csabam8_cla_h0_v6_fa2_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa1_6_xor1 = f_u_csabam8_cla_h0_v6_fa1_6_xor0 ^ f_u_csabam8_cla_h0_v6_ha1_5_and0;
  assign f_u_csabam8_cla_h0_v6_fa1_6_and1 = f_u_csabam8_cla_h0_v6_fa1_6_xor0 & f_u_csabam8_cla_h0_v6_ha1_5_and0;
  assign f_u_csabam8_cla_h0_v6_fa1_6_or0 = f_u_csabam8_cla_h0_v6_fa1_6_and0 | f_u_csabam8_cla_h0_v6_fa1_6_and1;
  assign f_u_csabam8_cla_h0_v6_and2_6 = a[2] & b[6];
  assign f_u_csabam8_cla_h0_v6_fa2_6_xor0 = f_u_csabam8_cla_h0_v6_and2_6 ^ f_u_csabam8_cla_h0_v6_fa3_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa2_6_and0 = f_u_csabam8_cla_h0_v6_and2_6 & f_u_csabam8_cla_h0_v6_fa3_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa2_6_xor1 = f_u_csabam8_cla_h0_v6_fa2_6_xor0 ^ f_u_csabam8_cla_h0_v6_fa2_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa2_6_and1 = f_u_csabam8_cla_h0_v6_fa2_6_xor0 & f_u_csabam8_cla_h0_v6_fa2_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa2_6_or0 = f_u_csabam8_cla_h0_v6_fa2_6_and0 | f_u_csabam8_cla_h0_v6_fa2_6_and1;
  assign f_u_csabam8_cla_h0_v6_and3_6 = a[3] & b[6];
  assign f_u_csabam8_cla_h0_v6_fa3_6_xor0 = f_u_csabam8_cla_h0_v6_and3_6 ^ f_u_csabam8_cla_h0_v6_fa4_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_6_and0 = f_u_csabam8_cla_h0_v6_and3_6 & f_u_csabam8_cla_h0_v6_fa4_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_6_xor1 = f_u_csabam8_cla_h0_v6_fa3_6_xor0 ^ f_u_csabam8_cla_h0_v6_fa3_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa3_6_and1 = f_u_csabam8_cla_h0_v6_fa3_6_xor0 & f_u_csabam8_cla_h0_v6_fa3_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa3_6_or0 = f_u_csabam8_cla_h0_v6_fa3_6_and0 | f_u_csabam8_cla_h0_v6_fa3_6_and1;
  assign f_u_csabam8_cla_h0_v6_and4_6 = a[4] & b[6];
  assign f_u_csabam8_cla_h0_v6_fa4_6_xor0 = f_u_csabam8_cla_h0_v6_and4_6 ^ f_u_csabam8_cla_h0_v6_fa5_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_6_and0 = f_u_csabam8_cla_h0_v6_and4_6 & f_u_csabam8_cla_h0_v6_fa5_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_6_xor1 = f_u_csabam8_cla_h0_v6_fa4_6_xor0 ^ f_u_csabam8_cla_h0_v6_fa4_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_6_and1 = f_u_csabam8_cla_h0_v6_fa4_6_xor0 & f_u_csabam8_cla_h0_v6_fa4_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_6_or0 = f_u_csabam8_cla_h0_v6_fa4_6_and0 | f_u_csabam8_cla_h0_v6_fa4_6_and1;
  assign f_u_csabam8_cla_h0_v6_and5_6 = a[5] & b[6];
  assign f_u_csabam8_cla_h0_v6_fa5_6_xor0 = f_u_csabam8_cla_h0_v6_and5_6 ^ f_u_csabam8_cla_h0_v6_fa6_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_6_and0 = f_u_csabam8_cla_h0_v6_and5_6 & f_u_csabam8_cla_h0_v6_fa6_5_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_6_xor1 = f_u_csabam8_cla_h0_v6_fa5_6_xor0 ^ f_u_csabam8_cla_h0_v6_fa5_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_6_and1 = f_u_csabam8_cla_h0_v6_fa5_6_xor0 & f_u_csabam8_cla_h0_v6_fa5_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_6_or0 = f_u_csabam8_cla_h0_v6_fa5_6_and0 | f_u_csabam8_cla_h0_v6_fa5_6_and1;
  assign f_u_csabam8_cla_h0_v6_and6_6 = a[6] & b[6];
  assign f_u_csabam8_cla_h0_v6_fa6_6_xor0 = f_u_csabam8_cla_h0_v6_and6_6 ^ f_u_csabam8_cla_h0_v6_and7_5;
  assign f_u_csabam8_cla_h0_v6_fa6_6_and0 = f_u_csabam8_cla_h0_v6_and6_6 & f_u_csabam8_cla_h0_v6_and7_5;
  assign f_u_csabam8_cla_h0_v6_fa6_6_xor1 = f_u_csabam8_cla_h0_v6_fa6_6_xor0 ^ f_u_csabam8_cla_h0_v6_fa6_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_6_and1 = f_u_csabam8_cla_h0_v6_fa6_6_xor0 & f_u_csabam8_cla_h0_v6_fa6_5_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_6_or0 = f_u_csabam8_cla_h0_v6_fa6_6_and0 | f_u_csabam8_cla_h0_v6_fa6_6_and1;
  assign f_u_csabam8_cla_h0_v6_and7_6 = a[7] & b[6];
  assign f_u_csabam8_cla_h0_v6_and0_7 = a[0] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa0_7_xor0 = f_u_csabam8_cla_h0_v6_and0_7 ^ f_u_csabam8_cla_h0_v6_fa1_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa0_7_and0 = f_u_csabam8_cla_h0_v6_and0_7 & f_u_csabam8_cla_h0_v6_fa1_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa0_7_xor1 = f_u_csabam8_cla_h0_v6_fa0_7_xor0 ^ f_u_csabam8_cla_h0_v6_ha0_6_and0;
  assign f_u_csabam8_cla_h0_v6_fa0_7_and1 = f_u_csabam8_cla_h0_v6_fa0_7_xor0 & f_u_csabam8_cla_h0_v6_ha0_6_and0;
  assign f_u_csabam8_cla_h0_v6_fa0_7_or0 = f_u_csabam8_cla_h0_v6_fa0_7_and0 | f_u_csabam8_cla_h0_v6_fa0_7_and1;
  assign f_u_csabam8_cla_h0_v6_and1_7 = a[1] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa1_7_xor0 = f_u_csabam8_cla_h0_v6_and1_7 ^ f_u_csabam8_cla_h0_v6_fa2_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa1_7_and0 = f_u_csabam8_cla_h0_v6_and1_7 & f_u_csabam8_cla_h0_v6_fa2_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa1_7_xor1 = f_u_csabam8_cla_h0_v6_fa1_7_xor0 ^ f_u_csabam8_cla_h0_v6_fa1_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa1_7_and1 = f_u_csabam8_cla_h0_v6_fa1_7_xor0 & f_u_csabam8_cla_h0_v6_fa1_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa1_7_or0 = f_u_csabam8_cla_h0_v6_fa1_7_and0 | f_u_csabam8_cla_h0_v6_fa1_7_and1;
  assign f_u_csabam8_cla_h0_v6_and2_7 = a[2] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa2_7_xor0 = f_u_csabam8_cla_h0_v6_and2_7 ^ f_u_csabam8_cla_h0_v6_fa3_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa2_7_and0 = f_u_csabam8_cla_h0_v6_and2_7 & f_u_csabam8_cla_h0_v6_fa3_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa2_7_xor1 = f_u_csabam8_cla_h0_v6_fa2_7_xor0 ^ f_u_csabam8_cla_h0_v6_fa2_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa2_7_and1 = f_u_csabam8_cla_h0_v6_fa2_7_xor0 & f_u_csabam8_cla_h0_v6_fa2_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa2_7_or0 = f_u_csabam8_cla_h0_v6_fa2_7_and0 | f_u_csabam8_cla_h0_v6_fa2_7_and1;
  assign f_u_csabam8_cla_h0_v6_and3_7 = a[3] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa3_7_xor0 = f_u_csabam8_cla_h0_v6_and3_7 ^ f_u_csabam8_cla_h0_v6_fa4_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_7_and0 = f_u_csabam8_cla_h0_v6_and3_7 & f_u_csabam8_cla_h0_v6_fa4_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa3_7_xor1 = f_u_csabam8_cla_h0_v6_fa3_7_xor0 ^ f_u_csabam8_cla_h0_v6_fa3_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa3_7_and1 = f_u_csabam8_cla_h0_v6_fa3_7_xor0 & f_u_csabam8_cla_h0_v6_fa3_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa3_7_or0 = f_u_csabam8_cla_h0_v6_fa3_7_and0 | f_u_csabam8_cla_h0_v6_fa3_7_and1;
  assign f_u_csabam8_cla_h0_v6_and4_7 = a[4] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa4_7_xor0 = f_u_csabam8_cla_h0_v6_and4_7 ^ f_u_csabam8_cla_h0_v6_fa5_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_7_and0 = f_u_csabam8_cla_h0_v6_and4_7 & f_u_csabam8_cla_h0_v6_fa5_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa4_7_xor1 = f_u_csabam8_cla_h0_v6_fa4_7_xor0 ^ f_u_csabam8_cla_h0_v6_fa4_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_7_and1 = f_u_csabam8_cla_h0_v6_fa4_7_xor0 & f_u_csabam8_cla_h0_v6_fa4_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa4_7_or0 = f_u_csabam8_cla_h0_v6_fa4_7_and0 | f_u_csabam8_cla_h0_v6_fa4_7_and1;
  assign f_u_csabam8_cla_h0_v6_and5_7 = a[5] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa5_7_xor0 = f_u_csabam8_cla_h0_v6_and5_7 ^ f_u_csabam8_cla_h0_v6_fa6_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_7_and0 = f_u_csabam8_cla_h0_v6_and5_7 & f_u_csabam8_cla_h0_v6_fa6_6_xor1;
  assign f_u_csabam8_cla_h0_v6_fa5_7_xor1 = f_u_csabam8_cla_h0_v6_fa5_7_xor0 ^ f_u_csabam8_cla_h0_v6_fa5_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_7_and1 = f_u_csabam8_cla_h0_v6_fa5_7_xor0 & f_u_csabam8_cla_h0_v6_fa5_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa5_7_or0 = f_u_csabam8_cla_h0_v6_fa5_7_and0 | f_u_csabam8_cla_h0_v6_fa5_7_and1;
  assign f_u_csabam8_cla_h0_v6_and6_7 = a[6] & b[7];
  assign f_u_csabam8_cla_h0_v6_fa6_7_xor0 = f_u_csabam8_cla_h0_v6_and6_7 ^ f_u_csabam8_cla_h0_v6_and7_6;
  assign f_u_csabam8_cla_h0_v6_fa6_7_and0 = f_u_csabam8_cla_h0_v6_and6_7 & f_u_csabam8_cla_h0_v6_and7_6;
  assign f_u_csabam8_cla_h0_v6_fa6_7_xor1 = f_u_csabam8_cla_h0_v6_fa6_7_xor0 ^ f_u_csabam8_cla_h0_v6_fa6_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_7_and1 = f_u_csabam8_cla_h0_v6_fa6_7_xor0 & f_u_csabam8_cla_h0_v6_fa6_6_or0;
  assign f_u_csabam8_cla_h0_v6_fa6_7_or0 = f_u_csabam8_cla_h0_v6_fa6_7_and0 | f_u_csabam8_cla_h0_v6_fa6_7_and1;
  assign f_u_csabam8_cla_h0_v6_and7_7 = a[7] & b[7];
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_or0 = f_u_csabam8_cla_h0_v6_fa1_7_xor1 | f_u_csabam8_cla_h0_v6_fa0_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_and0 = f_u_csabam8_cla_h0_v6_fa1_7_xor1 & f_u_csabam8_cla_h0_v6_fa0_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_xor0 = f_u_csabam8_cla_h0_v6_fa1_7_xor1 ^ f_u_csabam8_cla_h0_v6_fa0_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_or0 = f_u_csabam8_cla_h0_v6_fa2_7_xor1 | f_u_csabam8_cla_h0_v6_fa1_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_and0 = f_u_csabam8_cla_h0_v6_fa2_7_xor1 & f_u_csabam8_cla_h0_v6_fa1_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_xor0 = f_u_csabam8_cla_h0_v6_fa2_7_xor1 ^ f_u_csabam8_cla_h0_v6_fa1_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_xor1 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_xor0 ^ f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_and0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and0 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or0 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_and0 | f_u_csabam8_cla_h0_v6_u_cla8_and0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0 = f_u_csabam8_cla_h0_v6_fa3_7_xor1 | f_u_csabam8_cla_h0_v6_fa2_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_and0 = f_u_csabam8_cla_h0_v6_fa3_7_xor1 & f_u_csabam8_cla_h0_v6_fa2_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_xor0 = f_u_csabam8_cla_h0_v6_fa3_7_xor1 ^ f_u_csabam8_cla_h0_v6_fa2_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_xor2 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_xor0 ^ f_u_csabam8_cla_h0_v6_u_cla8_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and1 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and2 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and3 = f_u_csabam8_cla_h0_v6_u_cla8_and2 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and4 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or1 = f_u_csabam8_cla_h0_v6_u_cla8_and3 | f_u_csabam8_cla_h0_v6_u_cla8_and4;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or2 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_and0 | f_u_csabam8_cla_h0_v6_u_cla8_or1;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_or0 = f_u_csabam8_cla_h0_v6_fa4_7_xor1 | f_u_csabam8_cla_h0_v6_fa3_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_and0 = f_u_csabam8_cla_h0_v6_fa4_7_xor1 & f_u_csabam8_cla_h0_v6_fa3_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_xor0 = f_u_csabam8_cla_h0_v6_fa4_7_xor1 ^ f_u_csabam8_cla_h0_v6_fa3_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_xor3 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_xor0 ^ f_u_csabam8_cla_h0_v6_u_cla8_or2;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and5 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_or0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and6 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and7 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_or0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and8 = f_u_csabam8_cla_h0_v6_u_cla8_and6 & f_u_csabam8_cla_h0_v6_u_cla8_and7;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and9 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic1_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and10 = f_u_csabam8_cla_h0_v6_u_cla8_and9 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and11 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic2_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or3 = f_u_csabam8_cla_h0_v6_u_cla8_and8 | f_u_csabam8_cla_h0_v6_u_cla8_and11;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or4 = f_u_csabam8_cla_h0_v6_u_cla8_and10 | f_u_csabam8_cla_h0_v6_u_cla8_or3;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or5 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic3_and0 | f_u_csabam8_cla_h0_v6_u_cla8_or4;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_or0 = f_u_csabam8_cla_h0_v6_fa5_7_xor1 | f_u_csabam8_cla_h0_v6_fa4_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_and0 = f_u_csabam8_cla_h0_v6_fa5_7_xor1 & f_u_csabam8_cla_h0_v6_fa4_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_xor0 = f_u_csabam8_cla_h0_v6_fa5_7_xor1 ^ f_u_csabam8_cla_h0_v6_fa4_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_xor4 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_xor0 ^ f_u_csabam8_cla_h0_v6_u_cla8_or5;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and12 = f_u_csabam8_cla_h0_v6_u_cla8_or5 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or6 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_and0 | f_u_csabam8_cla_h0_v6_u_cla8_and12;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_or0 = f_u_csabam8_cla_h0_v6_fa6_7_xor1 | f_u_csabam8_cla_h0_v6_fa5_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_and0 = f_u_csabam8_cla_h0_v6_fa6_7_xor1 & f_u_csabam8_cla_h0_v6_fa5_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_xor0 = f_u_csabam8_cla_h0_v6_fa6_7_xor1 ^ f_u_csabam8_cla_h0_v6_fa5_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_xor5 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_xor0 ^ f_u_csabam8_cla_h0_v6_u_cla8_or6;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and13 = f_u_csabam8_cla_h0_v6_u_cla8_or5 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and14 = f_u_csabam8_cla_h0_v6_u_cla8_and13 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and15 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or7 = f_u_csabam8_cla_h0_v6_u_cla8_and14 | f_u_csabam8_cla_h0_v6_u_cla8_and15;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or8 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_and0 | f_u_csabam8_cla_h0_v6_u_cla8_or7;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0 = f_u_csabam8_cla_h0_v6_and7_7 | f_u_csabam8_cla_h0_v6_fa6_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_and0 = f_u_csabam8_cla_h0_v6_and7_7 & f_u_csabam8_cla_h0_v6_fa6_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_xor0 = f_u_csabam8_cla_h0_v6_and7_7 ^ f_u_csabam8_cla_h0_v6_fa6_7_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_xor6 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_xor0 ^ f_u_csabam8_cla_h0_v6_u_cla8_or8;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and16 = f_u_csabam8_cla_h0_v6_u_cla8_or5 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and17 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and18 = f_u_csabam8_cla_h0_v6_u_cla8_and16 & f_u_csabam8_cla_h0_v6_u_cla8_and17;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and19 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and20 = f_u_csabam8_cla_h0_v6_u_cla8_and19 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and21 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic5_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or9 = f_u_csabam8_cla_h0_v6_u_cla8_and18 | f_u_csabam8_cla_h0_v6_u_cla8_and20;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or10 = f_u_csabam8_cla_h0_v6_u_cla8_or9 | f_u_csabam8_cla_h0_v6_u_cla8_and21;
  assign f_u_csabam8_cla_h0_v6_u_cla8_or11 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_and0 | f_u_csabam8_cla_h0_v6_u_cla8_or10;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and22 = f_u_csabam8_cla_h0_v6_u_cla8_or5 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0;
  assign f_u_csabam8_cla_h0_v6_u_cla8_and23 = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic4_and0 & f_u_csabam8_cla_h0_v6_u_cla8_pg_logic6_or0;

  assign f_u_csabam8_cla_h0_v6_out[0] = 1'b0;
  assign f_u_csabam8_cla_h0_v6_out[1] = 1'b0;
  assign f_u_csabam8_cla_h0_v6_out[2] = 1'b0;
  assign f_u_csabam8_cla_h0_v6_out[3] = 1'b0;
  assign f_u_csabam8_cla_h0_v6_out[4] = 1'b0;
  assign f_u_csabam8_cla_h0_v6_out[5] = 1'b0;
  assign f_u_csabam8_cla_h0_v6_out[6] = f_u_csabam8_cla_h0_v6_ha0_6_xor0;
  assign f_u_csabam8_cla_h0_v6_out[7] = f_u_csabam8_cla_h0_v6_fa0_7_xor1;
  assign f_u_csabam8_cla_h0_v6_out[8] = f_u_csabam8_cla_h0_v6_u_cla8_pg_logic0_xor0;
  assign f_u_csabam8_cla_h0_v6_out[9] = f_u_csabam8_cla_h0_v6_u_cla8_xor1;
  assign f_u_csabam8_cla_h0_v6_out[10] = f_u_csabam8_cla_h0_v6_u_cla8_xor2;
  assign f_u_csabam8_cla_h0_v6_out[11] = f_u_csabam8_cla_h0_v6_u_cla8_xor3;
  assign f_u_csabam8_cla_h0_v6_out[12] = f_u_csabam8_cla_h0_v6_u_cla8_xor4;
  assign f_u_csabam8_cla_h0_v6_out[13] = f_u_csabam8_cla_h0_v6_u_cla8_xor5;
  assign f_u_csabam8_cla_h0_v6_out[14] = f_u_csabam8_cla_h0_v6_u_cla8_xor6;
  assign f_u_csabam8_cla_h0_v6_out[15] = f_u_csabam8_cla_h0_v6_u_cla8_or11;
endmodule