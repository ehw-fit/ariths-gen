module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;
  wire constant_wire_value_1_y0;
  wire constant_wire_value_1_y1;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_y0;
  wire fa_y1;
  wire fa_cin;
  wire fa_y3;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module h_s_arrmul12(input [11:0] a, input [11:0] b, output [23:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire constant_wire_1;
  wire h_s_arrmul12_and0_0_y0;
  wire h_s_arrmul12_and1_0_y0;
  wire h_s_arrmul12_and2_0_y0;
  wire h_s_arrmul12_and3_0_y0;
  wire h_s_arrmul12_and4_0_y0;
  wire h_s_arrmul12_and5_0_y0;
  wire h_s_arrmul12_and6_0_y0;
  wire h_s_arrmul12_and7_0_y0;
  wire h_s_arrmul12_and8_0_y0;
  wire h_s_arrmul12_and9_0_y0;
  wire h_s_arrmul12_and10_0_y0;
  wire h_s_arrmul12_nand11_0_y0;
  wire h_s_arrmul12_and0_1_y0;
  wire h_s_arrmul12_ha0_1_y0;
  wire h_s_arrmul12_ha0_1_y1;
  wire h_s_arrmul12_and1_1_y0;
  wire h_s_arrmul12_fa1_1_y2;
  wire h_s_arrmul12_fa1_1_y4;
  wire h_s_arrmul12_and2_1_y0;
  wire h_s_arrmul12_fa2_1_y2;
  wire h_s_arrmul12_fa2_1_y4;
  wire h_s_arrmul12_and3_1_y0;
  wire h_s_arrmul12_fa3_1_y2;
  wire h_s_arrmul12_fa3_1_y4;
  wire h_s_arrmul12_and4_1_y0;
  wire h_s_arrmul12_fa4_1_y2;
  wire h_s_arrmul12_fa4_1_y4;
  wire h_s_arrmul12_and5_1_y0;
  wire h_s_arrmul12_fa5_1_y2;
  wire h_s_arrmul12_fa5_1_y4;
  wire h_s_arrmul12_and6_1_y0;
  wire h_s_arrmul12_fa6_1_y2;
  wire h_s_arrmul12_fa6_1_y4;
  wire h_s_arrmul12_and7_1_y0;
  wire h_s_arrmul12_fa7_1_y2;
  wire h_s_arrmul12_fa7_1_y4;
  wire h_s_arrmul12_and8_1_y0;
  wire h_s_arrmul12_fa8_1_y2;
  wire h_s_arrmul12_fa8_1_y4;
  wire h_s_arrmul12_and9_1_y0;
  wire h_s_arrmul12_fa9_1_y2;
  wire h_s_arrmul12_fa9_1_y4;
  wire h_s_arrmul12_and10_1_y0;
  wire h_s_arrmul12_fa10_1_y2;
  wire h_s_arrmul12_fa10_1_y4;
  wire h_s_arrmul12_nand11_1_y0;
  wire h_s_arrmul12_fa11_1_y2;
  wire h_s_arrmul12_fa11_1_y4;
  wire h_s_arrmul12_and0_2_y0;
  wire h_s_arrmul12_ha0_2_y0;
  wire h_s_arrmul12_ha0_2_y1;
  wire h_s_arrmul12_and1_2_y0;
  wire h_s_arrmul12_fa1_2_y2;
  wire h_s_arrmul12_fa1_2_y4;
  wire h_s_arrmul12_and2_2_y0;
  wire h_s_arrmul12_fa2_2_y2;
  wire h_s_arrmul12_fa2_2_y4;
  wire h_s_arrmul12_and3_2_y0;
  wire h_s_arrmul12_fa3_2_y2;
  wire h_s_arrmul12_fa3_2_y4;
  wire h_s_arrmul12_and4_2_y0;
  wire h_s_arrmul12_fa4_2_y2;
  wire h_s_arrmul12_fa4_2_y4;
  wire h_s_arrmul12_and5_2_y0;
  wire h_s_arrmul12_fa5_2_y2;
  wire h_s_arrmul12_fa5_2_y4;
  wire h_s_arrmul12_and6_2_y0;
  wire h_s_arrmul12_fa6_2_y2;
  wire h_s_arrmul12_fa6_2_y4;
  wire h_s_arrmul12_and7_2_y0;
  wire h_s_arrmul12_fa7_2_y2;
  wire h_s_arrmul12_fa7_2_y4;
  wire h_s_arrmul12_and8_2_y0;
  wire h_s_arrmul12_fa8_2_y2;
  wire h_s_arrmul12_fa8_2_y4;
  wire h_s_arrmul12_and9_2_y0;
  wire h_s_arrmul12_fa9_2_y2;
  wire h_s_arrmul12_fa9_2_y4;
  wire h_s_arrmul12_and10_2_y0;
  wire h_s_arrmul12_fa10_2_y2;
  wire h_s_arrmul12_fa10_2_y4;
  wire h_s_arrmul12_nand11_2_y0;
  wire h_s_arrmul12_fa11_2_y2;
  wire h_s_arrmul12_fa11_2_y4;
  wire h_s_arrmul12_and0_3_y0;
  wire h_s_arrmul12_ha0_3_y0;
  wire h_s_arrmul12_ha0_3_y1;
  wire h_s_arrmul12_and1_3_y0;
  wire h_s_arrmul12_fa1_3_y2;
  wire h_s_arrmul12_fa1_3_y4;
  wire h_s_arrmul12_and2_3_y0;
  wire h_s_arrmul12_fa2_3_y2;
  wire h_s_arrmul12_fa2_3_y4;
  wire h_s_arrmul12_and3_3_y0;
  wire h_s_arrmul12_fa3_3_y2;
  wire h_s_arrmul12_fa3_3_y4;
  wire h_s_arrmul12_and4_3_y0;
  wire h_s_arrmul12_fa4_3_y2;
  wire h_s_arrmul12_fa4_3_y4;
  wire h_s_arrmul12_and5_3_y0;
  wire h_s_arrmul12_fa5_3_y2;
  wire h_s_arrmul12_fa5_3_y4;
  wire h_s_arrmul12_and6_3_y0;
  wire h_s_arrmul12_fa6_3_y2;
  wire h_s_arrmul12_fa6_3_y4;
  wire h_s_arrmul12_and7_3_y0;
  wire h_s_arrmul12_fa7_3_y2;
  wire h_s_arrmul12_fa7_3_y4;
  wire h_s_arrmul12_and8_3_y0;
  wire h_s_arrmul12_fa8_3_y2;
  wire h_s_arrmul12_fa8_3_y4;
  wire h_s_arrmul12_and9_3_y0;
  wire h_s_arrmul12_fa9_3_y2;
  wire h_s_arrmul12_fa9_3_y4;
  wire h_s_arrmul12_and10_3_y0;
  wire h_s_arrmul12_fa10_3_y2;
  wire h_s_arrmul12_fa10_3_y4;
  wire h_s_arrmul12_nand11_3_y0;
  wire h_s_arrmul12_fa11_3_y2;
  wire h_s_arrmul12_fa11_3_y4;
  wire h_s_arrmul12_and0_4_y0;
  wire h_s_arrmul12_ha0_4_y0;
  wire h_s_arrmul12_ha0_4_y1;
  wire h_s_arrmul12_and1_4_y0;
  wire h_s_arrmul12_fa1_4_y2;
  wire h_s_arrmul12_fa1_4_y4;
  wire h_s_arrmul12_and2_4_y0;
  wire h_s_arrmul12_fa2_4_y2;
  wire h_s_arrmul12_fa2_4_y4;
  wire h_s_arrmul12_and3_4_y0;
  wire h_s_arrmul12_fa3_4_y2;
  wire h_s_arrmul12_fa3_4_y4;
  wire h_s_arrmul12_and4_4_y0;
  wire h_s_arrmul12_fa4_4_y2;
  wire h_s_arrmul12_fa4_4_y4;
  wire h_s_arrmul12_and5_4_y0;
  wire h_s_arrmul12_fa5_4_y2;
  wire h_s_arrmul12_fa5_4_y4;
  wire h_s_arrmul12_and6_4_y0;
  wire h_s_arrmul12_fa6_4_y2;
  wire h_s_arrmul12_fa6_4_y4;
  wire h_s_arrmul12_and7_4_y0;
  wire h_s_arrmul12_fa7_4_y2;
  wire h_s_arrmul12_fa7_4_y4;
  wire h_s_arrmul12_and8_4_y0;
  wire h_s_arrmul12_fa8_4_y2;
  wire h_s_arrmul12_fa8_4_y4;
  wire h_s_arrmul12_and9_4_y0;
  wire h_s_arrmul12_fa9_4_y2;
  wire h_s_arrmul12_fa9_4_y4;
  wire h_s_arrmul12_and10_4_y0;
  wire h_s_arrmul12_fa10_4_y2;
  wire h_s_arrmul12_fa10_4_y4;
  wire h_s_arrmul12_nand11_4_y0;
  wire h_s_arrmul12_fa11_4_y2;
  wire h_s_arrmul12_fa11_4_y4;
  wire h_s_arrmul12_and0_5_y0;
  wire h_s_arrmul12_ha0_5_y0;
  wire h_s_arrmul12_ha0_5_y1;
  wire h_s_arrmul12_and1_5_y0;
  wire h_s_arrmul12_fa1_5_y2;
  wire h_s_arrmul12_fa1_5_y4;
  wire h_s_arrmul12_and2_5_y0;
  wire h_s_arrmul12_fa2_5_y2;
  wire h_s_arrmul12_fa2_5_y4;
  wire h_s_arrmul12_and3_5_y0;
  wire h_s_arrmul12_fa3_5_y2;
  wire h_s_arrmul12_fa3_5_y4;
  wire h_s_arrmul12_and4_5_y0;
  wire h_s_arrmul12_fa4_5_y2;
  wire h_s_arrmul12_fa4_5_y4;
  wire h_s_arrmul12_and5_5_y0;
  wire h_s_arrmul12_fa5_5_y2;
  wire h_s_arrmul12_fa5_5_y4;
  wire h_s_arrmul12_and6_5_y0;
  wire h_s_arrmul12_fa6_5_y2;
  wire h_s_arrmul12_fa6_5_y4;
  wire h_s_arrmul12_and7_5_y0;
  wire h_s_arrmul12_fa7_5_y2;
  wire h_s_arrmul12_fa7_5_y4;
  wire h_s_arrmul12_and8_5_y0;
  wire h_s_arrmul12_fa8_5_y2;
  wire h_s_arrmul12_fa8_5_y4;
  wire h_s_arrmul12_and9_5_y0;
  wire h_s_arrmul12_fa9_5_y2;
  wire h_s_arrmul12_fa9_5_y4;
  wire h_s_arrmul12_and10_5_y0;
  wire h_s_arrmul12_fa10_5_y2;
  wire h_s_arrmul12_fa10_5_y4;
  wire h_s_arrmul12_nand11_5_y0;
  wire h_s_arrmul12_fa11_5_y2;
  wire h_s_arrmul12_fa11_5_y4;
  wire h_s_arrmul12_and0_6_y0;
  wire h_s_arrmul12_ha0_6_y0;
  wire h_s_arrmul12_ha0_6_y1;
  wire h_s_arrmul12_and1_6_y0;
  wire h_s_arrmul12_fa1_6_y2;
  wire h_s_arrmul12_fa1_6_y4;
  wire h_s_arrmul12_and2_6_y0;
  wire h_s_arrmul12_fa2_6_y2;
  wire h_s_arrmul12_fa2_6_y4;
  wire h_s_arrmul12_and3_6_y0;
  wire h_s_arrmul12_fa3_6_y2;
  wire h_s_arrmul12_fa3_6_y4;
  wire h_s_arrmul12_and4_6_y0;
  wire h_s_arrmul12_fa4_6_y2;
  wire h_s_arrmul12_fa4_6_y4;
  wire h_s_arrmul12_and5_6_y0;
  wire h_s_arrmul12_fa5_6_y2;
  wire h_s_arrmul12_fa5_6_y4;
  wire h_s_arrmul12_and6_6_y0;
  wire h_s_arrmul12_fa6_6_y2;
  wire h_s_arrmul12_fa6_6_y4;
  wire h_s_arrmul12_and7_6_y0;
  wire h_s_arrmul12_fa7_6_y2;
  wire h_s_arrmul12_fa7_6_y4;
  wire h_s_arrmul12_and8_6_y0;
  wire h_s_arrmul12_fa8_6_y2;
  wire h_s_arrmul12_fa8_6_y4;
  wire h_s_arrmul12_and9_6_y0;
  wire h_s_arrmul12_fa9_6_y2;
  wire h_s_arrmul12_fa9_6_y4;
  wire h_s_arrmul12_and10_6_y0;
  wire h_s_arrmul12_fa10_6_y2;
  wire h_s_arrmul12_fa10_6_y4;
  wire h_s_arrmul12_nand11_6_y0;
  wire h_s_arrmul12_fa11_6_y2;
  wire h_s_arrmul12_fa11_6_y4;
  wire h_s_arrmul12_and0_7_y0;
  wire h_s_arrmul12_ha0_7_y0;
  wire h_s_arrmul12_ha0_7_y1;
  wire h_s_arrmul12_and1_7_y0;
  wire h_s_arrmul12_fa1_7_y2;
  wire h_s_arrmul12_fa1_7_y4;
  wire h_s_arrmul12_and2_7_y0;
  wire h_s_arrmul12_fa2_7_y2;
  wire h_s_arrmul12_fa2_7_y4;
  wire h_s_arrmul12_and3_7_y0;
  wire h_s_arrmul12_fa3_7_y2;
  wire h_s_arrmul12_fa3_7_y4;
  wire h_s_arrmul12_and4_7_y0;
  wire h_s_arrmul12_fa4_7_y2;
  wire h_s_arrmul12_fa4_7_y4;
  wire h_s_arrmul12_and5_7_y0;
  wire h_s_arrmul12_fa5_7_y2;
  wire h_s_arrmul12_fa5_7_y4;
  wire h_s_arrmul12_and6_7_y0;
  wire h_s_arrmul12_fa6_7_y2;
  wire h_s_arrmul12_fa6_7_y4;
  wire h_s_arrmul12_and7_7_y0;
  wire h_s_arrmul12_fa7_7_y2;
  wire h_s_arrmul12_fa7_7_y4;
  wire h_s_arrmul12_and8_7_y0;
  wire h_s_arrmul12_fa8_7_y2;
  wire h_s_arrmul12_fa8_7_y4;
  wire h_s_arrmul12_and9_7_y0;
  wire h_s_arrmul12_fa9_7_y2;
  wire h_s_arrmul12_fa9_7_y4;
  wire h_s_arrmul12_and10_7_y0;
  wire h_s_arrmul12_fa10_7_y2;
  wire h_s_arrmul12_fa10_7_y4;
  wire h_s_arrmul12_nand11_7_y0;
  wire h_s_arrmul12_fa11_7_y2;
  wire h_s_arrmul12_fa11_7_y4;
  wire h_s_arrmul12_and0_8_y0;
  wire h_s_arrmul12_ha0_8_y0;
  wire h_s_arrmul12_ha0_8_y1;
  wire h_s_arrmul12_and1_8_y0;
  wire h_s_arrmul12_fa1_8_y2;
  wire h_s_arrmul12_fa1_8_y4;
  wire h_s_arrmul12_and2_8_y0;
  wire h_s_arrmul12_fa2_8_y2;
  wire h_s_arrmul12_fa2_8_y4;
  wire h_s_arrmul12_and3_8_y0;
  wire h_s_arrmul12_fa3_8_y2;
  wire h_s_arrmul12_fa3_8_y4;
  wire h_s_arrmul12_and4_8_y0;
  wire h_s_arrmul12_fa4_8_y2;
  wire h_s_arrmul12_fa4_8_y4;
  wire h_s_arrmul12_and5_8_y0;
  wire h_s_arrmul12_fa5_8_y2;
  wire h_s_arrmul12_fa5_8_y4;
  wire h_s_arrmul12_and6_8_y0;
  wire h_s_arrmul12_fa6_8_y2;
  wire h_s_arrmul12_fa6_8_y4;
  wire h_s_arrmul12_and7_8_y0;
  wire h_s_arrmul12_fa7_8_y2;
  wire h_s_arrmul12_fa7_8_y4;
  wire h_s_arrmul12_and8_8_y0;
  wire h_s_arrmul12_fa8_8_y2;
  wire h_s_arrmul12_fa8_8_y4;
  wire h_s_arrmul12_and9_8_y0;
  wire h_s_arrmul12_fa9_8_y2;
  wire h_s_arrmul12_fa9_8_y4;
  wire h_s_arrmul12_and10_8_y0;
  wire h_s_arrmul12_fa10_8_y2;
  wire h_s_arrmul12_fa10_8_y4;
  wire h_s_arrmul12_nand11_8_y0;
  wire h_s_arrmul12_fa11_8_y2;
  wire h_s_arrmul12_fa11_8_y4;
  wire h_s_arrmul12_and0_9_y0;
  wire h_s_arrmul12_ha0_9_y0;
  wire h_s_arrmul12_ha0_9_y1;
  wire h_s_arrmul12_and1_9_y0;
  wire h_s_arrmul12_fa1_9_y2;
  wire h_s_arrmul12_fa1_9_y4;
  wire h_s_arrmul12_and2_9_y0;
  wire h_s_arrmul12_fa2_9_y2;
  wire h_s_arrmul12_fa2_9_y4;
  wire h_s_arrmul12_and3_9_y0;
  wire h_s_arrmul12_fa3_9_y2;
  wire h_s_arrmul12_fa3_9_y4;
  wire h_s_arrmul12_and4_9_y0;
  wire h_s_arrmul12_fa4_9_y2;
  wire h_s_arrmul12_fa4_9_y4;
  wire h_s_arrmul12_and5_9_y0;
  wire h_s_arrmul12_fa5_9_y2;
  wire h_s_arrmul12_fa5_9_y4;
  wire h_s_arrmul12_and6_9_y0;
  wire h_s_arrmul12_fa6_9_y2;
  wire h_s_arrmul12_fa6_9_y4;
  wire h_s_arrmul12_and7_9_y0;
  wire h_s_arrmul12_fa7_9_y2;
  wire h_s_arrmul12_fa7_9_y4;
  wire h_s_arrmul12_and8_9_y0;
  wire h_s_arrmul12_fa8_9_y2;
  wire h_s_arrmul12_fa8_9_y4;
  wire h_s_arrmul12_and9_9_y0;
  wire h_s_arrmul12_fa9_9_y2;
  wire h_s_arrmul12_fa9_9_y4;
  wire h_s_arrmul12_and10_9_y0;
  wire h_s_arrmul12_fa10_9_y2;
  wire h_s_arrmul12_fa10_9_y4;
  wire h_s_arrmul12_nand11_9_y0;
  wire h_s_arrmul12_fa11_9_y2;
  wire h_s_arrmul12_fa11_9_y4;
  wire h_s_arrmul12_and0_10_y0;
  wire h_s_arrmul12_ha0_10_y0;
  wire h_s_arrmul12_ha0_10_y1;
  wire h_s_arrmul12_and1_10_y0;
  wire h_s_arrmul12_fa1_10_y2;
  wire h_s_arrmul12_fa1_10_y4;
  wire h_s_arrmul12_and2_10_y0;
  wire h_s_arrmul12_fa2_10_y2;
  wire h_s_arrmul12_fa2_10_y4;
  wire h_s_arrmul12_and3_10_y0;
  wire h_s_arrmul12_fa3_10_y2;
  wire h_s_arrmul12_fa3_10_y4;
  wire h_s_arrmul12_and4_10_y0;
  wire h_s_arrmul12_fa4_10_y2;
  wire h_s_arrmul12_fa4_10_y4;
  wire h_s_arrmul12_and5_10_y0;
  wire h_s_arrmul12_fa5_10_y2;
  wire h_s_arrmul12_fa5_10_y4;
  wire h_s_arrmul12_and6_10_y0;
  wire h_s_arrmul12_fa6_10_y2;
  wire h_s_arrmul12_fa6_10_y4;
  wire h_s_arrmul12_and7_10_y0;
  wire h_s_arrmul12_fa7_10_y2;
  wire h_s_arrmul12_fa7_10_y4;
  wire h_s_arrmul12_and8_10_y0;
  wire h_s_arrmul12_fa8_10_y2;
  wire h_s_arrmul12_fa8_10_y4;
  wire h_s_arrmul12_and9_10_y0;
  wire h_s_arrmul12_fa9_10_y2;
  wire h_s_arrmul12_fa9_10_y4;
  wire h_s_arrmul12_and10_10_y0;
  wire h_s_arrmul12_fa10_10_y2;
  wire h_s_arrmul12_fa10_10_y4;
  wire h_s_arrmul12_nand11_10_y0;
  wire h_s_arrmul12_fa11_10_y2;
  wire h_s_arrmul12_fa11_10_y4;
  wire h_s_arrmul12_nand0_11_y0;
  wire h_s_arrmul12_ha0_11_y0;
  wire h_s_arrmul12_ha0_11_y1;
  wire h_s_arrmul12_nand1_11_y0;
  wire h_s_arrmul12_fa1_11_y2;
  wire h_s_arrmul12_fa1_11_y4;
  wire h_s_arrmul12_nand2_11_y0;
  wire h_s_arrmul12_fa2_11_y2;
  wire h_s_arrmul12_fa2_11_y4;
  wire h_s_arrmul12_nand3_11_y0;
  wire h_s_arrmul12_fa3_11_y2;
  wire h_s_arrmul12_fa3_11_y4;
  wire h_s_arrmul12_nand4_11_y0;
  wire h_s_arrmul12_fa4_11_y2;
  wire h_s_arrmul12_fa4_11_y4;
  wire h_s_arrmul12_nand5_11_y0;
  wire h_s_arrmul12_fa5_11_y2;
  wire h_s_arrmul12_fa5_11_y4;
  wire h_s_arrmul12_nand6_11_y0;
  wire h_s_arrmul12_fa6_11_y2;
  wire h_s_arrmul12_fa6_11_y4;
  wire h_s_arrmul12_nand7_11_y0;
  wire h_s_arrmul12_fa7_11_y2;
  wire h_s_arrmul12_fa7_11_y4;
  wire h_s_arrmul12_nand8_11_y0;
  wire h_s_arrmul12_fa8_11_y2;
  wire h_s_arrmul12_fa8_11_y4;
  wire h_s_arrmul12_nand9_11_y0;
  wire h_s_arrmul12_fa9_11_y2;
  wire h_s_arrmul12_fa9_11_y4;
  wire h_s_arrmul12_nand10_11_y0;
  wire h_s_arrmul12_fa10_11_y2;
  wire h_s_arrmul12_fa10_11_y4;
  wire h_s_arrmul12_and11_11_y0;
  wire h_s_arrmul12_fa11_11_y2;
  wire h_s_arrmul12_fa11_11_y4;
  wire h_s_arrmul12_xor12_11_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_arrmul12_and0_0_y0(a_0, b_0, h_s_arrmul12_and0_0_y0);
  and_gate and_gate_h_s_arrmul12_and1_0_y0(a_1, b_0, h_s_arrmul12_and1_0_y0);
  and_gate and_gate_h_s_arrmul12_and2_0_y0(a_2, b_0, h_s_arrmul12_and2_0_y0);
  and_gate and_gate_h_s_arrmul12_and3_0_y0(a_3, b_0, h_s_arrmul12_and3_0_y0);
  and_gate and_gate_h_s_arrmul12_and4_0_y0(a_4, b_0, h_s_arrmul12_and4_0_y0);
  and_gate and_gate_h_s_arrmul12_and5_0_y0(a_5, b_0, h_s_arrmul12_and5_0_y0);
  and_gate and_gate_h_s_arrmul12_and6_0_y0(a_6, b_0, h_s_arrmul12_and6_0_y0);
  and_gate and_gate_h_s_arrmul12_and7_0_y0(a_7, b_0, h_s_arrmul12_and7_0_y0);
  and_gate and_gate_h_s_arrmul12_and8_0_y0(a_8, b_0, h_s_arrmul12_and8_0_y0);
  and_gate and_gate_h_s_arrmul12_and9_0_y0(a_9, b_0, h_s_arrmul12_and9_0_y0);
  and_gate and_gate_h_s_arrmul12_and10_0_y0(a_10, b_0, h_s_arrmul12_and10_0_y0);
  nand_gate nand_gate_h_s_arrmul12_nand11_0_y0(a_11, b_0, h_s_arrmul12_nand11_0_y0);
  and_gate and_gate_h_s_arrmul12_and0_1_y0(a_0, b_1, h_s_arrmul12_and0_1_y0);
  ha ha_h_s_arrmul12_ha0_1_y0(h_s_arrmul12_and0_1_y0, h_s_arrmul12_and1_0_y0, h_s_arrmul12_ha0_1_y0, h_s_arrmul12_ha0_1_y1);
  and_gate and_gate_h_s_arrmul12_and1_1_y0(a_1, b_1, h_s_arrmul12_and1_1_y0);
  fa fa_h_s_arrmul12_fa1_1_y2(h_s_arrmul12_and1_1_y0, h_s_arrmul12_and2_0_y0, h_s_arrmul12_ha0_1_y1, h_s_arrmul12_fa1_1_y2, h_s_arrmul12_fa1_1_y4);
  and_gate and_gate_h_s_arrmul12_and2_1_y0(a_2, b_1, h_s_arrmul12_and2_1_y0);
  fa fa_h_s_arrmul12_fa2_1_y2(h_s_arrmul12_and2_1_y0, h_s_arrmul12_and3_0_y0, h_s_arrmul12_fa1_1_y4, h_s_arrmul12_fa2_1_y2, h_s_arrmul12_fa2_1_y4);
  and_gate and_gate_h_s_arrmul12_and3_1_y0(a_3, b_1, h_s_arrmul12_and3_1_y0);
  fa fa_h_s_arrmul12_fa3_1_y2(h_s_arrmul12_and3_1_y0, h_s_arrmul12_and4_0_y0, h_s_arrmul12_fa2_1_y4, h_s_arrmul12_fa3_1_y2, h_s_arrmul12_fa3_1_y4);
  and_gate and_gate_h_s_arrmul12_and4_1_y0(a_4, b_1, h_s_arrmul12_and4_1_y0);
  fa fa_h_s_arrmul12_fa4_1_y2(h_s_arrmul12_and4_1_y0, h_s_arrmul12_and5_0_y0, h_s_arrmul12_fa3_1_y4, h_s_arrmul12_fa4_1_y2, h_s_arrmul12_fa4_1_y4);
  and_gate and_gate_h_s_arrmul12_and5_1_y0(a_5, b_1, h_s_arrmul12_and5_1_y0);
  fa fa_h_s_arrmul12_fa5_1_y2(h_s_arrmul12_and5_1_y0, h_s_arrmul12_and6_0_y0, h_s_arrmul12_fa4_1_y4, h_s_arrmul12_fa5_1_y2, h_s_arrmul12_fa5_1_y4);
  and_gate and_gate_h_s_arrmul12_and6_1_y0(a_6, b_1, h_s_arrmul12_and6_1_y0);
  fa fa_h_s_arrmul12_fa6_1_y2(h_s_arrmul12_and6_1_y0, h_s_arrmul12_and7_0_y0, h_s_arrmul12_fa5_1_y4, h_s_arrmul12_fa6_1_y2, h_s_arrmul12_fa6_1_y4);
  and_gate and_gate_h_s_arrmul12_and7_1_y0(a_7, b_1, h_s_arrmul12_and7_1_y0);
  fa fa_h_s_arrmul12_fa7_1_y2(h_s_arrmul12_and7_1_y0, h_s_arrmul12_and8_0_y0, h_s_arrmul12_fa6_1_y4, h_s_arrmul12_fa7_1_y2, h_s_arrmul12_fa7_1_y4);
  and_gate and_gate_h_s_arrmul12_and8_1_y0(a_8, b_1, h_s_arrmul12_and8_1_y0);
  fa fa_h_s_arrmul12_fa8_1_y2(h_s_arrmul12_and8_1_y0, h_s_arrmul12_and9_0_y0, h_s_arrmul12_fa7_1_y4, h_s_arrmul12_fa8_1_y2, h_s_arrmul12_fa8_1_y4);
  and_gate and_gate_h_s_arrmul12_and9_1_y0(a_9, b_1, h_s_arrmul12_and9_1_y0);
  fa fa_h_s_arrmul12_fa9_1_y2(h_s_arrmul12_and9_1_y0, h_s_arrmul12_and10_0_y0, h_s_arrmul12_fa8_1_y4, h_s_arrmul12_fa9_1_y2, h_s_arrmul12_fa9_1_y4);
  and_gate and_gate_h_s_arrmul12_and10_1_y0(a_10, b_1, h_s_arrmul12_and10_1_y0);
  fa fa_h_s_arrmul12_fa10_1_y2(h_s_arrmul12_and10_1_y0, h_s_arrmul12_nand11_0_y0, h_s_arrmul12_fa9_1_y4, h_s_arrmul12_fa10_1_y2, h_s_arrmul12_fa10_1_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_1_y0(a_11, b_1, h_s_arrmul12_nand11_1_y0);
  fa fa_h_s_arrmul12_fa11_1_y2(h_s_arrmul12_nand11_1_y0, constant_wire_1, h_s_arrmul12_fa10_1_y4, h_s_arrmul12_fa11_1_y2, h_s_arrmul12_fa11_1_y4);
  and_gate and_gate_h_s_arrmul12_and0_2_y0(a_0, b_2, h_s_arrmul12_and0_2_y0);
  ha ha_h_s_arrmul12_ha0_2_y0(h_s_arrmul12_and0_2_y0, h_s_arrmul12_fa1_1_y2, h_s_arrmul12_ha0_2_y0, h_s_arrmul12_ha0_2_y1);
  and_gate and_gate_h_s_arrmul12_and1_2_y0(a_1, b_2, h_s_arrmul12_and1_2_y0);
  fa fa_h_s_arrmul12_fa1_2_y2(h_s_arrmul12_and1_2_y0, h_s_arrmul12_fa2_1_y2, h_s_arrmul12_ha0_2_y1, h_s_arrmul12_fa1_2_y2, h_s_arrmul12_fa1_2_y4);
  and_gate and_gate_h_s_arrmul12_and2_2_y0(a_2, b_2, h_s_arrmul12_and2_2_y0);
  fa fa_h_s_arrmul12_fa2_2_y2(h_s_arrmul12_and2_2_y0, h_s_arrmul12_fa3_1_y2, h_s_arrmul12_fa1_2_y4, h_s_arrmul12_fa2_2_y2, h_s_arrmul12_fa2_2_y4);
  and_gate and_gate_h_s_arrmul12_and3_2_y0(a_3, b_2, h_s_arrmul12_and3_2_y0);
  fa fa_h_s_arrmul12_fa3_2_y2(h_s_arrmul12_and3_2_y0, h_s_arrmul12_fa4_1_y2, h_s_arrmul12_fa2_2_y4, h_s_arrmul12_fa3_2_y2, h_s_arrmul12_fa3_2_y4);
  and_gate and_gate_h_s_arrmul12_and4_2_y0(a_4, b_2, h_s_arrmul12_and4_2_y0);
  fa fa_h_s_arrmul12_fa4_2_y2(h_s_arrmul12_and4_2_y0, h_s_arrmul12_fa5_1_y2, h_s_arrmul12_fa3_2_y4, h_s_arrmul12_fa4_2_y2, h_s_arrmul12_fa4_2_y4);
  and_gate and_gate_h_s_arrmul12_and5_2_y0(a_5, b_2, h_s_arrmul12_and5_2_y0);
  fa fa_h_s_arrmul12_fa5_2_y2(h_s_arrmul12_and5_2_y0, h_s_arrmul12_fa6_1_y2, h_s_arrmul12_fa4_2_y4, h_s_arrmul12_fa5_2_y2, h_s_arrmul12_fa5_2_y4);
  and_gate and_gate_h_s_arrmul12_and6_2_y0(a_6, b_2, h_s_arrmul12_and6_2_y0);
  fa fa_h_s_arrmul12_fa6_2_y2(h_s_arrmul12_and6_2_y0, h_s_arrmul12_fa7_1_y2, h_s_arrmul12_fa5_2_y4, h_s_arrmul12_fa6_2_y2, h_s_arrmul12_fa6_2_y4);
  and_gate and_gate_h_s_arrmul12_and7_2_y0(a_7, b_2, h_s_arrmul12_and7_2_y0);
  fa fa_h_s_arrmul12_fa7_2_y2(h_s_arrmul12_and7_2_y0, h_s_arrmul12_fa8_1_y2, h_s_arrmul12_fa6_2_y4, h_s_arrmul12_fa7_2_y2, h_s_arrmul12_fa7_2_y4);
  and_gate and_gate_h_s_arrmul12_and8_2_y0(a_8, b_2, h_s_arrmul12_and8_2_y0);
  fa fa_h_s_arrmul12_fa8_2_y2(h_s_arrmul12_and8_2_y0, h_s_arrmul12_fa9_1_y2, h_s_arrmul12_fa7_2_y4, h_s_arrmul12_fa8_2_y2, h_s_arrmul12_fa8_2_y4);
  and_gate and_gate_h_s_arrmul12_and9_2_y0(a_9, b_2, h_s_arrmul12_and9_2_y0);
  fa fa_h_s_arrmul12_fa9_2_y2(h_s_arrmul12_and9_2_y0, h_s_arrmul12_fa10_1_y2, h_s_arrmul12_fa8_2_y4, h_s_arrmul12_fa9_2_y2, h_s_arrmul12_fa9_2_y4);
  and_gate and_gate_h_s_arrmul12_and10_2_y0(a_10, b_2, h_s_arrmul12_and10_2_y0);
  fa fa_h_s_arrmul12_fa10_2_y2(h_s_arrmul12_and10_2_y0, h_s_arrmul12_fa11_1_y2, h_s_arrmul12_fa9_2_y4, h_s_arrmul12_fa10_2_y2, h_s_arrmul12_fa10_2_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_2_y0(a_11, b_2, h_s_arrmul12_nand11_2_y0);
  fa fa_h_s_arrmul12_fa11_2_y2(h_s_arrmul12_nand11_2_y0, h_s_arrmul12_fa11_1_y4, h_s_arrmul12_fa10_2_y4, h_s_arrmul12_fa11_2_y2, h_s_arrmul12_fa11_2_y4);
  and_gate and_gate_h_s_arrmul12_and0_3_y0(a_0, b_3, h_s_arrmul12_and0_3_y0);
  ha ha_h_s_arrmul12_ha0_3_y0(h_s_arrmul12_and0_3_y0, h_s_arrmul12_fa1_2_y2, h_s_arrmul12_ha0_3_y0, h_s_arrmul12_ha0_3_y1);
  and_gate and_gate_h_s_arrmul12_and1_3_y0(a_1, b_3, h_s_arrmul12_and1_3_y0);
  fa fa_h_s_arrmul12_fa1_3_y2(h_s_arrmul12_and1_3_y0, h_s_arrmul12_fa2_2_y2, h_s_arrmul12_ha0_3_y1, h_s_arrmul12_fa1_3_y2, h_s_arrmul12_fa1_3_y4);
  and_gate and_gate_h_s_arrmul12_and2_3_y0(a_2, b_3, h_s_arrmul12_and2_3_y0);
  fa fa_h_s_arrmul12_fa2_3_y2(h_s_arrmul12_and2_3_y0, h_s_arrmul12_fa3_2_y2, h_s_arrmul12_fa1_3_y4, h_s_arrmul12_fa2_3_y2, h_s_arrmul12_fa2_3_y4);
  and_gate and_gate_h_s_arrmul12_and3_3_y0(a_3, b_3, h_s_arrmul12_and3_3_y0);
  fa fa_h_s_arrmul12_fa3_3_y2(h_s_arrmul12_and3_3_y0, h_s_arrmul12_fa4_2_y2, h_s_arrmul12_fa2_3_y4, h_s_arrmul12_fa3_3_y2, h_s_arrmul12_fa3_3_y4);
  and_gate and_gate_h_s_arrmul12_and4_3_y0(a_4, b_3, h_s_arrmul12_and4_3_y0);
  fa fa_h_s_arrmul12_fa4_3_y2(h_s_arrmul12_and4_3_y0, h_s_arrmul12_fa5_2_y2, h_s_arrmul12_fa3_3_y4, h_s_arrmul12_fa4_3_y2, h_s_arrmul12_fa4_3_y4);
  and_gate and_gate_h_s_arrmul12_and5_3_y0(a_5, b_3, h_s_arrmul12_and5_3_y0);
  fa fa_h_s_arrmul12_fa5_3_y2(h_s_arrmul12_and5_3_y0, h_s_arrmul12_fa6_2_y2, h_s_arrmul12_fa4_3_y4, h_s_arrmul12_fa5_3_y2, h_s_arrmul12_fa5_3_y4);
  and_gate and_gate_h_s_arrmul12_and6_3_y0(a_6, b_3, h_s_arrmul12_and6_3_y0);
  fa fa_h_s_arrmul12_fa6_3_y2(h_s_arrmul12_and6_3_y0, h_s_arrmul12_fa7_2_y2, h_s_arrmul12_fa5_3_y4, h_s_arrmul12_fa6_3_y2, h_s_arrmul12_fa6_3_y4);
  and_gate and_gate_h_s_arrmul12_and7_3_y0(a_7, b_3, h_s_arrmul12_and7_3_y0);
  fa fa_h_s_arrmul12_fa7_3_y2(h_s_arrmul12_and7_3_y0, h_s_arrmul12_fa8_2_y2, h_s_arrmul12_fa6_3_y4, h_s_arrmul12_fa7_3_y2, h_s_arrmul12_fa7_3_y4);
  and_gate and_gate_h_s_arrmul12_and8_3_y0(a_8, b_3, h_s_arrmul12_and8_3_y0);
  fa fa_h_s_arrmul12_fa8_3_y2(h_s_arrmul12_and8_3_y0, h_s_arrmul12_fa9_2_y2, h_s_arrmul12_fa7_3_y4, h_s_arrmul12_fa8_3_y2, h_s_arrmul12_fa8_3_y4);
  and_gate and_gate_h_s_arrmul12_and9_3_y0(a_9, b_3, h_s_arrmul12_and9_3_y0);
  fa fa_h_s_arrmul12_fa9_3_y2(h_s_arrmul12_and9_3_y0, h_s_arrmul12_fa10_2_y2, h_s_arrmul12_fa8_3_y4, h_s_arrmul12_fa9_3_y2, h_s_arrmul12_fa9_3_y4);
  and_gate and_gate_h_s_arrmul12_and10_3_y0(a_10, b_3, h_s_arrmul12_and10_3_y0);
  fa fa_h_s_arrmul12_fa10_3_y2(h_s_arrmul12_and10_3_y0, h_s_arrmul12_fa11_2_y2, h_s_arrmul12_fa9_3_y4, h_s_arrmul12_fa10_3_y2, h_s_arrmul12_fa10_3_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_3_y0(a_11, b_3, h_s_arrmul12_nand11_3_y0);
  fa fa_h_s_arrmul12_fa11_3_y2(h_s_arrmul12_nand11_3_y0, h_s_arrmul12_fa11_2_y4, h_s_arrmul12_fa10_3_y4, h_s_arrmul12_fa11_3_y2, h_s_arrmul12_fa11_3_y4);
  and_gate and_gate_h_s_arrmul12_and0_4_y0(a_0, b_4, h_s_arrmul12_and0_4_y0);
  ha ha_h_s_arrmul12_ha0_4_y0(h_s_arrmul12_and0_4_y0, h_s_arrmul12_fa1_3_y2, h_s_arrmul12_ha0_4_y0, h_s_arrmul12_ha0_4_y1);
  and_gate and_gate_h_s_arrmul12_and1_4_y0(a_1, b_4, h_s_arrmul12_and1_4_y0);
  fa fa_h_s_arrmul12_fa1_4_y2(h_s_arrmul12_and1_4_y0, h_s_arrmul12_fa2_3_y2, h_s_arrmul12_ha0_4_y1, h_s_arrmul12_fa1_4_y2, h_s_arrmul12_fa1_4_y4);
  and_gate and_gate_h_s_arrmul12_and2_4_y0(a_2, b_4, h_s_arrmul12_and2_4_y0);
  fa fa_h_s_arrmul12_fa2_4_y2(h_s_arrmul12_and2_4_y0, h_s_arrmul12_fa3_3_y2, h_s_arrmul12_fa1_4_y4, h_s_arrmul12_fa2_4_y2, h_s_arrmul12_fa2_4_y4);
  and_gate and_gate_h_s_arrmul12_and3_4_y0(a_3, b_4, h_s_arrmul12_and3_4_y0);
  fa fa_h_s_arrmul12_fa3_4_y2(h_s_arrmul12_and3_4_y0, h_s_arrmul12_fa4_3_y2, h_s_arrmul12_fa2_4_y4, h_s_arrmul12_fa3_4_y2, h_s_arrmul12_fa3_4_y4);
  and_gate and_gate_h_s_arrmul12_and4_4_y0(a_4, b_4, h_s_arrmul12_and4_4_y0);
  fa fa_h_s_arrmul12_fa4_4_y2(h_s_arrmul12_and4_4_y0, h_s_arrmul12_fa5_3_y2, h_s_arrmul12_fa3_4_y4, h_s_arrmul12_fa4_4_y2, h_s_arrmul12_fa4_4_y4);
  and_gate and_gate_h_s_arrmul12_and5_4_y0(a_5, b_4, h_s_arrmul12_and5_4_y0);
  fa fa_h_s_arrmul12_fa5_4_y2(h_s_arrmul12_and5_4_y0, h_s_arrmul12_fa6_3_y2, h_s_arrmul12_fa4_4_y4, h_s_arrmul12_fa5_4_y2, h_s_arrmul12_fa5_4_y4);
  and_gate and_gate_h_s_arrmul12_and6_4_y0(a_6, b_4, h_s_arrmul12_and6_4_y0);
  fa fa_h_s_arrmul12_fa6_4_y2(h_s_arrmul12_and6_4_y0, h_s_arrmul12_fa7_3_y2, h_s_arrmul12_fa5_4_y4, h_s_arrmul12_fa6_4_y2, h_s_arrmul12_fa6_4_y4);
  and_gate and_gate_h_s_arrmul12_and7_4_y0(a_7, b_4, h_s_arrmul12_and7_4_y0);
  fa fa_h_s_arrmul12_fa7_4_y2(h_s_arrmul12_and7_4_y0, h_s_arrmul12_fa8_3_y2, h_s_arrmul12_fa6_4_y4, h_s_arrmul12_fa7_4_y2, h_s_arrmul12_fa7_4_y4);
  and_gate and_gate_h_s_arrmul12_and8_4_y0(a_8, b_4, h_s_arrmul12_and8_4_y0);
  fa fa_h_s_arrmul12_fa8_4_y2(h_s_arrmul12_and8_4_y0, h_s_arrmul12_fa9_3_y2, h_s_arrmul12_fa7_4_y4, h_s_arrmul12_fa8_4_y2, h_s_arrmul12_fa8_4_y4);
  and_gate and_gate_h_s_arrmul12_and9_4_y0(a_9, b_4, h_s_arrmul12_and9_4_y0);
  fa fa_h_s_arrmul12_fa9_4_y2(h_s_arrmul12_and9_4_y0, h_s_arrmul12_fa10_3_y2, h_s_arrmul12_fa8_4_y4, h_s_arrmul12_fa9_4_y2, h_s_arrmul12_fa9_4_y4);
  and_gate and_gate_h_s_arrmul12_and10_4_y0(a_10, b_4, h_s_arrmul12_and10_4_y0);
  fa fa_h_s_arrmul12_fa10_4_y2(h_s_arrmul12_and10_4_y0, h_s_arrmul12_fa11_3_y2, h_s_arrmul12_fa9_4_y4, h_s_arrmul12_fa10_4_y2, h_s_arrmul12_fa10_4_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_4_y0(a_11, b_4, h_s_arrmul12_nand11_4_y0);
  fa fa_h_s_arrmul12_fa11_4_y2(h_s_arrmul12_nand11_4_y0, h_s_arrmul12_fa11_3_y4, h_s_arrmul12_fa10_4_y4, h_s_arrmul12_fa11_4_y2, h_s_arrmul12_fa11_4_y4);
  and_gate and_gate_h_s_arrmul12_and0_5_y0(a_0, b_5, h_s_arrmul12_and0_5_y0);
  ha ha_h_s_arrmul12_ha0_5_y0(h_s_arrmul12_and0_5_y0, h_s_arrmul12_fa1_4_y2, h_s_arrmul12_ha0_5_y0, h_s_arrmul12_ha0_5_y1);
  and_gate and_gate_h_s_arrmul12_and1_5_y0(a_1, b_5, h_s_arrmul12_and1_5_y0);
  fa fa_h_s_arrmul12_fa1_5_y2(h_s_arrmul12_and1_5_y0, h_s_arrmul12_fa2_4_y2, h_s_arrmul12_ha0_5_y1, h_s_arrmul12_fa1_5_y2, h_s_arrmul12_fa1_5_y4);
  and_gate and_gate_h_s_arrmul12_and2_5_y0(a_2, b_5, h_s_arrmul12_and2_5_y0);
  fa fa_h_s_arrmul12_fa2_5_y2(h_s_arrmul12_and2_5_y0, h_s_arrmul12_fa3_4_y2, h_s_arrmul12_fa1_5_y4, h_s_arrmul12_fa2_5_y2, h_s_arrmul12_fa2_5_y4);
  and_gate and_gate_h_s_arrmul12_and3_5_y0(a_3, b_5, h_s_arrmul12_and3_5_y0);
  fa fa_h_s_arrmul12_fa3_5_y2(h_s_arrmul12_and3_5_y0, h_s_arrmul12_fa4_4_y2, h_s_arrmul12_fa2_5_y4, h_s_arrmul12_fa3_5_y2, h_s_arrmul12_fa3_5_y4);
  and_gate and_gate_h_s_arrmul12_and4_5_y0(a_4, b_5, h_s_arrmul12_and4_5_y0);
  fa fa_h_s_arrmul12_fa4_5_y2(h_s_arrmul12_and4_5_y0, h_s_arrmul12_fa5_4_y2, h_s_arrmul12_fa3_5_y4, h_s_arrmul12_fa4_5_y2, h_s_arrmul12_fa4_5_y4);
  and_gate and_gate_h_s_arrmul12_and5_5_y0(a_5, b_5, h_s_arrmul12_and5_5_y0);
  fa fa_h_s_arrmul12_fa5_5_y2(h_s_arrmul12_and5_5_y0, h_s_arrmul12_fa6_4_y2, h_s_arrmul12_fa4_5_y4, h_s_arrmul12_fa5_5_y2, h_s_arrmul12_fa5_5_y4);
  and_gate and_gate_h_s_arrmul12_and6_5_y0(a_6, b_5, h_s_arrmul12_and6_5_y0);
  fa fa_h_s_arrmul12_fa6_5_y2(h_s_arrmul12_and6_5_y0, h_s_arrmul12_fa7_4_y2, h_s_arrmul12_fa5_5_y4, h_s_arrmul12_fa6_5_y2, h_s_arrmul12_fa6_5_y4);
  and_gate and_gate_h_s_arrmul12_and7_5_y0(a_7, b_5, h_s_arrmul12_and7_5_y0);
  fa fa_h_s_arrmul12_fa7_5_y2(h_s_arrmul12_and7_5_y0, h_s_arrmul12_fa8_4_y2, h_s_arrmul12_fa6_5_y4, h_s_arrmul12_fa7_5_y2, h_s_arrmul12_fa7_5_y4);
  and_gate and_gate_h_s_arrmul12_and8_5_y0(a_8, b_5, h_s_arrmul12_and8_5_y0);
  fa fa_h_s_arrmul12_fa8_5_y2(h_s_arrmul12_and8_5_y0, h_s_arrmul12_fa9_4_y2, h_s_arrmul12_fa7_5_y4, h_s_arrmul12_fa8_5_y2, h_s_arrmul12_fa8_5_y4);
  and_gate and_gate_h_s_arrmul12_and9_5_y0(a_9, b_5, h_s_arrmul12_and9_5_y0);
  fa fa_h_s_arrmul12_fa9_5_y2(h_s_arrmul12_and9_5_y0, h_s_arrmul12_fa10_4_y2, h_s_arrmul12_fa8_5_y4, h_s_arrmul12_fa9_5_y2, h_s_arrmul12_fa9_5_y4);
  and_gate and_gate_h_s_arrmul12_and10_5_y0(a_10, b_5, h_s_arrmul12_and10_5_y0);
  fa fa_h_s_arrmul12_fa10_5_y2(h_s_arrmul12_and10_5_y0, h_s_arrmul12_fa11_4_y2, h_s_arrmul12_fa9_5_y4, h_s_arrmul12_fa10_5_y2, h_s_arrmul12_fa10_5_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_5_y0(a_11, b_5, h_s_arrmul12_nand11_5_y0);
  fa fa_h_s_arrmul12_fa11_5_y2(h_s_arrmul12_nand11_5_y0, h_s_arrmul12_fa11_4_y4, h_s_arrmul12_fa10_5_y4, h_s_arrmul12_fa11_5_y2, h_s_arrmul12_fa11_5_y4);
  and_gate and_gate_h_s_arrmul12_and0_6_y0(a_0, b_6, h_s_arrmul12_and0_6_y0);
  ha ha_h_s_arrmul12_ha0_6_y0(h_s_arrmul12_and0_6_y0, h_s_arrmul12_fa1_5_y2, h_s_arrmul12_ha0_6_y0, h_s_arrmul12_ha0_6_y1);
  and_gate and_gate_h_s_arrmul12_and1_6_y0(a_1, b_6, h_s_arrmul12_and1_6_y0);
  fa fa_h_s_arrmul12_fa1_6_y2(h_s_arrmul12_and1_6_y0, h_s_arrmul12_fa2_5_y2, h_s_arrmul12_ha0_6_y1, h_s_arrmul12_fa1_6_y2, h_s_arrmul12_fa1_6_y4);
  and_gate and_gate_h_s_arrmul12_and2_6_y0(a_2, b_6, h_s_arrmul12_and2_6_y0);
  fa fa_h_s_arrmul12_fa2_6_y2(h_s_arrmul12_and2_6_y0, h_s_arrmul12_fa3_5_y2, h_s_arrmul12_fa1_6_y4, h_s_arrmul12_fa2_6_y2, h_s_arrmul12_fa2_6_y4);
  and_gate and_gate_h_s_arrmul12_and3_6_y0(a_3, b_6, h_s_arrmul12_and3_6_y0);
  fa fa_h_s_arrmul12_fa3_6_y2(h_s_arrmul12_and3_6_y0, h_s_arrmul12_fa4_5_y2, h_s_arrmul12_fa2_6_y4, h_s_arrmul12_fa3_6_y2, h_s_arrmul12_fa3_6_y4);
  and_gate and_gate_h_s_arrmul12_and4_6_y0(a_4, b_6, h_s_arrmul12_and4_6_y0);
  fa fa_h_s_arrmul12_fa4_6_y2(h_s_arrmul12_and4_6_y0, h_s_arrmul12_fa5_5_y2, h_s_arrmul12_fa3_6_y4, h_s_arrmul12_fa4_6_y2, h_s_arrmul12_fa4_6_y4);
  and_gate and_gate_h_s_arrmul12_and5_6_y0(a_5, b_6, h_s_arrmul12_and5_6_y0);
  fa fa_h_s_arrmul12_fa5_6_y2(h_s_arrmul12_and5_6_y0, h_s_arrmul12_fa6_5_y2, h_s_arrmul12_fa4_6_y4, h_s_arrmul12_fa5_6_y2, h_s_arrmul12_fa5_6_y4);
  and_gate and_gate_h_s_arrmul12_and6_6_y0(a_6, b_6, h_s_arrmul12_and6_6_y0);
  fa fa_h_s_arrmul12_fa6_6_y2(h_s_arrmul12_and6_6_y0, h_s_arrmul12_fa7_5_y2, h_s_arrmul12_fa5_6_y4, h_s_arrmul12_fa6_6_y2, h_s_arrmul12_fa6_6_y4);
  and_gate and_gate_h_s_arrmul12_and7_6_y0(a_7, b_6, h_s_arrmul12_and7_6_y0);
  fa fa_h_s_arrmul12_fa7_6_y2(h_s_arrmul12_and7_6_y0, h_s_arrmul12_fa8_5_y2, h_s_arrmul12_fa6_6_y4, h_s_arrmul12_fa7_6_y2, h_s_arrmul12_fa7_6_y4);
  and_gate and_gate_h_s_arrmul12_and8_6_y0(a_8, b_6, h_s_arrmul12_and8_6_y0);
  fa fa_h_s_arrmul12_fa8_6_y2(h_s_arrmul12_and8_6_y0, h_s_arrmul12_fa9_5_y2, h_s_arrmul12_fa7_6_y4, h_s_arrmul12_fa8_6_y2, h_s_arrmul12_fa8_6_y4);
  and_gate and_gate_h_s_arrmul12_and9_6_y0(a_9, b_6, h_s_arrmul12_and9_6_y0);
  fa fa_h_s_arrmul12_fa9_6_y2(h_s_arrmul12_and9_6_y0, h_s_arrmul12_fa10_5_y2, h_s_arrmul12_fa8_6_y4, h_s_arrmul12_fa9_6_y2, h_s_arrmul12_fa9_6_y4);
  and_gate and_gate_h_s_arrmul12_and10_6_y0(a_10, b_6, h_s_arrmul12_and10_6_y0);
  fa fa_h_s_arrmul12_fa10_6_y2(h_s_arrmul12_and10_6_y0, h_s_arrmul12_fa11_5_y2, h_s_arrmul12_fa9_6_y4, h_s_arrmul12_fa10_6_y2, h_s_arrmul12_fa10_6_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_6_y0(a_11, b_6, h_s_arrmul12_nand11_6_y0);
  fa fa_h_s_arrmul12_fa11_6_y2(h_s_arrmul12_nand11_6_y0, h_s_arrmul12_fa11_5_y4, h_s_arrmul12_fa10_6_y4, h_s_arrmul12_fa11_6_y2, h_s_arrmul12_fa11_6_y4);
  and_gate and_gate_h_s_arrmul12_and0_7_y0(a_0, b_7, h_s_arrmul12_and0_7_y0);
  ha ha_h_s_arrmul12_ha0_7_y0(h_s_arrmul12_and0_7_y0, h_s_arrmul12_fa1_6_y2, h_s_arrmul12_ha0_7_y0, h_s_arrmul12_ha0_7_y1);
  and_gate and_gate_h_s_arrmul12_and1_7_y0(a_1, b_7, h_s_arrmul12_and1_7_y0);
  fa fa_h_s_arrmul12_fa1_7_y2(h_s_arrmul12_and1_7_y0, h_s_arrmul12_fa2_6_y2, h_s_arrmul12_ha0_7_y1, h_s_arrmul12_fa1_7_y2, h_s_arrmul12_fa1_7_y4);
  and_gate and_gate_h_s_arrmul12_and2_7_y0(a_2, b_7, h_s_arrmul12_and2_7_y0);
  fa fa_h_s_arrmul12_fa2_7_y2(h_s_arrmul12_and2_7_y0, h_s_arrmul12_fa3_6_y2, h_s_arrmul12_fa1_7_y4, h_s_arrmul12_fa2_7_y2, h_s_arrmul12_fa2_7_y4);
  and_gate and_gate_h_s_arrmul12_and3_7_y0(a_3, b_7, h_s_arrmul12_and3_7_y0);
  fa fa_h_s_arrmul12_fa3_7_y2(h_s_arrmul12_and3_7_y0, h_s_arrmul12_fa4_6_y2, h_s_arrmul12_fa2_7_y4, h_s_arrmul12_fa3_7_y2, h_s_arrmul12_fa3_7_y4);
  and_gate and_gate_h_s_arrmul12_and4_7_y0(a_4, b_7, h_s_arrmul12_and4_7_y0);
  fa fa_h_s_arrmul12_fa4_7_y2(h_s_arrmul12_and4_7_y0, h_s_arrmul12_fa5_6_y2, h_s_arrmul12_fa3_7_y4, h_s_arrmul12_fa4_7_y2, h_s_arrmul12_fa4_7_y4);
  and_gate and_gate_h_s_arrmul12_and5_7_y0(a_5, b_7, h_s_arrmul12_and5_7_y0);
  fa fa_h_s_arrmul12_fa5_7_y2(h_s_arrmul12_and5_7_y0, h_s_arrmul12_fa6_6_y2, h_s_arrmul12_fa4_7_y4, h_s_arrmul12_fa5_7_y2, h_s_arrmul12_fa5_7_y4);
  and_gate and_gate_h_s_arrmul12_and6_7_y0(a_6, b_7, h_s_arrmul12_and6_7_y0);
  fa fa_h_s_arrmul12_fa6_7_y2(h_s_arrmul12_and6_7_y0, h_s_arrmul12_fa7_6_y2, h_s_arrmul12_fa5_7_y4, h_s_arrmul12_fa6_7_y2, h_s_arrmul12_fa6_7_y4);
  and_gate and_gate_h_s_arrmul12_and7_7_y0(a_7, b_7, h_s_arrmul12_and7_7_y0);
  fa fa_h_s_arrmul12_fa7_7_y2(h_s_arrmul12_and7_7_y0, h_s_arrmul12_fa8_6_y2, h_s_arrmul12_fa6_7_y4, h_s_arrmul12_fa7_7_y2, h_s_arrmul12_fa7_7_y4);
  and_gate and_gate_h_s_arrmul12_and8_7_y0(a_8, b_7, h_s_arrmul12_and8_7_y0);
  fa fa_h_s_arrmul12_fa8_7_y2(h_s_arrmul12_and8_7_y0, h_s_arrmul12_fa9_6_y2, h_s_arrmul12_fa7_7_y4, h_s_arrmul12_fa8_7_y2, h_s_arrmul12_fa8_7_y4);
  and_gate and_gate_h_s_arrmul12_and9_7_y0(a_9, b_7, h_s_arrmul12_and9_7_y0);
  fa fa_h_s_arrmul12_fa9_7_y2(h_s_arrmul12_and9_7_y0, h_s_arrmul12_fa10_6_y2, h_s_arrmul12_fa8_7_y4, h_s_arrmul12_fa9_7_y2, h_s_arrmul12_fa9_7_y4);
  and_gate and_gate_h_s_arrmul12_and10_7_y0(a_10, b_7, h_s_arrmul12_and10_7_y0);
  fa fa_h_s_arrmul12_fa10_7_y2(h_s_arrmul12_and10_7_y0, h_s_arrmul12_fa11_6_y2, h_s_arrmul12_fa9_7_y4, h_s_arrmul12_fa10_7_y2, h_s_arrmul12_fa10_7_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_7_y0(a_11, b_7, h_s_arrmul12_nand11_7_y0);
  fa fa_h_s_arrmul12_fa11_7_y2(h_s_arrmul12_nand11_7_y0, h_s_arrmul12_fa11_6_y4, h_s_arrmul12_fa10_7_y4, h_s_arrmul12_fa11_7_y2, h_s_arrmul12_fa11_7_y4);
  and_gate and_gate_h_s_arrmul12_and0_8_y0(a_0, b_8, h_s_arrmul12_and0_8_y0);
  ha ha_h_s_arrmul12_ha0_8_y0(h_s_arrmul12_and0_8_y0, h_s_arrmul12_fa1_7_y2, h_s_arrmul12_ha0_8_y0, h_s_arrmul12_ha0_8_y1);
  and_gate and_gate_h_s_arrmul12_and1_8_y0(a_1, b_8, h_s_arrmul12_and1_8_y0);
  fa fa_h_s_arrmul12_fa1_8_y2(h_s_arrmul12_and1_8_y0, h_s_arrmul12_fa2_7_y2, h_s_arrmul12_ha0_8_y1, h_s_arrmul12_fa1_8_y2, h_s_arrmul12_fa1_8_y4);
  and_gate and_gate_h_s_arrmul12_and2_8_y0(a_2, b_8, h_s_arrmul12_and2_8_y0);
  fa fa_h_s_arrmul12_fa2_8_y2(h_s_arrmul12_and2_8_y0, h_s_arrmul12_fa3_7_y2, h_s_arrmul12_fa1_8_y4, h_s_arrmul12_fa2_8_y2, h_s_arrmul12_fa2_8_y4);
  and_gate and_gate_h_s_arrmul12_and3_8_y0(a_3, b_8, h_s_arrmul12_and3_8_y0);
  fa fa_h_s_arrmul12_fa3_8_y2(h_s_arrmul12_and3_8_y0, h_s_arrmul12_fa4_7_y2, h_s_arrmul12_fa2_8_y4, h_s_arrmul12_fa3_8_y2, h_s_arrmul12_fa3_8_y4);
  and_gate and_gate_h_s_arrmul12_and4_8_y0(a_4, b_8, h_s_arrmul12_and4_8_y0);
  fa fa_h_s_arrmul12_fa4_8_y2(h_s_arrmul12_and4_8_y0, h_s_arrmul12_fa5_7_y2, h_s_arrmul12_fa3_8_y4, h_s_arrmul12_fa4_8_y2, h_s_arrmul12_fa4_8_y4);
  and_gate and_gate_h_s_arrmul12_and5_8_y0(a_5, b_8, h_s_arrmul12_and5_8_y0);
  fa fa_h_s_arrmul12_fa5_8_y2(h_s_arrmul12_and5_8_y0, h_s_arrmul12_fa6_7_y2, h_s_arrmul12_fa4_8_y4, h_s_arrmul12_fa5_8_y2, h_s_arrmul12_fa5_8_y4);
  and_gate and_gate_h_s_arrmul12_and6_8_y0(a_6, b_8, h_s_arrmul12_and6_8_y0);
  fa fa_h_s_arrmul12_fa6_8_y2(h_s_arrmul12_and6_8_y0, h_s_arrmul12_fa7_7_y2, h_s_arrmul12_fa5_8_y4, h_s_arrmul12_fa6_8_y2, h_s_arrmul12_fa6_8_y4);
  and_gate and_gate_h_s_arrmul12_and7_8_y0(a_7, b_8, h_s_arrmul12_and7_8_y0);
  fa fa_h_s_arrmul12_fa7_8_y2(h_s_arrmul12_and7_8_y0, h_s_arrmul12_fa8_7_y2, h_s_arrmul12_fa6_8_y4, h_s_arrmul12_fa7_8_y2, h_s_arrmul12_fa7_8_y4);
  and_gate and_gate_h_s_arrmul12_and8_8_y0(a_8, b_8, h_s_arrmul12_and8_8_y0);
  fa fa_h_s_arrmul12_fa8_8_y2(h_s_arrmul12_and8_8_y0, h_s_arrmul12_fa9_7_y2, h_s_arrmul12_fa7_8_y4, h_s_arrmul12_fa8_8_y2, h_s_arrmul12_fa8_8_y4);
  and_gate and_gate_h_s_arrmul12_and9_8_y0(a_9, b_8, h_s_arrmul12_and9_8_y0);
  fa fa_h_s_arrmul12_fa9_8_y2(h_s_arrmul12_and9_8_y0, h_s_arrmul12_fa10_7_y2, h_s_arrmul12_fa8_8_y4, h_s_arrmul12_fa9_8_y2, h_s_arrmul12_fa9_8_y4);
  and_gate and_gate_h_s_arrmul12_and10_8_y0(a_10, b_8, h_s_arrmul12_and10_8_y0);
  fa fa_h_s_arrmul12_fa10_8_y2(h_s_arrmul12_and10_8_y0, h_s_arrmul12_fa11_7_y2, h_s_arrmul12_fa9_8_y4, h_s_arrmul12_fa10_8_y2, h_s_arrmul12_fa10_8_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_8_y0(a_11, b_8, h_s_arrmul12_nand11_8_y0);
  fa fa_h_s_arrmul12_fa11_8_y2(h_s_arrmul12_nand11_8_y0, h_s_arrmul12_fa11_7_y4, h_s_arrmul12_fa10_8_y4, h_s_arrmul12_fa11_8_y2, h_s_arrmul12_fa11_8_y4);
  and_gate and_gate_h_s_arrmul12_and0_9_y0(a_0, b_9, h_s_arrmul12_and0_9_y0);
  ha ha_h_s_arrmul12_ha0_9_y0(h_s_arrmul12_and0_9_y0, h_s_arrmul12_fa1_8_y2, h_s_arrmul12_ha0_9_y0, h_s_arrmul12_ha0_9_y1);
  and_gate and_gate_h_s_arrmul12_and1_9_y0(a_1, b_9, h_s_arrmul12_and1_9_y0);
  fa fa_h_s_arrmul12_fa1_9_y2(h_s_arrmul12_and1_9_y0, h_s_arrmul12_fa2_8_y2, h_s_arrmul12_ha0_9_y1, h_s_arrmul12_fa1_9_y2, h_s_arrmul12_fa1_9_y4);
  and_gate and_gate_h_s_arrmul12_and2_9_y0(a_2, b_9, h_s_arrmul12_and2_9_y0);
  fa fa_h_s_arrmul12_fa2_9_y2(h_s_arrmul12_and2_9_y0, h_s_arrmul12_fa3_8_y2, h_s_arrmul12_fa1_9_y4, h_s_arrmul12_fa2_9_y2, h_s_arrmul12_fa2_9_y4);
  and_gate and_gate_h_s_arrmul12_and3_9_y0(a_3, b_9, h_s_arrmul12_and3_9_y0);
  fa fa_h_s_arrmul12_fa3_9_y2(h_s_arrmul12_and3_9_y0, h_s_arrmul12_fa4_8_y2, h_s_arrmul12_fa2_9_y4, h_s_arrmul12_fa3_9_y2, h_s_arrmul12_fa3_9_y4);
  and_gate and_gate_h_s_arrmul12_and4_9_y0(a_4, b_9, h_s_arrmul12_and4_9_y0);
  fa fa_h_s_arrmul12_fa4_9_y2(h_s_arrmul12_and4_9_y0, h_s_arrmul12_fa5_8_y2, h_s_arrmul12_fa3_9_y4, h_s_arrmul12_fa4_9_y2, h_s_arrmul12_fa4_9_y4);
  and_gate and_gate_h_s_arrmul12_and5_9_y0(a_5, b_9, h_s_arrmul12_and5_9_y0);
  fa fa_h_s_arrmul12_fa5_9_y2(h_s_arrmul12_and5_9_y0, h_s_arrmul12_fa6_8_y2, h_s_arrmul12_fa4_9_y4, h_s_arrmul12_fa5_9_y2, h_s_arrmul12_fa5_9_y4);
  and_gate and_gate_h_s_arrmul12_and6_9_y0(a_6, b_9, h_s_arrmul12_and6_9_y0);
  fa fa_h_s_arrmul12_fa6_9_y2(h_s_arrmul12_and6_9_y0, h_s_arrmul12_fa7_8_y2, h_s_arrmul12_fa5_9_y4, h_s_arrmul12_fa6_9_y2, h_s_arrmul12_fa6_9_y4);
  and_gate and_gate_h_s_arrmul12_and7_9_y0(a_7, b_9, h_s_arrmul12_and7_9_y0);
  fa fa_h_s_arrmul12_fa7_9_y2(h_s_arrmul12_and7_9_y0, h_s_arrmul12_fa8_8_y2, h_s_arrmul12_fa6_9_y4, h_s_arrmul12_fa7_9_y2, h_s_arrmul12_fa7_9_y4);
  and_gate and_gate_h_s_arrmul12_and8_9_y0(a_8, b_9, h_s_arrmul12_and8_9_y0);
  fa fa_h_s_arrmul12_fa8_9_y2(h_s_arrmul12_and8_9_y0, h_s_arrmul12_fa9_8_y2, h_s_arrmul12_fa7_9_y4, h_s_arrmul12_fa8_9_y2, h_s_arrmul12_fa8_9_y4);
  and_gate and_gate_h_s_arrmul12_and9_9_y0(a_9, b_9, h_s_arrmul12_and9_9_y0);
  fa fa_h_s_arrmul12_fa9_9_y2(h_s_arrmul12_and9_9_y0, h_s_arrmul12_fa10_8_y2, h_s_arrmul12_fa8_9_y4, h_s_arrmul12_fa9_9_y2, h_s_arrmul12_fa9_9_y4);
  and_gate and_gate_h_s_arrmul12_and10_9_y0(a_10, b_9, h_s_arrmul12_and10_9_y0);
  fa fa_h_s_arrmul12_fa10_9_y2(h_s_arrmul12_and10_9_y0, h_s_arrmul12_fa11_8_y2, h_s_arrmul12_fa9_9_y4, h_s_arrmul12_fa10_9_y2, h_s_arrmul12_fa10_9_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_9_y0(a_11, b_9, h_s_arrmul12_nand11_9_y0);
  fa fa_h_s_arrmul12_fa11_9_y2(h_s_arrmul12_nand11_9_y0, h_s_arrmul12_fa11_8_y4, h_s_arrmul12_fa10_9_y4, h_s_arrmul12_fa11_9_y2, h_s_arrmul12_fa11_9_y4);
  and_gate and_gate_h_s_arrmul12_and0_10_y0(a_0, b_10, h_s_arrmul12_and0_10_y0);
  ha ha_h_s_arrmul12_ha0_10_y0(h_s_arrmul12_and0_10_y0, h_s_arrmul12_fa1_9_y2, h_s_arrmul12_ha0_10_y0, h_s_arrmul12_ha0_10_y1);
  and_gate and_gate_h_s_arrmul12_and1_10_y0(a_1, b_10, h_s_arrmul12_and1_10_y0);
  fa fa_h_s_arrmul12_fa1_10_y2(h_s_arrmul12_and1_10_y0, h_s_arrmul12_fa2_9_y2, h_s_arrmul12_ha0_10_y1, h_s_arrmul12_fa1_10_y2, h_s_arrmul12_fa1_10_y4);
  and_gate and_gate_h_s_arrmul12_and2_10_y0(a_2, b_10, h_s_arrmul12_and2_10_y0);
  fa fa_h_s_arrmul12_fa2_10_y2(h_s_arrmul12_and2_10_y0, h_s_arrmul12_fa3_9_y2, h_s_arrmul12_fa1_10_y4, h_s_arrmul12_fa2_10_y2, h_s_arrmul12_fa2_10_y4);
  and_gate and_gate_h_s_arrmul12_and3_10_y0(a_3, b_10, h_s_arrmul12_and3_10_y0);
  fa fa_h_s_arrmul12_fa3_10_y2(h_s_arrmul12_and3_10_y0, h_s_arrmul12_fa4_9_y2, h_s_arrmul12_fa2_10_y4, h_s_arrmul12_fa3_10_y2, h_s_arrmul12_fa3_10_y4);
  and_gate and_gate_h_s_arrmul12_and4_10_y0(a_4, b_10, h_s_arrmul12_and4_10_y0);
  fa fa_h_s_arrmul12_fa4_10_y2(h_s_arrmul12_and4_10_y0, h_s_arrmul12_fa5_9_y2, h_s_arrmul12_fa3_10_y4, h_s_arrmul12_fa4_10_y2, h_s_arrmul12_fa4_10_y4);
  and_gate and_gate_h_s_arrmul12_and5_10_y0(a_5, b_10, h_s_arrmul12_and5_10_y0);
  fa fa_h_s_arrmul12_fa5_10_y2(h_s_arrmul12_and5_10_y0, h_s_arrmul12_fa6_9_y2, h_s_arrmul12_fa4_10_y4, h_s_arrmul12_fa5_10_y2, h_s_arrmul12_fa5_10_y4);
  and_gate and_gate_h_s_arrmul12_and6_10_y0(a_6, b_10, h_s_arrmul12_and6_10_y0);
  fa fa_h_s_arrmul12_fa6_10_y2(h_s_arrmul12_and6_10_y0, h_s_arrmul12_fa7_9_y2, h_s_arrmul12_fa5_10_y4, h_s_arrmul12_fa6_10_y2, h_s_arrmul12_fa6_10_y4);
  and_gate and_gate_h_s_arrmul12_and7_10_y0(a_7, b_10, h_s_arrmul12_and7_10_y0);
  fa fa_h_s_arrmul12_fa7_10_y2(h_s_arrmul12_and7_10_y0, h_s_arrmul12_fa8_9_y2, h_s_arrmul12_fa6_10_y4, h_s_arrmul12_fa7_10_y2, h_s_arrmul12_fa7_10_y4);
  and_gate and_gate_h_s_arrmul12_and8_10_y0(a_8, b_10, h_s_arrmul12_and8_10_y0);
  fa fa_h_s_arrmul12_fa8_10_y2(h_s_arrmul12_and8_10_y0, h_s_arrmul12_fa9_9_y2, h_s_arrmul12_fa7_10_y4, h_s_arrmul12_fa8_10_y2, h_s_arrmul12_fa8_10_y4);
  and_gate and_gate_h_s_arrmul12_and9_10_y0(a_9, b_10, h_s_arrmul12_and9_10_y0);
  fa fa_h_s_arrmul12_fa9_10_y2(h_s_arrmul12_and9_10_y0, h_s_arrmul12_fa10_9_y2, h_s_arrmul12_fa8_10_y4, h_s_arrmul12_fa9_10_y2, h_s_arrmul12_fa9_10_y4);
  and_gate and_gate_h_s_arrmul12_and10_10_y0(a_10, b_10, h_s_arrmul12_and10_10_y0);
  fa fa_h_s_arrmul12_fa10_10_y2(h_s_arrmul12_and10_10_y0, h_s_arrmul12_fa11_9_y2, h_s_arrmul12_fa9_10_y4, h_s_arrmul12_fa10_10_y2, h_s_arrmul12_fa10_10_y4);
  nand_gate nand_gate_h_s_arrmul12_nand11_10_y0(a_11, b_10, h_s_arrmul12_nand11_10_y0);
  fa fa_h_s_arrmul12_fa11_10_y2(h_s_arrmul12_nand11_10_y0, h_s_arrmul12_fa11_9_y4, h_s_arrmul12_fa10_10_y4, h_s_arrmul12_fa11_10_y2, h_s_arrmul12_fa11_10_y4);
  nand_gate nand_gate_h_s_arrmul12_nand0_11_y0(a_0, b_11, h_s_arrmul12_nand0_11_y0);
  ha ha_h_s_arrmul12_ha0_11_y0(h_s_arrmul12_nand0_11_y0, h_s_arrmul12_fa1_10_y2, h_s_arrmul12_ha0_11_y0, h_s_arrmul12_ha0_11_y1);
  nand_gate nand_gate_h_s_arrmul12_nand1_11_y0(a_1, b_11, h_s_arrmul12_nand1_11_y0);
  fa fa_h_s_arrmul12_fa1_11_y2(h_s_arrmul12_nand1_11_y0, h_s_arrmul12_fa2_10_y2, h_s_arrmul12_ha0_11_y1, h_s_arrmul12_fa1_11_y2, h_s_arrmul12_fa1_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand2_11_y0(a_2, b_11, h_s_arrmul12_nand2_11_y0);
  fa fa_h_s_arrmul12_fa2_11_y2(h_s_arrmul12_nand2_11_y0, h_s_arrmul12_fa3_10_y2, h_s_arrmul12_fa1_11_y4, h_s_arrmul12_fa2_11_y2, h_s_arrmul12_fa2_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand3_11_y0(a_3, b_11, h_s_arrmul12_nand3_11_y0);
  fa fa_h_s_arrmul12_fa3_11_y2(h_s_arrmul12_nand3_11_y0, h_s_arrmul12_fa4_10_y2, h_s_arrmul12_fa2_11_y4, h_s_arrmul12_fa3_11_y2, h_s_arrmul12_fa3_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand4_11_y0(a_4, b_11, h_s_arrmul12_nand4_11_y0);
  fa fa_h_s_arrmul12_fa4_11_y2(h_s_arrmul12_nand4_11_y0, h_s_arrmul12_fa5_10_y2, h_s_arrmul12_fa3_11_y4, h_s_arrmul12_fa4_11_y2, h_s_arrmul12_fa4_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand5_11_y0(a_5, b_11, h_s_arrmul12_nand5_11_y0);
  fa fa_h_s_arrmul12_fa5_11_y2(h_s_arrmul12_nand5_11_y0, h_s_arrmul12_fa6_10_y2, h_s_arrmul12_fa4_11_y4, h_s_arrmul12_fa5_11_y2, h_s_arrmul12_fa5_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand6_11_y0(a_6, b_11, h_s_arrmul12_nand6_11_y0);
  fa fa_h_s_arrmul12_fa6_11_y2(h_s_arrmul12_nand6_11_y0, h_s_arrmul12_fa7_10_y2, h_s_arrmul12_fa5_11_y4, h_s_arrmul12_fa6_11_y2, h_s_arrmul12_fa6_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand7_11_y0(a_7, b_11, h_s_arrmul12_nand7_11_y0);
  fa fa_h_s_arrmul12_fa7_11_y2(h_s_arrmul12_nand7_11_y0, h_s_arrmul12_fa8_10_y2, h_s_arrmul12_fa6_11_y4, h_s_arrmul12_fa7_11_y2, h_s_arrmul12_fa7_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand8_11_y0(a_8, b_11, h_s_arrmul12_nand8_11_y0);
  fa fa_h_s_arrmul12_fa8_11_y2(h_s_arrmul12_nand8_11_y0, h_s_arrmul12_fa9_10_y2, h_s_arrmul12_fa7_11_y4, h_s_arrmul12_fa8_11_y2, h_s_arrmul12_fa8_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand9_11_y0(a_9, b_11, h_s_arrmul12_nand9_11_y0);
  fa fa_h_s_arrmul12_fa9_11_y2(h_s_arrmul12_nand9_11_y0, h_s_arrmul12_fa10_10_y2, h_s_arrmul12_fa8_11_y4, h_s_arrmul12_fa9_11_y2, h_s_arrmul12_fa9_11_y4);
  nand_gate nand_gate_h_s_arrmul12_nand10_11_y0(a_10, b_11, h_s_arrmul12_nand10_11_y0);
  fa fa_h_s_arrmul12_fa10_11_y2(h_s_arrmul12_nand10_11_y0, h_s_arrmul12_fa11_10_y2, h_s_arrmul12_fa9_11_y4, h_s_arrmul12_fa10_11_y2, h_s_arrmul12_fa10_11_y4);
  and_gate and_gate_h_s_arrmul12_and11_11_y0(a_11, b_11, h_s_arrmul12_and11_11_y0);
  fa fa_h_s_arrmul12_fa11_11_y2(h_s_arrmul12_and11_11_y0, h_s_arrmul12_fa11_10_y4, h_s_arrmul12_fa10_11_y4, h_s_arrmul12_fa11_11_y2, h_s_arrmul12_fa11_11_y4);
  xor_gate xor_gate_h_s_arrmul12_xor12_11_y0(h_s_arrmul12_fa11_11_y4, constant_wire_1, h_s_arrmul12_xor12_11_y0);

  assign out[0] = h_s_arrmul12_and0_0_y0;
  assign out[1] = h_s_arrmul12_ha0_1_y0;
  assign out[2] = h_s_arrmul12_ha0_2_y0;
  assign out[3] = h_s_arrmul12_ha0_3_y0;
  assign out[4] = h_s_arrmul12_ha0_4_y0;
  assign out[5] = h_s_arrmul12_ha0_5_y0;
  assign out[6] = h_s_arrmul12_ha0_6_y0;
  assign out[7] = h_s_arrmul12_ha0_7_y0;
  assign out[8] = h_s_arrmul12_ha0_8_y0;
  assign out[9] = h_s_arrmul12_ha0_9_y0;
  assign out[10] = h_s_arrmul12_ha0_10_y0;
  assign out[11] = h_s_arrmul12_ha0_11_y0;
  assign out[12] = h_s_arrmul12_fa1_11_y2;
  assign out[13] = h_s_arrmul12_fa2_11_y2;
  assign out[14] = h_s_arrmul12_fa3_11_y2;
  assign out[15] = h_s_arrmul12_fa4_11_y2;
  assign out[16] = h_s_arrmul12_fa5_11_y2;
  assign out[17] = h_s_arrmul12_fa6_11_y2;
  assign out[18] = h_s_arrmul12_fa7_11_y2;
  assign out[19] = h_s_arrmul12_fa8_11_y2;
  assign out[20] = h_s_arrmul12_fa9_11_y2;
  assign out[21] = h_s_arrmul12_fa10_11_y2;
  assign out[22] = h_s_arrmul12_fa11_11_y2;
  assign out[23] = h_s_arrmul12_xor12_11_y0;
endmodule