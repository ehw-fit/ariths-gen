module s_dadda_cska12(input [11:0] a, input [11:0] b, output [23:0] s_dadda_cska12_out);
  wire s_dadda_cska12_and_9_0;
  wire s_dadda_cska12_and_8_1;
  wire s_dadda_cska12_ha0_xor0;
  wire s_dadda_cska12_ha0_and0;
  wire s_dadda_cska12_and_10_0;
  wire s_dadda_cska12_and_9_1;
  wire s_dadda_cska12_fa0_xor0;
  wire s_dadda_cska12_fa0_and0;
  wire s_dadda_cska12_fa0_xor1;
  wire s_dadda_cska12_fa0_and1;
  wire s_dadda_cska12_fa0_or0;
  wire s_dadda_cska12_and_8_2;
  wire s_dadda_cska12_and_7_3;
  wire s_dadda_cska12_ha1_xor0;
  wire s_dadda_cska12_ha1_and0;
  wire s_dadda_cska12_nand_11_0;
  wire s_dadda_cska12_fa1_xor0;
  wire s_dadda_cska12_fa1_and0;
  wire s_dadda_cska12_fa1_xor1;
  wire s_dadda_cska12_fa1_and1;
  wire s_dadda_cska12_fa1_or0;
  wire s_dadda_cska12_and_10_1;
  wire s_dadda_cska12_and_9_2;
  wire s_dadda_cska12_and_8_3;
  wire s_dadda_cska12_fa2_xor0;
  wire s_dadda_cska12_fa2_and0;
  wire s_dadda_cska12_fa2_xor1;
  wire s_dadda_cska12_fa2_and1;
  wire s_dadda_cska12_fa2_or0;
  wire s_dadda_cska12_and_7_4;
  wire s_dadda_cska12_and_6_5;
  wire s_dadda_cska12_ha2_xor0;
  wire s_dadda_cska12_ha2_and0;
  wire s_dadda_cska12_fa3_xor0;
  wire s_dadda_cska12_fa3_and0;
  wire s_dadda_cska12_fa3_xor1;
  wire s_dadda_cska12_fa3_and1;
  wire s_dadda_cska12_fa3_or0;
  wire s_dadda_cska12_nand_11_1;
  wire s_dadda_cska12_and_10_2;
  wire s_dadda_cska12_fa4_xor0;
  wire s_dadda_cska12_fa4_xor1;
  wire s_dadda_cska12_fa4_and1;
  wire s_dadda_cska12_fa4_or0;
  wire s_dadda_cska12_and_9_3;
  wire s_dadda_cska12_and_8_4;
  wire s_dadda_cska12_and_7_5;
  wire s_dadda_cska12_fa5_xor0;
  wire s_dadda_cska12_fa5_and0;
  wire s_dadda_cska12_fa5_xor1;
  wire s_dadda_cska12_fa5_and1;
  wire s_dadda_cska12_fa5_or0;
  wire s_dadda_cska12_fa6_xor0;
  wire s_dadda_cska12_fa6_and0;
  wire s_dadda_cska12_fa6_xor1;
  wire s_dadda_cska12_fa6_and1;
  wire s_dadda_cska12_fa6_or0;
  wire s_dadda_cska12_nand_11_2;
  wire s_dadda_cska12_and_10_3;
  wire s_dadda_cska12_and_9_4;
  wire s_dadda_cska12_fa7_xor0;
  wire s_dadda_cska12_fa7_and0;
  wire s_dadda_cska12_fa7_xor1;
  wire s_dadda_cska12_fa7_and1;
  wire s_dadda_cska12_fa7_or0;
  wire s_dadda_cska12_nand_11_3;
  wire s_dadda_cska12_fa8_xor0;
  wire s_dadda_cska12_fa8_and0;
  wire s_dadda_cska12_fa8_xor1;
  wire s_dadda_cska12_fa8_and1;
  wire s_dadda_cska12_fa8_or0;
  wire s_dadda_cska12_and_4_0;
  wire s_dadda_cska12_and_3_1;
  wire s_dadda_cska12_ha3_xor0;
  wire s_dadda_cska12_ha3_and0;
  wire s_dadda_cska12_and_5_0;
  wire s_dadda_cska12_and_4_1;
  wire s_dadda_cska12_fa9_xor0;
  wire s_dadda_cska12_fa9_and0;
  wire s_dadda_cska12_fa9_xor1;
  wire s_dadda_cska12_fa9_and1;
  wire s_dadda_cska12_fa9_or0;
  wire s_dadda_cska12_and_3_2;
  wire s_dadda_cska12_and_2_3;
  wire s_dadda_cska12_ha4_xor0;
  wire s_dadda_cska12_ha4_and0;
  wire s_dadda_cska12_and_6_0;
  wire s_dadda_cska12_fa10_xor0;
  wire s_dadda_cska12_fa10_and0;
  wire s_dadda_cska12_fa10_xor1;
  wire s_dadda_cska12_fa10_and1;
  wire s_dadda_cska12_fa10_or0;
  wire s_dadda_cska12_and_5_1;
  wire s_dadda_cska12_and_4_2;
  wire s_dadda_cska12_and_3_3;
  wire s_dadda_cska12_fa11_xor0;
  wire s_dadda_cska12_fa11_and0;
  wire s_dadda_cska12_fa11_xor1;
  wire s_dadda_cska12_fa11_and1;
  wire s_dadda_cska12_fa11_or0;
  wire s_dadda_cska12_and_2_4;
  wire s_dadda_cska12_and_1_5;
  wire s_dadda_cska12_ha5_xor0;
  wire s_dadda_cska12_ha5_and0;
  wire s_dadda_cska12_fa12_xor0;
  wire s_dadda_cska12_fa12_and0;
  wire s_dadda_cska12_fa12_xor1;
  wire s_dadda_cska12_fa12_and1;
  wire s_dadda_cska12_fa12_or0;
  wire s_dadda_cska12_and_7_0;
  wire s_dadda_cska12_and_6_1;
  wire s_dadda_cska12_and_5_2;
  wire s_dadda_cska12_fa13_xor0;
  wire s_dadda_cska12_fa13_and0;
  wire s_dadda_cska12_fa13_xor1;
  wire s_dadda_cska12_fa13_and1;
  wire s_dadda_cska12_fa13_or0;
  wire s_dadda_cska12_and_4_3;
  wire s_dadda_cska12_and_3_4;
  wire s_dadda_cska12_and_2_5;
  wire s_dadda_cska12_fa14_xor0;
  wire s_dadda_cska12_fa14_and0;
  wire s_dadda_cska12_fa14_xor1;
  wire s_dadda_cska12_fa14_and1;
  wire s_dadda_cska12_fa14_or0;
  wire s_dadda_cska12_and_1_6;
  wire s_dadda_cska12_and_0_7;
  wire s_dadda_cska12_ha6_xor0;
  wire s_dadda_cska12_ha6_and0;
  wire s_dadda_cska12_fa15_xor0;
  wire s_dadda_cska12_fa15_and0;
  wire s_dadda_cska12_fa15_xor1;
  wire s_dadda_cska12_fa15_and1;
  wire s_dadda_cska12_fa15_or0;
  wire s_dadda_cska12_and_8_0;
  wire s_dadda_cska12_and_7_1;
  wire s_dadda_cska12_fa16_xor0;
  wire s_dadda_cska12_fa16_and0;
  wire s_dadda_cska12_fa16_xor1;
  wire s_dadda_cska12_fa16_and1;
  wire s_dadda_cska12_fa16_or0;
  wire s_dadda_cska12_and_6_2;
  wire s_dadda_cska12_and_5_3;
  wire s_dadda_cska12_and_4_4;
  wire s_dadda_cska12_fa17_xor0;
  wire s_dadda_cska12_fa17_and0;
  wire s_dadda_cska12_fa17_xor1;
  wire s_dadda_cska12_fa17_and1;
  wire s_dadda_cska12_fa17_or0;
  wire s_dadda_cska12_and_3_5;
  wire s_dadda_cska12_and_2_6;
  wire s_dadda_cska12_and_1_7;
  wire s_dadda_cska12_fa18_xor0;
  wire s_dadda_cska12_fa18_and0;
  wire s_dadda_cska12_fa18_xor1;
  wire s_dadda_cska12_fa18_and1;
  wire s_dadda_cska12_fa18_or0;
  wire s_dadda_cska12_and_0_8;
  wire s_dadda_cska12_ha7_xor0;
  wire s_dadda_cska12_ha7_and0;
  wire s_dadda_cska12_fa19_xor0;
  wire s_dadda_cska12_fa19_and0;
  wire s_dadda_cska12_fa19_xor1;
  wire s_dadda_cska12_fa19_and1;
  wire s_dadda_cska12_fa19_or0;
  wire s_dadda_cska12_and_7_2;
  wire s_dadda_cska12_fa20_xor0;
  wire s_dadda_cska12_fa20_and0;
  wire s_dadda_cska12_fa20_xor1;
  wire s_dadda_cska12_fa20_and1;
  wire s_dadda_cska12_fa20_or0;
  wire s_dadda_cska12_and_6_3;
  wire s_dadda_cska12_and_5_4;
  wire s_dadda_cska12_and_4_5;
  wire s_dadda_cska12_fa21_xor0;
  wire s_dadda_cska12_fa21_and0;
  wire s_dadda_cska12_fa21_xor1;
  wire s_dadda_cska12_fa21_and1;
  wire s_dadda_cska12_fa21_or0;
  wire s_dadda_cska12_and_3_6;
  wire s_dadda_cska12_and_2_7;
  wire s_dadda_cska12_and_1_8;
  wire s_dadda_cska12_fa22_xor0;
  wire s_dadda_cska12_fa22_and0;
  wire s_dadda_cska12_fa22_xor1;
  wire s_dadda_cska12_fa22_and1;
  wire s_dadda_cska12_fa22_or0;
  wire s_dadda_cska12_and_0_9;
  wire s_dadda_cska12_fa23_xor0;
  wire s_dadda_cska12_fa23_and0;
  wire s_dadda_cska12_fa23_xor1;
  wire s_dadda_cska12_fa23_and1;
  wire s_dadda_cska12_fa23_or0;
  wire s_dadda_cska12_fa24_xor0;
  wire s_dadda_cska12_fa24_and0;
  wire s_dadda_cska12_fa24_xor1;
  wire s_dadda_cska12_fa24_and1;
  wire s_dadda_cska12_fa24_or0;
  wire s_dadda_cska12_and_6_4;
  wire s_dadda_cska12_fa25_xor0;
  wire s_dadda_cska12_fa25_and0;
  wire s_dadda_cska12_fa25_xor1;
  wire s_dadda_cska12_fa25_and1;
  wire s_dadda_cska12_fa25_or0;
  wire s_dadda_cska12_and_5_5;
  wire s_dadda_cska12_and_4_6;
  wire s_dadda_cska12_and_3_7;
  wire s_dadda_cska12_fa26_xor0;
  wire s_dadda_cska12_fa26_and0;
  wire s_dadda_cska12_fa26_xor1;
  wire s_dadda_cska12_fa26_and1;
  wire s_dadda_cska12_fa26_or0;
  wire s_dadda_cska12_and_2_8;
  wire s_dadda_cska12_and_1_9;
  wire s_dadda_cska12_and_0_10;
  wire s_dadda_cska12_fa27_xor0;
  wire s_dadda_cska12_fa27_and0;
  wire s_dadda_cska12_fa27_xor1;
  wire s_dadda_cska12_fa27_and1;
  wire s_dadda_cska12_fa27_or0;
  wire s_dadda_cska12_fa28_xor0;
  wire s_dadda_cska12_fa28_and0;
  wire s_dadda_cska12_fa28_xor1;
  wire s_dadda_cska12_fa28_and1;
  wire s_dadda_cska12_fa28_or0;
  wire s_dadda_cska12_fa29_xor0;
  wire s_dadda_cska12_fa29_and0;
  wire s_dadda_cska12_fa29_xor1;
  wire s_dadda_cska12_fa29_and1;
  wire s_dadda_cska12_fa29_or0;
  wire s_dadda_cska12_and_5_6;
  wire s_dadda_cska12_fa30_xor0;
  wire s_dadda_cska12_fa30_and0;
  wire s_dadda_cska12_fa30_xor1;
  wire s_dadda_cska12_fa30_and1;
  wire s_dadda_cska12_fa30_or0;
  wire s_dadda_cska12_and_4_7;
  wire s_dadda_cska12_and_3_8;
  wire s_dadda_cska12_and_2_9;
  wire s_dadda_cska12_fa31_xor0;
  wire s_dadda_cska12_fa31_and0;
  wire s_dadda_cska12_fa31_xor1;
  wire s_dadda_cska12_fa31_and1;
  wire s_dadda_cska12_fa31_or0;
  wire s_dadda_cska12_and_1_10;
  wire s_dadda_cska12_nand_0_11;
  wire s_dadda_cska12_fa32_xor0;
  wire s_dadda_cska12_fa32_and0;
  wire s_dadda_cska12_fa32_xor1;
  wire s_dadda_cska12_fa32_and1;
  wire s_dadda_cska12_fa32_or0;
  wire s_dadda_cska12_fa33_xor0;
  wire s_dadda_cska12_fa33_and0;
  wire s_dadda_cska12_fa33_xor1;
  wire s_dadda_cska12_fa33_and1;
  wire s_dadda_cska12_fa33_or0;
  wire s_dadda_cska12_fa34_xor0;
  wire s_dadda_cska12_fa34_and0;
  wire s_dadda_cska12_fa34_xor1;
  wire s_dadda_cska12_fa34_and1;
  wire s_dadda_cska12_fa34_or0;
  wire s_dadda_cska12_and_6_6;
  wire s_dadda_cska12_fa35_xor0;
  wire s_dadda_cska12_fa35_and0;
  wire s_dadda_cska12_fa35_xor1;
  wire s_dadda_cska12_fa35_and1;
  wire s_dadda_cska12_fa35_or0;
  wire s_dadda_cska12_and_5_7;
  wire s_dadda_cska12_and_4_8;
  wire s_dadda_cska12_and_3_9;
  wire s_dadda_cska12_fa36_xor0;
  wire s_dadda_cska12_fa36_and0;
  wire s_dadda_cska12_fa36_xor1;
  wire s_dadda_cska12_fa36_and1;
  wire s_dadda_cska12_fa36_or0;
  wire s_dadda_cska12_and_2_10;
  wire s_dadda_cska12_nand_1_11;
  wire s_dadda_cska12_fa37_xor0;
  wire s_dadda_cska12_fa37_and0;
  wire s_dadda_cska12_fa37_xor1;
  wire s_dadda_cska12_fa37_and1;
  wire s_dadda_cska12_fa37_or0;
  wire s_dadda_cska12_fa38_xor0;
  wire s_dadda_cska12_fa38_and0;
  wire s_dadda_cska12_fa38_xor1;
  wire s_dadda_cska12_fa38_and1;
  wire s_dadda_cska12_fa38_or0;
  wire s_dadda_cska12_fa39_xor0;
  wire s_dadda_cska12_fa39_and0;
  wire s_dadda_cska12_fa39_xor1;
  wire s_dadda_cska12_fa39_and1;
  wire s_dadda_cska12_fa39_or0;
  wire s_dadda_cska12_and_8_5;
  wire s_dadda_cska12_fa40_xor0;
  wire s_dadda_cska12_fa40_and0;
  wire s_dadda_cska12_fa40_xor1;
  wire s_dadda_cska12_fa40_and1;
  wire s_dadda_cska12_fa40_or0;
  wire s_dadda_cska12_and_7_6;
  wire s_dadda_cska12_and_6_7;
  wire s_dadda_cska12_and_5_8;
  wire s_dadda_cska12_fa41_xor0;
  wire s_dadda_cska12_fa41_and0;
  wire s_dadda_cska12_fa41_xor1;
  wire s_dadda_cska12_fa41_and1;
  wire s_dadda_cska12_fa41_or0;
  wire s_dadda_cska12_and_4_9;
  wire s_dadda_cska12_and_3_10;
  wire s_dadda_cska12_nand_2_11;
  wire s_dadda_cska12_fa42_xor0;
  wire s_dadda_cska12_fa42_and0;
  wire s_dadda_cska12_fa42_xor1;
  wire s_dadda_cska12_fa42_and1;
  wire s_dadda_cska12_fa42_or0;
  wire s_dadda_cska12_fa43_xor0;
  wire s_dadda_cska12_fa43_and0;
  wire s_dadda_cska12_fa43_xor1;
  wire s_dadda_cska12_fa43_and1;
  wire s_dadda_cska12_fa43_or0;
  wire s_dadda_cska12_fa44_xor0;
  wire s_dadda_cska12_fa44_and0;
  wire s_dadda_cska12_fa44_xor1;
  wire s_dadda_cska12_fa44_and1;
  wire s_dadda_cska12_fa44_or0;
  wire s_dadda_cska12_and_10_4;
  wire s_dadda_cska12_fa45_xor0;
  wire s_dadda_cska12_fa45_and0;
  wire s_dadda_cska12_fa45_xor1;
  wire s_dadda_cska12_fa45_and1;
  wire s_dadda_cska12_fa45_or0;
  wire s_dadda_cska12_and_9_5;
  wire s_dadda_cska12_and_8_6;
  wire s_dadda_cska12_and_7_7;
  wire s_dadda_cska12_fa46_xor0;
  wire s_dadda_cska12_fa46_and0;
  wire s_dadda_cska12_fa46_xor1;
  wire s_dadda_cska12_fa46_and1;
  wire s_dadda_cska12_fa46_or0;
  wire s_dadda_cska12_and_6_8;
  wire s_dadda_cska12_and_5_9;
  wire s_dadda_cska12_and_4_10;
  wire s_dadda_cska12_fa47_xor0;
  wire s_dadda_cska12_fa47_and0;
  wire s_dadda_cska12_fa47_xor1;
  wire s_dadda_cska12_fa47_and1;
  wire s_dadda_cska12_fa47_or0;
  wire s_dadda_cska12_nand_3_11;
  wire s_dadda_cska12_fa48_xor0;
  wire s_dadda_cska12_fa48_and0;
  wire s_dadda_cska12_fa48_xor1;
  wire s_dadda_cska12_fa48_and1;
  wire s_dadda_cska12_fa48_or0;
  wire s_dadda_cska12_fa49_xor0;
  wire s_dadda_cska12_fa49_and0;
  wire s_dadda_cska12_fa49_xor1;
  wire s_dadda_cska12_fa49_and1;
  wire s_dadda_cska12_fa49_or0;
  wire s_dadda_cska12_fa50_xor0;
  wire s_dadda_cska12_fa50_and0;
  wire s_dadda_cska12_fa50_xor1;
  wire s_dadda_cska12_fa50_and1;
  wire s_dadda_cska12_fa50_or0;
  wire s_dadda_cska12_nand_11_4;
  wire s_dadda_cska12_and_10_5;
  wire s_dadda_cska12_and_9_6;
  wire s_dadda_cska12_fa51_xor0;
  wire s_dadda_cska12_fa51_and0;
  wire s_dadda_cska12_fa51_xor1;
  wire s_dadda_cska12_fa51_and1;
  wire s_dadda_cska12_fa51_or0;
  wire s_dadda_cska12_and_8_7;
  wire s_dadda_cska12_and_7_8;
  wire s_dadda_cska12_and_6_9;
  wire s_dadda_cska12_fa52_xor0;
  wire s_dadda_cska12_fa52_and0;
  wire s_dadda_cska12_fa52_xor1;
  wire s_dadda_cska12_fa52_and1;
  wire s_dadda_cska12_fa52_or0;
  wire s_dadda_cska12_and_5_10;
  wire s_dadda_cska12_nand_4_11;
  wire s_dadda_cska12_fa53_xor0;
  wire s_dadda_cska12_fa53_and0;
  wire s_dadda_cska12_fa53_xor1;
  wire s_dadda_cska12_fa53_and1;
  wire s_dadda_cska12_fa53_or0;
  wire s_dadda_cska12_fa54_xor0;
  wire s_dadda_cska12_fa54_and0;
  wire s_dadda_cska12_fa54_xor1;
  wire s_dadda_cska12_fa54_and1;
  wire s_dadda_cska12_fa54_or0;
  wire s_dadda_cska12_nand_11_5;
  wire s_dadda_cska12_fa55_xor0;
  wire s_dadda_cska12_fa55_and0;
  wire s_dadda_cska12_fa55_xor1;
  wire s_dadda_cska12_fa55_and1;
  wire s_dadda_cska12_fa55_or0;
  wire s_dadda_cska12_and_10_6;
  wire s_dadda_cska12_and_9_7;
  wire s_dadda_cska12_and_8_8;
  wire s_dadda_cska12_fa56_xor0;
  wire s_dadda_cska12_fa56_and0;
  wire s_dadda_cska12_fa56_xor1;
  wire s_dadda_cska12_fa56_and1;
  wire s_dadda_cska12_fa56_or0;
  wire s_dadda_cska12_and_7_9;
  wire s_dadda_cska12_and_6_10;
  wire s_dadda_cska12_nand_5_11;
  wire s_dadda_cska12_fa57_xor0;
  wire s_dadda_cska12_fa57_and0;
  wire s_dadda_cska12_fa57_xor1;
  wire s_dadda_cska12_fa57_and1;
  wire s_dadda_cska12_fa57_or0;
  wire s_dadda_cska12_fa58_xor0;
  wire s_dadda_cska12_fa58_and0;
  wire s_dadda_cska12_fa58_xor1;
  wire s_dadda_cska12_fa58_and1;
  wire s_dadda_cska12_fa58_or0;
  wire s_dadda_cska12_nand_11_6;
  wire s_dadda_cska12_and_10_7;
  wire s_dadda_cska12_fa59_xor0;
  wire s_dadda_cska12_fa59_and0;
  wire s_dadda_cska12_fa59_xor1;
  wire s_dadda_cska12_fa59_and1;
  wire s_dadda_cska12_fa59_or0;
  wire s_dadda_cska12_and_9_8;
  wire s_dadda_cska12_and_8_9;
  wire s_dadda_cska12_and_7_10;
  wire s_dadda_cska12_fa60_xor0;
  wire s_dadda_cska12_fa60_and0;
  wire s_dadda_cska12_fa60_xor1;
  wire s_dadda_cska12_fa60_and1;
  wire s_dadda_cska12_fa60_or0;
  wire s_dadda_cska12_fa61_xor0;
  wire s_dadda_cska12_fa61_and0;
  wire s_dadda_cska12_fa61_xor1;
  wire s_dadda_cska12_fa61_and1;
  wire s_dadda_cska12_fa61_or0;
  wire s_dadda_cska12_nand_11_7;
  wire s_dadda_cska12_and_10_8;
  wire s_dadda_cska12_and_9_9;
  wire s_dadda_cska12_fa62_xor0;
  wire s_dadda_cska12_fa62_and0;
  wire s_dadda_cska12_fa62_xor1;
  wire s_dadda_cska12_fa62_and1;
  wire s_dadda_cska12_fa62_or0;
  wire s_dadda_cska12_nand_11_8;
  wire s_dadda_cska12_fa63_xor0;
  wire s_dadda_cska12_fa63_and0;
  wire s_dadda_cska12_fa63_xor1;
  wire s_dadda_cska12_fa63_and1;
  wire s_dadda_cska12_fa63_or0;
  wire s_dadda_cska12_and_3_0;
  wire s_dadda_cska12_and_2_1;
  wire s_dadda_cska12_ha8_xor0;
  wire s_dadda_cska12_ha8_and0;
  wire s_dadda_cska12_and_2_2;
  wire s_dadda_cska12_and_1_3;
  wire s_dadda_cska12_fa64_xor0;
  wire s_dadda_cska12_fa64_and0;
  wire s_dadda_cska12_fa64_xor1;
  wire s_dadda_cska12_fa64_and1;
  wire s_dadda_cska12_fa64_or0;
  wire s_dadda_cska12_and_1_4;
  wire s_dadda_cska12_and_0_5;
  wire s_dadda_cska12_fa65_xor0;
  wire s_dadda_cska12_fa65_and0;
  wire s_dadda_cska12_fa65_xor1;
  wire s_dadda_cska12_fa65_and1;
  wire s_dadda_cska12_fa65_or0;
  wire s_dadda_cska12_and_0_6;
  wire s_dadda_cska12_fa66_xor0;
  wire s_dadda_cska12_fa66_and0;
  wire s_dadda_cska12_fa66_xor1;
  wire s_dadda_cska12_fa66_and1;
  wire s_dadda_cska12_fa66_or0;
  wire s_dadda_cska12_fa67_xor0;
  wire s_dadda_cska12_fa67_and0;
  wire s_dadda_cska12_fa67_xor1;
  wire s_dadda_cska12_fa67_and1;
  wire s_dadda_cska12_fa67_or0;
  wire s_dadda_cska12_fa68_xor0;
  wire s_dadda_cska12_fa68_and0;
  wire s_dadda_cska12_fa68_xor1;
  wire s_dadda_cska12_fa68_and1;
  wire s_dadda_cska12_fa68_or0;
  wire s_dadda_cska12_fa69_xor0;
  wire s_dadda_cska12_fa69_and0;
  wire s_dadda_cska12_fa69_xor1;
  wire s_dadda_cska12_fa69_and1;
  wire s_dadda_cska12_fa69_or0;
  wire s_dadda_cska12_fa70_xor0;
  wire s_dadda_cska12_fa70_and0;
  wire s_dadda_cska12_fa70_xor1;
  wire s_dadda_cska12_fa70_and1;
  wire s_dadda_cska12_fa70_or0;
  wire s_dadda_cska12_fa71_xor0;
  wire s_dadda_cska12_fa71_and0;
  wire s_dadda_cska12_fa71_xor1;
  wire s_dadda_cska12_fa71_and1;
  wire s_dadda_cska12_fa71_or0;
  wire s_dadda_cska12_fa72_xor0;
  wire s_dadda_cska12_fa72_and0;
  wire s_dadda_cska12_fa72_xor1;
  wire s_dadda_cska12_fa72_and1;
  wire s_dadda_cska12_fa72_or0;
  wire s_dadda_cska12_fa73_xor0;
  wire s_dadda_cska12_fa73_and0;
  wire s_dadda_cska12_fa73_xor1;
  wire s_dadda_cska12_fa73_and1;
  wire s_dadda_cska12_fa73_or0;
  wire s_dadda_cska12_fa74_xor0;
  wire s_dadda_cska12_fa74_and0;
  wire s_dadda_cska12_fa74_xor1;
  wire s_dadda_cska12_fa74_and1;
  wire s_dadda_cska12_fa74_or0;
  wire s_dadda_cska12_fa75_xor0;
  wire s_dadda_cska12_fa75_and0;
  wire s_dadda_cska12_fa75_xor1;
  wire s_dadda_cska12_fa75_and1;
  wire s_dadda_cska12_fa75_or0;
  wire s_dadda_cska12_fa76_xor0;
  wire s_dadda_cska12_fa76_and0;
  wire s_dadda_cska12_fa76_xor1;
  wire s_dadda_cska12_fa76_and1;
  wire s_dadda_cska12_fa76_or0;
  wire s_dadda_cska12_nand_6_11;
  wire s_dadda_cska12_fa77_xor0;
  wire s_dadda_cska12_fa77_and0;
  wire s_dadda_cska12_fa77_xor1;
  wire s_dadda_cska12_fa77_and1;
  wire s_dadda_cska12_fa77_or0;
  wire s_dadda_cska12_and_8_10;
  wire s_dadda_cska12_nand_7_11;
  wire s_dadda_cska12_fa78_xor0;
  wire s_dadda_cska12_fa78_and0;
  wire s_dadda_cska12_fa78_xor1;
  wire s_dadda_cska12_fa78_and1;
  wire s_dadda_cska12_fa78_or0;
  wire s_dadda_cska12_and_10_9;
  wire s_dadda_cska12_and_9_10;
  wire s_dadda_cska12_fa79_xor0;
  wire s_dadda_cska12_fa79_and0;
  wire s_dadda_cska12_fa79_xor1;
  wire s_dadda_cska12_fa79_and1;
  wire s_dadda_cska12_fa79_or0;
  wire s_dadda_cska12_nand_11_9;
  wire s_dadda_cska12_fa80_xor0;
  wire s_dadda_cska12_fa80_and0;
  wire s_dadda_cska12_fa80_xor1;
  wire s_dadda_cska12_fa80_and1;
  wire s_dadda_cska12_fa80_or0;
  wire s_dadda_cska12_and_2_0;
  wire s_dadda_cska12_and_1_1;
  wire s_dadda_cska12_ha9_xor0;
  wire s_dadda_cska12_ha9_and0;
  wire s_dadda_cska12_and_1_2;
  wire s_dadda_cska12_and_0_3;
  wire s_dadda_cska12_fa81_xor0;
  wire s_dadda_cska12_fa81_and0;
  wire s_dadda_cska12_fa81_xor1;
  wire s_dadda_cska12_fa81_and1;
  wire s_dadda_cska12_fa81_or0;
  wire s_dadda_cska12_and_0_4;
  wire s_dadda_cska12_fa82_xor0;
  wire s_dadda_cska12_fa82_and0;
  wire s_dadda_cska12_fa82_xor1;
  wire s_dadda_cska12_fa82_and1;
  wire s_dadda_cska12_fa82_or0;
  wire s_dadda_cska12_fa83_xor0;
  wire s_dadda_cska12_fa83_and0;
  wire s_dadda_cska12_fa83_xor1;
  wire s_dadda_cska12_fa83_and1;
  wire s_dadda_cska12_fa83_or0;
  wire s_dadda_cska12_fa84_xor0;
  wire s_dadda_cska12_fa84_and0;
  wire s_dadda_cska12_fa84_xor1;
  wire s_dadda_cska12_fa84_and1;
  wire s_dadda_cska12_fa84_or0;
  wire s_dadda_cska12_fa85_xor0;
  wire s_dadda_cska12_fa85_and0;
  wire s_dadda_cska12_fa85_xor1;
  wire s_dadda_cska12_fa85_and1;
  wire s_dadda_cska12_fa85_or0;
  wire s_dadda_cska12_fa86_xor0;
  wire s_dadda_cska12_fa86_and0;
  wire s_dadda_cska12_fa86_xor1;
  wire s_dadda_cska12_fa86_and1;
  wire s_dadda_cska12_fa86_or0;
  wire s_dadda_cska12_fa87_xor0;
  wire s_dadda_cska12_fa87_and0;
  wire s_dadda_cska12_fa87_xor1;
  wire s_dadda_cska12_fa87_and1;
  wire s_dadda_cska12_fa87_or0;
  wire s_dadda_cska12_fa88_xor0;
  wire s_dadda_cska12_fa88_and0;
  wire s_dadda_cska12_fa88_xor1;
  wire s_dadda_cska12_fa88_and1;
  wire s_dadda_cska12_fa88_or0;
  wire s_dadda_cska12_fa89_xor0;
  wire s_dadda_cska12_fa89_and0;
  wire s_dadda_cska12_fa89_xor1;
  wire s_dadda_cska12_fa89_and1;
  wire s_dadda_cska12_fa89_or0;
  wire s_dadda_cska12_fa90_xor0;
  wire s_dadda_cska12_fa90_and0;
  wire s_dadda_cska12_fa90_xor1;
  wire s_dadda_cska12_fa90_and1;
  wire s_dadda_cska12_fa90_or0;
  wire s_dadda_cska12_fa91_xor0;
  wire s_dadda_cska12_fa91_and0;
  wire s_dadda_cska12_fa91_xor1;
  wire s_dadda_cska12_fa91_and1;
  wire s_dadda_cska12_fa91_or0;
  wire s_dadda_cska12_fa92_xor0;
  wire s_dadda_cska12_fa92_and0;
  wire s_dadda_cska12_fa92_xor1;
  wire s_dadda_cska12_fa92_and1;
  wire s_dadda_cska12_fa92_or0;
  wire s_dadda_cska12_fa93_xor0;
  wire s_dadda_cska12_fa93_and0;
  wire s_dadda_cska12_fa93_xor1;
  wire s_dadda_cska12_fa93_and1;
  wire s_dadda_cska12_fa93_or0;
  wire s_dadda_cska12_fa94_xor0;
  wire s_dadda_cska12_fa94_and0;
  wire s_dadda_cska12_fa94_xor1;
  wire s_dadda_cska12_fa94_and1;
  wire s_dadda_cska12_fa94_or0;
  wire s_dadda_cska12_fa95_xor0;
  wire s_dadda_cska12_fa95_and0;
  wire s_dadda_cska12_fa95_xor1;
  wire s_dadda_cska12_fa95_and1;
  wire s_dadda_cska12_fa95_or0;
  wire s_dadda_cska12_fa96_xor0;
  wire s_dadda_cska12_fa96_and0;
  wire s_dadda_cska12_fa96_xor1;
  wire s_dadda_cska12_fa96_and1;
  wire s_dadda_cska12_fa96_or0;
  wire s_dadda_cska12_nand_8_11;
  wire s_dadda_cska12_fa97_xor0;
  wire s_dadda_cska12_fa97_and0;
  wire s_dadda_cska12_fa97_xor1;
  wire s_dadda_cska12_fa97_and1;
  wire s_dadda_cska12_fa97_or0;
  wire s_dadda_cska12_and_10_10;
  wire s_dadda_cska12_nand_9_11;
  wire s_dadda_cska12_fa98_xor0;
  wire s_dadda_cska12_fa98_and0;
  wire s_dadda_cska12_fa98_xor1;
  wire s_dadda_cska12_fa98_and1;
  wire s_dadda_cska12_fa98_or0;
  wire s_dadda_cska12_nand_11_10;
  wire s_dadda_cska12_fa99_xor0;
  wire s_dadda_cska12_fa99_and0;
  wire s_dadda_cska12_fa99_xor1;
  wire s_dadda_cska12_fa99_and1;
  wire s_dadda_cska12_fa99_or0;
  wire s_dadda_cska12_and_0_0;
  wire s_dadda_cska12_and_1_0;
  wire s_dadda_cska12_and_0_2;
  wire s_dadda_cska12_nand_10_11;
  wire s_dadda_cska12_and_0_1;
  wire s_dadda_cska12_and_11_11;
  wire s_dadda_cska12_u_cska22_xor0;
  wire s_dadda_cska12_u_cska22_ha0_xor0;
  wire s_dadda_cska12_u_cska22_ha0_and0;
  wire s_dadda_cska12_u_cska22_xor1;
  wire s_dadda_cska12_u_cska22_fa0_xor0;
  wire s_dadda_cska12_u_cska22_fa0_and0;
  wire s_dadda_cska12_u_cska22_fa0_xor1;
  wire s_dadda_cska12_u_cska22_fa0_and1;
  wire s_dadda_cska12_u_cska22_fa0_or0;
  wire s_dadda_cska12_u_cska22_xor2;
  wire s_dadda_cska12_u_cska22_fa1_xor0;
  wire s_dadda_cska12_u_cska22_fa1_and0;
  wire s_dadda_cska12_u_cska22_fa1_xor1;
  wire s_dadda_cska12_u_cska22_fa1_and1;
  wire s_dadda_cska12_u_cska22_fa1_or0;
  wire s_dadda_cska12_u_cska22_xor3;
  wire s_dadda_cska12_u_cska22_fa2_xor0;
  wire s_dadda_cska12_u_cska22_fa2_and0;
  wire s_dadda_cska12_u_cska22_fa2_xor1;
  wire s_dadda_cska12_u_cska22_fa2_and1;
  wire s_dadda_cska12_u_cska22_fa2_or0;
  wire s_dadda_cska12_u_cska22_and_propagate00;
  wire s_dadda_cska12_u_cska22_and_propagate01;
  wire s_dadda_cska12_u_cska22_and_propagate02;
  wire s_dadda_cska12_u_cska22_mux2to10_not0;
  wire s_dadda_cska12_u_cska22_mux2to10_and1;
  wire s_dadda_cska12_u_cska22_xor4;
  wire s_dadda_cska12_u_cska22_fa3_xor0;
  wire s_dadda_cska12_u_cska22_fa3_and0;
  wire s_dadda_cska12_u_cska22_fa3_xor1;
  wire s_dadda_cska12_u_cska22_fa3_and1;
  wire s_dadda_cska12_u_cska22_fa3_or0;
  wire s_dadda_cska12_u_cska22_xor5;
  wire s_dadda_cska12_u_cska22_fa4_xor0;
  wire s_dadda_cska12_u_cska22_fa4_and0;
  wire s_dadda_cska12_u_cska22_fa4_xor1;
  wire s_dadda_cska12_u_cska22_fa4_and1;
  wire s_dadda_cska12_u_cska22_fa4_or0;
  wire s_dadda_cska12_u_cska22_xor6;
  wire s_dadda_cska12_u_cska22_fa5_xor0;
  wire s_dadda_cska12_u_cska22_fa5_and0;
  wire s_dadda_cska12_u_cska22_fa5_xor1;
  wire s_dadda_cska12_u_cska22_fa5_and1;
  wire s_dadda_cska12_u_cska22_fa5_or0;
  wire s_dadda_cska12_u_cska22_xor7;
  wire s_dadda_cska12_u_cska22_fa6_xor0;
  wire s_dadda_cska12_u_cska22_fa6_and0;
  wire s_dadda_cska12_u_cska22_fa6_xor1;
  wire s_dadda_cska12_u_cska22_fa6_and1;
  wire s_dadda_cska12_u_cska22_fa6_or0;
  wire s_dadda_cska12_u_cska22_and_propagate13;
  wire s_dadda_cska12_u_cska22_and_propagate14;
  wire s_dadda_cska12_u_cska22_and_propagate15;
  wire s_dadda_cska12_u_cska22_mux2to11_and0;
  wire s_dadda_cska12_u_cska22_mux2to11_not0;
  wire s_dadda_cska12_u_cska22_mux2to11_and1;
  wire s_dadda_cska12_u_cska22_mux2to11_xor0;
  wire s_dadda_cska12_u_cska22_xor8;
  wire s_dadda_cska12_u_cska22_fa7_xor0;
  wire s_dadda_cska12_u_cska22_fa7_and0;
  wire s_dadda_cska12_u_cska22_fa7_xor1;
  wire s_dadda_cska12_u_cska22_fa7_and1;
  wire s_dadda_cska12_u_cska22_fa7_or0;
  wire s_dadda_cska12_u_cska22_xor9;
  wire s_dadda_cska12_u_cska22_fa8_xor0;
  wire s_dadda_cska12_u_cska22_fa8_and0;
  wire s_dadda_cska12_u_cska22_fa8_xor1;
  wire s_dadda_cska12_u_cska22_fa8_and1;
  wire s_dadda_cska12_u_cska22_fa8_or0;
  wire s_dadda_cska12_u_cska22_xor10;
  wire s_dadda_cska12_u_cska22_fa9_xor0;
  wire s_dadda_cska12_u_cska22_fa9_and0;
  wire s_dadda_cska12_u_cska22_fa9_xor1;
  wire s_dadda_cska12_u_cska22_fa9_and1;
  wire s_dadda_cska12_u_cska22_fa9_or0;
  wire s_dadda_cska12_u_cska22_xor11;
  wire s_dadda_cska12_u_cska22_fa10_xor0;
  wire s_dadda_cska12_u_cska22_fa10_and0;
  wire s_dadda_cska12_u_cska22_fa10_xor1;
  wire s_dadda_cska12_u_cska22_fa10_and1;
  wire s_dadda_cska12_u_cska22_fa10_or0;
  wire s_dadda_cska12_u_cska22_and_propagate26;
  wire s_dadda_cska12_u_cska22_and_propagate27;
  wire s_dadda_cska12_u_cska22_and_propagate28;
  wire s_dadda_cska12_u_cska22_mux2to12_and0;
  wire s_dadda_cska12_u_cska22_mux2to12_not0;
  wire s_dadda_cska12_u_cska22_mux2to12_and1;
  wire s_dadda_cska12_u_cska22_mux2to12_xor0;
  wire s_dadda_cska12_u_cska22_xor12;
  wire s_dadda_cska12_u_cska22_fa11_xor0;
  wire s_dadda_cska12_u_cska22_fa11_and0;
  wire s_dadda_cska12_u_cska22_fa11_xor1;
  wire s_dadda_cska12_u_cska22_fa11_and1;
  wire s_dadda_cska12_u_cska22_fa11_or0;
  wire s_dadda_cska12_u_cska22_xor13;
  wire s_dadda_cska12_u_cska22_fa12_xor0;
  wire s_dadda_cska12_u_cska22_fa12_and0;
  wire s_dadda_cska12_u_cska22_fa12_xor1;
  wire s_dadda_cska12_u_cska22_fa12_and1;
  wire s_dadda_cska12_u_cska22_fa12_or0;
  wire s_dadda_cska12_u_cska22_xor14;
  wire s_dadda_cska12_u_cska22_fa13_xor0;
  wire s_dadda_cska12_u_cska22_fa13_and0;
  wire s_dadda_cska12_u_cska22_fa13_xor1;
  wire s_dadda_cska12_u_cska22_fa13_and1;
  wire s_dadda_cska12_u_cska22_fa13_or0;
  wire s_dadda_cska12_u_cska22_xor15;
  wire s_dadda_cska12_u_cska22_fa14_xor0;
  wire s_dadda_cska12_u_cska22_fa14_and0;
  wire s_dadda_cska12_u_cska22_fa14_xor1;
  wire s_dadda_cska12_u_cska22_fa14_and1;
  wire s_dadda_cska12_u_cska22_fa14_or0;
  wire s_dadda_cska12_u_cska22_and_propagate39;
  wire s_dadda_cska12_u_cska22_and_propagate310;
  wire s_dadda_cska12_u_cska22_and_propagate311;
  wire s_dadda_cska12_u_cska22_mux2to13_and0;
  wire s_dadda_cska12_u_cska22_mux2to13_not0;
  wire s_dadda_cska12_u_cska22_mux2to13_and1;
  wire s_dadda_cska12_u_cska22_mux2to13_xor0;
  wire s_dadda_cska12_u_cska22_xor16;
  wire s_dadda_cska12_u_cska22_fa15_xor0;
  wire s_dadda_cska12_u_cska22_fa15_and0;
  wire s_dadda_cska12_u_cska22_fa15_xor1;
  wire s_dadda_cska12_u_cska22_fa15_and1;
  wire s_dadda_cska12_u_cska22_fa15_or0;
  wire s_dadda_cska12_u_cska22_xor17;
  wire s_dadda_cska12_u_cska22_fa16_xor0;
  wire s_dadda_cska12_u_cska22_fa16_and0;
  wire s_dadda_cska12_u_cska22_fa16_xor1;
  wire s_dadda_cska12_u_cska22_fa16_and1;
  wire s_dadda_cska12_u_cska22_fa16_or0;
  wire s_dadda_cska12_u_cska22_xor18;
  wire s_dadda_cska12_u_cska22_fa17_xor0;
  wire s_dadda_cska12_u_cska22_fa17_and0;
  wire s_dadda_cska12_u_cska22_fa17_xor1;
  wire s_dadda_cska12_u_cska22_fa17_and1;
  wire s_dadda_cska12_u_cska22_fa17_or0;
  wire s_dadda_cska12_u_cska22_xor19;
  wire s_dadda_cska12_u_cska22_fa18_xor0;
  wire s_dadda_cska12_u_cska22_fa18_and0;
  wire s_dadda_cska12_u_cska22_fa18_xor1;
  wire s_dadda_cska12_u_cska22_fa18_and1;
  wire s_dadda_cska12_u_cska22_fa18_or0;
  wire s_dadda_cska12_u_cska22_and_propagate412;
  wire s_dadda_cska12_u_cska22_and_propagate413;
  wire s_dadda_cska12_u_cska22_and_propagate414;
  wire s_dadda_cska12_u_cska22_mux2to14_and0;
  wire s_dadda_cska12_u_cska22_mux2to14_not0;
  wire s_dadda_cska12_u_cska22_mux2to14_and1;
  wire s_dadda_cska12_u_cska22_mux2to14_xor0;
  wire s_dadda_cska12_u_cska22_xor20;
  wire s_dadda_cska12_u_cska22_fa19_xor0;
  wire s_dadda_cska12_u_cska22_fa19_and0;
  wire s_dadda_cska12_u_cska22_fa19_xor1;
  wire s_dadda_cska12_u_cska22_fa19_and1;
  wire s_dadda_cska12_u_cska22_fa19_or0;
  wire s_dadda_cska12_u_cska22_xor21;
  wire s_dadda_cska12_u_cska22_fa20_xor0;
  wire s_dadda_cska12_u_cska22_fa20_and0;
  wire s_dadda_cska12_u_cska22_fa20_xor1;
  wire s_dadda_cska12_u_cska22_fa20_and1;
  wire s_dadda_cska12_u_cska22_fa20_or0;
  wire s_dadda_cska12_u_cska22_and_propagate515;
  wire s_dadda_cska12_u_cska22_mux2to15_and0;
  wire s_dadda_cska12_u_cska22_mux2to15_not0;
  wire s_dadda_cska12_u_cska22_mux2to15_and1;
  wire s_dadda_cska12_u_cska22_mux2to15_xor0;
  wire s_dadda_cska12_xor0;

  assign s_dadda_cska12_and_9_0 = a[9] & b[0];
  assign s_dadda_cska12_and_8_1 = a[8] & b[1];
  assign s_dadda_cska12_ha0_xor0 = s_dadda_cska12_and_9_0 ^ s_dadda_cska12_and_8_1;
  assign s_dadda_cska12_ha0_and0 = s_dadda_cska12_and_9_0 & s_dadda_cska12_and_8_1;
  assign s_dadda_cska12_and_10_0 = a[10] & b[0];
  assign s_dadda_cska12_and_9_1 = a[9] & b[1];
  assign s_dadda_cska12_fa0_xor0 = s_dadda_cska12_ha0_and0 ^ s_dadda_cska12_and_10_0;
  assign s_dadda_cska12_fa0_and0 = s_dadda_cska12_ha0_and0 & s_dadda_cska12_and_10_0;
  assign s_dadda_cska12_fa0_xor1 = s_dadda_cska12_fa0_xor0 ^ s_dadda_cska12_and_9_1;
  assign s_dadda_cska12_fa0_and1 = s_dadda_cska12_fa0_xor0 & s_dadda_cska12_and_9_1;
  assign s_dadda_cska12_fa0_or0 = s_dadda_cska12_fa0_and0 | s_dadda_cska12_fa0_and1;
  assign s_dadda_cska12_and_8_2 = a[8] & b[2];
  assign s_dadda_cska12_and_7_3 = a[7] & b[3];
  assign s_dadda_cska12_ha1_xor0 = s_dadda_cska12_and_8_2 ^ s_dadda_cska12_and_7_3;
  assign s_dadda_cska12_ha1_and0 = s_dadda_cska12_and_8_2 & s_dadda_cska12_and_7_3;
  assign s_dadda_cska12_nand_11_0 = ~(a[11] & b[0]);
  assign s_dadda_cska12_fa1_xor0 = s_dadda_cska12_ha1_and0 ^ s_dadda_cska12_fa0_or0;
  assign s_dadda_cska12_fa1_and0 = s_dadda_cska12_ha1_and0 & s_dadda_cska12_fa0_or0;
  assign s_dadda_cska12_fa1_xor1 = s_dadda_cska12_fa1_xor0 ^ s_dadda_cska12_nand_11_0;
  assign s_dadda_cska12_fa1_and1 = s_dadda_cska12_fa1_xor0 & s_dadda_cska12_nand_11_0;
  assign s_dadda_cska12_fa1_or0 = s_dadda_cska12_fa1_and0 | s_dadda_cska12_fa1_and1;
  assign s_dadda_cska12_and_10_1 = a[10] & b[1];
  assign s_dadda_cska12_and_9_2 = a[9] & b[2];
  assign s_dadda_cska12_and_8_3 = a[8] & b[3];
  assign s_dadda_cska12_fa2_xor0 = s_dadda_cska12_and_10_1 ^ s_dadda_cska12_and_9_2;
  assign s_dadda_cska12_fa2_and0 = s_dadda_cska12_and_10_1 & s_dadda_cska12_and_9_2;
  assign s_dadda_cska12_fa2_xor1 = s_dadda_cska12_fa2_xor0 ^ s_dadda_cska12_and_8_3;
  assign s_dadda_cska12_fa2_and1 = s_dadda_cska12_fa2_xor0 & s_dadda_cska12_and_8_3;
  assign s_dadda_cska12_fa2_or0 = s_dadda_cska12_fa2_and0 | s_dadda_cska12_fa2_and1;
  assign s_dadda_cska12_and_7_4 = a[7] & b[4];
  assign s_dadda_cska12_and_6_5 = a[6] & b[5];
  assign s_dadda_cska12_ha2_xor0 = s_dadda_cska12_and_7_4 ^ s_dadda_cska12_and_6_5;
  assign s_dadda_cska12_ha2_and0 = s_dadda_cska12_and_7_4 & s_dadda_cska12_and_6_5;
  assign s_dadda_cska12_fa3_xor0 = s_dadda_cska12_ha2_and0 ^ s_dadda_cska12_fa2_or0;
  assign s_dadda_cska12_fa3_and0 = s_dadda_cska12_ha2_and0 & s_dadda_cska12_fa2_or0;
  assign s_dadda_cska12_fa3_xor1 = s_dadda_cska12_fa3_xor0 ^ s_dadda_cska12_fa1_or0;
  assign s_dadda_cska12_fa3_and1 = s_dadda_cska12_fa3_xor0 & s_dadda_cska12_fa1_or0;
  assign s_dadda_cska12_fa3_or0 = s_dadda_cska12_fa3_and0 | s_dadda_cska12_fa3_and1;
  assign s_dadda_cska12_nand_11_1 = ~(a[11] & b[1]);
  assign s_dadda_cska12_and_10_2 = a[10] & b[2];
  assign s_dadda_cska12_fa4_xor0 = ~s_dadda_cska12_nand_11_1;
  assign s_dadda_cska12_fa4_xor1 = s_dadda_cska12_fa4_xor0 ^ s_dadda_cska12_and_10_2;
  assign s_dadda_cska12_fa4_and1 = s_dadda_cska12_fa4_xor0 & s_dadda_cska12_and_10_2;
  assign s_dadda_cska12_fa4_or0 = s_dadda_cska12_nand_11_1 | s_dadda_cska12_fa4_and1;
  assign s_dadda_cska12_and_9_3 = a[9] & b[3];
  assign s_dadda_cska12_and_8_4 = a[8] & b[4];
  assign s_dadda_cska12_and_7_5 = a[7] & b[5];
  assign s_dadda_cska12_fa5_xor0 = s_dadda_cska12_and_9_3 ^ s_dadda_cska12_and_8_4;
  assign s_dadda_cska12_fa5_and0 = s_dadda_cska12_and_9_3 & s_dadda_cska12_and_8_4;
  assign s_dadda_cska12_fa5_xor1 = s_dadda_cska12_fa5_xor0 ^ s_dadda_cska12_and_7_5;
  assign s_dadda_cska12_fa5_and1 = s_dadda_cska12_fa5_xor0 & s_dadda_cska12_and_7_5;
  assign s_dadda_cska12_fa5_or0 = s_dadda_cska12_fa5_and0 | s_dadda_cska12_fa5_and1;
  assign s_dadda_cska12_fa6_xor0 = s_dadda_cska12_fa5_or0 ^ s_dadda_cska12_fa4_or0;
  assign s_dadda_cska12_fa6_and0 = s_dadda_cska12_fa5_or0 & s_dadda_cska12_fa4_or0;
  assign s_dadda_cska12_fa6_xor1 = s_dadda_cska12_fa6_xor0 ^ s_dadda_cska12_fa3_or0;
  assign s_dadda_cska12_fa6_and1 = s_dadda_cska12_fa6_xor0 & s_dadda_cska12_fa3_or0;
  assign s_dadda_cska12_fa6_or0 = s_dadda_cska12_fa6_and0 | s_dadda_cska12_fa6_and1;
  assign s_dadda_cska12_nand_11_2 = ~(a[11] & b[2]);
  assign s_dadda_cska12_and_10_3 = a[10] & b[3];
  assign s_dadda_cska12_and_9_4 = a[9] & b[4];
  assign s_dadda_cska12_fa7_xor0 = s_dadda_cska12_nand_11_2 ^ s_dadda_cska12_and_10_3;
  assign s_dadda_cska12_fa7_and0 = s_dadda_cska12_nand_11_2 & s_dadda_cska12_and_10_3;
  assign s_dadda_cska12_fa7_xor1 = s_dadda_cska12_fa7_xor0 ^ s_dadda_cska12_and_9_4;
  assign s_dadda_cska12_fa7_and1 = s_dadda_cska12_fa7_xor0 & s_dadda_cska12_and_9_4;
  assign s_dadda_cska12_fa7_or0 = s_dadda_cska12_fa7_and0 | s_dadda_cska12_fa7_and1;
  assign s_dadda_cska12_nand_11_3 = ~(a[11] & b[3]);
  assign s_dadda_cska12_fa8_xor0 = s_dadda_cska12_fa7_or0 ^ s_dadda_cska12_fa6_or0;
  assign s_dadda_cska12_fa8_and0 = s_dadda_cska12_fa7_or0 & s_dadda_cska12_fa6_or0;
  assign s_dadda_cska12_fa8_xor1 = s_dadda_cska12_fa8_xor0 ^ s_dadda_cska12_nand_11_3;
  assign s_dadda_cska12_fa8_and1 = s_dadda_cska12_fa8_xor0 & s_dadda_cska12_nand_11_3;
  assign s_dadda_cska12_fa8_or0 = s_dadda_cska12_fa8_and0 | s_dadda_cska12_fa8_and1;
  assign s_dadda_cska12_and_4_0 = a[4] & b[0];
  assign s_dadda_cska12_and_3_1 = a[3] & b[1];
  assign s_dadda_cska12_ha3_xor0 = s_dadda_cska12_and_4_0 ^ s_dadda_cska12_and_3_1;
  assign s_dadda_cska12_ha3_and0 = s_dadda_cska12_and_4_0 & s_dadda_cska12_and_3_1;
  assign s_dadda_cska12_and_5_0 = a[5] & b[0];
  assign s_dadda_cska12_and_4_1 = a[4] & b[1];
  assign s_dadda_cska12_fa9_xor0 = s_dadda_cska12_ha3_and0 ^ s_dadda_cska12_and_5_0;
  assign s_dadda_cska12_fa9_and0 = s_dadda_cska12_ha3_and0 & s_dadda_cska12_and_5_0;
  assign s_dadda_cska12_fa9_xor1 = s_dadda_cska12_fa9_xor0 ^ s_dadda_cska12_and_4_1;
  assign s_dadda_cska12_fa9_and1 = s_dadda_cska12_fa9_xor0 & s_dadda_cska12_and_4_1;
  assign s_dadda_cska12_fa9_or0 = s_dadda_cska12_fa9_and0 | s_dadda_cska12_fa9_and1;
  assign s_dadda_cska12_and_3_2 = a[3] & b[2];
  assign s_dadda_cska12_and_2_3 = a[2] & b[3];
  assign s_dadda_cska12_ha4_xor0 = s_dadda_cska12_and_3_2 ^ s_dadda_cska12_and_2_3;
  assign s_dadda_cska12_ha4_and0 = s_dadda_cska12_and_3_2 & s_dadda_cska12_and_2_3;
  assign s_dadda_cska12_and_6_0 = a[6] & b[0];
  assign s_dadda_cska12_fa10_xor0 = s_dadda_cska12_ha4_and0 ^ s_dadda_cska12_fa9_or0;
  assign s_dadda_cska12_fa10_and0 = s_dadda_cska12_ha4_and0 & s_dadda_cska12_fa9_or0;
  assign s_dadda_cska12_fa10_xor1 = s_dadda_cska12_fa10_xor0 ^ s_dadda_cska12_and_6_0;
  assign s_dadda_cska12_fa10_and1 = s_dadda_cska12_fa10_xor0 & s_dadda_cska12_and_6_0;
  assign s_dadda_cska12_fa10_or0 = s_dadda_cska12_fa10_and0 | s_dadda_cska12_fa10_and1;
  assign s_dadda_cska12_and_5_1 = a[5] & b[1];
  assign s_dadda_cska12_and_4_2 = a[4] & b[2];
  assign s_dadda_cska12_and_3_3 = a[3] & b[3];
  assign s_dadda_cska12_fa11_xor0 = s_dadda_cska12_and_5_1 ^ s_dadda_cska12_and_4_2;
  assign s_dadda_cska12_fa11_and0 = s_dadda_cska12_and_5_1 & s_dadda_cska12_and_4_2;
  assign s_dadda_cska12_fa11_xor1 = s_dadda_cska12_fa11_xor0 ^ s_dadda_cska12_and_3_3;
  assign s_dadda_cska12_fa11_and1 = s_dadda_cska12_fa11_xor0 & s_dadda_cska12_and_3_3;
  assign s_dadda_cska12_fa11_or0 = s_dadda_cska12_fa11_and0 | s_dadda_cska12_fa11_and1;
  assign s_dadda_cska12_and_2_4 = a[2] & b[4];
  assign s_dadda_cska12_and_1_5 = a[1] & b[5];
  assign s_dadda_cska12_ha5_xor0 = s_dadda_cska12_and_2_4 ^ s_dadda_cska12_and_1_5;
  assign s_dadda_cska12_ha5_and0 = s_dadda_cska12_and_2_4 & s_dadda_cska12_and_1_5;
  assign s_dadda_cska12_fa12_xor0 = s_dadda_cska12_ha5_and0 ^ s_dadda_cska12_fa11_or0;
  assign s_dadda_cska12_fa12_and0 = s_dadda_cska12_ha5_and0 & s_dadda_cska12_fa11_or0;
  assign s_dadda_cska12_fa12_xor1 = s_dadda_cska12_fa12_xor0 ^ s_dadda_cska12_fa10_or0;
  assign s_dadda_cska12_fa12_and1 = s_dadda_cska12_fa12_xor0 & s_dadda_cska12_fa10_or0;
  assign s_dadda_cska12_fa12_or0 = s_dadda_cska12_fa12_and0 | s_dadda_cska12_fa12_and1;
  assign s_dadda_cska12_and_7_0 = a[7] & b[0];
  assign s_dadda_cska12_and_6_1 = a[6] & b[1];
  assign s_dadda_cska12_and_5_2 = a[5] & b[2];
  assign s_dadda_cska12_fa13_xor0 = s_dadda_cska12_and_7_0 ^ s_dadda_cska12_and_6_1;
  assign s_dadda_cska12_fa13_and0 = s_dadda_cska12_and_7_0 & s_dadda_cska12_and_6_1;
  assign s_dadda_cska12_fa13_xor1 = s_dadda_cska12_fa13_xor0 ^ s_dadda_cska12_and_5_2;
  assign s_dadda_cska12_fa13_and1 = s_dadda_cska12_fa13_xor0 & s_dadda_cska12_and_5_2;
  assign s_dadda_cska12_fa13_or0 = s_dadda_cska12_fa13_and0 | s_dadda_cska12_fa13_and1;
  assign s_dadda_cska12_and_4_3 = a[4] & b[3];
  assign s_dadda_cska12_and_3_4 = a[3] & b[4];
  assign s_dadda_cska12_and_2_5 = a[2] & b[5];
  assign s_dadda_cska12_fa14_xor0 = s_dadda_cska12_and_4_3 ^ s_dadda_cska12_and_3_4;
  assign s_dadda_cska12_fa14_and0 = s_dadda_cska12_and_4_3 & s_dadda_cska12_and_3_4;
  assign s_dadda_cska12_fa14_xor1 = s_dadda_cska12_fa14_xor0 ^ s_dadda_cska12_and_2_5;
  assign s_dadda_cska12_fa14_and1 = s_dadda_cska12_fa14_xor0 & s_dadda_cska12_and_2_5;
  assign s_dadda_cska12_fa14_or0 = s_dadda_cska12_fa14_and0 | s_dadda_cska12_fa14_and1;
  assign s_dadda_cska12_and_1_6 = a[1] & b[6];
  assign s_dadda_cska12_and_0_7 = a[0] & b[7];
  assign s_dadda_cska12_ha6_xor0 = s_dadda_cska12_and_1_6 ^ s_dadda_cska12_and_0_7;
  assign s_dadda_cska12_ha6_and0 = s_dadda_cska12_and_1_6 & s_dadda_cska12_and_0_7;
  assign s_dadda_cska12_fa15_xor0 = s_dadda_cska12_ha6_and0 ^ s_dadda_cska12_fa14_or0;
  assign s_dadda_cska12_fa15_and0 = s_dadda_cska12_ha6_and0 & s_dadda_cska12_fa14_or0;
  assign s_dadda_cska12_fa15_xor1 = s_dadda_cska12_fa15_xor0 ^ s_dadda_cska12_fa13_or0;
  assign s_dadda_cska12_fa15_and1 = s_dadda_cska12_fa15_xor0 & s_dadda_cska12_fa13_or0;
  assign s_dadda_cska12_fa15_or0 = s_dadda_cska12_fa15_and0 | s_dadda_cska12_fa15_and1;
  assign s_dadda_cska12_and_8_0 = a[8] & b[0];
  assign s_dadda_cska12_and_7_1 = a[7] & b[1];
  assign s_dadda_cska12_fa16_xor0 = s_dadda_cska12_fa12_or0 ^ s_dadda_cska12_and_8_0;
  assign s_dadda_cska12_fa16_and0 = s_dadda_cska12_fa12_or0 & s_dadda_cska12_and_8_0;
  assign s_dadda_cska12_fa16_xor1 = s_dadda_cska12_fa16_xor0 ^ s_dadda_cska12_and_7_1;
  assign s_dadda_cska12_fa16_and1 = s_dadda_cska12_fa16_xor0 & s_dadda_cska12_and_7_1;
  assign s_dadda_cska12_fa16_or0 = s_dadda_cska12_fa16_and0 | s_dadda_cska12_fa16_and1;
  assign s_dadda_cska12_and_6_2 = a[6] & b[2];
  assign s_dadda_cska12_and_5_3 = a[5] & b[3];
  assign s_dadda_cska12_and_4_4 = a[4] & b[4];
  assign s_dadda_cska12_fa17_xor0 = s_dadda_cska12_and_6_2 ^ s_dadda_cska12_and_5_3;
  assign s_dadda_cska12_fa17_and0 = s_dadda_cska12_and_6_2 & s_dadda_cska12_and_5_3;
  assign s_dadda_cska12_fa17_xor1 = s_dadda_cska12_fa17_xor0 ^ s_dadda_cska12_and_4_4;
  assign s_dadda_cska12_fa17_and1 = s_dadda_cska12_fa17_xor0 & s_dadda_cska12_and_4_4;
  assign s_dadda_cska12_fa17_or0 = s_dadda_cska12_fa17_and0 | s_dadda_cska12_fa17_and1;
  assign s_dadda_cska12_and_3_5 = a[3] & b[5];
  assign s_dadda_cska12_and_2_6 = a[2] & b[6];
  assign s_dadda_cska12_and_1_7 = a[1] & b[7];
  assign s_dadda_cska12_fa18_xor0 = s_dadda_cska12_and_3_5 ^ s_dadda_cska12_and_2_6;
  assign s_dadda_cska12_fa18_and0 = s_dadda_cska12_and_3_5 & s_dadda_cska12_and_2_6;
  assign s_dadda_cska12_fa18_xor1 = s_dadda_cska12_fa18_xor0 ^ s_dadda_cska12_and_1_7;
  assign s_dadda_cska12_fa18_and1 = s_dadda_cska12_fa18_xor0 & s_dadda_cska12_and_1_7;
  assign s_dadda_cska12_fa18_or0 = s_dadda_cska12_fa18_and0 | s_dadda_cska12_fa18_and1;
  assign s_dadda_cska12_and_0_8 = a[0] & b[8];
  assign s_dadda_cska12_ha7_xor0 = s_dadda_cska12_and_0_8 ^ s_dadda_cska12_fa15_xor1;
  assign s_dadda_cska12_ha7_and0 = s_dadda_cska12_and_0_8 & s_dadda_cska12_fa15_xor1;
  assign s_dadda_cska12_fa19_xor0 = s_dadda_cska12_ha7_and0 ^ s_dadda_cska12_fa18_or0;
  assign s_dadda_cska12_fa19_and0 = s_dadda_cska12_ha7_and0 & s_dadda_cska12_fa18_or0;
  assign s_dadda_cska12_fa19_xor1 = s_dadda_cska12_fa19_xor0 ^ s_dadda_cska12_fa17_or0;
  assign s_dadda_cska12_fa19_and1 = s_dadda_cska12_fa19_xor0 & s_dadda_cska12_fa17_or0;
  assign s_dadda_cska12_fa19_or0 = s_dadda_cska12_fa19_and0 | s_dadda_cska12_fa19_and1;
  assign s_dadda_cska12_and_7_2 = a[7] & b[2];
  assign s_dadda_cska12_fa20_xor0 = s_dadda_cska12_fa16_or0 ^ s_dadda_cska12_fa15_or0;
  assign s_dadda_cska12_fa20_and0 = s_dadda_cska12_fa16_or0 & s_dadda_cska12_fa15_or0;
  assign s_dadda_cska12_fa20_xor1 = s_dadda_cska12_fa20_xor0 ^ s_dadda_cska12_and_7_2;
  assign s_dadda_cska12_fa20_and1 = s_dadda_cska12_fa20_xor0 & s_dadda_cska12_and_7_2;
  assign s_dadda_cska12_fa20_or0 = s_dadda_cska12_fa20_and0 | s_dadda_cska12_fa20_and1;
  assign s_dadda_cska12_and_6_3 = a[6] & b[3];
  assign s_dadda_cska12_and_5_4 = a[5] & b[4];
  assign s_dadda_cska12_and_4_5 = a[4] & b[5];
  assign s_dadda_cska12_fa21_xor0 = s_dadda_cska12_and_6_3 ^ s_dadda_cska12_and_5_4;
  assign s_dadda_cska12_fa21_and0 = s_dadda_cska12_and_6_3 & s_dadda_cska12_and_5_4;
  assign s_dadda_cska12_fa21_xor1 = s_dadda_cska12_fa21_xor0 ^ s_dadda_cska12_and_4_5;
  assign s_dadda_cska12_fa21_and1 = s_dadda_cska12_fa21_xor0 & s_dadda_cska12_and_4_5;
  assign s_dadda_cska12_fa21_or0 = s_dadda_cska12_fa21_and0 | s_dadda_cska12_fa21_and1;
  assign s_dadda_cska12_and_3_6 = a[3] & b[6];
  assign s_dadda_cska12_and_2_7 = a[2] & b[7];
  assign s_dadda_cska12_and_1_8 = a[1] & b[8];
  assign s_dadda_cska12_fa22_xor0 = s_dadda_cska12_and_3_6 ^ s_dadda_cska12_and_2_7;
  assign s_dadda_cska12_fa22_and0 = s_dadda_cska12_and_3_6 & s_dadda_cska12_and_2_7;
  assign s_dadda_cska12_fa22_xor1 = s_dadda_cska12_fa22_xor0 ^ s_dadda_cska12_and_1_8;
  assign s_dadda_cska12_fa22_and1 = s_dadda_cska12_fa22_xor0 & s_dadda_cska12_and_1_8;
  assign s_dadda_cska12_fa22_or0 = s_dadda_cska12_fa22_and0 | s_dadda_cska12_fa22_and1;
  assign s_dadda_cska12_and_0_9 = a[0] & b[9];
  assign s_dadda_cska12_fa23_xor0 = s_dadda_cska12_and_0_9 ^ s_dadda_cska12_ha0_xor0;
  assign s_dadda_cska12_fa23_and0 = s_dadda_cska12_and_0_9 & s_dadda_cska12_ha0_xor0;
  assign s_dadda_cska12_fa23_xor1 = s_dadda_cska12_fa23_xor0 ^ s_dadda_cska12_fa19_xor1;
  assign s_dadda_cska12_fa23_and1 = s_dadda_cska12_fa23_xor0 & s_dadda_cska12_fa19_xor1;
  assign s_dadda_cska12_fa23_or0 = s_dadda_cska12_fa23_and0 | s_dadda_cska12_fa23_and1;
  assign s_dadda_cska12_fa24_xor0 = s_dadda_cska12_fa23_or0 ^ s_dadda_cska12_fa22_or0;
  assign s_dadda_cska12_fa24_and0 = s_dadda_cska12_fa23_or0 & s_dadda_cska12_fa22_or0;
  assign s_dadda_cska12_fa24_xor1 = s_dadda_cska12_fa24_xor0 ^ s_dadda_cska12_fa21_or0;
  assign s_dadda_cska12_fa24_and1 = s_dadda_cska12_fa24_xor0 & s_dadda_cska12_fa21_or0;
  assign s_dadda_cska12_fa24_or0 = s_dadda_cska12_fa24_and0 | s_dadda_cska12_fa24_and1;
  assign s_dadda_cska12_and_6_4 = a[6] & b[4];
  assign s_dadda_cska12_fa25_xor0 = s_dadda_cska12_fa20_or0 ^ s_dadda_cska12_fa19_or0;
  assign s_dadda_cska12_fa25_and0 = s_dadda_cska12_fa20_or0 & s_dadda_cska12_fa19_or0;
  assign s_dadda_cska12_fa25_xor1 = s_dadda_cska12_fa25_xor0 ^ s_dadda_cska12_and_6_4;
  assign s_dadda_cska12_fa25_and1 = s_dadda_cska12_fa25_xor0 & s_dadda_cska12_and_6_4;
  assign s_dadda_cska12_fa25_or0 = s_dadda_cska12_fa25_and0 | s_dadda_cska12_fa25_and1;
  assign s_dadda_cska12_and_5_5 = a[5] & b[5];
  assign s_dadda_cska12_and_4_6 = a[4] & b[6];
  assign s_dadda_cska12_and_3_7 = a[3] & b[7];
  assign s_dadda_cska12_fa26_xor0 = s_dadda_cska12_and_5_5 ^ s_dadda_cska12_and_4_6;
  assign s_dadda_cska12_fa26_and0 = s_dadda_cska12_and_5_5 & s_dadda_cska12_and_4_6;
  assign s_dadda_cska12_fa26_xor1 = s_dadda_cska12_fa26_xor0 ^ s_dadda_cska12_and_3_7;
  assign s_dadda_cska12_fa26_and1 = s_dadda_cska12_fa26_xor0 & s_dadda_cska12_and_3_7;
  assign s_dadda_cska12_fa26_or0 = s_dadda_cska12_fa26_and0 | s_dadda_cska12_fa26_and1;
  assign s_dadda_cska12_and_2_8 = a[2] & b[8];
  assign s_dadda_cska12_and_1_9 = a[1] & b[9];
  assign s_dadda_cska12_and_0_10 = a[0] & b[10];
  assign s_dadda_cska12_fa27_xor0 = s_dadda_cska12_and_2_8 ^ s_dadda_cska12_and_1_9;
  assign s_dadda_cska12_fa27_and0 = s_dadda_cska12_and_2_8 & s_dadda_cska12_and_1_9;
  assign s_dadda_cska12_fa27_xor1 = s_dadda_cska12_fa27_xor0 ^ s_dadda_cska12_and_0_10;
  assign s_dadda_cska12_fa27_and1 = s_dadda_cska12_fa27_xor0 & s_dadda_cska12_and_0_10;
  assign s_dadda_cska12_fa27_or0 = s_dadda_cska12_fa27_and0 | s_dadda_cska12_fa27_and1;
  assign s_dadda_cska12_fa28_xor0 = s_dadda_cska12_fa0_xor1 ^ s_dadda_cska12_ha1_xor0;
  assign s_dadda_cska12_fa28_and0 = s_dadda_cska12_fa0_xor1 & s_dadda_cska12_ha1_xor0;
  assign s_dadda_cska12_fa28_xor1 = s_dadda_cska12_fa28_xor0 ^ s_dadda_cska12_fa24_xor1;
  assign s_dadda_cska12_fa28_and1 = s_dadda_cska12_fa28_xor0 & s_dadda_cska12_fa24_xor1;
  assign s_dadda_cska12_fa28_or0 = s_dadda_cska12_fa28_and0 | s_dadda_cska12_fa28_and1;
  assign s_dadda_cska12_fa29_xor0 = s_dadda_cska12_fa28_or0 ^ s_dadda_cska12_fa27_or0;
  assign s_dadda_cska12_fa29_and0 = s_dadda_cska12_fa28_or0 & s_dadda_cska12_fa27_or0;
  assign s_dadda_cska12_fa29_xor1 = s_dadda_cska12_fa29_xor0 ^ s_dadda_cska12_fa26_or0;
  assign s_dadda_cska12_fa29_and1 = s_dadda_cska12_fa29_xor0 & s_dadda_cska12_fa26_or0;
  assign s_dadda_cska12_fa29_or0 = s_dadda_cska12_fa29_and0 | s_dadda_cska12_fa29_and1;
  assign s_dadda_cska12_and_5_6 = a[5] & b[6];
  assign s_dadda_cska12_fa30_xor0 = s_dadda_cska12_fa25_or0 ^ s_dadda_cska12_fa24_or0;
  assign s_dadda_cska12_fa30_and0 = s_dadda_cska12_fa25_or0 & s_dadda_cska12_fa24_or0;
  assign s_dadda_cska12_fa30_xor1 = s_dadda_cska12_fa30_xor0 ^ s_dadda_cska12_and_5_6;
  assign s_dadda_cska12_fa30_and1 = s_dadda_cska12_fa30_xor0 & s_dadda_cska12_and_5_6;
  assign s_dadda_cska12_fa30_or0 = s_dadda_cska12_fa30_and0 | s_dadda_cska12_fa30_and1;
  assign s_dadda_cska12_and_4_7 = a[4] & b[7];
  assign s_dadda_cska12_and_3_8 = a[3] & b[8];
  assign s_dadda_cska12_and_2_9 = a[2] & b[9];
  assign s_dadda_cska12_fa31_xor0 = s_dadda_cska12_and_4_7 ^ s_dadda_cska12_and_3_8;
  assign s_dadda_cska12_fa31_and0 = s_dadda_cska12_and_4_7 & s_dadda_cska12_and_3_8;
  assign s_dadda_cska12_fa31_xor1 = s_dadda_cska12_fa31_xor0 ^ s_dadda_cska12_and_2_9;
  assign s_dadda_cska12_fa31_and1 = s_dadda_cska12_fa31_xor0 & s_dadda_cska12_and_2_9;
  assign s_dadda_cska12_fa31_or0 = s_dadda_cska12_fa31_and0 | s_dadda_cska12_fa31_and1;
  assign s_dadda_cska12_and_1_10 = a[1] & b[10];
  assign s_dadda_cska12_nand_0_11 = ~(a[0] & b[11]);
  assign s_dadda_cska12_fa32_xor0 = s_dadda_cska12_and_1_10 ^ s_dadda_cska12_nand_0_11;
  assign s_dadda_cska12_fa32_and0 = s_dadda_cska12_and_1_10 & s_dadda_cska12_nand_0_11;
  assign s_dadda_cska12_fa32_xor1 = s_dadda_cska12_fa32_xor0 ^ s_dadda_cska12_fa1_xor1;
  assign s_dadda_cska12_fa32_and1 = s_dadda_cska12_fa32_xor0 & s_dadda_cska12_fa1_xor1;
  assign s_dadda_cska12_fa32_or0 = s_dadda_cska12_fa32_and0 | s_dadda_cska12_fa32_and1;
  assign s_dadda_cska12_fa33_xor0 = s_dadda_cska12_fa2_xor1 ^ s_dadda_cska12_ha2_xor0;
  assign s_dadda_cska12_fa33_and0 = s_dadda_cska12_fa2_xor1 & s_dadda_cska12_ha2_xor0;
  assign s_dadda_cska12_fa33_xor1 = s_dadda_cska12_fa33_xor0 ^ s_dadda_cska12_fa29_xor1;
  assign s_dadda_cska12_fa33_and1 = s_dadda_cska12_fa33_xor0 & s_dadda_cska12_fa29_xor1;
  assign s_dadda_cska12_fa33_or0 = s_dadda_cska12_fa33_and0 | s_dadda_cska12_fa33_and1;
  assign s_dadda_cska12_fa34_xor0 = s_dadda_cska12_fa33_or0 ^ s_dadda_cska12_fa32_or0;
  assign s_dadda_cska12_fa34_and0 = s_dadda_cska12_fa33_or0 & s_dadda_cska12_fa32_or0;
  assign s_dadda_cska12_fa34_xor1 = s_dadda_cska12_fa34_xor0 ^ s_dadda_cska12_fa31_or0;
  assign s_dadda_cska12_fa34_and1 = s_dadda_cska12_fa34_xor0 & s_dadda_cska12_fa31_or0;
  assign s_dadda_cska12_fa34_or0 = s_dadda_cska12_fa34_and0 | s_dadda_cska12_fa34_and1;
  assign s_dadda_cska12_and_6_6 = a[6] & b[6];
  assign s_dadda_cska12_fa35_xor0 = s_dadda_cska12_fa30_or0 ^ s_dadda_cska12_fa29_or0;
  assign s_dadda_cska12_fa35_and0 = s_dadda_cska12_fa30_or0 & s_dadda_cska12_fa29_or0;
  assign s_dadda_cska12_fa35_xor1 = s_dadda_cska12_fa35_xor0 ^ s_dadda_cska12_and_6_6;
  assign s_dadda_cska12_fa35_and1 = s_dadda_cska12_fa35_xor0 & s_dadda_cska12_and_6_6;
  assign s_dadda_cska12_fa35_or0 = s_dadda_cska12_fa35_and0 | s_dadda_cska12_fa35_and1;
  assign s_dadda_cska12_and_5_7 = a[5] & b[7];
  assign s_dadda_cska12_and_4_8 = a[4] & b[8];
  assign s_dadda_cska12_and_3_9 = a[3] & b[9];
  assign s_dadda_cska12_fa36_xor0 = s_dadda_cska12_and_5_7 ^ s_dadda_cska12_and_4_8;
  assign s_dadda_cska12_fa36_and0 = s_dadda_cska12_and_5_7 & s_dadda_cska12_and_4_8;
  assign s_dadda_cska12_fa36_xor1 = s_dadda_cska12_fa36_xor0 ^ s_dadda_cska12_and_3_9;
  assign s_dadda_cska12_fa36_and1 = s_dadda_cska12_fa36_xor0 & s_dadda_cska12_and_3_9;
  assign s_dadda_cska12_fa36_or0 = s_dadda_cska12_fa36_and0 | s_dadda_cska12_fa36_and1;
  assign s_dadda_cska12_and_2_10 = a[2] & b[10];
  assign s_dadda_cska12_nand_1_11 = ~(a[1] & b[11]);
  assign s_dadda_cska12_fa37_xor0 = s_dadda_cska12_and_2_10 ^ s_dadda_cska12_nand_1_11;
  assign s_dadda_cska12_fa37_and0 = s_dadda_cska12_and_2_10 & s_dadda_cska12_nand_1_11;
  assign s_dadda_cska12_fa37_xor1 = s_dadda_cska12_fa37_xor0 ^ s_dadda_cska12_fa3_xor1;
  assign s_dadda_cska12_fa37_and1 = s_dadda_cska12_fa37_xor0 & s_dadda_cska12_fa3_xor1;
  assign s_dadda_cska12_fa37_or0 = s_dadda_cska12_fa37_and0 | s_dadda_cska12_fa37_and1;
  assign s_dadda_cska12_fa38_xor0 = s_dadda_cska12_fa4_xor1 ^ s_dadda_cska12_fa5_xor1;
  assign s_dadda_cska12_fa38_and0 = s_dadda_cska12_fa4_xor1 & s_dadda_cska12_fa5_xor1;
  assign s_dadda_cska12_fa38_xor1 = s_dadda_cska12_fa38_xor0 ^ s_dadda_cska12_fa34_xor1;
  assign s_dadda_cska12_fa38_and1 = s_dadda_cska12_fa38_xor0 & s_dadda_cska12_fa34_xor1;
  assign s_dadda_cska12_fa38_or0 = s_dadda_cska12_fa38_and0 | s_dadda_cska12_fa38_and1;
  assign s_dadda_cska12_fa39_xor0 = s_dadda_cska12_fa38_or0 ^ s_dadda_cska12_fa37_or0;
  assign s_dadda_cska12_fa39_and0 = s_dadda_cska12_fa38_or0 & s_dadda_cska12_fa37_or0;
  assign s_dadda_cska12_fa39_xor1 = s_dadda_cska12_fa39_xor0 ^ s_dadda_cska12_fa36_or0;
  assign s_dadda_cska12_fa39_and1 = s_dadda_cska12_fa39_xor0 & s_dadda_cska12_fa36_or0;
  assign s_dadda_cska12_fa39_or0 = s_dadda_cska12_fa39_and0 | s_dadda_cska12_fa39_and1;
  assign s_dadda_cska12_and_8_5 = a[8] & b[5];
  assign s_dadda_cska12_fa40_xor0 = s_dadda_cska12_fa35_or0 ^ s_dadda_cska12_fa34_or0;
  assign s_dadda_cska12_fa40_and0 = s_dadda_cska12_fa35_or0 & s_dadda_cska12_fa34_or0;
  assign s_dadda_cska12_fa40_xor1 = s_dadda_cska12_fa40_xor0 ^ s_dadda_cska12_and_8_5;
  assign s_dadda_cska12_fa40_and1 = s_dadda_cska12_fa40_xor0 & s_dadda_cska12_and_8_5;
  assign s_dadda_cska12_fa40_or0 = s_dadda_cska12_fa40_and0 | s_dadda_cska12_fa40_and1;
  assign s_dadda_cska12_and_7_6 = a[7] & b[6];
  assign s_dadda_cska12_and_6_7 = a[6] & b[7];
  assign s_dadda_cska12_and_5_8 = a[5] & b[8];
  assign s_dadda_cska12_fa41_xor0 = s_dadda_cska12_and_7_6 ^ s_dadda_cska12_and_6_7;
  assign s_dadda_cska12_fa41_and0 = s_dadda_cska12_and_7_6 & s_dadda_cska12_and_6_7;
  assign s_dadda_cska12_fa41_xor1 = s_dadda_cska12_fa41_xor0 ^ s_dadda_cska12_and_5_8;
  assign s_dadda_cska12_fa41_and1 = s_dadda_cska12_fa41_xor0 & s_dadda_cska12_and_5_8;
  assign s_dadda_cska12_fa41_or0 = s_dadda_cska12_fa41_and0 | s_dadda_cska12_fa41_and1;
  assign s_dadda_cska12_and_4_9 = a[4] & b[9];
  assign s_dadda_cska12_and_3_10 = a[3] & b[10];
  assign s_dadda_cska12_nand_2_11 = ~(a[2] & b[11]);
  assign s_dadda_cska12_fa42_xor0 = s_dadda_cska12_and_4_9 ^ s_dadda_cska12_and_3_10;
  assign s_dadda_cska12_fa42_and0 = s_dadda_cska12_and_4_9 & s_dadda_cska12_and_3_10;
  assign s_dadda_cska12_fa42_xor1 = s_dadda_cska12_fa42_xor0 ^ s_dadda_cska12_nand_2_11;
  assign s_dadda_cska12_fa42_and1 = s_dadda_cska12_fa42_xor0 & s_dadda_cska12_nand_2_11;
  assign s_dadda_cska12_fa42_or0 = s_dadda_cska12_fa42_and0 | s_dadda_cska12_fa42_and1;
  assign s_dadda_cska12_fa43_xor0 = s_dadda_cska12_fa6_xor1 ^ s_dadda_cska12_fa7_xor1;
  assign s_dadda_cska12_fa43_and0 = s_dadda_cska12_fa6_xor1 & s_dadda_cska12_fa7_xor1;
  assign s_dadda_cska12_fa43_xor1 = s_dadda_cska12_fa43_xor0 ^ s_dadda_cska12_fa39_xor1;
  assign s_dadda_cska12_fa43_and1 = s_dadda_cska12_fa43_xor0 & s_dadda_cska12_fa39_xor1;
  assign s_dadda_cska12_fa43_or0 = s_dadda_cska12_fa43_and0 | s_dadda_cska12_fa43_and1;
  assign s_dadda_cska12_fa44_xor0 = s_dadda_cska12_fa43_or0 ^ s_dadda_cska12_fa42_or0;
  assign s_dadda_cska12_fa44_and0 = s_dadda_cska12_fa43_or0 & s_dadda_cska12_fa42_or0;
  assign s_dadda_cska12_fa44_xor1 = s_dadda_cska12_fa44_xor0 ^ s_dadda_cska12_fa41_or0;
  assign s_dadda_cska12_fa44_and1 = s_dadda_cska12_fa44_xor0 & s_dadda_cska12_fa41_or0;
  assign s_dadda_cska12_fa44_or0 = s_dadda_cska12_fa44_and0 | s_dadda_cska12_fa44_and1;
  assign s_dadda_cska12_and_10_4 = a[10] & b[4];
  assign s_dadda_cska12_fa45_xor0 = s_dadda_cska12_fa40_or0 ^ s_dadda_cska12_fa39_or0;
  assign s_dadda_cska12_fa45_and0 = s_dadda_cska12_fa40_or0 & s_dadda_cska12_fa39_or0;
  assign s_dadda_cska12_fa45_xor1 = s_dadda_cska12_fa45_xor0 ^ s_dadda_cska12_and_10_4;
  assign s_dadda_cska12_fa45_and1 = s_dadda_cska12_fa45_xor0 & s_dadda_cska12_and_10_4;
  assign s_dadda_cska12_fa45_or0 = s_dadda_cska12_fa45_and0 | s_dadda_cska12_fa45_and1;
  assign s_dadda_cska12_and_9_5 = a[9] & b[5];
  assign s_dadda_cska12_and_8_6 = a[8] & b[6];
  assign s_dadda_cska12_and_7_7 = a[7] & b[7];
  assign s_dadda_cska12_fa46_xor0 = s_dadda_cska12_and_9_5 ^ s_dadda_cska12_and_8_6;
  assign s_dadda_cska12_fa46_and0 = s_dadda_cska12_and_9_5 & s_dadda_cska12_and_8_6;
  assign s_dadda_cska12_fa46_xor1 = s_dadda_cska12_fa46_xor0 ^ s_dadda_cska12_and_7_7;
  assign s_dadda_cska12_fa46_and1 = s_dadda_cska12_fa46_xor0 & s_dadda_cska12_and_7_7;
  assign s_dadda_cska12_fa46_or0 = s_dadda_cska12_fa46_and0 | s_dadda_cska12_fa46_and1;
  assign s_dadda_cska12_and_6_8 = a[6] & b[8];
  assign s_dadda_cska12_and_5_9 = a[5] & b[9];
  assign s_dadda_cska12_and_4_10 = a[4] & b[10];
  assign s_dadda_cska12_fa47_xor0 = s_dadda_cska12_and_6_8 ^ s_dadda_cska12_and_5_9;
  assign s_dadda_cska12_fa47_and0 = s_dadda_cska12_and_6_8 & s_dadda_cska12_and_5_9;
  assign s_dadda_cska12_fa47_xor1 = s_dadda_cska12_fa47_xor0 ^ s_dadda_cska12_and_4_10;
  assign s_dadda_cska12_fa47_and1 = s_dadda_cska12_fa47_xor0 & s_dadda_cska12_and_4_10;
  assign s_dadda_cska12_fa47_or0 = s_dadda_cska12_fa47_and0 | s_dadda_cska12_fa47_and1;
  assign s_dadda_cska12_nand_3_11 = ~(a[3] & b[11]);
  assign s_dadda_cska12_fa48_xor0 = s_dadda_cska12_nand_3_11 ^ s_dadda_cska12_fa8_xor1;
  assign s_dadda_cska12_fa48_and0 = s_dadda_cska12_nand_3_11 & s_dadda_cska12_fa8_xor1;
  assign s_dadda_cska12_fa48_xor1 = s_dadda_cska12_fa48_xor0 ^ s_dadda_cska12_fa44_xor1;
  assign s_dadda_cska12_fa48_and1 = s_dadda_cska12_fa48_xor0 & s_dadda_cska12_fa44_xor1;
  assign s_dadda_cska12_fa48_or0 = s_dadda_cska12_fa48_and0 | s_dadda_cska12_fa48_and1;
  assign s_dadda_cska12_fa49_xor0 = s_dadda_cska12_fa48_or0 ^ s_dadda_cska12_fa47_or0;
  assign s_dadda_cska12_fa49_and0 = s_dadda_cska12_fa48_or0 & s_dadda_cska12_fa47_or0;
  assign s_dadda_cska12_fa49_xor1 = s_dadda_cska12_fa49_xor0 ^ s_dadda_cska12_fa46_or0;
  assign s_dadda_cska12_fa49_and1 = s_dadda_cska12_fa49_xor0 & s_dadda_cska12_fa46_or0;
  assign s_dadda_cska12_fa49_or0 = s_dadda_cska12_fa49_and0 | s_dadda_cska12_fa49_and1;
  assign s_dadda_cska12_fa50_xor0 = s_dadda_cska12_fa45_or0 ^ s_dadda_cska12_fa44_or0;
  assign s_dadda_cska12_fa50_and0 = s_dadda_cska12_fa45_or0 & s_dadda_cska12_fa44_or0;
  assign s_dadda_cska12_fa50_xor1 = s_dadda_cska12_fa50_xor0 ^ s_dadda_cska12_fa8_or0;
  assign s_dadda_cska12_fa50_and1 = s_dadda_cska12_fa50_xor0 & s_dadda_cska12_fa8_or0;
  assign s_dadda_cska12_fa50_or0 = s_dadda_cska12_fa50_and0 | s_dadda_cska12_fa50_and1;
  assign s_dadda_cska12_nand_11_4 = ~(a[11] & b[4]);
  assign s_dadda_cska12_and_10_5 = a[10] & b[5];
  assign s_dadda_cska12_and_9_6 = a[9] & b[6];
  assign s_dadda_cska12_fa51_xor0 = s_dadda_cska12_nand_11_4 ^ s_dadda_cska12_and_10_5;
  assign s_dadda_cska12_fa51_and0 = s_dadda_cska12_nand_11_4 & s_dadda_cska12_and_10_5;
  assign s_dadda_cska12_fa51_xor1 = s_dadda_cska12_fa51_xor0 ^ s_dadda_cska12_and_9_6;
  assign s_dadda_cska12_fa51_and1 = s_dadda_cska12_fa51_xor0 & s_dadda_cska12_and_9_6;
  assign s_dadda_cska12_fa51_or0 = s_dadda_cska12_fa51_and0 | s_dadda_cska12_fa51_and1;
  assign s_dadda_cska12_and_8_7 = a[8] & b[7];
  assign s_dadda_cska12_and_7_8 = a[7] & b[8];
  assign s_dadda_cska12_and_6_9 = a[6] & b[9];
  assign s_dadda_cska12_fa52_xor0 = s_dadda_cska12_and_8_7 ^ s_dadda_cska12_and_7_8;
  assign s_dadda_cska12_fa52_and0 = s_dadda_cska12_and_8_7 & s_dadda_cska12_and_7_8;
  assign s_dadda_cska12_fa52_xor1 = s_dadda_cska12_fa52_xor0 ^ s_dadda_cska12_and_6_9;
  assign s_dadda_cska12_fa52_and1 = s_dadda_cska12_fa52_xor0 & s_dadda_cska12_and_6_9;
  assign s_dadda_cska12_fa52_or0 = s_dadda_cska12_fa52_and0 | s_dadda_cska12_fa52_and1;
  assign s_dadda_cska12_and_5_10 = a[5] & b[10];
  assign s_dadda_cska12_nand_4_11 = ~(a[4] & b[11]);
  assign s_dadda_cska12_fa53_xor0 = s_dadda_cska12_and_5_10 ^ s_dadda_cska12_nand_4_11;
  assign s_dadda_cska12_fa53_and0 = s_dadda_cska12_and_5_10 & s_dadda_cska12_nand_4_11;
  assign s_dadda_cska12_fa53_xor1 = s_dadda_cska12_fa53_xor0 ^ s_dadda_cska12_fa49_xor1;
  assign s_dadda_cska12_fa53_and1 = s_dadda_cska12_fa53_xor0 & s_dadda_cska12_fa49_xor1;
  assign s_dadda_cska12_fa53_or0 = s_dadda_cska12_fa53_and0 | s_dadda_cska12_fa53_and1;
  assign s_dadda_cska12_fa54_xor0 = s_dadda_cska12_fa53_or0 ^ s_dadda_cska12_fa52_or0;
  assign s_dadda_cska12_fa54_and0 = s_dadda_cska12_fa53_or0 & s_dadda_cska12_fa52_or0;
  assign s_dadda_cska12_fa54_xor1 = s_dadda_cska12_fa54_xor0 ^ s_dadda_cska12_fa51_or0;
  assign s_dadda_cska12_fa54_and1 = s_dadda_cska12_fa54_xor0 & s_dadda_cska12_fa51_or0;
  assign s_dadda_cska12_fa54_or0 = s_dadda_cska12_fa54_and0 | s_dadda_cska12_fa54_and1;
  assign s_dadda_cska12_nand_11_5 = ~(a[11] & b[5]);
  assign s_dadda_cska12_fa55_xor0 = s_dadda_cska12_fa50_or0 ^ s_dadda_cska12_fa49_or0;
  assign s_dadda_cska12_fa55_and0 = s_dadda_cska12_fa50_or0 & s_dadda_cska12_fa49_or0;
  assign s_dadda_cska12_fa55_xor1 = s_dadda_cska12_fa55_xor0 ^ s_dadda_cska12_nand_11_5;
  assign s_dadda_cska12_fa55_and1 = s_dadda_cska12_fa55_xor0 & s_dadda_cska12_nand_11_5;
  assign s_dadda_cska12_fa55_or0 = s_dadda_cska12_fa55_and0 | s_dadda_cska12_fa55_and1;
  assign s_dadda_cska12_and_10_6 = a[10] & b[6];
  assign s_dadda_cska12_and_9_7 = a[9] & b[7];
  assign s_dadda_cska12_and_8_8 = a[8] & b[8];
  assign s_dadda_cska12_fa56_xor0 = s_dadda_cska12_and_10_6 ^ s_dadda_cska12_and_9_7;
  assign s_dadda_cska12_fa56_and0 = s_dadda_cska12_and_10_6 & s_dadda_cska12_and_9_7;
  assign s_dadda_cska12_fa56_xor1 = s_dadda_cska12_fa56_xor0 ^ s_dadda_cska12_and_8_8;
  assign s_dadda_cska12_fa56_and1 = s_dadda_cska12_fa56_xor0 & s_dadda_cska12_and_8_8;
  assign s_dadda_cska12_fa56_or0 = s_dadda_cska12_fa56_and0 | s_dadda_cska12_fa56_and1;
  assign s_dadda_cska12_and_7_9 = a[7] & b[9];
  assign s_dadda_cska12_and_6_10 = a[6] & b[10];
  assign s_dadda_cska12_nand_5_11 = ~(a[5] & b[11]);
  assign s_dadda_cska12_fa57_xor0 = s_dadda_cska12_and_7_9 ^ s_dadda_cska12_and_6_10;
  assign s_dadda_cska12_fa57_and0 = s_dadda_cska12_and_7_9 & s_dadda_cska12_and_6_10;
  assign s_dadda_cska12_fa57_xor1 = s_dadda_cska12_fa57_xor0 ^ s_dadda_cska12_nand_5_11;
  assign s_dadda_cska12_fa57_and1 = s_dadda_cska12_fa57_xor0 & s_dadda_cska12_nand_5_11;
  assign s_dadda_cska12_fa57_or0 = s_dadda_cska12_fa57_and0 | s_dadda_cska12_fa57_and1;
  assign s_dadda_cska12_fa58_xor0 = s_dadda_cska12_fa57_or0 ^ s_dadda_cska12_fa56_or0;
  assign s_dadda_cska12_fa58_and0 = s_dadda_cska12_fa57_or0 & s_dadda_cska12_fa56_or0;
  assign s_dadda_cska12_fa58_xor1 = s_dadda_cska12_fa58_xor0 ^ s_dadda_cska12_fa55_or0;
  assign s_dadda_cska12_fa58_and1 = s_dadda_cska12_fa58_xor0 & s_dadda_cska12_fa55_or0;
  assign s_dadda_cska12_fa58_or0 = s_dadda_cska12_fa58_and0 | s_dadda_cska12_fa58_and1;
  assign s_dadda_cska12_nand_11_6 = ~(a[11] & b[6]);
  assign s_dadda_cska12_and_10_7 = a[10] & b[7];
  assign s_dadda_cska12_fa59_xor0 = s_dadda_cska12_fa54_or0 ^ s_dadda_cska12_nand_11_6;
  assign s_dadda_cska12_fa59_and0 = s_dadda_cska12_fa54_or0 & s_dadda_cska12_nand_11_6;
  assign s_dadda_cska12_fa59_xor1 = s_dadda_cska12_fa59_xor0 ^ s_dadda_cska12_and_10_7;
  assign s_dadda_cska12_fa59_and1 = s_dadda_cska12_fa59_xor0 & s_dadda_cska12_and_10_7;
  assign s_dadda_cska12_fa59_or0 = s_dadda_cska12_fa59_and0 | s_dadda_cska12_fa59_and1;
  assign s_dadda_cska12_and_9_8 = a[9] & b[8];
  assign s_dadda_cska12_and_8_9 = a[8] & b[9];
  assign s_dadda_cska12_and_7_10 = a[7] & b[10];
  assign s_dadda_cska12_fa60_xor0 = s_dadda_cska12_and_9_8 ^ s_dadda_cska12_and_8_9;
  assign s_dadda_cska12_fa60_and0 = s_dadda_cska12_and_9_8 & s_dadda_cska12_and_8_9;
  assign s_dadda_cska12_fa60_xor1 = s_dadda_cska12_fa60_xor0 ^ s_dadda_cska12_and_7_10;
  assign s_dadda_cska12_fa60_and1 = s_dadda_cska12_fa60_xor0 & s_dadda_cska12_and_7_10;
  assign s_dadda_cska12_fa60_or0 = s_dadda_cska12_fa60_and0 | s_dadda_cska12_fa60_and1;
  assign s_dadda_cska12_fa61_xor0 = s_dadda_cska12_fa60_or0 ^ s_dadda_cska12_fa59_or0;
  assign s_dadda_cska12_fa61_and0 = s_dadda_cska12_fa60_or0 & s_dadda_cska12_fa59_or0;
  assign s_dadda_cska12_fa61_xor1 = s_dadda_cska12_fa61_xor0 ^ s_dadda_cska12_fa58_or0;
  assign s_dadda_cska12_fa61_and1 = s_dadda_cska12_fa61_xor0 & s_dadda_cska12_fa58_or0;
  assign s_dadda_cska12_fa61_or0 = s_dadda_cska12_fa61_and0 | s_dadda_cska12_fa61_and1;
  assign s_dadda_cska12_nand_11_7 = ~(a[11] & b[7]);
  assign s_dadda_cska12_and_10_8 = a[10] & b[8];
  assign s_dadda_cska12_and_9_9 = a[9] & b[9];
  assign s_dadda_cska12_fa62_xor0 = s_dadda_cska12_nand_11_7 ^ s_dadda_cska12_and_10_8;
  assign s_dadda_cska12_fa62_and0 = s_dadda_cska12_nand_11_7 & s_dadda_cska12_and_10_8;
  assign s_dadda_cska12_fa62_xor1 = s_dadda_cska12_fa62_xor0 ^ s_dadda_cska12_and_9_9;
  assign s_dadda_cska12_fa62_and1 = s_dadda_cska12_fa62_xor0 & s_dadda_cska12_and_9_9;
  assign s_dadda_cska12_fa62_or0 = s_dadda_cska12_fa62_and0 | s_dadda_cska12_fa62_and1;
  assign s_dadda_cska12_nand_11_8 = ~(a[11] & b[8]);
  assign s_dadda_cska12_fa63_xor0 = s_dadda_cska12_fa62_or0 ^ s_dadda_cska12_fa61_or0;
  assign s_dadda_cska12_fa63_and0 = s_dadda_cska12_fa62_or0 & s_dadda_cska12_fa61_or0;
  assign s_dadda_cska12_fa63_xor1 = s_dadda_cska12_fa63_xor0 ^ s_dadda_cska12_nand_11_8;
  assign s_dadda_cska12_fa63_and1 = s_dadda_cska12_fa63_xor0 & s_dadda_cska12_nand_11_8;
  assign s_dadda_cska12_fa63_or0 = s_dadda_cska12_fa63_and0 | s_dadda_cska12_fa63_and1;
  assign s_dadda_cska12_and_3_0 = a[3] & b[0];
  assign s_dadda_cska12_and_2_1 = a[2] & b[1];
  assign s_dadda_cska12_ha8_xor0 = s_dadda_cska12_and_3_0 ^ s_dadda_cska12_and_2_1;
  assign s_dadda_cska12_ha8_and0 = s_dadda_cska12_and_3_0 & s_dadda_cska12_and_2_1;
  assign s_dadda_cska12_and_2_2 = a[2] & b[2];
  assign s_dadda_cska12_and_1_3 = a[1] & b[3];
  assign s_dadda_cska12_fa64_xor0 = s_dadda_cska12_ha8_and0 ^ s_dadda_cska12_and_2_2;
  assign s_dadda_cska12_fa64_and0 = s_dadda_cska12_ha8_and0 & s_dadda_cska12_and_2_2;
  assign s_dadda_cska12_fa64_xor1 = s_dadda_cska12_fa64_xor0 ^ s_dadda_cska12_and_1_3;
  assign s_dadda_cska12_fa64_and1 = s_dadda_cska12_fa64_xor0 & s_dadda_cska12_and_1_3;
  assign s_dadda_cska12_fa64_or0 = s_dadda_cska12_fa64_and0 | s_dadda_cska12_fa64_and1;
  assign s_dadda_cska12_and_1_4 = a[1] & b[4];
  assign s_dadda_cska12_and_0_5 = a[0] & b[5];
  assign s_dadda_cska12_fa65_xor0 = s_dadda_cska12_fa64_or0 ^ s_dadda_cska12_and_1_4;
  assign s_dadda_cska12_fa65_and0 = s_dadda_cska12_fa64_or0 & s_dadda_cska12_and_1_4;
  assign s_dadda_cska12_fa65_xor1 = s_dadda_cska12_fa65_xor0 ^ s_dadda_cska12_and_0_5;
  assign s_dadda_cska12_fa65_and1 = s_dadda_cska12_fa65_xor0 & s_dadda_cska12_and_0_5;
  assign s_dadda_cska12_fa65_or0 = s_dadda_cska12_fa65_and0 | s_dadda_cska12_fa65_and1;
  assign s_dadda_cska12_and_0_6 = a[0] & b[6];
  assign s_dadda_cska12_fa66_xor0 = s_dadda_cska12_fa65_or0 ^ s_dadda_cska12_and_0_6;
  assign s_dadda_cska12_fa66_and0 = s_dadda_cska12_fa65_or0 & s_dadda_cska12_and_0_6;
  assign s_dadda_cska12_fa66_xor1 = s_dadda_cska12_fa66_xor0 ^ s_dadda_cska12_fa10_xor1;
  assign s_dadda_cska12_fa66_and1 = s_dadda_cska12_fa66_xor0 & s_dadda_cska12_fa10_xor1;
  assign s_dadda_cska12_fa66_or0 = s_dadda_cska12_fa66_and0 | s_dadda_cska12_fa66_and1;
  assign s_dadda_cska12_fa67_xor0 = s_dadda_cska12_fa66_or0 ^ s_dadda_cska12_fa12_xor1;
  assign s_dadda_cska12_fa67_and0 = s_dadda_cska12_fa66_or0 & s_dadda_cska12_fa12_xor1;
  assign s_dadda_cska12_fa67_xor1 = s_dadda_cska12_fa67_xor0 ^ s_dadda_cska12_fa13_xor1;
  assign s_dadda_cska12_fa67_and1 = s_dadda_cska12_fa67_xor0 & s_dadda_cska12_fa13_xor1;
  assign s_dadda_cska12_fa67_or0 = s_dadda_cska12_fa67_and0 | s_dadda_cska12_fa67_and1;
  assign s_dadda_cska12_fa68_xor0 = s_dadda_cska12_fa67_or0 ^ s_dadda_cska12_fa16_xor1;
  assign s_dadda_cska12_fa68_and0 = s_dadda_cska12_fa67_or0 & s_dadda_cska12_fa16_xor1;
  assign s_dadda_cska12_fa68_xor1 = s_dadda_cska12_fa68_xor0 ^ s_dadda_cska12_fa17_xor1;
  assign s_dadda_cska12_fa68_and1 = s_dadda_cska12_fa68_xor0 & s_dadda_cska12_fa17_xor1;
  assign s_dadda_cska12_fa68_or0 = s_dadda_cska12_fa68_and0 | s_dadda_cska12_fa68_and1;
  assign s_dadda_cska12_fa69_xor0 = s_dadda_cska12_fa68_or0 ^ s_dadda_cska12_fa20_xor1;
  assign s_dadda_cska12_fa69_and0 = s_dadda_cska12_fa68_or0 & s_dadda_cska12_fa20_xor1;
  assign s_dadda_cska12_fa69_xor1 = s_dadda_cska12_fa69_xor0 ^ s_dadda_cska12_fa21_xor1;
  assign s_dadda_cska12_fa69_and1 = s_dadda_cska12_fa69_xor0 & s_dadda_cska12_fa21_xor1;
  assign s_dadda_cska12_fa69_or0 = s_dadda_cska12_fa69_and0 | s_dadda_cska12_fa69_and1;
  assign s_dadda_cska12_fa70_xor0 = s_dadda_cska12_fa69_or0 ^ s_dadda_cska12_fa25_xor1;
  assign s_dadda_cska12_fa70_and0 = s_dadda_cska12_fa69_or0 & s_dadda_cska12_fa25_xor1;
  assign s_dadda_cska12_fa70_xor1 = s_dadda_cska12_fa70_xor0 ^ s_dadda_cska12_fa26_xor1;
  assign s_dadda_cska12_fa70_and1 = s_dadda_cska12_fa70_xor0 & s_dadda_cska12_fa26_xor1;
  assign s_dadda_cska12_fa70_or0 = s_dadda_cska12_fa70_and0 | s_dadda_cska12_fa70_and1;
  assign s_dadda_cska12_fa71_xor0 = s_dadda_cska12_fa70_or0 ^ s_dadda_cska12_fa30_xor1;
  assign s_dadda_cska12_fa71_and0 = s_dadda_cska12_fa70_or0 & s_dadda_cska12_fa30_xor1;
  assign s_dadda_cska12_fa71_xor1 = s_dadda_cska12_fa71_xor0 ^ s_dadda_cska12_fa31_xor1;
  assign s_dadda_cska12_fa71_and1 = s_dadda_cska12_fa71_xor0 & s_dadda_cska12_fa31_xor1;
  assign s_dadda_cska12_fa71_or0 = s_dadda_cska12_fa71_and0 | s_dadda_cska12_fa71_and1;
  assign s_dadda_cska12_fa72_xor0 = s_dadda_cska12_fa71_or0 ^ s_dadda_cska12_fa35_xor1;
  assign s_dadda_cska12_fa72_and0 = s_dadda_cska12_fa71_or0 & s_dadda_cska12_fa35_xor1;
  assign s_dadda_cska12_fa72_xor1 = s_dadda_cska12_fa72_xor0 ^ s_dadda_cska12_fa36_xor1;
  assign s_dadda_cska12_fa72_and1 = s_dadda_cska12_fa72_xor0 & s_dadda_cska12_fa36_xor1;
  assign s_dadda_cska12_fa72_or0 = s_dadda_cska12_fa72_and0 | s_dadda_cska12_fa72_and1;
  assign s_dadda_cska12_fa73_xor0 = s_dadda_cska12_fa72_or0 ^ s_dadda_cska12_fa40_xor1;
  assign s_dadda_cska12_fa73_and0 = s_dadda_cska12_fa72_or0 & s_dadda_cska12_fa40_xor1;
  assign s_dadda_cska12_fa73_xor1 = s_dadda_cska12_fa73_xor0 ^ s_dadda_cska12_fa41_xor1;
  assign s_dadda_cska12_fa73_and1 = s_dadda_cska12_fa73_xor0 & s_dadda_cska12_fa41_xor1;
  assign s_dadda_cska12_fa73_or0 = s_dadda_cska12_fa73_and0 | s_dadda_cska12_fa73_and1;
  assign s_dadda_cska12_fa74_xor0 = s_dadda_cska12_fa73_or0 ^ s_dadda_cska12_fa45_xor1;
  assign s_dadda_cska12_fa74_and0 = s_dadda_cska12_fa73_or0 & s_dadda_cska12_fa45_xor1;
  assign s_dadda_cska12_fa74_xor1 = s_dadda_cska12_fa74_xor0 ^ s_dadda_cska12_fa46_xor1;
  assign s_dadda_cska12_fa74_and1 = s_dadda_cska12_fa74_xor0 & s_dadda_cska12_fa46_xor1;
  assign s_dadda_cska12_fa74_or0 = s_dadda_cska12_fa74_and0 | s_dadda_cska12_fa74_and1;
  assign s_dadda_cska12_fa75_xor0 = s_dadda_cska12_fa74_or0 ^ s_dadda_cska12_fa50_xor1;
  assign s_dadda_cska12_fa75_and0 = s_dadda_cska12_fa74_or0 & s_dadda_cska12_fa50_xor1;
  assign s_dadda_cska12_fa75_xor1 = s_dadda_cska12_fa75_xor0 ^ s_dadda_cska12_fa51_xor1;
  assign s_dadda_cska12_fa75_and1 = s_dadda_cska12_fa75_xor0 & s_dadda_cska12_fa51_xor1;
  assign s_dadda_cska12_fa75_or0 = s_dadda_cska12_fa75_and0 | s_dadda_cska12_fa75_and1;
  assign s_dadda_cska12_fa76_xor0 = s_dadda_cska12_fa75_or0 ^ s_dadda_cska12_fa54_xor1;
  assign s_dadda_cska12_fa76_and0 = s_dadda_cska12_fa75_or0 & s_dadda_cska12_fa54_xor1;
  assign s_dadda_cska12_fa76_xor1 = s_dadda_cska12_fa76_xor0 ^ s_dadda_cska12_fa55_xor1;
  assign s_dadda_cska12_fa76_and1 = s_dadda_cska12_fa76_xor0 & s_dadda_cska12_fa55_xor1;
  assign s_dadda_cska12_fa76_or0 = s_dadda_cska12_fa76_and0 | s_dadda_cska12_fa76_and1;
  assign s_dadda_cska12_nand_6_11 = ~(a[6] & b[11]);
  assign s_dadda_cska12_fa77_xor0 = s_dadda_cska12_fa76_or0 ^ s_dadda_cska12_nand_6_11;
  assign s_dadda_cska12_fa77_and0 = s_dadda_cska12_fa76_or0 & s_dadda_cska12_nand_6_11;
  assign s_dadda_cska12_fa77_xor1 = s_dadda_cska12_fa77_xor0 ^ s_dadda_cska12_fa58_xor1;
  assign s_dadda_cska12_fa77_and1 = s_dadda_cska12_fa77_xor0 & s_dadda_cska12_fa58_xor1;
  assign s_dadda_cska12_fa77_or0 = s_dadda_cska12_fa77_and0 | s_dadda_cska12_fa77_and1;
  assign s_dadda_cska12_and_8_10 = a[8] & b[10];
  assign s_dadda_cska12_nand_7_11 = ~(a[7] & b[11]);
  assign s_dadda_cska12_fa78_xor0 = s_dadda_cska12_fa77_or0 ^ s_dadda_cska12_and_8_10;
  assign s_dadda_cska12_fa78_and0 = s_dadda_cska12_fa77_or0 & s_dadda_cska12_and_8_10;
  assign s_dadda_cska12_fa78_xor1 = s_dadda_cska12_fa78_xor0 ^ s_dadda_cska12_nand_7_11;
  assign s_dadda_cska12_fa78_and1 = s_dadda_cska12_fa78_xor0 & s_dadda_cska12_nand_7_11;
  assign s_dadda_cska12_fa78_or0 = s_dadda_cska12_fa78_and0 | s_dadda_cska12_fa78_and1;
  assign s_dadda_cska12_and_10_9 = a[10] & b[9];
  assign s_dadda_cska12_and_9_10 = a[9] & b[10];
  assign s_dadda_cska12_fa79_xor0 = s_dadda_cska12_fa78_or0 ^ s_dadda_cska12_and_10_9;
  assign s_dadda_cska12_fa79_and0 = s_dadda_cska12_fa78_or0 & s_dadda_cska12_and_10_9;
  assign s_dadda_cska12_fa79_xor1 = s_dadda_cska12_fa79_xor0 ^ s_dadda_cska12_and_9_10;
  assign s_dadda_cska12_fa79_and1 = s_dadda_cska12_fa79_xor0 & s_dadda_cska12_and_9_10;
  assign s_dadda_cska12_fa79_or0 = s_dadda_cska12_fa79_and0 | s_dadda_cska12_fa79_and1;
  assign s_dadda_cska12_nand_11_9 = ~(a[11] & b[9]);
  assign s_dadda_cska12_fa80_xor0 = s_dadda_cska12_fa79_or0 ^ s_dadda_cska12_fa63_or0;
  assign s_dadda_cska12_fa80_and0 = s_dadda_cska12_fa79_or0 & s_dadda_cska12_fa63_or0;
  assign s_dadda_cska12_fa80_xor1 = s_dadda_cska12_fa80_xor0 ^ s_dadda_cska12_nand_11_9;
  assign s_dadda_cska12_fa80_and1 = s_dadda_cska12_fa80_xor0 & s_dadda_cska12_nand_11_9;
  assign s_dadda_cska12_fa80_or0 = s_dadda_cska12_fa80_and0 | s_dadda_cska12_fa80_and1;
  assign s_dadda_cska12_and_2_0 = a[2] & b[0];
  assign s_dadda_cska12_and_1_1 = a[1] & b[1];
  assign s_dadda_cska12_ha9_xor0 = s_dadda_cska12_and_2_0 ^ s_dadda_cska12_and_1_1;
  assign s_dadda_cska12_ha9_and0 = s_dadda_cska12_and_2_0 & s_dadda_cska12_and_1_1;
  assign s_dadda_cska12_and_1_2 = a[1] & b[2];
  assign s_dadda_cska12_and_0_3 = a[0] & b[3];
  assign s_dadda_cska12_fa81_xor0 = s_dadda_cska12_ha9_and0 ^ s_dadda_cska12_and_1_2;
  assign s_dadda_cska12_fa81_and0 = s_dadda_cska12_ha9_and0 & s_dadda_cska12_and_1_2;
  assign s_dadda_cska12_fa81_xor1 = s_dadda_cska12_fa81_xor0 ^ s_dadda_cska12_and_0_3;
  assign s_dadda_cska12_fa81_and1 = s_dadda_cska12_fa81_xor0 & s_dadda_cska12_and_0_3;
  assign s_dadda_cska12_fa81_or0 = s_dadda_cska12_fa81_and0 | s_dadda_cska12_fa81_and1;
  assign s_dadda_cska12_and_0_4 = a[0] & b[4];
  assign s_dadda_cska12_fa82_xor0 = s_dadda_cska12_fa81_or0 ^ s_dadda_cska12_and_0_4;
  assign s_dadda_cska12_fa82_and0 = s_dadda_cska12_fa81_or0 & s_dadda_cska12_and_0_4;
  assign s_dadda_cska12_fa82_xor1 = s_dadda_cska12_fa82_xor0 ^ s_dadda_cska12_ha3_xor0;
  assign s_dadda_cska12_fa82_and1 = s_dadda_cska12_fa82_xor0 & s_dadda_cska12_ha3_xor0;
  assign s_dadda_cska12_fa82_or0 = s_dadda_cska12_fa82_and0 | s_dadda_cska12_fa82_and1;
  assign s_dadda_cska12_fa83_xor0 = s_dadda_cska12_fa82_or0 ^ s_dadda_cska12_fa9_xor1;
  assign s_dadda_cska12_fa83_and0 = s_dadda_cska12_fa82_or0 & s_dadda_cska12_fa9_xor1;
  assign s_dadda_cska12_fa83_xor1 = s_dadda_cska12_fa83_xor0 ^ s_dadda_cska12_ha4_xor0;
  assign s_dadda_cska12_fa83_and1 = s_dadda_cska12_fa83_xor0 & s_dadda_cska12_ha4_xor0;
  assign s_dadda_cska12_fa83_or0 = s_dadda_cska12_fa83_and0 | s_dadda_cska12_fa83_and1;
  assign s_dadda_cska12_fa84_xor0 = s_dadda_cska12_fa83_or0 ^ s_dadda_cska12_fa11_xor1;
  assign s_dadda_cska12_fa84_and0 = s_dadda_cska12_fa83_or0 & s_dadda_cska12_fa11_xor1;
  assign s_dadda_cska12_fa84_xor1 = s_dadda_cska12_fa84_xor0 ^ s_dadda_cska12_ha5_xor0;
  assign s_dadda_cska12_fa84_and1 = s_dadda_cska12_fa84_xor0 & s_dadda_cska12_ha5_xor0;
  assign s_dadda_cska12_fa84_or0 = s_dadda_cska12_fa84_and0 | s_dadda_cska12_fa84_and1;
  assign s_dadda_cska12_fa85_xor0 = s_dadda_cska12_fa84_or0 ^ s_dadda_cska12_fa14_xor1;
  assign s_dadda_cska12_fa85_and0 = s_dadda_cska12_fa84_or0 & s_dadda_cska12_fa14_xor1;
  assign s_dadda_cska12_fa85_xor1 = s_dadda_cska12_fa85_xor0 ^ s_dadda_cska12_ha6_xor0;
  assign s_dadda_cska12_fa85_and1 = s_dadda_cska12_fa85_xor0 & s_dadda_cska12_ha6_xor0;
  assign s_dadda_cska12_fa85_or0 = s_dadda_cska12_fa85_and0 | s_dadda_cska12_fa85_and1;
  assign s_dadda_cska12_fa86_xor0 = s_dadda_cska12_fa85_or0 ^ s_dadda_cska12_fa18_xor1;
  assign s_dadda_cska12_fa86_and0 = s_dadda_cska12_fa85_or0 & s_dadda_cska12_fa18_xor1;
  assign s_dadda_cska12_fa86_xor1 = s_dadda_cska12_fa86_xor0 ^ s_dadda_cska12_ha7_xor0;
  assign s_dadda_cska12_fa86_and1 = s_dadda_cska12_fa86_xor0 & s_dadda_cska12_ha7_xor0;
  assign s_dadda_cska12_fa86_or0 = s_dadda_cska12_fa86_and0 | s_dadda_cska12_fa86_and1;
  assign s_dadda_cska12_fa87_xor0 = s_dadda_cska12_fa86_or0 ^ s_dadda_cska12_fa22_xor1;
  assign s_dadda_cska12_fa87_and0 = s_dadda_cska12_fa86_or0 & s_dadda_cska12_fa22_xor1;
  assign s_dadda_cska12_fa87_xor1 = s_dadda_cska12_fa87_xor0 ^ s_dadda_cska12_fa23_xor1;
  assign s_dadda_cska12_fa87_and1 = s_dadda_cska12_fa87_xor0 & s_dadda_cska12_fa23_xor1;
  assign s_dadda_cska12_fa87_or0 = s_dadda_cska12_fa87_and0 | s_dadda_cska12_fa87_and1;
  assign s_dadda_cska12_fa88_xor0 = s_dadda_cska12_fa87_or0 ^ s_dadda_cska12_fa27_xor1;
  assign s_dadda_cska12_fa88_and0 = s_dadda_cska12_fa87_or0 & s_dadda_cska12_fa27_xor1;
  assign s_dadda_cska12_fa88_xor1 = s_dadda_cska12_fa88_xor0 ^ s_dadda_cska12_fa28_xor1;
  assign s_dadda_cska12_fa88_and1 = s_dadda_cska12_fa88_xor0 & s_dadda_cska12_fa28_xor1;
  assign s_dadda_cska12_fa88_or0 = s_dadda_cska12_fa88_and0 | s_dadda_cska12_fa88_and1;
  assign s_dadda_cska12_fa89_xor0 = s_dadda_cska12_fa88_or0 ^ s_dadda_cska12_fa32_xor1;
  assign s_dadda_cska12_fa89_and0 = s_dadda_cska12_fa88_or0 & s_dadda_cska12_fa32_xor1;
  assign s_dadda_cska12_fa89_xor1 = s_dadda_cska12_fa89_xor0 ^ s_dadda_cska12_fa33_xor1;
  assign s_dadda_cska12_fa89_and1 = s_dadda_cska12_fa89_xor0 & s_dadda_cska12_fa33_xor1;
  assign s_dadda_cska12_fa89_or0 = s_dadda_cska12_fa89_and0 | s_dadda_cska12_fa89_and1;
  assign s_dadda_cska12_fa90_xor0 = s_dadda_cska12_fa89_or0 ^ s_dadda_cska12_fa37_xor1;
  assign s_dadda_cska12_fa90_and0 = s_dadda_cska12_fa89_or0 & s_dadda_cska12_fa37_xor1;
  assign s_dadda_cska12_fa90_xor1 = s_dadda_cska12_fa90_xor0 ^ s_dadda_cska12_fa38_xor1;
  assign s_dadda_cska12_fa90_and1 = s_dadda_cska12_fa90_xor0 & s_dadda_cska12_fa38_xor1;
  assign s_dadda_cska12_fa90_or0 = s_dadda_cska12_fa90_and0 | s_dadda_cska12_fa90_and1;
  assign s_dadda_cska12_fa91_xor0 = s_dadda_cska12_fa90_or0 ^ s_dadda_cska12_fa42_xor1;
  assign s_dadda_cska12_fa91_and0 = s_dadda_cska12_fa90_or0 & s_dadda_cska12_fa42_xor1;
  assign s_dadda_cska12_fa91_xor1 = s_dadda_cska12_fa91_xor0 ^ s_dadda_cska12_fa43_xor1;
  assign s_dadda_cska12_fa91_and1 = s_dadda_cska12_fa91_xor0 & s_dadda_cska12_fa43_xor1;
  assign s_dadda_cska12_fa91_or0 = s_dadda_cska12_fa91_and0 | s_dadda_cska12_fa91_and1;
  assign s_dadda_cska12_fa92_xor0 = s_dadda_cska12_fa91_or0 ^ s_dadda_cska12_fa47_xor1;
  assign s_dadda_cska12_fa92_and0 = s_dadda_cska12_fa91_or0 & s_dadda_cska12_fa47_xor1;
  assign s_dadda_cska12_fa92_xor1 = s_dadda_cska12_fa92_xor0 ^ s_dadda_cska12_fa48_xor1;
  assign s_dadda_cska12_fa92_and1 = s_dadda_cska12_fa92_xor0 & s_dadda_cska12_fa48_xor1;
  assign s_dadda_cska12_fa92_or0 = s_dadda_cska12_fa92_and0 | s_dadda_cska12_fa92_and1;
  assign s_dadda_cska12_fa93_xor0 = s_dadda_cska12_fa92_or0 ^ s_dadda_cska12_fa52_xor1;
  assign s_dadda_cska12_fa93_and0 = s_dadda_cska12_fa92_or0 & s_dadda_cska12_fa52_xor1;
  assign s_dadda_cska12_fa93_xor1 = s_dadda_cska12_fa93_xor0 ^ s_dadda_cska12_fa53_xor1;
  assign s_dadda_cska12_fa93_and1 = s_dadda_cska12_fa93_xor0 & s_dadda_cska12_fa53_xor1;
  assign s_dadda_cska12_fa93_or0 = s_dadda_cska12_fa93_and0 | s_dadda_cska12_fa93_and1;
  assign s_dadda_cska12_fa94_xor0 = s_dadda_cska12_fa93_or0 ^ s_dadda_cska12_fa56_xor1;
  assign s_dadda_cska12_fa94_and0 = s_dadda_cska12_fa93_or0 & s_dadda_cska12_fa56_xor1;
  assign s_dadda_cska12_fa94_xor1 = s_dadda_cska12_fa94_xor0 ^ s_dadda_cska12_fa57_xor1;
  assign s_dadda_cska12_fa94_and1 = s_dadda_cska12_fa94_xor0 & s_dadda_cska12_fa57_xor1;
  assign s_dadda_cska12_fa94_or0 = s_dadda_cska12_fa94_and0 | s_dadda_cska12_fa94_and1;
  assign s_dadda_cska12_fa95_xor0 = s_dadda_cska12_fa94_or0 ^ s_dadda_cska12_fa59_xor1;
  assign s_dadda_cska12_fa95_and0 = s_dadda_cska12_fa94_or0 & s_dadda_cska12_fa59_xor1;
  assign s_dadda_cska12_fa95_xor1 = s_dadda_cska12_fa95_xor0 ^ s_dadda_cska12_fa60_xor1;
  assign s_dadda_cska12_fa95_and1 = s_dadda_cska12_fa95_xor0 & s_dadda_cska12_fa60_xor1;
  assign s_dadda_cska12_fa95_or0 = s_dadda_cska12_fa95_and0 | s_dadda_cska12_fa95_and1;
  assign s_dadda_cska12_fa96_xor0 = s_dadda_cska12_fa95_or0 ^ s_dadda_cska12_fa61_xor1;
  assign s_dadda_cska12_fa96_and0 = s_dadda_cska12_fa95_or0 & s_dadda_cska12_fa61_xor1;
  assign s_dadda_cska12_fa96_xor1 = s_dadda_cska12_fa96_xor0 ^ s_dadda_cska12_fa62_xor1;
  assign s_dadda_cska12_fa96_and1 = s_dadda_cska12_fa96_xor0 & s_dadda_cska12_fa62_xor1;
  assign s_dadda_cska12_fa96_or0 = s_dadda_cska12_fa96_and0 | s_dadda_cska12_fa96_and1;
  assign s_dadda_cska12_nand_8_11 = ~(a[8] & b[11]);
  assign s_dadda_cska12_fa97_xor0 = s_dadda_cska12_fa96_or0 ^ s_dadda_cska12_nand_8_11;
  assign s_dadda_cska12_fa97_and0 = s_dadda_cska12_fa96_or0 & s_dadda_cska12_nand_8_11;
  assign s_dadda_cska12_fa97_xor1 = s_dadda_cska12_fa97_xor0 ^ s_dadda_cska12_fa63_xor1;
  assign s_dadda_cska12_fa97_and1 = s_dadda_cska12_fa97_xor0 & s_dadda_cska12_fa63_xor1;
  assign s_dadda_cska12_fa97_or0 = s_dadda_cska12_fa97_and0 | s_dadda_cska12_fa97_and1;
  assign s_dadda_cska12_and_10_10 = a[10] & b[10];
  assign s_dadda_cska12_nand_9_11 = ~(a[9] & b[11]);
  assign s_dadda_cska12_fa98_xor0 = s_dadda_cska12_fa97_or0 ^ s_dadda_cska12_and_10_10;
  assign s_dadda_cska12_fa98_and0 = s_dadda_cska12_fa97_or0 & s_dadda_cska12_and_10_10;
  assign s_dadda_cska12_fa98_xor1 = s_dadda_cska12_fa98_xor0 ^ s_dadda_cska12_nand_9_11;
  assign s_dadda_cska12_fa98_and1 = s_dadda_cska12_fa98_xor0 & s_dadda_cska12_nand_9_11;
  assign s_dadda_cska12_fa98_or0 = s_dadda_cska12_fa98_and0 | s_dadda_cska12_fa98_and1;
  assign s_dadda_cska12_nand_11_10 = ~(a[11] & b[10]);
  assign s_dadda_cska12_fa99_xor0 = s_dadda_cska12_fa98_or0 ^ s_dadda_cska12_fa80_or0;
  assign s_dadda_cska12_fa99_and0 = s_dadda_cska12_fa98_or0 & s_dadda_cska12_fa80_or0;
  assign s_dadda_cska12_fa99_xor1 = s_dadda_cska12_fa99_xor0 ^ s_dadda_cska12_nand_11_10;
  assign s_dadda_cska12_fa99_and1 = s_dadda_cska12_fa99_xor0 & s_dadda_cska12_nand_11_10;
  assign s_dadda_cska12_fa99_or0 = s_dadda_cska12_fa99_and0 | s_dadda_cska12_fa99_and1;
  assign s_dadda_cska12_and_0_0 = a[0] & b[0];
  assign s_dadda_cska12_and_1_0 = a[1] & b[0];
  assign s_dadda_cska12_and_0_2 = a[0] & b[2];
  assign s_dadda_cska12_nand_10_11 = ~(a[10] & b[11]);
  assign s_dadda_cska12_and_0_1 = a[0] & b[1];
  assign s_dadda_cska12_and_11_11 = a[11] & b[11];
  assign s_dadda_cska12_u_cska22_xor0 = s_dadda_cska12_and_1_0 ^ s_dadda_cska12_and_0_1;
  assign s_dadda_cska12_u_cska22_ha0_xor0 = s_dadda_cska12_and_1_0 ^ s_dadda_cska12_and_0_1;
  assign s_dadda_cska12_u_cska22_ha0_and0 = s_dadda_cska12_and_1_0 & s_dadda_cska12_and_0_1;
  assign s_dadda_cska12_u_cska22_xor1 = s_dadda_cska12_and_0_2 ^ s_dadda_cska12_ha9_xor0;
  assign s_dadda_cska12_u_cska22_fa0_xor0 = s_dadda_cska12_and_0_2 ^ s_dadda_cska12_ha9_xor0;
  assign s_dadda_cska12_u_cska22_fa0_and0 = s_dadda_cska12_and_0_2 & s_dadda_cska12_ha9_xor0;
  assign s_dadda_cska12_u_cska22_fa0_xor1 = s_dadda_cska12_u_cska22_fa0_xor0 ^ s_dadda_cska12_u_cska22_ha0_and0;
  assign s_dadda_cska12_u_cska22_fa0_and1 = s_dadda_cska12_u_cska22_fa0_xor0 & s_dadda_cska12_u_cska22_ha0_and0;
  assign s_dadda_cska12_u_cska22_fa0_or0 = s_dadda_cska12_u_cska22_fa0_and0 | s_dadda_cska12_u_cska22_fa0_and1;
  assign s_dadda_cska12_u_cska22_xor2 = s_dadda_cska12_ha8_xor0 ^ s_dadda_cska12_fa81_xor1;
  assign s_dadda_cska12_u_cska22_fa1_xor0 = s_dadda_cska12_ha8_xor0 ^ s_dadda_cska12_fa81_xor1;
  assign s_dadda_cska12_u_cska22_fa1_and0 = s_dadda_cska12_ha8_xor0 & s_dadda_cska12_fa81_xor1;
  assign s_dadda_cska12_u_cska22_fa1_xor1 = s_dadda_cska12_u_cska22_fa1_xor0 ^ s_dadda_cska12_u_cska22_fa0_or0;
  assign s_dadda_cska12_u_cska22_fa1_and1 = s_dadda_cska12_u_cska22_fa1_xor0 & s_dadda_cska12_u_cska22_fa0_or0;
  assign s_dadda_cska12_u_cska22_fa1_or0 = s_dadda_cska12_u_cska22_fa1_and0 | s_dadda_cska12_u_cska22_fa1_and1;
  assign s_dadda_cska12_u_cska22_xor3 = s_dadda_cska12_fa64_xor1 ^ s_dadda_cska12_fa82_xor1;
  assign s_dadda_cska12_u_cska22_fa2_xor0 = s_dadda_cska12_fa64_xor1 ^ s_dadda_cska12_fa82_xor1;
  assign s_dadda_cska12_u_cska22_fa2_and0 = s_dadda_cska12_fa64_xor1 & s_dadda_cska12_fa82_xor1;
  assign s_dadda_cska12_u_cska22_fa2_xor1 = s_dadda_cska12_u_cska22_fa2_xor0 ^ s_dadda_cska12_u_cska22_fa1_or0;
  assign s_dadda_cska12_u_cska22_fa2_and1 = s_dadda_cska12_u_cska22_fa2_xor0 & s_dadda_cska12_u_cska22_fa1_or0;
  assign s_dadda_cska12_u_cska22_fa2_or0 = s_dadda_cska12_u_cska22_fa2_and0 | s_dadda_cska12_u_cska22_fa2_and1;
  assign s_dadda_cska12_u_cska22_and_propagate00 = s_dadda_cska12_u_cska22_xor0 & s_dadda_cska12_u_cska22_xor2;
  assign s_dadda_cska12_u_cska22_and_propagate01 = s_dadda_cska12_u_cska22_xor1 & s_dadda_cska12_u_cska22_xor3;
  assign s_dadda_cska12_u_cska22_and_propagate02 = s_dadda_cska12_u_cska22_and_propagate00 & s_dadda_cska12_u_cska22_and_propagate01;
  assign s_dadda_cska12_u_cska22_mux2to10_not0 = ~s_dadda_cska12_u_cska22_and_propagate02;
  assign s_dadda_cska12_u_cska22_mux2to10_and1 = s_dadda_cska12_u_cska22_fa2_or0 & s_dadda_cska12_u_cska22_mux2to10_not0;
  assign s_dadda_cska12_u_cska22_xor4 = s_dadda_cska12_fa65_xor1 ^ s_dadda_cska12_fa83_xor1;
  assign s_dadda_cska12_u_cska22_fa3_xor0 = s_dadda_cska12_fa65_xor1 ^ s_dadda_cska12_fa83_xor1;
  assign s_dadda_cska12_u_cska22_fa3_and0 = s_dadda_cska12_fa65_xor1 & s_dadda_cska12_fa83_xor1;
  assign s_dadda_cska12_u_cska22_fa3_xor1 = s_dadda_cska12_u_cska22_fa3_xor0 ^ s_dadda_cska12_u_cska22_mux2to10_and1;
  assign s_dadda_cska12_u_cska22_fa3_and1 = s_dadda_cska12_u_cska22_fa3_xor0 & s_dadda_cska12_u_cska22_mux2to10_and1;
  assign s_dadda_cska12_u_cska22_fa3_or0 = s_dadda_cska12_u_cska22_fa3_and0 | s_dadda_cska12_u_cska22_fa3_and1;
  assign s_dadda_cska12_u_cska22_xor5 = s_dadda_cska12_fa66_xor1 ^ s_dadda_cska12_fa84_xor1;
  assign s_dadda_cska12_u_cska22_fa4_xor0 = s_dadda_cska12_fa66_xor1 ^ s_dadda_cska12_fa84_xor1;
  assign s_dadda_cska12_u_cska22_fa4_and0 = s_dadda_cska12_fa66_xor1 & s_dadda_cska12_fa84_xor1;
  assign s_dadda_cska12_u_cska22_fa4_xor1 = s_dadda_cska12_u_cska22_fa4_xor0 ^ s_dadda_cska12_u_cska22_fa3_or0;
  assign s_dadda_cska12_u_cska22_fa4_and1 = s_dadda_cska12_u_cska22_fa4_xor0 & s_dadda_cska12_u_cska22_fa3_or0;
  assign s_dadda_cska12_u_cska22_fa4_or0 = s_dadda_cska12_u_cska22_fa4_and0 | s_dadda_cska12_u_cska22_fa4_and1;
  assign s_dadda_cska12_u_cska22_xor6 = s_dadda_cska12_fa67_xor1 ^ s_dadda_cska12_fa85_xor1;
  assign s_dadda_cska12_u_cska22_fa5_xor0 = s_dadda_cska12_fa67_xor1 ^ s_dadda_cska12_fa85_xor1;
  assign s_dadda_cska12_u_cska22_fa5_and0 = s_dadda_cska12_fa67_xor1 & s_dadda_cska12_fa85_xor1;
  assign s_dadda_cska12_u_cska22_fa5_xor1 = s_dadda_cska12_u_cska22_fa5_xor0 ^ s_dadda_cska12_u_cska22_fa4_or0;
  assign s_dadda_cska12_u_cska22_fa5_and1 = s_dadda_cska12_u_cska22_fa5_xor0 & s_dadda_cska12_u_cska22_fa4_or0;
  assign s_dadda_cska12_u_cska22_fa5_or0 = s_dadda_cska12_u_cska22_fa5_and0 | s_dadda_cska12_u_cska22_fa5_and1;
  assign s_dadda_cska12_u_cska22_xor7 = s_dadda_cska12_fa68_xor1 ^ s_dadda_cska12_fa86_xor1;
  assign s_dadda_cska12_u_cska22_fa6_xor0 = s_dadda_cska12_fa68_xor1 ^ s_dadda_cska12_fa86_xor1;
  assign s_dadda_cska12_u_cska22_fa6_and0 = s_dadda_cska12_fa68_xor1 & s_dadda_cska12_fa86_xor1;
  assign s_dadda_cska12_u_cska22_fa6_xor1 = s_dadda_cska12_u_cska22_fa6_xor0 ^ s_dadda_cska12_u_cska22_fa5_or0;
  assign s_dadda_cska12_u_cska22_fa6_and1 = s_dadda_cska12_u_cska22_fa6_xor0 & s_dadda_cska12_u_cska22_fa5_or0;
  assign s_dadda_cska12_u_cska22_fa6_or0 = s_dadda_cska12_u_cska22_fa6_and0 | s_dadda_cska12_u_cska22_fa6_and1;
  assign s_dadda_cska12_u_cska22_and_propagate13 = s_dadda_cska12_u_cska22_xor4 & s_dadda_cska12_u_cska22_xor6;
  assign s_dadda_cska12_u_cska22_and_propagate14 = s_dadda_cska12_u_cska22_xor5 & s_dadda_cska12_u_cska22_xor7;
  assign s_dadda_cska12_u_cska22_and_propagate15 = s_dadda_cska12_u_cska22_and_propagate13 & s_dadda_cska12_u_cska22_and_propagate14;
  assign s_dadda_cska12_u_cska22_mux2to11_and0 = s_dadda_cska12_u_cska22_mux2to10_and1 & s_dadda_cska12_u_cska22_and_propagate15;
  assign s_dadda_cska12_u_cska22_mux2to11_not0 = ~s_dadda_cska12_u_cska22_and_propagate15;
  assign s_dadda_cska12_u_cska22_mux2to11_and1 = s_dadda_cska12_u_cska22_fa6_or0 & s_dadda_cska12_u_cska22_mux2to11_not0;
  assign s_dadda_cska12_u_cska22_mux2to11_xor0 = s_dadda_cska12_u_cska22_mux2to11_and0 ^ s_dadda_cska12_u_cska22_mux2to11_and1;
  assign s_dadda_cska12_u_cska22_xor8 = s_dadda_cska12_fa69_xor1 ^ s_dadda_cska12_fa87_xor1;
  assign s_dadda_cska12_u_cska22_fa7_xor0 = s_dadda_cska12_fa69_xor1 ^ s_dadda_cska12_fa87_xor1;
  assign s_dadda_cska12_u_cska22_fa7_and0 = s_dadda_cska12_fa69_xor1 & s_dadda_cska12_fa87_xor1;
  assign s_dadda_cska12_u_cska22_fa7_xor1 = s_dadda_cska12_u_cska22_fa7_xor0 ^ s_dadda_cska12_u_cska22_mux2to11_xor0;
  assign s_dadda_cska12_u_cska22_fa7_and1 = s_dadda_cska12_u_cska22_fa7_xor0 & s_dadda_cska12_u_cska22_mux2to11_xor0;
  assign s_dadda_cska12_u_cska22_fa7_or0 = s_dadda_cska12_u_cska22_fa7_and0 | s_dadda_cska12_u_cska22_fa7_and1;
  assign s_dadda_cska12_u_cska22_xor9 = s_dadda_cska12_fa70_xor1 ^ s_dadda_cska12_fa88_xor1;
  assign s_dadda_cska12_u_cska22_fa8_xor0 = s_dadda_cska12_fa70_xor1 ^ s_dadda_cska12_fa88_xor1;
  assign s_dadda_cska12_u_cska22_fa8_and0 = s_dadda_cska12_fa70_xor1 & s_dadda_cska12_fa88_xor1;
  assign s_dadda_cska12_u_cska22_fa8_xor1 = s_dadda_cska12_u_cska22_fa8_xor0 ^ s_dadda_cska12_u_cska22_fa7_or0;
  assign s_dadda_cska12_u_cska22_fa8_and1 = s_dadda_cska12_u_cska22_fa8_xor0 & s_dadda_cska12_u_cska22_fa7_or0;
  assign s_dadda_cska12_u_cska22_fa8_or0 = s_dadda_cska12_u_cska22_fa8_and0 | s_dadda_cska12_u_cska22_fa8_and1;
  assign s_dadda_cska12_u_cska22_xor10 = s_dadda_cska12_fa71_xor1 ^ s_dadda_cska12_fa89_xor1;
  assign s_dadda_cska12_u_cska22_fa9_xor0 = s_dadda_cska12_fa71_xor1 ^ s_dadda_cska12_fa89_xor1;
  assign s_dadda_cska12_u_cska22_fa9_and0 = s_dadda_cska12_fa71_xor1 & s_dadda_cska12_fa89_xor1;
  assign s_dadda_cska12_u_cska22_fa9_xor1 = s_dadda_cska12_u_cska22_fa9_xor0 ^ s_dadda_cska12_u_cska22_fa8_or0;
  assign s_dadda_cska12_u_cska22_fa9_and1 = s_dadda_cska12_u_cska22_fa9_xor0 & s_dadda_cska12_u_cska22_fa8_or0;
  assign s_dadda_cska12_u_cska22_fa9_or0 = s_dadda_cska12_u_cska22_fa9_and0 | s_dadda_cska12_u_cska22_fa9_and1;
  assign s_dadda_cska12_u_cska22_xor11 = s_dadda_cska12_fa72_xor1 ^ s_dadda_cska12_fa90_xor1;
  assign s_dadda_cska12_u_cska22_fa10_xor0 = s_dadda_cska12_fa72_xor1 ^ s_dadda_cska12_fa90_xor1;
  assign s_dadda_cska12_u_cska22_fa10_and0 = s_dadda_cska12_fa72_xor1 & s_dadda_cska12_fa90_xor1;
  assign s_dadda_cska12_u_cska22_fa10_xor1 = s_dadda_cska12_u_cska22_fa10_xor0 ^ s_dadda_cska12_u_cska22_fa9_or0;
  assign s_dadda_cska12_u_cska22_fa10_and1 = s_dadda_cska12_u_cska22_fa10_xor0 & s_dadda_cska12_u_cska22_fa9_or0;
  assign s_dadda_cska12_u_cska22_fa10_or0 = s_dadda_cska12_u_cska22_fa10_and0 | s_dadda_cska12_u_cska22_fa10_and1;
  assign s_dadda_cska12_u_cska22_and_propagate26 = s_dadda_cska12_u_cska22_xor8 & s_dadda_cska12_u_cska22_xor10;
  assign s_dadda_cska12_u_cska22_and_propagate27 = s_dadda_cska12_u_cska22_xor9 & s_dadda_cska12_u_cska22_xor11;
  assign s_dadda_cska12_u_cska22_and_propagate28 = s_dadda_cska12_u_cska22_and_propagate26 & s_dadda_cska12_u_cska22_and_propagate27;
  assign s_dadda_cska12_u_cska22_mux2to12_and0 = s_dadda_cska12_u_cska22_mux2to11_xor0 & s_dadda_cska12_u_cska22_and_propagate28;
  assign s_dadda_cska12_u_cska22_mux2to12_not0 = ~s_dadda_cska12_u_cska22_and_propagate28;
  assign s_dadda_cska12_u_cska22_mux2to12_and1 = s_dadda_cska12_u_cska22_fa10_or0 & s_dadda_cska12_u_cska22_mux2to12_not0;
  assign s_dadda_cska12_u_cska22_mux2to12_xor0 = s_dadda_cska12_u_cska22_mux2to12_and0 ^ s_dadda_cska12_u_cska22_mux2to12_and1;
  assign s_dadda_cska12_u_cska22_xor12 = s_dadda_cska12_fa73_xor1 ^ s_dadda_cska12_fa91_xor1;
  assign s_dadda_cska12_u_cska22_fa11_xor0 = s_dadda_cska12_fa73_xor1 ^ s_dadda_cska12_fa91_xor1;
  assign s_dadda_cska12_u_cska22_fa11_and0 = s_dadda_cska12_fa73_xor1 & s_dadda_cska12_fa91_xor1;
  assign s_dadda_cska12_u_cska22_fa11_xor1 = s_dadda_cska12_u_cska22_fa11_xor0 ^ s_dadda_cska12_u_cska22_mux2to12_xor0;
  assign s_dadda_cska12_u_cska22_fa11_and1 = s_dadda_cska12_u_cska22_fa11_xor0 & s_dadda_cska12_u_cska22_mux2to12_xor0;
  assign s_dadda_cska12_u_cska22_fa11_or0 = s_dadda_cska12_u_cska22_fa11_and0 | s_dadda_cska12_u_cska22_fa11_and1;
  assign s_dadda_cska12_u_cska22_xor13 = s_dadda_cska12_fa74_xor1 ^ s_dadda_cska12_fa92_xor1;
  assign s_dadda_cska12_u_cska22_fa12_xor0 = s_dadda_cska12_fa74_xor1 ^ s_dadda_cska12_fa92_xor1;
  assign s_dadda_cska12_u_cska22_fa12_and0 = s_dadda_cska12_fa74_xor1 & s_dadda_cska12_fa92_xor1;
  assign s_dadda_cska12_u_cska22_fa12_xor1 = s_dadda_cska12_u_cska22_fa12_xor0 ^ s_dadda_cska12_u_cska22_fa11_or0;
  assign s_dadda_cska12_u_cska22_fa12_and1 = s_dadda_cska12_u_cska22_fa12_xor0 & s_dadda_cska12_u_cska22_fa11_or0;
  assign s_dadda_cska12_u_cska22_fa12_or0 = s_dadda_cska12_u_cska22_fa12_and0 | s_dadda_cska12_u_cska22_fa12_and1;
  assign s_dadda_cska12_u_cska22_xor14 = s_dadda_cska12_fa75_xor1 ^ s_dadda_cska12_fa93_xor1;
  assign s_dadda_cska12_u_cska22_fa13_xor0 = s_dadda_cska12_fa75_xor1 ^ s_dadda_cska12_fa93_xor1;
  assign s_dadda_cska12_u_cska22_fa13_and0 = s_dadda_cska12_fa75_xor1 & s_dadda_cska12_fa93_xor1;
  assign s_dadda_cska12_u_cska22_fa13_xor1 = s_dadda_cska12_u_cska22_fa13_xor0 ^ s_dadda_cska12_u_cska22_fa12_or0;
  assign s_dadda_cska12_u_cska22_fa13_and1 = s_dadda_cska12_u_cska22_fa13_xor0 & s_dadda_cska12_u_cska22_fa12_or0;
  assign s_dadda_cska12_u_cska22_fa13_or0 = s_dadda_cska12_u_cska22_fa13_and0 | s_dadda_cska12_u_cska22_fa13_and1;
  assign s_dadda_cska12_u_cska22_xor15 = s_dadda_cska12_fa76_xor1 ^ s_dadda_cska12_fa94_xor1;
  assign s_dadda_cska12_u_cska22_fa14_xor0 = s_dadda_cska12_fa76_xor1 ^ s_dadda_cska12_fa94_xor1;
  assign s_dadda_cska12_u_cska22_fa14_and0 = s_dadda_cska12_fa76_xor1 & s_dadda_cska12_fa94_xor1;
  assign s_dadda_cska12_u_cska22_fa14_xor1 = s_dadda_cska12_u_cska22_fa14_xor0 ^ s_dadda_cska12_u_cska22_fa13_or0;
  assign s_dadda_cska12_u_cska22_fa14_and1 = s_dadda_cska12_u_cska22_fa14_xor0 & s_dadda_cska12_u_cska22_fa13_or0;
  assign s_dadda_cska12_u_cska22_fa14_or0 = s_dadda_cska12_u_cska22_fa14_and0 | s_dadda_cska12_u_cska22_fa14_and1;
  assign s_dadda_cska12_u_cska22_and_propagate39 = s_dadda_cska12_u_cska22_xor12 & s_dadda_cska12_u_cska22_xor14;
  assign s_dadda_cska12_u_cska22_and_propagate310 = s_dadda_cska12_u_cska22_xor13 & s_dadda_cska12_u_cska22_xor15;
  assign s_dadda_cska12_u_cska22_and_propagate311 = s_dadda_cska12_u_cska22_and_propagate39 & s_dadda_cska12_u_cska22_and_propagate310;
  assign s_dadda_cska12_u_cska22_mux2to13_and0 = s_dadda_cska12_u_cska22_mux2to12_xor0 & s_dadda_cska12_u_cska22_and_propagate311;
  assign s_dadda_cska12_u_cska22_mux2to13_not0 = ~s_dadda_cska12_u_cska22_and_propagate311;
  assign s_dadda_cska12_u_cska22_mux2to13_and1 = s_dadda_cska12_u_cska22_fa14_or0 & s_dadda_cska12_u_cska22_mux2to13_not0;
  assign s_dadda_cska12_u_cska22_mux2to13_xor0 = s_dadda_cska12_u_cska22_mux2to13_and0 ^ s_dadda_cska12_u_cska22_mux2to13_and1;
  assign s_dadda_cska12_u_cska22_xor16 = s_dadda_cska12_fa77_xor1 ^ s_dadda_cska12_fa95_xor1;
  assign s_dadda_cska12_u_cska22_fa15_xor0 = s_dadda_cska12_fa77_xor1 ^ s_dadda_cska12_fa95_xor1;
  assign s_dadda_cska12_u_cska22_fa15_and0 = s_dadda_cska12_fa77_xor1 & s_dadda_cska12_fa95_xor1;
  assign s_dadda_cska12_u_cska22_fa15_xor1 = s_dadda_cska12_u_cska22_fa15_xor0 ^ s_dadda_cska12_u_cska22_mux2to13_xor0;
  assign s_dadda_cska12_u_cska22_fa15_and1 = s_dadda_cska12_u_cska22_fa15_xor0 & s_dadda_cska12_u_cska22_mux2to13_xor0;
  assign s_dadda_cska12_u_cska22_fa15_or0 = s_dadda_cska12_u_cska22_fa15_and0 | s_dadda_cska12_u_cska22_fa15_and1;
  assign s_dadda_cska12_u_cska22_xor17 = s_dadda_cska12_fa78_xor1 ^ s_dadda_cska12_fa96_xor1;
  assign s_dadda_cska12_u_cska22_fa16_xor0 = s_dadda_cska12_fa78_xor1 ^ s_dadda_cska12_fa96_xor1;
  assign s_dadda_cska12_u_cska22_fa16_and0 = s_dadda_cska12_fa78_xor1 & s_dadda_cska12_fa96_xor1;
  assign s_dadda_cska12_u_cska22_fa16_xor1 = s_dadda_cska12_u_cska22_fa16_xor0 ^ s_dadda_cska12_u_cska22_fa15_or0;
  assign s_dadda_cska12_u_cska22_fa16_and1 = s_dadda_cska12_u_cska22_fa16_xor0 & s_dadda_cska12_u_cska22_fa15_or0;
  assign s_dadda_cska12_u_cska22_fa16_or0 = s_dadda_cska12_u_cska22_fa16_and0 | s_dadda_cska12_u_cska22_fa16_and1;
  assign s_dadda_cska12_u_cska22_xor18 = s_dadda_cska12_fa79_xor1 ^ s_dadda_cska12_fa97_xor1;
  assign s_dadda_cska12_u_cska22_fa17_xor0 = s_dadda_cska12_fa79_xor1 ^ s_dadda_cska12_fa97_xor1;
  assign s_dadda_cska12_u_cska22_fa17_and0 = s_dadda_cska12_fa79_xor1 & s_dadda_cska12_fa97_xor1;
  assign s_dadda_cska12_u_cska22_fa17_xor1 = s_dadda_cska12_u_cska22_fa17_xor0 ^ s_dadda_cska12_u_cska22_fa16_or0;
  assign s_dadda_cska12_u_cska22_fa17_and1 = s_dadda_cska12_u_cska22_fa17_xor0 & s_dadda_cska12_u_cska22_fa16_or0;
  assign s_dadda_cska12_u_cska22_fa17_or0 = s_dadda_cska12_u_cska22_fa17_and0 | s_dadda_cska12_u_cska22_fa17_and1;
  assign s_dadda_cska12_u_cska22_xor19 = s_dadda_cska12_fa80_xor1 ^ s_dadda_cska12_fa98_xor1;
  assign s_dadda_cska12_u_cska22_fa18_xor0 = s_dadda_cska12_fa80_xor1 ^ s_dadda_cska12_fa98_xor1;
  assign s_dadda_cska12_u_cska22_fa18_and0 = s_dadda_cska12_fa80_xor1 & s_dadda_cska12_fa98_xor1;
  assign s_dadda_cska12_u_cska22_fa18_xor1 = s_dadda_cska12_u_cska22_fa18_xor0 ^ s_dadda_cska12_u_cska22_fa17_or0;
  assign s_dadda_cska12_u_cska22_fa18_and1 = s_dadda_cska12_u_cska22_fa18_xor0 & s_dadda_cska12_u_cska22_fa17_or0;
  assign s_dadda_cska12_u_cska22_fa18_or0 = s_dadda_cska12_u_cska22_fa18_and0 | s_dadda_cska12_u_cska22_fa18_and1;
  assign s_dadda_cska12_u_cska22_and_propagate412 = s_dadda_cska12_u_cska22_xor16 & s_dadda_cska12_u_cska22_xor18;
  assign s_dadda_cska12_u_cska22_and_propagate413 = s_dadda_cska12_u_cska22_xor17 & s_dadda_cska12_u_cska22_xor19;
  assign s_dadda_cska12_u_cska22_and_propagate414 = s_dadda_cska12_u_cska22_and_propagate412 & s_dadda_cska12_u_cska22_and_propagate413;
  assign s_dadda_cska12_u_cska22_mux2to14_and0 = s_dadda_cska12_u_cska22_mux2to13_xor0 & s_dadda_cska12_u_cska22_and_propagate414;
  assign s_dadda_cska12_u_cska22_mux2to14_not0 = ~s_dadda_cska12_u_cska22_and_propagate414;
  assign s_dadda_cska12_u_cska22_mux2to14_and1 = s_dadda_cska12_u_cska22_fa18_or0 & s_dadda_cska12_u_cska22_mux2to14_not0;
  assign s_dadda_cska12_u_cska22_mux2to14_xor0 = s_dadda_cska12_u_cska22_mux2to14_and0 ^ s_dadda_cska12_u_cska22_mux2to14_and1;
  assign s_dadda_cska12_u_cska22_xor20 = s_dadda_cska12_nand_10_11 ^ s_dadda_cska12_fa99_xor1;
  assign s_dadda_cska12_u_cska22_fa19_xor0 = s_dadda_cska12_nand_10_11 ^ s_dadda_cska12_fa99_xor1;
  assign s_dadda_cska12_u_cska22_fa19_and0 = s_dadda_cska12_nand_10_11 & s_dadda_cska12_fa99_xor1;
  assign s_dadda_cska12_u_cska22_fa19_xor1 = s_dadda_cska12_u_cska22_fa19_xor0 ^ s_dadda_cska12_u_cska22_mux2to14_xor0;
  assign s_dadda_cska12_u_cska22_fa19_and1 = s_dadda_cska12_u_cska22_fa19_xor0 & s_dadda_cska12_u_cska22_mux2to14_xor0;
  assign s_dadda_cska12_u_cska22_fa19_or0 = s_dadda_cska12_u_cska22_fa19_and0 | s_dadda_cska12_u_cska22_fa19_and1;
  assign s_dadda_cska12_u_cska22_xor21 = s_dadda_cska12_fa99_or0 ^ s_dadda_cska12_and_11_11;
  assign s_dadda_cska12_u_cska22_fa20_xor0 = s_dadda_cska12_fa99_or0 ^ s_dadda_cska12_and_11_11;
  assign s_dadda_cska12_u_cska22_fa20_and0 = s_dadda_cska12_fa99_or0 & s_dadda_cska12_and_11_11;
  assign s_dadda_cska12_u_cska22_fa20_xor1 = s_dadda_cska12_u_cska22_fa20_xor0 ^ s_dadda_cska12_u_cska22_fa19_or0;
  assign s_dadda_cska12_u_cska22_fa20_and1 = s_dadda_cska12_u_cska22_fa20_xor0 & s_dadda_cska12_u_cska22_fa19_or0;
  assign s_dadda_cska12_u_cska22_fa20_or0 = s_dadda_cska12_u_cska22_fa20_and0 | s_dadda_cska12_u_cska22_fa20_and1;
  assign s_dadda_cska12_u_cska22_and_propagate515 = s_dadda_cska12_u_cska22_xor20 & s_dadda_cska12_u_cska22_xor21;
  assign s_dadda_cska12_u_cska22_mux2to15_and0 = s_dadda_cska12_u_cska22_mux2to14_xor0 & s_dadda_cska12_u_cska22_and_propagate515;
  assign s_dadda_cska12_u_cska22_mux2to15_not0 = ~s_dadda_cska12_u_cska22_and_propagate515;
  assign s_dadda_cska12_u_cska22_mux2to15_and1 = s_dadda_cska12_u_cska22_fa20_or0 & s_dadda_cska12_u_cska22_mux2to15_not0;
  assign s_dadda_cska12_u_cska22_mux2to15_xor0 = s_dadda_cska12_u_cska22_mux2to15_and0 ^ s_dadda_cska12_u_cska22_mux2to15_and1;
  assign s_dadda_cska12_xor0 = ~s_dadda_cska12_u_cska22_mux2to15_xor0;

  assign s_dadda_cska12_out[0] = s_dadda_cska12_and_0_0;
  assign s_dadda_cska12_out[1] = s_dadda_cska12_u_cska22_ha0_xor0;
  assign s_dadda_cska12_out[2] = s_dadda_cska12_u_cska22_fa0_xor1;
  assign s_dadda_cska12_out[3] = s_dadda_cska12_u_cska22_fa1_xor1;
  assign s_dadda_cska12_out[4] = s_dadda_cska12_u_cska22_fa2_xor1;
  assign s_dadda_cska12_out[5] = s_dadda_cska12_u_cska22_fa3_xor1;
  assign s_dadda_cska12_out[6] = s_dadda_cska12_u_cska22_fa4_xor1;
  assign s_dadda_cska12_out[7] = s_dadda_cska12_u_cska22_fa5_xor1;
  assign s_dadda_cska12_out[8] = s_dadda_cska12_u_cska22_fa6_xor1;
  assign s_dadda_cska12_out[9] = s_dadda_cska12_u_cska22_fa7_xor1;
  assign s_dadda_cska12_out[10] = s_dadda_cska12_u_cska22_fa8_xor1;
  assign s_dadda_cska12_out[11] = s_dadda_cska12_u_cska22_fa9_xor1;
  assign s_dadda_cska12_out[12] = s_dadda_cska12_u_cska22_fa10_xor1;
  assign s_dadda_cska12_out[13] = s_dadda_cska12_u_cska22_fa11_xor1;
  assign s_dadda_cska12_out[14] = s_dadda_cska12_u_cska22_fa12_xor1;
  assign s_dadda_cska12_out[15] = s_dadda_cska12_u_cska22_fa13_xor1;
  assign s_dadda_cska12_out[16] = s_dadda_cska12_u_cska22_fa14_xor1;
  assign s_dadda_cska12_out[17] = s_dadda_cska12_u_cska22_fa15_xor1;
  assign s_dadda_cska12_out[18] = s_dadda_cska12_u_cska22_fa16_xor1;
  assign s_dadda_cska12_out[19] = s_dadda_cska12_u_cska22_fa17_xor1;
  assign s_dadda_cska12_out[20] = s_dadda_cska12_u_cska22_fa18_xor1;
  assign s_dadda_cska12_out[21] = s_dadda_cska12_u_cska22_fa19_xor1;
  assign s_dadda_cska12_out[22] = s_dadda_cska12_u_cska22_fa20_xor1;
  assign s_dadda_cska12_out[23] = s_dadda_cska12_xor0;
endmodule