module s_dadda_pg_rca24(input [23:0] a, input [23:0] b, output [47:0] s_dadda_pg_rca24_out);
  wire s_dadda_pg_rca24_and_19_0;
  wire s_dadda_pg_rca24_and_18_1;
  wire s_dadda_pg_rca24_ha0_xor0;
  wire s_dadda_pg_rca24_ha0_and0;
  wire s_dadda_pg_rca24_and_20_0;
  wire s_dadda_pg_rca24_and_19_1;
  wire s_dadda_pg_rca24_fa0_xor0;
  wire s_dadda_pg_rca24_fa0_and0;
  wire s_dadda_pg_rca24_fa0_xor1;
  wire s_dadda_pg_rca24_fa0_and1;
  wire s_dadda_pg_rca24_fa0_or0;
  wire s_dadda_pg_rca24_and_18_2;
  wire s_dadda_pg_rca24_and_17_3;
  wire s_dadda_pg_rca24_ha1_xor0;
  wire s_dadda_pg_rca24_ha1_and0;
  wire s_dadda_pg_rca24_and_21_0;
  wire s_dadda_pg_rca24_fa1_xor0;
  wire s_dadda_pg_rca24_fa1_and0;
  wire s_dadda_pg_rca24_fa1_xor1;
  wire s_dadda_pg_rca24_fa1_and1;
  wire s_dadda_pg_rca24_fa1_or0;
  wire s_dadda_pg_rca24_and_20_1;
  wire s_dadda_pg_rca24_and_19_2;
  wire s_dadda_pg_rca24_and_18_3;
  wire s_dadda_pg_rca24_fa2_xor0;
  wire s_dadda_pg_rca24_fa2_and0;
  wire s_dadda_pg_rca24_fa2_xor1;
  wire s_dadda_pg_rca24_fa2_and1;
  wire s_dadda_pg_rca24_fa2_or0;
  wire s_dadda_pg_rca24_and_17_4;
  wire s_dadda_pg_rca24_and_16_5;
  wire s_dadda_pg_rca24_ha2_xor0;
  wire s_dadda_pg_rca24_ha2_and0;
  wire s_dadda_pg_rca24_fa3_xor0;
  wire s_dadda_pg_rca24_fa3_and0;
  wire s_dadda_pg_rca24_fa3_xor1;
  wire s_dadda_pg_rca24_fa3_and1;
  wire s_dadda_pg_rca24_fa3_or0;
  wire s_dadda_pg_rca24_and_22_0;
  wire s_dadda_pg_rca24_and_21_1;
  wire s_dadda_pg_rca24_and_20_2;
  wire s_dadda_pg_rca24_fa4_xor0;
  wire s_dadda_pg_rca24_fa4_and0;
  wire s_dadda_pg_rca24_fa4_xor1;
  wire s_dadda_pg_rca24_fa4_and1;
  wire s_dadda_pg_rca24_fa4_or0;
  wire s_dadda_pg_rca24_and_19_3;
  wire s_dadda_pg_rca24_and_18_4;
  wire s_dadda_pg_rca24_and_17_5;
  wire s_dadda_pg_rca24_fa5_xor0;
  wire s_dadda_pg_rca24_fa5_and0;
  wire s_dadda_pg_rca24_fa5_xor1;
  wire s_dadda_pg_rca24_fa5_and1;
  wire s_dadda_pg_rca24_fa5_or0;
  wire s_dadda_pg_rca24_and_16_6;
  wire s_dadda_pg_rca24_and_15_7;
  wire s_dadda_pg_rca24_ha3_xor0;
  wire s_dadda_pg_rca24_ha3_and0;
  wire s_dadda_pg_rca24_fa6_xor0;
  wire s_dadda_pg_rca24_fa6_and0;
  wire s_dadda_pg_rca24_fa6_xor1;
  wire s_dadda_pg_rca24_fa6_and1;
  wire s_dadda_pg_rca24_fa6_or0;
  wire s_dadda_pg_rca24_nand_23_0;
  wire s_dadda_pg_rca24_and_22_1;
  wire s_dadda_pg_rca24_fa7_xor0;
  wire s_dadda_pg_rca24_fa7_and0;
  wire s_dadda_pg_rca24_fa7_xor1;
  wire s_dadda_pg_rca24_fa7_and1;
  wire s_dadda_pg_rca24_fa7_or0;
  wire s_dadda_pg_rca24_and_21_2;
  wire s_dadda_pg_rca24_and_20_3;
  wire s_dadda_pg_rca24_and_19_4;
  wire s_dadda_pg_rca24_fa8_xor0;
  wire s_dadda_pg_rca24_fa8_and0;
  wire s_dadda_pg_rca24_fa8_xor1;
  wire s_dadda_pg_rca24_fa8_and1;
  wire s_dadda_pg_rca24_fa8_or0;
  wire s_dadda_pg_rca24_and_18_5;
  wire s_dadda_pg_rca24_and_17_6;
  wire s_dadda_pg_rca24_and_16_7;
  wire s_dadda_pg_rca24_fa9_xor0;
  wire s_dadda_pg_rca24_fa9_and0;
  wire s_dadda_pg_rca24_fa9_xor1;
  wire s_dadda_pg_rca24_fa9_and1;
  wire s_dadda_pg_rca24_fa9_or0;
  wire s_dadda_pg_rca24_and_15_8;
  wire s_dadda_pg_rca24_and_14_9;
  wire s_dadda_pg_rca24_ha4_xor0;
  wire s_dadda_pg_rca24_ha4_and0;
  wire s_dadda_pg_rca24_fa10_xor0;
  wire s_dadda_pg_rca24_fa10_and0;
  wire s_dadda_pg_rca24_fa10_xor1;
  wire s_dadda_pg_rca24_fa10_and1;
  wire s_dadda_pg_rca24_fa10_or0;
  wire s_dadda_pg_rca24_fa11_xor0;
  wire s_dadda_pg_rca24_fa11_and0;
  wire s_dadda_pg_rca24_fa11_xor1;
  wire s_dadda_pg_rca24_fa11_or0;
  wire s_dadda_pg_rca24_nand_23_1;
  wire s_dadda_pg_rca24_and_22_2;
  wire s_dadda_pg_rca24_and_21_3;
  wire s_dadda_pg_rca24_fa12_xor0;
  wire s_dadda_pg_rca24_fa12_and0;
  wire s_dadda_pg_rca24_fa12_xor1;
  wire s_dadda_pg_rca24_fa12_and1;
  wire s_dadda_pg_rca24_fa12_or0;
  wire s_dadda_pg_rca24_and_20_4;
  wire s_dadda_pg_rca24_and_19_5;
  wire s_dadda_pg_rca24_and_18_6;
  wire s_dadda_pg_rca24_fa13_xor0;
  wire s_dadda_pg_rca24_fa13_and0;
  wire s_dadda_pg_rca24_fa13_xor1;
  wire s_dadda_pg_rca24_fa13_and1;
  wire s_dadda_pg_rca24_fa13_or0;
  wire s_dadda_pg_rca24_and_17_7;
  wire s_dadda_pg_rca24_and_16_8;
  wire s_dadda_pg_rca24_and_15_9;
  wire s_dadda_pg_rca24_fa14_xor0;
  wire s_dadda_pg_rca24_fa14_and0;
  wire s_dadda_pg_rca24_fa14_xor1;
  wire s_dadda_pg_rca24_fa14_and1;
  wire s_dadda_pg_rca24_fa14_or0;
  wire s_dadda_pg_rca24_fa15_xor0;
  wire s_dadda_pg_rca24_fa15_and0;
  wire s_dadda_pg_rca24_fa15_xor1;
  wire s_dadda_pg_rca24_fa15_and1;
  wire s_dadda_pg_rca24_fa15_or0;
  wire s_dadda_pg_rca24_nand_23_2;
  wire s_dadda_pg_rca24_fa16_xor0;
  wire s_dadda_pg_rca24_fa16_and0;
  wire s_dadda_pg_rca24_fa16_xor1;
  wire s_dadda_pg_rca24_fa16_and1;
  wire s_dadda_pg_rca24_fa16_or0;
  wire s_dadda_pg_rca24_and_22_3;
  wire s_dadda_pg_rca24_and_21_4;
  wire s_dadda_pg_rca24_and_20_5;
  wire s_dadda_pg_rca24_fa17_xor0;
  wire s_dadda_pg_rca24_fa17_and0;
  wire s_dadda_pg_rca24_fa17_xor1;
  wire s_dadda_pg_rca24_fa17_and1;
  wire s_dadda_pg_rca24_fa17_or0;
  wire s_dadda_pg_rca24_and_19_6;
  wire s_dadda_pg_rca24_and_18_7;
  wire s_dadda_pg_rca24_and_17_8;
  wire s_dadda_pg_rca24_fa18_xor0;
  wire s_dadda_pg_rca24_fa18_and0;
  wire s_dadda_pg_rca24_fa18_xor1;
  wire s_dadda_pg_rca24_fa18_and1;
  wire s_dadda_pg_rca24_fa18_or0;
  wire s_dadda_pg_rca24_fa19_xor0;
  wire s_dadda_pg_rca24_fa19_and0;
  wire s_dadda_pg_rca24_fa19_xor1;
  wire s_dadda_pg_rca24_fa19_and1;
  wire s_dadda_pg_rca24_fa19_or0;
  wire s_dadda_pg_rca24_nand_23_3;
  wire s_dadda_pg_rca24_and_22_4;
  wire s_dadda_pg_rca24_fa20_xor0;
  wire s_dadda_pg_rca24_fa20_and0;
  wire s_dadda_pg_rca24_fa20_xor1;
  wire s_dadda_pg_rca24_fa20_and1;
  wire s_dadda_pg_rca24_fa20_or0;
  wire s_dadda_pg_rca24_and_21_5;
  wire s_dadda_pg_rca24_and_20_6;
  wire s_dadda_pg_rca24_and_19_7;
  wire s_dadda_pg_rca24_fa21_xor0;
  wire s_dadda_pg_rca24_fa21_and0;
  wire s_dadda_pg_rca24_fa21_xor1;
  wire s_dadda_pg_rca24_fa21_and1;
  wire s_dadda_pg_rca24_fa21_or0;
  wire s_dadda_pg_rca24_fa22_xor0;
  wire s_dadda_pg_rca24_fa22_and0;
  wire s_dadda_pg_rca24_fa22_xor1;
  wire s_dadda_pg_rca24_fa22_and1;
  wire s_dadda_pg_rca24_fa22_or0;
  wire s_dadda_pg_rca24_nand_23_4;
  wire s_dadda_pg_rca24_and_22_5;
  wire s_dadda_pg_rca24_and_21_6;
  wire s_dadda_pg_rca24_fa23_xor0;
  wire s_dadda_pg_rca24_fa23_and0;
  wire s_dadda_pg_rca24_fa23_xor1;
  wire s_dadda_pg_rca24_fa23_and1;
  wire s_dadda_pg_rca24_fa23_or0;
  wire s_dadda_pg_rca24_nand_23_5;
  wire s_dadda_pg_rca24_fa24_xor0;
  wire s_dadda_pg_rca24_fa24_and0;
  wire s_dadda_pg_rca24_fa24_xor1;
  wire s_dadda_pg_rca24_fa24_and1;
  wire s_dadda_pg_rca24_fa24_or0;
  wire s_dadda_pg_rca24_and_6_0;
  wire s_dadda_pg_rca24_and_5_1;
  wire s_dadda_pg_rca24_ha5_xor0;
  wire s_dadda_pg_rca24_ha5_and0;
  wire s_dadda_pg_rca24_and_7_0;
  wire s_dadda_pg_rca24_and_6_1;
  wire s_dadda_pg_rca24_fa25_xor0;
  wire s_dadda_pg_rca24_fa25_and0;
  wire s_dadda_pg_rca24_fa25_xor1;
  wire s_dadda_pg_rca24_fa25_and1;
  wire s_dadda_pg_rca24_fa25_or0;
  wire s_dadda_pg_rca24_and_5_2;
  wire s_dadda_pg_rca24_and_4_3;
  wire s_dadda_pg_rca24_ha6_xor0;
  wire s_dadda_pg_rca24_ha6_and0;
  wire s_dadda_pg_rca24_and_8_0;
  wire s_dadda_pg_rca24_fa26_xor0;
  wire s_dadda_pg_rca24_fa26_and0;
  wire s_dadda_pg_rca24_fa26_xor1;
  wire s_dadda_pg_rca24_fa26_and1;
  wire s_dadda_pg_rca24_fa26_or0;
  wire s_dadda_pg_rca24_and_7_1;
  wire s_dadda_pg_rca24_and_6_2;
  wire s_dadda_pg_rca24_and_5_3;
  wire s_dadda_pg_rca24_fa27_xor0;
  wire s_dadda_pg_rca24_fa27_and0;
  wire s_dadda_pg_rca24_fa27_xor1;
  wire s_dadda_pg_rca24_fa27_and1;
  wire s_dadda_pg_rca24_fa27_or0;
  wire s_dadda_pg_rca24_and_4_4;
  wire s_dadda_pg_rca24_and_3_5;
  wire s_dadda_pg_rca24_ha7_xor0;
  wire s_dadda_pg_rca24_ha7_and0;
  wire s_dadda_pg_rca24_fa28_xor0;
  wire s_dadda_pg_rca24_fa28_and0;
  wire s_dadda_pg_rca24_fa28_xor1;
  wire s_dadda_pg_rca24_fa28_and1;
  wire s_dadda_pg_rca24_fa28_or0;
  wire s_dadda_pg_rca24_and_9_0;
  wire s_dadda_pg_rca24_and_8_1;
  wire s_dadda_pg_rca24_and_7_2;
  wire s_dadda_pg_rca24_fa29_xor0;
  wire s_dadda_pg_rca24_fa29_and0;
  wire s_dadda_pg_rca24_fa29_xor1;
  wire s_dadda_pg_rca24_fa29_and1;
  wire s_dadda_pg_rca24_fa29_or0;
  wire s_dadda_pg_rca24_and_6_3;
  wire s_dadda_pg_rca24_and_5_4;
  wire s_dadda_pg_rca24_and_4_5;
  wire s_dadda_pg_rca24_fa30_xor0;
  wire s_dadda_pg_rca24_fa30_and0;
  wire s_dadda_pg_rca24_fa30_xor1;
  wire s_dadda_pg_rca24_fa30_and1;
  wire s_dadda_pg_rca24_fa30_or0;
  wire s_dadda_pg_rca24_and_3_6;
  wire s_dadda_pg_rca24_and_2_7;
  wire s_dadda_pg_rca24_ha8_xor0;
  wire s_dadda_pg_rca24_ha8_and0;
  wire s_dadda_pg_rca24_fa31_xor0;
  wire s_dadda_pg_rca24_fa31_and0;
  wire s_dadda_pg_rca24_fa31_xor1;
  wire s_dadda_pg_rca24_fa31_and1;
  wire s_dadda_pg_rca24_fa31_or0;
  wire s_dadda_pg_rca24_and_10_0;
  wire s_dadda_pg_rca24_and_9_1;
  wire s_dadda_pg_rca24_fa32_xor0;
  wire s_dadda_pg_rca24_fa32_and0;
  wire s_dadda_pg_rca24_fa32_xor1;
  wire s_dadda_pg_rca24_fa32_and1;
  wire s_dadda_pg_rca24_fa32_or0;
  wire s_dadda_pg_rca24_and_8_2;
  wire s_dadda_pg_rca24_and_7_3;
  wire s_dadda_pg_rca24_and_6_4;
  wire s_dadda_pg_rca24_fa33_xor0;
  wire s_dadda_pg_rca24_fa33_and0;
  wire s_dadda_pg_rca24_fa33_xor1;
  wire s_dadda_pg_rca24_fa33_and1;
  wire s_dadda_pg_rca24_fa33_or0;
  wire s_dadda_pg_rca24_and_5_5;
  wire s_dadda_pg_rca24_and_4_6;
  wire s_dadda_pg_rca24_and_3_7;
  wire s_dadda_pg_rca24_fa34_xor0;
  wire s_dadda_pg_rca24_fa34_and0;
  wire s_dadda_pg_rca24_fa34_xor1;
  wire s_dadda_pg_rca24_fa34_and1;
  wire s_dadda_pg_rca24_fa34_or0;
  wire s_dadda_pg_rca24_and_2_8;
  wire s_dadda_pg_rca24_and_1_9;
  wire s_dadda_pg_rca24_ha9_xor0;
  wire s_dadda_pg_rca24_ha9_and0;
  wire s_dadda_pg_rca24_fa35_xor0;
  wire s_dadda_pg_rca24_fa35_and0;
  wire s_dadda_pg_rca24_fa35_xor1;
  wire s_dadda_pg_rca24_fa35_and1;
  wire s_dadda_pg_rca24_fa35_or0;
  wire s_dadda_pg_rca24_and_11_0;
  wire s_dadda_pg_rca24_fa36_xor0;
  wire s_dadda_pg_rca24_fa36_and0;
  wire s_dadda_pg_rca24_fa36_xor1;
  wire s_dadda_pg_rca24_fa36_and1;
  wire s_dadda_pg_rca24_fa36_or0;
  wire s_dadda_pg_rca24_and_10_1;
  wire s_dadda_pg_rca24_and_9_2;
  wire s_dadda_pg_rca24_and_8_3;
  wire s_dadda_pg_rca24_fa37_xor0;
  wire s_dadda_pg_rca24_fa37_and0;
  wire s_dadda_pg_rca24_fa37_xor1;
  wire s_dadda_pg_rca24_fa37_and1;
  wire s_dadda_pg_rca24_fa37_or0;
  wire s_dadda_pg_rca24_and_7_4;
  wire s_dadda_pg_rca24_and_6_5;
  wire s_dadda_pg_rca24_and_5_6;
  wire s_dadda_pg_rca24_fa38_xor0;
  wire s_dadda_pg_rca24_fa38_and0;
  wire s_dadda_pg_rca24_fa38_xor1;
  wire s_dadda_pg_rca24_fa38_and1;
  wire s_dadda_pg_rca24_fa38_or0;
  wire s_dadda_pg_rca24_and_4_7;
  wire s_dadda_pg_rca24_and_3_8;
  wire s_dadda_pg_rca24_and_2_9;
  wire s_dadda_pg_rca24_fa39_xor0;
  wire s_dadda_pg_rca24_fa39_and0;
  wire s_dadda_pg_rca24_fa39_xor1;
  wire s_dadda_pg_rca24_fa39_and1;
  wire s_dadda_pg_rca24_fa39_or0;
  wire s_dadda_pg_rca24_and_1_10;
  wire s_dadda_pg_rca24_and_0_11;
  wire s_dadda_pg_rca24_ha10_xor0;
  wire s_dadda_pg_rca24_ha10_and0;
  wire s_dadda_pg_rca24_fa40_xor0;
  wire s_dadda_pg_rca24_fa40_and0;
  wire s_dadda_pg_rca24_fa40_xor1;
  wire s_dadda_pg_rca24_fa40_and1;
  wire s_dadda_pg_rca24_fa40_or0;
  wire s_dadda_pg_rca24_fa41_xor0;
  wire s_dadda_pg_rca24_fa41_and0;
  wire s_dadda_pg_rca24_fa41_xor1;
  wire s_dadda_pg_rca24_fa41_and1;
  wire s_dadda_pg_rca24_fa41_or0;
  wire s_dadda_pg_rca24_and_12_0;
  wire s_dadda_pg_rca24_and_11_1;
  wire s_dadda_pg_rca24_and_10_2;
  wire s_dadda_pg_rca24_fa42_xor0;
  wire s_dadda_pg_rca24_fa42_and0;
  wire s_dadda_pg_rca24_fa42_xor1;
  wire s_dadda_pg_rca24_fa42_and1;
  wire s_dadda_pg_rca24_fa42_or0;
  wire s_dadda_pg_rca24_and_9_3;
  wire s_dadda_pg_rca24_and_8_4;
  wire s_dadda_pg_rca24_and_7_5;
  wire s_dadda_pg_rca24_fa43_xor0;
  wire s_dadda_pg_rca24_fa43_and0;
  wire s_dadda_pg_rca24_fa43_xor1;
  wire s_dadda_pg_rca24_fa43_and1;
  wire s_dadda_pg_rca24_fa43_or0;
  wire s_dadda_pg_rca24_and_6_6;
  wire s_dadda_pg_rca24_and_5_7;
  wire s_dadda_pg_rca24_and_4_8;
  wire s_dadda_pg_rca24_fa44_xor0;
  wire s_dadda_pg_rca24_fa44_and0;
  wire s_dadda_pg_rca24_fa44_xor1;
  wire s_dadda_pg_rca24_fa44_and1;
  wire s_dadda_pg_rca24_fa44_or0;
  wire s_dadda_pg_rca24_and_3_9;
  wire s_dadda_pg_rca24_and_2_10;
  wire s_dadda_pg_rca24_and_1_11;
  wire s_dadda_pg_rca24_fa45_xor0;
  wire s_dadda_pg_rca24_fa45_and0;
  wire s_dadda_pg_rca24_fa45_xor1;
  wire s_dadda_pg_rca24_fa45_and1;
  wire s_dadda_pg_rca24_fa45_or0;
  wire s_dadda_pg_rca24_and_0_12;
  wire s_dadda_pg_rca24_ha11_xor0;
  wire s_dadda_pg_rca24_ha11_and0;
  wire s_dadda_pg_rca24_fa46_xor0;
  wire s_dadda_pg_rca24_fa46_and0;
  wire s_dadda_pg_rca24_fa46_xor1;
  wire s_dadda_pg_rca24_fa46_and1;
  wire s_dadda_pg_rca24_fa46_or0;
  wire s_dadda_pg_rca24_fa47_xor0;
  wire s_dadda_pg_rca24_fa47_and0;
  wire s_dadda_pg_rca24_fa47_xor1;
  wire s_dadda_pg_rca24_fa47_and1;
  wire s_dadda_pg_rca24_fa47_or0;
  wire s_dadda_pg_rca24_and_13_0;
  wire s_dadda_pg_rca24_and_12_1;
  wire s_dadda_pg_rca24_fa48_xor0;
  wire s_dadda_pg_rca24_fa48_and0;
  wire s_dadda_pg_rca24_fa48_xor1;
  wire s_dadda_pg_rca24_fa48_and1;
  wire s_dadda_pg_rca24_fa48_or0;
  wire s_dadda_pg_rca24_and_11_2;
  wire s_dadda_pg_rca24_and_10_3;
  wire s_dadda_pg_rca24_and_9_4;
  wire s_dadda_pg_rca24_fa49_xor0;
  wire s_dadda_pg_rca24_fa49_and0;
  wire s_dadda_pg_rca24_fa49_xor1;
  wire s_dadda_pg_rca24_fa49_and1;
  wire s_dadda_pg_rca24_fa49_or0;
  wire s_dadda_pg_rca24_and_8_5;
  wire s_dadda_pg_rca24_and_7_6;
  wire s_dadda_pg_rca24_and_6_7;
  wire s_dadda_pg_rca24_fa50_xor0;
  wire s_dadda_pg_rca24_fa50_and0;
  wire s_dadda_pg_rca24_fa50_xor1;
  wire s_dadda_pg_rca24_fa50_and1;
  wire s_dadda_pg_rca24_fa50_or0;
  wire s_dadda_pg_rca24_and_5_8;
  wire s_dadda_pg_rca24_and_4_9;
  wire s_dadda_pg_rca24_and_3_10;
  wire s_dadda_pg_rca24_fa51_xor0;
  wire s_dadda_pg_rca24_fa51_and0;
  wire s_dadda_pg_rca24_fa51_xor1;
  wire s_dadda_pg_rca24_fa51_and1;
  wire s_dadda_pg_rca24_fa51_or0;
  wire s_dadda_pg_rca24_and_2_11;
  wire s_dadda_pg_rca24_and_1_12;
  wire s_dadda_pg_rca24_and_0_13;
  wire s_dadda_pg_rca24_fa52_xor0;
  wire s_dadda_pg_rca24_fa52_and0;
  wire s_dadda_pg_rca24_fa52_xor1;
  wire s_dadda_pg_rca24_fa52_and1;
  wire s_dadda_pg_rca24_fa52_or0;
  wire s_dadda_pg_rca24_ha12_xor0;
  wire s_dadda_pg_rca24_ha12_and0;
  wire s_dadda_pg_rca24_fa53_xor0;
  wire s_dadda_pg_rca24_fa53_and0;
  wire s_dadda_pg_rca24_fa53_xor1;
  wire s_dadda_pg_rca24_fa53_and1;
  wire s_dadda_pg_rca24_fa53_or0;
  wire s_dadda_pg_rca24_fa54_xor0;
  wire s_dadda_pg_rca24_fa54_and0;
  wire s_dadda_pg_rca24_fa54_xor1;
  wire s_dadda_pg_rca24_fa54_and1;
  wire s_dadda_pg_rca24_fa54_or0;
  wire s_dadda_pg_rca24_and_14_0;
  wire s_dadda_pg_rca24_fa55_xor0;
  wire s_dadda_pg_rca24_fa55_and0;
  wire s_dadda_pg_rca24_fa55_xor1;
  wire s_dadda_pg_rca24_fa55_and1;
  wire s_dadda_pg_rca24_fa55_or0;
  wire s_dadda_pg_rca24_and_13_1;
  wire s_dadda_pg_rca24_and_12_2;
  wire s_dadda_pg_rca24_and_11_3;
  wire s_dadda_pg_rca24_fa56_xor0;
  wire s_dadda_pg_rca24_fa56_and0;
  wire s_dadda_pg_rca24_fa56_xor1;
  wire s_dadda_pg_rca24_fa56_and1;
  wire s_dadda_pg_rca24_fa56_or0;
  wire s_dadda_pg_rca24_and_10_4;
  wire s_dadda_pg_rca24_and_9_5;
  wire s_dadda_pg_rca24_and_8_6;
  wire s_dadda_pg_rca24_fa57_xor0;
  wire s_dadda_pg_rca24_fa57_and0;
  wire s_dadda_pg_rca24_fa57_xor1;
  wire s_dadda_pg_rca24_fa57_and1;
  wire s_dadda_pg_rca24_fa57_or0;
  wire s_dadda_pg_rca24_and_7_7;
  wire s_dadda_pg_rca24_and_6_8;
  wire s_dadda_pg_rca24_and_5_9;
  wire s_dadda_pg_rca24_fa58_xor0;
  wire s_dadda_pg_rca24_fa58_and0;
  wire s_dadda_pg_rca24_fa58_xor1;
  wire s_dadda_pg_rca24_fa58_and1;
  wire s_dadda_pg_rca24_fa58_or0;
  wire s_dadda_pg_rca24_and_4_10;
  wire s_dadda_pg_rca24_and_3_11;
  wire s_dadda_pg_rca24_and_2_12;
  wire s_dadda_pg_rca24_fa59_xor0;
  wire s_dadda_pg_rca24_fa59_and0;
  wire s_dadda_pg_rca24_fa59_xor1;
  wire s_dadda_pg_rca24_fa59_and1;
  wire s_dadda_pg_rca24_fa59_or0;
  wire s_dadda_pg_rca24_and_1_13;
  wire s_dadda_pg_rca24_and_0_14;
  wire s_dadda_pg_rca24_fa60_xor0;
  wire s_dadda_pg_rca24_fa60_and0;
  wire s_dadda_pg_rca24_fa60_xor1;
  wire s_dadda_pg_rca24_fa60_and1;
  wire s_dadda_pg_rca24_fa60_or0;
  wire s_dadda_pg_rca24_ha13_xor0;
  wire s_dadda_pg_rca24_ha13_and0;
  wire s_dadda_pg_rca24_fa61_xor0;
  wire s_dadda_pg_rca24_fa61_and0;
  wire s_dadda_pg_rca24_fa61_xor1;
  wire s_dadda_pg_rca24_fa61_and1;
  wire s_dadda_pg_rca24_fa61_or0;
  wire s_dadda_pg_rca24_fa62_xor0;
  wire s_dadda_pg_rca24_fa62_and0;
  wire s_dadda_pg_rca24_fa62_xor1;
  wire s_dadda_pg_rca24_fa62_and1;
  wire s_dadda_pg_rca24_fa62_or0;
  wire s_dadda_pg_rca24_fa63_xor0;
  wire s_dadda_pg_rca24_fa63_and0;
  wire s_dadda_pg_rca24_fa63_xor1;
  wire s_dadda_pg_rca24_fa63_and1;
  wire s_dadda_pg_rca24_fa63_or0;
  wire s_dadda_pg_rca24_and_15_0;
  wire s_dadda_pg_rca24_and_14_1;
  wire s_dadda_pg_rca24_and_13_2;
  wire s_dadda_pg_rca24_fa64_xor0;
  wire s_dadda_pg_rca24_fa64_and0;
  wire s_dadda_pg_rca24_fa64_xor1;
  wire s_dadda_pg_rca24_fa64_and1;
  wire s_dadda_pg_rca24_fa64_or0;
  wire s_dadda_pg_rca24_and_12_3;
  wire s_dadda_pg_rca24_and_11_4;
  wire s_dadda_pg_rca24_and_10_5;
  wire s_dadda_pg_rca24_fa65_xor0;
  wire s_dadda_pg_rca24_fa65_and0;
  wire s_dadda_pg_rca24_fa65_xor1;
  wire s_dadda_pg_rca24_fa65_and1;
  wire s_dadda_pg_rca24_fa65_or0;
  wire s_dadda_pg_rca24_and_9_6;
  wire s_dadda_pg_rca24_and_8_7;
  wire s_dadda_pg_rca24_and_7_8;
  wire s_dadda_pg_rca24_fa66_xor0;
  wire s_dadda_pg_rca24_fa66_and0;
  wire s_dadda_pg_rca24_fa66_xor1;
  wire s_dadda_pg_rca24_fa66_and1;
  wire s_dadda_pg_rca24_fa66_or0;
  wire s_dadda_pg_rca24_and_6_9;
  wire s_dadda_pg_rca24_and_5_10;
  wire s_dadda_pg_rca24_and_4_11;
  wire s_dadda_pg_rca24_fa67_xor0;
  wire s_dadda_pg_rca24_fa67_and0;
  wire s_dadda_pg_rca24_fa67_xor1;
  wire s_dadda_pg_rca24_fa67_and1;
  wire s_dadda_pg_rca24_fa67_or0;
  wire s_dadda_pg_rca24_and_3_12;
  wire s_dadda_pg_rca24_and_2_13;
  wire s_dadda_pg_rca24_and_1_14;
  wire s_dadda_pg_rca24_fa68_xor0;
  wire s_dadda_pg_rca24_fa68_and0;
  wire s_dadda_pg_rca24_fa68_xor1;
  wire s_dadda_pg_rca24_fa68_and1;
  wire s_dadda_pg_rca24_fa68_or0;
  wire s_dadda_pg_rca24_and_0_15;
  wire s_dadda_pg_rca24_fa69_xor0;
  wire s_dadda_pg_rca24_fa69_and0;
  wire s_dadda_pg_rca24_fa69_xor1;
  wire s_dadda_pg_rca24_fa69_and1;
  wire s_dadda_pg_rca24_fa69_or0;
  wire s_dadda_pg_rca24_ha14_xor0;
  wire s_dadda_pg_rca24_ha14_and0;
  wire s_dadda_pg_rca24_fa70_xor0;
  wire s_dadda_pg_rca24_fa70_and0;
  wire s_dadda_pg_rca24_fa70_xor1;
  wire s_dadda_pg_rca24_fa70_and1;
  wire s_dadda_pg_rca24_fa70_or0;
  wire s_dadda_pg_rca24_fa71_xor0;
  wire s_dadda_pg_rca24_fa71_and0;
  wire s_dadda_pg_rca24_fa71_xor1;
  wire s_dadda_pg_rca24_fa71_and1;
  wire s_dadda_pg_rca24_fa71_or0;
  wire s_dadda_pg_rca24_fa72_xor0;
  wire s_dadda_pg_rca24_fa72_and0;
  wire s_dadda_pg_rca24_fa72_xor1;
  wire s_dadda_pg_rca24_fa72_and1;
  wire s_dadda_pg_rca24_fa72_or0;
  wire s_dadda_pg_rca24_and_16_0;
  wire s_dadda_pg_rca24_and_15_1;
  wire s_dadda_pg_rca24_fa73_xor0;
  wire s_dadda_pg_rca24_fa73_and0;
  wire s_dadda_pg_rca24_fa73_xor1;
  wire s_dadda_pg_rca24_fa73_and1;
  wire s_dadda_pg_rca24_fa73_or0;
  wire s_dadda_pg_rca24_and_14_2;
  wire s_dadda_pg_rca24_and_13_3;
  wire s_dadda_pg_rca24_and_12_4;
  wire s_dadda_pg_rca24_fa74_xor0;
  wire s_dadda_pg_rca24_fa74_and0;
  wire s_dadda_pg_rca24_fa74_xor1;
  wire s_dadda_pg_rca24_fa74_and1;
  wire s_dadda_pg_rca24_fa74_or0;
  wire s_dadda_pg_rca24_and_11_5;
  wire s_dadda_pg_rca24_and_10_6;
  wire s_dadda_pg_rca24_and_9_7;
  wire s_dadda_pg_rca24_fa75_xor0;
  wire s_dadda_pg_rca24_fa75_and0;
  wire s_dadda_pg_rca24_fa75_xor1;
  wire s_dadda_pg_rca24_fa75_and1;
  wire s_dadda_pg_rca24_fa75_or0;
  wire s_dadda_pg_rca24_and_8_8;
  wire s_dadda_pg_rca24_and_7_9;
  wire s_dadda_pg_rca24_and_6_10;
  wire s_dadda_pg_rca24_fa76_xor0;
  wire s_dadda_pg_rca24_fa76_and0;
  wire s_dadda_pg_rca24_fa76_xor1;
  wire s_dadda_pg_rca24_fa76_and1;
  wire s_dadda_pg_rca24_fa76_or0;
  wire s_dadda_pg_rca24_and_5_11;
  wire s_dadda_pg_rca24_and_4_12;
  wire s_dadda_pg_rca24_and_3_13;
  wire s_dadda_pg_rca24_fa77_xor0;
  wire s_dadda_pg_rca24_fa77_and0;
  wire s_dadda_pg_rca24_fa77_xor1;
  wire s_dadda_pg_rca24_fa77_and1;
  wire s_dadda_pg_rca24_fa77_or0;
  wire s_dadda_pg_rca24_and_2_14;
  wire s_dadda_pg_rca24_and_1_15;
  wire s_dadda_pg_rca24_and_0_16;
  wire s_dadda_pg_rca24_fa78_xor0;
  wire s_dadda_pg_rca24_fa78_and0;
  wire s_dadda_pg_rca24_fa78_xor1;
  wire s_dadda_pg_rca24_fa78_and1;
  wire s_dadda_pg_rca24_fa78_or0;
  wire s_dadda_pg_rca24_fa79_xor0;
  wire s_dadda_pg_rca24_fa79_and0;
  wire s_dadda_pg_rca24_fa79_xor1;
  wire s_dadda_pg_rca24_fa79_and1;
  wire s_dadda_pg_rca24_fa79_or0;
  wire s_dadda_pg_rca24_ha15_xor0;
  wire s_dadda_pg_rca24_ha15_and0;
  wire s_dadda_pg_rca24_fa80_xor0;
  wire s_dadda_pg_rca24_fa80_and0;
  wire s_dadda_pg_rca24_fa80_xor1;
  wire s_dadda_pg_rca24_fa80_and1;
  wire s_dadda_pg_rca24_fa80_or0;
  wire s_dadda_pg_rca24_fa81_xor0;
  wire s_dadda_pg_rca24_fa81_and0;
  wire s_dadda_pg_rca24_fa81_xor1;
  wire s_dadda_pg_rca24_fa81_and1;
  wire s_dadda_pg_rca24_fa81_or0;
  wire s_dadda_pg_rca24_fa82_xor0;
  wire s_dadda_pg_rca24_fa82_and0;
  wire s_dadda_pg_rca24_fa82_xor1;
  wire s_dadda_pg_rca24_fa82_and1;
  wire s_dadda_pg_rca24_fa82_or0;
  wire s_dadda_pg_rca24_and_17_0;
  wire s_dadda_pg_rca24_fa83_xor0;
  wire s_dadda_pg_rca24_fa83_and0;
  wire s_dadda_pg_rca24_fa83_xor1;
  wire s_dadda_pg_rca24_fa83_and1;
  wire s_dadda_pg_rca24_fa83_or0;
  wire s_dadda_pg_rca24_and_16_1;
  wire s_dadda_pg_rca24_and_15_2;
  wire s_dadda_pg_rca24_and_14_3;
  wire s_dadda_pg_rca24_fa84_xor0;
  wire s_dadda_pg_rca24_fa84_and0;
  wire s_dadda_pg_rca24_fa84_xor1;
  wire s_dadda_pg_rca24_fa84_and1;
  wire s_dadda_pg_rca24_fa84_or0;
  wire s_dadda_pg_rca24_and_13_4;
  wire s_dadda_pg_rca24_and_12_5;
  wire s_dadda_pg_rca24_and_11_6;
  wire s_dadda_pg_rca24_fa85_xor0;
  wire s_dadda_pg_rca24_fa85_and0;
  wire s_dadda_pg_rca24_fa85_xor1;
  wire s_dadda_pg_rca24_fa85_and1;
  wire s_dadda_pg_rca24_fa85_or0;
  wire s_dadda_pg_rca24_and_10_7;
  wire s_dadda_pg_rca24_and_9_8;
  wire s_dadda_pg_rca24_and_8_9;
  wire s_dadda_pg_rca24_fa86_xor0;
  wire s_dadda_pg_rca24_fa86_and0;
  wire s_dadda_pg_rca24_fa86_xor1;
  wire s_dadda_pg_rca24_fa86_and1;
  wire s_dadda_pg_rca24_fa86_or0;
  wire s_dadda_pg_rca24_and_7_10;
  wire s_dadda_pg_rca24_and_6_11;
  wire s_dadda_pg_rca24_and_5_12;
  wire s_dadda_pg_rca24_fa87_xor0;
  wire s_dadda_pg_rca24_fa87_and0;
  wire s_dadda_pg_rca24_fa87_xor1;
  wire s_dadda_pg_rca24_fa87_and1;
  wire s_dadda_pg_rca24_fa87_or0;
  wire s_dadda_pg_rca24_and_4_13;
  wire s_dadda_pg_rca24_and_3_14;
  wire s_dadda_pg_rca24_and_2_15;
  wire s_dadda_pg_rca24_fa88_xor0;
  wire s_dadda_pg_rca24_fa88_and0;
  wire s_dadda_pg_rca24_fa88_xor1;
  wire s_dadda_pg_rca24_fa88_and1;
  wire s_dadda_pg_rca24_fa88_or0;
  wire s_dadda_pg_rca24_and_1_16;
  wire s_dadda_pg_rca24_and_0_17;
  wire s_dadda_pg_rca24_fa89_xor0;
  wire s_dadda_pg_rca24_fa89_and0;
  wire s_dadda_pg_rca24_fa89_xor1;
  wire s_dadda_pg_rca24_fa89_and1;
  wire s_dadda_pg_rca24_fa89_or0;
  wire s_dadda_pg_rca24_fa90_xor0;
  wire s_dadda_pg_rca24_fa90_and0;
  wire s_dadda_pg_rca24_fa90_xor1;
  wire s_dadda_pg_rca24_fa90_and1;
  wire s_dadda_pg_rca24_fa90_or0;
  wire s_dadda_pg_rca24_ha16_xor0;
  wire s_dadda_pg_rca24_ha16_and0;
  wire s_dadda_pg_rca24_fa91_xor0;
  wire s_dadda_pg_rca24_fa91_and0;
  wire s_dadda_pg_rca24_fa91_xor1;
  wire s_dadda_pg_rca24_fa91_and1;
  wire s_dadda_pg_rca24_fa91_or0;
  wire s_dadda_pg_rca24_fa92_xor0;
  wire s_dadda_pg_rca24_fa92_and0;
  wire s_dadda_pg_rca24_fa92_xor1;
  wire s_dadda_pg_rca24_fa92_and1;
  wire s_dadda_pg_rca24_fa92_or0;
  wire s_dadda_pg_rca24_fa93_xor0;
  wire s_dadda_pg_rca24_fa93_and0;
  wire s_dadda_pg_rca24_fa93_xor1;
  wire s_dadda_pg_rca24_fa93_and1;
  wire s_dadda_pg_rca24_fa93_or0;
  wire s_dadda_pg_rca24_fa94_xor0;
  wire s_dadda_pg_rca24_fa94_and0;
  wire s_dadda_pg_rca24_fa94_xor1;
  wire s_dadda_pg_rca24_fa94_and1;
  wire s_dadda_pg_rca24_fa94_or0;
  wire s_dadda_pg_rca24_and_18_0;
  wire s_dadda_pg_rca24_and_17_1;
  wire s_dadda_pg_rca24_and_16_2;
  wire s_dadda_pg_rca24_fa95_xor0;
  wire s_dadda_pg_rca24_fa95_and0;
  wire s_dadda_pg_rca24_fa95_xor1;
  wire s_dadda_pg_rca24_fa95_and1;
  wire s_dadda_pg_rca24_fa95_or0;
  wire s_dadda_pg_rca24_and_15_3;
  wire s_dadda_pg_rca24_and_14_4;
  wire s_dadda_pg_rca24_and_13_5;
  wire s_dadda_pg_rca24_fa96_xor0;
  wire s_dadda_pg_rca24_fa96_and0;
  wire s_dadda_pg_rca24_fa96_xor1;
  wire s_dadda_pg_rca24_fa96_and1;
  wire s_dadda_pg_rca24_fa96_or0;
  wire s_dadda_pg_rca24_and_12_6;
  wire s_dadda_pg_rca24_and_11_7;
  wire s_dadda_pg_rca24_and_10_8;
  wire s_dadda_pg_rca24_fa97_xor0;
  wire s_dadda_pg_rca24_fa97_and0;
  wire s_dadda_pg_rca24_fa97_xor1;
  wire s_dadda_pg_rca24_fa97_and1;
  wire s_dadda_pg_rca24_fa97_or0;
  wire s_dadda_pg_rca24_and_9_9;
  wire s_dadda_pg_rca24_and_8_10;
  wire s_dadda_pg_rca24_and_7_11;
  wire s_dadda_pg_rca24_fa98_xor0;
  wire s_dadda_pg_rca24_fa98_and0;
  wire s_dadda_pg_rca24_fa98_xor1;
  wire s_dadda_pg_rca24_fa98_and1;
  wire s_dadda_pg_rca24_fa98_or0;
  wire s_dadda_pg_rca24_and_6_12;
  wire s_dadda_pg_rca24_and_5_13;
  wire s_dadda_pg_rca24_and_4_14;
  wire s_dadda_pg_rca24_fa99_xor0;
  wire s_dadda_pg_rca24_fa99_and0;
  wire s_dadda_pg_rca24_fa99_xor1;
  wire s_dadda_pg_rca24_fa99_and1;
  wire s_dadda_pg_rca24_fa99_or0;
  wire s_dadda_pg_rca24_and_3_15;
  wire s_dadda_pg_rca24_and_2_16;
  wire s_dadda_pg_rca24_and_1_17;
  wire s_dadda_pg_rca24_fa100_xor0;
  wire s_dadda_pg_rca24_fa100_and0;
  wire s_dadda_pg_rca24_fa100_xor1;
  wire s_dadda_pg_rca24_fa100_and1;
  wire s_dadda_pg_rca24_fa100_or0;
  wire s_dadda_pg_rca24_and_0_18;
  wire s_dadda_pg_rca24_fa101_xor0;
  wire s_dadda_pg_rca24_fa101_and0;
  wire s_dadda_pg_rca24_fa101_xor1;
  wire s_dadda_pg_rca24_fa101_and1;
  wire s_dadda_pg_rca24_fa101_or0;
  wire s_dadda_pg_rca24_fa102_xor0;
  wire s_dadda_pg_rca24_fa102_and0;
  wire s_dadda_pg_rca24_fa102_xor1;
  wire s_dadda_pg_rca24_fa102_and1;
  wire s_dadda_pg_rca24_fa102_or0;
  wire s_dadda_pg_rca24_ha17_xor0;
  wire s_dadda_pg_rca24_ha17_and0;
  wire s_dadda_pg_rca24_fa103_xor0;
  wire s_dadda_pg_rca24_fa103_and0;
  wire s_dadda_pg_rca24_fa103_xor1;
  wire s_dadda_pg_rca24_fa103_and1;
  wire s_dadda_pg_rca24_fa103_or0;
  wire s_dadda_pg_rca24_fa104_xor0;
  wire s_dadda_pg_rca24_fa104_and0;
  wire s_dadda_pg_rca24_fa104_xor1;
  wire s_dadda_pg_rca24_fa104_and1;
  wire s_dadda_pg_rca24_fa104_or0;
  wire s_dadda_pg_rca24_fa105_xor0;
  wire s_dadda_pg_rca24_fa105_and0;
  wire s_dadda_pg_rca24_fa105_xor1;
  wire s_dadda_pg_rca24_fa105_and1;
  wire s_dadda_pg_rca24_fa105_or0;
  wire s_dadda_pg_rca24_fa106_xor0;
  wire s_dadda_pg_rca24_fa106_and0;
  wire s_dadda_pg_rca24_fa106_xor1;
  wire s_dadda_pg_rca24_fa106_and1;
  wire s_dadda_pg_rca24_fa106_or0;
  wire s_dadda_pg_rca24_and_17_2;
  wire s_dadda_pg_rca24_and_16_3;
  wire s_dadda_pg_rca24_fa107_xor0;
  wire s_dadda_pg_rca24_fa107_and0;
  wire s_dadda_pg_rca24_fa107_xor1;
  wire s_dadda_pg_rca24_fa107_and1;
  wire s_dadda_pg_rca24_fa107_or0;
  wire s_dadda_pg_rca24_and_15_4;
  wire s_dadda_pg_rca24_and_14_5;
  wire s_dadda_pg_rca24_and_13_6;
  wire s_dadda_pg_rca24_fa108_xor0;
  wire s_dadda_pg_rca24_fa108_and0;
  wire s_dadda_pg_rca24_fa108_xor1;
  wire s_dadda_pg_rca24_fa108_and1;
  wire s_dadda_pg_rca24_fa108_or0;
  wire s_dadda_pg_rca24_and_12_7;
  wire s_dadda_pg_rca24_and_11_8;
  wire s_dadda_pg_rca24_and_10_9;
  wire s_dadda_pg_rca24_fa109_xor0;
  wire s_dadda_pg_rca24_fa109_and0;
  wire s_dadda_pg_rca24_fa109_xor1;
  wire s_dadda_pg_rca24_fa109_and1;
  wire s_dadda_pg_rca24_fa109_or0;
  wire s_dadda_pg_rca24_and_9_10;
  wire s_dadda_pg_rca24_and_8_11;
  wire s_dadda_pg_rca24_and_7_12;
  wire s_dadda_pg_rca24_fa110_xor0;
  wire s_dadda_pg_rca24_fa110_and0;
  wire s_dadda_pg_rca24_fa110_xor1;
  wire s_dadda_pg_rca24_fa110_and1;
  wire s_dadda_pg_rca24_fa110_or0;
  wire s_dadda_pg_rca24_and_6_13;
  wire s_dadda_pg_rca24_and_5_14;
  wire s_dadda_pg_rca24_and_4_15;
  wire s_dadda_pg_rca24_fa111_xor0;
  wire s_dadda_pg_rca24_fa111_and0;
  wire s_dadda_pg_rca24_fa111_xor1;
  wire s_dadda_pg_rca24_fa111_and1;
  wire s_dadda_pg_rca24_fa111_or0;
  wire s_dadda_pg_rca24_and_3_16;
  wire s_dadda_pg_rca24_and_2_17;
  wire s_dadda_pg_rca24_and_1_18;
  wire s_dadda_pg_rca24_fa112_xor0;
  wire s_dadda_pg_rca24_fa112_and0;
  wire s_dadda_pg_rca24_fa112_xor1;
  wire s_dadda_pg_rca24_fa112_and1;
  wire s_dadda_pg_rca24_fa112_or0;
  wire s_dadda_pg_rca24_and_0_19;
  wire s_dadda_pg_rca24_fa113_xor0;
  wire s_dadda_pg_rca24_fa113_and0;
  wire s_dadda_pg_rca24_fa113_xor1;
  wire s_dadda_pg_rca24_fa113_and1;
  wire s_dadda_pg_rca24_fa113_or0;
  wire s_dadda_pg_rca24_fa114_xor0;
  wire s_dadda_pg_rca24_fa114_and0;
  wire s_dadda_pg_rca24_fa114_xor1;
  wire s_dadda_pg_rca24_fa114_and1;
  wire s_dadda_pg_rca24_fa114_or0;
  wire s_dadda_pg_rca24_fa115_xor0;
  wire s_dadda_pg_rca24_fa115_and0;
  wire s_dadda_pg_rca24_fa115_xor1;
  wire s_dadda_pg_rca24_fa115_and1;
  wire s_dadda_pg_rca24_fa115_or0;
  wire s_dadda_pg_rca24_fa116_xor0;
  wire s_dadda_pg_rca24_fa116_and0;
  wire s_dadda_pg_rca24_fa116_xor1;
  wire s_dadda_pg_rca24_fa116_and1;
  wire s_dadda_pg_rca24_fa116_or0;
  wire s_dadda_pg_rca24_fa117_xor0;
  wire s_dadda_pg_rca24_fa117_and0;
  wire s_dadda_pg_rca24_fa117_xor1;
  wire s_dadda_pg_rca24_fa117_and1;
  wire s_dadda_pg_rca24_fa117_or0;
  wire s_dadda_pg_rca24_fa118_xor0;
  wire s_dadda_pg_rca24_fa118_and0;
  wire s_dadda_pg_rca24_fa118_xor1;
  wire s_dadda_pg_rca24_fa118_and1;
  wire s_dadda_pg_rca24_fa118_or0;
  wire s_dadda_pg_rca24_fa119_xor0;
  wire s_dadda_pg_rca24_fa119_and0;
  wire s_dadda_pg_rca24_fa119_xor1;
  wire s_dadda_pg_rca24_fa119_and1;
  wire s_dadda_pg_rca24_fa119_or0;
  wire s_dadda_pg_rca24_and_16_4;
  wire s_dadda_pg_rca24_and_15_5;
  wire s_dadda_pg_rca24_fa120_xor0;
  wire s_dadda_pg_rca24_fa120_and0;
  wire s_dadda_pg_rca24_fa120_xor1;
  wire s_dadda_pg_rca24_fa120_and1;
  wire s_dadda_pg_rca24_fa120_or0;
  wire s_dadda_pg_rca24_and_14_6;
  wire s_dadda_pg_rca24_and_13_7;
  wire s_dadda_pg_rca24_and_12_8;
  wire s_dadda_pg_rca24_fa121_xor0;
  wire s_dadda_pg_rca24_fa121_and0;
  wire s_dadda_pg_rca24_fa121_xor1;
  wire s_dadda_pg_rca24_fa121_and1;
  wire s_dadda_pg_rca24_fa121_or0;
  wire s_dadda_pg_rca24_and_11_9;
  wire s_dadda_pg_rca24_and_10_10;
  wire s_dadda_pg_rca24_and_9_11;
  wire s_dadda_pg_rca24_fa122_xor0;
  wire s_dadda_pg_rca24_fa122_and0;
  wire s_dadda_pg_rca24_fa122_xor1;
  wire s_dadda_pg_rca24_fa122_and1;
  wire s_dadda_pg_rca24_fa122_or0;
  wire s_dadda_pg_rca24_and_8_12;
  wire s_dadda_pg_rca24_and_7_13;
  wire s_dadda_pg_rca24_and_6_14;
  wire s_dadda_pg_rca24_fa123_xor0;
  wire s_dadda_pg_rca24_fa123_and0;
  wire s_dadda_pg_rca24_fa123_xor1;
  wire s_dadda_pg_rca24_fa123_and1;
  wire s_dadda_pg_rca24_fa123_or0;
  wire s_dadda_pg_rca24_and_5_15;
  wire s_dadda_pg_rca24_and_4_16;
  wire s_dadda_pg_rca24_and_3_17;
  wire s_dadda_pg_rca24_fa124_xor0;
  wire s_dadda_pg_rca24_fa124_and0;
  wire s_dadda_pg_rca24_fa124_xor1;
  wire s_dadda_pg_rca24_fa124_and1;
  wire s_dadda_pg_rca24_fa124_or0;
  wire s_dadda_pg_rca24_and_2_18;
  wire s_dadda_pg_rca24_and_1_19;
  wire s_dadda_pg_rca24_and_0_20;
  wire s_dadda_pg_rca24_fa125_xor0;
  wire s_dadda_pg_rca24_fa125_and0;
  wire s_dadda_pg_rca24_fa125_xor1;
  wire s_dadda_pg_rca24_fa125_and1;
  wire s_dadda_pg_rca24_fa125_or0;
  wire s_dadda_pg_rca24_fa126_xor0;
  wire s_dadda_pg_rca24_fa126_and0;
  wire s_dadda_pg_rca24_fa126_xor1;
  wire s_dadda_pg_rca24_fa126_and1;
  wire s_dadda_pg_rca24_fa126_or0;
  wire s_dadda_pg_rca24_fa127_xor0;
  wire s_dadda_pg_rca24_fa127_and0;
  wire s_dadda_pg_rca24_fa127_xor1;
  wire s_dadda_pg_rca24_fa127_and1;
  wire s_dadda_pg_rca24_fa127_or0;
  wire s_dadda_pg_rca24_fa128_xor0;
  wire s_dadda_pg_rca24_fa128_and0;
  wire s_dadda_pg_rca24_fa128_xor1;
  wire s_dadda_pg_rca24_fa128_and1;
  wire s_dadda_pg_rca24_fa128_or0;
  wire s_dadda_pg_rca24_fa129_xor0;
  wire s_dadda_pg_rca24_fa129_and0;
  wire s_dadda_pg_rca24_fa129_xor1;
  wire s_dadda_pg_rca24_fa129_and1;
  wire s_dadda_pg_rca24_fa129_or0;
  wire s_dadda_pg_rca24_fa130_xor0;
  wire s_dadda_pg_rca24_fa130_and0;
  wire s_dadda_pg_rca24_fa130_xor1;
  wire s_dadda_pg_rca24_fa130_and1;
  wire s_dadda_pg_rca24_fa130_or0;
  wire s_dadda_pg_rca24_fa131_xor0;
  wire s_dadda_pg_rca24_fa131_and0;
  wire s_dadda_pg_rca24_fa131_xor1;
  wire s_dadda_pg_rca24_fa131_and1;
  wire s_dadda_pg_rca24_fa131_or0;
  wire s_dadda_pg_rca24_fa132_xor0;
  wire s_dadda_pg_rca24_fa132_and0;
  wire s_dadda_pg_rca24_fa132_xor1;
  wire s_dadda_pg_rca24_fa132_and1;
  wire s_dadda_pg_rca24_fa132_or0;
  wire s_dadda_pg_rca24_and_15_6;
  wire s_dadda_pg_rca24_and_14_7;
  wire s_dadda_pg_rca24_fa133_xor0;
  wire s_dadda_pg_rca24_fa133_and0;
  wire s_dadda_pg_rca24_fa133_xor1;
  wire s_dadda_pg_rca24_fa133_and1;
  wire s_dadda_pg_rca24_fa133_or0;
  wire s_dadda_pg_rca24_and_13_8;
  wire s_dadda_pg_rca24_and_12_9;
  wire s_dadda_pg_rca24_and_11_10;
  wire s_dadda_pg_rca24_fa134_xor0;
  wire s_dadda_pg_rca24_fa134_and0;
  wire s_dadda_pg_rca24_fa134_xor1;
  wire s_dadda_pg_rca24_fa134_and1;
  wire s_dadda_pg_rca24_fa134_or0;
  wire s_dadda_pg_rca24_and_10_11;
  wire s_dadda_pg_rca24_and_9_12;
  wire s_dadda_pg_rca24_and_8_13;
  wire s_dadda_pg_rca24_fa135_xor0;
  wire s_dadda_pg_rca24_fa135_and0;
  wire s_dadda_pg_rca24_fa135_xor1;
  wire s_dadda_pg_rca24_fa135_and1;
  wire s_dadda_pg_rca24_fa135_or0;
  wire s_dadda_pg_rca24_and_7_14;
  wire s_dadda_pg_rca24_and_6_15;
  wire s_dadda_pg_rca24_and_5_16;
  wire s_dadda_pg_rca24_fa136_xor0;
  wire s_dadda_pg_rca24_fa136_and0;
  wire s_dadda_pg_rca24_fa136_xor1;
  wire s_dadda_pg_rca24_fa136_and1;
  wire s_dadda_pg_rca24_fa136_or0;
  wire s_dadda_pg_rca24_and_4_17;
  wire s_dadda_pg_rca24_and_3_18;
  wire s_dadda_pg_rca24_and_2_19;
  wire s_dadda_pg_rca24_fa137_xor0;
  wire s_dadda_pg_rca24_fa137_and0;
  wire s_dadda_pg_rca24_fa137_xor1;
  wire s_dadda_pg_rca24_fa137_and1;
  wire s_dadda_pg_rca24_fa137_or0;
  wire s_dadda_pg_rca24_and_1_20;
  wire s_dadda_pg_rca24_and_0_21;
  wire s_dadda_pg_rca24_fa138_xor0;
  wire s_dadda_pg_rca24_fa138_and0;
  wire s_dadda_pg_rca24_fa138_xor1;
  wire s_dadda_pg_rca24_fa138_and1;
  wire s_dadda_pg_rca24_fa138_or0;
  wire s_dadda_pg_rca24_fa139_xor0;
  wire s_dadda_pg_rca24_fa139_and0;
  wire s_dadda_pg_rca24_fa139_xor1;
  wire s_dadda_pg_rca24_fa139_and1;
  wire s_dadda_pg_rca24_fa139_or0;
  wire s_dadda_pg_rca24_fa140_xor0;
  wire s_dadda_pg_rca24_fa140_and0;
  wire s_dadda_pg_rca24_fa140_xor1;
  wire s_dadda_pg_rca24_fa140_and1;
  wire s_dadda_pg_rca24_fa140_or0;
  wire s_dadda_pg_rca24_fa141_xor0;
  wire s_dadda_pg_rca24_fa141_and0;
  wire s_dadda_pg_rca24_fa141_xor1;
  wire s_dadda_pg_rca24_fa141_and1;
  wire s_dadda_pg_rca24_fa141_or0;
  wire s_dadda_pg_rca24_fa142_xor0;
  wire s_dadda_pg_rca24_fa142_and0;
  wire s_dadda_pg_rca24_fa142_xor1;
  wire s_dadda_pg_rca24_fa142_and1;
  wire s_dadda_pg_rca24_fa142_or0;
  wire s_dadda_pg_rca24_fa143_xor0;
  wire s_dadda_pg_rca24_fa143_and0;
  wire s_dadda_pg_rca24_fa143_xor1;
  wire s_dadda_pg_rca24_fa143_and1;
  wire s_dadda_pg_rca24_fa143_or0;
  wire s_dadda_pg_rca24_fa144_xor0;
  wire s_dadda_pg_rca24_fa144_and0;
  wire s_dadda_pg_rca24_fa144_xor1;
  wire s_dadda_pg_rca24_fa144_and1;
  wire s_dadda_pg_rca24_fa144_or0;
  wire s_dadda_pg_rca24_fa145_xor0;
  wire s_dadda_pg_rca24_fa145_and0;
  wire s_dadda_pg_rca24_fa145_xor1;
  wire s_dadda_pg_rca24_fa145_and1;
  wire s_dadda_pg_rca24_fa145_or0;
  wire s_dadda_pg_rca24_and_14_8;
  wire s_dadda_pg_rca24_and_13_9;
  wire s_dadda_pg_rca24_fa146_xor0;
  wire s_dadda_pg_rca24_fa146_and0;
  wire s_dadda_pg_rca24_fa146_xor1;
  wire s_dadda_pg_rca24_fa146_and1;
  wire s_dadda_pg_rca24_fa146_or0;
  wire s_dadda_pg_rca24_and_12_10;
  wire s_dadda_pg_rca24_and_11_11;
  wire s_dadda_pg_rca24_and_10_12;
  wire s_dadda_pg_rca24_fa147_xor0;
  wire s_dadda_pg_rca24_fa147_and0;
  wire s_dadda_pg_rca24_fa147_xor1;
  wire s_dadda_pg_rca24_fa147_and1;
  wire s_dadda_pg_rca24_fa147_or0;
  wire s_dadda_pg_rca24_and_9_13;
  wire s_dadda_pg_rca24_and_8_14;
  wire s_dadda_pg_rca24_and_7_15;
  wire s_dadda_pg_rca24_fa148_xor0;
  wire s_dadda_pg_rca24_fa148_and0;
  wire s_dadda_pg_rca24_fa148_xor1;
  wire s_dadda_pg_rca24_fa148_and1;
  wire s_dadda_pg_rca24_fa148_or0;
  wire s_dadda_pg_rca24_and_6_16;
  wire s_dadda_pg_rca24_and_5_17;
  wire s_dadda_pg_rca24_and_4_18;
  wire s_dadda_pg_rca24_fa149_xor0;
  wire s_dadda_pg_rca24_fa149_and0;
  wire s_dadda_pg_rca24_fa149_xor1;
  wire s_dadda_pg_rca24_fa149_and1;
  wire s_dadda_pg_rca24_fa149_or0;
  wire s_dadda_pg_rca24_and_3_19;
  wire s_dadda_pg_rca24_and_2_20;
  wire s_dadda_pg_rca24_and_1_21;
  wire s_dadda_pg_rca24_fa150_xor0;
  wire s_dadda_pg_rca24_fa150_and0;
  wire s_dadda_pg_rca24_fa150_xor1;
  wire s_dadda_pg_rca24_fa150_and1;
  wire s_dadda_pg_rca24_fa150_or0;
  wire s_dadda_pg_rca24_and_0_22;
  wire s_dadda_pg_rca24_fa151_xor0;
  wire s_dadda_pg_rca24_fa151_and0;
  wire s_dadda_pg_rca24_fa151_xor1;
  wire s_dadda_pg_rca24_fa151_and1;
  wire s_dadda_pg_rca24_fa151_or0;
  wire s_dadda_pg_rca24_fa152_xor0;
  wire s_dadda_pg_rca24_fa152_and0;
  wire s_dadda_pg_rca24_fa152_xor1;
  wire s_dadda_pg_rca24_fa152_and1;
  wire s_dadda_pg_rca24_fa152_or0;
  wire s_dadda_pg_rca24_fa153_xor0;
  wire s_dadda_pg_rca24_fa153_and0;
  wire s_dadda_pg_rca24_fa153_xor1;
  wire s_dadda_pg_rca24_fa153_and1;
  wire s_dadda_pg_rca24_fa153_or0;
  wire s_dadda_pg_rca24_fa154_xor0;
  wire s_dadda_pg_rca24_fa154_and0;
  wire s_dadda_pg_rca24_fa154_xor1;
  wire s_dadda_pg_rca24_fa154_and1;
  wire s_dadda_pg_rca24_fa154_or0;
  wire s_dadda_pg_rca24_fa155_xor0;
  wire s_dadda_pg_rca24_fa155_and0;
  wire s_dadda_pg_rca24_fa155_xor1;
  wire s_dadda_pg_rca24_fa155_and1;
  wire s_dadda_pg_rca24_fa155_or0;
  wire s_dadda_pg_rca24_fa156_xor0;
  wire s_dadda_pg_rca24_fa156_and0;
  wire s_dadda_pg_rca24_fa156_xor1;
  wire s_dadda_pg_rca24_fa156_and1;
  wire s_dadda_pg_rca24_fa156_or0;
  wire s_dadda_pg_rca24_fa157_xor0;
  wire s_dadda_pg_rca24_fa157_and0;
  wire s_dadda_pg_rca24_fa157_xor1;
  wire s_dadda_pg_rca24_fa157_and1;
  wire s_dadda_pg_rca24_fa157_or0;
  wire s_dadda_pg_rca24_fa158_xor0;
  wire s_dadda_pg_rca24_fa158_and0;
  wire s_dadda_pg_rca24_fa158_xor1;
  wire s_dadda_pg_rca24_fa158_and1;
  wire s_dadda_pg_rca24_fa158_or0;
  wire s_dadda_pg_rca24_and_13_10;
  wire s_dadda_pg_rca24_and_12_11;
  wire s_dadda_pg_rca24_fa159_xor0;
  wire s_dadda_pg_rca24_fa159_and0;
  wire s_dadda_pg_rca24_fa159_xor1;
  wire s_dadda_pg_rca24_fa159_and1;
  wire s_dadda_pg_rca24_fa159_or0;
  wire s_dadda_pg_rca24_and_11_12;
  wire s_dadda_pg_rca24_and_10_13;
  wire s_dadda_pg_rca24_and_9_14;
  wire s_dadda_pg_rca24_fa160_xor0;
  wire s_dadda_pg_rca24_fa160_and0;
  wire s_dadda_pg_rca24_fa160_xor1;
  wire s_dadda_pg_rca24_fa160_and1;
  wire s_dadda_pg_rca24_fa160_or0;
  wire s_dadda_pg_rca24_and_8_15;
  wire s_dadda_pg_rca24_and_7_16;
  wire s_dadda_pg_rca24_and_6_17;
  wire s_dadda_pg_rca24_fa161_xor0;
  wire s_dadda_pg_rca24_fa161_and0;
  wire s_dadda_pg_rca24_fa161_xor1;
  wire s_dadda_pg_rca24_fa161_and1;
  wire s_dadda_pg_rca24_fa161_or0;
  wire s_dadda_pg_rca24_and_5_18;
  wire s_dadda_pg_rca24_and_4_19;
  wire s_dadda_pg_rca24_and_3_20;
  wire s_dadda_pg_rca24_fa162_xor0;
  wire s_dadda_pg_rca24_fa162_and0;
  wire s_dadda_pg_rca24_fa162_xor1;
  wire s_dadda_pg_rca24_fa162_and1;
  wire s_dadda_pg_rca24_fa162_or0;
  wire s_dadda_pg_rca24_and_2_21;
  wire s_dadda_pg_rca24_and_1_22;
  wire s_dadda_pg_rca24_nand_0_23;
  wire s_dadda_pg_rca24_fa163_xor0;
  wire s_dadda_pg_rca24_fa163_and0;
  wire s_dadda_pg_rca24_fa163_xor1;
  wire s_dadda_pg_rca24_fa163_and1;
  wire s_dadda_pg_rca24_fa163_or0;
  wire s_dadda_pg_rca24_fa164_xor0;
  wire s_dadda_pg_rca24_fa164_and0;
  wire s_dadda_pg_rca24_fa164_xor1;
  wire s_dadda_pg_rca24_fa164_and1;
  wire s_dadda_pg_rca24_fa164_or0;
  wire s_dadda_pg_rca24_fa165_xor0;
  wire s_dadda_pg_rca24_fa165_and0;
  wire s_dadda_pg_rca24_fa165_xor1;
  wire s_dadda_pg_rca24_fa165_and1;
  wire s_dadda_pg_rca24_fa165_or0;
  wire s_dadda_pg_rca24_fa166_xor0;
  wire s_dadda_pg_rca24_fa166_and0;
  wire s_dadda_pg_rca24_fa166_xor1;
  wire s_dadda_pg_rca24_fa166_and1;
  wire s_dadda_pg_rca24_fa166_or0;
  wire s_dadda_pg_rca24_fa167_xor0;
  wire s_dadda_pg_rca24_fa167_and0;
  wire s_dadda_pg_rca24_fa167_xor1;
  wire s_dadda_pg_rca24_fa167_and1;
  wire s_dadda_pg_rca24_fa167_or0;
  wire s_dadda_pg_rca24_fa168_xor0;
  wire s_dadda_pg_rca24_fa168_and0;
  wire s_dadda_pg_rca24_fa168_xor1;
  wire s_dadda_pg_rca24_fa168_and1;
  wire s_dadda_pg_rca24_fa168_or0;
  wire s_dadda_pg_rca24_fa169_xor0;
  wire s_dadda_pg_rca24_fa169_and0;
  wire s_dadda_pg_rca24_fa169_xor1;
  wire s_dadda_pg_rca24_fa169_and1;
  wire s_dadda_pg_rca24_fa169_or0;
  wire s_dadda_pg_rca24_fa170_xor0;
  wire s_dadda_pg_rca24_fa170_and0;
  wire s_dadda_pg_rca24_fa170_xor1;
  wire s_dadda_pg_rca24_fa170_and1;
  wire s_dadda_pg_rca24_fa170_or0;
  wire s_dadda_pg_rca24_fa171_xor0;
  wire s_dadda_pg_rca24_fa171_and0;
  wire s_dadda_pg_rca24_fa171_xor1;
  wire s_dadda_pg_rca24_fa171_and1;
  wire s_dadda_pg_rca24_fa171_or0;
  wire s_dadda_pg_rca24_and_14_10;
  wire s_dadda_pg_rca24_and_13_11;
  wire s_dadda_pg_rca24_fa172_xor0;
  wire s_dadda_pg_rca24_fa172_and0;
  wire s_dadda_pg_rca24_fa172_xor1;
  wire s_dadda_pg_rca24_fa172_and1;
  wire s_dadda_pg_rca24_fa172_or0;
  wire s_dadda_pg_rca24_and_12_12;
  wire s_dadda_pg_rca24_and_11_13;
  wire s_dadda_pg_rca24_and_10_14;
  wire s_dadda_pg_rca24_fa173_xor0;
  wire s_dadda_pg_rca24_fa173_and0;
  wire s_dadda_pg_rca24_fa173_xor1;
  wire s_dadda_pg_rca24_fa173_and1;
  wire s_dadda_pg_rca24_fa173_or0;
  wire s_dadda_pg_rca24_and_9_15;
  wire s_dadda_pg_rca24_and_8_16;
  wire s_dadda_pg_rca24_and_7_17;
  wire s_dadda_pg_rca24_fa174_xor0;
  wire s_dadda_pg_rca24_fa174_and0;
  wire s_dadda_pg_rca24_fa174_xor1;
  wire s_dadda_pg_rca24_fa174_and1;
  wire s_dadda_pg_rca24_fa174_or0;
  wire s_dadda_pg_rca24_and_6_18;
  wire s_dadda_pg_rca24_and_5_19;
  wire s_dadda_pg_rca24_and_4_20;
  wire s_dadda_pg_rca24_fa175_xor0;
  wire s_dadda_pg_rca24_fa175_and0;
  wire s_dadda_pg_rca24_fa175_xor1;
  wire s_dadda_pg_rca24_fa175_and1;
  wire s_dadda_pg_rca24_fa175_or0;
  wire s_dadda_pg_rca24_and_3_21;
  wire s_dadda_pg_rca24_and_2_22;
  wire s_dadda_pg_rca24_nand_1_23;
  wire s_dadda_pg_rca24_fa176_xor0;
  wire s_dadda_pg_rca24_fa176_and0;
  wire s_dadda_pg_rca24_fa176_xor1;
  wire s_dadda_pg_rca24_fa176_and1;
  wire s_dadda_pg_rca24_fa176_or0;
  wire s_dadda_pg_rca24_fa177_xor0;
  wire s_dadda_pg_rca24_fa177_and0;
  wire s_dadda_pg_rca24_fa177_xor1;
  wire s_dadda_pg_rca24_fa177_and1;
  wire s_dadda_pg_rca24_fa177_or0;
  wire s_dadda_pg_rca24_fa178_xor0;
  wire s_dadda_pg_rca24_fa178_and0;
  wire s_dadda_pg_rca24_fa178_xor1;
  wire s_dadda_pg_rca24_fa178_and1;
  wire s_dadda_pg_rca24_fa178_or0;
  wire s_dadda_pg_rca24_fa179_xor0;
  wire s_dadda_pg_rca24_fa179_and0;
  wire s_dadda_pg_rca24_fa179_xor1;
  wire s_dadda_pg_rca24_fa179_and1;
  wire s_dadda_pg_rca24_fa179_or0;
  wire s_dadda_pg_rca24_fa180_xor0;
  wire s_dadda_pg_rca24_fa180_and0;
  wire s_dadda_pg_rca24_fa180_xor1;
  wire s_dadda_pg_rca24_fa180_and1;
  wire s_dadda_pg_rca24_fa180_or0;
  wire s_dadda_pg_rca24_fa181_xor0;
  wire s_dadda_pg_rca24_fa181_and0;
  wire s_dadda_pg_rca24_fa181_xor1;
  wire s_dadda_pg_rca24_fa181_and1;
  wire s_dadda_pg_rca24_fa181_or0;
  wire s_dadda_pg_rca24_fa182_xor0;
  wire s_dadda_pg_rca24_fa182_and0;
  wire s_dadda_pg_rca24_fa182_xor1;
  wire s_dadda_pg_rca24_fa182_and1;
  wire s_dadda_pg_rca24_fa182_or0;
  wire s_dadda_pg_rca24_fa183_xor0;
  wire s_dadda_pg_rca24_fa183_and0;
  wire s_dadda_pg_rca24_fa183_xor1;
  wire s_dadda_pg_rca24_fa183_and1;
  wire s_dadda_pg_rca24_fa183_or0;
  wire s_dadda_pg_rca24_fa184_xor0;
  wire s_dadda_pg_rca24_fa184_and0;
  wire s_dadda_pg_rca24_fa184_xor1;
  wire s_dadda_pg_rca24_fa184_and1;
  wire s_dadda_pg_rca24_fa184_or0;
  wire s_dadda_pg_rca24_and_16_9;
  wire s_dadda_pg_rca24_and_15_10;
  wire s_dadda_pg_rca24_fa185_xor0;
  wire s_dadda_pg_rca24_fa185_and0;
  wire s_dadda_pg_rca24_fa185_xor1;
  wire s_dadda_pg_rca24_fa185_and1;
  wire s_dadda_pg_rca24_fa185_or0;
  wire s_dadda_pg_rca24_and_14_11;
  wire s_dadda_pg_rca24_and_13_12;
  wire s_dadda_pg_rca24_and_12_13;
  wire s_dadda_pg_rca24_fa186_xor0;
  wire s_dadda_pg_rca24_fa186_and0;
  wire s_dadda_pg_rca24_fa186_xor1;
  wire s_dadda_pg_rca24_fa186_and1;
  wire s_dadda_pg_rca24_fa186_or0;
  wire s_dadda_pg_rca24_and_11_14;
  wire s_dadda_pg_rca24_and_10_15;
  wire s_dadda_pg_rca24_and_9_16;
  wire s_dadda_pg_rca24_fa187_xor0;
  wire s_dadda_pg_rca24_fa187_and0;
  wire s_dadda_pg_rca24_fa187_xor1;
  wire s_dadda_pg_rca24_fa187_and1;
  wire s_dadda_pg_rca24_fa187_or0;
  wire s_dadda_pg_rca24_and_8_17;
  wire s_dadda_pg_rca24_and_7_18;
  wire s_dadda_pg_rca24_and_6_19;
  wire s_dadda_pg_rca24_fa188_xor0;
  wire s_dadda_pg_rca24_fa188_and0;
  wire s_dadda_pg_rca24_fa188_xor1;
  wire s_dadda_pg_rca24_fa188_and1;
  wire s_dadda_pg_rca24_fa188_or0;
  wire s_dadda_pg_rca24_and_5_20;
  wire s_dadda_pg_rca24_and_4_21;
  wire s_dadda_pg_rca24_and_3_22;
  wire s_dadda_pg_rca24_fa189_xor0;
  wire s_dadda_pg_rca24_fa189_and0;
  wire s_dadda_pg_rca24_fa189_xor1;
  wire s_dadda_pg_rca24_fa189_and1;
  wire s_dadda_pg_rca24_fa189_or0;
  wire s_dadda_pg_rca24_nand_2_23;
  wire s_dadda_pg_rca24_fa190_xor0;
  wire s_dadda_pg_rca24_fa190_and0;
  wire s_dadda_pg_rca24_fa190_xor1;
  wire s_dadda_pg_rca24_fa190_and1;
  wire s_dadda_pg_rca24_fa190_or0;
  wire s_dadda_pg_rca24_fa191_xor0;
  wire s_dadda_pg_rca24_fa191_and0;
  wire s_dadda_pg_rca24_fa191_xor1;
  wire s_dadda_pg_rca24_fa191_and1;
  wire s_dadda_pg_rca24_fa191_or0;
  wire s_dadda_pg_rca24_fa192_xor0;
  wire s_dadda_pg_rca24_fa192_and0;
  wire s_dadda_pg_rca24_fa192_xor1;
  wire s_dadda_pg_rca24_fa192_and1;
  wire s_dadda_pg_rca24_fa192_or0;
  wire s_dadda_pg_rca24_fa193_xor0;
  wire s_dadda_pg_rca24_fa193_and0;
  wire s_dadda_pg_rca24_fa193_xor1;
  wire s_dadda_pg_rca24_fa193_and1;
  wire s_dadda_pg_rca24_fa193_or0;
  wire s_dadda_pg_rca24_fa194_xor0;
  wire s_dadda_pg_rca24_fa194_and0;
  wire s_dadda_pg_rca24_fa194_xor1;
  wire s_dadda_pg_rca24_fa194_and1;
  wire s_dadda_pg_rca24_fa194_or0;
  wire s_dadda_pg_rca24_fa195_xor0;
  wire s_dadda_pg_rca24_fa195_and0;
  wire s_dadda_pg_rca24_fa195_xor1;
  wire s_dadda_pg_rca24_fa195_and1;
  wire s_dadda_pg_rca24_fa195_or0;
  wire s_dadda_pg_rca24_fa196_xor0;
  wire s_dadda_pg_rca24_fa196_and0;
  wire s_dadda_pg_rca24_fa196_xor1;
  wire s_dadda_pg_rca24_fa196_and1;
  wire s_dadda_pg_rca24_fa196_or0;
  wire s_dadda_pg_rca24_fa197_xor0;
  wire s_dadda_pg_rca24_fa197_and0;
  wire s_dadda_pg_rca24_fa197_xor1;
  wire s_dadda_pg_rca24_fa197_and1;
  wire s_dadda_pg_rca24_fa197_or0;
  wire s_dadda_pg_rca24_and_18_8;
  wire s_dadda_pg_rca24_and_17_9;
  wire s_dadda_pg_rca24_fa198_xor0;
  wire s_dadda_pg_rca24_fa198_and0;
  wire s_dadda_pg_rca24_fa198_xor1;
  wire s_dadda_pg_rca24_fa198_and1;
  wire s_dadda_pg_rca24_fa198_or0;
  wire s_dadda_pg_rca24_and_16_10;
  wire s_dadda_pg_rca24_and_15_11;
  wire s_dadda_pg_rca24_and_14_12;
  wire s_dadda_pg_rca24_fa199_xor0;
  wire s_dadda_pg_rca24_fa199_and0;
  wire s_dadda_pg_rca24_fa199_xor1;
  wire s_dadda_pg_rca24_fa199_and1;
  wire s_dadda_pg_rca24_fa199_or0;
  wire s_dadda_pg_rca24_and_13_13;
  wire s_dadda_pg_rca24_and_12_14;
  wire s_dadda_pg_rca24_and_11_15;
  wire s_dadda_pg_rca24_fa200_xor0;
  wire s_dadda_pg_rca24_fa200_and0;
  wire s_dadda_pg_rca24_fa200_xor1;
  wire s_dadda_pg_rca24_fa200_and1;
  wire s_dadda_pg_rca24_fa200_or0;
  wire s_dadda_pg_rca24_and_10_16;
  wire s_dadda_pg_rca24_and_9_17;
  wire s_dadda_pg_rca24_and_8_18;
  wire s_dadda_pg_rca24_fa201_xor0;
  wire s_dadda_pg_rca24_fa201_and0;
  wire s_dadda_pg_rca24_fa201_xor1;
  wire s_dadda_pg_rca24_fa201_and1;
  wire s_dadda_pg_rca24_fa201_or0;
  wire s_dadda_pg_rca24_and_7_19;
  wire s_dadda_pg_rca24_and_6_20;
  wire s_dadda_pg_rca24_and_5_21;
  wire s_dadda_pg_rca24_fa202_xor0;
  wire s_dadda_pg_rca24_fa202_and0;
  wire s_dadda_pg_rca24_fa202_xor1;
  wire s_dadda_pg_rca24_fa202_and1;
  wire s_dadda_pg_rca24_fa202_or0;
  wire s_dadda_pg_rca24_and_4_22;
  wire s_dadda_pg_rca24_nand_3_23;
  wire s_dadda_pg_rca24_fa203_xor0;
  wire s_dadda_pg_rca24_fa203_and0;
  wire s_dadda_pg_rca24_fa203_xor1;
  wire s_dadda_pg_rca24_fa203_and1;
  wire s_dadda_pg_rca24_fa203_or0;
  wire s_dadda_pg_rca24_fa204_xor0;
  wire s_dadda_pg_rca24_fa204_and0;
  wire s_dadda_pg_rca24_fa204_xor1;
  wire s_dadda_pg_rca24_fa204_and1;
  wire s_dadda_pg_rca24_fa204_or0;
  wire s_dadda_pg_rca24_fa205_xor0;
  wire s_dadda_pg_rca24_fa205_and0;
  wire s_dadda_pg_rca24_fa205_xor1;
  wire s_dadda_pg_rca24_fa205_and1;
  wire s_dadda_pg_rca24_fa205_or0;
  wire s_dadda_pg_rca24_fa206_xor0;
  wire s_dadda_pg_rca24_fa206_and0;
  wire s_dadda_pg_rca24_fa206_xor1;
  wire s_dadda_pg_rca24_fa206_and1;
  wire s_dadda_pg_rca24_fa206_or0;
  wire s_dadda_pg_rca24_fa207_xor0;
  wire s_dadda_pg_rca24_fa207_and0;
  wire s_dadda_pg_rca24_fa207_xor1;
  wire s_dadda_pg_rca24_fa207_and1;
  wire s_dadda_pg_rca24_fa207_or0;
  wire s_dadda_pg_rca24_fa208_xor0;
  wire s_dadda_pg_rca24_fa208_and0;
  wire s_dadda_pg_rca24_fa208_xor1;
  wire s_dadda_pg_rca24_fa208_and1;
  wire s_dadda_pg_rca24_fa208_or0;
  wire s_dadda_pg_rca24_fa209_xor0;
  wire s_dadda_pg_rca24_fa209_and0;
  wire s_dadda_pg_rca24_fa209_xor1;
  wire s_dadda_pg_rca24_fa209_and1;
  wire s_dadda_pg_rca24_fa209_or0;
  wire s_dadda_pg_rca24_fa210_xor0;
  wire s_dadda_pg_rca24_fa210_and0;
  wire s_dadda_pg_rca24_fa210_xor1;
  wire s_dadda_pg_rca24_fa210_and1;
  wire s_dadda_pg_rca24_fa210_or0;
  wire s_dadda_pg_rca24_and_20_7;
  wire s_dadda_pg_rca24_and_19_8;
  wire s_dadda_pg_rca24_fa211_xor0;
  wire s_dadda_pg_rca24_fa211_and0;
  wire s_dadda_pg_rca24_fa211_xor1;
  wire s_dadda_pg_rca24_fa211_and1;
  wire s_dadda_pg_rca24_fa211_or0;
  wire s_dadda_pg_rca24_and_18_9;
  wire s_dadda_pg_rca24_and_17_10;
  wire s_dadda_pg_rca24_and_16_11;
  wire s_dadda_pg_rca24_fa212_xor0;
  wire s_dadda_pg_rca24_fa212_and0;
  wire s_dadda_pg_rca24_fa212_xor1;
  wire s_dadda_pg_rca24_fa212_and1;
  wire s_dadda_pg_rca24_fa212_or0;
  wire s_dadda_pg_rca24_and_15_12;
  wire s_dadda_pg_rca24_and_14_13;
  wire s_dadda_pg_rca24_and_13_14;
  wire s_dadda_pg_rca24_fa213_xor0;
  wire s_dadda_pg_rca24_fa213_and0;
  wire s_dadda_pg_rca24_fa213_xor1;
  wire s_dadda_pg_rca24_fa213_and1;
  wire s_dadda_pg_rca24_fa213_or0;
  wire s_dadda_pg_rca24_and_12_15;
  wire s_dadda_pg_rca24_and_11_16;
  wire s_dadda_pg_rca24_and_10_17;
  wire s_dadda_pg_rca24_fa214_xor0;
  wire s_dadda_pg_rca24_fa214_and0;
  wire s_dadda_pg_rca24_fa214_xor1;
  wire s_dadda_pg_rca24_fa214_and1;
  wire s_dadda_pg_rca24_fa214_or0;
  wire s_dadda_pg_rca24_and_9_18;
  wire s_dadda_pg_rca24_and_8_19;
  wire s_dadda_pg_rca24_and_7_20;
  wire s_dadda_pg_rca24_fa215_xor0;
  wire s_dadda_pg_rca24_fa215_and0;
  wire s_dadda_pg_rca24_fa215_xor1;
  wire s_dadda_pg_rca24_fa215_and1;
  wire s_dadda_pg_rca24_fa215_or0;
  wire s_dadda_pg_rca24_and_6_21;
  wire s_dadda_pg_rca24_and_5_22;
  wire s_dadda_pg_rca24_nand_4_23;
  wire s_dadda_pg_rca24_fa216_xor0;
  wire s_dadda_pg_rca24_fa216_and0;
  wire s_dadda_pg_rca24_fa216_xor1;
  wire s_dadda_pg_rca24_fa216_and1;
  wire s_dadda_pg_rca24_fa216_or0;
  wire s_dadda_pg_rca24_fa217_xor0;
  wire s_dadda_pg_rca24_fa217_and0;
  wire s_dadda_pg_rca24_fa217_xor1;
  wire s_dadda_pg_rca24_fa217_and1;
  wire s_dadda_pg_rca24_fa217_or0;
  wire s_dadda_pg_rca24_fa218_xor0;
  wire s_dadda_pg_rca24_fa218_and0;
  wire s_dadda_pg_rca24_fa218_xor1;
  wire s_dadda_pg_rca24_fa218_and1;
  wire s_dadda_pg_rca24_fa218_or0;
  wire s_dadda_pg_rca24_fa219_xor0;
  wire s_dadda_pg_rca24_fa219_and0;
  wire s_dadda_pg_rca24_fa219_xor1;
  wire s_dadda_pg_rca24_fa219_and1;
  wire s_dadda_pg_rca24_fa219_or0;
  wire s_dadda_pg_rca24_fa220_xor0;
  wire s_dadda_pg_rca24_fa220_and0;
  wire s_dadda_pg_rca24_fa220_xor1;
  wire s_dadda_pg_rca24_fa220_and1;
  wire s_dadda_pg_rca24_fa220_or0;
  wire s_dadda_pg_rca24_fa221_xor0;
  wire s_dadda_pg_rca24_fa221_and0;
  wire s_dadda_pg_rca24_fa221_xor1;
  wire s_dadda_pg_rca24_fa221_and1;
  wire s_dadda_pg_rca24_fa221_or0;
  wire s_dadda_pg_rca24_fa222_xor0;
  wire s_dadda_pg_rca24_fa222_and0;
  wire s_dadda_pg_rca24_fa222_xor1;
  wire s_dadda_pg_rca24_fa222_and1;
  wire s_dadda_pg_rca24_fa222_or0;
  wire s_dadda_pg_rca24_fa223_xor0;
  wire s_dadda_pg_rca24_fa223_and0;
  wire s_dadda_pg_rca24_fa223_xor1;
  wire s_dadda_pg_rca24_fa223_and1;
  wire s_dadda_pg_rca24_fa223_or0;
  wire s_dadda_pg_rca24_and_22_6;
  wire s_dadda_pg_rca24_and_21_7;
  wire s_dadda_pg_rca24_fa224_xor0;
  wire s_dadda_pg_rca24_fa224_and0;
  wire s_dadda_pg_rca24_fa224_xor1;
  wire s_dadda_pg_rca24_fa224_and1;
  wire s_dadda_pg_rca24_fa224_or0;
  wire s_dadda_pg_rca24_and_20_8;
  wire s_dadda_pg_rca24_and_19_9;
  wire s_dadda_pg_rca24_and_18_10;
  wire s_dadda_pg_rca24_fa225_xor0;
  wire s_dadda_pg_rca24_fa225_and0;
  wire s_dadda_pg_rca24_fa225_xor1;
  wire s_dadda_pg_rca24_fa225_and1;
  wire s_dadda_pg_rca24_fa225_or0;
  wire s_dadda_pg_rca24_and_17_11;
  wire s_dadda_pg_rca24_and_16_12;
  wire s_dadda_pg_rca24_and_15_13;
  wire s_dadda_pg_rca24_fa226_xor0;
  wire s_dadda_pg_rca24_fa226_and0;
  wire s_dadda_pg_rca24_fa226_xor1;
  wire s_dadda_pg_rca24_fa226_and1;
  wire s_dadda_pg_rca24_fa226_or0;
  wire s_dadda_pg_rca24_and_14_14;
  wire s_dadda_pg_rca24_and_13_15;
  wire s_dadda_pg_rca24_and_12_16;
  wire s_dadda_pg_rca24_fa227_xor0;
  wire s_dadda_pg_rca24_fa227_and0;
  wire s_dadda_pg_rca24_fa227_xor1;
  wire s_dadda_pg_rca24_fa227_and1;
  wire s_dadda_pg_rca24_fa227_or0;
  wire s_dadda_pg_rca24_and_11_17;
  wire s_dadda_pg_rca24_and_10_18;
  wire s_dadda_pg_rca24_and_9_19;
  wire s_dadda_pg_rca24_fa228_xor0;
  wire s_dadda_pg_rca24_fa228_and0;
  wire s_dadda_pg_rca24_fa228_xor1;
  wire s_dadda_pg_rca24_fa228_and1;
  wire s_dadda_pg_rca24_fa228_or0;
  wire s_dadda_pg_rca24_and_8_20;
  wire s_dadda_pg_rca24_and_7_21;
  wire s_dadda_pg_rca24_and_6_22;
  wire s_dadda_pg_rca24_fa229_xor0;
  wire s_dadda_pg_rca24_fa229_and0;
  wire s_dadda_pg_rca24_fa229_xor1;
  wire s_dadda_pg_rca24_fa229_and1;
  wire s_dadda_pg_rca24_fa229_or0;
  wire s_dadda_pg_rca24_nand_5_23;
  wire s_dadda_pg_rca24_fa230_xor0;
  wire s_dadda_pg_rca24_fa230_and0;
  wire s_dadda_pg_rca24_fa230_xor1;
  wire s_dadda_pg_rca24_fa230_and1;
  wire s_dadda_pg_rca24_fa230_or0;
  wire s_dadda_pg_rca24_fa231_xor0;
  wire s_dadda_pg_rca24_fa231_and0;
  wire s_dadda_pg_rca24_fa231_xor1;
  wire s_dadda_pg_rca24_fa231_and1;
  wire s_dadda_pg_rca24_fa231_or0;
  wire s_dadda_pg_rca24_fa232_xor0;
  wire s_dadda_pg_rca24_fa232_and0;
  wire s_dadda_pg_rca24_fa232_xor1;
  wire s_dadda_pg_rca24_fa232_and1;
  wire s_dadda_pg_rca24_fa232_or0;
  wire s_dadda_pg_rca24_fa233_xor0;
  wire s_dadda_pg_rca24_fa233_and0;
  wire s_dadda_pg_rca24_fa233_xor1;
  wire s_dadda_pg_rca24_fa233_and1;
  wire s_dadda_pg_rca24_fa233_or0;
  wire s_dadda_pg_rca24_fa234_xor0;
  wire s_dadda_pg_rca24_fa234_and0;
  wire s_dadda_pg_rca24_fa234_xor1;
  wire s_dadda_pg_rca24_fa234_and1;
  wire s_dadda_pg_rca24_fa234_or0;
  wire s_dadda_pg_rca24_fa235_xor0;
  wire s_dadda_pg_rca24_fa235_and0;
  wire s_dadda_pg_rca24_fa235_xor1;
  wire s_dadda_pg_rca24_fa235_and1;
  wire s_dadda_pg_rca24_fa235_or0;
  wire s_dadda_pg_rca24_fa236_xor0;
  wire s_dadda_pg_rca24_fa236_and0;
  wire s_dadda_pg_rca24_fa236_xor1;
  wire s_dadda_pg_rca24_fa236_and1;
  wire s_dadda_pg_rca24_fa236_or0;
  wire s_dadda_pg_rca24_nand_23_6;
  wire s_dadda_pg_rca24_fa237_xor0;
  wire s_dadda_pg_rca24_fa237_and0;
  wire s_dadda_pg_rca24_fa237_xor1;
  wire s_dadda_pg_rca24_fa237_and1;
  wire s_dadda_pg_rca24_fa237_or0;
  wire s_dadda_pg_rca24_and_22_7;
  wire s_dadda_pg_rca24_and_21_8;
  wire s_dadda_pg_rca24_and_20_9;
  wire s_dadda_pg_rca24_fa238_xor0;
  wire s_dadda_pg_rca24_fa238_and0;
  wire s_dadda_pg_rca24_fa238_xor1;
  wire s_dadda_pg_rca24_fa238_and1;
  wire s_dadda_pg_rca24_fa238_or0;
  wire s_dadda_pg_rca24_and_19_10;
  wire s_dadda_pg_rca24_and_18_11;
  wire s_dadda_pg_rca24_and_17_12;
  wire s_dadda_pg_rca24_fa239_xor0;
  wire s_dadda_pg_rca24_fa239_and0;
  wire s_dadda_pg_rca24_fa239_xor1;
  wire s_dadda_pg_rca24_fa239_and1;
  wire s_dadda_pg_rca24_fa239_or0;
  wire s_dadda_pg_rca24_and_16_13;
  wire s_dadda_pg_rca24_and_15_14;
  wire s_dadda_pg_rca24_and_14_15;
  wire s_dadda_pg_rca24_fa240_xor0;
  wire s_dadda_pg_rca24_fa240_and0;
  wire s_dadda_pg_rca24_fa240_xor1;
  wire s_dadda_pg_rca24_fa240_and1;
  wire s_dadda_pg_rca24_fa240_or0;
  wire s_dadda_pg_rca24_and_13_16;
  wire s_dadda_pg_rca24_and_12_17;
  wire s_dadda_pg_rca24_and_11_18;
  wire s_dadda_pg_rca24_fa241_xor0;
  wire s_dadda_pg_rca24_fa241_and0;
  wire s_dadda_pg_rca24_fa241_xor1;
  wire s_dadda_pg_rca24_fa241_and1;
  wire s_dadda_pg_rca24_fa241_or0;
  wire s_dadda_pg_rca24_and_10_19;
  wire s_dadda_pg_rca24_and_9_20;
  wire s_dadda_pg_rca24_and_8_21;
  wire s_dadda_pg_rca24_fa242_xor0;
  wire s_dadda_pg_rca24_fa242_and0;
  wire s_dadda_pg_rca24_fa242_xor1;
  wire s_dadda_pg_rca24_fa242_and1;
  wire s_dadda_pg_rca24_fa242_or0;
  wire s_dadda_pg_rca24_and_7_22;
  wire s_dadda_pg_rca24_nand_6_23;
  wire s_dadda_pg_rca24_fa243_xor0;
  wire s_dadda_pg_rca24_fa243_and0;
  wire s_dadda_pg_rca24_fa243_xor1;
  wire s_dadda_pg_rca24_fa243_and1;
  wire s_dadda_pg_rca24_fa243_or0;
  wire s_dadda_pg_rca24_fa244_xor0;
  wire s_dadda_pg_rca24_fa244_and0;
  wire s_dadda_pg_rca24_fa244_xor1;
  wire s_dadda_pg_rca24_fa244_and1;
  wire s_dadda_pg_rca24_fa244_or0;
  wire s_dadda_pg_rca24_fa245_xor0;
  wire s_dadda_pg_rca24_fa245_and0;
  wire s_dadda_pg_rca24_fa245_xor1;
  wire s_dadda_pg_rca24_fa245_and1;
  wire s_dadda_pg_rca24_fa245_or0;
  wire s_dadda_pg_rca24_fa246_xor0;
  wire s_dadda_pg_rca24_fa246_and0;
  wire s_dadda_pg_rca24_fa246_xor1;
  wire s_dadda_pg_rca24_fa246_and1;
  wire s_dadda_pg_rca24_fa246_or0;
  wire s_dadda_pg_rca24_fa247_xor0;
  wire s_dadda_pg_rca24_fa247_and0;
  wire s_dadda_pg_rca24_fa247_xor1;
  wire s_dadda_pg_rca24_fa247_and1;
  wire s_dadda_pg_rca24_fa247_or0;
  wire s_dadda_pg_rca24_fa248_xor0;
  wire s_dadda_pg_rca24_fa248_and0;
  wire s_dadda_pg_rca24_fa248_xor1;
  wire s_dadda_pg_rca24_fa248_and1;
  wire s_dadda_pg_rca24_fa248_or0;
  wire s_dadda_pg_rca24_fa249_xor0;
  wire s_dadda_pg_rca24_fa249_and0;
  wire s_dadda_pg_rca24_fa249_xor1;
  wire s_dadda_pg_rca24_fa249_and1;
  wire s_dadda_pg_rca24_fa249_or0;
  wire s_dadda_pg_rca24_nand_23_7;
  wire s_dadda_pg_rca24_and_22_8;
  wire s_dadda_pg_rca24_fa250_xor0;
  wire s_dadda_pg_rca24_fa250_and0;
  wire s_dadda_pg_rca24_fa250_xor1;
  wire s_dadda_pg_rca24_fa250_and1;
  wire s_dadda_pg_rca24_fa250_or0;
  wire s_dadda_pg_rca24_and_21_9;
  wire s_dadda_pg_rca24_and_20_10;
  wire s_dadda_pg_rca24_and_19_11;
  wire s_dadda_pg_rca24_fa251_xor0;
  wire s_dadda_pg_rca24_fa251_and0;
  wire s_dadda_pg_rca24_fa251_xor1;
  wire s_dadda_pg_rca24_fa251_and1;
  wire s_dadda_pg_rca24_fa251_or0;
  wire s_dadda_pg_rca24_and_18_12;
  wire s_dadda_pg_rca24_and_17_13;
  wire s_dadda_pg_rca24_and_16_14;
  wire s_dadda_pg_rca24_fa252_xor0;
  wire s_dadda_pg_rca24_fa252_and0;
  wire s_dadda_pg_rca24_fa252_xor1;
  wire s_dadda_pg_rca24_fa252_and1;
  wire s_dadda_pg_rca24_fa252_or0;
  wire s_dadda_pg_rca24_and_15_15;
  wire s_dadda_pg_rca24_and_14_16;
  wire s_dadda_pg_rca24_and_13_17;
  wire s_dadda_pg_rca24_fa253_xor0;
  wire s_dadda_pg_rca24_fa253_and0;
  wire s_dadda_pg_rca24_fa253_xor1;
  wire s_dadda_pg_rca24_fa253_and1;
  wire s_dadda_pg_rca24_fa253_or0;
  wire s_dadda_pg_rca24_and_12_18;
  wire s_dadda_pg_rca24_and_11_19;
  wire s_dadda_pg_rca24_and_10_20;
  wire s_dadda_pg_rca24_fa254_xor0;
  wire s_dadda_pg_rca24_fa254_and0;
  wire s_dadda_pg_rca24_fa254_xor1;
  wire s_dadda_pg_rca24_fa254_and1;
  wire s_dadda_pg_rca24_fa254_or0;
  wire s_dadda_pg_rca24_and_9_21;
  wire s_dadda_pg_rca24_and_8_22;
  wire s_dadda_pg_rca24_nand_7_23;
  wire s_dadda_pg_rca24_fa255_xor0;
  wire s_dadda_pg_rca24_fa255_and0;
  wire s_dadda_pg_rca24_fa255_xor1;
  wire s_dadda_pg_rca24_fa255_and1;
  wire s_dadda_pg_rca24_fa255_or0;
  wire s_dadda_pg_rca24_fa256_xor0;
  wire s_dadda_pg_rca24_fa256_and0;
  wire s_dadda_pg_rca24_fa256_xor1;
  wire s_dadda_pg_rca24_fa256_and1;
  wire s_dadda_pg_rca24_fa256_or0;
  wire s_dadda_pg_rca24_fa257_xor0;
  wire s_dadda_pg_rca24_fa257_and0;
  wire s_dadda_pg_rca24_fa257_xor1;
  wire s_dadda_pg_rca24_fa257_and1;
  wire s_dadda_pg_rca24_fa257_or0;
  wire s_dadda_pg_rca24_fa258_xor0;
  wire s_dadda_pg_rca24_fa258_and0;
  wire s_dadda_pg_rca24_fa258_xor1;
  wire s_dadda_pg_rca24_fa258_and1;
  wire s_dadda_pg_rca24_fa258_or0;
  wire s_dadda_pg_rca24_fa259_xor0;
  wire s_dadda_pg_rca24_fa259_and0;
  wire s_dadda_pg_rca24_fa259_xor1;
  wire s_dadda_pg_rca24_fa259_and1;
  wire s_dadda_pg_rca24_fa259_or0;
  wire s_dadda_pg_rca24_fa260_xor0;
  wire s_dadda_pg_rca24_fa260_and0;
  wire s_dadda_pg_rca24_fa260_xor1;
  wire s_dadda_pg_rca24_fa260_and1;
  wire s_dadda_pg_rca24_fa260_or0;
  wire s_dadda_pg_rca24_fa261_xor0;
  wire s_dadda_pg_rca24_fa261_and0;
  wire s_dadda_pg_rca24_fa261_xor1;
  wire s_dadda_pg_rca24_fa261_and1;
  wire s_dadda_pg_rca24_fa261_or0;
  wire s_dadda_pg_rca24_nand_23_8;
  wire s_dadda_pg_rca24_and_22_9;
  wire s_dadda_pg_rca24_and_21_10;
  wire s_dadda_pg_rca24_fa262_xor0;
  wire s_dadda_pg_rca24_fa262_and0;
  wire s_dadda_pg_rca24_fa262_xor1;
  wire s_dadda_pg_rca24_fa262_and1;
  wire s_dadda_pg_rca24_fa262_or0;
  wire s_dadda_pg_rca24_and_20_11;
  wire s_dadda_pg_rca24_and_19_12;
  wire s_dadda_pg_rca24_and_18_13;
  wire s_dadda_pg_rca24_fa263_xor0;
  wire s_dadda_pg_rca24_fa263_and0;
  wire s_dadda_pg_rca24_fa263_xor1;
  wire s_dadda_pg_rca24_fa263_and1;
  wire s_dadda_pg_rca24_fa263_or0;
  wire s_dadda_pg_rca24_and_17_14;
  wire s_dadda_pg_rca24_and_16_15;
  wire s_dadda_pg_rca24_and_15_16;
  wire s_dadda_pg_rca24_fa264_xor0;
  wire s_dadda_pg_rca24_fa264_and0;
  wire s_dadda_pg_rca24_fa264_xor1;
  wire s_dadda_pg_rca24_fa264_and1;
  wire s_dadda_pg_rca24_fa264_or0;
  wire s_dadda_pg_rca24_and_14_17;
  wire s_dadda_pg_rca24_and_13_18;
  wire s_dadda_pg_rca24_and_12_19;
  wire s_dadda_pg_rca24_fa265_xor0;
  wire s_dadda_pg_rca24_fa265_and0;
  wire s_dadda_pg_rca24_fa265_xor1;
  wire s_dadda_pg_rca24_fa265_and1;
  wire s_dadda_pg_rca24_fa265_or0;
  wire s_dadda_pg_rca24_and_11_20;
  wire s_dadda_pg_rca24_and_10_21;
  wire s_dadda_pg_rca24_and_9_22;
  wire s_dadda_pg_rca24_fa266_xor0;
  wire s_dadda_pg_rca24_fa266_and0;
  wire s_dadda_pg_rca24_fa266_xor1;
  wire s_dadda_pg_rca24_fa266_and1;
  wire s_dadda_pg_rca24_fa266_or0;
  wire s_dadda_pg_rca24_nand_8_23;
  wire s_dadda_pg_rca24_fa267_xor0;
  wire s_dadda_pg_rca24_fa267_and0;
  wire s_dadda_pg_rca24_fa267_xor1;
  wire s_dadda_pg_rca24_fa267_and1;
  wire s_dadda_pg_rca24_fa267_or0;
  wire s_dadda_pg_rca24_fa268_xor0;
  wire s_dadda_pg_rca24_fa268_and0;
  wire s_dadda_pg_rca24_fa268_xor1;
  wire s_dadda_pg_rca24_fa268_and1;
  wire s_dadda_pg_rca24_fa268_or0;
  wire s_dadda_pg_rca24_fa269_xor0;
  wire s_dadda_pg_rca24_fa269_and0;
  wire s_dadda_pg_rca24_fa269_xor1;
  wire s_dadda_pg_rca24_fa269_and1;
  wire s_dadda_pg_rca24_fa269_or0;
  wire s_dadda_pg_rca24_fa270_xor0;
  wire s_dadda_pg_rca24_fa270_and0;
  wire s_dadda_pg_rca24_fa270_xor1;
  wire s_dadda_pg_rca24_fa270_and1;
  wire s_dadda_pg_rca24_fa270_or0;
  wire s_dadda_pg_rca24_fa271_xor0;
  wire s_dadda_pg_rca24_fa271_and0;
  wire s_dadda_pg_rca24_fa271_xor1;
  wire s_dadda_pg_rca24_fa271_and1;
  wire s_dadda_pg_rca24_fa271_or0;
  wire s_dadda_pg_rca24_nand_23_9;
  wire s_dadda_pg_rca24_fa272_xor0;
  wire s_dadda_pg_rca24_fa272_and0;
  wire s_dadda_pg_rca24_fa272_xor1;
  wire s_dadda_pg_rca24_fa272_and1;
  wire s_dadda_pg_rca24_fa272_or0;
  wire s_dadda_pg_rca24_and_22_10;
  wire s_dadda_pg_rca24_and_21_11;
  wire s_dadda_pg_rca24_and_20_12;
  wire s_dadda_pg_rca24_fa273_xor0;
  wire s_dadda_pg_rca24_fa273_and0;
  wire s_dadda_pg_rca24_fa273_xor1;
  wire s_dadda_pg_rca24_fa273_and1;
  wire s_dadda_pg_rca24_fa273_or0;
  wire s_dadda_pg_rca24_and_19_13;
  wire s_dadda_pg_rca24_and_18_14;
  wire s_dadda_pg_rca24_and_17_15;
  wire s_dadda_pg_rca24_fa274_xor0;
  wire s_dadda_pg_rca24_fa274_and0;
  wire s_dadda_pg_rca24_fa274_xor1;
  wire s_dadda_pg_rca24_fa274_and1;
  wire s_dadda_pg_rca24_fa274_or0;
  wire s_dadda_pg_rca24_and_16_16;
  wire s_dadda_pg_rca24_and_15_17;
  wire s_dadda_pg_rca24_and_14_18;
  wire s_dadda_pg_rca24_fa275_xor0;
  wire s_dadda_pg_rca24_fa275_and0;
  wire s_dadda_pg_rca24_fa275_xor1;
  wire s_dadda_pg_rca24_fa275_and1;
  wire s_dadda_pg_rca24_fa275_or0;
  wire s_dadda_pg_rca24_and_13_19;
  wire s_dadda_pg_rca24_and_12_20;
  wire s_dadda_pg_rca24_and_11_21;
  wire s_dadda_pg_rca24_fa276_xor0;
  wire s_dadda_pg_rca24_fa276_and0;
  wire s_dadda_pg_rca24_fa276_xor1;
  wire s_dadda_pg_rca24_fa276_and1;
  wire s_dadda_pg_rca24_fa276_or0;
  wire s_dadda_pg_rca24_and_10_22;
  wire s_dadda_pg_rca24_nand_9_23;
  wire s_dadda_pg_rca24_fa277_xor0;
  wire s_dadda_pg_rca24_fa277_and0;
  wire s_dadda_pg_rca24_fa277_xor1;
  wire s_dadda_pg_rca24_fa277_and1;
  wire s_dadda_pg_rca24_fa277_or0;
  wire s_dadda_pg_rca24_fa278_xor0;
  wire s_dadda_pg_rca24_fa278_and0;
  wire s_dadda_pg_rca24_fa278_xor1;
  wire s_dadda_pg_rca24_fa278_and1;
  wire s_dadda_pg_rca24_fa278_or0;
  wire s_dadda_pg_rca24_fa279_xor0;
  wire s_dadda_pg_rca24_fa279_and0;
  wire s_dadda_pg_rca24_fa279_xor1;
  wire s_dadda_pg_rca24_fa279_and1;
  wire s_dadda_pg_rca24_fa279_or0;
  wire s_dadda_pg_rca24_fa280_xor0;
  wire s_dadda_pg_rca24_fa280_and0;
  wire s_dadda_pg_rca24_fa280_xor1;
  wire s_dadda_pg_rca24_fa280_and1;
  wire s_dadda_pg_rca24_fa280_or0;
  wire s_dadda_pg_rca24_fa281_xor0;
  wire s_dadda_pg_rca24_fa281_and0;
  wire s_dadda_pg_rca24_fa281_xor1;
  wire s_dadda_pg_rca24_fa281_and1;
  wire s_dadda_pg_rca24_fa281_or0;
  wire s_dadda_pg_rca24_nand_23_10;
  wire s_dadda_pg_rca24_and_22_11;
  wire s_dadda_pg_rca24_fa282_xor0;
  wire s_dadda_pg_rca24_fa282_and0;
  wire s_dadda_pg_rca24_fa282_xor1;
  wire s_dadda_pg_rca24_fa282_and1;
  wire s_dadda_pg_rca24_fa282_or0;
  wire s_dadda_pg_rca24_and_21_12;
  wire s_dadda_pg_rca24_and_20_13;
  wire s_dadda_pg_rca24_and_19_14;
  wire s_dadda_pg_rca24_fa283_xor0;
  wire s_dadda_pg_rca24_fa283_and0;
  wire s_dadda_pg_rca24_fa283_xor1;
  wire s_dadda_pg_rca24_fa283_and1;
  wire s_dadda_pg_rca24_fa283_or0;
  wire s_dadda_pg_rca24_and_18_15;
  wire s_dadda_pg_rca24_and_17_16;
  wire s_dadda_pg_rca24_and_16_17;
  wire s_dadda_pg_rca24_fa284_xor0;
  wire s_dadda_pg_rca24_fa284_and0;
  wire s_dadda_pg_rca24_fa284_xor1;
  wire s_dadda_pg_rca24_fa284_and1;
  wire s_dadda_pg_rca24_fa284_or0;
  wire s_dadda_pg_rca24_and_15_18;
  wire s_dadda_pg_rca24_and_14_19;
  wire s_dadda_pg_rca24_and_13_20;
  wire s_dadda_pg_rca24_fa285_xor0;
  wire s_dadda_pg_rca24_fa285_and0;
  wire s_dadda_pg_rca24_fa285_xor1;
  wire s_dadda_pg_rca24_fa285_and1;
  wire s_dadda_pg_rca24_fa285_or0;
  wire s_dadda_pg_rca24_and_12_21;
  wire s_dadda_pg_rca24_and_11_22;
  wire s_dadda_pg_rca24_nand_10_23;
  wire s_dadda_pg_rca24_fa286_xor0;
  wire s_dadda_pg_rca24_fa286_and0;
  wire s_dadda_pg_rca24_fa286_xor1;
  wire s_dadda_pg_rca24_fa286_and1;
  wire s_dadda_pg_rca24_fa286_or0;
  wire s_dadda_pg_rca24_fa287_xor0;
  wire s_dadda_pg_rca24_fa287_and0;
  wire s_dadda_pg_rca24_fa287_xor1;
  wire s_dadda_pg_rca24_fa287_and1;
  wire s_dadda_pg_rca24_fa287_or0;
  wire s_dadda_pg_rca24_fa288_xor0;
  wire s_dadda_pg_rca24_fa288_and0;
  wire s_dadda_pg_rca24_fa288_xor1;
  wire s_dadda_pg_rca24_fa288_and1;
  wire s_dadda_pg_rca24_fa288_or0;
  wire s_dadda_pg_rca24_fa289_xor0;
  wire s_dadda_pg_rca24_fa289_and0;
  wire s_dadda_pg_rca24_fa289_xor1;
  wire s_dadda_pg_rca24_fa289_and1;
  wire s_dadda_pg_rca24_fa289_or0;
  wire s_dadda_pg_rca24_fa290_xor0;
  wire s_dadda_pg_rca24_fa290_and0;
  wire s_dadda_pg_rca24_fa290_xor1;
  wire s_dadda_pg_rca24_fa290_and1;
  wire s_dadda_pg_rca24_fa290_or0;
  wire s_dadda_pg_rca24_nand_23_11;
  wire s_dadda_pg_rca24_and_22_12;
  wire s_dadda_pg_rca24_and_21_13;
  wire s_dadda_pg_rca24_fa291_xor0;
  wire s_dadda_pg_rca24_fa291_and0;
  wire s_dadda_pg_rca24_fa291_xor1;
  wire s_dadda_pg_rca24_fa291_and1;
  wire s_dadda_pg_rca24_fa291_or0;
  wire s_dadda_pg_rca24_and_20_14;
  wire s_dadda_pg_rca24_and_19_15;
  wire s_dadda_pg_rca24_and_18_16;
  wire s_dadda_pg_rca24_fa292_xor0;
  wire s_dadda_pg_rca24_fa292_and0;
  wire s_dadda_pg_rca24_fa292_xor1;
  wire s_dadda_pg_rca24_fa292_and1;
  wire s_dadda_pg_rca24_fa292_or0;
  wire s_dadda_pg_rca24_and_17_17;
  wire s_dadda_pg_rca24_and_16_18;
  wire s_dadda_pg_rca24_and_15_19;
  wire s_dadda_pg_rca24_fa293_xor0;
  wire s_dadda_pg_rca24_fa293_and0;
  wire s_dadda_pg_rca24_fa293_xor1;
  wire s_dadda_pg_rca24_fa293_and1;
  wire s_dadda_pg_rca24_fa293_or0;
  wire s_dadda_pg_rca24_and_14_20;
  wire s_dadda_pg_rca24_and_13_21;
  wire s_dadda_pg_rca24_and_12_22;
  wire s_dadda_pg_rca24_fa294_xor0;
  wire s_dadda_pg_rca24_fa294_and0;
  wire s_dadda_pg_rca24_fa294_xor1;
  wire s_dadda_pg_rca24_fa294_and1;
  wire s_dadda_pg_rca24_fa294_or0;
  wire s_dadda_pg_rca24_nand_11_23;
  wire s_dadda_pg_rca24_fa295_xor0;
  wire s_dadda_pg_rca24_fa295_and0;
  wire s_dadda_pg_rca24_fa295_xor1;
  wire s_dadda_pg_rca24_fa295_and1;
  wire s_dadda_pg_rca24_fa295_or0;
  wire s_dadda_pg_rca24_fa296_xor0;
  wire s_dadda_pg_rca24_fa296_and0;
  wire s_dadda_pg_rca24_fa296_xor1;
  wire s_dadda_pg_rca24_fa296_and1;
  wire s_dadda_pg_rca24_fa296_or0;
  wire s_dadda_pg_rca24_fa297_xor0;
  wire s_dadda_pg_rca24_fa297_and0;
  wire s_dadda_pg_rca24_fa297_xor1;
  wire s_dadda_pg_rca24_fa297_and1;
  wire s_dadda_pg_rca24_fa297_or0;
  wire s_dadda_pg_rca24_nand_23_12;
  wire s_dadda_pg_rca24_fa298_xor0;
  wire s_dadda_pg_rca24_fa298_and0;
  wire s_dadda_pg_rca24_fa298_xor1;
  wire s_dadda_pg_rca24_fa298_and1;
  wire s_dadda_pg_rca24_fa298_or0;
  wire s_dadda_pg_rca24_and_22_13;
  wire s_dadda_pg_rca24_and_21_14;
  wire s_dadda_pg_rca24_and_20_15;
  wire s_dadda_pg_rca24_fa299_xor0;
  wire s_dadda_pg_rca24_fa299_and0;
  wire s_dadda_pg_rca24_fa299_xor1;
  wire s_dadda_pg_rca24_fa299_and1;
  wire s_dadda_pg_rca24_fa299_or0;
  wire s_dadda_pg_rca24_and_19_16;
  wire s_dadda_pg_rca24_and_18_17;
  wire s_dadda_pg_rca24_and_17_18;
  wire s_dadda_pg_rca24_fa300_xor0;
  wire s_dadda_pg_rca24_fa300_and0;
  wire s_dadda_pg_rca24_fa300_xor1;
  wire s_dadda_pg_rca24_fa300_and1;
  wire s_dadda_pg_rca24_fa300_or0;
  wire s_dadda_pg_rca24_and_16_19;
  wire s_dadda_pg_rca24_and_15_20;
  wire s_dadda_pg_rca24_and_14_21;
  wire s_dadda_pg_rca24_fa301_xor0;
  wire s_dadda_pg_rca24_fa301_and0;
  wire s_dadda_pg_rca24_fa301_xor1;
  wire s_dadda_pg_rca24_fa301_and1;
  wire s_dadda_pg_rca24_fa301_or0;
  wire s_dadda_pg_rca24_and_13_22;
  wire s_dadda_pg_rca24_nand_12_23;
  wire s_dadda_pg_rca24_fa302_xor0;
  wire s_dadda_pg_rca24_fa302_and0;
  wire s_dadda_pg_rca24_fa302_xor1;
  wire s_dadda_pg_rca24_fa302_and1;
  wire s_dadda_pg_rca24_fa302_or0;
  wire s_dadda_pg_rca24_fa303_xor0;
  wire s_dadda_pg_rca24_fa303_and0;
  wire s_dadda_pg_rca24_fa303_xor1;
  wire s_dadda_pg_rca24_fa303_and1;
  wire s_dadda_pg_rca24_fa303_or0;
  wire s_dadda_pg_rca24_fa304_xor0;
  wire s_dadda_pg_rca24_fa304_and0;
  wire s_dadda_pg_rca24_fa304_xor1;
  wire s_dadda_pg_rca24_fa304_and1;
  wire s_dadda_pg_rca24_fa304_or0;
  wire s_dadda_pg_rca24_nand_23_13;
  wire s_dadda_pg_rca24_and_22_14;
  wire s_dadda_pg_rca24_fa305_xor0;
  wire s_dadda_pg_rca24_fa305_and0;
  wire s_dadda_pg_rca24_fa305_xor1;
  wire s_dadda_pg_rca24_fa305_and1;
  wire s_dadda_pg_rca24_fa305_or0;
  wire s_dadda_pg_rca24_and_21_15;
  wire s_dadda_pg_rca24_and_20_16;
  wire s_dadda_pg_rca24_and_19_17;
  wire s_dadda_pg_rca24_fa306_xor0;
  wire s_dadda_pg_rca24_fa306_and0;
  wire s_dadda_pg_rca24_fa306_xor1;
  wire s_dadda_pg_rca24_fa306_and1;
  wire s_dadda_pg_rca24_fa306_or0;
  wire s_dadda_pg_rca24_and_18_18;
  wire s_dadda_pg_rca24_and_17_19;
  wire s_dadda_pg_rca24_and_16_20;
  wire s_dadda_pg_rca24_fa307_xor0;
  wire s_dadda_pg_rca24_fa307_and0;
  wire s_dadda_pg_rca24_fa307_xor1;
  wire s_dadda_pg_rca24_fa307_and1;
  wire s_dadda_pg_rca24_fa307_or0;
  wire s_dadda_pg_rca24_and_15_21;
  wire s_dadda_pg_rca24_and_14_22;
  wire s_dadda_pg_rca24_nand_13_23;
  wire s_dadda_pg_rca24_fa308_xor0;
  wire s_dadda_pg_rca24_fa308_and0;
  wire s_dadda_pg_rca24_fa308_xor1;
  wire s_dadda_pg_rca24_fa308_and1;
  wire s_dadda_pg_rca24_fa308_or0;
  wire s_dadda_pg_rca24_fa309_xor0;
  wire s_dadda_pg_rca24_fa309_and0;
  wire s_dadda_pg_rca24_fa309_xor1;
  wire s_dadda_pg_rca24_fa309_and1;
  wire s_dadda_pg_rca24_fa309_or0;
  wire s_dadda_pg_rca24_fa310_xor0;
  wire s_dadda_pg_rca24_fa310_and0;
  wire s_dadda_pg_rca24_fa310_xor1;
  wire s_dadda_pg_rca24_fa310_and1;
  wire s_dadda_pg_rca24_fa310_or0;
  wire s_dadda_pg_rca24_nand_23_14;
  wire s_dadda_pg_rca24_and_22_15;
  wire s_dadda_pg_rca24_and_21_16;
  wire s_dadda_pg_rca24_fa311_xor0;
  wire s_dadda_pg_rca24_fa311_and0;
  wire s_dadda_pg_rca24_fa311_xor1;
  wire s_dadda_pg_rca24_fa311_and1;
  wire s_dadda_pg_rca24_fa311_or0;
  wire s_dadda_pg_rca24_and_20_17;
  wire s_dadda_pg_rca24_and_19_18;
  wire s_dadda_pg_rca24_and_18_19;
  wire s_dadda_pg_rca24_fa312_xor0;
  wire s_dadda_pg_rca24_fa312_and0;
  wire s_dadda_pg_rca24_fa312_xor1;
  wire s_dadda_pg_rca24_fa312_and1;
  wire s_dadda_pg_rca24_fa312_or0;
  wire s_dadda_pg_rca24_and_17_20;
  wire s_dadda_pg_rca24_and_16_21;
  wire s_dadda_pg_rca24_and_15_22;
  wire s_dadda_pg_rca24_fa313_xor0;
  wire s_dadda_pg_rca24_fa313_and0;
  wire s_dadda_pg_rca24_fa313_xor1;
  wire s_dadda_pg_rca24_fa313_and1;
  wire s_dadda_pg_rca24_fa313_or0;
  wire s_dadda_pg_rca24_fa314_xor0;
  wire s_dadda_pg_rca24_fa314_and0;
  wire s_dadda_pg_rca24_fa314_xor1;
  wire s_dadda_pg_rca24_fa314_and1;
  wire s_dadda_pg_rca24_fa314_or0;
  wire s_dadda_pg_rca24_nand_23_15;
  wire s_dadda_pg_rca24_fa315_xor0;
  wire s_dadda_pg_rca24_fa315_and0;
  wire s_dadda_pg_rca24_fa315_xor1;
  wire s_dadda_pg_rca24_fa315_and1;
  wire s_dadda_pg_rca24_fa315_or0;
  wire s_dadda_pg_rca24_and_22_16;
  wire s_dadda_pg_rca24_and_21_17;
  wire s_dadda_pg_rca24_and_20_18;
  wire s_dadda_pg_rca24_fa316_xor0;
  wire s_dadda_pg_rca24_fa316_and0;
  wire s_dadda_pg_rca24_fa316_xor1;
  wire s_dadda_pg_rca24_fa316_and1;
  wire s_dadda_pg_rca24_fa316_or0;
  wire s_dadda_pg_rca24_and_19_19;
  wire s_dadda_pg_rca24_and_18_20;
  wire s_dadda_pg_rca24_and_17_21;
  wire s_dadda_pg_rca24_fa317_xor0;
  wire s_dadda_pg_rca24_fa317_and0;
  wire s_dadda_pg_rca24_fa317_xor1;
  wire s_dadda_pg_rca24_fa317_and1;
  wire s_dadda_pg_rca24_fa317_or0;
  wire s_dadda_pg_rca24_fa318_xor0;
  wire s_dadda_pg_rca24_fa318_and0;
  wire s_dadda_pg_rca24_fa318_xor1;
  wire s_dadda_pg_rca24_fa318_and1;
  wire s_dadda_pg_rca24_fa318_or0;
  wire s_dadda_pg_rca24_nand_23_16;
  wire s_dadda_pg_rca24_and_22_17;
  wire s_dadda_pg_rca24_fa319_xor0;
  wire s_dadda_pg_rca24_fa319_and0;
  wire s_dadda_pg_rca24_fa319_xor1;
  wire s_dadda_pg_rca24_fa319_and1;
  wire s_dadda_pg_rca24_fa319_or0;
  wire s_dadda_pg_rca24_and_21_18;
  wire s_dadda_pg_rca24_and_20_19;
  wire s_dadda_pg_rca24_and_19_20;
  wire s_dadda_pg_rca24_fa320_xor0;
  wire s_dadda_pg_rca24_fa320_and0;
  wire s_dadda_pg_rca24_fa320_xor1;
  wire s_dadda_pg_rca24_fa320_and1;
  wire s_dadda_pg_rca24_fa320_or0;
  wire s_dadda_pg_rca24_fa321_xor0;
  wire s_dadda_pg_rca24_fa321_and0;
  wire s_dadda_pg_rca24_fa321_xor1;
  wire s_dadda_pg_rca24_fa321_and1;
  wire s_dadda_pg_rca24_fa321_or0;
  wire s_dadda_pg_rca24_nand_23_17;
  wire s_dadda_pg_rca24_and_22_18;
  wire s_dadda_pg_rca24_and_21_19;
  wire s_dadda_pg_rca24_fa322_xor0;
  wire s_dadda_pg_rca24_fa322_and0;
  wire s_dadda_pg_rca24_fa322_xor1;
  wire s_dadda_pg_rca24_fa322_and1;
  wire s_dadda_pg_rca24_fa322_or0;
  wire s_dadda_pg_rca24_nand_23_18;
  wire s_dadda_pg_rca24_fa323_xor0;
  wire s_dadda_pg_rca24_fa323_and0;
  wire s_dadda_pg_rca24_fa323_xor1;
  wire s_dadda_pg_rca24_fa323_and1;
  wire s_dadda_pg_rca24_fa323_or0;
  wire s_dadda_pg_rca24_and_4_0;
  wire s_dadda_pg_rca24_and_3_1;
  wire s_dadda_pg_rca24_ha18_xor0;
  wire s_dadda_pg_rca24_ha18_and0;
  wire s_dadda_pg_rca24_and_5_0;
  wire s_dadda_pg_rca24_and_4_1;
  wire s_dadda_pg_rca24_fa324_xor0;
  wire s_dadda_pg_rca24_fa324_and0;
  wire s_dadda_pg_rca24_fa324_xor1;
  wire s_dadda_pg_rca24_fa324_and1;
  wire s_dadda_pg_rca24_fa324_or0;
  wire s_dadda_pg_rca24_and_3_2;
  wire s_dadda_pg_rca24_and_2_3;
  wire s_dadda_pg_rca24_ha19_xor0;
  wire s_dadda_pg_rca24_ha19_and0;
  wire s_dadda_pg_rca24_and_4_2;
  wire s_dadda_pg_rca24_fa325_xor0;
  wire s_dadda_pg_rca24_fa325_and0;
  wire s_dadda_pg_rca24_fa325_xor1;
  wire s_dadda_pg_rca24_fa325_and1;
  wire s_dadda_pg_rca24_fa325_or0;
  wire s_dadda_pg_rca24_and_3_3;
  wire s_dadda_pg_rca24_and_2_4;
  wire s_dadda_pg_rca24_and_1_5;
  wire s_dadda_pg_rca24_fa326_xor0;
  wire s_dadda_pg_rca24_fa326_and0;
  wire s_dadda_pg_rca24_fa326_xor1;
  wire s_dadda_pg_rca24_fa326_and1;
  wire s_dadda_pg_rca24_fa326_or0;
  wire s_dadda_pg_rca24_and_3_4;
  wire s_dadda_pg_rca24_fa327_xor0;
  wire s_dadda_pg_rca24_fa327_and0;
  wire s_dadda_pg_rca24_fa327_xor1;
  wire s_dadda_pg_rca24_fa327_and1;
  wire s_dadda_pg_rca24_fa327_or0;
  wire s_dadda_pg_rca24_and_2_5;
  wire s_dadda_pg_rca24_and_1_6;
  wire s_dadda_pg_rca24_and_0_7;
  wire s_dadda_pg_rca24_fa328_xor0;
  wire s_dadda_pg_rca24_fa328_and0;
  wire s_dadda_pg_rca24_fa328_xor1;
  wire s_dadda_pg_rca24_fa328_and1;
  wire s_dadda_pg_rca24_fa328_or0;
  wire s_dadda_pg_rca24_and_2_6;
  wire s_dadda_pg_rca24_fa329_xor0;
  wire s_dadda_pg_rca24_fa329_and0;
  wire s_dadda_pg_rca24_fa329_xor1;
  wire s_dadda_pg_rca24_fa329_and1;
  wire s_dadda_pg_rca24_fa329_or0;
  wire s_dadda_pg_rca24_and_1_7;
  wire s_dadda_pg_rca24_and_0_8;
  wire s_dadda_pg_rca24_fa330_xor0;
  wire s_dadda_pg_rca24_fa330_and0;
  wire s_dadda_pg_rca24_fa330_xor1;
  wire s_dadda_pg_rca24_fa330_and1;
  wire s_dadda_pg_rca24_fa330_or0;
  wire s_dadda_pg_rca24_and_1_8;
  wire s_dadda_pg_rca24_fa331_xor0;
  wire s_dadda_pg_rca24_fa331_and0;
  wire s_dadda_pg_rca24_fa331_xor1;
  wire s_dadda_pg_rca24_fa331_and1;
  wire s_dadda_pg_rca24_fa331_or0;
  wire s_dadda_pg_rca24_and_0_9;
  wire s_dadda_pg_rca24_fa332_xor0;
  wire s_dadda_pg_rca24_fa332_and0;
  wire s_dadda_pg_rca24_fa332_xor1;
  wire s_dadda_pg_rca24_fa332_and1;
  wire s_dadda_pg_rca24_fa332_or0;
  wire s_dadda_pg_rca24_and_0_10;
  wire s_dadda_pg_rca24_fa333_xor0;
  wire s_dadda_pg_rca24_fa333_and0;
  wire s_dadda_pg_rca24_fa333_xor1;
  wire s_dadda_pg_rca24_fa333_and1;
  wire s_dadda_pg_rca24_fa333_or0;
  wire s_dadda_pg_rca24_fa334_xor0;
  wire s_dadda_pg_rca24_fa334_and0;
  wire s_dadda_pg_rca24_fa334_xor1;
  wire s_dadda_pg_rca24_fa334_and1;
  wire s_dadda_pg_rca24_fa334_or0;
  wire s_dadda_pg_rca24_fa335_xor0;
  wire s_dadda_pg_rca24_fa335_and0;
  wire s_dadda_pg_rca24_fa335_xor1;
  wire s_dadda_pg_rca24_fa335_and1;
  wire s_dadda_pg_rca24_fa335_or0;
  wire s_dadda_pg_rca24_fa336_xor0;
  wire s_dadda_pg_rca24_fa336_and0;
  wire s_dadda_pg_rca24_fa336_xor1;
  wire s_dadda_pg_rca24_fa336_and1;
  wire s_dadda_pg_rca24_fa336_or0;
  wire s_dadda_pg_rca24_fa337_xor0;
  wire s_dadda_pg_rca24_fa337_and0;
  wire s_dadda_pg_rca24_fa337_xor1;
  wire s_dadda_pg_rca24_fa337_and1;
  wire s_dadda_pg_rca24_fa337_or0;
  wire s_dadda_pg_rca24_fa338_xor0;
  wire s_dadda_pg_rca24_fa338_and0;
  wire s_dadda_pg_rca24_fa338_xor1;
  wire s_dadda_pg_rca24_fa338_and1;
  wire s_dadda_pg_rca24_fa338_or0;
  wire s_dadda_pg_rca24_fa339_xor0;
  wire s_dadda_pg_rca24_fa339_and0;
  wire s_dadda_pg_rca24_fa339_xor1;
  wire s_dadda_pg_rca24_fa339_and1;
  wire s_dadda_pg_rca24_fa339_or0;
  wire s_dadda_pg_rca24_fa340_xor0;
  wire s_dadda_pg_rca24_fa340_and0;
  wire s_dadda_pg_rca24_fa340_xor1;
  wire s_dadda_pg_rca24_fa340_and1;
  wire s_dadda_pg_rca24_fa340_or0;
  wire s_dadda_pg_rca24_fa341_xor0;
  wire s_dadda_pg_rca24_fa341_and0;
  wire s_dadda_pg_rca24_fa341_xor1;
  wire s_dadda_pg_rca24_fa341_and1;
  wire s_dadda_pg_rca24_fa341_or0;
  wire s_dadda_pg_rca24_fa342_xor0;
  wire s_dadda_pg_rca24_fa342_and0;
  wire s_dadda_pg_rca24_fa342_xor1;
  wire s_dadda_pg_rca24_fa342_and1;
  wire s_dadda_pg_rca24_fa342_or0;
  wire s_dadda_pg_rca24_fa343_xor0;
  wire s_dadda_pg_rca24_fa343_and0;
  wire s_dadda_pg_rca24_fa343_xor1;
  wire s_dadda_pg_rca24_fa343_and1;
  wire s_dadda_pg_rca24_fa343_or0;
  wire s_dadda_pg_rca24_fa344_xor0;
  wire s_dadda_pg_rca24_fa344_and0;
  wire s_dadda_pg_rca24_fa344_xor1;
  wire s_dadda_pg_rca24_fa344_and1;
  wire s_dadda_pg_rca24_fa344_or0;
  wire s_dadda_pg_rca24_fa345_xor0;
  wire s_dadda_pg_rca24_fa345_and0;
  wire s_dadda_pg_rca24_fa345_xor1;
  wire s_dadda_pg_rca24_fa345_and1;
  wire s_dadda_pg_rca24_fa345_or0;
  wire s_dadda_pg_rca24_fa346_xor0;
  wire s_dadda_pg_rca24_fa346_and0;
  wire s_dadda_pg_rca24_fa346_xor1;
  wire s_dadda_pg_rca24_fa346_and1;
  wire s_dadda_pg_rca24_fa346_or0;
  wire s_dadda_pg_rca24_fa347_xor0;
  wire s_dadda_pg_rca24_fa347_and0;
  wire s_dadda_pg_rca24_fa347_xor1;
  wire s_dadda_pg_rca24_fa347_and1;
  wire s_dadda_pg_rca24_fa347_or0;
  wire s_dadda_pg_rca24_fa348_xor0;
  wire s_dadda_pg_rca24_fa348_and0;
  wire s_dadda_pg_rca24_fa348_xor1;
  wire s_dadda_pg_rca24_fa348_and1;
  wire s_dadda_pg_rca24_fa348_or0;
  wire s_dadda_pg_rca24_fa349_xor0;
  wire s_dadda_pg_rca24_fa349_and0;
  wire s_dadda_pg_rca24_fa349_xor1;
  wire s_dadda_pg_rca24_fa349_and1;
  wire s_dadda_pg_rca24_fa349_or0;
  wire s_dadda_pg_rca24_fa350_xor0;
  wire s_dadda_pg_rca24_fa350_and0;
  wire s_dadda_pg_rca24_fa350_xor1;
  wire s_dadda_pg_rca24_fa350_and1;
  wire s_dadda_pg_rca24_fa350_or0;
  wire s_dadda_pg_rca24_fa351_xor0;
  wire s_dadda_pg_rca24_fa351_and0;
  wire s_dadda_pg_rca24_fa351_xor1;
  wire s_dadda_pg_rca24_fa351_and1;
  wire s_dadda_pg_rca24_fa351_or0;
  wire s_dadda_pg_rca24_fa352_xor0;
  wire s_dadda_pg_rca24_fa352_and0;
  wire s_dadda_pg_rca24_fa352_xor1;
  wire s_dadda_pg_rca24_fa352_and1;
  wire s_dadda_pg_rca24_fa352_or0;
  wire s_dadda_pg_rca24_fa353_xor0;
  wire s_dadda_pg_rca24_fa353_and0;
  wire s_dadda_pg_rca24_fa353_xor1;
  wire s_dadda_pg_rca24_fa353_and1;
  wire s_dadda_pg_rca24_fa353_or0;
  wire s_dadda_pg_rca24_fa354_xor0;
  wire s_dadda_pg_rca24_fa354_and0;
  wire s_dadda_pg_rca24_fa354_xor1;
  wire s_dadda_pg_rca24_fa354_and1;
  wire s_dadda_pg_rca24_fa354_or0;
  wire s_dadda_pg_rca24_fa355_xor0;
  wire s_dadda_pg_rca24_fa355_and0;
  wire s_dadda_pg_rca24_fa355_xor1;
  wire s_dadda_pg_rca24_fa355_and1;
  wire s_dadda_pg_rca24_fa355_or0;
  wire s_dadda_pg_rca24_fa356_xor0;
  wire s_dadda_pg_rca24_fa356_and0;
  wire s_dadda_pg_rca24_fa356_xor1;
  wire s_dadda_pg_rca24_fa356_and1;
  wire s_dadda_pg_rca24_fa356_or0;
  wire s_dadda_pg_rca24_fa357_xor0;
  wire s_dadda_pg_rca24_fa357_and0;
  wire s_dadda_pg_rca24_fa357_xor1;
  wire s_dadda_pg_rca24_fa357_and1;
  wire s_dadda_pg_rca24_fa357_or0;
  wire s_dadda_pg_rca24_fa358_xor0;
  wire s_dadda_pg_rca24_fa358_and0;
  wire s_dadda_pg_rca24_fa358_xor1;
  wire s_dadda_pg_rca24_fa358_and1;
  wire s_dadda_pg_rca24_fa358_or0;
  wire s_dadda_pg_rca24_fa359_xor0;
  wire s_dadda_pg_rca24_fa359_and0;
  wire s_dadda_pg_rca24_fa359_xor1;
  wire s_dadda_pg_rca24_fa359_and1;
  wire s_dadda_pg_rca24_fa359_or0;
  wire s_dadda_pg_rca24_fa360_xor0;
  wire s_dadda_pg_rca24_fa360_and0;
  wire s_dadda_pg_rca24_fa360_xor1;
  wire s_dadda_pg_rca24_fa360_and1;
  wire s_dadda_pg_rca24_fa360_or0;
  wire s_dadda_pg_rca24_fa361_xor0;
  wire s_dadda_pg_rca24_fa361_and0;
  wire s_dadda_pg_rca24_fa361_xor1;
  wire s_dadda_pg_rca24_fa361_and1;
  wire s_dadda_pg_rca24_fa361_or0;
  wire s_dadda_pg_rca24_fa362_xor0;
  wire s_dadda_pg_rca24_fa362_and0;
  wire s_dadda_pg_rca24_fa362_xor1;
  wire s_dadda_pg_rca24_fa362_and1;
  wire s_dadda_pg_rca24_fa362_or0;
  wire s_dadda_pg_rca24_fa363_xor0;
  wire s_dadda_pg_rca24_fa363_and0;
  wire s_dadda_pg_rca24_fa363_xor1;
  wire s_dadda_pg_rca24_fa363_and1;
  wire s_dadda_pg_rca24_fa363_or0;
  wire s_dadda_pg_rca24_fa364_xor0;
  wire s_dadda_pg_rca24_fa364_and0;
  wire s_dadda_pg_rca24_fa364_xor1;
  wire s_dadda_pg_rca24_fa364_and1;
  wire s_dadda_pg_rca24_fa364_or0;
  wire s_dadda_pg_rca24_fa365_xor0;
  wire s_dadda_pg_rca24_fa365_and0;
  wire s_dadda_pg_rca24_fa365_xor1;
  wire s_dadda_pg_rca24_fa365_and1;
  wire s_dadda_pg_rca24_fa365_or0;
  wire s_dadda_pg_rca24_fa366_xor0;
  wire s_dadda_pg_rca24_fa366_and0;
  wire s_dadda_pg_rca24_fa366_xor1;
  wire s_dadda_pg_rca24_fa366_and1;
  wire s_dadda_pg_rca24_fa366_or0;
  wire s_dadda_pg_rca24_fa367_xor0;
  wire s_dadda_pg_rca24_fa367_and0;
  wire s_dadda_pg_rca24_fa367_xor1;
  wire s_dadda_pg_rca24_fa367_and1;
  wire s_dadda_pg_rca24_fa367_or0;
  wire s_dadda_pg_rca24_fa368_xor0;
  wire s_dadda_pg_rca24_fa368_and0;
  wire s_dadda_pg_rca24_fa368_xor1;
  wire s_dadda_pg_rca24_fa368_and1;
  wire s_dadda_pg_rca24_fa368_or0;
  wire s_dadda_pg_rca24_fa369_xor0;
  wire s_dadda_pg_rca24_fa369_and0;
  wire s_dadda_pg_rca24_fa369_xor1;
  wire s_dadda_pg_rca24_fa369_and1;
  wire s_dadda_pg_rca24_fa369_or0;
  wire s_dadda_pg_rca24_fa370_xor0;
  wire s_dadda_pg_rca24_fa370_and0;
  wire s_dadda_pg_rca24_fa370_xor1;
  wire s_dadda_pg_rca24_fa370_and1;
  wire s_dadda_pg_rca24_fa370_or0;
  wire s_dadda_pg_rca24_fa371_xor0;
  wire s_dadda_pg_rca24_fa371_and0;
  wire s_dadda_pg_rca24_fa371_xor1;
  wire s_dadda_pg_rca24_fa371_and1;
  wire s_dadda_pg_rca24_fa371_or0;
  wire s_dadda_pg_rca24_fa372_xor0;
  wire s_dadda_pg_rca24_fa372_and0;
  wire s_dadda_pg_rca24_fa372_xor1;
  wire s_dadda_pg_rca24_fa372_and1;
  wire s_dadda_pg_rca24_fa372_or0;
  wire s_dadda_pg_rca24_fa373_xor0;
  wire s_dadda_pg_rca24_fa373_and0;
  wire s_dadda_pg_rca24_fa373_xor1;
  wire s_dadda_pg_rca24_fa373_and1;
  wire s_dadda_pg_rca24_fa373_or0;
  wire s_dadda_pg_rca24_fa374_xor0;
  wire s_dadda_pg_rca24_fa374_and0;
  wire s_dadda_pg_rca24_fa374_xor1;
  wire s_dadda_pg_rca24_fa374_and1;
  wire s_dadda_pg_rca24_fa374_or0;
  wire s_dadda_pg_rca24_fa375_xor0;
  wire s_dadda_pg_rca24_fa375_and0;
  wire s_dadda_pg_rca24_fa375_xor1;
  wire s_dadda_pg_rca24_fa375_and1;
  wire s_dadda_pg_rca24_fa375_or0;
  wire s_dadda_pg_rca24_fa376_xor0;
  wire s_dadda_pg_rca24_fa376_and0;
  wire s_dadda_pg_rca24_fa376_xor1;
  wire s_dadda_pg_rca24_fa376_and1;
  wire s_dadda_pg_rca24_fa376_or0;
  wire s_dadda_pg_rca24_fa377_xor0;
  wire s_dadda_pg_rca24_fa377_and0;
  wire s_dadda_pg_rca24_fa377_xor1;
  wire s_dadda_pg_rca24_fa377_and1;
  wire s_dadda_pg_rca24_fa377_or0;
  wire s_dadda_pg_rca24_fa378_xor0;
  wire s_dadda_pg_rca24_fa378_and0;
  wire s_dadda_pg_rca24_fa378_xor1;
  wire s_dadda_pg_rca24_fa378_and1;
  wire s_dadda_pg_rca24_fa378_or0;
  wire s_dadda_pg_rca24_fa379_xor0;
  wire s_dadda_pg_rca24_fa379_and0;
  wire s_dadda_pg_rca24_fa379_xor1;
  wire s_dadda_pg_rca24_fa379_and1;
  wire s_dadda_pg_rca24_fa379_or0;
  wire s_dadda_pg_rca24_fa380_xor0;
  wire s_dadda_pg_rca24_fa380_and0;
  wire s_dadda_pg_rca24_fa380_xor1;
  wire s_dadda_pg_rca24_fa380_and1;
  wire s_dadda_pg_rca24_fa380_or0;
  wire s_dadda_pg_rca24_fa381_xor0;
  wire s_dadda_pg_rca24_fa381_and0;
  wire s_dadda_pg_rca24_fa381_xor1;
  wire s_dadda_pg_rca24_fa381_and1;
  wire s_dadda_pg_rca24_fa381_or0;
  wire s_dadda_pg_rca24_fa382_xor0;
  wire s_dadda_pg_rca24_fa382_and0;
  wire s_dadda_pg_rca24_fa382_xor1;
  wire s_dadda_pg_rca24_fa382_and1;
  wire s_dadda_pg_rca24_fa382_or0;
  wire s_dadda_pg_rca24_fa383_xor0;
  wire s_dadda_pg_rca24_fa383_and0;
  wire s_dadda_pg_rca24_fa383_xor1;
  wire s_dadda_pg_rca24_fa383_and1;
  wire s_dadda_pg_rca24_fa383_or0;
  wire s_dadda_pg_rca24_fa384_xor0;
  wire s_dadda_pg_rca24_fa384_and0;
  wire s_dadda_pg_rca24_fa384_xor1;
  wire s_dadda_pg_rca24_fa384_and1;
  wire s_dadda_pg_rca24_fa384_or0;
  wire s_dadda_pg_rca24_fa385_xor0;
  wire s_dadda_pg_rca24_fa385_and0;
  wire s_dadda_pg_rca24_fa385_xor1;
  wire s_dadda_pg_rca24_fa385_and1;
  wire s_dadda_pg_rca24_fa385_or0;
  wire s_dadda_pg_rca24_fa386_xor0;
  wire s_dadda_pg_rca24_fa386_and0;
  wire s_dadda_pg_rca24_fa386_xor1;
  wire s_dadda_pg_rca24_fa386_and1;
  wire s_dadda_pg_rca24_fa386_or0;
  wire s_dadda_pg_rca24_nand_14_23;
  wire s_dadda_pg_rca24_fa387_xor0;
  wire s_dadda_pg_rca24_fa387_and0;
  wire s_dadda_pg_rca24_fa387_xor1;
  wire s_dadda_pg_rca24_fa387_and1;
  wire s_dadda_pg_rca24_fa387_or0;
  wire s_dadda_pg_rca24_fa388_xor0;
  wire s_dadda_pg_rca24_fa388_and0;
  wire s_dadda_pg_rca24_fa388_xor1;
  wire s_dadda_pg_rca24_fa388_and1;
  wire s_dadda_pg_rca24_fa388_or0;
  wire s_dadda_pg_rca24_and_16_22;
  wire s_dadda_pg_rca24_fa389_xor0;
  wire s_dadda_pg_rca24_fa389_and0;
  wire s_dadda_pg_rca24_fa389_xor1;
  wire s_dadda_pg_rca24_fa389_and1;
  wire s_dadda_pg_rca24_fa389_or0;
  wire s_dadda_pg_rca24_nand_15_23;
  wire s_dadda_pg_rca24_fa390_xor0;
  wire s_dadda_pg_rca24_fa390_and0;
  wire s_dadda_pg_rca24_fa390_xor1;
  wire s_dadda_pg_rca24_fa390_and1;
  wire s_dadda_pg_rca24_fa390_or0;
  wire s_dadda_pg_rca24_and_18_21;
  wire s_dadda_pg_rca24_fa391_xor0;
  wire s_dadda_pg_rca24_fa391_and0;
  wire s_dadda_pg_rca24_fa391_xor1;
  wire s_dadda_pg_rca24_fa391_and1;
  wire s_dadda_pg_rca24_fa391_or0;
  wire s_dadda_pg_rca24_and_17_22;
  wire s_dadda_pg_rca24_nand_16_23;
  wire s_dadda_pg_rca24_fa392_xor0;
  wire s_dadda_pg_rca24_fa392_and0;
  wire s_dadda_pg_rca24_fa392_xor1;
  wire s_dadda_pg_rca24_fa392_and1;
  wire s_dadda_pg_rca24_fa392_or0;
  wire s_dadda_pg_rca24_and_20_20;
  wire s_dadda_pg_rca24_fa393_xor0;
  wire s_dadda_pg_rca24_fa393_and0;
  wire s_dadda_pg_rca24_fa393_xor1;
  wire s_dadda_pg_rca24_fa393_and1;
  wire s_dadda_pg_rca24_fa393_or0;
  wire s_dadda_pg_rca24_and_19_21;
  wire s_dadda_pg_rca24_and_18_22;
  wire s_dadda_pg_rca24_nand_17_23;
  wire s_dadda_pg_rca24_fa394_xor0;
  wire s_dadda_pg_rca24_fa394_and0;
  wire s_dadda_pg_rca24_fa394_xor1;
  wire s_dadda_pg_rca24_fa394_and1;
  wire s_dadda_pg_rca24_fa394_or0;
  wire s_dadda_pg_rca24_and_22_19;
  wire s_dadda_pg_rca24_fa395_xor0;
  wire s_dadda_pg_rca24_fa395_and0;
  wire s_dadda_pg_rca24_fa395_xor1;
  wire s_dadda_pg_rca24_fa395_and1;
  wire s_dadda_pg_rca24_fa395_or0;
  wire s_dadda_pg_rca24_and_21_20;
  wire s_dadda_pg_rca24_and_20_21;
  wire s_dadda_pg_rca24_and_19_22;
  wire s_dadda_pg_rca24_fa396_xor0;
  wire s_dadda_pg_rca24_fa396_and0;
  wire s_dadda_pg_rca24_fa396_xor1;
  wire s_dadda_pg_rca24_fa396_and1;
  wire s_dadda_pg_rca24_fa396_or0;
  wire s_dadda_pg_rca24_fa397_xor0;
  wire s_dadda_pg_rca24_fa397_and0;
  wire s_dadda_pg_rca24_fa397_xor1;
  wire s_dadda_pg_rca24_fa397_and1;
  wire s_dadda_pg_rca24_fa397_or0;
  wire s_dadda_pg_rca24_nand_23_19;
  wire s_dadda_pg_rca24_and_22_20;
  wire s_dadda_pg_rca24_and_21_21;
  wire s_dadda_pg_rca24_fa398_xor0;
  wire s_dadda_pg_rca24_fa398_and0;
  wire s_dadda_pg_rca24_fa398_xor1;
  wire s_dadda_pg_rca24_fa398_and1;
  wire s_dadda_pg_rca24_fa398_or0;
  wire s_dadda_pg_rca24_nand_23_20;
  wire s_dadda_pg_rca24_fa399_xor0;
  wire s_dadda_pg_rca24_fa399_and0;
  wire s_dadda_pg_rca24_fa399_xor1;
  wire s_dadda_pg_rca24_fa399_and1;
  wire s_dadda_pg_rca24_fa399_or0;
  wire s_dadda_pg_rca24_and_3_0;
  wire s_dadda_pg_rca24_and_2_1;
  wire s_dadda_pg_rca24_ha20_xor0;
  wire s_dadda_pg_rca24_ha20_and0;
  wire s_dadda_pg_rca24_and_2_2;
  wire s_dadda_pg_rca24_and_1_3;
  wire s_dadda_pg_rca24_fa400_xor0;
  wire s_dadda_pg_rca24_fa400_and0;
  wire s_dadda_pg_rca24_fa400_xor1;
  wire s_dadda_pg_rca24_fa400_and1;
  wire s_dadda_pg_rca24_fa400_or0;
  wire s_dadda_pg_rca24_and_1_4;
  wire s_dadda_pg_rca24_and_0_5;
  wire s_dadda_pg_rca24_fa401_xor0;
  wire s_dadda_pg_rca24_fa401_and0;
  wire s_dadda_pg_rca24_fa401_xor1;
  wire s_dadda_pg_rca24_fa401_and1;
  wire s_dadda_pg_rca24_fa401_or0;
  wire s_dadda_pg_rca24_and_0_6;
  wire s_dadda_pg_rca24_fa402_xor0;
  wire s_dadda_pg_rca24_fa402_and0;
  wire s_dadda_pg_rca24_fa402_xor1;
  wire s_dadda_pg_rca24_fa402_and1;
  wire s_dadda_pg_rca24_fa402_or0;
  wire s_dadda_pg_rca24_fa403_xor0;
  wire s_dadda_pg_rca24_fa403_and0;
  wire s_dadda_pg_rca24_fa403_xor1;
  wire s_dadda_pg_rca24_fa403_and1;
  wire s_dadda_pg_rca24_fa403_or0;
  wire s_dadda_pg_rca24_fa404_xor0;
  wire s_dadda_pg_rca24_fa404_and0;
  wire s_dadda_pg_rca24_fa404_xor1;
  wire s_dadda_pg_rca24_fa404_and1;
  wire s_dadda_pg_rca24_fa404_or0;
  wire s_dadda_pg_rca24_fa405_xor0;
  wire s_dadda_pg_rca24_fa405_and0;
  wire s_dadda_pg_rca24_fa405_xor1;
  wire s_dadda_pg_rca24_fa405_and1;
  wire s_dadda_pg_rca24_fa405_or0;
  wire s_dadda_pg_rca24_fa406_xor0;
  wire s_dadda_pg_rca24_fa406_and0;
  wire s_dadda_pg_rca24_fa406_xor1;
  wire s_dadda_pg_rca24_fa406_and1;
  wire s_dadda_pg_rca24_fa406_or0;
  wire s_dadda_pg_rca24_fa407_xor0;
  wire s_dadda_pg_rca24_fa407_and0;
  wire s_dadda_pg_rca24_fa407_xor1;
  wire s_dadda_pg_rca24_fa407_and1;
  wire s_dadda_pg_rca24_fa407_or0;
  wire s_dadda_pg_rca24_fa408_xor0;
  wire s_dadda_pg_rca24_fa408_and0;
  wire s_dadda_pg_rca24_fa408_xor1;
  wire s_dadda_pg_rca24_fa408_and1;
  wire s_dadda_pg_rca24_fa408_or0;
  wire s_dadda_pg_rca24_fa409_xor0;
  wire s_dadda_pg_rca24_fa409_and0;
  wire s_dadda_pg_rca24_fa409_xor1;
  wire s_dadda_pg_rca24_fa409_and1;
  wire s_dadda_pg_rca24_fa409_or0;
  wire s_dadda_pg_rca24_fa410_xor0;
  wire s_dadda_pg_rca24_fa410_and0;
  wire s_dadda_pg_rca24_fa410_xor1;
  wire s_dadda_pg_rca24_fa410_and1;
  wire s_dadda_pg_rca24_fa410_or0;
  wire s_dadda_pg_rca24_fa411_xor0;
  wire s_dadda_pg_rca24_fa411_and0;
  wire s_dadda_pg_rca24_fa411_xor1;
  wire s_dadda_pg_rca24_fa411_and1;
  wire s_dadda_pg_rca24_fa411_or0;
  wire s_dadda_pg_rca24_fa412_xor0;
  wire s_dadda_pg_rca24_fa412_and0;
  wire s_dadda_pg_rca24_fa412_xor1;
  wire s_dadda_pg_rca24_fa412_and1;
  wire s_dadda_pg_rca24_fa412_or0;
  wire s_dadda_pg_rca24_fa413_xor0;
  wire s_dadda_pg_rca24_fa413_and0;
  wire s_dadda_pg_rca24_fa413_xor1;
  wire s_dadda_pg_rca24_fa413_and1;
  wire s_dadda_pg_rca24_fa413_or0;
  wire s_dadda_pg_rca24_fa414_xor0;
  wire s_dadda_pg_rca24_fa414_and0;
  wire s_dadda_pg_rca24_fa414_xor1;
  wire s_dadda_pg_rca24_fa414_and1;
  wire s_dadda_pg_rca24_fa414_or0;
  wire s_dadda_pg_rca24_fa415_xor0;
  wire s_dadda_pg_rca24_fa415_and0;
  wire s_dadda_pg_rca24_fa415_xor1;
  wire s_dadda_pg_rca24_fa415_and1;
  wire s_dadda_pg_rca24_fa415_or0;
  wire s_dadda_pg_rca24_fa416_xor0;
  wire s_dadda_pg_rca24_fa416_and0;
  wire s_dadda_pg_rca24_fa416_xor1;
  wire s_dadda_pg_rca24_fa416_and1;
  wire s_dadda_pg_rca24_fa416_or0;
  wire s_dadda_pg_rca24_fa417_xor0;
  wire s_dadda_pg_rca24_fa417_and0;
  wire s_dadda_pg_rca24_fa417_xor1;
  wire s_dadda_pg_rca24_fa417_and1;
  wire s_dadda_pg_rca24_fa417_or0;
  wire s_dadda_pg_rca24_fa418_xor0;
  wire s_dadda_pg_rca24_fa418_and0;
  wire s_dadda_pg_rca24_fa418_xor1;
  wire s_dadda_pg_rca24_fa418_and1;
  wire s_dadda_pg_rca24_fa418_or0;
  wire s_dadda_pg_rca24_fa419_xor0;
  wire s_dadda_pg_rca24_fa419_and0;
  wire s_dadda_pg_rca24_fa419_xor1;
  wire s_dadda_pg_rca24_fa419_and1;
  wire s_dadda_pg_rca24_fa419_or0;
  wire s_dadda_pg_rca24_fa420_xor0;
  wire s_dadda_pg_rca24_fa420_and0;
  wire s_dadda_pg_rca24_fa420_xor1;
  wire s_dadda_pg_rca24_fa420_and1;
  wire s_dadda_pg_rca24_fa420_or0;
  wire s_dadda_pg_rca24_fa421_xor0;
  wire s_dadda_pg_rca24_fa421_and0;
  wire s_dadda_pg_rca24_fa421_xor1;
  wire s_dadda_pg_rca24_fa421_and1;
  wire s_dadda_pg_rca24_fa421_or0;
  wire s_dadda_pg_rca24_fa422_xor0;
  wire s_dadda_pg_rca24_fa422_and0;
  wire s_dadda_pg_rca24_fa422_xor1;
  wire s_dadda_pg_rca24_fa422_and1;
  wire s_dadda_pg_rca24_fa422_or0;
  wire s_dadda_pg_rca24_fa423_xor0;
  wire s_dadda_pg_rca24_fa423_and0;
  wire s_dadda_pg_rca24_fa423_xor1;
  wire s_dadda_pg_rca24_fa423_and1;
  wire s_dadda_pg_rca24_fa423_or0;
  wire s_dadda_pg_rca24_fa424_xor0;
  wire s_dadda_pg_rca24_fa424_and0;
  wire s_dadda_pg_rca24_fa424_xor1;
  wire s_dadda_pg_rca24_fa424_and1;
  wire s_dadda_pg_rca24_fa424_or0;
  wire s_dadda_pg_rca24_fa425_xor0;
  wire s_dadda_pg_rca24_fa425_and0;
  wire s_dadda_pg_rca24_fa425_xor1;
  wire s_dadda_pg_rca24_fa425_and1;
  wire s_dadda_pg_rca24_fa425_or0;
  wire s_dadda_pg_rca24_fa426_xor0;
  wire s_dadda_pg_rca24_fa426_and0;
  wire s_dadda_pg_rca24_fa426_xor1;
  wire s_dadda_pg_rca24_fa426_and1;
  wire s_dadda_pg_rca24_fa426_or0;
  wire s_dadda_pg_rca24_fa427_xor0;
  wire s_dadda_pg_rca24_fa427_and0;
  wire s_dadda_pg_rca24_fa427_xor1;
  wire s_dadda_pg_rca24_fa427_and1;
  wire s_dadda_pg_rca24_fa427_or0;
  wire s_dadda_pg_rca24_fa428_xor0;
  wire s_dadda_pg_rca24_fa428_and0;
  wire s_dadda_pg_rca24_fa428_xor1;
  wire s_dadda_pg_rca24_fa428_and1;
  wire s_dadda_pg_rca24_fa428_or0;
  wire s_dadda_pg_rca24_fa429_xor0;
  wire s_dadda_pg_rca24_fa429_and0;
  wire s_dadda_pg_rca24_fa429_xor1;
  wire s_dadda_pg_rca24_fa429_and1;
  wire s_dadda_pg_rca24_fa429_or0;
  wire s_dadda_pg_rca24_fa430_xor0;
  wire s_dadda_pg_rca24_fa430_and0;
  wire s_dadda_pg_rca24_fa430_xor1;
  wire s_dadda_pg_rca24_fa430_and1;
  wire s_dadda_pg_rca24_fa430_or0;
  wire s_dadda_pg_rca24_fa431_xor0;
  wire s_dadda_pg_rca24_fa431_and0;
  wire s_dadda_pg_rca24_fa431_xor1;
  wire s_dadda_pg_rca24_fa431_and1;
  wire s_dadda_pg_rca24_fa431_or0;
  wire s_dadda_pg_rca24_fa432_xor0;
  wire s_dadda_pg_rca24_fa432_and0;
  wire s_dadda_pg_rca24_fa432_xor1;
  wire s_dadda_pg_rca24_fa432_and1;
  wire s_dadda_pg_rca24_fa432_or0;
  wire s_dadda_pg_rca24_fa433_xor0;
  wire s_dadda_pg_rca24_fa433_and0;
  wire s_dadda_pg_rca24_fa433_xor1;
  wire s_dadda_pg_rca24_fa433_and1;
  wire s_dadda_pg_rca24_fa433_or0;
  wire s_dadda_pg_rca24_fa434_xor0;
  wire s_dadda_pg_rca24_fa434_and0;
  wire s_dadda_pg_rca24_fa434_xor1;
  wire s_dadda_pg_rca24_fa434_and1;
  wire s_dadda_pg_rca24_fa434_or0;
  wire s_dadda_pg_rca24_fa435_xor0;
  wire s_dadda_pg_rca24_fa435_and0;
  wire s_dadda_pg_rca24_fa435_xor1;
  wire s_dadda_pg_rca24_fa435_and1;
  wire s_dadda_pg_rca24_fa435_or0;
  wire s_dadda_pg_rca24_fa436_xor0;
  wire s_dadda_pg_rca24_fa436_and0;
  wire s_dadda_pg_rca24_fa436_xor1;
  wire s_dadda_pg_rca24_fa436_and1;
  wire s_dadda_pg_rca24_fa436_or0;
  wire s_dadda_pg_rca24_nand_18_23;
  wire s_dadda_pg_rca24_fa437_xor0;
  wire s_dadda_pg_rca24_fa437_and0;
  wire s_dadda_pg_rca24_fa437_xor1;
  wire s_dadda_pg_rca24_fa437_and1;
  wire s_dadda_pg_rca24_fa437_or0;
  wire s_dadda_pg_rca24_and_20_22;
  wire s_dadda_pg_rca24_nand_19_23;
  wire s_dadda_pg_rca24_fa438_xor0;
  wire s_dadda_pg_rca24_fa438_and0;
  wire s_dadda_pg_rca24_fa438_xor1;
  wire s_dadda_pg_rca24_fa438_and1;
  wire s_dadda_pg_rca24_fa438_or0;
  wire s_dadda_pg_rca24_and_22_21;
  wire s_dadda_pg_rca24_and_21_22;
  wire s_dadda_pg_rca24_fa439_xor0;
  wire s_dadda_pg_rca24_fa439_and0;
  wire s_dadda_pg_rca24_fa439_xor1;
  wire s_dadda_pg_rca24_fa439_and1;
  wire s_dadda_pg_rca24_fa439_or0;
  wire s_dadda_pg_rca24_nand_23_21;
  wire s_dadda_pg_rca24_fa440_xor0;
  wire s_dadda_pg_rca24_fa440_and0;
  wire s_dadda_pg_rca24_fa440_xor1;
  wire s_dadda_pg_rca24_fa440_and1;
  wire s_dadda_pg_rca24_fa440_or0;
  wire s_dadda_pg_rca24_and_2_0;
  wire s_dadda_pg_rca24_and_1_1;
  wire s_dadda_pg_rca24_ha21_xor0;
  wire s_dadda_pg_rca24_ha21_and0;
  wire s_dadda_pg_rca24_and_1_2;
  wire s_dadda_pg_rca24_and_0_3;
  wire s_dadda_pg_rca24_fa441_xor0;
  wire s_dadda_pg_rca24_fa441_and0;
  wire s_dadda_pg_rca24_fa441_xor1;
  wire s_dadda_pg_rca24_fa441_and1;
  wire s_dadda_pg_rca24_fa441_or0;
  wire s_dadda_pg_rca24_and_0_4;
  wire s_dadda_pg_rca24_fa442_xor0;
  wire s_dadda_pg_rca24_fa442_and0;
  wire s_dadda_pg_rca24_fa442_xor1;
  wire s_dadda_pg_rca24_fa442_and1;
  wire s_dadda_pg_rca24_fa442_or0;
  wire s_dadda_pg_rca24_fa443_xor0;
  wire s_dadda_pg_rca24_fa443_and0;
  wire s_dadda_pg_rca24_fa443_xor1;
  wire s_dadda_pg_rca24_fa443_and1;
  wire s_dadda_pg_rca24_fa443_or0;
  wire s_dadda_pg_rca24_fa444_xor0;
  wire s_dadda_pg_rca24_fa444_and0;
  wire s_dadda_pg_rca24_fa444_xor1;
  wire s_dadda_pg_rca24_fa444_and1;
  wire s_dadda_pg_rca24_fa444_or0;
  wire s_dadda_pg_rca24_fa445_xor0;
  wire s_dadda_pg_rca24_fa445_and0;
  wire s_dadda_pg_rca24_fa445_xor1;
  wire s_dadda_pg_rca24_fa445_and1;
  wire s_dadda_pg_rca24_fa445_or0;
  wire s_dadda_pg_rca24_fa446_xor0;
  wire s_dadda_pg_rca24_fa446_and0;
  wire s_dadda_pg_rca24_fa446_xor1;
  wire s_dadda_pg_rca24_fa446_and1;
  wire s_dadda_pg_rca24_fa446_or0;
  wire s_dadda_pg_rca24_fa447_xor0;
  wire s_dadda_pg_rca24_fa447_and0;
  wire s_dadda_pg_rca24_fa447_xor1;
  wire s_dadda_pg_rca24_fa447_and1;
  wire s_dadda_pg_rca24_fa447_or0;
  wire s_dadda_pg_rca24_fa448_xor0;
  wire s_dadda_pg_rca24_fa448_and0;
  wire s_dadda_pg_rca24_fa448_xor1;
  wire s_dadda_pg_rca24_fa448_and1;
  wire s_dadda_pg_rca24_fa448_or0;
  wire s_dadda_pg_rca24_fa449_xor0;
  wire s_dadda_pg_rca24_fa449_and0;
  wire s_dadda_pg_rca24_fa449_xor1;
  wire s_dadda_pg_rca24_fa449_and1;
  wire s_dadda_pg_rca24_fa449_or0;
  wire s_dadda_pg_rca24_fa450_xor0;
  wire s_dadda_pg_rca24_fa450_and0;
  wire s_dadda_pg_rca24_fa450_xor1;
  wire s_dadda_pg_rca24_fa450_and1;
  wire s_dadda_pg_rca24_fa450_or0;
  wire s_dadda_pg_rca24_fa451_xor0;
  wire s_dadda_pg_rca24_fa451_and0;
  wire s_dadda_pg_rca24_fa451_xor1;
  wire s_dadda_pg_rca24_fa451_and1;
  wire s_dadda_pg_rca24_fa451_or0;
  wire s_dadda_pg_rca24_fa452_xor0;
  wire s_dadda_pg_rca24_fa452_and0;
  wire s_dadda_pg_rca24_fa452_xor1;
  wire s_dadda_pg_rca24_fa452_and1;
  wire s_dadda_pg_rca24_fa452_or0;
  wire s_dadda_pg_rca24_fa453_xor0;
  wire s_dadda_pg_rca24_fa453_and0;
  wire s_dadda_pg_rca24_fa453_xor1;
  wire s_dadda_pg_rca24_fa453_and1;
  wire s_dadda_pg_rca24_fa453_or0;
  wire s_dadda_pg_rca24_fa454_xor0;
  wire s_dadda_pg_rca24_fa454_and0;
  wire s_dadda_pg_rca24_fa454_xor1;
  wire s_dadda_pg_rca24_fa454_and1;
  wire s_dadda_pg_rca24_fa454_or0;
  wire s_dadda_pg_rca24_fa455_xor0;
  wire s_dadda_pg_rca24_fa455_and0;
  wire s_dadda_pg_rca24_fa455_xor1;
  wire s_dadda_pg_rca24_fa455_and1;
  wire s_dadda_pg_rca24_fa455_or0;
  wire s_dadda_pg_rca24_fa456_xor0;
  wire s_dadda_pg_rca24_fa456_and0;
  wire s_dadda_pg_rca24_fa456_xor1;
  wire s_dadda_pg_rca24_fa456_and1;
  wire s_dadda_pg_rca24_fa456_or0;
  wire s_dadda_pg_rca24_fa457_xor0;
  wire s_dadda_pg_rca24_fa457_and0;
  wire s_dadda_pg_rca24_fa457_xor1;
  wire s_dadda_pg_rca24_fa457_and1;
  wire s_dadda_pg_rca24_fa457_or0;
  wire s_dadda_pg_rca24_fa458_xor0;
  wire s_dadda_pg_rca24_fa458_and0;
  wire s_dadda_pg_rca24_fa458_xor1;
  wire s_dadda_pg_rca24_fa458_and1;
  wire s_dadda_pg_rca24_fa458_or0;
  wire s_dadda_pg_rca24_fa459_xor0;
  wire s_dadda_pg_rca24_fa459_and0;
  wire s_dadda_pg_rca24_fa459_xor1;
  wire s_dadda_pg_rca24_fa459_and1;
  wire s_dadda_pg_rca24_fa459_or0;
  wire s_dadda_pg_rca24_fa460_xor0;
  wire s_dadda_pg_rca24_fa460_and0;
  wire s_dadda_pg_rca24_fa460_xor1;
  wire s_dadda_pg_rca24_fa460_and1;
  wire s_dadda_pg_rca24_fa460_or0;
  wire s_dadda_pg_rca24_fa461_xor0;
  wire s_dadda_pg_rca24_fa461_and0;
  wire s_dadda_pg_rca24_fa461_xor1;
  wire s_dadda_pg_rca24_fa461_and1;
  wire s_dadda_pg_rca24_fa461_or0;
  wire s_dadda_pg_rca24_fa462_xor0;
  wire s_dadda_pg_rca24_fa462_and0;
  wire s_dadda_pg_rca24_fa462_xor1;
  wire s_dadda_pg_rca24_fa462_and1;
  wire s_dadda_pg_rca24_fa462_or0;
  wire s_dadda_pg_rca24_fa463_xor0;
  wire s_dadda_pg_rca24_fa463_and0;
  wire s_dadda_pg_rca24_fa463_xor1;
  wire s_dadda_pg_rca24_fa463_and1;
  wire s_dadda_pg_rca24_fa463_or0;
  wire s_dadda_pg_rca24_fa464_xor0;
  wire s_dadda_pg_rca24_fa464_and0;
  wire s_dadda_pg_rca24_fa464_xor1;
  wire s_dadda_pg_rca24_fa464_and1;
  wire s_dadda_pg_rca24_fa464_or0;
  wire s_dadda_pg_rca24_fa465_xor0;
  wire s_dadda_pg_rca24_fa465_and0;
  wire s_dadda_pg_rca24_fa465_xor1;
  wire s_dadda_pg_rca24_fa465_and1;
  wire s_dadda_pg_rca24_fa465_or0;
  wire s_dadda_pg_rca24_fa466_xor0;
  wire s_dadda_pg_rca24_fa466_and0;
  wire s_dadda_pg_rca24_fa466_xor1;
  wire s_dadda_pg_rca24_fa466_and1;
  wire s_dadda_pg_rca24_fa466_or0;
  wire s_dadda_pg_rca24_fa467_xor0;
  wire s_dadda_pg_rca24_fa467_and0;
  wire s_dadda_pg_rca24_fa467_xor1;
  wire s_dadda_pg_rca24_fa467_and1;
  wire s_dadda_pg_rca24_fa467_or0;
  wire s_dadda_pg_rca24_fa468_xor0;
  wire s_dadda_pg_rca24_fa468_and0;
  wire s_dadda_pg_rca24_fa468_xor1;
  wire s_dadda_pg_rca24_fa468_and1;
  wire s_dadda_pg_rca24_fa468_or0;
  wire s_dadda_pg_rca24_fa469_xor0;
  wire s_dadda_pg_rca24_fa469_and0;
  wire s_dadda_pg_rca24_fa469_xor1;
  wire s_dadda_pg_rca24_fa469_and1;
  wire s_dadda_pg_rca24_fa469_or0;
  wire s_dadda_pg_rca24_fa470_xor0;
  wire s_dadda_pg_rca24_fa470_and0;
  wire s_dadda_pg_rca24_fa470_xor1;
  wire s_dadda_pg_rca24_fa470_and1;
  wire s_dadda_pg_rca24_fa470_or0;
  wire s_dadda_pg_rca24_fa471_xor0;
  wire s_dadda_pg_rca24_fa471_and0;
  wire s_dadda_pg_rca24_fa471_xor1;
  wire s_dadda_pg_rca24_fa471_and1;
  wire s_dadda_pg_rca24_fa471_or0;
  wire s_dadda_pg_rca24_fa472_xor0;
  wire s_dadda_pg_rca24_fa472_and0;
  wire s_dadda_pg_rca24_fa472_xor1;
  wire s_dadda_pg_rca24_fa472_and1;
  wire s_dadda_pg_rca24_fa472_or0;
  wire s_dadda_pg_rca24_fa473_xor0;
  wire s_dadda_pg_rca24_fa473_and0;
  wire s_dadda_pg_rca24_fa473_xor1;
  wire s_dadda_pg_rca24_fa473_and1;
  wire s_dadda_pg_rca24_fa473_or0;
  wire s_dadda_pg_rca24_fa474_xor0;
  wire s_dadda_pg_rca24_fa474_and0;
  wire s_dadda_pg_rca24_fa474_xor1;
  wire s_dadda_pg_rca24_fa474_and1;
  wire s_dadda_pg_rca24_fa474_or0;
  wire s_dadda_pg_rca24_fa475_xor0;
  wire s_dadda_pg_rca24_fa475_and0;
  wire s_dadda_pg_rca24_fa475_xor1;
  wire s_dadda_pg_rca24_fa475_and1;
  wire s_dadda_pg_rca24_fa475_or0;
  wire s_dadda_pg_rca24_fa476_xor0;
  wire s_dadda_pg_rca24_fa476_and0;
  wire s_dadda_pg_rca24_fa476_xor1;
  wire s_dadda_pg_rca24_fa476_and1;
  wire s_dadda_pg_rca24_fa476_or0;
  wire s_dadda_pg_rca24_fa477_xor0;
  wire s_dadda_pg_rca24_fa477_and0;
  wire s_dadda_pg_rca24_fa477_xor1;
  wire s_dadda_pg_rca24_fa477_and1;
  wire s_dadda_pg_rca24_fa477_or0;
  wire s_dadda_pg_rca24_fa478_xor0;
  wire s_dadda_pg_rca24_fa478_and0;
  wire s_dadda_pg_rca24_fa478_xor1;
  wire s_dadda_pg_rca24_fa478_and1;
  wire s_dadda_pg_rca24_fa478_or0;
  wire s_dadda_pg_rca24_fa479_xor0;
  wire s_dadda_pg_rca24_fa479_and0;
  wire s_dadda_pg_rca24_fa479_xor1;
  wire s_dadda_pg_rca24_fa479_and1;
  wire s_dadda_pg_rca24_fa479_or0;
  wire s_dadda_pg_rca24_fa480_xor0;
  wire s_dadda_pg_rca24_fa480_and0;
  wire s_dadda_pg_rca24_fa480_xor1;
  wire s_dadda_pg_rca24_fa480_and1;
  wire s_dadda_pg_rca24_fa480_or0;
  wire s_dadda_pg_rca24_nand_20_23;
  wire s_dadda_pg_rca24_fa481_xor0;
  wire s_dadda_pg_rca24_fa481_and0;
  wire s_dadda_pg_rca24_fa481_xor1;
  wire s_dadda_pg_rca24_fa481_and1;
  wire s_dadda_pg_rca24_fa481_or0;
  wire s_dadda_pg_rca24_and_22_22;
  wire s_dadda_pg_rca24_nand_21_23;
  wire s_dadda_pg_rca24_fa482_xor0;
  wire s_dadda_pg_rca24_fa482_and0;
  wire s_dadda_pg_rca24_fa482_xor1;
  wire s_dadda_pg_rca24_fa482_and1;
  wire s_dadda_pg_rca24_fa482_or0;
  wire s_dadda_pg_rca24_nand_23_22;
  wire s_dadda_pg_rca24_fa483_xor0;
  wire s_dadda_pg_rca24_fa483_and0;
  wire s_dadda_pg_rca24_fa483_xor1;
  wire s_dadda_pg_rca24_fa483_and1;
  wire s_dadda_pg_rca24_fa483_or0;
  wire s_dadda_pg_rca24_and_0_0;
  wire s_dadda_pg_rca24_and_1_0;
  wire s_dadda_pg_rca24_and_0_2;
  wire s_dadda_pg_rca24_nand_22_23;
  wire s_dadda_pg_rca24_and_0_1;
  wire s_dadda_pg_rca24_and_23_23;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa0_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa0_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa1_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and1;
  wire s_dadda_pg_rca24_u_pg_rca46_or1;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa2_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and2;
  wire s_dadda_pg_rca24_u_pg_rca46_or2;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa3_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and3;
  wire s_dadda_pg_rca24_u_pg_rca46_or3;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa4_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and4;
  wire s_dadda_pg_rca24_u_pg_rca46_or4;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa5_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and5;
  wire s_dadda_pg_rca24_u_pg_rca46_or5;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa6_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and6;
  wire s_dadda_pg_rca24_u_pg_rca46_or6;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa7_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and7;
  wire s_dadda_pg_rca24_u_pg_rca46_or7;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa8_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and8;
  wire s_dadda_pg_rca24_u_pg_rca46_or8;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa9_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and9;
  wire s_dadda_pg_rca24_u_pg_rca46_or9;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa10_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and10;
  wire s_dadda_pg_rca24_u_pg_rca46_or10;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa11_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and11;
  wire s_dadda_pg_rca24_u_pg_rca46_or11;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa12_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and12;
  wire s_dadda_pg_rca24_u_pg_rca46_or12;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa13_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and13;
  wire s_dadda_pg_rca24_u_pg_rca46_or13;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa14_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and14;
  wire s_dadda_pg_rca24_u_pg_rca46_or14;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa15_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and15;
  wire s_dadda_pg_rca24_u_pg_rca46_or15;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa16_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and16;
  wire s_dadda_pg_rca24_u_pg_rca46_or16;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa17_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and17;
  wire s_dadda_pg_rca24_u_pg_rca46_or17;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa18_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and18;
  wire s_dadda_pg_rca24_u_pg_rca46_or18;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa19_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and19;
  wire s_dadda_pg_rca24_u_pg_rca46_or19;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa20_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and20;
  wire s_dadda_pg_rca24_u_pg_rca46_or20;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa21_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and21;
  wire s_dadda_pg_rca24_u_pg_rca46_or21;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa22_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and22;
  wire s_dadda_pg_rca24_u_pg_rca46_or22;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa23_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and23;
  wire s_dadda_pg_rca24_u_pg_rca46_or23;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa24_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and24;
  wire s_dadda_pg_rca24_u_pg_rca46_or24;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa25_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and25;
  wire s_dadda_pg_rca24_u_pg_rca46_or25;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa26_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and26;
  wire s_dadda_pg_rca24_u_pg_rca46_or26;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa27_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and27;
  wire s_dadda_pg_rca24_u_pg_rca46_or27;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa28_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and28;
  wire s_dadda_pg_rca24_u_pg_rca46_or28;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa29_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and29;
  wire s_dadda_pg_rca24_u_pg_rca46_or29;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa30_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and30;
  wire s_dadda_pg_rca24_u_pg_rca46_or30;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa31_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and31;
  wire s_dadda_pg_rca24_u_pg_rca46_or31;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa32_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and32;
  wire s_dadda_pg_rca24_u_pg_rca46_or32;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa33_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and33;
  wire s_dadda_pg_rca24_u_pg_rca46_or33;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa34_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and34;
  wire s_dadda_pg_rca24_u_pg_rca46_or34;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa35_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and35;
  wire s_dadda_pg_rca24_u_pg_rca46_or35;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa36_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and36;
  wire s_dadda_pg_rca24_u_pg_rca46_or36;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa37_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and37;
  wire s_dadda_pg_rca24_u_pg_rca46_or37;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa38_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and38;
  wire s_dadda_pg_rca24_u_pg_rca46_or38;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa39_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and39;
  wire s_dadda_pg_rca24_u_pg_rca46_or39;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa40_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and40;
  wire s_dadda_pg_rca24_u_pg_rca46_or40;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa41_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and41;
  wire s_dadda_pg_rca24_u_pg_rca46_or41;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa42_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and42;
  wire s_dadda_pg_rca24_u_pg_rca46_or42;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa43_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and43;
  wire s_dadda_pg_rca24_u_pg_rca46_or43;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa44_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and44;
  wire s_dadda_pg_rca24_u_pg_rca46_or44;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa45_and0;
  wire s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor1;
  wire s_dadda_pg_rca24_u_pg_rca46_and45;
  wire s_dadda_pg_rca24_u_pg_rca46_or45;
  wire s_dadda_pg_rca24_xor0;

  assign s_dadda_pg_rca24_and_19_0 = a[19] & b[0];
  assign s_dadda_pg_rca24_and_18_1 = a[18] & b[1];
  assign s_dadda_pg_rca24_ha0_xor0 = s_dadda_pg_rca24_and_19_0 ^ s_dadda_pg_rca24_and_18_1;
  assign s_dadda_pg_rca24_ha0_and0 = s_dadda_pg_rca24_and_19_0 & s_dadda_pg_rca24_and_18_1;
  assign s_dadda_pg_rca24_and_20_0 = a[20] & b[0];
  assign s_dadda_pg_rca24_and_19_1 = a[19] & b[1];
  assign s_dadda_pg_rca24_fa0_xor0 = s_dadda_pg_rca24_ha0_and0 ^ s_dadda_pg_rca24_and_20_0;
  assign s_dadda_pg_rca24_fa0_and0 = s_dadda_pg_rca24_ha0_and0 & s_dadda_pg_rca24_and_20_0;
  assign s_dadda_pg_rca24_fa0_xor1 = s_dadda_pg_rca24_fa0_xor0 ^ s_dadda_pg_rca24_and_19_1;
  assign s_dadda_pg_rca24_fa0_and1 = s_dadda_pg_rca24_fa0_xor0 & s_dadda_pg_rca24_and_19_1;
  assign s_dadda_pg_rca24_fa0_or0 = s_dadda_pg_rca24_fa0_and0 | s_dadda_pg_rca24_fa0_and1;
  assign s_dadda_pg_rca24_and_18_2 = a[18] & b[2];
  assign s_dadda_pg_rca24_and_17_3 = a[17] & b[3];
  assign s_dadda_pg_rca24_ha1_xor0 = s_dadda_pg_rca24_and_18_2 ^ s_dadda_pg_rca24_and_17_3;
  assign s_dadda_pg_rca24_ha1_and0 = s_dadda_pg_rca24_and_18_2 & s_dadda_pg_rca24_and_17_3;
  assign s_dadda_pg_rca24_and_21_0 = a[21] & b[0];
  assign s_dadda_pg_rca24_fa1_xor0 = s_dadda_pg_rca24_ha1_and0 ^ s_dadda_pg_rca24_fa0_or0;
  assign s_dadda_pg_rca24_fa1_and0 = s_dadda_pg_rca24_ha1_and0 & s_dadda_pg_rca24_fa0_or0;
  assign s_dadda_pg_rca24_fa1_xor1 = s_dadda_pg_rca24_fa1_xor0 ^ s_dadda_pg_rca24_and_21_0;
  assign s_dadda_pg_rca24_fa1_and1 = s_dadda_pg_rca24_fa1_xor0 & s_dadda_pg_rca24_and_21_0;
  assign s_dadda_pg_rca24_fa1_or0 = s_dadda_pg_rca24_fa1_and0 | s_dadda_pg_rca24_fa1_and1;
  assign s_dadda_pg_rca24_and_20_1 = a[20] & b[1];
  assign s_dadda_pg_rca24_and_19_2 = a[19] & b[2];
  assign s_dadda_pg_rca24_and_18_3 = a[18] & b[3];
  assign s_dadda_pg_rca24_fa2_xor0 = s_dadda_pg_rca24_and_20_1 ^ s_dadda_pg_rca24_and_19_2;
  assign s_dadda_pg_rca24_fa2_and0 = s_dadda_pg_rca24_and_20_1 & s_dadda_pg_rca24_and_19_2;
  assign s_dadda_pg_rca24_fa2_xor1 = s_dadda_pg_rca24_fa2_xor0 ^ s_dadda_pg_rca24_and_18_3;
  assign s_dadda_pg_rca24_fa2_and1 = s_dadda_pg_rca24_fa2_xor0 & s_dadda_pg_rca24_and_18_3;
  assign s_dadda_pg_rca24_fa2_or0 = s_dadda_pg_rca24_fa2_and0 | s_dadda_pg_rca24_fa2_and1;
  assign s_dadda_pg_rca24_and_17_4 = a[17] & b[4];
  assign s_dadda_pg_rca24_and_16_5 = a[16] & b[5];
  assign s_dadda_pg_rca24_ha2_xor0 = s_dadda_pg_rca24_and_17_4 ^ s_dadda_pg_rca24_and_16_5;
  assign s_dadda_pg_rca24_ha2_and0 = s_dadda_pg_rca24_and_17_4 & s_dadda_pg_rca24_and_16_5;
  assign s_dadda_pg_rca24_fa3_xor0 = s_dadda_pg_rca24_ha2_and0 ^ s_dadda_pg_rca24_fa2_or0;
  assign s_dadda_pg_rca24_fa3_and0 = s_dadda_pg_rca24_ha2_and0 & s_dadda_pg_rca24_fa2_or0;
  assign s_dadda_pg_rca24_fa3_xor1 = s_dadda_pg_rca24_fa3_xor0 ^ s_dadda_pg_rca24_fa1_or0;
  assign s_dadda_pg_rca24_fa3_and1 = s_dadda_pg_rca24_fa3_xor0 & s_dadda_pg_rca24_fa1_or0;
  assign s_dadda_pg_rca24_fa3_or0 = s_dadda_pg_rca24_fa3_and0 | s_dadda_pg_rca24_fa3_and1;
  assign s_dadda_pg_rca24_and_22_0 = a[22] & b[0];
  assign s_dadda_pg_rca24_and_21_1 = a[21] & b[1];
  assign s_dadda_pg_rca24_and_20_2 = a[20] & b[2];
  assign s_dadda_pg_rca24_fa4_xor0 = s_dadda_pg_rca24_and_22_0 ^ s_dadda_pg_rca24_and_21_1;
  assign s_dadda_pg_rca24_fa4_and0 = s_dadda_pg_rca24_and_22_0 & s_dadda_pg_rca24_and_21_1;
  assign s_dadda_pg_rca24_fa4_xor1 = s_dadda_pg_rca24_fa4_xor0 ^ s_dadda_pg_rca24_and_20_2;
  assign s_dadda_pg_rca24_fa4_and1 = s_dadda_pg_rca24_fa4_xor0 & s_dadda_pg_rca24_and_20_2;
  assign s_dadda_pg_rca24_fa4_or0 = s_dadda_pg_rca24_fa4_and0 | s_dadda_pg_rca24_fa4_and1;
  assign s_dadda_pg_rca24_and_19_3 = a[19] & b[3];
  assign s_dadda_pg_rca24_and_18_4 = a[18] & b[4];
  assign s_dadda_pg_rca24_and_17_5 = a[17] & b[5];
  assign s_dadda_pg_rca24_fa5_xor0 = s_dadda_pg_rca24_and_19_3 ^ s_dadda_pg_rca24_and_18_4;
  assign s_dadda_pg_rca24_fa5_and0 = s_dadda_pg_rca24_and_19_3 & s_dadda_pg_rca24_and_18_4;
  assign s_dadda_pg_rca24_fa5_xor1 = s_dadda_pg_rca24_fa5_xor0 ^ s_dadda_pg_rca24_and_17_5;
  assign s_dadda_pg_rca24_fa5_and1 = s_dadda_pg_rca24_fa5_xor0 & s_dadda_pg_rca24_and_17_5;
  assign s_dadda_pg_rca24_fa5_or0 = s_dadda_pg_rca24_fa5_and0 | s_dadda_pg_rca24_fa5_and1;
  assign s_dadda_pg_rca24_and_16_6 = a[16] & b[6];
  assign s_dadda_pg_rca24_and_15_7 = a[15] & b[7];
  assign s_dadda_pg_rca24_ha3_xor0 = s_dadda_pg_rca24_and_16_6 ^ s_dadda_pg_rca24_and_15_7;
  assign s_dadda_pg_rca24_ha3_and0 = s_dadda_pg_rca24_and_16_6 & s_dadda_pg_rca24_and_15_7;
  assign s_dadda_pg_rca24_fa6_xor0 = s_dadda_pg_rca24_ha3_and0 ^ s_dadda_pg_rca24_fa5_or0;
  assign s_dadda_pg_rca24_fa6_and0 = s_dadda_pg_rca24_ha3_and0 & s_dadda_pg_rca24_fa5_or0;
  assign s_dadda_pg_rca24_fa6_xor1 = s_dadda_pg_rca24_fa6_xor0 ^ s_dadda_pg_rca24_fa4_or0;
  assign s_dadda_pg_rca24_fa6_and1 = s_dadda_pg_rca24_fa6_xor0 & s_dadda_pg_rca24_fa4_or0;
  assign s_dadda_pg_rca24_fa6_or0 = s_dadda_pg_rca24_fa6_and0 | s_dadda_pg_rca24_fa6_and1;
  assign s_dadda_pg_rca24_nand_23_0 = ~(a[23] & b[0]);
  assign s_dadda_pg_rca24_and_22_1 = a[22] & b[1];
  assign s_dadda_pg_rca24_fa7_xor0 = s_dadda_pg_rca24_fa3_or0 ^ s_dadda_pg_rca24_nand_23_0;
  assign s_dadda_pg_rca24_fa7_and0 = s_dadda_pg_rca24_fa3_or0 & s_dadda_pg_rca24_nand_23_0;
  assign s_dadda_pg_rca24_fa7_xor1 = s_dadda_pg_rca24_fa7_xor0 ^ s_dadda_pg_rca24_and_22_1;
  assign s_dadda_pg_rca24_fa7_and1 = s_dadda_pg_rca24_fa7_xor0 & s_dadda_pg_rca24_and_22_1;
  assign s_dadda_pg_rca24_fa7_or0 = s_dadda_pg_rca24_fa7_and0 | s_dadda_pg_rca24_fa7_and1;
  assign s_dadda_pg_rca24_and_21_2 = a[21] & b[2];
  assign s_dadda_pg_rca24_and_20_3 = a[20] & b[3];
  assign s_dadda_pg_rca24_and_19_4 = a[19] & b[4];
  assign s_dadda_pg_rca24_fa8_xor0 = s_dadda_pg_rca24_and_21_2 ^ s_dadda_pg_rca24_and_20_3;
  assign s_dadda_pg_rca24_fa8_and0 = s_dadda_pg_rca24_and_21_2 & s_dadda_pg_rca24_and_20_3;
  assign s_dadda_pg_rca24_fa8_xor1 = s_dadda_pg_rca24_fa8_xor0 ^ s_dadda_pg_rca24_and_19_4;
  assign s_dadda_pg_rca24_fa8_and1 = s_dadda_pg_rca24_fa8_xor0 & s_dadda_pg_rca24_and_19_4;
  assign s_dadda_pg_rca24_fa8_or0 = s_dadda_pg_rca24_fa8_and0 | s_dadda_pg_rca24_fa8_and1;
  assign s_dadda_pg_rca24_and_18_5 = a[18] & b[5];
  assign s_dadda_pg_rca24_and_17_6 = a[17] & b[6];
  assign s_dadda_pg_rca24_and_16_7 = a[16] & b[7];
  assign s_dadda_pg_rca24_fa9_xor0 = s_dadda_pg_rca24_and_18_5 ^ s_dadda_pg_rca24_and_17_6;
  assign s_dadda_pg_rca24_fa9_and0 = s_dadda_pg_rca24_and_18_5 & s_dadda_pg_rca24_and_17_6;
  assign s_dadda_pg_rca24_fa9_xor1 = s_dadda_pg_rca24_fa9_xor0 ^ s_dadda_pg_rca24_and_16_7;
  assign s_dadda_pg_rca24_fa9_and1 = s_dadda_pg_rca24_fa9_xor0 & s_dadda_pg_rca24_and_16_7;
  assign s_dadda_pg_rca24_fa9_or0 = s_dadda_pg_rca24_fa9_and0 | s_dadda_pg_rca24_fa9_and1;
  assign s_dadda_pg_rca24_and_15_8 = a[15] & b[8];
  assign s_dadda_pg_rca24_and_14_9 = a[14] & b[9];
  assign s_dadda_pg_rca24_ha4_xor0 = s_dadda_pg_rca24_and_15_8 ^ s_dadda_pg_rca24_and_14_9;
  assign s_dadda_pg_rca24_ha4_and0 = s_dadda_pg_rca24_and_15_8 & s_dadda_pg_rca24_and_14_9;
  assign s_dadda_pg_rca24_fa10_xor0 = s_dadda_pg_rca24_ha4_and0 ^ s_dadda_pg_rca24_fa9_or0;
  assign s_dadda_pg_rca24_fa10_and0 = s_dadda_pg_rca24_ha4_and0 & s_dadda_pg_rca24_fa9_or0;
  assign s_dadda_pg_rca24_fa10_xor1 = s_dadda_pg_rca24_fa10_xor0 ^ s_dadda_pg_rca24_fa8_or0;
  assign s_dadda_pg_rca24_fa10_and1 = s_dadda_pg_rca24_fa10_xor0 & s_dadda_pg_rca24_fa8_or0;
  assign s_dadda_pg_rca24_fa10_or0 = s_dadda_pg_rca24_fa10_and0 | s_dadda_pg_rca24_fa10_and1;
  assign s_dadda_pg_rca24_fa11_xor0 = s_dadda_pg_rca24_fa7_or0 ^ s_dadda_pg_rca24_fa6_or0;
  assign s_dadda_pg_rca24_fa11_and0 = s_dadda_pg_rca24_fa7_or0 & s_dadda_pg_rca24_fa6_or0;
  assign s_dadda_pg_rca24_fa11_xor1 = ~s_dadda_pg_rca24_fa11_xor0;
  assign s_dadda_pg_rca24_fa11_or0 = s_dadda_pg_rca24_fa11_and0 | s_dadda_pg_rca24_fa11_xor0;
  assign s_dadda_pg_rca24_nand_23_1 = ~(a[23] & b[1]);
  assign s_dadda_pg_rca24_and_22_2 = a[22] & b[2];
  assign s_dadda_pg_rca24_and_21_3 = a[21] & b[3];
  assign s_dadda_pg_rca24_fa12_xor0 = s_dadda_pg_rca24_nand_23_1 ^ s_dadda_pg_rca24_and_22_2;
  assign s_dadda_pg_rca24_fa12_and0 = s_dadda_pg_rca24_nand_23_1 & s_dadda_pg_rca24_and_22_2;
  assign s_dadda_pg_rca24_fa12_xor1 = s_dadda_pg_rca24_fa12_xor0 ^ s_dadda_pg_rca24_and_21_3;
  assign s_dadda_pg_rca24_fa12_and1 = s_dadda_pg_rca24_fa12_xor0 & s_dadda_pg_rca24_and_21_3;
  assign s_dadda_pg_rca24_fa12_or0 = s_dadda_pg_rca24_fa12_and0 | s_dadda_pg_rca24_fa12_and1;
  assign s_dadda_pg_rca24_and_20_4 = a[20] & b[4];
  assign s_dadda_pg_rca24_and_19_5 = a[19] & b[5];
  assign s_dadda_pg_rca24_and_18_6 = a[18] & b[6];
  assign s_dadda_pg_rca24_fa13_xor0 = s_dadda_pg_rca24_and_20_4 ^ s_dadda_pg_rca24_and_19_5;
  assign s_dadda_pg_rca24_fa13_and0 = s_dadda_pg_rca24_and_20_4 & s_dadda_pg_rca24_and_19_5;
  assign s_dadda_pg_rca24_fa13_xor1 = s_dadda_pg_rca24_fa13_xor0 ^ s_dadda_pg_rca24_and_18_6;
  assign s_dadda_pg_rca24_fa13_and1 = s_dadda_pg_rca24_fa13_xor0 & s_dadda_pg_rca24_and_18_6;
  assign s_dadda_pg_rca24_fa13_or0 = s_dadda_pg_rca24_fa13_and0 | s_dadda_pg_rca24_fa13_and1;
  assign s_dadda_pg_rca24_and_17_7 = a[17] & b[7];
  assign s_dadda_pg_rca24_and_16_8 = a[16] & b[8];
  assign s_dadda_pg_rca24_and_15_9 = a[15] & b[9];
  assign s_dadda_pg_rca24_fa14_xor0 = s_dadda_pg_rca24_and_17_7 ^ s_dadda_pg_rca24_and_16_8;
  assign s_dadda_pg_rca24_fa14_and0 = s_dadda_pg_rca24_and_17_7 & s_dadda_pg_rca24_and_16_8;
  assign s_dadda_pg_rca24_fa14_xor1 = s_dadda_pg_rca24_fa14_xor0 ^ s_dadda_pg_rca24_and_15_9;
  assign s_dadda_pg_rca24_fa14_and1 = s_dadda_pg_rca24_fa14_xor0 & s_dadda_pg_rca24_and_15_9;
  assign s_dadda_pg_rca24_fa14_or0 = s_dadda_pg_rca24_fa14_and0 | s_dadda_pg_rca24_fa14_and1;
  assign s_dadda_pg_rca24_fa15_xor0 = s_dadda_pg_rca24_fa14_or0 ^ s_dadda_pg_rca24_fa13_or0;
  assign s_dadda_pg_rca24_fa15_and0 = s_dadda_pg_rca24_fa14_or0 & s_dadda_pg_rca24_fa13_or0;
  assign s_dadda_pg_rca24_fa15_xor1 = s_dadda_pg_rca24_fa15_xor0 ^ s_dadda_pg_rca24_fa12_or0;
  assign s_dadda_pg_rca24_fa15_and1 = s_dadda_pg_rca24_fa15_xor0 & s_dadda_pg_rca24_fa12_or0;
  assign s_dadda_pg_rca24_fa15_or0 = s_dadda_pg_rca24_fa15_and0 | s_dadda_pg_rca24_fa15_and1;
  assign s_dadda_pg_rca24_nand_23_2 = ~(a[23] & b[2]);
  assign s_dadda_pg_rca24_fa16_xor0 = s_dadda_pg_rca24_fa11_or0 ^ s_dadda_pg_rca24_fa10_or0;
  assign s_dadda_pg_rca24_fa16_and0 = s_dadda_pg_rca24_fa11_or0 & s_dadda_pg_rca24_fa10_or0;
  assign s_dadda_pg_rca24_fa16_xor1 = s_dadda_pg_rca24_fa16_xor0 ^ s_dadda_pg_rca24_nand_23_2;
  assign s_dadda_pg_rca24_fa16_and1 = s_dadda_pg_rca24_fa16_xor0 & s_dadda_pg_rca24_nand_23_2;
  assign s_dadda_pg_rca24_fa16_or0 = s_dadda_pg_rca24_fa16_and0 | s_dadda_pg_rca24_fa16_and1;
  assign s_dadda_pg_rca24_and_22_3 = a[22] & b[3];
  assign s_dadda_pg_rca24_and_21_4 = a[21] & b[4];
  assign s_dadda_pg_rca24_and_20_5 = a[20] & b[5];
  assign s_dadda_pg_rca24_fa17_xor0 = s_dadda_pg_rca24_and_22_3 ^ s_dadda_pg_rca24_and_21_4;
  assign s_dadda_pg_rca24_fa17_and0 = s_dadda_pg_rca24_and_22_3 & s_dadda_pg_rca24_and_21_4;
  assign s_dadda_pg_rca24_fa17_xor1 = s_dadda_pg_rca24_fa17_xor0 ^ s_dadda_pg_rca24_and_20_5;
  assign s_dadda_pg_rca24_fa17_and1 = s_dadda_pg_rca24_fa17_xor0 & s_dadda_pg_rca24_and_20_5;
  assign s_dadda_pg_rca24_fa17_or0 = s_dadda_pg_rca24_fa17_and0 | s_dadda_pg_rca24_fa17_and1;
  assign s_dadda_pg_rca24_and_19_6 = a[19] & b[6];
  assign s_dadda_pg_rca24_and_18_7 = a[18] & b[7];
  assign s_dadda_pg_rca24_and_17_8 = a[17] & b[8];
  assign s_dadda_pg_rca24_fa18_xor0 = s_dadda_pg_rca24_and_19_6 ^ s_dadda_pg_rca24_and_18_7;
  assign s_dadda_pg_rca24_fa18_and0 = s_dadda_pg_rca24_and_19_6 & s_dadda_pg_rca24_and_18_7;
  assign s_dadda_pg_rca24_fa18_xor1 = s_dadda_pg_rca24_fa18_xor0 ^ s_dadda_pg_rca24_and_17_8;
  assign s_dadda_pg_rca24_fa18_and1 = s_dadda_pg_rca24_fa18_xor0 & s_dadda_pg_rca24_and_17_8;
  assign s_dadda_pg_rca24_fa18_or0 = s_dadda_pg_rca24_fa18_and0 | s_dadda_pg_rca24_fa18_and1;
  assign s_dadda_pg_rca24_fa19_xor0 = s_dadda_pg_rca24_fa18_or0 ^ s_dadda_pg_rca24_fa17_or0;
  assign s_dadda_pg_rca24_fa19_and0 = s_dadda_pg_rca24_fa18_or0 & s_dadda_pg_rca24_fa17_or0;
  assign s_dadda_pg_rca24_fa19_xor1 = s_dadda_pg_rca24_fa19_xor0 ^ s_dadda_pg_rca24_fa16_or0;
  assign s_dadda_pg_rca24_fa19_and1 = s_dadda_pg_rca24_fa19_xor0 & s_dadda_pg_rca24_fa16_or0;
  assign s_dadda_pg_rca24_fa19_or0 = s_dadda_pg_rca24_fa19_and0 | s_dadda_pg_rca24_fa19_and1;
  assign s_dadda_pg_rca24_nand_23_3 = ~(a[23] & b[3]);
  assign s_dadda_pg_rca24_and_22_4 = a[22] & b[4];
  assign s_dadda_pg_rca24_fa20_xor0 = s_dadda_pg_rca24_fa15_or0 ^ s_dadda_pg_rca24_nand_23_3;
  assign s_dadda_pg_rca24_fa20_and0 = s_dadda_pg_rca24_fa15_or0 & s_dadda_pg_rca24_nand_23_3;
  assign s_dadda_pg_rca24_fa20_xor1 = s_dadda_pg_rca24_fa20_xor0 ^ s_dadda_pg_rca24_and_22_4;
  assign s_dadda_pg_rca24_fa20_and1 = s_dadda_pg_rca24_fa20_xor0 & s_dadda_pg_rca24_and_22_4;
  assign s_dadda_pg_rca24_fa20_or0 = s_dadda_pg_rca24_fa20_and0 | s_dadda_pg_rca24_fa20_and1;
  assign s_dadda_pg_rca24_and_21_5 = a[21] & b[5];
  assign s_dadda_pg_rca24_and_20_6 = a[20] & b[6];
  assign s_dadda_pg_rca24_and_19_7 = a[19] & b[7];
  assign s_dadda_pg_rca24_fa21_xor0 = s_dadda_pg_rca24_and_21_5 ^ s_dadda_pg_rca24_and_20_6;
  assign s_dadda_pg_rca24_fa21_and0 = s_dadda_pg_rca24_and_21_5 & s_dadda_pg_rca24_and_20_6;
  assign s_dadda_pg_rca24_fa21_xor1 = s_dadda_pg_rca24_fa21_xor0 ^ s_dadda_pg_rca24_and_19_7;
  assign s_dadda_pg_rca24_fa21_and1 = s_dadda_pg_rca24_fa21_xor0 & s_dadda_pg_rca24_and_19_7;
  assign s_dadda_pg_rca24_fa21_or0 = s_dadda_pg_rca24_fa21_and0 | s_dadda_pg_rca24_fa21_and1;
  assign s_dadda_pg_rca24_fa22_xor0 = s_dadda_pg_rca24_fa21_or0 ^ s_dadda_pg_rca24_fa20_or0;
  assign s_dadda_pg_rca24_fa22_and0 = s_dadda_pg_rca24_fa21_or0 & s_dadda_pg_rca24_fa20_or0;
  assign s_dadda_pg_rca24_fa22_xor1 = s_dadda_pg_rca24_fa22_xor0 ^ s_dadda_pg_rca24_fa19_or0;
  assign s_dadda_pg_rca24_fa22_and1 = s_dadda_pg_rca24_fa22_xor0 & s_dadda_pg_rca24_fa19_or0;
  assign s_dadda_pg_rca24_fa22_or0 = s_dadda_pg_rca24_fa22_and0 | s_dadda_pg_rca24_fa22_and1;
  assign s_dadda_pg_rca24_nand_23_4 = ~(a[23] & b[4]);
  assign s_dadda_pg_rca24_and_22_5 = a[22] & b[5];
  assign s_dadda_pg_rca24_and_21_6 = a[21] & b[6];
  assign s_dadda_pg_rca24_fa23_xor0 = s_dadda_pg_rca24_nand_23_4 ^ s_dadda_pg_rca24_and_22_5;
  assign s_dadda_pg_rca24_fa23_and0 = s_dadda_pg_rca24_nand_23_4 & s_dadda_pg_rca24_and_22_5;
  assign s_dadda_pg_rca24_fa23_xor1 = s_dadda_pg_rca24_fa23_xor0 ^ s_dadda_pg_rca24_and_21_6;
  assign s_dadda_pg_rca24_fa23_and1 = s_dadda_pg_rca24_fa23_xor0 & s_dadda_pg_rca24_and_21_6;
  assign s_dadda_pg_rca24_fa23_or0 = s_dadda_pg_rca24_fa23_and0 | s_dadda_pg_rca24_fa23_and1;
  assign s_dadda_pg_rca24_nand_23_5 = ~(a[23] & b[5]);
  assign s_dadda_pg_rca24_fa24_xor0 = s_dadda_pg_rca24_fa23_or0 ^ s_dadda_pg_rca24_fa22_or0;
  assign s_dadda_pg_rca24_fa24_and0 = s_dadda_pg_rca24_fa23_or0 & s_dadda_pg_rca24_fa22_or0;
  assign s_dadda_pg_rca24_fa24_xor1 = s_dadda_pg_rca24_fa24_xor0 ^ s_dadda_pg_rca24_nand_23_5;
  assign s_dadda_pg_rca24_fa24_and1 = s_dadda_pg_rca24_fa24_xor0 & s_dadda_pg_rca24_nand_23_5;
  assign s_dadda_pg_rca24_fa24_or0 = s_dadda_pg_rca24_fa24_and0 | s_dadda_pg_rca24_fa24_and1;
  assign s_dadda_pg_rca24_and_6_0 = a[6] & b[0];
  assign s_dadda_pg_rca24_and_5_1 = a[5] & b[1];
  assign s_dadda_pg_rca24_ha5_xor0 = s_dadda_pg_rca24_and_6_0 ^ s_dadda_pg_rca24_and_5_1;
  assign s_dadda_pg_rca24_ha5_and0 = s_dadda_pg_rca24_and_6_0 & s_dadda_pg_rca24_and_5_1;
  assign s_dadda_pg_rca24_and_7_0 = a[7] & b[0];
  assign s_dadda_pg_rca24_and_6_1 = a[6] & b[1];
  assign s_dadda_pg_rca24_fa25_xor0 = s_dadda_pg_rca24_ha5_and0 ^ s_dadda_pg_rca24_and_7_0;
  assign s_dadda_pg_rca24_fa25_and0 = s_dadda_pg_rca24_ha5_and0 & s_dadda_pg_rca24_and_7_0;
  assign s_dadda_pg_rca24_fa25_xor1 = s_dadda_pg_rca24_fa25_xor0 ^ s_dadda_pg_rca24_and_6_1;
  assign s_dadda_pg_rca24_fa25_and1 = s_dadda_pg_rca24_fa25_xor0 & s_dadda_pg_rca24_and_6_1;
  assign s_dadda_pg_rca24_fa25_or0 = s_dadda_pg_rca24_fa25_and0 | s_dadda_pg_rca24_fa25_and1;
  assign s_dadda_pg_rca24_and_5_2 = a[5] & b[2];
  assign s_dadda_pg_rca24_and_4_3 = a[4] & b[3];
  assign s_dadda_pg_rca24_ha6_xor0 = s_dadda_pg_rca24_and_5_2 ^ s_dadda_pg_rca24_and_4_3;
  assign s_dadda_pg_rca24_ha6_and0 = s_dadda_pg_rca24_and_5_2 & s_dadda_pg_rca24_and_4_3;
  assign s_dadda_pg_rca24_and_8_0 = a[8] & b[0];
  assign s_dadda_pg_rca24_fa26_xor0 = s_dadda_pg_rca24_ha6_and0 ^ s_dadda_pg_rca24_fa25_or0;
  assign s_dadda_pg_rca24_fa26_and0 = s_dadda_pg_rca24_ha6_and0 & s_dadda_pg_rca24_fa25_or0;
  assign s_dadda_pg_rca24_fa26_xor1 = s_dadda_pg_rca24_fa26_xor0 ^ s_dadda_pg_rca24_and_8_0;
  assign s_dadda_pg_rca24_fa26_and1 = s_dadda_pg_rca24_fa26_xor0 & s_dadda_pg_rca24_and_8_0;
  assign s_dadda_pg_rca24_fa26_or0 = s_dadda_pg_rca24_fa26_and0 | s_dadda_pg_rca24_fa26_and1;
  assign s_dadda_pg_rca24_and_7_1 = a[7] & b[1];
  assign s_dadda_pg_rca24_and_6_2 = a[6] & b[2];
  assign s_dadda_pg_rca24_and_5_3 = a[5] & b[3];
  assign s_dadda_pg_rca24_fa27_xor0 = s_dadda_pg_rca24_and_7_1 ^ s_dadda_pg_rca24_and_6_2;
  assign s_dadda_pg_rca24_fa27_and0 = s_dadda_pg_rca24_and_7_1 & s_dadda_pg_rca24_and_6_2;
  assign s_dadda_pg_rca24_fa27_xor1 = s_dadda_pg_rca24_fa27_xor0 ^ s_dadda_pg_rca24_and_5_3;
  assign s_dadda_pg_rca24_fa27_and1 = s_dadda_pg_rca24_fa27_xor0 & s_dadda_pg_rca24_and_5_3;
  assign s_dadda_pg_rca24_fa27_or0 = s_dadda_pg_rca24_fa27_and0 | s_dadda_pg_rca24_fa27_and1;
  assign s_dadda_pg_rca24_and_4_4 = a[4] & b[4];
  assign s_dadda_pg_rca24_and_3_5 = a[3] & b[5];
  assign s_dadda_pg_rca24_ha7_xor0 = s_dadda_pg_rca24_and_4_4 ^ s_dadda_pg_rca24_and_3_5;
  assign s_dadda_pg_rca24_ha7_and0 = s_dadda_pg_rca24_and_4_4 & s_dadda_pg_rca24_and_3_5;
  assign s_dadda_pg_rca24_fa28_xor0 = s_dadda_pg_rca24_ha7_and0 ^ s_dadda_pg_rca24_fa27_or0;
  assign s_dadda_pg_rca24_fa28_and0 = s_dadda_pg_rca24_ha7_and0 & s_dadda_pg_rca24_fa27_or0;
  assign s_dadda_pg_rca24_fa28_xor1 = s_dadda_pg_rca24_fa28_xor0 ^ s_dadda_pg_rca24_fa26_or0;
  assign s_dadda_pg_rca24_fa28_and1 = s_dadda_pg_rca24_fa28_xor0 & s_dadda_pg_rca24_fa26_or0;
  assign s_dadda_pg_rca24_fa28_or0 = s_dadda_pg_rca24_fa28_and0 | s_dadda_pg_rca24_fa28_and1;
  assign s_dadda_pg_rca24_and_9_0 = a[9] & b[0];
  assign s_dadda_pg_rca24_and_8_1 = a[8] & b[1];
  assign s_dadda_pg_rca24_and_7_2 = a[7] & b[2];
  assign s_dadda_pg_rca24_fa29_xor0 = s_dadda_pg_rca24_and_9_0 ^ s_dadda_pg_rca24_and_8_1;
  assign s_dadda_pg_rca24_fa29_and0 = s_dadda_pg_rca24_and_9_0 & s_dadda_pg_rca24_and_8_1;
  assign s_dadda_pg_rca24_fa29_xor1 = s_dadda_pg_rca24_fa29_xor0 ^ s_dadda_pg_rca24_and_7_2;
  assign s_dadda_pg_rca24_fa29_and1 = s_dadda_pg_rca24_fa29_xor0 & s_dadda_pg_rca24_and_7_2;
  assign s_dadda_pg_rca24_fa29_or0 = s_dadda_pg_rca24_fa29_and0 | s_dadda_pg_rca24_fa29_and1;
  assign s_dadda_pg_rca24_and_6_3 = a[6] & b[3];
  assign s_dadda_pg_rca24_and_5_4 = a[5] & b[4];
  assign s_dadda_pg_rca24_and_4_5 = a[4] & b[5];
  assign s_dadda_pg_rca24_fa30_xor0 = s_dadda_pg_rca24_and_6_3 ^ s_dadda_pg_rca24_and_5_4;
  assign s_dadda_pg_rca24_fa30_and0 = s_dadda_pg_rca24_and_6_3 & s_dadda_pg_rca24_and_5_4;
  assign s_dadda_pg_rca24_fa30_xor1 = s_dadda_pg_rca24_fa30_xor0 ^ s_dadda_pg_rca24_and_4_5;
  assign s_dadda_pg_rca24_fa30_and1 = s_dadda_pg_rca24_fa30_xor0 & s_dadda_pg_rca24_and_4_5;
  assign s_dadda_pg_rca24_fa30_or0 = s_dadda_pg_rca24_fa30_and0 | s_dadda_pg_rca24_fa30_and1;
  assign s_dadda_pg_rca24_and_3_6 = a[3] & b[6];
  assign s_dadda_pg_rca24_and_2_7 = a[2] & b[7];
  assign s_dadda_pg_rca24_ha8_xor0 = s_dadda_pg_rca24_and_3_6 ^ s_dadda_pg_rca24_and_2_7;
  assign s_dadda_pg_rca24_ha8_and0 = s_dadda_pg_rca24_and_3_6 & s_dadda_pg_rca24_and_2_7;
  assign s_dadda_pg_rca24_fa31_xor0 = s_dadda_pg_rca24_ha8_and0 ^ s_dadda_pg_rca24_fa30_or0;
  assign s_dadda_pg_rca24_fa31_and0 = s_dadda_pg_rca24_ha8_and0 & s_dadda_pg_rca24_fa30_or0;
  assign s_dadda_pg_rca24_fa31_xor1 = s_dadda_pg_rca24_fa31_xor0 ^ s_dadda_pg_rca24_fa29_or0;
  assign s_dadda_pg_rca24_fa31_and1 = s_dadda_pg_rca24_fa31_xor0 & s_dadda_pg_rca24_fa29_or0;
  assign s_dadda_pg_rca24_fa31_or0 = s_dadda_pg_rca24_fa31_and0 | s_dadda_pg_rca24_fa31_and1;
  assign s_dadda_pg_rca24_and_10_0 = a[10] & b[0];
  assign s_dadda_pg_rca24_and_9_1 = a[9] & b[1];
  assign s_dadda_pg_rca24_fa32_xor0 = s_dadda_pg_rca24_fa28_or0 ^ s_dadda_pg_rca24_and_10_0;
  assign s_dadda_pg_rca24_fa32_and0 = s_dadda_pg_rca24_fa28_or0 & s_dadda_pg_rca24_and_10_0;
  assign s_dadda_pg_rca24_fa32_xor1 = s_dadda_pg_rca24_fa32_xor0 ^ s_dadda_pg_rca24_and_9_1;
  assign s_dadda_pg_rca24_fa32_and1 = s_dadda_pg_rca24_fa32_xor0 & s_dadda_pg_rca24_and_9_1;
  assign s_dadda_pg_rca24_fa32_or0 = s_dadda_pg_rca24_fa32_and0 | s_dadda_pg_rca24_fa32_and1;
  assign s_dadda_pg_rca24_and_8_2 = a[8] & b[2];
  assign s_dadda_pg_rca24_and_7_3 = a[7] & b[3];
  assign s_dadda_pg_rca24_and_6_4 = a[6] & b[4];
  assign s_dadda_pg_rca24_fa33_xor0 = s_dadda_pg_rca24_and_8_2 ^ s_dadda_pg_rca24_and_7_3;
  assign s_dadda_pg_rca24_fa33_and0 = s_dadda_pg_rca24_and_8_2 & s_dadda_pg_rca24_and_7_3;
  assign s_dadda_pg_rca24_fa33_xor1 = s_dadda_pg_rca24_fa33_xor0 ^ s_dadda_pg_rca24_and_6_4;
  assign s_dadda_pg_rca24_fa33_and1 = s_dadda_pg_rca24_fa33_xor0 & s_dadda_pg_rca24_and_6_4;
  assign s_dadda_pg_rca24_fa33_or0 = s_dadda_pg_rca24_fa33_and0 | s_dadda_pg_rca24_fa33_and1;
  assign s_dadda_pg_rca24_and_5_5 = a[5] & b[5];
  assign s_dadda_pg_rca24_and_4_6 = a[4] & b[6];
  assign s_dadda_pg_rca24_and_3_7 = a[3] & b[7];
  assign s_dadda_pg_rca24_fa34_xor0 = s_dadda_pg_rca24_and_5_5 ^ s_dadda_pg_rca24_and_4_6;
  assign s_dadda_pg_rca24_fa34_and0 = s_dadda_pg_rca24_and_5_5 & s_dadda_pg_rca24_and_4_6;
  assign s_dadda_pg_rca24_fa34_xor1 = s_dadda_pg_rca24_fa34_xor0 ^ s_dadda_pg_rca24_and_3_7;
  assign s_dadda_pg_rca24_fa34_and1 = s_dadda_pg_rca24_fa34_xor0 & s_dadda_pg_rca24_and_3_7;
  assign s_dadda_pg_rca24_fa34_or0 = s_dadda_pg_rca24_fa34_and0 | s_dadda_pg_rca24_fa34_and1;
  assign s_dadda_pg_rca24_and_2_8 = a[2] & b[8];
  assign s_dadda_pg_rca24_and_1_9 = a[1] & b[9];
  assign s_dadda_pg_rca24_ha9_xor0 = s_dadda_pg_rca24_and_2_8 ^ s_dadda_pg_rca24_and_1_9;
  assign s_dadda_pg_rca24_ha9_and0 = s_dadda_pg_rca24_and_2_8 & s_dadda_pg_rca24_and_1_9;
  assign s_dadda_pg_rca24_fa35_xor0 = s_dadda_pg_rca24_ha9_and0 ^ s_dadda_pg_rca24_fa34_or0;
  assign s_dadda_pg_rca24_fa35_and0 = s_dadda_pg_rca24_ha9_and0 & s_dadda_pg_rca24_fa34_or0;
  assign s_dadda_pg_rca24_fa35_xor1 = s_dadda_pg_rca24_fa35_xor0 ^ s_dadda_pg_rca24_fa33_or0;
  assign s_dadda_pg_rca24_fa35_and1 = s_dadda_pg_rca24_fa35_xor0 & s_dadda_pg_rca24_fa33_or0;
  assign s_dadda_pg_rca24_fa35_or0 = s_dadda_pg_rca24_fa35_and0 | s_dadda_pg_rca24_fa35_and1;
  assign s_dadda_pg_rca24_and_11_0 = a[11] & b[0];
  assign s_dadda_pg_rca24_fa36_xor0 = s_dadda_pg_rca24_fa32_or0 ^ s_dadda_pg_rca24_fa31_or0;
  assign s_dadda_pg_rca24_fa36_and0 = s_dadda_pg_rca24_fa32_or0 & s_dadda_pg_rca24_fa31_or0;
  assign s_dadda_pg_rca24_fa36_xor1 = s_dadda_pg_rca24_fa36_xor0 ^ s_dadda_pg_rca24_and_11_0;
  assign s_dadda_pg_rca24_fa36_and1 = s_dadda_pg_rca24_fa36_xor0 & s_dadda_pg_rca24_and_11_0;
  assign s_dadda_pg_rca24_fa36_or0 = s_dadda_pg_rca24_fa36_and0 | s_dadda_pg_rca24_fa36_and1;
  assign s_dadda_pg_rca24_and_10_1 = a[10] & b[1];
  assign s_dadda_pg_rca24_and_9_2 = a[9] & b[2];
  assign s_dadda_pg_rca24_and_8_3 = a[8] & b[3];
  assign s_dadda_pg_rca24_fa37_xor0 = s_dadda_pg_rca24_and_10_1 ^ s_dadda_pg_rca24_and_9_2;
  assign s_dadda_pg_rca24_fa37_and0 = s_dadda_pg_rca24_and_10_1 & s_dadda_pg_rca24_and_9_2;
  assign s_dadda_pg_rca24_fa37_xor1 = s_dadda_pg_rca24_fa37_xor0 ^ s_dadda_pg_rca24_and_8_3;
  assign s_dadda_pg_rca24_fa37_and1 = s_dadda_pg_rca24_fa37_xor0 & s_dadda_pg_rca24_and_8_3;
  assign s_dadda_pg_rca24_fa37_or0 = s_dadda_pg_rca24_fa37_and0 | s_dadda_pg_rca24_fa37_and1;
  assign s_dadda_pg_rca24_and_7_4 = a[7] & b[4];
  assign s_dadda_pg_rca24_and_6_5 = a[6] & b[5];
  assign s_dadda_pg_rca24_and_5_6 = a[5] & b[6];
  assign s_dadda_pg_rca24_fa38_xor0 = s_dadda_pg_rca24_and_7_4 ^ s_dadda_pg_rca24_and_6_5;
  assign s_dadda_pg_rca24_fa38_and0 = s_dadda_pg_rca24_and_7_4 & s_dadda_pg_rca24_and_6_5;
  assign s_dadda_pg_rca24_fa38_xor1 = s_dadda_pg_rca24_fa38_xor0 ^ s_dadda_pg_rca24_and_5_6;
  assign s_dadda_pg_rca24_fa38_and1 = s_dadda_pg_rca24_fa38_xor0 & s_dadda_pg_rca24_and_5_6;
  assign s_dadda_pg_rca24_fa38_or0 = s_dadda_pg_rca24_fa38_and0 | s_dadda_pg_rca24_fa38_and1;
  assign s_dadda_pg_rca24_and_4_7 = a[4] & b[7];
  assign s_dadda_pg_rca24_and_3_8 = a[3] & b[8];
  assign s_dadda_pg_rca24_and_2_9 = a[2] & b[9];
  assign s_dadda_pg_rca24_fa39_xor0 = s_dadda_pg_rca24_and_4_7 ^ s_dadda_pg_rca24_and_3_8;
  assign s_dadda_pg_rca24_fa39_and0 = s_dadda_pg_rca24_and_4_7 & s_dadda_pg_rca24_and_3_8;
  assign s_dadda_pg_rca24_fa39_xor1 = s_dadda_pg_rca24_fa39_xor0 ^ s_dadda_pg_rca24_and_2_9;
  assign s_dadda_pg_rca24_fa39_and1 = s_dadda_pg_rca24_fa39_xor0 & s_dadda_pg_rca24_and_2_9;
  assign s_dadda_pg_rca24_fa39_or0 = s_dadda_pg_rca24_fa39_and0 | s_dadda_pg_rca24_fa39_and1;
  assign s_dadda_pg_rca24_and_1_10 = a[1] & b[10];
  assign s_dadda_pg_rca24_and_0_11 = a[0] & b[11];
  assign s_dadda_pg_rca24_ha10_xor0 = s_dadda_pg_rca24_and_1_10 ^ s_dadda_pg_rca24_and_0_11;
  assign s_dadda_pg_rca24_ha10_and0 = s_dadda_pg_rca24_and_1_10 & s_dadda_pg_rca24_and_0_11;
  assign s_dadda_pg_rca24_fa40_xor0 = s_dadda_pg_rca24_ha10_and0 ^ s_dadda_pg_rca24_fa39_or0;
  assign s_dadda_pg_rca24_fa40_and0 = s_dadda_pg_rca24_ha10_and0 & s_dadda_pg_rca24_fa39_or0;
  assign s_dadda_pg_rca24_fa40_xor1 = s_dadda_pg_rca24_fa40_xor0 ^ s_dadda_pg_rca24_fa38_or0;
  assign s_dadda_pg_rca24_fa40_and1 = s_dadda_pg_rca24_fa40_xor0 & s_dadda_pg_rca24_fa38_or0;
  assign s_dadda_pg_rca24_fa40_or0 = s_dadda_pg_rca24_fa40_and0 | s_dadda_pg_rca24_fa40_and1;
  assign s_dadda_pg_rca24_fa41_xor0 = s_dadda_pg_rca24_fa37_or0 ^ s_dadda_pg_rca24_fa36_or0;
  assign s_dadda_pg_rca24_fa41_and0 = s_dadda_pg_rca24_fa37_or0 & s_dadda_pg_rca24_fa36_or0;
  assign s_dadda_pg_rca24_fa41_xor1 = s_dadda_pg_rca24_fa41_xor0 ^ s_dadda_pg_rca24_fa35_or0;
  assign s_dadda_pg_rca24_fa41_and1 = s_dadda_pg_rca24_fa41_xor0 & s_dadda_pg_rca24_fa35_or0;
  assign s_dadda_pg_rca24_fa41_or0 = s_dadda_pg_rca24_fa41_and0 | s_dadda_pg_rca24_fa41_and1;
  assign s_dadda_pg_rca24_and_12_0 = a[12] & b[0];
  assign s_dadda_pg_rca24_and_11_1 = a[11] & b[1];
  assign s_dadda_pg_rca24_and_10_2 = a[10] & b[2];
  assign s_dadda_pg_rca24_fa42_xor0 = s_dadda_pg_rca24_and_12_0 ^ s_dadda_pg_rca24_and_11_1;
  assign s_dadda_pg_rca24_fa42_and0 = s_dadda_pg_rca24_and_12_0 & s_dadda_pg_rca24_and_11_1;
  assign s_dadda_pg_rca24_fa42_xor1 = s_dadda_pg_rca24_fa42_xor0 ^ s_dadda_pg_rca24_and_10_2;
  assign s_dadda_pg_rca24_fa42_and1 = s_dadda_pg_rca24_fa42_xor0 & s_dadda_pg_rca24_and_10_2;
  assign s_dadda_pg_rca24_fa42_or0 = s_dadda_pg_rca24_fa42_and0 | s_dadda_pg_rca24_fa42_and1;
  assign s_dadda_pg_rca24_and_9_3 = a[9] & b[3];
  assign s_dadda_pg_rca24_and_8_4 = a[8] & b[4];
  assign s_dadda_pg_rca24_and_7_5 = a[7] & b[5];
  assign s_dadda_pg_rca24_fa43_xor0 = s_dadda_pg_rca24_and_9_3 ^ s_dadda_pg_rca24_and_8_4;
  assign s_dadda_pg_rca24_fa43_and0 = s_dadda_pg_rca24_and_9_3 & s_dadda_pg_rca24_and_8_4;
  assign s_dadda_pg_rca24_fa43_xor1 = s_dadda_pg_rca24_fa43_xor0 ^ s_dadda_pg_rca24_and_7_5;
  assign s_dadda_pg_rca24_fa43_and1 = s_dadda_pg_rca24_fa43_xor0 & s_dadda_pg_rca24_and_7_5;
  assign s_dadda_pg_rca24_fa43_or0 = s_dadda_pg_rca24_fa43_and0 | s_dadda_pg_rca24_fa43_and1;
  assign s_dadda_pg_rca24_and_6_6 = a[6] & b[6];
  assign s_dadda_pg_rca24_and_5_7 = a[5] & b[7];
  assign s_dadda_pg_rca24_and_4_8 = a[4] & b[8];
  assign s_dadda_pg_rca24_fa44_xor0 = s_dadda_pg_rca24_and_6_6 ^ s_dadda_pg_rca24_and_5_7;
  assign s_dadda_pg_rca24_fa44_and0 = s_dadda_pg_rca24_and_6_6 & s_dadda_pg_rca24_and_5_7;
  assign s_dadda_pg_rca24_fa44_xor1 = s_dadda_pg_rca24_fa44_xor0 ^ s_dadda_pg_rca24_and_4_8;
  assign s_dadda_pg_rca24_fa44_and1 = s_dadda_pg_rca24_fa44_xor0 & s_dadda_pg_rca24_and_4_8;
  assign s_dadda_pg_rca24_fa44_or0 = s_dadda_pg_rca24_fa44_and0 | s_dadda_pg_rca24_fa44_and1;
  assign s_dadda_pg_rca24_and_3_9 = a[3] & b[9];
  assign s_dadda_pg_rca24_and_2_10 = a[2] & b[10];
  assign s_dadda_pg_rca24_and_1_11 = a[1] & b[11];
  assign s_dadda_pg_rca24_fa45_xor0 = s_dadda_pg_rca24_and_3_9 ^ s_dadda_pg_rca24_and_2_10;
  assign s_dadda_pg_rca24_fa45_and0 = s_dadda_pg_rca24_and_3_9 & s_dadda_pg_rca24_and_2_10;
  assign s_dadda_pg_rca24_fa45_xor1 = s_dadda_pg_rca24_fa45_xor0 ^ s_dadda_pg_rca24_and_1_11;
  assign s_dadda_pg_rca24_fa45_and1 = s_dadda_pg_rca24_fa45_xor0 & s_dadda_pg_rca24_and_1_11;
  assign s_dadda_pg_rca24_fa45_or0 = s_dadda_pg_rca24_fa45_and0 | s_dadda_pg_rca24_fa45_and1;
  assign s_dadda_pg_rca24_and_0_12 = a[0] & b[12];
  assign s_dadda_pg_rca24_ha11_xor0 = s_dadda_pg_rca24_and_0_12 ^ s_dadda_pg_rca24_fa40_xor1;
  assign s_dadda_pg_rca24_ha11_and0 = s_dadda_pg_rca24_and_0_12 & s_dadda_pg_rca24_fa40_xor1;
  assign s_dadda_pg_rca24_fa46_xor0 = s_dadda_pg_rca24_ha11_and0 ^ s_dadda_pg_rca24_fa45_or0;
  assign s_dadda_pg_rca24_fa46_and0 = s_dadda_pg_rca24_ha11_and0 & s_dadda_pg_rca24_fa45_or0;
  assign s_dadda_pg_rca24_fa46_xor1 = s_dadda_pg_rca24_fa46_xor0 ^ s_dadda_pg_rca24_fa44_or0;
  assign s_dadda_pg_rca24_fa46_and1 = s_dadda_pg_rca24_fa46_xor0 & s_dadda_pg_rca24_fa44_or0;
  assign s_dadda_pg_rca24_fa46_or0 = s_dadda_pg_rca24_fa46_and0 | s_dadda_pg_rca24_fa46_and1;
  assign s_dadda_pg_rca24_fa47_xor0 = s_dadda_pg_rca24_fa43_or0 ^ s_dadda_pg_rca24_fa42_or0;
  assign s_dadda_pg_rca24_fa47_and0 = s_dadda_pg_rca24_fa43_or0 & s_dadda_pg_rca24_fa42_or0;
  assign s_dadda_pg_rca24_fa47_xor1 = s_dadda_pg_rca24_fa47_xor0 ^ s_dadda_pg_rca24_fa41_or0;
  assign s_dadda_pg_rca24_fa47_and1 = s_dadda_pg_rca24_fa47_xor0 & s_dadda_pg_rca24_fa41_or0;
  assign s_dadda_pg_rca24_fa47_or0 = s_dadda_pg_rca24_fa47_and0 | s_dadda_pg_rca24_fa47_and1;
  assign s_dadda_pg_rca24_and_13_0 = a[13] & b[0];
  assign s_dadda_pg_rca24_and_12_1 = a[12] & b[1];
  assign s_dadda_pg_rca24_fa48_xor0 = s_dadda_pg_rca24_fa40_or0 ^ s_dadda_pg_rca24_and_13_0;
  assign s_dadda_pg_rca24_fa48_and0 = s_dadda_pg_rca24_fa40_or0 & s_dadda_pg_rca24_and_13_0;
  assign s_dadda_pg_rca24_fa48_xor1 = s_dadda_pg_rca24_fa48_xor0 ^ s_dadda_pg_rca24_and_12_1;
  assign s_dadda_pg_rca24_fa48_and1 = s_dadda_pg_rca24_fa48_xor0 & s_dadda_pg_rca24_and_12_1;
  assign s_dadda_pg_rca24_fa48_or0 = s_dadda_pg_rca24_fa48_and0 | s_dadda_pg_rca24_fa48_and1;
  assign s_dadda_pg_rca24_and_11_2 = a[11] & b[2];
  assign s_dadda_pg_rca24_and_10_3 = a[10] & b[3];
  assign s_dadda_pg_rca24_and_9_4 = a[9] & b[4];
  assign s_dadda_pg_rca24_fa49_xor0 = s_dadda_pg_rca24_and_11_2 ^ s_dadda_pg_rca24_and_10_3;
  assign s_dadda_pg_rca24_fa49_and0 = s_dadda_pg_rca24_and_11_2 & s_dadda_pg_rca24_and_10_3;
  assign s_dadda_pg_rca24_fa49_xor1 = s_dadda_pg_rca24_fa49_xor0 ^ s_dadda_pg_rca24_and_9_4;
  assign s_dadda_pg_rca24_fa49_and1 = s_dadda_pg_rca24_fa49_xor0 & s_dadda_pg_rca24_and_9_4;
  assign s_dadda_pg_rca24_fa49_or0 = s_dadda_pg_rca24_fa49_and0 | s_dadda_pg_rca24_fa49_and1;
  assign s_dadda_pg_rca24_and_8_5 = a[8] & b[5];
  assign s_dadda_pg_rca24_and_7_6 = a[7] & b[6];
  assign s_dadda_pg_rca24_and_6_7 = a[6] & b[7];
  assign s_dadda_pg_rca24_fa50_xor0 = s_dadda_pg_rca24_and_8_5 ^ s_dadda_pg_rca24_and_7_6;
  assign s_dadda_pg_rca24_fa50_and0 = s_dadda_pg_rca24_and_8_5 & s_dadda_pg_rca24_and_7_6;
  assign s_dadda_pg_rca24_fa50_xor1 = s_dadda_pg_rca24_fa50_xor0 ^ s_dadda_pg_rca24_and_6_7;
  assign s_dadda_pg_rca24_fa50_and1 = s_dadda_pg_rca24_fa50_xor0 & s_dadda_pg_rca24_and_6_7;
  assign s_dadda_pg_rca24_fa50_or0 = s_dadda_pg_rca24_fa50_and0 | s_dadda_pg_rca24_fa50_and1;
  assign s_dadda_pg_rca24_and_5_8 = a[5] & b[8];
  assign s_dadda_pg_rca24_and_4_9 = a[4] & b[9];
  assign s_dadda_pg_rca24_and_3_10 = a[3] & b[10];
  assign s_dadda_pg_rca24_fa51_xor0 = s_dadda_pg_rca24_and_5_8 ^ s_dadda_pg_rca24_and_4_9;
  assign s_dadda_pg_rca24_fa51_and0 = s_dadda_pg_rca24_and_5_8 & s_dadda_pg_rca24_and_4_9;
  assign s_dadda_pg_rca24_fa51_xor1 = s_dadda_pg_rca24_fa51_xor0 ^ s_dadda_pg_rca24_and_3_10;
  assign s_dadda_pg_rca24_fa51_and1 = s_dadda_pg_rca24_fa51_xor0 & s_dadda_pg_rca24_and_3_10;
  assign s_dadda_pg_rca24_fa51_or0 = s_dadda_pg_rca24_fa51_and0 | s_dadda_pg_rca24_fa51_and1;
  assign s_dadda_pg_rca24_and_2_11 = a[2] & b[11];
  assign s_dadda_pg_rca24_and_1_12 = a[1] & b[12];
  assign s_dadda_pg_rca24_and_0_13 = a[0] & b[13];
  assign s_dadda_pg_rca24_fa52_xor0 = s_dadda_pg_rca24_and_2_11 ^ s_dadda_pg_rca24_and_1_12;
  assign s_dadda_pg_rca24_fa52_and0 = s_dadda_pg_rca24_and_2_11 & s_dadda_pg_rca24_and_1_12;
  assign s_dadda_pg_rca24_fa52_xor1 = s_dadda_pg_rca24_fa52_xor0 ^ s_dadda_pg_rca24_and_0_13;
  assign s_dadda_pg_rca24_fa52_and1 = s_dadda_pg_rca24_fa52_xor0 & s_dadda_pg_rca24_and_0_13;
  assign s_dadda_pg_rca24_fa52_or0 = s_dadda_pg_rca24_fa52_and0 | s_dadda_pg_rca24_fa52_and1;
  assign s_dadda_pg_rca24_ha12_xor0 = s_dadda_pg_rca24_fa46_xor1 ^ s_dadda_pg_rca24_fa47_xor1;
  assign s_dadda_pg_rca24_ha12_and0 = s_dadda_pg_rca24_fa46_xor1 & s_dadda_pg_rca24_fa47_xor1;
  assign s_dadda_pg_rca24_fa53_xor0 = s_dadda_pg_rca24_ha12_and0 ^ s_dadda_pg_rca24_fa52_or0;
  assign s_dadda_pg_rca24_fa53_and0 = s_dadda_pg_rca24_ha12_and0 & s_dadda_pg_rca24_fa52_or0;
  assign s_dadda_pg_rca24_fa53_xor1 = s_dadda_pg_rca24_fa53_xor0 ^ s_dadda_pg_rca24_fa51_or0;
  assign s_dadda_pg_rca24_fa53_and1 = s_dadda_pg_rca24_fa53_xor0 & s_dadda_pg_rca24_fa51_or0;
  assign s_dadda_pg_rca24_fa53_or0 = s_dadda_pg_rca24_fa53_and0 | s_dadda_pg_rca24_fa53_and1;
  assign s_dadda_pg_rca24_fa54_xor0 = s_dadda_pg_rca24_fa50_or0 ^ s_dadda_pg_rca24_fa49_or0;
  assign s_dadda_pg_rca24_fa54_and0 = s_dadda_pg_rca24_fa50_or0 & s_dadda_pg_rca24_fa49_or0;
  assign s_dadda_pg_rca24_fa54_xor1 = s_dadda_pg_rca24_fa54_xor0 ^ s_dadda_pg_rca24_fa48_or0;
  assign s_dadda_pg_rca24_fa54_and1 = s_dadda_pg_rca24_fa54_xor0 & s_dadda_pg_rca24_fa48_or0;
  assign s_dadda_pg_rca24_fa54_or0 = s_dadda_pg_rca24_fa54_and0 | s_dadda_pg_rca24_fa54_and1;
  assign s_dadda_pg_rca24_and_14_0 = a[14] & b[0];
  assign s_dadda_pg_rca24_fa55_xor0 = s_dadda_pg_rca24_fa47_or0 ^ s_dadda_pg_rca24_fa46_or0;
  assign s_dadda_pg_rca24_fa55_and0 = s_dadda_pg_rca24_fa47_or0 & s_dadda_pg_rca24_fa46_or0;
  assign s_dadda_pg_rca24_fa55_xor1 = s_dadda_pg_rca24_fa55_xor0 ^ s_dadda_pg_rca24_and_14_0;
  assign s_dadda_pg_rca24_fa55_and1 = s_dadda_pg_rca24_fa55_xor0 & s_dadda_pg_rca24_and_14_0;
  assign s_dadda_pg_rca24_fa55_or0 = s_dadda_pg_rca24_fa55_and0 | s_dadda_pg_rca24_fa55_and1;
  assign s_dadda_pg_rca24_and_13_1 = a[13] & b[1];
  assign s_dadda_pg_rca24_and_12_2 = a[12] & b[2];
  assign s_dadda_pg_rca24_and_11_3 = a[11] & b[3];
  assign s_dadda_pg_rca24_fa56_xor0 = s_dadda_pg_rca24_and_13_1 ^ s_dadda_pg_rca24_and_12_2;
  assign s_dadda_pg_rca24_fa56_and0 = s_dadda_pg_rca24_and_13_1 & s_dadda_pg_rca24_and_12_2;
  assign s_dadda_pg_rca24_fa56_xor1 = s_dadda_pg_rca24_fa56_xor0 ^ s_dadda_pg_rca24_and_11_3;
  assign s_dadda_pg_rca24_fa56_and1 = s_dadda_pg_rca24_fa56_xor0 & s_dadda_pg_rca24_and_11_3;
  assign s_dadda_pg_rca24_fa56_or0 = s_dadda_pg_rca24_fa56_and0 | s_dadda_pg_rca24_fa56_and1;
  assign s_dadda_pg_rca24_and_10_4 = a[10] & b[4];
  assign s_dadda_pg_rca24_and_9_5 = a[9] & b[5];
  assign s_dadda_pg_rca24_and_8_6 = a[8] & b[6];
  assign s_dadda_pg_rca24_fa57_xor0 = s_dadda_pg_rca24_and_10_4 ^ s_dadda_pg_rca24_and_9_5;
  assign s_dadda_pg_rca24_fa57_and0 = s_dadda_pg_rca24_and_10_4 & s_dadda_pg_rca24_and_9_5;
  assign s_dadda_pg_rca24_fa57_xor1 = s_dadda_pg_rca24_fa57_xor0 ^ s_dadda_pg_rca24_and_8_6;
  assign s_dadda_pg_rca24_fa57_and1 = s_dadda_pg_rca24_fa57_xor0 & s_dadda_pg_rca24_and_8_6;
  assign s_dadda_pg_rca24_fa57_or0 = s_dadda_pg_rca24_fa57_and0 | s_dadda_pg_rca24_fa57_and1;
  assign s_dadda_pg_rca24_and_7_7 = a[7] & b[7];
  assign s_dadda_pg_rca24_and_6_8 = a[6] & b[8];
  assign s_dadda_pg_rca24_and_5_9 = a[5] & b[9];
  assign s_dadda_pg_rca24_fa58_xor0 = s_dadda_pg_rca24_and_7_7 ^ s_dadda_pg_rca24_and_6_8;
  assign s_dadda_pg_rca24_fa58_and0 = s_dadda_pg_rca24_and_7_7 & s_dadda_pg_rca24_and_6_8;
  assign s_dadda_pg_rca24_fa58_xor1 = s_dadda_pg_rca24_fa58_xor0 ^ s_dadda_pg_rca24_and_5_9;
  assign s_dadda_pg_rca24_fa58_and1 = s_dadda_pg_rca24_fa58_xor0 & s_dadda_pg_rca24_and_5_9;
  assign s_dadda_pg_rca24_fa58_or0 = s_dadda_pg_rca24_fa58_and0 | s_dadda_pg_rca24_fa58_and1;
  assign s_dadda_pg_rca24_and_4_10 = a[4] & b[10];
  assign s_dadda_pg_rca24_and_3_11 = a[3] & b[11];
  assign s_dadda_pg_rca24_and_2_12 = a[2] & b[12];
  assign s_dadda_pg_rca24_fa59_xor0 = s_dadda_pg_rca24_and_4_10 ^ s_dadda_pg_rca24_and_3_11;
  assign s_dadda_pg_rca24_fa59_and0 = s_dadda_pg_rca24_and_4_10 & s_dadda_pg_rca24_and_3_11;
  assign s_dadda_pg_rca24_fa59_xor1 = s_dadda_pg_rca24_fa59_xor0 ^ s_dadda_pg_rca24_and_2_12;
  assign s_dadda_pg_rca24_fa59_and1 = s_dadda_pg_rca24_fa59_xor0 & s_dadda_pg_rca24_and_2_12;
  assign s_dadda_pg_rca24_fa59_or0 = s_dadda_pg_rca24_fa59_and0 | s_dadda_pg_rca24_fa59_and1;
  assign s_dadda_pg_rca24_and_1_13 = a[1] & b[13];
  assign s_dadda_pg_rca24_and_0_14 = a[0] & b[14];
  assign s_dadda_pg_rca24_fa60_xor0 = s_dadda_pg_rca24_and_1_13 ^ s_dadda_pg_rca24_and_0_14;
  assign s_dadda_pg_rca24_fa60_and0 = s_dadda_pg_rca24_and_1_13 & s_dadda_pg_rca24_and_0_14;
  assign s_dadda_pg_rca24_fa60_xor1 = s_dadda_pg_rca24_fa60_xor0 ^ s_dadda_pg_rca24_fa53_xor1;
  assign s_dadda_pg_rca24_fa60_and1 = s_dadda_pg_rca24_fa60_xor0 & s_dadda_pg_rca24_fa53_xor1;
  assign s_dadda_pg_rca24_fa60_or0 = s_dadda_pg_rca24_fa60_and0 | s_dadda_pg_rca24_fa60_and1;
  assign s_dadda_pg_rca24_ha13_xor0 = s_dadda_pg_rca24_fa54_xor1 ^ s_dadda_pg_rca24_fa55_xor1;
  assign s_dadda_pg_rca24_ha13_and0 = s_dadda_pg_rca24_fa54_xor1 & s_dadda_pg_rca24_fa55_xor1;
  assign s_dadda_pg_rca24_fa61_xor0 = s_dadda_pg_rca24_ha13_and0 ^ s_dadda_pg_rca24_fa60_or0;
  assign s_dadda_pg_rca24_fa61_and0 = s_dadda_pg_rca24_ha13_and0 & s_dadda_pg_rca24_fa60_or0;
  assign s_dadda_pg_rca24_fa61_xor1 = s_dadda_pg_rca24_fa61_xor0 ^ s_dadda_pg_rca24_fa59_or0;
  assign s_dadda_pg_rca24_fa61_and1 = s_dadda_pg_rca24_fa61_xor0 & s_dadda_pg_rca24_fa59_or0;
  assign s_dadda_pg_rca24_fa61_or0 = s_dadda_pg_rca24_fa61_and0 | s_dadda_pg_rca24_fa61_and1;
  assign s_dadda_pg_rca24_fa62_xor0 = s_dadda_pg_rca24_fa58_or0 ^ s_dadda_pg_rca24_fa57_or0;
  assign s_dadda_pg_rca24_fa62_and0 = s_dadda_pg_rca24_fa58_or0 & s_dadda_pg_rca24_fa57_or0;
  assign s_dadda_pg_rca24_fa62_xor1 = s_dadda_pg_rca24_fa62_xor0 ^ s_dadda_pg_rca24_fa56_or0;
  assign s_dadda_pg_rca24_fa62_and1 = s_dadda_pg_rca24_fa62_xor0 & s_dadda_pg_rca24_fa56_or0;
  assign s_dadda_pg_rca24_fa62_or0 = s_dadda_pg_rca24_fa62_and0 | s_dadda_pg_rca24_fa62_and1;
  assign s_dadda_pg_rca24_fa63_xor0 = s_dadda_pg_rca24_fa55_or0 ^ s_dadda_pg_rca24_fa54_or0;
  assign s_dadda_pg_rca24_fa63_and0 = s_dadda_pg_rca24_fa55_or0 & s_dadda_pg_rca24_fa54_or0;
  assign s_dadda_pg_rca24_fa63_xor1 = s_dadda_pg_rca24_fa63_xor0 ^ s_dadda_pg_rca24_fa53_or0;
  assign s_dadda_pg_rca24_fa63_and1 = s_dadda_pg_rca24_fa63_xor0 & s_dadda_pg_rca24_fa53_or0;
  assign s_dadda_pg_rca24_fa63_or0 = s_dadda_pg_rca24_fa63_and0 | s_dadda_pg_rca24_fa63_and1;
  assign s_dadda_pg_rca24_and_15_0 = a[15] & b[0];
  assign s_dadda_pg_rca24_and_14_1 = a[14] & b[1];
  assign s_dadda_pg_rca24_and_13_2 = a[13] & b[2];
  assign s_dadda_pg_rca24_fa64_xor0 = s_dadda_pg_rca24_and_15_0 ^ s_dadda_pg_rca24_and_14_1;
  assign s_dadda_pg_rca24_fa64_and0 = s_dadda_pg_rca24_and_15_0 & s_dadda_pg_rca24_and_14_1;
  assign s_dadda_pg_rca24_fa64_xor1 = s_dadda_pg_rca24_fa64_xor0 ^ s_dadda_pg_rca24_and_13_2;
  assign s_dadda_pg_rca24_fa64_and1 = s_dadda_pg_rca24_fa64_xor0 & s_dadda_pg_rca24_and_13_2;
  assign s_dadda_pg_rca24_fa64_or0 = s_dadda_pg_rca24_fa64_and0 | s_dadda_pg_rca24_fa64_and1;
  assign s_dadda_pg_rca24_and_12_3 = a[12] & b[3];
  assign s_dadda_pg_rca24_and_11_4 = a[11] & b[4];
  assign s_dadda_pg_rca24_and_10_5 = a[10] & b[5];
  assign s_dadda_pg_rca24_fa65_xor0 = s_dadda_pg_rca24_and_12_3 ^ s_dadda_pg_rca24_and_11_4;
  assign s_dadda_pg_rca24_fa65_and0 = s_dadda_pg_rca24_and_12_3 & s_dadda_pg_rca24_and_11_4;
  assign s_dadda_pg_rca24_fa65_xor1 = s_dadda_pg_rca24_fa65_xor0 ^ s_dadda_pg_rca24_and_10_5;
  assign s_dadda_pg_rca24_fa65_and1 = s_dadda_pg_rca24_fa65_xor0 & s_dadda_pg_rca24_and_10_5;
  assign s_dadda_pg_rca24_fa65_or0 = s_dadda_pg_rca24_fa65_and0 | s_dadda_pg_rca24_fa65_and1;
  assign s_dadda_pg_rca24_and_9_6 = a[9] & b[6];
  assign s_dadda_pg_rca24_and_8_7 = a[8] & b[7];
  assign s_dadda_pg_rca24_and_7_8 = a[7] & b[8];
  assign s_dadda_pg_rca24_fa66_xor0 = s_dadda_pg_rca24_and_9_6 ^ s_dadda_pg_rca24_and_8_7;
  assign s_dadda_pg_rca24_fa66_and0 = s_dadda_pg_rca24_and_9_6 & s_dadda_pg_rca24_and_8_7;
  assign s_dadda_pg_rca24_fa66_xor1 = s_dadda_pg_rca24_fa66_xor0 ^ s_dadda_pg_rca24_and_7_8;
  assign s_dadda_pg_rca24_fa66_and1 = s_dadda_pg_rca24_fa66_xor0 & s_dadda_pg_rca24_and_7_8;
  assign s_dadda_pg_rca24_fa66_or0 = s_dadda_pg_rca24_fa66_and0 | s_dadda_pg_rca24_fa66_and1;
  assign s_dadda_pg_rca24_and_6_9 = a[6] & b[9];
  assign s_dadda_pg_rca24_and_5_10 = a[5] & b[10];
  assign s_dadda_pg_rca24_and_4_11 = a[4] & b[11];
  assign s_dadda_pg_rca24_fa67_xor0 = s_dadda_pg_rca24_and_6_9 ^ s_dadda_pg_rca24_and_5_10;
  assign s_dadda_pg_rca24_fa67_and0 = s_dadda_pg_rca24_and_6_9 & s_dadda_pg_rca24_and_5_10;
  assign s_dadda_pg_rca24_fa67_xor1 = s_dadda_pg_rca24_fa67_xor0 ^ s_dadda_pg_rca24_and_4_11;
  assign s_dadda_pg_rca24_fa67_and1 = s_dadda_pg_rca24_fa67_xor0 & s_dadda_pg_rca24_and_4_11;
  assign s_dadda_pg_rca24_fa67_or0 = s_dadda_pg_rca24_fa67_and0 | s_dadda_pg_rca24_fa67_and1;
  assign s_dadda_pg_rca24_and_3_12 = a[3] & b[12];
  assign s_dadda_pg_rca24_and_2_13 = a[2] & b[13];
  assign s_dadda_pg_rca24_and_1_14 = a[1] & b[14];
  assign s_dadda_pg_rca24_fa68_xor0 = s_dadda_pg_rca24_and_3_12 ^ s_dadda_pg_rca24_and_2_13;
  assign s_dadda_pg_rca24_fa68_and0 = s_dadda_pg_rca24_and_3_12 & s_dadda_pg_rca24_and_2_13;
  assign s_dadda_pg_rca24_fa68_xor1 = s_dadda_pg_rca24_fa68_xor0 ^ s_dadda_pg_rca24_and_1_14;
  assign s_dadda_pg_rca24_fa68_and1 = s_dadda_pg_rca24_fa68_xor0 & s_dadda_pg_rca24_and_1_14;
  assign s_dadda_pg_rca24_fa68_or0 = s_dadda_pg_rca24_fa68_and0 | s_dadda_pg_rca24_fa68_and1;
  assign s_dadda_pg_rca24_and_0_15 = a[0] & b[15];
  assign s_dadda_pg_rca24_fa69_xor0 = s_dadda_pg_rca24_and_0_15 ^ s_dadda_pg_rca24_fa61_xor1;
  assign s_dadda_pg_rca24_fa69_and0 = s_dadda_pg_rca24_and_0_15 & s_dadda_pg_rca24_fa61_xor1;
  assign s_dadda_pg_rca24_fa69_xor1 = s_dadda_pg_rca24_fa69_xor0 ^ s_dadda_pg_rca24_fa62_xor1;
  assign s_dadda_pg_rca24_fa69_and1 = s_dadda_pg_rca24_fa69_xor0 & s_dadda_pg_rca24_fa62_xor1;
  assign s_dadda_pg_rca24_fa69_or0 = s_dadda_pg_rca24_fa69_and0 | s_dadda_pg_rca24_fa69_and1;
  assign s_dadda_pg_rca24_ha14_xor0 = s_dadda_pg_rca24_fa63_xor1 ^ s_dadda_pg_rca24_fa64_xor1;
  assign s_dadda_pg_rca24_ha14_and0 = s_dadda_pg_rca24_fa63_xor1 & s_dadda_pg_rca24_fa64_xor1;
  assign s_dadda_pg_rca24_fa70_xor0 = s_dadda_pg_rca24_ha14_and0 ^ s_dadda_pg_rca24_fa69_or0;
  assign s_dadda_pg_rca24_fa70_and0 = s_dadda_pg_rca24_ha14_and0 & s_dadda_pg_rca24_fa69_or0;
  assign s_dadda_pg_rca24_fa70_xor1 = s_dadda_pg_rca24_fa70_xor0 ^ s_dadda_pg_rca24_fa68_or0;
  assign s_dadda_pg_rca24_fa70_and1 = s_dadda_pg_rca24_fa70_xor0 & s_dadda_pg_rca24_fa68_or0;
  assign s_dadda_pg_rca24_fa70_or0 = s_dadda_pg_rca24_fa70_and0 | s_dadda_pg_rca24_fa70_and1;
  assign s_dadda_pg_rca24_fa71_xor0 = s_dadda_pg_rca24_fa67_or0 ^ s_dadda_pg_rca24_fa66_or0;
  assign s_dadda_pg_rca24_fa71_and0 = s_dadda_pg_rca24_fa67_or0 & s_dadda_pg_rca24_fa66_or0;
  assign s_dadda_pg_rca24_fa71_xor1 = s_dadda_pg_rca24_fa71_xor0 ^ s_dadda_pg_rca24_fa65_or0;
  assign s_dadda_pg_rca24_fa71_and1 = s_dadda_pg_rca24_fa71_xor0 & s_dadda_pg_rca24_fa65_or0;
  assign s_dadda_pg_rca24_fa71_or0 = s_dadda_pg_rca24_fa71_and0 | s_dadda_pg_rca24_fa71_and1;
  assign s_dadda_pg_rca24_fa72_xor0 = s_dadda_pg_rca24_fa64_or0 ^ s_dadda_pg_rca24_fa63_or0;
  assign s_dadda_pg_rca24_fa72_and0 = s_dadda_pg_rca24_fa64_or0 & s_dadda_pg_rca24_fa63_or0;
  assign s_dadda_pg_rca24_fa72_xor1 = s_dadda_pg_rca24_fa72_xor0 ^ s_dadda_pg_rca24_fa62_or0;
  assign s_dadda_pg_rca24_fa72_and1 = s_dadda_pg_rca24_fa72_xor0 & s_dadda_pg_rca24_fa62_or0;
  assign s_dadda_pg_rca24_fa72_or0 = s_dadda_pg_rca24_fa72_and0 | s_dadda_pg_rca24_fa72_and1;
  assign s_dadda_pg_rca24_and_16_0 = a[16] & b[0];
  assign s_dadda_pg_rca24_and_15_1 = a[15] & b[1];
  assign s_dadda_pg_rca24_fa73_xor0 = s_dadda_pg_rca24_fa61_or0 ^ s_dadda_pg_rca24_and_16_0;
  assign s_dadda_pg_rca24_fa73_and0 = s_dadda_pg_rca24_fa61_or0 & s_dadda_pg_rca24_and_16_0;
  assign s_dadda_pg_rca24_fa73_xor1 = s_dadda_pg_rca24_fa73_xor0 ^ s_dadda_pg_rca24_and_15_1;
  assign s_dadda_pg_rca24_fa73_and1 = s_dadda_pg_rca24_fa73_xor0 & s_dadda_pg_rca24_and_15_1;
  assign s_dadda_pg_rca24_fa73_or0 = s_dadda_pg_rca24_fa73_and0 | s_dadda_pg_rca24_fa73_and1;
  assign s_dadda_pg_rca24_and_14_2 = a[14] & b[2];
  assign s_dadda_pg_rca24_and_13_3 = a[13] & b[3];
  assign s_dadda_pg_rca24_and_12_4 = a[12] & b[4];
  assign s_dadda_pg_rca24_fa74_xor0 = s_dadda_pg_rca24_and_14_2 ^ s_dadda_pg_rca24_and_13_3;
  assign s_dadda_pg_rca24_fa74_and0 = s_dadda_pg_rca24_and_14_2 & s_dadda_pg_rca24_and_13_3;
  assign s_dadda_pg_rca24_fa74_xor1 = s_dadda_pg_rca24_fa74_xor0 ^ s_dadda_pg_rca24_and_12_4;
  assign s_dadda_pg_rca24_fa74_and1 = s_dadda_pg_rca24_fa74_xor0 & s_dadda_pg_rca24_and_12_4;
  assign s_dadda_pg_rca24_fa74_or0 = s_dadda_pg_rca24_fa74_and0 | s_dadda_pg_rca24_fa74_and1;
  assign s_dadda_pg_rca24_and_11_5 = a[11] & b[5];
  assign s_dadda_pg_rca24_and_10_6 = a[10] & b[6];
  assign s_dadda_pg_rca24_and_9_7 = a[9] & b[7];
  assign s_dadda_pg_rca24_fa75_xor0 = s_dadda_pg_rca24_and_11_5 ^ s_dadda_pg_rca24_and_10_6;
  assign s_dadda_pg_rca24_fa75_and0 = s_dadda_pg_rca24_and_11_5 & s_dadda_pg_rca24_and_10_6;
  assign s_dadda_pg_rca24_fa75_xor1 = s_dadda_pg_rca24_fa75_xor0 ^ s_dadda_pg_rca24_and_9_7;
  assign s_dadda_pg_rca24_fa75_and1 = s_dadda_pg_rca24_fa75_xor0 & s_dadda_pg_rca24_and_9_7;
  assign s_dadda_pg_rca24_fa75_or0 = s_dadda_pg_rca24_fa75_and0 | s_dadda_pg_rca24_fa75_and1;
  assign s_dadda_pg_rca24_and_8_8 = a[8] & b[8];
  assign s_dadda_pg_rca24_and_7_9 = a[7] & b[9];
  assign s_dadda_pg_rca24_and_6_10 = a[6] & b[10];
  assign s_dadda_pg_rca24_fa76_xor0 = s_dadda_pg_rca24_and_8_8 ^ s_dadda_pg_rca24_and_7_9;
  assign s_dadda_pg_rca24_fa76_and0 = s_dadda_pg_rca24_and_8_8 & s_dadda_pg_rca24_and_7_9;
  assign s_dadda_pg_rca24_fa76_xor1 = s_dadda_pg_rca24_fa76_xor0 ^ s_dadda_pg_rca24_and_6_10;
  assign s_dadda_pg_rca24_fa76_and1 = s_dadda_pg_rca24_fa76_xor0 & s_dadda_pg_rca24_and_6_10;
  assign s_dadda_pg_rca24_fa76_or0 = s_dadda_pg_rca24_fa76_and0 | s_dadda_pg_rca24_fa76_and1;
  assign s_dadda_pg_rca24_and_5_11 = a[5] & b[11];
  assign s_dadda_pg_rca24_and_4_12 = a[4] & b[12];
  assign s_dadda_pg_rca24_and_3_13 = a[3] & b[13];
  assign s_dadda_pg_rca24_fa77_xor0 = s_dadda_pg_rca24_and_5_11 ^ s_dadda_pg_rca24_and_4_12;
  assign s_dadda_pg_rca24_fa77_and0 = s_dadda_pg_rca24_and_5_11 & s_dadda_pg_rca24_and_4_12;
  assign s_dadda_pg_rca24_fa77_xor1 = s_dadda_pg_rca24_fa77_xor0 ^ s_dadda_pg_rca24_and_3_13;
  assign s_dadda_pg_rca24_fa77_and1 = s_dadda_pg_rca24_fa77_xor0 & s_dadda_pg_rca24_and_3_13;
  assign s_dadda_pg_rca24_fa77_or0 = s_dadda_pg_rca24_fa77_and0 | s_dadda_pg_rca24_fa77_and1;
  assign s_dadda_pg_rca24_and_2_14 = a[2] & b[14];
  assign s_dadda_pg_rca24_and_1_15 = a[1] & b[15];
  assign s_dadda_pg_rca24_and_0_16 = a[0] & b[16];
  assign s_dadda_pg_rca24_fa78_xor0 = s_dadda_pg_rca24_and_2_14 ^ s_dadda_pg_rca24_and_1_15;
  assign s_dadda_pg_rca24_fa78_and0 = s_dadda_pg_rca24_and_2_14 & s_dadda_pg_rca24_and_1_15;
  assign s_dadda_pg_rca24_fa78_xor1 = s_dadda_pg_rca24_fa78_xor0 ^ s_dadda_pg_rca24_and_0_16;
  assign s_dadda_pg_rca24_fa78_and1 = s_dadda_pg_rca24_fa78_xor0 & s_dadda_pg_rca24_and_0_16;
  assign s_dadda_pg_rca24_fa78_or0 = s_dadda_pg_rca24_fa78_and0 | s_dadda_pg_rca24_fa78_and1;
  assign s_dadda_pg_rca24_fa79_xor0 = s_dadda_pg_rca24_fa70_xor1 ^ s_dadda_pg_rca24_fa71_xor1;
  assign s_dadda_pg_rca24_fa79_and0 = s_dadda_pg_rca24_fa70_xor1 & s_dadda_pg_rca24_fa71_xor1;
  assign s_dadda_pg_rca24_fa79_xor1 = s_dadda_pg_rca24_fa79_xor0 ^ s_dadda_pg_rca24_fa72_xor1;
  assign s_dadda_pg_rca24_fa79_and1 = s_dadda_pg_rca24_fa79_xor0 & s_dadda_pg_rca24_fa72_xor1;
  assign s_dadda_pg_rca24_fa79_or0 = s_dadda_pg_rca24_fa79_and0 | s_dadda_pg_rca24_fa79_and1;
  assign s_dadda_pg_rca24_ha15_xor0 = s_dadda_pg_rca24_fa73_xor1 ^ s_dadda_pg_rca24_fa74_xor1;
  assign s_dadda_pg_rca24_ha15_and0 = s_dadda_pg_rca24_fa73_xor1 & s_dadda_pg_rca24_fa74_xor1;
  assign s_dadda_pg_rca24_fa80_xor0 = s_dadda_pg_rca24_ha15_and0 ^ s_dadda_pg_rca24_fa79_or0;
  assign s_dadda_pg_rca24_fa80_and0 = s_dadda_pg_rca24_ha15_and0 & s_dadda_pg_rca24_fa79_or0;
  assign s_dadda_pg_rca24_fa80_xor1 = s_dadda_pg_rca24_fa80_xor0 ^ s_dadda_pg_rca24_fa78_or0;
  assign s_dadda_pg_rca24_fa80_and1 = s_dadda_pg_rca24_fa80_xor0 & s_dadda_pg_rca24_fa78_or0;
  assign s_dadda_pg_rca24_fa80_or0 = s_dadda_pg_rca24_fa80_and0 | s_dadda_pg_rca24_fa80_and1;
  assign s_dadda_pg_rca24_fa81_xor0 = s_dadda_pg_rca24_fa77_or0 ^ s_dadda_pg_rca24_fa76_or0;
  assign s_dadda_pg_rca24_fa81_and0 = s_dadda_pg_rca24_fa77_or0 & s_dadda_pg_rca24_fa76_or0;
  assign s_dadda_pg_rca24_fa81_xor1 = s_dadda_pg_rca24_fa81_xor0 ^ s_dadda_pg_rca24_fa75_or0;
  assign s_dadda_pg_rca24_fa81_and1 = s_dadda_pg_rca24_fa81_xor0 & s_dadda_pg_rca24_fa75_or0;
  assign s_dadda_pg_rca24_fa81_or0 = s_dadda_pg_rca24_fa81_and0 | s_dadda_pg_rca24_fa81_and1;
  assign s_dadda_pg_rca24_fa82_xor0 = s_dadda_pg_rca24_fa74_or0 ^ s_dadda_pg_rca24_fa73_or0;
  assign s_dadda_pg_rca24_fa82_and0 = s_dadda_pg_rca24_fa74_or0 & s_dadda_pg_rca24_fa73_or0;
  assign s_dadda_pg_rca24_fa82_xor1 = s_dadda_pg_rca24_fa82_xor0 ^ s_dadda_pg_rca24_fa72_or0;
  assign s_dadda_pg_rca24_fa82_and1 = s_dadda_pg_rca24_fa82_xor0 & s_dadda_pg_rca24_fa72_or0;
  assign s_dadda_pg_rca24_fa82_or0 = s_dadda_pg_rca24_fa82_and0 | s_dadda_pg_rca24_fa82_and1;
  assign s_dadda_pg_rca24_and_17_0 = a[17] & b[0];
  assign s_dadda_pg_rca24_fa83_xor0 = s_dadda_pg_rca24_fa71_or0 ^ s_dadda_pg_rca24_fa70_or0;
  assign s_dadda_pg_rca24_fa83_and0 = s_dadda_pg_rca24_fa71_or0 & s_dadda_pg_rca24_fa70_or0;
  assign s_dadda_pg_rca24_fa83_xor1 = s_dadda_pg_rca24_fa83_xor0 ^ s_dadda_pg_rca24_and_17_0;
  assign s_dadda_pg_rca24_fa83_and1 = s_dadda_pg_rca24_fa83_xor0 & s_dadda_pg_rca24_and_17_0;
  assign s_dadda_pg_rca24_fa83_or0 = s_dadda_pg_rca24_fa83_and0 | s_dadda_pg_rca24_fa83_and1;
  assign s_dadda_pg_rca24_and_16_1 = a[16] & b[1];
  assign s_dadda_pg_rca24_and_15_2 = a[15] & b[2];
  assign s_dadda_pg_rca24_and_14_3 = a[14] & b[3];
  assign s_dadda_pg_rca24_fa84_xor0 = s_dadda_pg_rca24_and_16_1 ^ s_dadda_pg_rca24_and_15_2;
  assign s_dadda_pg_rca24_fa84_and0 = s_dadda_pg_rca24_and_16_1 & s_dadda_pg_rca24_and_15_2;
  assign s_dadda_pg_rca24_fa84_xor1 = s_dadda_pg_rca24_fa84_xor0 ^ s_dadda_pg_rca24_and_14_3;
  assign s_dadda_pg_rca24_fa84_and1 = s_dadda_pg_rca24_fa84_xor0 & s_dadda_pg_rca24_and_14_3;
  assign s_dadda_pg_rca24_fa84_or0 = s_dadda_pg_rca24_fa84_and0 | s_dadda_pg_rca24_fa84_and1;
  assign s_dadda_pg_rca24_and_13_4 = a[13] & b[4];
  assign s_dadda_pg_rca24_and_12_5 = a[12] & b[5];
  assign s_dadda_pg_rca24_and_11_6 = a[11] & b[6];
  assign s_dadda_pg_rca24_fa85_xor0 = s_dadda_pg_rca24_and_13_4 ^ s_dadda_pg_rca24_and_12_5;
  assign s_dadda_pg_rca24_fa85_and0 = s_dadda_pg_rca24_and_13_4 & s_dadda_pg_rca24_and_12_5;
  assign s_dadda_pg_rca24_fa85_xor1 = s_dadda_pg_rca24_fa85_xor0 ^ s_dadda_pg_rca24_and_11_6;
  assign s_dadda_pg_rca24_fa85_and1 = s_dadda_pg_rca24_fa85_xor0 & s_dadda_pg_rca24_and_11_6;
  assign s_dadda_pg_rca24_fa85_or0 = s_dadda_pg_rca24_fa85_and0 | s_dadda_pg_rca24_fa85_and1;
  assign s_dadda_pg_rca24_and_10_7 = a[10] & b[7];
  assign s_dadda_pg_rca24_and_9_8 = a[9] & b[8];
  assign s_dadda_pg_rca24_and_8_9 = a[8] & b[9];
  assign s_dadda_pg_rca24_fa86_xor0 = s_dadda_pg_rca24_and_10_7 ^ s_dadda_pg_rca24_and_9_8;
  assign s_dadda_pg_rca24_fa86_and0 = s_dadda_pg_rca24_and_10_7 & s_dadda_pg_rca24_and_9_8;
  assign s_dadda_pg_rca24_fa86_xor1 = s_dadda_pg_rca24_fa86_xor0 ^ s_dadda_pg_rca24_and_8_9;
  assign s_dadda_pg_rca24_fa86_and1 = s_dadda_pg_rca24_fa86_xor0 & s_dadda_pg_rca24_and_8_9;
  assign s_dadda_pg_rca24_fa86_or0 = s_dadda_pg_rca24_fa86_and0 | s_dadda_pg_rca24_fa86_and1;
  assign s_dadda_pg_rca24_and_7_10 = a[7] & b[10];
  assign s_dadda_pg_rca24_and_6_11 = a[6] & b[11];
  assign s_dadda_pg_rca24_and_5_12 = a[5] & b[12];
  assign s_dadda_pg_rca24_fa87_xor0 = s_dadda_pg_rca24_and_7_10 ^ s_dadda_pg_rca24_and_6_11;
  assign s_dadda_pg_rca24_fa87_and0 = s_dadda_pg_rca24_and_7_10 & s_dadda_pg_rca24_and_6_11;
  assign s_dadda_pg_rca24_fa87_xor1 = s_dadda_pg_rca24_fa87_xor0 ^ s_dadda_pg_rca24_and_5_12;
  assign s_dadda_pg_rca24_fa87_and1 = s_dadda_pg_rca24_fa87_xor0 & s_dadda_pg_rca24_and_5_12;
  assign s_dadda_pg_rca24_fa87_or0 = s_dadda_pg_rca24_fa87_and0 | s_dadda_pg_rca24_fa87_and1;
  assign s_dadda_pg_rca24_and_4_13 = a[4] & b[13];
  assign s_dadda_pg_rca24_and_3_14 = a[3] & b[14];
  assign s_dadda_pg_rca24_and_2_15 = a[2] & b[15];
  assign s_dadda_pg_rca24_fa88_xor0 = s_dadda_pg_rca24_and_4_13 ^ s_dadda_pg_rca24_and_3_14;
  assign s_dadda_pg_rca24_fa88_and0 = s_dadda_pg_rca24_and_4_13 & s_dadda_pg_rca24_and_3_14;
  assign s_dadda_pg_rca24_fa88_xor1 = s_dadda_pg_rca24_fa88_xor0 ^ s_dadda_pg_rca24_and_2_15;
  assign s_dadda_pg_rca24_fa88_and1 = s_dadda_pg_rca24_fa88_xor0 & s_dadda_pg_rca24_and_2_15;
  assign s_dadda_pg_rca24_fa88_or0 = s_dadda_pg_rca24_fa88_and0 | s_dadda_pg_rca24_fa88_and1;
  assign s_dadda_pg_rca24_and_1_16 = a[1] & b[16];
  assign s_dadda_pg_rca24_and_0_17 = a[0] & b[17];
  assign s_dadda_pg_rca24_fa89_xor0 = s_dadda_pg_rca24_and_1_16 ^ s_dadda_pg_rca24_and_0_17;
  assign s_dadda_pg_rca24_fa89_and0 = s_dadda_pg_rca24_and_1_16 & s_dadda_pg_rca24_and_0_17;
  assign s_dadda_pg_rca24_fa89_xor1 = s_dadda_pg_rca24_fa89_xor0 ^ s_dadda_pg_rca24_fa80_xor1;
  assign s_dadda_pg_rca24_fa89_and1 = s_dadda_pg_rca24_fa89_xor0 & s_dadda_pg_rca24_fa80_xor1;
  assign s_dadda_pg_rca24_fa89_or0 = s_dadda_pg_rca24_fa89_and0 | s_dadda_pg_rca24_fa89_and1;
  assign s_dadda_pg_rca24_fa90_xor0 = s_dadda_pg_rca24_fa81_xor1 ^ s_dadda_pg_rca24_fa82_xor1;
  assign s_dadda_pg_rca24_fa90_and0 = s_dadda_pg_rca24_fa81_xor1 & s_dadda_pg_rca24_fa82_xor1;
  assign s_dadda_pg_rca24_fa90_xor1 = s_dadda_pg_rca24_fa90_xor0 ^ s_dadda_pg_rca24_fa83_xor1;
  assign s_dadda_pg_rca24_fa90_and1 = s_dadda_pg_rca24_fa90_xor0 & s_dadda_pg_rca24_fa83_xor1;
  assign s_dadda_pg_rca24_fa90_or0 = s_dadda_pg_rca24_fa90_and0 | s_dadda_pg_rca24_fa90_and1;
  assign s_dadda_pg_rca24_ha16_xor0 = s_dadda_pg_rca24_fa84_xor1 ^ s_dadda_pg_rca24_fa85_xor1;
  assign s_dadda_pg_rca24_ha16_and0 = s_dadda_pg_rca24_fa84_xor1 & s_dadda_pg_rca24_fa85_xor1;
  assign s_dadda_pg_rca24_fa91_xor0 = s_dadda_pg_rca24_ha16_and0 ^ s_dadda_pg_rca24_fa90_or0;
  assign s_dadda_pg_rca24_fa91_and0 = s_dadda_pg_rca24_ha16_and0 & s_dadda_pg_rca24_fa90_or0;
  assign s_dadda_pg_rca24_fa91_xor1 = s_dadda_pg_rca24_fa91_xor0 ^ s_dadda_pg_rca24_fa89_or0;
  assign s_dadda_pg_rca24_fa91_and1 = s_dadda_pg_rca24_fa91_xor0 & s_dadda_pg_rca24_fa89_or0;
  assign s_dadda_pg_rca24_fa91_or0 = s_dadda_pg_rca24_fa91_and0 | s_dadda_pg_rca24_fa91_and1;
  assign s_dadda_pg_rca24_fa92_xor0 = s_dadda_pg_rca24_fa88_or0 ^ s_dadda_pg_rca24_fa87_or0;
  assign s_dadda_pg_rca24_fa92_and0 = s_dadda_pg_rca24_fa88_or0 & s_dadda_pg_rca24_fa87_or0;
  assign s_dadda_pg_rca24_fa92_xor1 = s_dadda_pg_rca24_fa92_xor0 ^ s_dadda_pg_rca24_fa86_or0;
  assign s_dadda_pg_rca24_fa92_and1 = s_dadda_pg_rca24_fa92_xor0 & s_dadda_pg_rca24_fa86_or0;
  assign s_dadda_pg_rca24_fa92_or0 = s_dadda_pg_rca24_fa92_and0 | s_dadda_pg_rca24_fa92_and1;
  assign s_dadda_pg_rca24_fa93_xor0 = s_dadda_pg_rca24_fa85_or0 ^ s_dadda_pg_rca24_fa84_or0;
  assign s_dadda_pg_rca24_fa93_and0 = s_dadda_pg_rca24_fa85_or0 & s_dadda_pg_rca24_fa84_or0;
  assign s_dadda_pg_rca24_fa93_xor1 = s_dadda_pg_rca24_fa93_xor0 ^ s_dadda_pg_rca24_fa83_or0;
  assign s_dadda_pg_rca24_fa93_and1 = s_dadda_pg_rca24_fa93_xor0 & s_dadda_pg_rca24_fa83_or0;
  assign s_dadda_pg_rca24_fa93_or0 = s_dadda_pg_rca24_fa93_and0 | s_dadda_pg_rca24_fa93_and1;
  assign s_dadda_pg_rca24_fa94_xor0 = s_dadda_pg_rca24_fa82_or0 ^ s_dadda_pg_rca24_fa81_or0;
  assign s_dadda_pg_rca24_fa94_and0 = s_dadda_pg_rca24_fa82_or0 & s_dadda_pg_rca24_fa81_or0;
  assign s_dadda_pg_rca24_fa94_xor1 = s_dadda_pg_rca24_fa94_xor0 ^ s_dadda_pg_rca24_fa80_or0;
  assign s_dadda_pg_rca24_fa94_and1 = s_dadda_pg_rca24_fa94_xor0 & s_dadda_pg_rca24_fa80_or0;
  assign s_dadda_pg_rca24_fa94_or0 = s_dadda_pg_rca24_fa94_and0 | s_dadda_pg_rca24_fa94_and1;
  assign s_dadda_pg_rca24_and_18_0 = a[18] & b[0];
  assign s_dadda_pg_rca24_and_17_1 = a[17] & b[1];
  assign s_dadda_pg_rca24_and_16_2 = a[16] & b[2];
  assign s_dadda_pg_rca24_fa95_xor0 = s_dadda_pg_rca24_and_18_0 ^ s_dadda_pg_rca24_and_17_1;
  assign s_dadda_pg_rca24_fa95_and0 = s_dadda_pg_rca24_and_18_0 & s_dadda_pg_rca24_and_17_1;
  assign s_dadda_pg_rca24_fa95_xor1 = s_dadda_pg_rca24_fa95_xor0 ^ s_dadda_pg_rca24_and_16_2;
  assign s_dadda_pg_rca24_fa95_and1 = s_dadda_pg_rca24_fa95_xor0 & s_dadda_pg_rca24_and_16_2;
  assign s_dadda_pg_rca24_fa95_or0 = s_dadda_pg_rca24_fa95_and0 | s_dadda_pg_rca24_fa95_and1;
  assign s_dadda_pg_rca24_and_15_3 = a[15] & b[3];
  assign s_dadda_pg_rca24_and_14_4 = a[14] & b[4];
  assign s_dadda_pg_rca24_and_13_5 = a[13] & b[5];
  assign s_dadda_pg_rca24_fa96_xor0 = s_dadda_pg_rca24_and_15_3 ^ s_dadda_pg_rca24_and_14_4;
  assign s_dadda_pg_rca24_fa96_and0 = s_dadda_pg_rca24_and_15_3 & s_dadda_pg_rca24_and_14_4;
  assign s_dadda_pg_rca24_fa96_xor1 = s_dadda_pg_rca24_fa96_xor0 ^ s_dadda_pg_rca24_and_13_5;
  assign s_dadda_pg_rca24_fa96_and1 = s_dadda_pg_rca24_fa96_xor0 & s_dadda_pg_rca24_and_13_5;
  assign s_dadda_pg_rca24_fa96_or0 = s_dadda_pg_rca24_fa96_and0 | s_dadda_pg_rca24_fa96_and1;
  assign s_dadda_pg_rca24_and_12_6 = a[12] & b[6];
  assign s_dadda_pg_rca24_and_11_7 = a[11] & b[7];
  assign s_dadda_pg_rca24_and_10_8 = a[10] & b[8];
  assign s_dadda_pg_rca24_fa97_xor0 = s_dadda_pg_rca24_and_12_6 ^ s_dadda_pg_rca24_and_11_7;
  assign s_dadda_pg_rca24_fa97_and0 = s_dadda_pg_rca24_and_12_6 & s_dadda_pg_rca24_and_11_7;
  assign s_dadda_pg_rca24_fa97_xor1 = s_dadda_pg_rca24_fa97_xor0 ^ s_dadda_pg_rca24_and_10_8;
  assign s_dadda_pg_rca24_fa97_and1 = s_dadda_pg_rca24_fa97_xor0 & s_dadda_pg_rca24_and_10_8;
  assign s_dadda_pg_rca24_fa97_or0 = s_dadda_pg_rca24_fa97_and0 | s_dadda_pg_rca24_fa97_and1;
  assign s_dadda_pg_rca24_and_9_9 = a[9] & b[9];
  assign s_dadda_pg_rca24_and_8_10 = a[8] & b[10];
  assign s_dadda_pg_rca24_and_7_11 = a[7] & b[11];
  assign s_dadda_pg_rca24_fa98_xor0 = s_dadda_pg_rca24_and_9_9 ^ s_dadda_pg_rca24_and_8_10;
  assign s_dadda_pg_rca24_fa98_and0 = s_dadda_pg_rca24_and_9_9 & s_dadda_pg_rca24_and_8_10;
  assign s_dadda_pg_rca24_fa98_xor1 = s_dadda_pg_rca24_fa98_xor0 ^ s_dadda_pg_rca24_and_7_11;
  assign s_dadda_pg_rca24_fa98_and1 = s_dadda_pg_rca24_fa98_xor0 & s_dadda_pg_rca24_and_7_11;
  assign s_dadda_pg_rca24_fa98_or0 = s_dadda_pg_rca24_fa98_and0 | s_dadda_pg_rca24_fa98_and1;
  assign s_dadda_pg_rca24_and_6_12 = a[6] & b[12];
  assign s_dadda_pg_rca24_and_5_13 = a[5] & b[13];
  assign s_dadda_pg_rca24_and_4_14 = a[4] & b[14];
  assign s_dadda_pg_rca24_fa99_xor0 = s_dadda_pg_rca24_and_6_12 ^ s_dadda_pg_rca24_and_5_13;
  assign s_dadda_pg_rca24_fa99_and0 = s_dadda_pg_rca24_and_6_12 & s_dadda_pg_rca24_and_5_13;
  assign s_dadda_pg_rca24_fa99_xor1 = s_dadda_pg_rca24_fa99_xor0 ^ s_dadda_pg_rca24_and_4_14;
  assign s_dadda_pg_rca24_fa99_and1 = s_dadda_pg_rca24_fa99_xor0 & s_dadda_pg_rca24_and_4_14;
  assign s_dadda_pg_rca24_fa99_or0 = s_dadda_pg_rca24_fa99_and0 | s_dadda_pg_rca24_fa99_and1;
  assign s_dadda_pg_rca24_and_3_15 = a[3] & b[15];
  assign s_dadda_pg_rca24_and_2_16 = a[2] & b[16];
  assign s_dadda_pg_rca24_and_1_17 = a[1] & b[17];
  assign s_dadda_pg_rca24_fa100_xor0 = s_dadda_pg_rca24_and_3_15 ^ s_dadda_pg_rca24_and_2_16;
  assign s_dadda_pg_rca24_fa100_and0 = s_dadda_pg_rca24_and_3_15 & s_dadda_pg_rca24_and_2_16;
  assign s_dadda_pg_rca24_fa100_xor1 = s_dadda_pg_rca24_fa100_xor0 ^ s_dadda_pg_rca24_and_1_17;
  assign s_dadda_pg_rca24_fa100_and1 = s_dadda_pg_rca24_fa100_xor0 & s_dadda_pg_rca24_and_1_17;
  assign s_dadda_pg_rca24_fa100_or0 = s_dadda_pg_rca24_fa100_and0 | s_dadda_pg_rca24_fa100_and1;
  assign s_dadda_pg_rca24_and_0_18 = a[0] & b[18];
  assign s_dadda_pg_rca24_fa101_xor0 = s_dadda_pg_rca24_and_0_18 ^ s_dadda_pg_rca24_fa91_xor1;
  assign s_dadda_pg_rca24_fa101_and0 = s_dadda_pg_rca24_and_0_18 & s_dadda_pg_rca24_fa91_xor1;
  assign s_dadda_pg_rca24_fa101_xor1 = s_dadda_pg_rca24_fa101_xor0 ^ s_dadda_pg_rca24_fa92_xor1;
  assign s_dadda_pg_rca24_fa101_and1 = s_dadda_pg_rca24_fa101_xor0 & s_dadda_pg_rca24_fa92_xor1;
  assign s_dadda_pg_rca24_fa101_or0 = s_dadda_pg_rca24_fa101_and0 | s_dadda_pg_rca24_fa101_and1;
  assign s_dadda_pg_rca24_fa102_xor0 = s_dadda_pg_rca24_fa93_xor1 ^ s_dadda_pg_rca24_fa94_xor1;
  assign s_dadda_pg_rca24_fa102_and0 = s_dadda_pg_rca24_fa93_xor1 & s_dadda_pg_rca24_fa94_xor1;
  assign s_dadda_pg_rca24_fa102_xor1 = s_dadda_pg_rca24_fa102_xor0 ^ s_dadda_pg_rca24_fa95_xor1;
  assign s_dadda_pg_rca24_fa102_and1 = s_dadda_pg_rca24_fa102_xor0 & s_dadda_pg_rca24_fa95_xor1;
  assign s_dadda_pg_rca24_fa102_or0 = s_dadda_pg_rca24_fa102_and0 | s_dadda_pg_rca24_fa102_and1;
  assign s_dadda_pg_rca24_ha17_xor0 = s_dadda_pg_rca24_fa96_xor1 ^ s_dadda_pg_rca24_fa97_xor1;
  assign s_dadda_pg_rca24_ha17_and0 = s_dadda_pg_rca24_fa96_xor1 & s_dadda_pg_rca24_fa97_xor1;
  assign s_dadda_pg_rca24_fa103_xor0 = s_dadda_pg_rca24_ha17_and0 ^ s_dadda_pg_rca24_fa102_or0;
  assign s_dadda_pg_rca24_fa103_and0 = s_dadda_pg_rca24_ha17_and0 & s_dadda_pg_rca24_fa102_or0;
  assign s_dadda_pg_rca24_fa103_xor1 = s_dadda_pg_rca24_fa103_xor0 ^ s_dadda_pg_rca24_fa101_or0;
  assign s_dadda_pg_rca24_fa103_and1 = s_dadda_pg_rca24_fa103_xor0 & s_dadda_pg_rca24_fa101_or0;
  assign s_dadda_pg_rca24_fa103_or0 = s_dadda_pg_rca24_fa103_and0 | s_dadda_pg_rca24_fa103_and1;
  assign s_dadda_pg_rca24_fa104_xor0 = s_dadda_pg_rca24_fa100_or0 ^ s_dadda_pg_rca24_fa99_or0;
  assign s_dadda_pg_rca24_fa104_and0 = s_dadda_pg_rca24_fa100_or0 & s_dadda_pg_rca24_fa99_or0;
  assign s_dadda_pg_rca24_fa104_xor1 = s_dadda_pg_rca24_fa104_xor0 ^ s_dadda_pg_rca24_fa98_or0;
  assign s_dadda_pg_rca24_fa104_and1 = s_dadda_pg_rca24_fa104_xor0 & s_dadda_pg_rca24_fa98_or0;
  assign s_dadda_pg_rca24_fa104_or0 = s_dadda_pg_rca24_fa104_and0 | s_dadda_pg_rca24_fa104_and1;
  assign s_dadda_pg_rca24_fa105_xor0 = s_dadda_pg_rca24_fa97_or0 ^ s_dadda_pg_rca24_fa96_or0;
  assign s_dadda_pg_rca24_fa105_and0 = s_dadda_pg_rca24_fa97_or0 & s_dadda_pg_rca24_fa96_or0;
  assign s_dadda_pg_rca24_fa105_xor1 = s_dadda_pg_rca24_fa105_xor0 ^ s_dadda_pg_rca24_fa95_or0;
  assign s_dadda_pg_rca24_fa105_and1 = s_dadda_pg_rca24_fa105_xor0 & s_dadda_pg_rca24_fa95_or0;
  assign s_dadda_pg_rca24_fa105_or0 = s_dadda_pg_rca24_fa105_and0 | s_dadda_pg_rca24_fa105_and1;
  assign s_dadda_pg_rca24_fa106_xor0 = s_dadda_pg_rca24_fa94_or0 ^ s_dadda_pg_rca24_fa93_or0;
  assign s_dadda_pg_rca24_fa106_and0 = s_dadda_pg_rca24_fa94_or0 & s_dadda_pg_rca24_fa93_or0;
  assign s_dadda_pg_rca24_fa106_xor1 = s_dadda_pg_rca24_fa106_xor0 ^ s_dadda_pg_rca24_fa92_or0;
  assign s_dadda_pg_rca24_fa106_and1 = s_dadda_pg_rca24_fa106_xor0 & s_dadda_pg_rca24_fa92_or0;
  assign s_dadda_pg_rca24_fa106_or0 = s_dadda_pg_rca24_fa106_and0 | s_dadda_pg_rca24_fa106_and1;
  assign s_dadda_pg_rca24_and_17_2 = a[17] & b[2];
  assign s_dadda_pg_rca24_and_16_3 = a[16] & b[3];
  assign s_dadda_pg_rca24_fa107_xor0 = s_dadda_pg_rca24_fa91_or0 ^ s_dadda_pg_rca24_and_17_2;
  assign s_dadda_pg_rca24_fa107_and0 = s_dadda_pg_rca24_fa91_or0 & s_dadda_pg_rca24_and_17_2;
  assign s_dadda_pg_rca24_fa107_xor1 = s_dadda_pg_rca24_fa107_xor0 ^ s_dadda_pg_rca24_and_16_3;
  assign s_dadda_pg_rca24_fa107_and1 = s_dadda_pg_rca24_fa107_xor0 & s_dadda_pg_rca24_and_16_3;
  assign s_dadda_pg_rca24_fa107_or0 = s_dadda_pg_rca24_fa107_and0 | s_dadda_pg_rca24_fa107_and1;
  assign s_dadda_pg_rca24_and_15_4 = a[15] & b[4];
  assign s_dadda_pg_rca24_and_14_5 = a[14] & b[5];
  assign s_dadda_pg_rca24_and_13_6 = a[13] & b[6];
  assign s_dadda_pg_rca24_fa108_xor0 = s_dadda_pg_rca24_and_15_4 ^ s_dadda_pg_rca24_and_14_5;
  assign s_dadda_pg_rca24_fa108_and0 = s_dadda_pg_rca24_and_15_4 & s_dadda_pg_rca24_and_14_5;
  assign s_dadda_pg_rca24_fa108_xor1 = s_dadda_pg_rca24_fa108_xor0 ^ s_dadda_pg_rca24_and_13_6;
  assign s_dadda_pg_rca24_fa108_and1 = s_dadda_pg_rca24_fa108_xor0 & s_dadda_pg_rca24_and_13_6;
  assign s_dadda_pg_rca24_fa108_or0 = s_dadda_pg_rca24_fa108_and0 | s_dadda_pg_rca24_fa108_and1;
  assign s_dadda_pg_rca24_and_12_7 = a[12] & b[7];
  assign s_dadda_pg_rca24_and_11_8 = a[11] & b[8];
  assign s_dadda_pg_rca24_and_10_9 = a[10] & b[9];
  assign s_dadda_pg_rca24_fa109_xor0 = s_dadda_pg_rca24_and_12_7 ^ s_dadda_pg_rca24_and_11_8;
  assign s_dadda_pg_rca24_fa109_and0 = s_dadda_pg_rca24_and_12_7 & s_dadda_pg_rca24_and_11_8;
  assign s_dadda_pg_rca24_fa109_xor1 = s_dadda_pg_rca24_fa109_xor0 ^ s_dadda_pg_rca24_and_10_9;
  assign s_dadda_pg_rca24_fa109_and1 = s_dadda_pg_rca24_fa109_xor0 & s_dadda_pg_rca24_and_10_9;
  assign s_dadda_pg_rca24_fa109_or0 = s_dadda_pg_rca24_fa109_and0 | s_dadda_pg_rca24_fa109_and1;
  assign s_dadda_pg_rca24_and_9_10 = a[9] & b[10];
  assign s_dadda_pg_rca24_and_8_11 = a[8] & b[11];
  assign s_dadda_pg_rca24_and_7_12 = a[7] & b[12];
  assign s_dadda_pg_rca24_fa110_xor0 = s_dadda_pg_rca24_and_9_10 ^ s_dadda_pg_rca24_and_8_11;
  assign s_dadda_pg_rca24_fa110_and0 = s_dadda_pg_rca24_and_9_10 & s_dadda_pg_rca24_and_8_11;
  assign s_dadda_pg_rca24_fa110_xor1 = s_dadda_pg_rca24_fa110_xor0 ^ s_dadda_pg_rca24_and_7_12;
  assign s_dadda_pg_rca24_fa110_and1 = s_dadda_pg_rca24_fa110_xor0 & s_dadda_pg_rca24_and_7_12;
  assign s_dadda_pg_rca24_fa110_or0 = s_dadda_pg_rca24_fa110_and0 | s_dadda_pg_rca24_fa110_and1;
  assign s_dadda_pg_rca24_and_6_13 = a[6] & b[13];
  assign s_dadda_pg_rca24_and_5_14 = a[5] & b[14];
  assign s_dadda_pg_rca24_and_4_15 = a[4] & b[15];
  assign s_dadda_pg_rca24_fa111_xor0 = s_dadda_pg_rca24_and_6_13 ^ s_dadda_pg_rca24_and_5_14;
  assign s_dadda_pg_rca24_fa111_and0 = s_dadda_pg_rca24_and_6_13 & s_dadda_pg_rca24_and_5_14;
  assign s_dadda_pg_rca24_fa111_xor1 = s_dadda_pg_rca24_fa111_xor0 ^ s_dadda_pg_rca24_and_4_15;
  assign s_dadda_pg_rca24_fa111_and1 = s_dadda_pg_rca24_fa111_xor0 & s_dadda_pg_rca24_and_4_15;
  assign s_dadda_pg_rca24_fa111_or0 = s_dadda_pg_rca24_fa111_and0 | s_dadda_pg_rca24_fa111_and1;
  assign s_dadda_pg_rca24_and_3_16 = a[3] & b[16];
  assign s_dadda_pg_rca24_and_2_17 = a[2] & b[17];
  assign s_dadda_pg_rca24_and_1_18 = a[1] & b[18];
  assign s_dadda_pg_rca24_fa112_xor0 = s_dadda_pg_rca24_and_3_16 ^ s_dadda_pg_rca24_and_2_17;
  assign s_dadda_pg_rca24_fa112_and0 = s_dadda_pg_rca24_and_3_16 & s_dadda_pg_rca24_and_2_17;
  assign s_dadda_pg_rca24_fa112_xor1 = s_dadda_pg_rca24_fa112_xor0 ^ s_dadda_pg_rca24_and_1_18;
  assign s_dadda_pg_rca24_fa112_and1 = s_dadda_pg_rca24_fa112_xor0 & s_dadda_pg_rca24_and_1_18;
  assign s_dadda_pg_rca24_fa112_or0 = s_dadda_pg_rca24_fa112_and0 | s_dadda_pg_rca24_fa112_and1;
  assign s_dadda_pg_rca24_and_0_19 = a[0] & b[19];
  assign s_dadda_pg_rca24_fa113_xor0 = s_dadda_pg_rca24_and_0_19 ^ s_dadda_pg_rca24_ha0_xor0;
  assign s_dadda_pg_rca24_fa113_and0 = s_dadda_pg_rca24_and_0_19 & s_dadda_pg_rca24_ha0_xor0;
  assign s_dadda_pg_rca24_fa113_xor1 = s_dadda_pg_rca24_fa113_xor0 ^ s_dadda_pg_rca24_fa103_xor1;
  assign s_dadda_pg_rca24_fa113_and1 = s_dadda_pg_rca24_fa113_xor0 & s_dadda_pg_rca24_fa103_xor1;
  assign s_dadda_pg_rca24_fa113_or0 = s_dadda_pg_rca24_fa113_and0 | s_dadda_pg_rca24_fa113_and1;
  assign s_dadda_pg_rca24_fa114_xor0 = s_dadda_pg_rca24_fa104_xor1 ^ s_dadda_pg_rca24_fa105_xor1;
  assign s_dadda_pg_rca24_fa114_and0 = s_dadda_pg_rca24_fa104_xor1 & s_dadda_pg_rca24_fa105_xor1;
  assign s_dadda_pg_rca24_fa114_xor1 = s_dadda_pg_rca24_fa114_xor0 ^ s_dadda_pg_rca24_fa106_xor1;
  assign s_dadda_pg_rca24_fa114_and1 = s_dadda_pg_rca24_fa114_xor0 & s_dadda_pg_rca24_fa106_xor1;
  assign s_dadda_pg_rca24_fa114_or0 = s_dadda_pg_rca24_fa114_and0 | s_dadda_pg_rca24_fa114_and1;
  assign s_dadda_pg_rca24_fa115_xor0 = s_dadda_pg_rca24_fa107_xor1 ^ s_dadda_pg_rca24_fa108_xor1;
  assign s_dadda_pg_rca24_fa115_and0 = s_dadda_pg_rca24_fa107_xor1 & s_dadda_pg_rca24_fa108_xor1;
  assign s_dadda_pg_rca24_fa115_xor1 = s_dadda_pg_rca24_fa115_xor0 ^ s_dadda_pg_rca24_fa109_xor1;
  assign s_dadda_pg_rca24_fa115_and1 = s_dadda_pg_rca24_fa115_xor0 & s_dadda_pg_rca24_fa109_xor1;
  assign s_dadda_pg_rca24_fa115_or0 = s_dadda_pg_rca24_fa115_and0 | s_dadda_pg_rca24_fa115_and1;
  assign s_dadda_pg_rca24_fa116_xor0 = s_dadda_pg_rca24_fa115_or0 ^ s_dadda_pg_rca24_fa114_or0;
  assign s_dadda_pg_rca24_fa116_and0 = s_dadda_pg_rca24_fa115_or0 & s_dadda_pg_rca24_fa114_or0;
  assign s_dadda_pg_rca24_fa116_xor1 = s_dadda_pg_rca24_fa116_xor0 ^ s_dadda_pg_rca24_fa113_or0;
  assign s_dadda_pg_rca24_fa116_and1 = s_dadda_pg_rca24_fa116_xor0 & s_dadda_pg_rca24_fa113_or0;
  assign s_dadda_pg_rca24_fa116_or0 = s_dadda_pg_rca24_fa116_and0 | s_dadda_pg_rca24_fa116_and1;
  assign s_dadda_pg_rca24_fa117_xor0 = s_dadda_pg_rca24_fa112_or0 ^ s_dadda_pg_rca24_fa111_or0;
  assign s_dadda_pg_rca24_fa117_and0 = s_dadda_pg_rca24_fa112_or0 & s_dadda_pg_rca24_fa111_or0;
  assign s_dadda_pg_rca24_fa117_xor1 = s_dadda_pg_rca24_fa117_xor0 ^ s_dadda_pg_rca24_fa110_or0;
  assign s_dadda_pg_rca24_fa117_and1 = s_dadda_pg_rca24_fa117_xor0 & s_dadda_pg_rca24_fa110_or0;
  assign s_dadda_pg_rca24_fa117_or0 = s_dadda_pg_rca24_fa117_and0 | s_dadda_pg_rca24_fa117_and1;
  assign s_dadda_pg_rca24_fa118_xor0 = s_dadda_pg_rca24_fa109_or0 ^ s_dadda_pg_rca24_fa108_or0;
  assign s_dadda_pg_rca24_fa118_and0 = s_dadda_pg_rca24_fa109_or0 & s_dadda_pg_rca24_fa108_or0;
  assign s_dadda_pg_rca24_fa118_xor1 = s_dadda_pg_rca24_fa118_xor0 ^ s_dadda_pg_rca24_fa107_or0;
  assign s_dadda_pg_rca24_fa118_and1 = s_dadda_pg_rca24_fa118_xor0 & s_dadda_pg_rca24_fa107_or0;
  assign s_dadda_pg_rca24_fa118_or0 = s_dadda_pg_rca24_fa118_and0 | s_dadda_pg_rca24_fa118_and1;
  assign s_dadda_pg_rca24_fa119_xor0 = s_dadda_pg_rca24_fa106_or0 ^ s_dadda_pg_rca24_fa105_or0;
  assign s_dadda_pg_rca24_fa119_and0 = s_dadda_pg_rca24_fa106_or0 & s_dadda_pg_rca24_fa105_or0;
  assign s_dadda_pg_rca24_fa119_xor1 = s_dadda_pg_rca24_fa119_xor0 ^ s_dadda_pg_rca24_fa104_or0;
  assign s_dadda_pg_rca24_fa119_and1 = s_dadda_pg_rca24_fa119_xor0 & s_dadda_pg_rca24_fa104_or0;
  assign s_dadda_pg_rca24_fa119_or0 = s_dadda_pg_rca24_fa119_and0 | s_dadda_pg_rca24_fa119_and1;
  assign s_dadda_pg_rca24_and_16_4 = a[16] & b[4];
  assign s_dadda_pg_rca24_and_15_5 = a[15] & b[5];
  assign s_dadda_pg_rca24_fa120_xor0 = s_dadda_pg_rca24_fa103_or0 ^ s_dadda_pg_rca24_and_16_4;
  assign s_dadda_pg_rca24_fa120_and0 = s_dadda_pg_rca24_fa103_or0 & s_dadda_pg_rca24_and_16_4;
  assign s_dadda_pg_rca24_fa120_xor1 = s_dadda_pg_rca24_fa120_xor0 ^ s_dadda_pg_rca24_and_15_5;
  assign s_dadda_pg_rca24_fa120_and1 = s_dadda_pg_rca24_fa120_xor0 & s_dadda_pg_rca24_and_15_5;
  assign s_dadda_pg_rca24_fa120_or0 = s_dadda_pg_rca24_fa120_and0 | s_dadda_pg_rca24_fa120_and1;
  assign s_dadda_pg_rca24_and_14_6 = a[14] & b[6];
  assign s_dadda_pg_rca24_and_13_7 = a[13] & b[7];
  assign s_dadda_pg_rca24_and_12_8 = a[12] & b[8];
  assign s_dadda_pg_rca24_fa121_xor0 = s_dadda_pg_rca24_and_14_6 ^ s_dadda_pg_rca24_and_13_7;
  assign s_dadda_pg_rca24_fa121_and0 = s_dadda_pg_rca24_and_14_6 & s_dadda_pg_rca24_and_13_7;
  assign s_dadda_pg_rca24_fa121_xor1 = s_dadda_pg_rca24_fa121_xor0 ^ s_dadda_pg_rca24_and_12_8;
  assign s_dadda_pg_rca24_fa121_and1 = s_dadda_pg_rca24_fa121_xor0 & s_dadda_pg_rca24_and_12_8;
  assign s_dadda_pg_rca24_fa121_or0 = s_dadda_pg_rca24_fa121_and0 | s_dadda_pg_rca24_fa121_and1;
  assign s_dadda_pg_rca24_and_11_9 = a[11] & b[9];
  assign s_dadda_pg_rca24_and_10_10 = a[10] & b[10];
  assign s_dadda_pg_rca24_and_9_11 = a[9] & b[11];
  assign s_dadda_pg_rca24_fa122_xor0 = s_dadda_pg_rca24_and_11_9 ^ s_dadda_pg_rca24_and_10_10;
  assign s_dadda_pg_rca24_fa122_and0 = s_dadda_pg_rca24_and_11_9 & s_dadda_pg_rca24_and_10_10;
  assign s_dadda_pg_rca24_fa122_xor1 = s_dadda_pg_rca24_fa122_xor0 ^ s_dadda_pg_rca24_and_9_11;
  assign s_dadda_pg_rca24_fa122_and1 = s_dadda_pg_rca24_fa122_xor0 & s_dadda_pg_rca24_and_9_11;
  assign s_dadda_pg_rca24_fa122_or0 = s_dadda_pg_rca24_fa122_and0 | s_dadda_pg_rca24_fa122_and1;
  assign s_dadda_pg_rca24_and_8_12 = a[8] & b[12];
  assign s_dadda_pg_rca24_and_7_13 = a[7] & b[13];
  assign s_dadda_pg_rca24_and_6_14 = a[6] & b[14];
  assign s_dadda_pg_rca24_fa123_xor0 = s_dadda_pg_rca24_and_8_12 ^ s_dadda_pg_rca24_and_7_13;
  assign s_dadda_pg_rca24_fa123_and0 = s_dadda_pg_rca24_and_8_12 & s_dadda_pg_rca24_and_7_13;
  assign s_dadda_pg_rca24_fa123_xor1 = s_dadda_pg_rca24_fa123_xor0 ^ s_dadda_pg_rca24_and_6_14;
  assign s_dadda_pg_rca24_fa123_and1 = s_dadda_pg_rca24_fa123_xor0 & s_dadda_pg_rca24_and_6_14;
  assign s_dadda_pg_rca24_fa123_or0 = s_dadda_pg_rca24_fa123_and0 | s_dadda_pg_rca24_fa123_and1;
  assign s_dadda_pg_rca24_and_5_15 = a[5] & b[15];
  assign s_dadda_pg_rca24_and_4_16 = a[4] & b[16];
  assign s_dadda_pg_rca24_and_3_17 = a[3] & b[17];
  assign s_dadda_pg_rca24_fa124_xor0 = s_dadda_pg_rca24_and_5_15 ^ s_dadda_pg_rca24_and_4_16;
  assign s_dadda_pg_rca24_fa124_and0 = s_dadda_pg_rca24_and_5_15 & s_dadda_pg_rca24_and_4_16;
  assign s_dadda_pg_rca24_fa124_xor1 = s_dadda_pg_rca24_fa124_xor0 ^ s_dadda_pg_rca24_and_3_17;
  assign s_dadda_pg_rca24_fa124_and1 = s_dadda_pg_rca24_fa124_xor0 & s_dadda_pg_rca24_and_3_17;
  assign s_dadda_pg_rca24_fa124_or0 = s_dadda_pg_rca24_fa124_and0 | s_dadda_pg_rca24_fa124_and1;
  assign s_dadda_pg_rca24_and_2_18 = a[2] & b[18];
  assign s_dadda_pg_rca24_and_1_19 = a[1] & b[19];
  assign s_dadda_pg_rca24_and_0_20 = a[0] & b[20];
  assign s_dadda_pg_rca24_fa125_xor0 = s_dadda_pg_rca24_and_2_18 ^ s_dadda_pg_rca24_and_1_19;
  assign s_dadda_pg_rca24_fa125_and0 = s_dadda_pg_rca24_and_2_18 & s_dadda_pg_rca24_and_1_19;
  assign s_dadda_pg_rca24_fa125_xor1 = s_dadda_pg_rca24_fa125_xor0 ^ s_dadda_pg_rca24_and_0_20;
  assign s_dadda_pg_rca24_fa125_and1 = s_dadda_pg_rca24_fa125_xor0 & s_dadda_pg_rca24_and_0_20;
  assign s_dadda_pg_rca24_fa125_or0 = s_dadda_pg_rca24_fa125_and0 | s_dadda_pg_rca24_fa125_and1;
  assign s_dadda_pg_rca24_fa126_xor0 = s_dadda_pg_rca24_fa0_xor1 ^ s_dadda_pg_rca24_ha1_xor0;
  assign s_dadda_pg_rca24_fa126_and0 = s_dadda_pg_rca24_fa0_xor1 & s_dadda_pg_rca24_ha1_xor0;
  assign s_dadda_pg_rca24_fa126_xor1 = s_dadda_pg_rca24_fa126_xor0 ^ s_dadda_pg_rca24_fa116_xor1;
  assign s_dadda_pg_rca24_fa126_and1 = s_dadda_pg_rca24_fa126_xor0 & s_dadda_pg_rca24_fa116_xor1;
  assign s_dadda_pg_rca24_fa126_or0 = s_dadda_pg_rca24_fa126_and0 | s_dadda_pg_rca24_fa126_and1;
  assign s_dadda_pg_rca24_fa127_xor0 = s_dadda_pg_rca24_fa117_xor1 ^ s_dadda_pg_rca24_fa118_xor1;
  assign s_dadda_pg_rca24_fa127_and0 = s_dadda_pg_rca24_fa117_xor1 & s_dadda_pg_rca24_fa118_xor1;
  assign s_dadda_pg_rca24_fa127_xor1 = s_dadda_pg_rca24_fa127_xor0 ^ s_dadda_pg_rca24_fa119_xor1;
  assign s_dadda_pg_rca24_fa127_and1 = s_dadda_pg_rca24_fa127_xor0 & s_dadda_pg_rca24_fa119_xor1;
  assign s_dadda_pg_rca24_fa127_or0 = s_dadda_pg_rca24_fa127_and0 | s_dadda_pg_rca24_fa127_and1;
  assign s_dadda_pg_rca24_fa128_xor0 = s_dadda_pg_rca24_fa120_xor1 ^ s_dadda_pg_rca24_fa121_xor1;
  assign s_dadda_pg_rca24_fa128_and0 = s_dadda_pg_rca24_fa120_xor1 & s_dadda_pg_rca24_fa121_xor1;
  assign s_dadda_pg_rca24_fa128_xor1 = s_dadda_pg_rca24_fa128_xor0 ^ s_dadda_pg_rca24_fa122_xor1;
  assign s_dadda_pg_rca24_fa128_and1 = s_dadda_pg_rca24_fa128_xor0 & s_dadda_pg_rca24_fa122_xor1;
  assign s_dadda_pg_rca24_fa128_or0 = s_dadda_pg_rca24_fa128_and0 | s_dadda_pg_rca24_fa128_and1;
  assign s_dadda_pg_rca24_fa129_xor0 = s_dadda_pg_rca24_fa128_or0 ^ s_dadda_pg_rca24_fa127_or0;
  assign s_dadda_pg_rca24_fa129_and0 = s_dadda_pg_rca24_fa128_or0 & s_dadda_pg_rca24_fa127_or0;
  assign s_dadda_pg_rca24_fa129_xor1 = s_dadda_pg_rca24_fa129_xor0 ^ s_dadda_pg_rca24_fa126_or0;
  assign s_dadda_pg_rca24_fa129_and1 = s_dadda_pg_rca24_fa129_xor0 & s_dadda_pg_rca24_fa126_or0;
  assign s_dadda_pg_rca24_fa129_or0 = s_dadda_pg_rca24_fa129_and0 | s_dadda_pg_rca24_fa129_and1;
  assign s_dadda_pg_rca24_fa130_xor0 = s_dadda_pg_rca24_fa125_or0 ^ s_dadda_pg_rca24_fa124_or0;
  assign s_dadda_pg_rca24_fa130_and0 = s_dadda_pg_rca24_fa125_or0 & s_dadda_pg_rca24_fa124_or0;
  assign s_dadda_pg_rca24_fa130_xor1 = s_dadda_pg_rca24_fa130_xor0 ^ s_dadda_pg_rca24_fa123_or0;
  assign s_dadda_pg_rca24_fa130_and1 = s_dadda_pg_rca24_fa130_xor0 & s_dadda_pg_rca24_fa123_or0;
  assign s_dadda_pg_rca24_fa130_or0 = s_dadda_pg_rca24_fa130_and0 | s_dadda_pg_rca24_fa130_and1;
  assign s_dadda_pg_rca24_fa131_xor0 = s_dadda_pg_rca24_fa122_or0 ^ s_dadda_pg_rca24_fa121_or0;
  assign s_dadda_pg_rca24_fa131_and0 = s_dadda_pg_rca24_fa122_or0 & s_dadda_pg_rca24_fa121_or0;
  assign s_dadda_pg_rca24_fa131_xor1 = s_dadda_pg_rca24_fa131_xor0 ^ s_dadda_pg_rca24_fa120_or0;
  assign s_dadda_pg_rca24_fa131_and1 = s_dadda_pg_rca24_fa131_xor0 & s_dadda_pg_rca24_fa120_or0;
  assign s_dadda_pg_rca24_fa131_or0 = s_dadda_pg_rca24_fa131_and0 | s_dadda_pg_rca24_fa131_and1;
  assign s_dadda_pg_rca24_fa132_xor0 = s_dadda_pg_rca24_fa119_or0 ^ s_dadda_pg_rca24_fa118_or0;
  assign s_dadda_pg_rca24_fa132_and0 = s_dadda_pg_rca24_fa119_or0 & s_dadda_pg_rca24_fa118_or0;
  assign s_dadda_pg_rca24_fa132_xor1 = s_dadda_pg_rca24_fa132_xor0 ^ s_dadda_pg_rca24_fa117_or0;
  assign s_dadda_pg_rca24_fa132_and1 = s_dadda_pg_rca24_fa132_xor0 & s_dadda_pg_rca24_fa117_or0;
  assign s_dadda_pg_rca24_fa132_or0 = s_dadda_pg_rca24_fa132_and0 | s_dadda_pg_rca24_fa132_and1;
  assign s_dadda_pg_rca24_and_15_6 = a[15] & b[6];
  assign s_dadda_pg_rca24_and_14_7 = a[14] & b[7];
  assign s_dadda_pg_rca24_fa133_xor0 = s_dadda_pg_rca24_fa116_or0 ^ s_dadda_pg_rca24_and_15_6;
  assign s_dadda_pg_rca24_fa133_and0 = s_dadda_pg_rca24_fa116_or0 & s_dadda_pg_rca24_and_15_6;
  assign s_dadda_pg_rca24_fa133_xor1 = s_dadda_pg_rca24_fa133_xor0 ^ s_dadda_pg_rca24_and_14_7;
  assign s_dadda_pg_rca24_fa133_and1 = s_dadda_pg_rca24_fa133_xor0 & s_dadda_pg_rca24_and_14_7;
  assign s_dadda_pg_rca24_fa133_or0 = s_dadda_pg_rca24_fa133_and0 | s_dadda_pg_rca24_fa133_and1;
  assign s_dadda_pg_rca24_and_13_8 = a[13] & b[8];
  assign s_dadda_pg_rca24_and_12_9 = a[12] & b[9];
  assign s_dadda_pg_rca24_and_11_10 = a[11] & b[10];
  assign s_dadda_pg_rca24_fa134_xor0 = s_dadda_pg_rca24_and_13_8 ^ s_dadda_pg_rca24_and_12_9;
  assign s_dadda_pg_rca24_fa134_and0 = s_dadda_pg_rca24_and_13_8 & s_dadda_pg_rca24_and_12_9;
  assign s_dadda_pg_rca24_fa134_xor1 = s_dadda_pg_rca24_fa134_xor0 ^ s_dadda_pg_rca24_and_11_10;
  assign s_dadda_pg_rca24_fa134_and1 = s_dadda_pg_rca24_fa134_xor0 & s_dadda_pg_rca24_and_11_10;
  assign s_dadda_pg_rca24_fa134_or0 = s_dadda_pg_rca24_fa134_and0 | s_dadda_pg_rca24_fa134_and1;
  assign s_dadda_pg_rca24_and_10_11 = a[10] & b[11];
  assign s_dadda_pg_rca24_and_9_12 = a[9] & b[12];
  assign s_dadda_pg_rca24_and_8_13 = a[8] & b[13];
  assign s_dadda_pg_rca24_fa135_xor0 = s_dadda_pg_rca24_and_10_11 ^ s_dadda_pg_rca24_and_9_12;
  assign s_dadda_pg_rca24_fa135_and0 = s_dadda_pg_rca24_and_10_11 & s_dadda_pg_rca24_and_9_12;
  assign s_dadda_pg_rca24_fa135_xor1 = s_dadda_pg_rca24_fa135_xor0 ^ s_dadda_pg_rca24_and_8_13;
  assign s_dadda_pg_rca24_fa135_and1 = s_dadda_pg_rca24_fa135_xor0 & s_dadda_pg_rca24_and_8_13;
  assign s_dadda_pg_rca24_fa135_or0 = s_dadda_pg_rca24_fa135_and0 | s_dadda_pg_rca24_fa135_and1;
  assign s_dadda_pg_rca24_and_7_14 = a[7] & b[14];
  assign s_dadda_pg_rca24_and_6_15 = a[6] & b[15];
  assign s_dadda_pg_rca24_and_5_16 = a[5] & b[16];
  assign s_dadda_pg_rca24_fa136_xor0 = s_dadda_pg_rca24_and_7_14 ^ s_dadda_pg_rca24_and_6_15;
  assign s_dadda_pg_rca24_fa136_and0 = s_dadda_pg_rca24_and_7_14 & s_dadda_pg_rca24_and_6_15;
  assign s_dadda_pg_rca24_fa136_xor1 = s_dadda_pg_rca24_fa136_xor0 ^ s_dadda_pg_rca24_and_5_16;
  assign s_dadda_pg_rca24_fa136_and1 = s_dadda_pg_rca24_fa136_xor0 & s_dadda_pg_rca24_and_5_16;
  assign s_dadda_pg_rca24_fa136_or0 = s_dadda_pg_rca24_fa136_and0 | s_dadda_pg_rca24_fa136_and1;
  assign s_dadda_pg_rca24_and_4_17 = a[4] & b[17];
  assign s_dadda_pg_rca24_and_3_18 = a[3] & b[18];
  assign s_dadda_pg_rca24_and_2_19 = a[2] & b[19];
  assign s_dadda_pg_rca24_fa137_xor0 = s_dadda_pg_rca24_and_4_17 ^ s_dadda_pg_rca24_and_3_18;
  assign s_dadda_pg_rca24_fa137_and0 = s_dadda_pg_rca24_and_4_17 & s_dadda_pg_rca24_and_3_18;
  assign s_dadda_pg_rca24_fa137_xor1 = s_dadda_pg_rca24_fa137_xor0 ^ s_dadda_pg_rca24_and_2_19;
  assign s_dadda_pg_rca24_fa137_and1 = s_dadda_pg_rca24_fa137_xor0 & s_dadda_pg_rca24_and_2_19;
  assign s_dadda_pg_rca24_fa137_or0 = s_dadda_pg_rca24_fa137_and0 | s_dadda_pg_rca24_fa137_and1;
  assign s_dadda_pg_rca24_and_1_20 = a[1] & b[20];
  assign s_dadda_pg_rca24_and_0_21 = a[0] & b[21];
  assign s_dadda_pg_rca24_fa138_xor0 = s_dadda_pg_rca24_and_1_20 ^ s_dadda_pg_rca24_and_0_21;
  assign s_dadda_pg_rca24_fa138_and0 = s_dadda_pg_rca24_and_1_20 & s_dadda_pg_rca24_and_0_21;
  assign s_dadda_pg_rca24_fa138_xor1 = s_dadda_pg_rca24_fa138_xor0 ^ s_dadda_pg_rca24_fa1_xor1;
  assign s_dadda_pg_rca24_fa138_and1 = s_dadda_pg_rca24_fa138_xor0 & s_dadda_pg_rca24_fa1_xor1;
  assign s_dadda_pg_rca24_fa138_or0 = s_dadda_pg_rca24_fa138_and0 | s_dadda_pg_rca24_fa138_and1;
  assign s_dadda_pg_rca24_fa139_xor0 = s_dadda_pg_rca24_fa2_xor1 ^ s_dadda_pg_rca24_ha2_xor0;
  assign s_dadda_pg_rca24_fa139_and0 = s_dadda_pg_rca24_fa2_xor1 & s_dadda_pg_rca24_ha2_xor0;
  assign s_dadda_pg_rca24_fa139_xor1 = s_dadda_pg_rca24_fa139_xor0 ^ s_dadda_pg_rca24_fa129_xor1;
  assign s_dadda_pg_rca24_fa139_and1 = s_dadda_pg_rca24_fa139_xor0 & s_dadda_pg_rca24_fa129_xor1;
  assign s_dadda_pg_rca24_fa139_or0 = s_dadda_pg_rca24_fa139_and0 | s_dadda_pg_rca24_fa139_and1;
  assign s_dadda_pg_rca24_fa140_xor0 = s_dadda_pg_rca24_fa130_xor1 ^ s_dadda_pg_rca24_fa131_xor1;
  assign s_dadda_pg_rca24_fa140_and0 = s_dadda_pg_rca24_fa130_xor1 & s_dadda_pg_rca24_fa131_xor1;
  assign s_dadda_pg_rca24_fa140_xor1 = s_dadda_pg_rca24_fa140_xor0 ^ s_dadda_pg_rca24_fa132_xor1;
  assign s_dadda_pg_rca24_fa140_and1 = s_dadda_pg_rca24_fa140_xor0 & s_dadda_pg_rca24_fa132_xor1;
  assign s_dadda_pg_rca24_fa140_or0 = s_dadda_pg_rca24_fa140_and0 | s_dadda_pg_rca24_fa140_and1;
  assign s_dadda_pg_rca24_fa141_xor0 = s_dadda_pg_rca24_fa133_xor1 ^ s_dadda_pg_rca24_fa134_xor1;
  assign s_dadda_pg_rca24_fa141_and0 = s_dadda_pg_rca24_fa133_xor1 & s_dadda_pg_rca24_fa134_xor1;
  assign s_dadda_pg_rca24_fa141_xor1 = s_dadda_pg_rca24_fa141_xor0 ^ s_dadda_pg_rca24_fa135_xor1;
  assign s_dadda_pg_rca24_fa141_and1 = s_dadda_pg_rca24_fa141_xor0 & s_dadda_pg_rca24_fa135_xor1;
  assign s_dadda_pg_rca24_fa141_or0 = s_dadda_pg_rca24_fa141_and0 | s_dadda_pg_rca24_fa141_and1;
  assign s_dadda_pg_rca24_fa142_xor0 = s_dadda_pg_rca24_fa141_or0 ^ s_dadda_pg_rca24_fa140_or0;
  assign s_dadda_pg_rca24_fa142_and0 = s_dadda_pg_rca24_fa141_or0 & s_dadda_pg_rca24_fa140_or0;
  assign s_dadda_pg_rca24_fa142_xor1 = s_dadda_pg_rca24_fa142_xor0 ^ s_dadda_pg_rca24_fa139_or0;
  assign s_dadda_pg_rca24_fa142_and1 = s_dadda_pg_rca24_fa142_xor0 & s_dadda_pg_rca24_fa139_or0;
  assign s_dadda_pg_rca24_fa142_or0 = s_dadda_pg_rca24_fa142_and0 | s_dadda_pg_rca24_fa142_and1;
  assign s_dadda_pg_rca24_fa143_xor0 = s_dadda_pg_rca24_fa138_or0 ^ s_dadda_pg_rca24_fa137_or0;
  assign s_dadda_pg_rca24_fa143_and0 = s_dadda_pg_rca24_fa138_or0 & s_dadda_pg_rca24_fa137_or0;
  assign s_dadda_pg_rca24_fa143_xor1 = s_dadda_pg_rca24_fa143_xor0 ^ s_dadda_pg_rca24_fa136_or0;
  assign s_dadda_pg_rca24_fa143_and1 = s_dadda_pg_rca24_fa143_xor0 & s_dadda_pg_rca24_fa136_or0;
  assign s_dadda_pg_rca24_fa143_or0 = s_dadda_pg_rca24_fa143_and0 | s_dadda_pg_rca24_fa143_and1;
  assign s_dadda_pg_rca24_fa144_xor0 = s_dadda_pg_rca24_fa135_or0 ^ s_dadda_pg_rca24_fa134_or0;
  assign s_dadda_pg_rca24_fa144_and0 = s_dadda_pg_rca24_fa135_or0 & s_dadda_pg_rca24_fa134_or0;
  assign s_dadda_pg_rca24_fa144_xor1 = s_dadda_pg_rca24_fa144_xor0 ^ s_dadda_pg_rca24_fa133_or0;
  assign s_dadda_pg_rca24_fa144_and1 = s_dadda_pg_rca24_fa144_xor0 & s_dadda_pg_rca24_fa133_or0;
  assign s_dadda_pg_rca24_fa144_or0 = s_dadda_pg_rca24_fa144_and0 | s_dadda_pg_rca24_fa144_and1;
  assign s_dadda_pg_rca24_fa145_xor0 = s_dadda_pg_rca24_fa132_or0 ^ s_dadda_pg_rca24_fa131_or0;
  assign s_dadda_pg_rca24_fa145_and0 = s_dadda_pg_rca24_fa132_or0 & s_dadda_pg_rca24_fa131_or0;
  assign s_dadda_pg_rca24_fa145_xor1 = s_dadda_pg_rca24_fa145_xor0 ^ s_dadda_pg_rca24_fa130_or0;
  assign s_dadda_pg_rca24_fa145_and1 = s_dadda_pg_rca24_fa145_xor0 & s_dadda_pg_rca24_fa130_or0;
  assign s_dadda_pg_rca24_fa145_or0 = s_dadda_pg_rca24_fa145_and0 | s_dadda_pg_rca24_fa145_and1;
  assign s_dadda_pg_rca24_and_14_8 = a[14] & b[8];
  assign s_dadda_pg_rca24_and_13_9 = a[13] & b[9];
  assign s_dadda_pg_rca24_fa146_xor0 = s_dadda_pg_rca24_fa129_or0 ^ s_dadda_pg_rca24_and_14_8;
  assign s_dadda_pg_rca24_fa146_and0 = s_dadda_pg_rca24_fa129_or0 & s_dadda_pg_rca24_and_14_8;
  assign s_dadda_pg_rca24_fa146_xor1 = s_dadda_pg_rca24_fa146_xor0 ^ s_dadda_pg_rca24_and_13_9;
  assign s_dadda_pg_rca24_fa146_and1 = s_dadda_pg_rca24_fa146_xor0 & s_dadda_pg_rca24_and_13_9;
  assign s_dadda_pg_rca24_fa146_or0 = s_dadda_pg_rca24_fa146_and0 | s_dadda_pg_rca24_fa146_and1;
  assign s_dadda_pg_rca24_and_12_10 = a[12] & b[10];
  assign s_dadda_pg_rca24_and_11_11 = a[11] & b[11];
  assign s_dadda_pg_rca24_and_10_12 = a[10] & b[12];
  assign s_dadda_pg_rca24_fa147_xor0 = s_dadda_pg_rca24_and_12_10 ^ s_dadda_pg_rca24_and_11_11;
  assign s_dadda_pg_rca24_fa147_and0 = s_dadda_pg_rca24_and_12_10 & s_dadda_pg_rca24_and_11_11;
  assign s_dadda_pg_rca24_fa147_xor1 = s_dadda_pg_rca24_fa147_xor0 ^ s_dadda_pg_rca24_and_10_12;
  assign s_dadda_pg_rca24_fa147_and1 = s_dadda_pg_rca24_fa147_xor0 & s_dadda_pg_rca24_and_10_12;
  assign s_dadda_pg_rca24_fa147_or0 = s_dadda_pg_rca24_fa147_and0 | s_dadda_pg_rca24_fa147_and1;
  assign s_dadda_pg_rca24_and_9_13 = a[9] & b[13];
  assign s_dadda_pg_rca24_and_8_14 = a[8] & b[14];
  assign s_dadda_pg_rca24_and_7_15 = a[7] & b[15];
  assign s_dadda_pg_rca24_fa148_xor0 = s_dadda_pg_rca24_and_9_13 ^ s_dadda_pg_rca24_and_8_14;
  assign s_dadda_pg_rca24_fa148_and0 = s_dadda_pg_rca24_and_9_13 & s_dadda_pg_rca24_and_8_14;
  assign s_dadda_pg_rca24_fa148_xor1 = s_dadda_pg_rca24_fa148_xor0 ^ s_dadda_pg_rca24_and_7_15;
  assign s_dadda_pg_rca24_fa148_and1 = s_dadda_pg_rca24_fa148_xor0 & s_dadda_pg_rca24_and_7_15;
  assign s_dadda_pg_rca24_fa148_or0 = s_dadda_pg_rca24_fa148_and0 | s_dadda_pg_rca24_fa148_and1;
  assign s_dadda_pg_rca24_and_6_16 = a[6] & b[16];
  assign s_dadda_pg_rca24_and_5_17 = a[5] & b[17];
  assign s_dadda_pg_rca24_and_4_18 = a[4] & b[18];
  assign s_dadda_pg_rca24_fa149_xor0 = s_dadda_pg_rca24_and_6_16 ^ s_dadda_pg_rca24_and_5_17;
  assign s_dadda_pg_rca24_fa149_and0 = s_dadda_pg_rca24_and_6_16 & s_dadda_pg_rca24_and_5_17;
  assign s_dadda_pg_rca24_fa149_xor1 = s_dadda_pg_rca24_fa149_xor0 ^ s_dadda_pg_rca24_and_4_18;
  assign s_dadda_pg_rca24_fa149_and1 = s_dadda_pg_rca24_fa149_xor0 & s_dadda_pg_rca24_and_4_18;
  assign s_dadda_pg_rca24_fa149_or0 = s_dadda_pg_rca24_fa149_and0 | s_dadda_pg_rca24_fa149_and1;
  assign s_dadda_pg_rca24_and_3_19 = a[3] & b[19];
  assign s_dadda_pg_rca24_and_2_20 = a[2] & b[20];
  assign s_dadda_pg_rca24_and_1_21 = a[1] & b[21];
  assign s_dadda_pg_rca24_fa150_xor0 = s_dadda_pg_rca24_and_3_19 ^ s_dadda_pg_rca24_and_2_20;
  assign s_dadda_pg_rca24_fa150_and0 = s_dadda_pg_rca24_and_3_19 & s_dadda_pg_rca24_and_2_20;
  assign s_dadda_pg_rca24_fa150_xor1 = s_dadda_pg_rca24_fa150_xor0 ^ s_dadda_pg_rca24_and_1_21;
  assign s_dadda_pg_rca24_fa150_and1 = s_dadda_pg_rca24_fa150_xor0 & s_dadda_pg_rca24_and_1_21;
  assign s_dadda_pg_rca24_fa150_or0 = s_dadda_pg_rca24_fa150_and0 | s_dadda_pg_rca24_fa150_and1;
  assign s_dadda_pg_rca24_and_0_22 = a[0] & b[22];
  assign s_dadda_pg_rca24_fa151_xor0 = s_dadda_pg_rca24_and_0_22 ^ s_dadda_pg_rca24_fa3_xor1;
  assign s_dadda_pg_rca24_fa151_and0 = s_dadda_pg_rca24_and_0_22 & s_dadda_pg_rca24_fa3_xor1;
  assign s_dadda_pg_rca24_fa151_xor1 = s_dadda_pg_rca24_fa151_xor0 ^ s_dadda_pg_rca24_fa4_xor1;
  assign s_dadda_pg_rca24_fa151_and1 = s_dadda_pg_rca24_fa151_xor0 & s_dadda_pg_rca24_fa4_xor1;
  assign s_dadda_pg_rca24_fa151_or0 = s_dadda_pg_rca24_fa151_and0 | s_dadda_pg_rca24_fa151_and1;
  assign s_dadda_pg_rca24_fa152_xor0 = s_dadda_pg_rca24_fa5_xor1 ^ s_dadda_pg_rca24_ha3_xor0;
  assign s_dadda_pg_rca24_fa152_and0 = s_dadda_pg_rca24_fa5_xor1 & s_dadda_pg_rca24_ha3_xor0;
  assign s_dadda_pg_rca24_fa152_xor1 = s_dadda_pg_rca24_fa152_xor0 ^ s_dadda_pg_rca24_fa142_xor1;
  assign s_dadda_pg_rca24_fa152_and1 = s_dadda_pg_rca24_fa152_xor0 & s_dadda_pg_rca24_fa142_xor1;
  assign s_dadda_pg_rca24_fa152_or0 = s_dadda_pg_rca24_fa152_and0 | s_dadda_pg_rca24_fa152_and1;
  assign s_dadda_pg_rca24_fa153_xor0 = s_dadda_pg_rca24_fa143_xor1 ^ s_dadda_pg_rca24_fa144_xor1;
  assign s_dadda_pg_rca24_fa153_and0 = s_dadda_pg_rca24_fa143_xor1 & s_dadda_pg_rca24_fa144_xor1;
  assign s_dadda_pg_rca24_fa153_xor1 = s_dadda_pg_rca24_fa153_xor0 ^ s_dadda_pg_rca24_fa145_xor1;
  assign s_dadda_pg_rca24_fa153_and1 = s_dadda_pg_rca24_fa153_xor0 & s_dadda_pg_rca24_fa145_xor1;
  assign s_dadda_pg_rca24_fa153_or0 = s_dadda_pg_rca24_fa153_and0 | s_dadda_pg_rca24_fa153_and1;
  assign s_dadda_pg_rca24_fa154_xor0 = s_dadda_pg_rca24_fa146_xor1 ^ s_dadda_pg_rca24_fa147_xor1;
  assign s_dadda_pg_rca24_fa154_and0 = s_dadda_pg_rca24_fa146_xor1 & s_dadda_pg_rca24_fa147_xor1;
  assign s_dadda_pg_rca24_fa154_xor1 = s_dadda_pg_rca24_fa154_xor0 ^ s_dadda_pg_rca24_fa148_xor1;
  assign s_dadda_pg_rca24_fa154_and1 = s_dadda_pg_rca24_fa154_xor0 & s_dadda_pg_rca24_fa148_xor1;
  assign s_dadda_pg_rca24_fa154_or0 = s_dadda_pg_rca24_fa154_and0 | s_dadda_pg_rca24_fa154_and1;
  assign s_dadda_pg_rca24_fa155_xor0 = s_dadda_pg_rca24_fa154_or0 ^ s_dadda_pg_rca24_fa153_or0;
  assign s_dadda_pg_rca24_fa155_and0 = s_dadda_pg_rca24_fa154_or0 & s_dadda_pg_rca24_fa153_or0;
  assign s_dadda_pg_rca24_fa155_xor1 = s_dadda_pg_rca24_fa155_xor0 ^ s_dadda_pg_rca24_fa152_or0;
  assign s_dadda_pg_rca24_fa155_and1 = s_dadda_pg_rca24_fa155_xor0 & s_dadda_pg_rca24_fa152_or0;
  assign s_dadda_pg_rca24_fa155_or0 = s_dadda_pg_rca24_fa155_and0 | s_dadda_pg_rca24_fa155_and1;
  assign s_dadda_pg_rca24_fa156_xor0 = s_dadda_pg_rca24_fa151_or0 ^ s_dadda_pg_rca24_fa150_or0;
  assign s_dadda_pg_rca24_fa156_and0 = s_dadda_pg_rca24_fa151_or0 & s_dadda_pg_rca24_fa150_or0;
  assign s_dadda_pg_rca24_fa156_xor1 = s_dadda_pg_rca24_fa156_xor0 ^ s_dadda_pg_rca24_fa149_or0;
  assign s_dadda_pg_rca24_fa156_and1 = s_dadda_pg_rca24_fa156_xor0 & s_dadda_pg_rca24_fa149_or0;
  assign s_dadda_pg_rca24_fa156_or0 = s_dadda_pg_rca24_fa156_and0 | s_dadda_pg_rca24_fa156_and1;
  assign s_dadda_pg_rca24_fa157_xor0 = s_dadda_pg_rca24_fa148_or0 ^ s_dadda_pg_rca24_fa147_or0;
  assign s_dadda_pg_rca24_fa157_and0 = s_dadda_pg_rca24_fa148_or0 & s_dadda_pg_rca24_fa147_or0;
  assign s_dadda_pg_rca24_fa157_xor1 = s_dadda_pg_rca24_fa157_xor0 ^ s_dadda_pg_rca24_fa146_or0;
  assign s_dadda_pg_rca24_fa157_and1 = s_dadda_pg_rca24_fa157_xor0 & s_dadda_pg_rca24_fa146_or0;
  assign s_dadda_pg_rca24_fa157_or0 = s_dadda_pg_rca24_fa157_and0 | s_dadda_pg_rca24_fa157_and1;
  assign s_dadda_pg_rca24_fa158_xor0 = s_dadda_pg_rca24_fa145_or0 ^ s_dadda_pg_rca24_fa144_or0;
  assign s_dadda_pg_rca24_fa158_and0 = s_dadda_pg_rca24_fa145_or0 & s_dadda_pg_rca24_fa144_or0;
  assign s_dadda_pg_rca24_fa158_xor1 = s_dadda_pg_rca24_fa158_xor0 ^ s_dadda_pg_rca24_fa143_or0;
  assign s_dadda_pg_rca24_fa158_and1 = s_dadda_pg_rca24_fa158_xor0 & s_dadda_pg_rca24_fa143_or0;
  assign s_dadda_pg_rca24_fa158_or0 = s_dadda_pg_rca24_fa158_and0 | s_dadda_pg_rca24_fa158_and1;
  assign s_dadda_pg_rca24_and_13_10 = a[13] & b[10];
  assign s_dadda_pg_rca24_and_12_11 = a[12] & b[11];
  assign s_dadda_pg_rca24_fa159_xor0 = s_dadda_pg_rca24_fa142_or0 ^ s_dadda_pg_rca24_and_13_10;
  assign s_dadda_pg_rca24_fa159_and0 = s_dadda_pg_rca24_fa142_or0 & s_dadda_pg_rca24_and_13_10;
  assign s_dadda_pg_rca24_fa159_xor1 = s_dadda_pg_rca24_fa159_xor0 ^ s_dadda_pg_rca24_and_12_11;
  assign s_dadda_pg_rca24_fa159_and1 = s_dadda_pg_rca24_fa159_xor0 & s_dadda_pg_rca24_and_12_11;
  assign s_dadda_pg_rca24_fa159_or0 = s_dadda_pg_rca24_fa159_and0 | s_dadda_pg_rca24_fa159_and1;
  assign s_dadda_pg_rca24_and_11_12 = a[11] & b[12];
  assign s_dadda_pg_rca24_and_10_13 = a[10] & b[13];
  assign s_dadda_pg_rca24_and_9_14 = a[9] & b[14];
  assign s_dadda_pg_rca24_fa160_xor0 = s_dadda_pg_rca24_and_11_12 ^ s_dadda_pg_rca24_and_10_13;
  assign s_dadda_pg_rca24_fa160_and0 = s_dadda_pg_rca24_and_11_12 & s_dadda_pg_rca24_and_10_13;
  assign s_dadda_pg_rca24_fa160_xor1 = s_dadda_pg_rca24_fa160_xor0 ^ s_dadda_pg_rca24_and_9_14;
  assign s_dadda_pg_rca24_fa160_and1 = s_dadda_pg_rca24_fa160_xor0 & s_dadda_pg_rca24_and_9_14;
  assign s_dadda_pg_rca24_fa160_or0 = s_dadda_pg_rca24_fa160_and0 | s_dadda_pg_rca24_fa160_and1;
  assign s_dadda_pg_rca24_and_8_15 = a[8] & b[15];
  assign s_dadda_pg_rca24_and_7_16 = a[7] & b[16];
  assign s_dadda_pg_rca24_and_6_17 = a[6] & b[17];
  assign s_dadda_pg_rca24_fa161_xor0 = s_dadda_pg_rca24_and_8_15 ^ s_dadda_pg_rca24_and_7_16;
  assign s_dadda_pg_rca24_fa161_and0 = s_dadda_pg_rca24_and_8_15 & s_dadda_pg_rca24_and_7_16;
  assign s_dadda_pg_rca24_fa161_xor1 = s_dadda_pg_rca24_fa161_xor0 ^ s_dadda_pg_rca24_and_6_17;
  assign s_dadda_pg_rca24_fa161_and1 = s_dadda_pg_rca24_fa161_xor0 & s_dadda_pg_rca24_and_6_17;
  assign s_dadda_pg_rca24_fa161_or0 = s_dadda_pg_rca24_fa161_and0 | s_dadda_pg_rca24_fa161_and1;
  assign s_dadda_pg_rca24_and_5_18 = a[5] & b[18];
  assign s_dadda_pg_rca24_and_4_19 = a[4] & b[19];
  assign s_dadda_pg_rca24_and_3_20 = a[3] & b[20];
  assign s_dadda_pg_rca24_fa162_xor0 = s_dadda_pg_rca24_and_5_18 ^ s_dadda_pg_rca24_and_4_19;
  assign s_dadda_pg_rca24_fa162_and0 = s_dadda_pg_rca24_and_5_18 & s_dadda_pg_rca24_and_4_19;
  assign s_dadda_pg_rca24_fa162_xor1 = s_dadda_pg_rca24_fa162_xor0 ^ s_dadda_pg_rca24_and_3_20;
  assign s_dadda_pg_rca24_fa162_and1 = s_dadda_pg_rca24_fa162_xor0 & s_dadda_pg_rca24_and_3_20;
  assign s_dadda_pg_rca24_fa162_or0 = s_dadda_pg_rca24_fa162_and0 | s_dadda_pg_rca24_fa162_and1;
  assign s_dadda_pg_rca24_and_2_21 = a[2] & b[21];
  assign s_dadda_pg_rca24_and_1_22 = a[1] & b[22];
  assign s_dadda_pg_rca24_nand_0_23 = ~(a[0] & b[23]);
  assign s_dadda_pg_rca24_fa163_xor0 = s_dadda_pg_rca24_and_2_21 ^ s_dadda_pg_rca24_and_1_22;
  assign s_dadda_pg_rca24_fa163_and0 = s_dadda_pg_rca24_and_2_21 & s_dadda_pg_rca24_and_1_22;
  assign s_dadda_pg_rca24_fa163_xor1 = s_dadda_pg_rca24_fa163_xor0 ^ s_dadda_pg_rca24_nand_0_23;
  assign s_dadda_pg_rca24_fa163_and1 = s_dadda_pg_rca24_fa163_xor0 & s_dadda_pg_rca24_nand_0_23;
  assign s_dadda_pg_rca24_fa163_or0 = s_dadda_pg_rca24_fa163_and0 | s_dadda_pg_rca24_fa163_and1;
  assign s_dadda_pg_rca24_fa164_xor0 = s_dadda_pg_rca24_fa6_xor1 ^ s_dadda_pg_rca24_fa7_xor1;
  assign s_dadda_pg_rca24_fa164_and0 = s_dadda_pg_rca24_fa6_xor1 & s_dadda_pg_rca24_fa7_xor1;
  assign s_dadda_pg_rca24_fa164_xor1 = s_dadda_pg_rca24_fa164_xor0 ^ s_dadda_pg_rca24_fa8_xor1;
  assign s_dadda_pg_rca24_fa164_and1 = s_dadda_pg_rca24_fa164_xor0 & s_dadda_pg_rca24_fa8_xor1;
  assign s_dadda_pg_rca24_fa164_or0 = s_dadda_pg_rca24_fa164_and0 | s_dadda_pg_rca24_fa164_and1;
  assign s_dadda_pg_rca24_fa165_xor0 = s_dadda_pg_rca24_fa9_xor1 ^ s_dadda_pg_rca24_ha4_xor0;
  assign s_dadda_pg_rca24_fa165_and0 = s_dadda_pg_rca24_fa9_xor1 & s_dadda_pg_rca24_ha4_xor0;
  assign s_dadda_pg_rca24_fa165_xor1 = s_dadda_pg_rca24_fa165_xor0 ^ s_dadda_pg_rca24_fa155_xor1;
  assign s_dadda_pg_rca24_fa165_and1 = s_dadda_pg_rca24_fa165_xor0 & s_dadda_pg_rca24_fa155_xor1;
  assign s_dadda_pg_rca24_fa165_or0 = s_dadda_pg_rca24_fa165_and0 | s_dadda_pg_rca24_fa165_and1;
  assign s_dadda_pg_rca24_fa166_xor0 = s_dadda_pg_rca24_fa156_xor1 ^ s_dadda_pg_rca24_fa157_xor1;
  assign s_dadda_pg_rca24_fa166_and0 = s_dadda_pg_rca24_fa156_xor1 & s_dadda_pg_rca24_fa157_xor1;
  assign s_dadda_pg_rca24_fa166_xor1 = s_dadda_pg_rca24_fa166_xor0 ^ s_dadda_pg_rca24_fa158_xor1;
  assign s_dadda_pg_rca24_fa166_and1 = s_dadda_pg_rca24_fa166_xor0 & s_dadda_pg_rca24_fa158_xor1;
  assign s_dadda_pg_rca24_fa166_or0 = s_dadda_pg_rca24_fa166_and0 | s_dadda_pg_rca24_fa166_and1;
  assign s_dadda_pg_rca24_fa167_xor0 = s_dadda_pg_rca24_fa159_xor1 ^ s_dadda_pg_rca24_fa160_xor1;
  assign s_dadda_pg_rca24_fa167_and0 = s_dadda_pg_rca24_fa159_xor1 & s_dadda_pg_rca24_fa160_xor1;
  assign s_dadda_pg_rca24_fa167_xor1 = s_dadda_pg_rca24_fa167_xor0 ^ s_dadda_pg_rca24_fa161_xor1;
  assign s_dadda_pg_rca24_fa167_and1 = s_dadda_pg_rca24_fa167_xor0 & s_dadda_pg_rca24_fa161_xor1;
  assign s_dadda_pg_rca24_fa167_or0 = s_dadda_pg_rca24_fa167_and0 | s_dadda_pg_rca24_fa167_and1;
  assign s_dadda_pg_rca24_fa168_xor0 = s_dadda_pg_rca24_fa167_or0 ^ s_dadda_pg_rca24_fa166_or0;
  assign s_dadda_pg_rca24_fa168_and0 = s_dadda_pg_rca24_fa167_or0 & s_dadda_pg_rca24_fa166_or0;
  assign s_dadda_pg_rca24_fa168_xor1 = s_dadda_pg_rca24_fa168_xor0 ^ s_dadda_pg_rca24_fa165_or0;
  assign s_dadda_pg_rca24_fa168_and1 = s_dadda_pg_rca24_fa168_xor0 & s_dadda_pg_rca24_fa165_or0;
  assign s_dadda_pg_rca24_fa168_or0 = s_dadda_pg_rca24_fa168_and0 | s_dadda_pg_rca24_fa168_and1;
  assign s_dadda_pg_rca24_fa169_xor0 = s_dadda_pg_rca24_fa164_or0 ^ s_dadda_pg_rca24_fa163_or0;
  assign s_dadda_pg_rca24_fa169_and0 = s_dadda_pg_rca24_fa164_or0 & s_dadda_pg_rca24_fa163_or0;
  assign s_dadda_pg_rca24_fa169_xor1 = s_dadda_pg_rca24_fa169_xor0 ^ s_dadda_pg_rca24_fa162_or0;
  assign s_dadda_pg_rca24_fa169_and1 = s_dadda_pg_rca24_fa169_xor0 & s_dadda_pg_rca24_fa162_or0;
  assign s_dadda_pg_rca24_fa169_or0 = s_dadda_pg_rca24_fa169_and0 | s_dadda_pg_rca24_fa169_and1;
  assign s_dadda_pg_rca24_fa170_xor0 = s_dadda_pg_rca24_fa161_or0 ^ s_dadda_pg_rca24_fa160_or0;
  assign s_dadda_pg_rca24_fa170_and0 = s_dadda_pg_rca24_fa161_or0 & s_dadda_pg_rca24_fa160_or0;
  assign s_dadda_pg_rca24_fa170_xor1 = s_dadda_pg_rca24_fa170_xor0 ^ s_dadda_pg_rca24_fa159_or0;
  assign s_dadda_pg_rca24_fa170_and1 = s_dadda_pg_rca24_fa170_xor0 & s_dadda_pg_rca24_fa159_or0;
  assign s_dadda_pg_rca24_fa170_or0 = s_dadda_pg_rca24_fa170_and0 | s_dadda_pg_rca24_fa170_and1;
  assign s_dadda_pg_rca24_fa171_xor0 = s_dadda_pg_rca24_fa158_or0 ^ s_dadda_pg_rca24_fa157_or0;
  assign s_dadda_pg_rca24_fa171_and0 = s_dadda_pg_rca24_fa158_or0 & s_dadda_pg_rca24_fa157_or0;
  assign s_dadda_pg_rca24_fa171_xor1 = s_dadda_pg_rca24_fa171_xor0 ^ s_dadda_pg_rca24_fa156_or0;
  assign s_dadda_pg_rca24_fa171_and1 = s_dadda_pg_rca24_fa171_xor0 & s_dadda_pg_rca24_fa156_or0;
  assign s_dadda_pg_rca24_fa171_or0 = s_dadda_pg_rca24_fa171_and0 | s_dadda_pg_rca24_fa171_and1;
  assign s_dadda_pg_rca24_and_14_10 = a[14] & b[10];
  assign s_dadda_pg_rca24_and_13_11 = a[13] & b[11];
  assign s_dadda_pg_rca24_fa172_xor0 = s_dadda_pg_rca24_fa155_or0 ^ s_dadda_pg_rca24_and_14_10;
  assign s_dadda_pg_rca24_fa172_and0 = s_dadda_pg_rca24_fa155_or0 & s_dadda_pg_rca24_and_14_10;
  assign s_dadda_pg_rca24_fa172_xor1 = s_dadda_pg_rca24_fa172_xor0 ^ s_dadda_pg_rca24_and_13_11;
  assign s_dadda_pg_rca24_fa172_and1 = s_dadda_pg_rca24_fa172_xor0 & s_dadda_pg_rca24_and_13_11;
  assign s_dadda_pg_rca24_fa172_or0 = s_dadda_pg_rca24_fa172_and0 | s_dadda_pg_rca24_fa172_and1;
  assign s_dadda_pg_rca24_and_12_12 = a[12] & b[12];
  assign s_dadda_pg_rca24_and_11_13 = a[11] & b[13];
  assign s_dadda_pg_rca24_and_10_14 = a[10] & b[14];
  assign s_dadda_pg_rca24_fa173_xor0 = s_dadda_pg_rca24_and_12_12 ^ s_dadda_pg_rca24_and_11_13;
  assign s_dadda_pg_rca24_fa173_and0 = s_dadda_pg_rca24_and_12_12 & s_dadda_pg_rca24_and_11_13;
  assign s_dadda_pg_rca24_fa173_xor1 = s_dadda_pg_rca24_fa173_xor0 ^ s_dadda_pg_rca24_and_10_14;
  assign s_dadda_pg_rca24_fa173_and1 = s_dadda_pg_rca24_fa173_xor0 & s_dadda_pg_rca24_and_10_14;
  assign s_dadda_pg_rca24_fa173_or0 = s_dadda_pg_rca24_fa173_and0 | s_dadda_pg_rca24_fa173_and1;
  assign s_dadda_pg_rca24_and_9_15 = a[9] & b[15];
  assign s_dadda_pg_rca24_and_8_16 = a[8] & b[16];
  assign s_dadda_pg_rca24_and_7_17 = a[7] & b[17];
  assign s_dadda_pg_rca24_fa174_xor0 = s_dadda_pg_rca24_and_9_15 ^ s_dadda_pg_rca24_and_8_16;
  assign s_dadda_pg_rca24_fa174_and0 = s_dadda_pg_rca24_and_9_15 & s_dadda_pg_rca24_and_8_16;
  assign s_dadda_pg_rca24_fa174_xor1 = s_dadda_pg_rca24_fa174_xor0 ^ s_dadda_pg_rca24_and_7_17;
  assign s_dadda_pg_rca24_fa174_and1 = s_dadda_pg_rca24_fa174_xor0 & s_dadda_pg_rca24_and_7_17;
  assign s_dadda_pg_rca24_fa174_or0 = s_dadda_pg_rca24_fa174_and0 | s_dadda_pg_rca24_fa174_and1;
  assign s_dadda_pg_rca24_and_6_18 = a[6] & b[18];
  assign s_dadda_pg_rca24_and_5_19 = a[5] & b[19];
  assign s_dadda_pg_rca24_and_4_20 = a[4] & b[20];
  assign s_dadda_pg_rca24_fa175_xor0 = s_dadda_pg_rca24_and_6_18 ^ s_dadda_pg_rca24_and_5_19;
  assign s_dadda_pg_rca24_fa175_and0 = s_dadda_pg_rca24_and_6_18 & s_dadda_pg_rca24_and_5_19;
  assign s_dadda_pg_rca24_fa175_xor1 = s_dadda_pg_rca24_fa175_xor0 ^ s_dadda_pg_rca24_and_4_20;
  assign s_dadda_pg_rca24_fa175_and1 = s_dadda_pg_rca24_fa175_xor0 & s_dadda_pg_rca24_and_4_20;
  assign s_dadda_pg_rca24_fa175_or0 = s_dadda_pg_rca24_fa175_and0 | s_dadda_pg_rca24_fa175_and1;
  assign s_dadda_pg_rca24_and_3_21 = a[3] & b[21];
  assign s_dadda_pg_rca24_and_2_22 = a[2] & b[22];
  assign s_dadda_pg_rca24_nand_1_23 = ~(a[1] & b[23]);
  assign s_dadda_pg_rca24_fa176_xor0 = s_dadda_pg_rca24_and_3_21 ^ s_dadda_pg_rca24_and_2_22;
  assign s_dadda_pg_rca24_fa176_and0 = s_dadda_pg_rca24_and_3_21 & s_dadda_pg_rca24_and_2_22;
  assign s_dadda_pg_rca24_fa176_xor1 = s_dadda_pg_rca24_fa176_xor0 ^ s_dadda_pg_rca24_nand_1_23;
  assign s_dadda_pg_rca24_fa176_and1 = s_dadda_pg_rca24_fa176_xor0 & s_dadda_pg_rca24_nand_1_23;
  assign s_dadda_pg_rca24_fa176_or0 = s_dadda_pg_rca24_fa176_and0 | s_dadda_pg_rca24_fa176_and1;
  assign s_dadda_pg_rca24_fa177_xor0 = s_dadda_pg_rca24_fa10_xor1 ^ s_dadda_pg_rca24_fa11_xor1;
  assign s_dadda_pg_rca24_fa177_and0 = s_dadda_pg_rca24_fa10_xor1 & s_dadda_pg_rca24_fa11_xor1;
  assign s_dadda_pg_rca24_fa177_xor1 = s_dadda_pg_rca24_fa177_xor0 ^ s_dadda_pg_rca24_fa12_xor1;
  assign s_dadda_pg_rca24_fa177_and1 = s_dadda_pg_rca24_fa177_xor0 & s_dadda_pg_rca24_fa12_xor1;
  assign s_dadda_pg_rca24_fa177_or0 = s_dadda_pg_rca24_fa177_and0 | s_dadda_pg_rca24_fa177_and1;
  assign s_dadda_pg_rca24_fa178_xor0 = s_dadda_pg_rca24_fa13_xor1 ^ s_dadda_pg_rca24_fa14_xor1;
  assign s_dadda_pg_rca24_fa178_and0 = s_dadda_pg_rca24_fa13_xor1 & s_dadda_pg_rca24_fa14_xor1;
  assign s_dadda_pg_rca24_fa178_xor1 = s_dadda_pg_rca24_fa178_xor0 ^ s_dadda_pg_rca24_fa168_xor1;
  assign s_dadda_pg_rca24_fa178_and1 = s_dadda_pg_rca24_fa178_xor0 & s_dadda_pg_rca24_fa168_xor1;
  assign s_dadda_pg_rca24_fa178_or0 = s_dadda_pg_rca24_fa178_and0 | s_dadda_pg_rca24_fa178_and1;
  assign s_dadda_pg_rca24_fa179_xor0 = s_dadda_pg_rca24_fa169_xor1 ^ s_dadda_pg_rca24_fa170_xor1;
  assign s_dadda_pg_rca24_fa179_and0 = s_dadda_pg_rca24_fa169_xor1 & s_dadda_pg_rca24_fa170_xor1;
  assign s_dadda_pg_rca24_fa179_xor1 = s_dadda_pg_rca24_fa179_xor0 ^ s_dadda_pg_rca24_fa171_xor1;
  assign s_dadda_pg_rca24_fa179_and1 = s_dadda_pg_rca24_fa179_xor0 & s_dadda_pg_rca24_fa171_xor1;
  assign s_dadda_pg_rca24_fa179_or0 = s_dadda_pg_rca24_fa179_and0 | s_dadda_pg_rca24_fa179_and1;
  assign s_dadda_pg_rca24_fa180_xor0 = s_dadda_pg_rca24_fa172_xor1 ^ s_dadda_pg_rca24_fa173_xor1;
  assign s_dadda_pg_rca24_fa180_and0 = s_dadda_pg_rca24_fa172_xor1 & s_dadda_pg_rca24_fa173_xor1;
  assign s_dadda_pg_rca24_fa180_xor1 = s_dadda_pg_rca24_fa180_xor0 ^ s_dadda_pg_rca24_fa174_xor1;
  assign s_dadda_pg_rca24_fa180_and1 = s_dadda_pg_rca24_fa180_xor0 & s_dadda_pg_rca24_fa174_xor1;
  assign s_dadda_pg_rca24_fa180_or0 = s_dadda_pg_rca24_fa180_and0 | s_dadda_pg_rca24_fa180_and1;
  assign s_dadda_pg_rca24_fa181_xor0 = s_dadda_pg_rca24_fa180_or0 ^ s_dadda_pg_rca24_fa179_or0;
  assign s_dadda_pg_rca24_fa181_and0 = s_dadda_pg_rca24_fa180_or0 & s_dadda_pg_rca24_fa179_or0;
  assign s_dadda_pg_rca24_fa181_xor1 = s_dadda_pg_rca24_fa181_xor0 ^ s_dadda_pg_rca24_fa178_or0;
  assign s_dadda_pg_rca24_fa181_and1 = s_dadda_pg_rca24_fa181_xor0 & s_dadda_pg_rca24_fa178_or0;
  assign s_dadda_pg_rca24_fa181_or0 = s_dadda_pg_rca24_fa181_and0 | s_dadda_pg_rca24_fa181_and1;
  assign s_dadda_pg_rca24_fa182_xor0 = s_dadda_pg_rca24_fa177_or0 ^ s_dadda_pg_rca24_fa176_or0;
  assign s_dadda_pg_rca24_fa182_and0 = s_dadda_pg_rca24_fa177_or0 & s_dadda_pg_rca24_fa176_or0;
  assign s_dadda_pg_rca24_fa182_xor1 = s_dadda_pg_rca24_fa182_xor0 ^ s_dadda_pg_rca24_fa175_or0;
  assign s_dadda_pg_rca24_fa182_and1 = s_dadda_pg_rca24_fa182_xor0 & s_dadda_pg_rca24_fa175_or0;
  assign s_dadda_pg_rca24_fa182_or0 = s_dadda_pg_rca24_fa182_and0 | s_dadda_pg_rca24_fa182_and1;
  assign s_dadda_pg_rca24_fa183_xor0 = s_dadda_pg_rca24_fa174_or0 ^ s_dadda_pg_rca24_fa173_or0;
  assign s_dadda_pg_rca24_fa183_and0 = s_dadda_pg_rca24_fa174_or0 & s_dadda_pg_rca24_fa173_or0;
  assign s_dadda_pg_rca24_fa183_xor1 = s_dadda_pg_rca24_fa183_xor0 ^ s_dadda_pg_rca24_fa172_or0;
  assign s_dadda_pg_rca24_fa183_and1 = s_dadda_pg_rca24_fa183_xor0 & s_dadda_pg_rca24_fa172_or0;
  assign s_dadda_pg_rca24_fa183_or0 = s_dadda_pg_rca24_fa183_and0 | s_dadda_pg_rca24_fa183_and1;
  assign s_dadda_pg_rca24_fa184_xor0 = s_dadda_pg_rca24_fa171_or0 ^ s_dadda_pg_rca24_fa170_or0;
  assign s_dadda_pg_rca24_fa184_and0 = s_dadda_pg_rca24_fa171_or0 & s_dadda_pg_rca24_fa170_or0;
  assign s_dadda_pg_rca24_fa184_xor1 = s_dadda_pg_rca24_fa184_xor0 ^ s_dadda_pg_rca24_fa169_or0;
  assign s_dadda_pg_rca24_fa184_and1 = s_dadda_pg_rca24_fa184_xor0 & s_dadda_pg_rca24_fa169_or0;
  assign s_dadda_pg_rca24_fa184_or0 = s_dadda_pg_rca24_fa184_and0 | s_dadda_pg_rca24_fa184_and1;
  assign s_dadda_pg_rca24_and_16_9 = a[16] & b[9];
  assign s_dadda_pg_rca24_and_15_10 = a[15] & b[10];
  assign s_dadda_pg_rca24_fa185_xor0 = s_dadda_pg_rca24_fa168_or0 ^ s_dadda_pg_rca24_and_16_9;
  assign s_dadda_pg_rca24_fa185_and0 = s_dadda_pg_rca24_fa168_or0 & s_dadda_pg_rca24_and_16_9;
  assign s_dadda_pg_rca24_fa185_xor1 = s_dadda_pg_rca24_fa185_xor0 ^ s_dadda_pg_rca24_and_15_10;
  assign s_dadda_pg_rca24_fa185_and1 = s_dadda_pg_rca24_fa185_xor0 & s_dadda_pg_rca24_and_15_10;
  assign s_dadda_pg_rca24_fa185_or0 = s_dadda_pg_rca24_fa185_and0 | s_dadda_pg_rca24_fa185_and1;
  assign s_dadda_pg_rca24_and_14_11 = a[14] & b[11];
  assign s_dadda_pg_rca24_and_13_12 = a[13] & b[12];
  assign s_dadda_pg_rca24_and_12_13 = a[12] & b[13];
  assign s_dadda_pg_rca24_fa186_xor0 = s_dadda_pg_rca24_and_14_11 ^ s_dadda_pg_rca24_and_13_12;
  assign s_dadda_pg_rca24_fa186_and0 = s_dadda_pg_rca24_and_14_11 & s_dadda_pg_rca24_and_13_12;
  assign s_dadda_pg_rca24_fa186_xor1 = s_dadda_pg_rca24_fa186_xor0 ^ s_dadda_pg_rca24_and_12_13;
  assign s_dadda_pg_rca24_fa186_and1 = s_dadda_pg_rca24_fa186_xor0 & s_dadda_pg_rca24_and_12_13;
  assign s_dadda_pg_rca24_fa186_or0 = s_dadda_pg_rca24_fa186_and0 | s_dadda_pg_rca24_fa186_and1;
  assign s_dadda_pg_rca24_and_11_14 = a[11] & b[14];
  assign s_dadda_pg_rca24_and_10_15 = a[10] & b[15];
  assign s_dadda_pg_rca24_and_9_16 = a[9] & b[16];
  assign s_dadda_pg_rca24_fa187_xor0 = s_dadda_pg_rca24_and_11_14 ^ s_dadda_pg_rca24_and_10_15;
  assign s_dadda_pg_rca24_fa187_and0 = s_dadda_pg_rca24_and_11_14 & s_dadda_pg_rca24_and_10_15;
  assign s_dadda_pg_rca24_fa187_xor1 = s_dadda_pg_rca24_fa187_xor0 ^ s_dadda_pg_rca24_and_9_16;
  assign s_dadda_pg_rca24_fa187_and1 = s_dadda_pg_rca24_fa187_xor0 & s_dadda_pg_rca24_and_9_16;
  assign s_dadda_pg_rca24_fa187_or0 = s_dadda_pg_rca24_fa187_and0 | s_dadda_pg_rca24_fa187_and1;
  assign s_dadda_pg_rca24_and_8_17 = a[8] & b[17];
  assign s_dadda_pg_rca24_and_7_18 = a[7] & b[18];
  assign s_dadda_pg_rca24_and_6_19 = a[6] & b[19];
  assign s_dadda_pg_rca24_fa188_xor0 = s_dadda_pg_rca24_and_8_17 ^ s_dadda_pg_rca24_and_7_18;
  assign s_dadda_pg_rca24_fa188_and0 = s_dadda_pg_rca24_and_8_17 & s_dadda_pg_rca24_and_7_18;
  assign s_dadda_pg_rca24_fa188_xor1 = s_dadda_pg_rca24_fa188_xor0 ^ s_dadda_pg_rca24_and_6_19;
  assign s_dadda_pg_rca24_fa188_and1 = s_dadda_pg_rca24_fa188_xor0 & s_dadda_pg_rca24_and_6_19;
  assign s_dadda_pg_rca24_fa188_or0 = s_dadda_pg_rca24_fa188_and0 | s_dadda_pg_rca24_fa188_and1;
  assign s_dadda_pg_rca24_and_5_20 = a[5] & b[20];
  assign s_dadda_pg_rca24_and_4_21 = a[4] & b[21];
  assign s_dadda_pg_rca24_and_3_22 = a[3] & b[22];
  assign s_dadda_pg_rca24_fa189_xor0 = s_dadda_pg_rca24_and_5_20 ^ s_dadda_pg_rca24_and_4_21;
  assign s_dadda_pg_rca24_fa189_and0 = s_dadda_pg_rca24_and_5_20 & s_dadda_pg_rca24_and_4_21;
  assign s_dadda_pg_rca24_fa189_xor1 = s_dadda_pg_rca24_fa189_xor0 ^ s_dadda_pg_rca24_and_3_22;
  assign s_dadda_pg_rca24_fa189_and1 = s_dadda_pg_rca24_fa189_xor0 & s_dadda_pg_rca24_and_3_22;
  assign s_dadda_pg_rca24_fa189_or0 = s_dadda_pg_rca24_fa189_and0 | s_dadda_pg_rca24_fa189_and1;
  assign s_dadda_pg_rca24_nand_2_23 = ~(a[2] & b[23]);
  assign s_dadda_pg_rca24_fa190_xor0 = s_dadda_pg_rca24_nand_2_23 ^ s_dadda_pg_rca24_fa15_xor1;
  assign s_dadda_pg_rca24_fa190_and0 = s_dadda_pg_rca24_nand_2_23 & s_dadda_pg_rca24_fa15_xor1;
  assign s_dadda_pg_rca24_fa190_xor1 = s_dadda_pg_rca24_fa190_xor0 ^ s_dadda_pg_rca24_fa16_xor1;
  assign s_dadda_pg_rca24_fa190_and1 = s_dadda_pg_rca24_fa190_xor0 & s_dadda_pg_rca24_fa16_xor1;
  assign s_dadda_pg_rca24_fa190_or0 = s_dadda_pg_rca24_fa190_and0 | s_dadda_pg_rca24_fa190_and1;
  assign s_dadda_pg_rca24_fa191_xor0 = s_dadda_pg_rca24_fa17_xor1 ^ s_dadda_pg_rca24_fa18_xor1;
  assign s_dadda_pg_rca24_fa191_and0 = s_dadda_pg_rca24_fa17_xor1 & s_dadda_pg_rca24_fa18_xor1;
  assign s_dadda_pg_rca24_fa191_xor1 = s_dadda_pg_rca24_fa191_xor0 ^ s_dadda_pg_rca24_fa181_xor1;
  assign s_dadda_pg_rca24_fa191_and1 = s_dadda_pg_rca24_fa191_xor0 & s_dadda_pg_rca24_fa181_xor1;
  assign s_dadda_pg_rca24_fa191_or0 = s_dadda_pg_rca24_fa191_and0 | s_dadda_pg_rca24_fa191_and1;
  assign s_dadda_pg_rca24_fa192_xor0 = s_dadda_pg_rca24_fa182_xor1 ^ s_dadda_pg_rca24_fa183_xor1;
  assign s_dadda_pg_rca24_fa192_and0 = s_dadda_pg_rca24_fa182_xor1 & s_dadda_pg_rca24_fa183_xor1;
  assign s_dadda_pg_rca24_fa192_xor1 = s_dadda_pg_rca24_fa192_xor0 ^ s_dadda_pg_rca24_fa184_xor1;
  assign s_dadda_pg_rca24_fa192_and1 = s_dadda_pg_rca24_fa192_xor0 & s_dadda_pg_rca24_fa184_xor1;
  assign s_dadda_pg_rca24_fa192_or0 = s_dadda_pg_rca24_fa192_and0 | s_dadda_pg_rca24_fa192_and1;
  assign s_dadda_pg_rca24_fa193_xor0 = s_dadda_pg_rca24_fa185_xor1 ^ s_dadda_pg_rca24_fa186_xor1;
  assign s_dadda_pg_rca24_fa193_and0 = s_dadda_pg_rca24_fa185_xor1 & s_dadda_pg_rca24_fa186_xor1;
  assign s_dadda_pg_rca24_fa193_xor1 = s_dadda_pg_rca24_fa193_xor0 ^ s_dadda_pg_rca24_fa187_xor1;
  assign s_dadda_pg_rca24_fa193_and1 = s_dadda_pg_rca24_fa193_xor0 & s_dadda_pg_rca24_fa187_xor1;
  assign s_dadda_pg_rca24_fa193_or0 = s_dadda_pg_rca24_fa193_and0 | s_dadda_pg_rca24_fa193_and1;
  assign s_dadda_pg_rca24_fa194_xor0 = s_dadda_pg_rca24_fa193_or0 ^ s_dadda_pg_rca24_fa192_or0;
  assign s_dadda_pg_rca24_fa194_and0 = s_dadda_pg_rca24_fa193_or0 & s_dadda_pg_rca24_fa192_or0;
  assign s_dadda_pg_rca24_fa194_xor1 = s_dadda_pg_rca24_fa194_xor0 ^ s_dadda_pg_rca24_fa191_or0;
  assign s_dadda_pg_rca24_fa194_and1 = s_dadda_pg_rca24_fa194_xor0 & s_dadda_pg_rca24_fa191_or0;
  assign s_dadda_pg_rca24_fa194_or0 = s_dadda_pg_rca24_fa194_and0 | s_dadda_pg_rca24_fa194_and1;
  assign s_dadda_pg_rca24_fa195_xor0 = s_dadda_pg_rca24_fa190_or0 ^ s_dadda_pg_rca24_fa189_or0;
  assign s_dadda_pg_rca24_fa195_and0 = s_dadda_pg_rca24_fa190_or0 & s_dadda_pg_rca24_fa189_or0;
  assign s_dadda_pg_rca24_fa195_xor1 = s_dadda_pg_rca24_fa195_xor0 ^ s_dadda_pg_rca24_fa188_or0;
  assign s_dadda_pg_rca24_fa195_and1 = s_dadda_pg_rca24_fa195_xor0 & s_dadda_pg_rca24_fa188_or0;
  assign s_dadda_pg_rca24_fa195_or0 = s_dadda_pg_rca24_fa195_and0 | s_dadda_pg_rca24_fa195_and1;
  assign s_dadda_pg_rca24_fa196_xor0 = s_dadda_pg_rca24_fa187_or0 ^ s_dadda_pg_rca24_fa186_or0;
  assign s_dadda_pg_rca24_fa196_and0 = s_dadda_pg_rca24_fa187_or0 & s_dadda_pg_rca24_fa186_or0;
  assign s_dadda_pg_rca24_fa196_xor1 = s_dadda_pg_rca24_fa196_xor0 ^ s_dadda_pg_rca24_fa185_or0;
  assign s_dadda_pg_rca24_fa196_and1 = s_dadda_pg_rca24_fa196_xor0 & s_dadda_pg_rca24_fa185_or0;
  assign s_dadda_pg_rca24_fa196_or0 = s_dadda_pg_rca24_fa196_and0 | s_dadda_pg_rca24_fa196_and1;
  assign s_dadda_pg_rca24_fa197_xor0 = s_dadda_pg_rca24_fa184_or0 ^ s_dadda_pg_rca24_fa183_or0;
  assign s_dadda_pg_rca24_fa197_and0 = s_dadda_pg_rca24_fa184_or0 & s_dadda_pg_rca24_fa183_or0;
  assign s_dadda_pg_rca24_fa197_xor1 = s_dadda_pg_rca24_fa197_xor0 ^ s_dadda_pg_rca24_fa182_or0;
  assign s_dadda_pg_rca24_fa197_and1 = s_dadda_pg_rca24_fa197_xor0 & s_dadda_pg_rca24_fa182_or0;
  assign s_dadda_pg_rca24_fa197_or0 = s_dadda_pg_rca24_fa197_and0 | s_dadda_pg_rca24_fa197_and1;
  assign s_dadda_pg_rca24_and_18_8 = a[18] & b[8];
  assign s_dadda_pg_rca24_and_17_9 = a[17] & b[9];
  assign s_dadda_pg_rca24_fa198_xor0 = s_dadda_pg_rca24_fa181_or0 ^ s_dadda_pg_rca24_and_18_8;
  assign s_dadda_pg_rca24_fa198_and0 = s_dadda_pg_rca24_fa181_or0 & s_dadda_pg_rca24_and_18_8;
  assign s_dadda_pg_rca24_fa198_xor1 = s_dadda_pg_rca24_fa198_xor0 ^ s_dadda_pg_rca24_and_17_9;
  assign s_dadda_pg_rca24_fa198_and1 = s_dadda_pg_rca24_fa198_xor0 & s_dadda_pg_rca24_and_17_9;
  assign s_dadda_pg_rca24_fa198_or0 = s_dadda_pg_rca24_fa198_and0 | s_dadda_pg_rca24_fa198_and1;
  assign s_dadda_pg_rca24_and_16_10 = a[16] & b[10];
  assign s_dadda_pg_rca24_and_15_11 = a[15] & b[11];
  assign s_dadda_pg_rca24_and_14_12 = a[14] & b[12];
  assign s_dadda_pg_rca24_fa199_xor0 = s_dadda_pg_rca24_and_16_10 ^ s_dadda_pg_rca24_and_15_11;
  assign s_dadda_pg_rca24_fa199_and0 = s_dadda_pg_rca24_and_16_10 & s_dadda_pg_rca24_and_15_11;
  assign s_dadda_pg_rca24_fa199_xor1 = s_dadda_pg_rca24_fa199_xor0 ^ s_dadda_pg_rca24_and_14_12;
  assign s_dadda_pg_rca24_fa199_and1 = s_dadda_pg_rca24_fa199_xor0 & s_dadda_pg_rca24_and_14_12;
  assign s_dadda_pg_rca24_fa199_or0 = s_dadda_pg_rca24_fa199_and0 | s_dadda_pg_rca24_fa199_and1;
  assign s_dadda_pg_rca24_and_13_13 = a[13] & b[13];
  assign s_dadda_pg_rca24_and_12_14 = a[12] & b[14];
  assign s_dadda_pg_rca24_and_11_15 = a[11] & b[15];
  assign s_dadda_pg_rca24_fa200_xor0 = s_dadda_pg_rca24_and_13_13 ^ s_dadda_pg_rca24_and_12_14;
  assign s_dadda_pg_rca24_fa200_and0 = s_dadda_pg_rca24_and_13_13 & s_dadda_pg_rca24_and_12_14;
  assign s_dadda_pg_rca24_fa200_xor1 = s_dadda_pg_rca24_fa200_xor0 ^ s_dadda_pg_rca24_and_11_15;
  assign s_dadda_pg_rca24_fa200_and1 = s_dadda_pg_rca24_fa200_xor0 & s_dadda_pg_rca24_and_11_15;
  assign s_dadda_pg_rca24_fa200_or0 = s_dadda_pg_rca24_fa200_and0 | s_dadda_pg_rca24_fa200_and1;
  assign s_dadda_pg_rca24_and_10_16 = a[10] & b[16];
  assign s_dadda_pg_rca24_and_9_17 = a[9] & b[17];
  assign s_dadda_pg_rca24_and_8_18 = a[8] & b[18];
  assign s_dadda_pg_rca24_fa201_xor0 = s_dadda_pg_rca24_and_10_16 ^ s_dadda_pg_rca24_and_9_17;
  assign s_dadda_pg_rca24_fa201_and0 = s_dadda_pg_rca24_and_10_16 & s_dadda_pg_rca24_and_9_17;
  assign s_dadda_pg_rca24_fa201_xor1 = s_dadda_pg_rca24_fa201_xor0 ^ s_dadda_pg_rca24_and_8_18;
  assign s_dadda_pg_rca24_fa201_and1 = s_dadda_pg_rca24_fa201_xor0 & s_dadda_pg_rca24_and_8_18;
  assign s_dadda_pg_rca24_fa201_or0 = s_dadda_pg_rca24_fa201_and0 | s_dadda_pg_rca24_fa201_and1;
  assign s_dadda_pg_rca24_and_7_19 = a[7] & b[19];
  assign s_dadda_pg_rca24_and_6_20 = a[6] & b[20];
  assign s_dadda_pg_rca24_and_5_21 = a[5] & b[21];
  assign s_dadda_pg_rca24_fa202_xor0 = s_dadda_pg_rca24_and_7_19 ^ s_dadda_pg_rca24_and_6_20;
  assign s_dadda_pg_rca24_fa202_and0 = s_dadda_pg_rca24_and_7_19 & s_dadda_pg_rca24_and_6_20;
  assign s_dadda_pg_rca24_fa202_xor1 = s_dadda_pg_rca24_fa202_xor0 ^ s_dadda_pg_rca24_and_5_21;
  assign s_dadda_pg_rca24_fa202_and1 = s_dadda_pg_rca24_fa202_xor0 & s_dadda_pg_rca24_and_5_21;
  assign s_dadda_pg_rca24_fa202_or0 = s_dadda_pg_rca24_fa202_and0 | s_dadda_pg_rca24_fa202_and1;
  assign s_dadda_pg_rca24_and_4_22 = a[4] & b[22];
  assign s_dadda_pg_rca24_nand_3_23 = ~(a[3] & b[23]);
  assign s_dadda_pg_rca24_fa203_xor0 = s_dadda_pg_rca24_and_4_22 ^ s_dadda_pg_rca24_nand_3_23;
  assign s_dadda_pg_rca24_fa203_and0 = s_dadda_pg_rca24_and_4_22 & s_dadda_pg_rca24_nand_3_23;
  assign s_dadda_pg_rca24_fa203_xor1 = s_dadda_pg_rca24_fa203_xor0 ^ s_dadda_pg_rca24_fa19_xor1;
  assign s_dadda_pg_rca24_fa203_and1 = s_dadda_pg_rca24_fa203_xor0 & s_dadda_pg_rca24_fa19_xor1;
  assign s_dadda_pg_rca24_fa203_or0 = s_dadda_pg_rca24_fa203_and0 | s_dadda_pg_rca24_fa203_and1;
  assign s_dadda_pg_rca24_fa204_xor0 = s_dadda_pg_rca24_fa20_xor1 ^ s_dadda_pg_rca24_fa21_xor1;
  assign s_dadda_pg_rca24_fa204_and0 = s_dadda_pg_rca24_fa20_xor1 & s_dadda_pg_rca24_fa21_xor1;
  assign s_dadda_pg_rca24_fa204_xor1 = s_dadda_pg_rca24_fa204_xor0 ^ s_dadda_pg_rca24_fa194_xor1;
  assign s_dadda_pg_rca24_fa204_and1 = s_dadda_pg_rca24_fa204_xor0 & s_dadda_pg_rca24_fa194_xor1;
  assign s_dadda_pg_rca24_fa204_or0 = s_dadda_pg_rca24_fa204_and0 | s_dadda_pg_rca24_fa204_and1;
  assign s_dadda_pg_rca24_fa205_xor0 = s_dadda_pg_rca24_fa195_xor1 ^ s_dadda_pg_rca24_fa196_xor1;
  assign s_dadda_pg_rca24_fa205_and0 = s_dadda_pg_rca24_fa195_xor1 & s_dadda_pg_rca24_fa196_xor1;
  assign s_dadda_pg_rca24_fa205_xor1 = s_dadda_pg_rca24_fa205_xor0 ^ s_dadda_pg_rca24_fa197_xor1;
  assign s_dadda_pg_rca24_fa205_and1 = s_dadda_pg_rca24_fa205_xor0 & s_dadda_pg_rca24_fa197_xor1;
  assign s_dadda_pg_rca24_fa205_or0 = s_dadda_pg_rca24_fa205_and0 | s_dadda_pg_rca24_fa205_and1;
  assign s_dadda_pg_rca24_fa206_xor0 = s_dadda_pg_rca24_fa198_xor1 ^ s_dadda_pg_rca24_fa199_xor1;
  assign s_dadda_pg_rca24_fa206_and0 = s_dadda_pg_rca24_fa198_xor1 & s_dadda_pg_rca24_fa199_xor1;
  assign s_dadda_pg_rca24_fa206_xor1 = s_dadda_pg_rca24_fa206_xor0 ^ s_dadda_pg_rca24_fa200_xor1;
  assign s_dadda_pg_rca24_fa206_and1 = s_dadda_pg_rca24_fa206_xor0 & s_dadda_pg_rca24_fa200_xor1;
  assign s_dadda_pg_rca24_fa206_or0 = s_dadda_pg_rca24_fa206_and0 | s_dadda_pg_rca24_fa206_and1;
  assign s_dadda_pg_rca24_fa207_xor0 = s_dadda_pg_rca24_fa206_or0 ^ s_dadda_pg_rca24_fa205_or0;
  assign s_dadda_pg_rca24_fa207_and0 = s_dadda_pg_rca24_fa206_or0 & s_dadda_pg_rca24_fa205_or0;
  assign s_dadda_pg_rca24_fa207_xor1 = s_dadda_pg_rca24_fa207_xor0 ^ s_dadda_pg_rca24_fa204_or0;
  assign s_dadda_pg_rca24_fa207_and1 = s_dadda_pg_rca24_fa207_xor0 & s_dadda_pg_rca24_fa204_or0;
  assign s_dadda_pg_rca24_fa207_or0 = s_dadda_pg_rca24_fa207_and0 | s_dadda_pg_rca24_fa207_and1;
  assign s_dadda_pg_rca24_fa208_xor0 = s_dadda_pg_rca24_fa203_or0 ^ s_dadda_pg_rca24_fa202_or0;
  assign s_dadda_pg_rca24_fa208_and0 = s_dadda_pg_rca24_fa203_or0 & s_dadda_pg_rca24_fa202_or0;
  assign s_dadda_pg_rca24_fa208_xor1 = s_dadda_pg_rca24_fa208_xor0 ^ s_dadda_pg_rca24_fa201_or0;
  assign s_dadda_pg_rca24_fa208_and1 = s_dadda_pg_rca24_fa208_xor0 & s_dadda_pg_rca24_fa201_or0;
  assign s_dadda_pg_rca24_fa208_or0 = s_dadda_pg_rca24_fa208_and0 | s_dadda_pg_rca24_fa208_and1;
  assign s_dadda_pg_rca24_fa209_xor0 = s_dadda_pg_rca24_fa200_or0 ^ s_dadda_pg_rca24_fa199_or0;
  assign s_dadda_pg_rca24_fa209_and0 = s_dadda_pg_rca24_fa200_or0 & s_dadda_pg_rca24_fa199_or0;
  assign s_dadda_pg_rca24_fa209_xor1 = s_dadda_pg_rca24_fa209_xor0 ^ s_dadda_pg_rca24_fa198_or0;
  assign s_dadda_pg_rca24_fa209_and1 = s_dadda_pg_rca24_fa209_xor0 & s_dadda_pg_rca24_fa198_or0;
  assign s_dadda_pg_rca24_fa209_or0 = s_dadda_pg_rca24_fa209_and0 | s_dadda_pg_rca24_fa209_and1;
  assign s_dadda_pg_rca24_fa210_xor0 = s_dadda_pg_rca24_fa197_or0 ^ s_dadda_pg_rca24_fa196_or0;
  assign s_dadda_pg_rca24_fa210_and0 = s_dadda_pg_rca24_fa197_or0 & s_dadda_pg_rca24_fa196_or0;
  assign s_dadda_pg_rca24_fa210_xor1 = s_dadda_pg_rca24_fa210_xor0 ^ s_dadda_pg_rca24_fa195_or0;
  assign s_dadda_pg_rca24_fa210_and1 = s_dadda_pg_rca24_fa210_xor0 & s_dadda_pg_rca24_fa195_or0;
  assign s_dadda_pg_rca24_fa210_or0 = s_dadda_pg_rca24_fa210_and0 | s_dadda_pg_rca24_fa210_and1;
  assign s_dadda_pg_rca24_and_20_7 = a[20] & b[7];
  assign s_dadda_pg_rca24_and_19_8 = a[19] & b[8];
  assign s_dadda_pg_rca24_fa211_xor0 = s_dadda_pg_rca24_fa194_or0 ^ s_dadda_pg_rca24_and_20_7;
  assign s_dadda_pg_rca24_fa211_and0 = s_dadda_pg_rca24_fa194_or0 & s_dadda_pg_rca24_and_20_7;
  assign s_dadda_pg_rca24_fa211_xor1 = s_dadda_pg_rca24_fa211_xor0 ^ s_dadda_pg_rca24_and_19_8;
  assign s_dadda_pg_rca24_fa211_and1 = s_dadda_pg_rca24_fa211_xor0 & s_dadda_pg_rca24_and_19_8;
  assign s_dadda_pg_rca24_fa211_or0 = s_dadda_pg_rca24_fa211_and0 | s_dadda_pg_rca24_fa211_and1;
  assign s_dadda_pg_rca24_and_18_9 = a[18] & b[9];
  assign s_dadda_pg_rca24_and_17_10 = a[17] & b[10];
  assign s_dadda_pg_rca24_and_16_11 = a[16] & b[11];
  assign s_dadda_pg_rca24_fa212_xor0 = s_dadda_pg_rca24_and_18_9 ^ s_dadda_pg_rca24_and_17_10;
  assign s_dadda_pg_rca24_fa212_and0 = s_dadda_pg_rca24_and_18_9 & s_dadda_pg_rca24_and_17_10;
  assign s_dadda_pg_rca24_fa212_xor1 = s_dadda_pg_rca24_fa212_xor0 ^ s_dadda_pg_rca24_and_16_11;
  assign s_dadda_pg_rca24_fa212_and1 = s_dadda_pg_rca24_fa212_xor0 & s_dadda_pg_rca24_and_16_11;
  assign s_dadda_pg_rca24_fa212_or0 = s_dadda_pg_rca24_fa212_and0 | s_dadda_pg_rca24_fa212_and1;
  assign s_dadda_pg_rca24_and_15_12 = a[15] & b[12];
  assign s_dadda_pg_rca24_and_14_13 = a[14] & b[13];
  assign s_dadda_pg_rca24_and_13_14 = a[13] & b[14];
  assign s_dadda_pg_rca24_fa213_xor0 = s_dadda_pg_rca24_and_15_12 ^ s_dadda_pg_rca24_and_14_13;
  assign s_dadda_pg_rca24_fa213_and0 = s_dadda_pg_rca24_and_15_12 & s_dadda_pg_rca24_and_14_13;
  assign s_dadda_pg_rca24_fa213_xor1 = s_dadda_pg_rca24_fa213_xor0 ^ s_dadda_pg_rca24_and_13_14;
  assign s_dadda_pg_rca24_fa213_and1 = s_dadda_pg_rca24_fa213_xor0 & s_dadda_pg_rca24_and_13_14;
  assign s_dadda_pg_rca24_fa213_or0 = s_dadda_pg_rca24_fa213_and0 | s_dadda_pg_rca24_fa213_and1;
  assign s_dadda_pg_rca24_and_12_15 = a[12] & b[15];
  assign s_dadda_pg_rca24_and_11_16 = a[11] & b[16];
  assign s_dadda_pg_rca24_and_10_17 = a[10] & b[17];
  assign s_dadda_pg_rca24_fa214_xor0 = s_dadda_pg_rca24_and_12_15 ^ s_dadda_pg_rca24_and_11_16;
  assign s_dadda_pg_rca24_fa214_and0 = s_dadda_pg_rca24_and_12_15 & s_dadda_pg_rca24_and_11_16;
  assign s_dadda_pg_rca24_fa214_xor1 = s_dadda_pg_rca24_fa214_xor0 ^ s_dadda_pg_rca24_and_10_17;
  assign s_dadda_pg_rca24_fa214_and1 = s_dadda_pg_rca24_fa214_xor0 & s_dadda_pg_rca24_and_10_17;
  assign s_dadda_pg_rca24_fa214_or0 = s_dadda_pg_rca24_fa214_and0 | s_dadda_pg_rca24_fa214_and1;
  assign s_dadda_pg_rca24_and_9_18 = a[9] & b[18];
  assign s_dadda_pg_rca24_and_8_19 = a[8] & b[19];
  assign s_dadda_pg_rca24_and_7_20 = a[7] & b[20];
  assign s_dadda_pg_rca24_fa215_xor0 = s_dadda_pg_rca24_and_9_18 ^ s_dadda_pg_rca24_and_8_19;
  assign s_dadda_pg_rca24_fa215_and0 = s_dadda_pg_rca24_and_9_18 & s_dadda_pg_rca24_and_8_19;
  assign s_dadda_pg_rca24_fa215_xor1 = s_dadda_pg_rca24_fa215_xor0 ^ s_dadda_pg_rca24_and_7_20;
  assign s_dadda_pg_rca24_fa215_and1 = s_dadda_pg_rca24_fa215_xor0 & s_dadda_pg_rca24_and_7_20;
  assign s_dadda_pg_rca24_fa215_or0 = s_dadda_pg_rca24_fa215_and0 | s_dadda_pg_rca24_fa215_and1;
  assign s_dadda_pg_rca24_and_6_21 = a[6] & b[21];
  assign s_dadda_pg_rca24_and_5_22 = a[5] & b[22];
  assign s_dadda_pg_rca24_nand_4_23 = ~(a[4] & b[23]);
  assign s_dadda_pg_rca24_fa216_xor0 = s_dadda_pg_rca24_and_6_21 ^ s_dadda_pg_rca24_and_5_22;
  assign s_dadda_pg_rca24_fa216_and0 = s_dadda_pg_rca24_and_6_21 & s_dadda_pg_rca24_and_5_22;
  assign s_dadda_pg_rca24_fa216_xor1 = s_dadda_pg_rca24_fa216_xor0 ^ s_dadda_pg_rca24_nand_4_23;
  assign s_dadda_pg_rca24_fa216_and1 = s_dadda_pg_rca24_fa216_xor0 & s_dadda_pg_rca24_nand_4_23;
  assign s_dadda_pg_rca24_fa216_or0 = s_dadda_pg_rca24_fa216_and0 | s_dadda_pg_rca24_fa216_and1;
  assign s_dadda_pg_rca24_fa217_xor0 = s_dadda_pg_rca24_fa22_xor1 ^ s_dadda_pg_rca24_fa23_xor1;
  assign s_dadda_pg_rca24_fa217_and0 = s_dadda_pg_rca24_fa22_xor1 & s_dadda_pg_rca24_fa23_xor1;
  assign s_dadda_pg_rca24_fa217_xor1 = s_dadda_pg_rca24_fa217_xor0 ^ s_dadda_pg_rca24_fa207_xor1;
  assign s_dadda_pg_rca24_fa217_and1 = s_dadda_pg_rca24_fa217_xor0 & s_dadda_pg_rca24_fa207_xor1;
  assign s_dadda_pg_rca24_fa217_or0 = s_dadda_pg_rca24_fa217_and0 | s_dadda_pg_rca24_fa217_and1;
  assign s_dadda_pg_rca24_fa218_xor0 = s_dadda_pg_rca24_fa208_xor1 ^ s_dadda_pg_rca24_fa209_xor1;
  assign s_dadda_pg_rca24_fa218_and0 = s_dadda_pg_rca24_fa208_xor1 & s_dadda_pg_rca24_fa209_xor1;
  assign s_dadda_pg_rca24_fa218_xor1 = s_dadda_pg_rca24_fa218_xor0 ^ s_dadda_pg_rca24_fa210_xor1;
  assign s_dadda_pg_rca24_fa218_and1 = s_dadda_pg_rca24_fa218_xor0 & s_dadda_pg_rca24_fa210_xor1;
  assign s_dadda_pg_rca24_fa218_or0 = s_dadda_pg_rca24_fa218_and0 | s_dadda_pg_rca24_fa218_and1;
  assign s_dadda_pg_rca24_fa219_xor0 = s_dadda_pg_rca24_fa211_xor1 ^ s_dadda_pg_rca24_fa212_xor1;
  assign s_dadda_pg_rca24_fa219_and0 = s_dadda_pg_rca24_fa211_xor1 & s_dadda_pg_rca24_fa212_xor1;
  assign s_dadda_pg_rca24_fa219_xor1 = s_dadda_pg_rca24_fa219_xor0 ^ s_dadda_pg_rca24_fa213_xor1;
  assign s_dadda_pg_rca24_fa219_and1 = s_dadda_pg_rca24_fa219_xor0 & s_dadda_pg_rca24_fa213_xor1;
  assign s_dadda_pg_rca24_fa219_or0 = s_dadda_pg_rca24_fa219_and0 | s_dadda_pg_rca24_fa219_and1;
  assign s_dadda_pg_rca24_fa220_xor0 = s_dadda_pg_rca24_fa219_or0 ^ s_dadda_pg_rca24_fa218_or0;
  assign s_dadda_pg_rca24_fa220_and0 = s_dadda_pg_rca24_fa219_or0 & s_dadda_pg_rca24_fa218_or0;
  assign s_dadda_pg_rca24_fa220_xor1 = s_dadda_pg_rca24_fa220_xor0 ^ s_dadda_pg_rca24_fa217_or0;
  assign s_dadda_pg_rca24_fa220_and1 = s_dadda_pg_rca24_fa220_xor0 & s_dadda_pg_rca24_fa217_or0;
  assign s_dadda_pg_rca24_fa220_or0 = s_dadda_pg_rca24_fa220_and0 | s_dadda_pg_rca24_fa220_and1;
  assign s_dadda_pg_rca24_fa221_xor0 = s_dadda_pg_rca24_fa216_or0 ^ s_dadda_pg_rca24_fa215_or0;
  assign s_dadda_pg_rca24_fa221_and0 = s_dadda_pg_rca24_fa216_or0 & s_dadda_pg_rca24_fa215_or0;
  assign s_dadda_pg_rca24_fa221_xor1 = s_dadda_pg_rca24_fa221_xor0 ^ s_dadda_pg_rca24_fa214_or0;
  assign s_dadda_pg_rca24_fa221_and1 = s_dadda_pg_rca24_fa221_xor0 & s_dadda_pg_rca24_fa214_or0;
  assign s_dadda_pg_rca24_fa221_or0 = s_dadda_pg_rca24_fa221_and0 | s_dadda_pg_rca24_fa221_and1;
  assign s_dadda_pg_rca24_fa222_xor0 = s_dadda_pg_rca24_fa213_or0 ^ s_dadda_pg_rca24_fa212_or0;
  assign s_dadda_pg_rca24_fa222_and0 = s_dadda_pg_rca24_fa213_or0 & s_dadda_pg_rca24_fa212_or0;
  assign s_dadda_pg_rca24_fa222_xor1 = s_dadda_pg_rca24_fa222_xor0 ^ s_dadda_pg_rca24_fa211_or0;
  assign s_dadda_pg_rca24_fa222_and1 = s_dadda_pg_rca24_fa222_xor0 & s_dadda_pg_rca24_fa211_or0;
  assign s_dadda_pg_rca24_fa222_or0 = s_dadda_pg_rca24_fa222_and0 | s_dadda_pg_rca24_fa222_and1;
  assign s_dadda_pg_rca24_fa223_xor0 = s_dadda_pg_rca24_fa210_or0 ^ s_dadda_pg_rca24_fa209_or0;
  assign s_dadda_pg_rca24_fa223_and0 = s_dadda_pg_rca24_fa210_or0 & s_dadda_pg_rca24_fa209_or0;
  assign s_dadda_pg_rca24_fa223_xor1 = s_dadda_pg_rca24_fa223_xor0 ^ s_dadda_pg_rca24_fa208_or0;
  assign s_dadda_pg_rca24_fa223_and1 = s_dadda_pg_rca24_fa223_xor0 & s_dadda_pg_rca24_fa208_or0;
  assign s_dadda_pg_rca24_fa223_or0 = s_dadda_pg_rca24_fa223_and0 | s_dadda_pg_rca24_fa223_and1;
  assign s_dadda_pg_rca24_and_22_6 = a[22] & b[6];
  assign s_dadda_pg_rca24_and_21_7 = a[21] & b[7];
  assign s_dadda_pg_rca24_fa224_xor0 = s_dadda_pg_rca24_fa207_or0 ^ s_dadda_pg_rca24_and_22_6;
  assign s_dadda_pg_rca24_fa224_and0 = s_dadda_pg_rca24_fa207_or0 & s_dadda_pg_rca24_and_22_6;
  assign s_dadda_pg_rca24_fa224_xor1 = s_dadda_pg_rca24_fa224_xor0 ^ s_dadda_pg_rca24_and_21_7;
  assign s_dadda_pg_rca24_fa224_and1 = s_dadda_pg_rca24_fa224_xor0 & s_dadda_pg_rca24_and_21_7;
  assign s_dadda_pg_rca24_fa224_or0 = s_dadda_pg_rca24_fa224_and0 | s_dadda_pg_rca24_fa224_and1;
  assign s_dadda_pg_rca24_and_20_8 = a[20] & b[8];
  assign s_dadda_pg_rca24_and_19_9 = a[19] & b[9];
  assign s_dadda_pg_rca24_and_18_10 = a[18] & b[10];
  assign s_dadda_pg_rca24_fa225_xor0 = s_dadda_pg_rca24_and_20_8 ^ s_dadda_pg_rca24_and_19_9;
  assign s_dadda_pg_rca24_fa225_and0 = s_dadda_pg_rca24_and_20_8 & s_dadda_pg_rca24_and_19_9;
  assign s_dadda_pg_rca24_fa225_xor1 = s_dadda_pg_rca24_fa225_xor0 ^ s_dadda_pg_rca24_and_18_10;
  assign s_dadda_pg_rca24_fa225_and1 = s_dadda_pg_rca24_fa225_xor0 & s_dadda_pg_rca24_and_18_10;
  assign s_dadda_pg_rca24_fa225_or0 = s_dadda_pg_rca24_fa225_and0 | s_dadda_pg_rca24_fa225_and1;
  assign s_dadda_pg_rca24_and_17_11 = a[17] & b[11];
  assign s_dadda_pg_rca24_and_16_12 = a[16] & b[12];
  assign s_dadda_pg_rca24_and_15_13 = a[15] & b[13];
  assign s_dadda_pg_rca24_fa226_xor0 = s_dadda_pg_rca24_and_17_11 ^ s_dadda_pg_rca24_and_16_12;
  assign s_dadda_pg_rca24_fa226_and0 = s_dadda_pg_rca24_and_17_11 & s_dadda_pg_rca24_and_16_12;
  assign s_dadda_pg_rca24_fa226_xor1 = s_dadda_pg_rca24_fa226_xor0 ^ s_dadda_pg_rca24_and_15_13;
  assign s_dadda_pg_rca24_fa226_and1 = s_dadda_pg_rca24_fa226_xor0 & s_dadda_pg_rca24_and_15_13;
  assign s_dadda_pg_rca24_fa226_or0 = s_dadda_pg_rca24_fa226_and0 | s_dadda_pg_rca24_fa226_and1;
  assign s_dadda_pg_rca24_and_14_14 = a[14] & b[14];
  assign s_dadda_pg_rca24_and_13_15 = a[13] & b[15];
  assign s_dadda_pg_rca24_and_12_16 = a[12] & b[16];
  assign s_dadda_pg_rca24_fa227_xor0 = s_dadda_pg_rca24_and_14_14 ^ s_dadda_pg_rca24_and_13_15;
  assign s_dadda_pg_rca24_fa227_and0 = s_dadda_pg_rca24_and_14_14 & s_dadda_pg_rca24_and_13_15;
  assign s_dadda_pg_rca24_fa227_xor1 = s_dadda_pg_rca24_fa227_xor0 ^ s_dadda_pg_rca24_and_12_16;
  assign s_dadda_pg_rca24_fa227_and1 = s_dadda_pg_rca24_fa227_xor0 & s_dadda_pg_rca24_and_12_16;
  assign s_dadda_pg_rca24_fa227_or0 = s_dadda_pg_rca24_fa227_and0 | s_dadda_pg_rca24_fa227_and1;
  assign s_dadda_pg_rca24_and_11_17 = a[11] & b[17];
  assign s_dadda_pg_rca24_and_10_18 = a[10] & b[18];
  assign s_dadda_pg_rca24_and_9_19 = a[9] & b[19];
  assign s_dadda_pg_rca24_fa228_xor0 = s_dadda_pg_rca24_and_11_17 ^ s_dadda_pg_rca24_and_10_18;
  assign s_dadda_pg_rca24_fa228_and0 = s_dadda_pg_rca24_and_11_17 & s_dadda_pg_rca24_and_10_18;
  assign s_dadda_pg_rca24_fa228_xor1 = s_dadda_pg_rca24_fa228_xor0 ^ s_dadda_pg_rca24_and_9_19;
  assign s_dadda_pg_rca24_fa228_and1 = s_dadda_pg_rca24_fa228_xor0 & s_dadda_pg_rca24_and_9_19;
  assign s_dadda_pg_rca24_fa228_or0 = s_dadda_pg_rca24_fa228_and0 | s_dadda_pg_rca24_fa228_and1;
  assign s_dadda_pg_rca24_and_8_20 = a[8] & b[20];
  assign s_dadda_pg_rca24_and_7_21 = a[7] & b[21];
  assign s_dadda_pg_rca24_and_6_22 = a[6] & b[22];
  assign s_dadda_pg_rca24_fa229_xor0 = s_dadda_pg_rca24_and_8_20 ^ s_dadda_pg_rca24_and_7_21;
  assign s_dadda_pg_rca24_fa229_and0 = s_dadda_pg_rca24_and_8_20 & s_dadda_pg_rca24_and_7_21;
  assign s_dadda_pg_rca24_fa229_xor1 = s_dadda_pg_rca24_fa229_xor0 ^ s_dadda_pg_rca24_and_6_22;
  assign s_dadda_pg_rca24_fa229_and1 = s_dadda_pg_rca24_fa229_xor0 & s_dadda_pg_rca24_and_6_22;
  assign s_dadda_pg_rca24_fa229_or0 = s_dadda_pg_rca24_fa229_and0 | s_dadda_pg_rca24_fa229_and1;
  assign s_dadda_pg_rca24_nand_5_23 = ~(a[5] & b[23]);
  assign s_dadda_pg_rca24_fa230_xor0 = s_dadda_pg_rca24_nand_5_23 ^ s_dadda_pg_rca24_fa24_xor1;
  assign s_dadda_pg_rca24_fa230_and0 = s_dadda_pg_rca24_nand_5_23 & s_dadda_pg_rca24_fa24_xor1;
  assign s_dadda_pg_rca24_fa230_xor1 = s_dadda_pg_rca24_fa230_xor0 ^ s_dadda_pg_rca24_fa220_xor1;
  assign s_dadda_pg_rca24_fa230_and1 = s_dadda_pg_rca24_fa230_xor0 & s_dadda_pg_rca24_fa220_xor1;
  assign s_dadda_pg_rca24_fa230_or0 = s_dadda_pg_rca24_fa230_and0 | s_dadda_pg_rca24_fa230_and1;
  assign s_dadda_pg_rca24_fa231_xor0 = s_dadda_pg_rca24_fa221_xor1 ^ s_dadda_pg_rca24_fa222_xor1;
  assign s_dadda_pg_rca24_fa231_and0 = s_dadda_pg_rca24_fa221_xor1 & s_dadda_pg_rca24_fa222_xor1;
  assign s_dadda_pg_rca24_fa231_xor1 = s_dadda_pg_rca24_fa231_xor0 ^ s_dadda_pg_rca24_fa223_xor1;
  assign s_dadda_pg_rca24_fa231_and1 = s_dadda_pg_rca24_fa231_xor0 & s_dadda_pg_rca24_fa223_xor1;
  assign s_dadda_pg_rca24_fa231_or0 = s_dadda_pg_rca24_fa231_and0 | s_dadda_pg_rca24_fa231_and1;
  assign s_dadda_pg_rca24_fa232_xor0 = s_dadda_pg_rca24_fa224_xor1 ^ s_dadda_pg_rca24_fa225_xor1;
  assign s_dadda_pg_rca24_fa232_and0 = s_dadda_pg_rca24_fa224_xor1 & s_dadda_pg_rca24_fa225_xor1;
  assign s_dadda_pg_rca24_fa232_xor1 = s_dadda_pg_rca24_fa232_xor0 ^ s_dadda_pg_rca24_fa226_xor1;
  assign s_dadda_pg_rca24_fa232_and1 = s_dadda_pg_rca24_fa232_xor0 & s_dadda_pg_rca24_fa226_xor1;
  assign s_dadda_pg_rca24_fa232_or0 = s_dadda_pg_rca24_fa232_and0 | s_dadda_pg_rca24_fa232_and1;
  assign s_dadda_pg_rca24_fa233_xor0 = s_dadda_pg_rca24_fa232_or0 ^ s_dadda_pg_rca24_fa231_or0;
  assign s_dadda_pg_rca24_fa233_and0 = s_dadda_pg_rca24_fa232_or0 & s_dadda_pg_rca24_fa231_or0;
  assign s_dadda_pg_rca24_fa233_xor1 = s_dadda_pg_rca24_fa233_xor0 ^ s_dadda_pg_rca24_fa230_or0;
  assign s_dadda_pg_rca24_fa233_and1 = s_dadda_pg_rca24_fa233_xor0 & s_dadda_pg_rca24_fa230_or0;
  assign s_dadda_pg_rca24_fa233_or0 = s_dadda_pg_rca24_fa233_and0 | s_dadda_pg_rca24_fa233_and1;
  assign s_dadda_pg_rca24_fa234_xor0 = s_dadda_pg_rca24_fa229_or0 ^ s_dadda_pg_rca24_fa228_or0;
  assign s_dadda_pg_rca24_fa234_and0 = s_dadda_pg_rca24_fa229_or0 & s_dadda_pg_rca24_fa228_or0;
  assign s_dadda_pg_rca24_fa234_xor1 = s_dadda_pg_rca24_fa234_xor0 ^ s_dadda_pg_rca24_fa227_or0;
  assign s_dadda_pg_rca24_fa234_and1 = s_dadda_pg_rca24_fa234_xor0 & s_dadda_pg_rca24_fa227_or0;
  assign s_dadda_pg_rca24_fa234_or0 = s_dadda_pg_rca24_fa234_and0 | s_dadda_pg_rca24_fa234_and1;
  assign s_dadda_pg_rca24_fa235_xor0 = s_dadda_pg_rca24_fa226_or0 ^ s_dadda_pg_rca24_fa225_or0;
  assign s_dadda_pg_rca24_fa235_and0 = s_dadda_pg_rca24_fa226_or0 & s_dadda_pg_rca24_fa225_or0;
  assign s_dadda_pg_rca24_fa235_xor1 = s_dadda_pg_rca24_fa235_xor0 ^ s_dadda_pg_rca24_fa224_or0;
  assign s_dadda_pg_rca24_fa235_and1 = s_dadda_pg_rca24_fa235_xor0 & s_dadda_pg_rca24_fa224_or0;
  assign s_dadda_pg_rca24_fa235_or0 = s_dadda_pg_rca24_fa235_and0 | s_dadda_pg_rca24_fa235_and1;
  assign s_dadda_pg_rca24_fa236_xor0 = s_dadda_pg_rca24_fa223_or0 ^ s_dadda_pg_rca24_fa222_or0;
  assign s_dadda_pg_rca24_fa236_and0 = s_dadda_pg_rca24_fa223_or0 & s_dadda_pg_rca24_fa222_or0;
  assign s_dadda_pg_rca24_fa236_xor1 = s_dadda_pg_rca24_fa236_xor0 ^ s_dadda_pg_rca24_fa221_or0;
  assign s_dadda_pg_rca24_fa236_and1 = s_dadda_pg_rca24_fa236_xor0 & s_dadda_pg_rca24_fa221_or0;
  assign s_dadda_pg_rca24_fa236_or0 = s_dadda_pg_rca24_fa236_and0 | s_dadda_pg_rca24_fa236_and1;
  assign s_dadda_pg_rca24_nand_23_6 = ~(a[23] & b[6]);
  assign s_dadda_pg_rca24_fa237_xor0 = s_dadda_pg_rca24_fa220_or0 ^ s_dadda_pg_rca24_fa24_or0;
  assign s_dadda_pg_rca24_fa237_and0 = s_dadda_pg_rca24_fa220_or0 & s_dadda_pg_rca24_fa24_or0;
  assign s_dadda_pg_rca24_fa237_xor1 = s_dadda_pg_rca24_fa237_xor0 ^ s_dadda_pg_rca24_nand_23_6;
  assign s_dadda_pg_rca24_fa237_and1 = s_dadda_pg_rca24_fa237_xor0 & s_dadda_pg_rca24_nand_23_6;
  assign s_dadda_pg_rca24_fa237_or0 = s_dadda_pg_rca24_fa237_and0 | s_dadda_pg_rca24_fa237_and1;
  assign s_dadda_pg_rca24_and_22_7 = a[22] & b[7];
  assign s_dadda_pg_rca24_and_21_8 = a[21] & b[8];
  assign s_dadda_pg_rca24_and_20_9 = a[20] & b[9];
  assign s_dadda_pg_rca24_fa238_xor0 = s_dadda_pg_rca24_and_22_7 ^ s_dadda_pg_rca24_and_21_8;
  assign s_dadda_pg_rca24_fa238_and0 = s_dadda_pg_rca24_and_22_7 & s_dadda_pg_rca24_and_21_8;
  assign s_dadda_pg_rca24_fa238_xor1 = s_dadda_pg_rca24_fa238_xor0 ^ s_dadda_pg_rca24_and_20_9;
  assign s_dadda_pg_rca24_fa238_and1 = s_dadda_pg_rca24_fa238_xor0 & s_dadda_pg_rca24_and_20_9;
  assign s_dadda_pg_rca24_fa238_or0 = s_dadda_pg_rca24_fa238_and0 | s_dadda_pg_rca24_fa238_and1;
  assign s_dadda_pg_rca24_and_19_10 = a[19] & b[10];
  assign s_dadda_pg_rca24_and_18_11 = a[18] & b[11];
  assign s_dadda_pg_rca24_and_17_12 = a[17] & b[12];
  assign s_dadda_pg_rca24_fa239_xor0 = s_dadda_pg_rca24_and_19_10 ^ s_dadda_pg_rca24_and_18_11;
  assign s_dadda_pg_rca24_fa239_and0 = s_dadda_pg_rca24_and_19_10 & s_dadda_pg_rca24_and_18_11;
  assign s_dadda_pg_rca24_fa239_xor1 = s_dadda_pg_rca24_fa239_xor0 ^ s_dadda_pg_rca24_and_17_12;
  assign s_dadda_pg_rca24_fa239_and1 = s_dadda_pg_rca24_fa239_xor0 & s_dadda_pg_rca24_and_17_12;
  assign s_dadda_pg_rca24_fa239_or0 = s_dadda_pg_rca24_fa239_and0 | s_dadda_pg_rca24_fa239_and1;
  assign s_dadda_pg_rca24_and_16_13 = a[16] & b[13];
  assign s_dadda_pg_rca24_and_15_14 = a[15] & b[14];
  assign s_dadda_pg_rca24_and_14_15 = a[14] & b[15];
  assign s_dadda_pg_rca24_fa240_xor0 = s_dadda_pg_rca24_and_16_13 ^ s_dadda_pg_rca24_and_15_14;
  assign s_dadda_pg_rca24_fa240_and0 = s_dadda_pg_rca24_and_16_13 & s_dadda_pg_rca24_and_15_14;
  assign s_dadda_pg_rca24_fa240_xor1 = s_dadda_pg_rca24_fa240_xor0 ^ s_dadda_pg_rca24_and_14_15;
  assign s_dadda_pg_rca24_fa240_and1 = s_dadda_pg_rca24_fa240_xor0 & s_dadda_pg_rca24_and_14_15;
  assign s_dadda_pg_rca24_fa240_or0 = s_dadda_pg_rca24_fa240_and0 | s_dadda_pg_rca24_fa240_and1;
  assign s_dadda_pg_rca24_and_13_16 = a[13] & b[16];
  assign s_dadda_pg_rca24_and_12_17 = a[12] & b[17];
  assign s_dadda_pg_rca24_and_11_18 = a[11] & b[18];
  assign s_dadda_pg_rca24_fa241_xor0 = s_dadda_pg_rca24_and_13_16 ^ s_dadda_pg_rca24_and_12_17;
  assign s_dadda_pg_rca24_fa241_and0 = s_dadda_pg_rca24_and_13_16 & s_dadda_pg_rca24_and_12_17;
  assign s_dadda_pg_rca24_fa241_xor1 = s_dadda_pg_rca24_fa241_xor0 ^ s_dadda_pg_rca24_and_11_18;
  assign s_dadda_pg_rca24_fa241_and1 = s_dadda_pg_rca24_fa241_xor0 & s_dadda_pg_rca24_and_11_18;
  assign s_dadda_pg_rca24_fa241_or0 = s_dadda_pg_rca24_fa241_and0 | s_dadda_pg_rca24_fa241_and1;
  assign s_dadda_pg_rca24_and_10_19 = a[10] & b[19];
  assign s_dadda_pg_rca24_and_9_20 = a[9] & b[20];
  assign s_dadda_pg_rca24_and_8_21 = a[8] & b[21];
  assign s_dadda_pg_rca24_fa242_xor0 = s_dadda_pg_rca24_and_10_19 ^ s_dadda_pg_rca24_and_9_20;
  assign s_dadda_pg_rca24_fa242_and0 = s_dadda_pg_rca24_and_10_19 & s_dadda_pg_rca24_and_9_20;
  assign s_dadda_pg_rca24_fa242_xor1 = s_dadda_pg_rca24_fa242_xor0 ^ s_dadda_pg_rca24_and_8_21;
  assign s_dadda_pg_rca24_fa242_and1 = s_dadda_pg_rca24_fa242_xor0 & s_dadda_pg_rca24_and_8_21;
  assign s_dadda_pg_rca24_fa242_or0 = s_dadda_pg_rca24_fa242_and0 | s_dadda_pg_rca24_fa242_and1;
  assign s_dadda_pg_rca24_and_7_22 = a[7] & b[22];
  assign s_dadda_pg_rca24_nand_6_23 = ~(a[6] & b[23]);
  assign s_dadda_pg_rca24_fa243_xor0 = s_dadda_pg_rca24_and_7_22 ^ s_dadda_pg_rca24_nand_6_23;
  assign s_dadda_pg_rca24_fa243_and0 = s_dadda_pg_rca24_and_7_22 & s_dadda_pg_rca24_nand_6_23;
  assign s_dadda_pg_rca24_fa243_xor1 = s_dadda_pg_rca24_fa243_xor0 ^ s_dadda_pg_rca24_fa233_xor1;
  assign s_dadda_pg_rca24_fa243_and1 = s_dadda_pg_rca24_fa243_xor0 & s_dadda_pg_rca24_fa233_xor1;
  assign s_dadda_pg_rca24_fa243_or0 = s_dadda_pg_rca24_fa243_and0 | s_dadda_pg_rca24_fa243_and1;
  assign s_dadda_pg_rca24_fa244_xor0 = s_dadda_pg_rca24_fa234_xor1 ^ s_dadda_pg_rca24_fa235_xor1;
  assign s_dadda_pg_rca24_fa244_and0 = s_dadda_pg_rca24_fa234_xor1 & s_dadda_pg_rca24_fa235_xor1;
  assign s_dadda_pg_rca24_fa244_xor1 = s_dadda_pg_rca24_fa244_xor0 ^ s_dadda_pg_rca24_fa236_xor1;
  assign s_dadda_pg_rca24_fa244_and1 = s_dadda_pg_rca24_fa244_xor0 & s_dadda_pg_rca24_fa236_xor1;
  assign s_dadda_pg_rca24_fa244_or0 = s_dadda_pg_rca24_fa244_and0 | s_dadda_pg_rca24_fa244_and1;
  assign s_dadda_pg_rca24_fa245_xor0 = s_dadda_pg_rca24_fa237_xor1 ^ s_dadda_pg_rca24_fa238_xor1;
  assign s_dadda_pg_rca24_fa245_and0 = s_dadda_pg_rca24_fa237_xor1 & s_dadda_pg_rca24_fa238_xor1;
  assign s_dadda_pg_rca24_fa245_xor1 = s_dadda_pg_rca24_fa245_xor0 ^ s_dadda_pg_rca24_fa239_xor1;
  assign s_dadda_pg_rca24_fa245_and1 = s_dadda_pg_rca24_fa245_xor0 & s_dadda_pg_rca24_fa239_xor1;
  assign s_dadda_pg_rca24_fa245_or0 = s_dadda_pg_rca24_fa245_and0 | s_dadda_pg_rca24_fa245_and1;
  assign s_dadda_pg_rca24_fa246_xor0 = s_dadda_pg_rca24_fa245_or0 ^ s_dadda_pg_rca24_fa244_or0;
  assign s_dadda_pg_rca24_fa246_and0 = s_dadda_pg_rca24_fa245_or0 & s_dadda_pg_rca24_fa244_or0;
  assign s_dadda_pg_rca24_fa246_xor1 = s_dadda_pg_rca24_fa246_xor0 ^ s_dadda_pg_rca24_fa243_or0;
  assign s_dadda_pg_rca24_fa246_and1 = s_dadda_pg_rca24_fa246_xor0 & s_dadda_pg_rca24_fa243_or0;
  assign s_dadda_pg_rca24_fa246_or0 = s_dadda_pg_rca24_fa246_and0 | s_dadda_pg_rca24_fa246_and1;
  assign s_dadda_pg_rca24_fa247_xor0 = s_dadda_pg_rca24_fa242_or0 ^ s_dadda_pg_rca24_fa241_or0;
  assign s_dadda_pg_rca24_fa247_and0 = s_dadda_pg_rca24_fa242_or0 & s_dadda_pg_rca24_fa241_or0;
  assign s_dadda_pg_rca24_fa247_xor1 = s_dadda_pg_rca24_fa247_xor0 ^ s_dadda_pg_rca24_fa240_or0;
  assign s_dadda_pg_rca24_fa247_and1 = s_dadda_pg_rca24_fa247_xor0 & s_dadda_pg_rca24_fa240_or0;
  assign s_dadda_pg_rca24_fa247_or0 = s_dadda_pg_rca24_fa247_and0 | s_dadda_pg_rca24_fa247_and1;
  assign s_dadda_pg_rca24_fa248_xor0 = s_dadda_pg_rca24_fa239_or0 ^ s_dadda_pg_rca24_fa238_or0;
  assign s_dadda_pg_rca24_fa248_and0 = s_dadda_pg_rca24_fa239_or0 & s_dadda_pg_rca24_fa238_or0;
  assign s_dadda_pg_rca24_fa248_xor1 = s_dadda_pg_rca24_fa248_xor0 ^ s_dadda_pg_rca24_fa237_or0;
  assign s_dadda_pg_rca24_fa248_and1 = s_dadda_pg_rca24_fa248_xor0 & s_dadda_pg_rca24_fa237_or0;
  assign s_dadda_pg_rca24_fa248_or0 = s_dadda_pg_rca24_fa248_and0 | s_dadda_pg_rca24_fa248_and1;
  assign s_dadda_pg_rca24_fa249_xor0 = s_dadda_pg_rca24_fa236_or0 ^ s_dadda_pg_rca24_fa235_or0;
  assign s_dadda_pg_rca24_fa249_and0 = s_dadda_pg_rca24_fa236_or0 & s_dadda_pg_rca24_fa235_or0;
  assign s_dadda_pg_rca24_fa249_xor1 = s_dadda_pg_rca24_fa249_xor0 ^ s_dadda_pg_rca24_fa234_or0;
  assign s_dadda_pg_rca24_fa249_and1 = s_dadda_pg_rca24_fa249_xor0 & s_dadda_pg_rca24_fa234_or0;
  assign s_dadda_pg_rca24_fa249_or0 = s_dadda_pg_rca24_fa249_and0 | s_dadda_pg_rca24_fa249_and1;
  assign s_dadda_pg_rca24_nand_23_7 = ~(a[23] & b[7]);
  assign s_dadda_pg_rca24_and_22_8 = a[22] & b[8];
  assign s_dadda_pg_rca24_fa250_xor0 = s_dadda_pg_rca24_fa233_or0 ^ s_dadda_pg_rca24_nand_23_7;
  assign s_dadda_pg_rca24_fa250_and0 = s_dadda_pg_rca24_fa233_or0 & s_dadda_pg_rca24_nand_23_7;
  assign s_dadda_pg_rca24_fa250_xor1 = s_dadda_pg_rca24_fa250_xor0 ^ s_dadda_pg_rca24_and_22_8;
  assign s_dadda_pg_rca24_fa250_and1 = s_dadda_pg_rca24_fa250_xor0 & s_dadda_pg_rca24_and_22_8;
  assign s_dadda_pg_rca24_fa250_or0 = s_dadda_pg_rca24_fa250_and0 | s_dadda_pg_rca24_fa250_and1;
  assign s_dadda_pg_rca24_and_21_9 = a[21] & b[9];
  assign s_dadda_pg_rca24_and_20_10 = a[20] & b[10];
  assign s_dadda_pg_rca24_and_19_11 = a[19] & b[11];
  assign s_dadda_pg_rca24_fa251_xor0 = s_dadda_pg_rca24_and_21_9 ^ s_dadda_pg_rca24_and_20_10;
  assign s_dadda_pg_rca24_fa251_and0 = s_dadda_pg_rca24_and_21_9 & s_dadda_pg_rca24_and_20_10;
  assign s_dadda_pg_rca24_fa251_xor1 = s_dadda_pg_rca24_fa251_xor0 ^ s_dadda_pg_rca24_and_19_11;
  assign s_dadda_pg_rca24_fa251_and1 = s_dadda_pg_rca24_fa251_xor0 & s_dadda_pg_rca24_and_19_11;
  assign s_dadda_pg_rca24_fa251_or0 = s_dadda_pg_rca24_fa251_and0 | s_dadda_pg_rca24_fa251_and1;
  assign s_dadda_pg_rca24_and_18_12 = a[18] & b[12];
  assign s_dadda_pg_rca24_and_17_13 = a[17] & b[13];
  assign s_dadda_pg_rca24_and_16_14 = a[16] & b[14];
  assign s_dadda_pg_rca24_fa252_xor0 = s_dadda_pg_rca24_and_18_12 ^ s_dadda_pg_rca24_and_17_13;
  assign s_dadda_pg_rca24_fa252_and0 = s_dadda_pg_rca24_and_18_12 & s_dadda_pg_rca24_and_17_13;
  assign s_dadda_pg_rca24_fa252_xor1 = s_dadda_pg_rca24_fa252_xor0 ^ s_dadda_pg_rca24_and_16_14;
  assign s_dadda_pg_rca24_fa252_and1 = s_dadda_pg_rca24_fa252_xor0 & s_dadda_pg_rca24_and_16_14;
  assign s_dadda_pg_rca24_fa252_or0 = s_dadda_pg_rca24_fa252_and0 | s_dadda_pg_rca24_fa252_and1;
  assign s_dadda_pg_rca24_and_15_15 = a[15] & b[15];
  assign s_dadda_pg_rca24_and_14_16 = a[14] & b[16];
  assign s_dadda_pg_rca24_and_13_17 = a[13] & b[17];
  assign s_dadda_pg_rca24_fa253_xor0 = s_dadda_pg_rca24_and_15_15 ^ s_dadda_pg_rca24_and_14_16;
  assign s_dadda_pg_rca24_fa253_and0 = s_dadda_pg_rca24_and_15_15 & s_dadda_pg_rca24_and_14_16;
  assign s_dadda_pg_rca24_fa253_xor1 = s_dadda_pg_rca24_fa253_xor0 ^ s_dadda_pg_rca24_and_13_17;
  assign s_dadda_pg_rca24_fa253_and1 = s_dadda_pg_rca24_fa253_xor0 & s_dadda_pg_rca24_and_13_17;
  assign s_dadda_pg_rca24_fa253_or0 = s_dadda_pg_rca24_fa253_and0 | s_dadda_pg_rca24_fa253_and1;
  assign s_dadda_pg_rca24_and_12_18 = a[12] & b[18];
  assign s_dadda_pg_rca24_and_11_19 = a[11] & b[19];
  assign s_dadda_pg_rca24_and_10_20 = a[10] & b[20];
  assign s_dadda_pg_rca24_fa254_xor0 = s_dadda_pg_rca24_and_12_18 ^ s_dadda_pg_rca24_and_11_19;
  assign s_dadda_pg_rca24_fa254_and0 = s_dadda_pg_rca24_and_12_18 & s_dadda_pg_rca24_and_11_19;
  assign s_dadda_pg_rca24_fa254_xor1 = s_dadda_pg_rca24_fa254_xor0 ^ s_dadda_pg_rca24_and_10_20;
  assign s_dadda_pg_rca24_fa254_and1 = s_dadda_pg_rca24_fa254_xor0 & s_dadda_pg_rca24_and_10_20;
  assign s_dadda_pg_rca24_fa254_or0 = s_dadda_pg_rca24_fa254_and0 | s_dadda_pg_rca24_fa254_and1;
  assign s_dadda_pg_rca24_and_9_21 = a[9] & b[21];
  assign s_dadda_pg_rca24_and_8_22 = a[8] & b[22];
  assign s_dadda_pg_rca24_nand_7_23 = ~(a[7] & b[23]);
  assign s_dadda_pg_rca24_fa255_xor0 = s_dadda_pg_rca24_and_9_21 ^ s_dadda_pg_rca24_and_8_22;
  assign s_dadda_pg_rca24_fa255_and0 = s_dadda_pg_rca24_and_9_21 & s_dadda_pg_rca24_and_8_22;
  assign s_dadda_pg_rca24_fa255_xor1 = s_dadda_pg_rca24_fa255_xor0 ^ s_dadda_pg_rca24_nand_7_23;
  assign s_dadda_pg_rca24_fa255_and1 = s_dadda_pg_rca24_fa255_xor0 & s_dadda_pg_rca24_nand_7_23;
  assign s_dadda_pg_rca24_fa255_or0 = s_dadda_pg_rca24_fa255_and0 | s_dadda_pg_rca24_fa255_and1;
  assign s_dadda_pg_rca24_fa256_xor0 = s_dadda_pg_rca24_fa246_xor1 ^ s_dadda_pg_rca24_fa247_xor1;
  assign s_dadda_pg_rca24_fa256_and0 = s_dadda_pg_rca24_fa246_xor1 & s_dadda_pg_rca24_fa247_xor1;
  assign s_dadda_pg_rca24_fa256_xor1 = s_dadda_pg_rca24_fa256_xor0 ^ s_dadda_pg_rca24_fa248_xor1;
  assign s_dadda_pg_rca24_fa256_and1 = s_dadda_pg_rca24_fa256_xor0 & s_dadda_pg_rca24_fa248_xor1;
  assign s_dadda_pg_rca24_fa256_or0 = s_dadda_pg_rca24_fa256_and0 | s_dadda_pg_rca24_fa256_and1;
  assign s_dadda_pg_rca24_fa257_xor0 = s_dadda_pg_rca24_fa249_xor1 ^ s_dadda_pg_rca24_fa250_xor1;
  assign s_dadda_pg_rca24_fa257_and0 = s_dadda_pg_rca24_fa249_xor1 & s_dadda_pg_rca24_fa250_xor1;
  assign s_dadda_pg_rca24_fa257_xor1 = s_dadda_pg_rca24_fa257_xor0 ^ s_dadda_pg_rca24_fa251_xor1;
  assign s_dadda_pg_rca24_fa257_and1 = s_dadda_pg_rca24_fa257_xor0 & s_dadda_pg_rca24_fa251_xor1;
  assign s_dadda_pg_rca24_fa257_or0 = s_dadda_pg_rca24_fa257_and0 | s_dadda_pg_rca24_fa257_and1;
  assign s_dadda_pg_rca24_fa258_xor0 = s_dadda_pg_rca24_fa257_or0 ^ s_dadda_pg_rca24_fa256_or0;
  assign s_dadda_pg_rca24_fa258_and0 = s_dadda_pg_rca24_fa257_or0 & s_dadda_pg_rca24_fa256_or0;
  assign s_dadda_pg_rca24_fa258_xor1 = s_dadda_pg_rca24_fa258_xor0 ^ s_dadda_pg_rca24_fa255_or0;
  assign s_dadda_pg_rca24_fa258_and1 = s_dadda_pg_rca24_fa258_xor0 & s_dadda_pg_rca24_fa255_or0;
  assign s_dadda_pg_rca24_fa258_or0 = s_dadda_pg_rca24_fa258_and0 | s_dadda_pg_rca24_fa258_and1;
  assign s_dadda_pg_rca24_fa259_xor0 = s_dadda_pg_rca24_fa254_or0 ^ s_dadda_pg_rca24_fa253_or0;
  assign s_dadda_pg_rca24_fa259_and0 = s_dadda_pg_rca24_fa254_or0 & s_dadda_pg_rca24_fa253_or0;
  assign s_dadda_pg_rca24_fa259_xor1 = s_dadda_pg_rca24_fa259_xor0 ^ s_dadda_pg_rca24_fa252_or0;
  assign s_dadda_pg_rca24_fa259_and1 = s_dadda_pg_rca24_fa259_xor0 & s_dadda_pg_rca24_fa252_or0;
  assign s_dadda_pg_rca24_fa259_or0 = s_dadda_pg_rca24_fa259_and0 | s_dadda_pg_rca24_fa259_and1;
  assign s_dadda_pg_rca24_fa260_xor0 = s_dadda_pg_rca24_fa251_or0 ^ s_dadda_pg_rca24_fa250_or0;
  assign s_dadda_pg_rca24_fa260_and0 = s_dadda_pg_rca24_fa251_or0 & s_dadda_pg_rca24_fa250_or0;
  assign s_dadda_pg_rca24_fa260_xor1 = s_dadda_pg_rca24_fa260_xor0 ^ s_dadda_pg_rca24_fa249_or0;
  assign s_dadda_pg_rca24_fa260_and1 = s_dadda_pg_rca24_fa260_xor0 & s_dadda_pg_rca24_fa249_or0;
  assign s_dadda_pg_rca24_fa260_or0 = s_dadda_pg_rca24_fa260_and0 | s_dadda_pg_rca24_fa260_and1;
  assign s_dadda_pg_rca24_fa261_xor0 = s_dadda_pg_rca24_fa248_or0 ^ s_dadda_pg_rca24_fa247_or0;
  assign s_dadda_pg_rca24_fa261_and0 = s_dadda_pg_rca24_fa248_or0 & s_dadda_pg_rca24_fa247_or0;
  assign s_dadda_pg_rca24_fa261_xor1 = s_dadda_pg_rca24_fa261_xor0 ^ s_dadda_pg_rca24_fa246_or0;
  assign s_dadda_pg_rca24_fa261_and1 = s_dadda_pg_rca24_fa261_xor0 & s_dadda_pg_rca24_fa246_or0;
  assign s_dadda_pg_rca24_fa261_or0 = s_dadda_pg_rca24_fa261_and0 | s_dadda_pg_rca24_fa261_and1;
  assign s_dadda_pg_rca24_nand_23_8 = ~(a[23] & b[8]);
  assign s_dadda_pg_rca24_and_22_9 = a[22] & b[9];
  assign s_dadda_pg_rca24_and_21_10 = a[21] & b[10];
  assign s_dadda_pg_rca24_fa262_xor0 = s_dadda_pg_rca24_nand_23_8 ^ s_dadda_pg_rca24_and_22_9;
  assign s_dadda_pg_rca24_fa262_and0 = s_dadda_pg_rca24_nand_23_8 & s_dadda_pg_rca24_and_22_9;
  assign s_dadda_pg_rca24_fa262_xor1 = s_dadda_pg_rca24_fa262_xor0 ^ s_dadda_pg_rca24_and_21_10;
  assign s_dadda_pg_rca24_fa262_and1 = s_dadda_pg_rca24_fa262_xor0 & s_dadda_pg_rca24_and_21_10;
  assign s_dadda_pg_rca24_fa262_or0 = s_dadda_pg_rca24_fa262_and0 | s_dadda_pg_rca24_fa262_and1;
  assign s_dadda_pg_rca24_and_20_11 = a[20] & b[11];
  assign s_dadda_pg_rca24_and_19_12 = a[19] & b[12];
  assign s_dadda_pg_rca24_and_18_13 = a[18] & b[13];
  assign s_dadda_pg_rca24_fa263_xor0 = s_dadda_pg_rca24_and_20_11 ^ s_dadda_pg_rca24_and_19_12;
  assign s_dadda_pg_rca24_fa263_and0 = s_dadda_pg_rca24_and_20_11 & s_dadda_pg_rca24_and_19_12;
  assign s_dadda_pg_rca24_fa263_xor1 = s_dadda_pg_rca24_fa263_xor0 ^ s_dadda_pg_rca24_and_18_13;
  assign s_dadda_pg_rca24_fa263_and1 = s_dadda_pg_rca24_fa263_xor0 & s_dadda_pg_rca24_and_18_13;
  assign s_dadda_pg_rca24_fa263_or0 = s_dadda_pg_rca24_fa263_and0 | s_dadda_pg_rca24_fa263_and1;
  assign s_dadda_pg_rca24_and_17_14 = a[17] & b[14];
  assign s_dadda_pg_rca24_and_16_15 = a[16] & b[15];
  assign s_dadda_pg_rca24_and_15_16 = a[15] & b[16];
  assign s_dadda_pg_rca24_fa264_xor0 = s_dadda_pg_rca24_and_17_14 ^ s_dadda_pg_rca24_and_16_15;
  assign s_dadda_pg_rca24_fa264_and0 = s_dadda_pg_rca24_and_17_14 & s_dadda_pg_rca24_and_16_15;
  assign s_dadda_pg_rca24_fa264_xor1 = s_dadda_pg_rca24_fa264_xor0 ^ s_dadda_pg_rca24_and_15_16;
  assign s_dadda_pg_rca24_fa264_and1 = s_dadda_pg_rca24_fa264_xor0 & s_dadda_pg_rca24_and_15_16;
  assign s_dadda_pg_rca24_fa264_or0 = s_dadda_pg_rca24_fa264_and0 | s_dadda_pg_rca24_fa264_and1;
  assign s_dadda_pg_rca24_and_14_17 = a[14] & b[17];
  assign s_dadda_pg_rca24_and_13_18 = a[13] & b[18];
  assign s_dadda_pg_rca24_and_12_19 = a[12] & b[19];
  assign s_dadda_pg_rca24_fa265_xor0 = s_dadda_pg_rca24_and_14_17 ^ s_dadda_pg_rca24_and_13_18;
  assign s_dadda_pg_rca24_fa265_and0 = s_dadda_pg_rca24_and_14_17 & s_dadda_pg_rca24_and_13_18;
  assign s_dadda_pg_rca24_fa265_xor1 = s_dadda_pg_rca24_fa265_xor0 ^ s_dadda_pg_rca24_and_12_19;
  assign s_dadda_pg_rca24_fa265_and1 = s_dadda_pg_rca24_fa265_xor0 & s_dadda_pg_rca24_and_12_19;
  assign s_dadda_pg_rca24_fa265_or0 = s_dadda_pg_rca24_fa265_and0 | s_dadda_pg_rca24_fa265_and1;
  assign s_dadda_pg_rca24_and_11_20 = a[11] & b[20];
  assign s_dadda_pg_rca24_and_10_21 = a[10] & b[21];
  assign s_dadda_pg_rca24_and_9_22 = a[9] & b[22];
  assign s_dadda_pg_rca24_fa266_xor0 = s_dadda_pg_rca24_and_11_20 ^ s_dadda_pg_rca24_and_10_21;
  assign s_dadda_pg_rca24_fa266_and0 = s_dadda_pg_rca24_and_11_20 & s_dadda_pg_rca24_and_10_21;
  assign s_dadda_pg_rca24_fa266_xor1 = s_dadda_pg_rca24_fa266_xor0 ^ s_dadda_pg_rca24_and_9_22;
  assign s_dadda_pg_rca24_fa266_and1 = s_dadda_pg_rca24_fa266_xor0 & s_dadda_pg_rca24_and_9_22;
  assign s_dadda_pg_rca24_fa266_or0 = s_dadda_pg_rca24_fa266_and0 | s_dadda_pg_rca24_fa266_and1;
  assign s_dadda_pg_rca24_nand_8_23 = ~(a[8] & b[23]);
  assign s_dadda_pg_rca24_fa267_xor0 = s_dadda_pg_rca24_nand_8_23 ^ s_dadda_pg_rca24_fa258_xor1;
  assign s_dadda_pg_rca24_fa267_and0 = s_dadda_pg_rca24_nand_8_23 & s_dadda_pg_rca24_fa258_xor1;
  assign s_dadda_pg_rca24_fa267_xor1 = s_dadda_pg_rca24_fa267_xor0 ^ s_dadda_pg_rca24_fa259_xor1;
  assign s_dadda_pg_rca24_fa267_and1 = s_dadda_pg_rca24_fa267_xor0 & s_dadda_pg_rca24_fa259_xor1;
  assign s_dadda_pg_rca24_fa267_or0 = s_dadda_pg_rca24_fa267_and0 | s_dadda_pg_rca24_fa267_and1;
  assign s_dadda_pg_rca24_fa268_xor0 = s_dadda_pg_rca24_fa260_xor1 ^ s_dadda_pg_rca24_fa261_xor1;
  assign s_dadda_pg_rca24_fa268_and0 = s_dadda_pg_rca24_fa260_xor1 & s_dadda_pg_rca24_fa261_xor1;
  assign s_dadda_pg_rca24_fa268_xor1 = s_dadda_pg_rca24_fa268_xor0 ^ s_dadda_pg_rca24_fa262_xor1;
  assign s_dadda_pg_rca24_fa268_and1 = s_dadda_pg_rca24_fa268_xor0 & s_dadda_pg_rca24_fa262_xor1;
  assign s_dadda_pg_rca24_fa268_or0 = s_dadda_pg_rca24_fa268_and0 | s_dadda_pg_rca24_fa268_and1;
  assign s_dadda_pg_rca24_fa269_xor0 = s_dadda_pg_rca24_fa268_or0 ^ s_dadda_pg_rca24_fa267_or0;
  assign s_dadda_pg_rca24_fa269_and0 = s_dadda_pg_rca24_fa268_or0 & s_dadda_pg_rca24_fa267_or0;
  assign s_dadda_pg_rca24_fa269_xor1 = s_dadda_pg_rca24_fa269_xor0 ^ s_dadda_pg_rca24_fa266_or0;
  assign s_dadda_pg_rca24_fa269_and1 = s_dadda_pg_rca24_fa269_xor0 & s_dadda_pg_rca24_fa266_or0;
  assign s_dadda_pg_rca24_fa269_or0 = s_dadda_pg_rca24_fa269_and0 | s_dadda_pg_rca24_fa269_and1;
  assign s_dadda_pg_rca24_fa270_xor0 = s_dadda_pg_rca24_fa265_or0 ^ s_dadda_pg_rca24_fa264_or0;
  assign s_dadda_pg_rca24_fa270_and0 = s_dadda_pg_rca24_fa265_or0 & s_dadda_pg_rca24_fa264_or0;
  assign s_dadda_pg_rca24_fa270_xor1 = s_dadda_pg_rca24_fa270_xor0 ^ s_dadda_pg_rca24_fa263_or0;
  assign s_dadda_pg_rca24_fa270_and1 = s_dadda_pg_rca24_fa270_xor0 & s_dadda_pg_rca24_fa263_or0;
  assign s_dadda_pg_rca24_fa270_or0 = s_dadda_pg_rca24_fa270_and0 | s_dadda_pg_rca24_fa270_and1;
  assign s_dadda_pg_rca24_fa271_xor0 = s_dadda_pg_rca24_fa262_or0 ^ s_dadda_pg_rca24_fa261_or0;
  assign s_dadda_pg_rca24_fa271_and0 = s_dadda_pg_rca24_fa262_or0 & s_dadda_pg_rca24_fa261_or0;
  assign s_dadda_pg_rca24_fa271_xor1 = s_dadda_pg_rca24_fa271_xor0 ^ s_dadda_pg_rca24_fa260_or0;
  assign s_dadda_pg_rca24_fa271_and1 = s_dadda_pg_rca24_fa271_xor0 & s_dadda_pg_rca24_fa260_or0;
  assign s_dadda_pg_rca24_fa271_or0 = s_dadda_pg_rca24_fa271_and0 | s_dadda_pg_rca24_fa271_and1;
  assign s_dadda_pg_rca24_nand_23_9 = ~(a[23] & b[9]);
  assign s_dadda_pg_rca24_fa272_xor0 = s_dadda_pg_rca24_fa259_or0 ^ s_dadda_pg_rca24_fa258_or0;
  assign s_dadda_pg_rca24_fa272_and0 = s_dadda_pg_rca24_fa259_or0 & s_dadda_pg_rca24_fa258_or0;
  assign s_dadda_pg_rca24_fa272_xor1 = s_dadda_pg_rca24_fa272_xor0 ^ s_dadda_pg_rca24_nand_23_9;
  assign s_dadda_pg_rca24_fa272_and1 = s_dadda_pg_rca24_fa272_xor0 & s_dadda_pg_rca24_nand_23_9;
  assign s_dadda_pg_rca24_fa272_or0 = s_dadda_pg_rca24_fa272_and0 | s_dadda_pg_rca24_fa272_and1;
  assign s_dadda_pg_rca24_and_22_10 = a[22] & b[10];
  assign s_dadda_pg_rca24_and_21_11 = a[21] & b[11];
  assign s_dadda_pg_rca24_and_20_12 = a[20] & b[12];
  assign s_dadda_pg_rca24_fa273_xor0 = s_dadda_pg_rca24_and_22_10 ^ s_dadda_pg_rca24_and_21_11;
  assign s_dadda_pg_rca24_fa273_and0 = s_dadda_pg_rca24_and_22_10 & s_dadda_pg_rca24_and_21_11;
  assign s_dadda_pg_rca24_fa273_xor1 = s_dadda_pg_rca24_fa273_xor0 ^ s_dadda_pg_rca24_and_20_12;
  assign s_dadda_pg_rca24_fa273_and1 = s_dadda_pg_rca24_fa273_xor0 & s_dadda_pg_rca24_and_20_12;
  assign s_dadda_pg_rca24_fa273_or0 = s_dadda_pg_rca24_fa273_and0 | s_dadda_pg_rca24_fa273_and1;
  assign s_dadda_pg_rca24_and_19_13 = a[19] & b[13];
  assign s_dadda_pg_rca24_and_18_14 = a[18] & b[14];
  assign s_dadda_pg_rca24_and_17_15 = a[17] & b[15];
  assign s_dadda_pg_rca24_fa274_xor0 = s_dadda_pg_rca24_and_19_13 ^ s_dadda_pg_rca24_and_18_14;
  assign s_dadda_pg_rca24_fa274_and0 = s_dadda_pg_rca24_and_19_13 & s_dadda_pg_rca24_and_18_14;
  assign s_dadda_pg_rca24_fa274_xor1 = s_dadda_pg_rca24_fa274_xor0 ^ s_dadda_pg_rca24_and_17_15;
  assign s_dadda_pg_rca24_fa274_and1 = s_dadda_pg_rca24_fa274_xor0 & s_dadda_pg_rca24_and_17_15;
  assign s_dadda_pg_rca24_fa274_or0 = s_dadda_pg_rca24_fa274_and0 | s_dadda_pg_rca24_fa274_and1;
  assign s_dadda_pg_rca24_and_16_16 = a[16] & b[16];
  assign s_dadda_pg_rca24_and_15_17 = a[15] & b[17];
  assign s_dadda_pg_rca24_and_14_18 = a[14] & b[18];
  assign s_dadda_pg_rca24_fa275_xor0 = s_dadda_pg_rca24_and_16_16 ^ s_dadda_pg_rca24_and_15_17;
  assign s_dadda_pg_rca24_fa275_and0 = s_dadda_pg_rca24_and_16_16 & s_dadda_pg_rca24_and_15_17;
  assign s_dadda_pg_rca24_fa275_xor1 = s_dadda_pg_rca24_fa275_xor0 ^ s_dadda_pg_rca24_and_14_18;
  assign s_dadda_pg_rca24_fa275_and1 = s_dadda_pg_rca24_fa275_xor0 & s_dadda_pg_rca24_and_14_18;
  assign s_dadda_pg_rca24_fa275_or0 = s_dadda_pg_rca24_fa275_and0 | s_dadda_pg_rca24_fa275_and1;
  assign s_dadda_pg_rca24_and_13_19 = a[13] & b[19];
  assign s_dadda_pg_rca24_and_12_20 = a[12] & b[20];
  assign s_dadda_pg_rca24_and_11_21 = a[11] & b[21];
  assign s_dadda_pg_rca24_fa276_xor0 = s_dadda_pg_rca24_and_13_19 ^ s_dadda_pg_rca24_and_12_20;
  assign s_dadda_pg_rca24_fa276_and0 = s_dadda_pg_rca24_and_13_19 & s_dadda_pg_rca24_and_12_20;
  assign s_dadda_pg_rca24_fa276_xor1 = s_dadda_pg_rca24_fa276_xor0 ^ s_dadda_pg_rca24_and_11_21;
  assign s_dadda_pg_rca24_fa276_and1 = s_dadda_pg_rca24_fa276_xor0 & s_dadda_pg_rca24_and_11_21;
  assign s_dadda_pg_rca24_fa276_or0 = s_dadda_pg_rca24_fa276_and0 | s_dadda_pg_rca24_fa276_and1;
  assign s_dadda_pg_rca24_and_10_22 = a[10] & b[22];
  assign s_dadda_pg_rca24_nand_9_23 = ~(a[9] & b[23]);
  assign s_dadda_pg_rca24_fa277_xor0 = s_dadda_pg_rca24_and_10_22 ^ s_dadda_pg_rca24_nand_9_23;
  assign s_dadda_pg_rca24_fa277_and0 = s_dadda_pg_rca24_and_10_22 & s_dadda_pg_rca24_nand_9_23;
  assign s_dadda_pg_rca24_fa277_xor1 = s_dadda_pg_rca24_fa277_xor0 ^ s_dadda_pg_rca24_fa269_xor1;
  assign s_dadda_pg_rca24_fa277_and1 = s_dadda_pg_rca24_fa277_xor0 & s_dadda_pg_rca24_fa269_xor1;
  assign s_dadda_pg_rca24_fa277_or0 = s_dadda_pg_rca24_fa277_and0 | s_dadda_pg_rca24_fa277_and1;
  assign s_dadda_pg_rca24_fa278_xor0 = s_dadda_pg_rca24_fa270_xor1 ^ s_dadda_pg_rca24_fa271_xor1;
  assign s_dadda_pg_rca24_fa278_and0 = s_dadda_pg_rca24_fa270_xor1 & s_dadda_pg_rca24_fa271_xor1;
  assign s_dadda_pg_rca24_fa278_xor1 = s_dadda_pg_rca24_fa278_xor0 ^ s_dadda_pg_rca24_fa272_xor1;
  assign s_dadda_pg_rca24_fa278_and1 = s_dadda_pg_rca24_fa278_xor0 & s_dadda_pg_rca24_fa272_xor1;
  assign s_dadda_pg_rca24_fa278_or0 = s_dadda_pg_rca24_fa278_and0 | s_dadda_pg_rca24_fa278_and1;
  assign s_dadda_pg_rca24_fa279_xor0 = s_dadda_pg_rca24_fa278_or0 ^ s_dadda_pg_rca24_fa277_or0;
  assign s_dadda_pg_rca24_fa279_and0 = s_dadda_pg_rca24_fa278_or0 & s_dadda_pg_rca24_fa277_or0;
  assign s_dadda_pg_rca24_fa279_xor1 = s_dadda_pg_rca24_fa279_xor0 ^ s_dadda_pg_rca24_fa276_or0;
  assign s_dadda_pg_rca24_fa279_and1 = s_dadda_pg_rca24_fa279_xor0 & s_dadda_pg_rca24_fa276_or0;
  assign s_dadda_pg_rca24_fa279_or0 = s_dadda_pg_rca24_fa279_and0 | s_dadda_pg_rca24_fa279_and1;
  assign s_dadda_pg_rca24_fa280_xor0 = s_dadda_pg_rca24_fa275_or0 ^ s_dadda_pg_rca24_fa274_or0;
  assign s_dadda_pg_rca24_fa280_and0 = s_dadda_pg_rca24_fa275_or0 & s_dadda_pg_rca24_fa274_or0;
  assign s_dadda_pg_rca24_fa280_xor1 = s_dadda_pg_rca24_fa280_xor0 ^ s_dadda_pg_rca24_fa273_or0;
  assign s_dadda_pg_rca24_fa280_and1 = s_dadda_pg_rca24_fa280_xor0 & s_dadda_pg_rca24_fa273_or0;
  assign s_dadda_pg_rca24_fa280_or0 = s_dadda_pg_rca24_fa280_and0 | s_dadda_pg_rca24_fa280_and1;
  assign s_dadda_pg_rca24_fa281_xor0 = s_dadda_pg_rca24_fa272_or0 ^ s_dadda_pg_rca24_fa271_or0;
  assign s_dadda_pg_rca24_fa281_and0 = s_dadda_pg_rca24_fa272_or0 & s_dadda_pg_rca24_fa271_or0;
  assign s_dadda_pg_rca24_fa281_xor1 = s_dadda_pg_rca24_fa281_xor0 ^ s_dadda_pg_rca24_fa270_or0;
  assign s_dadda_pg_rca24_fa281_and1 = s_dadda_pg_rca24_fa281_xor0 & s_dadda_pg_rca24_fa270_or0;
  assign s_dadda_pg_rca24_fa281_or0 = s_dadda_pg_rca24_fa281_and0 | s_dadda_pg_rca24_fa281_and1;
  assign s_dadda_pg_rca24_nand_23_10 = ~(a[23] & b[10]);
  assign s_dadda_pg_rca24_and_22_11 = a[22] & b[11];
  assign s_dadda_pg_rca24_fa282_xor0 = s_dadda_pg_rca24_fa269_or0 ^ s_dadda_pg_rca24_nand_23_10;
  assign s_dadda_pg_rca24_fa282_and0 = s_dadda_pg_rca24_fa269_or0 & s_dadda_pg_rca24_nand_23_10;
  assign s_dadda_pg_rca24_fa282_xor1 = s_dadda_pg_rca24_fa282_xor0 ^ s_dadda_pg_rca24_and_22_11;
  assign s_dadda_pg_rca24_fa282_and1 = s_dadda_pg_rca24_fa282_xor0 & s_dadda_pg_rca24_and_22_11;
  assign s_dadda_pg_rca24_fa282_or0 = s_dadda_pg_rca24_fa282_and0 | s_dadda_pg_rca24_fa282_and1;
  assign s_dadda_pg_rca24_and_21_12 = a[21] & b[12];
  assign s_dadda_pg_rca24_and_20_13 = a[20] & b[13];
  assign s_dadda_pg_rca24_and_19_14 = a[19] & b[14];
  assign s_dadda_pg_rca24_fa283_xor0 = s_dadda_pg_rca24_and_21_12 ^ s_dadda_pg_rca24_and_20_13;
  assign s_dadda_pg_rca24_fa283_and0 = s_dadda_pg_rca24_and_21_12 & s_dadda_pg_rca24_and_20_13;
  assign s_dadda_pg_rca24_fa283_xor1 = s_dadda_pg_rca24_fa283_xor0 ^ s_dadda_pg_rca24_and_19_14;
  assign s_dadda_pg_rca24_fa283_and1 = s_dadda_pg_rca24_fa283_xor0 & s_dadda_pg_rca24_and_19_14;
  assign s_dadda_pg_rca24_fa283_or0 = s_dadda_pg_rca24_fa283_and0 | s_dadda_pg_rca24_fa283_and1;
  assign s_dadda_pg_rca24_and_18_15 = a[18] & b[15];
  assign s_dadda_pg_rca24_and_17_16 = a[17] & b[16];
  assign s_dadda_pg_rca24_and_16_17 = a[16] & b[17];
  assign s_dadda_pg_rca24_fa284_xor0 = s_dadda_pg_rca24_and_18_15 ^ s_dadda_pg_rca24_and_17_16;
  assign s_dadda_pg_rca24_fa284_and0 = s_dadda_pg_rca24_and_18_15 & s_dadda_pg_rca24_and_17_16;
  assign s_dadda_pg_rca24_fa284_xor1 = s_dadda_pg_rca24_fa284_xor0 ^ s_dadda_pg_rca24_and_16_17;
  assign s_dadda_pg_rca24_fa284_and1 = s_dadda_pg_rca24_fa284_xor0 & s_dadda_pg_rca24_and_16_17;
  assign s_dadda_pg_rca24_fa284_or0 = s_dadda_pg_rca24_fa284_and0 | s_dadda_pg_rca24_fa284_and1;
  assign s_dadda_pg_rca24_and_15_18 = a[15] & b[18];
  assign s_dadda_pg_rca24_and_14_19 = a[14] & b[19];
  assign s_dadda_pg_rca24_and_13_20 = a[13] & b[20];
  assign s_dadda_pg_rca24_fa285_xor0 = s_dadda_pg_rca24_and_15_18 ^ s_dadda_pg_rca24_and_14_19;
  assign s_dadda_pg_rca24_fa285_and0 = s_dadda_pg_rca24_and_15_18 & s_dadda_pg_rca24_and_14_19;
  assign s_dadda_pg_rca24_fa285_xor1 = s_dadda_pg_rca24_fa285_xor0 ^ s_dadda_pg_rca24_and_13_20;
  assign s_dadda_pg_rca24_fa285_and1 = s_dadda_pg_rca24_fa285_xor0 & s_dadda_pg_rca24_and_13_20;
  assign s_dadda_pg_rca24_fa285_or0 = s_dadda_pg_rca24_fa285_and0 | s_dadda_pg_rca24_fa285_and1;
  assign s_dadda_pg_rca24_and_12_21 = a[12] & b[21];
  assign s_dadda_pg_rca24_and_11_22 = a[11] & b[22];
  assign s_dadda_pg_rca24_nand_10_23 = ~(a[10] & b[23]);
  assign s_dadda_pg_rca24_fa286_xor0 = s_dadda_pg_rca24_and_12_21 ^ s_dadda_pg_rca24_and_11_22;
  assign s_dadda_pg_rca24_fa286_and0 = s_dadda_pg_rca24_and_12_21 & s_dadda_pg_rca24_and_11_22;
  assign s_dadda_pg_rca24_fa286_xor1 = s_dadda_pg_rca24_fa286_xor0 ^ s_dadda_pg_rca24_nand_10_23;
  assign s_dadda_pg_rca24_fa286_and1 = s_dadda_pg_rca24_fa286_xor0 & s_dadda_pg_rca24_nand_10_23;
  assign s_dadda_pg_rca24_fa286_or0 = s_dadda_pg_rca24_fa286_and0 | s_dadda_pg_rca24_fa286_and1;
  assign s_dadda_pg_rca24_fa287_xor0 = s_dadda_pg_rca24_fa279_xor1 ^ s_dadda_pg_rca24_fa280_xor1;
  assign s_dadda_pg_rca24_fa287_and0 = s_dadda_pg_rca24_fa279_xor1 & s_dadda_pg_rca24_fa280_xor1;
  assign s_dadda_pg_rca24_fa287_xor1 = s_dadda_pg_rca24_fa287_xor0 ^ s_dadda_pg_rca24_fa281_xor1;
  assign s_dadda_pg_rca24_fa287_and1 = s_dadda_pg_rca24_fa287_xor0 & s_dadda_pg_rca24_fa281_xor1;
  assign s_dadda_pg_rca24_fa287_or0 = s_dadda_pg_rca24_fa287_and0 | s_dadda_pg_rca24_fa287_and1;
  assign s_dadda_pg_rca24_fa288_xor0 = s_dadda_pg_rca24_fa287_or0 ^ s_dadda_pg_rca24_fa286_or0;
  assign s_dadda_pg_rca24_fa288_and0 = s_dadda_pg_rca24_fa287_or0 & s_dadda_pg_rca24_fa286_or0;
  assign s_dadda_pg_rca24_fa288_xor1 = s_dadda_pg_rca24_fa288_xor0 ^ s_dadda_pg_rca24_fa285_or0;
  assign s_dadda_pg_rca24_fa288_and1 = s_dadda_pg_rca24_fa288_xor0 & s_dadda_pg_rca24_fa285_or0;
  assign s_dadda_pg_rca24_fa288_or0 = s_dadda_pg_rca24_fa288_and0 | s_dadda_pg_rca24_fa288_and1;
  assign s_dadda_pg_rca24_fa289_xor0 = s_dadda_pg_rca24_fa284_or0 ^ s_dadda_pg_rca24_fa283_or0;
  assign s_dadda_pg_rca24_fa289_and0 = s_dadda_pg_rca24_fa284_or0 & s_dadda_pg_rca24_fa283_or0;
  assign s_dadda_pg_rca24_fa289_xor1 = s_dadda_pg_rca24_fa289_xor0 ^ s_dadda_pg_rca24_fa282_or0;
  assign s_dadda_pg_rca24_fa289_and1 = s_dadda_pg_rca24_fa289_xor0 & s_dadda_pg_rca24_fa282_or0;
  assign s_dadda_pg_rca24_fa289_or0 = s_dadda_pg_rca24_fa289_and0 | s_dadda_pg_rca24_fa289_and1;
  assign s_dadda_pg_rca24_fa290_xor0 = s_dadda_pg_rca24_fa281_or0 ^ s_dadda_pg_rca24_fa280_or0;
  assign s_dadda_pg_rca24_fa290_and0 = s_dadda_pg_rca24_fa281_or0 & s_dadda_pg_rca24_fa280_or0;
  assign s_dadda_pg_rca24_fa290_xor1 = s_dadda_pg_rca24_fa290_xor0 ^ s_dadda_pg_rca24_fa279_or0;
  assign s_dadda_pg_rca24_fa290_and1 = s_dadda_pg_rca24_fa290_xor0 & s_dadda_pg_rca24_fa279_or0;
  assign s_dadda_pg_rca24_fa290_or0 = s_dadda_pg_rca24_fa290_and0 | s_dadda_pg_rca24_fa290_and1;
  assign s_dadda_pg_rca24_nand_23_11 = ~(a[23] & b[11]);
  assign s_dadda_pg_rca24_and_22_12 = a[22] & b[12];
  assign s_dadda_pg_rca24_and_21_13 = a[21] & b[13];
  assign s_dadda_pg_rca24_fa291_xor0 = s_dadda_pg_rca24_nand_23_11 ^ s_dadda_pg_rca24_and_22_12;
  assign s_dadda_pg_rca24_fa291_and0 = s_dadda_pg_rca24_nand_23_11 & s_dadda_pg_rca24_and_22_12;
  assign s_dadda_pg_rca24_fa291_xor1 = s_dadda_pg_rca24_fa291_xor0 ^ s_dadda_pg_rca24_and_21_13;
  assign s_dadda_pg_rca24_fa291_and1 = s_dadda_pg_rca24_fa291_xor0 & s_dadda_pg_rca24_and_21_13;
  assign s_dadda_pg_rca24_fa291_or0 = s_dadda_pg_rca24_fa291_and0 | s_dadda_pg_rca24_fa291_and1;
  assign s_dadda_pg_rca24_and_20_14 = a[20] & b[14];
  assign s_dadda_pg_rca24_and_19_15 = a[19] & b[15];
  assign s_dadda_pg_rca24_and_18_16 = a[18] & b[16];
  assign s_dadda_pg_rca24_fa292_xor0 = s_dadda_pg_rca24_and_20_14 ^ s_dadda_pg_rca24_and_19_15;
  assign s_dadda_pg_rca24_fa292_and0 = s_dadda_pg_rca24_and_20_14 & s_dadda_pg_rca24_and_19_15;
  assign s_dadda_pg_rca24_fa292_xor1 = s_dadda_pg_rca24_fa292_xor0 ^ s_dadda_pg_rca24_and_18_16;
  assign s_dadda_pg_rca24_fa292_and1 = s_dadda_pg_rca24_fa292_xor0 & s_dadda_pg_rca24_and_18_16;
  assign s_dadda_pg_rca24_fa292_or0 = s_dadda_pg_rca24_fa292_and0 | s_dadda_pg_rca24_fa292_and1;
  assign s_dadda_pg_rca24_and_17_17 = a[17] & b[17];
  assign s_dadda_pg_rca24_and_16_18 = a[16] & b[18];
  assign s_dadda_pg_rca24_and_15_19 = a[15] & b[19];
  assign s_dadda_pg_rca24_fa293_xor0 = s_dadda_pg_rca24_and_17_17 ^ s_dadda_pg_rca24_and_16_18;
  assign s_dadda_pg_rca24_fa293_and0 = s_dadda_pg_rca24_and_17_17 & s_dadda_pg_rca24_and_16_18;
  assign s_dadda_pg_rca24_fa293_xor1 = s_dadda_pg_rca24_fa293_xor0 ^ s_dadda_pg_rca24_and_15_19;
  assign s_dadda_pg_rca24_fa293_and1 = s_dadda_pg_rca24_fa293_xor0 & s_dadda_pg_rca24_and_15_19;
  assign s_dadda_pg_rca24_fa293_or0 = s_dadda_pg_rca24_fa293_and0 | s_dadda_pg_rca24_fa293_and1;
  assign s_dadda_pg_rca24_and_14_20 = a[14] & b[20];
  assign s_dadda_pg_rca24_and_13_21 = a[13] & b[21];
  assign s_dadda_pg_rca24_and_12_22 = a[12] & b[22];
  assign s_dadda_pg_rca24_fa294_xor0 = s_dadda_pg_rca24_and_14_20 ^ s_dadda_pg_rca24_and_13_21;
  assign s_dadda_pg_rca24_fa294_and0 = s_dadda_pg_rca24_and_14_20 & s_dadda_pg_rca24_and_13_21;
  assign s_dadda_pg_rca24_fa294_xor1 = s_dadda_pg_rca24_fa294_xor0 ^ s_dadda_pg_rca24_and_12_22;
  assign s_dadda_pg_rca24_fa294_and1 = s_dadda_pg_rca24_fa294_xor0 & s_dadda_pg_rca24_and_12_22;
  assign s_dadda_pg_rca24_fa294_or0 = s_dadda_pg_rca24_fa294_and0 | s_dadda_pg_rca24_fa294_and1;
  assign s_dadda_pg_rca24_nand_11_23 = ~(a[11] & b[23]);
  assign s_dadda_pg_rca24_fa295_xor0 = s_dadda_pg_rca24_nand_11_23 ^ s_dadda_pg_rca24_fa288_xor1;
  assign s_dadda_pg_rca24_fa295_and0 = s_dadda_pg_rca24_nand_11_23 & s_dadda_pg_rca24_fa288_xor1;
  assign s_dadda_pg_rca24_fa295_xor1 = s_dadda_pg_rca24_fa295_xor0 ^ s_dadda_pg_rca24_fa289_xor1;
  assign s_dadda_pg_rca24_fa295_and1 = s_dadda_pg_rca24_fa295_xor0 & s_dadda_pg_rca24_fa289_xor1;
  assign s_dadda_pg_rca24_fa295_or0 = s_dadda_pg_rca24_fa295_and0 | s_dadda_pg_rca24_fa295_and1;
  assign s_dadda_pg_rca24_fa296_xor0 = s_dadda_pg_rca24_fa295_or0 ^ s_dadda_pg_rca24_fa294_or0;
  assign s_dadda_pg_rca24_fa296_and0 = s_dadda_pg_rca24_fa295_or0 & s_dadda_pg_rca24_fa294_or0;
  assign s_dadda_pg_rca24_fa296_xor1 = s_dadda_pg_rca24_fa296_xor0 ^ s_dadda_pg_rca24_fa293_or0;
  assign s_dadda_pg_rca24_fa296_and1 = s_dadda_pg_rca24_fa296_xor0 & s_dadda_pg_rca24_fa293_or0;
  assign s_dadda_pg_rca24_fa296_or0 = s_dadda_pg_rca24_fa296_and0 | s_dadda_pg_rca24_fa296_and1;
  assign s_dadda_pg_rca24_fa297_xor0 = s_dadda_pg_rca24_fa292_or0 ^ s_dadda_pg_rca24_fa291_or0;
  assign s_dadda_pg_rca24_fa297_and0 = s_dadda_pg_rca24_fa292_or0 & s_dadda_pg_rca24_fa291_or0;
  assign s_dadda_pg_rca24_fa297_xor1 = s_dadda_pg_rca24_fa297_xor0 ^ s_dadda_pg_rca24_fa290_or0;
  assign s_dadda_pg_rca24_fa297_and1 = s_dadda_pg_rca24_fa297_xor0 & s_dadda_pg_rca24_fa290_or0;
  assign s_dadda_pg_rca24_fa297_or0 = s_dadda_pg_rca24_fa297_and0 | s_dadda_pg_rca24_fa297_and1;
  assign s_dadda_pg_rca24_nand_23_12 = ~(a[23] & b[12]);
  assign s_dadda_pg_rca24_fa298_xor0 = s_dadda_pg_rca24_fa289_or0 ^ s_dadda_pg_rca24_fa288_or0;
  assign s_dadda_pg_rca24_fa298_and0 = s_dadda_pg_rca24_fa289_or0 & s_dadda_pg_rca24_fa288_or0;
  assign s_dadda_pg_rca24_fa298_xor1 = s_dadda_pg_rca24_fa298_xor0 ^ s_dadda_pg_rca24_nand_23_12;
  assign s_dadda_pg_rca24_fa298_and1 = s_dadda_pg_rca24_fa298_xor0 & s_dadda_pg_rca24_nand_23_12;
  assign s_dadda_pg_rca24_fa298_or0 = s_dadda_pg_rca24_fa298_and0 | s_dadda_pg_rca24_fa298_and1;
  assign s_dadda_pg_rca24_and_22_13 = a[22] & b[13];
  assign s_dadda_pg_rca24_and_21_14 = a[21] & b[14];
  assign s_dadda_pg_rca24_and_20_15 = a[20] & b[15];
  assign s_dadda_pg_rca24_fa299_xor0 = s_dadda_pg_rca24_and_22_13 ^ s_dadda_pg_rca24_and_21_14;
  assign s_dadda_pg_rca24_fa299_and0 = s_dadda_pg_rca24_and_22_13 & s_dadda_pg_rca24_and_21_14;
  assign s_dadda_pg_rca24_fa299_xor1 = s_dadda_pg_rca24_fa299_xor0 ^ s_dadda_pg_rca24_and_20_15;
  assign s_dadda_pg_rca24_fa299_and1 = s_dadda_pg_rca24_fa299_xor0 & s_dadda_pg_rca24_and_20_15;
  assign s_dadda_pg_rca24_fa299_or0 = s_dadda_pg_rca24_fa299_and0 | s_dadda_pg_rca24_fa299_and1;
  assign s_dadda_pg_rca24_and_19_16 = a[19] & b[16];
  assign s_dadda_pg_rca24_and_18_17 = a[18] & b[17];
  assign s_dadda_pg_rca24_and_17_18 = a[17] & b[18];
  assign s_dadda_pg_rca24_fa300_xor0 = s_dadda_pg_rca24_and_19_16 ^ s_dadda_pg_rca24_and_18_17;
  assign s_dadda_pg_rca24_fa300_and0 = s_dadda_pg_rca24_and_19_16 & s_dadda_pg_rca24_and_18_17;
  assign s_dadda_pg_rca24_fa300_xor1 = s_dadda_pg_rca24_fa300_xor0 ^ s_dadda_pg_rca24_and_17_18;
  assign s_dadda_pg_rca24_fa300_and1 = s_dadda_pg_rca24_fa300_xor0 & s_dadda_pg_rca24_and_17_18;
  assign s_dadda_pg_rca24_fa300_or0 = s_dadda_pg_rca24_fa300_and0 | s_dadda_pg_rca24_fa300_and1;
  assign s_dadda_pg_rca24_and_16_19 = a[16] & b[19];
  assign s_dadda_pg_rca24_and_15_20 = a[15] & b[20];
  assign s_dadda_pg_rca24_and_14_21 = a[14] & b[21];
  assign s_dadda_pg_rca24_fa301_xor0 = s_dadda_pg_rca24_and_16_19 ^ s_dadda_pg_rca24_and_15_20;
  assign s_dadda_pg_rca24_fa301_and0 = s_dadda_pg_rca24_and_16_19 & s_dadda_pg_rca24_and_15_20;
  assign s_dadda_pg_rca24_fa301_xor1 = s_dadda_pg_rca24_fa301_xor0 ^ s_dadda_pg_rca24_and_14_21;
  assign s_dadda_pg_rca24_fa301_and1 = s_dadda_pg_rca24_fa301_xor0 & s_dadda_pg_rca24_and_14_21;
  assign s_dadda_pg_rca24_fa301_or0 = s_dadda_pg_rca24_fa301_and0 | s_dadda_pg_rca24_fa301_and1;
  assign s_dadda_pg_rca24_and_13_22 = a[13] & b[22];
  assign s_dadda_pg_rca24_nand_12_23 = ~(a[12] & b[23]);
  assign s_dadda_pg_rca24_fa302_xor0 = s_dadda_pg_rca24_and_13_22 ^ s_dadda_pg_rca24_nand_12_23;
  assign s_dadda_pg_rca24_fa302_and0 = s_dadda_pg_rca24_and_13_22 & s_dadda_pg_rca24_nand_12_23;
  assign s_dadda_pg_rca24_fa302_xor1 = s_dadda_pg_rca24_fa302_xor0 ^ s_dadda_pg_rca24_fa296_xor1;
  assign s_dadda_pg_rca24_fa302_and1 = s_dadda_pg_rca24_fa302_xor0 & s_dadda_pg_rca24_fa296_xor1;
  assign s_dadda_pg_rca24_fa302_or0 = s_dadda_pg_rca24_fa302_and0 | s_dadda_pg_rca24_fa302_and1;
  assign s_dadda_pg_rca24_fa303_xor0 = s_dadda_pg_rca24_fa302_or0 ^ s_dadda_pg_rca24_fa301_or0;
  assign s_dadda_pg_rca24_fa303_and0 = s_dadda_pg_rca24_fa302_or0 & s_dadda_pg_rca24_fa301_or0;
  assign s_dadda_pg_rca24_fa303_xor1 = s_dadda_pg_rca24_fa303_xor0 ^ s_dadda_pg_rca24_fa300_or0;
  assign s_dadda_pg_rca24_fa303_and1 = s_dadda_pg_rca24_fa303_xor0 & s_dadda_pg_rca24_fa300_or0;
  assign s_dadda_pg_rca24_fa303_or0 = s_dadda_pg_rca24_fa303_and0 | s_dadda_pg_rca24_fa303_and1;
  assign s_dadda_pg_rca24_fa304_xor0 = s_dadda_pg_rca24_fa299_or0 ^ s_dadda_pg_rca24_fa298_or0;
  assign s_dadda_pg_rca24_fa304_and0 = s_dadda_pg_rca24_fa299_or0 & s_dadda_pg_rca24_fa298_or0;
  assign s_dadda_pg_rca24_fa304_xor1 = s_dadda_pg_rca24_fa304_xor0 ^ s_dadda_pg_rca24_fa297_or0;
  assign s_dadda_pg_rca24_fa304_and1 = s_dadda_pg_rca24_fa304_xor0 & s_dadda_pg_rca24_fa297_or0;
  assign s_dadda_pg_rca24_fa304_or0 = s_dadda_pg_rca24_fa304_and0 | s_dadda_pg_rca24_fa304_and1;
  assign s_dadda_pg_rca24_nand_23_13 = ~(a[23] & b[13]);
  assign s_dadda_pg_rca24_and_22_14 = a[22] & b[14];
  assign s_dadda_pg_rca24_fa305_xor0 = s_dadda_pg_rca24_fa296_or0 ^ s_dadda_pg_rca24_nand_23_13;
  assign s_dadda_pg_rca24_fa305_and0 = s_dadda_pg_rca24_fa296_or0 & s_dadda_pg_rca24_nand_23_13;
  assign s_dadda_pg_rca24_fa305_xor1 = s_dadda_pg_rca24_fa305_xor0 ^ s_dadda_pg_rca24_and_22_14;
  assign s_dadda_pg_rca24_fa305_and1 = s_dadda_pg_rca24_fa305_xor0 & s_dadda_pg_rca24_and_22_14;
  assign s_dadda_pg_rca24_fa305_or0 = s_dadda_pg_rca24_fa305_and0 | s_dadda_pg_rca24_fa305_and1;
  assign s_dadda_pg_rca24_and_21_15 = a[21] & b[15];
  assign s_dadda_pg_rca24_and_20_16 = a[20] & b[16];
  assign s_dadda_pg_rca24_and_19_17 = a[19] & b[17];
  assign s_dadda_pg_rca24_fa306_xor0 = s_dadda_pg_rca24_and_21_15 ^ s_dadda_pg_rca24_and_20_16;
  assign s_dadda_pg_rca24_fa306_and0 = s_dadda_pg_rca24_and_21_15 & s_dadda_pg_rca24_and_20_16;
  assign s_dadda_pg_rca24_fa306_xor1 = s_dadda_pg_rca24_fa306_xor0 ^ s_dadda_pg_rca24_and_19_17;
  assign s_dadda_pg_rca24_fa306_and1 = s_dadda_pg_rca24_fa306_xor0 & s_dadda_pg_rca24_and_19_17;
  assign s_dadda_pg_rca24_fa306_or0 = s_dadda_pg_rca24_fa306_and0 | s_dadda_pg_rca24_fa306_and1;
  assign s_dadda_pg_rca24_and_18_18 = a[18] & b[18];
  assign s_dadda_pg_rca24_and_17_19 = a[17] & b[19];
  assign s_dadda_pg_rca24_and_16_20 = a[16] & b[20];
  assign s_dadda_pg_rca24_fa307_xor0 = s_dadda_pg_rca24_and_18_18 ^ s_dadda_pg_rca24_and_17_19;
  assign s_dadda_pg_rca24_fa307_and0 = s_dadda_pg_rca24_and_18_18 & s_dadda_pg_rca24_and_17_19;
  assign s_dadda_pg_rca24_fa307_xor1 = s_dadda_pg_rca24_fa307_xor0 ^ s_dadda_pg_rca24_and_16_20;
  assign s_dadda_pg_rca24_fa307_and1 = s_dadda_pg_rca24_fa307_xor0 & s_dadda_pg_rca24_and_16_20;
  assign s_dadda_pg_rca24_fa307_or0 = s_dadda_pg_rca24_fa307_and0 | s_dadda_pg_rca24_fa307_and1;
  assign s_dadda_pg_rca24_and_15_21 = a[15] & b[21];
  assign s_dadda_pg_rca24_and_14_22 = a[14] & b[22];
  assign s_dadda_pg_rca24_nand_13_23 = ~(a[13] & b[23]);
  assign s_dadda_pg_rca24_fa308_xor0 = s_dadda_pg_rca24_and_15_21 ^ s_dadda_pg_rca24_and_14_22;
  assign s_dadda_pg_rca24_fa308_and0 = s_dadda_pg_rca24_and_15_21 & s_dadda_pg_rca24_and_14_22;
  assign s_dadda_pg_rca24_fa308_xor1 = s_dadda_pg_rca24_fa308_xor0 ^ s_dadda_pg_rca24_nand_13_23;
  assign s_dadda_pg_rca24_fa308_and1 = s_dadda_pg_rca24_fa308_xor0 & s_dadda_pg_rca24_nand_13_23;
  assign s_dadda_pg_rca24_fa308_or0 = s_dadda_pg_rca24_fa308_and0 | s_dadda_pg_rca24_fa308_and1;
  assign s_dadda_pg_rca24_fa309_xor0 = s_dadda_pg_rca24_fa308_or0 ^ s_dadda_pg_rca24_fa307_or0;
  assign s_dadda_pg_rca24_fa309_and0 = s_dadda_pg_rca24_fa308_or0 & s_dadda_pg_rca24_fa307_or0;
  assign s_dadda_pg_rca24_fa309_xor1 = s_dadda_pg_rca24_fa309_xor0 ^ s_dadda_pg_rca24_fa306_or0;
  assign s_dadda_pg_rca24_fa309_and1 = s_dadda_pg_rca24_fa309_xor0 & s_dadda_pg_rca24_fa306_or0;
  assign s_dadda_pg_rca24_fa309_or0 = s_dadda_pg_rca24_fa309_and0 | s_dadda_pg_rca24_fa309_and1;
  assign s_dadda_pg_rca24_fa310_xor0 = s_dadda_pg_rca24_fa305_or0 ^ s_dadda_pg_rca24_fa304_or0;
  assign s_dadda_pg_rca24_fa310_and0 = s_dadda_pg_rca24_fa305_or0 & s_dadda_pg_rca24_fa304_or0;
  assign s_dadda_pg_rca24_fa310_xor1 = s_dadda_pg_rca24_fa310_xor0 ^ s_dadda_pg_rca24_fa303_or0;
  assign s_dadda_pg_rca24_fa310_and1 = s_dadda_pg_rca24_fa310_xor0 & s_dadda_pg_rca24_fa303_or0;
  assign s_dadda_pg_rca24_fa310_or0 = s_dadda_pg_rca24_fa310_and0 | s_dadda_pg_rca24_fa310_and1;
  assign s_dadda_pg_rca24_nand_23_14 = ~(a[23] & b[14]);
  assign s_dadda_pg_rca24_and_22_15 = a[22] & b[15];
  assign s_dadda_pg_rca24_and_21_16 = a[21] & b[16];
  assign s_dadda_pg_rca24_fa311_xor0 = s_dadda_pg_rca24_nand_23_14 ^ s_dadda_pg_rca24_and_22_15;
  assign s_dadda_pg_rca24_fa311_and0 = s_dadda_pg_rca24_nand_23_14 & s_dadda_pg_rca24_and_22_15;
  assign s_dadda_pg_rca24_fa311_xor1 = s_dadda_pg_rca24_fa311_xor0 ^ s_dadda_pg_rca24_and_21_16;
  assign s_dadda_pg_rca24_fa311_and1 = s_dadda_pg_rca24_fa311_xor0 & s_dadda_pg_rca24_and_21_16;
  assign s_dadda_pg_rca24_fa311_or0 = s_dadda_pg_rca24_fa311_and0 | s_dadda_pg_rca24_fa311_and1;
  assign s_dadda_pg_rca24_and_20_17 = a[20] & b[17];
  assign s_dadda_pg_rca24_and_19_18 = a[19] & b[18];
  assign s_dadda_pg_rca24_and_18_19 = a[18] & b[19];
  assign s_dadda_pg_rca24_fa312_xor0 = s_dadda_pg_rca24_and_20_17 ^ s_dadda_pg_rca24_and_19_18;
  assign s_dadda_pg_rca24_fa312_and0 = s_dadda_pg_rca24_and_20_17 & s_dadda_pg_rca24_and_19_18;
  assign s_dadda_pg_rca24_fa312_xor1 = s_dadda_pg_rca24_fa312_xor0 ^ s_dadda_pg_rca24_and_18_19;
  assign s_dadda_pg_rca24_fa312_and1 = s_dadda_pg_rca24_fa312_xor0 & s_dadda_pg_rca24_and_18_19;
  assign s_dadda_pg_rca24_fa312_or0 = s_dadda_pg_rca24_fa312_and0 | s_dadda_pg_rca24_fa312_and1;
  assign s_dadda_pg_rca24_and_17_20 = a[17] & b[20];
  assign s_dadda_pg_rca24_and_16_21 = a[16] & b[21];
  assign s_dadda_pg_rca24_and_15_22 = a[15] & b[22];
  assign s_dadda_pg_rca24_fa313_xor0 = s_dadda_pg_rca24_and_17_20 ^ s_dadda_pg_rca24_and_16_21;
  assign s_dadda_pg_rca24_fa313_and0 = s_dadda_pg_rca24_and_17_20 & s_dadda_pg_rca24_and_16_21;
  assign s_dadda_pg_rca24_fa313_xor1 = s_dadda_pg_rca24_fa313_xor0 ^ s_dadda_pg_rca24_and_15_22;
  assign s_dadda_pg_rca24_fa313_and1 = s_dadda_pg_rca24_fa313_xor0 & s_dadda_pg_rca24_and_15_22;
  assign s_dadda_pg_rca24_fa313_or0 = s_dadda_pg_rca24_fa313_and0 | s_dadda_pg_rca24_fa313_and1;
  assign s_dadda_pg_rca24_fa314_xor0 = s_dadda_pg_rca24_fa313_or0 ^ s_dadda_pg_rca24_fa312_or0;
  assign s_dadda_pg_rca24_fa314_and0 = s_dadda_pg_rca24_fa313_or0 & s_dadda_pg_rca24_fa312_or0;
  assign s_dadda_pg_rca24_fa314_xor1 = s_dadda_pg_rca24_fa314_xor0 ^ s_dadda_pg_rca24_fa311_or0;
  assign s_dadda_pg_rca24_fa314_and1 = s_dadda_pg_rca24_fa314_xor0 & s_dadda_pg_rca24_fa311_or0;
  assign s_dadda_pg_rca24_fa314_or0 = s_dadda_pg_rca24_fa314_and0 | s_dadda_pg_rca24_fa314_and1;
  assign s_dadda_pg_rca24_nand_23_15 = ~(a[23] & b[15]);
  assign s_dadda_pg_rca24_fa315_xor0 = s_dadda_pg_rca24_fa310_or0 ^ s_dadda_pg_rca24_fa309_or0;
  assign s_dadda_pg_rca24_fa315_and0 = s_dadda_pg_rca24_fa310_or0 & s_dadda_pg_rca24_fa309_or0;
  assign s_dadda_pg_rca24_fa315_xor1 = s_dadda_pg_rca24_fa315_xor0 ^ s_dadda_pg_rca24_nand_23_15;
  assign s_dadda_pg_rca24_fa315_and1 = s_dadda_pg_rca24_fa315_xor0 & s_dadda_pg_rca24_nand_23_15;
  assign s_dadda_pg_rca24_fa315_or0 = s_dadda_pg_rca24_fa315_and0 | s_dadda_pg_rca24_fa315_and1;
  assign s_dadda_pg_rca24_and_22_16 = a[22] & b[16];
  assign s_dadda_pg_rca24_and_21_17 = a[21] & b[17];
  assign s_dadda_pg_rca24_and_20_18 = a[20] & b[18];
  assign s_dadda_pg_rca24_fa316_xor0 = s_dadda_pg_rca24_and_22_16 ^ s_dadda_pg_rca24_and_21_17;
  assign s_dadda_pg_rca24_fa316_and0 = s_dadda_pg_rca24_and_22_16 & s_dadda_pg_rca24_and_21_17;
  assign s_dadda_pg_rca24_fa316_xor1 = s_dadda_pg_rca24_fa316_xor0 ^ s_dadda_pg_rca24_and_20_18;
  assign s_dadda_pg_rca24_fa316_and1 = s_dadda_pg_rca24_fa316_xor0 & s_dadda_pg_rca24_and_20_18;
  assign s_dadda_pg_rca24_fa316_or0 = s_dadda_pg_rca24_fa316_and0 | s_dadda_pg_rca24_fa316_and1;
  assign s_dadda_pg_rca24_and_19_19 = a[19] & b[19];
  assign s_dadda_pg_rca24_and_18_20 = a[18] & b[20];
  assign s_dadda_pg_rca24_and_17_21 = a[17] & b[21];
  assign s_dadda_pg_rca24_fa317_xor0 = s_dadda_pg_rca24_and_19_19 ^ s_dadda_pg_rca24_and_18_20;
  assign s_dadda_pg_rca24_fa317_and0 = s_dadda_pg_rca24_and_19_19 & s_dadda_pg_rca24_and_18_20;
  assign s_dadda_pg_rca24_fa317_xor1 = s_dadda_pg_rca24_fa317_xor0 ^ s_dadda_pg_rca24_and_17_21;
  assign s_dadda_pg_rca24_fa317_and1 = s_dadda_pg_rca24_fa317_xor0 & s_dadda_pg_rca24_and_17_21;
  assign s_dadda_pg_rca24_fa317_or0 = s_dadda_pg_rca24_fa317_and0 | s_dadda_pg_rca24_fa317_and1;
  assign s_dadda_pg_rca24_fa318_xor0 = s_dadda_pg_rca24_fa317_or0 ^ s_dadda_pg_rca24_fa316_or0;
  assign s_dadda_pg_rca24_fa318_and0 = s_dadda_pg_rca24_fa317_or0 & s_dadda_pg_rca24_fa316_or0;
  assign s_dadda_pg_rca24_fa318_xor1 = s_dadda_pg_rca24_fa318_xor0 ^ s_dadda_pg_rca24_fa315_or0;
  assign s_dadda_pg_rca24_fa318_and1 = s_dadda_pg_rca24_fa318_xor0 & s_dadda_pg_rca24_fa315_or0;
  assign s_dadda_pg_rca24_fa318_or0 = s_dadda_pg_rca24_fa318_and0 | s_dadda_pg_rca24_fa318_and1;
  assign s_dadda_pg_rca24_nand_23_16 = ~(a[23] & b[16]);
  assign s_dadda_pg_rca24_and_22_17 = a[22] & b[17];
  assign s_dadda_pg_rca24_fa319_xor0 = s_dadda_pg_rca24_fa314_or0 ^ s_dadda_pg_rca24_nand_23_16;
  assign s_dadda_pg_rca24_fa319_and0 = s_dadda_pg_rca24_fa314_or0 & s_dadda_pg_rca24_nand_23_16;
  assign s_dadda_pg_rca24_fa319_xor1 = s_dadda_pg_rca24_fa319_xor0 ^ s_dadda_pg_rca24_and_22_17;
  assign s_dadda_pg_rca24_fa319_and1 = s_dadda_pg_rca24_fa319_xor0 & s_dadda_pg_rca24_and_22_17;
  assign s_dadda_pg_rca24_fa319_or0 = s_dadda_pg_rca24_fa319_and0 | s_dadda_pg_rca24_fa319_and1;
  assign s_dadda_pg_rca24_and_21_18 = a[21] & b[18];
  assign s_dadda_pg_rca24_and_20_19 = a[20] & b[19];
  assign s_dadda_pg_rca24_and_19_20 = a[19] & b[20];
  assign s_dadda_pg_rca24_fa320_xor0 = s_dadda_pg_rca24_and_21_18 ^ s_dadda_pg_rca24_and_20_19;
  assign s_dadda_pg_rca24_fa320_and0 = s_dadda_pg_rca24_and_21_18 & s_dadda_pg_rca24_and_20_19;
  assign s_dadda_pg_rca24_fa320_xor1 = s_dadda_pg_rca24_fa320_xor0 ^ s_dadda_pg_rca24_and_19_20;
  assign s_dadda_pg_rca24_fa320_and1 = s_dadda_pg_rca24_fa320_xor0 & s_dadda_pg_rca24_and_19_20;
  assign s_dadda_pg_rca24_fa320_or0 = s_dadda_pg_rca24_fa320_and0 | s_dadda_pg_rca24_fa320_and1;
  assign s_dadda_pg_rca24_fa321_xor0 = s_dadda_pg_rca24_fa320_or0 ^ s_dadda_pg_rca24_fa319_or0;
  assign s_dadda_pg_rca24_fa321_and0 = s_dadda_pg_rca24_fa320_or0 & s_dadda_pg_rca24_fa319_or0;
  assign s_dadda_pg_rca24_fa321_xor1 = s_dadda_pg_rca24_fa321_xor0 ^ s_dadda_pg_rca24_fa318_or0;
  assign s_dadda_pg_rca24_fa321_and1 = s_dadda_pg_rca24_fa321_xor0 & s_dadda_pg_rca24_fa318_or0;
  assign s_dadda_pg_rca24_fa321_or0 = s_dadda_pg_rca24_fa321_and0 | s_dadda_pg_rca24_fa321_and1;
  assign s_dadda_pg_rca24_nand_23_17 = ~(a[23] & b[17]);
  assign s_dadda_pg_rca24_and_22_18 = a[22] & b[18];
  assign s_dadda_pg_rca24_and_21_19 = a[21] & b[19];
  assign s_dadda_pg_rca24_fa322_xor0 = s_dadda_pg_rca24_nand_23_17 ^ s_dadda_pg_rca24_and_22_18;
  assign s_dadda_pg_rca24_fa322_and0 = s_dadda_pg_rca24_nand_23_17 & s_dadda_pg_rca24_and_22_18;
  assign s_dadda_pg_rca24_fa322_xor1 = s_dadda_pg_rca24_fa322_xor0 ^ s_dadda_pg_rca24_and_21_19;
  assign s_dadda_pg_rca24_fa322_and1 = s_dadda_pg_rca24_fa322_xor0 & s_dadda_pg_rca24_and_21_19;
  assign s_dadda_pg_rca24_fa322_or0 = s_dadda_pg_rca24_fa322_and0 | s_dadda_pg_rca24_fa322_and1;
  assign s_dadda_pg_rca24_nand_23_18 = ~(a[23] & b[18]);
  assign s_dadda_pg_rca24_fa323_xor0 = s_dadda_pg_rca24_fa322_or0 ^ s_dadda_pg_rca24_fa321_or0;
  assign s_dadda_pg_rca24_fa323_and0 = s_dadda_pg_rca24_fa322_or0 & s_dadda_pg_rca24_fa321_or0;
  assign s_dadda_pg_rca24_fa323_xor1 = s_dadda_pg_rca24_fa323_xor0 ^ s_dadda_pg_rca24_nand_23_18;
  assign s_dadda_pg_rca24_fa323_and1 = s_dadda_pg_rca24_fa323_xor0 & s_dadda_pg_rca24_nand_23_18;
  assign s_dadda_pg_rca24_fa323_or0 = s_dadda_pg_rca24_fa323_and0 | s_dadda_pg_rca24_fa323_and1;
  assign s_dadda_pg_rca24_and_4_0 = a[4] & b[0];
  assign s_dadda_pg_rca24_and_3_1 = a[3] & b[1];
  assign s_dadda_pg_rca24_ha18_xor0 = s_dadda_pg_rca24_and_4_0 ^ s_dadda_pg_rca24_and_3_1;
  assign s_dadda_pg_rca24_ha18_and0 = s_dadda_pg_rca24_and_4_0 & s_dadda_pg_rca24_and_3_1;
  assign s_dadda_pg_rca24_and_5_0 = a[5] & b[0];
  assign s_dadda_pg_rca24_and_4_1 = a[4] & b[1];
  assign s_dadda_pg_rca24_fa324_xor0 = s_dadda_pg_rca24_ha18_and0 ^ s_dadda_pg_rca24_and_5_0;
  assign s_dadda_pg_rca24_fa324_and0 = s_dadda_pg_rca24_ha18_and0 & s_dadda_pg_rca24_and_5_0;
  assign s_dadda_pg_rca24_fa324_xor1 = s_dadda_pg_rca24_fa324_xor0 ^ s_dadda_pg_rca24_and_4_1;
  assign s_dadda_pg_rca24_fa324_and1 = s_dadda_pg_rca24_fa324_xor0 & s_dadda_pg_rca24_and_4_1;
  assign s_dadda_pg_rca24_fa324_or0 = s_dadda_pg_rca24_fa324_and0 | s_dadda_pg_rca24_fa324_and1;
  assign s_dadda_pg_rca24_and_3_2 = a[3] & b[2];
  assign s_dadda_pg_rca24_and_2_3 = a[2] & b[3];
  assign s_dadda_pg_rca24_ha19_xor0 = s_dadda_pg_rca24_and_3_2 ^ s_dadda_pg_rca24_and_2_3;
  assign s_dadda_pg_rca24_ha19_and0 = s_dadda_pg_rca24_and_3_2 & s_dadda_pg_rca24_and_2_3;
  assign s_dadda_pg_rca24_and_4_2 = a[4] & b[2];
  assign s_dadda_pg_rca24_fa325_xor0 = s_dadda_pg_rca24_ha19_and0 ^ s_dadda_pg_rca24_fa324_or0;
  assign s_dadda_pg_rca24_fa325_and0 = s_dadda_pg_rca24_ha19_and0 & s_dadda_pg_rca24_fa324_or0;
  assign s_dadda_pg_rca24_fa325_xor1 = s_dadda_pg_rca24_fa325_xor0 ^ s_dadda_pg_rca24_and_4_2;
  assign s_dadda_pg_rca24_fa325_and1 = s_dadda_pg_rca24_fa325_xor0 & s_dadda_pg_rca24_and_4_2;
  assign s_dadda_pg_rca24_fa325_or0 = s_dadda_pg_rca24_fa325_and0 | s_dadda_pg_rca24_fa325_and1;
  assign s_dadda_pg_rca24_and_3_3 = a[3] & b[3];
  assign s_dadda_pg_rca24_and_2_4 = a[2] & b[4];
  assign s_dadda_pg_rca24_and_1_5 = a[1] & b[5];
  assign s_dadda_pg_rca24_fa326_xor0 = s_dadda_pg_rca24_and_3_3 ^ s_dadda_pg_rca24_and_2_4;
  assign s_dadda_pg_rca24_fa326_and0 = s_dadda_pg_rca24_and_3_3 & s_dadda_pg_rca24_and_2_4;
  assign s_dadda_pg_rca24_fa326_xor1 = s_dadda_pg_rca24_fa326_xor0 ^ s_dadda_pg_rca24_and_1_5;
  assign s_dadda_pg_rca24_fa326_and1 = s_dadda_pg_rca24_fa326_xor0 & s_dadda_pg_rca24_and_1_5;
  assign s_dadda_pg_rca24_fa326_or0 = s_dadda_pg_rca24_fa326_and0 | s_dadda_pg_rca24_fa326_and1;
  assign s_dadda_pg_rca24_and_3_4 = a[3] & b[4];
  assign s_dadda_pg_rca24_fa327_xor0 = s_dadda_pg_rca24_fa326_or0 ^ s_dadda_pg_rca24_fa325_or0;
  assign s_dadda_pg_rca24_fa327_and0 = s_dadda_pg_rca24_fa326_or0 & s_dadda_pg_rca24_fa325_or0;
  assign s_dadda_pg_rca24_fa327_xor1 = s_dadda_pg_rca24_fa327_xor0 ^ s_dadda_pg_rca24_and_3_4;
  assign s_dadda_pg_rca24_fa327_and1 = s_dadda_pg_rca24_fa327_xor0 & s_dadda_pg_rca24_and_3_4;
  assign s_dadda_pg_rca24_fa327_or0 = s_dadda_pg_rca24_fa327_and0 | s_dadda_pg_rca24_fa327_and1;
  assign s_dadda_pg_rca24_and_2_5 = a[2] & b[5];
  assign s_dadda_pg_rca24_and_1_6 = a[1] & b[6];
  assign s_dadda_pg_rca24_and_0_7 = a[0] & b[7];
  assign s_dadda_pg_rca24_fa328_xor0 = s_dadda_pg_rca24_and_2_5 ^ s_dadda_pg_rca24_and_1_6;
  assign s_dadda_pg_rca24_fa328_and0 = s_dadda_pg_rca24_and_2_5 & s_dadda_pg_rca24_and_1_6;
  assign s_dadda_pg_rca24_fa328_xor1 = s_dadda_pg_rca24_fa328_xor0 ^ s_dadda_pg_rca24_and_0_7;
  assign s_dadda_pg_rca24_fa328_and1 = s_dadda_pg_rca24_fa328_xor0 & s_dadda_pg_rca24_and_0_7;
  assign s_dadda_pg_rca24_fa328_or0 = s_dadda_pg_rca24_fa328_and0 | s_dadda_pg_rca24_fa328_and1;
  assign s_dadda_pg_rca24_and_2_6 = a[2] & b[6];
  assign s_dadda_pg_rca24_fa329_xor0 = s_dadda_pg_rca24_fa328_or0 ^ s_dadda_pg_rca24_fa327_or0;
  assign s_dadda_pg_rca24_fa329_and0 = s_dadda_pg_rca24_fa328_or0 & s_dadda_pg_rca24_fa327_or0;
  assign s_dadda_pg_rca24_fa329_xor1 = s_dadda_pg_rca24_fa329_xor0 ^ s_dadda_pg_rca24_and_2_6;
  assign s_dadda_pg_rca24_fa329_and1 = s_dadda_pg_rca24_fa329_xor0 & s_dadda_pg_rca24_and_2_6;
  assign s_dadda_pg_rca24_fa329_or0 = s_dadda_pg_rca24_fa329_and0 | s_dadda_pg_rca24_fa329_and1;
  assign s_dadda_pg_rca24_and_1_7 = a[1] & b[7];
  assign s_dadda_pg_rca24_and_0_8 = a[0] & b[8];
  assign s_dadda_pg_rca24_fa330_xor0 = s_dadda_pg_rca24_and_1_7 ^ s_dadda_pg_rca24_and_0_8;
  assign s_dadda_pg_rca24_fa330_and0 = s_dadda_pg_rca24_and_1_7 & s_dadda_pg_rca24_and_0_8;
  assign s_dadda_pg_rca24_fa330_xor1 = s_dadda_pg_rca24_fa330_xor0 ^ s_dadda_pg_rca24_fa26_xor1;
  assign s_dadda_pg_rca24_fa330_and1 = s_dadda_pg_rca24_fa330_xor0 & s_dadda_pg_rca24_fa26_xor1;
  assign s_dadda_pg_rca24_fa330_or0 = s_dadda_pg_rca24_fa330_and0 | s_dadda_pg_rca24_fa330_and1;
  assign s_dadda_pg_rca24_and_1_8 = a[1] & b[8];
  assign s_dadda_pg_rca24_fa331_xor0 = s_dadda_pg_rca24_fa330_or0 ^ s_dadda_pg_rca24_fa329_or0;
  assign s_dadda_pg_rca24_fa331_and0 = s_dadda_pg_rca24_fa330_or0 & s_dadda_pg_rca24_fa329_or0;
  assign s_dadda_pg_rca24_fa331_xor1 = s_dadda_pg_rca24_fa331_xor0 ^ s_dadda_pg_rca24_and_1_8;
  assign s_dadda_pg_rca24_fa331_and1 = s_dadda_pg_rca24_fa331_xor0 & s_dadda_pg_rca24_and_1_8;
  assign s_dadda_pg_rca24_fa331_or0 = s_dadda_pg_rca24_fa331_and0 | s_dadda_pg_rca24_fa331_and1;
  assign s_dadda_pg_rca24_and_0_9 = a[0] & b[9];
  assign s_dadda_pg_rca24_fa332_xor0 = s_dadda_pg_rca24_and_0_9 ^ s_dadda_pg_rca24_fa28_xor1;
  assign s_dadda_pg_rca24_fa332_and0 = s_dadda_pg_rca24_and_0_9 & s_dadda_pg_rca24_fa28_xor1;
  assign s_dadda_pg_rca24_fa332_xor1 = s_dadda_pg_rca24_fa332_xor0 ^ s_dadda_pg_rca24_fa29_xor1;
  assign s_dadda_pg_rca24_fa332_and1 = s_dadda_pg_rca24_fa332_xor0 & s_dadda_pg_rca24_fa29_xor1;
  assign s_dadda_pg_rca24_fa332_or0 = s_dadda_pg_rca24_fa332_and0 | s_dadda_pg_rca24_fa332_and1;
  assign s_dadda_pg_rca24_and_0_10 = a[0] & b[10];
  assign s_dadda_pg_rca24_fa333_xor0 = s_dadda_pg_rca24_fa332_or0 ^ s_dadda_pg_rca24_fa331_or0;
  assign s_dadda_pg_rca24_fa333_and0 = s_dadda_pg_rca24_fa332_or0 & s_dadda_pg_rca24_fa331_or0;
  assign s_dadda_pg_rca24_fa333_xor1 = s_dadda_pg_rca24_fa333_xor0 ^ s_dadda_pg_rca24_and_0_10;
  assign s_dadda_pg_rca24_fa333_and1 = s_dadda_pg_rca24_fa333_xor0 & s_dadda_pg_rca24_and_0_10;
  assign s_dadda_pg_rca24_fa333_or0 = s_dadda_pg_rca24_fa333_and0 | s_dadda_pg_rca24_fa333_and1;
  assign s_dadda_pg_rca24_fa334_xor0 = s_dadda_pg_rca24_fa31_xor1 ^ s_dadda_pg_rca24_fa32_xor1;
  assign s_dadda_pg_rca24_fa334_and0 = s_dadda_pg_rca24_fa31_xor1 & s_dadda_pg_rca24_fa32_xor1;
  assign s_dadda_pg_rca24_fa334_xor1 = s_dadda_pg_rca24_fa334_xor0 ^ s_dadda_pg_rca24_fa33_xor1;
  assign s_dadda_pg_rca24_fa334_and1 = s_dadda_pg_rca24_fa334_xor0 & s_dadda_pg_rca24_fa33_xor1;
  assign s_dadda_pg_rca24_fa334_or0 = s_dadda_pg_rca24_fa334_and0 | s_dadda_pg_rca24_fa334_and1;
  assign s_dadda_pg_rca24_fa335_xor0 = s_dadda_pg_rca24_fa334_or0 ^ s_dadda_pg_rca24_fa333_or0;
  assign s_dadda_pg_rca24_fa335_and0 = s_dadda_pg_rca24_fa334_or0 & s_dadda_pg_rca24_fa333_or0;
  assign s_dadda_pg_rca24_fa335_xor1 = s_dadda_pg_rca24_fa335_xor0 ^ s_dadda_pg_rca24_fa35_xor1;
  assign s_dadda_pg_rca24_fa335_and1 = s_dadda_pg_rca24_fa335_xor0 & s_dadda_pg_rca24_fa35_xor1;
  assign s_dadda_pg_rca24_fa335_or0 = s_dadda_pg_rca24_fa335_and0 | s_dadda_pg_rca24_fa335_and1;
  assign s_dadda_pg_rca24_fa336_xor0 = s_dadda_pg_rca24_fa36_xor1 ^ s_dadda_pg_rca24_fa37_xor1;
  assign s_dadda_pg_rca24_fa336_and0 = s_dadda_pg_rca24_fa36_xor1 & s_dadda_pg_rca24_fa37_xor1;
  assign s_dadda_pg_rca24_fa336_xor1 = s_dadda_pg_rca24_fa336_xor0 ^ s_dadda_pg_rca24_fa38_xor1;
  assign s_dadda_pg_rca24_fa336_and1 = s_dadda_pg_rca24_fa336_xor0 & s_dadda_pg_rca24_fa38_xor1;
  assign s_dadda_pg_rca24_fa336_or0 = s_dadda_pg_rca24_fa336_and0 | s_dadda_pg_rca24_fa336_and1;
  assign s_dadda_pg_rca24_fa337_xor0 = s_dadda_pg_rca24_fa336_or0 ^ s_dadda_pg_rca24_fa335_or0;
  assign s_dadda_pg_rca24_fa337_and0 = s_dadda_pg_rca24_fa336_or0 & s_dadda_pg_rca24_fa335_or0;
  assign s_dadda_pg_rca24_fa337_xor1 = s_dadda_pg_rca24_fa337_xor0 ^ s_dadda_pg_rca24_fa41_xor1;
  assign s_dadda_pg_rca24_fa337_and1 = s_dadda_pg_rca24_fa337_xor0 & s_dadda_pg_rca24_fa41_xor1;
  assign s_dadda_pg_rca24_fa337_or0 = s_dadda_pg_rca24_fa337_and0 | s_dadda_pg_rca24_fa337_and1;
  assign s_dadda_pg_rca24_fa338_xor0 = s_dadda_pg_rca24_fa42_xor1 ^ s_dadda_pg_rca24_fa43_xor1;
  assign s_dadda_pg_rca24_fa338_and0 = s_dadda_pg_rca24_fa42_xor1 & s_dadda_pg_rca24_fa43_xor1;
  assign s_dadda_pg_rca24_fa338_xor1 = s_dadda_pg_rca24_fa338_xor0 ^ s_dadda_pg_rca24_fa44_xor1;
  assign s_dadda_pg_rca24_fa338_and1 = s_dadda_pg_rca24_fa338_xor0 & s_dadda_pg_rca24_fa44_xor1;
  assign s_dadda_pg_rca24_fa338_or0 = s_dadda_pg_rca24_fa338_and0 | s_dadda_pg_rca24_fa338_and1;
  assign s_dadda_pg_rca24_fa339_xor0 = s_dadda_pg_rca24_fa338_or0 ^ s_dadda_pg_rca24_fa337_or0;
  assign s_dadda_pg_rca24_fa339_and0 = s_dadda_pg_rca24_fa338_or0 & s_dadda_pg_rca24_fa337_or0;
  assign s_dadda_pg_rca24_fa339_xor1 = s_dadda_pg_rca24_fa339_xor0 ^ s_dadda_pg_rca24_fa48_xor1;
  assign s_dadda_pg_rca24_fa339_and1 = s_dadda_pg_rca24_fa339_xor0 & s_dadda_pg_rca24_fa48_xor1;
  assign s_dadda_pg_rca24_fa339_or0 = s_dadda_pg_rca24_fa339_and0 | s_dadda_pg_rca24_fa339_and1;
  assign s_dadda_pg_rca24_fa340_xor0 = s_dadda_pg_rca24_fa49_xor1 ^ s_dadda_pg_rca24_fa50_xor1;
  assign s_dadda_pg_rca24_fa340_and0 = s_dadda_pg_rca24_fa49_xor1 & s_dadda_pg_rca24_fa50_xor1;
  assign s_dadda_pg_rca24_fa340_xor1 = s_dadda_pg_rca24_fa340_xor0 ^ s_dadda_pg_rca24_fa51_xor1;
  assign s_dadda_pg_rca24_fa340_and1 = s_dadda_pg_rca24_fa340_xor0 & s_dadda_pg_rca24_fa51_xor1;
  assign s_dadda_pg_rca24_fa340_or0 = s_dadda_pg_rca24_fa340_and0 | s_dadda_pg_rca24_fa340_and1;
  assign s_dadda_pg_rca24_fa341_xor0 = s_dadda_pg_rca24_fa340_or0 ^ s_dadda_pg_rca24_fa339_or0;
  assign s_dadda_pg_rca24_fa341_and0 = s_dadda_pg_rca24_fa340_or0 & s_dadda_pg_rca24_fa339_or0;
  assign s_dadda_pg_rca24_fa341_xor1 = s_dadda_pg_rca24_fa341_xor0 ^ s_dadda_pg_rca24_fa56_xor1;
  assign s_dadda_pg_rca24_fa341_and1 = s_dadda_pg_rca24_fa341_xor0 & s_dadda_pg_rca24_fa56_xor1;
  assign s_dadda_pg_rca24_fa341_or0 = s_dadda_pg_rca24_fa341_and0 | s_dadda_pg_rca24_fa341_and1;
  assign s_dadda_pg_rca24_fa342_xor0 = s_dadda_pg_rca24_fa57_xor1 ^ s_dadda_pg_rca24_fa58_xor1;
  assign s_dadda_pg_rca24_fa342_and0 = s_dadda_pg_rca24_fa57_xor1 & s_dadda_pg_rca24_fa58_xor1;
  assign s_dadda_pg_rca24_fa342_xor1 = s_dadda_pg_rca24_fa342_xor0 ^ s_dadda_pg_rca24_fa59_xor1;
  assign s_dadda_pg_rca24_fa342_and1 = s_dadda_pg_rca24_fa342_xor0 & s_dadda_pg_rca24_fa59_xor1;
  assign s_dadda_pg_rca24_fa342_or0 = s_dadda_pg_rca24_fa342_and0 | s_dadda_pg_rca24_fa342_and1;
  assign s_dadda_pg_rca24_fa343_xor0 = s_dadda_pg_rca24_fa342_or0 ^ s_dadda_pg_rca24_fa341_or0;
  assign s_dadda_pg_rca24_fa343_and0 = s_dadda_pg_rca24_fa342_or0 & s_dadda_pg_rca24_fa341_or0;
  assign s_dadda_pg_rca24_fa343_xor1 = s_dadda_pg_rca24_fa343_xor0 ^ s_dadda_pg_rca24_fa65_xor1;
  assign s_dadda_pg_rca24_fa343_and1 = s_dadda_pg_rca24_fa343_xor0 & s_dadda_pg_rca24_fa65_xor1;
  assign s_dadda_pg_rca24_fa343_or0 = s_dadda_pg_rca24_fa343_and0 | s_dadda_pg_rca24_fa343_and1;
  assign s_dadda_pg_rca24_fa344_xor0 = s_dadda_pg_rca24_fa66_xor1 ^ s_dadda_pg_rca24_fa67_xor1;
  assign s_dadda_pg_rca24_fa344_and0 = s_dadda_pg_rca24_fa66_xor1 & s_dadda_pg_rca24_fa67_xor1;
  assign s_dadda_pg_rca24_fa344_xor1 = s_dadda_pg_rca24_fa344_xor0 ^ s_dadda_pg_rca24_fa68_xor1;
  assign s_dadda_pg_rca24_fa344_and1 = s_dadda_pg_rca24_fa344_xor0 & s_dadda_pg_rca24_fa68_xor1;
  assign s_dadda_pg_rca24_fa344_or0 = s_dadda_pg_rca24_fa344_and0 | s_dadda_pg_rca24_fa344_and1;
  assign s_dadda_pg_rca24_fa345_xor0 = s_dadda_pg_rca24_fa344_or0 ^ s_dadda_pg_rca24_fa343_or0;
  assign s_dadda_pg_rca24_fa345_and0 = s_dadda_pg_rca24_fa344_or0 & s_dadda_pg_rca24_fa343_or0;
  assign s_dadda_pg_rca24_fa345_xor1 = s_dadda_pg_rca24_fa345_xor0 ^ s_dadda_pg_rca24_fa75_xor1;
  assign s_dadda_pg_rca24_fa345_and1 = s_dadda_pg_rca24_fa345_xor0 & s_dadda_pg_rca24_fa75_xor1;
  assign s_dadda_pg_rca24_fa345_or0 = s_dadda_pg_rca24_fa345_and0 | s_dadda_pg_rca24_fa345_and1;
  assign s_dadda_pg_rca24_fa346_xor0 = s_dadda_pg_rca24_fa76_xor1 ^ s_dadda_pg_rca24_fa77_xor1;
  assign s_dadda_pg_rca24_fa346_and0 = s_dadda_pg_rca24_fa76_xor1 & s_dadda_pg_rca24_fa77_xor1;
  assign s_dadda_pg_rca24_fa346_xor1 = s_dadda_pg_rca24_fa346_xor0 ^ s_dadda_pg_rca24_fa78_xor1;
  assign s_dadda_pg_rca24_fa346_and1 = s_dadda_pg_rca24_fa346_xor0 & s_dadda_pg_rca24_fa78_xor1;
  assign s_dadda_pg_rca24_fa346_or0 = s_dadda_pg_rca24_fa346_and0 | s_dadda_pg_rca24_fa346_and1;
  assign s_dadda_pg_rca24_fa347_xor0 = s_dadda_pg_rca24_fa346_or0 ^ s_dadda_pg_rca24_fa345_or0;
  assign s_dadda_pg_rca24_fa347_and0 = s_dadda_pg_rca24_fa346_or0 & s_dadda_pg_rca24_fa345_or0;
  assign s_dadda_pg_rca24_fa347_xor1 = s_dadda_pg_rca24_fa347_xor0 ^ s_dadda_pg_rca24_fa86_xor1;
  assign s_dadda_pg_rca24_fa347_and1 = s_dadda_pg_rca24_fa347_xor0 & s_dadda_pg_rca24_fa86_xor1;
  assign s_dadda_pg_rca24_fa347_or0 = s_dadda_pg_rca24_fa347_and0 | s_dadda_pg_rca24_fa347_and1;
  assign s_dadda_pg_rca24_fa348_xor0 = s_dadda_pg_rca24_fa87_xor1 ^ s_dadda_pg_rca24_fa88_xor1;
  assign s_dadda_pg_rca24_fa348_and0 = s_dadda_pg_rca24_fa87_xor1 & s_dadda_pg_rca24_fa88_xor1;
  assign s_dadda_pg_rca24_fa348_xor1 = s_dadda_pg_rca24_fa348_xor0 ^ s_dadda_pg_rca24_fa89_xor1;
  assign s_dadda_pg_rca24_fa348_and1 = s_dadda_pg_rca24_fa348_xor0 & s_dadda_pg_rca24_fa89_xor1;
  assign s_dadda_pg_rca24_fa348_or0 = s_dadda_pg_rca24_fa348_and0 | s_dadda_pg_rca24_fa348_and1;
  assign s_dadda_pg_rca24_fa349_xor0 = s_dadda_pg_rca24_fa348_or0 ^ s_dadda_pg_rca24_fa347_or0;
  assign s_dadda_pg_rca24_fa349_and0 = s_dadda_pg_rca24_fa348_or0 & s_dadda_pg_rca24_fa347_or0;
  assign s_dadda_pg_rca24_fa349_xor1 = s_dadda_pg_rca24_fa349_xor0 ^ s_dadda_pg_rca24_fa98_xor1;
  assign s_dadda_pg_rca24_fa349_and1 = s_dadda_pg_rca24_fa349_xor0 & s_dadda_pg_rca24_fa98_xor1;
  assign s_dadda_pg_rca24_fa349_or0 = s_dadda_pg_rca24_fa349_and0 | s_dadda_pg_rca24_fa349_and1;
  assign s_dadda_pg_rca24_fa350_xor0 = s_dadda_pg_rca24_fa99_xor1 ^ s_dadda_pg_rca24_fa100_xor1;
  assign s_dadda_pg_rca24_fa350_and0 = s_dadda_pg_rca24_fa99_xor1 & s_dadda_pg_rca24_fa100_xor1;
  assign s_dadda_pg_rca24_fa350_xor1 = s_dadda_pg_rca24_fa350_xor0 ^ s_dadda_pg_rca24_fa101_xor1;
  assign s_dadda_pg_rca24_fa350_and1 = s_dadda_pg_rca24_fa350_xor0 & s_dadda_pg_rca24_fa101_xor1;
  assign s_dadda_pg_rca24_fa350_or0 = s_dadda_pg_rca24_fa350_and0 | s_dadda_pg_rca24_fa350_and1;
  assign s_dadda_pg_rca24_fa351_xor0 = s_dadda_pg_rca24_fa350_or0 ^ s_dadda_pg_rca24_fa349_or0;
  assign s_dadda_pg_rca24_fa351_and0 = s_dadda_pg_rca24_fa350_or0 & s_dadda_pg_rca24_fa349_or0;
  assign s_dadda_pg_rca24_fa351_xor1 = s_dadda_pg_rca24_fa351_xor0 ^ s_dadda_pg_rca24_fa110_xor1;
  assign s_dadda_pg_rca24_fa351_and1 = s_dadda_pg_rca24_fa351_xor0 & s_dadda_pg_rca24_fa110_xor1;
  assign s_dadda_pg_rca24_fa351_or0 = s_dadda_pg_rca24_fa351_and0 | s_dadda_pg_rca24_fa351_and1;
  assign s_dadda_pg_rca24_fa352_xor0 = s_dadda_pg_rca24_fa111_xor1 ^ s_dadda_pg_rca24_fa112_xor1;
  assign s_dadda_pg_rca24_fa352_and0 = s_dadda_pg_rca24_fa111_xor1 & s_dadda_pg_rca24_fa112_xor1;
  assign s_dadda_pg_rca24_fa352_xor1 = s_dadda_pg_rca24_fa352_xor0 ^ s_dadda_pg_rca24_fa113_xor1;
  assign s_dadda_pg_rca24_fa352_and1 = s_dadda_pg_rca24_fa352_xor0 & s_dadda_pg_rca24_fa113_xor1;
  assign s_dadda_pg_rca24_fa352_or0 = s_dadda_pg_rca24_fa352_and0 | s_dadda_pg_rca24_fa352_and1;
  assign s_dadda_pg_rca24_fa353_xor0 = s_dadda_pg_rca24_fa352_or0 ^ s_dadda_pg_rca24_fa351_or0;
  assign s_dadda_pg_rca24_fa353_and0 = s_dadda_pg_rca24_fa352_or0 & s_dadda_pg_rca24_fa351_or0;
  assign s_dadda_pg_rca24_fa353_xor1 = s_dadda_pg_rca24_fa353_xor0 ^ s_dadda_pg_rca24_fa123_xor1;
  assign s_dadda_pg_rca24_fa353_and1 = s_dadda_pg_rca24_fa353_xor0 & s_dadda_pg_rca24_fa123_xor1;
  assign s_dadda_pg_rca24_fa353_or0 = s_dadda_pg_rca24_fa353_and0 | s_dadda_pg_rca24_fa353_and1;
  assign s_dadda_pg_rca24_fa354_xor0 = s_dadda_pg_rca24_fa124_xor1 ^ s_dadda_pg_rca24_fa125_xor1;
  assign s_dadda_pg_rca24_fa354_and0 = s_dadda_pg_rca24_fa124_xor1 & s_dadda_pg_rca24_fa125_xor1;
  assign s_dadda_pg_rca24_fa354_xor1 = s_dadda_pg_rca24_fa354_xor0 ^ s_dadda_pg_rca24_fa126_xor1;
  assign s_dadda_pg_rca24_fa354_and1 = s_dadda_pg_rca24_fa354_xor0 & s_dadda_pg_rca24_fa126_xor1;
  assign s_dadda_pg_rca24_fa354_or0 = s_dadda_pg_rca24_fa354_and0 | s_dadda_pg_rca24_fa354_and1;
  assign s_dadda_pg_rca24_fa355_xor0 = s_dadda_pg_rca24_fa354_or0 ^ s_dadda_pg_rca24_fa353_or0;
  assign s_dadda_pg_rca24_fa355_and0 = s_dadda_pg_rca24_fa354_or0 & s_dadda_pg_rca24_fa353_or0;
  assign s_dadda_pg_rca24_fa355_xor1 = s_dadda_pg_rca24_fa355_xor0 ^ s_dadda_pg_rca24_fa136_xor1;
  assign s_dadda_pg_rca24_fa355_and1 = s_dadda_pg_rca24_fa355_xor0 & s_dadda_pg_rca24_fa136_xor1;
  assign s_dadda_pg_rca24_fa355_or0 = s_dadda_pg_rca24_fa355_and0 | s_dadda_pg_rca24_fa355_and1;
  assign s_dadda_pg_rca24_fa356_xor0 = s_dadda_pg_rca24_fa137_xor1 ^ s_dadda_pg_rca24_fa138_xor1;
  assign s_dadda_pg_rca24_fa356_and0 = s_dadda_pg_rca24_fa137_xor1 & s_dadda_pg_rca24_fa138_xor1;
  assign s_dadda_pg_rca24_fa356_xor1 = s_dadda_pg_rca24_fa356_xor0 ^ s_dadda_pg_rca24_fa139_xor1;
  assign s_dadda_pg_rca24_fa356_and1 = s_dadda_pg_rca24_fa356_xor0 & s_dadda_pg_rca24_fa139_xor1;
  assign s_dadda_pg_rca24_fa356_or0 = s_dadda_pg_rca24_fa356_and0 | s_dadda_pg_rca24_fa356_and1;
  assign s_dadda_pg_rca24_fa357_xor0 = s_dadda_pg_rca24_fa356_or0 ^ s_dadda_pg_rca24_fa355_or0;
  assign s_dadda_pg_rca24_fa357_and0 = s_dadda_pg_rca24_fa356_or0 & s_dadda_pg_rca24_fa355_or0;
  assign s_dadda_pg_rca24_fa357_xor1 = s_dadda_pg_rca24_fa357_xor0 ^ s_dadda_pg_rca24_fa149_xor1;
  assign s_dadda_pg_rca24_fa357_and1 = s_dadda_pg_rca24_fa357_xor0 & s_dadda_pg_rca24_fa149_xor1;
  assign s_dadda_pg_rca24_fa357_or0 = s_dadda_pg_rca24_fa357_and0 | s_dadda_pg_rca24_fa357_and1;
  assign s_dadda_pg_rca24_fa358_xor0 = s_dadda_pg_rca24_fa150_xor1 ^ s_dadda_pg_rca24_fa151_xor1;
  assign s_dadda_pg_rca24_fa358_and0 = s_dadda_pg_rca24_fa150_xor1 & s_dadda_pg_rca24_fa151_xor1;
  assign s_dadda_pg_rca24_fa358_xor1 = s_dadda_pg_rca24_fa358_xor0 ^ s_dadda_pg_rca24_fa152_xor1;
  assign s_dadda_pg_rca24_fa358_and1 = s_dadda_pg_rca24_fa358_xor0 & s_dadda_pg_rca24_fa152_xor1;
  assign s_dadda_pg_rca24_fa358_or0 = s_dadda_pg_rca24_fa358_and0 | s_dadda_pg_rca24_fa358_and1;
  assign s_dadda_pg_rca24_fa359_xor0 = s_dadda_pg_rca24_fa358_or0 ^ s_dadda_pg_rca24_fa357_or0;
  assign s_dadda_pg_rca24_fa359_and0 = s_dadda_pg_rca24_fa358_or0 & s_dadda_pg_rca24_fa357_or0;
  assign s_dadda_pg_rca24_fa359_xor1 = s_dadda_pg_rca24_fa359_xor0 ^ s_dadda_pg_rca24_fa162_xor1;
  assign s_dadda_pg_rca24_fa359_and1 = s_dadda_pg_rca24_fa359_xor0 & s_dadda_pg_rca24_fa162_xor1;
  assign s_dadda_pg_rca24_fa359_or0 = s_dadda_pg_rca24_fa359_and0 | s_dadda_pg_rca24_fa359_and1;
  assign s_dadda_pg_rca24_fa360_xor0 = s_dadda_pg_rca24_fa163_xor1 ^ s_dadda_pg_rca24_fa164_xor1;
  assign s_dadda_pg_rca24_fa360_and0 = s_dadda_pg_rca24_fa163_xor1 & s_dadda_pg_rca24_fa164_xor1;
  assign s_dadda_pg_rca24_fa360_xor1 = s_dadda_pg_rca24_fa360_xor0 ^ s_dadda_pg_rca24_fa165_xor1;
  assign s_dadda_pg_rca24_fa360_and1 = s_dadda_pg_rca24_fa360_xor0 & s_dadda_pg_rca24_fa165_xor1;
  assign s_dadda_pg_rca24_fa360_or0 = s_dadda_pg_rca24_fa360_and0 | s_dadda_pg_rca24_fa360_and1;
  assign s_dadda_pg_rca24_fa361_xor0 = s_dadda_pg_rca24_fa360_or0 ^ s_dadda_pg_rca24_fa359_or0;
  assign s_dadda_pg_rca24_fa361_and0 = s_dadda_pg_rca24_fa360_or0 & s_dadda_pg_rca24_fa359_or0;
  assign s_dadda_pg_rca24_fa361_xor1 = s_dadda_pg_rca24_fa361_xor0 ^ s_dadda_pg_rca24_fa175_xor1;
  assign s_dadda_pg_rca24_fa361_and1 = s_dadda_pg_rca24_fa361_xor0 & s_dadda_pg_rca24_fa175_xor1;
  assign s_dadda_pg_rca24_fa361_or0 = s_dadda_pg_rca24_fa361_and0 | s_dadda_pg_rca24_fa361_and1;
  assign s_dadda_pg_rca24_fa362_xor0 = s_dadda_pg_rca24_fa176_xor1 ^ s_dadda_pg_rca24_fa177_xor1;
  assign s_dadda_pg_rca24_fa362_and0 = s_dadda_pg_rca24_fa176_xor1 & s_dadda_pg_rca24_fa177_xor1;
  assign s_dadda_pg_rca24_fa362_xor1 = s_dadda_pg_rca24_fa362_xor0 ^ s_dadda_pg_rca24_fa178_xor1;
  assign s_dadda_pg_rca24_fa362_and1 = s_dadda_pg_rca24_fa362_xor0 & s_dadda_pg_rca24_fa178_xor1;
  assign s_dadda_pg_rca24_fa362_or0 = s_dadda_pg_rca24_fa362_and0 | s_dadda_pg_rca24_fa362_and1;
  assign s_dadda_pg_rca24_fa363_xor0 = s_dadda_pg_rca24_fa362_or0 ^ s_dadda_pg_rca24_fa361_or0;
  assign s_dadda_pg_rca24_fa363_and0 = s_dadda_pg_rca24_fa362_or0 & s_dadda_pg_rca24_fa361_or0;
  assign s_dadda_pg_rca24_fa363_xor1 = s_dadda_pg_rca24_fa363_xor0 ^ s_dadda_pg_rca24_fa188_xor1;
  assign s_dadda_pg_rca24_fa363_and1 = s_dadda_pg_rca24_fa363_xor0 & s_dadda_pg_rca24_fa188_xor1;
  assign s_dadda_pg_rca24_fa363_or0 = s_dadda_pg_rca24_fa363_and0 | s_dadda_pg_rca24_fa363_and1;
  assign s_dadda_pg_rca24_fa364_xor0 = s_dadda_pg_rca24_fa189_xor1 ^ s_dadda_pg_rca24_fa190_xor1;
  assign s_dadda_pg_rca24_fa364_and0 = s_dadda_pg_rca24_fa189_xor1 & s_dadda_pg_rca24_fa190_xor1;
  assign s_dadda_pg_rca24_fa364_xor1 = s_dadda_pg_rca24_fa364_xor0 ^ s_dadda_pg_rca24_fa191_xor1;
  assign s_dadda_pg_rca24_fa364_and1 = s_dadda_pg_rca24_fa364_xor0 & s_dadda_pg_rca24_fa191_xor1;
  assign s_dadda_pg_rca24_fa364_or0 = s_dadda_pg_rca24_fa364_and0 | s_dadda_pg_rca24_fa364_and1;
  assign s_dadda_pg_rca24_fa365_xor0 = s_dadda_pg_rca24_fa364_or0 ^ s_dadda_pg_rca24_fa363_or0;
  assign s_dadda_pg_rca24_fa365_and0 = s_dadda_pg_rca24_fa364_or0 & s_dadda_pg_rca24_fa363_or0;
  assign s_dadda_pg_rca24_fa365_xor1 = s_dadda_pg_rca24_fa365_xor0 ^ s_dadda_pg_rca24_fa201_xor1;
  assign s_dadda_pg_rca24_fa365_and1 = s_dadda_pg_rca24_fa365_xor0 & s_dadda_pg_rca24_fa201_xor1;
  assign s_dadda_pg_rca24_fa365_or0 = s_dadda_pg_rca24_fa365_and0 | s_dadda_pg_rca24_fa365_and1;
  assign s_dadda_pg_rca24_fa366_xor0 = s_dadda_pg_rca24_fa202_xor1 ^ s_dadda_pg_rca24_fa203_xor1;
  assign s_dadda_pg_rca24_fa366_and0 = s_dadda_pg_rca24_fa202_xor1 & s_dadda_pg_rca24_fa203_xor1;
  assign s_dadda_pg_rca24_fa366_xor1 = s_dadda_pg_rca24_fa366_xor0 ^ s_dadda_pg_rca24_fa204_xor1;
  assign s_dadda_pg_rca24_fa366_and1 = s_dadda_pg_rca24_fa366_xor0 & s_dadda_pg_rca24_fa204_xor1;
  assign s_dadda_pg_rca24_fa366_or0 = s_dadda_pg_rca24_fa366_and0 | s_dadda_pg_rca24_fa366_and1;
  assign s_dadda_pg_rca24_fa367_xor0 = s_dadda_pg_rca24_fa366_or0 ^ s_dadda_pg_rca24_fa365_or0;
  assign s_dadda_pg_rca24_fa367_and0 = s_dadda_pg_rca24_fa366_or0 & s_dadda_pg_rca24_fa365_or0;
  assign s_dadda_pg_rca24_fa367_xor1 = s_dadda_pg_rca24_fa367_xor0 ^ s_dadda_pg_rca24_fa214_xor1;
  assign s_dadda_pg_rca24_fa367_and1 = s_dadda_pg_rca24_fa367_xor0 & s_dadda_pg_rca24_fa214_xor1;
  assign s_dadda_pg_rca24_fa367_or0 = s_dadda_pg_rca24_fa367_and0 | s_dadda_pg_rca24_fa367_and1;
  assign s_dadda_pg_rca24_fa368_xor0 = s_dadda_pg_rca24_fa215_xor1 ^ s_dadda_pg_rca24_fa216_xor1;
  assign s_dadda_pg_rca24_fa368_and0 = s_dadda_pg_rca24_fa215_xor1 & s_dadda_pg_rca24_fa216_xor1;
  assign s_dadda_pg_rca24_fa368_xor1 = s_dadda_pg_rca24_fa368_xor0 ^ s_dadda_pg_rca24_fa217_xor1;
  assign s_dadda_pg_rca24_fa368_and1 = s_dadda_pg_rca24_fa368_xor0 & s_dadda_pg_rca24_fa217_xor1;
  assign s_dadda_pg_rca24_fa368_or0 = s_dadda_pg_rca24_fa368_and0 | s_dadda_pg_rca24_fa368_and1;
  assign s_dadda_pg_rca24_fa369_xor0 = s_dadda_pg_rca24_fa368_or0 ^ s_dadda_pg_rca24_fa367_or0;
  assign s_dadda_pg_rca24_fa369_and0 = s_dadda_pg_rca24_fa368_or0 & s_dadda_pg_rca24_fa367_or0;
  assign s_dadda_pg_rca24_fa369_xor1 = s_dadda_pg_rca24_fa369_xor0 ^ s_dadda_pg_rca24_fa227_xor1;
  assign s_dadda_pg_rca24_fa369_and1 = s_dadda_pg_rca24_fa369_xor0 & s_dadda_pg_rca24_fa227_xor1;
  assign s_dadda_pg_rca24_fa369_or0 = s_dadda_pg_rca24_fa369_and0 | s_dadda_pg_rca24_fa369_and1;
  assign s_dadda_pg_rca24_fa370_xor0 = s_dadda_pg_rca24_fa228_xor1 ^ s_dadda_pg_rca24_fa229_xor1;
  assign s_dadda_pg_rca24_fa370_and0 = s_dadda_pg_rca24_fa228_xor1 & s_dadda_pg_rca24_fa229_xor1;
  assign s_dadda_pg_rca24_fa370_xor1 = s_dadda_pg_rca24_fa370_xor0 ^ s_dadda_pg_rca24_fa230_xor1;
  assign s_dadda_pg_rca24_fa370_and1 = s_dadda_pg_rca24_fa370_xor0 & s_dadda_pg_rca24_fa230_xor1;
  assign s_dadda_pg_rca24_fa370_or0 = s_dadda_pg_rca24_fa370_and0 | s_dadda_pg_rca24_fa370_and1;
  assign s_dadda_pg_rca24_fa371_xor0 = s_dadda_pg_rca24_fa370_or0 ^ s_dadda_pg_rca24_fa369_or0;
  assign s_dadda_pg_rca24_fa371_and0 = s_dadda_pg_rca24_fa370_or0 & s_dadda_pg_rca24_fa369_or0;
  assign s_dadda_pg_rca24_fa371_xor1 = s_dadda_pg_rca24_fa371_xor0 ^ s_dadda_pg_rca24_fa240_xor1;
  assign s_dadda_pg_rca24_fa371_and1 = s_dadda_pg_rca24_fa371_xor0 & s_dadda_pg_rca24_fa240_xor1;
  assign s_dadda_pg_rca24_fa371_or0 = s_dadda_pg_rca24_fa371_and0 | s_dadda_pg_rca24_fa371_and1;
  assign s_dadda_pg_rca24_fa372_xor0 = s_dadda_pg_rca24_fa241_xor1 ^ s_dadda_pg_rca24_fa242_xor1;
  assign s_dadda_pg_rca24_fa372_and0 = s_dadda_pg_rca24_fa241_xor1 & s_dadda_pg_rca24_fa242_xor1;
  assign s_dadda_pg_rca24_fa372_xor1 = s_dadda_pg_rca24_fa372_xor0 ^ s_dadda_pg_rca24_fa243_xor1;
  assign s_dadda_pg_rca24_fa372_and1 = s_dadda_pg_rca24_fa372_xor0 & s_dadda_pg_rca24_fa243_xor1;
  assign s_dadda_pg_rca24_fa372_or0 = s_dadda_pg_rca24_fa372_and0 | s_dadda_pg_rca24_fa372_and1;
  assign s_dadda_pg_rca24_fa373_xor0 = s_dadda_pg_rca24_fa372_or0 ^ s_dadda_pg_rca24_fa371_or0;
  assign s_dadda_pg_rca24_fa373_and0 = s_dadda_pg_rca24_fa372_or0 & s_dadda_pg_rca24_fa371_or0;
  assign s_dadda_pg_rca24_fa373_xor1 = s_dadda_pg_rca24_fa373_xor0 ^ s_dadda_pg_rca24_fa252_xor1;
  assign s_dadda_pg_rca24_fa373_and1 = s_dadda_pg_rca24_fa373_xor0 & s_dadda_pg_rca24_fa252_xor1;
  assign s_dadda_pg_rca24_fa373_or0 = s_dadda_pg_rca24_fa373_and0 | s_dadda_pg_rca24_fa373_and1;
  assign s_dadda_pg_rca24_fa374_xor0 = s_dadda_pg_rca24_fa253_xor1 ^ s_dadda_pg_rca24_fa254_xor1;
  assign s_dadda_pg_rca24_fa374_and0 = s_dadda_pg_rca24_fa253_xor1 & s_dadda_pg_rca24_fa254_xor1;
  assign s_dadda_pg_rca24_fa374_xor1 = s_dadda_pg_rca24_fa374_xor0 ^ s_dadda_pg_rca24_fa255_xor1;
  assign s_dadda_pg_rca24_fa374_and1 = s_dadda_pg_rca24_fa374_xor0 & s_dadda_pg_rca24_fa255_xor1;
  assign s_dadda_pg_rca24_fa374_or0 = s_dadda_pg_rca24_fa374_and0 | s_dadda_pg_rca24_fa374_and1;
  assign s_dadda_pg_rca24_fa375_xor0 = s_dadda_pg_rca24_fa374_or0 ^ s_dadda_pg_rca24_fa373_or0;
  assign s_dadda_pg_rca24_fa375_and0 = s_dadda_pg_rca24_fa374_or0 & s_dadda_pg_rca24_fa373_or0;
  assign s_dadda_pg_rca24_fa375_xor1 = s_dadda_pg_rca24_fa375_xor0 ^ s_dadda_pg_rca24_fa263_xor1;
  assign s_dadda_pg_rca24_fa375_and1 = s_dadda_pg_rca24_fa375_xor0 & s_dadda_pg_rca24_fa263_xor1;
  assign s_dadda_pg_rca24_fa375_or0 = s_dadda_pg_rca24_fa375_and0 | s_dadda_pg_rca24_fa375_and1;
  assign s_dadda_pg_rca24_fa376_xor0 = s_dadda_pg_rca24_fa264_xor1 ^ s_dadda_pg_rca24_fa265_xor1;
  assign s_dadda_pg_rca24_fa376_and0 = s_dadda_pg_rca24_fa264_xor1 & s_dadda_pg_rca24_fa265_xor1;
  assign s_dadda_pg_rca24_fa376_xor1 = s_dadda_pg_rca24_fa376_xor0 ^ s_dadda_pg_rca24_fa266_xor1;
  assign s_dadda_pg_rca24_fa376_and1 = s_dadda_pg_rca24_fa376_xor0 & s_dadda_pg_rca24_fa266_xor1;
  assign s_dadda_pg_rca24_fa376_or0 = s_dadda_pg_rca24_fa376_and0 | s_dadda_pg_rca24_fa376_and1;
  assign s_dadda_pg_rca24_fa377_xor0 = s_dadda_pg_rca24_fa376_or0 ^ s_dadda_pg_rca24_fa375_or0;
  assign s_dadda_pg_rca24_fa377_and0 = s_dadda_pg_rca24_fa376_or0 & s_dadda_pg_rca24_fa375_or0;
  assign s_dadda_pg_rca24_fa377_xor1 = s_dadda_pg_rca24_fa377_xor0 ^ s_dadda_pg_rca24_fa273_xor1;
  assign s_dadda_pg_rca24_fa377_and1 = s_dadda_pg_rca24_fa377_xor0 & s_dadda_pg_rca24_fa273_xor1;
  assign s_dadda_pg_rca24_fa377_or0 = s_dadda_pg_rca24_fa377_and0 | s_dadda_pg_rca24_fa377_and1;
  assign s_dadda_pg_rca24_fa378_xor0 = s_dadda_pg_rca24_fa274_xor1 ^ s_dadda_pg_rca24_fa275_xor1;
  assign s_dadda_pg_rca24_fa378_and0 = s_dadda_pg_rca24_fa274_xor1 & s_dadda_pg_rca24_fa275_xor1;
  assign s_dadda_pg_rca24_fa378_xor1 = s_dadda_pg_rca24_fa378_xor0 ^ s_dadda_pg_rca24_fa276_xor1;
  assign s_dadda_pg_rca24_fa378_and1 = s_dadda_pg_rca24_fa378_xor0 & s_dadda_pg_rca24_fa276_xor1;
  assign s_dadda_pg_rca24_fa378_or0 = s_dadda_pg_rca24_fa378_and0 | s_dadda_pg_rca24_fa378_and1;
  assign s_dadda_pg_rca24_fa379_xor0 = s_dadda_pg_rca24_fa378_or0 ^ s_dadda_pg_rca24_fa377_or0;
  assign s_dadda_pg_rca24_fa379_and0 = s_dadda_pg_rca24_fa378_or0 & s_dadda_pg_rca24_fa377_or0;
  assign s_dadda_pg_rca24_fa379_xor1 = s_dadda_pg_rca24_fa379_xor0 ^ s_dadda_pg_rca24_fa282_xor1;
  assign s_dadda_pg_rca24_fa379_and1 = s_dadda_pg_rca24_fa379_xor0 & s_dadda_pg_rca24_fa282_xor1;
  assign s_dadda_pg_rca24_fa379_or0 = s_dadda_pg_rca24_fa379_and0 | s_dadda_pg_rca24_fa379_and1;
  assign s_dadda_pg_rca24_fa380_xor0 = s_dadda_pg_rca24_fa283_xor1 ^ s_dadda_pg_rca24_fa284_xor1;
  assign s_dadda_pg_rca24_fa380_and0 = s_dadda_pg_rca24_fa283_xor1 & s_dadda_pg_rca24_fa284_xor1;
  assign s_dadda_pg_rca24_fa380_xor1 = s_dadda_pg_rca24_fa380_xor0 ^ s_dadda_pg_rca24_fa285_xor1;
  assign s_dadda_pg_rca24_fa380_and1 = s_dadda_pg_rca24_fa380_xor0 & s_dadda_pg_rca24_fa285_xor1;
  assign s_dadda_pg_rca24_fa380_or0 = s_dadda_pg_rca24_fa380_and0 | s_dadda_pg_rca24_fa380_and1;
  assign s_dadda_pg_rca24_fa381_xor0 = s_dadda_pg_rca24_fa380_or0 ^ s_dadda_pg_rca24_fa379_or0;
  assign s_dadda_pg_rca24_fa381_and0 = s_dadda_pg_rca24_fa380_or0 & s_dadda_pg_rca24_fa379_or0;
  assign s_dadda_pg_rca24_fa381_xor1 = s_dadda_pg_rca24_fa381_xor0 ^ s_dadda_pg_rca24_fa290_xor1;
  assign s_dadda_pg_rca24_fa381_and1 = s_dadda_pg_rca24_fa381_xor0 & s_dadda_pg_rca24_fa290_xor1;
  assign s_dadda_pg_rca24_fa381_or0 = s_dadda_pg_rca24_fa381_and0 | s_dadda_pg_rca24_fa381_and1;
  assign s_dadda_pg_rca24_fa382_xor0 = s_dadda_pg_rca24_fa291_xor1 ^ s_dadda_pg_rca24_fa292_xor1;
  assign s_dadda_pg_rca24_fa382_and0 = s_dadda_pg_rca24_fa291_xor1 & s_dadda_pg_rca24_fa292_xor1;
  assign s_dadda_pg_rca24_fa382_xor1 = s_dadda_pg_rca24_fa382_xor0 ^ s_dadda_pg_rca24_fa293_xor1;
  assign s_dadda_pg_rca24_fa382_and1 = s_dadda_pg_rca24_fa382_xor0 & s_dadda_pg_rca24_fa293_xor1;
  assign s_dadda_pg_rca24_fa382_or0 = s_dadda_pg_rca24_fa382_and0 | s_dadda_pg_rca24_fa382_and1;
  assign s_dadda_pg_rca24_fa383_xor0 = s_dadda_pg_rca24_fa382_or0 ^ s_dadda_pg_rca24_fa381_or0;
  assign s_dadda_pg_rca24_fa383_and0 = s_dadda_pg_rca24_fa382_or0 & s_dadda_pg_rca24_fa381_or0;
  assign s_dadda_pg_rca24_fa383_xor1 = s_dadda_pg_rca24_fa383_xor0 ^ s_dadda_pg_rca24_fa297_xor1;
  assign s_dadda_pg_rca24_fa383_and1 = s_dadda_pg_rca24_fa383_xor0 & s_dadda_pg_rca24_fa297_xor1;
  assign s_dadda_pg_rca24_fa383_or0 = s_dadda_pg_rca24_fa383_and0 | s_dadda_pg_rca24_fa383_and1;
  assign s_dadda_pg_rca24_fa384_xor0 = s_dadda_pg_rca24_fa298_xor1 ^ s_dadda_pg_rca24_fa299_xor1;
  assign s_dadda_pg_rca24_fa384_and0 = s_dadda_pg_rca24_fa298_xor1 & s_dadda_pg_rca24_fa299_xor1;
  assign s_dadda_pg_rca24_fa384_xor1 = s_dadda_pg_rca24_fa384_xor0 ^ s_dadda_pg_rca24_fa300_xor1;
  assign s_dadda_pg_rca24_fa384_and1 = s_dadda_pg_rca24_fa384_xor0 & s_dadda_pg_rca24_fa300_xor1;
  assign s_dadda_pg_rca24_fa384_or0 = s_dadda_pg_rca24_fa384_and0 | s_dadda_pg_rca24_fa384_and1;
  assign s_dadda_pg_rca24_fa385_xor0 = s_dadda_pg_rca24_fa384_or0 ^ s_dadda_pg_rca24_fa383_or0;
  assign s_dadda_pg_rca24_fa385_and0 = s_dadda_pg_rca24_fa384_or0 & s_dadda_pg_rca24_fa383_or0;
  assign s_dadda_pg_rca24_fa385_xor1 = s_dadda_pg_rca24_fa385_xor0 ^ s_dadda_pg_rca24_fa303_xor1;
  assign s_dadda_pg_rca24_fa385_and1 = s_dadda_pg_rca24_fa385_xor0 & s_dadda_pg_rca24_fa303_xor1;
  assign s_dadda_pg_rca24_fa385_or0 = s_dadda_pg_rca24_fa385_and0 | s_dadda_pg_rca24_fa385_and1;
  assign s_dadda_pg_rca24_fa386_xor0 = s_dadda_pg_rca24_fa304_xor1 ^ s_dadda_pg_rca24_fa305_xor1;
  assign s_dadda_pg_rca24_fa386_and0 = s_dadda_pg_rca24_fa304_xor1 & s_dadda_pg_rca24_fa305_xor1;
  assign s_dadda_pg_rca24_fa386_xor1 = s_dadda_pg_rca24_fa386_xor0 ^ s_dadda_pg_rca24_fa306_xor1;
  assign s_dadda_pg_rca24_fa386_and1 = s_dadda_pg_rca24_fa386_xor0 & s_dadda_pg_rca24_fa306_xor1;
  assign s_dadda_pg_rca24_fa386_or0 = s_dadda_pg_rca24_fa386_and0 | s_dadda_pg_rca24_fa386_and1;
  assign s_dadda_pg_rca24_nand_14_23 = ~(a[14] & b[23]);
  assign s_dadda_pg_rca24_fa387_xor0 = s_dadda_pg_rca24_fa386_or0 ^ s_dadda_pg_rca24_fa385_or0;
  assign s_dadda_pg_rca24_fa387_and0 = s_dadda_pg_rca24_fa386_or0 & s_dadda_pg_rca24_fa385_or0;
  assign s_dadda_pg_rca24_fa387_xor1 = s_dadda_pg_rca24_fa387_xor0 ^ s_dadda_pg_rca24_nand_14_23;
  assign s_dadda_pg_rca24_fa387_and1 = s_dadda_pg_rca24_fa387_xor0 & s_dadda_pg_rca24_nand_14_23;
  assign s_dadda_pg_rca24_fa387_or0 = s_dadda_pg_rca24_fa387_and0 | s_dadda_pg_rca24_fa387_and1;
  assign s_dadda_pg_rca24_fa388_xor0 = s_dadda_pg_rca24_fa309_xor1 ^ s_dadda_pg_rca24_fa310_xor1;
  assign s_dadda_pg_rca24_fa388_and0 = s_dadda_pg_rca24_fa309_xor1 & s_dadda_pg_rca24_fa310_xor1;
  assign s_dadda_pg_rca24_fa388_xor1 = s_dadda_pg_rca24_fa388_xor0 ^ s_dadda_pg_rca24_fa311_xor1;
  assign s_dadda_pg_rca24_fa388_and1 = s_dadda_pg_rca24_fa388_xor0 & s_dadda_pg_rca24_fa311_xor1;
  assign s_dadda_pg_rca24_fa388_or0 = s_dadda_pg_rca24_fa388_and0 | s_dadda_pg_rca24_fa388_and1;
  assign s_dadda_pg_rca24_and_16_22 = a[16] & b[22];
  assign s_dadda_pg_rca24_fa389_xor0 = s_dadda_pg_rca24_fa388_or0 ^ s_dadda_pg_rca24_fa387_or0;
  assign s_dadda_pg_rca24_fa389_and0 = s_dadda_pg_rca24_fa388_or0 & s_dadda_pg_rca24_fa387_or0;
  assign s_dadda_pg_rca24_fa389_xor1 = s_dadda_pg_rca24_fa389_xor0 ^ s_dadda_pg_rca24_and_16_22;
  assign s_dadda_pg_rca24_fa389_and1 = s_dadda_pg_rca24_fa389_xor0 & s_dadda_pg_rca24_and_16_22;
  assign s_dadda_pg_rca24_fa389_or0 = s_dadda_pg_rca24_fa389_and0 | s_dadda_pg_rca24_fa389_and1;
  assign s_dadda_pg_rca24_nand_15_23 = ~(a[15] & b[23]);
  assign s_dadda_pg_rca24_fa390_xor0 = s_dadda_pg_rca24_nand_15_23 ^ s_dadda_pg_rca24_fa314_xor1;
  assign s_dadda_pg_rca24_fa390_and0 = s_dadda_pg_rca24_nand_15_23 & s_dadda_pg_rca24_fa314_xor1;
  assign s_dadda_pg_rca24_fa390_xor1 = s_dadda_pg_rca24_fa390_xor0 ^ s_dadda_pg_rca24_fa315_xor1;
  assign s_dadda_pg_rca24_fa390_and1 = s_dadda_pg_rca24_fa390_xor0 & s_dadda_pg_rca24_fa315_xor1;
  assign s_dadda_pg_rca24_fa390_or0 = s_dadda_pg_rca24_fa390_and0 | s_dadda_pg_rca24_fa390_and1;
  assign s_dadda_pg_rca24_and_18_21 = a[18] & b[21];
  assign s_dadda_pg_rca24_fa391_xor0 = s_dadda_pg_rca24_fa390_or0 ^ s_dadda_pg_rca24_fa389_or0;
  assign s_dadda_pg_rca24_fa391_and0 = s_dadda_pg_rca24_fa390_or0 & s_dadda_pg_rca24_fa389_or0;
  assign s_dadda_pg_rca24_fa391_xor1 = s_dadda_pg_rca24_fa391_xor0 ^ s_dadda_pg_rca24_and_18_21;
  assign s_dadda_pg_rca24_fa391_and1 = s_dadda_pg_rca24_fa391_xor0 & s_dadda_pg_rca24_and_18_21;
  assign s_dadda_pg_rca24_fa391_or0 = s_dadda_pg_rca24_fa391_and0 | s_dadda_pg_rca24_fa391_and1;
  assign s_dadda_pg_rca24_and_17_22 = a[17] & b[22];
  assign s_dadda_pg_rca24_nand_16_23 = ~(a[16] & b[23]);
  assign s_dadda_pg_rca24_fa392_xor0 = s_dadda_pg_rca24_and_17_22 ^ s_dadda_pg_rca24_nand_16_23;
  assign s_dadda_pg_rca24_fa392_and0 = s_dadda_pg_rca24_and_17_22 & s_dadda_pg_rca24_nand_16_23;
  assign s_dadda_pg_rca24_fa392_xor1 = s_dadda_pg_rca24_fa392_xor0 ^ s_dadda_pg_rca24_fa318_xor1;
  assign s_dadda_pg_rca24_fa392_and1 = s_dadda_pg_rca24_fa392_xor0 & s_dadda_pg_rca24_fa318_xor1;
  assign s_dadda_pg_rca24_fa392_or0 = s_dadda_pg_rca24_fa392_and0 | s_dadda_pg_rca24_fa392_and1;
  assign s_dadda_pg_rca24_and_20_20 = a[20] & b[20];
  assign s_dadda_pg_rca24_fa393_xor0 = s_dadda_pg_rca24_fa392_or0 ^ s_dadda_pg_rca24_fa391_or0;
  assign s_dadda_pg_rca24_fa393_and0 = s_dadda_pg_rca24_fa392_or0 & s_dadda_pg_rca24_fa391_or0;
  assign s_dadda_pg_rca24_fa393_xor1 = s_dadda_pg_rca24_fa393_xor0 ^ s_dadda_pg_rca24_and_20_20;
  assign s_dadda_pg_rca24_fa393_and1 = s_dadda_pg_rca24_fa393_xor0 & s_dadda_pg_rca24_and_20_20;
  assign s_dadda_pg_rca24_fa393_or0 = s_dadda_pg_rca24_fa393_and0 | s_dadda_pg_rca24_fa393_and1;
  assign s_dadda_pg_rca24_and_19_21 = a[19] & b[21];
  assign s_dadda_pg_rca24_and_18_22 = a[18] & b[22];
  assign s_dadda_pg_rca24_nand_17_23 = ~(a[17] & b[23]);
  assign s_dadda_pg_rca24_fa394_xor0 = s_dadda_pg_rca24_and_19_21 ^ s_dadda_pg_rca24_and_18_22;
  assign s_dadda_pg_rca24_fa394_and0 = s_dadda_pg_rca24_and_19_21 & s_dadda_pg_rca24_and_18_22;
  assign s_dadda_pg_rca24_fa394_xor1 = s_dadda_pg_rca24_fa394_xor0 ^ s_dadda_pg_rca24_nand_17_23;
  assign s_dadda_pg_rca24_fa394_and1 = s_dadda_pg_rca24_fa394_xor0 & s_dadda_pg_rca24_nand_17_23;
  assign s_dadda_pg_rca24_fa394_or0 = s_dadda_pg_rca24_fa394_and0 | s_dadda_pg_rca24_fa394_and1;
  assign s_dadda_pg_rca24_and_22_19 = a[22] & b[19];
  assign s_dadda_pg_rca24_fa395_xor0 = s_dadda_pg_rca24_fa394_or0 ^ s_dadda_pg_rca24_fa393_or0;
  assign s_dadda_pg_rca24_fa395_and0 = s_dadda_pg_rca24_fa394_or0 & s_dadda_pg_rca24_fa393_or0;
  assign s_dadda_pg_rca24_fa395_xor1 = s_dadda_pg_rca24_fa395_xor0 ^ s_dadda_pg_rca24_and_22_19;
  assign s_dadda_pg_rca24_fa395_and1 = s_dadda_pg_rca24_fa395_xor0 & s_dadda_pg_rca24_and_22_19;
  assign s_dadda_pg_rca24_fa395_or0 = s_dadda_pg_rca24_fa395_and0 | s_dadda_pg_rca24_fa395_and1;
  assign s_dadda_pg_rca24_and_21_20 = a[21] & b[20];
  assign s_dadda_pg_rca24_and_20_21 = a[20] & b[21];
  assign s_dadda_pg_rca24_and_19_22 = a[19] & b[22];
  assign s_dadda_pg_rca24_fa396_xor0 = s_dadda_pg_rca24_and_21_20 ^ s_dadda_pg_rca24_and_20_21;
  assign s_dadda_pg_rca24_fa396_and0 = s_dadda_pg_rca24_and_21_20 & s_dadda_pg_rca24_and_20_21;
  assign s_dadda_pg_rca24_fa396_xor1 = s_dadda_pg_rca24_fa396_xor0 ^ s_dadda_pg_rca24_and_19_22;
  assign s_dadda_pg_rca24_fa396_and1 = s_dadda_pg_rca24_fa396_xor0 & s_dadda_pg_rca24_and_19_22;
  assign s_dadda_pg_rca24_fa396_or0 = s_dadda_pg_rca24_fa396_and0 | s_dadda_pg_rca24_fa396_and1;
  assign s_dadda_pg_rca24_fa397_xor0 = s_dadda_pg_rca24_fa396_or0 ^ s_dadda_pg_rca24_fa395_or0;
  assign s_dadda_pg_rca24_fa397_and0 = s_dadda_pg_rca24_fa396_or0 & s_dadda_pg_rca24_fa395_or0;
  assign s_dadda_pg_rca24_fa397_xor1 = s_dadda_pg_rca24_fa397_xor0 ^ s_dadda_pg_rca24_fa323_or0;
  assign s_dadda_pg_rca24_fa397_and1 = s_dadda_pg_rca24_fa397_xor0 & s_dadda_pg_rca24_fa323_or0;
  assign s_dadda_pg_rca24_fa397_or0 = s_dadda_pg_rca24_fa397_and0 | s_dadda_pg_rca24_fa397_and1;
  assign s_dadda_pg_rca24_nand_23_19 = ~(a[23] & b[19]);
  assign s_dadda_pg_rca24_and_22_20 = a[22] & b[20];
  assign s_dadda_pg_rca24_and_21_21 = a[21] & b[21];
  assign s_dadda_pg_rca24_fa398_xor0 = s_dadda_pg_rca24_nand_23_19 ^ s_dadda_pg_rca24_and_22_20;
  assign s_dadda_pg_rca24_fa398_and0 = s_dadda_pg_rca24_nand_23_19 & s_dadda_pg_rca24_and_22_20;
  assign s_dadda_pg_rca24_fa398_xor1 = s_dadda_pg_rca24_fa398_xor0 ^ s_dadda_pg_rca24_and_21_21;
  assign s_dadda_pg_rca24_fa398_and1 = s_dadda_pg_rca24_fa398_xor0 & s_dadda_pg_rca24_and_21_21;
  assign s_dadda_pg_rca24_fa398_or0 = s_dadda_pg_rca24_fa398_and0 | s_dadda_pg_rca24_fa398_and1;
  assign s_dadda_pg_rca24_nand_23_20 = ~(a[23] & b[20]);
  assign s_dadda_pg_rca24_fa399_xor0 = s_dadda_pg_rca24_fa398_or0 ^ s_dadda_pg_rca24_fa397_or0;
  assign s_dadda_pg_rca24_fa399_and0 = s_dadda_pg_rca24_fa398_or0 & s_dadda_pg_rca24_fa397_or0;
  assign s_dadda_pg_rca24_fa399_xor1 = s_dadda_pg_rca24_fa399_xor0 ^ s_dadda_pg_rca24_nand_23_20;
  assign s_dadda_pg_rca24_fa399_and1 = s_dadda_pg_rca24_fa399_xor0 & s_dadda_pg_rca24_nand_23_20;
  assign s_dadda_pg_rca24_fa399_or0 = s_dadda_pg_rca24_fa399_and0 | s_dadda_pg_rca24_fa399_and1;
  assign s_dadda_pg_rca24_and_3_0 = a[3] & b[0];
  assign s_dadda_pg_rca24_and_2_1 = a[2] & b[1];
  assign s_dadda_pg_rca24_ha20_xor0 = s_dadda_pg_rca24_and_3_0 ^ s_dadda_pg_rca24_and_2_1;
  assign s_dadda_pg_rca24_ha20_and0 = s_dadda_pg_rca24_and_3_0 & s_dadda_pg_rca24_and_2_1;
  assign s_dadda_pg_rca24_and_2_2 = a[2] & b[2];
  assign s_dadda_pg_rca24_and_1_3 = a[1] & b[3];
  assign s_dadda_pg_rca24_fa400_xor0 = s_dadda_pg_rca24_ha20_and0 ^ s_dadda_pg_rca24_and_2_2;
  assign s_dadda_pg_rca24_fa400_and0 = s_dadda_pg_rca24_ha20_and0 & s_dadda_pg_rca24_and_2_2;
  assign s_dadda_pg_rca24_fa400_xor1 = s_dadda_pg_rca24_fa400_xor0 ^ s_dadda_pg_rca24_and_1_3;
  assign s_dadda_pg_rca24_fa400_and1 = s_dadda_pg_rca24_fa400_xor0 & s_dadda_pg_rca24_and_1_3;
  assign s_dadda_pg_rca24_fa400_or0 = s_dadda_pg_rca24_fa400_and0 | s_dadda_pg_rca24_fa400_and1;
  assign s_dadda_pg_rca24_and_1_4 = a[1] & b[4];
  assign s_dadda_pg_rca24_and_0_5 = a[0] & b[5];
  assign s_dadda_pg_rca24_fa401_xor0 = s_dadda_pg_rca24_fa400_or0 ^ s_dadda_pg_rca24_and_1_4;
  assign s_dadda_pg_rca24_fa401_and0 = s_dadda_pg_rca24_fa400_or0 & s_dadda_pg_rca24_and_1_4;
  assign s_dadda_pg_rca24_fa401_xor1 = s_dadda_pg_rca24_fa401_xor0 ^ s_dadda_pg_rca24_and_0_5;
  assign s_dadda_pg_rca24_fa401_and1 = s_dadda_pg_rca24_fa401_xor0 & s_dadda_pg_rca24_and_0_5;
  assign s_dadda_pg_rca24_fa401_or0 = s_dadda_pg_rca24_fa401_and0 | s_dadda_pg_rca24_fa401_and1;
  assign s_dadda_pg_rca24_and_0_6 = a[0] & b[6];
  assign s_dadda_pg_rca24_fa402_xor0 = s_dadda_pg_rca24_fa401_or0 ^ s_dadda_pg_rca24_and_0_6;
  assign s_dadda_pg_rca24_fa402_and0 = s_dadda_pg_rca24_fa401_or0 & s_dadda_pg_rca24_and_0_6;
  assign s_dadda_pg_rca24_fa402_xor1 = s_dadda_pg_rca24_fa402_xor0 ^ s_dadda_pg_rca24_ha5_xor0;
  assign s_dadda_pg_rca24_fa402_and1 = s_dadda_pg_rca24_fa402_xor0 & s_dadda_pg_rca24_ha5_xor0;
  assign s_dadda_pg_rca24_fa402_or0 = s_dadda_pg_rca24_fa402_and0 | s_dadda_pg_rca24_fa402_and1;
  assign s_dadda_pg_rca24_fa403_xor0 = s_dadda_pg_rca24_fa402_or0 ^ s_dadda_pg_rca24_fa25_xor1;
  assign s_dadda_pg_rca24_fa403_and0 = s_dadda_pg_rca24_fa402_or0 & s_dadda_pg_rca24_fa25_xor1;
  assign s_dadda_pg_rca24_fa403_xor1 = s_dadda_pg_rca24_fa403_xor0 ^ s_dadda_pg_rca24_ha6_xor0;
  assign s_dadda_pg_rca24_fa403_and1 = s_dadda_pg_rca24_fa403_xor0 & s_dadda_pg_rca24_ha6_xor0;
  assign s_dadda_pg_rca24_fa403_or0 = s_dadda_pg_rca24_fa403_and0 | s_dadda_pg_rca24_fa403_and1;
  assign s_dadda_pg_rca24_fa404_xor0 = s_dadda_pg_rca24_fa403_or0 ^ s_dadda_pg_rca24_fa27_xor1;
  assign s_dadda_pg_rca24_fa404_and0 = s_dadda_pg_rca24_fa403_or0 & s_dadda_pg_rca24_fa27_xor1;
  assign s_dadda_pg_rca24_fa404_xor1 = s_dadda_pg_rca24_fa404_xor0 ^ s_dadda_pg_rca24_ha7_xor0;
  assign s_dadda_pg_rca24_fa404_and1 = s_dadda_pg_rca24_fa404_xor0 & s_dadda_pg_rca24_ha7_xor0;
  assign s_dadda_pg_rca24_fa404_or0 = s_dadda_pg_rca24_fa404_and0 | s_dadda_pg_rca24_fa404_and1;
  assign s_dadda_pg_rca24_fa405_xor0 = s_dadda_pg_rca24_fa404_or0 ^ s_dadda_pg_rca24_fa30_xor1;
  assign s_dadda_pg_rca24_fa405_and0 = s_dadda_pg_rca24_fa404_or0 & s_dadda_pg_rca24_fa30_xor1;
  assign s_dadda_pg_rca24_fa405_xor1 = s_dadda_pg_rca24_fa405_xor0 ^ s_dadda_pg_rca24_ha8_xor0;
  assign s_dadda_pg_rca24_fa405_and1 = s_dadda_pg_rca24_fa405_xor0 & s_dadda_pg_rca24_ha8_xor0;
  assign s_dadda_pg_rca24_fa405_or0 = s_dadda_pg_rca24_fa405_and0 | s_dadda_pg_rca24_fa405_and1;
  assign s_dadda_pg_rca24_fa406_xor0 = s_dadda_pg_rca24_fa405_or0 ^ s_dadda_pg_rca24_fa34_xor1;
  assign s_dadda_pg_rca24_fa406_and0 = s_dadda_pg_rca24_fa405_or0 & s_dadda_pg_rca24_fa34_xor1;
  assign s_dadda_pg_rca24_fa406_xor1 = s_dadda_pg_rca24_fa406_xor0 ^ s_dadda_pg_rca24_ha9_xor0;
  assign s_dadda_pg_rca24_fa406_and1 = s_dadda_pg_rca24_fa406_xor0 & s_dadda_pg_rca24_ha9_xor0;
  assign s_dadda_pg_rca24_fa406_or0 = s_dadda_pg_rca24_fa406_and0 | s_dadda_pg_rca24_fa406_and1;
  assign s_dadda_pg_rca24_fa407_xor0 = s_dadda_pg_rca24_fa406_or0 ^ s_dadda_pg_rca24_fa39_xor1;
  assign s_dadda_pg_rca24_fa407_and0 = s_dadda_pg_rca24_fa406_or0 & s_dadda_pg_rca24_fa39_xor1;
  assign s_dadda_pg_rca24_fa407_xor1 = s_dadda_pg_rca24_fa407_xor0 ^ s_dadda_pg_rca24_ha10_xor0;
  assign s_dadda_pg_rca24_fa407_and1 = s_dadda_pg_rca24_fa407_xor0 & s_dadda_pg_rca24_ha10_xor0;
  assign s_dadda_pg_rca24_fa407_or0 = s_dadda_pg_rca24_fa407_and0 | s_dadda_pg_rca24_fa407_and1;
  assign s_dadda_pg_rca24_fa408_xor0 = s_dadda_pg_rca24_fa407_or0 ^ s_dadda_pg_rca24_fa45_xor1;
  assign s_dadda_pg_rca24_fa408_and0 = s_dadda_pg_rca24_fa407_or0 & s_dadda_pg_rca24_fa45_xor1;
  assign s_dadda_pg_rca24_fa408_xor1 = s_dadda_pg_rca24_fa408_xor0 ^ s_dadda_pg_rca24_ha11_xor0;
  assign s_dadda_pg_rca24_fa408_and1 = s_dadda_pg_rca24_fa408_xor0 & s_dadda_pg_rca24_ha11_xor0;
  assign s_dadda_pg_rca24_fa408_or0 = s_dadda_pg_rca24_fa408_and0 | s_dadda_pg_rca24_fa408_and1;
  assign s_dadda_pg_rca24_fa409_xor0 = s_dadda_pg_rca24_fa408_or0 ^ s_dadda_pg_rca24_fa52_xor1;
  assign s_dadda_pg_rca24_fa409_and0 = s_dadda_pg_rca24_fa408_or0 & s_dadda_pg_rca24_fa52_xor1;
  assign s_dadda_pg_rca24_fa409_xor1 = s_dadda_pg_rca24_fa409_xor0 ^ s_dadda_pg_rca24_ha12_xor0;
  assign s_dadda_pg_rca24_fa409_and1 = s_dadda_pg_rca24_fa409_xor0 & s_dadda_pg_rca24_ha12_xor0;
  assign s_dadda_pg_rca24_fa409_or0 = s_dadda_pg_rca24_fa409_and0 | s_dadda_pg_rca24_fa409_and1;
  assign s_dadda_pg_rca24_fa410_xor0 = s_dadda_pg_rca24_fa409_or0 ^ s_dadda_pg_rca24_fa60_xor1;
  assign s_dadda_pg_rca24_fa410_and0 = s_dadda_pg_rca24_fa409_or0 & s_dadda_pg_rca24_fa60_xor1;
  assign s_dadda_pg_rca24_fa410_xor1 = s_dadda_pg_rca24_fa410_xor0 ^ s_dadda_pg_rca24_ha13_xor0;
  assign s_dadda_pg_rca24_fa410_and1 = s_dadda_pg_rca24_fa410_xor0 & s_dadda_pg_rca24_ha13_xor0;
  assign s_dadda_pg_rca24_fa410_or0 = s_dadda_pg_rca24_fa410_and0 | s_dadda_pg_rca24_fa410_and1;
  assign s_dadda_pg_rca24_fa411_xor0 = s_dadda_pg_rca24_fa410_or0 ^ s_dadda_pg_rca24_fa69_xor1;
  assign s_dadda_pg_rca24_fa411_and0 = s_dadda_pg_rca24_fa410_or0 & s_dadda_pg_rca24_fa69_xor1;
  assign s_dadda_pg_rca24_fa411_xor1 = s_dadda_pg_rca24_fa411_xor0 ^ s_dadda_pg_rca24_ha14_xor0;
  assign s_dadda_pg_rca24_fa411_and1 = s_dadda_pg_rca24_fa411_xor0 & s_dadda_pg_rca24_ha14_xor0;
  assign s_dadda_pg_rca24_fa411_or0 = s_dadda_pg_rca24_fa411_and0 | s_dadda_pg_rca24_fa411_and1;
  assign s_dadda_pg_rca24_fa412_xor0 = s_dadda_pg_rca24_fa411_or0 ^ s_dadda_pg_rca24_fa79_xor1;
  assign s_dadda_pg_rca24_fa412_and0 = s_dadda_pg_rca24_fa411_or0 & s_dadda_pg_rca24_fa79_xor1;
  assign s_dadda_pg_rca24_fa412_xor1 = s_dadda_pg_rca24_fa412_xor0 ^ s_dadda_pg_rca24_ha15_xor0;
  assign s_dadda_pg_rca24_fa412_and1 = s_dadda_pg_rca24_fa412_xor0 & s_dadda_pg_rca24_ha15_xor0;
  assign s_dadda_pg_rca24_fa412_or0 = s_dadda_pg_rca24_fa412_and0 | s_dadda_pg_rca24_fa412_and1;
  assign s_dadda_pg_rca24_fa413_xor0 = s_dadda_pg_rca24_fa412_or0 ^ s_dadda_pg_rca24_fa90_xor1;
  assign s_dadda_pg_rca24_fa413_and0 = s_dadda_pg_rca24_fa412_or0 & s_dadda_pg_rca24_fa90_xor1;
  assign s_dadda_pg_rca24_fa413_xor1 = s_dadda_pg_rca24_fa413_xor0 ^ s_dadda_pg_rca24_ha16_xor0;
  assign s_dadda_pg_rca24_fa413_and1 = s_dadda_pg_rca24_fa413_xor0 & s_dadda_pg_rca24_ha16_xor0;
  assign s_dadda_pg_rca24_fa413_or0 = s_dadda_pg_rca24_fa413_and0 | s_dadda_pg_rca24_fa413_and1;
  assign s_dadda_pg_rca24_fa414_xor0 = s_dadda_pg_rca24_fa413_or0 ^ s_dadda_pg_rca24_fa102_xor1;
  assign s_dadda_pg_rca24_fa414_and0 = s_dadda_pg_rca24_fa413_or0 & s_dadda_pg_rca24_fa102_xor1;
  assign s_dadda_pg_rca24_fa414_xor1 = s_dadda_pg_rca24_fa414_xor0 ^ s_dadda_pg_rca24_ha17_xor0;
  assign s_dadda_pg_rca24_fa414_and1 = s_dadda_pg_rca24_fa414_xor0 & s_dadda_pg_rca24_ha17_xor0;
  assign s_dadda_pg_rca24_fa414_or0 = s_dadda_pg_rca24_fa414_and0 | s_dadda_pg_rca24_fa414_and1;
  assign s_dadda_pg_rca24_fa415_xor0 = s_dadda_pg_rca24_fa414_or0 ^ s_dadda_pg_rca24_fa114_xor1;
  assign s_dadda_pg_rca24_fa415_and0 = s_dadda_pg_rca24_fa414_or0 & s_dadda_pg_rca24_fa114_xor1;
  assign s_dadda_pg_rca24_fa415_xor1 = s_dadda_pg_rca24_fa415_xor0 ^ s_dadda_pg_rca24_fa115_xor1;
  assign s_dadda_pg_rca24_fa415_and1 = s_dadda_pg_rca24_fa415_xor0 & s_dadda_pg_rca24_fa115_xor1;
  assign s_dadda_pg_rca24_fa415_or0 = s_dadda_pg_rca24_fa415_and0 | s_dadda_pg_rca24_fa415_and1;
  assign s_dadda_pg_rca24_fa416_xor0 = s_dadda_pg_rca24_fa415_or0 ^ s_dadda_pg_rca24_fa127_xor1;
  assign s_dadda_pg_rca24_fa416_and0 = s_dadda_pg_rca24_fa415_or0 & s_dadda_pg_rca24_fa127_xor1;
  assign s_dadda_pg_rca24_fa416_xor1 = s_dadda_pg_rca24_fa416_xor0 ^ s_dadda_pg_rca24_fa128_xor1;
  assign s_dadda_pg_rca24_fa416_and1 = s_dadda_pg_rca24_fa416_xor0 & s_dadda_pg_rca24_fa128_xor1;
  assign s_dadda_pg_rca24_fa416_or0 = s_dadda_pg_rca24_fa416_and0 | s_dadda_pg_rca24_fa416_and1;
  assign s_dadda_pg_rca24_fa417_xor0 = s_dadda_pg_rca24_fa416_or0 ^ s_dadda_pg_rca24_fa140_xor1;
  assign s_dadda_pg_rca24_fa417_and0 = s_dadda_pg_rca24_fa416_or0 & s_dadda_pg_rca24_fa140_xor1;
  assign s_dadda_pg_rca24_fa417_xor1 = s_dadda_pg_rca24_fa417_xor0 ^ s_dadda_pg_rca24_fa141_xor1;
  assign s_dadda_pg_rca24_fa417_and1 = s_dadda_pg_rca24_fa417_xor0 & s_dadda_pg_rca24_fa141_xor1;
  assign s_dadda_pg_rca24_fa417_or0 = s_dadda_pg_rca24_fa417_and0 | s_dadda_pg_rca24_fa417_and1;
  assign s_dadda_pg_rca24_fa418_xor0 = s_dadda_pg_rca24_fa417_or0 ^ s_dadda_pg_rca24_fa153_xor1;
  assign s_dadda_pg_rca24_fa418_and0 = s_dadda_pg_rca24_fa417_or0 & s_dadda_pg_rca24_fa153_xor1;
  assign s_dadda_pg_rca24_fa418_xor1 = s_dadda_pg_rca24_fa418_xor0 ^ s_dadda_pg_rca24_fa154_xor1;
  assign s_dadda_pg_rca24_fa418_and1 = s_dadda_pg_rca24_fa418_xor0 & s_dadda_pg_rca24_fa154_xor1;
  assign s_dadda_pg_rca24_fa418_or0 = s_dadda_pg_rca24_fa418_and0 | s_dadda_pg_rca24_fa418_and1;
  assign s_dadda_pg_rca24_fa419_xor0 = s_dadda_pg_rca24_fa418_or0 ^ s_dadda_pg_rca24_fa166_xor1;
  assign s_dadda_pg_rca24_fa419_and0 = s_dadda_pg_rca24_fa418_or0 & s_dadda_pg_rca24_fa166_xor1;
  assign s_dadda_pg_rca24_fa419_xor1 = s_dadda_pg_rca24_fa419_xor0 ^ s_dadda_pg_rca24_fa167_xor1;
  assign s_dadda_pg_rca24_fa419_and1 = s_dadda_pg_rca24_fa419_xor0 & s_dadda_pg_rca24_fa167_xor1;
  assign s_dadda_pg_rca24_fa419_or0 = s_dadda_pg_rca24_fa419_and0 | s_dadda_pg_rca24_fa419_and1;
  assign s_dadda_pg_rca24_fa420_xor0 = s_dadda_pg_rca24_fa419_or0 ^ s_dadda_pg_rca24_fa179_xor1;
  assign s_dadda_pg_rca24_fa420_and0 = s_dadda_pg_rca24_fa419_or0 & s_dadda_pg_rca24_fa179_xor1;
  assign s_dadda_pg_rca24_fa420_xor1 = s_dadda_pg_rca24_fa420_xor0 ^ s_dadda_pg_rca24_fa180_xor1;
  assign s_dadda_pg_rca24_fa420_and1 = s_dadda_pg_rca24_fa420_xor0 & s_dadda_pg_rca24_fa180_xor1;
  assign s_dadda_pg_rca24_fa420_or0 = s_dadda_pg_rca24_fa420_and0 | s_dadda_pg_rca24_fa420_and1;
  assign s_dadda_pg_rca24_fa421_xor0 = s_dadda_pg_rca24_fa420_or0 ^ s_dadda_pg_rca24_fa192_xor1;
  assign s_dadda_pg_rca24_fa421_and0 = s_dadda_pg_rca24_fa420_or0 & s_dadda_pg_rca24_fa192_xor1;
  assign s_dadda_pg_rca24_fa421_xor1 = s_dadda_pg_rca24_fa421_xor0 ^ s_dadda_pg_rca24_fa193_xor1;
  assign s_dadda_pg_rca24_fa421_and1 = s_dadda_pg_rca24_fa421_xor0 & s_dadda_pg_rca24_fa193_xor1;
  assign s_dadda_pg_rca24_fa421_or0 = s_dadda_pg_rca24_fa421_and0 | s_dadda_pg_rca24_fa421_and1;
  assign s_dadda_pg_rca24_fa422_xor0 = s_dadda_pg_rca24_fa421_or0 ^ s_dadda_pg_rca24_fa205_xor1;
  assign s_dadda_pg_rca24_fa422_and0 = s_dadda_pg_rca24_fa421_or0 & s_dadda_pg_rca24_fa205_xor1;
  assign s_dadda_pg_rca24_fa422_xor1 = s_dadda_pg_rca24_fa422_xor0 ^ s_dadda_pg_rca24_fa206_xor1;
  assign s_dadda_pg_rca24_fa422_and1 = s_dadda_pg_rca24_fa422_xor0 & s_dadda_pg_rca24_fa206_xor1;
  assign s_dadda_pg_rca24_fa422_or0 = s_dadda_pg_rca24_fa422_and0 | s_dadda_pg_rca24_fa422_and1;
  assign s_dadda_pg_rca24_fa423_xor0 = s_dadda_pg_rca24_fa422_or0 ^ s_dadda_pg_rca24_fa218_xor1;
  assign s_dadda_pg_rca24_fa423_and0 = s_dadda_pg_rca24_fa422_or0 & s_dadda_pg_rca24_fa218_xor1;
  assign s_dadda_pg_rca24_fa423_xor1 = s_dadda_pg_rca24_fa423_xor0 ^ s_dadda_pg_rca24_fa219_xor1;
  assign s_dadda_pg_rca24_fa423_and1 = s_dadda_pg_rca24_fa423_xor0 & s_dadda_pg_rca24_fa219_xor1;
  assign s_dadda_pg_rca24_fa423_or0 = s_dadda_pg_rca24_fa423_and0 | s_dadda_pg_rca24_fa423_and1;
  assign s_dadda_pg_rca24_fa424_xor0 = s_dadda_pg_rca24_fa423_or0 ^ s_dadda_pg_rca24_fa231_xor1;
  assign s_dadda_pg_rca24_fa424_and0 = s_dadda_pg_rca24_fa423_or0 & s_dadda_pg_rca24_fa231_xor1;
  assign s_dadda_pg_rca24_fa424_xor1 = s_dadda_pg_rca24_fa424_xor0 ^ s_dadda_pg_rca24_fa232_xor1;
  assign s_dadda_pg_rca24_fa424_and1 = s_dadda_pg_rca24_fa424_xor0 & s_dadda_pg_rca24_fa232_xor1;
  assign s_dadda_pg_rca24_fa424_or0 = s_dadda_pg_rca24_fa424_and0 | s_dadda_pg_rca24_fa424_and1;
  assign s_dadda_pg_rca24_fa425_xor0 = s_dadda_pg_rca24_fa424_or0 ^ s_dadda_pg_rca24_fa244_xor1;
  assign s_dadda_pg_rca24_fa425_and0 = s_dadda_pg_rca24_fa424_or0 & s_dadda_pg_rca24_fa244_xor1;
  assign s_dadda_pg_rca24_fa425_xor1 = s_dadda_pg_rca24_fa425_xor0 ^ s_dadda_pg_rca24_fa245_xor1;
  assign s_dadda_pg_rca24_fa425_and1 = s_dadda_pg_rca24_fa425_xor0 & s_dadda_pg_rca24_fa245_xor1;
  assign s_dadda_pg_rca24_fa425_or0 = s_dadda_pg_rca24_fa425_and0 | s_dadda_pg_rca24_fa425_and1;
  assign s_dadda_pg_rca24_fa426_xor0 = s_dadda_pg_rca24_fa425_or0 ^ s_dadda_pg_rca24_fa256_xor1;
  assign s_dadda_pg_rca24_fa426_and0 = s_dadda_pg_rca24_fa425_or0 & s_dadda_pg_rca24_fa256_xor1;
  assign s_dadda_pg_rca24_fa426_xor1 = s_dadda_pg_rca24_fa426_xor0 ^ s_dadda_pg_rca24_fa257_xor1;
  assign s_dadda_pg_rca24_fa426_and1 = s_dadda_pg_rca24_fa426_xor0 & s_dadda_pg_rca24_fa257_xor1;
  assign s_dadda_pg_rca24_fa426_or0 = s_dadda_pg_rca24_fa426_and0 | s_dadda_pg_rca24_fa426_and1;
  assign s_dadda_pg_rca24_fa427_xor0 = s_dadda_pg_rca24_fa426_or0 ^ s_dadda_pg_rca24_fa267_xor1;
  assign s_dadda_pg_rca24_fa427_and0 = s_dadda_pg_rca24_fa426_or0 & s_dadda_pg_rca24_fa267_xor1;
  assign s_dadda_pg_rca24_fa427_xor1 = s_dadda_pg_rca24_fa427_xor0 ^ s_dadda_pg_rca24_fa268_xor1;
  assign s_dadda_pg_rca24_fa427_and1 = s_dadda_pg_rca24_fa427_xor0 & s_dadda_pg_rca24_fa268_xor1;
  assign s_dadda_pg_rca24_fa427_or0 = s_dadda_pg_rca24_fa427_and0 | s_dadda_pg_rca24_fa427_and1;
  assign s_dadda_pg_rca24_fa428_xor0 = s_dadda_pg_rca24_fa427_or0 ^ s_dadda_pg_rca24_fa277_xor1;
  assign s_dadda_pg_rca24_fa428_and0 = s_dadda_pg_rca24_fa427_or0 & s_dadda_pg_rca24_fa277_xor1;
  assign s_dadda_pg_rca24_fa428_xor1 = s_dadda_pg_rca24_fa428_xor0 ^ s_dadda_pg_rca24_fa278_xor1;
  assign s_dadda_pg_rca24_fa428_and1 = s_dadda_pg_rca24_fa428_xor0 & s_dadda_pg_rca24_fa278_xor1;
  assign s_dadda_pg_rca24_fa428_or0 = s_dadda_pg_rca24_fa428_and0 | s_dadda_pg_rca24_fa428_and1;
  assign s_dadda_pg_rca24_fa429_xor0 = s_dadda_pg_rca24_fa428_or0 ^ s_dadda_pg_rca24_fa286_xor1;
  assign s_dadda_pg_rca24_fa429_and0 = s_dadda_pg_rca24_fa428_or0 & s_dadda_pg_rca24_fa286_xor1;
  assign s_dadda_pg_rca24_fa429_xor1 = s_dadda_pg_rca24_fa429_xor0 ^ s_dadda_pg_rca24_fa287_xor1;
  assign s_dadda_pg_rca24_fa429_and1 = s_dadda_pg_rca24_fa429_xor0 & s_dadda_pg_rca24_fa287_xor1;
  assign s_dadda_pg_rca24_fa429_or0 = s_dadda_pg_rca24_fa429_and0 | s_dadda_pg_rca24_fa429_and1;
  assign s_dadda_pg_rca24_fa430_xor0 = s_dadda_pg_rca24_fa429_or0 ^ s_dadda_pg_rca24_fa294_xor1;
  assign s_dadda_pg_rca24_fa430_and0 = s_dadda_pg_rca24_fa429_or0 & s_dadda_pg_rca24_fa294_xor1;
  assign s_dadda_pg_rca24_fa430_xor1 = s_dadda_pg_rca24_fa430_xor0 ^ s_dadda_pg_rca24_fa295_xor1;
  assign s_dadda_pg_rca24_fa430_and1 = s_dadda_pg_rca24_fa430_xor0 & s_dadda_pg_rca24_fa295_xor1;
  assign s_dadda_pg_rca24_fa430_or0 = s_dadda_pg_rca24_fa430_and0 | s_dadda_pg_rca24_fa430_and1;
  assign s_dadda_pg_rca24_fa431_xor0 = s_dadda_pg_rca24_fa430_or0 ^ s_dadda_pg_rca24_fa301_xor1;
  assign s_dadda_pg_rca24_fa431_and0 = s_dadda_pg_rca24_fa430_or0 & s_dadda_pg_rca24_fa301_xor1;
  assign s_dadda_pg_rca24_fa431_xor1 = s_dadda_pg_rca24_fa431_xor0 ^ s_dadda_pg_rca24_fa302_xor1;
  assign s_dadda_pg_rca24_fa431_and1 = s_dadda_pg_rca24_fa431_xor0 & s_dadda_pg_rca24_fa302_xor1;
  assign s_dadda_pg_rca24_fa431_or0 = s_dadda_pg_rca24_fa431_and0 | s_dadda_pg_rca24_fa431_and1;
  assign s_dadda_pg_rca24_fa432_xor0 = s_dadda_pg_rca24_fa431_or0 ^ s_dadda_pg_rca24_fa307_xor1;
  assign s_dadda_pg_rca24_fa432_and0 = s_dadda_pg_rca24_fa431_or0 & s_dadda_pg_rca24_fa307_xor1;
  assign s_dadda_pg_rca24_fa432_xor1 = s_dadda_pg_rca24_fa432_xor0 ^ s_dadda_pg_rca24_fa308_xor1;
  assign s_dadda_pg_rca24_fa432_and1 = s_dadda_pg_rca24_fa432_xor0 & s_dadda_pg_rca24_fa308_xor1;
  assign s_dadda_pg_rca24_fa432_or0 = s_dadda_pg_rca24_fa432_and0 | s_dadda_pg_rca24_fa432_and1;
  assign s_dadda_pg_rca24_fa433_xor0 = s_dadda_pg_rca24_fa432_or0 ^ s_dadda_pg_rca24_fa312_xor1;
  assign s_dadda_pg_rca24_fa433_and0 = s_dadda_pg_rca24_fa432_or0 & s_dadda_pg_rca24_fa312_xor1;
  assign s_dadda_pg_rca24_fa433_xor1 = s_dadda_pg_rca24_fa433_xor0 ^ s_dadda_pg_rca24_fa313_xor1;
  assign s_dadda_pg_rca24_fa433_and1 = s_dadda_pg_rca24_fa433_xor0 & s_dadda_pg_rca24_fa313_xor1;
  assign s_dadda_pg_rca24_fa433_or0 = s_dadda_pg_rca24_fa433_and0 | s_dadda_pg_rca24_fa433_and1;
  assign s_dadda_pg_rca24_fa434_xor0 = s_dadda_pg_rca24_fa433_or0 ^ s_dadda_pg_rca24_fa316_xor1;
  assign s_dadda_pg_rca24_fa434_and0 = s_dadda_pg_rca24_fa433_or0 & s_dadda_pg_rca24_fa316_xor1;
  assign s_dadda_pg_rca24_fa434_xor1 = s_dadda_pg_rca24_fa434_xor0 ^ s_dadda_pg_rca24_fa317_xor1;
  assign s_dadda_pg_rca24_fa434_and1 = s_dadda_pg_rca24_fa434_xor0 & s_dadda_pg_rca24_fa317_xor1;
  assign s_dadda_pg_rca24_fa434_or0 = s_dadda_pg_rca24_fa434_and0 | s_dadda_pg_rca24_fa434_and1;
  assign s_dadda_pg_rca24_fa435_xor0 = s_dadda_pg_rca24_fa434_or0 ^ s_dadda_pg_rca24_fa319_xor1;
  assign s_dadda_pg_rca24_fa435_and0 = s_dadda_pg_rca24_fa434_or0 & s_dadda_pg_rca24_fa319_xor1;
  assign s_dadda_pg_rca24_fa435_xor1 = s_dadda_pg_rca24_fa435_xor0 ^ s_dadda_pg_rca24_fa320_xor1;
  assign s_dadda_pg_rca24_fa435_and1 = s_dadda_pg_rca24_fa435_xor0 & s_dadda_pg_rca24_fa320_xor1;
  assign s_dadda_pg_rca24_fa435_or0 = s_dadda_pg_rca24_fa435_and0 | s_dadda_pg_rca24_fa435_and1;
  assign s_dadda_pg_rca24_fa436_xor0 = s_dadda_pg_rca24_fa435_or0 ^ s_dadda_pg_rca24_fa321_xor1;
  assign s_dadda_pg_rca24_fa436_and0 = s_dadda_pg_rca24_fa435_or0 & s_dadda_pg_rca24_fa321_xor1;
  assign s_dadda_pg_rca24_fa436_xor1 = s_dadda_pg_rca24_fa436_xor0 ^ s_dadda_pg_rca24_fa322_xor1;
  assign s_dadda_pg_rca24_fa436_and1 = s_dadda_pg_rca24_fa436_xor0 & s_dadda_pg_rca24_fa322_xor1;
  assign s_dadda_pg_rca24_fa436_or0 = s_dadda_pg_rca24_fa436_and0 | s_dadda_pg_rca24_fa436_and1;
  assign s_dadda_pg_rca24_nand_18_23 = ~(a[18] & b[23]);
  assign s_dadda_pg_rca24_fa437_xor0 = s_dadda_pg_rca24_fa436_or0 ^ s_dadda_pg_rca24_nand_18_23;
  assign s_dadda_pg_rca24_fa437_and0 = s_dadda_pg_rca24_fa436_or0 & s_dadda_pg_rca24_nand_18_23;
  assign s_dadda_pg_rca24_fa437_xor1 = s_dadda_pg_rca24_fa437_xor0 ^ s_dadda_pg_rca24_fa323_xor1;
  assign s_dadda_pg_rca24_fa437_and1 = s_dadda_pg_rca24_fa437_xor0 & s_dadda_pg_rca24_fa323_xor1;
  assign s_dadda_pg_rca24_fa437_or0 = s_dadda_pg_rca24_fa437_and0 | s_dadda_pg_rca24_fa437_and1;
  assign s_dadda_pg_rca24_and_20_22 = a[20] & b[22];
  assign s_dadda_pg_rca24_nand_19_23 = ~(a[19] & b[23]);
  assign s_dadda_pg_rca24_fa438_xor0 = s_dadda_pg_rca24_fa437_or0 ^ s_dadda_pg_rca24_and_20_22;
  assign s_dadda_pg_rca24_fa438_and0 = s_dadda_pg_rca24_fa437_or0 & s_dadda_pg_rca24_and_20_22;
  assign s_dadda_pg_rca24_fa438_xor1 = s_dadda_pg_rca24_fa438_xor0 ^ s_dadda_pg_rca24_nand_19_23;
  assign s_dadda_pg_rca24_fa438_and1 = s_dadda_pg_rca24_fa438_xor0 & s_dadda_pg_rca24_nand_19_23;
  assign s_dadda_pg_rca24_fa438_or0 = s_dadda_pg_rca24_fa438_and0 | s_dadda_pg_rca24_fa438_and1;
  assign s_dadda_pg_rca24_and_22_21 = a[22] & b[21];
  assign s_dadda_pg_rca24_and_21_22 = a[21] & b[22];
  assign s_dadda_pg_rca24_fa439_xor0 = s_dadda_pg_rca24_fa438_or0 ^ s_dadda_pg_rca24_and_22_21;
  assign s_dadda_pg_rca24_fa439_and0 = s_dadda_pg_rca24_fa438_or0 & s_dadda_pg_rca24_and_22_21;
  assign s_dadda_pg_rca24_fa439_xor1 = s_dadda_pg_rca24_fa439_xor0 ^ s_dadda_pg_rca24_and_21_22;
  assign s_dadda_pg_rca24_fa439_and1 = s_dadda_pg_rca24_fa439_xor0 & s_dadda_pg_rca24_and_21_22;
  assign s_dadda_pg_rca24_fa439_or0 = s_dadda_pg_rca24_fa439_and0 | s_dadda_pg_rca24_fa439_and1;
  assign s_dadda_pg_rca24_nand_23_21 = ~(a[23] & b[21]);
  assign s_dadda_pg_rca24_fa440_xor0 = s_dadda_pg_rca24_fa439_or0 ^ s_dadda_pg_rca24_fa399_or0;
  assign s_dadda_pg_rca24_fa440_and0 = s_dadda_pg_rca24_fa439_or0 & s_dadda_pg_rca24_fa399_or0;
  assign s_dadda_pg_rca24_fa440_xor1 = s_dadda_pg_rca24_fa440_xor0 ^ s_dadda_pg_rca24_nand_23_21;
  assign s_dadda_pg_rca24_fa440_and1 = s_dadda_pg_rca24_fa440_xor0 & s_dadda_pg_rca24_nand_23_21;
  assign s_dadda_pg_rca24_fa440_or0 = s_dadda_pg_rca24_fa440_and0 | s_dadda_pg_rca24_fa440_and1;
  assign s_dadda_pg_rca24_and_2_0 = a[2] & b[0];
  assign s_dadda_pg_rca24_and_1_1 = a[1] & b[1];
  assign s_dadda_pg_rca24_ha21_xor0 = s_dadda_pg_rca24_and_2_0 ^ s_dadda_pg_rca24_and_1_1;
  assign s_dadda_pg_rca24_ha21_and0 = s_dadda_pg_rca24_and_2_0 & s_dadda_pg_rca24_and_1_1;
  assign s_dadda_pg_rca24_and_1_2 = a[1] & b[2];
  assign s_dadda_pg_rca24_and_0_3 = a[0] & b[3];
  assign s_dadda_pg_rca24_fa441_xor0 = s_dadda_pg_rca24_ha21_and0 ^ s_dadda_pg_rca24_and_1_2;
  assign s_dadda_pg_rca24_fa441_and0 = s_dadda_pg_rca24_ha21_and0 & s_dadda_pg_rca24_and_1_2;
  assign s_dadda_pg_rca24_fa441_xor1 = s_dadda_pg_rca24_fa441_xor0 ^ s_dadda_pg_rca24_and_0_3;
  assign s_dadda_pg_rca24_fa441_and1 = s_dadda_pg_rca24_fa441_xor0 & s_dadda_pg_rca24_and_0_3;
  assign s_dadda_pg_rca24_fa441_or0 = s_dadda_pg_rca24_fa441_and0 | s_dadda_pg_rca24_fa441_and1;
  assign s_dadda_pg_rca24_and_0_4 = a[0] & b[4];
  assign s_dadda_pg_rca24_fa442_xor0 = s_dadda_pg_rca24_fa441_or0 ^ s_dadda_pg_rca24_and_0_4;
  assign s_dadda_pg_rca24_fa442_and0 = s_dadda_pg_rca24_fa441_or0 & s_dadda_pg_rca24_and_0_4;
  assign s_dadda_pg_rca24_fa442_xor1 = s_dadda_pg_rca24_fa442_xor0 ^ s_dadda_pg_rca24_ha18_xor0;
  assign s_dadda_pg_rca24_fa442_and1 = s_dadda_pg_rca24_fa442_xor0 & s_dadda_pg_rca24_ha18_xor0;
  assign s_dadda_pg_rca24_fa442_or0 = s_dadda_pg_rca24_fa442_and0 | s_dadda_pg_rca24_fa442_and1;
  assign s_dadda_pg_rca24_fa443_xor0 = s_dadda_pg_rca24_fa442_or0 ^ s_dadda_pg_rca24_fa324_xor1;
  assign s_dadda_pg_rca24_fa443_and0 = s_dadda_pg_rca24_fa442_or0 & s_dadda_pg_rca24_fa324_xor1;
  assign s_dadda_pg_rca24_fa443_xor1 = s_dadda_pg_rca24_fa443_xor0 ^ s_dadda_pg_rca24_ha19_xor0;
  assign s_dadda_pg_rca24_fa443_and1 = s_dadda_pg_rca24_fa443_xor0 & s_dadda_pg_rca24_ha19_xor0;
  assign s_dadda_pg_rca24_fa443_or0 = s_dadda_pg_rca24_fa443_and0 | s_dadda_pg_rca24_fa443_and1;
  assign s_dadda_pg_rca24_fa444_xor0 = s_dadda_pg_rca24_fa443_or0 ^ s_dadda_pg_rca24_fa325_xor1;
  assign s_dadda_pg_rca24_fa444_and0 = s_dadda_pg_rca24_fa443_or0 & s_dadda_pg_rca24_fa325_xor1;
  assign s_dadda_pg_rca24_fa444_xor1 = s_dadda_pg_rca24_fa444_xor0 ^ s_dadda_pg_rca24_fa326_xor1;
  assign s_dadda_pg_rca24_fa444_and1 = s_dadda_pg_rca24_fa444_xor0 & s_dadda_pg_rca24_fa326_xor1;
  assign s_dadda_pg_rca24_fa444_or0 = s_dadda_pg_rca24_fa444_and0 | s_dadda_pg_rca24_fa444_and1;
  assign s_dadda_pg_rca24_fa445_xor0 = s_dadda_pg_rca24_fa444_or0 ^ s_dadda_pg_rca24_fa327_xor1;
  assign s_dadda_pg_rca24_fa445_and0 = s_dadda_pg_rca24_fa444_or0 & s_dadda_pg_rca24_fa327_xor1;
  assign s_dadda_pg_rca24_fa445_xor1 = s_dadda_pg_rca24_fa445_xor0 ^ s_dadda_pg_rca24_fa328_xor1;
  assign s_dadda_pg_rca24_fa445_and1 = s_dadda_pg_rca24_fa445_xor0 & s_dadda_pg_rca24_fa328_xor1;
  assign s_dadda_pg_rca24_fa445_or0 = s_dadda_pg_rca24_fa445_and0 | s_dadda_pg_rca24_fa445_and1;
  assign s_dadda_pg_rca24_fa446_xor0 = s_dadda_pg_rca24_fa445_or0 ^ s_dadda_pg_rca24_fa329_xor1;
  assign s_dadda_pg_rca24_fa446_and0 = s_dadda_pg_rca24_fa445_or0 & s_dadda_pg_rca24_fa329_xor1;
  assign s_dadda_pg_rca24_fa446_xor1 = s_dadda_pg_rca24_fa446_xor0 ^ s_dadda_pg_rca24_fa330_xor1;
  assign s_dadda_pg_rca24_fa446_and1 = s_dadda_pg_rca24_fa446_xor0 & s_dadda_pg_rca24_fa330_xor1;
  assign s_dadda_pg_rca24_fa446_or0 = s_dadda_pg_rca24_fa446_and0 | s_dadda_pg_rca24_fa446_and1;
  assign s_dadda_pg_rca24_fa447_xor0 = s_dadda_pg_rca24_fa446_or0 ^ s_dadda_pg_rca24_fa331_xor1;
  assign s_dadda_pg_rca24_fa447_and0 = s_dadda_pg_rca24_fa446_or0 & s_dadda_pg_rca24_fa331_xor1;
  assign s_dadda_pg_rca24_fa447_xor1 = s_dadda_pg_rca24_fa447_xor0 ^ s_dadda_pg_rca24_fa332_xor1;
  assign s_dadda_pg_rca24_fa447_and1 = s_dadda_pg_rca24_fa447_xor0 & s_dadda_pg_rca24_fa332_xor1;
  assign s_dadda_pg_rca24_fa447_or0 = s_dadda_pg_rca24_fa447_and0 | s_dadda_pg_rca24_fa447_and1;
  assign s_dadda_pg_rca24_fa448_xor0 = s_dadda_pg_rca24_fa447_or0 ^ s_dadda_pg_rca24_fa333_xor1;
  assign s_dadda_pg_rca24_fa448_and0 = s_dadda_pg_rca24_fa447_or0 & s_dadda_pg_rca24_fa333_xor1;
  assign s_dadda_pg_rca24_fa448_xor1 = s_dadda_pg_rca24_fa448_xor0 ^ s_dadda_pg_rca24_fa334_xor1;
  assign s_dadda_pg_rca24_fa448_and1 = s_dadda_pg_rca24_fa448_xor0 & s_dadda_pg_rca24_fa334_xor1;
  assign s_dadda_pg_rca24_fa448_or0 = s_dadda_pg_rca24_fa448_and0 | s_dadda_pg_rca24_fa448_and1;
  assign s_dadda_pg_rca24_fa449_xor0 = s_dadda_pg_rca24_fa448_or0 ^ s_dadda_pg_rca24_fa335_xor1;
  assign s_dadda_pg_rca24_fa449_and0 = s_dadda_pg_rca24_fa448_or0 & s_dadda_pg_rca24_fa335_xor1;
  assign s_dadda_pg_rca24_fa449_xor1 = s_dadda_pg_rca24_fa449_xor0 ^ s_dadda_pg_rca24_fa336_xor1;
  assign s_dadda_pg_rca24_fa449_and1 = s_dadda_pg_rca24_fa449_xor0 & s_dadda_pg_rca24_fa336_xor1;
  assign s_dadda_pg_rca24_fa449_or0 = s_dadda_pg_rca24_fa449_and0 | s_dadda_pg_rca24_fa449_and1;
  assign s_dadda_pg_rca24_fa450_xor0 = s_dadda_pg_rca24_fa449_or0 ^ s_dadda_pg_rca24_fa337_xor1;
  assign s_dadda_pg_rca24_fa450_and0 = s_dadda_pg_rca24_fa449_or0 & s_dadda_pg_rca24_fa337_xor1;
  assign s_dadda_pg_rca24_fa450_xor1 = s_dadda_pg_rca24_fa450_xor0 ^ s_dadda_pg_rca24_fa338_xor1;
  assign s_dadda_pg_rca24_fa450_and1 = s_dadda_pg_rca24_fa450_xor0 & s_dadda_pg_rca24_fa338_xor1;
  assign s_dadda_pg_rca24_fa450_or0 = s_dadda_pg_rca24_fa450_and0 | s_dadda_pg_rca24_fa450_and1;
  assign s_dadda_pg_rca24_fa451_xor0 = s_dadda_pg_rca24_fa450_or0 ^ s_dadda_pg_rca24_fa339_xor1;
  assign s_dadda_pg_rca24_fa451_and0 = s_dadda_pg_rca24_fa450_or0 & s_dadda_pg_rca24_fa339_xor1;
  assign s_dadda_pg_rca24_fa451_xor1 = s_dadda_pg_rca24_fa451_xor0 ^ s_dadda_pg_rca24_fa340_xor1;
  assign s_dadda_pg_rca24_fa451_and1 = s_dadda_pg_rca24_fa451_xor0 & s_dadda_pg_rca24_fa340_xor1;
  assign s_dadda_pg_rca24_fa451_or0 = s_dadda_pg_rca24_fa451_and0 | s_dadda_pg_rca24_fa451_and1;
  assign s_dadda_pg_rca24_fa452_xor0 = s_dadda_pg_rca24_fa451_or0 ^ s_dadda_pg_rca24_fa341_xor1;
  assign s_dadda_pg_rca24_fa452_and0 = s_dadda_pg_rca24_fa451_or0 & s_dadda_pg_rca24_fa341_xor1;
  assign s_dadda_pg_rca24_fa452_xor1 = s_dadda_pg_rca24_fa452_xor0 ^ s_dadda_pg_rca24_fa342_xor1;
  assign s_dadda_pg_rca24_fa452_and1 = s_dadda_pg_rca24_fa452_xor0 & s_dadda_pg_rca24_fa342_xor1;
  assign s_dadda_pg_rca24_fa452_or0 = s_dadda_pg_rca24_fa452_and0 | s_dadda_pg_rca24_fa452_and1;
  assign s_dadda_pg_rca24_fa453_xor0 = s_dadda_pg_rca24_fa452_or0 ^ s_dadda_pg_rca24_fa343_xor1;
  assign s_dadda_pg_rca24_fa453_and0 = s_dadda_pg_rca24_fa452_or0 & s_dadda_pg_rca24_fa343_xor1;
  assign s_dadda_pg_rca24_fa453_xor1 = s_dadda_pg_rca24_fa453_xor0 ^ s_dadda_pg_rca24_fa344_xor1;
  assign s_dadda_pg_rca24_fa453_and1 = s_dadda_pg_rca24_fa453_xor0 & s_dadda_pg_rca24_fa344_xor1;
  assign s_dadda_pg_rca24_fa453_or0 = s_dadda_pg_rca24_fa453_and0 | s_dadda_pg_rca24_fa453_and1;
  assign s_dadda_pg_rca24_fa454_xor0 = s_dadda_pg_rca24_fa453_or0 ^ s_dadda_pg_rca24_fa345_xor1;
  assign s_dadda_pg_rca24_fa454_and0 = s_dadda_pg_rca24_fa453_or0 & s_dadda_pg_rca24_fa345_xor1;
  assign s_dadda_pg_rca24_fa454_xor1 = s_dadda_pg_rca24_fa454_xor0 ^ s_dadda_pg_rca24_fa346_xor1;
  assign s_dadda_pg_rca24_fa454_and1 = s_dadda_pg_rca24_fa454_xor0 & s_dadda_pg_rca24_fa346_xor1;
  assign s_dadda_pg_rca24_fa454_or0 = s_dadda_pg_rca24_fa454_and0 | s_dadda_pg_rca24_fa454_and1;
  assign s_dadda_pg_rca24_fa455_xor0 = s_dadda_pg_rca24_fa454_or0 ^ s_dadda_pg_rca24_fa347_xor1;
  assign s_dadda_pg_rca24_fa455_and0 = s_dadda_pg_rca24_fa454_or0 & s_dadda_pg_rca24_fa347_xor1;
  assign s_dadda_pg_rca24_fa455_xor1 = s_dadda_pg_rca24_fa455_xor0 ^ s_dadda_pg_rca24_fa348_xor1;
  assign s_dadda_pg_rca24_fa455_and1 = s_dadda_pg_rca24_fa455_xor0 & s_dadda_pg_rca24_fa348_xor1;
  assign s_dadda_pg_rca24_fa455_or0 = s_dadda_pg_rca24_fa455_and0 | s_dadda_pg_rca24_fa455_and1;
  assign s_dadda_pg_rca24_fa456_xor0 = s_dadda_pg_rca24_fa455_or0 ^ s_dadda_pg_rca24_fa349_xor1;
  assign s_dadda_pg_rca24_fa456_and0 = s_dadda_pg_rca24_fa455_or0 & s_dadda_pg_rca24_fa349_xor1;
  assign s_dadda_pg_rca24_fa456_xor1 = s_dadda_pg_rca24_fa456_xor0 ^ s_dadda_pg_rca24_fa350_xor1;
  assign s_dadda_pg_rca24_fa456_and1 = s_dadda_pg_rca24_fa456_xor0 & s_dadda_pg_rca24_fa350_xor1;
  assign s_dadda_pg_rca24_fa456_or0 = s_dadda_pg_rca24_fa456_and0 | s_dadda_pg_rca24_fa456_and1;
  assign s_dadda_pg_rca24_fa457_xor0 = s_dadda_pg_rca24_fa456_or0 ^ s_dadda_pg_rca24_fa351_xor1;
  assign s_dadda_pg_rca24_fa457_and0 = s_dadda_pg_rca24_fa456_or0 & s_dadda_pg_rca24_fa351_xor1;
  assign s_dadda_pg_rca24_fa457_xor1 = s_dadda_pg_rca24_fa457_xor0 ^ s_dadda_pg_rca24_fa352_xor1;
  assign s_dadda_pg_rca24_fa457_and1 = s_dadda_pg_rca24_fa457_xor0 & s_dadda_pg_rca24_fa352_xor1;
  assign s_dadda_pg_rca24_fa457_or0 = s_dadda_pg_rca24_fa457_and0 | s_dadda_pg_rca24_fa457_and1;
  assign s_dadda_pg_rca24_fa458_xor0 = s_dadda_pg_rca24_fa457_or0 ^ s_dadda_pg_rca24_fa353_xor1;
  assign s_dadda_pg_rca24_fa458_and0 = s_dadda_pg_rca24_fa457_or0 & s_dadda_pg_rca24_fa353_xor1;
  assign s_dadda_pg_rca24_fa458_xor1 = s_dadda_pg_rca24_fa458_xor0 ^ s_dadda_pg_rca24_fa354_xor1;
  assign s_dadda_pg_rca24_fa458_and1 = s_dadda_pg_rca24_fa458_xor0 & s_dadda_pg_rca24_fa354_xor1;
  assign s_dadda_pg_rca24_fa458_or0 = s_dadda_pg_rca24_fa458_and0 | s_dadda_pg_rca24_fa458_and1;
  assign s_dadda_pg_rca24_fa459_xor0 = s_dadda_pg_rca24_fa458_or0 ^ s_dadda_pg_rca24_fa355_xor1;
  assign s_dadda_pg_rca24_fa459_and0 = s_dadda_pg_rca24_fa458_or0 & s_dadda_pg_rca24_fa355_xor1;
  assign s_dadda_pg_rca24_fa459_xor1 = s_dadda_pg_rca24_fa459_xor0 ^ s_dadda_pg_rca24_fa356_xor1;
  assign s_dadda_pg_rca24_fa459_and1 = s_dadda_pg_rca24_fa459_xor0 & s_dadda_pg_rca24_fa356_xor1;
  assign s_dadda_pg_rca24_fa459_or0 = s_dadda_pg_rca24_fa459_and0 | s_dadda_pg_rca24_fa459_and1;
  assign s_dadda_pg_rca24_fa460_xor0 = s_dadda_pg_rca24_fa459_or0 ^ s_dadda_pg_rca24_fa357_xor1;
  assign s_dadda_pg_rca24_fa460_and0 = s_dadda_pg_rca24_fa459_or0 & s_dadda_pg_rca24_fa357_xor1;
  assign s_dadda_pg_rca24_fa460_xor1 = s_dadda_pg_rca24_fa460_xor0 ^ s_dadda_pg_rca24_fa358_xor1;
  assign s_dadda_pg_rca24_fa460_and1 = s_dadda_pg_rca24_fa460_xor0 & s_dadda_pg_rca24_fa358_xor1;
  assign s_dadda_pg_rca24_fa460_or0 = s_dadda_pg_rca24_fa460_and0 | s_dadda_pg_rca24_fa460_and1;
  assign s_dadda_pg_rca24_fa461_xor0 = s_dadda_pg_rca24_fa460_or0 ^ s_dadda_pg_rca24_fa359_xor1;
  assign s_dadda_pg_rca24_fa461_and0 = s_dadda_pg_rca24_fa460_or0 & s_dadda_pg_rca24_fa359_xor1;
  assign s_dadda_pg_rca24_fa461_xor1 = s_dadda_pg_rca24_fa461_xor0 ^ s_dadda_pg_rca24_fa360_xor1;
  assign s_dadda_pg_rca24_fa461_and1 = s_dadda_pg_rca24_fa461_xor0 & s_dadda_pg_rca24_fa360_xor1;
  assign s_dadda_pg_rca24_fa461_or0 = s_dadda_pg_rca24_fa461_and0 | s_dadda_pg_rca24_fa461_and1;
  assign s_dadda_pg_rca24_fa462_xor0 = s_dadda_pg_rca24_fa461_or0 ^ s_dadda_pg_rca24_fa361_xor1;
  assign s_dadda_pg_rca24_fa462_and0 = s_dadda_pg_rca24_fa461_or0 & s_dadda_pg_rca24_fa361_xor1;
  assign s_dadda_pg_rca24_fa462_xor1 = s_dadda_pg_rca24_fa462_xor0 ^ s_dadda_pg_rca24_fa362_xor1;
  assign s_dadda_pg_rca24_fa462_and1 = s_dadda_pg_rca24_fa462_xor0 & s_dadda_pg_rca24_fa362_xor1;
  assign s_dadda_pg_rca24_fa462_or0 = s_dadda_pg_rca24_fa462_and0 | s_dadda_pg_rca24_fa462_and1;
  assign s_dadda_pg_rca24_fa463_xor0 = s_dadda_pg_rca24_fa462_or0 ^ s_dadda_pg_rca24_fa363_xor1;
  assign s_dadda_pg_rca24_fa463_and0 = s_dadda_pg_rca24_fa462_or0 & s_dadda_pg_rca24_fa363_xor1;
  assign s_dadda_pg_rca24_fa463_xor1 = s_dadda_pg_rca24_fa463_xor0 ^ s_dadda_pg_rca24_fa364_xor1;
  assign s_dadda_pg_rca24_fa463_and1 = s_dadda_pg_rca24_fa463_xor0 & s_dadda_pg_rca24_fa364_xor1;
  assign s_dadda_pg_rca24_fa463_or0 = s_dadda_pg_rca24_fa463_and0 | s_dadda_pg_rca24_fa463_and1;
  assign s_dadda_pg_rca24_fa464_xor0 = s_dadda_pg_rca24_fa463_or0 ^ s_dadda_pg_rca24_fa365_xor1;
  assign s_dadda_pg_rca24_fa464_and0 = s_dadda_pg_rca24_fa463_or0 & s_dadda_pg_rca24_fa365_xor1;
  assign s_dadda_pg_rca24_fa464_xor1 = s_dadda_pg_rca24_fa464_xor0 ^ s_dadda_pg_rca24_fa366_xor1;
  assign s_dadda_pg_rca24_fa464_and1 = s_dadda_pg_rca24_fa464_xor0 & s_dadda_pg_rca24_fa366_xor1;
  assign s_dadda_pg_rca24_fa464_or0 = s_dadda_pg_rca24_fa464_and0 | s_dadda_pg_rca24_fa464_and1;
  assign s_dadda_pg_rca24_fa465_xor0 = s_dadda_pg_rca24_fa464_or0 ^ s_dadda_pg_rca24_fa367_xor1;
  assign s_dadda_pg_rca24_fa465_and0 = s_dadda_pg_rca24_fa464_or0 & s_dadda_pg_rca24_fa367_xor1;
  assign s_dadda_pg_rca24_fa465_xor1 = s_dadda_pg_rca24_fa465_xor0 ^ s_dadda_pg_rca24_fa368_xor1;
  assign s_dadda_pg_rca24_fa465_and1 = s_dadda_pg_rca24_fa465_xor0 & s_dadda_pg_rca24_fa368_xor1;
  assign s_dadda_pg_rca24_fa465_or0 = s_dadda_pg_rca24_fa465_and0 | s_dadda_pg_rca24_fa465_and1;
  assign s_dadda_pg_rca24_fa466_xor0 = s_dadda_pg_rca24_fa465_or0 ^ s_dadda_pg_rca24_fa369_xor1;
  assign s_dadda_pg_rca24_fa466_and0 = s_dadda_pg_rca24_fa465_or0 & s_dadda_pg_rca24_fa369_xor1;
  assign s_dadda_pg_rca24_fa466_xor1 = s_dadda_pg_rca24_fa466_xor0 ^ s_dadda_pg_rca24_fa370_xor1;
  assign s_dadda_pg_rca24_fa466_and1 = s_dadda_pg_rca24_fa466_xor0 & s_dadda_pg_rca24_fa370_xor1;
  assign s_dadda_pg_rca24_fa466_or0 = s_dadda_pg_rca24_fa466_and0 | s_dadda_pg_rca24_fa466_and1;
  assign s_dadda_pg_rca24_fa467_xor0 = s_dadda_pg_rca24_fa466_or0 ^ s_dadda_pg_rca24_fa371_xor1;
  assign s_dadda_pg_rca24_fa467_and0 = s_dadda_pg_rca24_fa466_or0 & s_dadda_pg_rca24_fa371_xor1;
  assign s_dadda_pg_rca24_fa467_xor1 = s_dadda_pg_rca24_fa467_xor0 ^ s_dadda_pg_rca24_fa372_xor1;
  assign s_dadda_pg_rca24_fa467_and1 = s_dadda_pg_rca24_fa467_xor0 & s_dadda_pg_rca24_fa372_xor1;
  assign s_dadda_pg_rca24_fa467_or0 = s_dadda_pg_rca24_fa467_and0 | s_dadda_pg_rca24_fa467_and1;
  assign s_dadda_pg_rca24_fa468_xor0 = s_dadda_pg_rca24_fa467_or0 ^ s_dadda_pg_rca24_fa373_xor1;
  assign s_dadda_pg_rca24_fa468_and0 = s_dadda_pg_rca24_fa467_or0 & s_dadda_pg_rca24_fa373_xor1;
  assign s_dadda_pg_rca24_fa468_xor1 = s_dadda_pg_rca24_fa468_xor0 ^ s_dadda_pg_rca24_fa374_xor1;
  assign s_dadda_pg_rca24_fa468_and1 = s_dadda_pg_rca24_fa468_xor0 & s_dadda_pg_rca24_fa374_xor1;
  assign s_dadda_pg_rca24_fa468_or0 = s_dadda_pg_rca24_fa468_and0 | s_dadda_pg_rca24_fa468_and1;
  assign s_dadda_pg_rca24_fa469_xor0 = s_dadda_pg_rca24_fa468_or0 ^ s_dadda_pg_rca24_fa375_xor1;
  assign s_dadda_pg_rca24_fa469_and0 = s_dadda_pg_rca24_fa468_or0 & s_dadda_pg_rca24_fa375_xor1;
  assign s_dadda_pg_rca24_fa469_xor1 = s_dadda_pg_rca24_fa469_xor0 ^ s_dadda_pg_rca24_fa376_xor1;
  assign s_dadda_pg_rca24_fa469_and1 = s_dadda_pg_rca24_fa469_xor0 & s_dadda_pg_rca24_fa376_xor1;
  assign s_dadda_pg_rca24_fa469_or0 = s_dadda_pg_rca24_fa469_and0 | s_dadda_pg_rca24_fa469_and1;
  assign s_dadda_pg_rca24_fa470_xor0 = s_dadda_pg_rca24_fa469_or0 ^ s_dadda_pg_rca24_fa377_xor1;
  assign s_dadda_pg_rca24_fa470_and0 = s_dadda_pg_rca24_fa469_or0 & s_dadda_pg_rca24_fa377_xor1;
  assign s_dadda_pg_rca24_fa470_xor1 = s_dadda_pg_rca24_fa470_xor0 ^ s_dadda_pg_rca24_fa378_xor1;
  assign s_dadda_pg_rca24_fa470_and1 = s_dadda_pg_rca24_fa470_xor0 & s_dadda_pg_rca24_fa378_xor1;
  assign s_dadda_pg_rca24_fa470_or0 = s_dadda_pg_rca24_fa470_and0 | s_dadda_pg_rca24_fa470_and1;
  assign s_dadda_pg_rca24_fa471_xor0 = s_dadda_pg_rca24_fa470_or0 ^ s_dadda_pg_rca24_fa379_xor1;
  assign s_dadda_pg_rca24_fa471_and0 = s_dadda_pg_rca24_fa470_or0 & s_dadda_pg_rca24_fa379_xor1;
  assign s_dadda_pg_rca24_fa471_xor1 = s_dadda_pg_rca24_fa471_xor0 ^ s_dadda_pg_rca24_fa380_xor1;
  assign s_dadda_pg_rca24_fa471_and1 = s_dadda_pg_rca24_fa471_xor0 & s_dadda_pg_rca24_fa380_xor1;
  assign s_dadda_pg_rca24_fa471_or0 = s_dadda_pg_rca24_fa471_and0 | s_dadda_pg_rca24_fa471_and1;
  assign s_dadda_pg_rca24_fa472_xor0 = s_dadda_pg_rca24_fa471_or0 ^ s_dadda_pg_rca24_fa381_xor1;
  assign s_dadda_pg_rca24_fa472_and0 = s_dadda_pg_rca24_fa471_or0 & s_dadda_pg_rca24_fa381_xor1;
  assign s_dadda_pg_rca24_fa472_xor1 = s_dadda_pg_rca24_fa472_xor0 ^ s_dadda_pg_rca24_fa382_xor1;
  assign s_dadda_pg_rca24_fa472_and1 = s_dadda_pg_rca24_fa472_xor0 & s_dadda_pg_rca24_fa382_xor1;
  assign s_dadda_pg_rca24_fa472_or0 = s_dadda_pg_rca24_fa472_and0 | s_dadda_pg_rca24_fa472_and1;
  assign s_dadda_pg_rca24_fa473_xor0 = s_dadda_pg_rca24_fa472_or0 ^ s_dadda_pg_rca24_fa383_xor1;
  assign s_dadda_pg_rca24_fa473_and0 = s_dadda_pg_rca24_fa472_or0 & s_dadda_pg_rca24_fa383_xor1;
  assign s_dadda_pg_rca24_fa473_xor1 = s_dadda_pg_rca24_fa473_xor0 ^ s_dadda_pg_rca24_fa384_xor1;
  assign s_dadda_pg_rca24_fa473_and1 = s_dadda_pg_rca24_fa473_xor0 & s_dadda_pg_rca24_fa384_xor1;
  assign s_dadda_pg_rca24_fa473_or0 = s_dadda_pg_rca24_fa473_and0 | s_dadda_pg_rca24_fa473_and1;
  assign s_dadda_pg_rca24_fa474_xor0 = s_dadda_pg_rca24_fa473_or0 ^ s_dadda_pg_rca24_fa385_xor1;
  assign s_dadda_pg_rca24_fa474_and0 = s_dadda_pg_rca24_fa473_or0 & s_dadda_pg_rca24_fa385_xor1;
  assign s_dadda_pg_rca24_fa474_xor1 = s_dadda_pg_rca24_fa474_xor0 ^ s_dadda_pg_rca24_fa386_xor1;
  assign s_dadda_pg_rca24_fa474_and1 = s_dadda_pg_rca24_fa474_xor0 & s_dadda_pg_rca24_fa386_xor1;
  assign s_dadda_pg_rca24_fa474_or0 = s_dadda_pg_rca24_fa474_and0 | s_dadda_pg_rca24_fa474_and1;
  assign s_dadda_pg_rca24_fa475_xor0 = s_dadda_pg_rca24_fa474_or0 ^ s_dadda_pg_rca24_fa387_xor1;
  assign s_dadda_pg_rca24_fa475_and0 = s_dadda_pg_rca24_fa474_or0 & s_dadda_pg_rca24_fa387_xor1;
  assign s_dadda_pg_rca24_fa475_xor1 = s_dadda_pg_rca24_fa475_xor0 ^ s_dadda_pg_rca24_fa388_xor1;
  assign s_dadda_pg_rca24_fa475_and1 = s_dadda_pg_rca24_fa475_xor0 & s_dadda_pg_rca24_fa388_xor1;
  assign s_dadda_pg_rca24_fa475_or0 = s_dadda_pg_rca24_fa475_and0 | s_dadda_pg_rca24_fa475_and1;
  assign s_dadda_pg_rca24_fa476_xor0 = s_dadda_pg_rca24_fa475_or0 ^ s_dadda_pg_rca24_fa389_xor1;
  assign s_dadda_pg_rca24_fa476_and0 = s_dadda_pg_rca24_fa475_or0 & s_dadda_pg_rca24_fa389_xor1;
  assign s_dadda_pg_rca24_fa476_xor1 = s_dadda_pg_rca24_fa476_xor0 ^ s_dadda_pg_rca24_fa390_xor1;
  assign s_dadda_pg_rca24_fa476_and1 = s_dadda_pg_rca24_fa476_xor0 & s_dadda_pg_rca24_fa390_xor1;
  assign s_dadda_pg_rca24_fa476_or0 = s_dadda_pg_rca24_fa476_and0 | s_dadda_pg_rca24_fa476_and1;
  assign s_dadda_pg_rca24_fa477_xor0 = s_dadda_pg_rca24_fa476_or0 ^ s_dadda_pg_rca24_fa391_xor1;
  assign s_dadda_pg_rca24_fa477_and0 = s_dadda_pg_rca24_fa476_or0 & s_dadda_pg_rca24_fa391_xor1;
  assign s_dadda_pg_rca24_fa477_xor1 = s_dadda_pg_rca24_fa477_xor0 ^ s_dadda_pg_rca24_fa392_xor1;
  assign s_dadda_pg_rca24_fa477_and1 = s_dadda_pg_rca24_fa477_xor0 & s_dadda_pg_rca24_fa392_xor1;
  assign s_dadda_pg_rca24_fa477_or0 = s_dadda_pg_rca24_fa477_and0 | s_dadda_pg_rca24_fa477_and1;
  assign s_dadda_pg_rca24_fa478_xor0 = s_dadda_pg_rca24_fa477_or0 ^ s_dadda_pg_rca24_fa393_xor1;
  assign s_dadda_pg_rca24_fa478_and0 = s_dadda_pg_rca24_fa477_or0 & s_dadda_pg_rca24_fa393_xor1;
  assign s_dadda_pg_rca24_fa478_xor1 = s_dadda_pg_rca24_fa478_xor0 ^ s_dadda_pg_rca24_fa394_xor1;
  assign s_dadda_pg_rca24_fa478_and1 = s_dadda_pg_rca24_fa478_xor0 & s_dadda_pg_rca24_fa394_xor1;
  assign s_dadda_pg_rca24_fa478_or0 = s_dadda_pg_rca24_fa478_and0 | s_dadda_pg_rca24_fa478_and1;
  assign s_dadda_pg_rca24_fa479_xor0 = s_dadda_pg_rca24_fa478_or0 ^ s_dadda_pg_rca24_fa395_xor1;
  assign s_dadda_pg_rca24_fa479_and0 = s_dadda_pg_rca24_fa478_or0 & s_dadda_pg_rca24_fa395_xor1;
  assign s_dadda_pg_rca24_fa479_xor1 = s_dadda_pg_rca24_fa479_xor0 ^ s_dadda_pg_rca24_fa396_xor1;
  assign s_dadda_pg_rca24_fa479_and1 = s_dadda_pg_rca24_fa479_xor0 & s_dadda_pg_rca24_fa396_xor1;
  assign s_dadda_pg_rca24_fa479_or0 = s_dadda_pg_rca24_fa479_and0 | s_dadda_pg_rca24_fa479_and1;
  assign s_dadda_pg_rca24_fa480_xor0 = s_dadda_pg_rca24_fa479_or0 ^ s_dadda_pg_rca24_fa397_xor1;
  assign s_dadda_pg_rca24_fa480_and0 = s_dadda_pg_rca24_fa479_or0 & s_dadda_pg_rca24_fa397_xor1;
  assign s_dadda_pg_rca24_fa480_xor1 = s_dadda_pg_rca24_fa480_xor0 ^ s_dadda_pg_rca24_fa398_xor1;
  assign s_dadda_pg_rca24_fa480_and1 = s_dadda_pg_rca24_fa480_xor0 & s_dadda_pg_rca24_fa398_xor1;
  assign s_dadda_pg_rca24_fa480_or0 = s_dadda_pg_rca24_fa480_and0 | s_dadda_pg_rca24_fa480_and1;
  assign s_dadda_pg_rca24_nand_20_23 = ~(a[20] & b[23]);
  assign s_dadda_pg_rca24_fa481_xor0 = s_dadda_pg_rca24_fa480_or0 ^ s_dadda_pg_rca24_nand_20_23;
  assign s_dadda_pg_rca24_fa481_and0 = s_dadda_pg_rca24_fa480_or0 & s_dadda_pg_rca24_nand_20_23;
  assign s_dadda_pg_rca24_fa481_xor1 = s_dadda_pg_rca24_fa481_xor0 ^ s_dadda_pg_rca24_fa399_xor1;
  assign s_dadda_pg_rca24_fa481_and1 = s_dadda_pg_rca24_fa481_xor0 & s_dadda_pg_rca24_fa399_xor1;
  assign s_dadda_pg_rca24_fa481_or0 = s_dadda_pg_rca24_fa481_and0 | s_dadda_pg_rca24_fa481_and1;
  assign s_dadda_pg_rca24_and_22_22 = a[22] & b[22];
  assign s_dadda_pg_rca24_nand_21_23 = ~(a[21] & b[23]);
  assign s_dadda_pg_rca24_fa482_xor0 = s_dadda_pg_rca24_fa481_or0 ^ s_dadda_pg_rca24_and_22_22;
  assign s_dadda_pg_rca24_fa482_and0 = s_dadda_pg_rca24_fa481_or0 & s_dadda_pg_rca24_and_22_22;
  assign s_dadda_pg_rca24_fa482_xor1 = s_dadda_pg_rca24_fa482_xor0 ^ s_dadda_pg_rca24_nand_21_23;
  assign s_dadda_pg_rca24_fa482_and1 = s_dadda_pg_rca24_fa482_xor0 & s_dadda_pg_rca24_nand_21_23;
  assign s_dadda_pg_rca24_fa482_or0 = s_dadda_pg_rca24_fa482_and0 | s_dadda_pg_rca24_fa482_and1;
  assign s_dadda_pg_rca24_nand_23_22 = ~(a[23] & b[22]);
  assign s_dadda_pg_rca24_fa483_xor0 = s_dadda_pg_rca24_fa482_or0 ^ s_dadda_pg_rca24_fa440_or0;
  assign s_dadda_pg_rca24_fa483_and0 = s_dadda_pg_rca24_fa482_or0 & s_dadda_pg_rca24_fa440_or0;
  assign s_dadda_pg_rca24_fa483_xor1 = s_dadda_pg_rca24_fa483_xor0 ^ s_dadda_pg_rca24_nand_23_22;
  assign s_dadda_pg_rca24_fa483_and1 = s_dadda_pg_rca24_fa483_xor0 & s_dadda_pg_rca24_nand_23_22;
  assign s_dadda_pg_rca24_fa483_or0 = s_dadda_pg_rca24_fa483_and0 | s_dadda_pg_rca24_fa483_and1;
  assign s_dadda_pg_rca24_and_0_0 = a[0] & b[0];
  assign s_dadda_pg_rca24_and_1_0 = a[1] & b[0];
  assign s_dadda_pg_rca24_and_0_2 = a[0] & b[2];
  assign s_dadda_pg_rca24_nand_22_23 = ~(a[22] & b[23]);
  assign s_dadda_pg_rca24_and_0_1 = a[0] & b[1];
  assign s_dadda_pg_rca24_and_23_23 = a[23] & b[23];
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa0_xor0 = s_dadda_pg_rca24_and_1_0 ^ s_dadda_pg_rca24_and_0_1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa0_and0 = s_dadda_pg_rca24_and_1_0 & s_dadda_pg_rca24_and_0_1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor0 = s_dadda_pg_rca24_and_0_2 ^ s_dadda_pg_rca24_ha21_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa1_and0 = s_dadda_pg_rca24_and_0_2 & s_dadda_pg_rca24_ha21_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_pg_fa0_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_and1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa0_and0 & s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or1 = s_dadda_pg_rca24_u_pg_rca46_and1 | s_dadda_pg_rca24_u_pg_rca46_pg_fa1_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor0 = s_dadda_pg_rca24_ha20_xor0 ^ s_dadda_pg_rca24_fa441_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa2_and0 = s_dadda_pg_rca24_ha20_xor0 & s_dadda_pg_rca24_fa441_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or1;
  assign s_dadda_pg_rca24_u_pg_rca46_and2 = s_dadda_pg_rca24_u_pg_rca46_or1 & s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or2 = s_dadda_pg_rca24_u_pg_rca46_and2 | s_dadda_pg_rca24_u_pg_rca46_pg_fa2_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor0 = s_dadda_pg_rca24_fa400_xor1 ^ s_dadda_pg_rca24_fa442_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa3_and0 = s_dadda_pg_rca24_fa400_xor1 & s_dadda_pg_rca24_fa442_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or2;
  assign s_dadda_pg_rca24_u_pg_rca46_and3 = s_dadda_pg_rca24_u_pg_rca46_or2 & s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or3 = s_dadda_pg_rca24_u_pg_rca46_and3 | s_dadda_pg_rca24_u_pg_rca46_pg_fa3_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor0 = s_dadda_pg_rca24_fa401_xor1 ^ s_dadda_pg_rca24_fa443_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa4_and0 = s_dadda_pg_rca24_fa401_xor1 & s_dadda_pg_rca24_fa443_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or3;
  assign s_dadda_pg_rca24_u_pg_rca46_and4 = s_dadda_pg_rca24_u_pg_rca46_or3 & s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or4 = s_dadda_pg_rca24_u_pg_rca46_and4 | s_dadda_pg_rca24_u_pg_rca46_pg_fa4_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor0 = s_dadda_pg_rca24_fa402_xor1 ^ s_dadda_pg_rca24_fa444_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa5_and0 = s_dadda_pg_rca24_fa402_xor1 & s_dadda_pg_rca24_fa444_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or4;
  assign s_dadda_pg_rca24_u_pg_rca46_and5 = s_dadda_pg_rca24_u_pg_rca46_or4 & s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or5 = s_dadda_pg_rca24_u_pg_rca46_and5 | s_dadda_pg_rca24_u_pg_rca46_pg_fa5_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor0 = s_dadda_pg_rca24_fa403_xor1 ^ s_dadda_pg_rca24_fa445_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa6_and0 = s_dadda_pg_rca24_fa403_xor1 & s_dadda_pg_rca24_fa445_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or5;
  assign s_dadda_pg_rca24_u_pg_rca46_and6 = s_dadda_pg_rca24_u_pg_rca46_or5 & s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or6 = s_dadda_pg_rca24_u_pg_rca46_and6 | s_dadda_pg_rca24_u_pg_rca46_pg_fa6_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor0 = s_dadda_pg_rca24_fa404_xor1 ^ s_dadda_pg_rca24_fa446_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa7_and0 = s_dadda_pg_rca24_fa404_xor1 & s_dadda_pg_rca24_fa446_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or6;
  assign s_dadda_pg_rca24_u_pg_rca46_and7 = s_dadda_pg_rca24_u_pg_rca46_or6 & s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or7 = s_dadda_pg_rca24_u_pg_rca46_and7 | s_dadda_pg_rca24_u_pg_rca46_pg_fa7_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor0 = s_dadda_pg_rca24_fa405_xor1 ^ s_dadda_pg_rca24_fa447_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa8_and0 = s_dadda_pg_rca24_fa405_xor1 & s_dadda_pg_rca24_fa447_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or7;
  assign s_dadda_pg_rca24_u_pg_rca46_and8 = s_dadda_pg_rca24_u_pg_rca46_or7 & s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or8 = s_dadda_pg_rca24_u_pg_rca46_and8 | s_dadda_pg_rca24_u_pg_rca46_pg_fa8_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor0 = s_dadda_pg_rca24_fa406_xor1 ^ s_dadda_pg_rca24_fa448_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa9_and0 = s_dadda_pg_rca24_fa406_xor1 & s_dadda_pg_rca24_fa448_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or8;
  assign s_dadda_pg_rca24_u_pg_rca46_and9 = s_dadda_pg_rca24_u_pg_rca46_or8 & s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or9 = s_dadda_pg_rca24_u_pg_rca46_and9 | s_dadda_pg_rca24_u_pg_rca46_pg_fa9_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor0 = s_dadda_pg_rca24_fa407_xor1 ^ s_dadda_pg_rca24_fa449_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa10_and0 = s_dadda_pg_rca24_fa407_xor1 & s_dadda_pg_rca24_fa449_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or9;
  assign s_dadda_pg_rca24_u_pg_rca46_and10 = s_dadda_pg_rca24_u_pg_rca46_or9 & s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or10 = s_dadda_pg_rca24_u_pg_rca46_and10 | s_dadda_pg_rca24_u_pg_rca46_pg_fa10_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor0 = s_dadda_pg_rca24_fa408_xor1 ^ s_dadda_pg_rca24_fa450_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa11_and0 = s_dadda_pg_rca24_fa408_xor1 & s_dadda_pg_rca24_fa450_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or10;
  assign s_dadda_pg_rca24_u_pg_rca46_and11 = s_dadda_pg_rca24_u_pg_rca46_or10 & s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or11 = s_dadda_pg_rca24_u_pg_rca46_and11 | s_dadda_pg_rca24_u_pg_rca46_pg_fa11_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor0 = s_dadda_pg_rca24_fa409_xor1 ^ s_dadda_pg_rca24_fa451_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa12_and0 = s_dadda_pg_rca24_fa409_xor1 & s_dadda_pg_rca24_fa451_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or11;
  assign s_dadda_pg_rca24_u_pg_rca46_and12 = s_dadda_pg_rca24_u_pg_rca46_or11 & s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or12 = s_dadda_pg_rca24_u_pg_rca46_and12 | s_dadda_pg_rca24_u_pg_rca46_pg_fa12_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor0 = s_dadda_pg_rca24_fa410_xor1 ^ s_dadda_pg_rca24_fa452_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa13_and0 = s_dadda_pg_rca24_fa410_xor1 & s_dadda_pg_rca24_fa452_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or12;
  assign s_dadda_pg_rca24_u_pg_rca46_and13 = s_dadda_pg_rca24_u_pg_rca46_or12 & s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or13 = s_dadda_pg_rca24_u_pg_rca46_and13 | s_dadda_pg_rca24_u_pg_rca46_pg_fa13_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor0 = s_dadda_pg_rca24_fa411_xor1 ^ s_dadda_pg_rca24_fa453_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa14_and0 = s_dadda_pg_rca24_fa411_xor1 & s_dadda_pg_rca24_fa453_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or13;
  assign s_dadda_pg_rca24_u_pg_rca46_and14 = s_dadda_pg_rca24_u_pg_rca46_or13 & s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or14 = s_dadda_pg_rca24_u_pg_rca46_and14 | s_dadda_pg_rca24_u_pg_rca46_pg_fa14_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor0 = s_dadda_pg_rca24_fa412_xor1 ^ s_dadda_pg_rca24_fa454_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa15_and0 = s_dadda_pg_rca24_fa412_xor1 & s_dadda_pg_rca24_fa454_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or14;
  assign s_dadda_pg_rca24_u_pg_rca46_and15 = s_dadda_pg_rca24_u_pg_rca46_or14 & s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or15 = s_dadda_pg_rca24_u_pg_rca46_and15 | s_dadda_pg_rca24_u_pg_rca46_pg_fa15_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor0 = s_dadda_pg_rca24_fa413_xor1 ^ s_dadda_pg_rca24_fa455_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa16_and0 = s_dadda_pg_rca24_fa413_xor1 & s_dadda_pg_rca24_fa455_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or15;
  assign s_dadda_pg_rca24_u_pg_rca46_and16 = s_dadda_pg_rca24_u_pg_rca46_or15 & s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or16 = s_dadda_pg_rca24_u_pg_rca46_and16 | s_dadda_pg_rca24_u_pg_rca46_pg_fa16_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor0 = s_dadda_pg_rca24_fa414_xor1 ^ s_dadda_pg_rca24_fa456_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa17_and0 = s_dadda_pg_rca24_fa414_xor1 & s_dadda_pg_rca24_fa456_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or16;
  assign s_dadda_pg_rca24_u_pg_rca46_and17 = s_dadda_pg_rca24_u_pg_rca46_or16 & s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or17 = s_dadda_pg_rca24_u_pg_rca46_and17 | s_dadda_pg_rca24_u_pg_rca46_pg_fa17_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor0 = s_dadda_pg_rca24_fa415_xor1 ^ s_dadda_pg_rca24_fa457_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa18_and0 = s_dadda_pg_rca24_fa415_xor1 & s_dadda_pg_rca24_fa457_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or17;
  assign s_dadda_pg_rca24_u_pg_rca46_and18 = s_dadda_pg_rca24_u_pg_rca46_or17 & s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or18 = s_dadda_pg_rca24_u_pg_rca46_and18 | s_dadda_pg_rca24_u_pg_rca46_pg_fa18_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor0 = s_dadda_pg_rca24_fa416_xor1 ^ s_dadda_pg_rca24_fa458_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa19_and0 = s_dadda_pg_rca24_fa416_xor1 & s_dadda_pg_rca24_fa458_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or18;
  assign s_dadda_pg_rca24_u_pg_rca46_and19 = s_dadda_pg_rca24_u_pg_rca46_or18 & s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or19 = s_dadda_pg_rca24_u_pg_rca46_and19 | s_dadda_pg_rca24_u_pg_rca46_pg_fa19_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor0 = s_dadda_pg_rca24_fa417_xor1 ^ s_dadda_pg_rca24_fa459_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa20_and0 = s_dadda_pg_rca24_fa417_xor1 & s_dadda_pg_rca24_fa459_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or19;
  assign s_dadda_pg_rca24_u_pg_rca46_and20 = s_dadda_pg_rca24_u_pg_rca46_or19 & s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or20 = s_dadda_pg_rca24_u_pg_rca46_and20 | s_dadda_pg_rca24_u_pg_rca46_pg_fa20_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor0 = s_dadda_pg_rca24_fa418_xor1 ^ s_dadda_pg_rca24_fa460_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa21_and0 = s_dadda_pg_rca24_fa418_xor1 & s_dadda_pg_rca24_fa460_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or20;
  assign s_dadda_pg_rca24_u_pg_rca46_and21 = s_dadda_pg_rca24_u_pg_rca46_or20 & s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or21 = s_dadda_pg_rca24_u_pg_rca46_and21 | s_dadda_pg_rca24_u_pg_rca46_pg_fa21_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor0 = s_dadda_pg_rca24_fa419_xor1 ^ s_dadda_pg_rca24_fa461_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa22_and0 = s_dadda_pg_rca24_fa419_xor1 & s_dadda_pg_rca24_fa461_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or21;
  assign s_dadda_pg_rca24_u_pg_rca46_and22 = s_dadda_pg_rca24_u_pg_rca46_or21 & s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or22 = s_dadda_pg_rca24_u_pg_rca46_and22 | s_dadda_pg_rca24_u_pg_rca46_pg_fa22_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor0 = s_dadda_pg_rca24_fa420_xor1 ^ s_dadda_pg_rca24_fa462_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa23_and0 = s_dadda_pg_rca24_fa420_xor1 & s_dadda_pg_rca24_fa462_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or22;
  assign s_dadda_pg_rca24_u_pg_rca46_and23 = s_dadda_pg_rca24_u_pg_rca46_or22 & s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or23 = s_dadda_pg_rca24_u_pg_rca46_and23 | s_dadda_pg_rca24_u_pg_rca46_pg_fa23_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor0 = s_dadda_pg_rca24_fa421_xor1 ^ s_dadda_pg_rca24_fa463_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa24_and0 = s_dadda_pg_rca24_fa421_xor1 & s_dadda_pg_rca24_fa463_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or23;
  assign s_dadda_pg_rca24_u_pg_rca46_and24 = s_dadda_pg_rca24_u_pg_rca46_or23 & s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or24 = s_dadda_pg_rca24_u_pg_rca46_and24 | s_dadda_pg_rca24_u_pg_rca46_pg_fa24_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor0 = s_dadda_pg_rca24_fa422_xor1 ^ s_dadda_pg_rca24_fa464_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa25_and0 = s_dadda_pg_rca24_fa422_xor1 & s_dadda_pg_rca24_fa464_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or24;
  assign s_dadda_pg_rca24_u_pg_rca46_and25 = s_dadda_pg_rca24_u_pg_rca46_or24 & s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or25 = s_dadda_pg_rca24_u_pg_rca46_and25 | s_dadda_pg_rca24_u_pg_rca46_pg_fa25_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor0 = s_dadda_pg_rca24_fa423_xor1 ^ s_dadda_pg_rca24_fa465_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa26_and0 = s_dadda_pg_rca24_fa423_xor1 & s_dadda_pg_rca24_fa465_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or25;
  assign s_dadda_pg_rca24_u_pg_rca46_and26 = s_dadda_pg_rca24_u_pg_rca46_or25 & s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or26 = s_dadda_pg_rca24_u_pg_rca46_and26 | s_dadda_pg_rca24_u_pg_rca46_pg_fa26_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor0 = s_dadda_pg_rca24_fa424_xor1 ^ s_dadda_pg_rca24_fa466_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa27_and0 = s_dadda_pg_rca24_fa424_xor1 & s_dadda_pg_rca24_fa466_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or26;
  assign s_dadda_pg_rca24_u_pg_rca46_and27 = s_dadda_pg_rca24_u_pg_rca46_or26 & s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or27 = s_dadda_pg_rca24_u_pg_rca46_and27 | s_dadda_pg_rca24_u_pg_rca46_pg_fa27_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor0 = s_dadda_pg_rca24_fa425_xor1 ^ s_dadda_pg_rca24_fa467_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa28_and0 = s_dadda_pg_rca24_fa425_xor1 & s_dadda_pg_rca24_fa467_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or27;
  assign s_dadda_pg_rca24_u_pg_rca46_and28 = s_dadda_pg_rca24_u_pg_rca46_or27 & s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or28 = s_dadda_pg_rca24_u_pg_rca46_and28 | s_dadda_pg_rca24_u_pg_rca46_pg_fa28_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor0 = s_dadda_pg_rca24_fa426_xor1 ^ s_dadda_pg_rca24_fa468_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa29_and0 = s_dadda_pg_rca24_fa426_xor1 & s_dadda_pg_rca24_fa468_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or28;
  assign s_dadda_pg_rca24_u_pg_rca46_and29 = s_dadda_pg_rca24_u_pg_rca46_or28 & s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or29 = s_dadda_pg_rca24_u_pg_rca46_and29 | s_dadda_pg_rca24_u_pg_rca46_pg_fa29_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor0 = s_dadda_pg_rca24_fa427_xor1 ^ s_dadda_pg_rca24_fa469_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa30_and0 = s_dadda_pg_rca24_fa427_xor1 & s_dadda_pg_rca24_fa469_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or29;
  assign s_dadda_pg_rca24_u_pg_rca46_and30 = s_dadda_pg_rca24_u_pg_rca46_or29 & s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or30 = s_dadda_pg_rca24_u_pg_rca46_and30 | s_dadda_pg_rca24_u_pg_rca46_pg_fa30_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor0 = s_dadda_pg_rca24_fa428_xor1 ^ s_dadda_pg_rca24_fa470_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa31_and0 = s_dadda_pg_rca24_fa428_xor1 & s_dadda_pg_rca24_fa470_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or30;
  assign s_dadda_pg_rca24_u_pg_rca46_and31 = s_dadda_pg_rca24_u_pg_rca46_or30 & s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or31 = s_dadda_pg_rca24_u_pg_rca46_and31 | s_dadda_pg_rca24_u_pg_rca46_pg_fa31_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor0 = s_dadda_pg_rca24_fa429_xor1 ^ s_dadda_pg_rca24_fa471_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa32_and0 = s_dadda_pg_rca24_fa429_xor1 & s_dadda_pg_rca24_fa471_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or31;
  assign s_dadda_pg_rca24_u_pg_rca46_and32 = s_dadda_pg_rca24_u_pg_rca46_or31 & s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or32 = s_dadda_pg_rca24_u_pg_rca46_and32 | s_dadda_pg_rca24_u_pg_rca46_pg_fa32_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor0 = s_dadda_pg_rca24_fa430_xor1 ^ s_dadda_pg_rca24_fa472_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa33_and0 = s_dadda_pg_rca24_fa430_xor1 & s_dadda_pg_rca24_fa472_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or32;
  assign s_dadda_pg_rca24_u_pg_rca46_and33 = s_dadda_pg_rca24_u_pg_rca46_or32 & s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or33 = s_dadda_pg_rca24_u_pg_rca46_and33 | s_dadda_pg_rca24_u_pg_rca46_pg_fa33_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor0 = s_dadda_pg_rca24_fa431_xor1 ^ s_dadda_pg_rca24_fa473_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa34_and0 = s_dadda_pg_rca24_fa431_xor1 & s_dadda_pg_rca24_fa473_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or33;
  assign s_dadda_pg_rca24_u_pg_rca46_and34 = s_dadda_pg_rca24_u_pg_rca46_or33 & s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or34 = s_dadda_pg_rca24_u_pg_rca46_and34 | s_dadda_pg_rca24_u_pg_rca46_pg_fa34_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor0 = s_dadda_pg_rca24_fa432_xor1 ^ s_dadda_pg_rca24_fa474_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa35_and0 = s_dadda_pg_rca24_fa432_xor1 & s_dadda_pg_rca24_fa474_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or34;
  assign s_dadda_pg_rca24_u_pg_rca46_and35 = s_dadda_pg_rca24_u_pg_rca46_or34 & s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or35 = s_dadda_pg_rca24_u_pg_rca46_and35 | s_dadda_pg_rca24_u_pg_rca46_pg_fa35_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor0 = s_dadda_pg_rca24_fa433_xor1 ^ s_dadda_pg_rca24_fa475_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa36_and0 = s_dadda_pg_rca24_fa433_xor1 & s_dadda_pg_rca24_fa475_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or35;
  assign s_dadda_pg_rca24_u_pg_rca46_and36 = s_dadda_pg_rca24_u_pg_rca46_or35 & s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or36 = s_dadda_pg_rca24_u_pg_rca46_and36 | s_dadda_pg_rca24_u_pg_rca46_pg_fa36_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor0 = s_dadda_pg_rca24_fa434_xor1 ^ s_dadda_pg_rca24_fa476_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa37_and0 = s_dadda_pg_rca24_fa434_xor1 & s_dadda_pg_rca24_fa476_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or36;
  assign s_dadda_pg_rca24_u_pg_rca46_and37 = s_dadda_pg_rca24_u_pg_rca46_or36 & s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or37 = s_dadda_pg_rca24_u_pg_rca46_and37 | s_dadda_pg_rca24_u_pg_rca46_pg_fa37_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor0 = s_dadda_pg_rca24_fa435_xor1 ^ s_dadda_pg_rca24_fa477_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa38_and0 = s_dadda_pg_rca24_fa435_xor1 & s_dadda_pg_rca24_fa477_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or37;
  assign s_dadda_pg_rca24_u_pg_rca46_and38 = s_dadda_pg_rca24_u_pg_rca46_or37 & s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or38 = s_dadda_pg_rca24_u_pg_rca46_and38 | s_dadda_pg_rca24_u_pg_rca46_pg_fa38_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor0 = s_dadda_pg_rca24_fa436_xor1 ^ s_dadda_pg_rca24_fa478_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa39_and0 = s_dadda_pg_rca24_fa436_xor1 & s_dadda_pg_rca24_fa478_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or38;
  assign s_dadda_pg_rca24_u_pg_rca46_and39 = s_dadda_pg_rca24_u_pg_rca46_or38 & s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or39 = s_dadda_pg_rca24_u_pg_rca46_and39 | s_dadda_pg_rca24_u_pg_rca46_pg_fa39_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor0 = s_dadda_pg_rca24_fa437_xor1 ^ s_dadda_pg_rca24_fa479_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa40_and0 = s_dadda_pg_rca24_fa437_xor1 & s_dadda_pg_rca24_fa479_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or39;
  assign s_dadda_pg_rca24_u_pg_rca46_and40 = s_dadda_pg_rca24_u_pg_rca46_or39 & s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or40 = s_dadda_pg_rca24_u_pg_rca46_and40 | s_dadda_pg_rca24_u_pg_rca46_pg_fa40_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor0 = s_dadda_pg_rca24_fa438_xor1 ^ s_dadda_pg_rca24_fa480_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa41_and0 = s_dadda_pg_rca24_fa438_xor1 & s_dadda_pg_rca24_fa480_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or40;
  assign s_dadda_pg_rca24_u_pg_rca46_and41 = s_dadda_pg_rca24_u_pg_rca46_or40 & s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or41 = s_dadda_pg_rca24_u_pg_rca46_and41 | s_dadda_pg_rca24_u_pg_rca46_pg_fa41_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor0 = s_dadda_pg_rca24_fa439_xor1 ^ s_dadda_pg_rca24_fa481_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa42_and0 = s_dadda_pg_rca24_fa439_xor1 & s_dadda_pg_rca24_fa481_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or41;
  assign s_dadda_pg_rca24_u_pg_rca46_and42 = s_dadda_pg_rca24_u_pg_rca46_or41 & s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or42 = s_dadda_pg_rca24_u_pg_rca46_and42 | s_dadda_pg_rca24_u_pg_rca46_pg_fa42_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor0 = s_dadda_pg_rca24_fa440_xor1 ^ s_dadda_pg_rca24_fa482_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa43_and0 = s_dadda_pg_rca24_fa440_xor1 & s_dadda_pg_rca24_fa482_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or42;
  assign s_dadda_pg_rca24_u_pg_rca46_and43 = s_dadda_pg_rca24_u_pg_rca46_or42 & s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or43 = s_dadda_pg_rca24_u_pg_rca46_and43 | s_dadda_pg_rca24_u_pg_rca46_pg_fa43_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor0 = s_dadda_pg_rca24_nand_22_23 ^ s_dadda_pg_rca24_fa483_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa44_and0 = s_dadda_pg_rca24_nand_22_23 & s_dadda_pg_rca24_fa483_xor1;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or43;
  assign s_dadda_pg_rca24_u_pg_rca46_and44 = s_dadda_pg_rca24_u_pg_rca46_or43 & s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or44 = s_dadda_pg_rca24_u_pg_rca46_and44 | s_dadda_pg_rca24_u_pg_rca46_pg_fa44_and0;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor0 = s_dadda_pg_rca24_fa483_or0 ^ s_dadda_pg_rca24_and_23_23;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa45_and0 = s_dadda_pg_rca24_fa483_or0 & s_dadda_pg_rca24_and_23_23;
  assign s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor1 = s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor0 ^ s_dadda_pg_rca24_u_pg_rca46_or44;
  assign s_dadda_pg_rca24_u_pg_rca46_and45 = s_dadda_pg_rca24_u_pg_rca46_or44 & s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor0;
  assign s_dadda_pg_rca24_u_pg_rca46_or45 = s_dadda_pg_rca24_u_pg_rca46_and45 | s_dadda_pg_rca24_u_pg_rca46_pg_fa45_and0;
  assign s_dadda_pg_rca24_xor0 = ~s_dadda_pg_rca24_u_pg_rca46_or45;

  assign s_dadda_pg_rca24_out[0] = s_dadda_pg_rca24_and_0_0;
  assign s_dadda_pg_rca24_out[1] = s_dadda_pg_rca24_u_pg_rca46_pg_fa0_xor0;
  assign s_dadda_pg_rca24_out[2] = s_dadda_pg_rca24_u_pg_rca46_pg_fa1_xor1;
  assign s_dadda_pg_rca24_out[3] = s_dadda_pg_rca24_u_pg_rca46_pg_fa2_xor1;
  assign s_dadda_pg_rca24_out[4] = s_dadda_pg_rca24_u_pg_rca46_pg_fa3_xor1;
  assign s_dadda_pg_rca24_out[5] = s_dadda_pg_rca24_u_pg_rca46_pg_fa4_xor1;
  assign s_dadda_pg_rca24_out[6] = s_dadda_pg_rca24_u_pg_rca46_pg_fa5_xor1;
  assign s_dadda_pg_rca24_out[7] = s_dadda_pg_rca24_u_pg_rca46_pg_fa6_xor1;
  assign s_dadda_pg_rca24_out[8] = s_dadda_pg_rca24_u_pg_rca46_pg_fa7_xor1;
  assign s_dadda_pg_rca24_out[9] = s_dadda_pg_rca24_u_pg_rca46_pg_fa8_xor1;
  assign s_dadda_pg_rca24_out[10] = s_dadda_pg_rca24_u_pg_rca46_pg_fa9_xor1;
  assign s_dadda_pg_rca24_out[11] = s_dadda_pg_rca24_u_pg_rca46_pg_fa10_xor1;
  assign s_dadda_pg_rca24_out[12] = s_dadda_pg_rca24_u_pg_rca46_pg_fa11_xor1;
  assign s_dadda_pg_rca24_out[13] = s_dadda_pg_rca24_u_pg_rca46_pg_fa12_xor1;
  assign s_dadda_pg_rca24_out[14] = s_dadda_pg_rca24_u_pg_rca46_pg_fa13_xor1;
  assign s_dadda_pg_rca24_out[15] = s_dadda_pg_rca24_u_pg_rca46_pg_fa14_xor1;
  assign s_dadda_pg_rca24_out[16] = s_dadda_pg_rca24_u_pg_rca46_pg_fa15_xor1;
  assign s_dadda_pg_rca24_out[17] = s_dadda_pg_rca24_u_pg_rca46_pg_fa16_xor1;
  assign s_dadda_pg_rca24_out[18] = s_dadda_pg_rca24_u_pg_rca46_pg_fa17_xor1;
  assign s_dadda_pg_rca24_out[19] = s_dadda_pg_rca24_u_pg_rca46_pg_fa18_xor1;
  assign s_dadda_pg_rca24_out[20] = s_dadda_pg_rca24_u_pg_rca46_pg_fa19_xor1;
  assign s_dadda_pg_rca24_out[21] = s_dadda_pg_rca24_u_pg_rca46_pg_fa20_xor1;
  assign s_dadda_pg_rca24_out[22] = s_dadda_pg_rca24_u_pg_rca46_pg_fa21_xor1;
  assign s_dadda_pg_rca24_out[23] = s_dadda_pg_rca24_u_pg_rca46_pg_fa22_xor1;
  assign s_dadda_pg_rca24_out[24] = s_dadda_pg_rca24_u_pg_rca46_pg_fa23_xor1;
  assign s_dadda_pg_rca24_out[25] = s_dadda_pg_rca24_u_pg_rca46_pg_fa24_xor1;
  assign s_dadda_pg_rca24_out[26] = s_dadda_pg_rca24_u_pg_rca46_pg_fa25_xor1;
  assign s_dadda_pg_rca24_out[27] = s_dadda_pg_rca24_u_pg_rca46_pg_fa26_xor1;
  assign s_dadda_pg_rca24_out[28] = s_dadda_pg_rca24_u_pg_rca46_pg_fa27_xor1;
  assign s_dadda_pg_rca24_out[29] = s_dadda_pg_rca24_u_pg_rca46_pg_fa28_xor1;
  assign s_dadda_pg_rca24_out[30] = s_dadda_pg_rca24_u_pg_rca46_pg_fa29_xor1;
  assign s_dadda_pg_rca24_out[31] = s_dadda_pg_rca24_u_pg_rca46_pg_fa30_xor1;
  assign s_dadda_pg_rca24_out[32] = s_dadda_pg_rca24_u_pg_rca46_pg_fa31_xor1;
  assign s_dadda_pg_rca24_out[33] = s_dadda_pg_rca24_u_pg_rca46_pg_fa32_xor1;
  assign s_dadda_pg_rca24_out[34] = s_dadda_pg_rca24_u_pg_rca46_pg_fa33_xor1;
  assign s_dadda_pg_rca24_out[35] = s_dadda_pg_rca24_u_pg_rca46_pg_fa34_xor1;
  assign s_dadda_pg_rca24_out[36] = s_dadda_pg_rca24_u_pg_rca46_pg_fa35_xor1;
  assign s_dadda_pg_rca24_out[37] = s_dadda_pg_rca24_u_pg_rca46_pg_fa36_xor1;
  assign s_dadda_pg_rca24_out[38] = s_dadda_pg_rca24_u_pg_rca46_pg_fa37_xor1;
  assign s_dadda_pg_rca24_out[39] = s_dadda_pg_rca24_u_pg_rca46_pg_fa38_xor1;
  assign s_dadda_pg_rca24_out[40] = s_dadda_pg_rca24_u_pg_rca46_pg_fa39_xor1;
  assign s_dadda_pg_rca24_out[41] = s_dadda_pg_rca24_u_pg_rca46_pg_fa40_xor1;
  assign s_dadda_pg_rca24_out[42] = s_dadda_pg_rca24_u_pg_rca46_pg_fa41_xor1;
  assign s_dadda_pg_rca24_out[43] = s_dadda_pg_rca24_u_pg_rca46_pg_fa42_xor1;
  assign s_dadda_pg_rca24_out[44] = s_dadda_pg_rca24_u_pg_rca46_pg_fa43_xor1;
  assign s_dadda_pg_rca24_out[45] = s_dadda_pg_rca24_u_pg_rca46_pg_fa44_xor1;
  assign s_dadda_pg_rca24_out[46] = s_dadda_pg_rca24_u_pg_rca46_pg_fa45_xor1;
  assign s_dadda_pg_rca24_out[47] = s_dadda_pg_rca24_xor0;
endmodule