module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_cin;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module h_u_arrmul32(input [31:0] a, input [31:0] b, output [63:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire a_30;
  wire a_31;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire b_30;
  wire b_31;
  wire h_u_arrmul32_and0_0_y0;
  wire h_u_arrmul32_and1_0_y0;
  wire h_u_arrmul32_and2_0_y0;
  wire h_u_arrmul32_and3_0_y0;
  wire h_u_arrmul32_and4_0_y0;
  wire h_u_arrmul32_and5_0_y0;
  wire h_u_arrmul32_and6_0_y0;
  wire h_u_arrmul32_and7_0_y0;
  wire h_u_arrmul32_and8_0_y0;
  wire h_u_arrmul32_and9_0_y0;
  wire h_u_arrmul32_and10_0_y0;
  wire h_u_arrmul32_and11_0_y0;
  wire h_u_arrmul32_and12_0_y0;
  wire h_u_arrmul32_and13_0_y0;
  wire h_u_arrmul32_and14_0_y0;
  wire h_u_arrmul32_and15_0_y0;
  wire h_u_arrmul32_and16_0_y0;
  wire h_u_arrmul32_and17_0_y0;
  wire h_u_arrmul32_and18_0_y0;
  wire h_u_arrmul32_and19_0_y0;
  wire h_u_arrmul32_and20_0_y0;
  wire h_u_arrmul32_and21_0_y0;
  wire h_u_arrmul32_and22_0_y0;
  wire h_u_arrmul32_and23_0_y0;
  wire h_u_arrmul32_and24_0_y0;
  wire h_u_arrmul32_and25_0_y0;
  wire h_u_arrmul32_and26_0_y0;
  wire h_u_arrmul32_and27_0_y0;
  wire h_u_arrmul32_and28_0_y0;
  wire h_u_arrmul32_and29_0_y0;
  wire h_u_arrmul32_and30_0_y0;
  wire h_u_arrmul32_and31_0_y0;
  wire h_u_arrmul32_and0_1_y0;
  wire h_u_arrmul32_ha0_1_y0;
  wire h_u_arrmul32_ha0_1_y1;
  wire h_u_arrmul32_and1_1_y0;
  wire h_u_arrmul32_fa1_1_y2;
  wire h_u_arrmul32_fa1_1_y4;
  wire h_u_arrmul32_and2_1_y0;
  wire h_u_arrmul32_fa2_1_y2;
  wire h_u_arrmul32_fa2_1_y4;
  wire h_u_arrmul32_and3_1_y0;
  wire h_u_arrmul32_fa3_1_y2;
  wire h_u_arrmul32_fa3_1_y4;
  wire h_u_arrmul32_and4_1_y0;
  wire h_u_arrmul32_fa4_1_y2;
  wire h_u_arrmul32_fa4_1_y4;
  wire h_u_arrmul32_and5_1_y0;
  wire h_u_arrmul32_fa5_1_y2;
  wire h_u_arrmul32_fa5_1_y4;
  wire h_u_arrmul32_and6_1_y0;
  wire h_u_arrmul32_fa6_1_y2;
  wire h_u_arrmul32_fa6_1_y4;
  wire h_u_arrmul32_and7_1_y0;
  wire h_u_arrmul32_fa7_1_y2;
  wire h_u_arrmul32_fa7_1_y4;
  wire h_u_arrmul32_and8_1_y0;
  wire h_u_arrmul32_fa8_1_y2;
  wire h_u_arrmul32_fa8_1_y4;
  wire h_u_arrmul32_and9_1_y0;
  wire h_u_arrmul32_fa9_1_y2;
  wire h_u_arrmul32_fa9_1_y4;
  wire h_u_arrmul32_and10_1_y0;
  wire h_u_arrmul32_fa10_1_y2;
  wire h_u_arrmul32_fa10_1_y4;
  wire h_u_arrmul32_and11_1_y0;
  wire h_u_arrmul32_fa11_1_y2;
  wire h_u_arrmul32_fa11_1_y4;
  wire h_u_arrmul32_and12_1_y0;
  wire h_u_arrmul32_fa12_1_y2;
  wire h_u_arrmul32_fa12_1_y4;
  wire h_u_arrmul32_and13_1_y0;
  wire h_u_arrmul32_fa13_1_y2;
  wire h_u_arrmul32_fa13_1_y4;
  wire h_u_arrmul32_and14_1_y0;
  wire h_u_arrmul32_fa14_1_y2;
  wire h_u_arrmul32_fa14_1_y4;
  wire h_u_arrmul32_and15_1_y0;
  wire h_u_arrmul32_fa15_1_y2;
  wire h_u_arrmul32_fa15_1_y4;
  wire h_u_arrmul32_and16_1_y0;
  wire h_u_arrmul32_fa16_1_y2;
  wire h_u_arrmul32_fa16_1_y4;
  wire h_u_arrmul32_and17_1_y0;
  wire h_u_arrmul32_fa17_1_y2;
  wire h_u_arrmul32_fa17_1_y4;
  wire h_u_arrmul32_and18_1_y0;
  wire h_u_arrmul32_fa18_1_y2;
  wire h_u_arrmul32_fa18_1_y4;
  wire h_u_arrmul32_and19_1_y0;
  wire h_u_arrmul32_fa19_1_y2;
  wire h_u_arrmul32_fa19_1_y4;
  wire h_u_arrmul32_and20_1_y0;
  wire h_u_arrmul32_fa20_1_y2;
  wire h_u_arrmul32_fa20_1_y4;
  wire h_u_arrmul32_and21_1_y0;
  wire h_u_arrmul32_fa21_1_y2;
  wire h_u_arrmul32_fa21_1_y4;
  wire h_u_arrmul32_and22_1_y0;
  wire h_u_arrmul32_fa22_1_y2;
  wire h_u_arrmul32_fa22_1_y4;
  wire h_u_arrmul32_and23_1_y0;
  wire h_u_arrmul32_fa23_1_y2;
  wire h_u_arrmul32_fa23_1_y4;
  wire h_u_arrmul32_and24_1_y0;
  wire h_u_arrmul32_fa24_1_y2;
  wire h_u_arrmul32_fa24_1_y4;
  wire h_u_arrmul32_and25_1_y0;
  wire h_u_arrmul32_fa25_1_y2;
  wire h_u_arrmul32_fa25_1_y4;
  wire h_u_arrmul32_and26_1_y0;
  wire h_u_arrmul32_fa26_1_y2;
  wire h_u_arrmul32_fa26_1_y4;
  wire h_u_arrmul32_and27_1_y0;
  wire h_u_arrmul32_fa27_1_y2;
  wire h_u_arrmul32_fa27_1_y4;
  wire h_u_arrmul32_and28_1_y0;
  wire h_u_arrmul32_fa28_1_y2;
  wire h_u_arrmul32_fa28_1_y4;
  wire h_u_arrmul32_and29_1_y0;
  wire h_u_arrmul32_fa29_1_y2;
  wire h_u_arrmul32_fa29_1_y4;
  wire h_u_arrmul32_and30_1_y0;
  wire h_u_arrmul32_fa30_1_y2;
  wire h_u_arrmul32_fa30_1_y4;
  wire h_u_arrmul32_and31_1_y0;
  wire h_u_arrmul32_ha31_1_y0;
  wire h_u_arrmul32_ha31_1_y1;
  wire h_u_arrmul32_and0_2_y0;
  wire h_u_arrmul32_ha0_2_y0;
  wire h_u_arrmul32_ha0_2_y1;
  wire h_u_arrmul32_and1_2_y0;
  wire h_u_arrmul32_fa1_2_y2;
  wire h_u_arrmul32_fa1_2_y4;
  wire h_u_arrmul32_and2_2_y0;
  wire h_u_arrmul32_fa2_2_y2;
  wire h_u_arrmul32_fa2_2_y4;
  wire h_u_arrmul32_and3_2_y0;
  wire h_u_arrmul32_fa3_2_y2;
  wire h_u_arrmul32_fa3_2_y4;
  wire h_u_arrmul32_and4_2_y0;
  wire h_u_arrmul32_fa4_2_y2;
  wire h_u_arrmul32_fa4_2_y4;
  wire h_u_arrmul32_and5_2_y0;
  wire h_u_arrmul32_fa5_2_y2;
  wire h_u_arrmul32_fa5_2_y4;
  wire h_u_arrmul32_and6_2_y0;
  wire h_u_arrmul32_fa6_2_y2;
  wire h_u_arrmul32_fa6_2_y4;
  wire h_u_arrmul32_and7_2_y0;
  wire h_u_arrmul32_fa7_2_y2;
  wire h_u_arrmul32_fa7_2_y4;
  wire h_u_arrmul32_and8_2_y0;
  wire h_u_arrmul32_fa8_2_y2;
  wire h_u_arrmul32_fa8_2_y4;
  wire h_u_arrmul32_and9_2_y0;
  wire h_u_arrmul32_fa9_2_y2;
  wire h_u_arrmul32_fa9_2_y4;
  wire h_u_arrmul32_and10_2_y0;
  wire h_u_arrmul32_fa10_2_y2;
  wire h_u_arrmul32_fa10_2_y4;
  wire h_u_arrmul32_and11_2_y0;
  wire h_u_arrmul32_fa11_2_y2;
  wire h_u_arrmul32_fa11_2_y4;
  wire h_u_arrmul32_and12_2_y0;
  wire h_u_arrmul32_fa12_2_y2;
  wire h_u_arrmul32_fa12_2_y4;
  wire h_u_arrmul32_and13_2_y0;
  wire h_u_arrmul32_fa13_2_y2;
  wire h_u_arrmul32_fa13_2_y4;
  wire h_u_arrmul32_and14_2_y0;
  wire h_u_arrmul32_fa14_2_y2;
  wire h_u_arrmul32_fa14_2_y4;
  wire h_u_arrmul32_and15_2_y0;
  wire h_u_arrmul32_fa15_2_y2;
  wire h_u_arrmul32_fa15_2_y4;
  wire h_u_arrmul32_and16_2_y0;
  wire h_u_arrmul32_fa16_2_y2;
  wire h_u_arrmul32_fa16_2_y4;
  wire h_u_arrmul32_and17_2_y0;
  wire h_u_arrmul32_fa17_2_y2;
  wire h_u_arrmul32_fa17_2_y4;
  wire h_u_arrmul32_and18_2_y0;
  wire h_u_arrmul32_fa18_2_y2;
  wire h_u_arrmul32_fa18_2_y4;
  wire h_u_arrmul32_and19_2_y0;
  wire h_u_arrmul32_fa19_2_y2;
  wire h_u_arrmul32_fa19_2_y4;
  wire h_u_arrmul32_and20_2_y0;
  wire h_u_arrmul32_fa20_2_y2;
  wire h_u_arrmul32_fa20_2_y4;
  wire h_u_arrmul32_and21_2_y0;
  wire h_u_arrmul32_fa21_2_y2;
  wire h_u_arrmul32_fa21_2_y4;
  wire h_u_arrmul32_and22_2_y0;
  wire h_u_arrmul32_fa22_2_y2;
  wire h_u_arrmul32_fa22_2_y4;
  wire h_u_arrmul32_and23_2_y0;
  wire h_u_arrmul32_fa23_2_y2;
  wire h_u_arrmul32_fa23_2_y4;
  wire h_u_arrmul32_and24_2_y0;
  wire h_u_arrmul32_fa24_2_y2;
  wire h_u_arrmul32_fa24_2_y4;
  wire h_u_arrmul32_and25_2_y0;
  wire h_u_arrmul32_fa25_2_y2;
  wire h_u_arrmul32_fa25_2_y4;
  wire h_u_arrmul32_and26_2_y0;
  wire h_u_arrmul32_fa26_2_y2;
  wire h_u_arrmul32_fa26_2_y4;
  wire h_u_arrmul32_and27_2_y0;
  wire h_u_arrmul32_fa27_2_y2;
  wire h_u_arrmul32_fa27_2_y4;
  wire h_u_arrmul32_and28_2_y0;
  wire h_u_arrmul32_fa28_2_y2;
  wire h_u_arrmul32_fa28_2_y4;
  wire h_u_arrmul32_and29_2_y0;
  wire h_u_arrmul32_fa29_2_y2;
  wire h_u_arrmul32_fa29_2_y4;
  wire h_u_arrmul32_and30_2_y0;
  wire h_u_arrmul32_fa30_2_y2;
  wire h_u_arrmul32_fa30_2_y4;
  wire h_u_arrmul32_and31_2_y0;
  wire h_u_arrmul32_fa31_2_y2;
  wire h_u_arrmul32_fa31_2_y4;
  wire h_u_arrmul32_and0_3_y0;
  wire h_u_arrmul32_ha0_3_y0;
  wire h_u_arrmul32_ha0_3_y1;
  wire h_u_arrmul32_and1_3_y0;
  wire h_u_arrmul32_fa1_3_y2;
  wire h_u_arrmul32_fa1_3_y4;
  wire h_u_arrmul32_and2_3_y0;
  wire h_u_arrmul32_fa2_3_y2;
  wire h_u_arrmul32_fa2_3_y4;
  wire h_u_arrmul32_and3_3_y0;
  wire h_u_arrmul32_fa3_3_y2;
  wire h_u_arrmul32_fa3_3_y4;
  wire h_u_arrmul32_and4_3_y0;
  wire h_u_arrmul32_fa4_3_y2;
  wire h_u_arrmul32_fa4_3_y4;
  wire h_u_arrmul32_and5_3_y0;
  wire h_u_arrmul32_fa5_3_y2;
  wire h_u_arrmul32_fa5_3_y4;
  wire h_u_arrmul32_and6_3_y0;
  wire h_u_arrmul32_fa6_3_y2;
  wire h_u_arrmul32_fa6_3_y4;
  wire h_u_arrmul32_and7_3_y0;
  wire h_u_arrmul32_fa7_3_y2;
  wire h_u_arrmul32_fa7_3_y4;
  wire h_u_arrmul32_and8_3_y0;
  wire h_u_arrmul32_fa8_3_y2;
  wire h_u_arrmul32_fa8_3_y4;
  wire h_u_arrmul32_and9_3_y0;
  wire h_u_arrmul32_fa9_3_y2;
  wire h_u_arrmul32_fa9_3_y4;
  wire h_u_arrmul32_and10_3_y0;
  wire h_u_arrmul32_fa10_3_y2;
  wire h_u_arrmul32_fa10_3_y4;
  wire h_u_arrmul32_and11_3_y0;
  wire h_u_arrmul32_fa11_3_y2;
  wire h_u_arrmul32_fa11_3_y4;
  wire h_u_arrmul32_and12_3_y0;
  wire h_u_arrmul32_fa12_3_y2;
  wire h_u_arrmul32_fa12_3_y4;
  wire h_u_arrmul32_and13_3_y0;
  wire h_u_arrmul32_fa13_3_y2;
  wire h_u_arrmul32_fa13_3_y4;
  wire h_u_arrmul32_and14_3_y0;
  wire h_u_arrmul32_fa14_3_y2;
  wire h_u_arrmul32_fa14_3_y4;
  wire h_u_arrmul32_and15_3_y0;
  wire h_u_arrmul32_fa15_3_y2;
  wire h_u_arrmul32_fa15_3_y4;
  wire h_u_arrmul32_and16_3_y0;
  wire h_u_arrmul32_fa16_3_y2;
  wire h_u_arrmul32_fa16_3_y4;
  wire h_u_arrmul32_and17_3_y0;
  wire h_u_arrmul32_fa17_3_y2;
  wire h_u_arrmul32_fa17_3_y4;
  wire h_u_arrmul32_and18_3_y0;
  wire h_u_arrmul32_fa18_3_y2;
  wire h_u_arrmul32_fa18_3_y4;
  wire h_u_arrmul32_and19_3_y0;
  wire h_u_arrmul32_fa19_3_y2;
  wire h_u_arrmul32_fa19_3_y4;
  wire h_u_arrmul32_and20_3_y0;
  wire h_u_arrmul32_fa20_3_y2;
  wire h_u_arrmul32_fa20_3_y4;
  wire h_u_arrmul32_and21_3_y0;
  wire h_u_arrmul32_fa21_3_y2;
  wire h_u_arrmul32_fa21_3_y4;
  wire h_u_arrmul32_and22_3_y0;
  wire h_u_arrmul32_fa22_3_y2;
  wire h_u_arrmul32_fa22_3_y4;
  wire h_u_arrmul32_and23_3_y0;
  wire h_u_arrmul32_fa23_3_y2;
  wire h_u_arrmul32_fa23_3_y4;
  wire h_u_arrmul32_and24_3_y0;
  wire h_u_arrmul32_fa24_3_y2;
  wire h_u_arrmul32_fa24_3_y4;
  wire h_u_arrmul32_and25_3_y0;
  wire h_u_arrmul32_fa25_3_y2;
  wire h_u_arrmul32_fa25_3_y4;
  wire h_u_arrmul32_and26_3_y0;
  wire h_u_arrmul32_fa26_3_y2;
  wire h_u_arrmul32_fa26_3_y4;
  wire h_u_arrmul32_and27_3_y0;
  wire h_u_arrmul32_fa27_3_y2;
  wire h_u_arrmul32_fa27_3_y4;
  wire h_u_arrmul32_and28_3_y0;
  wire h_u_arrmul32_fa28_3_y2;
  wire h_u_arrmul32_fa28_3_y4;
  wire h_u_arrmul32_and29_3_y0;
  wire h_u_arrmul32_fa29_3_y2;
  wire h_u_arrmul32_fa29_3_y4;
  wire h_u_arrmul32_and30_3_y0;
  wire h_u_arrmul32_fa30_3_y2;
  wire h_u_arrmul32_fa30_3_y4;
  wire h_u_arrmul32_and31_3_y0;
  wire h_u_arrmul32_fa31_3_y2;
  wire h_u_arrmul32_fa31_3_y4;
  wire h_u_arrmul32_and0_4_y0;
  wire h_u_arrmul32_ha0_4_y0;
  wire h_u_arrmul32_ha0_4_y1;
  wire h_u_arrmul32_and1_4_y0;
  wire h_u_arrmul32_fa1_4_y2;
  wire h_u_arrmul32_fa1_4_y4;
  wire h_u_arrmul32_and2_4_y0;
  wire h_u_arrmul32_fa2_4_y2;
  wire h_u_arrmul32_fa2_4_y4;
  wire h_u_arrmul32_and3_4_y0;
  wire h_u_arrmul32_fa3_4_y2;
  wire h_u_arrmul32_fa3_4_y4;
  wire h_u_arrmul32_and4_4_y0;
  wire h_u_arrmul32_fa4_4_y2;
  wire h_u_arrmul32_fa4_4_y4;
  wire h_u_arrmul32_and5_4_y0;
  wire h_u_arrmul32_fa5_4_y2;
  wire h_u_arrmul32_fa5_4_y4;
  wire h_u_arrmul32_and6_4_y0;
  wire h_u_arrmul32_fa6_4_y2;
  wire h_u_arrmul32_fa6_4_y4;
  wire h_u_arrmul32_and7_4_y0;
  wire h_u_arrmul32_fa7_4_y2;
  wire h_u_arrmul32_fa7_4_y4;
  wire h_u_arrmul32_and8_4_y0;
  wire h_u_arrmul32_fa8_4_y2;
  wire h_u_arrmul32_fa8_4_y4;
  wire h_u_arrmul32_and9_4_y0;
  wire h_u_arrmul32_fa9_4_y2;
  wire h_u_arrmul32_fa9_4_y4;
  wire h_u_arrmul32_and10_4_y0;
  wire h_u_arrmul32_fa10_4_y2;
  wire h_u_arrmul32_fa10_4_y4;
  wire h_u_arrmul32_and11_4_y0;
  wire h_u_arrmul32_fa11_4_y2;
  wire h_u_arrmul32_fa11_4_y4;
  wire h_u_arrmul32_and12_4_y0;
  wire h_u_arrmul32_fa12_4_y2;
  wire h_u_arrmul32_fa12_4_y4;
  wire h_u_arrmul32_and13_4_y0;
  wire h_u_arrmul32_fa13_4_y2;
  wire h_u_arrmul32_fa13_4_y4;
  wire h_u_arrmul32_and14_4_y0;
  wire h_u_arrmul32_fa14_4_y2;
  wire h_u_arrmul32_fa14_4_y4;
  wire h_u_arrmul32_and15_4_y0;
  wire h_u_arrmul32_fa15_4_y2;
  wire h_u_arrmul32_fa15_4_y4;
  wire h_u_arrmul32_and16_4_y0;
  wire h_u_arrmul32_fa16_4_y2;
  wire h_u_arrmul32_fa16_4_y4;
  wire h_u_arrmul32_and17_4_y0;
  wire h_u_arrmul32_fa17_4_y2;
  wire h_u_arrmul32_fa17_4_y4;
  wire h_u_arrmul32_and18_4_y0;
  wire h_u_arrmul32_fa18_4_y2;
  wire h_u_arrmul32_fa18_4_y4;
  wire h_u_arrmul32_and19_4_y0;
  wire h_u_arrmul32_fa19_4_y2;
  wire h_u_arrmul32_fa19_4_y4;
  wire h_u_arrmul32_and20_4_y0;
  wire h_u_arrmul32_fa20_4_y2;
  wire h_u_arrmul32_fa20_4_y4;
  wire h_u_arrmul32_and21_4_y0;
  wire h_u_arrmul32_fa21_4_y2;
  wire h_u_arrmul32_fa21_4_y4;
  wire h_u_arrmul32_and22_4_y0;
  wire h_u_arrmul32_fa22_4_y2;
  wire h_u_arrmul32_fa22_4_y4;
  wire h_u_arrmul32_and23_4_y0;
  wire h_u_arrmul32_fa23_4_y2;
  wire h_u_arrmul32_fa23_4_y4;
  wire h_u_arrmul32_and24_4_y0;
  wire h_u_arrmul32_fa24_4_y2;
  wire h_u_arrmul32_fa24_4_y4;
  wire h_u_arrmul32_and25_4_y0;
  wire h_u_arrmul32_fa25_4_y2;
  wire h_u_arrmul32_fa25_4_y4;
  wire h_u_arrmul32_and26_4_y0;
  wire h_u_arrmul32_fa26_4_y2;
  wire h_u_arrmul32_fa26_4_y4;
  wire h_u_arrmul32_and27_4_y0;
  wire h_u_arrmul32_fa27_4_y2;
  wire h_u_arrmul32_fa27_4_y4;
  wire h_u_arrmul32_and28_4_y0;
  wire h_u_arrmul32_fa28_4_y2;
  wire h_u_arrmul32_fa28_4_y4;
  wire h_u_arrmul32_and29_4_y0;
  wire h_u_arrmul32_fa29_4_y2;
  wire h_u_arrmul32_fa29_4_y4;
  wire h_u_arrmul32_and30_4_y0;
  wire h_u_arrmul32_fa30_4_y2;
  wire h_u_arrmul32_fa30_4_y4;
  wire h_u_arrmul32_and31_4_y0;
  wire h_u_arrmul32_fa31_4_y2;
  wire h_u_arrmul32_fa31_4_y4;
  wire h_u_arrmul32_and0_5_y0;
  wire h_u_arrmul32_ha0_5_y0;
  wire h_u_arrmul32_ha0_5_y1;
  wire h_u_arrmul32_and1_5_y0;
  wire h_u_arrmul32_fa1_5_y2;
  wire h_u_arrmul32_fa1_5_y4;
  wire h_u_arrmul32_and2_5_y0;
  wire h_u_arrmul32_fa2_5_y2;
  wire h_u_arrmul32_fa2_5_y4;
  wire h_u_arrmul32_and3_5_y0;
  wire h_u_arrmul32_fa3_5_y2;
  wire h_u_arrmul32_fa3_5_y4;
  wire h_u_arrmul32_and4_5_y0;
  wire h_u_arrmul32_fa4_5_y2;
  wire h_u_arrmul32_fa4_5_y4;
  wire h_u_arrmul32_and5_5_y0;
  wire h_u_arrmul32_fa5_5_y2;
  wire h_u_arrmul32_fa5_5_y4;
  wire h_u_arrmul32_and6_5_y0;
  wire h_u_arrmul32_fa6_5_y2;
  wire h_u_arrmul32_fa6_5_y4;
  wire h_u_arrmul32_and7_5_y0;
  wire h_u_arrmul32_fa7_5_y2;
  wire h_u_arrmul32_fa7_5_y4;
  wire h_u_arrmul32_and8_5_y0;
  wire h_u_arrmul32_fa8_5_y2;
  wire h_u_arrmul32_fa8_5_y4;
  wire h_u_arrmul32_and9_5_y0;
  wire h_u_arrmul32_fa9_5_y2;
  wire h_u_arrmul32_fa9_5_y4;
  wire h_u_arrmul32_and10_5_y0;
  wire h_u_arrmul32_fa10_5_y2;
  wire h_u_arrmul32_fa10_5_y4;
  wire h_u_arrmul32_and11_5_y0;
  wire h_u_arrmul32_fa11_5_y2;
  wire h_u_arrmul32_fa11_5_y4;
  wire h_u_arrmul32_and12_5_y0;
  wire h_u_arrmul32_fa12_5_y2;
  wire h_u_arrmul32_fa12_5_y4;
  wire h_u_arrmul32_and13_5_y0;
  wire h_u_arrmul32_fa13_5_y2;
  wire h_u_arrmul32_fa13_5_y4;
  wire h_u_arrmul32_and14_5_y0;
  wire h_u_arrmul32_fa14_5_y2;
  wire h_u_arrmul32_fa14_5_y4;
  wire h_u_arrmul32_and15_5_y0;
  wire h_u_arrmul32_fa15_5_y2;
  wire h_u_arrmul32_fa15_5_y4;
  wire h_u_arrmul32_and16_5_y0;
  wire h_u_arrmul32_fa16_5_y2;
  wire h_u_arrmul32_fa16_5_y4;
  wire h_u_arrmul32_and17_5_y0;
  wire h_u_arrmul32_fa17_5_y2;
  wire h_u_arrmul32_fa17_5_y4;
  wire h_u_arrmul32_and18_5_y0;
  wire h_u_arrmul32_fa18_5_y2;
  wire h_u_arrmul32_fa18_5_y4;
  wire h_u_arrmul32_and19_5_y0;
  wire h_u_arrmul32_fa19_5_y2;
  wire h_u_arrmul32_fa19_5_y4;
  wire h_u_arrmul32_and20_5_y0;
  wire h_u_arrmul32_fa20_5_y2;
  wire h_u_arrmul32_fa20_5_y4;
  wire h_u_arrmul32_and21_5_y0;
  wire h_u_arrmul32_fa21_5_y2;
  wire h_u_arrmul32_fa21_5_y4;
  wire h_u_arrmul32_and22_5_y0;
  wire h_u_arrmul32_fa22_5_y2;
  wire h_u_arrmul32_fa22_5_y4;
  wire h_u_arrmul32_and23_5_y0;
  wire h_u_arrmul32_fa23_5_y2;
  wire h_u_arrmul32_fa23_5_y4;
  wire h_u_arrmul32_and24_5_y0;
  wire h_u_arrmul32_fa24_5_y2;
  wire h_u_arrmul32_fa24_5_y4;
  wire h_u_arrmul32_and25_5_y0;
  wire h_u_arrmul32_fa25_5_y2;
  wire h_u_arrmul32_fa25_5_y4;
  wire h_u_arrmul32_and26_5_y0;
  wire h_u_arrmul32_fa26_5_y2;
  wire h_u_arrmul32_fa26_5_y4;
  wire h_u_arrmul32_and27_5_y0;
  wire h_u_arrmul32_fa27_5_y2;
  wire h_u_arrmul32_fa27_5_y4;
  wire h_u_arrmul32_and28_5_y0;
  wire h_u_arrmul32_fa28_5_y2;
  wire h_u_arrmul32_fa28_5_y4;
  wire h_u_arrmul32_and29_5_y0;
  wire h_u_arrmul32_fa29_5_y2;
  wire h_u_arrmul32_fa29_5_y4;
  wire h_u_arrmul32_and30_5_y0;
  wire h_u_arrmul32_fa30_5_y2;
  wire h_u_arrmul32_fa30_5_y4;
  wire h_u_arrmul32_and31_5_y0;
  wire h_u_arrmul32_fa31_5_y2;
  wire h_u_arrmul32_fa31_5_y4;
  wire h_u_arrmul32_and0_6_y0;
  wire h_u_arrmul32_ha0_6_y0;
  wire h_u_arrmul32_ha0_6_y1;
  wire h_u_arrmul32_and1_6_y0;
  wire h_u_arrmul32_fa1_6_y2;
  wire h_u_arrmul32_fa1_6_y4;
  wire h_u_arrmul32_and2_6_y0;
  wire h_u_arrmul32_fa2_6_y2;
  wire h_u_arrmul32_fa2_6_y4;
  wire h_u_arrmul32_and3_6_y0;
  wire h_u_arrmul32_fa3_6_y2;
  wire h_u_arrmul32_fa3_6_y4;
  wire h_u_arrmul32_and4_6_y0;
  wire h_u_arrmul32_fa4_6_y2;
  wire h_u_arrmul32_fa4_6_y4;
  wire h_u_arrmul32_and5_6_y0;
  wire h_u_arrmul32_fa5_6_y2;
  wire h_u_arrmul32_fa5_6_y4;
  wire h_u_arrmul32_and6_6_y0;
  wire h_u_arrmul32_fa6_6_y2;
  wire h_u_arrmul32_fa6_6_y4;
  wire h_u_arrmul32_and7_6_y0;
  wire h_u_arrmul32_fa7_6_y2;
  wire h_u_arrmul32_fa7_6_y4;
  wire h_u_arrmul32_and8_6_y0;
  wire h_u_arrmul32_fa8_6_y2;
  wire h_u_arrmul32_fa8_6_y4;
  wire h_u_arrmul32_and9_6_y0;
  wire h_u_arrmul32_fa9_6_y2;
  wire h_u_arrmul32_fa9_6_y4;
  wire h_u_arrmul32_and10_6_y0;
  wire h_u_arrmul32_fa10_6_y2;
  wire h_u_arrmul32_fa10_6_y4;
  wire h_u_arrmul32_and11_6_y0;
  wire h_u_arrmul32_fa11_6_y2;
  wire h_u_arrmul32_fa11_6_y4;
  wire h_u_arrmul32_and12_6_y0;
  wire h_u_arrmul32_fa12_6_y2;
  wire h_u_arrmul32_fa12_6_y4;
  wire h_u_arrmul32_and13_6_y0;
  wire h_u_arrmul32_fa13_6_y2;
  wire h_u_arrmul32_fa13_6_y4;
  wire h_u_arrmul32_and14_6_y0;
  wire h_u_arrmul32_fa14_6_y2;
  wire h_u_arrmul32_fa14_6_y4;
  wire h_u_arrmul32_and15_6_y0;
  wire h_u_arrmul32_fa15_6_y2;
  wire h_u_arrmul32_fa15_6_y4;
  wire h_u_arrmul32_and16_6_y0;
  wire h_u_arrmul32_fa16_6_y2;
  wire h_u_arrmul32_fa16_6_y4;
  wire h_u_arrmul32_and17_6_y0;
  wire h_u_arrmul32_fa17_6_y2;
  wire h_u_arrmul32_fa17_6_y4;
  wire h_u_arrmul32_and18_6_y0;
  wire h_u_arrmul32_fa18_6_y2;
  wire h_u_arrmul32_fa18_6_y4;
  wire h_u_arrmul32_and19_6_y0;
  wire h_u_arrmul32_fa19_6_y2;
  wire h_u_arrmul32_fa19_6_y4;
  wire h_u_arrmul32_and20_6_y0;
  wire h_u_arrmul32_fa20_6_y2;
  wire h_u_arrmul32_fa20_6_y4;
  wire h_u_arrmul32_and21_6_y0;
  wire h_u_arrmul32_fa21_6_y2;
  wire h_u_arrmul32_fa21_6_y4;
  wire h_u_arrmul32_and22_6_y0;
  wire h_u_arrmul32_fa22_6_y2;
  wire h_u_arrmul32_fa22_6_y4;
  wire h_u_arrmul32_and23_6_y0;
  wire h_u_arrmul32_fa23_6_y2;
  wire h_u_arrmul32_fa23_6_y4;
  wire h_u_arrmul32_and24_6_y0;
  wire h_u_arrmul32_fa24_6_y2;
  wire h_u_arrmul32_fa24_6_y4;
  wire h_u_arrmul32_and25_6_y0;
  wire h_u_arrmul32_fa25_6_y2;
  wire h_u_arrmul32_fa25_6_y4;
  wire h_u_arrmul32_and26_6_y0;
  wire h_u_arrmul32_fa26_6_y2;
  wire h_u_arrmul32_fa26_6_y4;
  wire h_u_arrmul32_and27_6_y0;
  wire h_u_arrmul32_fa27_6_y2;
  wire h_u_arrmul32_fa27_6_y4;
  wire h_u_arrmul32_and28_6_y0;
  wire h_u_arrmul32_fa28_6_y2;
  wire h_u_arrmul32_fa28_6_y4;
  wire h_u_arrmul32_and29_6_y0;
  wire h_u_arrmul32_fa29_6_y2;
  wire h_u_arrmul32_fa29_6_y4;
  wire h_u_arrmul32_and30_6_y0;
  wire h_u_arrmul32_fa30_6_y2;
  wire h_u_arrmul32_fa30_6_y4;
  wire h_u_arrmul32_and31_6_y0;
  wire h_u_arrmul32_fa31_6_y2;
  wire h_u_arrmul32_fa31_6_y4;
  wire h_u_arrmul32_and0_7_y0;
  wire h_u_arrmul32_ha0_7_y0;
  wire h_u_arrmul32_ha0_7_y1;
  wire h_u_arrmul32_and1_7_y0;
  wire h_u_arrmul32_fa1_7_y2;
  wire h_u_arrmul32_fa1_7_y4;
  wire h_u_arrmul32_and2_7_y0;
  wire h_u_arrmul32_fa2_7_y2;
  wire h_u_arrmul32_fa2_7_y4;
  wire h_u_arrmul32_and3_7_y0;
  wire h_u_arrmul32_fa3_7_y2;
  wire h_u_arrmul32_fa3_7_y4;
  wire h_u_arrmul32_and4_7_y0;
  wire h_u_arrmul32_fa4_7_y2;
  wire h_u_arrmul32_fa4_7_y4;
  wire h_u_arrmul32_and5_7_y0;
  wire h_u_arrmul32_fa5_7_y2;
  wire h_u_arrmul32_fa5_7_y4;
  wire h_u_arrmul32_and6_7_y0;
  wire h_u_arrmul32_fa6_7_y2;
  wire h_u_arrmul32_fa6_7_y4;
  wire h_u_arrmul32_and7_7_y0;
  wire h_u_arrmul32_fa7_7_y2;
  wire h_u_arrmul32_fa7_7_y4;
  wire h_u_arrmul32_and8_7_y0;
  wire h_u_arrmul32_fa8_7_y2;
  wire h_u_arrmul32_fa8_7_y4;
  wire h_u_arrmul32_and9_7_y0;
  wire h_u_arrmul32_fa9_7_y2;
  wire h_u_arrmul32_fa9_7_y4;
  wire h_u_arrmul32_and10_7_y0;
  wire h_u_arrmul32_fa10_7_y2;
  wire h_u_arrmul32_fa10_7_y4;
  wire h_u_arrmul32_and11_7_y0;
  wire h_u_arrmul32_fa11_7_y2;
  wire h_u_arrmul32_fa11_7_y4;
  wire h_u_arrmul32_and12_7_y0;
  wire h_u_arrmul32_fa12_7_y2;
  wire h_u_arrmul32_fa12_7_y4;
  wire h_u_arrmul32_and13_7_y0;
  wire h_u_arrmul32_fa13_7_y2;
  wire h_u_arrmul32_fa13_7_y4;
  wire h_u_arrmul32_and14_7_y0;
  wire h_u_arrmul32_fa14_7_y2;
  wire h_u_arrmul32_fa14_7_y4;
  wire h_u_arrmul32_and15_7_y0;
  wire h_u_arrmul32_fa15_7_y2;
  wire h_u_arrmul32_fa15_7_y4;
  wire h_u_arrmul32_and16_7_y0;
  wire h_u_arrmul32_fa16_7_y2;
  wire h_u_arrmul32_fa16_7_y4;
  wire h_u_arrmul32_and17_7_y0;
  wire h_u_arrmul32_fa17_7_y2;
  wire h_u_arrmul32_fa17_7_y4;
  wire h_u_arrmul32_and18_7_y0;
  wire h_u_arrmul32_fa18_7_y2;
  wire h_u_arrmul32_fa18_7_y4;
  wire h_u_arrmul32_and19_7_y0;
  wire h_u_arrmul32_fa19_7_y2;
  wire h_u_arrmul32_fa19_7_y4;
  wire h_u_arrmul32_and20_7_y0;
  wire h_u_arrmul32_fa20_7_y2;
  wire h_u_arrmul32_fa20_7_y4;
  wire h_u_arrmul32_and21_7_y0;
  wire h_u_arrmul32_fa21_7_y2;
  wire h_u_arrmul32_fa21_7_y4;
  wire h_u_arrmul32_and22_7_y0;
  wire h_u_arrmul32_fa22_7_y2;
  wire h_u_arrmul32_fa22_7_y4;
  wire h_u_arrmul32_and23_7_y0;
  wire h_u_arrmul32_fa23_7_y2;
  wire h_u_arrmul32_fa23_7_y4;
  wire h_u_arrmul32_and24_7_y0;
  wire h_u_arrmul32_fa24_7_y2;
  wire h_u_arrmul32_fa24_7_y4;
  wire h_u_arrmul32_and25_7_y0;
  wire h_u_arrmul32_fa25_7_y2;
  wire h_u_arrmul32_fa25_7_y4;
  wire h_u_arrmul32_and26_7_y0;
  wire h_u_arrmul32_fa26_7_y2;
  wire h_u_arrmul32_fa26_7_y4;
  wire h_u_arrmul32_and27_7_y0;
  wire h_u_arrmul32_fa27_7_y2;
  wire h_u_arrmul32_fa27_7_y4;
  wire h_u_arrmul32_and28_7_y0;
  wire h_u_arrmul32_fa28_7_y2;
  wire h_u_arrmul32_fa28_7_y4;
  wire h_u_arrmul32_and29_7_y0;
  wire h_u_arrmul32_fa29_7_y2;
  wire h_u_arrmul32_fa29_7_y4;
  wire h_u_arrmul32_and30_7_y0;
  wire h_u_arrmul32_fa30_7_y2;
  wire h_u_arrmul32_fa30_7_y4;
  wire h_u_arrmul32_and31_7_y0;
  wire h_u_arrmul32_fa31_7_y2;
  wire h_u_arrmul32_fa31_7_y4;
  wire h_u_arrmul32_and0_8_y0;
  wire h_u_arrmul32_ha0_8_y0;
  wire h_u_arrmul32_ha0_8_y1;
  wire h_u_arrmul32_and1_8_y0;
  wire h_u_arrmul32_fa1_8_y2;
  wire h_u_arrmul32_fa1_8_y4;
  wire h_u_arrmul32_and2_8_y0;
  wire h_u_arrmul32_fa2_8_y2;
  wire h_u_arrmul32_fa2_8_y4;
  wire h_u_arrmul32_and3_8_y0;
  wire h_u_arrmul32_fa3_8_y2;
  wire h_u_arrmul32_fa3_8_y4;
  wire h_u_arrmul32_and4_8_y0;
  wire h_u_arrmul32_fa4_8_y2;
  wire h_u_arrmul32_fa4_8_y4;
  wire h_u_arrmul32_and5_8_y0;
  wire h_u_arrmul32_fa5_8_y2;
  wire h_u_arrmul32_fa5_8_y4;
  wire h_u_arrmul32_and6_8_y0;
  wire h_u_arrmul32_fa6_8_y2;
  wire h_u_arrmul32_fa6_8_y4;
  wire h_u_arrmul32_and7_8_y0;
  wire h_u_arrmul32_fa7_8_y2;
  wire h_u_arrmul32_fa7_8_y4;
  wire h_u_arrmul32_and8_8_y0;
  wire h_u_arrmul32_fa8_8_y2;
  wire h_u_arrmul32_fa8_8_y4;
  wire h_u_arrmul32_and9_8_y0;
  wire h_u_arrmul32_fa9_8_y2;
  wire h_u_arrmul32_fa9_8_y4;
  wire h_u_arrmul32_and10_8_y0;
  wire h_u_arrmul32_fa10_8_y2;
  wire h_u_arrmul32_fa10_8_y4;
  wire h_u_arrmul32_and11_8_y0;
  wire h_u_arrmul32_fa11_8_y2;
  wire h_u_arrmul32_fa11_8_y4;
  wire h_u_arrmul32_and12_8_y0;
  wire h_u_arrmul32_fa12_8_y2;
  wire h_u_arrmul32_fa12_8_y4;
  wire h_u_arrmul32_and13_8_y0;
  wire h_u_arrmul32_fa13_8_y2;
  wire h_u_arrmul32_fa13_8_y4;
  wire h_u_arrmul32_and14_8_y0;
  wire h_u_arrmul32_fa14_8_y2;
  wire h_u_arrmul32_fa14_8_y4;
  wire h_u_arrmul32_and15_8_y0;
  wire h_u_arrmul32_fa15_8_y2;
  wire h_u_arrmul32_fa15_8_y4;
  wire h_u_arrmul32_and16_8_y0;
  wire h_u_arrmul32_fa16_8_y2;
  wire h_u_arrmul32_fa16_8_y4;
  wire h_u_arrmul32_and17_8_y0;
  wire h_u_arrmul32_fa17_8_y2;
  wire h_u_arrmul32_fa17_8_y4;
  wire h_u_arrmul32_and18_8_y0;
  wire h_u_arrmul32_fa18_8_y2;
  wire h_u_arrmul32_fa18_8_y4;
  wire h_u_arrmul32_and19_8_y0;
  wire h_u_arrmul32_fa19_8_y2;
  wire h_u_arrmul32_fa19_8_y4;
  wire h_u_arrmul32_and20_8_y0;
  wire h_u_arrmul32_fa20_8_y2;
  wire h_u_arrmul32_fa20_8_y4;
  wire h_u_arrmul32_and21_8_y0;
  wire h_u_arrmul32_fa21_8_y2;
  wire h_u_arrmul32_fa21_8_y4;
  wire h_u_arrmul32_and22_8_y0;
  wire h_u_arrmul32_fa22_8_y2;
  wire h_u_arrmul32_fa22_8_y4;
  wire h_u_arrmul32_and23_8_y0;
  wire h_u_arrmul32_fa23_8_y2;
  wire h_u_arrmul32_fa23_8_y4;
  wire h_u_arrmul32_and24_8_y0;
  wire h_u_arrmul32_fa24_8_y2;
  wire h_u_arrmul32_fa24_8_y4;
  wire h_u_arrmul32_and25_8_y0;
  wire h_u_arrmul32_fa25_8_y2;
  wire h_u_arrmul32_fa25_8_y4;
  wire h_u_arrmul32_and26_8_y0;
  wire h_u_arrmul32_fa26_8_y2;
  wire h_u_arrmul32_fa26_8_y4;
  wire h_u_arrmul32_and27_8_y0;
  wire h_u_arrmul32_fa27_8_y2;
  wire h_u_arrmul32_fa27_8_y4;
  wire h_u_arrmul32_and28_8_y0;
  wire h_u_arrmul32_fa28_8_y2;
  wire h_u_arrmul32_fa28_8_y4;
  wire h_u_arrmul32_and29_8_y0;
  wire h_u_arrmul32_fa29_8_y2;
  wire h_u_arrmul32_fa29_8_y4;
  wire h_u_arrmul32_and30_8_y0;
  wire h_u_arrmul32_fa30_8_y2;
  wire h_u_arrmul32_fa30_8_y4;
  wire h_u_arrmul32_and31_8_y0;
  wire h_u_arrmul32_fa31_8_y2;
  wire h_u_arrmul32_fa31_8_y4;
  wire h_u_arrmul32_and0_9_y0;
  wire h_u_arrmul32_ha0_9_y0;
  wire h_u_arrmul32_ha0_9_y1;
  wire h_u_arrmul32_and1_9_y0;
  wire h_u_arrmul32_fa1_9_y2;
  wire h_u_arrmul32_fa1_9_y4;
  wire h_u_arrmul32_and2_9_y0;
  wire h_u_arrmul32_fa2_9_y2;
  wire h_u_arrmul32_fa2_9_y4;
  wire h_u_arrmul32_and3_9_y0;
  wire h_u_arrmul32_fa3_9_y2;
  wire h_u_arrmul32_fa3_9_y4;
  wire h_u_arrmul32_and4_9_y0;
  wire h_u_arrmul32_fa4_9_y2;
  wire h_u_arrmul32_fa4_9_y4;
  wire h_u_arrmul32_and5_9_y0;
  wire h_u_arrmul32_fa5_9_y2;
  wire h_u_arrmul32_fa5_9_y4;
  wire h_u_arrmul32_and6_9_y0;
  wire h_u_arrmul32_fa6_9_y2;
  wire h_u_arrmul32_fa6_9_y4;
  wire h_u_arrmul32_and7_9_y0;
  wire h_u_arrmul32_fa7_9_y2;
  wire h_u_arrmul32_fa7_9_y4;
  wire h_u_arrmul32_and8_9_y0;
  wire h_u_arrmul32_fa8_9_y2;
  wire h_u_arrmul32_fa8_9_y4;
  wire h_u_arrmul32_and9_9_y0;
  wire h_u_arrmul32_fa9_9_y2;
  wire h_u_arrmul32_fa9_9_y4;
  wire h_u_arrmul32_and10_9_y0;
  wire h_u_arrmul32_fa10_9_y2;
  wire h_u_arrmul32_fa10_9_y4;
  wire h_u_arrmul32_and11_9_y0;
  wire h_u_arrmul32_fa11_9_y2;
  wire h_u_arrmul32_fa11_9_y4;
  wire h_u_arrmul32_and12_9_y0;
  wire h_u_arrmul32_fa12_9_y2;
  wire h_u_arrmul32_fa12_9_y4;
  wire h_u_arrmul32_and13_9_y0;
  wire h_u_arrmul32_fa13_9_y2;
  wire h_u_arrmul32_fa13_9_y4;
  wire h_u_arrmul32_and14_9_y0;
  wire h_u_arrmul32_fa14_9_y2;
  wire h_u_arrmul32_fa14_9_y4;
  wire h_u_arrmul32_and15_9_y0;
  wire h_u_arrmul32_fa15_9_y2;
  wire h_u_arrmul32_fa15_9_y4;
  wire h_u_arrmul32_and16_9_y0;
  wire h_u_arrmul32_fa16_9_y2;
  wire h_u_arrmul32_fa16_9_y4;
  wire h_u_arrmul32_and17_9_y0;
  wire h_u_arrmul32_fa17_9_y2;
  wire h_u_arrmul32_fa17_9_y4;
  wire h_u_arrmul32_and18_9_y0;
  wire h_u_arrmul32_fa18_9_y2;
  wire h_u_arrmul32_fa18_9_y4;
  wire h_u_arrmul32_and19_9_y0;
  wire h_u_arrmul32_fa19_9_y2;
  wire h_u_arrmul32_fa19_9_y4;
  wire h_u_arrmul32_and20_9_y0;
  wire h_u_arrmul32_fa20_9_y2;
  wire h_u_arrmul32_fa20_9_y4;
  wire h_u_arrmul32_and21_9_y0;
  wire h_u_arrmul32_fa21_9_y2;
  wire h_u_arrmul32_fa21_9_y4;
  wire h_u_arrmul32_and22_9_y0;
  wire h_u_arrmul32_fa22_9_y2;
  wire h_u_arrmul32_fa22_9_y4;
  wire h_u_arrmul32_and23_9_y0;
  wire h_u_arrmul32_fa23_9_y2;
  wire h_u_arrmul32_fa23_9_y4;
  wire h_u_arrmul32_and24_9_y0;
  wire h_u_arrmul32_fa24_9_y2;
  wire h_u_arrmul32_fa24_9_y4;
  wire h_u_arrmul32_and25_9_y0;
  wire h_u_arrmul32_fa25_9_y2;
  wire h_u_arrmul32_fa25_9_y4;
  wire h_u_arrmul32_and26_9_y0;
  wire h_u_arrmul32_fa26_9_y2;
  wire h_u_arrmul32_fa26_9_y4;
  wire h_u_arrmul32_and27_9_y0;
  wire h_u_arrmul32_fa27_9_y2;
  wire h_u_arrmul32_fa27_9_y4;
  wire h_u_arrmul32_and28_9_y0;
  wire h_u_arrmul32_fa28_9_y2;
  wire h_u_arrmul32_fa28_9_y4;
  wire h_u_arrmul32_and29_9_y0;
  wire h_u_arrmul32_fa29_9_y2;
  wire h_u_arrmul32_fa29_9_y4;
  wire h_u_arrmul32_and30_9_y0;
  wire h_u_arrmul32_fa30_9_y2;
  wire h_u_arrmul32_fa30_9_y4;
  wire h_u_arrmul32_and31_9_y0;
  wire h_u_arrmul32_fa31_9_y2;
  wire h_u_arrmul32_fa31_9_y4;
  wire h_u_arrmul32_and0_10_y0;
  wire h_u_arrmul32_ha0_10_y0;
  wire h_u_arrmul32_ha0_10_y1;
  wire h_u_arrmul32_and1_10_y0;
  wire h_u_arrmul32_fa1_10_y2;
  wire h_u_arrmul32_fa1_10_y4;
  wire h_u_arrmul32_and2_10_y0;
  wire h_u_arrmul32_fa2_10_y2;
  wire h_u_arrmul32_fa2_10_y4;
  wire h_u_arrmul32_and3_10_y0;
  wire h_u_arrmul32_fa3_10_y2;
  wire h_u_arrmul32_fa3_10_y4;
  wire h_u_arrmul32_and4_10_y0;
  wire h_u_arrmul32_fa4_10_y2;
  wire h_u_arrmul32_fa4_10_y4;
  wire h_u_arrmul32_and5_10_y0;
  wire h_u_arrmul32_fa5_10_y2;
  wire h_u_arrmul32_fa5_10_y4;
  wire h_u_arrmul32_and6_10_y0;
  wire h_u_arrmul32_fa6_10_y2;
  wire h_u_arrmul32_fa6_10_y4;
  wire h_u_arrmul32_and7_10_y0;
  wire h_u_arrmul32_fa7_10_y2;
  wire h_u_arrmul32_fa7_10_y4;
  wire h_u_arrmul32_and8_10_y0;
  wire h_u_arrmul32_fa8_10_y2;
  wire h_u_arrmul32_fa8_10_y4;
  wire h_u_arrmul32_and9_10_y0;
  wire h_u_arrmul32_fa9_10_y2;
  wire h_u_arrmul32_fa9_10_y4;
  wire h_u_arrmul32_and10_10_y0;
  wire h_u_arrmul32_fa10_10_y2;
  wire h_u_arrmul32_fa10_10_y4;
  wire h_u_arrmul32_and11_10_y0;
  wire h_u_arrmul32_fa11_10_y2;
  wire h_u_arrmul32_fa11_10_y4;
  wire h_u_arrmul32_and12_10_y0;
  wire h_u_arrmul32_fa12_10_y2;
  wire h_u_arrmul32_fa12_10_y4;
  wire h_u_arrmul32_and13_10_y0;
  wire h_u_arrmul32_fa13_10_y2;
  wire h_u_arrmul32_fa13_10_y4;
  wire h_u_arrmul32_and14_10_y0;
  wire h_u_arrmul32_fa14_10_y2;
  wire h_u_arrmul32_fa14_10_y4;
  wire h_u_arrmul32_and15_10_y0;
  wire h_u_arrmul32_fa15_10_y2;
  wire h_u_arrmul32_fa15_10_y4;
  wire h_u_arrmul32_and16_10_y0;
  wire h_u_arrmul32_fa16_10_y2;
  wire h_u_arrmul32_fa16_10_y4;
  wire h_u_arrmul32_and17_10_y0;
  wire h_u_arrmul32_fa17_10_y2;
  wire h_u_arrmul32_fa17_10_y4;
  wire h_u_arrmul32_and18_10_y0;
  wire h_u_arrmul32_fa18_10_y2;
  wire h_u_arrmul32_fa18_10_y4;
  wire h_u_arrmul32_and19_10_y0;
  wire h_u_arrmul32_fa19_10_y2;
  wire h_u_arrmul32_fa19_10_y4;
  wire h_u_arrmul32_and20_10_y0;
  wire h_u_arrmul32_fa20_10_y2;
  wire h_u_arrmul32_fa20_10_y4;
  wire h_u_arrmul32_and21_10_y0;
  wire h_u_arrmul32_fa21_10_y2;
  wire h_u_arrmul32_fa21_10_y4;
  wire h_u_arrmul32_and22_10_y0;
  wire h_u_arrmul32_fa22_10_y2;
  wire h_u_arrmul32_fa22_10_y4;
  wire h_u_arrmul32_and23_10_y0;
  wire h_u_arrmul32_fa23_10_y2;
  wire h_u_arrmul32_fa23_10_y4;
  wire h_u_arrmul32_and24_10_y0;
  wire h_u_arrmul32_fa24_10_y2;
  wire h_u_arrmul32_fa24_10_y4;
  wire h_u_arrmul32_and25_10_y0;
  wire h_u_arrmul32_fa25_10_y2;
  wire h_u_arrmul32_fa25_10_y4;
  wire h_u_arrmul32_and26_10_y0;
  wire h_u_arrmul32_fa26_10_y2;
  wire h_u_arrmul32_fa26_10_y4;
  wire h_u_arrmul32_and27_10_y0;
  wire h_u_arrmul32_fa27_10_y2;
  wire h_u_arrmul32_fa27_10_y4;
  wire h_u_arrmul32_and28_10_y0;
  wire h_u_arrmul32_fa28_10_y2;
  wire h_u_arrmul32_fa28_10_y4;
  wire h_u_arrmul32_and29_10_y0;
  wire h_u_arrmul32_fa29_10_y2;
  wire h_u_arrmul32_fa29_10_y4;
  wire h_u_arrmul32_and30_10_y0;
  wire h_u_arrmul32_fa30_10_y2;
  wire h_u_arrmul32_fa30_10_y4;
  wire h_u_arrmul32_and31_10_y0;
  wire h_u_arrmul32_fa31_10_y2;
  wire h_u_arrmul32_fa31_10_y4;
  wire h_u_arrmul32_and0_11_y0;
  wire h_u_arrmul32_ha0_11_y0;
  wire h_u_arrmul32_ha0_11_y1;
  wire h_u_arrmul32_and1_11_y0;
  wire h_u_arrmul32_fa1_11_y2;
  wire h_u_arrmul32_fa1_11_y4;
  wire h_u_arrmul32_and2_11_y0;
  wire h_u_arrmul32_fa2_11_y2;
  wire h_u_arrmul32_fa2_11_y4;
  wire h_u_arrmul32_and3_11_y0;
  wire h_u_arrmul32_fa3_11_y2;
  wire h_u_arrmul32_fa3_11_y4;
  wire h_u_arrmul32_and4_11_y0;
  wire h_u_arrmul32_fa4_11_y2;
  wire h_u_arrmul32_fa4_11_y4;
  wire h_u_arrmul32_and5_11_y0;
  wire h_u_arrmul32_fa5_11_y2;
  wire h_u_arrmul32_fa5_11_y4;
  wire h_u_arrmul32_and6_11_y0;
  wire h_u_arrmul32_fa6_11_y2;
  wire h_u_arrmul32_fa6_11_y4;
  wire h_u_arrmul32_and7_11_y0;
  wire h_u_arrmul32_fa7_11_y2;
  wire h_u_arrmul32_fa7_11_y4;
  wire h_u_arrmul32_and8_11_y0;
  wire h_u_arrmul32_fa8_11_y2;
  wire h_u_arrmul32_fa8_11_y4;
  wire h_u_arrmul32_and9_11_y0;
  wire h_u_arrmul32_fa9_11_y2;
  wire h_u_arrmul32_fa9_11_y4;
  wire h_u_arrmul32_and10_11_y0;
  wire h_u_arrmul32_fa10_11_y2;
  wire h_u_arrmul32_fa10_11_y4;
  wire h_u_arrmul32_and11_11_y0;
  wire h_u_arrmul32_fa11_11_y2;
  wire h_u_arrmul32_fa11_11_y4;
  wire h_u_arrmul32_and12_11_y0;
  wire h_u_arrmul32_fa12_11_y2;
  wire h_u_arrmul32_fa12_11_y4;
  wire h_u_arrmul32_and13_11_y0;
  wire h_u_arrmul32_fa13_11_y2;
  wire h_u_arrmul32_fa13_11_y4;
  wire h_u_arrmul32_and14_11_y0;
  wire h_u_arrmul32_fa14_11_y2;
  wire h_u_arrmul32_fa14_11_y4;
  wire h_u_arrmul32_and15_11_y0;
  wire h_u_arrmul32_fa15_11_y2;
  wire h_u_arrmul32_fa15_11_y4;
  wire h_u_arrmul32_and16_11_y0;
  wire h_u_arrmul32_fa16_11_y2;
  wire h_u_arrmul32_fa16_11_y4;
  wire h_u_arrmul32_and17_11_y0;
  wire h_u_arrmul32_fa17_11_y2;
  wire h_u_arrmul32_fa17_11_y4;
  wire h_u_arrmul32_and18_11_y0;
  wire h_u_arrmul32_fa18_11_y2;
  wire h_u_arrmul32_fa18_11_y4;
  wire h_u_arrmul32_and19_11_y0;
  wire h_u_arrmul32_fa19_11_y2;
  wire h_u_arrmul32_fa19_11_y4;
  wire h_u_arrmul32_and20_11_y0;
  wire h_u_arrmul32_fa20_11_y2;
  wire h_u_arrmul32_fa20_11_y4;
  wire h_u_arrmul32_and21_11_y0;
  wire h_u_arrmul32_fa21_11_y2;
  wire h_u_arrmul32_fa21_11_y4;
  wire h_u_arrmul32_and22_11_y0;
  wire h_u_arrmul32_fa22_11_y2;
  wire h_u_arrmul32_fa22_11_y4;
  wire h_u_arrmul32_and23_11_y0;
  wire h_u_arrmul32_fa23_11_y2;
  wire h_u_arrmul32_fa23_11_y4;
  wire h_u_arrmul32_and24_11_y0;
  wire h_u_arrmul32_fa24_11_y2;
  wire h_u_arrmul32_fa24_11_y4;
  wire h_u_arrmul32_and25_11_y0;
  wire h_u_arrmul32_fa25_11_y2;
  wire h_u_arrmul32_fa25_11_y4;
  wire h_u_arrmul32_and26_11_y0;
  wire h_u_arrmul32_fa26_11_y2;
  wire h_u_arrmul32_fa26_11_y4;
  wire h_u_arrmul32_and27_11_y0;
  wire h_u_arrmul32_fa27_11_y2;
  wire h_u_arrmul32_fa27_11_y4;
  wire h_u_arrmul32_and28_11_y0;
  wire h_u_arrmul32_fa28_11_y2;
  wire h_u_arrmul32_fa28_11_y4;
  wire h_u_arrmul32_and29_11_y0;
  wire h_u_arrmul32_fa29_11_y2;
  wire h_u_arrmul32_fa29_11_y4;
  wire h_u_arrmul32_and30_11_y0;
  wire h_u_arrmul32_fa30_11_y2;
  wire h_u_arrmul32_fa30_11_y4;
  wire h_u_arrmul32_and31_11_y0;
  wire h_u_arrmul32_fa31_11_y2;
  wire h_u_arrmul32_fa31_11_y4;
  wire h_u_arrmul32_and0_12_y0;
  wire h_u_arrmul32_ha0_12_y0;
  wire h_u_arrmul32_ha0_12_y1;
  wire h_u_arrmul32_and1_12_y0;
  wire h_u_arrmul32_fa1_12_y2;
  wire h_u_arrmul32_fa1_12_y4;
  wire h_u_arrmul32_and2_12_y0;
  wire h_u_arrmul32_fa2_12_y2;
  wire h_u_arrmul32_fa2_12_y4;
  wire h_u_arrmul32_and3_12_y0;
  wire h_u_arrmul32_fa3_12_y2;
  wire h_u_arrmul32_fa3_12_y4;
  wire h_u_arrmul32_and4_12_y0;
  wire h_u_arrmul32_fa4_12_y2;
  wire h_u_arrmul32_fa4_12_y4;
  wire h_u_arrmul32_and5_12_y0;
  wire h_u_arrmul32_fa5_12_y2;
  wire h_u_arrmul32_fa5_12_y4;
  wire h_u_arrmul32_and6_12_y0;
  wire h_u_arrmul32_fa6_12_y2;
  wire h_u_arrmul32_fa6_12_y4;
  wire h_u_arrmul32_and7_12_y0;
  wire h_u_arrmul32_fa7_12_y2;
  wire h_u_arrmul32_fa7_12_y4;
  wire h_u_arrmul32_and8_12_y0;
  wire h_u_arrmul32_fa8_12_y2;
  wire h_u_arrmul32_fa8_12_y4;
  wire h_u_arrmul32_and9_12_y0;
  wire h_u_arrmul32_fa9_12_y2;
  wire h_u_arrmul32_fa9_12_y4;
  wire h_u_arrmul32_and10_12_y0;
  wire h_u_arrmul32_fa10_12_y2;
  wire h_u_arrmul32_fa10_12_y4;
  wire h_u_arrmul32_and11_12_y0;
  wire h_u_arrmul32_fa11_12_y2;
  wire h_u_arrmul32_fa11_12_y4;
  wire h_u_arrmul32_and12_12_y0;
  wire h_u_arrmul32_fa12_12_y2;
  wire h_u_arrmul32_fa12_12_y4;
  wire h_u_arrmul32_and13_12_y0;
  wire h_u_arrmul32_fa13_12_y2;
  wire h_u_arrmul32_fa13_12_y4;
  wire h_u_arrmul32_and14_12_y0;
  wire h_u_arrmul32_fa14_12_y2;
  wire h_u_arrmul32_fa14_12_y4;
  wire h_u_arrmul32_and15_12_y0;
  wire h_u_arrmul32_fa15_12_y2;
  wire h_u_arrmul32_fa15_12_y4;
  wire h_u_arrmul32_and16_12_y0;
  wire h_u_arrmul32_fa16_12_y2;
  wire h_u_arrmul32_fa16_12_y4;
  wire h_u_arrmul32_and17_12_y0;
  wire h_u_arrmul32_fa17_12_y2;
  wire h_u_arrmul32_fa17_12_y4;
  wire h_u_arrmul32_and18_12_y0;
  wire h_u_arrmul32_fa18_12_y2;
  wire h_u_arrmul32_fa18_12_y4;
  wire h_u_arrmul32_and19_12_y0;
  wire h_u_arrmul32_fa19_12_y2;
  wire h_u_arrmul32_fa19_12_y4;
  wire h_u_arrmul32_and20_12_y0;
  wire h_u_arrmul32_fa20_12_y2;
  wire h_u_arrmul32_fa20_12_y4;
  wire h_u_arrmul32_and21_12_y0;
  wire h_u_arrmul32_fa21_12_y2;
  wire h_u_arrmul32_fa21_12_y4;
  wire h_u_arrmul32_and22_12_y0;
  wire h_u_arrmul32_fa22_12_y2;
  wire h_u_arrmul32_fa22_12_y4;
  wire h_u_arrmul32_and23_12_y0;
  wire h_u_arrmul32_fa23_12_y2;
  wire h_u_arrmul32_fa23_12_y4;
  wire h_u_arrmul32_and24_12_y0;
  wire h_u_arrmul32_fa24_12_y2;
  wire h_u_arrmul32_fa24_12_y4;
  wire h_u_arrmul32_and25_12_y0;
  wire h_u_arrmul32_fa25_12_y2;
  wire h_u_arrmul32_fa25_12_y4;
  wire h_u_arrmul32_and26_12_y0;
  wire h_u_arrmul32_fa26_12_y2;
  wire h_u_arrmul32_fa26_12_y4;
  wire h_u_arrmul32_and27_12_y0;
  wire h_u_arrmul32_fa27_12_y2;
  wire h_u_arrmul32_fa27_12_y4;
  wire h_u_arrmul32_and28_12_y0;
  wire h_u_arrmul32_fa28_12_y2;
  wire h_u_arrmul32_fa28_12_y4;
  wire h_u_arrmul32_and29_12_y0;
  wire h_u_arrmul32_fa29_12_y2;
  wire h_u_arrmul32_fa29_12_y4;
  wire h_u_arrmul32_and30_12_y0;
  wire h_u_arrmul32_fa30_12_y2;
  wire h_u_arrmul32_fa30_12_y4;
  wire h_u_arrmul32_and31_12_y0;
  wire h_u_arrmul32_fa31_12_y2;
  wire h_u_arrmul32_fa31_12_y4;
  wire h_u_arrmul32_and0_13_y0;
  wire h_u_arrmul32_ha0_13_y0;
  wire h_u_arrmul32_ha0_13_y1;
  wire h_u_arrmul32_and1_13_y0;
  wire h_u_arrmul32_fa1_13_y2;
  wire h_u_arrmul32_fa1_13_y4;
  wire h_u_arrmul32_and2_13_y0;
  wire h_u_arrmul32_fa2_13_y2;
  wire h_u_arrmul32_fa2_13_y4;
  wire h_u_arrmul32_and3_13_y0;
  wire h_u_arrmul32_fa3_13_y2;
  wire h_u_arrmul32_fa3_13_y4;
  wire h_u_arrmul32_and4_13_y0;
  wire h_u_arrmul32_fa4_13_y2;
  wire h_u_arrmul32_fa4_13_y4;
  wire h_u_arrmul32_and5_13_y0;
  wire h_u_arrmul32_fa5_13_y2;
  wire h_u_arrmul32_fa5_13_y4;
  wire h_u_arrmul32_and6_13_y0;
  wire h_u_arrmul32_fa6_13_y2;
  wire h_u_arrmul32_fa6_13_y4;
  wire h_u_arrmul32_and7_13_y0;
  wire h_u_arrmul32_fa7_13_y2;
  wire h_u_arrmul32_fa7_13_y4;
  wire h_u_arrmul32_and8_13_y0;
  wire h_u_arrmul32_fa8_13_y2;
  wire h_u_arrmul32_fa8_13_y4;
  wire h_u_arrmul32_and9_13_y0;
  wire h_u_arrmul32_fa9_13_y2;
  wire h_u_arrmul32_fa9_13_y4;
  wire h_u_arrmul32_and10_13_y0;
  wire h_u_arrmul32_fa10_13_y2;
  wire h_u_arrmul32_fa10_13_y4;
  wire h_u_arrmul32_and11_13_y0;
  wire h_u_arrmul32_fa11_13_y2;
  wire h_u_arrmul32_fa11_13_y4;
  wire h_u_arrmul32_and12_13_y0;
  wire h_u_arrmul32_fa12_13_y2;
  wire h_u_arrmul32_fa12_13_y4;
  wire h_u_arrmul32_and13_13_y0;
  wire h_u_arrmul32_fa13_13_y2;
  wire h_u_arrmul32_fa13_13_y4;
  wire h_u_arrmul32_and14_13_y0;
  wire h_u_arrmul32_fa14_13_y2;
  wire h_u_arrmul32_fa14_13_y4;
  wire h_u_arrmul32_and15_13_y0;
  wire h_u_arrmul32_fa15_13_y2;
  wire h_u_arrmul32_fa15_13_y4;
  wire h_u_arrmul32_and16_13_y0;
  wire h_u_arrmul32_fa16_13_y2;
  wire h_u_arrmul32_fa16_13_y4;
  wire h_u_arrmul32_and17_13_y0;
  wire h_u_arrmul32_fa17_13_y2;
  wire h_u_arrmul32_fa17_13_y4;
  wire h_u_arrmul32_and18_13_y0;
  wire h_u_arrmul32_fa18_13_y2;
  wire h_u_arrmul32_fa18_13_y4;
  wire h_u_arrmul32_and19_13_y0;
  wire h_u_arrmul32_fa19_13_y2;
  wire h_u_arrmul32_fa19_13_y4;
  wire h_u_arrmul32_and20_13_y0;
  wire h_u_arrmul32_fa20_13_y2;
  wire h_u_arrmul32_fa20_13_y4;
  wire h_u_arrmul32_and21_13_y0;
  wire h_u_arrmul32_fa21_13_y2;
  wire h_u_arrmul32_fa21_13_y4;
  wire h_u_arrmul32_and22_13_y0;
  wire h_u_arrmul32_fa22_13_y2;
  wire h_u_arrmul32_fa22_13_y4;
  wire h_u_arrmul32_and23_13_y0;
  wire h_u_arrmul32_fa23_13_y2;
  wire h_u_arrmul32_fa23_13_y4;
  wire h_u_arrmul32_and24_13_y0;
  wire h_u_arrmul32_fa24_13_y2;
  wire h_u_arrmul32_fa24_13_y4;
  wire h_u_arrmul32_and25_13_y0;
  wire h_u_arrmul32_fa25_13_y2;
  wire h_u_arrmul32_fa25_13_y4;
  wire h_u_arrmul32_and26_13_y0;
  wire h_u_arrmul32_fa26_13_y2;
  wire h_u_arrmul32_fa26_13_y4;
  wire h_u_arrmul32_and27_13_y0;
  wire h_u_arrmul32_fa27_13_y2;
  wire h_u_arrmul32_fa27_13_y4;
  wire h_u_arrmul32_and28_13_y0;
  wire h_u_arrmul32_fa28_13_y2;
  wire h_u_arrmul32_fa28_13_y4;
  wire h_u_arrmul32_and29_13_y0;
  wire h_u_arrmul32_fa29_13_y2;
  wire h_u_arrmul32_fa29_13_y4;
  wire h_u_arrmul32_and30_13_y0;
  wire h_u_arrmul32_fa30_13_y2;
  wire h_u_arrmul32_fa30_13_y4;
  wire h_u_arrmul32_and31_13_y0;
  wire h_u_arrmul32_fa31_13_y2;
  wire h_u_arrmul32_fa31_13_y4;
  wire h_u_arrmul32_and0_14_y0;
  wire h_u_arrmul32_ha0_14_y0;
  wire h_u_arrmul32_ha0_14_y1;
  wire h_u_arrmul32_and1_14_y0;
  wire h_u_arrmul32_fa1_14_y2;
  wire h_u_arrmul32_fa1_14_y4;
  wire h_u_arrmul32_and2_14_y0;
  wire h_u_arrmul32_fa2_14_y2;
  wire h_u_arrmul32_fa2_14_y4;
  wire h_u_arrmul32_and3_14_y0;
  wire h_u_arrmul32_fa3_14_y2;
  wire h_u_arrmul32_fa3_14_y4;
  wire h_u_arrmul32_and4_14_y0;
  wire h_u_arrmul32_fa4_14_y2;
  wire h_u_arrmul32_fa4_14_y4;
  wire h_u_arrmul32_and5_14_y0;
  wire h_u_arrmul32_fa5_14_y2;
  wire h_u_arrmul32_fa5_14_y4;
  wire h_u_arrmul32_and6_14_y0;
  wire h_u_arrmul32_fa6_14_y2;
  wire h_u_arrmul32_fa6_14_y4;
  wire h_u_arrmul32_and7_14_y0;
  wire h_u_arrmul32_fa7_14_y2;
  wire h_u_arrmul32_fa7_14_y4;
  wire h_u_arrmul32_and8_14_y0;
  wire h_u_arrmul32_fa8_14_y2;
  wire h_u_arrmul32_fa8_14_y4;
  wire h_u_arrmul32_and9_14_y0;
  wire h_u_arrmul32_fa9_14_y2;
  wire h_u_arrmul32_fa9_14_y4;
  wire h_u_arrmul32_and10_14_y0;
  wire h_u_arrmul32_fa10_14_y2;
  wire h_u_arrmul32_fa10_14_y4;
  wire h_u_arrmul32_and11_14_y0;
  wire h_u_arrmul32_fa11_14_y2;
  wire h_u_arrmul32_fa11_14_y4;
  wire h_u_arrmul32_and12_14_y0;
  wire h_u_arrmul32_fa12_14_y2;
  wire h_u_arrmul32_fa12_14_y4;
  wire h_u_arrmul32_and13_14_y0;
  wire h_u_arrmul32_fa13_14_y2;
  wire h_u_arrmul32_fa13_14_y4;
  wire h_u_arrmul32_and14_14_y0;
  wire h_u_arrmul32_fa14_14_y2;
  wire h_u_arrmul32_fa14_14_y4;
  wire h_u_arrmul32_and15_14_y0;
  wire h_u_arrmul32_fa15_14_y2;
  wire h_u_arrmul32_fa15_14_y4;
  wire h_u_arrmul32_and16_14_y0;
  wire h_u_arrmul32_fa16_14_y2;
  wire h_u_arrmul32_fa16_14_y4;
  wire h_u_arrmul32_and17_14_y0;
  wire h_u_arrmul32_fa17_14_y2;
  wire h_u_arrmul32_fa17_14_y4;
  wire h_u_arrmul32_and18_14_y0;
  wire h_u_arrmul32_fa18_14_y2;
  wire h_u_arrmul32_fa18_14_y4;
  wire h_u_arrmul32_and19_14_y0;
  wire h_u_arrmul32_fa19_14_y2;
  wire h_u_arrmul32_fa19_14_y4;
  wire h_u_arrmul32_and20_14_y0;
  wire h_u_arrmul32_fa20_14_y2;
  wire h_u_arrmul32_fa20_14_y4;
  wire h_u_arrmul32_and21_14_y0;
  wire h_u_arrmul32_fa21_14_y2;
  wire h_u_arrmul32_fa21_14_y4;
  wire h_u_arrmul32_and22_14_y0;
  wire h_u_arrmul32_fa22_14_y2;
  wire h_u_arrmul32_fa22_14_y4;
  wire h_u_arrmul32_and23_14_y0;
  wire h_u_arrmul32_fa23_14_y2;
  wire h_u_arrmul32_fa23_14_y4;
  wire h_u_arrmul32_and24_14_y0;
  wire h_u_arrmul32_fa24_14_y2;
  wire h_u_arrmul32_fa24_14_y4;
  wire h_u_arrmul32_and25_14_y0;
  wire h_u_arrmul32_fa25_14_y2;
  wire h_u_arrmul32_fa25_14_y4;
  wire h_u_arrmul32_and26_14_y0;
  wire h_u_arrmul32_fa26_14_y2;
  wire h_u_arrmul32_fa26_14_y4;
  wire h_u_arrmul32_and27_14_y0;
  wire h_u_arrmul32_fa27_14_y2;
  wire h_u_arrmul32_fa27_14_y4;
  wire h_u_arrmul32_and28_14_y0;
  wire h_u_arrmul32_fa28_14_y2;
  wire h_u_arrmul32_fa28_14_y4;
  wire h_u_arrmul32_and29_14_y0;
  wire h_u_arrmul32_fa29_14_y2;
  wire h_u_arrmul32_fa29_14_y4;
  wire h_u_arrmul32_and30_14_y0;
  wire h_u_arrmul32_fa30_14_y2;
  wire h_u_arrmul32_fa30_14_y4;
  wire h_u_arrmul32_and31_14_y0;
  wire h_u_arrmul32_fa31_14_y2;
  wire h_u_arrmul32_fa31_14_y4;
  wire h_u_arrmul32_and0_15_y0;
  wire h_u_arrmul32_ha0_15_y0;
  wire h_u_arrmul32_ha0_15_y1;
  wire h_u_arrmul32_and1_15_y0;
  wire h_u_arrmul32_fa1_15_y2;
  wire h_u_arrmul32_fa1_15_y4;
  wire h_u_arrmul32_and2_15_y0;
  wire h_u_arrmul32_fa2_15_y2;
  wire h_u_arrmul32_fa2_15_y4;
  wire h_u_arrmul32_and3_15_y0;
  wire h_u_arrmul32_fa3_15_y2;
  wire h_u_arrmul32_fa3_15_y4;
  wire h_u_arrmul32_and4_15_y0;
  wire h_u_arrmul32_fa4_15_y2;
  wire h_u_arrmul32_fa4_15_y4;
  wire h_u_arrmul32_and5_15_y0;
  wire h_u_arrmul32_fa5_15_y2;
  wire h_u_arrmul32_fa5_15_y4;
  wire h_u_arrmul32_and6_15_y0;
  wire h_u_arrmul32_fa6_15_y2;
  wire h_u_arrmul32_fa6_15_y4;
  wire h_u_arrmul32_and7_15_y0;
  wire h_u_arrmul32_fa7_15_y2;
  wire h_u_arrmul32_fa7_15_y4;
  wire h_u_arrmul32_and8_15_y0;
  wire h_u_arrmul32_fa8_15_y2;
  wire h_u_arrmul32_fa8_15_y4;
  wire h_u_arrmul32_and9_15_y0;
  wire h_u_arrmul32_fa9_15_y2;
  wire h_u_arrmul32_fa9_15_y4;
  wire h_u_arrmul32_and10_15_y0;
  wire h_u_arrmul32_fa10_15_y2;
  wire h_u_arrmul32_fa10_15_y4;
  wire h_u_arrmul32_and11_15_y0;
  wire h_u_arrmul32_fa11_15_y2;
  wire h_u_arrmul32_fa11_15_y4;
  wire h_u_arrmul32_and12_15_y0;
  wire h_u_arrmul32_fa12_15_y2;
  wire h_u_arrmul32_fa12_15_y4;
  wire h_u_arrmul32_and13_15_y0;
  wire h_u_arrmul32_fa13_15_y2;
  wire h_u_arrmul32_fa13_15_y4;
  wire h_u_arrmul32_and14_15_y0;
  wire h_u_arrmul32_fa14_15_y2;
  wire h_u_arrmul32_fa14_15_y4;
  wire h_u_arrmul32_and15_15_y0;
  wire h_u_arrmul32_fa15_15_y2;
  wire h_u_arrmul32_fa15_15_y4;
  wire h_u_arrmul32_and16_15_y0;
  wire h_u_arrmul32_fa16_15_y2;
  wire h_u_arrmul32_fa16_15_y4;
  wire h_u_arrmul32_and17_15_y0;
  wire h_u_arrmul32_fa17_15_y2;
  wire h_u_arrmul32_fa17_15_y4;
  wire h_u_arrmul32_and18_15_y0;
  wire h_u_arrmul32_fa18_15_y2;
  wire h_u_arrmul32_fa18_15_y4;
  wire h_u_arrmul32_and19_15_y0;
  wire h_u_arrmul32_fa19_15_y2;
  wire h_u_arrmul32_fa19_15_y4;
  wire h_u_arrmul32_and20_15_y0;
  wire h_u_arrmul32_fa20_15_y2;
  wire h_u_arrmul32_fa20_15_y4;
  wire h_u_arrmul32_and21_15_y0;
  wire h_u_arrmul32_fa21_15_y2;
  wire h_u_arrmul32_fa21_15_y4;
  wire h_u_arrmul32_and22_15_y0;
  wire h_u_arrmul32_fa22_15_y2;
  wire h_u_arrmul32_fa22_15_y4;
  wire h_u_arrmul32_and23_15_y0;
  wire h_u_arrmul32_fa23_15_y2;
  wire h_u_arrmul32_fa23_15_y4;
  wire h_u_arrmul32_and24_15_y0;
  wire h_u_arrmul32_fa24_15_y2;
  wire h_u_arrmul32_fa24_15_y4;
  wire h_u_arrmul32_and25_15_y0;
  wire h_u_arrmul32_fa25_15_y2;
  wire h_u_arrmul32_fa25_15_y4;
  wire h_u_arrmul32_and26_15_y0;
  wire h_u_arrmul32_fa26_15_y2;
  wire h_u_arrmul32_fa26_15_y4;
  wire h_u_arrmul32_and27_15_y0;
  wire h_u_arrmul32_fa27_15_y2;
  wire h_u_arrmul32_fa27_15_y4;
  wire h_u_arrmul32_and28_15_y0;
  wire h_u_arrmul32_fa28_15_y2;
  wire h_u_arrmul32_fa28_15_y4;
  wire h_u_arrmul32_and29_15_y0;
  wire h_u_arrmul32_fa29_15_y2;
  wire h_u_arrmul32_fa29_15_y4;
  wire h_u_arrmul32_and30_15_y0;
  wire h_u_arrmul32_fa30_15_y2;
  wire h_u_arrmul32_fa30_15_y4;
  wire h_u_arrmul32_and31_15_y0;
  wire h_u_arrmul32_fa31_15_y2;
  wire h_u_arrmul32_fa31_15_y4;
  wire h_u_arrmul32_and0_16_y0;
  wire h_u_arrmul32_ha0_16_y0;
  wire h_u_arrmul32_ha0_16_y1;
  wire h_u_arrmul32_and1_16_y0;
  wire h_u_arrmul32_fa1_16_y2;
  wire h_u_arrmul32_fa1_16_y4;
  wire h_u_arrmul32_and2_16_y0;
  wire h_u_arrmul32_fa2_16_y2;
  wire h_u_arrmul32_fa2_16_y4;
  wire h_u_arrmul32_and3_16_y0;
  wire h_u_arrmul32_fa3_16_y2;
  wire h_u_arrmul32_fa3_16_y4;
  wire h_u_arrmul32_and4_16_y0;
  wire h_u_arrmul32_fa4_16_y2;
  wire h_u_arrmul32_fa4_16_y4;
  wire h_u_arrmul32_and5_16_y0;
  wire h_u_arrmul32_fa5_16_y2;
  wire h_u_arrmul32_fa5_16_y4;
  wire h_u_arrmul32_and6_16_y0;
  wire h_u_arrmul32_fa6_16_y2;
  wire h_u_arrmul32_fa6_16_y4;
  wire h_u_arrmul32_and7_16_y0;
  wire h_u_arrmul32_fa7_16_y2;
  wire h_u_arrmul32_fa7_16_y4;
  wire h_u_arrmul32_and8_16_y0;
  wire h_u_arrmul32_fa8_16_y2;
  wire h_u_arrmul32_fa8_16_y4;
  wire h_u_arrmul32_and9_16_y0;
  wire h_u_arrmul32_fa9_16_y2;
  wire h_u_arrmul32_fa9_16_y4;
  wire h_u_arrmul32_and10_16_y0;
  wire h_u_arrmul32_fa10_16_y2;
  wire h_u_arrmul32_fa10_16_y4;
  wire h_u_arrmul32_and11_16_y0;
  wire h_u_arrmul32_fa11_16_y2;
  wire h_u_arrmul32_fa11_16_y4;
  wire h_u_arrmul32_and12_16_y0;
  wire h_u_arrmul32_fa12_16_y2;
  wire h_u_arrmul32_fa12_16_y4;
  wire h_u_arrmul32_and13_16_y0;
  wire h_u_arrmul32_fa13_16_y2;
  wire h_u_arrmul32_fa13_16_y4;
  wire h_u_arrmul32_and14_16_y0;
  wire h_u_arrmul32_fa14_16_y2;
  wire h_u_arrmul32_fa14_16_y4;
  wire h_u_arrmul32_and15_16_y0;
  wire h_u_arrmul32_fa15_16_y2;
  wire h_u_arrmul32_fa15_16_y4;
  wire h_u_arrmul32_and16_16_y0;
  wire h_u_arrmul32_fa16_16_y2;
  wire h_u_arrmul32_fa16_16_y4;
  wire h_u_arrmul32_and17_16_y0;
  wire h_u_arrmul32_fa17_16_y2;
  wire h_u_arrmul32_fa17_16_y4;
  wire h_u_arrmul32_and18_16_y0;
  wire h_u_arrmul32_fa18_16_y2;
  wire h_u_arrmul32_fa18_16_y4;
  wire h_u_arrmul32_and19_16_y0;
  wire h_u_arrmul32_fa19_16_y2;
  wire h_u_arrmul32_fa19_16_y4;
  wire h_u_arrmul32_and20_16_y0;
  wire h_u_arrmul32_fa20_16_y2;
  wire h_u_arrmul32_fa20_16_y4;
  wire h_u_arrmul32_and21_16_y0;
  wire h_u_arrmul32_fa21_16_y2;
  wire h_u_arrmul32_fa21_16_y4;
  wire h_u_arrmul32_and22_16_y0;
  wire h_u_arrmul32_fa22_16_y2;
  wire h_u_arrmul32_fa22_16_y4;
  wire h_u_arrmul32_and23_16_y0;
  wire h_u_arrmul32_fa23_16_y2;
  wire h_u_arrmul32_fa23_16_y4;
  wire h_u_arrmul32_and24_16_y0;
  wire h_u_arrmul32_fa24_16_y2;
  wire h_u_arrmul32_fa24_16_y4;
  wire h_u_arrmul32_and25_16_y0;
  wire h_u_arrmul32_fa25_16_y2;
  wire h_u_arrmul32_fa25_16_y4;
  wire h_u_arrmul32_and26_16_y0;
  wire h_u_arrmul32_fa26_16_y2;
  wire h_u_arrmul32_fa26_16_y4;
  wire h_u_arrmul32_and27_16_y0;
  wire h_u_arrmul32_fa27_16_y2;
  wire h_u_arrmul32_fa27_16_y4;
  wire h_u_arrmul32_and28_16_y0;
  wire h_u_arrmul32_fa28_16_y2;
  wire h_u_arrmul32_fa28_16_y4;
  wire h_u_arrmul32_and29_16_y0;
  wire h_u_arrmul32_fa29_16_y2;
  wire h_u_arrmul32_fa29_16_y4;
  wire h_u_arrmul32_and30_16_y0;
  wire h_u_arrmul32_fa30_16_y2;
  wire h_u_arrmul32_fa30_16_y4;
  wire h_u_arrmul32_and31_16_y0;
  wire h_u_arrmul32_fa31_16_y2;
  wire h_u_arrmul32_fa31_16_y4;
  wire h_u_arrmul32_and0_17_y0;
  wire h_u_arrmul32_ha0_17_y0;
  wire h_u_arrmul32_ha0_17_y1;
  wire h_u_arrmul32_and1_17_y0;
  wire h_u_arrmul32_fa1_17_y2;
  wire h_u_arrmul32_fa1_17_y4;
  wire h_u_arrmul32_and2_17_y0;
  wire h_u_arrmul32_fa2_17_y2;
  wire h_u_arrmul32_fa2_17_y4;
  wire h_u_arrmul32_and3_17_y0;
  wire h_u_arrmul32_fa3_17_y2;
  wire h_u_arrmul32_fa3_17_y4;
  wire h_u_arrmul32_and4_17_y0;
  wire h_u_arrmul32_fa4_17_y2;
  wire h_u_arrmul32_fa4_17_y4;
  wire h_u_arrmul32_and5_17_y0;
  wire h_u_arrmul32_fa5_17_y2;
  wire h_u_arrmul32_fa5_17_y4;
  wire h_u_arrmul32_and6_17_y0;
  wire h_u_arrmul32_fa6_17_y2;
  wire h_u_arrmul32_fa6_17_y4;
  wire h_u_arrmul32_and7_17_y0;
  wire h_u_arrmul32_fa7_17_y2;
  wire h_u_arrmul32_fa7_17_y4;
  wire h_u_arrmul32_and8_17_y0;
  wire h_u_arrmul32_fa8_17_y2;
  wire h_u_arrmul32_fa8_17_y4;
  wire h_u_arrmul32_and9_17_y0;
  wire h_u_arrmul32_fa9_17_y2;
  wire h_u_arrmul32_fa9_17_y4;
  wire h_u_arrmul32_and10_17_y0;
  wire h_u_arrmul32_fa10_17_y2;
  wire h_u_arrmul32_fa10_17_y4;
  wire h_u_arrmul32_and11_17_y0;
  wire h_u_arrmul32_fa11_17_y2;
  wire h_u_arrmul32_fa11_17_y4;
  wire h_u_arrmul32_and12_17_y0;
  wire h_u_arrmul32_fa12_17_y2;
  wire h_u_arrmul32_fa12_17_y4;
  wire h_u_arrmul32_and13_17_y0;
  wire h_u_arrmul32_fa13_17_y2;
  wire h_u_arrmul32_fa13_17_y4;
  wire h_u_arrmul32_and14_17_y0;
  wire h_u_arrmul32_fa14_17_y2;
  wire h_u_arrmul32_fa14_17_y4;
  wire h_u_arrmul32_and15_17_y0;
  wire h_u_arrmul32_fa15_17_y2;
  wire h_u_arrmul32_fa15_17_y4;
  wire h_u_arrmul32_and16_17_y0;
  wire h_u_arrmul32_fa16_17_y2;
  wire h_u_arrmul32_fa16_17_y4;
  wire h_u_arrmul32_and17_17_y0;
  wire h_u_arrmul32_fa17_17_y2;
  wire h_u_arrmul32_fa17_17_y4;
  wire h_u_arrmul32_and18_17_y0;
  wire h_u_arrmul32_fa18_17_y2;
  wire h_u_arrmul32_fa18_17_y4;
  wire h_u_arrmul32_and19_17_y0;
  wire h_u_arrmul32_fa19_17_y2;
  wire h_u_arrmul32_fa19_17_y4;
  wire h_u_arrmul32_and20_17_y0;
  wire h_u_arrmul32_fa20_17_y2;
  wire h_u_arrmul32_fa20_17_y4;
  wire h_u_arrmul32_and21_17_y0;
  wire h_u_arrmul32_fa21_17_y2;
  wire h_u_arrmul32_fa21_17_y4;
  wire h_u_arrmul32_and22_17_y0;
  wire h_u_arrmul32_fa22_17_y2;
  wire h_u_arrmul32_fa22_17_y4;
  wire h_u_arrmul32_and23_17_y0;
  wire h_u_arrmul32_fa23_17_y2;
  wire h_u_arrmul32_fa23_17_y4;
  wire h_u_arrmul32_and24_17_y0;
  wire h_u_arrmul32_fa24_17_y2;
  wire h_u_arrmul32_fa24_17_y4;
  wire h_u_arrmul32_and25_17_y0;
  wire h_u_arrmul32_fa25_17_y2;
  wire h_u_arrmul32_fa25_17_y4;
  wire h_u_arrmul32_and26_17_y0;
  wire h_u_arrmul32_fa26_17_y2;
  wire h_u_arrmul32_fa26_17_y4;
  wire h_u_arrmul32_and27_17_y0;
  wire h_u_arrmul32_fa27_17_y2;
  wire h_u_arrmul32_fa27_17_y4;
  wire h_u_arrmul32_and28_17_y0;
  wire h_u_arrmul32_fa28_17_y2;
  wire h_u_arrmul32_fa28_17_y4;
  wire h_u_arrmul32_and29_17_y0;
  wire h_u_arrmul32_fa29_17_y2;
  wire h_u_arrmul32_fa29_17_y4;
  wire h_u_arrmul32_and30_17_y0;
  wire h_u_arrmul32_fa30_17_y2;
  wire h_u_arrmul32_fa30_17_y4;
  wire h_u_arrmul32_and31_17_y0;
  wire h_u_arrmul32_fa31_17_y2;
  wire h_u_arrmul32_fa31_17_y4;
  wire h_u_arrmul32_and0_18_y0;
  wire h_u_arrmul32_ha0_18_y0;
  wire h_u_arrmul32_ha0_18_y1;
  wire h_u_arrmul32_and1_18_y0;
  wire h_u_arrmul32_fa1_18_y2;
  wire h_u_arrmul32_fa1_18_y4;
  wire h_u_arrmul32_and2_18_y0;
  wire h_u_arrmul32_fa2_18_y2;
  wire h_u_arrmul32_fa2_18_y4;
  wire h_u_arrmul32_and3_18_y0;
  wire h_u_arrmul32_fa3_18_y2;
  wire h_u_arrmul32_fa3_18_y4;
  wire h_u_arrmul32_and4_18_y0;
  wire h_u_arrmul32_fa4_18_y2;
  wire h_u_arrmul32_fa4_18_y4;
  wire h_u_arrmul32_and5_18_y0;
  wire h_u_arrmul32_fa5_18_y2;
  wire h_u_arrmul32_fa5_18_y4;
  wire h_u_arrmul32_and6_18_y0;
  wire h_u_arrmul32_fa6_18_y2;
  wire h_u_arrmul32_fa6_18_y4;
  wire h_u_arrmul32_and7_18_y0;
  wire h_u_arrmul32_fa7_18_y2;
  wire h_u_arrmul32_fa7_18_y4;
  wire h_u_arrmul32_and8_18_y0;
  wire h_u_arrmul32_fa8_18_y2;
  wire h_u_arrmul32_fa8_18_y4;
  wire h_u_arrmul32_and9_18_y0;
  wire h_u_arrmul32_fa9_18_y2;
  wire h_u_arrmul32_fa9_18_y4;
  wire h_u_arrmul32_and10_18_y0;
  wire h_u_arrmul32_fa10_18_y2;
  wire h_u_arrmul32_fa10_18_y4;
  wire h_u_arrmul32_and11_18_y0;
  wire h_u_arrmul32_fa11_18_y2;
  wire h_u_arrmul32_fa11_18_y4;
  wire h_u_arrmul32_and12_18_y0;
  wire h_u_arrmul32_fa12_18_y2;
  wire h_u_arrmul32_fa12_18_y4;
  wire h_u_arrmul32_and13_18_y0;
  wire h_u_arrmul32_fa13_18_y2;
  wire h_u_arrmul32_fa13_18_y4;
  wire h_u_arrmul32_and14_18_y0;
  wire h_u_arrmul32_fa14_18_y2;
  wire h_u_arrmul32_fa14_18_y4;
  wire h_u_arrmul32_and15_18_y0;
  wire h_u_arrmul32_fa15_18_y2;
  wire h_u_arrmul32_fa15_18_y4;
  wire h_u_arrmul32_and16_18_y0;
  wire h_u_arrmul32_fa16_18_y2;
  wire h_u_arrmul32_fa16_18_y4;
  wire h_u_arrmul32_and17_18_y0;
  wire h_u_arrmul32_fa17_18_y2;
  wire h_u_arrmul32_fa17_18_y4;
  wire h_u_arrmul32_and18_18_y0;
  wire h_u_arrmul32_fa18_18_y2;
  wire h_u_arrmul32_fa18_18_y4;
  wire h_u_arrmul32_and19_18_y0;
  wire h_u_arrmul32_fa19_18_y2;
  wire h_u_arrmul32_fa19_18_y4;
  wire h_u_arrmul32_and20_18_y0;
  wire h_u_arrmul32_fa20_18_y2;
  wire h_u_arrmul32_fa20_18_y4;
  wire h_u_arrmul32_and21_18_y0;
  wire h_u_arrmul32_fa21_18_y2;
  wire h_u_arrmul32_fa21_18_y4;
  wire h_u_arrmul32_and22_18_y0;
  wire h_u_arrmul32_fa22_18_y2;
  wire h_u_arrmul32_fa22_18_y4;
  wire h_u_arrmul32_and23_18_y0;
  wire h_u_arrmul32_fa23_18_y2;
  wire h_u_arrmul32_fa23_18_y4;
  wire h_u_arrmul32_and24_18_y0;
  wire h_u_arrmul32_fa24_18_y2;
  wire h_u_arrmul32_fa24_18_y4;
  wire h_u_arrmul32_and25_18_y0;
  wire h_u_arrmul32_fa25_18_y2;
  wire h_u_arrmul32_fa25_18_y4;
  wire h_u_arrmul32_and26_18_y0;
  wire h_u_arrmul32_fa26_18_y2;
  wire h_u_arrmul32_fa26_18_y4;
  wire h_u_arrmul32_and27_18_y0;
  wire h_u_arrmul32_fa27_18_y2;
  wire h_u_arrmul32_fa27_18_y4;
  wire h_u_arrmul32_and28_18_y0;
  wire h_u_arrmul32_fa28_18_y2;
  wire h_u_arrmul32_fa28_18_y4;
  wire h_u_arrmul32_and29_18_y0;
  wire h_u_arrmul32_fa29_18_y2;
  wire h_u_arrmul32_fa29_18_y4;
  wire h_u_arrmul32_and30_18_y0;
  wire h_u_arrmul32_fa30_18_y2;
  wire h_u_arrmul32_fa30_18_y4;
  wire h_u_arrmul32_and31_18_y0;
  wire h_u_arrmul32_fa31_18_y2;
  wire h_u_arrmul32_fa31_18_y4;
  wire h_u_arrmul32_and0_19_y0;
  wire h_u_arrmul32_ha0_19_y0;
  wire h_u_arrmul32_ha0_19_y1;
  wire h_u_arrmul32_and1_19_y0;
  wire h_u_arrmul32_fa1_19_y2;
  wire h_u_arrmul32_fa1_19_y4;
  wire h_u_arrmul32_and2_19_y0;
  wire h_u_arrmul32_fa2_19_y2;
  wire h_u_arrmul32_fa2_19_y4;
  wire h_u_arrmul32_and3_19_y0;
  wire h_u_arrmul32_fa3_19_y2;
  wire h_u_arrmul32_fa3_19_y4;
  wire h_u_arrmul32_and4_19_y0;
  wire h_u_arrmul32_fa4_19_y2;
  wire h_u_arrmul32_fa4_19_y4;
  wire h_u_arrmul32_and5_19_y0;
  wire h_u_arrmul32_fa5_19_y2;
  wire h_u_arrmul32_fa5_19_y4;
  wire h_u_arrmul32_and6_19_y0;
  wire h_u_arrmul32_fa6_19_y2;
  wire h_u_arrmul32_fa6_19_y4;
  wire h_u_arrmul32_and7_19_y0;
  wire h_u_arrmul32_fa7_19_y2;
  wire h_u_arrmul32_fa7_19_y4;
  wire h_u_arrmul32_and8_19_y0;
  wire h_u_arrmul32_fa8_19_y2;
  wire h_u_arrmul32_fa8_19_y4;
  wire h_u_arrmul32_and9_19_y0;
  wire h_u_arrmul32_fa9_19_y2;
  wire h_u_arrmul32_fa9_19_y4;
  wire h_u_arrmul32_and10_19_y0;
  wire h_u_arrmul32_fa10_19_y2;
  wire h_u_arrmul32_fa10_19_y4;
  wire h_u_arrmul32_and11_19_y0;
  wire h_u_arrmul32_fa11_19_y2;
  wire h_u_arrmul32_fa11_19_y4;
  wire h_u_arrmul32_and12_19_y0;
  wire h_u_arrmul32_fa12_19_y2;
  wire h_u_arrmul32_fa12_19_y4;
  wire h_u_arrmul32_and13_19_y0;
  wire h_u_arrmul32_fa13_19_y2;
  wire h_u_arrmul32_fa13_19_y4;
  wire h_u_arrmul32_and14_19_y0;
  wire h_u_arrmul32_fa14_19_y2;
  wire h_u_arrmul32_fa14_19_y4;
  wire h_u_arrmul32_and15_19_y0;
  wire h_u_arrmul32_fa15_19_y2;
  wire h_u_arrmul32_fa15_19_y4;
  wire h_u_arrmul32_and16_19_y0;
  wire h_u_arrmul32_fa16_19_y2;
  wire h_u_arrmul32_fa16_19_y4;
  wire h_u_arrmul32_and17_19_y0;
  wire h_u_arrmul32_fa17_19_y2;
  wire h_u_arrmul32_fa17_19_y4;
  wire h_u_arrmul32_and18_19_y0;
  wire h_u_arrmul32_fa18_19_y2;
  wire h_u_arrmul32_fa18_19_y4;
  wire h_u_arrmul32_and19_19_y0;
  wire h_u_arrmul32_fa19_19_y2;
  wire h_u_arrmul32_fa19_19_y4;
  wire h_u_arrmul32_and20_19_y0;
  wire h_u_arrmul32_fa20_19_y2;
  wire h_u_arrmul32_fa20_19_y4;
  wire h_u_arrmul32_and21_19_y0;
  wire h_u_arrmul32_fa21_19_y2;
  wire h_u_arrmul32_fa21_19_y4;
  wire h_u_arrmul32_and22_19_y0;
  wire h_u_arrmul32_fa22_19_y2;
  wire h_u_arrmul32_fa22_19_y4;
  wire h_u_arrmul32_and23_19_y0;
  wire h_u_arrmul32_fa23_19_y2;
  wire h_u_arrmul32_fa23_19_y4;
  wire h_u_arrmul32_and24_19_y0;
  wire h_u_arrmul32_fa24_19_y2;
  wire h_u_arrmul32_fa24_19_y4;
  wire h_u_arrmul32_and25_19_y0;
  wire h_u_arrmul32_fa25_19_y2;
  wire h_u_arrmul32_fa25_19_y4;
  wire h_u_arrmul32_and26_19_y0;
  wire h_u_arrmul32_fa26_19_y2;
  wire h_u_arrmul32_fa26_19_y4;
  wire h_u_arrmul32_and27_19_y0;
  wire h_u_arrmul32_fa27_19_y2;
  wire h_u_arrmul32_fa27_19_y4;
  wire h_u_arrmul32_and28_19_y0;
  wire h_u_arrmul32_fa28_19_y2;
  wire h_u_arrmul32_fa28_19_y4;
  wire h_u_arrmul32_and29_19_y0;
  wire h_u_arrmul32_fa29_19_y2;
  wire h_u_arrmul32_fa29_19_y4;
  wire h_u_arrmul32_and30_19_y0;
  wire h_u_arrmul32_fa30_19_y2;
  wire h_u_arrmul32_fa30_19_y4;
  wire h_u_arrmul32_and31_19_y0;
  wire h_u_arrmul32_fa31_19_y2;
  wire h_u_arrmul32_fa31_19_y4;
  wire h_u_arrmul32_and0_20_y0;
  wire h_u_arrmul32_ha0_20_y0;
  wire h_u_arrmul32_ha0_20_y1;
  wire h_u_arrmul32_and1_20_y0;
  wire h_u_arrmul32_fa1_20_y2;
  wire h_u_arrmul32_fa1_20_y4;
  wire h_u_arrmul32_and2_20_y0;
  wire h_u_arrmul32_fa2_20_y2;
  wire h_u_arrmul32_fa2_20_y4;
  wire h_u_arrmul32_and3_20_y0;
  wire h_u_arrmul32_fa3_20_y2;
  wire h_u_arrmul32_fa3_20_y4;
  wire h_u_arrmul32_and4_20_y0;
  wire h_u_arrmul32_fa4_20_y2;
  wire h_u_arrmul32_fa4_20_y4;
  wire h_u_arrmul32_and5_20_y0;
  wire h_u_arrmul32_fa5_20_y2;
  wire h_u_arrmul32_fa5_20_y4;
  wire h_u_arrmul32_and6_20_y0;
  wire h_u_arrmul32_fa6_20_y2;
  wire h_u_arrmul32_fa6_20_y4;
  wire h_u_arrmul32_and7_20_y0;
  wire h_u_arrmul32_fa7_20_y2;
  wire h_u_arrmul32_fa7_20_y4;
  wire h_u_arrmul32_and8_20_y0;
  wire h_u_arrmul32_fa8_20_y2;
  wire h_u_arrmul32_fa8_20_y4;
  wire h_u_arrmul32_and9_20_y0;
  wire h_u_arrmul32_fa9_20_y2;
  wire h_u_arrmul32_fa9_20_y4;
  wire h_u_arrmul32_and10_20_y0;
  wire h_u_arrmul32_fa10_20_y2;
  wire h_u_arrmul32_fa10_20_y4;
  wire h_u_arrmul32_and11_20_y0;
  wire h_u_arrmul32_fa11_20_y2;
  wire h_u_arrmul32_fa11_20_y4;
  wire h_u_arrmul32_and12_20_y0;
  wire h_u_arrmul32_fa12_20_y2;
  wire h_u_arrmul32_fa12_20_y4;
  wire h_u_arrmul32_and13_20_y0;
  wire h_u_arrmul32_fa13_20_y2;
  wire h_u_arrmul32_fa13_20_y4;
  wire h_u_arrmul32_and14_20_y0;
  wire h_u_arrmul32_fa14_20_y2;
  wire h_u_arrmul32_fa14_20_y4;
  wire h_u_arrmul32_and15_20_y0;
  wire h_u_arrmul32_fa15_20_y2;
  wire h_u_arrmul32_fa15_20_y4;
  wire h_u_arrmul32_and16_20_y0;
  wire h_u_arrmul32_fa16_20_y2;
  wire h_u_arrmul32_fa16_20_y4;
  wire h_u_arrmul32_and17_20_y0;
  wire h_u_arrmul32_fa17_20_y2;
  wire h_u_arrmul32_fa17_20_y4;
  wire h_u_arrmul32_and18_20_y0;
  wire h_u_arrmul32_fa18_20_y2;
  wire h_u_arrmul32_fa18_20_y4;
  wire h_u_arrmul32_and19_20_y0;
  wire h_u_arrmul32_fa19_20_y2;
  wire h_u_arrmul32_fa19_20_y4;
  wire h_u_arrmul32_and20_20_y0;
  wire h_u_arrmul32_fa20_20_y2;
  wire h_u_arrmul32_fa20_20_y4;
  wire h_u_arrmul32_and21_20_y0;
  wire h_u_arrmul32_fa21_20_y2;
  wire h_u_arrmul32_fa21_20_y4;
  wire h_u_arrmul32_and22_20_y0;
  wire h_u_arrmul32_fa22_20_y2;
  wire h_u_arrmul32_fa22_20_y4;
  wire h_u_arrmul32_and23_20_y0;
  wire h_u_arrmul32_fa23_20_y2;
  wire h_u_arrmul32_fa23_20_y4;
  wire h_u_arrmul32_and24_20_y0;
  wire h_u_arrmul32_fa24_20_y2;
  wire h_u_arrmul32_fa24_20_y4;
  wire h_u_arrmul32_and25_20_y0;
  wire h_u_arrmul32_fa25_20_y2;
  wire h_u_arrmul32_fa25_20_y4;
  wire h_u_arrmul32_and26_20_y0;
  wire h_u_arrmul32_fa26_20_y2;
  wire h_u_arrmul32_fa26_20_y4;
  wire h_u_arrmul32_and27_20_y0;
  wire h_u_arrmul32_fa27_20_y2;
  wire h_u_arrmul32_fa27_20_y4;
  wire h_u_arrmul32_and28_20_y0;
  wire h_u_arrmul32_fa28_20_y2;
  wire h_u_arrmul32_fa28_20_y4;
  wire h_u_arrmul32_and29_20_y0;
  wire h_u_arrmul32_fa29_20_y2;
  wire h_u_arrmul32_fa29_20_y4;
  wire h_u_arrmul32_and30_20_y0;
  wire h_u_arrmul32_fa30_20_y2;
  wire h_u_arrmul32_fa30_20_y4;
  wire h_u_arrmul32_and31_20_y0;
  wire h_u_arrmul32_fa31_20_y2;
  wire h_u_arrmul32_fa31_20_y4;
  wire h_u_arrmul32_and0_21_y0;
  wire h_u_arrmul32_ha0_21_y0;
  wire h_u_arrmul32_ha0_21_y1;
  wire h_u_arrmul32_and1_21_y0;
  wire h_u_arrmul32_fa1_21_y2;
  wire h_u_arrmul32_fa1_21_y4;
  wire h_u_arrmul32_and2_21_y0;
  wire h_u_arrmul32_fa2_21_y2;
  wire h_u_arrmul32_fa2_21_y4;
  wire h_u_arrmul32_and3_21_y0;
  wire h_u_arrmul32_fa3_21_y2;
  wire h_u_arrmul32_fa3_21_y4;
  wire h_u_arrmul32_and4_21_y0;
  wire h_u_arrmul32_fa4_21_y2;
  wire h_u_arrmul32_fa4_21_y4;
  wire h_u_arrmul32_and5_21_y0;
  wire h_u_arrmul32_fa5_21_y2;
  wire h_u_arrmul32_fa5_21_y4;
  wire h_u_arrmul32_and6_21_y0;
  wire h_u_arrmul32_fa6_21_y2;
  wire h_u_arrmul32_fa6_21_y4;
  wire h_u_arrmul32_and7_21_y0;
  wire h_u_arrmul32_fa7_21_y2;
  wire h_u_arrmul32_fa7_21_y4;
  wire h_u_arrmul32_and8_21_y0;
  wire h_u_arrmul32_fa8_21_y2;
  wire h_u_arrmul32_fa8_21_y4;
  wire h_u_arrmul32_and9_21_y0;
  wire h_u_arrmul32_fa9_21_y2;
  wire h_u_arrmul32_fa9_21_y4;
  wire h_u_arrmul32_and10_21_y0;
  wire h_u_arrmul32_fa10_21_y2;
  wire h_u_arrmul32_fa10_21_y4;
  wire h_u_arrmul32_and11_21_y0;
  wire h_u_arrmul32_fa11_21_y2;
  wire h_u_arrmul32_fa11_21_y4;
  wire h_u_arrmul32_and12_21_y0;
  wire h_u_arrmul32_fa12_21_y2;
  wire h_u_arrmul32_fa12_21_y4;
  wire h_u_arrmul32_and13_21_y0;
  wire h_u_arrmul32_fa13_21_y2;
  wire h_u_arrmul32_fa13_21_y4;
  wire h_u_arrmul32_and14_21_y0;
  wire h_u_arrmul32_fa14_21_y2;
  wire h_u_arrmul32_fa14_21_y4;
  wire h_u_arrmul32_and15_21_y0;
  wire h_u_arrmul32_fa15_21_y2;
  wire h_u_arrmul32_fa15_21_y4;
  wire h_u_arrmul32_and16_21_y0;
  wire h_u_arrmul32_fa16_21_y2;
  wire h_u_arrmul32_fa16_21_y4;
  wire h_u_arrmul32_and17_21_y0;
  wire h_u_arrmul32_fa17_21_y2;
  wire h_u_arrmul32_fa17_21_y4;
  wire h_u_arrmul32_and18_21_y0;
  wire h_u_arrmul32_fa18_21_y2;
  wire h_u_arrmul32_fa18_21_y4;
  wire h_u_arrmul32_and19_21_y0;
  wire h_u_arrmul32_fa19_21_y2;
  wire h_u_arrmul32_fa19_21_y4;
  wire h_u_arrmul32_and20_21_y0;
  wire h_u_arrmul32_fa20_21_y2;
  wire h_u_arrmul32_fa20_21_y4;
  wire h_u_arrmul32_and21_21_y0;
  wire h_u_arrmul32_fa21_21_y2;
  wire h_u_arrmul32_fa21_21_y4;
  wire h_u_arrmul32_and22_21_y0;
  wire h_u_arrmul32_fa22_21_y2;
  wire h_u_arrmul32_fa22_21_y4;
  wire h_u_arrmul32_and23_21_y0;
  wire h_u_arrmul32_fa23_21_y2;
  wire h_u_arrmul32_fa23_21_y4;
  wire h_u_arrmul32_and24_21_y0;
  wire h_u_arrmul32_fa24_21_y2;
  wire h_u_arrmul32_fa24_21_y4;
  wire h_u_arrmul32_and25_21_y0;
  wire h_u_arrmul32_fa25_21_y2;
  wire h_u_arrmul32_fa25_21_y4;
  wire h_u_arrmul32_and26_21_y0;
  wire h_u_arrmul32_fa26_21_y2;
  wire h_u_arrmul32_fa26_21_y4;
  wire h_u_arrmul32_and27_21_y0;
  wire h_u_arrmul32_fa27_21_y2;
  wire h_u_arrmul32_fa27_21_y4;
  wire h_u_arrmul32_and28_21_y0;
  wire h_u_arrmul32_fa28_21_y2;
  wire h_u_arrmul32_fa28_21_y4;
  wire h_u_arrmul32_and29_21_y0;
  wire h_u_arrmul32_fa29_21_y2;
  wire h_u_arrmul32_fa29_21_y4;
  wire h_u_arrmul32_and30_21_y0;
  wire h_u_arrmul32_fa30_21_y2;
  wire h_u_arrmul32_fa30_21_y4;
  wire h_u_arrmul32_and31_21_y0;
  wire h_u_arrmul32_fa31_21_y2;
  wire h_u_arrmul32_fa31_21_y4;
  wire h_u_arrmul32_and0_22_y0;
  wire h_u_arrmul32_ha0_22_y0;
  wire h_u_arrmul32_ha0_22_y1;
  wire h_u_arrmul32_and1_22_y0;
  wire h_u_arrmul32_fa1_22_y2;
  wire h_u_arrmul32_fa1_22_y4;
  wire h_u_arrmul32_and2_22_y0;
  wire h_u_arrmul32_fa2_22_y2;
  wire h_u_arrmul32_fa2_22_y4;
  wire h_u_arrmul32_and3_22_y0;
  wire h_u_arrmul32_fa3_22_y2;
  wire h_u_arrmul32_fa3_22_y4;
  wire h_u_arrmul32_and4_22_y0;
  wire h_u_arrmul32_fa4_22_y2;
  wire h_u_arrmul32_fa4_22_y4;
  wire h_u_arrmul32_and5_22_y0;
  wire h_u_arrmul32_fa5_22_y2;
  wire h_u_arrmul32_fa5_22_y4;
  wire h_u_arrmul32_and6_22_y0;
  wire h_u_arrmul32_fa6_22_y2;
  wire h_u_arrmul32_fa6_22_y4;
  wire h_u_arrmul32_and7_22_y0;
  wire h_u_arrmul32_fa7_22_y2;
  wire h_u_arrmul32_fa7_22_y4;
  wire h_u_arrmul32_and8_22_y0;
  wire h_u_arrmul32_fa8_22_y2;
  wire h_u_arrmul32_fa8_22_y4;
  wire h_u_arrmul32_and9_22_y0;
  wire h_u_arrmul32_fa9_22_y2;
  wire h_u_arrmul32_fa9_22_y4;
  wire h_u_arrmul32_and10_22_y0;
  wire h_u_arrmul32_fa10_22_y2;
  wire h_u_arrmul32_fa10_22_y4;
  wire h_u_arrmul32_and11_22_y0;
  wire h_u_arrmul32_fa11_22_y2;
  wire h_u_arrmul32_fa11_22_y4;
  wire h_u_arrmul32_and12_22_y0;
  wire h_u_arrmul32_fa12_22_y2;
  wire h_u_arrmul32_fa12_22_y4;
  wire h_u_arrmul32_and13_22_y0;
  wire h_u_arrmul32_fa13_22_y2;
  wire h_u_arrmul32_fa13_22_y4;
  wire h_u_arrmul32_and14_22_y0;
  wire h_u_arrmul32_fa14_22_y2;
  wire h_u_arrmul32_fa14_22_y4;
  wire h_u_arrmul32_and15_22_y0;
  wire h_u_arrmul32_fa15_22_y2;
  wire h_u_arrmul32_fa15_22_y4;
  wire h_u_arrmul32_and16_22_y0;
  wire h_u_arrmul32_fa16_22_y2;
  wire h_u_arrmul32_fa16_22_y4;
  wire h_u_arrmul32_and17_22_y0;
  wire h_u_arrmul32_fa17_22_y2;
  wire h_u_arrmul32_fa17_22_y4;
  wire h_u_arrmul32_and18_22_y0;
  wire h_u_arrmul32_fa18_22_y2;
  wire h_u_arrmul32_fa18_22_y4;
  wire h_u_arrmul32_and19_22_y0;
  wire h_u_arrmul32_fa19_22_y2;
  wire h_u_arrmul32_fa19_22_y4;
  wire h_u_arrmul32_and20_22_y0;
  wire h_u_arrmul32_fa20_22_y2;
  wire h_u_arrmul32_fa20_22_y4;
  wire h_u_arrmul32_and21_22_y0;
  wire h_u_arrmul32_fa21_22_y2;
  wire h_u_arrmul32_fa21_22_y4;
  wire h_u_arrmul32_and22_22_y0;
  wire h_u_arrmul32_fa22_22_y2;
  wire h_u_arrmul32_fa22_22_y4;
  wire h_u_arrmul32_and23_22_y0;
  wire h_u_arrmul32_fa23_22_y2;
  wire h_u_arrmul32_fa23_22_y4;
  wire h_u_arrmul32_and24_22_y0;
  wire h_u_arrmul32_fa24_22_y2;
  wire h_u_arrmul32_fa24_22_y4;
  wire h_u_arrmul32_and25_22_y0;
  wire h_u_arrmul32_fa25_22_y2;
  wire h_u_arrmul32_fa25_22_y4;
  wire h_u_arrmul32_and26_22_y0;
  wire h_u_arrmul32_fa26_22_y2;
  wire h_u_arrmul32_fa26_22_y4;
  wire h_u_arrmul32_and27_22_y0;
  wire h_u_arrmul32_fa27_22_y2;
  wire h_u_arrmul32_fa27_22_y4;
  wire h_u_arrmul32_and28_22_y0;
  wire h_u_arrmul32_fa28_22_y2;
  wire h_u_arrmul32_fa28_22_y4;
  wire h_u_arrmul32_and29_22_y0;
  wire h_u_arrmul32_fa29_22_y2;
  wire h_u_arrmul32_fa29_22_y4;
  wire h_u_arrmul32_and30_22_y0;
  wire h_u_arrmul32_fa30_22_y2;
  wire h_u_arrmul32_fa30_22_y4;
  wire h_u_arrmul32_and31_22_y0;
  wire h_u_arrmul32_fa31_22_y2;
  wire h_u_arrmul32_fa31_22_y4;
  wire h_u_arrmul32_and0_23_y0;
  wire h_u_arrmul32_ha0_23_y0;
  wire h_u_arrmul32_ha0_23_y1;
  wire h_u_arrmul32_and1_23_y0;
  wire h_u_arrmul32_fa1_23_y2;
  wire h_u_arrmul32_fa1_23_y4;
  wire h_u_arrmul32_and2_23_y0;
  wire h_u_arrmul32_fa2_23_y2;
  wire h_u_arrmul32_fa2_23_y4;
  wire h_u_arrmul32_and3_23_y0;
  wire h_u_arrmul32_fa3_23_y2;
  wire h_u_arrmul32_fa3_23_y4;
  wire h_u_arrmul32_and4_23_y0;
  wire h_u_arrmul32_fa4_23_y2;
  wire h_u_arrmul32_fa4_23_y4;
  wire h_u_arrmul32_and5_23_y0;
  wire h_u_arrmul32_fa5_23_y2;
  wire h_u_arrmul32_fa5_23_y4;
  wire h_u_arrmul32_and6_23_y0;
  wire h_u_arrmul32_fa6_23_y2;
  wire h_u_arrmul32_fa6_23_y4;
  wire h_u_arrmul32_and7_23_y0;
  wire h_u_arrmul32_fa7_23_y2;
  wire h_u_arrmul32_fa7_23_y4;
  wire h_u_arrmul32_and8_23_y0;
  wire h_u_arrmul32_fa8_23_y2;
  wire h_u_arrmul32_fa8_23_y4;
  wire h_u_arrmul32_and9_23_y0;
  wire h_u_arrmul32_fa9_23_y2;
  wire h_u_arrmul32_fa9_23_y4;
  wire h_u_arrmul32_and10_23_y0;
  wire h_u_arrmul32_fa10_23_y2;
  wire h_u_arrmul32_fa10_23_y4;
  wire h_u_arrmul32_and11_23_y0;
  wire h_u_arrmul32_fa11_23_y2;
  wire h_u_arrmul32_fa11_23_y4;
  wire h_u_arrmul32_and12_23_y0;
  wire h_u_arrmul32_fa12_23_y2;
  wire h_u_arrmul32_fa12_23_y4;
  wire h_u_arrmul32_and13_23_y0;
  wire h_u_arrmul32_fa13_23_y2;
  wire h_u_arrmul32_fa13_23_y4;
  wire h_u_arrmul32_and14_23_y0;
  wire h_u_arrmul32_fa14_23_y2;
  wire h_u_arrmul32_fa14_23_y4;
  wire h_u_arrmul32_and15_23_y0;
  wire h_u_arrmul32_fa15_23_y2;
  wire h_u_arrmul32_fa15_23_y4;
  wire h_u_arrmul32_and16_23_y0;
  wire h_u_arrmul32_fa16_23_y2;
  wire h_u_arrmul32_fa16_23_y4;
  wire h_u_arrmul32_and17_23_y0;
  wire h_u_arrmul32_fa17_23_y2;
  wire h_u_arrmul32_fa17_23_y4;
  wire h_u_arrmul32_and18_23_y0;
  wire h_u_arrmul32_fa18_23_y2;
  wire h_u_arrmul32_fa18_23_y4;
  wire h_u_arrmul32_and19_23_y0;
  wire h_u_arrmul32_fa19_23_y2;
  wire h_u_arrmul32_fa19_23_y4;
  wire h_u_arrmul32_and20_23_y0;
  wire h_u_arrmul32_fa20_23_y2;
  wire h_u_arrmul32_fa20_23_y4;
  wire h_u_arrmul32_and21_23_y0;
  wire h_u_arrmul32_fa21_23_y2;
  wire h_u_arrmul32_fa21_23_y4;
  wire h_u_arrmul32_and22_23_y0;
  wire h_u_arrmul32_fa22_23_y2;
  wire h_u_arrmul32_fa22_23_y4;
  wire h_u_arrmul32_and23_23_y0;
  wire h_u_arrmul32_fa23_23_y2;
  wire h_u_arrmul32_fa23_23_y4;
  wire h_u_arrmul32_and24_23_y0;
  wire h_u_arrmul32_fa24_23_y2;
  wire h_u_arrmul32_fa24_23_y4;
  wire h_u_arrmul32_and25_23_y0;
  wire h_u_arrmul32_fa25_23_y2;
  wire h_u_arrmul32_fa25_23_y4;
  wire h_u_arrmul32_and26_23_y0;
  wire h_u_arrmul32_fa26_23_y2;
  wire h_u_arrmul32_fa26_23_y4;
  wire h_u_arrmul32_and27_23_y0;
  wire h_u_arrmul32_fa27_23_y2;
  wire h_u_arrmul32_fa27_23_y4;
  wire h_u_arrmul32_and28_23_y0;
  wire h_u_arrmul32_fa28_23_y2;
  wire h_u_arrmul32_fa28_23_y4;
  wire h_u_arrmul32_and29_23_y0;
  wire h_u_arrmul32_fa29_23_y2;
  wire h_u_arrmul32_fa29_23_y4;
  wire h_u_arrmul32_and30_23_y0;
  wire h_u_arrmul32_fa30_23_y2;
  wire h_u_arrmul32_fa30_23_y4;
  wire h_u_arrmul32_and31_23_y0;
  wire h_u_arrmul32_fa31_23_y2;
  wire h_u_arrmul32_fa31_23_y4;
  wire h_u_arrmul32_and0_24_y0;
  wire h_u_arrmul32_ha0_24_y0;
  wire h_u_arrmul32_ha0_24_y1;
  wire h_u_arrmul32_and1_24_y0;
  wire h_u_arrmul32_fa1_24_y2;
  wire h_u_arrmul32_fa1_24_y4;
  wire h_u_arrmul32_and2_24_y0;
  wire h_u_arrmul32_fa2_24_y2;
  wire h_u_arrmul32_fa2_24_y4;
  wire h_u_arrmul32_and3_24_y0;
  wire h_u_arrmul32_fa3_24_y2;
  wire h_u_arrmul32_fa3_24_y4;
  wire h_u_arrmul32_and4_24_y0;
  wire h_u_arrmul32_fa4_24_y2;
  wire h_u_arrmul32_fa4_24_y4;
  wire h_u_arrmul32_and5_24_y0;
  wire h_u_arrmul32_fa5_24_y2;
  wire h_u_arrmul32_fa5_24_y4;
  wire h_u_arrmul32_and6_24_y0;
  wire h_u_arrmul32_fa6_24_y2;
  wire h_u_arrmul32_fa6_24_y4;
  wire h_u_arrmul32_and7_24_y0;
  wire h_u_arrmul32_fa7_24_y2;
  wire h_u_arrmul32_fa7_24_y4;
  wire h_u_arrmul32_and8_24_y0;
  wire h_u_arrmul32_fa8_24_y2;
  wire h_u_arrmul32_fa8_24_y4;
  wire h_u_arrmul32_and9_24_y0;
  wire h_u_arrmul32_fa9_24_y2;
  wire h_u_arrmul32_fa9_24_y4;
  wire h_u_arrmul32_and10_24_y0;
  wire h_u_arrmul32_fa10_24_y2;
  wire h_u_arrmul32_fa10_24_y4;
  wire h_u_arrmul32_and11_24_y0;
  wire h_u_arrmul32_fa11_24_y2;
  wire h_u_arrmul32_fa11_24_y4;
  wire h_u_arrmul32_and12_24_y0;
  wire h_u_arrmul32_fa12_24_y2;
  wire h_u_arrmul32_fa12_24_y4;
  wire h_u_arrmul32_and13_24_y0;
  wire h_u_arrmul32_fa13_24_y2;
  wire h_u_arrmul32_fa13_24_y4;
  wire h_u_arrmul32_and14_24_y0;
  wire h_u_arrmul32_fa14_24_y2;
  wire h_u_arrmul32_fa14_24_y4;
  wire h_u_arrmul32_and15_24_y0;
  wire h_u_arrmul32_fa15_24_y2;
  wire h_u_arrmul32_fa15_24_y4;
  wire h_u_arrmul32_and16_24_y0;
  wire h_u_arrmul32_fa16_24_y2;
  wire h_u_arrmul32_fa16_24_y4;
  wire h_u_arrmul32_and17_24_y0;
  wire h_u_arrmul32_fa17_24_y2;
  wire h_u_arrmul32_fa17_24_y4;
  wire h_u_arrmul32_and18_24_y0;
  wire h_u_arrmul32_fa18_24_y2;
  wire h_u_arrmul32_fa18_24_y4;
  wire h_u_arrmul32_and19_24_y0;
  wire h_u_arrmul32_fa19_24_y2;
  wire h_u_arrmul32_fa19_24_y4;
  wire h_u_arrmul32_and20_24_y0;
  wire h_u_arrmul32_fa20_24_y2;
  wire h_u_arrmul32_fa20_24_y4;
  wire h_u_arrmul32_and21_24_y0;
  wire h_u_arrmul32_fa21_24_y2;
  wire h_u_arrmul32_fa21_24_y4;
  wire h_u_arrmul32_and22_24_y0;
  wire h_u_arrmul32_fa22_24_y2;
  wire h_u_arrmul32_fa22_24_y4;
  wire h_u_arrmul32_and23_24_y0;
  wire h_u_arrmul32_fa23_24_y2;
  wire h_u_arrmul32_fa23_24_y4;
  wire h_u_arrmul32_and24_24_y0;
  wire h_u_arrmul32_fa24_24_y2;
  wire h_u_arrmul32_fa24_24_y4;
  wire h_u_arrmul32_and25_24_y0;
  wire h_u_arrmul32_fa25_24_y2;
  wire h_u_arrmul32_fa25_24_y4;
  wire h_u_arrmul32_and26_24_y0;
  wire h_u_arrmul32_fa26_24_y2;
  wire h_u_arrmul32_fa26_24_y4;
  wire h_u_arrmul32_and27_24_y0;
  wire h_u_arrmul32_fa27_24_y2;
  wire h_u_arrmul32_fa27_24_y4;
  wire h_u_arrmul32_and28_24_y0;
  wire h_u_arrmul32_fa28_24_y2;
  wire h_u_arrmul32_fa28_24_y4;
  wire h_u_arrmul32_and29_24_y0;
  wire h_u_arrmul32_fa29_24_y2;
  wire h_u_arrmul32_fa29_24_y4;
  wire h_u_arrmul32_and30_24_y0;
  wire h_u_arrmul32_fa30_24_y2;
  wire h_u_arrmul32_fa30_24_y4;
  wire h_u_arrmul32_and31_24_y0;
  wire h_u_arrmul32_fa31_24_y2;
  wire h_u_arrmul32_fa31_24_y4;
  wire h_u_arrmul32_and0_25_y0;
  wire h_u_arrmul32_ha0_25_y0;
  wire h_u_arrmul32_ha0_25_y1;
  wire h_u_arrmul32_and1_25_y0;
  wire h_u_arrmul32_fa1_25_y2;
  wire h_u_arrmul32_fa1_25_y4;
  wire h_u_arrmul32_and2_25_y0;
  wire h_u_arrmul32_fa2_25_y2;
  wire h_u_arrmul32_fa2_25_y4;
  wire h_u_arrmul32_and3_25_y0;
  wire h_u_arrmul32_fa3_25_y2;
  wire h_u_arrmul32_fa3_25_y4;
  wire h_u_arrmul32_and4_25_y0;
  wire h_u_arrmul32_fa4_25_y2;
  wire h_u_arrmul32_fa4_25_y4;
  wire h_u_arrmul32_and5_25_y0;
  wire h_u_arrmul32_fa5_25_y2;
  wire h_u_arrmul32_fa5_25_y4;
  wire h_u_arrmul32_and6_25_y0;
  wire h_u_arrmul32_fa6_25_y2;
  wire h_u_arrmul32_fa6_25_y4;
  wire h_u_arrmul32_and7_25_y0;
  wire h_u_arrmul32_fa7_25_y2;
  wire h_u_arrmul32_fa7_25_y4;
  wire h_u_arrmul32_and8_25_y0;
  wire h_u_arrmul32_fa8_25_y2;
  wire h_u_arrmul32_fa8_25_y4;
  wire h_u_arrmul32_and9_25_y0;
  wire h_u_arrmul32_fa9_25_y2;
  wire h_u_arrmul32_fa9_25_y4;
  wire h_u_arrmul32_and10_25_y0;
  wire h_u_arrmul32_fa10_25_y2;
  wire h_u_arrmul32_fa10_25_y4;
  wire h_u_arrmul32_and11_25_y0;
  wire h_u_arrmul32_fa11_25_y2;
  wire h_u_arrmul32_fa11_25_y4;
  wire h_u_arrmul32_and12_25_y0;
  wire h_u_arrmul32_fa12_25_y2;
  wire h_u_arrmul32_fa12_25_y4;
  wire h_u_arrmul32_and13_25_y0;
  wire h_u_arrmul32_fa13_25_y2;
  wire h_u_arrmul32_fa13_25_y4;
  wire h_u_arrmul32_and14_25_y0;
  wire h_u_arrmul32_fa14_25_y2;
  wire h_u_arrmul32_fa14_25_y4;
  wire h_u_arrmul32_and15_25_y0;
  wire h_u_arrmul32_fa15_25_y2;
  wire h_u_arrmul32_fa15_25_y4;
  wire h_u_arrmul32_and16_25_y0;
  wire h_u_arrmul32_fa16_25_y2;
  wire h_u_arrmul32_fa16_25_y4;
  wire h_u_arrmul32_and17_25_y0;
  wire h_u_arrmul32_fa17_25_y2;
  wire h_u_arrmul32_fa17_25_y4;
  wire h_u_arrmul32_and18_25_y0;
  wire h_u_arrmul32_fa18_25_y2;
  wire h_u_arrmul32_fa18_25_y4;
  wire h_u_arrmul32_and19_25_y0;
  wire h_u_arrmul32_fa19_25_y2;
  wire h_u_arrmul32_fa19_25_y4;
  wire h_u_arrmul32_and20_25_y0;
  wire h_u_arrmul32_fa20_25_y2;
  wire h_u_arrmul32_fa20_25_y4;
  wire h_u_arrmul32_and21_25_y0;
  wire h_u_arrmul32_fa21_25_y2;
  wire h_u_arrmul32_fa21_25_y4;
  wire h_u_arrmul32_and22_25_y0;
  wire h_u_arrmul32_fa22_25_y2;
  wire h_u_arrmul32_fa22_25_y4;
  wire h_u_arrmul32_and23_25_y0;
  wire h_u_arrmul32_fa23_25_y2;
  wire h_u_arrmul32_fa23_25_y4;
  wire h_u_arrmul32_and24_25_y0;
  wire h_u_arrmul32_fa24_25_y2;
  wire h_u_arrmul32_fa24_25_y4;
  wire h_u_arrmul32_and25_25_y0;
  wire h_u_arrmul32_fa25_25_y2;
  wire h_u_arrmul32_fa25_25_y4;
  wire h_u_arrmul32_and26_25_y0;
  wire h_u_arrmul32_fa26_25_y2;
  wire h_u_arrmul32_fa26_25_y4;
  wire h_u_arrmul32_and27_25_y0;
  wire h_u_arrmul32_fa27_25_y2;
  wire h_u_arrmul32_fa27_25_y4;
  wire h_u_arrmul32_and28_25_y0;
  wire h_u_arrmul32_fa28_25_y2;
  wire h_u_arrmul32_fa28_25_y4;
  wire h_u_arrmul32_and29_25_y0;
  wire h_u_arrmul32_fa29_25_y2;
  wire h_u_arrmul32_fa29_25_y4;
  wire h_u_arrmul32_and30_25_y0;
  wire h_u_arrmul32_fa30_25_y2;
  wire h_u_arrmul32_fa30_25_y4;
  wire h_u_arrmul32_and31_25_y0;
  wire h_u_arrmul32_fa31_25_y2;
  wire h_u_arrmul32_fa31_25_y4;
  wire h_u_arrmul32_and0_26_y0;
  wire h_u_arrmul32_ha0_26_y0;
  wire h_u_arrmul32_ha0_26_y1;
  wire h_u_arrmul32_and1_26_y0;
  wire h_u_arrmul32_fa1_26_y2;
  wire h_u_arrmul32_fa1_26_y4;
  wire h_u_arrmul32_and2_26_y0;
  wire h_u_arrmul32_fa2_26_y2;
  wire h_u_arrmul32_fa2_26_y4;
  wire h_u_arrmul32_and3_26_y0;
  wire h_u_arrmul32_fa3_26_y2;
  wire h_u_arrmul32_fa3_26_y4;
  wire h_u_arrmul32_and4_26_y0;
  wire h_u_arrmul32_fa4_26_y2;
  wire h_u_arrmul32_fa4_26_y4;
  wire h_u_arrmul32_and5_26_y0;
  wire h_u_arrmul32_fa5_26_y2;
  wire h_u_arrmul32_fa5_26_y4;
  wire h_u_arrmul32_and6_26_y0;
  wire h_u_arrmul32_fa6_26_y2;
  wire h_u_arrmul32_fa6_26_y4;
  wire h_u_arrmul32_and7_26_y0;
  wire h_u_arrmul32_fa7_26_y2;
  wire h_u_arrmul32_fa7_26_y4;
  wire h_u_arrmul32_and8_26_y0;
  wire h_u_arrmul32_fa8_26_y2;
  wire h_u_arrmul32_fa8_26_y4;
  wire h_u_arrmul32_and9_26_y0;
  wire h_u_arrmul32_fa9_26_y2;
  wire h_u_arrmul32_fa9_26_y4;
  wire h_u_arrmul32_and10_26_y0;
  wire h_u_arrmul32_fa10_26_y2;
  wire h_u_arrmul32_fa10_26_y4;
  wire h_u_arrmul32_and11_26_y0;
  wire h_u_arrmul32_fa11_26_y2;
  wire h_u_arrmul32_fa11_26_y4;
  wire h_u_arrmul32_and12_26_y0;
  wire h_u_arrmul32_fa12_26_y2;
  wire h_u_arrmul32_fa12_26_y4;
  wire h_u_arrmul32_and13_26_y0;
  wire h_u_arrmul32_fa13_26_y2;
  wire h_u_arrmul32_fa13_26_y4;
  wire h_u_arrmul32_and14_26_y0;
  wire h_u_arrmul32_fa14_26_y2;
  wire h_u_arrmul32_fa14_26_y4;
  wire h_u_arrmul32_and15_26_y0;
  wire h_u_arrmul32_fa15_26_y2;
  wire h_u_arrmul32_fa15_26_y4;
  wire h_u_arrmul32_and16_26_y0;
  wire h_u_arrmul32_fa16_26_y2;
  wire h_u_arrmul32_fa16_26_y4;
  wire h_u_arrmul32_and17_26_y0;
  wire h_u_arrmul32_fa17_26_y2;
  wire h_u_arrmul32_fa17_26_y4;
  wire h_u_arrmul32_and18_26_y0;
  wire h_u_arrmul32_fa18_26_y2;
  wire h_u_arrmul32_fa18_26_y4;
  wire h_u_arrmul32_and19_26_y0;
  wire h_u_arrmul32_fa19_26_y2;
  wire h_u_arrmul32_fa19_26_y4;
  wire h_u_arrmul32_and20_26_y0;
  wire h_u_arrmul32_fa20_26_y2;
  wire h_u_arrmul32_fa20_26_y4;
  wire h_u_arrmul32_and21_26_y0;
  wire h_u_arrmul32_fa21_26_y2;
  wire h_u_arrmul32_fa21_26_y4;
  wire h_u_arrmul32_and22_26_y0;
  wire h_u_arrmul32_fa22_26_y2;
  wire h_u_arrmul32_fa22_26_y4;
  wire h_u_arrmul32_and23_26_y0;
  wire h_u_arrmul32_fa23_26_y2;
  wire h_u_arrmul32_fa23_26_y4;
  wire h_u_arrmul32_and24_26_y0;
  wire h_u_arrmul32_fa24_26_y2;
  wire h_u_arrmul32_fa24_26_y4;
  wire h_u_arrmul32_and25_26_y0;
  wire h_u_arrmul32_fa25_26_y2;
  wire h_u_arrmul32_fa25_26_y4;
  wire h_u_arrmul32_and26_26_y0;
  wire h_u_arrmul32_fa26_26_y2;
  wire h_u_arrmul32_fa26_26_y4;
  wire h_u_arrmul32_and27_26_y0;
  wire h_u_arrmul32_fa27_26_y2;
  wire h_u_arrmul32_fa27_26_y4;
  wire h_u_arrmul32_and28_26_y0;
  wire h_u_arrmul32_fa28_26_y2;
  wire h_u_arrmul32_fa28_26_y4;
  wire h_u_arrmul32_and29_26_y0;
  wire h_u_arrmul32_fa29_26_y2;
  wire h_u_arrmul32_fa29_26_y4;
  wire h_u_arrmul32_and30_26_y0;
  wire h_u_arrmul32_fa30_26_y2;
  wire h_u_arrmul32_fa30_26_y4;
  wire h_u_arrmul32_and31_26_y0;
  wire h_u_arrmul32_fa31_26_y2;
  wire h_u_arrmul32_fa31_26_y4;
  wire h_u_arrmul32_and0_27_y0;
  wire h_u_arrmul32_ha0_27_y0;
  wire h_u_arrmul32_ha0_27_y1;
  wire h_u_arrmul32_and1_27_y0;
  wire h_u_arrmul32_fa1_27_y2;
  wire h_u_arrmul32_fa1_27_y4;
  wire h_u_arrmul32_and2_27_y0;
  wire h_u_arrmul32_fa2_27_y2;
  wire h_u_arrmul32_fa2_27_y4;
  wire h_u_arrmul32_and3_27_y0;
  wire h_u_arrmul32_fa3_27_y2;
  wire h_u_arrmul32_fa3_27_y4;
  wire h_u_arrmul32_and4_27_y0;
  wire h_u_arrmul32_fa4_27_y2;
  wire h_u_arrmul32_fa4_27_y4;
  wire h_u_arrmul32_and5_27_y0;
  wire h_u_arrmul32_fa5_27_y2;
  wire h_u_arrmul32_fa5_27_y4;
  wire h_u_arrmul32_and6_27_y0;
  wire h_u_arrmul32_fa6_27_y2;
  wire h_u_arrmul32_fa6_27_y4;
  wire h_u_arrmul32_and7_27_y0;
  wire h_u_arrmul32_fa7_27_y2;
  wire h_u_arrmul32_fa7_27_y4;
  wire h_u_arrmul32_and8_27_y0;
  wire h_u_arrmul32_fa8_27_y2;
  wire h_u_arrmul32_fa8_27_y4;
  wire h_u_arrmul32_and9_27_y0;
  wire h_u_arrmul32_fa9_27_y2;
  wire h_u_arrmul32_fa9_27_y4;
  wire h_u_arrmul32_and10_27_y0;
  wire h_u_arrmul32_fa10_27_y2;
  wire h_u_arrmul32_fa10_27_y4;
  wire h_u_arrmul32_and11_27_y0;
  wire h_u_arrmul32_fa11_27_y2;
  wire h_u_arrmul32_fa11_27_y4;
  wire h_u_arrmul32_and12_27_y0;
  wire h_u_arrmul32_fa12_27_y2;
  wire h_u_arrmul32_fa12_27_y4;
  wire h_u_arrmul32_and13_27_y0;
  wire h_u_arrmul32_fa13_27_y2;
  wire h_u_arrmul32_fa13_27_y4;
  wire h_u_arrmul32_and14_27_y0;
  wire h_u_arrmul32_fa14_27_y2;
  wire h_u_arrmul32_fa14_27_y4;
  wire h_u_arrmul32_and15_27_y0;
  wire h_u_arrmul32_fa15_27_y2;
  wire h_u_arrmul32_fa15_27_y4;
  wire h_u_arrmul32_and16_27_y0;
  wire h_u_arrmul32_fa16_27_y2;
  wire h_u_arrmul32_fa16_27_y4;
  wire h_u_arrmul32_and17_27_y0;
  wire h_u_arrmul32_fa17_27_y2;
  wire h_u_arrmul32_fa17_27_y4;
  wire h_u_arrmul32_and18_27_y0;
  wire h_u_arrmul32_fa18_27_y2;
  wire h_u_arrmul32_fa18_27_y4;
  wire h_u_arrmul32_and19_27_y0;
  wire h_u_arrmul32_fa19_27_y2;
  wire h_u_arrmul32_fa19_27_y4;
  wire h_u_arrmul32_and20_27_y0;
  wire h_u_arrmul32_fa20_27_y2;
  wire h_u_arrmul32_fa20_27_y4;
  wire h_u_arrmul32_and21_27_y0;
  wire h_u_arrmul32_fa21_27_y2;
  wire h_u_arrmul32_fa21_27_y4;
  wire h_u_arrmul32_and22_27_y0;
  wire h_u_arrmul32_fa22_27_y2;
  wire h_u_arrmul32_fa22_27_y4;
  wire h_u_arrmul32_and23_27_y0;
  wire h_u_arrmul32_fa23_27_y2;
  wire h_u_arrmul32_fa23_27_y4;
  wire h_u_arrmul32_and24_27_y0;
  wire h_u_arrmul32_fa24_27_y2;
  wire h_u_arrmul32_fa24_27_y4;
  wire h_u_arrmul32_and25_27_y0;
  wire h_u_arrmul32_fa25_27_y2;
  wire h_u_arrmul32_fa25_27_y4;
  wire h_u_arrmul32_and26_27_y0;
  wire h_u_arrmul32_fa26_27_y2;
  wire h_u_arrmul32_fa26_27_y4;
  wire h_u_arrmul32_and27_27_y0;
  wire h_u_arrmul32_fa27_27_y2;
  wire h_u_arrmul32_fa27_27_y4;
  wire h_u_arrmul32_and28_27_y0;
  wire h_u_arrmul32_fa28_27_y2;
  wire h_u_arrmul32_fa28_27_y4;
  wire h_u_arrmul32_and29_27_y0;
  wire h_u_arrmul32_fa29_27_y2;
  wire h_u_arrmul32_fa29_27_y4;
  wire h_u_arrmul32_and30_27_y0;
  wire h_u_arrmul32_fa30_27_y2;
  wire h_u_arrmul32_fa30_27_y4;
  wire h_u_arrmul32_and31_27_y0;
  wire h_u_arrmul32_fa31_27_y2;
  wire h_u_arrmul32_fa31_27_y4;
  wire h_u_arrmul32_and0_28_y0;
  wire h_u_arrmul32_ha0_28_y0;
  wire h_u_arrmul32_ha0_28_y1;
  wire h_u_arrmul32_and1_28_y0;
  wire h_u_arrmul32_fa1_28_y2;
  wire h_u_arrmul32_fa1_28_y4;
  wire h_u_arrmul32_and2_28_y0;
  wire h_u_arrmul32_fa2_28_y2;
  wire h_u_arrmul32_fa2_28_y4;
  wire h_u_arrmul32_and3_28_y0;
  wire h_u_arrmul32_fa3_28_y2;
  wire h_u_arrmul32_fa3_28_y4;
  wire h_u_arrmul32_and4_28_y0;
  wire h_u_arrmul32_fa4_28_y2;
  wire h_u_arrmul32_fa4_28_y4;
  wire h_u_arrmul32_and5_28_y0;
  wire h_u_arrmul32_fa5_28_y2;
  wire h_u_arrmul32_fa5_28_y4;
  wire h_u_arrmul32_and6_28_y0;
  wire h_u_arrmul32_fa6_28_y2;
  wire h_u_arrmul32_fa6_28_y4;
  wire h_u_arrmul32_and7_28_y0;
  wire h_u_arrmul32_fa7_28_y2;
  wire h_u_arrmul32_fa7_28_y4;
  wire h_u_arrmul32_and8_28_y0;
  wire h_u_arrmul32_fa8_28_y2;
  wire h_u_arrmul32_fa8_28_y4;
  wire h_u_arrmul32_and9_28_y0;
  wire h_u_arrmul32_fa9_28_y2;
  wire h_u_arrmul32_fa9_28_y4;
  wire h_u_arrmul32_and10_28_y0;
  wire h_u_arrmul32_fa10_28_y2;
  wire h_u_arrmul32_fa10_28_y4;
  wire h_u_arrmul32_and11_28_y0;
  wire h_u_arrmul32_fa11_28_y2;
  wire h_u_arrmul32_fa11_28_y4;
  wire h_u_arrmul32_and12_28_y0;
  wire h_u_arrmul32_fa12_28_y2;
  wire h_u_arrmul32_fa12_28_y4;
  wire h_u_arrmul32_and13_28_y0;
  wire h_u_arrmul32_fa13_28_y2;
  wire h_u_arrmul32_fa13_28_y4;
  wire h_u_arrmul32_and14_28_y0;
  wire h_u_arrmul32_fa14_28_y2;
  wire h_u_arrmul32_fa14_28_y4;
  wire h_u_arrmul32_and15_28_y0;
  wire h_u_arrmul32_fa15_28_y2;
  wire h_u_arrmul32_fa15_28_y4;
  wire h_u_arrmul32_and16_28_y0;
  wire h_u_arrmul32_fa16_28_y2;
  wire h_u_arrmul32_fa16_28_y4;
  wire h_u_arrmul32_and17_28_y0;
  wire h_u_arrmul32_fa17_28_y2;
  wire h_u_arrmul32_fa17_28_y4;
  wire h_u_arrmul32_and18_28_y0;
  wire h_u_arrmul32_fa18_28_y2;
  wire h_u_arrmul32_fa18_28_y4;
  wire h_u_arrmul32_and19_28_y0;
  wire h_u_arrmul32_fa19_28_y2;
  wire h_u_arrmul32_fa19_28_y4;
  wire h_u_arrmul32_and20_28_y0;
  wire h_u_arrmul32_fa20_28_y2;
  wire h_u_arrmul32_fa20_28_y4;
  wire h_u_arrmul32_and21_28_y0;
  wire h_u_arrmul32_fa21_28_y2;
  wire h_u_arrmul32_fa21_28_y4;
  wire h_u_arrmul32_and22_28_y0;
  wire h_u_arrmul32_fa22_28_y2;
  wire h_u_arrmul32_fa22_28_y4;
  wire h_u_arrmul32_and23_28_y0;
  wire h_u_arrmul32_fa23_28_y2;
  wire h_u_arrmul32_fa23_28_y4;
  wire h_u_arrmul32_and24_28_y0;
  wire h_u_arrmul32_fa24_28_y2;
  wire h_u_arrmul32_fa24_28_y4;
  wire h_u_arrmul32_and25_28_y0;
  wire h_u_arrmul32_fa25_28_y2;
  wire h_u_arrmul32_fa25_28_y4;
  wire h_u_arrmul32_and26_28_y0;
  wire h_u_arrmul32_fa26_28_y2;
  wire h_u_arrmul32_fa26_28_y4;
  wire h_u_arrmul32_and27_28_y0;
  wire h_u_arrmul32_fa27_28_y2;
  wire h_u_arrmul32_fa27_28_y4;
  wire h_u_arrmul32_and28_28_y0;
  wire h_u_arrmul32_fa28_28_y2;
  wire h_u_arrmul32_fa28_28_y4;
  wire h_u_arrmul32_and29_28_y0;
  wire h_u_arrmul32_fa29_28_y2;
  wire h_u_arrmul32_fa29_28_y4;
  wire h_u_arrmul32_and30_28_y0;
  wire h_u_arrmul32_fa30_28_y2;
  wire h_u_arrmul32_fa30_28_y4;
  wire h_u_arrmul32_and31_28_y0;
  wire h_u_arrmul32_fa31_28_y2;
  wire h_u_arrmul32_fa31_28_y4;
  wire h_u_arrmul32_and0_29_y0;
  wire h_u_arrmul32_ha0_29_y0;
  wire h_u_arrmul32_ha0_29_y1;
  wire h_u_arrmul32_and1_29_y0;
  wire h_u_arrmul32_fa1_29_y2;
  wire h_u_arrmul32_fa1_29_y4;
  wire h_u_arrmul32_and2_29_y0;
  wire h_u_arrmul32_fa2_29_y2;
  wire h_u_arrmul32_fa2_29_y4;
  wire h_u_arrmul32_and3_29_y0;
  wire h_u_arrmul32_fa3_29_y2;
  wire h_u_arrmul32_fa3_29_y4;
  wire h_u_arrmul32_and4_29_y0;
  wire h_u_arrmul32_fa4_29_y2;
  wire h_u_arrmul32_fa4_29_y4;
  wire h_u_arrmul32_and5_29_y0;
  wire h_u_arrmul32_fa5_29_y2;
  wire h_u_arrmul32_fa5_29_y4;
  wire h_u_arrmul32_and6_29_y0;
  wire h_u_arrmul32_fa6_29_y2;
  wire h_u_arrmul32_fa6_29_y4;
  wire h_u_arrmul32_and7_29_y0;
  wire h_u_arrmul32_fa7_29_y2;
  wire h_u_arrmul32_fa7_29_y4;
  wire h_u_arrmul32_and8_29_y0;
  wire h_u_arrmul32_fa8_29_y2;
  wire h_u_arrmul32_fa8_29_y4;
  wire h_u_arrmul32_and9_29_y0;
  wire h_u_arrmul32_fa9_29_y2;
  wire h_u_arrmul32_fa9_29_y4;
  wire h_u_arrmul32_and10_29_y0;
  wire h_u_arrmul32_fa10_29_y2;
  wire h_u_arrmul32_fa10_29_y4;
  wire h_u_arrmul32_and11_29_y0;
  wire h_u_arrmul32_fa11_29_y2;
  wire h_u_arrmul32_fa11_29_y4;
  wire h_u_arrmul32_and12_29_y0;
  wire h_u_arrmul32_fa12_29_y2;
  wire h_u_arrmul32_fa12_29_y4;
  wire h_u_arrmul32_and13_29_y0;
  wire h_u_arrmul32_fa13_29_y2;
  wire h_u_arrmul32_fa13_29_y4;
  wire h_u_arrmul32_and14_29_y0;
  wire h_u_arrmul32_fa14_29_y2;
  wire h_u_arrmul32_fa14_29_y4;
  wire h_u_arrmul32_and15_29_y0;
  wire h_u_arrmul32_fa15_29_y2;
  wire h_u_arrmul32_fa15_29_y4;
  wire h_u_arrmul32_and16_29_y0;
  wire h_u_arrmul32_fa16_29_y2;
  wire h_u_arrmul32_fa16_29_y4;
  wire h_u_arrmul32_and17_29_y0;
  wire h_u_arrmul32_fa17_29_y2;
  wire h_u_arrmul32_fa17_29_y4;
  wire h_u_arrmul32_and18_29_y0;
  wire h_u_arrmul32_fa18_29_y2;
  wire h_u_arrmul32_fa18_29_y4;
  wire h_u_arrmul32_and19_29_y0;
  wire h_u_arrmul32_fa19_29_y2;
  wire h_u_arrmul32_fa19_29_y4;
  wire h_u_arrmul32_and20_29_y0;
  wire h_u_arrmul32_fa20_29_y2;
  wire h_u_arrmul32_fa20_29_y4;
  wire h_u_arrmul32_and21_29_y0;
  wire h_u_arrmul32_fa21_29_y2;
  wire h_u_arrmul32_fa21_29_y4;
  wire h_u_arrmul32_and22_29_y0;
  wire h_u_arrmul32_fa22_29_y2;
  wire h_u_arrmul32_fa22_29_y4;
  wire h_u_arrmul32_and23_29_y0;
  wire h_u_arrmul32_fa23_29_y2;
  wire h_u_arrmul32_fa23_29_y4;
  wire h_u_arrmul32_and24_29_y0;
  wire h_u_arrmul32_fa24_29_y2;
  wire h_u_arrmul32_fa24_29_y4;
  wire h_u_arrmul32_and25_29_y0;
  wire h_u_arrmul32_fa25_29_y2;
  wire h_u_arrmul32_fa25_29_y4;
  wire h_u_arrmul32_and26_29_y0;
  wire h_u_arrmul32_fa26_29_y2;
  wire h_u_arrmul32_fa26_29_y4;
  wire h_u_arrmul32_and27_29_y0;
  wire h_u_arrmul32_fa27_29_y2;
  wire h_u_arrmul32_fa27_29_y4;
  wire h_u_arrmul32_and28_29_y0;
  wire h_u_arrmul32_fa28_29_y2;
  wire h_u_arrmul32_fa28_29_y4;
  wire h_u_arrmul32_and29_29_y0;
  wire h_u_arrmul32_fa29_29_y2;
  wire h_u_arrmul32_fa29_29_y4;
  wire h_u_arrmul32_and30_29_y0;
  wire h_u_arrmul32_fa30_29_y2;
  wire h_u_arrmul32_fa30_29_y4;
  wire h_u_arrmul32_and31_29_y0;
  wire h_u_arrmul32_fa31_29_y2;
  wire h_u_arrmul32_fa31_29_y4;
  wire h_u_arrmul32_and0_30_y0;
  wire h_u_arrmul32_ha0_30_y0;
  wire h_u_arrmul32_ha0_30_y1;
  wire h_u_arrmul32_and1_30_y0;
  wire h_u_arrmul32_fa1_30_y2;
  wire h_u_arrmul32_fa1_30_y4;
  wire h_u_arrmul32_and2_30_y0;
  wire h_u_arrmul32_fa2_30_y2;
  wire h_u_arrmul32_fa2_30_y4;
  wire h_u_arrmul32_and3_30_y0;
  wire h_u_arrmul32_fa3_30_y2;
  wire h_u_arrmul32_fa3_30_y4;
  wire h_u_arrmul32_and4_30_y0;
  wire h_u_arrmul32_fa4_30_y2;
  wire h_u_arrmul32_fa4_30_y4;
  wire h_u_arrmul32_and5_30_y0;
  wire h_u_arrmul32_fa5_30_y2;
  wire h_u_arrmul32_fa5_30_y4;
  wire h_u_arrmul32_and6_30_y0;
  wire h_u_arrmul32_fa6_30_y2;
  wire h_u_arrmul32_fa6_30_y4;
  wire h_u_arrmul32_and7_30_y0;
  wire h_u_arrmul32_fa7_30_y2;
  wire h_u_arrmul32_fa7_30_y4;
  wire h_u_arrmul32_and8_30_y0;
  wire h_u_arrmul32_fa8_30_y2;
  wire h_u_arrmul32_fa8_30_y4;
  wire h_u_arrmul32_and9_30_y0;
  wire h_u_arrmul32_fa9_30_y2;
  wire h_u_arrmul32_fa9_30_y4;
  wire h_u_arrmul32_and10_30_y0;
  wire h_u_arrmul32_fa10_30_y2;
  wire h_u_arrmul32_fa10_30_y4;
  wire h_u_arrmul32_and11_30_y0;
  wire h_u_arrmul32_fa11_30_y2;
  wire h_u_arrmul32_fa11_30_y4;
  wire h_u_arrmul32_and12_30_y0;
  wire h_u_arrmul32_fa12_30_y2;
  wire h_u_arrmul32_fa12_30_y4;
  wire h_u_arrmul32_and13_30_y0;
  wire h_u_arrmul32_fa13_30_y2;
  wire h_u_arrmul32_fa13_30_y4;
  wire h_u_arrmul32_and14_30_y0;
  wire h_u_arrmul32_fa14_30_y2;
  wire h_u_arrmul32_fa14_30_y4;
  wire h_u_arrmul32_and15_30_y0;
  wire h_u_arrmul32_fa15_30_y2;
  wire h_u_arrmul32_fa15_30_y4;
  wire h_u_arrmul32_and16_30_y0;
  wire h_u_arrmul32_fa16_30_y2;
  wire h_u_arrmul32_fa16_30_y4;
  wire h_u_arrmul32_and17_30_y0;
  wire h_u_arrmul32_fa17_30_y2;
  wire h_u_arrmul32_fa17_30_y4;
  wire h_u_arrmul32_and18_30_y0;
  wire h_u_arrmul32_fa18_30_y2;
  wire h_u_arrmul32_fa18_30_y4;
  wire h_u_arrmul32_and19_30_y0;
  wire h_u_arrmul32_fa19_30_y2;
  wire h_u_arrmul32_fa19_30_y4;
  wire h_u_arrmul32_and20_30_y0;
  wire h_u_arrmul32_fa20_30_y2;
  wire h_u_arrmul32_fa20_30_y4;
  wire h_u_arrmul32_and21_30_y0;
  wire h_u_arrmul32_fa21_30_y2;
  wire h_u_arrmul32_fa21_30_y4;
  wire h_u_arrmul32_and22_30_y0;
  wire h_u_arrmul32_fa22_30_y2;
  wire h_u_arrmul32_fa22_30_y4;
  wire h_u_arrmul32_and23_30_y0;
  wire h_u_arrmul32_fa23_30_y2;
  wire h_u_arrmul32_fa23_30_y4;
  wire h_u_arrmul32_and24_30_y0;
  wire h_u_arrmul32_fa24_30_y2;
  wire h_u_arrmul32_fa24_30_y4;
  wire h_u_arrmul32_and25_30_y0;
  wire h_u_arrmul32_fa25_30_y2;
  wire h_u_arrmul32_fa25_30_y4;
  wire h_u_arrmul32_and26_30_y0;
  wire h_u_arrmul32_fa26_30_y2;
  wire h_u_arrmul32_fa26_30_y4;
  wire h_u_arrmul32_and27_30_y0;
  wire h_u_arrmul32_fa27_30_y2;
  wire h_u_arrmul32_fa27_30_y4;
  wire h_u_arrmul32_and28_30_y0;
  wire h_u_arrmul32_fa28_30_y2;
  wire h_u_arrmul32_fa28_30_y4;
  wire h_u_arrmul32_and29_30_y0;
  wire h_u_arrmul32_fa29_30_y2;
  wire h_u_arrmul32_fa29_30_y4;
  wire h_u_arrmul32_and30_30_y0;
  wire h_u_arrmul32_fa30_30_y2;
  wire h_u_arrmul32_fa30_30_y4;
  wire h_u_arrmul32_and31_30_y0;
  wire h_u_arrmul32_fa31_30_y2;
  wire h_u_arrmul32_fa31_30_y4;
  wire h_u_arrmul32_and0_31_y0;
  wire h_u_arrmul32_ha0_31_y0;
  wire h_u_arrmul32_ha0_31_y1;
  wire h_u_arrmul32_and1_31_y0;
  wire h_u_arrmul32_fa1_31_y2;
  wire h_u_arrmul32_fa1_31_y4;
  wire h_u_arrmul32_and2_31_y0;
  wire h_u_arrmul32_fa2_31_y2;
  wire h_u_arrmul32_fa2_31_y4;
  wire h_u_arrmul32_and3_31_y0;
  wire h_u_arrmul32_fa3_31_y2;
  wire h_u_arrmul32_fa3_31_y4;
  wire h_u_arrmul32_and4_31_y0;
  wire h_u_arrmul32_fa4_31_y2;
  wire h_u_arrmul32_fa4_31_y4;
  wire h_u_arrmul32_and5_31_y0;
  wire h_u_arrmul32_fa5_31_y2;
  wire h_u_arrmul32_fa5_31_y4;
  wire h_u_arrmul32_and6_31_y0;
  wire h_u_arrmul32_fa6_31_y2;
  wire h_u_arrmul32_fa6_31_y4;
  wire h_u_arrmul32_and7_31_y0;
  wire h_u_arrmul32_fa7_31_y2;
  wire h_u_arrmul32_fa7_31_y4;
  wire h_u_arrmul32_and8_31_y0;
  wire h_u_arrmul32_fa8_31_y2;
  wire h_u_arrmul32_fa8_31_y4;
  wire h_u_arrmul32_and9_31_y0;
  wire h_u_arrmul32_fa9_31_y2;
  wire h_u_arrmul32_fa9_31_y4;
  wire h_u_arrmul32_and10_31_y0;
  wire h_u_arrmul32_fa10_31_y2;
  wire h_u_arrmul32_fa10_31_y4;
  wire h_u_arrmul32_and11_31_y0;
  wire h_u_arrmul32_fa11_31_y2;
  wire h_u_arrmul32_fa11_31_y4;
  wire h_u_arrmul32_and12_31_y0;
  wire h_u_arrmul32_fa12_31_y2;
  wire h_u_arrmul32_fa12_31_y4;
  wire h_u_arrmul32_and13_31_y0;
  wire h_u_arrmul32_fa13_31_y2;
  wire h_u_arrmul32_fa13_31_y4;
  wire h_u_arrmul32_and14_31_y0;
  wire h_u_arrmul32_fa14_31_y2;
  wire h_u_arrmul32_fa14_31_y4;
  wire h_u_arrmul32_and15_31_y0;
  wire h_u_arrmul32_fa15_31_y2;
  wire h_u_arrmul32_fa15_31_y4;
  wire h_u_arrmul32_and16_31_y0;
  wire h_u_arrmul32_fa16_31_y2;
  wire h_u_arrmul32_fa16_31_y4;
  wire h_u_arrmul32_and17_31_y0;
  wire h_u_arrmul32_fa17_31_y2;
  wire h_u_arrmul32_fa17_31_y4;
  wire h_u_arrmul32_and18_31_y0;
  wire h_u_arrmul32_fa18_31_y2;
  wire h_u_arrmul32_fa18_31_y4;
  wire h_u_arrmul32_and19_31_y0;
  wire h_u_arrmul32_fa19_31_y2;
  wire h_u_arrmul32_fa19_31_y4;
  wire h_u_arrmul32_and20_31_y0;
  wire h_u_arrmul32_fa20_31_y2;
  wire h_u_arrmul32_fa20_31_y4;
  wire h_u_arrmul32_and21_31_y0;
  wire h_u_arrmul32_fa21_31_y2;
  wire h_u_arrmul32_fa21_31_y4;
  wire h_u_arrmul32_and22_31_y0;
  wire h_u_arrmul32_fa22_31_y2;
  wire h_u_arrmul32_fa22_31_y4;
  wire h_u_arrmul32_and23_31_y0;
  wire h_u_arrmul32_fa23_31_y2;
  wire h_u_arrmul32_fa23_31_y4;
  wire h_u_arrmul32_and24_31_y0;
  wire h_u_arrmul32_fa24_31_y2;
  wire h_u_arrmul32_fa24_31_y4;
  wire h_u_arrmul32_and25_31_y0;
  wire h_u_arrmul32_fa25_31_y2;
  wire h_u_arrmul32_fa25_31_y4;
  wire h_u_arrmul32_and26_31_y0;
  wire h_u_arrmul32_fa26_31_y2;
  wire h_u_arrmul32_fa26_31_y4;
  wire h_u_arrmul32_and27_31_y0;
  wire h_u_arrmul32_fa27_31_y2;
  wire h_u_arrmul32_fa27_31_y4;
  wire h_u_arrmul32_and28_31_y0;
  wire h_u_arrmul32_fa28_31_y2;
  wire h_u_arrmul32_fa28_31_y4;
  wire h_u_arrmul32_and29_31_y0;
  wire h_u_arrmul32_fa29_31_y2;
  wire h_u_arrmul32_fa29_31_y4;
  wire h_u_arrmul32_and30_31_y0;
  wire h_u_arrmul32_fa30_31_y2;
  wire h_u_arrmul32_fa30_31_y4;
  wire h_u_arrmul32_and31_31_y0;
  wire h_u_arrmul32_fa31_31_y2;
  wire h_u_arrmul32_fa31_31_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign a_30 = a[30];
  assign a_31 = a[31];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  assign b_30 = b[30];
  assign b_31 = b[31];
  and_gate and_gate_h_u_arrmul32_and0_0_y0(a_0, b_0, h_u_arrmul32_and0_0_y0);
  and_gate and_gate_h_u_arrmul32_and1_0_y0(a_1, b_0, h_u_arrmul32_and1_0_y0);
  and_gate and_gate_h_u_arrmul32_and2_0_y0(a_2, b_0, h_u_arrmul32_and2_0_y0);
  and_gate and_gate_h_u_arrmul32_and3_0_y0(a_3, b_0, h_u_arrmul32_and3_0_y0);
  and_gate and_gate_h_u_arrmul32_and4_0_y0(a_4, b_0, h_u_arrmul32_and4_0_y0);
  and_gate and_gate_h_u_arrmul32_and5_0_y0(a_5, b_0, h_u_arrmul32_and5_0_y0);
  and_gate and_gate_h_u_arrmul32_and6_0_y0(a_6, b_0, h_u_arrmul32_and6_0_y0);
  and_gate and_gate_h_u_arrmul32_and7_0_y0(a_7, b_0, h_u_arrmul32_and7_0_y0);
  and_gate and_gate_h_u_arrmul32_and8_0_y0(a_8, b_0, h_u_arrmul32_and8_0_y0);
  and_gate and_gate_h_u_arrmul32_and9_0_y0(a_9, b_0, h_u_arrmul32_and9_0_y0);
  and_gate and_gate_h_u_arrmul32_and10_0_y0(a_10, b_0, h_u_arrmul32_and10_0_y0);
  and_gate and_gate_h_u_arrmul32_and11_0_y0(a_11, b_0, h_u_arrmul32_and11_0_y0);
  and_gate and_gate_h_u_arrmul32_and12_0_y0(a_12, b_0, h_u_arrmul32_and12_0_y0);
  and_gate and_gate_h_u_arrmul32_and13_0_y0(a_13, b_0, h_u_arrmul32_and13_0_y0);
  and_gate and_gate_h_u_arrmul32_and14_0_y0(a_14, b_0, h_u_arrmul32_and14_0_y0);
  and_gate and_gate_h_u_arrmul32_and15_0_y0(a_15, b_0, h_u_arrmul32_and15_0_y0);
  and_gate and_gate_h_u_arrmul32_and16_0_y0(a_16, b_0, h_u_arrmul32_and16_0_y0);
  and_gate and_gate_h_u_arrmul32_and17_0_y0(a_17, b_0, h_u_arrmul32_and17_0_y0);
  and_gate and_gate_h_u_arrmul32_and18_0_y0(a_18, b_0, h_u_arrmul32_and18_0_y0);
  and_gate and_gate_h_u_arrmul32_and19_0_y0(a_19, b_0, h_u_arrmul32_and19_0_y0);
  and_gate and_gate_h_u_arrmul32_and20_0_y0(a_20, b_0, h_u_arrmul32_and20_0_y0);
  and_gate and_gate_h_u_arrmul32_and21_0_y0(a_21, b_0, h_u_arrmul32_and21_0_y0);
  and_gate and_gate_h_u_arrmul32_and22_0_y0(a_22, b_0, h_u_arrmul32_and22_0_y0);
  and_gate and_gate_h_u_arrmul32_and23_0_y0(a_23, b_0, h_u_arrmul32_and23_0_y0);
  and_gate and_gate_h_u_arrmul32_and24_0_y0(a_24, b_0, h_u_arrmul32_and24_0_y0);
  and_gate and_gate_h_u_arrmul32_and25_0_y0(a_25, b_0, h_u_arrmul32_and25_0_y0);
  and_gate and_gate_h_u_arrmul32_and26_0_y0(a_26, b_0, h_u_arrmul32_and26_0_y0);
  and_gate and_gate_h_u_arrmul32_and27_0_y0(a_27, b_0, h_u_arrmul32_and27_0_y0);
  and_gate and_gate_h_u_arrmul32_and28_0_y0(a_28, b_0, h_u_arrmul32_and28_0_y0);
  and_gate and_gate_h_u_arrmul32_and29_0_y0(a_29, b_0, h_u_arrmul32_and29_0_y0);
  and_gate and_gate_h_u_arrmul32_and30_0_y0(a_30, b_0, h_u_arrmul32_and30_0_y0);
  and_gate and_gate_h_u_arrmul32_and31_0_y0(a_31, b_0, h_u_arrmul32_and31_0_y0);
  and_gate and_gate_h_u_arrmul32_and0_1_y0(a_0, b_1, h_u_arrmul32_and0_1_y0);
  ha ha_h_u_arrmul32_ha0_1_y0(h_u_arrmul32_and0_1_y0, h_u_arrmul32_and1_0_y0, h_u_arrmul32_ha0_1_y0, h_u_arrmul32_ha0_1_y1);
  and_gate and_gate_h_u_arrmul32_and1_1_y0(a_1, b_1, h_u_arrmul32_and1_1_y0);
  fa fa_h_u_arrmul32_fa1_1_y2(h_u_arrmul32_and1_1_y0, h_u_arrmul32_and2_0_y0, h_u_arrmul32_ha0_1_y1, h_u_arrmul32_fa1_1_y2, h_u_arrmul32_fa1_1_y4);
  and_gate and_gate_h_u_arrmul32_and2_1_y0(a_2, b_1, h_u_arrmul32_and2_1_y0);
  fa fa_h_u_arrmul32_fa2_1_y2(h_u_arrmul32_and2_1_y0, h_u_arrmul32_and3_0_y0, h_u_arrmul32_fa1_1_y4, h_u_arrmul32_fa2_1_y2, h_u_arrmul32_fa2_1_y4);
  and_gate and_gate_h_u_arrmul32_and3_1_y0(a_3, b_1, h_u_arrmul32_and3_1_y0);
  fa fa_h_u_arrmul32_fa3_1_y2(h_u_arrmul32_and3_1_y0, h_u_arrmul32_and4_0_y0, h_u_arrmul32_fa2_1_y4, h_u_arrmul32_fa3_1_y2, h_u_arrmul32_fa3_1_y4);
  and_gate and_gate_h_u_arrmul32_and4_1_y0(a_4, b_1, h_u_arrmul32_and4_1_y0);
  fa fa_h_u_arrmul32_fa4_1_y2(h_u_arrmul32_and4_1_y0, h_u_arrmul32_and5_0_y0, h_u_arrmul32_fa3_1_y4, h_u_arrmul32_fa4_1_y2, h_u_arrmul32_fa4_1_y4);
  and_gate and_gate_h_u_arrmul32_and5_1_y0(a_5, b_1, h_u_arrmul32_and5_1_y0);
  fa fa_h_u_arrmul32_fa5_1_y2(h_u_arrmul32_and5_1_y0, h_u_arrmul32_and6_0_y0, h_u_arrmul32_fa4_1_y4, h_u_arrmul32_fa5_1_y2, h_u_arrmul32_fa5_1_y4);
  and_gate and_gate_h_u_arrmul32_and6_1_y0(a_6, b_1, h_u_arrmul32_and6_1_y0);
  fa fa_h_u_arrmul32_fa6_1_y2(h_u_arrmul32_and6_1_y0, h_u_arrmul32_and7_0_y0, h_u_arrmul32_fa5_1_y4, h_u_arrmul32_fa6_1_y2, h_u_arrmul32_fa6_1_y4);
  and_gate and_gate_h_u_arrmul32_and7_1_y0(a_7, b_1, h_u_arrmul32_and7_1_y0);
  fa fa_h_u_arrmul32_fa7_1_y2(h_u_arrmul32_and7_1_y0, h_u_arrmul32_and8_0_y0, h_u_arrmul32_fa6_1_y4, h_u_arrmul32_fa7_1_y2, h_u_arrmul32_fa7_1_y4);
  and_gate and_gate_h_u_arrmul32_and8_1_y0(a_8, b_1, h_u_arrmul32_and8_1_y0);
  fa fa_h_u_arrmul32_fa8_1_y2(h_u_arrmul32_and8_1_y0, h_u_arrmul32_and9_0_y0, h_u_arrmul32_fa7_1_y4, h_u_arrmul32_fa8_1_y2, h_u_arrmul32_fa8_1_y4);
  and_gate and_gate_h_u_arrmul32_and9_1_y0(a_9, b_1, h_u_arrmul32_and9_1_y0);
  fa fa_h_u_arrmul32_fa9_1_y2(h_u_arrmul32_and9_1_y0, h_u_arrmul32_and10_0_y0, h_u_arrmul32_fa8_1_y4, h_u_arrmul32_fa9_1_y2, h_u_arrmul32_fa9_1_y4);
  and_gate and_gate_h_u_arrmul32_and10_1_y0(a_10, b_1, h_u_arrmul32_and10_1_y0);
  fa fa_h_u_arrmul32_fa10_1_y2(h_u_arrmul32_and10_1_y0, h_u_arrmul32_and11_0_y0, h_u_arrmul32_fa9_1_y4, h_u_arrmul32_fa10_1_y2, h_u_arrmul32_fa10_1_y4);
  and_gate and_gate_h_u_arrmul32_and11_1_y0(a_11, b_1, h_u_arrmul32_and11_1_y0);
  fa fa_h_u_arrmul32_fa11_1_y2(h_u_arrmul32_and11_1_y0, h_u_arrmul32_and12_0_y0, h_u_arrmul32_fa10_1_y4, h_u_arrmul32_fa11_1_y2, h_u_arrmul32_fa11_1_y4);
  and_gate and_gate_h_u_arrmul32_and12_1_y0(a_12, b_1, h_u_arrmul32_and12_1_y0);
  fa fa_h_u_arrmul32_fa12_1_y2(h_u_arrmul32_and12_1_y0, h_u_arrmul32_and13_0_y0, h_u_arrmul32_fa11_1_y4, h_u_arrmul32_fa12_1_y2, h_u_arrmul32_fa12_1_y4);
  and_gate and_gate_h_u_arrmul32_and13_1_y0(a_13, b_1, h_u_arrmul32_and13_1_y0);
  fa fa_h_u_arrmul32_fa13_1_y2(h_u_arrmul32_and13_1_y0, h_u_arrmul32_and14_0_y0, h_u_arrmul32_fa12_1_y4, h_u_arrmul32_fa13_1_y2, h_u_arrmul32_fa13_1_y4);
  and_gate and_gate_h_u_arrmul32_and14_1_y0(a_14, b_1, h_u_arrmul32_and14_1_y0);
  fa fa_h_u_arrmul32_fa14_1_y2(h_u_arrmul32_and14_1_y0, h_u_arrmul32_and15_0_y0, h_u_arrmul32_fa13_1_y4, h_u_arrmul32_fa14_1_y2, h_u_arrmul32_fa14_1_y4);
  and_gate and_gate_h_u_arrmul32_and15_1_y0(a_15, b_1, h_u_arrmul32_and15_1_y0);
  fa fa_h_u_arrmul32_fa15_1_y2(h_u_arrmul32_and15_1_y0, h_u_arrmul32_and16_0_y0, h_u_arrmul32_fa14_1_y4, h_u_arrmul32_fa15_1_y2, h_u_arrmul32_fa15_1_y4);
  and_gate and_gate_h_u_arrmul32_and16_1_y0(a_16, b_1, h_u_arrmul32_and16_1_y0);
  fa fa_h_u_arrmul32_fa16_1_y2(h_u_arrmul32_and16_1_y0, h_u_arrmul32_and17_0_y0, h_u_arrmul32_fa15_1_y4, h_u_arrmul32_fa16_1_y2, h_u_arrmul32_fa16_1_y4);
  and_gate and_gate_h_u_arrmul32_and17_1_y0(a_17, b_1, h_u_arrmul32_and17_1_y0);
  fa fa_h_u_arrmul32_fa17_1_y2(h_u_arrmul32_and17_1_y0, h_u_arrmul32_and18_0_y0, h_u_arrmul32_fa16_1_y4, h_u_arrmul32_fa17_1_y2, h_u_arrmul32_fa17_1_y4);
  and_gate and_gate_h_u_arrmul32_and18_1_y0(a_18, b_1, h_u_arrmul32_and18_1_y0);
  fa fa_h_u_arrmul32_fa18_1_y2(h_u_arrmul32_and18_1_y0, h_u_arrmul32_and19_0_y0, h_u_arrmul32_fa17_1_y4, h_u_arrmul32_fa18_1_y2, h_u_arrmul32_fa18_1_y4);
  and_gate and_gate_h_u_arrmul32_and19_1_y0(a_19, b_1, h_u_arrmul32_and19_1_y0);
  fa fa_h_u_arrmul32_fa19_1_y2(h_u_arrmul32_and19_1_y0, h_u_arrmul32_and20_0_y0, h_u_arrmul32_fa18_1_y4, h_u_arrmul32_fa19_1_y2, h_u_arrmul32_fa19_1_y4);
  and_gate and_gate_h_u_arrmul32_and20_1_y0(a_20, b_1, h_u_arrmul32_and20_1_y0);
  fa fa_h_u_arrmul32_fa20_1_y2(h_u_arrmul32_and20_1_y0, h_u_arrmul32_and21_0_y0, h_u_arrmul32_fa19_1_y4, h_u_arrmul32_fa20_1_y2, h_u_arrmul32_fa20_1_y4);
  and_gate and_gate_h_u_arrmul32_and21_1_y0(a_21, b_1, h_u_arrmul32_and21_1_y0);
  fa fa_h_u_arrmul32_fa21_1_y2(h_u_arrmul32_and21_1_y0, h_u_arrmul32_and22_0_y0, h_u_arrmul32_fa20_1_y4, h_u_arrmul32_fa21_1_y2, h_u_arrmul32_fa21_1_y4);
  and_gate and_gate_h_u_arrmul32_and22_1_y0(a_22, b_1, h_u_arrmul32_and22_1_y0);
  fa fa_h_u_arrmul32_fa22_1_y2(h_u_arrmul32_and22_1_y0, h_u_arrmul32_and23_0_y0, h_u_arrmul32_fa21_1_y4, h_u_arrmul32_fa22_1_y2, h_u_arrmul32_fa22_1_y4);
  and_gate and_gate_h_u_arrmul32_and23_1_y0(a_23, b_1, h_u_arrmul32_and23_1_y0);
  fa fa_h_u_arrmul32_fa23_1_y2(h_u_arrmul32_and23_1_y0, h_u_arrmul32_and24_0_y0, h_u_arrmul32_fa22_1_y4, h_u_arrmul32_fa23_1_y2, h_u_arrmul32_fa23_1_y4);
  and_gate and_gate_h_u_arrmul32_and24_1_y0(a_24, b_1, h_u_arrmul32_and24_1_y0);
  fa fa_h_u_arrmul32_fa24_1_y2(h_u_arrmul32_and24_1_y0, h_u_arrmul32_and25_0_y0, h_u_arrmul32_fa23_1_y4, h_u_arrmul32_fa24_1_y2, h_u_arrmul32_fa24_1_y4);
  and_gate and_gate_h_u_arrmul32_and25_1_y0(a_25, b_1, h_u_arrmul32_and25_1_y0);
  fa fa_h_u_arrmul32_fa25_1_y2(h_u_arrmul32_and25_1_y0, h_u_arrmul32_and26_0_y0, h_u_arrmul32_fa24_1_y4, h_u_arrmul32_fa25_1_y2, h_u_arrmul32_fa25_1_y4);
  and_gate and_gate_h_u_arrmul32_and26_1_y0(a_26, b_1, h_u_arrmul32_and26_1_y0);
  fa fa_h_u_arrmul32_fa26_1_y2(h_u_arrmul32_and26_1_y0, h_u_arrmul32_and27_0_y0, h_u_arrmul32_fa25_1_y4, h_u_arrmul32_fa26_1_y2, h_u_arrmul32_fa26_1_y4);
  and_gate and_gate_h_u_arrmul32_and27_1_y0(a_27, b_1, h_u_arrmul32_and27_1_y0);
  fa fa_h_u_arrmul32_fa27_1_y2(h_u_arrmul32_and27_1_y0, h_u_arrmul32_and28_0_y0, h_u_arrmul32_fa26_1_y4, h_u_arrmul32_fa27_1_y2, h_u_arrmul32_fa27_1_y4);
  and_gate and_gate_h_u_arrmul32_and28_1_y0(a_28, b_1, h_u_arrmul32_and28_1_y0);
  fa fa_h_u_arrmul32_fa28_1_y2(h_u_arrmul32_and28_1_y0, h_u_arrmul32_and29_0_y0, h_u_arrmul32_fa27_1_y4, h_u_arrmul32_fa28_1_y2, h_u_arrmul32_fa28_1_y4);
  and_gate and_gate_h_u_arrmul32_and29_1_y0(a_29, b_1, h_u_arrmul32_and29_1_y0);
  fa fa_h_u_arrmul32_fa29_1_y2(h_u_arrmul32_and29_1_y0, h_u_arrmul32_and30_0_y0, h_u_arrmul32_fa28_1_y4, h_u_arrmul32_fa29_1_y2, h_u_arrmul32_fa29_1_y4);
  and_gate and_gate_h_u_arrmul32_and30_1_y0(a_30, b_1, h_u_arrmul32_and30_1_y0);
  fa fa_h_u_arrmul32_fa30_1_y2(h_u_arrmul32_and30_1_y0, h_u_arrmul32_and31_0_y0, h_u_arrmul32_fa29_1_y4, h_u_arrmul32_fa30_1_y2, h_u_arrmul32_fa30_1_y4);
  and_gate and_gate_h_u_arrmul32_and31_1_y0(a_31, b_1, h_u_arrmul32_and31_1_y0);
  ha ha_h_u_arrmul32_ha31_1_y0(h_u_arrmul32_and31_1_y0, h_u_arrmul32_fa30_1_y4, h_u_arrmul32_ha31_1_y0, h_u_arrmul32_ha31_1_y1);
  and_gate and_gate_h_u_arrmul32_and0_2_y0(a_0, b_2, h_u_arrmul32_and0_2_y0);
  ha ha_h_u_arrmul32_ha0_2_y0(h_u_arrmul32_and0_2_y0, h_u_arrmul32_fa1_1_y2, h_u_arrmul32_ha0_2_y0, h_u_arrmul32_ha0_2_y1);
  and_gate and_gate_h_u_arrmul32_and1_2_y0(a_1, b_2, h_u_arrmul32_and1_2_y0);
  fa fa_h_u_arrmul32_fa1_2_y2(h_u_arrmul32_and1_2_y0, h_u_arrmul32_fa2_1_y2, h_u_arrmul32_ha0_2_y1, h_u_arrmul32_fa1_2_y2, h_u_arrmul32_fa1_2_y4);
  and_gate and_gate_h_u_arrmul32_and2_2_y0(a_2, b_2, h_u_arrmul32_and2_2_y0);
  fa fa_h_u_arrmul32_fa2_2_y2(h_u_arrmul32_and2_2_y0, h_u_arrmul32_fa3_1_y2, h_u_arrmul32_fa1_2_y4, h_u_arrmul32_fa2_2_y2, h_u_arrmul32_fa2_2_y4);
  and_gate and_gate_h_u_arrmul32_and3_2_y0(a_3, b_2, h_u_arrmul32_and3_2_y0);
  fa fa_h_u_arrmul32_fa3_2_y2(h_u_arrmul32_and3_2_y0, h_u_arrmul32_fa4_1_y2, h_u_arrmul32_fa2_2_y4, h_u_arrmul32_fa3_2_y2, h_u_arrmul32_fa3_2_y4);
  and_gate and_gate_h_u_arrmul32_and4_2_y0(a_4, b_2, h_u_arrmul32_and4_2_y0);
  fa fa_h_u_arrmul32_fa4_2_y2(h_u_arrmul32_and4_2_y0, h_u_arrmul32_fa5_1_y2, h_u_arrmul32_fa3_2_y4, h_u_arrmul32_fa4_2_y2, h_u_arrmul32_fa4_2_y4);
  and_gate and_gate_h_u_arrmul32_and5_2_y0(a_5, b_2, h_u_arrmul32_and5_2_y0);
  fa fa_h_u_arrmul32_fa5_2_y2(h_u_arrmul32_and5_2_y0, h_u_arrmul32_fa6_1_y2, h_u_arrmul32_fa4_2_y4, h_u_arrmul32_fa5_2_y2, h_u_arrmul32_fa5_2_y4);
  and_gate and_gate_h_u_arrmul32_and6_2_y0(a_6, b_2, h_u_arrmul32_and6_2_y0);
  fa fa_h_u_arrmul32_fa6_2_y2(h_u_arrmul32_and6_2_y0, h_u_arrmul32_fa7_1_y2, h_u_arrmul32_fa5_2_y4, h_u_arrmul32_fa6_2_y2, h_u_arrmul32_fa6_2_y4);
  and_gate and_gate_h_u_arrmul32_and7_2_y0(a_7, b_2, h_u_arrmul32_and7_2_y0);
  fa fa_h_u_arrmul32_fa7_2_y2(h_u_arrmul32_and7_2_y0, h_u_arrmul32_fa8_1_y2, h_u_arrmul32_fa6_2_y4, h_u_arrmul32_fa7_2_y2, h_u_arrmul32_fa7_2_y4);
  and_gate and_gate_h_u_arrmul32_and8_2_y0(a_8, b_2, h_u_arrmul32_and8_2_y0);
  fa fa_h_u_arrmul32_fa8_2_y2(h_u_arrmul32_and8_2_y0, h_u_arrmul32_fa9_1_y2, h_u_arrmul32_fa7_2_y4, h_u_arrmul32_fa8_2_y2, h_u_arrmul32_fa8_2_y4);
  and_gate and_gate_h_u_arrmul32_and9_2_y0(a_9, b_2, h_u_arrmul32_and9_2_y0);
  fa fa_h_u_arrmul32_fa9_2_y2(h_u_arrmul32_and9_2_y0, h_u_arrmul32_fa10_1_y2, h_u_arrmul32_fa8_2_y4, h_u_arrmul32_fa9_2_y2, h_u_arrmul32_fa9_2_y4);
  and_gate and_gate_h_u_arrmul32_and10_2_y0(a_10, b_2, h_u_arrmul32_and10_2_y0);
  fa fa_h_u_arrmul32_fa10_2_y2(h_u_arrmul32_and10_2_y0, h_u_arrmul32_fa11_1_y2, h_u_arrmul32_fa9_2_y4, h_u_arrmul32_fa10_2_y2, h_u_arrmul32_fa10_2_y4);
  and_gate and_gate_h_u_arrmul32_and11_2_y0(a_11, b_2, h_u_arrmul32_and11_2_y0);
  fa fa_h_u_arrmul32_fa11_2_y2(h_u_arrmul32_and11_2_y0, h_u_arrmul32_fa12_1_y2, h_u_arrmul32_fa10_2_y4, h_u_arrmul32_fa11_2_y2, h_u_arrmul32_fa11_2_y4);
  and_gate and_gate_h_u_arrmul32_and12_2_y0(a_12, b_2, h_u_arrmul32_and12_2_y0);
  fa fa_h_u_arrmul32_fa12_2_y2(h_u_arrmul32_and12_2_y0, h_u_arrmul32_fa13_1_y2, h_u_arrmul32_fa11_2_y4, h_u_arrmul32_fa12_2_y2, h_u_arrmul32_fa12_2_y4);
  and_gate and_gate_h_u_arrmul32_and13_2_y0(a_13, b_2, h_u_arrmul32_and13_2_y0);
  fa fa_h_u_arrmul32_fa13_2_y2(h_u_arrmul32_and13_2_y0, h_u_arrmul32_fa14_1_y2, h_u_arrmul32_fa12_2_y4, h_u_arrmul32_fa13_2_y2, h_u_arrmul32_fa13_2_y4);
  and_gate and_gate_h_u_arrmul32_and14_2_y0(a_14, b_2, h_u_arrmul32_and14_2_y0);
  fa fa_h_u_arrmul32_fa14_2_y2(h_u_arrmul32_and14_2_y0, h_u_arrmul32_fa15_1_y2, h_u_arrmul32_fa13_2_y4, h_u_arrmul32_fa14_2_y2, h_u_arrmul32_fa14_2_y4);
  and_gate and_gate_h_u_arrmul32_and15_2_y0(a_15, b_2, h_u_arrmul32_and15_2_y0);
  fa fa_h_u_arrmul32_fa15_2_y2(h_u_arrmul32_and15_2_y0, h_u_arrmul32_fa16_1_y2, h_u_arrmul32_fa14_2_y4, h_u_arrmul32_fa15_2_y2, h_u_arrmul32_fa15_2_y4);
  and_gate and_gate_h_u_arrmul32_and16_2_y0(a_16, b_2, h_u_arrmul32_and16_2_y0);
  fa fa_h_u_arrmul32_fa16_2_y2(h_u_arrmul32_and16_2_y0, h_u_arrmul32_fa17_1_y2, h_u_arrmul32_fa15_2_y4, h_u_arrmul32_fa16_2_y2, h_u_arrmul32_fa16_2_y4);
  and_gate and_gate_h_u_arrmul32_and17_2_y0(a_17, b_2, h_u_arrmul32_and17_2_y0);
  fa fa_h_u_arrmul32_fa17_2_y2(h_u_arrmul32_and17_2_y0, h_u_arrmul32_fa18_1_y2, h_u_arrmul32_fa16_2_y4, h_u_arrmul32_fa17_2_y2, h_u_arrmul32_fa17_2_y4);
  and_gate and_gate_h_u_arrmul32_and18_2_y0(a_18, b_2, h_u_arrmul32_and18_2_y0);
  fa fa_h_u_arrmul32_fa18_2_y2(h_u_arrmul32_and18_2_y0, h_u_arrmul32_fa19_1_y2, h_u_arrmul32_fa17_2_y4, h_u_arrmul32_fa18_2_y2, h_u_arrmul32_fa18_2_y4);
  and_gate and_gate_h_u_arrmul32_and19_2_y0(a_19, b_2, h_u_arrmul32_and19_2_y0);
  fa fa_h_u_arrmul32_fa19_2_y2(h_u_arrmul32_and19_2_y0, h_u_arrmul32_fa20_1_y2, h_u_arrmul32_fa18_2_y4, h_u_arrmul32_fa19_2_y2, h_u_arrmul32_fa19_2_y4);
  and_gate and_gate_h_u_arrmul32_and20_2_y0(a_20, b_2, h_u_arrmul32_and20_2_y0);
  fa fa_h_u_arrmul32_fa20_2_y2(h_u_arrmul32_and20_2_y0, h_u_arrmul32_fa21_1_y2, h_u_arrmul32_fa19_2_y4, h_u_arrmul32_fa20_2_y2, h_u_arrmul32_fa20_2_y4);
  and_gate and_gate_h_u_arrmul32_and21_2_y0(a_21, b_2, h_u_arrmul32_and21_2_y0);
  fa fa_h_u_arrmul32_fa21_2_y2(h_u_arrmul32_and21_2_y0, h_u_arrmul32_fa22_1_y2, h_u_arrmul32_fa20_2_y4, h_u_arrmul32_fa21_2_y2, h_u_arrmul32_fa21_2_y4);
  and_gate and_gate_h_u_arrmul32_and22_2_y0(a_22, b_2, h_u_arrmul32_and22_2_y0);
  fa fa_h_u_arrmul32_fa22_2_y2(h_u_arrmul32_and22_2_y0, h_u_arrmul32_fa23_1_y2, h_u_arrmul32_fa21_2_y4, h_u_arrmul32_fa22_2_y2, h_u_arrmul32_fa22_2_y4);
  and_gate and_gate_h_u_arrmul32_and23_2_y0(a_23, b_2, h_u_arrmul32_and23_2_y0);
  fa fa_h_u_arrmul32_fa23_2_y2(h_u_arrmul32_and23_2_y0, h_u_arrmul32_fa24_1_y2, h_u_arrmul32_fa22_2_y4, h_u_arrmul32_fa23_2_y2, h_u_arrmul32_fa23_2_y4);
  and_gate and_gate_h_u_arrmul32_and24_2_y0(a_24, b_2, h_u_arrmul32_and24_2_y0);
  fa fa_h_u_arrmul32_fa24_2_y2(h_u_arrmul32_and24_2_y0, h_u_arrmul32_fa25_1_y2, h_u_arrmul32_fa23_2_y4, h_u_arrmul32_fa24_2_y2, h_u_arrmul32_fa24_2_y4);
  and_gate and_gate_h_u_arrmul32_and25_2_y0(a_25, b_2, h_u_arrmul32_and25_2_y0);
  fa fa_h_u_arrmul32_fa25_2_y2(h_u_arrmul32_and25_2_y0, h_u_arrmul32_fa26_1_y2, h_u_arrmul32_fa24_2_y4, h_u_arrmul32_fa25_2_y2, h_u_arrmul32_fa25_2_y4);
  and_gate and_gate_h_u_arrmul32_and26_2_y0(a_26, b_2, h_u_arrmul32_and26_2_y0);
  fa fa_h_u_arrmul32_fa26_2_y2(h_u_arrmul32_and26_2_y0, h_u_arrmul32_fa27_1_y2, h_u_arrmul32_fa25_2_y4, h_u_arrmul32_fa26_2_y2, h_u_arrmul32_fa26_2_y4);
  and_gate and_gate_h_u_arrmul32_and27_2_y0(a_27, b_2, h_u_arrmul32_and27_2_y0);
  fa fa_h_u_arrmul32_fa27_2_y2(h_u_arrmul32_and27_2_y0, h_u_arrmul32_fa28_1_y2, h_u_arrmul32_fa26_2_y4, h_u_arrmul32_fa27_2_y2, h_u_arrmul32_fa27_2_y4);
  and_gate and_gate_h_u_arrmul32_and28_2_y0(a_28, b_2, h_u_arrmul32_and28_2_y0);
  fa fa_h_u_arrmul32_fa28_2_y2(h_u_arrmul32_and28_2_y0, h_u_arrmul32_fa29_1_y2, h_u_arrmul32_fa27_2_y4, h_u_arrmul32_fa28_2_y2, h_u_arrmul32_fa28_2_y4);
  and_gate and_gate_h_u_arrmul32_and29_2_y0(a_29, b_2, h_u_arrmul32_and29_2_y0);
  fa fa_h_u_arrmul32_fa29_2_y2(h_u_arrmul32_and29_2_y0, h_u_arrmul32_fa30_1_y2, h_u_arrmul32_fa28_2_y4, h_u_arrmul32_fa29_2_y2, h_u_arrmul32_fa29_2_y4);
  and_gate and_gate_h_u_arrmul32_and30_2_y0(a_30, b_2, h_u_arrmul32_and30_2_y0);
  fa fa_h_u_arrmul32_fa30_2_y2(h_u_arrmul32_and30_2_y0, h_u_arrmul32_ha31_1_y0, h_u_arrmul32_fa29_2_y4, h_u_arrmul32_fa30_2_y2, h_u_arrmul32_fa30_2_y4);
  and_gate and_gate_h_u_arrmul32_and31_2_y0(a_31, b_2, h_u_arrmul32_and31_2_y0);
  fa fa_h_u_arrmul32_fa31_2_y2(h_u_arrmul32_and31_2_y0, h_u_arrmul32_ha31_1_y1, h_u_arrmul32_fa30_2_y4, h_u_arrmul32_fa31_2_y2, h_u_arrmul32_fa31_2_y4);
  and_gate and_gate_h_u_arrmul32_and0_3_y0(a_0, b_3, h_u_arrmul32_and0_3_y0);
  ha ha_h_u_arrmul32_ha0_3_y0(h_u_arrmul32_and0_3_y0, h_u_arrmul32_fa1_2_y2, h_u_arrmul32_ha0_3_y0, h_u_arrmul32_ha0_3_y1);
  and_gate and_gate_h_u_arrmul32_and1_3_y0(a_1, b_3, h_u_arrmul32_and1_3_y0);
  fa fa_h_u_arrmul32_fa1_3_y2(h_u_arrmul32_and1_3_y0, h_u_arrmul32_fa2_2_y2, h_u_arrmul32_ha0_3_y1, h_u_arrmul32_fa1_3_y2, h_u_arrmul32_fa1_3_y4);
  and_gate and_gate_h_u_arrmul32_and2_3_y0(a_2, b_3, h_u_arrmul32_and2_3_y0);
  fa fa_h_u_arrmul32_fa2_3_y2(h_u_arrmul32_and2_3_y0, h_u_arrmul32_fa3_2_y2, h_u_arrmul32_fa1_3_y4, h_u_arrmul32_fa2_3_y2, h_u_arrmul32_fa2_3_y4);
  and_gate and_gate_h_u_arrmul32_and3_3_y0(a_3, b_3, h_u_arrmul32_and3_3_y0);
  fa fa_h_u_arrmul32_fa3_3_y2(h_u_arrmul32_and3_3_y0, h_u_arrmul32_fa4_2_y2, h_u_arrmul32_fa2_3_y4, h_u_arrmul32_fa3_3_y2, h_u_arrmul32_fa3_3_y4);
  and_gate and_gate_h_u_arrmul32_and4_3_y0(a_4, b_3, h_u_arrmul32_and4_3_y0);
  fa fa_h_u_arrmul32_fa4_3_y2(h_u_arrmul32_and4_3_y0, h_u_arrmul32_fa5_2_y2, h_u_arrmul32_fa3_3_y4, h_u_arrmul32_fa4_3_y2, h_u_arrmul32_fa4_3_y4);
  and_gate and_gate_h_u_arrmul32_and5_3_y0(a_5, b_3, h_u_arrmul32_and5_3_y0);
  fa fa_h_u_arrmul32_fa5_3_y2(h_u_arrmul32_and5_3_y0, h_u_arrmul32_fa6_2_y2, h_u_arrmul32_fa4_3_y4, h_u_arrmul32_fa5_3_y2, h_u_arrmul32_fa5_3_y4);
  and_gate and_gate_h_u_arrmul32_and6_3_y0(a_6, b_3, h_u_arrmul32_and6_3_y0);
  fa fa_h_u_arrmul32_fa6_3_y2(h_u_arrmul32_and6_3_y0, h_u_arrmul32_fa7_2_y2, h_u_arrmul32_fa5_3_y4, h_u_arrmul32_fa6_3_y2, h_u_arrmul32_fa6_3_y4);
  and_gate and_gate_h_u_arrmul32_and7_3_y0(a_7, b_3, h_u_arrmul32_and7_3_y0);
  fa fa_h_u_arrmul32_fa7_3_y2(h_u_arrmul32_and7_3_y0, h_u_arrmul32_fa8_2_y2, h_u_arrmul32_fa6_3_y4, h_u_arrmul32_fa7_3_y2, h_u_arrmul32_fa7_3_y4);
  and_gate and_gate_h_u_arrmul32_and8_3_y0(a_8, b_3, h_u_arrmul32_and8_3_y0);
  fa fa_h_u_arrmul32_fa8_3_y2(h_u_arrmul32_and8_3_y0, h_u_arrmul32_fa9_2_y2, h_u_arrmul32_fa7_3_y4, h_u_arrmul32_fa8_3_y2, h_u_arrmul32_fa8_3_y4);
  and_gate and_gate_h_u_arrmul32_and9_3_y0(a_9, b_3, h_u_arrmul32_and9_3_y0);
  fa fa_h_u_arrmul32_fa9_3_y2(h_u_arrmul32_and9_3_y0, h_u_arrmul32_fa10_2_y2, h_u_arrmul32_fa8_3_y4, h_u_arrmul32_fa9_3_y2, h_u_arrmul32_fa9_3_y4);
  and_gate and_gate_h_u_arrmul32_and10_3_y0(a_10, b_3, h_u_arrmul32_and10_3_y0);
  fa fa_h_u_arrmul32_fa10_3_y2(h_u_arrmul32_and10_3_y0, h_u_arrmul32_fa11_2_y2, h_u_arrmul32_fa9_3_y4, h_u_arrmul32_fa10_3_y2, h_u_arrmul32_fa10_3_y4);
  and_gate and_gate_h_u_arrmul32_and11_3_y0(a_11, b_3, h_u_arrmul32_and11_3_y0);
  fa fa_h_u_arrmul32_fa11_3_y2(h_u_arrmul32_and11_3_y0, h_u_arrmul32_fa12_2_y2, h_u_arrmul32_fa10_3_y4, h_u_arrmul32_fa11_3_y2, h_u_arrmul32_fa11_3_y4);
  and_gate and_gate_h_u_arrmul32_and12_3_y0(a_12, b_3, h_u_arrmul32_and12_3_y0);
  fa fa_h_u_arrmul32_fa12_3_y2(h_u_arrmul32_and12_3_y0, h_u_arrmul32_fa13_2_y2, h_u_arrmul32_fa11_3_y4, h_u_arrmul32_fa12_3_y2, h_u_arrmul32_fa12_3_y4);
  and_gate and_gate_h_u_arrmul32_and13_3_y0(a_13, b_3, h_u_arrmul32_and13_3_y0);
  fa fa_h_u_arrmul32_fa13_3_y2(h_u_arrmul32_and13_3_y0, h_u_arrmul32_fa14_2_y2, h_u_arrmul32_fa12_3_y4, h_u_arrmul32_fa13_3_y2, h_u_arrmul32_fa13_3_y4);
  and_gate and_gate_h_u_arrmul32_and14_3_y0(a_14, b_3, h_u_arrmul32_and14_3_y0);
  fa fa_h_u_arrmul32_fa14_3_y2(h_u_arrmul32_and14_3_y0, h_u_arrmul32_fa15_2_y2, h_u_arrmul32_fa13_3_y4, h_u_arrmul32_fa14_3_y2, h_u_arrmul32_fa14_3_y4);
  and_gate and_gate_h_u_arrmul32_and15_3_y0(a_15, b_3, h_u_arrmul32_and15_3_y0);
  fa fa_h_u_arrmul32_fa15_3_y2(h_u_arrmul32_and15_3_y0, h_u_arrmul32_fa16_2_y2, h_u_arrmul32_fa14_3_y4, h_u_arrmul32_fa15_3_y2, h_u_arrmul32_fa15_3_y4);
  and_gate and_gate_h_u_arrmul32_and16_3_y0(a_16, b_3, h_u_arrmul32_and16_3_y0);
  fa fa_h_u_arrmul32_fa16_3_y2(h_u_arrmul32_and16_3_y0, h_u_arrmul32_fa17_2_y2, h_u_arrmul32_fa15_3_y4, h_u_arrmul32_fa16_3_y2, h_u_arrmul32_fa16_3_y4);
  and_gate and_gate_h_u_arrmul32_and17_3_y0(a_17, b_3, h_u_arrmul32_and17_3_y0);
  fa fa_h_u_arrmul32_fa17_3_y2(h_u_arrmul32_and17_3_y0, h_u_arrmul32_fa18_2_y2, h_u_arrmul32_fa16_3_y4, h_u_arrmul32_fa17_3_y2, h_u_arrmul32_fa17_3_y4);
  and_gate and_gate_h_u_arrmul32_and18_3_y0(a_18, b_3, h_u_arrmul32_and18_3_y0);
  fa fa_h_u_arrmul32_fa18_3_y2(h_u_arrmul32_and18_3_y0, h_u_arrmul32_fa19_2_y2, h_u_arrmul32_fa17_3_y4, h_u_arrmul32_fa18_3_y2, h_u_arrmul32_fa18_3_y4);
  and_gate and_gate_h_u_arrmul32_and19_3_y0(a_19, b_3, h_u_arrmul32_and19_3_y0);
  fa fa_h_u_arrmul32_fa19_3_y2(h_u_arrmul32_and19_3_y0, h_u_arrmul32_fa20_2_y2, h_u_arrmul32_fa18_3_y4, h_u_arrmul32_fa19_3_y2, h_u_arrmul32_fa19_3_y4);
  and_gate and_gate_h_u_arrmul32_and20_3_y0(a_20, b_3, h_u_arrmul32_and20_3_y0);
  fa fa_h_u_arrmul32_fa20_3_y2(h_u_arrmul32_and20_3_y0, h_u_arrmul32_fa21_2_y2, h_u_arrmul32_fa19_3_y4, h_u_arrmul32_fa20_3_y2, h_u_arrmul32_fa20_3_y4);
  and_gate and_gate_h_u_arrmul32_and21_3_y0(a_21, b_3, h_u_arrmul32_and21_3_y0);
  fa fa_h_u_arrmul32_fa21_3_y2(h_u_arrmul32_and21_3_y0, h_u_arrmul32_fa22_2_y2, h_u_arrmul32_fa20_3_y4, h_u_arrmul32_fa21_3_y2, h_u_arrmul32_fa21_3_y4);
  and_gate and_gate_h_u_arrmul32_and22_3_y0(a_22, b_3, h_u_arrmul32_and22_3_y0);
  fa fa_h_u_arrmul32_fa22_3_y2(h_u_arrmul32_and22_3_y0, h_u_arrmul32_fa23_2_y2, h_u_arrmul32_fa21_3_y4, h_u_arrmul32_fa22_3_y2, h_u_arrmul32_fa22_3_y4);
  and_gate and_gate_h_u_arrmul32_and23_3_y0(a_23, b_3, h_u_arrmul32_and23_3_y0);
  fa fa_h_u_arrmul32_fa23_3_y2(h_u_arrmul32_and23_3_y0, h_u_arrmul32_fa24_2_y2, h_u_arrmul32_fa22_3_y4, h_u_arrmul32_fa23_3_y2, h_u_arrmul32_fa23_3_y4);
  and_gate and_gate_h_u_arrmul32_and24_3_y0(a_24, b_3, h_u_arrmul32_and24_3_y0);
  fa fa_h_u_arrmul32_fa24_3_y2(h_u_arrmul32_and24_3_y0, h_u_arrmul32_fa25_2_y2, h_u_arrmul32_fa23_3_y4, h_u_arrmul32_fa24_3_y2, h_u_arrmul32_fa24_3_y4);
  and_gate and_gate_h_u_arrmul32_and25_3_y0(a_25, b_3, h_u_arrmul32_and25_3_y0);
  fa fa_h_u_arrmul32_fa25_3_y2(h_u_arrmul32_and25_3_y0, h_u_arrmul32_fa26_2_y2, h_u_arrmul32_fa24_3_y4, h_u_arrmul32_fa25_3_y2, h_u_arrmul32_fa25_3_y4);
  and_gate and_gate_h_u_arrmul32_and26_3_y0(a_26, b_3, h_u_arrmul32_and26_3_y0);
  fa fa_h_u_arrmul32_fa26_3_y2(h_u_arrmul32_and26_3_y0, h_u_arrmul32_fa27_2_y2, h_u_arrmul32_fa25_3_y4, h_u_arrmul32_fa26_3_y2, h_u_arrmul32_fa26_3_y4);
  and_gate and_gate_h_u_arrmul32_and27_3_y0(a_27, b_3, h_u_arrmul32_and27_3_y0);
  fa fa_h_u_arrmul32_fa27_3_y2(h_u_arrmul32_and27_3_y0, h_u_arrmul32_fa28_2_y2, h_u_arrmul32_fa26_3_y4, h_u_arrmul32_fa27_3_y2, h_u_arrmul32_fa27_3_y4);
  and_gate and_gate_h_u_arrmul32_and28_3_y0(a_28, b_3, h_u_arrmul32_and28_3_y0);
  fa fa_h_u_arrmul32_fa28_3_y2(h_u_arrmul32_and28_3_y0, h_u_arrmul32_fa29_2_y2, h_u_arrmul32_fa27_3_y4, h_u_arrmul32_fa28_3_y2, h_u_arrmul32_fa28_3_y4);
  and_gate and_gate_h_u_arrmul32_and29_3_y0(a_29, b_3, h_u_arrmul32_and29_3_y0);
  fa fa_h_u_arrmul32_fa29_3_y2(h_u_arrmul32_and29_3_y0, h_u_arrmul32_fa30_2_y2, h_u_arrmul32_fa28_3_y4, h_u_arrmul32_fa29_3_y2, h_u_arrmul32_fa29_3_y4);
  and_gate and_gate_h_u_arrmul32_and30_3_y0(a_30, b_3, h_u_arrmul32_and30_3_y0);
  fa fa_h_u_arrmul32_fa30_3_y2(h_u_arrmul32_and30_3_y0, h_u_arrmul32_fa31_2_y2, h_u_arrmul32_fa29_3_y4, h_u_arrmul32_fa30_3_y2, h_u_arrmul32_fa30_3_y4);
  and_gate and_gate_h_u_arrmul32_and31_3_y0(a_31, b_3, h_u_arrmul32_and31_3_y0);
  fa fa_h_u_arrmul32_fa31_3_y2(h_u_arrmul32_and31_3_y0, h_u_arrmul32_fa31_2_y4, h_u_arrmul32_fa30_3_y4, h_u_arrmul32_fa31_3_y2, h_u_arrmul32_fa31_3_y4);
  and_gate and_gate_h_u_arrmul32_and0_4_y0(a_0, b_4, h_u_arrmul32_and0_4_y0);
  ha ha_h_u_arrmul32_ha0_4_y0(h_u_arrmul32_and0_4_y0, h_u_arrmul32_fa1_3_y2, h_u_arrmul32_ha0_4_y0, h_u_arrmul32_ha0_4_y1);
  and_gate and_gate_h_u_arrmul32_and1_4_y0(a_1, b_4, h_u_arrmul32_and1_4_y0);
  fa fa_h_u_arrmul32_fa1_4_y2(h_u_arrmul32_and1_4_y0, h_u_arrmul32_fa2_3_y2, h_u_arrmul32_ha0_4_y1, h_u_arrmul32_fa1_4_y2, h_u_arrmul32_fa1_4_y4);
  and_gate and_gate_h_u_arrmul32_and2_4_y0(a_2, b_4, h_u_arrmul32_and2_4_y0);
  fa fa_h_u_arrmul32_fa2_4_y2(h_u_arrmul32_and2_4_y0, h_u_arrmul32_fa3_3_y2, h_u_arrmul32_fa1_4_y4, h_u_arrmul32_fa2_4_y2, h_u_arrmul32_fa2_4_y4);
  and_gate and_gate_h_u_arrmul32_and3_4_y0(a_3, b_4, h_u_arrmul32_and3_4_y0);
  fa fa_h_u_arrmul32_fa3_4_y2(h_u_arrmul32_and3_4_y0, h_u_arrmul32_fa4_3_y2, h_u_arrmul32_fa2_4_y4, h_u_arrmul32_fa3_4_y2, h_u_arrmul32_fa3_4_y4);
  and_gate and_gate_h_u_arrmul32_and4_4_y0(a_4, b_4, h_u_arrmul32_and4_4_y0);
  fa fa_h_u_arrmul32_fa4_4_y2(h_u_arrmul32_and4_4_y0, h_u_arrmul32_fa5_3_y2, h_u_arrmul32_fa3_4_y4, h_u_arrmul32_fa4_4_y2, h_u_arrmul32_fa4_4_y4);
  and_gate and_gate_h_u_arrmul32_and5_4_y0(a_5, b_4, h_u_arrmul32_and5_4_y0);
  fa fa_h_u_arrmul32_fa5_4_y2(h_u_arrmul32_and5_4_y0, h_u_arrmul32_fa6_3_y2, h_u_arrmul32_fa4_4_y4, h_u_arrmul32_fa5_4_y2, h_u_arrmul32_fa5_4_y4);
  and_gate and_gate_h_u_arrmul32_and6_4_y0(a_6, b_4, h_u_arrmul32_and6_4_y0);
  fa fa_h_u_arrmul32_fa6_4_y2(h_u_arrmul32_and6_4_y0, h_u_arrmul32_fa7_3_y2, h_u_arrmul32_fa5_4_y4, h_u_arrmul32_fa6_4_y2, h_u_arrmul32_fa6_4_y4);
  and_gate and_gate_h_u_arrmul32_and7_4_y0(a_7, b_4, h_u_arrmul32_and7_4_y0);
  fa fa_h_u_arrmul32_fa7_4_y2(h_u_arrmul32_and7_4_y0, h_u_arrmul32_fa8_3_y2, h_u_arrmul32_fa6_4_y4, h_u_arrmul32_fa7_4_y2, h_u_arrmul32_fa7_4_y4);
  and_gate and_gate_h_u_arrmul32_and8_4_y0(a_8, b_4, h_u_arrmul32_and8_4_y0);
  fa fa_h_u_arrmul32_fa8_4_y2(h_u_arrmul32_and8_4_y0, h_u_arrmul32_fa9_3_y2, h_u_arrmul32_fa7_4_y4, h_u_arrmul32_fa8_4_y2, h_u_arrmul32_fa8_4_y4);
  and_gate and_gate_h_u_arrmul32_and9_4_y0(a_9, b_4, h_u_arrmul32_and9_4_y0);
  fa fa_h_u_arrmul32_fa9_4_y2(h_u_arrmul32_and9_4_y0, h_u_arrmul32_fa10_3_y2, h_u_arrmul32_fa8_4_y4, h_u_arrmul32_fa9_4_y2, h_u_arrmul32_fa9_4_y4);
  and_gate and_gate_h_u_arrmul32_and10_4_y0(a_10, b_4, h_u_arrmul32_and10_4_y0);
  fa fa_h_u_arrmul32_fa10_4_y2(h_u_arrmul32_and10_4_y0, h_u_arrmul32_fa11_3_y2, h_u_arrmul32_fa9_4_y4, h_u_arrmul32_fa10_4_y2, h_u_arrmul32_fa10_4_y4);
  and_gate and_gate_h_u_arrmul32_and11_4_y0(a_11, b_4, h_u_arrmul32_and11_4_y0);
  fa fa_h_u_arrmul32_fa11_4_y2(h_u_arrmul32_and11_4_y0, h_u_arrmul32_fa12_3_y2, h_u_arrmul32_fa10_4_y4, h_u_arrmul32_fa11_4_y2, h_u_arrmul32_fa11_4_y4);
  and_gate and_gate_h_u_arrmul32_and12_4_y0(a_12, b_4, h_u_arrmul32_and12_4_y0);
  fa fa_h_u_arrmul32_fa12_4_y2(h_u_arrmul32_and12_4_y0, h_u_arrmul32_fa13_3_y2, h_u_arrmul32_fa11_4_y4, h_u_arrmul32_fa12_4_y2, h_u_arrmul32_fa12_4_y4);
  and_gate and_gate_h_u_arrmul32_and13_4_y0(a_13, b_4, h_u_arrmul32_and13_4_y0);
  fa fa_h_u_arrmul32_fa13_4_y2(h_u_arrmul32_and13_4_y0, h_u_arrmul32_fa14_3_y2, h_u_arrmul32_fa12_4_y4, h_u_arrmul32_fa13_4_y2, h_u_arrmul32_fa13_4_y4);
  and_gate and_gate_h_u_arrmul32_and14_4_y0(a_14, b_4, h_u_arrmul32_and14_4_y0);
  fa fa_h_u_arrmul32_fa14_4_y2(h_u_arrmul32_and14_4_y0, h_u_arrmul32_fa15_3_y2, h_u_arrmul32_fa13_4_y4, h_u_arrmul32_fa14_4_y2, h_u_arrmul32_fa14_4_y4);
  and_gate and_gate_h_u_arrmul32_and15_4_y0(a_15, b_4, h_u_arrmul32_and15_4_y0);
  fa fa_h_u_arrmul32_fa15_4_y2(h_u_arrmul32_and15_4_y0, h_u_arrmul32_fa16_3_y2, h_u_arrmul32_fa14_4_y4, h_u_arrmul32_fa15_4_y2, h_u_arrmul32_fa15_4_y4);
  and_gate and_gate_h_u_arrmul32_and16_4_y0(a_16, b_4, h_u_arrmul32_and16_4_y0);
  fa fa_h_u_arrmul32_fa16_4_y2(h_u_arrmul32_and16_4_y0, h_u_arrmul32_fa17_3_y2, h_u_arrmul32_fa15_4_y4, h_u_arrmul32_fa16_4_y2, h_u_arrmul32_fa16_4_y4);
  and_gate and_gate_h_u_arrmul32_and17_4_y0(a_17, b_4, h_u_arrmul32_and17_4_y0);
  fa fa_h_u_arrmul32_fa17_4_y2(h_u_arrmul32_and17_4_y0, h_u_arrmul32_fa18_3_y2, h_u_arrmul32_fa16_4_y4, h_u_arrmul32_fa17_4_y2, h_u_arrmul32_fa17_4_y4);
  and_gate and_gate_h_u_arrmul32_and18_4_y0(a_18, b_4, h_u_arrmul32_and18_4_y0);
  fa fa_h_u_arrmul32_fa18_4_y2(h_u_arrmul32_and18_4_y0, h_u_arrmul32_fa19_3_y2, h_u_arrmul32_fa17_4_y4, h_u_arrmul32_fa18_4_y2, h_u_arrmul32_fa18_4_y4);
  and_gate and_gate_h_u_arrmul32_and19_4_y0(a_19, b_4, h_u_arrmul32_and19_4_y0);
  fa fa_h_u_arrmul32_fa19_4_y2(h_u_arrmul32_and19_4_y0, h_u_arrmul32_fa20_3_y2, h_u_arrmul32_fa18_4_y4, h_u_arrmul32_fa19_4_y2, h_u_arrmul32_fa19_4_y4);
  and_gate and_gate_h_u_arrmul32_and20_4_y0(a_20, b_4, h_u_arrmul32_and20_4_y0);
  fa fa_h_u_arrmul32_fa20_4_y2(h_u_arrmul32_and20_4_y0, h_u_arrmul32_fa21_3_y2, h_u_arrmul32_fa19_4_y4, h_u_arrmul32_fa20_4_y2, h_u_arrmul32_fa20_4_y4);
  and_gate and_gate_h_u_arrmul32_and21_4_y0(a_21, b_4, h_u_arrmul32_and21_4_y0);
  fa fa_h_u_arrmul32_fa21_4_y2(h_u_arrmul32_and21_4_y0, h_u_arrmul32_fa22_3_y2, h_u_arrmul32_fa20_4_y4, h_u_arrmul32_fa21_4_y2, h_u_arrmul32_fa21_4_y4);
  and_gate and_gate_h_u_arrmul32_and22_4_y0(a_22, b_4, h_u_arrmul32_and22_4_y0);
  fa fa_h_u_arrmul32_fa22_4_y2(h_u_arrmul32_and22_4_y0, h_u_arrmul32_fa23_3_y2, h_u_arrmul32_fa21_4_y4, h_u_arrmul32_fa22_4_y2, h_u_arrmul32_fa22_4_y4);
  and_gate and_gate_h_u_arrmul32_and23_4_y0(a_23, b_4, h_u_arrmul32_and23_4_y0);
  fa fa_h_u_arrmul32_fa23_4_y2(h_u_arrmul32_and23_4_y0, h_u_arrmul32_fa24_3_y2, h_u_arrmul32_fa22_4_y4, h_u_arrmul32_fa23_4_y2, h_u_arrmul32_fa23_4_y4);
  and_gate and_gate_h_u_arrmul32_and24_4_y0(a_24, b_4, h_u_arrmul32_and24_4_y0);
  fa fa_h_u_arrmul32_fa24_4_y2(h_u_arrmul32_and24_4_y0, h_u_arrmul32_fa25_3_y2, h_u_arrmul32_fa23_4_y4, h_u_arrmul32_fa24_4_y2, h_u_arrmul32_fa24_4_y4);
  and_gate and_gate_h_u_arrmul32_and25_4_y0(a_25, b_4, h_u_arrmul32_and25_4_y0);
  fa fa_h_u_arrmul32_fa25_4_y2(h_u_arrmul32_and25_4_y0, h_u_arrmul32_fa26_3_y2, h_u_arrmul32_fa24_4_y4, h_u_arrmul32_fa25_4_y2, h_u_arrmul32_fa25_4_y4);
  and_gate and_gate_h_u_arrmul32_and26_4_y0(a_26, b_4, h_u_arrmul32_and26_4_y0);
  fa fa_h_u_arrmul32_fa26_4_y2(h_u_arrmul32_and26_4_y0, h_u_arrmul32_fa27_3_y2, h_u_arrmul32_fa25_4_y4, h_u_arrmul32_fa26_4_y2, h_u_arrmul32_fa26_4_y4);
  and_gate and_gate_h_u_arrmul32_and27_4_y0(a_27, b_4, h_u_arrmul32_and27_4_y0);
  fa fa_h_u_arrmul32_fa27_4_y2(h_u_arrmul32_and27_4_y0, h_u_arrmul32_fa28_3_y2, h_u_arrmul32_fa26_4_y4, h_u_arrmul32_fa27_4_y2, h_u_arrmul32_fa27_4_y4);
  and_gate and_gate_h_u_arrmul32_and28_4_y0(a_28, b_4, h_u_arrmul32_and28_4_y0);
  fa fa_h_u_arrmul32_fa28_4_y2(h_u_arrmul32_and28_4_y0, h_u_arrmul32_fa29_3_y2, h_u_arrmul32_fa27_4_y4, h_u_arrmul32_fa28_4_y2, h_u_arrmul32_fa28_4_y4);
  and_gate and_gate_h_u_arrmul32_and29_4_y0(a_29, b_4, h_u_arrmul32_and29_4_y0);
  fa fa_h_u_arrmul32_fa29_4_y2(h_u_arrmul32_and29_4_y0, h_u_arrmul32_fa30_3_y2, h_u_arrmul32_fa28_4_y4, h_u_arrmul32_fa29_4_y2, h_u_arrmul32_fa29_4_y4);
  and_gate and_gate_h_u_arrmul32_and30_4_y0(a_30, b_4, h_u_arrmul32_and30_4_y0);
  fa fa_h_u_arrmul32_fa30_4_y2(h_u_arrmul32_and30_4_y0, h_u_arrmul32_fa31_3_y2, h_u_arrmul32_fa29_4_y4, h_u_arrmul32_fa30_4_y2, h_u_arrmul32_fa30_4_y4);
  and_gate and_gate_h_u_arrmul32_and31_4_y0(a_31, b_4, h_u_arrmul32_and31_4_y0);
  fa fa_h_u_arrmul32_fa31_4_y2(h_u_arrmul32_and31_4_y0, h_u_arrmul32_fa31_3_y4, h_u_arrmul32_fa30_4_y4, h_u_arrmul32_fa31_4_y2, h_u_arrmul32_fa31_4_y4);
  and_gate and_gate_h_u_arrmul32_and0_5_y0(a_0, b_5, h_u_arrmul32_and0_5_y0);
  ha ha_h_u_arrmul32_ha0_5_y0(h_u_arrmul32_and0_5_y0, h_u_arrmul32_fa1_4_y2, h_u_arrmul32_ha0_5_y0, h_u_arrmul32_ha0_5_y1);
  and_gate and_gate_h_u_arrmul32_and1_5_y0(a_1, b_5, h_u_arrmul32_and1_5_y0);
  fa fa_h_u_arrmul32_fa1_5_y2(h_u_arrmul32_and1_5_y0, h_u_arrmul32_fa2_4_y2, h_u_arrmul32_ha0_5_y1, h_u_arrmul32_fa1_5_y2, h_u_arrmul32_fa1_5_y4);
  and_gate and_gate_h_u_arrmul32_and2_5_y0(a_2, b_5, h_u_arrmul32_and2_5_y0);
  fa fa_h_u_arrmul32_fa2_5_y2(h_u_arrmul32_and2_5_y0, h_u_arrmul32_fa3_4_y2, h_u_arrmul32_fa1_5_y4, h_u_arrmul32_fa2_5_y2, h_u_arrmul32_fa2_5_y4);
  and_gate and_gate_h_u_arrmul32_and3_5_y0(a_3, b_5, h_u_arrmul32_and3_5_y0);
  fa fa_h_u_arrmul32_fa3_5_y2(h_u_arrmul32_and3_5_y0, h_u_arrmul32_fa4_4_y2, h_u_arrmul32_fa2_5_y4, h_u_arrmul32_fa3_5_y2, h_u_arrmul32_fa3_5_y4);
  and_gate and_gate_h_u_arrmul32_and4_5_y0(a_4, b_5, h_u_arrmul32_and4_5_y0);
  fa fa_h_u_arrmul32_fa4_5_y2(h_u_arrmul32_and4_5_y0, h_u_arrmul32_fa5_4_y2, h_u_arrmul32_fa3_5_y4, h_u_arrmul32_fa4_5_y2, h_u_arrmul32_fa4_5_y4);
  and_gate and_gate_h_u_arrmul32_and5_5_y0(a_5, b_5, h_u_arrmul32_and5_5_y0);
  fa fa_h_u_arrmul32_fa5_5_y2(h_u_arrmul32_and5_5_y0, h_u_arrmul32_fa6_4_y2, h_u_arrmul32_fa4_5_y4, h_u_arrmul32_fa5_5_y2, h_u_arrmul32_fa5_5_y4);
  and_gate and_gate_h_u_arrmul32_and6_5_y0(a_6, b_5, h_u_arrmul32_and6_5_y0);
  fa fa_h_u_arrmul32_fa6_5_y2(h_u_arrmul32_and6_5_y0, h_u_arrmul32_fa7_4_y2, h_u_arrmul32_fa5_5_y4, h_u_arrmul32_fa6_5_y2, h_u_arrmul32_fa6_5_y4);
  and_gate and_gate_h_u_arrmul32_and7_5_y0(a_7, b_5, h_u_arrmul32_and7_5_y0);
  fa fa_h_u_arrmul32_fa7_5_y2(h_u_arrmul32_and7_5_y0, h_u_arrmul32_fa8_4_y2, h_u_arrmul32_fa6_5_y4, h_u_arrmul32_fa7_5_y2, h_u_arrmul32_fa7_5_y4);
  and_gate and_gate_h_u_arrmul32_and8_5_y0(a_8, b_5, h_u_arrmul32_and8_5_y0);
  fa fa_h_u_arrmul32_fa8_5_y2(h_u_arrmul32_and8_5_y0, h_u_arrmul32_fa9_4_y2, h_u_arrmul32_fa7_5_y4, h_u_arrmul32_fa8_5_y2, h_u_arrmul32_fa8_5_y4);
  and_gate and_gate_h_u_arrmul32_and9_5_y0(a_9, b_5, h_u_arrmul32_and9_5_y0);
  fa fa_h_u_arrmul32_fa9_5_y2(h_u_arrmul32_and9_5_y0, h_u_arrmul32_fa10_4_y2, h_u_arrmul32_fa8_5_y4, h_u_arrmul32_fa9_5_y2, h_u_arrmul32_fa9_5_y4);
  and_gate and_gate_h_u_arrmul32_and10_5_y0(a_10, b_5, h_u_arrmul32_and10_5_y0);
  fa fa_h_u_arrmul32_fa10_5_y2(h_u_arrmul32_and10_5_y0, h_u_arrmul32_fa11_4_y2, h_u_arrmul32_fa9_5_y4, h_u_arrmul32_fa10_5_y2, h_u_arrmul32_fa10_5_y4);
  and_gate and_gate_h_u_arrmul32_and11_5_y0(a_11, b_5, h_u_arrmul32_and11_5_y0);
  fa fa_h_u_arrmul32_fa11_5_y2(h_u_arrmul32_and11_5_y0, h_u_arrmul32_fa12_4_y2, h_u_arrmul32_fa10_5_y4, h_u_arrmul32_fa11_5_y2, h_u_arrmul32_fa11_5_y4);
  and_gate and_gate_h_u_arrmul32_and12_5_y0(a_12, b_5, h_u_arrmul32_and12_5_y0);
  fa fa_h_u_arrmul32_fa12_5_y2(h_u_arrmul32_and12_5_y0, h_u_arrmul32_fa13_4_y2, h_u_arrmul32_fa11_5_y4, h_u_arrmul32_fa12_5_y2, h_u_arrmul32_fa12_5_y4);
  and_gate and_gate_h_u_arrmul32_and13_5_y0(a_13, b_5, h_u_arrmul32_and13_5_y0);
  fa fa_h_u_arrmul32_fa13_5_y2(h_u_arrmul32_and13_5_y0, h_u_arrmul32_fa14_4_y2, h_u_arrmul32_fa12_5_y4, h_u_arrmul32_fa13_5_y2, h_u_arrmul32_fa13_5_y4);
  and_gate and_gate_h_u_arrmul32_and14_5_y0(a_14, b_5, h_u_arrmul32_and14_5_y0);
  fa fa_h_u_arrmul32_fa14_5_y2(h_u_arrmul32_and14_5_y0, h_u_arrmul32_fa15_4_y2, h_u_arrmul32_fa13_5_y4, h_u_arrmul32_fa14_5_y2, h_u_arrmul32_fa14_5_y4);
  and_gate and_gate_h_u_arrmul32_and15_5_y0(a_15, b_5, h_u_arrmul32_and15_5_y0);
  fa fa_h_u_arrmul32_fa15_5_y2(h_u_arrmul32_and15_5_y0, h_u_arrmul32_fa16_4_y2, h_u_arrmul32_fa14_5_y4, h_u_arrmul32_fa15_5_y2, h_u_arrmul32_fa15_5_y4);
  and_gate and_gate_h_u_arrmul32_and16_5_y0(a_16, b_5, h_u_arrmul32_and16_5_y0);
  fa fa_h_u_arrmul32_fa16_5_y2(h_u_arrmul32_and16_5_y0, h_u_arrmul32_fa17_4_y2, h_u_arrmul32_fa15_5_y4, h_u_arrmul32_fa16_5_y2, h_u_arrmul32_fa16_5_y4);
  and_gate and_gate_h_u_arrmul32_and17_5_y0(a_17, b_5, h_u_arrmul32_and17_5_y0);
  fa fa_h_u_arrmul32_fa17_5_y2(h_u_arrmul32_and17_5_y0, h_u_arrmul32_fa18_4_y2, h_u_arrmul32_fa16_5_y4, h_u_arrmul32_fa17_5_y2, h_u_arrmul32_fa17_5_y4);
  and_gate and_gate_h_u_arrmul32_and18_5_y0(a_18, b_5, h_u_arrmul32_and18_5_y0);
  fa fa_h_u_arrmul32_fa18_5_y2(h_u_arrmul32_and18_5_y0, h_u_arrmul32_fa19_4_y2, h_u_arrmul32_fa17_5_y4, h_u_arrmul32_fa18_5_y2, h_u_arrmul32_fa18_5_y4);
  and_gate and_gate_h_u_arrmul32_and19_5_y0(a_19, b_5, h_u_arrmul32_and19_5_y0);
  fa fa_h_u_arrmul32_fa19_5_y2(h_u_arrmul32_and19_5_y0, h_u_arrmul32_fa20_4_y2, h_u_arrmul32_fa18_5_y4, h_u_arrmul32_fa19_5_y2, h_u_arrmul32_fa19_5_y4);
  and_gate and_gate_h_u_arrmul32_and20_5_y0(a_20, b_5, h_u_arrmul32_and20_5_y0);
  fa fa_h_u_arrmul32_fa20_5_y2(h_u_arrmul32_and20_5_y0, h_u_arrmul32_fa21_4_y2, h_u_arrmul32_fa19_5_y4, h_u_arrmul32_fa20_5_y2, h_u_arrmul32_fa20_5_y4);
  and_gate and_gate_h_u_arrmul32_and21_5_y0(a_21, b_5, h_u_arrmul32_and21_5_y0);
  fa fa_h_u_arrmul32_fa21_5_y2(h_u_arrmul32_and21_5_y0, h_u_arrmul32_fa22_4_y2, h_u_arrmul32_fa20_5_y4, h_u_arrmul32_fa21_5_y2, h_u_arrmul32_fa21_5_y4);
  and_gate and_gate_h_u_arrmul32_and22_5_y0(a_22, b_5, h_u_arrmul32_and22_5_y0);
  fa fa_h_u_arrmul32_fa22_5_y2(h_u_arrmul32_and22_5_y0, h_u_arrmul32_fa23_4_y2, h_u_arrmul32_fa21_5_y4, h_u_arrmul32_fa22_5_y2, h_u_arrmul32_fa22_5_y4);
  and_gate and_gate_h_u_arrmul32_and23_5_y0(a_23, b_5, h_u_arrmul32_and23_5_y0);
  fa fa_h_u_arrmul32_fa23_5_y2(h_u_arrmul32_and23_5_y0, h_u_arrmul32_fa24_4_y2, h_u_arrmul32_fa22_5_y4, h_u_arrmul32_fa23_5_y2, h_u_arrmul32_fa23_5_y4);
  and_gate and_gate_h_u_arrmul32_and24_5_y0(a_24, b_5, h_u_arrmul32_and24_5_y0);
  fa fa_h_u_arrmul32_fa24_5_y2(h_u_arrmul32_and24_5_y0, h_u_arrmul32_fa25_4_y2, h_u_arrmul32_fa23_5_y4, h_u_arrmul32_fa24_5_y2, h_u_arrmul32_fa24_5_y4);
  and_gate and_gate_h_u_arrmul32_and25_5_y0(a_25, b_5, h_u_arrmul32_and25_5_y0);
  fa fa_h_u_arrmul32_fa25_5_y2(h_u_arrmul32_and25_5_y0, h_u_arrmul32_fa26_4_y2, h_u_arrmul32_fa24_5_y4, h_u_arrmul32_fa25_5_y2, h_u_arrmul32_fa25_5_y4);
  and_gate and_gate_h_u_arrmul32_and26_5_y0(a_26, b_5, h_u_arrmul32_and26_5_y0);
  fa fa_h_u_arrmul32_fa26_5_y2(h_u_arrmul32_and26_5_y0, h_u_arrmul32_fa27_4_y2, h_u_arrmul32_fa25_5_y4, h_u_arrmul32_fa26_5_y2, h_u_arrmul32_fa26_5_y4);
  and_gate and_gate_h_u_arrmul32_and27_5_y0(a_27, b_5, h_u_arrmul32_and27_5_y0);
  fa fa_h_u_arrmul32_fa27_5_y2(h_u_arrmul32_and27_5_y0, h_u_arrmul32_fa28_4_y2, h_u_arrmul32_fa26_5_y4, h_u_arrmul32_fa27_5_y2, h_u_arrmul32_fa27_5_y4);
  and_gate and_gate_h_u_arrmul32_and28_5_y0(a_28, b_5, h_u_arrmul32_and28_5_y0);
  fa fa_h_u_arrmul32_fa28_5_y2(h_u_arrmul32_and28_5_y0, h_u_arrmul32_fa29_4_y2, h_u_arrmul32_fa27_5_y4, h_u_arrmul32_fa28_5_y2, h_u_arrmul32_fa28_5_y4);
  and_gate and_gate_h_u_arrmul32_and29_5_y0(a_29, b_5, h_u_arrmul32_and29_5_y0);
  fa fa_h_u_arrmul32_fa29_5_y2(h_u_arrmul32_and29_5_y0, h_u_arrmul32_fa30_4_y2, h_u_arrmul32_fa28_5_y4, h_u_arrmul32_fa29_5_y2, h_u_arrmul32_fa29_5_y4);
  and_gate and_gate_h_u_arrmul32_and30_5_y0(a_30, b_5, h_u_arrmul32_and30_5_y0);
  fa fa_h_u_arrmul32_fa30_5_y2(h_u_arrmul32_and30_5_y0, h_u_arrmul32_fa31_4_y2, h_u_arrmul32_fa29_5_y4, h_u_arrmul32_fa30_5_y2, h_u_arrmul32_fa30_5_y4);
  and_gate and_gate_h_u_arrmul32_and31_5_y0(a_31, b_5, h_u_arrmul32_and31_5_y0);
  fa fa_h_u_arrmul32_fa31_5_y2(h_u_arrmul32_and31_5_y0, h_u_arrmul32_fa31_4_y4, h_u_arrmul32_fa30_5_y4, h_u_arrmul32_fa31_5_y2, h_u_arrmul32_fa31_5_y4);
  and_gate and_gate_h_u_arrmul32_and0_6_y0(a_0, b_6, h_u_arrmul32_and0_6_y0);
  ha ha_h_u_arrmul32_ha0_6_y0(h_u_arrmul32_and0_6_y0, h_u_arrmul32_fa1_5_y2, h_u_arrmul32_ha0_6_y0, h_u_arrmul32_ha0_6_y1);
  and_gate and_gate_h_u_arrmul32_and1_6_y0(a_1, b_6, h_u_arrmul32_and1_6_y0);
  fa fa_h_u_arrmul32_fa1_6_y2(h_u_arrmul32_and1_6_y0, h_u_arrmul32_fa2_5_y2, h_u_arrmul32_ha0_6_y1, h_u_arrmul32_fa1_6_y2, h_u_arrmul32_fa1_6_y4);
  and_gate and_gate_h_u_arrmul32_and2_6_y0(a_2, b_6, h_u_arrmul32_and2_6_y0);
  fa fa_h_u_arrmul32_fa2_6_y2(h_u_arrmul32_and2_6_y0, h_u_arrmul32_fa3_5_y2, h_u_arrmul32_fa1_6_y4, h_u_arrmul32_fa2_6_y2, h_u_arrmul32_fa2_6_y4);
  and_gate and_gate_h_u_arrmul32_and3_6_y0(a_3, b_6, h_u_arrmul32_and3_6_y0);
  fa fa_h_u_arrmul32_fa3_6_y2(h_u_arrmul32_and3_6_y0, h_u_arrmul32_fa4_5_y2, h_u_arrmul32_fa2_6_y4, h_u_arrmul32_fa3_6_y2, h_u_arrmul32_fa3_6_y4);
  and_gate and_gate_h_u_arrmul32_and4_6_y0(a_4, b_6, h_u_arrmul32_and4_6_y0);
  fa fa_h_u_arrmul32_fa4_6_y2(h_u_arrmul32_and4_6_y0, h_u_arrmul32_fa5_5_y2, h_u_arrmul32_fa3_6_y4, h_u_arrmul32_fa4_6_y2, h_u_arrmul32_fa4_6_y4);
  and_gate and_gate_h_u_arrmul32_and5_6_y0(a_5, b_6, h_u_arrmul32_and5_6_y0);
  fa fa_h_u_arrmul32_fa5_6_y2(h_u_arrmul32_and5_6_y0, h_u_arrmul32_fa6_5_y2, h_u_arrmul32_fa4_6_y4, h_u_arrmul32_fa5_6_y2, h_u_arrmul32_fa5_6_y4);
  and_gate and_gate_h_u_arrmul32_and6_6_y0(a_6, b_6, h_u_arrmul32_and6_6_y0);
  fa fa_h_u_arrmul32_fa6_6_y2(h_u_arrmul32_and6_6_y0, h_u_arrmul32_fa7_5_y2, h_u_arrmul32_fa5_6_y4, h_u_arrmul32_fa6_6_y2, h_u_arrmul32_fa6_6_y4);
  and_gate and_gate_h_u_arrmul32_and7_6_y0(a_7, b_6, h_u_arrmul32_and7_6_y0);
  fa fa_h_u_arrmul32_fa7_6_y2(h_u_arrmul32_and7_6_y0, h_u_arrmul32_fa8_5_y2, h_u_arrmul32_fa6_6_y4, h_u_arrmul32_fa7_6_y2, h_u_arrmul32_fa7_6_y4);
  and_gate and_gate_h_u_arrmul32_and8_6_y0(a_8, b_6, h_u_arrmul32_and8_6_y0);
  fa fa_h_u_arrmul32_fa8_6_y2(h_u_arrmul32_and8_6_y0, h_u_arrmul32_fa9_5_y2, h_u_arrmul32_fa7_6_y4, h_u_arrmul32_fa8_6_y2, h_u_arrmul32_fa8_6_y4);
  and_gate and_gate_h_u_arrmul32_and9_6_y0(a_9, b_6, h_u_arrmul32_and9_6_y0);
  fa fa_h_u_arrmul32_fa9_6_y2(h_u_arrmul32_and9_6_y0, h_u_arrmul32_fa10_5_y2, h_u_arrmul32_fa8_6_y4, h_u_arrmul32_fa9_6_y2, h_u_arrmul32_fa9_6_y4);
  and_gate and_gate_h_u_arrmul32_and10_6_y0(a_10, b_6, h_u_arrmul32_and10_6_y0);
  fa fa_h_u_arrmul32_fa10_6_y2(h_u_arrmul32_and10_6_y0, h_u_arrmul32_fa11_5_y2, h_u_arrmul32_fa9_6_y4, h_u_arrmul32_fa10_6_y2, h_u_arrmul32_fa10_6_y4);
  and_gate and_gate_h_u_arrmul32_and11_6_y0(a_11, b_6, h_u_arrmul32_and11_6_y0);
  fa fa_h_u_arrmul32_fa11_6_y2(h_u_arrmul32_and11_6_y0, h_u_arrmul32_fa12_5_y2, h_u_arrmul32_fa10_6_y4, h_u_arrmul32_fa11_6_y2, h_u_arrmul32_fa11_6_y4);
  and_gate and_gate_h_u_arrmul32_and12_6_y0(a_12, b_6, h_u_arrmul32_and12_6_y0);
  fa fa_h_u_arrmul32_fa12_6_y2(h_u_arrmul32_and12_6_y0, h_u_arrmul32_fa13_5_y2, h_u_arrmul32_fa11_6_y4, h_u_arrmul32_fa12_6_y2, h_u_arrmul32_fa12_6_y4);
  and_gate and_gate_h_u_arrmul32_and13_6_y0(a_13, b_6, h_u_arrmul32_and13_6_y0);
  fa fa_h_u_arrmul32_fa13_6_y2(h_u_arrmul32_and13_6_y0, h_u_arrmul32_fa14_5_y2, h_u_arrmul32_fa12_6_y4, h_u_arrmul32_fa13_6_y2, h_u_arrmul32_fa13_6_y4);
  and_gate and_gate_h_u_arrmul32_and14_6_y0(a_14, b_6, h_u_arrmul32_and14_6_y0);
  fa fa_h_u_arrmul32_fa14_6_y2(h_u_arrmul32_and14_6_y0, h_u_arrmul32_fa15_5_y2, h_u_arrmul32_fa13_6_y4, h_u_arrmul32_fa14_6_y2, h_u_arrmul32_fa14_6_y4);
  and_gate and_gate_h_u_arrmul32_and15_6_y0(a_15, b_6, h_u_arrmul32_and15_6_y0);
  fa fa_h_u_arrmul32_fa15_6_y2(h_u_arrmul32_and15_6_y0, h_u_arrmul32_fa16_5_y2, h_u_arrmul32_fa14_6_y4, h_u_arrmul32_fa15_6_y2, h_u_arrmul32_fa15_6_y4);
  and_gate and_gate_h_u_arrmul32_and16_6_y0(a_16, b_6, h_u_arrmul32_and16_6_y0);
  fa fa_h_u_arrmul32_fa16_6_y2(h_u_arrmul32_and16_6_y0, h_u_arrmul32_fa17_5_y2, h_u_arrmul32_fa15_6_y4, h_u_arrmul32_fa16_6_y2, h_u_arrmul32_fa16_6_y4);
  and_gate and_gate_h_u_arrmul32_and17_6_y0(a_17, b_6, h_u_arrmul32_and17_6_y0);
  fa fa_h_u_arrmul32_fa17_6_y2(h_u_arrmul32_and17_6_y0, h_u_arrmul32_fa18_5_y2, h_u_arrmul32_fa16_6_y4, h_u_arrmul32_fa17_6_y2, h_u_arrmul32_fa17_6_y4);
  and_gate and_gate_h_u_arrmul32_and18_6_y0(a_18, b_6, h_u_arrmul32_and18_6_y0);
  fa fa_h_u_arrmul32_fa18_6_y2(h_u_arrmul32_and18_6_y0, h_u_arrmul32_fa19_5_y2, h_u_arrmul32_fa17_6_y4, h_u_arrmul32_fa18_6_y2, h_u_arrmul32_fa18_6_y4);
  and_gate and_gate_h_u_arrmul32_and19_6_y0(a_19, b_6, h_u_arrmul32_and19_6_y0);
  fa fa_h_u_arrmul32_fa19_6_y2(h_u_arrmul32_and19_6_y0, h_u_arrmul32_fa20_5_y2, h_u_arrmul32_fa18_6_y4, h_u_arrmul32_fa19_6_y2, h_u_arrmul32_fa19_6_y4);
  and_gate and_gate_h_u_arrmul32_and20_6_y0(a_20, b_6, h_u_arrmul32_and20_6_y0);
  fa fa_h_u_arrmul32_fa20_6_y2(h_u_arrmul32_and20_6_y0, h_u_arrmul32_fa21_5_y2, h_u_arrmul32_fa19_6_y4, h_u_arrmul32_fa20_6_y2, h_u_arrmul32_fa20_6_y4);
  and_gate and_gate_h_u_arrmul32_and21_6_y0(a_21, b_6, h_u_arrmul32_and21_6_y0);
  fa fa_h_u_arrmul32_fa21_6_y2(h_u_arrmul32_and21_6_y0, h_u_arrmul32_fa22_5_y2, h_u_arrmul32_fa20_6_y4, h_u_arrmul32_fa21_6_y2, h_u_arrmul32_fa21_6_y4);
  and_gate and_gate_h_u_arrmul32_and22_6_y0(a_22, b_6, h_u_arrmul32_and22_6_y0);
  fa fa_h_u_arrmul32_fa22_6_y2(h_u_arrmul32_and22_6_y0, h_u_arrmul32_fa23_5_y2, h_u_arrmul32_fa21_6_y4, h_u_arrmul32_fa22_6_y2, h_u_arrmul32_fa22_6_y4);
  and_gate and_gate_h_u_arrmul32_and23_6_y0(a_23, b_6, h_u_arrmul32_and23_6_y0);
  fa fa_h_u_arrmul32_fa23_6_y2(h_u_arrmul32_and23_6_y0, h_u_arrmul32_fa24_5_y2, h_u_arrmul32_fa22_6_y4, h_u_arrmul32_fa23_6_y2, h_u_arrmul32_fa23_6_y4);
  and_gate and_gate_h_u_arrmul32_and24_6_y0(a_24, b_6, h_u_arrmul32_and24_6_y0);
  fa fa_h_u_arrmul32_fa24_6_y2(h_u_arrmul32_and24_6_y0, h_u_arrmul32_fa25_5_y2, h_u_arrmul32_fa23_6_y4, h_u_arrmul32_fa24_6_y2, h_u_arrmul32_fa24_6_y4);
  and_gate and_gate_h_u_arrmul32_and25_6_y0(a_25, b_6, h_u_arrmul32_and25_6_y0);
  fa fa_h_u_arrmul32_fa25_6_y2(h_u_arrmul32_and25_6_y0, h_u_arrmul32_fa26_5_y2, h_u_arrmul32_fa24_6_y4, h_u_arrmul32_fa25_6_y2, h_u_arrmul32_fa25_6_y4);
  and_gate and_gate_h_u_arrmul32_and26_6_y0(a_26, b_6, h_u_arrmul32_and26_6_y0);
  fa fa_h_u_arrmul32_fa26_6_y2(h_u_arrmul32_and26_6_y0, h_u_arrmul32_fa27_5_y2, h_u_arrmul32_fa25_6_y4, h_u_arrmul32_fa26_6_y2, h_u_arrmul32_fa26_6_y4);
  and_gate and_gate_h_u_arrmul32_and27_6_y0(a_27, b_6, h_u_arrmul32_and27_6_y0);
  fa fa_h_u_arrmul32_fa27_6_y2(h_u_arrmul32_and27_6_y0, h_u_arrmul32_fa28_5_y2, h_u_arrmul32_fa26_6_y4, h_u_arrmul32_fa27_6_y2, h_u_arrmul32_fa27_6_y4);
  and_gate and_gate_h_u_arrmul32_and28_6_y0(a_28, b_6, h_u_arrmul32_and28_6_y0);
  fa fa_h_u_arrmul32_fa28_6_y2(h_u_arrmul32_and28_6_y0, h_u_arrmul32_fa29_5_y2, h_u_arrmul32_fa27_6_y4, h_u_arrmul32_fa28_6_y2, h_u_arrmul32_fa28_6_y4);
  and_gate and_gate_h_u_arrmul32_and29_6_y0(a_29, b_6, h_u_arrmul32_and29_6_y0);
  fa fa_h_u_arrmul32_fa29_6_y2(h_u_arrmul32_and29_6_y0, h_u_arrmul32_fa30_5_y2, h_u_arrmul32_fa28_6_y4, h_u_arrmul32_fa29_6_y2, h_u_arrmul32_fa29_6_y4);
  and_gate and_gate_h_u_arrmul32_and30_6_y0(a_30, b_6, h_u_arrmul32_and30_6_y0);
  fa fa_h_u_arrmul32_fa30_6_y2(h_u_arrmul32_and30_6_y0, h_u_arrmul32_fa31_5_y2, h_u_arrmul32_fa29_6_y4, h_u_arrmul32_fa30_6_y2, h_u_arrmul32_fa30_6_y4);
  and_gate and_gate_h_u_arrmul32_and31_6_y0(a_31, b_6, h_u_arrmul32_and31_6_y0);
  fa fa_h_u_arrmul32_fa31_6_y2(h_u_arrmul32_and31_6_y0, h_u_arrmul32_fa31_5_y4, h_u_arrmul32_fa30_6_y4, h_u_arrmul32_fa31_6_y2, h_u_arrmul32_fa31_6_y4);
  and_gate and_gate_h_u_arrmul32_and0_7_y0(a_0, b_7, h_u_arrmul32_and0_7_y0);
  ha ha_h_u_arrmul32_ha0_7_y0(h_u_arrmul32_and0_7_y0, h_u_arrmul32_fa1_6_y2, h_u_arrmul32_ha0_7_y0, h_u_arrmul32_ha0_7_y1);
  and_gate and_gate_h_u_arrmul32_and1_7_y0(a_1, b_7, h_u_arrmul32_and1_7_y0);
  fa fa_h_u_arrmul32_fa1_7_y2(h_u_arrmul32_and1_7_y0, h_u_arrmul32_fa2_6_y2, h_u_arrmul32_ha0_7_y1, h_u_arrmul32_fa1_7_y2, h_u_arrmul32_fa1_7_y4);
  and_gate and_gate_h_u_arrmul32_and2_7_y0(a_2, b_7, h_u_arrmul32_and2_7_y0);
  fa fa_h_u_arrmul32_fa2_7_y2(h_u_arrmul32_and2_7_y0, h_u_arrmul32_fa3_6_y2, h_u_arrmul32_fa1_7_y4, h_u_arrmul32_fa2_7_y2, h_u_arrmul32_fa2_7_y4);
  and_gate and_gate_h_u_arrmul32_and3_7_y0(a_3, b_7, h_u_arrmul32_and3_7_y0);
  fa fa_h_u_arrmul32_fa3_7_y2(h_u_arrmul32_and3_7_y0, h_u_arrmul32_fa4_6_y2, h_u_arrmul32_fa2_7_y4, h_u_arrmul32_fa3_7_y2, h_u_arrmul32_fa3_7_y4);
  and_gate and_gate_h_u_arrmul32_and4_7_y0(a_4, b_7, h_u_arrmul32_and4_7_y0);
  fa fa_h_u_arrmul32_fa4_7_y2(h_u_arrmul32_and4_7_y0, h_u_arrmul32_fa5_6_y2, h_u_arrmul32_fa3_7_y4, h_u_arrmul32_fa4_7_y2, h_u_arrmul32_fa4_7_y4);
  and_gate and_gate_h_u_arrmul32_and5_7_y0(a_5, b_7, h_u_arrmul32_and5_7_y0);
  fa fa_h_u_arrmul32_fa5_7_y2(h_u_arrmul32_and5_7_y0, h_u_arrmul32_fa6_6_y2, h_u_arrmul32_fa4_7_y4, h_u_arrmul32_fa5_7_y2, h_u_arrmul32_fa5_7_y4);
  and_gate and_gate_h_u_arrmul32_and6_7_y0(a_6, b_7, h_u_arrmul32_and6_7_y0);
  fa fa_h_u_arrmul32_fa6_7_y2(h_u_arrmul32_and6_7_y0, h_u_arrmul32_fa7_6_y2, h_u_arrmul32_fa5_7_y4, h_u_arrmul32_fa6_7_y2, h_u_arrmul32_fa6_7_y4);
  and_gate and_gate_h_u_arrmul32_and7_7_y0(a_7, b_7, h_u_arrmul32_and7_7_y0);
  fa fa_h_u_arrmul32_fa7_7_y2(h_u_arrmul32_and7_7_y0, h_u_arrmul32_fa8_6_y2, h_u_arrmul32_fa6_7_y4, h_u_arrmul32_fa7_7_y2, h_u_arrmul32_fa7_7_y4);
  and_gate and_gate_h_u_arrmul32_and8_7_y0(a_8, b_7, h_u_arrmul32_and8_7_y0);
  fa fa_h_u_arrmul32_fa8_7_y2(h_u_arrmul32_and8_7_y0, h_u_arrmul32_fa9_6_y2, h_u_arrmul32_fa7_7_y4, h_u_arrmul32_fa8_7_y2, h_u_arrmul32_fa8_7_y4);
  and_gate and_gate_h_u_arrmul32_and9_7_y0(a_9, b_7, h_u_arrmul32_and9_7_y0);
  fa fa_h_u_arrmul32_fa9_7_y2(h_u_arrmul32_and9_7_y0, h_u_arrmul32_fa10_6_y2, h_u_arrmul32_fa8_7_y4, h_u_arrmul32_fa9_7_y2, h_u_arrmul32_fa9_7_y4);
  and_gate and_gate_h_u_arrmul32_and10_7_y0(a_10, b_7, h_u_arrmul32_and10_7_y0);
  fa fa_h_u_arrmul32_fa10_7_y2(h_u_arrmul32_and10_7_y0, h_u_arrmul32_fa11_6_y2, h_u_arrmul32_fa9_7_y4, h_u_arrmul32_fa10_7_y2, h_u_arrmul32_fa10_7_y4);
  and_gate and_gate_h_u_arrmul32_and11_7_y0(a_11, b_7, h_u_arrmul32_and11_7_y0);
  fa fa_h_u_arrmul32_fa11_7_y2(h_u_arrmul32_and11_7_y0, h_u_arrmul32_fa12_6_y2, h_u_arrmul32_fa10_7_y4, h_u_arrmul32_fa11_7_y2, h_u_arrmul32_fa11_7_y4);
  and_gate and_gate_h_u_arrmul32_and12_7_y0(a_12, b_7, h_u_arrmul32_and12_7_y0);
  fa fa_h_u_arrmul32_fa12_7_y2(h_u_arrmul32_and12_7_y0, h_u_arrmul32_fa13_6_y2, h_u_arrmul32_fa11_7_y4, h_u_arrmul32_fa12_7_y2, h_u_arrmul32_fa12_7_y4);
  and_gate and_gate_h_u_arrmul32_and13_7_y0(a_13, b_7, h_u_arrmul32_and13_7_y0);
  fa fa_h_u_arrmul32_fa13_7_y2(h_u_arrmul32_and13_7_y0, h_u_arrmul32_fa14_6_y2, h_u_arrmul32_fa12_7_y4, h_u_arrmul32_fa13_7_y2, h_u_arrmul32_fa13_7_y4);
  and_gate and_gate_h_u_arrmul32_and14_7_y0(a_14, b_7, h_u_arrmul32_and14_7_y0);
  fa fa_h_u_arrmul32_fa14_7_y2(h_u_arrmul32_and14_7_y0, h_u_arrmul32_fa15_6_y2, h_u_arrmul32_fa13_7_y4, h_u_arrmul32_fa14_7_y2, h_u_arrmul32_fa14_7_y4);
  and_gate and_gate_h_u_arrmul32_and15_7_y0(a_15, b_7, h_u_arrmul32_and15_7_y0);
  fa fa_h_u_arrmul32_fa15_7_y2(h_u_arrmul32_and15_7_y0, h_u_arrmul32_fa16_6_y2, h_u_arrmul32_fa14_7_y4, h_u_arrmul32_fa15_7_y2, h_u_arrmul32_fa15_7_y4);
  and_gate and_gate_h_u_arrmul32_and16_7_y0(a_16, b_7, h_u_arrmul32_and16_7_y0);
  fa fa_h_u_arrmul32_fa16_7_y2(h_u_arrmul32_and16_7_y0, h_u_arrmul32_fa17_6_y2, h_u_arrmul32_fa15_7_y4, h_u_arrmul32_fa16_7_y2, h_u_arrmul32_fa16_7_y4);
  and_gate and_gate_h_u_arrmul32_and17_7_y0(a_17, b_7, h_u_arrmul32_and17_7_y0);
  fa fa_h_u_arrmul32_fa17_7_y2(h_u_arrmul32_and17_7_y0, h_u_arrmul32_fa18_6_y2, h_u_arrmul32_fa16_7_y4, h_u_arrmul32_fa17_7_y2, h_u_arrmul32_fa17_7_y4);
  and_gate and_gate_h_u_arrmul32_and18_7_y0(a_18, b_7, h_u_arrmul32_and18_7_y0);
  fa fa_h_u_arrmul32_fa18_7_y2(h_u_arrmul32_and18_7_y0, h_u_arrmul32_fa19_6_y2, h_u_arrmul32_fa17_7_y4, h_u_arrmul32_fa18_7_y2, h_u_arrmul32_fa18_7_y4);
  and_gate and_gate_h_u_arrmul32_and19_7_y0(a_19, b_7, h_u_arrmul32_and19_7_y0);
  fa fa_h_u_arrmul32_fa19_7_y2(h_u_arrmul32_and19_7_y0, h_u_arrmul32_fa20_6_y2, h_u_arrmul32_fa18_7_y4, h_u_arrmul32_fa19_7_y2, h_u_arrmul32_fa19_7_y4);
  and_gate and_gate_h_u_arrmul32_and20_7_y0(a_20, b_7, h_u_arrmul32_and20_7_y0);
  fa fa_h_u_arrmul32_fa20_7_y2(h_u_arrmul32_and20_7_y0, h_u_arrmul32_fa21_6_y2, h_u_arrmul32_fa19_7_y4, h_u_arrmul32_fa20_7_y2, h_u_arrmul32_fa20_7_y4);
  and_gate and_gate_h_u_arrmul32_and21_7_y0(a_21, b_7, h_u_arrmul32_and21_7_y0);
  fa fa_h_u_arrmul32_fa21_7_y2(h_u_arrmul32_and21_7_y0, h_u_arrmul32_fa22_6_y2, h_u_arrmul32_fa20_7_y4, h_u_arrmul32_fa21_7_y2, h_u_arrmul32_fa21_7_y4);
  and_gate and_gate_h_u_arrmul32_and22_7_y0(a_22, b_7, h_u_arrmul32_and22_7_y0);
  fa fa_h_u_arrmul32_fa22_7_y2(h_u_arrmul32_and22_7_y0, h_u_arrmul32_fa23_6_y2, h_u_arrmul32_fa21_7_y4, h_u_arrmul32_fa22_7_y2, h_u_arrmul32_fa22_7_y4);
  and_gate and_gate_h_u_arrmul32_and23_7_y0(a_23, b_7, h_u_arrmul32_and23_7_y0);
  fa fa_h_u_arrmul32_fa23_7_y2(h_u_arrmul32_and23_7_y0, h_u_arrmul32_fa24_6_y2, h_u_arrmul32_fa22_7_y4, h_u_arrmul32_fa23_7_y2, h_u_arrmul32_fa23_7_y4);
  and_gate and_gate_h_u_arrmul32_and24_7_y0(a_24, b_7, h_u_arrmul32_and24_7_y0);
  fa fa_h_u_arrmul32_fa24_7_y2(h_u_arrmul32_and24_7_y0, h_u_arrmul32_fa25_6_y2, h_u_arrmul32_fa23_7_y4, h_u_arrmul32_fa24_7_y2, h_u_arrmul32_fa24_7_y4);
  and_gate and_gate_h_u_arrmul32_and25_7_y0(a_25, b_7, h_u_arrmul32_and25_7_y0);
  fa fa_h_u_arrmul32_fa25_7_y2(h_u_arrmul32_and25_7_y0, h_u_arrmul32_fa26_6_y2, h_u_arrmul32_fa24_7_y4, h_u_arrmul32_fa25_7_y2, h_u_arrmul32_fa25_7_y4);
  and_gate and_gate_h_u_arrmul32_and26_7_y0(a_26, b_7, h_u_arrmul32_and26_7_y0);
  fa fa_h_u_arrmul32_fa26_7_y2(h_u_arrmul32_and26_7_y0, h_u_arrmul32_fa27_6_y2, h_u_arrmul32_fa25_7_y4, h_u_arrmul32_fa26_7_y2, h_u_arrmul32_fa26_7_y4);
  and_gate and_gate_h_u_arrmul32_and27_7_y0(a_27, b_7, h_u_arrmul32_and27_7_y0);
  fa fa_h_u_arrmul32_fa27_7_y2(h_u_arrmul32_and27_7_y0, h_u_arrmul32_fa28_6_y2, h_u_arrmul32_fa26_7_y4, h_u_arrmul32_fa27_7_y2, h_u_arrmul32_fa27_7_y4);
  and_gate and_gate_h_u_arrmul32_and28_7_y0(a_28, b_7, h_u_arrmul32_and28_7_y0);
  fa fa_h_u_arrmul32_fa28_7_y2(h_u_arrmul32_and28_7_y0, h_u_arrmul32_fa29_6_y2, h_u_arrmul32_fa27_7_y4, h_u_arrmul32_fa28_7_y2, h_u_arrmul32_fa28_7_y4);
  and_gate and_gate_h_u_arrmul32_and29_7_y0(a_29, b_7, h_u_arrmul32_and29_7_y0);
  fa fa_h_u_arrmul32_fa29_7_y2(h_u_arrmul32_and29_7_y0, h_u_arrmul32_fa30_6_y2, h_u_arrmul32_fa28_7_y4, h_u_arrmul32_fa29_7_y2, h_u_arrmul32_fa29_7_y4);
  and_gate and_gate_h_u_arrmul32_and30_7_y0(a_30, b_7, h_u_arrmul32_and30_7_y0);
  fa fa_h_u_arrmul32_fa30_7_y2(h_u_arrmul32_and30_7_y0, h_u_arrmul32_fa31_6_y2, h_u_arrmul32_fa29_7_y4, h_u_arrmul32_fa30_7_y2, h_u_arrmul32_fa30_7_y4);
  and_gate and_gate_h_u_arrmul32_and31_7_y0(a_31, b_7, h_u_arrmul32_and31_7_y0);
  fa fa_h_u_arrmul32_fa31_7_y2(h_u_arrmul32_and31_7_y0, h_u_arrmul32_fa31_6_y4, h_u_arrmul32_fa30_7_y4, h_u_arrmul32_fa31_7_y2, h_u_arrmul32_fa31_7_y4);
  and_gate and_gate_h_u_arrmul32_and0_8_y0(a_0, b_8, h_u_arrmul32_and0_8_y0);
  ha ha_h_u_arrmul32_ha0_8_y0(h_u_arrmul32_and0_8_y0, h_u_arrmul32_fa1_7_y2, h_u_arrmul32_ha0_8_y0, h_u_arrmul32_ha0_8_y1);
  and_gate and_gate_h_u_arrmul32_and1_8_y0(a_1, b_8, h_u_arrmul32_and1_8_y0);
  fa fa_h_u_arrmul32_fa1_8_y2(h_u_arrmul32_and1_8_y0, h_u_arrmul32_fa2_7_y2, h_u_arrmul32_ha0_8_y1, h_u_arrmul32_fa1_8_y2, h_u_arrmul32_fa1_8_y4);
  and_gate and_gate_h_u_arrmul32_and2_8_y0(a_2, b_8, h_u_arrmul32_and2_8_y0);
  fa fa_h_u_arrmul32_fa2_8_y2(h_u_arrmul32_and2_8_y0, h_u_arrmul32_fa3_7_y2, h_u_arrmul32_fa1_8_y4, h_u_arrmul32_fa2_8_y2, h_u_arrmul32_fa2_8_y4);
  and_gate and_gate_h_u_arrmul32_and3_8_y0(a_3, b_8, h_u_arrmul32_and3_8_y0);
  fa fa_h_u_arrmul32_fa3_8_y2(h_u_arrmul32_and3_8_y0, h_u_arrmul32_fa4_7_y2, h_u_arrmul32_fa2_8_y4, h_u_arrmul32_fa3_8_y2, h_u_arrmul32_fa3_8_y4);
  and_gate and_gate_h_u_arrmul32_and4_8_y0(a_4, b_8, h_u_arrmul32_and4_8_y0);
  fa fa_h_u_arrmul32_fa4_8_y2(h_u_arrmul32_and4_8_y0, h_u_arrmul32_fa5_7_y2, h_u_arrmul32_fa3_8_y4, h_u_arrmul32_fa4_8_y2, h_u_arrmul32_fa4_8_y4);
  and_gate and_gate_h_u_arrmul32_and5_8_y0(a_5, b_8, h_u_arrmul32_and5_8_y0);
  fa fa_h_u_arrmul32_fa5_8_y2(h_u_arrmul32_and5_8_y0, h_u_arrmul32_fa6_7_y2, h_u_arrmul32_fa4_8_y4, h_u_arrmul32_fa5_8_y2, h_u_arrmul32_fa5_8_y4);
  and_gate and_gate_h_u_arrmul32_and6_8_y0(a_6, b_8, h_u_arrmul32_and6_8_y0);
  fa fa_h_u_arrmul32_fa6_8_y2(h_u_arrmul32_and6_8_y0, h_u_arrmul32_fa7_7_y2, h_u_arrmul32_fa5_8_y4, h_u_arrmul32_fa6_8_y2, h_u_arrmul32_fa6_8_y4);
  and_gate and_gate_h_u_arrmul32_and7_8_y0(a_7, b_8, h_u_arrmul32_and7_8_y0);
  fa fa_h_u_arrmul32_fa7_8_y2(h_u_arrmul32_and7_8_y0, h_u_arrmul32_fa8_7_y2, h_u_arrmul32_fa6_8_y4, h_u_arrmul32_fa7_8_y2, h_u_arrmul32_fa7_8_y4);
  and_gate and_gate_h_u_arrmul32_and8_8_y0(a_8, b_8, h_u_arrmul32_and8_8_y0);
  fa fa_h_u_arrmul32_fa8_8_y2(h_u_arrmul32_and8_8_y0, h_u_arrmul32_fa9_7_y2, h_u_arrmul32_fa7_8_y4, h_u_arrmul32_fa8_8_y2, h_u_arrmul32_fa8_8_y4);
  and_gate and_gate_h_u_arrmul32_and9_8_y0(a_9, b_8, h_u_arrmul32_and9_8_y0);
  fa fa_h_u_arrmul32_fa9_8_y2(h_u_arrmul32_and9_8_y0, h_u_arrmul32_fa10_7_y2, h_u_arrmul32_fa8_8_y4, h_u_arrmul32_fa9_8_y2, h_u_arrmul32_fa9_8_y4);
  and_gate and_gate_h_u_arrmul32_and10_8_y0(a_10, b_8, h_u_arrmul32_and10_8_y0);
  fa fa_h_u_arrmul32_fa10_8_y2(h_u_arrmul32_and10_8_y0, h_u_arrmul32_fa11_7_y2, h_u_arrmul32_fa9_8_y4, h_u_arrmul32_fa10_8_y2, h_u_arrmul32_fa10_8_y4);
  and_gate and_gate_h_u_arrmul32_and11_8_y0(a_11, b_8, h_u_arrmul32_and11_8_y0);
  fa fa_h_u_arrmul32_fa11_8_y2(h_u_arrmul32_and11_8_y0, h_u_arrmul32_fa12_7_y2, h_u_arrmul32_fa10_8_y4, h_u_arrmul32_fa11_8_y2, h_u_arrmul32_fa11_8_y4);
  and_gate and_gate_h_u_arrmul32_and12_8_y0(a_12, b_8, h_u_arrmul32_and12_8_y0);
  fa fa_h_u_arrmul32_fa12_8_y2(h_u_arrmul32_and12_8_y0, h_u_arrmul32_fa13_7_y2, h_u_arrmul32_fa11_8_y4, h_u_arrmul32_fa12_8_y2, h_u_arrmul32_fa12_8_y4);
  and_gate and_gate_h_u_arrmul32_and13_8_y0(a_13, b_8, h_u_arrmul32_and13_8_y0);
  fa fa_h_u_arrmul32_fa13_8_y2(h_u_arrmul32_and13_8_y0, h_u_arrmul32_fa14_7_y2, h_u_arrmul32_fa12_8_y4, h_u_arrmul32_fa13_8_y2, h_u_arrmul32_fa13_8_y4);
  and_gate and_gate_h_u_arrmul32_and14_8_y0(a_14, b_8, h_u_arrmul32_and14_8_y0);
  fa fa_h_u_arrmul32_fa14_8_y2(h_u_arrmul32_and14_8_y0, h_u_arrmul32_fa15_7_y2, h_u_arrmul32_fa13_8_y4, h_u_arrmul32_fa14_8_y2, h_u_arrmul32_fa14_8_y4);
  and_gate and_gate_h_u_arrmul32_and15_8_y0(a_15, b_8, h_u_arrmul32_and15_8_y0);
  fa fa_h_u_arrmul32_fa15_8_y2(h_u_arrmul32_and15_8_y0, h_u_arrmul32_fa16_7_y2, h_u_arrmul32_fa14_8_y4, h_u_arrmul32_fa15_8_y2, h_u_arrmul32_fa15_8_y4);
  and_gate and_gate_h_u_arrmul32_and16_8_y0(a_16, b_8, h_u_arrmul32_and16_8_y0);
  fa fa_h_u_arrmul32_fa16_8_y2(h_u_arrmul32_and16_8_y0, h_u_arrmul32_fa17_7_y2, h_u_arrmul32_fa15_8_y4, h_u_arrmul32_fa16_8_y2, h_u_arrmul32_fa16_8_y4);
  and_gate and_gate_h_u_arrmul32_and17_8_y0(a_17, b_8, h_u_arrmul32_and17_8_y0);
  fa fa_h_u_arrmul32_fa17_8_y2(h_u_arrmul32_and17_8_y0, h_u_arrmul32_fa18_7_y2, h_u_arrmul32_fa16_8_y4, h_u_arrmul32_fa17_8_y2, h_u_arrmul32_fa17_8_y4);
  and_gate and_gate_h_u_arrmul32_and18_8_y0(a_18, b_8, h_u_arrmul32_and18_8_y0);
  fa fa_h_u_arrmul32_fa18_8_y2(h_u_arrmul32_and18_8_y0, h_u_arrmul32_fa19_7_y2, h_u_arrmul32_fa17_8_y4, h_u_arrmul32_fa18_8_y2, h_u_arrmul32_fa18_8_y4);
  and_gate and_gate_h_u_arrmul32_and19_8_y0(a_19, b_8, h_u_arrmul32_and19_8_y0);
  fa fa_h_u_arrmul32_fa19_8_y2(h_u_arrmul32_and19_8_y0, h_u_arrmul32_fa20_7_y2, h_u_arrmul32_fa18_8_y4, h_u_arrmul32_fa19_8_y2, h_u_arrmul32_fa19_8_y4);
  and_gate and_gate_h_u_arrmul32_and20_8_y0(a_20, b_8, h_u_arrmul32_and20_8_y0);
  fa fa_h_u_arrmul32_fa20_8_y2(h_u_arrmul32_and20_8_y0, h_u_arrmul32_fa21_7_y2, h_u_arrmul32_fa19_8_y4, h_u_arrmul32_fa20_8_y2, h_u_arrmul32_fa20_8_y4);
  and_gate and_gate_h_u_arrmul32_and21_8_y0(a_21, b_8, h_u_arrmul32_and21_8_y0);
  fa fa_h_u_arrmul32_fa21_8_y2(h_u_arrmul32_and21_8_y0, h_u_arrmul32_fa22_7_y2, h_u_arrmul32_fa20_8_y4, h_u_arrmul32_fa21_8_y2, h_u_arrmul32_fa21_8_y4);
  and_gate and_gate_h_u_arrmul32_and22_8_y0(a_22, b_8, h_u_arrmul32_and22_8_y0);
  fa fa_h_u_arrmul32_fa22_8_y2(h_u_arrmul32_and22_8_y0, h_u_arrmul32_fa23_7_y2, h_u_arrmul32_fa21_8_y4, h_u_arrmul32_fa22_8_y2, h_u_arrmul32_fa22_8_y4);
  and_gate and_gate_h_u_arrmul32_and23_8_y0(a_23, b_8, h_u_arrmul32_and23_8_y0);
  fa fa_h_u_arrmul32_fa23_8_y2(h_u_arrmul32_and23_8_y0, h_u_arrmul32_fa24_7_y2, h_u_arrmul32_fa22_8_y4, h_u_arrmul32_fa23_8_y2, h_u_arrmul32_fa23_8_y4);
  and_gate and_gate_h_u_arrmul32_and24_8_y0(a_24, b_8, h_u_arrmul32_and24_8_y0);
  fa fa_h_u_arrmul32_fa24_8_y2(h_u_arrmul32_and24_8_y0, h_u_arrmul32_fa25_7_y2, h_u_arrmul32_fa23_8_y4, h_u_arrmul32_fa24_8_y2, h_u_arrmul32_fa24_8_y4);
  and_gate and_gate_h_u_arrmul32_and25_8_y0(a_25, b_8, h_u_arrmul32_and25_8_y0);
  fa fa_h_u_arrmul32_fa25_8_y2(h_u_arrmul32_and25_8_y0, h_u_arrmul32_fa26_7_y2, h_u_arrmul32_fa24_8_y4, h_u_arrmul32_fa25_8_y2, h_u_arrmul32_fa25_8_y4);
  and_gate and_gate_h_u_arrmul32_and26_8_y0(a_26, b_8, h_u_arrmul32_and26_8_y0);
  fa fa_h_u_arrmul32_fa26_8_y2(h_u_arrmul32_and26_8_y0, h_u_arrmul32_fa27_7_y2, h_u_arrmul32_fa25_8_y4, h_u_arrmul32_fa26_8_y2, h_u_arrmul32_fa26_8_y4);
  and_gate and_gate_h_u_arrmul32_and27_8_y0(a_27, b_8, h_u_arrmul32_and27_8_y0);
  fa fa_h_u_arrmul32_fa27_8_y2(h_u_arrmul32_and27_8_y0, h_u_arrmul32_fa28_7_y2, h_u_arrmul32_fa26_8_y4, h_u_arrmul32_fa27_8_y2, h_u_arrmul32_fa27_8_y4);
  and_gate and_gate_h_u_arrmul32_and28_8_y0(a_28, b_8, h_u_arrmul32_and28_8_y0);
  fa fa_h_u_arrmul32_fa28_8_y2(h_u_arrmul32_and28_8_y0, h_u_arrmul32_fa29_7_y2, h_u_arrmul32_fa27_8_y4, h_u_arrmul32_fa28_8_y2, h_u_arrmul32_fa28_8_y4);
  and_gate and_gate_h_u_arrmul32_and29_8_y0(a_29, b_8, h_u_arrmul32_and29_8_y0);
  fa fa_h_u_arrmul32_fa29_8_y2(h_u_arrmul32_and29_8_y0, h_u_arrmul32_fa30_7_y2, h_u_arrmul32_fa28_8_y4, h_u_arrmul32_fa29_8_y2, h_u_arrmul32_fa29_8_y4);
  and_gate and_gate_h_u_arrmul32_and30_8_y0(a_30, b_8, h_u_arrmul32_and30_8_y0);
  fa fa_h_u_arrmul32_fa30_8_y2(h_u_arrmul32_and30_8_y0, h_u_arrmul32_fa31_7_y2, h_u_arrmul32_fa29_8_y4, h_u_arrmul32_fa30_8_y2, h_u_arrmul32_fa30_8_y4);
  and_gate and_gate_h_u_arrmul32_and31_8_y0(a_31, b_8, h_u_arrmul32_and31_8_y0);
  fa fa_h_u_arrmul32_fa31_8_y2(h_u_arrmul32_and31_8_y0, h_u_arrmul32_fa31_7_y4, h_u_arrmul32_fa30_8_y4, h_u_arrmul32_fa31_8_y2, h_u_arrmul32_fa31_8_y4);
  and_gate and_gate_h_u_arrmul32_and0_9_y0(a_0, b_9, h_u_arrmul32_and0_9_y0);
  ha ha_h_u_arrmul32_ha0_9_y0(h_u_arrmul32_and0_9_y0, h_u_arrmul32_fa1_8_y2, h_u_arrmul32_ha0_9_y0, h_u_arrmul32_ha0_9_y1);
  and_gate and_gate_h_u_arrmul32_and1_9_y0(a_1, b_9, h_u_arrmul32_and1_9_y0);
  fa fa_h_u_arrmul32_fa1_9_y2(h_u_arrmul32_and1_9_y0, h_u_arrmul32_fa2_8_y2, h_u_arrmul32_ha0_9_y1, h_u_arrmul32_fa1_9_y2, h_u_arrmul32_fa1_9_y4);
  and_gate and_gate_h_u_arrmul32_and2_9_y0(a_2, b_9, h_u_arrmul32_and2_9_y0);
  fa fa_h_u_arrmul32_fa2_9_y2(h_u_arrmul32_and2_9_y0, h_u_arrmul32_fa3_8_y2, h_u_arrmul32_fa1_9_y4, h_u_arrmul32_fa2_9_y2, h_u_arrmul32_fa2_9_y4);
  and_gate and_gate_h_u_arrmul32_and3_9_y0(a_3, b_9, h_u_arrmul32_and3_9_y0);
  fa fa_h_u_arrmul32_fa3_9_y2(h_u_arrmul32_and3_9_y0, h_u_arrmul32_fa4_8_y2, h_u_arrmul32_fa2_9_y4, h_u_arrmul32_fa3_9_y2, h_u_arrmul32_fa3_9_y4);
  and_gate and_gate_h_u_arrmul32_and4_9_y0(a_4, b_9, h_u_arrmul32_and4_9_y0);
  fa fa_h_u_arrmul32_fa4_9_y2(h_u_arrmul32_and4_9_y0, h_u_arrmul32_fa5_8_y2, h_u_arrmul32_fa3_9_y4, h_u_arrmul32_fa4_9_y2, h_u_arrmul32_fa4_9_y4);
  and_gate and_gate_h_u_arrmul32_and5_9_y0(a_5, b_9, h_u_arrmul32_and5_9_y0);
  fa fa_h_u_arrmul32_fa5_9_y2(h_u_arrmul32_and5_9_y0, h_u_arrmul32_fa6_8_y2, h_u_arrmul32_fa4_9_y4, h_u_arrmul32_fa5_9_y2, h_u_arrmul32_fa5_9_y4);
  and_gate and_gate_h_u_arrmul32_and6_9_y0(a_6, b_9, h_u_arrmul32_and6_9_y0);
  fa fa_h_u_arrmul32_fa6_9_y2(h_u_arrmul32_and6_9_y0, h_u_arrmul32_fa7_8_y2, h_u_arrmul32_fa5_9_y4, h_u_arrmul32_fa6_9_y2, h_u_arrmul32_fa6_9_y4);
  and_gate and_gate_h_u_arrmul32_and7_9_y0(a_7, b_9, h_u_arrmul32_and7_9_y0);
  fa fa_h_u_arrmul32_fa7_9_y2(h_u_arrmul32_and7_9_y0, h_u_arrmul32_fa8_8_y2, h_u_arrmul32_fa6_9_y4, h_u_arrmul32_fa7_9_y2, h_u_arrmul32_fa7_9_y4);
  and_gate and_gate_h_u_arrmul32_and8_9_y0(a_8, b_9, h_u_arrmul32_and8_9_y0);
  fa fa_h_u_arrmul32_fa8_9_y2(h_u_arrmul32_and8_9_y0, h_u_arrmul32_fa9_8_y2, h_u_arrmul32_fa7_9_y4, h_u_arrmul32_fa8_9_y2, h_u_arrmul32_fa8_9_y4);
  and_gate and_gate_h_u_arrmul32_and9_9_y0(a_9, b_9, h_u_arrmul32_and9_9_y0);
  fa fa_h_u_arrmul32_fa9_9_y2(h_u_arrmul32_and9_9_y0, h_u_arrmul32_fa10_8_y2, h_u_arrmul32_fa8_9_y4, h_u_arrmul32_fa9_9_y2, h_u_arrmul32_fa9_9_y4);
  and_gate and_gate_h_u_arrmul32_and10_9_y0(a_10, b_9, h_u_arrmul32_and10_9_y0);
  fa fa_h_u_arrmul32_fa10_9_y2(h_u_arrmul32_and10_9_y0, h_u_arrmul32_fa11_8_y2, h_u_arrmul32_fa9_9_y4, h_u_arrmul32_fa10_9_y2, h_u_arrmul32_fa10_9_y4);
  and_gate and_gate_h_u_arrmul32_and11_9_y0(a_11, b_9, h_u_arrmul32_and11_9_y0);
  fa fa_h_u_arrmul32_fa11_9_y2(h_u_arrmul32_and11_9_y0, h_u_arrmul32_fa12_8_y2, h_u_arrmul32_fa10_9_y4, h_u_arrmul32_fa11_9_y2, h_u_arrmul32_fa11_9_y4);
  and_gate and_gate_h_u_arrmul32_and12_9_y0(a_12, b_9, h_u_arrmul32_and12_9_y0);
  fa fa_h_u_arrmul32_fa12_9_y2(h_u_arrmul32_and12_9_y0, h_u_arrmul32_fa13_8_y2, h_u_arrmul32_fa11_9_y4, h_u_arrmul32_fa12_9_y2, h_u_arrmul32_fa12_9_y4);
  and_gate and_gate_h_u_arrmul32_and13_9_y0(a_13, b_9, h_u_arrmul32_and13_9_y0);
  fa fa_h_u_arrmul32_fa13_9_y2(h_u_arrmul32_and13_9_y0, h_u_arrmul32_fa14_8_y2, h_u_arrmul32_fa12_9_y4, h_u_arrmul32_fa13_9_y2, h_u_arrmul32_fa13_9_y4);
  and_gate and_gate_h_u_arrmul32_and14_9_y0(a_14, b_9, h_u_arrmul32_and14_9_y0);
  fa fa_h_u_arrmul32_fa14_9_y2(h_u_arrmul32_and14_9_y0, h_u_arrmul32_fa15_8_y2, h_u_arrmul32_fa13_9_y4, h_u_arrmul32_fa14_9_y2, h_u_arrmul32_fa14_9_y4);
  and_gate and_gate_h_u_arrmul32_and15_9_y0(a_15, b_9, h_u_arrmul32_and15_9_y0);
  fa fa_h_u_arrmul32_fa15_9_y2(h_u_arrmul32_and15_9_y0, h_u_arrmul32_fa16_8_y2, h_u_arrmul32_fa14_9_y4, h_u_arrmul32_fa15_9_y2, h_u_arrmul32_fa15_9_y4);
  and_gate and_gate_h_u_arrmul32_and16_9_y0(a_16, b_9, h_u_arrmul32_and16_9_y0);
  fa fa_h_u_arrmul32_fa16_9_y2(h_u_arrmul32_and16_9_y0, h_u_arrmul32_fa17_8_y2, h_u_arrmul32_fa15_9_y4, h_u_arrmul32_fa16_9_y2, h_u_arrmul32_fa16_9_y4);
  and_gate and_gate_h_u_arrmul32_and17_9_y0(a_17, b_9, h_u_arrmul32_and17_9_y0);
  fa fa_h_u_arrmul32_fa17_9_y2(h_u_arrmul32_and17_9_y0, h_u_arrmul32_fa18_8_y2, h_u_arrmul32_fa16_9_y4, h_u_arrmul32_fa17_9_y2, h_u_arrmul32_fa17_9_y4);
  and_gate and_gate_h_u_arrmul32_and18_9_y0(a_18, b_9, h_u_arrmul32_and18_9_y0);
  fa fa_h_u_arrmul32_fa18_9_y2(h_u_arrmul32_and18_9_y0, h_u_arrmul32_fa19_8_y2, h_u_arrmul32_fa17_9_y4, h_u_arrmul32_fa18_9_y2, h_u_arrmul32_fa18_9_y4);
  and_gate and_gate_h_u_arrmul32_and19_9_y0(a_19, b_9, h_u_arrmul32_and19_9_y0);
  fa fa_h_u_arrmul32_fa19_9_y2(h_u_arrmul32_and19_9_y0, h_u_arrmul32_fa20_8_y2, h_u_arrmul32_fa18_9_y4, h_u_arrmul32_fa19_9_y2, h_u_arrmul32_fa19_9_y4);
  and_gate and_gate_h_u_arrmul32_and20_9_y0(a_20, b_9, h_u_arrmul32_and20_9_y0);
  fa fa_h_u_arrmul32_fa20_9_y2(h_u_arrmul32_and20_9_y0, h_u_arrmul32_fa21_8_y2, h_u_arrmul32_fa19_9_y4, h_u_arrmul32_fa20_9_y2, h_u_arrmul32_fa20_9_y4);
  and_gate and_gate_h_u_arrmul32_and21_9_y0(a_21, b_9, h_u_arrmul32_and21_9_y0);
  fa fa_h_u_arrmul32_fa21_9_y2(h_u_arrmul32_and21_9_y0, h_u_arrmul32_fa22_8_y2, h_u_arrmul32_fa20_9_y4, h_u_arrmul32_fa21_9_y2, h_u_arrmul32_fa21_9_y4);
  and_gate and_gate_h_u_arrmul32_and22_9_y0(a_22, b_9, h_u_arrmul32_and22_9_y0);
  fa fa_h_u_arrmul32_fa22_9_y2(h_u_arrmul32_and22_9_y0, h_u_arrmul32_fa23_8_y2, h_u_arrmul32_fa21_9_y4, h_u_arrmul32_fa22_9_y2, h_u_arrmul32_fa22_9_y4);
  and_gate and_gate_h_u_arrmul32_and23_9_y0(a_23, b_9, h_u_arrmul32_and23_9_y0);
  fa fa_h_u_arrmul32_fa23_9_y2(h_u_arrmul32_and23_9_y0, h_u_arrmul32_fa24_8_y2, h_u_arrmul32_fa22_9_y4, h_u_arrmul32_fa23_9_y2, h_u_arrmul32_fa23_9_y4);
  and_gate and_gate_h_u_arrmul32_and24_9_y0(a_24, b_9, h_u_arrmul32_and24_9_y0);
  fa fa_h_u_arrmul32_fa24_9_y2(h_u_arrmul32_and24_9_y0, h_u_arrmul32_fa25_8_y2, h_u_arrmul32_fa23_9_y4, h_u_arrmul32_fa24_9_y2, h_u_arrmul32_fa24_9_y4);
  and_gate and_gate_h_u_arrmul32_and25_9_y0(a_25, b_9, h_u_arrmul32_and25_9_y0);
  fa fa_h_u_arrmul32_fa25_9_y2(h_u_arrmul32_and25_9_y0, h_u_arrmul32_fa26_8_y2, h_u_arrmul32_fa24_9_y4, h_u_arrmul32_fa25_9_y2, h_u_arrmul32_fa25_9_y4);
  and_gate and_gate_h_u_arrmul32_and26_9_y0(a_26, b_9, h_u_arrmul32_and26_9_y0);
  fa fa_h_u_arrmul32_fa26_9_y2(h_u_arrmul32_and26_9_y0, h_u_arrmul32_fa27_8_y2, h_u_arrmul32_fa25_9_y4, h_u_arrmul32_fa26_9_y2, h_u_arrmul32_fa26_9_y4);
  and_gate and_gate_h_u_arrmul32_and27_9_y0(a_27, b_9, h_u_arrmul32_and27_9_y0);
  fa fa_h_u_arrmul32_fa27_9_y2(h_u_arrmul32_and27_9_y0, h_u_arrmul32_fa28_8_y2, h_u_arrmul32_fa26_9_y4, h_u_arrmul32_fa27_9_y2, h_u_arrmul32_fa27_9_y4);
  and_gate and_gate_h_u_arrmul32_and28_9_y0(a_28, b_9, h_u_arrmul32_and28_9_y0);
  fa fa_h_u_arrmul32_fa28_9_y2(h_u_arrmul32_and28_9_y0, h_u_arrmul32_fa29_8_y2, h_u_arrmul32_fa27_9_y4, h_u_arrmul32_fa28_9_y2, h_u_arrmul32_fa28_9_y4);
  and_gate and_gate_h_u_arrmul32_and29_9_y0(a_29, b_9, h_u_arrmul32_and29_9_y0);
  fa fa_h_u_arrmul32_fa29_9_y2(h_u_arrmul32_and29_9_y0, h_u_arrmul32_fa30_8_y2, h_u_arrmul32_fa28_9_y4, h_u_arrmul32_fa29_9_y2, h_u_arrmul32_fa29_9_y4);
  and_gate and_gate_h_u_arrmul32_and30_9_y0(a_30, b_9, h_u_arrmul32_and30_9_y0);
  fa fa_h_u_arrmul32_fa30_9_y2(h_u_arrmul32_and30_9_y0, h_u_arrmul32_fa31_8_y2, h_u_arrmul32_fa29_9_y4, h_u_arrmul32_fa30_9_y2, h_u_arrmul32_fa30_9_y4);
  and_gate and_gate_h_u_arrmul32_and31_9_y0(a_31, b_9, h_u_arrmul32_and31_9_y0);
  fa fa_h_u_arrmul32_fa31_9_y2(h_u_arrmul32_and31_9_y0, h_u_arrmul32_fa31_8_y4, h_u_arrmul32_fa30_9_y4, h_u_arrmul32_fa31_9_y2, h_u_arrmul32_fa31_9_y4);
  and_gate and_gate_h_u_arrmul32_and0_10_y0(a_0, b_10, h_u_arrmul32_and0_10_y0);
  ha ha_h_u_arrmul32_ha0_10_y0(h_u_arrmul32_and0_10_y0, h_u_arrmul32_fa1_9_y2, h_u_arrmul32_ha0_10_y0, h_u_arrmul32_ha0_10_y1);
  and_gate and_gate_h_u_arrmul32_and1_10_y0(a_1, b_10, h_u_arrmul32_and1_10_y0);
  fa fa_h_u_arrmul32_fa1_10_y2(h_u_arrmul32_and1_10_y0, h_u_arrmul32_fa2_9_y2, h_u_arrmul32_ha0_10_y1, h_u_arrmul32_fa1_10_y2, h_u_arrmul32_fa1_10_y4);
  and_gate and_gate_h_u_arrmul32_and2_10_y0(a_2, b_10, h_u_arrmul32_and2_10_y0);
  fa fa_h_u_arrmul32_fa2_10_y2(h_u_arrmul32_and2_10_y0, h_u_arrmul32_fa3_9_y2, h_u_arrmul32_fa1_10_y4, h_u_arrmul32_fa2_10_y2, h_u_arrmul32_fa2_10_y4);
  and_gate and_gate_h_u_arrmul32_and3_10_y0(a_3, b_10, h_u_arrmul32_and3_10_y0);
  fa fa_h_u_arrmul32_fa3_10_y2(h_u_arrmul32_and3_10_y0, h_u_arrmul32_fa4_9_y2, h_u_arrmul32_fa2_10_y4, h_u_arrmul32_fa3_10_y2, h_u_arrmul32_fa3_10_y4);
  and_gate and_gate_h_u_arrmul32_and4_10_y0(a_4, b_10, h_u_arrmul32_and4_10_y0);
  fa fa_h_u_arrmul32_fa4_10_y2(h_u_arrmul32_and4_10_y0, h_u_arrmul32_fa5_9_y2, h_u_arrmul32_fa3_10_y4, h_u_arrmul32_fa4_10_y2, h_u_arrmul32_fa4_10_y4);
  and_gate and_gate_h_u_arrmul32_and5_10_y0(a_5, b_10, h_u_arrmul32_and5_10_y0);
  fa fa_h_u_arrmul32_fa5_10_y2(h_u_arrmul32_and5_10_y0, h_u_arrmul32_fa6_9_y2, h_u_arrmul32_fa4_10_y4, h_u_arrmul32_fa5_10_y2, h_u_arrmul32_fa5_10_y4);
  and_gate and_gate_h_u_arrmul32_and6_10_y0(a_6, b_10, h_u_arrmul32_and6_10_y0);
  fa fa_h_u_arrmul32_fa6_10_y2(h_u_arrmul32_and6_10_y0, h_u_arrmul32_fa7_9_y2, h_u_arrmul32_fa5_10_y4, h_u_arrmul32_fa6_10_y2, h_u_arrmul32_fa6_10_y4);
  and_gate and_gate_h_u_arrmul32_and7_10_y0(a_7, b_10, h_u_arrmul32_and7_10_y0);
  fa fa_h_u_arrmul32_fa7_10_y2(h_u_arrmul32_and7_10_y0, h_u_arrmul32_fa8_9_y2, h_u_arrmul32_fa6_10_y4, h_u_arrmul32_fa7_10_y2, h_u_arrmul32_fa7_10_y4);
  and_gate and_gate_h_u_arrmul32_and8_10_y0(a_8, b_10, h_u_arrmul32_and8_10_y0);
  fa fa_h_u_arrmul32_fa8_10_y2(h_u_arrmul32_and8_10_y0, h_u_arrmul32_fa9_9_y2, h_u_arrmul32_fa7_10_y4, h_u_arrmul32_fa8_10_y2, h_u_arrmul32_fa8_10_y4);
  and_gate and_gate_h_u_arrmul32_and9_10_y0(a_9, b_10, h_u_arrmul32_and9_10_y0);
  fa fa_h_u_arrmul32_fa9_10_y2(h_u_arrmul32_and9_10_y0, h_u_arrmul32_fa10_9_y2, h_u_arrmul32_fa8_10_y4, h_u_arrmul32_fa9_10_y2, h_u_arrmul32_fa9_10_y4);
  and_gate and_gate_h_u_arrmul32_and10_10_y0(a_10, b_10, h_u_arrmul32_and10_10_y0);
  fa fa_h_u_arrmul32_fa10_10_y2(h_u_arrmul32_and10_10_y0, h_u_arrmul32_fa11_9_y2, h_u_arrmul32_fa9_10_y4, h_u_arrmul32_fa10_10_y2, h_u_arrmul32_fa10_10_y4);
  and_gate and_gate_h_u_arrmul32_and11_10_y0(a_11, b_10, h_u_arrmul32_and11_10_y0);
  fa fa_h_u_arrmul32_fa11_10_y2(h_u_arrmul32_and11_10_y0, h_u_arrmul32_fa12_9_y2, h_u_arrmul32_fa10_10_y4, h_u_arrmul32_fa11_10_y2, h_u_arrmul32_fa11_10_y4);
  and_gate and_gate_h_u_arrmul32_and12_10_y0(a_12, b_10, h_u_arrmul32_and12_10_y0);
  fa fa_h_u_arrmul32_fa12_10_y2(h_u_arrmul32_and12_10_y0, h_u_arrmul32_fa13_9_y2, h_u_arrmul32_fa11_10_y4, h_u_arrmul32_fa12_10_y2, h_u_arrmul32_fa12_10_y4);
  and_gate and_gate_h_u_arrmul32_and13_10_y0(a_13, b_10, h_u_arrmul32_and13_10_y0);
  fa fa_h_u_arrmul32_fa13_10_y2(h_u_arrmul32_and13_10_y0, h_u_arrmul32_fa14_9_y2, h_u_arrmul32_fa12_10_y4, h_u_arrmul32_fa13_10_y2, h_u_arrmul32_fa13_10_y4);
  and_gate and_gate_h_u_arrmul32_and14_10_y0(a_14, b_10, h_u_arrmul32_and14_10_y0);
  fa fa_h_u_arrmul32_fa14_10_y2(h_u_arrmul32_and14_10_y0, h_u_arrmul32_fa15_9_y2, h_u_arrmul32_fa13_10_y4, h_u_arrmul32_fa14_10_y2, h_u_arrmul32_fa14_10_y4);
  and_gate and_gate_h_u_arrmul32_and15_10_y0(a_15, b_10, h_u_arrmul32_and15_10_y0);
  fa fa_h_u_arrmul32_fa15_10_y2(h_u_arrmul32_and15_10_y0, h_u_arrmul32_fa16_9_y2, h_u_arrmul32_fa14_10_y4, h_u_arrmul32_fa15_10_y2, h_u_arrmul32_fa15_10_y4);
  and_gate and_gate_h_u_arrmul32_and16_10_y0(a_16, b_10, h_u_arrmul32_and16_10_y0);
  fa fa_h_u_arrmul32_fa16_10_y2(h_u_arrmul32_and16_10_y0, h_u_arrmul32_fa17_9_y2, h_u_arrmul32_fa15_10_y4, h_u_arrmul32_fa16_10_y2, h_u_arrmul32_fa16_10_y4);
  and_gate and_gate_h_u_arrmul32_and17_10_y0(a_17, b_10, h_u_arrmul32_and17_10_y0);
  fa fa_h_u_arrmul32_fa17_10_y2(h_u_arrmul32_and17_10_y0, h_u_arrmul32_fa18_9_y2, h_u_arrmul32_fa16_10_y4, h_u_arrmul32_fa17_10_y2, h_u_arrmul32_fa17_10_y4);
  and_gate and_gate_h_u_arrmul32_and18_10_y0(a_18, b_10, h_u_arrmul32_and18_10_y0);
  fa fa_h_u_arrmul32_fa18_10_y2(h_u_arrmul32_and18_10_y0, h_u_arrmul32_fa19_9_y2, h_u_arrmul32_fa17_10_y4, h_u_arrmul32_fa18_10_y2, h_u_arrmul32_fa18_10_y4);
  and_gate and_gate_h_u_arrmul32_and19_10_y0(a_19, b_10, h_u_arrmul32_and19_10_y0);
  fa fa_h_u_arrmul32_fa19_10_y2(h_u_arrmul32_and19_10_y0, h_u_arrmul32_fa20_9_y2, h_u_arrmul32_fa18_10_y4, h_u_arrmul32_fa19_10_y2, h_u_arrmul32_fa19_10_y4);
  and_gate and_gate_h_u_arrmul32_and20_10_y0(a_20, b_10, h_u_arrmul32_and20_10_y0);
  fa fa_h_u_arrmul32_fa20_10_y2(h_u_arrmul32_and20_10_y0, h_u_arrmul32_fa21_9_y2, h_u_arrmul32_fa19_10_y4, h_u_arrmul32_fa20_10_y2, h_u_arrmul32_fa20_10_y4);
  and_gate and_gate_h_u_arrmul32_and21_10_y0(a_21, b_10, h_u_arrmul32_and21_10_y0);
  fa fa_h_u_arrmul32_fa21_10_y2(h_u_arrmul32_and21_10_y0, h_u_arrmul32_fa22_9_y2, h_u_arrmul32_fa20_10_y4, h_u_arrmul32_fa21_10_y2, h_u_arrmul32_fa21_10_y4);
  and_gate and_gate_h_u_arrmul32_and22_10_y0(a_22, b_10, h_u_arrmul32_and22_10_y0);
  fa fa_h_u_arrmul32_fa22_10_y2(h_u_arrmul32_and22_10_y0, h_u_arrmul32_fa23_9_y2, h_u_arrmul32_fa21_10_y4, h_u_arrmul32_fa22_10_y2, h_u_arrmul32_fa22_10_y4);
  and_gate and_gate_h_u_arrmul32_and23_10_y0(a_23, b_10, h_u_arrmul32_and23_10_y0);
  fa fa_h_u_arrmul32_fa23_10_y2(h_u_arrmul32_and23_10_y0, h_u_arrmul32_fa24_9_y2, h_u_arrmul32_fa22_10_y4, h_u_arrmul32_fa23_10_y2, h_u_arrmul32_fa23_10_y4);
  and_gate and_gate_h_u_arrmul32_and24_10_y0(a_24, b_10, h_u_arrmul32_and24_10_y0);
  fa fa_h_u_arrmul32_fa24_10_y2(h_u_arrmul32_and24_10_y0, h_u_arrmul32_fa25_9_y2, h_u_arrmul32_fa23_10_y4, h_u_arrmul32_fa24_10_y2, h_u_arrmul32_fa24_10_y4);
  and_gate and_gate_h_u_arrmul32_and25_10_y0(a_25, b_10, h_u_arrmul32_and25_10_y0);
  fa fa_h_u_arrmul32_fa25_10_y2(h_u_arrmul32_and25_10_y0, h_u_arrmul32_fa26_9_y2, h_u_arrmul32_fa24_10_y4, h_u_arrmul32_fa25_10_y2, h_u_arrmul32_fa25_10_y4);
  and_gate and_gate_h_u_arrmul32_and26_10_y0(a_26, b_10, h_u_arrmul32_and26_10_y0);
  fa fa_h_u_arrmul32_fa26_10_y2(h_u_arrmul32_and26_10_y0, h_u_arrmul32_fa27_9_y2, h_u_arrmul32_fa25_10_y4, h_u_arrmul32_fa26_10_y2, h_u_arrmul32_fa26_10_y4);
  and_gate and_gate_h_u_arrmul32_and27_10_y0(a_27, b_10, h_u_arrmul32_and27_10_y0);
  fa fa_h_u_arrmul32_fa27_10_y2(h_u_arrmul32_and27_10_y0, h_u_arrmul32_fa28_9_y2, h_u_arrmul32_fa26_10_y4, h_u_arrmul32_fa27_10_y2, h_u_arrmul32_fa27_10_y4);
  and_gate and_gate_h_u_arrmul32_and28_10_y0(a_28, b_10, h_u_arrmul32_and28_10_y0);
  fa fa_h_u_arrmul32_fa28_10_y2(h_u_arrmul32_and28_10_y0, h_u_arrmul32_fa29_9_y2, h_u_arrmul32_fa27_10_y4, h_u_arrmul32_fa28_10_y2, h_u_arrmul32_fa28_10_y4);
  and_gate and_gate_h_u_arrmul32_and29_10_y0(a_29, b_10, h_u_arrmul32_and29_10_y0);
  fa fa_h_u_arrmul32_fa29_10_y2(h_u_arrmul32_and29_10_y0, h_u_arrmul32_fa30_9_y2, h_u_arrmul32_fa28_10_y4, h_u_arrmul32_fa29_10_y2, h_u_arrmul32_fa29_10_y4);
  and_gate and_gate_h_u_arrmul32_and30_10_y0(a_30, b_10, h_u_arrmul32_and30_10_y0);
  fa fa_h_u_arrmul32_fa30_10_y2(h_u_arrmul32_and30_10_y0, h_u_arrmul32_fa31_9_y2, h_u_arrmul32_fa29_10_y4, h_u_arrmul32_fa30_10_y2, h_u_arrmul32_fa30_10_y4);
  and_gate and_gate_h_u_arrmul32_and31_10_y0(a_31, b_10, h_u_arrmul32_and31_10_y0);
  fa fa_h_u_arrmul32_fa31_10_y2(h_u_arrmul32_and31_10_y0, h_u_arrmul32_fa31_9_y4, h_u_arrmul32_fa30_10_y4, h_u_arrmul32_fa31_10_y2, h_u_arrmul32_fa31_10_y4);
  and_gate and_gate_h_u_arrmul32_and0_11_y0(a_0, b_11, h_u_arrmul32_and0_11_y0);
  ha ha_h_u_arrmul32_ha0_11_y0(h_u_arrmul32_and0_11_y0, h_u_arrmul32_fa1_10_y2, h_u_arrmul32_ha0_11_y0, h_u_arrmul32_ha0_11_y1);
  and_gate and_gate_h_u_arrmul32_and1_11_y0(a_1, b_11, h_u_arrmul32_and1_11_y0);
  fa fa_h_u_arrmul32_fa1_11_y2(h_u_arrmul32_and1_11_y0, h_u_arrmul32_fa2_10_y2, h_u_arrmul32_ha0_11_y1, h_u_arrmul32_fa1_11_y2, h_u_arrmul32_fa1_11_y4);
  and_gate and_gate_h_u_arrmul32_and2_11_y0(a_2, b_11, h_u_arrmul32_and2_11_y0);
  fa fa_h_u_arrmul32_fa2_11_y2(h_u_arrmul32_and2_11_y0, h_u_arrmul32_fa3_10_y2, h_u_arrmul32_fa1_11_y4, h_u_arrmul32_fa2_11_y2, h_u_arrmul32_fa2_11_y4);
  and_gate and_gate_h_u_arrmul32_and3_11_y0(a_3, b_11, h_u_arrmul32_and3_11_y0);
  fa fa_h_u_arrmul32_fa3_11_y2(h_u_arrmul32_and3_11_y0, h_u_arrmul32_fa4_10_y2, h_u_arrmul32_fa2_11_y4, h_u_arrmul32_fa3_11_y2, h_u_arrmul32_fa3_11_y4);
  and_gate and_gate_h_u_arrmul32_and4_11_y0(a_4, b_11, h_u_arrmul32_and4_11_y0);
  fa fa_h_u_arrmul32_fa4_11_y2(h_u_arrmul32_and4_11_y0, h_u_arrmul32_fa5_10_y2, h_u_arrmul32_fa3_11_y4, h_u_arrmul32_fa4_11_y2, h_u_arrmul32_fa4_11_y4);
  and_gate and_gate_h_u_arrmul32_and5_11_y0(a_5, b_11, h_u_arrmul32_and5_11_y0);
  fa fa_h_u_arrmul32_fa5_11_y2(h_u_arrmul32_and5_11_y0, h_u_arrmul32_fa6_10_y2, h_u_arrmul32_fa4_11_y4, h_u_arrmul32_fa5_11_y2, h_u_arrmul32_fa5_11_y4);
  and_gate and_gate_h_u_arrmul32_and6_11_y0(a_6, b_11, h_u_arrmul32_and6_11_y0);
  fa fa_h_u_arrmul32_fa6_11_y2(h_u_arrmul32_and6_11_y0, h_u_arrmul32_fa7_10_y2, h_u_arrmul32_fa5_11_y4, h_u_arrmul32_fa6_11_y2, h_u_arrmul32_fa6_11_y4);
  and_gate and_gate_h_u_arrmul32_and7_11_y0(a_7, b_11, h_u_arrmul32_and7_11_y0);
  fa fa_h_u_arrmul32_fa7_11_y2(h_u_arrmul32_and7_11_y0, h_u_arrmul32_fa8_10_y2, h_u_arrmul32_fa6_11_y4, h_u_arrmul32_fa7_11_y2, h_u_arrmul32_fa7_11_y4);
  and_gate and_gate_h_u_arrmul32_and8_11_y0(a_8, b_11, h_u_arrmul32_and8_11_y0);
  fa fa_h_u_arrmul32_fa8_11_y2(h_u_arrmul32_and8_11_y0, h_u_arrmul32_fa9_10_y2, h_u_arrmul32_fa7_11_y4, h_u_arrmul32_fa8_11_y2, h_u_arrmul32_fa8_11_y4);
  and_gate and_gate_h_u_arrmul32_and9_11_y0(a_9, b_11, h_u_arrmul32_and9_11_y0);
  fa fa_h_u_arrmul32_fa9_11_y2(h_u_arrmul32_and9_11_y0, h_u_arrmul32_fa10_10_y2, h_u_arrmul32_fa8_11_y4, h_u_arrmul32_fa9_11_y2, h_u_arrmul32_fa9_11_y4);
  and_gate and_gate_h_u_arrmul32_and10_11_y0(a_10, b_11, h_u_arrmul32_and10_11_y0);
  fa fa_h_u_arrmul32_fa10_11_y2(h_u_arrmul32_and10_11_y0, h_u_arrmul32_fa11_10_y2, h_u_arrmul32_fa9_11_y4, h_u_arrmul32_fa10_11_y2, h_u_arrmul32_fa10_11_y4);
  and_gate and_gate_h_u_arrmul32_and11_11_y0(a_11, b_11, h_u_arrmul32_and11_11_y0);
  fa fa_h_u_arrmul32_fa11_11_y2(h_u_arrmul32_and11_11_y0, h_u_arrmul32_fa12_10_y2, h_u_arrmul32_fa10_11_y4, h_u_arrmul32_fa11_11_y2, h_u_arrmul32_fa11_11_y4);
  and_gate and_gate_h_u_arrmul32_and12_11_y0(a_12, b_11, h_u_arrmul32_and12_11_y0);
  fa fa_h_u_arrmul32_fa12_11_y2(h_u_arrmul32_and12_11_y0, h_u_arrmul32_fa13_10_y2, h_u_arrmul32_fa11_11_y4, h_u_arrmul32_fa12_11_y2, h_u_arrmul32_fa12_11_y4);
  and_gate and_gate_h_u_arrmul32_and13_11_y0(a_13, b_11, h_u_arrmul32_and13_11_y0);
  fa fa_h_u_arrmul32_fa13_11_y2(h_u_arrmul32_and13_11_y0, h_u_arrmul32_fa14_10_y2, h_u_arrmul32_fa12_11_y4, h_u_arrmul32_fa13_11_y2, h_u_arrmul32_fa13_11_y4);
  and_gate and_gate_h_u_arrmul32_and14_11_y0(a_14, b_11, h_u_arrmul32_and14_11_y0);
  fa fa_h_u_arrmul32_fa14_11_y2(h_u_arrmul32_and14_11_y0, h_u_arrmul32_fa15_10_y2, h_u_arrmul32_fa13_11_y4, h_u_arrmul32_fa14_11_y2, h_u_arrmul32_fa14_11_y4);
  and_gate and_gate_h_u_arrmul32_and15_11_y0(a_15, b_11, h_u_arrmul32_and15_11_y0);
  fa fa_h_u_arrmul32_fa15_11_y2(h_u_arrmul32_and15_11_y0, h_u_arrmul32_fa16_10_y2, h_u_arrmul32_fa14_11_y4, h_u_arrmul32_fa15_11_y2, h_u_arrmul32_fa15_11_y4);
  and_gate and_gate_h_u_arrmul32_and16_11_y0(a_16, b_11, h_u_arrmul32_and16_11_y0);
  fa fa_h_u_arrmul32_fa16_11_y2(h_u_arrmul32_and16_11_y0, h_u_arrmul32_fa17_10_y2, h_u_arrmul32_fa15_11_y4, h_u_arrmul32_fa16_11_y2, h_u_arrmul32_fa16_11_y4);
  and_gate and_gate_h_u_arrmul32_and17_11_y0(a_17, b_11, h_u_arrmul32_and17_11_y0);
  fa fa_h_u_arrmul32_fa17_11_y2(h_u_arrmul32_and17_11_y0, h_u_arrmul32_fa18_10_y2, h_u_arrmul32_fa16_11_y4, h_u_arrmul32_fa17_11_y2, h_u_arrmul32_fa17_11_y4);
  and_gate and_gate_h_u_arrmul32_and18_11_y0(a_18, b_11, h_u_arrmul32_and18_11_y0);
  fa fa_h_u_arrmul32_fa18_11_y2(h_u_arrmul32_and18_11_y0, h_u_arrmul32_fa19_10_y2, h_u_arrmul32_fa17_11_y4, h_u_arrmul32_fa18_11_y2, h_u_arrmul32_fa18_11_y4);
  and_gate and_gate_h_u_arrmul32_and19_11_y0(a_19, b_11, h_u_arrmul32_and19_11_y0);
  fa fa_h_u_arrmul32_fa19_11_y2(h_u_arrmul32_and19_11_y0, h_u_arrmul32_fa20_10_y2, h_u_arrmul32_fa18_11_y4, h_u_arrmul32_fa19_11_y2, h_u_arrmul32_fa19_11_y4);
  and_gate and_gate_h_u_arrmul32_and20_11_y0(a_20, b_11, h_u_arrmul32_and20_11_y0);
  fa fa_h_u_arrmul32_fa20_11_y2(h_u_arrmul32_and20_11_y0, h_u_arrmul32_fa21_10_y2, h_u_arrmul32_fa19_11_y4, h_u_arrmul32_fa20_11_y2, h_u_arrmul32_fa20_11_y4);
  and_gate and_gate_h_u_arrmul32_and21_11_y0(a_21, b_11, h_u_arrmul32_and21_11_y0);
  fa fa_h_u_arrmul32_fa21_11_y2(h_u_arrmul32_and21_11_y0, h_u_arrmul32_fa22_10_y2, h_u_arrmul32_fa20_11_y4, h_u_arrmul32_fa21_11_y2, h_u_arrmul32_fa21_11_y4);
  and_gate and_gate_h_u_arrmul32_and22_11_y0(a_22, b_11, h_u_arrmul32_and22_11_y0);
  fa fa_h_u_arrmul32_fa22_11_y2(h_u_arrmul32_and22_11_y0, h_u_arrmul32_fa23_10_y2, h_u_arrmul32_fa21_11_y4, h_u_arrmul32_fa22_11_y2, h_u_arrmul32_fa22_11_y4);
  and_gate and_gate_h_u_arrmul32_and23_11_y0(a_23, b_11, h_u_arrmul32_and23_11_y0);
  fa fa_h_u_arrmul32_fa23_11_y2(h_u_arrmul32_and23_11_y0, h_u_arrmul32_fa24_10_y2, h_u_arrmul32_fa22_11_y4, h_u_arrmul32_fa23_11_y2, h_u_arrmul32_fa23_11_y4);
  and_gate and_gate_h_u_arrmul32_and24_11_y0(a_24, b_11, h_u_arrmul32_and24_11_y0);
  fa fa_h_u_arrmul32_fa24_11_y2(h_u_arrmul32_and24_11_y0, h_u_arrmul32_fa25_10_y2, h_u_arrmul32_fa23_11_y4, h_u_arrmul32_fa24_11_y2, h_u_arrmul32_fa24_11_y4);
  and_gate and_gate_h_u_arrmul32_and25_11_y0(a_25, b_11, h_u_arrmul32_and25_11_y0);
  fa fa_h_u_arrmul32_fa25_11_y2(h_u_arrmul32_and25_11_y0, h_u_arrmul32_fa26_10_y2, h_u_arrmul32_fa24_11_y4, h_u_arrmul32_fa25_11_y2, h_u_arrmul32_fa25_11_y4);
  and_gate and_gate_h_u_arrmul32_and26_11_y0(a_26, b_11, h_u_arrmul32_and26_11_y0);
  fa fa_h_u_arrmul32_fa26_11_y2(h_u_arrmul32_and26_11_y0, h_u_arrmul32_fa27_10_y2, h_u_arrmul32_fa25_11_y4, h_u_arrmul32_fa26_11_y2, h_u_arrmul32_fa26_11_y4);
  and_gate and_gate_h_u_arrmul32_and27_11_y0(a_27, b_11, h_u_arrmul32_and27_11_y0);
  fa fa_h_u_arrmul32_fa27_11_y2(h_u_arrmul32_and27_11_y0, h_u_arrmul32_fa28_10_y2, h_u_arrmul32_fa26_11_y4, h_u_arrmul32_fa27_11_y2, h_u_arrmul32_fa27_11_y4);
  and_gate and_gate_h_u_arrmul32_and28_11_y0(a_28, b_11, h_u_arrmul32_and28_11_y0);
  fa fa_h_u_arrmul32_fa28_11_y2(h_u_arrmul32_and28_11_y0, h_u_arrmul32_fa29_10_y2, h_u_arrmul32_fa27_11_y4, h_u_arrmul32_fa28_11_y2, h_u_arrmul32_fa28_11_y4);
  and_gate and_gate_h_u_arrmul32_and29_11_y0(a_29, b_11, h_u_arrmul32_and29_11_y0);
  fa fa_h_u_arrmul32_fa29_11_y2(h_u_arrmul32_and29_11_y0, h_u_arrmul32_fa30_10_y2, h_u_arrmul32_fa28_11_y4, h_u_arrmul32_fa29_11_y2, h_u_arrmul32_fa29_11_y4);
  and_gate and_gate_h_u_arrmul32_and30_11_y0(a_30, b_11, h_u_arrmul32_and30_11_y0);
  fa fa_h_u_arrmul32_fa30_11_y2(h_u_arrmul32_and30_11_y0, h_u_arrmul32_fa31_10_y2, h_u_arrmul32_fa29_11_y4, h_u_arrmul32_fa30_11_y2, h_u_arrmul32_fa30_11_y4);
  and_gate and_gate_h_u_arrmul32_and31_11_y0(a_31, b_11, h_u_arrmul32_and31_11_y0);
  fa fa_h_u_arrmul32_fa31_11_y2(h_u_arrmul32_and31_11_y0, h_u_arrmul32_fa31_10_y4, h_u_arrmul32_fa30_11_y4, h_u_arrmul32_fa31_11_y2, h_u_arrmul32_fa31_11_y4);
  and_gate and_gate_h_u_arrmul32_and0_12_y0(a_0, b_12, h_u_arrmul32_and0_12_y0);
  ha ha_h_u_arrmul32_ha0_12_y0(h_u_arrmul32_and0_12_y0, h_u_arrmul32_fa1_11_y2, h_u_arrmul32_ha0_12_y0, h_u_arrmul32_ha0_12_y1);
  and_gate and_gate_h_u_arrmul32_and1_12_y0(a_1, b_12, h_u_arrmul32_and1_12_y0);
  fa fa_h_u_arrmul32_fa1_12_y2(h_u_arrmul32_and1_12_y0, h_u_arrmul32_fa2_11_y2, h_u_arrmul32_ha0_12_y1, h_u_arrmul32_fa1_12_y2, h_u_arrmul32_fa1_12_y4);
  and_gate and_gate_h_u_arrmul32_and2_12_y0(a_2, b_12, h_u_arrmul32_and2_12_y0);
  fa fa_h_u_arrmul32_fa2_12_y2(h_u_arrmul32_and2_12_y0, h_u_arrmul32_fa3_11_y2, h_u_arrmul32_fa1_12_y4, h_u_arrmul32_fa2_12_y2, h_u_arrmul32_fa2_12_y4);
  and_gate and_gate_h_u_arrmul32_and3_12_y0(a_3, b_12, h_u_arrmul32_and3_12_y0);
  fa fa_h_u_arrmul32_fa3_12_y2(h_u_arrmul32_and3_12_y0, h_u_arrmul32_fa4_11_y2, h_u_arrmul32_fa2_12_y4, h_u_arrmul32_fa3_12_y2, h_u_arrmul32_fa3_12_y4);
  and_gate and_gate_h_u_arrmul32_and4_12_y0(a_4, b_12, h_u_arrmul32_and4_12_y0);
  fa fa_h_u_arrmul32_fa4_12_y2(h_u_arrmul32_and4_12_y0, h_u_arrmul32_fa5_11_y2, h_u_arrmul32_fa3_12_y4, h_u_arrmul32_fa4_12_y2, h_u_arrmul32_fa4_12_y4);
  and_gate and_gate_h_u_arrmul32_and5_12_y0(a_5, b_12, h_u_arrmul32_and5_12_y0);
  fa fa_h_u_arrmul32_fa5_12_y2(h_u_arrmul32_and5_12_y0, h_u_arrmul32_fa6_11_y2, h_u_arrmul32_fa4_12_y4, h_u_arrmul32_fa5_12_y2, h_u_arrmul32_fa5_12_y4);
  and_gate and_gate_h_u_arrmul32_and6_12_y0(a_6, b_12, h_u_arrmul32_and6_12_y0);
  fa fa_h_u_arrmul32_fa6_12_y2(h_u_arrmul32_and6_12_y0, h_u_arrmul32_fa7_11_y2, h_u_arrmul32_fa5_12_y4, h_u_arrmul32_fa6_12_y2, h_u_arrmul32_fa6_12_y4);
  and_gate and_gate_h_u_arrmul32_and7_12_y0(a_7, b_12, h_u_arrmul32_and7_12_y0);
  fa fa_h_u_arrmul32_fa7_12_y2(h_u_arrmul32_and7_12_y0, h_u_arrmul32_fa8_11_y2, h_u_arrmul32_fa6_12_y4, h_u_arrmul32_fa7_12_y2, h_u_arrmul32_fa7_12_y4);
  and_gate and_gate_h_u_arrmul32_and8_12_y0(a_8, b_12, h_u_arrmul32_and8_12_y0);
  fa fa_h_u_arrmul32_fa8_12_y2(h_u_arrmul32_and8_12_y0, h_u_arrmul32_fa9_11_y2, h_u_arrmul32_fa7_12_y4, h_u_arrmul32_fa8_12_y2, h_u_arrmul32_fa8_12_y4);
  and_gate and_gate_h_u_arrmul32_and9_12_y0(a_9, b_12, h_u_arrmul32_and9_12_y0);
  fa fa_h_u_arrmul32_fa9_12_y2(h_u_arrmul32_and9_12_y0, h_u_arrmul32_fa10_11_y2, h_u_arrmul32_fa8_12_y4, h_u_arrmul32_fa9_12_y2, h_u_arrmul32_fa9_12_y4);
  and_gate and_gate_h_u_arrmul32_and10_12_y0(a_10, b_12, h_u_arrmul32_and10_12_y0);
  fa fa_h_u_arrmul32_fa10_12_y2(h_u_arrmul32_and10_12_y0, h_u_arrmul32_fa11_11_y2, h_u_arrmul32_fa9_12_y4, h_u_arrmul32_fa10_12_y2, h_u_arrmul32_fa10_12_y4);
  and_gate and_gate_h_u_arrmul32_and11_12_y0(a_11, b_12, h_u_arrmul32_and11_12_y0);
  fa fa_h_u_arrmul32_fa11_12_y2(h_u_arrmul32_and11_12_y0, h_u_arrmul32_fa12_11_y2, h_u_arrmul32_fa10_12_y4, h_u_arrmul32_fa11_12_y2, h_u_arrmul32_fa11_12_y4);
  and_gate and_gate_h_u_arrmul32_and12_12_y0(a_12, b_12, h_u_arrmul32_and12_12_y0);
  fa fa_h_u_arrmul32_fa12_12_y2(h_u_arrmul32_and12_12_y0, h_u_arrmul32_fa13_11_y2, h_u_arrmul32_fa11_12_y4, h_u_arrmul32_fa12_12_y2, h_u_arrmul32_fa12_12_y4);
  and_gate and_gate_h_u_arrmul32_and13_12_y0(a_13, b_12, h_u_arrmul32_and13_12_y0);
  fa fa_h_u_arrmul32_fa13_12_y2(h_u_arrmul32_and13_12_y0, h_u_arrmul32_fa14_11_y2, h_u_arrmul32_fa12_12_y4, h_u_arrmul32_fa13_12_y2, h_u_arrmul32_fa13_12_y4);
  and_gate and_gate_h_u_arrmul32_and14_12_y0(a_14, b_12, h_u_arrmul32_and14_12_y0);
  fa fa_h_u_arrmul32_fa14_12_y2(h_u_arrmul32_and14_12_y0, h_u_arrmul32_fa15_11_y2, h_u_arrmul32_fa13_12_y4, h_u_arrmul32_fa14_12_y2, h_u_arrmul32_fa14_12_y4);
  and_gate and_gate_h_u_arrmul32_and15_12_y0(a_15, b_12, h_u_arrmul32_and15_12_y0);
  fa fa_h_u_arrmul32_fa15_12_y2(h_u_arrmul32_and15_12_y0, h_u_arrmul32_fa16_11_y2, h_u_arrmul32_fa14_12_y4, h_u_arrmul32_fa15_12_y2, h_u_arrmul32_fa15_12_y4);
  and_gate and_gate_h_u_arrmul32_and16_12_y0(a_16, b_12, h_u_arrmul32_and16_12_y0);
  fa fa_h_u_arrmul32_fa16_12_y2(h_u_arrmul32_and16_12_y0, h_u_arrmul32_fa17_11_y2, h_u_arrmul32_fa15_12_y4, h_u_arrmul32_fa16_12_y2, h_u_arrmul32_fa16_12_y4);
  and_gate and_gate_h_u_arrmul32_and17_12_y0(a_17, b_12, h_u_arrmul32_and17_12_y0);
  fa fa_h_u_arrmul32_fa17_12_y2(h_u_arrmul32_and17_12_y0, h_u_arrmul32_fa18_11_y2, h_u_arrmul32_fa16_12_y4, h_u_arrmul32_fa17_12_y2, h_u_arrmul32_fa17_12_y4);
  and_gate and_gate_h_u_arrmul32_and18_12_y0(a_18, b_12, h_u_arrmul32_and18_12_y0);
  fa fa_h_u_arrmul32_fa18_12_y2(h_u_arrmul32_and18_12_y0, h_u_arrmul32_fa19_11_y2, h_u_arrmul32_fa17_12_y4, h_u_arrmul32_fa18_12_y2, h_u_arrmul32_fa18_12_y4);
  and_gate and_gate_h_u_arrmul32_and19_12_y0(a_19, b_12, h_u_arrmul32_and19_12_y0);
  fa fa_h_u_arrmul32_fa19_12_y2(h_u_arrmul32_and19_12_y0, h_u_arrmul32_fa20_11_y2, h_u_arrmul32_fa18_12_y4, h_u_arrmul32_fa19_12_y2, h_u_arrmul32_fa19_12_y4);
  and_gate and_gate_h_u_arrmul32_and20_12_y0(a_20, b_12, h_u_arrmul32_and20_12_y0);
  fa fa_h_u_arrmul32_fa20_12_y2(h_u_arrmul32_and20_12_y0, h_u_arrmul32_fa21_11_y2, h_u_arrmul32_fa19_12_y4, h_u_arrmul32_fa20_12_y2, h_u_arrmul32_fa20_12_y4);
  and_gate and_gate_h_u_arrmul32_and21_12_y0(a_21, b_12, h_u_arrmul32_and21_12_y0);
  fa fa_h_u_arrmul32_fa21_12_y2(h_u_arrmul32_and21_12_y0, h_u_arrmul32_fa22_11_y2, h_u_arrmul32_fa20_12_y4, h_u_arrmul32_fa21_12_y2, h_u_arrmul32_fa21_12_y4);
  and_gate and_gate_h_u_arrmul32_and22_12_y0(a_22, b_12, h_u_arrmul32_and22_12_y0);
  fa fa_h_u_arrmul32_fa22_12_y2(h_u_arrmul32_and22_12_y0, h_u_arrmul32_fa23_11_y2, h_u_arrmul32_fa21_12_y4, h_u_arrmul32_fa22_12_y2, h_u_arrmul32_fa22_12_y4);
  and_gate and_gate_h_u_arrmul32_and23_12_y0(a_23, b_12, h_u_arrmul32_and23_12_y0);
  fa fa_h_u_arrmul32_fa23_12_y2(h_u_arrmul32_and23_12_y0, h_u_arrmul32_fa24_11_y2, h_u_arrmul32_fa22_12_y4, h_u_arrmul32_fa23_12_y2, h_u_arrmul32_fa23_12_y4);
  and_gate and_gate_h_u_arrmul32_and24_12_y0(a_24, b_12, h_u_arrmul32_and24_12_y0);
  fa fa_h_u_arrmul32_fa24_12_y2(h_u_arrmul32_and24_12_y0, h_u_arrmul32_fa25_11_y2, h_u_arrmul32_fa23_12_y4, h_u_arrmul32_fa24_12_y2, h_u_arrmul32_fa24_12_y4);
  and_gate and_gate_h_u_arrmul32_and25_12_y0(a_25, b_12, h_u_arrmul32_and25_12_y0);
  fa fa_h_u_arrmul32_fa25_12_y2(h_u_arrmul32_and25_12_y0, h_u_arrmul32_fa26_11_y2, h_u_arrmul32_fa24_12_y4, h_u_arrmul32_fa25_12_y2, h_u_arrmul32_fa25_12_y4);
  and_gate and_gate_h_u_arrmul32_and26_12_y0(a_26, b_12, h_u_arrmul32_and26_12_y0);
  fa fa_h_u_arrmul32_fa26_12_y2(h_u_arrmul32_and26_12_y0, h_u_arrmul32_fa27_11_y2, h_u_arrmul32_fa25_12_y4, h_u_arrmul32_fa26_12_y2, h_u_arrmul32_fa26_12_y4);
  and_gate and_gate_h_u_arrmul32_and27_12_y0(a_27, b_12, h_u_arrmul32_and27_12_y0);
  fa fa_h_u_arrmul32_fa27_12_y2(h_u_arrmul32_and27_12_y0, h_u_arrmul32_fa28_11_y2, h_u_arrmul32_fa26_12_y4, h_u_arrmul32_fa27_12_y2, h_u_arrmul32_fa27_12_y4);
  and_gate and_gate_h_u_arrmul32_and28_12_y0(a_28, b_12, h_u_arrmul32_and28_12_y0);
  fa fa_h_u_arrmul32_fa28_12_y2(h_u_arrmul32_and28_12_y0, h_u_arrmul32_fa29_11_y2, h_u_arrmul32_fa27_12_y4, h_u_arrmul32_fa28_12_y2, h_u_arrmul32_fa28_12_y4);
  and_gate and_gate_h_u_arrmul32_and29_12_y0(a_29, b_12, h_u_arrmul32_and29_12_y0);
  fa fa_h_u_arrmul32_fa29_12_y2(h_u_arrmul32_and29_12_y0, h_u_arrmul32_fa30_11_y2, h_u_arrmul32_fa28_12_y4, h_u_arrmul32_fa29_12_y2, h_u_arrmul32_fa29_12_y4);
  and_gate and_gate_h_u_arrmul32_and30_12_y0(a_30, b_12, h_u_arrmul32_and30_12_y0);
  fa fa_h_u_arrmul32_fa30_12_y2(h_u_arrmul32_and30_12_y0, h_u_arrmul32_fa31_11_y2, h_u_arrmul32_fa29_12_y4, h_u_arrmul32_fa30_12_y2, h_u_arrmul32_fa30_12_y4);
  and_gate and_gate_h_u_arrmul32_and31_12_y0(a_31, b_12, h_u_arrmul32_and31_12_y0);
  fa fa_h_u_arrmul32_fa31_12_y2(h_u_arrmul32_and31_12_y0, h_u_arrmul32_fa31_11_y4, h_u_arrmul32_fa30_12_y4, h_u_arrmul32_fa31_12_y2, h_u_arrmul32_fa31_12_y4);
  and_gate and_gate_h_u_arrmul32_and0_13_y0(a_0, b_13, h_u_arrmul32_and0_13_y0);
  ha ha_h_u_arrmul32_ha0_13_y0(h_u_arrmul32_and0_13_y0, h_u_arrmul32_fa1_12_y2, h_u_arrmul32_ha0_13_y0, h_u_arrmul32_ha0_13_y1);
  and_gate and_gate_h_u_arrmul32_and1_13_y0(a_1, b_13, h_u_arrmul32_and1_13_y0);
  fa fa_h_u_arrmul32_fa1_13_y2(h_u_arrmul32_and1_13_y0, h_u_arrmul32_fa2_12_y2, h_u_arrmul32_ha0_13_y1, h_u_arrmul32_fa1_13_y2, h_u_arrmul32_fa1_13_y4);
  and_gate and_gate_h_u_arrmul32_and2_13_y0(a_2, b_13, h_u_arrmul32_and2_13_y0);
  fa fa_h_u_arrmul32_fa2_13_y2(h_u_arrmul32_and2_13_y0, h_u_arrmul32_fa3_12_y2, h_u_arrmul32_fa1_13_y4, h_u_arrmul32_fa2_13_y2, h_u_arrmul32_fa2_13_y4);
  and_gate and_gate_h_u_arrmul32_and3_13_y0(a_3, b_13, h_u_arrmul32_and3_13_y0);
  fa fa_h_u_arrmul32_fa3_13_y2(h_u_arrmul32_and3_13_y0, h_u_arrmul32_fa4_12_y2, h_u_arrmul32_fa2_13_y4, h_u_arrmul32_fa3_13_y2, h_u_arrmul32_fa3_13_y4);
  and_gate and_gate_h_u_arrmul32_and4_13_y0(a_4, b_13, h_u_arrmul32_and4_13_y0);
  fa fa_h_u_arrmul32_fa4_13_y2(h_u_arrmul32_and4_13_y0, h_u_arrmul32_fa5_12_y2, h_u_arrmul32_fa3_13_y4, h_u_arrmul32_fa4_13_y2, h_u_arrmul32_fa4_13_y4);
  and_gate and_gate_h_u_arrmul32_and5_13_y0(a_5, b_13, h_u_arrmul32_and5_13_y0);
  fa fa_h_u_arrmul32_fa5_13_y2(h_u_arrmul32_and5_13_y0, h_u_arrmul32_fa6_12_y2, h_u_arrmul32_fa4_13_y4, h_u_arrmul32_fa5_13_y2, h_u_arrmul32_fa5_13_y4);
  and_gate and_gate_h_u_arrmul32_and6_13_y0(a_6, b_13, h_u_arrmul32_and6_13_y0);
  fa fa_h_u_arrmul32_fa6_13_y2(h_u_arrmul32_and6_13_y0, h_u_arrmul32_fa7_12_y2, h_u_arrmul32_fa5_13_y4, h_u_arrmul32_fa6_13_y2, h_u_arrmul32_fa6_13_y4);
  and_gate and_gate_h_u_arrmul32_and7_13_y0(a_7, b_13, h_u_arrmul32_and7_13_y0);
  fa fa_h_u_arrmul32_fa7_13_y2(h_u_arrmul32_and7_13_y0, h_u_arrmul32_fa8_12_y2, h_u_arrmul32_fa6_13_y4, h_u_arrmul32_fa7_13_y2, h_u_arrmul32_fa7_13_y4);
  and_gate and_gate_h_u_arrmul32_and8_13_y0(a_8, b_13, h_u_arrmul32_and8_13_y0);
  fa fa_h_u_arrmul32_fa8_13_y2(h_u_arrmul32_and8_13_y0, h_u_arrmul32_fa9_12_y2, h_u_arrmul32_fa7_13_y4, h_u_arrmul32_fa8_13_y2, h_u_arrmul32_fa8_13_y4);
  and_gate and_gate_h_u_arrmul32_and9_13_y0(a_9, b_13, h_u_arrmul32_and9_13_y0);
  fa fa_h_u_arrmul32_fa9_13_y2(h_u_arrmul32_and9_13_y0, h_u_arrmul32_fa10_12_y2, h_u_arrmul32_fa8_13_y4, h_u_arrmul32_fa9_13_y2, h_u_arrmul32_fa9_13_y4);
  and_gate and_gate_h_u_arrmul32_and10_13_y0(a_10, b_13, h_u_arrmul32_and10_13_y0);
  fa fa_h_u_arrmul32_fa10_13_y2(h_u_arrmul32_and10_13_y0, h_u_arrmul32_fa11_12_y2, h_u_arrmul32_fa9_13_y4, h_u_arrmul32_fa10_13_y2, h_u_arrmul32_fa10_13_y4);
  and_gate and_gate_h_u_arrmul32_and11_13_y0(a_11, b_13, h_u_arrmul32_and11_13_y0);
  fa fa_h_u_arrmul32_fa11_13_y2(h_u_arrmul32_and11_13_y0, h_u_arrmul32_fa12_12_y2, h_u_arrmul32_fa10_13_y4, h_u_arrmul32_fa11_13_y2, h_u_arrmul32_fa11_13_y4);
  and_gate and_gate_h_u_arrmul32_and12_13_y0(a_12, b_13, h_u_arrmul32_and12_13_y0);
  fa fa_h_u_arrmul32_fa12_13_y2(h_u_arrmul32_and12_13_y0, h_u_arrmul32_fa13_12_y2, h_u_arrmul32_fa11_13_y4, h_u_arrmul32_fa12_13_y2, h_u_arrmul32_fa12_13_y4);
  and_gate and_gate_h_u_arrmul32_and13_13_y0(a_13, b_13, h_u_arrmul32_and13_13_y0);
  fa fa_h_u_arrmul32_fa13_13_y2(h_u_arrmul32_and13_13_y0, h_u_arrmul32_fa14_12_y2, h_u_arrmul32_fa12_13_y4, h_u_arrmul32_fa13_13_y2, h_u_arrmul32_fa13_13_y4);
  and_gate and_gate_h_u_arrmul32_and14_13_y0(a_14, b_13, h_u_arrmul32_and14_13_y0);
  fa fa_h_u_arrmul32_fa14_13_y2(h_u_arrmul32_and14_13_y0, h_u_arrmul32_fa15_12_y2, h_u_arrmul32_fa13_13_y4, h_u_arrmul32_fa14_13_y2, h_u_arrmul32_fa14_13_y4);
  and_gate and_gate_h_u_arrmul32_and15_13_y0(a_15, b_13, h_u_arrmul32_and15_13_y0);
  fa fa_h_u_arrmul32_fa15_13_y2(h_u_arrmul32_and15_13_y0, h_u_arrmul32_fa16_12_y2, h_u_arrmul32_fa14_13_y4, h_u_arrmul32_fa15_13_y2, h_u_arrmul32_fa15_13_y4);
  and_gate and_gate_h_u_arrmul32_and16_13_y0(a_16, b_13, h_u_arrmul32_and16_13_y0);
  fa fa_h_u_arrmul32_fa16_13_y2(h_u_arrmul32_and16_13_y0, h_u_arrmul32_fa17_12_y2, h_u_arrmul32_fa15_13_y4, h_u_arrmul32_fa16_13_y2, h_u_arrmul32_fa16_13_y4);
  and_gate and_gate_h_u_arrmul32_and17_13_y0(a_17, b_13, h_u_arrmul32_and17_13_y0);
  fa fa_h_u_arrmul32_fa17_13_y2(h_u_arrmul32_and17_13_y0, h_u_arrmul32_fa18_12_y2, h_u_arrmul32_fa16_13_y4, h_u_arrmul32_fa17_13_y2, h_u_arrmul32_fa17_13_y4);
  and_gate and_gate_h_u_arrmul32_and18_13_y0(a_18, b_13, h_u_arrmul32_and18_13_y0);
  fa fa_h_u_arrmul32_fa18_13_y2(h_u_arrmul32_and18_13_y0, h_u_arrmul32_fa19_12_y2, h_u_arrmul32_fa17_13_y4, h_u_arrmul32_fa18_13_y2, h_u_arrmul32_fa18_13_y4);
  and_gate and_gate_h_u_arrmul32_and19_13_y0(a_19, b_13, h_u_arrmul32_and19_13_y0);
  fa fa_h_u_arrmul32_fa19_13_y2(h_u_arrmul32_and19_13_y0, h_u_arrmul32_fa20_12_y2, h_u_arrmul32_fa18_13_y4, h_u_arrmul32_fa19_13_y2, h_u_arrmul32_fa19_13_y4);
  and_gate and_gate_h_u_arrmul32_and20_13_y0(a_20, b_13, h_u_arrmul32_and20_13_y0);
  fa fa_h_u_arrmul32_fa20_13_y2(h_u_arrmul32_and20_13_y0, h_u_arrmul32_fa21_12_y2, h_u_arrmul32_fa19_13_y4, h_u_arrmul32_fa20_13_y2, h_u_arrmul32_fa20_13_y4);
  and_gate and_gate_h_u_arrmul32_and21_13_y0(a_21, b_13, h_u_arrmul32_and21_13_y0);
  fa fa_h_u_arrmul32_fa21_13_y2(h_u_arrmul32_and21_13_y0, h_u_arrmul32_fa22_12_y2, h_u_arrmul32_fa20_13_y4, h_u_arrmul32_fa21_13_y2, h_u_arrmul32_fa21_13_y4);
  and_gate and_gate_h_u_arrmul32_and22_13_y0(a_22, b_13, h_u_arrmul32_and22_13_y0);
  fa fa_h_u_arrmul32_fa22_13_y2(h_u_arrmul32_and22_13_y0, h_u_arrmul32_fa23_12_y2, h_u_arrmul32_fa21_13_y4, h_u_arrmul32_fa22_13_y2, h_u_arrmul32_fa22_13_y4);
  and_gate and_gate_h_u_arrmul32_and23_13_y0(a_23, b_13, h_u_arrmul32_and23_13_y0);
  fa fa_h_u_arrmul32_fa23_13_y2(h_u_arrmul32_and23_13_y0, h_u_arrmul32_fa24_12_y2, h_u_arrmul32_fa22_13_y4, h_u_arrmul32_fa23_13_y2, h_u_arrmul32_fa23_13_y4);
  and_gate and_gate_h_u_arrmul32_and24_13_y0(a_24, b_13, h_u_arrmul32_and24_13_y0);
  fa fa_h_u_arrmul32_fa24_13_y2(h_u_arrmul32_and24_13_y0, h_u_arrmul32_fa25_12_y2, h_u_arrmul32_fa23_13_y4, h_u_arrmul32_fa24_13_y2, h_u_arrmul32_fa24_13_y4);
  and_gate and_gate_h_u_arrmul32_and25_13_y0(a_25, b_13, h_u_arrmul32_and25_13_y0);
  fa fa_h_u_arrmul32_fa25_13_y2(h_u_arrmul32_and25_13_y0, h_u_arrmul32_fa26_12_y2, h_u_arrmul32_fa24_13_y4, h_u_arrmul32_fa25_13_y2, h_u_arrmul32_fa25_13_y4);
  and_gate and_gate_h_u_arrmul32_and26_13_y0(a_26, b_13, h_u_arrmul32_and26_13_y0);
  fa fa_h_u_arrmul32_fa26_13_y2(h_u_arrmul32_and26_13_y0, h_u_arrmul32_fa27_12_y2, h_u_arrmul32_fa25_13_y4, h_u_arrmul32_fa26_13_y2, h_u_arrmul32_fa26_13_y4);
  and_gate and_gate_h_u_arrmul32_and27_13_y0(a_27, b_13, h_u_arrmul32_and27_13_y0);
  fa fa_h_u_arrmul32_fa27_13_y2(h_u_arrmul32_and27_13_y0, h_u_arrmul32_fa28_12_y2, h_u_arrmul32_fa26_13_y4, h_u_arrmul32_fa27_13_y2, h_u_arrmul32_fa27_13_y4);
  and_gate and_gate_h_u_arrmul32_and28_13_y0(a_28, b_13, h_u_arrmul32_and28_13_y0);
  fa fa_h_u_arrmul32_fa28_13_y2(h_u_arrmul32_and28_13_y0, h_u_arrmul32_fa29_12_y2, h_u_arrmul32_fa27_13_y4, h_u_arrmul32_fa28_13_y2, h_u_arrmul32_fa28_13_y4);
  and_gate and_gate_h_u_arrmul32_and29_13_y0(a_29, b_13, h_u_arrmul32_and29_13_y0);
  fa fa_h_u_arrmul32_fa29_13_y2(h_u_arrmul32_and29_13_y0, h_u_arrmul32_fa30_12_y2, h_u_arrmul32_fa28_13_y4, h_u_arrmul32_fa29_13_y2, h_u_arrmul32_fa29_13_y4);
  and_gate and_gate_h_u_arrmul32_and30_13_y0(a_30, b_13, h_u_arrmul32_and30_13_y0);
  fa fa_h_u_arrmul32_fa30_13_y2(h_u_arrmul32_and30_13_y0, h_u_arrmul32_fa31_12_y2, h_u_arrmul32_fa29_13_y4, h_u_arrmul32_fa30_13_y2, h_u_arrmul32_fa30_13_y4);
  and_gate and_gate_h_u_arrmul32_and31_13_y0(a_31, b_13, h_u_arrmul32_and31_13_y0);
  fa fa_h_u_arrmul32_fa31_13_y2(h_u_arrmul32_and31_13_y0, h_u_arrmul32_fa31_12_y4, h_u_arrmul32_fa30_13_y4, h_u_arrmul32_fa31_13_y2, h_u_arrmul32_fa31_13_y4);
  and_gate and_gate_h_u_arrmul32_and0_14_y0(a_0, b_14, h_u_arrmul32_and0_14_y0);
  ha ha_h_u_arrmul32_ha0_14_y0(h_u_arrmul32_and0_14_y0, h_u_arrmul32_fa1_13_y2, h_u_arrmul32_ha0_14_y0, h_u_arrmul32_ha0_14_y1);
  and_gate and_gate_h_u_arrmul32_and1_14_y0(a_1, b_14, h_u_arrmul32_and1_14_y0);
  fa fa_h_u_arrmul32_fa1_14_y2(h_u_arrmul32_and1_14_y0, h_u_arrmul32_fa2_13_y2, h_u_arrmul32_ha0_14_y1, h_u_arrmul32_fa1_14_y2, h_u_arrmul32_fa1_14_y4);
  and_gate and_gate_h_u_arrmul32_and2_14_y0(a_2, b_14, h_u_arrmul32_and2_14_y0);
  fa fa_h_u_arrmul32_fa2_14_y2(h_u_arrmul32_and2_14_y0, h_u_arrmul32_fa3_13_y2, h_u_arrmul32_fa1_14_y4, h_u_arrmul32_fa2_14_y2, h_u_arrmul32_fa2_14_y4);
  and_gate and_gate_h_u_arrmul32_and3_14_y0(a_3, b_14, h_u_arrmul32_and3_14_y0);
  fa fa_h_u_arrmul32_fa3_14_y2(h_u_arrmul32_and3_14_y0, h_u_arrmul32_fa4_13_y2, h_u_arrmul32_fa2_14_y4, h_u_arrmul32_fa3_14_y2, h_u_arrmul32_fa3_14_y4);
  and_gate and_gate_h_u_arrmul32_and4_14_y0(a_4, b_14, h_u_arrmul32_and4_14_y0);
  fa fa_h_u_arrmul32_fa4_14_y2(h_u_arrmul32_and4_14_y0, h_u_arrmul32_fa5_13_y2, h_u_arrmul32_fa3_14_y4, h_u_arrmul32_fa4_14_y2, h_u_arrmul32_fa4_14_y4);
  and_gate and_gate_h_u_arrmul32_and5_14_y0(a_5, b_14, h_u_arrmul32_and5_14_y0);
  fa fa_h_u_arrmul32_fa5_14_y2(h_u_arrmul32_and5_14_y0, h_u_arrmul32_fa6_13_y2, h_u_arrmul32_fa4_14_y4, h_u_arrmul32_fa5_14_y2, h_u_arrmul32_fa5_14_y4);
  and_gate and_gate_h_u_arrmul32_and6_14_y0(a_6, b_14, h_u_arrmul32_and6_14_y0);
  fa fa_h_u_arrmul32_fa6_14_y2(h_u_arrmul32_and6_14_y0, h_u_arrmul32_fa7_13_y2, h_u_arrmul32_fa5_14_y4, h_u_arrmul32_fa6_14_y2, h_u_arrmul32_fa6_14_y4);
  and_gate and_gate_h_u_arrmul32_and7_14_y0(a_7, b_14, h_u_arrmul32_and7_14_y0);
  fa fa_h_u_arrmul32_fa7_14_y2(h_u_arrmul32_and7_14_y0, h_u_arrmul32_fa8_13_y2, h_u_arrmul32_fa6_14_y4, h_u_arrmul32_fa7_14_y2, h_u_arrmul32_fa7_14_y4);
  and_gate and_gate_h_u_arrmul32_and8_14_y0(a_8, b_14, h_u_arrmul32_and8_14_y0);
  fa fa_h_u_arrmul32_fa8_14_y2(h_u_arrmul32_and8_14_y0, h_u_arrmul32_fa9_13_y2, h_u_arrmul32_fa7_14_y4, h_u_arrmul32_fa8_14_y2, h_u_arrmul32_fa8_14_y4);
  and_gate and_gate_h_u_arrmul32_and9_14_y0(a_9, b_14, h_u_arrmul32_and9_14_y0);
  fa fa_h_u_arrmul32_fa9_14_y2(h_u_arrmul32_and9_14_y0, h_u_arrmul32_fa10_13_y2, h_u_arrmul32_fa8_14_y4, h_u_arrmul32_fa9_14_y2, h_u_arrmul32_fa9_14_y4);
  and_gate and_gate_h_u_arrmul32_and10_14_y0(a_10, b_14, h_u_arrmul32_and10_14_y0);
  fa fa_h_u_arrmul32_fa10_14_y2(h_u_arrmul32_and10_14_y0, h_u_arrmul32_fa11_13_y2, h_u_arrmul32_fa9_14_y4, h_u_arrmul32_fa10_14_y2, h_u_arrmul32_fa10_14_y4);
  and_gate and_gate_h_u_arrmul32_and11_14_y0(a_11, b_14, h_u_arrmul32_and11_14_y0);
  fa fa_h_u_arrmul32_fa11_14_y2(h_u_arrmul32_and11_14_y0, h_u_arrmul32_fa12_13_y2, h_u_arrmul32_fa10_14_y4, h_u_arrmul32_fa11_14_y2, h_u_arrmul32_fa11_14_y4);
  and_gate and_gate_h_u_arrmul32_and12_14_y0(a_12, b_14, h_u_arrmul32_and12_14_y0);
  fa fa_h_u_arrmul32_fa12_14_y2(h_u_arrmul32_and12_14_y0, h_u_arrmul32_fa13_13_y2, h_u_arrmul32_fa11_14_y4, h_u_arrmul32_fa12_14_y2, h_u_arrmul32_fa12_14_y4);
  and_gate and_gate_h_u_arrmul32_and13_14_y0(a_13, b_14, h_u_arrmul32_and13_14_y0);
  fa fa_h_u_arrmul32_fa13_14_y2(h_u_arrmul32_and13_14_y0, h_u_arrmul32_fa14_13_y2, h_u_arrmul32_fa12_14_y4, h_u_arrmul32_fa13_14_y2, h_u_arrmul32_fa13_14_y4);
  and_gate and_gate_h_u_arrmul32_and14_14_y0(a_14, b_14, h_u_arrmul32_and14_14_y0);
  fa fa_h_u_arrmul32_fa14_14_y2(h_u_arrmul32_and14_14_y0, h_u_arrmul32_fa15_13_y2, h_u_arrmul32_fa13_14_y4, h_u_arrmul32_fa14_14_y2, h_u_arrmul32_fa14_14_y4);
  and_gate and_gate_h_u_arrmul32_and15_14_y0(a_15, b_14, h_u_arrmul32_and15_14_y0);
  fa fa_h_u_arrmul32_fa15_14_y2(h_u_arrmul32_and15_14_y0, h_u_arrmul32_fa16_13_y2, h_u_arrmul32_fa14_14_y4, h_u_arrmul32_fa15_14_y2, h_u_arrmul32_fa15_14_y4);
  and_gate and_gate_h_u_arrmul32_and16_14_y0(a_16, b_14, h_u_arrmul32_and16_14_y0);
  fa fa_h_u_arrmul32_fa16_14_y2(h_u_arrmul32_and16_14_y0, h_u_arrmul32_fa17_13_y2, h_u_arrmul32_fa15_14_y4, h_u_arrmul32_fa16_14_y2, h_u_arrmul32_fa16_14_y4);
  and_gate and_gate_h_u_arrmul32_and17_14_y0(a_17, b_14, h_u_arrmul32_and17_14_y0);
  fa fa_h_u_arrmul32_fa17_14_y2(h_u_arrmul32_and17_14_y0, h_u_arrmul32_fa18_13_y2, h_u_arrmul32_fa16_14_y4, h_u_arrmul32_fa17_14_y2, h_u_arrmul32_fa17_14_y4);
  and_gate and_gate_h_u_arrmul32_and18_14_y0(a_18, b_14, h_u_arrmul32_and18_14_y0);
  fa fa_h_u_arrmul32_fa18_14_y2(h_u_arrmul32_and18_14_y0, h_u_arrmul32_fa19_13_y2, h_u_arrmul32_fa17_14_y4, h_u_arrmul32_fa18_14_y2, h_u_arrmul32_fa18_14_y4);
  and_gate and_gate_h_u_arrmul32_and19_14_y0(a_19, b_14, h_u_arrmul32_and19_14_y0);
  fa fa_h_u_arrmul32_fa19_14_y2(h_u_arrmul32_and19_14_y0, h_u_arrmul32_fa20_13_y2, h_u_arrmul32_fa18_14_y4, h_u_arrmul32_fa19_14_y2, h_u_arrmul32_fa19_14_y4);
  and_gate and_gate_h_u_arrmul32_and20_14_y0(a_20, b_14, h_u_arrmul32_and20_14_y0);
  fa fa_h_u_arrmul32_fa20_14_y2(h_u_arrmul32_and20_14_y0, h_u_arrmul32_fa21_13_y2, h_u_arrmul32_fa19_14_y4, h_u_arrmul32_fa20_14_y2, h_u_arrmul32_fa20_14_y4);
  and_gate and_gate_h_u_arrmul32_and21_14_y0(a_21, b_14, h_u_arrmul32_and21_14_y0);
  fa fa_h_u_arrmul32_fa21_14_y2(h_u_arrmul32_and21_14_y0, h_u_arrmul32_fa22_13_y2, h_u_arrmul32_fa20_14_y4, h_u_arrmul32_fa21_14_y2, h_u_arrmul32_fa21_14_y4);
  and_gate and_gate_h_u_arrmul32_and22_14_y0(a_22, b_14, h_u_arrmul32_and22_14_y0);
  fa fa_h_u_arrmul32_fa22_14_y2(h_u_arrmul32_and22_14_y0, h_u_arrmul32_fa23_13_y2, h_u_arrmul32_fa21_14_y4, h_u_arrmul32_fa22_14_y2, h_u_arrmul32_fa22_14_y4);
  and_gate and_gate_h_u_arrmul32_and23_14_y0(a_23, b_14, h_u_arrmul32_and23_14_y0);
  fa fa_h_u_arrmul32_fa23_14_y2(h_u_arrmul32_and23_14_y0, h_u_arrmul32_fa24_13_y2, h_u_arrmul32_fa22_14_y4, h_u_arrmul32_fa23_14_y2, h_u_arrmul32_fa23_14_y4);
  and_gate and_gate_h_u_arrmul32_and24_14_y0(a_24, b_14, h_u_arrmul32_and24_14_y0);
  fa fa_h_u_arrmul32_fa24_14_y2(h_u_arrmul32_and24_14_y0, h_u_arrmul32_fa25_13_y2, h_u_arrmul32_fa23_14_y4, h_u_arrmul32_fa24_14_y2, h_u_arrmul32_fa24_14_y4);
  and_gate and_gate_h_u_arrmul32_and25_14_y0(a_25, b_14, h_u_arrmul32_and25_14_y0);
  fa fa_h_u_arrmul32_fa25_14_y2(h_u_arrmul32_and25_14_y0, h_u_arrmul32_fa26_13_y2, h_u_arrmul32_fa24_14_y4, h_u_arrmul32_fa25_14_y2, h_u_arrmul32_fa25_14_y4);
  and_gate and_gate_h_u_arrmul32_and26_14_y0(a_26, b_14, h_u_arrmul32_and26_14_y0);
  fa fa_h_u_arrmul32_fa26_14_y2(h_u_arrmul32_and26_14_y0, h_u_arrmul32_fa27_13_y2, h_u_arrmul32_fa25_14_y4, h_u_arrmul32_fa26_14_y2, h_u_arrmul32_fa26_14_y4);
  and_gate and_gate_h_u_arrmul32_and27_14_y0(a_27, b_14, h_u_arrmul32_and27_14_y0);
  fa fa_h_u_arrmul32_fa27_14_y2(h_u_arrmul32_and27_14_y0, h_u_arrmul32_fa28_13_y2, h_u_arrmul32_fa26_14_y4, h_u_arrmul32_fa27_14_y2, h_u_arrmul32_fa27_14_y4);
  and_gate and_gate_h_u_arrmul32_and28_14_y0(a_28, b_14, h_u_arrmul32_and28_14_y0);
  fa fa_h_u_arrmul32_fa28_14_y2(h_u_arrmul32_and28_14_y0, h_u_arrmul32_fa29_13_y2, h_u_arrmul32_fa27_14_y4, h_u_arrmul32_fa28_14_y2, h_u_arrmul32_fa28_14_y4);
  and_gate and_gate_h_u_arrmul32_and29_14_y0(a_29, b_14, h_u_arrmul32_and29_14_y0);
  fa fa_h_u_arrmul32_fa29_14_y2(h_u_arrmul32_and29_14_y0, h_u_arrmul32_fa30_13_y2, h_u_arrmul32_fa28_14_y4, h_u_arrmul32_fa29_14_y2, h_u_arrmul32_fa29_14_y4);
  and_gate and_gate_h_u_arrmul32_and30_14_y0(a_30, b_14, h_u_arrmul32_and30_14_y0);
  fa fa_h_u_arrmul32_fa30_14_y2(h_u_arrmul32_and30_14_y0, h_u_arrmul32_fa31_13_y2, h_u_arrmul32_fa29_14_y4, h_u_arrmul32_fa30_14_y2, h_u_arrmul32_fa30_14_y4);
  and_gate and_gate_h_u_arrmul32_and31_14_y0(a_31, b_14, h_u_arrmul32_and31_14_y0);
  fa fa_h_u_arrmul32_fa31_14_y2(h_u_arrmul32_and31_14_y0, h_u_arrmul32_fa31_13_y4, h_u_arrmul32_fa30_14_y4, h_u_arrmul32_fa31_14_y2, h_u_arrmul32_fa31_14_y4);
  and_gate and_gate_h_u_arrmul32_and0_15_y0(a_0, b_15, h_u_arrmul32_and0_15_y0);
  ha ha_h_u_arrmul32_ha0_15_y0(h_u_arrmul32_and0_15_y0, h_u_arrmul32_fa1_14_y2, h_u_arrmul32_ha0_15_y0, h_u_arrmul32_ha0_15_y1);
  and_gate and_gate_h_u_arrmul32_and1_15_y0(a_1, b_15, h_u_arrmul32_and1_15_y0);
  fa fa_h_u_arrmul32_fa1_15_y2(h_u_arrmul32_and1_15_y0, h_u_arrmul32_fa2_14_y2, h_u_arrmul32_ha0_15_y1, h_u_arrmul32_fa1_15_y2, h_u_arrmul32_fa1_15_y4);
  and_gate and_gate_h_u_arrmul32_and2_15_y0(a_2, b_15, h_u_arrmul32_and2_15_y0);
  fa fa_h_u_arrmul32_fa2_15_y2(h_u_arrmul32_and2_15_y0, h_u_arrmul32_fa3_14_y2, h_u_arrmul32_fa1_15_y4, h_u_arrmul32_fa2_15_y2, h_u_arrmul32_fa2_15_y4);
  and_gate and_gate_h_u_arrmul32_and3_15_y0(a_3, b_15, h_u_arrmul32_and3_15_y0);
  fa fa_h_u_arrmul32_fa3_15_y2(h_u_arrmul32_and3_15_y0, h_u_arrmul32_fa4_14_y2, h_u_arrmul32_fa2_15_y4, h_u_arrmul32_fa3_15_y2, h_u_arrmul32_fa3_15_y4);
  and_gate and_gate_h_u_arrmul32_and4_15_y0(a_4, b_15, h_u_arrmul32_and4_15_y0);
  fa fa_h_u_arrmul32_fa4_15_y2(h_u_arrmul32_and4_15_y0, h_u_arrmul32_fa5_14_y2, h_u_arrmul32_fa3_15_y4, h_u_arrmul32_fa4_15_y2, h_u_arrmul32_fa4_15_y4);
  and_gate and_gate_h_u_arrmul32_and5_15_y0(a_5, b_15, h_u_arrmul32_and5_15_y0);
  fa fa_h_u_arrmul32_fa5_15_y2(h_u_arrmul32_and5_15_y0, h_u_arrmul32_fa6_14_y2, h_u_arrmul32_fa4_15_y4, h_u_arrmul32_fa5_15_y2, h_u_arrmul32_fa5_15_y4);
  and_gate and_gate_h_u_arrmul32_and6_15_y0(a_6, b_15, h_u_arrmul32_and6_15_y0);
  fa fa_h_u_arrmul32_fa6_15_y2(h_u_arrmul32_and6_15_y0, h_u_arrmul32_fa7_14_y2, h_u_arrmul32_fa5_15_y4, h_u_arrmul32_fa6_15_y2, h_u_arrmul32_fa6_15_y4);
  and_gate and_gate_h_u_arrmul32_and7_15_y0(a_7, b_15, h_u_arrmul32_and7_15_y0);
  fa fa_h_u_arrmul32_fa7_15_y2(h_u_arrmul32_and7_15_y0, h_u_arrmul32_fa8_14_y2, h_u_arrmul32_fa6_15_y4, h_u_arrmul32_fa7_15_y2, h_u_arrmul32_fa7_15_y4);
  and_gate and_gate_h_u_arrmul32_and8_15_y0(a_8, b_15, h_u_arrmul32_and8_15_y0);
  fa fa_h_u_arrmul32_fa8_15_y2(h_u_arrmul32_and8_15_y0, h_u_arrmul32_fa9_14_y2, h_u_arrmul32_fa7_15_y4, h_u_arrmul32_fa8_15_y2, h_u_arrmul32_fa8_15_y4);
  and_gate and_gate_h_u_arrmul32_and9_15_y0(a_9, b_15, h_u_arrmul32_and9_15_y0);
  fa fa_h_u_arrmul32_fa9_15_y2(h_u_arrmul32_and9_15_y0, h_u_arrmul32_fa10_14_y2, h_u_arrmul32_fa8_15_y4, h_u_arrmul32_fa9_15_y2, h_u_arrmul32_fa9_15_y4);
  and_gate and_gate_h_u_arrmul32_and10_15_y0(a_10, b_15, h_u_arrmul32_and10_15_y0);
  fa fa_h_u_arrmul32_fa10_15_y2(h_u_arrmul32_and10_15_y0, h_u_arrmul32_fa11_14_y2, h_u_arrmul32_fa9_15_y4, h_u_arrmul32_fa10_15_y2, h_u_arrmul32_fa10_15_y4);
  and_gate and_gate_h_u_arrmul32_and11_15_y0(a_11, b_15, h_u_arrmul32_and11_15_y0);
  fa fa_h_u_arrmul32_fa11_15_y2(h_u_arrmul32_and11_15_y0, h_u_arrmul32_fa12_14_y2, h_u_arrmul32_fa10_15_y4, h_u_arrmul32_fa11_15_y2, h_u_arrmul32_fa11_15_y4);
  and_gate and_gate_h_u_arrmul32_and12_15_y0(a_12, b_15, h_u_arrmul32_and12_15_y0);
  fa fa_h_u_arrmul32_fa12_15_y2(h_u_arrmul32_and12_15_y0, h_u_arrmul32_fa13_14_y2, h_u_arrmul32_fa11_15_y4, h_u_arrmul32_fa12_15_y2, h_u_arrmul32_fa12_15_y4);
  and_gate and_gate_h_u_arrmul32_and13_15_y0(a_13, b_15, h_u_arrmul32_and13_15_y0);
  fa fa_h_u_arrmul32_fa13_15_y2(h_u_arrmul32_and13_15_y0, h_u_arrmul32_fa14_14_y2, h_u_arrmul32_fa12_15_y4, h_u_arrmul32_fa13_15_y2, h_u_arrmul32_fa13_15_y4);
  and_gate and_gate_h_u_arrmul32_and14_15_y0(a_14, b_15, h_u_arrmul32_and14_15_y0);
  fa fa_h_u_arrmul32_fa14_15_y2(h_u_arrmul32_and14_15_y0, h_u_arrmul32_fa15_14_y2, h_u_arrmul32_fa13_15_y4, h_u_arrmul32_fa14_15_y2, h_u_arrmul32_fa14_15_y4);
  and_gate and_gate_h_u_arrmul32_and15_15_y0(a_15, b_15, h_u_arrmul32_and15_15_y0);
  fa fa_h_u_arrmul32_fa15_15_y2(h_u_arrmul32_and15_15_y0, h_u_arrmul32_fa16_14_y2, h_u_arrmul32_fa14_15_y4, h_u_arrmul32_fa15_15_y2, h_u_arrmul32_fa15_15_y4);
  and_gate and_gate_h_u_arrmul32_and16_15_y0(a_16, b_15, h_u_arrmul32_and16_15_y0);
  fa fa_h_u_arrmul32_fa16_15_y2(h_u_arrmul32_and16_15_y0, h_u_arrmul32_fa17_14_y2, h_u_arrmul32_fa15_15_y4, h_u_arrmul32_fa16_15_y2, h_u_arrmul32_fa16_15_y4);
  and_gate and_gate_h_u_arrmul32_and17_15_y0(a_17, b_15, h_u_arrmul32_and17_15_y0);
  fa fa_h_u_arrmul32_fa17_15_y2(h_u_arrmul32_and17_15_y0, h_u_arrmul32_fa18_14_y2, h_u_arrmul32_fa16_15_y4, h_u_arrmul32_fa17_15_y2, h_u_arrmul32_fa17_15_y4);
  and_gate and_gate_h_u_arrmul32_and18_15_y0(a_18, b_15, h_u_arrmul32_and18_15_y0);
  fa fa_h_u_arrmul32_fa18_15_y2(h_u_arrmul32_and18_15_y0, h_u_arrmul32_fa19_14_y2, h_u_arrmul32_fa17_15_y4, h_u_arrmul32_fa18_15_y2, h_u_arrmul32_fa18_15_y4);
  and_gate and_gate_h_u_arrmul32_and19_15_y0(a_19, b_15, h_u_arrmul32_and19_15_y0);
  fa fa_h_u_arrmul32_fa19_15_y2(h_u_arrmul32_and19_15_y0, h_u_arrmul32_fa20_14_y2, h_u_arrmul32_fa18_15_y4, h_u_arrmul32_fa19_15_y2, h_u_arrmul32_fa19_15_y4);
  and_gate and_gate_h_u_arrmul32_and20_15_y0(a_20, b_15, h_u_arrmul32_and20_15_y0);
  fa fa_h_u_arrmul32_fa20_15_y2(h_u_arrmul32_and20_15_y0, h_u_arrmul32_fa21_14_y2, h_u_arrmul32_fa19_15_y4, h_u_arrmul32_fa20_15_y2, h_u_arrmul32_fa20_15_y4);
  and_gate and_gate_h_u_arrmul32_and21_15_y0(a_21, b_15, h_u_arrmul32_and21_15_y0);
  fa fa_h_u_arrmul32_fa21_15_y2(h_u_arrmul32_and21_15_y0, h_u_arrmul32_fa22_14_y2, h_u_arrmul32_fa20_15_y4, h_u_arrmul32_fa21_15_y2, h_u_arrmul32_fa21_15_y4);
  and_gate and_gate_h_u_arrmul32_and22_15_y0(a_22, b_15, h_u_arrmul32_and22_15_y0);
  fa fa_h_u_arrmul32_fa22_15_y2(h_u_arrmul32_and22_15_y0, h_u_arrmul32_fa23_14_y2, h_u_arrmul32_fa21_15_y4, h_u_arrmul32_fa22_15_y2, h_u_arrmul32_fa22_15_y4);
  and_gate and_gate_h_u_arrmul32_and23_15_y0(a_23, b_15, h_u_arrmul32_and23_15_y0);
  fa fa_h_u_arrmul32_fa23_15_y2(h_u_arrmul32_and23_15_y0, h_u_arrmul32_fa24_14_y2, h_u_arrmul32_fa22_15_y4, h_u_arrmul32_fa23_15_y2, h_u_arrmul32_fa23_15_y4);
  and_gate and_gate_h_u_arrmul32_and24_15_y0(a_24, b_15, h_u_arrmul32_and24_15_y0);
  fa fa_h_u_arrmul32_fa24_15_y2(h_u_arrmul32_and24_15_y0, h_u_arrmul32_fa25_14_y2, h_u_arrmul32_fa23_15_y4, h_u_arrmul32_fa24_15_y2, h_u_arrmul32_fa24_15_y4);
  and_gate and_gate_h_u_arrmul32_and25_15_y0(a_25, b_15, h_u_arrmul32_and25_15_y0);
  fa fa_h_u_arrmul32_fa25_15_y2(h_u_arrmul32_and25_15_y0, h_u_arrmul32_fa26_14_y2, h_u_arrmul32_fa24_15_y4, h_u_arrmul32_fa25_15_y2, h_u_arrmul32_fa25_15_y4);
  and_gate and_gate_h_u_arrmul32_and26_15_y0(a_26, b_15, h_u_arrmul32_and26_15_y0);
  fa fa_h_u_arrmul32_fa26_15_y2(h_u_arrmul32_and26_15_y0, h_u_arrmul32_fa27_14_y2, h_u_arrmul32_fa25_15_y4, h_u_arrmul32_fa26_15_y2, h_u_arrmul32_fa26_15_y4);
  and_gate and_gate_h_u_arrmul32_and27_15_y0(a_27, b_15, h_u_arrmul32_and27_15_y0);
  fa fa_h_u_arrmul32_fa27_15_y2(h_u_arrmul32_and27_15_y0, h_u_arrmul32_fa28_14_y2, h_u_arrmul32_fa26_15_y4, h_u_arrmul32_fa27_15_y2, h_u_arrmul32_fa27_15_y4);
  and_gate and_gate_h_u_arrmul32_and28_15_y0(a_28, b_15, h_u_arrmul32_and28_15_y0);
  fa fa_h_u_arrmul32_fa28_15_y2(h_u_arrmul32_and28_15_y0, h_u_arrmul32_fa29_14_y2, h_u_arrmul32_fa27_15_y4, h_u_arrmul32_fa28_15_y2, h_u_arrmul32_fa28_15_y4);
  and_gate and_gate_h_u_arrmul32_and29_15_y0(a_29, b_15, h_u_arrmul32_and29_15_y0);
  fa fa_h_u_arrmul32_fa29_15_y2(h_u_arrmul32_and29_15_y0, h_u_arrmul32_fa30_14_y2, h_u_arrmul32_fa28_15_y4, h_u_arrmul32_fa29_15_y2, h_u_arrmul32_fa29_15_y4);
  and_gate and_gate_h_u_arrmul32_and30_15_y0(a_30, b_15, h_u_arrmul32_and30_15_y0);
  fa fa_h_u_arrmul32_fa30_15_y2(h_u_arrmul32_and30_15_y0, h_u_arrmul32_fa31_14_y2, h_u_arrmul32_fa29_15_y4, h_u_arrmul32_fa30_15_y2, h_u_arrmul32_fa30_15_y4);
  and_gate and_gate_h_u_arrmul32_and31_15_y0(a_31, b_15, h_u_arrmul32_and31_15_y0);
  fa fa_h_u_arrmul32_fa31_15_y2(h_u_arrmul32_and31_15_y0, h_u_arrmul32_fa31_14_y4, h_u_arrmul32_fa30_15_y4, h_u_arrmul32_fa31_15_y2, h_u_arrmul32_fa31_15_y4);
  and_gate and_gate_h_u_arrmul32_and0_16_y0(a_0, b_16, h_u_arrmul32_and0_16_y0);
  ha ha_h_u_arrmul32_ha0_16_y0(h_u_arrmul32_and0_16_y0, h_u_arrmul32_fa1_15_y2, h_u_arrmul32_ha0_16_y0, h_u_arrmul32_ha0_16_y1);
  and_gate and_gate_h_u_arrmul32_and1_16_y0(a_1, b_16, h_u_arrmul32_and1_16_y0);
  fa fa_h_u_arrmul32_fa1_16_y2(h_u_arrmul32_and1_16_y0, h_u_arrmul32_fa2_15_y2, h_u_arrmul32_ha0_16_y1, h_u_arrmul32_fa1_16_y2, h_u_arrmul32_fa1_16_y4);
  and_gate and_gate_h_u_arrmul32_and2_16_y0(a_2, b_16, h_u_arrmul32_and2_16_y0);
  fa fa_h_u_arrmul32_fa2_16_y2(h_u_arrmul32_and2_16_y0, h_u_arrmul32_fa3_15_y2, h_u_arrmul32_fa1_16_y4, h_u_arrmul32_fa2_16_y2, h_u_arrmul32_fa2_16_y4);
  and_gate and_gate_h_u_arrmul32_and3_16_y0(a_3, b_16, h_u_arrmul32_and3_16_y0);
  fa fa_h_u_arrmul32_fa3_16_y2(h_u_arrmul32_and3_16_y0, h_u_arrmul32_fa4_15_y2, h_u_arrmul32_fa2_16_y4, h_u_arrmul32_fa3_16_y2, h_u_arrmul32_fa3_16_y4);
  and_gate and_gate_h_u_arrmul32_and4_16_y0(a_4, b_16, h_u_arrmul32_and4_16_y0);
  fa fa_h_u_arrmul32_fa4_16_y2(h_u_arrmul32_and4_16_y0, h_u_arrmul32_fa5_15_y2, h_u_arrmul32_fa3_16_y4, h_u_arrmul32_fa4_16_y2, h_u_arrmul32_fa4_16_y4);
  and_gate and_gate_h_u_arrmul32_and5_16_y0(a_5, b_16, h_u_arrmul32_and5_16_y0);
  fa fa_h_u_arrmul32_fa5_16_y2(h_u_arrmul32_and5_16_y0, h_u_arrmul32_fa6_15_y2, h_u_arrmul32_fa4_16_y4, h_u_arrmul32_fa5_16_y2, h_u_arrmul32_fa5_16_y4);
  and_gate and_gate_h_u_arrmul32_and6_16_y0(a_6, b_16, h_u_arrmul32_and6_16_y0);
  fa fa_h_u_arrmul32_fa6_16_y2(h_u_arrmul32_and6_16_y0, h_u_arrmul32_fa7_15_y2, h_u_arrmul32_fa5_16_y4, h_u_arrmul32_fa6_16_y2, h_u_arrmul32_fa6_16_y4);
  and_gate and_gate_h_u_arrmul32_and7_16_y0(a_7, b_16, h_u_arrmul32_and7_16_y0);
  fa fa_h_u_arrmul32_fa7_16_y2(h_u_arrmul32_and7_16_y0, h_u_arrmul32_fa8_15_y2, h_u_arrmul32_fa6_16_y4, h_u_arrmul32_fa7_16_y2, h_u_arrmul32_fa7_16_y4);
  and_gate and_gate_h_u_arrmul32_and8_16_y0(a_8, b_16, h_u_arrmul32_and8_16_y0);
  fa fa_h_u_arrmul32_fa8_16_y2(h_u_arrmul32_and8_16_y0, h_u_arrmul32_fa9_15_y2, h_u_arrmul32_fa7_16_y4, h_u_arrmul32_fa8_16_y2, h_u_arrmul32_fa8_16_y4);
  and_gate and_gate_h_u_arrmul32_and9_16_y0(a_9, b_16, h_u_arrmul32_and9_16_y0);
  fa fa_h_u_arrmul32_fa9_16_y2(h_u_arrmul32_and9_16_y0, h_u_arrmul32_fa10_15_y2, h_u_arrmul32_fa8_16_y4, h_u_arrmul32_fa9_16_y2, h_u_arrmul32_fa9_16_y4);
  and_gate and_gate_h_u_arrmul32_and10_16_y0(a_10, b_16, h_u_arrmul32_and10_16_y0);
  fa fa_h_u_arrmul32_fa10_16_y2(h_u_arrmul32_and10_16_y0, h_u_arrmul32_fa11_15_y2, h_u_arrmul32_fa9_16_y4, h_u_arrmul32_fa10_16_y2, h_u_arrmul32_fa10_16_y4);
  and_gate and_gate_h_u_arrmul32_and11_16_y0(a_11, b_16, h_u_arrmul32_and11_16_y0);
  fa fa_h_u_arrmul32_fa11_16_y2(h_u_arrmul32_and11_16_y0, h_u_arrmul32_fa12_15_y2, h_u_arrmul32_fa10_16_y4, h_u_arrmul32_fa11_16_y2, h_u_arrmul32_fa11_16_y4);
  and_gate and_gate_h_u_arrmul32_and12_16_y0(a_12, b_16, h_u_arrmul32_and12_16_y0);
  fa fa_h_u_arrmul32_fa12_16_y2(h_u_arrmul32_and12_16_y0, h_u_arrmul32_fa13_15_y2, h_u_arrmul32_fa11_16_y4, h_u_arrmul32_fa12_16_y2, h_u_arrmul32_fa12_16_y4);
  and_gate and_gate_h_u_arrmul32_and13_16_y0(a_13, b_16, h_u_arrmul32_and13_16_y0);
  fa fa_h_u_arrmul32_fa13_16_y2(h_u_arrmul32_and13_16_y0, h_u_arrmul32_fa14_15_y2, h_u_arrmul32_fa12_16_y4, h_u_arrmul32_fa13_16_y2, h_u_arrmul32_fa13_16_y4);
  and_gate and_gate_h_u_arrmul32_and14_16_y0(a_14, b_16, h_u_arrmul32_and14_16_y0);
  fa fa_h_u_arrmul32_fa14_16_y2(h_u_arrmul32_and14_16_y0, h_u_arrmul32_fa15_15_y2, h_u_arrmul32_fa13_16_y4, h_u_arrmul32_fa14_16_y2, h_u_arrmul32_fa14_16_y4);
  and_gate and_gate_h_u_arrmul32_and15_16_y0(a_15, b_16, h_u_arrmul32_and15_16_y0);
  fa fa_h_u_arrmul32_fa15_16_y2(h_u_arrmul32_and15_16_y0, h_u_arrmul32_fa16_15_y2, h_u_arrmul32_fa14_16_y4, h_u_arrmul32_fa15_16_y2, h_u_arrmul32_fa15_16_y4);
  and_gate and_gate_h_u_arrmul32_and16_16_y0(a_16, b_16, h_u_arrmul32_and16_16_y0);
  fa fa_h_u_arrmul32_fa16_16_y2(h_u_arrmul32_and16_16_y0, h_u_arrmul32_fa17_15_y2, h_u_arrmul32_fa15_16_y4, h_u_arrmul32_fa16_16_y2, h_u_arrmul32_fa16_16_y4);
  and_gate and_gate_h_u_arrmul32_and17_16_y0(a_17, b_16, h_u_arrmul32_and17_16_y0);
  fa fa_h_u_arrmul32_fa17_16_y2(h_u_arrmul32_and17_16_y0, h_u_arrmul32_fa18_15_y2, h_u_arrmul32_fa16_16_y4, h_u_arrmul32_fa17_16_y2, h_u_arrmul32_fa17_16_y4);
  and_gate and_gate_h_u_arrmul32_and18_16_y0(a_18, b_16, h_u_arrmul32_and18_16_y0);
  fa fa_h_u_arrmul32_fa18_16_y2(h_u_arrmul32_and18_16_y0, h_u_arrmul32_fa19_15_y2, h_u_arrmul32_fa17_16_y4, h_u_arrmul32_fa18_16_y2, h_u_arrmul32_fa18_16_y4);
  and_gate and_gate_h_u_arrmul32_and19_16_y0(a_19, b_16, h_u_arrmul32_and19_16_y0);
  fa fa_h_u_arrmul32_fa19_16_y2(h_u_arrmul32_and19_16_y0, h_u_arrmul32_fa20_15_y2, h_u_arrmul32_fa18_16_y4, h_u_arrmul32_fa19_16_y2, h_u_arrmul32_fa19_16_y4);
  and_gate and_gate_h_u_arrmul32_and20_16_y0(a_20, b_16, h_u_arrmul32_and20_16_y0);
  fa fa_h_u_arrmul32_fa20_16_y2(h_u_arrmul32_and20_16_y0, h_u_arrmul32_fa21_15_y2, h_u_arrmul32_fa19_16_y4, h_u_arrmul32_fa20_16_y2, h_u_arrmul32_fa20_16_y4);
  and_gate and_gate_h_u_arrmul32_and21_16_y0(a_21, b_16, h_u_arrmul32_and21_16_y0);
  fa fa_h_u_arrmul32_fa21_16_y2(h_u_arrmul32_and21_16_y0, h_u_arrmul32_fa22_15_y2, h_u_arrmul32_fa20_16_y4, h_u_arrmul32_fa21_16_y2, h_u_arrmul32_fa21_16_y4);
  and_gate and_gate_h_u_arrmul32_and22_16_y0(a_22, b_16, h_u_arrmul32_and22_16_y0);
  fa fa_h_u_arrmul32_fa22_16_y2(h_u_arrmul32_and22_16_y0, h_u_arrmul32_fa23_15_y2, h_u_arrmul32_fa21_16_y4, h_u_arrmul32_fa22_16_y2, h_u_arrmul32_fa22_16_y4);
  and_gate and_gate_h_u_arrmul32_and23_16_y0(a_23, b_16, h_u_arrmul32_and23_16_y0);
  fa fa_h_u_arrmul32_fa23_16_y2(h_u_arrmul32_and23_16_y0, h_u_arrmul32_fa24_15_y2, h_u_arrmul32_fa22_16_y4, h_u_arrmul32_fa23_16_y2, h_u_arrmul32_fa23_16_y4);
  and_gate and_gate_h_u_arrmul32_and24_16_y0(a_24, b_16, h_u_arrmul32_and24_16_y0);
  fa fa_h_u_arrmul32_fa24_16_y2(h_u_arrmul32_and24_16_y0, h_u_arrmul32_fa25_15_y2, h_u_arrmul32_fa23_16_y4, h_u_arrmul32_fa24_16_y2, h_u_arrmul32_fa24_16_y4);
  and_gate and_gate_h_u_arrmul32_and25_16_y0(a_25, b_16, h_u_arrmul32_and25_16_y0);
  fa fa_h_u_arrmul32_fa25_16_y2(h_u_arrmul32_and25_16_y0, h_u_arrmul32_fa26_15_y2, h_u_arrmul32_fa24_16_y4, h_u_arrmul32_fa25_16_y2, h_u_arrmul32_fa25_16_y4);
  and_gate and_gate_h_u_arrmul32_and26_16_y0(a_26, b_16, h_u_arrmul32_and26_16_y0);
  fa fa_h_u_arrmul32_fa26_16_y2(h_u_arrmul32_and26_16_y0, h_u_arrmul32_fa27_15_y2, h_u_arrmul32_fa25_16_y4, h_u_arrmul32_fa26_16_y2, h_u_arrmul32_fa26_16_y4);
  and_gate and_gate_h_u_arrmul32_and27_16_y0(a_27, b_16, h_u_arrmul32_and27_16_y0);
  fa fa_h_u_arrmul32_fa27_16_y2(h_u_arrmul32_and27_16_y0, h_u_arrmul32_fa28_15_y2, h_u_arrmul32_fa26_16_y4, h_u_arrmul32_fa27_16_y2, h_u_arrmul32_fa27_16_y4);
  and_gate and_gate_h_u_arrmul32_and28_16_y0(a_28, b_16, h_u_arrmul32_and28_16_y0);
  fa fa_h_u_arrmul32_fa28_16_y2(h_u_arrmul32_and28_16_y0, h_u_arrmul32_fa29_15_y2, h_u_arrmul32_fa27_16_y4, h_u_arrmul32_fa28_16_y2, h_u_arrmul32_fa28_16_y4);
  and_gate and_gate_h_u_arrmul32_and29_16_y0(a_29, b_16, h_u_arrmul32_and29_16_y0);
  fa fa_h_u_arrmul32_fa29_16_y2(h_u_arrmul32_and29_16_y0, h_u_arrmul32_fa30_15_y2, h_u_arrmul32_fa28_16_y4, h_u_arrmul32_fa29_16_y2, h_u_arrmul32_fa29_16_y4);
  and_gate and_gate_h_u_arrmul32_and30_16_y0(a_30, b_16, h_u_arrmul32_and30_16_y0);
  fa fa_h_u_arrmul32_fa30_16_y2(h_u_arrmul32_and30_16_y0, h_u_arrmul32_fa31_15_y2, h_u_arrmul32_fa29_16_y4, h_u_arrmul32_fa30_16_y2, h_u_arrmul32_fa30_16_y4);
  and_gate and_gate_h_u_arrmul32_and31_16_y0(a_31, b_16, h_u_arrmul32_and31_16_y0);
  fa fa_h_u_arrmul32_fa31_16_y2(h_u_arrmul32_and31_16_y0, h_u_arrmul32_fa31_15_y4, h_u_arrmul32_fa30_16_y4, h_u_arrmul32_fa31_16_y2, h_u_arrmul32_fa31_16_y4);
  and_gate and_gate_h_u_arrmul32_and0_17_y0(a_0, b_17, h_u_arrmul32_and0_17_y0);
  ha ha_h_u_arrmul32_ha0_17_y0(h_u_arrmul32_and0_17_y0, h_u_arrmul32_fa1_16_y2, h_u_arrmul32_ha0_17_y0, h_u_arrmul32_ha0_17_y1);
  and_gate and_gate_h_u_arrmul32_and1_17_y0(a_1, b_17, h_u_arrmul32_and1_17_y0);
  fa fa_h_u_arrmul32_fa1_17_y2(h_u_arrmul32_and1_17_y0, h_u_arrmul32_fa2_16_y2, h_u_arrmul32_ha0_17_y1, h_u_arrmul32_fa1_17_y2, h_u_arrmul32_fa1_17_y4);
  and_gate and_gate_h_u_arrmul32_and2_17_y0(a_2, b_17, h_u_arrmul32_and2_17_y0);
  fa fa_h_u_arrmul32_fa2_17_y2(h_u_arrmul32_and2_17_y0, h_u_arrmul32_fa3_16_y2, h_u_arrmul32_fa1_17_y4, h_u_arrmul32_fa2_17_y2, h_u_arrmul32_fa2_17_y4);
  and_gate and_gate_h_u_arrmul32_and3_17_y0(a_3, b_17, h_u_arrmul32_and3_17_y0);
  fa fa_h_u_arrmul32_fa3_17_y2(h_u_arrmul32_and3_17_y0, h_u_arrmul32_fa4_16_y2, h_u_arrmul32_fa2_17_y4, h_u_arrmul32_fa3_17_y2, h_u_arrmul32_fa3_17_y4);
  and_gate and_gate_h_u_arrmul32_and4_17_y0(a_4, b_17, h_u_arrmul32_and4_17_y0);
  fa fa_h_u_arrmul32_fa4_17_y2(h_u_arrmul32_and4_17_y0, h_u_arrmul32_fa5_16_y2, h_u_arrmul32_fa3_17_y4, h_u_arrmul32_fa4_17_y2, h_u_arrmul32_fa4_17_y4);
  and_gate and_gate_h_u_arrmul32_and5_17_y0(a_5, b_17, h_u_arrmul32_and5_17_y0);
  fa fa_h_u_arrmul32_fa5_17_y2(h_u_arrmul32_and5_17_y0, h_u_arrmul32_fa6_16_y2, h_u_arrmul32_fa4_17_y4, h_u_arrmul32_fa5_17_y2, h_u_arrmul32_fa5_17_y4);
  and_gate and_gate_h_u_arrmul32_and6_17_y0(a_6, b_17, h_u_arrmul32_and6_17_y0);
  fa fa_h_u_arrmul32_fa6_17_y2(h_u_arrmul32_and6_17_y0, h_u_arrmul32_fa7_16_y2, h_u_arrmul32_fa5_17_y4, h_u_arrmul32_fa6_17_y2, h_u_arrmul32_fa6_17_y4);
  and_gate and_gate_h_u_arrmul32_and7_17_y0(a_7, b_17, h_u_arrmul32_and7_17_y0);
  fa fa_h_u_arrmul32_fa7_17_y2(h_u_arrmul32_and7_17_y0, h_u_arrmul32_fa8_16_y2, h_u_arrmul32_fa6_17_y4, h_u_arrmul32_fa7_17_y2, h_u_arrmul32_fa7_17_y4);
  and_gate and_gate_h_u_arrmul32_and8_17_y0(a_8, b_17, h_u_arrmul32_and8_17_y0);
  fa fa_h_u_arrmul32_fa8_17_y2(h_u_arrmul32_and8_17_y0, h_u_arrmul32_fa9_16_y2, h_u_arrmul32_fa7_17_y4, h_u_arrmul32_fa8_17_y2, h_u_arrmul32_fa8_17_y4);
  and_gate and_gate_h_u_arrmul32_and9_17_y0(a_9, b_17, h_u_arrmul32_and9_17_y0);
  fa fa_h_u_arrmul32_fa9_17_y2(h_u_arrmul32_and9_17_y0, h_u_arrmul32_fa10_16_y2, h_u_arrmul32_fa8_17_y4, h_u_arrmul32_fa9_17_y2, h_u_arrmul32_fa9_17_y4);
  and_gate and_gate_h_u_arrmul32_and10_17_y0(a_10, b_17, h_u_arrmul32_and10_17_y0);
  fa fa_h_u_arrmul32_fa10_17_y2(h_u_arrmul32_and10_17_y0, h_u_arrmul32_fa11_16_y2, h_u_arrmul32_fa9_17_y4, h_u_arrmul32_fa10_17_y2, h_u_arrmul32_fa10_17_y4);
  and_gate and_gate_h_u_arrmul32_and11_17_y0(a_11, b_17, h_u_arrmul32_and11_17_y0);
  fa fa_h_u_arrmul32_fa11_17_y2(h_u_arrmul32_and11_17_y0, h_u_arrmul32_fa12_16_y2, h_u_arrmul32_fa10_17_y4, h_u_arrmul32_fa11_17_y2, h_u_arrmul32_fa11_17_y4);
  and_gate and_gate_h_u_arrmul32_and12_17_y0(a_12, b_17, h_u_arrmul32_and12_17_y0);
  fa fa_h_u_arrmul32_fa12_17_y2(h_u_arrmul32_and12_17_y0, h_u_arrmul32_fa13_16_y2, h_u_arrmul32_fa11_17_y4, h_u_arrmul32_fa12_17_y2, h_u_arrmul32_fa12_17_y4);
  and_gate and_gate_h_u_arrmul32_and13_17_y0(a_13, b_17, h_u_arrmul32_and13_17_y0);
  fa fa_h_u_arrmul32_fa13_17_y2(h_u_arrmul32_and13_17_y0, h_u_arrmul32_fa14_16_y2, h_u_arrmul32_fa12_17_y4, h_u_arrmul32_fa13_17_y2, h_u_arrmul32_fa13_17_y4);
  and_gate and_gate_h_u_arrmul32_and14_17_y0(a_14, b_17, h_u_arrmul32_and14_17_y0);
  fa fa_h_u_arrmul32_fa14_17_y2(h_u_arrmul32_and14_17_y0, h_u_arrmul32_fa15_16_y2, h_u_arrmul32_fa13_17_y4, h_u_arrmul32_fa14_17_y2, h_u_arrmul32_fa14_17_y4);
  and_gate and_gate_h_u_arrmul32_and15_17_y0(a_15, b_17, h_u_arrmul32_and15_17_y0);
  fa fa_h_u_arrmul32_fa15_17_y2(h_u_arrmul32_and15_17_y0, h_u_arrmul32_fa16_16_y2, h_u_arrmul32_fa14_17_y4, h_u_arrmul32_fa15_17_y2, h_u_arrmul32_fa15_17_y4);
  and_gate and_gate_h_u_arrmul32_and16_17_y0(a_16, b_17, h_u_arrmul32_and16_17_y0);
  fa fa_h_u_arrmul32_fa16_17_y2(h_u_arrmul32_and16_17_y0, h_u_arrmul32_fa17_16_y2, h_u_arrmul32_fa15_17_y4, h_u_arrmul32_fa16_17_y2, h_u_arrmul32_fa16_17_y4);
  and_gate and_gate_h_u_arrmul32_and17_17_y0(a_17, b_17, h_u_arrmul32_and17_17_y0);
  fa fa_h_u_arrmul32_fa17_17_y2(h_u_arrmul32_and17_17_y0, h_u_arrmul32_fa18_16_y2, h_u_arrmul32_fa16_17_y4, h_u_arrmul32_fa17_17_y2, h_u_arrmul32_fa17_17_y4);
  and_gate and_gate_h_u_arrmul32_and18_17_y0(a_18, b_17, h_u_arrmul32_and18_17_y0);
  fa fa_h_u_arrmul32_fa18_17_y2(h_u_arrmul32_and18_17_y0, h_u_arrmul32_fa19_16_y2, h_u_arrmul32_fa17_17_y4, h_u_arrmul32_fa18_17_y2, h_u_arrmul32_fa18_17_y4);
  and_gate and_gate_h_u_arrmul32_and19_17_y0(a_19, b_17, h_u_arrmul32_and19_17_y0);
  fa fa_h_u_arrmul32_fa19_17_y2(h_u_arrmul32_and19_17_y0, h_u_arrmul32_fa20_16_y2, h_u_arrmul32_fa18_17_y4, h_u_arrmul32_fa19_17_y2, h_u_arrmul32_fa19_17_y4);
  and_gate and_gate_h_u_arrmul32_and20_17_y0(a_20, b_17, h_u_arrmul32_and20_17_y0);
  fa fa_h_u_arrmul32_fa20_17_y2(h_u_arrmul32_and20_17_y0, h_u_arrmul32_fa21_16_y2, h_u_arrmul32_fa19_17_y4, h_u_arrmul32_fa20_17_y2, h_u_arrmul32_fa20_17_y4);
  and_gate and_gate_h_u_arrmul32_and21_17_y0(a_21, b_17, h_u_arrmul32_and21_17_y0);
  fa fa_h_u_arrmul32_fa21_17_y2(h_u_arrmul32_and21_17_y0, h_u_arrmul32_fa22_16_y2, h_u_arrmul32_fa20_17_y4, h_u_arrmul32_fa21_17_y2, h_u_arrmul32_fa21_17_y4);
  and_gate and_gate_h_u_arrmul32_and22_17_y0(a_22, b_17, h_u_arrmul32_and22_17_y0);
  fa fa_h_u_arrmul32_fa22_17_y2(h_u_arrmul32_and22_17_y0, h_u_arrmul32_fa23_16_y2, h_u_arrmul32_fa21_17_y4, h_u_arrmul32_fa22_17_y2, h_u_arrmul32_fa22_17_y4);
  and_gate and_gate_h_u_arrmul32_and23_17_y0(a_23, b_17, h_u_arrmul32_and23_17_y0);
  fa fa_h_u_arrmul32_fa23_17_y2(h_u_arrmul32_and23_17_y0, h_u_arrmul32_fa24_16_y2, h_u_arrmul32_fa22_17_y4, h_u_arrmul32_fa23_17_y2, h_u_arrmul32_fa23_17_y4);
  and_gate and_gate_h_u_arrmul32_and24_17_y0(a_24, b_17, h_u_arrmul32_and24_17_y0);
  fa fa_h_u_arrmul32_fa24_17_y2(h_u_arrmul32_and24_17_y0, h_u_arrmul32_fa25_16_y2, h_u_arrmul32_fa23_17_y4, h_u_arrmul32_fa24_17_y2, h_u_arrmul32_fa24_17_y4);
  and_gate and_gate_h_u_arrmul32_and25_17_y0(a_25, b_17, h_u_arrmul32_and25_17_y0);
  fa fa_h_u_arrmul32_fa25_17_y2(h_u_arrmul32_and25_17_y0, h_u_arrmul32_fa26_16_y2, h_u_arrmul32_fa24_17_y4, h_u_arrmul32_fa25_17_y2, h_u_arrmul32_fa25_17_y4);
  and_gate and_gate_h_u_arrmul32_and26_17_y0(a_26, b_17, h_u_arrmul32_and26_17_y0);
  fa fa_h_u_arrmul32_fa26_17_y2(h_u_arrmul32_and26_17_y0, h_u_arrmul32_fa27_16_y2, h_u_arrmul32_fa25_17_y4, h_u_arrmul32_fa26_17_y2, h_u_arrmul32_fa26_17_y4);
  and_gate and_gate_h_u_arrmul32_and27_17_y0(a_27, b_17, h_u_arrmul32_and27_17_y0);
  fa fa_h_u_arrmul32_fa27_17_y2(h_u_arrmul32_and27_17_y0, h_u_arrmul32_fa28_16_y2, h_u_arrmul32_fa26_17_y4, h_u_arrmul32_fa27_17_y2, h_u_arrmul32_fa27_17_y4);
  and_gate and_gate_h_u_arrmul32_and28_17_y0(a_28, b_17, h_u_arrmul32_and28_17_y0);
  fa fa_h_u_arrmul32_fa28_17_y2(h_u_arrmul32_and28_17_y0, h_u_arrmul32_fa29_16_y2, h_u_arrmul32_fa27_17_y4, h_u_arrmul32_fa28_17_y2, h_u_arrmul32_fa28_17_y4);
  and_gate and_gate_h_u_arrmul32_and29_17_y0(a_29, b_17, h_u_arrmul32_and29_17_y0);
  fa fa_h_u_arrmul32_fa29_17_y2(h_u_arrmul32_and29_17_y0, h_u_arrmul32_fa30_16_y2, h_u_arrmul32_fa28_17_y4, h_u_arrmul32_fa29_17_y2, h_u_arrmul32_fa29_17_y4);
  and_gate and_gate_h_u_arrmul32_and30_17_y0(a_30, b_17, h_u_arrmul32_and30_17_y0);
  fa fa_h_u_arrmul32_fa30_17_y2(h_u_arrmul32_and30_17_y0, h_u_arrmul32_fa31_16_y2, h_u_arrmul32_fa29_17_y4, h_u_arrmul32_fa30_17_y2, h_u_arrmul32_fa30_17_y4);
  and_gate and_gate_h_u_arrmul32_and31_17_y0(a_31, b_17, h_u_arrmul32_and31_17_y0);
  fa fa_h_u_arrmul32_fa31_17_y2(h_u_arrmul32_and31_17_y0, h_u_arrmul32_fa31_16_y4, h_u_arrmul32_fa30_17_y4, h_u_arrmul32_fa31_17_y2, h_u_arrmul32_fa31_17_y4);
  and_gate and_gate_h_u_arrmul32_and0_18_y0(a_0, b_18, h_u_arrmul32_and0_18_y0);
  ha ha_h_u_arrmul32_ha0_18_y0(h_u_arrmul32_and0_18_y0, h_u_arrmul32_fa1_17_y2, h_u_arrmul32_ha0_18_y0, h_u_arrmul32_ha0_18_y1);
  and_gate and_gate_h_u_arrmul32_and1_18_y0(a_1, b_18, h_u_arrmul32_and1_18_y0);
  fa fa_h_u_arrmul32_fa1_18_y2(h_u_arrmul32_and1_18_y0, h_u_arrmul32_fa2_17_y2, h_u_arrmul32_ha0_18_y1, h_u_arrmul32_fa1_18_y2, h_u_arrmul32_fa1_18_y4);
  and_gate and_gate_h_u_arrmul32_and2_18_y0(a_2, b_18, h_u_arrmul32_and2_18_y0);
  fa fa_h_u_arrmul32_fa2_18_y2(h_u_arrmul32_and2_18_y0, h_u_arrmul32_fa3_17_y2, h_u_arrmul32_fa1_18_y4, h_u_arrmul32_fa2_18_y2, h_u_arrmul32_fa2_18_y4);
  and_gate and_gate_h_u_arrmul32_and3_18_y0(a_3, b_18, h_u_arrmul32_and3_18_y0);
  fa fa_h_u_arrmul32_fa3_18_y2(h_u_arrmul32_and3_18_y0, h_u_arrmul32_fa4_17_y2, h_u_arrmul32_fa2_18_y4, h_u_arrmul32_fa3_18_y2, h_u_arrmul32_fa3_18_y4);
  and_gate and_gate_h_u_arrmul32_and4_18_y0(a_4, b_18, h_u_arrmul32_and4_18_y0);
  fa fa_h_u_arrmul32_fa4_18_y2(h_u_arrmul32_and4_18_y0, h_u_arrmul32_fa5_17_y2, h_u_arrmul32_fa3_18_y4, h_u_arrmul32_fa4_18_y2, h_u_arrmul32_fa4_18_y4);
  and_gate and_gate_h_u_arrmul32_and5_18_y0(a_5, b_18, h_u_arrmul32_and5_18_y0);
  fa fa_h_u_arrmul32_fa5_18_y2(h_u_arrmul32_and5_18_y0, h_u_arrmul32_fa6_17_y2, h_u_arrmul32_fa4_18_y4, h_u_arrmul32_fa5_18_y2, h_u_arrmul32_fa5_18_y4);
  and_gate and_gate_h_u_arrmul32_and6_18_y0(a_6, b_18, h_u_arrmul32_and6_18_y0);
  fa fa_h_u_arrmul32_fa6_18_y2(h_u_arrmul32_and6_18_y0, h_u_arrmul32_fa7_17_y2, h_u_arrmul32_fa5_18_y4, h_u_arrmul32_fa6_18_y2, h_u_arrmul32_fa6_18_y4);
  and_gate and_gate_h_u_arrmul32_and7_18_y0(a_7, b_18, h_u_arrmul32_and7_18_y0);
  fa fa_h_u_arrmul32_fa7_18_y2(h_u_arrmul32_and7_18_y0, h_u_arrmul32_fa8_17_y2, h_u_arrmul32_fa6_18_y4, h_u_arrmul32_fa7_18_y2, h_u_arrmul32_fa7_18_y4);
  and_gate and_gate_h_u_arrmul32_and8_18_y0(a_8, b_18, h_u_arrmul32_and8_18_y0);
  fa fa_h_u_arrmul32_fa8_18_y2(h_u_arrmul32_and8_18_y0, h_u_arrmul32_fa9_17_y2, h_u_arrmul32_fa7_18_y4, h_u_arrmul32_fa8_18_y2, h_u_arrmul32_fa8_18_y4);
  and_gate and_gate_h_u_arrmul32_and9_18_y0(a_9, b_18, h_u_arrmul32_and9_18_y0);
  fa fa_h_u_arrmul32_fa9_18_y2(h_u_arrmul32_and9_18_y0, h_u_arrmul32_fa10_17_y2, h_u_arrmul32_fa8_18_y4, h_u_arrmul32_fa9_18_y2, h_u_arrmul32_fa9_18_y4);
  and_gate and_gate_h_u_arrmul32_and10_18_y0(a_10, b_18, h_u_arrmul32_and10_18_y0);
  fa fa_h_u_arrmul32_fa10_18_y2(h_u_arrmul32_and10_18_y0, h_u_arrmul32_fa11_17_y2, h_u_arrmul32_fa9_18_y4, h_u_arrmul32_fa10_18_y2, h_u_arrmul32_fa10_18_y4);
  and_gate and_gate_h_u_arrmul32_and11_18_y0(a_11, b_18, h_u_arrmul32_and11_18_y0);
  fa fa_h_u_arrmul32_fa11_18_y2(h_u_arrmul32_and11_18_y0, h_u_arrmul32_fa12_17_y2, h_u_arrmul32_fa10_18_y4, h_u_arrmul32_fa11_18_y2, h_u_arrmul32_fa11_18_y4);
  and_gate and_gate_h_u_arrmul32_and12_18_y0(a_12, b_18, h_u_arrmul32_and12_18_y0);
  fa fa_h_u_arrmul32_fa12_18_y2(h_u_arrmul32_and12_18_y0, h_u_arrmul32_fa13_17_y2, h_u_arrmul32_fa11_18_y4, h_u_arrmul32_fa12_18_y2, h_u_arrmul32_fa12_18_y4);
  and_gate and_gate_h_u_arrmul32_and13_18_y0(a_13, b_18, h_u_arrmul32_and13_18_y0);
  fa fa_h_u_arrmul32_fa13_18_y2(h_u_arrmul32_and13_18_y0, h_u_arrmul32_fa14_17_y2, h_u_arrmul32_fa12_18_y4, h_u_arrmul32_fa13_18_y2, h_u_arrmul32_fa13_18_y4);
  and_gate and_gate_h_u_arrmul32_and14_18_y0(a_14, b_18, h_u_arrmul32_and14_18_y0);
  fa fa_h_u_arrmul32_fa14_18_y2(h_u_arrmul32_and14_18_y0, h_u_arrmul32_fa15_17_y2, h_u_arrmul32_fa13_18_y4, h_u_arrmul32_fa14_18_y2, h_u_arrmul32_fa14_18_y4);
  and_gate and_gate_h_u_arrmul32_and15_18_y0(a_15, b_18, h_u_arrmul32_and15_18_y0);
  fa fa_h_u_arrmul32_fa15_18_y2(h_u_arrmul32_and15_18_y0, h_u_arrmul32_fa16_17_y2, h_u_arrmul32_fa14_18_y4, h_u_arrmul32_fa15_18_y2, h_u_arrmul32_fa15_18_y4);
  and_gate and_gate_h_u_arrmul32_and16_18_y0(a_16, b_18, h_u_arrmul32_and16_18_y0);
  fa fa_h_u_arrmul32_fa16_18_y2(h_u_arrmul32_and16_18_y0, h_u_arrmul32_fa17_17_y2, h_u_arrmul32_fa15_18_y4, h_u_arrmul32_fa16_18_y2, h_u_arrmul32_fa16_18_y4);
  and_gate and_gate_h_u_arrmul32_and17_18_y0(a_17, b_18, h_u_arrmul32_and17_18_y0);
  fa fa_h_u_arrmul32_fa17_18_y2(h_u_arrmul32_and17_18_y0, h_u_arrmul32_fa18_17_y2, h_u_arrmul32_fa16_18_y4, h_u_arrmul32_fa17_18_y2, h_u_arrmul32_fa17_18_y4);
  and_gate and_gate_h_u_arrmul32_and18_18_y0(a_18, b_18, h_u_arrmul32_and18_18_y0);
  fa fa_h_u_arrmul32_fa18_18_y2(h_u_arrmul32_and18_18_y0, h_u_arrmul32_fa19_17_y2, h_u_arrmul32_fa17_18_y4, h_u_arrmul32_fa18_18_y2, h_u_arrmul32_fa18_18_y4);
  and_gate and_gate_h_u_arrmul32_and19_18_y0(a_19, b_18, h_u_arrmul32_and19_18_y0);
  fa fa_h_u_arrmul32_fa19_18_y2(h_u_arrmul32_and19_18_y0, h_u_arrmul32_fa20_17_y2, h_u_arrmul32_fa18_18_y4, h_u_arrmul32_fa19_18_y2, h_u_arrmul32_fa19_18_y4);
  and_gate and_gate_h_u_arrmul32_and20_18_y0(a_20, b_18, h_u_arrmul32_and20_18_y0);
  fa fa_h_u_arrmul32_fa20_18_y2(h_u_arrmul32_and20_18_y0, h_u_arrmul32_fa21_17_y2, h_u_arrmul32_fa19_18_y4, h_u_arrmul32_fa20_18_y2, h_u_arrmul32_fa20_18_y4);
  and_gate and_gate_h_u_arrmul32_and21_18_y0(a_21, b_18, h_u_arrmul32_and21_18_y0);
  fa fa_h_u_arrmul32_fa21_18_y2(h_u_arrmul32_and21_18_y0, h_u_arrmul32_fa22_17_y2, h_u_arrmul32_fa20_18_y4, h_u_arrmul32_fa21_18_y2, h_u_arrmul32_fa21_18_y4);
  and_gate and_gate_h_u_arrmul32_and22_18_y0(a_22, b_18, h_u_arrmul32_and22_18_y0);
  fa fa_h_u_arrmul32_fa22_18_y2(h_u_arrmul32_and22_18_y0, h_u_arrmul32_fa23_17_y2, h_u_arrmul32_fa21_18_y4, h_u_arrmul32_fa22_18_y2, h_u_arrmul32_fa22_18_y4);
  and_gate and_gate_h_u_arrmul32_and23_18_y0(a_23, b_18, h_u_arrmul32_and23_18_y0);
  fa fa_h_u_arrmul32_fa23_18_y2(h_u_arrmul32_and23_18_y0, h_u_arrmul32_fa24_17_y2, h_u_arrmul32_fa22_18_y4, h_u_arrmul32_fa23_18_y2, h_u_arrmul32_fa23_18_y4);
  and_gate and_gate_h_u_arrmul32_and24_18_y0(a_24, b_18, h_u_arrmul32_and24_18_y0);
  fa fa_h_u_arrmul32_fa24_18_y2(h_u_arrmul32_and24_18_y0, h_u_arrmul32_fa25_17_y2, h_u_arrmul32_fa23_18_y4, h_u_arrmul32_fa24_18_y2, h_u_arrmul32_fa24_18_y4);
  and_gate and_gate_h_u_arrmul32_and25_18_y0(a_25, b_18, h_u_arrmul32_and25_18_y0);
  fa fa_h_u_arrmul32_fa25_18_y2(h_u_arrmul32_and25_18_y0, h_u_arrmul32_fa26_17_y2, h_u_arrmul32_fa24_18_y4, h_u_arrmul32_fa25_18_y2, h_u_arrmul32_fa25_18_y4);
  and_gate and_gate_h_u_arrmul32_and26_18_y0(a_26, b_18, h_u_arrmul32_and26_18_y0);
  fa fa_h_u_arrmul32_fa26_18_y2(h_u_arrmul32_and26_18_y0, h_u_arrmul32_fa27_17_y2, h_u_arrmul32_fa25_18_y4, h_u_arrmul32_fa26_18_y2, h_u_arrmul32_fa26_18_y4);
  and_gate and_gate_h_u_arrmul32_and27_18_y0(a_27, b_18, h_u_arrmul32_and27_18_y0);
  fa fa_h_u_arrmul32_fa27_18_y2(h_u_arrmul32_and27_18_y0, h_u_arrmul32_fa28_17_y2, h_u_arrmul32_fa26_18_y4, h_u_arrmul32_fa27_18_y2, h_u_arrmul32_fa27_18_y4);
  and_gate and_gate_h_u_arrmul32_and28_18_y0(a_28, b_18, h_u_arrmul32_and28_18_y0);
  fa fa_h_u_arrmul32_fa28_18_y2(h_u_arrmul32_and28_18_y0, h_u_arrmul32_fa29_17_y2, h_u_arrmul32_fa27_18_y4, h_u_arrmul32_fa28_18_y2, h_u_arrmul32_fa28_18_y4);
  and_gate and_gate_h_u_arrmul32_and29_18_y0(a_29, b_18, h_u_arrmul32_and29_18_y0);
  fa fa_h_u_arrmul32_fa29_18_y2(h_u_arrmul32_and29_18_y0, h_u_arrmul32_fa30_17_y2, h_u_arrmul32_fa28_18_y4, h_u_arrmul32_fa29_18_y2, h_u_arrmul32_fa29_18_y4);
  and_gate and_gate_h_u_arrmul32_and30_18_y0(a_30, b_18, h_u_arrmul32_and30_18_y0);
  fa fa_h_u_arrmul32_fa30_18_y2(h_u_arrmul32_and30_18_y0, h_u_arrmul32_fa31_17_y2, h_u_arrmul32_fa29_18_y4, h_u_arrmul32_fa30_18_y2, h_u_arrmul32_fa30_18_y4);
  and_gate and_gate_h_u_arrmul32_and31_18_y0(a_31, b_18, h_u_arrmul32_and31_18_y0);
  fa fa_h_u_arrmul32_fa31_18_y2(h_u_arrmul32_and31_18_y0, h_u_arrmul32_fa31_17_y4, h_u_arrmul32_fa30_18_y4, h_u_arrmul32_fa31_18_y2, h_u_arrmul32_fa31_18_y4);
  and_gate and_gate_h_u_arrmul32_and0_19_y0(a_0, b_19, h_u_arrmul32_and0_19_y0);
  ha ha_h_u_arrmul32_ha0_19_y0(h_u_arrmul32_and0_19_y0, h_u_arrmul32_fa1_18_y2, h_u_arrmul32_ha0_19_y0, h_u_arrmul32_ha0_19_y1);
  and_gate and_gate_h_u_arrmul32_and1_19_y0(a_1, b_19, h_u_arrmul32_and1_19_y0);
  fa fa_h_u_arrmul32_fa1_19_y2(h_u_arrmul32_and1_19_y0, h_u_arrmul32_fa2_18_y2, h_u_arrmul32_ha0_19_y1, h_u_arrmul32_fa1_19_y2, h_u_arrmul32_fa1_19_y4);
  and_gate and_gate_h_u_arrmul32_and2_19_y0(a_2, b_19, h_u_arrmul32_and2_19_y0);
  fa fa_h_u_arrmul32_fa2_19_y2(h_u_arrmul32_and2_19_y0, h_u_arrmul32_fa3_18_y2, h_u_arrmul32_fa1_19_y4, h_u_arrmul32_fa2_19_y2, h_u_arrmul32_fa2_19_y4);
  and_gate and_gate_h_u_arrmul32_and3_19_y0(a_3, b_19, h_u_arrmul32_and3_19_y0);
  fa fa_h_u_arrmul32_fa3_19_y2(h_u_arrmul32_and3_19_y0, h_u_arrmul32_fa4_18_y2, h_u_arrmul32_fa2_19_y4, h_u_arrmul32_fa3_19_y2, h_u_arrmul32_fa3_19_y4);
  and_gate and_gate_h_u_arrmul32_and4_19_y0(a_4, b_19, h_u_arrmul32_and4_19_y0);
  fa fa_h_u_arrmul32_fa4_19_y2(h_u_arrmul32_and4_19_y0, h_u_arrmul32_fa5_18_y2, h_u_arrmul32_fa3_19_y4, h_u_arrmul32_fa4_19_y2, h_u_arrmul32_fa4_19_y4);
  and_gate and_gate_h_u_arrmul32_and5_19_y0(a_5, b_19, h_u_arrmul32_and5_19_y0);
  fa fa_h_u_arrmul32_fa5_19_y2(h_u_arrmul32_and5_19_y0, h_u_arrmul32_fa6_18_y2, h_u_arrmul32_fa4_19_y4, h_u_arrmul32_fa5_19_y2, h_u_arrmul32_fa5_19_y4);
  and_gate and_gate_h_u_arrmul32_and6_19_y0(a_6, b_19, h_u_arrmul32_and6_19_y0);
  fa fa_h_u_arrmul32_fa6_19_y2(h_u_arrmul32_and6_19_y0, h_u_arrmul32_fa7_18_y2, h_u_arrmul32_fa5_19_y4, h_u_arrmul32_fa6_19_y2, h_u_arrmul32_fa6_19_y4);
  and_gate and_gate_h_u_arrmul32_and7_19_y0(a_7, b_19, h_u_arrmul32_and7_19_y0);
  fa fa_h_u_arrmul32_fa7_19_y2(h_u_arrmul32_and7_19_y0, h_u_arrmul32_fa8_18_y2, h_u_arrmul32_fa6_19_y4, h_u_arrmul32_fa7_19_y2, h_u_arrmul32_fa7_19_y4);
  and_gate and_gate_h_u_arrmul32_and8_19_y0(a_8, b_19, h_u_arrmul32_and8_19_y0);
  fa fa_h_u_arrmul32_fa8_19_y2(h_u_arrmul32_and8_19_y0, h_u_arrmul32_fa9_18_y2, h_u_arrmul32_fa7_19_y4, h_u_arrmul32_fa8_19_y2, h_u_arrmul32_fa8_19_y4);
  and_gate and_gate_h_u_arrmul32_and9_19_y0(a_9, b_19, h_u_arrmul32_and9_19_y0);
  fa fa_h_u_arrmul32_fa9_19_y2(h_u_arrmul32_and9_19_y0, h_u_arrmul32_fa10_18_y2, h_u_arrmul32_fa8_19_y4, h_u_arrmul32_fa9_19_y2, h_u_arrmul32_fa9_19_y4);
  and_gate and_gate_h_u_arrmul32_and10_19_y0(a_10, b_19, h_u_arrmul32_and10_19_y0);
  fa fa_h_u_arrmul32_fa10_19_y2(h_u_arrmul32_and10_19_y0, h_u_arrmul32_fa11_18_y2, h_u_arrmul32_fa9_19_y4, h_u_arrmul32_fa10_19_y2, h_u_arrmul32_fa10_19_y4);
  and_gate and_gate_h_u_arrmul32_and11_19_y0(a_11, b_19, h_u_arrmul32_and11_19_y0);
  fa fa_h_u_arrmul32_fa11_19_y2(h_u_arrmul32_and11_19_y0, h_u_arrmul32_fa12_18_y2, h_u_arrmul32_fa10_19_y4, h_u_arrmul32_fa11_19_y2, h_u_arrmul32_fa11_19_y4);
  and_gate and_gate_h_u_arrmul32_and12_19_y0(a_12, b_19, h_u_arrmul32_and12_19_y0);
  fa fa_h_u_arrmul32_fa12_19_y2(h_u_arrmul32_and12_19_y0, h_u_arrmul32_fa13_18_y2, h_u_arrmul32_fa11_19_y4, h_u_arrmul32_fa12_19_y2, h_u_arrmul32_fa12_19_y4);
  and_gate and_gate_h_u_arrmul32_and13_19_y0(a_13, b_19, h_u_arrmul32_and13_19_y0);
  fa fa_h_u_arrmul32_fa13_19_y2(h_u_arrmul32_and13_19_y0, h_u_arrmul32_fa14_18_y2, h_u_arrmul32_fa12_19_y4, h_u_arrmul32_fa13_19_y2, h_u_arrmul32_fa13_19_y4);
  and_gate and_gate_h_u_arrmul32_and14_19_y0(a_14, b_19, h_u_arrmul32_and14_19_y0);
  fa fa_h_u_arrmul32_fa14_19_y2(h_u_arrmul32_and14_19_y0, h_u_arrmul32_fa15_18_y2, h_u_arrmul32_fa13_19_y4, h_u_arrmul32_fa14_19_y2, h_u_arrmul32_fa14_19_y4);
  and_gate and_gate_h_u_arrmul32_and15_19_y0(a_15, b_19, h_u_arrmul32_and15_19_y0);
  fa fa_h_u_arrmul32_fa15_19_y2(h_u_arrmul32_and15_19_y0, h_u_arrmul32_fa16_18_y2, h_u_arrmul32_fa14_19_y4, h_u_arrmul32_fa15_19_y2, h_u_arrmul32_fa15_19_y4);
  and_gate and_gate_h_u_arrmul32_and16_19_y0(a_16, b_19, h_u_arrmul32_and16_19_y0);
  fa fa_h_u_arrmul32_fa16_19_y2(h_u_arrmul32_and16_19_y0, h_u_arrmul32_fa17_18_y2, h_u_arrmul32_fa15_19_y4, h_u_arrmul32_fa16_19_y2, h_u_arrmul32_fa16_19_y4);
  and_gate and_gate_h_u_arrmul32_and17_19_y0(a_17, b_19, h_u_arrmul32_and17_19_y0);
  fa fa_h_u_arrmul32_fa17_19_y2(h_u_arrmul32_and17_19_y0, h_u_arrmul32_fa18_18_y2, h_u_arrmul32_fa16_19_y4, h_u_arrmul32_fa17_19_y2, h_u_arrmul32_fa17_19_y4);
  and_gate and_gate_h_u_arrmul32_and18_19_y0(a_18, b_19, h_u_arrmul32_and18_19_y0);
  fa fa_h_u_arrmul32_fa18_19_y2(h_u_arrmul32_and18_19_y0, h_u_arrmul32_fa19_18_y2, h_u_arrmul32_fa17_19_y4, h_u_arrmul32_fa18_19_y2, h_u_arrmul32_fa18_19_y4);
  and_gate and_gate_h_u_arrmul32_and19_19_y0(a_19, b_19, h_u_arrmul32_and19_19_y0);
  fa fa_h_u_arrmul32_fa19_19_y2(h_u_arrmul32_and19_19_y0, h_u_arrmul32_fa20_18_y2, h_u_arrmul32_fa18_19_y4, h_u_arrmul32_fa19_19_y2, h_u_arrmul32_fa19_19_y4);
  and_gate and_gate_h_u_arrmul32_and20_19_y0(a_20, b_19, h_u_arrmul32_and20_19_y0);
  fa fa_h_u_arrmul32_fa20_19_y2(h_u_arrmul32_and20_19_y0, h_u_arrmul32_fa21_18_y2, h_u_arrmul32_fa19_19_y4, h_u_arrmul32_fa20_19_y2, h_u_arrmul32_fa20_19_y4);
  and_gate and_gate_h_u_arrmul32_and21_19_y0(a_21, b_19, h_u_arrmul32_and21_19_y0);
  fa fa_h_u_arrmul32_fa21_19_y2(h_u_arrmul32_and21_19_y0, h_u_arrmul32_fa22_18_y2, h_u_arrmul32_fa20_19_y4, h_u_arrmul32_fa21_19_y2, h_u_arrmul32_fa21_19_y4);
  and_gate and_gate_h_u_arrmul32_and22_19_y0(a_22, b_19, h_u_arrmul32_and22_19_y0);
  fa fa_h_u_arrmul32_fa22_19_y2(h_u_arrmul32_and22_19_y0, h_u_arrmul32_fa23_18_y2, h_u_arrmul32_fa21_19_y4, h_u_arrmul32_fa22_19_y2, h_u_arrmul32_fa22_19_y4);
  and_gate and_gate_h_u_arrmul32_and23_19_y0(a_23, b_19, h_u_arrmul32_and23_19_y0);
  fa fa_h_u_arrmul32_fa23_19_y2(h_u_arrmul32_and23_19_y0, h_u_arrmul32_fa24_18_y2, h_u_arrmul32_fa22_19_y4, h_u_arrmul32_fa23_19_y2, h_u_arrmul32_fa23_19_y4);
  and_gate and_gate_h_u_arrmul32_and24_19_y0(a_24, b_19, h_u_arrmul32_and24_19_y0);
  fa fa_h_u_arrmul32_fa24_19_y2(h_u_arrmul32_and24_19_y0, h_u_arrmul32_fa25_18_y2, h_u_arrmul32_fa23_19_y4, h_u_arrmul32_fa24_19_y2, h_u_arrmul32_fa24_19_y4);
  and_gate and_gate_h_u_arrmul32_and25_19_y0(a_25, b_19, h_u_arrmul32_and25_19_y0);
  fa fa_h_u_arrmul32_fa25_19_y2(h_u_arrmul32_and25_19_y0, h_u_arrmul32_fa26_18_y2, h_u_arrmul32_fa24_19_y4, h_u_arrmul32_fa25_19_y2, h_u_arrmul32_fa25_19_y4);
  and_gate and_gate_h_u_arrmul32_and26_19_y0(a_26, b_19, h_u_arrmul32_and26_19_y0);
  fa fa_h_u_arrmul32_fa26_19_y2(h_u_arrmul32_and26_19_y0, h_u_arrmul32_fa27_18_y2, h_u_arrmul32_fa25_19_y4, h_u_arrmul32_fa26_19_y2, h_u_arrmul32_fa26_19_y4);
  and_gate and_gate_h_u_arrmul32_and27_19_y0(a_27, b_19, h_u_arrmul32_and27_19_y0);
  fa fa_h_u_arrmul32_fa27_19_y2(h_u_arrmul32_and27_19_y0, h_u_arrmul32_fa28_18_y2, h_u_arrmul32_fa26_19_y4, h_u_arrmul32_fa27_19_y2, h_u_arrmul32_fa27_19_y4);
  and_gate and_gate_h_u_arrmul32_and28_19_y0(a_28, b_19, h_u_arrmul32_and28_19_y0);
  fa fa_h_u_arrmul32_fa28_19_y2(h_u_arrmul32_and28_19_y0, h_u_arrmul32_fa29_18_y2, h_u_arrmul32_fa27_19_y4, h_u_arrmul32_fa28_19_y2, h_u_arrmul32_fa28_19_y4);
  and_gate and_gate_h_u_arrmul32_and29_19_y0(a_29, b_19, h_u_arrmul32_and29_19_y0);
  fa fa_h_u_arrmul32_fa29_19_y2(h_u_arrmul32_and29_19_y0, h_u_arrmul32_fa30_18_y2, h_u_arrmul32_fa28_19_y4, h_u_arrmul32_fa29_19_y2, h_u_arrmul32_fa29_19_y4);
  and_gate and_gate_h_u_arrmul32_and30_19_y0(a_30, b_19, h_u_arrmul32_and30_19_y0);
  fa fa_h_u_arrmul32_fa30_19_y2(h_u_arrmul32_and30_19_y0, h_u_arrmul32_fa31_18_y2, h_u_arrmul32_fa29_19_y4, h_u_arrmul32_fa30_19_y2, h_u_arrmul32_fa30_19_y4);
  and_gate and_gate_h_u_arrmul32_and31_19_y0(a_31, b_19, h_u_arrmul32_and31_19_y0);
  fa fa_h_u_arrmul32_fa31_19_y2(h_u_arrmul32_and31_19_y0, h_u_arrmul32_fa31_18_y4, h_u_arrmul32_fa30_19_y4, h_u_arrmul32_fa31_19_y2, h_u_arrmul32_fa31_19_y4);
  and_gate and_gate_h_u_arrmul32_and0_20_y0(a_0, b_20, h_u_arrmul32_and0_20_y0);
  ha ha_h_u_arrmul32_ha0_20_y0(h_u_arrmul32_and0_20_y0, h_u_arrmul32_fa1_19_y2, h_u_arrmul32_ha0_20_y0, h_u_arrmul32_ha0_20_y1);
  and_gate and_gate_h_u_arrmul32_and1_20_y0(a_1, b_20, h_u_arrmul32_and1_20_y0);
  fa fa_h_u_arrmul32_fa1_20_y2(h_u_arrmul32_and1_20_y0, h_u_arrmul32_fa2_19_y2, h_u_arrmul32_ha0_20_y1, h_u_arrmul32_fa1_20_y2, h_u_arrmul32_fa1_20_y4);
  and_gate and_gate_h_u_arrmul32_and2_20_y0(a_2, b_20, h_u_arrmul32_and2_20_y0);
  fa fa_h_u_arrmul32_fa2_20_y2(h_u_arrmul32_and2_20_y0, h_u_arrmul32_fa3_19_y2, h_u_arrmul32_fa1_20_y4, h_u_arrmul32_fa2_20_y2, h_u_arrmul32_fa2_20_y4);
  and_gate and_gate_h_u_arrmul32_and3_20_y0(a_3, b_20, h_u_arrmul32_and3_20_y0);
  fa fa_h_u_arrmul32_fa3_20_y2(h_u_arrmul32_and3_20_y0, h_u_arrmul32_fa4_19_y2, h_u_arrmul32_fa2_20_y4, h_u_arrmul32_fa3_20_y2, h_u_arrmul32_fa3_20_y4);
  and_gate and_gate_h_u_arrmul32_and4_20_y0(a_4, b_20, h_u_arrmul32_and4_20_y0);
  fa fa_h_u_arrmul32_fa4_20_y2(h_u_arrmul32_and4_20_y0, h_u_arrmul32_fa5_19_y2, h_u_arrmul32_fa3_20_y4, h_u_arrmul32_fa4_20_y2, h_u_arrmul32_fa4_20_y4);
  and_gate and_gate_h_u_arrmul32_and5_20_y0(a_5, b_20, h_u_arrmul32_and5_20_y0);
  fa fa_h_u_arrmul32_fa5_20_y2(h_u_arrmul32_and5_20_y0, h_u_arrmul32_fa6_19_y2, h_u_arrmul32_fa4_20_y4, h_u_arrmul32_fa5_20_y2, h_u_arrmul32_fa5_20_y4);
  and_gate and_gate_h_u_arrmul32_and6_20_y0(a_6, b_20, h_u_arrmul32_and6_20_y0);
  fa fa_h_u_arrmul32_fa6_20_y2(h_u_arrmul32_and6_20_y0, h_u_arrmul32_fa7_19_y2, h_u_arrmul32_fa5_20_y4, h_u_arrmul32_fa6_20_y2, h_u_arrmul32_fa6_20_y4);
  and_gate and_gate_h_u_arrmul32_and7_20_y0(a_7, b_20, h_u_arrmul32_and7_20_y0);
  fa fa_h_u_arrmul32_fa7_20_y2(h_u_arrmul32_and7_20_y0, h_u_arrmul32_fa8_19_y2, h_u_arrmul32_fa6_20_y4, h_u_arrmul32_fa7_20_y2, h_u_arrmul32_fa7_20_y4);
  and_gate and_gate_h_u_arrmul32_and8_20_y0(a_8, b_20, h_u_arrmul32_and8_20_y0);
  fa fa_h_u_arrmul32_fa8_20_y2(h_u_arrmul32_and8_20_y0, h_u_arrmul32_fa9_19_y2, h_u_arrmul32_fa7_20_y4, h_u_arrmul32_fa8_20_y2, h_u_arrmul32_fa8_20_y4);
  and_gate and_gate_h_u_arrmul32_and9_20_y0(a_9, b_20, h_u_arrmul32_and9_20_y0);
  fa fa_h_u_arrmul32_fa9_20_y2(h_u_arrmul32_and9_20_y0, h_u_arrmul32_fa10_19_y2, h_u_arrmul32_fa8_20_y4, h_u_arrmul32_fa9_20_y2, h_u_arrmul32_fa9_20_y4);
  and_gate and_gate_h_u_arrmul32_and10_20_y0(a_10, b_20, h_u_arrmul32_and10_20_y0);
  fa fa_h_u_arrmul32_fa10_20_y2(h_u_arrmul32_and10_20_y0, h_u_arrmul32_fa11_19_y2, h_u_arrmul32_fa9_20_y4, h_u_arrmul32_fa10_20_y2, h_u_arrmul32_fa10_20_y4);
  and_gate and_gate_h_u_arrmul32_and11_20_y0(a_11, b_20, h_u_arrmul32_and11_20_y0);
  fa fa_h_u_arrmul32_fa11_20_y2(h_u_arrmul32_and11_20_y0, h_u_arrmul32_fa12_19_y2, h_u_arrmul32_fa10_20_y4, h_u_arrmul32_fa11_20_y2, h_u_arrmul32_fa11_20_y4);
  and_gate and_gate_h_u_arrmul32_and12_20_y0(a_12, b_20, h_u_arrmul32_and12_20_y0);
  fa fa_h_u_arrmul32_fa12_20_y2(h_u_arrmul32_and12_20_y0, h_u_arrmul32_fa13_19_y2, h_u_arrmul32_fa11_20_y4, h_u_arrmul32_fa12_20_y2, h_u_arrmul32_fa12_20_y4);
  and_gate and_gate_h_u_arrmul32_and13_20_y0(a_13, b_20, h_u_arrmul32_and13_20_y0);
  fa fa_h_u_arrmul32_fa13_20_y2(h_u_arrmul32_and13_20_y0, h_u_arrmul32_fa14_19_y2, h_u_arrmul32_fa12_20_y4, h_u_arrmul32_fa13_20_y2, h_u_arrmul32_fa13_20_y4);
  and_gate and_gate_h_u_arrmul32_and14_20_y0(a_14, b_20, h_u_arrmul32_and14_20_y0);
  fa fa_h_u_arrmul32_fa14_20_y2(h_u_arrmul32_and14_20_y0, h_u_arrmul32_fa15_19_y2, h_u_arrmul32_fa13_20_y4, h_u_arrmul32_fa14_20_y2, h_u_arrmul32_fa14_20_y4);
  and_gate and_gate_h_u_arrmul32_and15_20_y0(a_15, b_20, h_u_arrmul32_and15_20_y0);
  fa fa_h_u_arrmul32_fa15_20_y2(h_u_arrmul32_and15_20_y0, h_u_arrmul32_fa16_19_y2, h_u_arrmul32_fa14_20_y4, h_u_arrmul32_fa15_20_y2, h_u_arrmul32_fa15_20_y4);
  and_gate and_gate_h_u_arrmul32_and16_20_y0(a_16, b_20, h_u_arrmul32_and16_20_y0);
  fa fa_h_u_arrmul32_fa16_20_y2(h_u_arrmul32_and16_20_y0, h_u_arrmul32_fa17_19_y2, h_u_arrmul32_fa15_20_y4, h_u_arrmul32_fa16_20_y2, h_u_arrmul32_fa16_20_y4);
  and_gate and_gate_h_u_arrmul32_and17_20_y0(a_17, b_20, h_u_arrmul32_and17_20_y0);
  fa fa_h_u_arrmul32_fa17_20_y2(h_u_arrmul32_and17_20_y0, h_u_arrmul32_fa18_19_y2, h_u_arrmul32_fa16_20_y4, h_u_arrmul32_fa17_20_y2, h_u_arrmul32_fa17_20_y4);
  and_gate and_gate_h_u_arrmul32_and18_20_y0(a_18, b_20, h_u_arrmul32_and18_20_y0);
  fa fa_h_u_arrmul32_fa18_20_y2(h_u_arrmul32_and18_20_y0, h_u_arrmul32_fa19_19_y2, h_u_arrmul32_fa17_20_y4, h_u_arrmul32_fa18_20_y2, h_u_arrmul32_fa18_20_y4);
  and_gate and_gate_h_u_arrmul32_and19_20_y0(a_19, b_20, h_u_arrmul32_and19_20_y0);
  fa fa_h_u_arrmul32_fa19_20_y2(h_u_arrmul32_and19_20_y0, h_u_arrmul32_fa20_19_y2, h_u_arrmul32_fa18_20_y4, h_u_arrmul32_fa19_20_y2, h_u_arrmul32_fa19_20_y4);
  and_gate and_gate_h_u_arrmul32_and20_20_y0(a_20, b_20, h_u_arrmul32_and20_20_y0);
  fa fa_h_u_arrmul32_fa20_20_y2(h_u_arrmul32_and20_20_y0, h_u_arrmul32_fa21_19_y2, h_u_arrmul32_fa19_20_y4, h_u_arrmul32_fa20_20_y2, h_u_arrmul32_fa20_20_y4);
  and_gate and_gate_h_u_arrmul32_and21_20_y0(a_21, b_20, h_u_arrmul32_and21_20_y0);
  fa fa_h_u_arrmul32_fa21_20_y2(h_u_arrmul32_and21_20_y0, h_u_arrmul32_fa22_19_y2, h_u_arrmul32_fa20_20_y4, h_u_arrmul32_fa21_20_y2, h_u_arrmul32_fa21_20_y4);
  and_gate and_gate_h_u_arrmul32_and22_20_y0(a_22, b_20, h_u_arrmul32_and22_20_y0);
  fa fa_h_u_arrmul32_fa22_20_y2(h_u_arrmul32_and22_20_y0, h_u_arrmul32_fa23_19_y2, h_u_arrmul32_fa21_20_y4, h_u_arrmul32_fa22_20_y2, h_u_arrmul32_fa22_20_y4);
  and_gate and_gate_h_u_arrmul32_and23_20_y0(a_23, b_20, h_u_arrmul32_and23_20_y0);
  fa fa_h_u_arrmul32_fa23_20_y2(h_u_arrmul32_and23_20_y0, h_u_arrmul32_fa24_19_y2, h_u_arrmul32_fa22_20_y4, h_u_arrmul32_fa23_20_y2, h_u_arrmul32_fa23_20_y4);
  and_gate and_gate_h_u_arrmul32_and24_20_y0(a_24, b_20, h_u_arrmul32_and24_20_y0);
  fa fa_h_u_arrmul32_fa24_20_y2(h_u_arrmul32_and24_20_y0, h_u_arrmul32_fa25_19_y2, h_u_arrmul32_fa23_20_y4, h_u_arrmul32_fa24_20_y2, h_u_arrmul32_fa24_20_y4);
  and_gate and_gate_h_u_arrmul32_and25_20_y0(a_25, b_20, h_u_arrmul32_and25_20_y0);
  fa fa_h_u_arrmul32_fa25_20_y2(h_u_arrmul32_and25_20_y0, h_u_arrmul32_fa26_19_y2, h_u_arrmul32_fa24_20_y4, h_u_arrmul32_fa25_20_y2, h_u_arrmul32_fa25_20_y4);
  and_gate and_gate_h_u_arrmul32_and26_20_y0(a_26, b_20, h_u_arrmul32_and26_20_y0);
  fa fa_h_u_arrmul32_fa26_20_y2(h_u_arrmul32_and26_20_y0, h_u_arrmul32_fa27_19_y2, h_u_arrmul32_fa25_20_y4, h_u_arrmul32_fa26_20_y2, h_u_arrmul32_fa26_20_y4);
  and_gate and_gate_h_u_arrmul32_and27_20_y0(a_27, b_20, h_u_arrmul32_and27_20_y0);
  fa fa_h_u_arrmul32_fa27_20_y2(h_u_arrmul32_and27_20_y0, h_u_arrmul32_fa28_19_y2, h_u_arrmul32_fa26_20_y4, h_u_arrmul32_fa27_20_y2, h_u_arrmul32_fa27_20_y4);
  and_gate and_gate_h_u_arrmul32_and28_20_y0(a_28, b_20, h_u_arrmul32_and28_20_y0);
  fa fa_h_u_arrmul32_fa28_20_y2(h_u_arrmul32_and28_20_y0, h_u_arrmul32_fa29_19_y2, h_u_arrmul32_fa27_20_y4, h_u_arrmul32_fa28_20_y2, h_u_arrmul32_fa28_20_y4);
  and_gate and_gate_h_u_arrmul32_and29_20_y0(a_29, b_20, h_u_arrmul32_and29_20_y0);
  fa fa_h_u_arrmul32_fa29_20_y2(h_u_arrmul32_and29_20_y0, h_u_arrmul32_fa30_19_y2, h_u_arrmul32_fa28_20_y4, h_u_arrmul32_fa29_20_y2, h_u_arrmul32_fa29_20_y4);
  and_gate and_gate_h_u_arrmul32_and30_20_y0(a_30, b_20, h_u_arrmul32_and30_20_y0);
  fa fa_h_u_arrmul32_fa30_20_y2(h_u_arrmul32_and30_20_y0, h_u_arrmul32_fa31_19_y2, h_u_arrmul32_fa29_20_y4, h_u_arrmul32_fa30_20_y2, h_u_arrmul32_fa30_20_y4);
  and_gate and_gate_h_u_arrmul32_and31_20_y0(a_31, b_20, h_u_arrmul32_and31_20_y0);
  fa fa_h_u_arrmul32_fa31_20_y2(h_u_arrmul32_and31_20_y0, h_u_arrmul32_fa31_19_y4, h_u_arrmul32_fa30_20_y4, h_u_arrmul32_fa31_20_y2, h_u_arrmul32_fa31_20_y4);
  and_gate and_gate_h_u_arrmul32_and0_21_y0(a_0, b_21, h_u_arrmul32_and0_21_y0);
  ha ha_h_u_arrmul32_ha0_21_y0(h_u_arrmul32_and0_21_y0, h_u_arrmul32_fa1_20_y2, h_u_arrmul32_ha0_21_y0, h_u_arrmul32_ha0_21_y1);
  and_gate and_gate_h_u_arrmul32_and1_21_y0(a_1, b_21, h_u_arrmul32_and1_21_y0);
  fa fa_h_u_arrmul32_fa1_21_y2(h_u_arrmul32_and1_21_y0, h_u_arrmul32_fa2_20_y2, h_u_arrmul32_ha0_21_y1, h_u_arrmul32_fa1_21_y2, h_u_arrmul32_fa1_21_y4);
  and_gate and_gate_h_u_arrmul32_and2_21_y0(a_2, b_21, h_u_arrmul32_and2_21_y0);
  fa fa_h_u_arrmul32_fa2_21_y2(h_u_arrmul32_and2_21_y0, h_u_arrmul32_fa3_20_y2, h_u_arrmul32_fa1_21_y4, h_u_arrmul32_fa2_21_y2, h_u_arrmul32_fa2_21_y4);
  and_gate and_gate_h_u_arrmul32_and3_21_y0(a_3, b_21, h_u_arrmul32_and3_21_y0);
  fa fa_h_u_arrmul32_fa3_21_y2(h_u_arrmul32_and3_21_y0, h_u_arrmul32_fa4_20_y2, h_u_arrmul32_fa2_21_y4, h_u_arrmul32_fa3_21_y2, h_u_arrmul32_fa3_21_y4);
  and_gate and_gate_h_u_arrmul32_and4_21_y0(a_4, b_21, h_u_arrmul32_and4_21_y0);
  fa fa_h_u_arrmul32_fa4_21_y2(h_u_arrmul32_and4_21_y0, h_u_arrmul32_fa5_20_y2, h_u_arrmul32_fa3_21_y4, h_u_arrmul32_fa4_21_y2, h_u_arrmul32_fa4_21_y4);
  and_gate and_gate_h_u_arrmul32_and5_21_y0(a_5, b_21, h_u_arrmul32_and5_21_y0);
  fa fa_h_u_arrmul32_fa5_21_y2(h_u_arrmul32_and5_21_y0, h_u_arrmul32_fa6_20_y2, h_u_arrmul32_fa4_21_y4, h_u_arrmul32_fa5_21_y2, h_u_arrmul32_fa5_21_y4);
  and_gate and_gate_h_u_arrmul32_and6_21_y0(a_6, b_21, h_u_arrmul32_and6_21_y0);
  fa fa_h_u_arrmul32_fa6_21_y2(h_u_arrmul32_and6_21_y0, h_u_arrmul32_fa7_20_y2, h_u_arrmul32_fa5_21_y4, h_u_arrmul32_fa6_21_y2, h_u_arrmul32_fa6_21_y4);
  and_gate and_gate_h_u_arrmul32_and7_21_y0(a_7, b_21, h_u_arrmul32_and7_21_y0);
  fa fa_h_u_arrmul32_fa7_21_y2(h_u_arrmul32_and7_21_y0, h_u_arrmul32_fa8_20_y2, h_u_arrmul32_fa6_21_y4, h_u_arrmul32_fa7_21_y2, h_u_arrmul32_fa7_21_y4);
  and_gate and_gate_h_u_arrmul32_and8_21_y0(a_8, b_21, h_u_arrmul32_and8_21_y0);
  fa fa_h_u_arrmul32_fa8_21_y2(h_u_arrmul32_and8_21_y0, h_u_arrmul32_fa9_20_y2, h_u_arrmul32_fa7_21_y4, h_u_arrmul32_fa8_21_y2, h_u_arrmul32_fa8_21_y4);
  and_gate and_gate_h_u_arrmul32_and9_21_y0(a_9, b_21, h_u_arrmul32_and9_21_y0);
  fa fa_h_u_arrmul32_fa9_21_y2(h_u_arrmul32_and9_21_y0, h_u_arrmul32_fa10_20_y2, h_u_arrmul32_fa8_21_y4, h_u_arrmul32_fa9_21_y2, h_u_arrmul32_fa9_21_y4);
  and_gate and_gate_h_u_arrmul32_and10_21_y0(a_10, b_21, h_u_arrmul32_and10_21_y0);
  fa fa_h_u_arrmul32_fa10_21_y2(h_u_arrmul32_and10_21_y0, h_u_arrmul32_fa11_20_y2, h_u_arrmul32_fa9_21_y4, h_u_arrmul32_fa10_21_y2, h_u_arrmul32_fa10_21_y4);
  and_gate and_gate_h_u_arrmul32_and11_21_y0(a_11, b_21, h_u_arrmul32_and11_21_y0);
  fa fa_h_u_arrmul32_fa11_21_y2(h_u_arrmul32_and11_21_y0, h_u_arrmul32_fa12_20_y2, h_u_arrmul32_fa10_21_y4, h_u_arrmul32_fa11_21_y2, h_u_arrmul32_fa11_21_y4);
  and_gate and_gate_h_u_arrmul32_and12_21_y0(a_12, b_21, h_u_arrmul32_and12_21_y0);
  fa fa_h_u_arrmul32_fa12_21_y2(h_u_arrmul32_and12_21_y0, h_u_arrmul32_fa13_20_y2, h_u_arrmul32_fa11_21_y4, h_u_arrmul32_fa12_21_y2, h_u_arrmul32_fa12_21_y4);
  and_gate and_gate_h_u_arrmul32_and13_21_y0(a_13, b_21, h_u_arrmul32_and13_21_y0);
  fa fa_h_u_arrmul32_fa13_21_y2(h_u_arrmul32_and13_21_y0, h_u_arrmul32_fa14_20_y2, h_u_arrmul32_fa12_21_y4, h_u_arrmul32_fa13_21_y2, h_u_arrmul32_fa13_21_y4);
  and_gate and_gate_h_u_arrmul32_and14_21_y0(a_14, b_21, h_u_arrmul32_and14_21_y0);
  fa fa_h_u_arrmul32_fa14_21_y2(h_u_arrmul32_and14_21_y0, h_u_arrmul32_fa15_20_y2, h_u_arrmul32_fa13_21_y4, h_u_arrmul32_fa14_21_y2, h_u_arrmul32_fa14_21_y4);
  and_gate and_gate_h_u_arrmul32_and15_21_y0(a_15, b_21, h_u_arrmul32_and15_21_y0);
  fa fa_h_u_arrmul32_fa15_21_y2(h_u_arrmul32_and15_21_y0, h_u_arrmul32_fa16_20_y2, h_u_arrmul32_fa14_21_y4, h_u_arrmul32_fa15_21_y2, h_u_arrmul32_fa15_21_y4);
  and_gate and_gate_h_u_arrmul32_and16_21_y0(a_16, b_21, h_u_arrmul32_and16_21_y0);
  fa fa_h_u_arrmul32_fa16_21_y2(h_u_arrmul32_and16_21_y0, h_u_arrmul32_fa17_20_y2, h_u_arrmul32_fa15_21_y4, h_u_arrmul32_fa16_21_y2, h_u_arrmul32_fa16_21_y4);
  and_gate and_gate_h_u_arrmul32_and17_21_y0(a_17, b_21, h_u_arrmul32_and17_21_y0);
  fa fa_h_u_arrmul32_fa17_21_y2(h_u_arrmul32_and17_21_y0, h_u_arrmul32_fa18_20_y2, h_u_arrmul32_fa16_21_y4, h_u_arrmul32_fa17_21_y2, h_u_arrmul32_fa17_21_y4);
  and_gate and_gate_h_u_arrmul32_and18_21_y0(a_18, b_21, h_u_arrmul32_and18_21_y0);
  fa fa_h_u_arrmul32_fa18_21_y2(h_u_arrmul32_and18_21_y0, h_u_arrmul32_fa19_20_y2, h_u_arrmul32_fa17_21_y4, h_u_arrmul32_fa18_21_y2, h_u_arrmul32_fa18_21_y4);
  and_gate and_gate_h_u_arrmul32_and19_21_y0(a_19, b_21, h_u_arrmul32_and19_21_y0);
  fa fa_h_u_arrmul32_fa19_21_y2(h_u_arrmul32_and19_21_y0, h_u_arrmul32_fa20_20_y2, h_u_arrmul32_fa18_21_y4, h_u_arrmul32_fa19_21_y2, h_u_arrmul32_fa19_21_y4);
  and_gate and_gate_h_u_arrmul32_and20_21_y0(a_20, b_21, h_u_arrmul32_and20_21_y0);
  fa fa_h_u_arrmul32_fa20_21_y2(h_u_arrmul32_and20_21_y0, h_u_arrmul32_fa21_20_y2, h_u_arrmul32_fa19_21_y4, h_u_arrmul32_fa20_21_y2, h_u_arrmul32_fa20_21_y4);
  and_gate and_gate_h_u_arrmul32_and21_21_y0(a_21, b_21, h_u_arrmul32_and21_21_y0);
  fa fa_h_u_arrmul32_fa21_21_y2(h_u_arrmul32_and21_21_y0, h_u_arrmul32_fa22_20_y2, h_u_arrmul32_fa20_21_y4, h_u_arrmul32_fa21_21_y2, h_u_arrmul32_fa21_21_y4);
  and_gate and_gate_h_u_arrmul32_and22_21_y0(a_22, b_21, h_u_arrmul32_and22_21_y0);
  fa fa_h_u_arrmul32_fa22_21_y2(h_u_arrmul32_and22_21_y0, h_u_arrmul32_fa23_20_y2, h_u_arrmul32_fa21_21_y4, h_u_arrmul32_fa22_21_y2, h_u_arrmul32_fa22_21_y4);
  and_gate and_gate_h_u_arrmul32_and23_21_y0(a_23, b_21, h_u_arrmul32_and23_21_y0);
  fa fa_h_u_arrmul32_fa23_21_y2(h_u_arrmul32_and23_21_y0, h_u_arrmul32_fa24_20_y2, h_u_arrmul32_fa22_21_y4, h_u_arrmul32_fa23_21_y2, h_u_arrmul32_fa23_21_y4);
  and_gate and_gate_h_u_arrmul32_and24_21_y0(a_24, b_21, h_u_arrmul32_and24_21_y0);
  fa fa_h_u_arrmul32_fa24_21_y2(h_u_arrmul32_and24_21_y0, h_u_arrmul32_fa25_20_y2, h_u_arrmul32_fa23_21_y4, h_u_arrmul32_fa24_21_y2, h_u_arrmul32_fa24_21_y4);
  and_gate and_gate_h_u_arrmul32_and25_21_y0(a_25, b_21, h_u_arrmul32_and25_21_y0);
  fa fa_h_u_arrmul32_fa25_21_y2(h_u_arrmul32_and25_21_y0, h_u_arrmul32_fa26_20_y2, h_u_arrmul32_fa24_21_y4, h_u_arrmul32_fa25_21_y2, h_u_arrmul32_fa25_21_y4);
  and_gate and_gate_h_u_arrmul32_and26_21_y0(a_26, b_21, h_u_arrmul32_and26_21_y0);
  fa fa_h_u_arrmul32_fa26_21_y2(h_u_arrmul32_and26_21_y0, h_u_arrmul32_fa27_20_y2, h_u_arrmul32_fa25_21_y4, h_u_arrmul32_fa26_21_y2, h_u_arrmul32_fa26_21_y4);
  and_gate and_gate_h_u_arrmul32_and27_21_y0(a_27, b_21, h_u_arrmul32_and27_21_y0);
  fa fa_h_u_arrmul32_fa27_21_y2(h_u_arrmul32_and27_21_y0, h_u_arrmul32_fa28_20_y2, h_u_arrmul32_fa26_21_y4, h_u_arrmul32_fa27_21_y2, h_u_arrmul32_fa27_21_y4);
  and_gate and_gate_h_u_arrmul32_and28_21_y0(a_28, b_21, h_u_arrmul32_and28_21_y0);
  fa fa_h_u_arrmul32_fa28_21_y2(h_u_arrmul32_and28_21_y0, h_u_arrmul32_fa29_20_y2, h_u_arrmul32_fa27_21_y4, h_u_arrmul32_fa28_21_y2, h_u_arrmul32_fa28_21_y4);
  and_gate and_gate_h_u_arrmul32_and29_21_y0(a_29, b_21, h_u_arrmul32_and29_21_y0);
  fa fa_h_u_arrmul32_fa29_21_y2(h_u_arrmul32_and29_21_y0, h_u_arrmul32_fa30_20_y2, h_u_arrmul32_fa28_21_y4, h_u_arrmul32_fa29_21_y2, h_u_arrmul32_fa29_21_y4);
  and_gate and_gate_h_u_arrmul32_and30_21_y0(a_30, b_21, h_u_arrmul32_and30_21_y0);
  fa fa_h_u_arrmul32_fa30_21_y2(h_u_arrmul32_and30_21_y0, h_u_arrmul32_fa31_20_y2, h_u_arrmul32_fa29_21_y4, h_u_arrmul32_fa30_21_y2, h_u_arrmul32_fa30_21_y4);
  and_gate and_gate_h_u_arrmul32_and31_21_y0(a_31, b_21, h_u_arrmul32_and31_21_y0);
  fa fa_h_u_arrmul32_fa31_21_y2(h_u_arrmul32_and31_21_y0, h_u_arrmul32_fa31_20_y4, h_u_arrmul32_fa30_21_y4, h_u_arrmul32_fa31_21_y2, h_u_arrmul32_fa31_21_y4);
  and_gate and_gate_h_u_arrmul32_and0_22_y0(a_0, b_22, h_u_arrmul32_and0_22_y0);
  ha ha_h_u_arrmul32_ha0_22_y0(h_u_arrmul32_and0_22_y0, h_u_arrmul32_fa1_21_y2, h_u_arrmul32_ha0_22_y0, h_u_arrmul32_ha0_22_y1);
  and_gate and_gate_h_u_arrmul32_and1_22_y0(a_1, b_22, h_u_arrmul32_and1_22_y0);
  fa fa_h_u_arrmul32_fa1_22_y2(h_u_arrmul32_and1_22_y0, h_u_arrmul32_fa2_21_y2, h_u_arrmul32_ha0_22_y1, h_u_arrmul32_fa1_22_y2, h_u_arrmul32_fa1_22_y4);
  and_gate and_gate_h_u_arrmul32_and2_22_y0(a_2, b_22, h_u_arrmul32_and2_22_y0);
  fa fa_h_u_arrmul32_fa2_22_y2(h_u_arrmul32_and2_22_y0, h_u_arrmul32_fa3_21_y2, h_u_arrmul32_fa1_22_y4, h_u_arrmul32_fa2_22_y2, h_u_arrmul32_fa2_22_y4);
  and_gate and_gate_h_u_arrmul32_and3_22_y0(a_3, b_22, h_u_arrmul32_and3_22_y0);
  fa fa_h_u_arrmul32_fa3_22_y2(h_u_arrmul32_and3_22_y0, h_u_arrmul32_fa4_21_y2, h_u_arrmul32_fa2_22_y4, h_u_arrmul32_fa3_22_y2, h_u_arrmul32_fa3_22_y4);
  and_gate and_gate_h_u_arrmul32_and4_22_y0(a_4, b_22, h_u_arrmul32_and4_22_y0);
  fa fa_h_u_arrmul32_fa4_22_y2(h_u_arrmul32_and4_22_y0, h_u_arrmul32_fa5_21_y2, h_u_arrmul32_fa3_22_y4, h_u_arrmul32_fa4_22_y2, h_u_arrmul32_fa4_22_y4);
  and_gate and_gate_h_u_arrmul32_and5_22_y0(a_5, b_22, h_u_arrmul32_and5_22_y0);
  fa fa_h_u_arrmul32_fa5_22_y2(h_u_arrmul32_and5_22_y0, h_u_arrmul32_fa6_21_y2, h_u_arrmul32_fa4_22_y4, h_u_arrmul32_fa5_22_y2, h_u_arrmul32_fa5_22_y4);
  and_gate and_gate_h_u_arrmul32_and6_22_y0(a_6, b_22, h_u_arrmul32_and6_22_y0);
  fa fa_h_u_arrmul32_fa6_22_y2(h_u_arrmul32_and6_22_y0, h_u_arrmul32_fa7_21_y2, h_u_arrmul32_fa5_22_y4, h_u_arrmul32_fa6_22_y2, h_u_arrmul32_fa6_22_y4);
  and_gate and_gate_h_u_arrmul32_and7_22_y0(a_7, b_22, h_u_arrmul32_and7_22_y0);
  fa fa_h_u_arrmul32_fa7_22_y2(h_u_arrmul32_and7_22_y0, h_u_arrmul32_fa8_21_y2, h_u_arrmul32_fa6_22_y4, h_u_arrmul32_fa7_22_y2, h_u_arrmul32_fa7_22_y4);
  and_gate and_gate_h_u_arrmul32_and8_22_y0(a_8, b_22, h_u_arrmul32_and8_22_y0);
  fa fa_h_u_arrmul32_fa8_22_y2(h_u_arrmul32_and8_22_y0, h_u_arrmul32_fa9_21_y2, h_u_arrmul32_fa7_22_y4, h_u_arrmul32_fa8_22_y2, h_u_arrmul32_fa8_22_y4);
  and_gate and_gate_h_u_arrmul32_and9_22_y0(a_9, b_22, h_u_arrmul32_and9_22_y0);
  fa fa_h_u_arrmul32_fa9_22_y2(h_u_arrmul32_and9_22_y0, h_u_arrmul32_fa10_21_y2, h_u_arrmul32_fa8_22_y4, h_u_arrmul32_fa9_22_y2, h_u_arrmul32_fa9_22_y4);
  and_gate and_gate_h_u_arrmul32_and10_22_y0(a_10, b_22, h_u_arrmul32_and10_22_y0);
  fa fa_h_u_arrmul32_fa10_22_y2(h_u_arrmul32_and10_22_y0, h_u_arrmul32_fa11_21_y2, h_u_arrmul32_fa9_22_y4, h_u_arrmul32_fa10_22_y2, h_u_arrmul32_fa10_22_y4);
  and_gate and_gate_h_u_arrmul32_and11_22_y0(a_11, b_22, h_u_arrmul32_and11_22_y0);
  fa fa_h_u_arrmul32_fa11_22_y2(h_u_arrmul32_and11_22_y0, h_u_arrmul32_fa12_21_y2, h_u_arrmul32_fa10_22_y4, h_u_arrmul32_fa11_22_y2, h_u_arrmul32_fa11_22_y4);
  and_gate and_gate_h_u_arrmul32_and12_22_y0(a_12, b_22, h_u_arrmul32_and12_22_y0);
  fa fa_h_u_arrmul32_fa12_22_y2(h_u_arrmul32_and12_22_y0, h_u_arrmul32_fa13_21_y2, h_u_arrmul32_fa11_22_y4, h_u_arrmul32_fa12_22_y2, h_u_arrmul32_fa12_22_y4);
  and_gate and_gate_h_u_arrmul32_and13_22_y0(a_13, b_22, h_u_arrmul32_and13_22_y0);
  fa fa_h_u_arrmul32_fa13_22_y2(h_u_arrmul32_and13_22_y0, h_u_arrmul32_fa14_21_y2, h_u_arrmul32_fa12_22_y4, h_u_arrmul32_fa13_22_y2, h_u_arrmul32_fa13_22_y4);
  and_gate and_gate_h_u_arrmul32_and14_22_y0(a_14, b_22, h_u_arrmul32_and14_22_y0);
  fa fa_h_u_arrmul32_fa14_22_y2(h_u_arrmul32_and14_22_y0, h_u_arrmul32_fa15_21_y2, h_u_arrmul32_fa13_22_y4, h_u_arrmul32_fa14_22_y2, h_u_arrmul32_fa14_22_y4);
  and_gate and_gate_h_u_arrmul32_and15_22_y0(a_15, b_22, h_u_arrmul32_and15_22_y0);
  fa fa_h_u_arrmul32_fa15_22_y2(h_u_arrmul32_and15_22_y0, h_u_arrmul32_fa16_21_y2, h_u_arrmul32_fa14_22_y4, h_u_arrmul32_fa15_22_y2, h_u_arrmul32_fa15_22_y4);
  and_gate and_gate_h_u_arrmul32_and16_22_y0(a_16, b_22, h_u_arrmul32_and16_22_y0);
  fa fa_h_u_arrmul32_fa16_22_y2(h_u_arrmul32_and16_22_y0, h_u_arrmul32_fa17_21_y2, h_u_arrmul32_fa15_22_y4, h_u_arrmul32_fa16_22_y2, h_u_arrmul32_fa16_22_y4);
  and_gate and_gate_h_u_arrmul32_and17_22_y0(a_17, b_22, h_u_arrmul32_and17_22_y0);
  fa fa_h_u_arrmul32_fa17_22_y2(h_u_arrmul32_and17_22_y0, h_u_arrmul32_fa18_21_y2, h_u_arrmul32_fa16_22_y4, h_u_arrmul32_fa17_22_y2, h_u_arrmul32_fa17_22_y4);
  and_gate and_gate_h_u_arrmul32_and18_22_y0(a_18, b_22, h_u_arrmul32_and18_22_y0);
  fa fa_h_u_arrmul32_fa18_22_y2(h_u_arrmul32_and18_22_y0, h_u_arrmul32_fa19_21_y2, h_u_arrmul32_fa17_22_y4, h_u_arrmul32_fa18_22_y2, h_u_arrmul32_fa18_22_y4);
  and_gate and_gate_h_u_arrmul32_and19_22_y0(a_19, b_22, h_u_arrmul32_and19_22_y0);
  fa fa_h_u_arrmul32_fa19_22_y2(h_u_arrmul32_and19_22_y0, h_u_arrmul32_fa20_21_y2, h_u_arrmul32_fa18_22_y4, h_u_arrmul32_fa19_22_y2, h_u_arrmul32_fa19_22_y4);
  and_gate and_gate_h_u_arrmul32_and20_22_y0(a_20, b_22, h_u_arrmul32_and20_22_y0);
  fa fa_h_u_arrmul32_fa20_22_y2(h_u_arrmul32_and20_22_y0, h_u_arrmul32_fa21_21_y2, h_u_arrmul32_fa19_22_y4, h_u_arrmul32_fa20_22_y2, h_u_arrmul32_fa20_22_y4);
  and_gate and_gate_h_u_arrmul32_and21_22_y0(a_21, b_22, h_u_arrmul32_and21_22_y0);
  fa fa_h_u_arrmul32_fa21_22_y2(h_u_arrmul32_and21_22_y0, h_u_arrmul32_fa22_21_y2, h_u_arrmul32_fa20_22_y4, h_u_arrmul32_fa21_22_y2, h_u_arrmul32_fa21_22_y4);
  and_gate and_gate_h_u_arrmul32_and22_22_y0(a_22, b_22, h_u_arrmul32_and22_22_y0);
  fa fa_h_u_arrmul32_fa22_22_y2(h_u_arrmul32_and22_22_y0, h_u_arrmul32_fa23_21_y2, h_u_arrmul32_fa21_22_y4, h_u_arrmul32_fa22_22_y2, h_u_arrmul32_fa22_22_y4);
  and_gate and_gate_h_u_arrmul32_and23_22_y0(a_23, b_22, h_u_arrmul32_and23_22_y0);
  fa fa_h_u_arrmul32_fa23_22_y2(h_u_arrmul32_and23_22_y0, h_u_arrmul32_fa24_21_y2, h_u_arrmul32_fa22_22_y4, h_u_arrmul32_fa23_22_y2, h_u_arrmul32_fa23_22_y4);
  and_gate and_gate_h_u_arrmul32_and24_22_y0(a_24, b_22, h_u_arrmul32_and24_22_y0);
  fa fa_h_u_arrmul32_fa24_22_y2(h_u_arrmul32_and24_22_y0, h_u_arrmul32_fa25_21_y2, h_u_arrmul32_fa23_22_y4, h_u_arrmul32_fa24_22_y2, h_u_arrmul32_fa24_22_y4);
  and_gate and_gate_h_u_arrmul32_and25_22_y0(a_25, b_22, h_u_arrmul32_and25_22_y0);
  fa fa_h_u_arrmul32_fa25_22_y2(h_u_arrmul32_and25_22_y0, h_u_arrmul32_fa26_21_y2, h_u_arrmul32_fa24_22_y4, h_u_arrmul32_fa25_22_y2, h_u_arrmul32_fa25_22_y4);
  and_gate and_gate_h_u_arrmul32_and26_22_y0(a_26, b_22, h_u_arrmul32_and26_22_y0);
  fa fa_h_u_arrmul32_fa26_22_y2(h_u_arrmul32_and26_22_y0, h_u_arrmul32_fa27_21_y2, h_u_arrmul32_fa25_22_y4, h_u_arrmul32_fa26_22_y2, h_u_arrmul32_fa26_22_y4);
  and_gate and_gate_h_u_arrmul32_and27_22_y0(a_27, b_22, h_u_arrmul32_and27_22_y0);
  fa fa_h_u_arrmul32_fa27_22_y2(h_u_arrmul32_and27_22_y0, h_u_arrmul32_fa28_21_y2, h_u_arrmul32_fa26_22_y4, h_u_arrmul32_fa27_22_y2, h_u_arrmul32_fa27_22_y4);
  and_gate and_gate_h_u_arrmul32_and28_22_y0(a_28, b_22, h_u_arrmul32_and28_22_y0);
  fa fa_h_u_arrmul32_fa28_22_y2(h_u_arrmul32_and28_22_y0, h_u_arrmul32_fa29_21_y2, h_u_arrmul32_fa27_22_y4, h_u_arrmul32_fa28_22_y2, h_u_arrmul32_fa28_22_y4);
  and_gate and_gate_h_u_arrmul32_and29_22_y0(a_29, b_22, h_u_arrmul32_and29_22_y0);
  fa fa_h_u_arrmul32_fa29_22_y2(h_u_arrmul32_and29_22_y0, h_u_arrmul32_fa30_21_y2, h_u_arrmul32_fa28_22_y4, h_u_arrmul32_fa29_22_y2, h_u_arrmul32_fa29_22_y4);
  and_gate and_gate_h_u_arrmul32_and30_22_y0(a_30, b_22, h_u_arrmul32_and30_22_y0);
  fa fa_h_u_arrmul32_fa30_22_y2(h_u_arrmul32_and30_22_y0, h_u_arrmul32_fa31_21_y2, h_u_arrmul32_fa29_22_y4, h_u_arrmul32_fa30_22_y2, h_u_arrmul32_fa30_22_y4);
  and_gate and_gate_h_u_arrmul32_and31_22_y0(a_31, b_22, h_u_arrmul32_and31_22_y0);
  fa fa_h_u_arrmul32_fa31_22_y2(h_u_arrmul32_and31_22_y0, h_u_arrmul32_fa31_21_y4, h_u_arrmul32_fa30_22_y4, h_u_arrmul32_fa31_22_y2, h_u_arrmul32_fa31_22_y4);
  and_gate and_gate_h_u_arrmul32_and0_23_y0(a_0, b_23, h_u_arrmul32_and0_23_y0);
  ha ha_h_u_arrmul32_ha0_23_y0(h_u_arrmul32_and0_23_y0, h_u_arrmul32_fa1_22_y2, h_u_arrmul32_ha0_23_y0, h_u_arrmul32_ha0_23_y1);
  and_gate and_gate_h_u_arrmul32_and1_23_y0(a_1, b_23, h_u_arrmul32_and1_23_y0);
  fa fa_h_u_arrmul32_fa1_23_y2(h_u_arrmul32_and1_23_y0, h_u_arrmul32_fa2_22_y2, h_u_arrmul32_ha0_23_y1, h_u_arrmul32_fa1_23_y2, h_u_arrmul32_fa1_23_y4);
  and_gate and_gate_h_u_arrmul32_and2_23_y0(a_2, b_23, h_u_arrmul32_and2_23_y0);
  fa fa_h_u_arrmul32_fa2_23_y2(h_u_arrmul32_and2_23_y0, h_u_arrmul32_fa3_22_y2, h_u_arrmul32_fa1_23_y4, h_u_arrmul32_fa2_23_y2, h_u_arrmul32_fa2_23_y4);
  and_gate and_gate_h_u_arrmul32_and3_23_y0(a_3, b_23, h_u_arrmul32_and3_23_y0);
  fa fa_h_u_arrmul32_fa3_23_y2(h_u_arrmul32_and3_23_y0, h_u_arrmul32_fa4_22_y2, h_u_arrmul32_fa2_23_y4, h_u_arrmul32_fa3_23_y2, h_u_arrmul32_fa3_23_y4);
  and_gate and_gate_h_u_arrmul32_and4_23_y0(a_4, b_23, h_u_arrmul32_and4_23_y0);
  fa fa_h_u_arrmul32_fa4_23_y2(h_u_arrmul32_and4_23_y0, h_u_arrmul32_fa5_22_y2, h_u_arrmul32_fa3_23_y4, h_u_arrmul32_fa4_23_y2, h_u_arrmul32_fa4_23_y4);
  and_gate and_gate_h_u_arrmul32_and5_23_y0(a_5, b_23, h_u_arrmul32_and5_23_y0);
  fa fa_h_u_arrmul32_fa5_23_y2(h_u_arrmul32_and5_23_y0, h_u_arrmul32_fa6_22_y2, h_u_arrmul32_fa4_23_y4, h_u_arrmul32_fa5_23_y2, h_u_arrmul32_fa5_23_y4);
  and_gate and_gate_h_u_arrmul32_and6_23_y0(a_6, b_23, h_u_arrmul32_and6_23_y0);
  fa fa_h_u_arrmul32_fa6_23_y2(h_u_arrmul32_and6_23_y0, h_u_arrmul32_fa7_22_y2, h_u_arrmul32_fa5_23_y4, h_u_arrmul32_fa6_23_y2, h_u_arrmul32_fa6_23_y4);
  and_gate and_gate_h_u_arrmul32_and7_23_y0(a_7, b_23, h_u_arrmul32_and7_23_y0);
  fa fa_h_u_arrmul32_fa7_23_y2(h_u_arrmul32_and7_23_y0, h_u_arrmul32_fa8_22_y2, h_u_arrmul32_fa6_23_y4, h_u_arrmul32_fa7_23_y2, h_u_arrmul32_fa7_23_y4);
  and_gate and_gate_h_u_arrmul32_and8_23_y0(a_8, b_23, h_u_arrmul32_and8_23_y0);
  fa fa_h_u_arrmul32_fa8_23_y2(h_u_arrmul32_and8_23_y0, h_u_arrmul32_fa9_22_y2, h_u_arrmul32_fa7_23_y4, h_u_arrmul32_fa8_23_y2, h_u_arrmul32_fa8_23_y4);
  and_gate and_gate_h_u_arrmul32_and9_23_y0(a_9, b_23, h_u_arrmul32_and9_23_y0);
  fa fa_h_u_arrmul32_fa9_23_y2(h_u_arrmul32_and9_23_y0, h_u_arrmul32_fa10_22_y2, h_u_arrmul32_fa8_23_y4, h_u_arrmul32_fa9_23_y2, h_u_arrmul32_fa9_23_y4);
  and_gate and_gate_h_u_arrmul32_and10_23_y0(a_10, b_23, h_u_arrmul32_and10_23_y0);
  fa fa_h_u_arrmul32_fa10_23_y2(h_u_arrmul32_and10_23_y0, h_u_arrmul32_fa11_22_y2, h_u_arrmul32_fa9_23_y4, h_u_arrmul32_fa10_23_y2, h_u_arrmul32_fa10_23_y4);
  and_gate and_gate_h_u_arrmul32_and11_23_y0(a_11, b_23, h_u_arrmul32_and11_23_y0);
  fa fa_h_u_arrmul32_fa11_23_y2(h_u_arrmul32_and11_23_y0, h_u_arrmul32_fa12_22_y2, h_u_arrmul32_fa10_23_y4, h_u_arrmul32_fa11_23_y2, h_u_arrmul32_fa11_23_y4);
  and_gate and_gate_h_u_arrmul32_and12_23_y0(a_12, b_23, h_u_arrmul32_and12_23_y0);
  fa fa_h_u_arrmul32_fa12_23_y2(h_u_arrmul32_and12_23_y0, h_u_arrmul32_fa13_22_y2, h_u_arrmul32_fa11_23_y4, h_u_arrmul32_fa12_23_y2, h_u_arrmul32_fa12_23_y4);
  and_gate and_gate_h_u_arrmul32_and13_23_y0(a_13, b_23, h_u_arrmul32_and13_23_y0);
  fa fa_h_u_arrmul32_fa13_23_y2(h_u_arrmul32_and13_23_y0, h_u_arrmul32_fa14_22_y2, h_u_arrmul32_fa12_23_y4, h_u_arrmul32_fa13_23_y2, h_u_arrmul32_fa13_23_y4);
  and_gate and_gate_h_u_arrmul32_and14_23_y0(a_14, b_23, h_u_arrmul32_and14_23_y0);
  fa fa_h_u_arrmul32_fa14_23_y2(h_u_arrmul32_and14_23_y0, h_u_arrmul32_fa15_22_y2, h_u_arrmul32_fa13_23_y4, h_u_arrmul32_fa14_23_y2, h_u_arrmul32_fa14_23_y4);
  and_gate and_gate_h_u_arrmul32_and15_23_y0(a_15, b_23, h_u_arrmul32_and15_23_y0);
  fa fa_h_u_arrmul32_fa15_23_y2(h_u_arrmul32_and15_23_y0, h_u_arrmul32_fa16_22_y2, h_u_arrmul32_fa14_23_y4, h_u_arrmul32_fa15_23_y2, h_u_arrmul32_fa15_23_y4);
  and_gate and_gate_h_u_arrmul32_and16_23_y0(a_16, b_23, h_u_arrmul32_and16_23_y0);
  fa fa_h_u_arrmul32_fa16_23_y2(h_u_arrmul32_and16_23_y0, h_u_arrmul32_fa17_22_y2, h_u_arrmul32_fa15_23_y4, h_u_arrmul32_fa16_23_y2, h_u_arrmul32_fa16_23_y4);
  and_gate and_gate_h_u_arrmul32_and17_23_y0(a_17, b_23, h_u_arrmul32_and17_23_y0);
  fa fa_h_u_arrmul32_fa17_23_y2(h_u_arrmul32_and17_23_y0, h_u_arrmul32_fa18_22_y2, h_u_arrmul32_fa16_23_y4, h_u_arrmul32_fa17_23_y2, h_u_arrmul32_fa17_23_y4);
  and_gate and_gate_h_u_arrmul32_and18_23_y0(a_18, b_23, h_u_arrmul32_and18_23_y0);
  fa fa_h_u_arrmul32_fa18_23_y2(h_u_arrmul32_and18_23_y0, h_u_arrmul32_fa19_22_y2, h_u_arrmul32_fa17_23_y4, h_u_arrmul32_fa18_23_y2, h_u_arrmul32_fa18_23_y4);
  and_gate and_gate_h_u_arrmul32_and19_23_y0(a_19, b_23, h_u_arrmul32_and19_23_y0);
  fa fa_h_u_arrmul32_fa19_23_y2(h_u_arrmul32_and19_23_y0, h_u_arrmul32_fa20_22_y2, h_u_arrmul32_fa18_23_y4, h_u_arrmul32_fa19_23_y2, h_u_arrmul32_fa19_23_y4);
  and_gate and_gate_h_u_arrmul32_and20_23_y0(a_20, b_23, h_u_arrmul32_and20_23_y0);
  fa fa_h_u_arrmul32_fa20_23_y2(h_u_arrmul32_and20_23_y0, h_u_arrmul32_fa21_22_y2, h_u_arrmul32_fa19_23_y4, h_u_arrmul32_fa20_23_y2, h_u_arrmul32_fa20_23_y4);
  and_gate and_gate_h_u_arrmul32_and21_23_y0(a_21, b_23, h_u_arrmul32_and21_23_y0);
  fa fa_h_u_arrmul32_fa21_23_y2(h_u_arrmul32_and21_23_y0, h_u_arrmul32_fa22_22_y2, h_u_arrmul32_fa20_23_y4, h_u_arrmul32_fa21_23_y2, h_u_arrmul32_fa21_23_y4);
  and_gate and_gate_h_u_arrmul32_and22_23_y0(a_22, b_23, h_u_arrmul32_and22_23_y0);
  fa fa_h_u_arrmul32_fa22_23_y2(h_u_arrmul32_and22_23_y0, h_u_arrmul32_fa23_22_y2, h_u_arrmul32_fa21_23_y4, h_u_arrmul32_fa22_23_y2, h_u_arrmul32_fa22_23_y4);
  and_gate and_gate_h_u_arrmul32_and23_23_y0(a_23, b_23, h_u_arrmul32_and23_23_y0);
  fa fa_h_u_arrmul32_fa23_23_y2(h_u_arrmul32_and23_23_y0, h_u_arrmul32_fa24_22_y2, h_u_arrmul32_fa22_23_y4, h_u_arrmul32_fa23_23_y2, h_u_arrmul32_fa23_23_y4);
  and_gate and_gate_h_u_arrmul32_and24_23_y0(a_24, b_23, h_u_arrmul32_and24_23_y0);
  fa fa_h_u_arrmul32_fa24_23_y2(h_u_arrmul32_and24_23_y0, h_u_arrmul32_fa25_22_y2, h_u_arrmul32_fa23_23_y4, h_u_arrmul32_fa24_23_y2, h_u_arrmul32_fa24_23_y4);
  and_gate and_gate_h_u_arrmul32_and25_23_y0(a_25, b_23, h_u_arrmul32_and25_23_y0);
  fa fa_h_u_arrmul32_fa25_23_y2(h_u_arrmul32_and25_23_y0, h_u_arrmul32_fa26_22_y2, h_u_arrmul32_fa24_23_y4, h_u_arrmul32_fa25_23_y2, h_u_arrmul32_fa25_23_y4);
  and_gate and_gate_h_u_arrmul32_and26_23_y0(a_26, b_23, h_u_arrmul32_and26_23_y0);
  fa fa_h_u_arrmul32_fa26_23_y2(h_u_arrmul32_and26_23_y0, h_u_arrmul32_fa27_22_y2, h_u_arrmul32_fa25_23_y4, h_u_arrmul32_fa26_23_y2, h_u_arrmul32_fa26_23_y4);
  and_gate and_gate_h_u_arrmul32_and27_23_y0(a_27, b_23, h_u_arrmul32_and27_23_y0);
  fa fa_h_u_arrmul32_fa27_23_y2(h_u_arrmul32_and27_23_y0, h_u_arrmul32_fa28_22_y2, h_u_arrmul32_fa26_23_y4, h_u_arrmul32_fa27_23_y2, h_u_arrmul32_fa27_23_y4);
  and_gate and_gate_h_u_arrmul32_and28_23_y0(a_28, b_23, h_u_arrmul32_and28_23_y0);
  fa fa_h_u_arrmul32_fa28_23_y2(h_u_arrmul32_and28_23_y0, h_u_arrmul32_fa29_22_y2, h_u_arrmul32_fa27_23_y4, h_u_arrmul32_fa28_23_y2, h_u_arrmul32_fa28_23_y4);
  and_gate and_gate_h_u_arrmul32_and29_23_y0(a_29, b_23, h_u_arrmul32_and29_23_y0);
  fa fa_h_u_arrmul32_fa29_23_y2(h_u_arrmul32_and29_23_y0, h_u_arrmul32_fa30_22_y2, h_u_arrmul32_fa28_23_y4, h_u_arrmul32_fa29_23_y2, h_u_arrmul32_fa29_23_y4);
  and_gate and_gate_h_u_arrmul32_and30_23_y0(a_30, b_23, h_u_arrmul32_and30_23_y0);
  fa fa_h_u_arrmul32_fa30_23_y2(h_u_arrmul32_and30_23_y0, h_u_arrmul32_fa31_22_y2, h_u_arrmul32_fa29_23_y4, h_u_arrmul32_fa30_23_y2, h_u_arrmul32_fa30_23_y4);
  and_gate and_gate_h_u_arrmul32_and31_23_y0(a_31, b_23, h_u_arrmul32_and31_23_y0);
  fa fa_h_u_arrmul32_fa31_23_y2(h_u_arrmul32_and31_23_y0, h_u_arrmul32_fa31_22_y4, h_u_arrmul32_fa30_23_y4, h_u_arrmul32_fa31_23_y2, h_u_arrmul32_fa31_23_y4);
  and_gate and_gate_h_u_arrmul32_and0_24_y0(a_0, b_24, h_u_arrmul32_and0_24_y0);
  ha ha_h_u_arrmul32_ha0_24_y0(h_u_arrmul32_and0_24_y0, h_u_arrmul32_fa1_23_y2, h_u_arrmul32_ha0_24_y0, h_u_arrmul32_ha0_24_y1);
  and_gate and_gate_h_u_arrmul32_and1_24_y0(a_1, b_24, h_u_arrmul32_and1_24_y0);
  fa fa_h_u_arrmul32_fa1_24_y2(h_u_arrmul32_and1_24_y0, h_u_arrmul32_fa2_23_y2, h_u_arrmul32_ha0_24_y1, h_u_arrmul32_fa1_24_y2, h_u_arrmul32_fa1_24_y4);
  and_gate and_gate_h_u_arrmul32_and2_24_y0(a_2, b_24, h_u_arrmul32_and2_24_y0);
  fa fa_h_u_arrmul32_fa2_24_y2(h_u_arrmul32_and2_24_y0, h_u_arrmul32_fa3_23_y2, h_u_arrmul32_fa1_24_y4, h_u_arrmul32_fa2_24_y2, h_u_arrmul32_fa2_24_y4);
  and_gate and_gate_h_u_arrmul32_and3_24_y0(a_3, b_24, h_u_arrmul32_and3_24_y0);
  fa fa_h_u_arrmul32_fa3_24_y2(h_u_arrmul32_and3_24_y0, h_u_arrmul32_fa4_23_y2, h_u_arrmul32_fa2_24_y4, h_u_arrmul32_fa3_24_y2, h_u_arrmul32_fa3_24_y4);
  and_gate and_gate_h_u_arrmul32_and4_24_y0(a_4, b_24, h_u_arrmul32_and4_24_y0);
  fa fa_h_u_arrmul32_fa4_24_y2(h_u_arrmul32_and4_24_y0, h_u_arrmul32_fa5_23_y2, h_u_arrmul32_fa3_24_y4, h_u_arrmul32_fa4_24_y2, h_u_arrmul32_fa4_24_y4);
  and_gate and_gate_h_u_arrmul32_and5_24_y0(a_5, b_24, h_u_arrmul32_and5_24_y0);
  fa fa_h_u_arrmul32_fa5_24_y2(h_u_arrmul32_and5_24_y0, h_u_arrmul32_fa6_23_y2, h_u_arrmul32_fa4_24_y4, h_u_arrmul32_fa5_24_y2, h_u_arrmul32_fa5_24_y4);
  and_gate and_gate_h_u_arrmul32_and6_24_y0(a_6, b_24, h_u_arrmul32_and6_24_y0);
  fa fa_h_u_arrmul32_fa6_24_y2(h_u_arrmul32_and6_24_y0, h_u_arrmul32_fa7_23_y2, h_u_arrmul32_fa5_24_y4, h_u_arrmul32_fa6_24_y2, h_u_arrmul32_fa6_24_y4);
  and_gate and_gate_h_u_arrmul32_and7_24_y0(a_7, b_24, h_u_arrmul32_and7_24_y0);
  fa fa_h_u_arrmul32_fa7_24_y2(h_u_arrmul32_and7_24_y0, h_u_arrmul32_fa8_23_y2, h_u_arrmul32_fa6_24_y4, h_u_arrmul32_fa7_24_y2, h_u_arrmul32_fa7_24_y4);
  and_gate and_gate_h_u_arrmul32_and8_24_y0(a_8, b_24, h_u_arrmul32_and8_24_y0);
  fa fa_h_u_arrmul32_fa8_24_y2(h_u_arrmul32_and8_24_y0, h_u_arrmul32_fa9_23_y2, h_u_arrmul32_fa7_24_y4, h_u_arrmul32_fa8_24_y2, h_u_arrmul32_fa8_24_y4);
  and_gate and_gate_h_u_arrmul32_and9_24_y0(a_9, b_24, h_u_arrmul32_and9_24_y0);
  fa fa_h_u_arrmul32_fa9_24_y2(h_u_arrmul32_and9_24_y0, h_u_arrmul32_fa10_23_y2, h_u_arrmul32_fa8_24_y4, h_u_arrmul32_fa9_24_y2, h_u_arrmul32_fa9_24_y4);
  and_gate and_gate_h_u_arrmul32_and10_24_y0(a_10, b_24, h_u_arrmul32_and10_24_y0);
  fa fa_h_u_arrmul32_fa10_24_y2(h_u_arrmul32_and10_24_y0, h_u_arrmul32_fa11_23_y2, h_u_arrmul32_fa9_24_y4, h_u_arrmul32_fa10_24_y2, h_u_arrmul32_fa10_24_y4);
  and_gate and_gate_h_u_arrmul32_and11_24_y0(a_11, b_24, h_u_arrmul32_and11_24_y0);
  fa fa_h_u_arrmul32_fa11_24_y2(h_u_arrmul32_and11_24_y0, h_u_arrmul32_fa12_23_y2, h_u_arrmul32_fa10_24_y4, h_u_arrmul32_fa11_24_y2, h_u_arrmul32_fa11_24_y4);
  and_gate and_gate_h_u_arrmul32_and12_24_y0(a_12, b_24, h_u_arrmul32_and12_24_y0);
  fa fa_h_u_arrmul32_fa12_24_y2(h_u_arrmul32_and12_24_y0, h_u_arrmul32_fa13_23_y2, h_u_arrmul32_fa11_24_y4, h_u_arrmul32_fa12_24_y2, h_u_arrmul32_fa12_24_y4);
  and_gate and_gate_h_u_arrmul32_and13_24_y0(a_13, b_24, h_u_arrmul32_and13_24_y0);
  fa fa_h_u_arrmul32_fa13_24_y2(h_u_arrmul32_and13_24_y0, h_u_arrmul32_fa14_23_y2, h_u_arrmul32_fa12_24_y4, h_u_arrmul32_fa13_24_y2, h_u_arrmul32_fa13_24_y4);
  and_gate and_gate_h_u_arrmul32_and14_24_y0(a_14, b_24, h_u_arrmul32_and14_24_y0);
  fa fa_h_u_arrmul32_fa14_24_y2(h_u_arrmul32_and14_24_y0, h_u_arrmul32_fa15_23_y2, h_u_arrmul32_fa13_24_y4, h_u_arrmul32_fa14_24_y2, h_u_arrmul32_fa14_24_y4);
  and_gate and_gate_h_u_arrmul32_and15_24_y0(a_15, b_24, h_u_arrmul32_and15_24_y0);
  fa fa_h_u_arrmul32_fa15_24_y2(h_u_arrmul32_and15_24_y0, h_u_arrmul32_fa16_23_y2, h_u_arrmul32_fa14_24_y4, h_u_arrmul32_fa15_24_y2, h_u_arrmul32_fa15_24_y4);
  and_gate and_gate_h_u_arrmul32_and16_24_y0(a_16, b_24, h_u_arrmul32_and16_24_y0);
  fa fa_h_u_arrmul32_fa16_24_y2(h_u_arrmul32_and16_24_y0, h_u_arrmul32_fa17_23_y2, h_u_arrmul32_fa15_24_y4, h_u_arrmul32_fa16_24_y2, h_u_arrmul32_fa16_24_y4);
  and_gate and_gate_h_u_arrmul32_and17_24_y0(a_17, b_24, h_u_arrmul32_and17_24_y0);
  fa fa_h_u_arrmul32_fa17_24_y2(h_u_arrmul32_and17_24_y0, h_u_arrmul32_fa18_23_y2, h_u_arrmul32_fa16_24_y4, h_u_arrmul32_fa17_24_y2, h_u_arrmul32_fa17_24_y4);
  and_gate and_gate_h_u_arrmul32_and18_24_y0(a_18, b_24, h_u_arrmul32_and18_24_y0);
  fa fa_h_u_arrmul32_fa18_24_y2(h_u_arrmul32_and18_24_y0, h_u_arrmul32_fa19_23_y2, h_u_arrmul32_fa17_24_y4, h_u_arrmul32_fa18_24_y2, h_u_arrmul32_fa18_24_y4);
  and_gate and_gate_h_u_arrmul32_and19_24_y0(a_19, b_24, h_u_arrmul32_and19_24_y0);
  fa fa_h_u_arrmul32_fa19_24_y2(h_u_arrmul32_and19_24_y0, h_u_arrmul32_fa20_23_y2, h_u_arrmul32_fa18_24_y4, h_u_arrmul32_fa19_24_y2, h_u_arrmul32_fa19_24_y4);
  and_gate and_gate_h_u_arrmul32_and20_24_y0(a_20, b_24, h_u_arrmul32_and20_24_y0);
  fa fa_h_u_arrmul32_fa20_24_y2(h_u_arrmul32_and20_24_y0, h_u_arrmul32_fa21_23_y2, h_u_arrmul32_fa19_24_y4, h_u_arrmul32_fa20_24_y2, h_u_arrmul32_fa20_24_y4);
  and_gate and_gate_h_u_arrmul32_and21_24_y0(a_21, b_24, h_u_arrmul32_and21_24_y0);
  fa fa_h_u_arrmul32_fa21_24_y2(h_u_arrmul32_and21_24_y0, h_u_arrmul32_fa22_23_y2, h_u_arrmul32_fa20_24_y4, h_u_arrmul32_fa21_24_y2, h_u_arrmul32_fa21_24_y4);
  and_gate and_gate_h_u_arrmul32_and22_24_y0(a_22, b_24, h_u_arrmul32_and22_24_y0);
  fa fa_h_u_arrmul32_fa22_24_y2(h_u_arrmul32_and22_24_y0, h_u_arrmul32_fa23_23_y2, h_u_arrmul32_fa21_24_y4, h_u_arrmul32_fa22_24_y2, h_u_arrmul32_fa22_24_y4);
  and_gate and_gate_h_u_arrmul32_and23_24_y0(a_23, b_24, h_u_arrmul32_and23_24_y0);
  fa fa_h_u_arrmul32_fa23_24_y2(h_u_arrmul32_and23_24_y0, h_u_arrmul32_fa24_23_y2, h_u_arrmul32_fa22_24_y4, h_u_arrmul32_fa23_24_y2, h_u_arrmul32_fa23_24_y4);
  and_gate and_gate_h_u_arrmul32_and24_24_y0(a_24, b_24, h_u_arrmul32_and24_24_y0);
  fa fa_h_u_arrmul32_fa24_24_y2(h_u_arrmul32_and24_24_y0, h_u_arrmul32_fa25_23_y2, h_u_arrmul32_fa23_24_y4, h_u_arrmul32_fa24_24_y2, h_u_arrmul32_fa24_24_y4);
  and_gate and_gate_h_u_arrmul32_and25_24_y0(a_25, b_24, h_u_arrmul32_and25_24_y0);
  fa fa_h_u_arrmul32_fa25_24_y2(h_u_arrmul32_and25_24_y0, h_u_arrmul32_fa26_23_y2, h_u_arrmul32_fa24_24_y4, h_u_arrmul32_fa25_24_y2, h_u_arrmul32_fa25_24_y4);
  and_gate and_gate_h_u_arrmul32_and26_24_y0(a_26, b_24, h_u_arrmul32_and26_24_y0);
  fa fa_h_u_arrmul32_fa26_24_y2(h_u_arrmul32_and26_24_y0, h_u_arrmul32_fa27_23_y2, h_u_arrmul32_fa25_24_y4, h_u_arrmul32_fa26_24_y2, h_u_arrmul32_fa26_24_y4);
  and_gate and_gate_h_u_arrmul32_and27_24_y0(a_27, b_24, h_u_arrmul32_and27_24_y0);
  fa fa_h_u_arrmul32_fa27_24_y2(h_u_arrmul32_and27_24_y0, h_u_arrmul32_fa28_23_y2, h_u_arrmul32_fa26_24_y4, h_u_arrmul32_fa27_24_y2, h_u_arrmul32_fa27_24_y4);
  and_gate and_gate_h_u_arrmul32_and28_24_y0(a_28, b_24, h_u_arrmul32_and28_24_y0);
  fa fa_h_u_arrmul32_fa28_24_y2(h_u_arrmul32_and28_24_y0, h_u_arrmul32_fa29_23_y2, h_u_arrmul32_fa27_24_y4, h_u_arrmul32_fa28_24_y2, h_u_arrmul32_fa28_24_y4);
  and_gate and_gate_h_u_arrmul32_and29_24_y0(a_29, b_24, h_u_arrmul32_and29_24_y0);
  fa fa_h_u_arrmul32_fa29_24_y2(h_u_arrmul32_and29_24_y0, h_u_arrmul32_fa30_23_y2, h_u_arrmul32_fa28_24_y4, h_u_arrmul32_fa29_24_y2, h_u_arrmul32_fa29_24_y4);
  and_gate and_gate_h_u_arrmul32_and30_24_y0(a_30, b_24, h_u_arrmul32_and30_24_y0);
  fa fa_h_u_arrmul32_fa30_24_y2(h_u_arrmul32_and30_24_y0, h_u_arrmul32_fa31_23_y2, h_u_arrmul32_fa29_24_y4, h_u_arrmul32_fa30_24_y2, h_u_arrmul32_fa30_24_y4);
  and_gate and_gate_h_u_arrmul32_and31_24_y0(a_31, b_24, h_u_arrmul32_and31_24_y0);
  fa fa_h_u_arrmul32_fa31_24_y2(h_u_arrmul32_and31_24_y0, h_u_arrmul32_fa31_23_y4, h_u_arrmul32_fa30_24_y4, h_u_arrmul32_fa31_24_y2, h_u_arrmul32_fa31_24_y4);
  and_gate and_gate_h_u_arrmul32_and0_25_y0(a_0, b_25, h_u_arrmul32_and0_25_y0);
  ha ha_h_u_arrmul32_ha0_25_y0(h_u_arrmul32_and0_25_y0, h_u_arrmul32_fa1_24_y2, h_u_arrmul32_ha0_25_y0, h_u_arrmul32_ha0_25_y1);
  and_gate and_gate_h_u_arrmul32_and1_25_y0(a_1, b_25, h_u_arrmul32_and1_25_y0);
  fa fa_h_u_arrmul32_fa1_25_y2(h_u_arrmul32_and1_25_y0, h_u_arrmul32_fa2_24_y2, h_u_arrmul32_ha0_25_y1, h_u_arrmul32_fa1_25_y2, h_u_arrmul32_fa1_25_y4);
  and_gate and_gate_h_u_arrmul32_and2_25_y0(a_2, b_25, h_u_arrmul32_and2_25_y0);
  fa fa_h_u_arrmul32_fa2_25_y2(h_u_arrmul32_and2_25_y0, h_u_arrmul32_fa3_24_y2, h_u_arrmul32_fa1_25_y4, h_u_arrmul32_fa2_25_y2, h_u_arrmul32_fa2_25_y4);
  and_gate and_gate_h_u_arrmul32_and3_25_y0(a_3, b_25, h_u_arrmul32_and3_25_y0);
  fa fa_h_u_arrmul32_fa3_25_y2(h_u_arrmul32_and3_25_y0, h_u_arrmul32_fa4_24_y2, h_u_arrmul32_fa2_25_y4, h_u_arrmul32_fa3_25_y2, h_u_arrmul32_fa3_25_y4);
  and_gate and_gate_h_u_arrmul32_and4_25_y0(a_4, b_25, h_u_arrmul32_and4_25_y0);
  fa fa_h_u_arrmul32_fa4_25_y2(h_u_arrmul32_and4_25_y0, h_u_arrmul32_fa5_24_y2, h_u_arrmul32_fa3_25_y4, h_u_arrmul32_fa4_25_y2, h_u_arrmul32_fa4_25_y4);
  and_gate and_gate_h_u_arrmul32_and5_25_y0(a_5, b_25, h_u_arrmul32_and5_25_y0);
  fa fa_h_u_arrmul32_fa5_25_y2(h_u_arrmul32_and5_25_y0, h_u_arrmul32_fa6_24_y2, h_u_arrmul32_fa4_25_y4, h_u_arrmul32_fa5_25_y2, h_u_arrmul32_fa5_25_y4);
  and_gate and_gate_h_u_arrmul32_and6_25_y0(a_6, b_25, h_u_arrmul32_and6_25_y0);
  fa fa_h_u_arrmul32_fa6_25_y2(h_u_arrmul32_and6_25_y0, h_u_arrmul32_fa7_24_y2, h_u_arrmul32_fa5_25_y4, h_u_arrmul32_fa6_25_y2, h_u_arrmul32_fa6_25_y4);
  and_gate and_gate_h_u_arrmul32_and7_25_y0(a_7, b_25, h_u_arrmul32_and7_25_y0);
  fa fa_h_u_arrmul32_fa7_25_y2(h_u_arrmul32_and7_25_y0, h_u_arrmul32_fa8_24_y2, h_u_arrmul32_fa6_25_y4, h_u_arrmul32_fa7_25_y2, h_u_arrmul32_fa7_25_y4);
  and_gate and_gate_h_u_arrmul32_and8_25_y0(a_8, b_25, h_u_arrmul32_and8_25_y0);
  fa fa_h_u_arrmul32_fa8_25_y2(h_u_arrmul32_and8_25_y0, h_u_arrmul32_fa9_24_y2, h_u_arrmul32_fa7_25_y4, h_u_arrmul32_fa8_25_y2, h_u_arrmul32_fa8_25_y4);
  and_gate and_gate_h_u_arrmul32_and9_25_y0(a_9, b_25, h_u_arrmul32_and9_25_y0);
  fa fa_h_u_arrmul32_fa9_25_y2(h_u_arrmul32_and9_25_y0, h_u_arrmul32_fa10_24_y2, h_u_arrmul32_fa8_25_y4, h_u_arrmul32_fa9_25_y2, h_u_arrmul32_fa9_25_y4);
  and_gate and_gate_h_u_arrmul32_and10_25_y0(a_10, b_25, h_u_arrmul32_and10_25_y0);
  fa fa_h_u_arrmul32_fa10_25_y2(h_u_arrmul32_and10_25_y0, h_u_arrmul32_fa11_24_y2, h_u_arrmul32_fa9_25_y4, h_u_arrmul32_fa10_25_y2, h_u_arrmul32_fa10_25_y4);
  and_gate and_gate_h_u_arrmul32_and11_25_y0(a_11, b_25, h_u_arrmul32_and11_25_y0);
  fa fa_h_u_arrmul32_fa11_25_y2(h_u_arrmul32_and11_25_y0, h_u_arrmul32_fa12_24_y2, h_u_arrmul32_fa10_25_y4, h_u_arrmul32_fa11_25_y2, h_u_arrmul32_fa11_25_y4);
  and_gate and_gate_h_u_arrmul32_and12_25_y0(a_12, b_25, h_u_arrmul32_and12_25_y0);
  fa fa_h_u_arrmul32_fa12_25_y2(h_u_arrmul32_and12_25_y0, h_u_arrmul32_fa13_24_y2, h_u_arrmul32_fa11_25_y4, h_u_arrmul32_fa12_25_y2, h_u_arrmul32_fa12_25_y4);
  and_gate and_gate_h_u_arrmul32_and13_25_y0(a_13, b_25, h_u_arrmul32_and13_25_y0);
  fa fa_h_u_arrmul32_fa13_25_y2(h_u_arrmul32_and13_25_y0, h_u_arrmul32_fa14_24_y2, h_u_arrmul32_fa12_25_y4, h_u_arrmul32_fa13_25_y2, h_u_arrmul32_fa13_25_y4);
  and_gate and_gate_h_u_arrmul32_and14_25_y0(a_14, b_25, h_u_arrmul32_and14_25_y0);
  fa fa_h_u_arrmul32_fa14_25_y2(h_u_arrmul32_and14_25_y0, h_u_arrmul32_fa15_24_y2, h_u_arrmul32_fa13_25_y4, h_u_arrmul32_fa14_25_y2, h_u_arrmul32_fa14_25_y4);
  and_gate and_gate_h_u_arrmul32_and15_25_y0(a_15, b_25, h_u_arrmul32_and15_25_y0);
  fa fa_h_u_arrmul32_fa15_25_y2(h_u_arrmul32_and15_25_y0, h_u_arrmul32_fa16_24_y2, h_u_arrmul32_fa14_25_y4, h_u_arrmul32_fa15_25_y2, h_u_arrmul32_fa15_25_y4);
  and_gate and_gate_h_u_arrmul32_and16_25_y0(a_16, b_25, h_u_arrmul32_and16_25_y0);
  fa fa_h_u_arrmul32_fa16_25_y2(h_u_arrmul32_and16_25_y0, h_u_arrmul32_fa17_24_y2, h_u_arrmul32_fa15_25_y4, h_u_arrmul32_fa16_25_y2, h_u_arrmul32_fa16_25_y4);
  and_gate and_gate_h_u_arrmul32_and17_25_y0(a_17, b_25, h_u_arrmul32_and17_25_y0);
  fa fa_h_u_arrmul32_fa17_25_y2(h_u_arrmul32_and17_25_y0, h_u_arrmul32_fa18_24_y2, h_u_arrmul32_fa16_25_y4, h_u_arrmul32_fa17_25_y2, h_u_arrmul32_fa17_25_y4);
  and_gate and_gate_h_u_arrmul32_and18_25_y0(a_18, b_25, h_u_arrmul32_and18_25_y0);
  fa fa_h_u_arrmul32_fa18_25_y2(h_u_arrmul32_and18_25_y0, h_u_arrmul32_fa19_24_y2, h_u_arrmul32_fa17_25_y4, h_u_arrmul32_fa18_25_y2, h_u_arrmul32_fa18_25_y4);
  and_gate and_gate_h_u_arrmul32_and19_25_y0(a_19, b_25, h_u_arrmul32_and19_25_y0);
  fa fa_h_u_arrmul32_fa19_25_y2(h_u_arrmul32_and19_25_y0, h_u_arrmul32_fa20_24_y2, h_u_arrmul32_fa18_25_y4, h_u_arrmul32_fa19_25_y2, h_u_arrmul32_fa19_25_y4);
  and_gate and_gate_h_u_arrmul32_and20_25_y0(a_20, b_25, h_u_arrmul32_and20_25_y0);
  fa fa_h_u_arrmul32_fa20_25_y2(h_u_arrmul32_and20_25_y0, h_u_arrmul32_fa21_24_y2, h_u_arrmul32_fa19_25_y4, h_u_arrmul32_fa20_25_y2, h_u_arrmul32_fa20_25_y4);
  and_gate and_gate_h_u_arrmul32_and21_25_y0(a_21, b_25, h_u_arrmul32_and21_25_y0);
  fa fa_h_u_arrmul32_fa21_25_y2(h_u_arrmul32_and21_25_y0, h_u_arrmul32_fa22_24_y2, h_u_arrmul32_fa20_25_y4, h_u_arrmul32_fa21_25_y2, h_u_arrmul32_fa21_25_y4);
  and_gate and_gate_h_u_arrmul32_and22_25_y0(a_22, b_25, h_u_arrmul32_and22_25_y0);
  fa fa_h_u_arrmul32_fa22_25_y2(h_u_arrmul32_and22_25_y0, h_u_arrmul32_fa23_24_y2, h_u_arrmul32_fa21_25_y4, h_u_arrmul32_fa22_25_y2, h_u_arrmul32_fa22_25_y4);
  and_gate and_gate_h_u_arrmul32_and23_25_y0(a_23, b_25, h_u_arrmul32_and23_25_y0);
  fa fa_h_u_arrmul32_fa23_25_y2(h_u_arrmul32_and23_25_y0, h_u_arrmul32_fa24_24_y2, h_u_arrmul32_fa22_25_y4, h_u_arrmul32_fa23_25_y2, h_u_arrmul32_fa23_25_y4);
  and_gate and_gate_h_u_arrmul32_and24_25_y0(a_24, b_25, h_u_arrmul32_and24_25_y0);
  fa fa_h_u_arrmul32_fa24_25_y2(h_u_arrmul32_and24_25_y0, h_u_arrmul32_fa25_24_y2, h_u_arrmul32_fa23_25_y4, h_u_arrmul32_fa24_25_y2, h_u_arrmul32_fa24_25_y4);
  and_gate and_gate_h_u_arrmul32_and25_25_y0(a_25, b_25, h_u_arrmul32_and25_25_y0);
  fa fa_h_u_arrmul32_fa25_25_y2(h_u_arrmul32_and25_25_y0, h_u_arrmul32_fa26_24_y2, h_u_arrmul32_fa24_25_y4, h_u_arrmul32_fa25_25_y2, h_u_arrmul32_fa25_25_y4);
  and_gate and_gate_h_u_arrmul32_and26_25_y0(a_26, b_25, h_u_arrmul32_and26_25_y0);
  fa fa_h_u_arrmul32_fa26_25_y2(h_u_arrmul32_and26_25_y0, h_u_arrmul32_fa27_24_y2, h_u_arrmul32_fa25_25_y4, h_u_arrmul32_fa26_25_y2, h_u_arrmul32_fa26_25_y4);
  and_gate and_gate_h_u_arrmul32_and27_25_y0(a_27, b_25, h_u_arrmul32_and27_25_y0);
  fa fa_h_u_arrmul32_fa27_25_y2(h_u_arrmul32_and27_25_y0, h_u_arrmul32_fa28_24_y2, h_u_arrmul32_fa26_25_y4, h_u_arrmul32_fa27_25_y2, h_u_arrmul32_fa27_25_y4);
  and_gate and_gate_h_u_arrmul32_and28_25_y0(a_28, b_25, h_u_arrmul32_and28_25_y0);
  fa fa_h_u_arrmul32_fa28_25_y2(h_u_arrmul32_and28_25_y0, h_u_arrmul32_fa29_24_y2, h_u_arrmul32_fa27_25_y4, h_u_arrmul32_fa28_25_y2, h_u_arrmul32_fa28_25_y4);
  and_gate and_gate_h_u_arrmul32_and29_25_y0(a_29, b_25, h_u_arrmul32_and29_25_y0);
  fa fa_h_u_arrmul32_fa29_25_y2(h_u_arrmul32_and29_25_y0, h_u_arrmul32_fa30_24_y2, h_u_arrmul32_fa28_25_y4, h_u_arrmul32_fa29_25_y2, h_u_arrmul32_fa29_25_y4);
  and_gate and_gate_h_u_arrmul32_and30_25_y0(a_30, b_25, h_u_arrmul32_and30_25_y0);
  fa fa_h_u_arrmul32_fa30_25_y2(h_u_arrmul32_and30_25_y0, h_u_arrmul32_fa31_24_y2, h_u_arrmul32_fa29_25_y4, h_u_arrmul32_fa30_25_y2, h_u_arrmul32_fa30_25_y4);
  and_gate and_gate_h_u_arrmul32_and31_25_y0(a_31, b_25, h_u_arrmul32_and31_25_y0);
  fa fa_h_u_arrmul32_fa31_25_y2(h_u_arrmul32_and31_25_y0, h_u_arrmul32_fa31_24_y4, h_u_arrmul32_fa30_25_y4, h_u_arrmul32_fa31_25_y2, h_u_arrmul32_fa31_25_y4);
  and_gate and_gate_h_u_arrmul32_and0_26_y0(a_0, b_26, h_u_arrmul32_and0_26_y0);
  ha ha_h_u_arrmul32_ha0_26_y0(h_u_arrmul32_and0_26_y0, h_u_arrmul32_fa1_25_y2, h_u_arrmul32_ha0_26_y0, h_u_arrmul32_ha0_26_y1);
  and_gate and_gate_h_u_arrmul32_and1_26_y0(a_1, b_26, h_u_arrmul32_and1_26_y0);
  fa fa_h_u_arrmul32_fa1_26_y2(h_u_arrmul32_and1_26_y0, h_u_arrmul32_fa2_25_y2, h_u_arrmul32_ha0_26_y1, h_u_arrmul32_fa1_26_y2, h_u_arrmul32_fa1_26_y4);
  and_gate and_gate_h_u_arrmul32_and2_26_y0(a_2, b_26, h_u_arrmul32_and2_26_y0);
  fa fa_h_u_arrmul32_fa2_26_y2(h_u_arrmul32_and2_26_y0, h_u_arrmul32_fa3_25_y2, h_u_arrmul32_fa1_26_y4, h_u_arrmul32_fa2_26_y2, h_u_arrmul32_fa2_26_y4);
  and_gate and_gate_h_u_arrmul32_and3_26_y0(a_3, b_26, h_u_arrmul32_and3_26_y0);
  fa fa_h_u_arrmul32_fa3_26_y2(h_u_arrmul32_and3_26_y0, h_u_arrmul32_fa4_25_y2, h_u_arrmul32_fa2_26_y4, h_u_arrmul32_fa3_26_y2, h_u_arrmul32_fa3_26_y4);
  and_gate and_gate_h_u_arrmul32_and4_26_y0(a_4, b_26, h_u_arrmul32_and4_26_y0);
  fa fa_h_u_arrmul32_fa4_26_y2(h_u_arrmul32_and4_26_y0, h_u_arrmul32_fa5_25_y2, h_u_arrmul32_fa3_26_y4, h_u_arrmul32_fa4_26_y2, h_u_arrmul32_fa4_26_y4);
  and_gate and_gate_h_u_arrmul32_and5_26_y0(a_5, b_26, h_u_arrmul32_and5_26_y0);
  fa fa_h_u_arrmul32_fa5_26_y2(h_u_arrmul32_and5_26_y0, h_u_arrmul32_fa6_25_y2, h_u_arrmul32_fa4_26_y4, h_u_arrmul32_fa5_26_y2, h_u_arrmul32_fa5_26_y4);
  and_gate and_gate_h_u_arrmul32_and6_26_y0(a_6, b_26, h_u_arrmul32_and6_26_y0);
  fa fa_h_u_arrmul32_fa6_26_y2(h_u_arrmul32_and6_26_y0, h_u_arrmul32_fa7_25_y2, h_u_arrmul32_fa5_26_y4, h_u_arrmul32_fa6_26_y2, h_u_arrmul32_fa6_26_y4);
  and_gate and_gate_h_u_arrmul32_and7_26_y0(a_7, b_26, h_u_arrmul32_and7_26_y0);
  fa fa_h_u_arrmul32_fa7_26_y2(h_u_arrmul32_and7_26_y0, h_u_arrmul32_fa8_25_y2, h_u_arrmul32_fa6_26_y4, h_u_arrmul32_fa7_26_y2, h_u_arrmul32_fa7_26_y4);
  and_gate and_gate_h_u_arrmul32_and8_26_y0(a_8, b_26, h_u_arrmul32_and8_26_y0);
  fa fa_h_u_arrmul32_fa8_26_y2(h_u_arrmul32_and8_26_y0, h_u_arrmul32_fa9_25_y2, h_u_arrmul32_fa7_26_y4, h_u_arrmul32_fa8_26_y2, h_u_arrmul32_fa8_26_y4);
  and_gate and_gate_h_u_arrmul32_and9_26_y0(a_9, b_26, h_u_arrmul32_and9_26_y0);
  fa fa_h_u_arrmul32_fa9_26_y2(h_u_arrmul32_and9_26_y0, h_u_arrmul32_fa10_25_y2, h_u_arrmul32_fa8_26_y4, h_u_arrmul32_fa9_26_y2, h_u_arrmul32_fa9_26_y4);
  and_gate and_gate_h_u_arrmul32_and10_26_y0(a_10, b_26, h_u_arrmul32_and10_26_y0);
  fa fa_h_u_arrmul32_fa10_26_y2(h_u_arrmul32_and10_26_y0, h_u_arrmul32_fa11_25_y2, h_u_arrmul32_fa9_26_y4, h_u_arrmul32_fa10_26_y2, h_u_arrmul32_fa10_26_y4);
  and_gate and_gate_h_u_arrmul32_and11_26_y0(a_11, b_26, h_u_arrmul32_and11_26_y0);
  fa fa_h_u_arrmul32_fa11_26_y2(h_u_arrmul32_and11_26_y0, h_u_arrmul32_fa12_25_y2, h_u_arrmul32_fa10_26_y4, h_u_arrmul32_fa11_26_y2, h_u_arrmul32_fa11_26_y4);
  and_gate and_gate_h_u_arrmul32_and12_26_y0(a_12, b_26, h_u_arrmul32_and12_26_y0);
  fa fa_h_u_arrmul32_fa12_26_y2(h_u_arrmul32_and12_26_y0, h_u_arrmul32_fa13_25_y2, h_u_arrmul32_fa11_26_y4, h_u_arrmul32_fa12_26_y2, h_u_arrmul32_fa12_26_y4);
  and_gate and_gate_h_u_arrmul32_and13_26_y0(a_13, b_26, h_u_arrmul32_and13_26_y0);
  fa fa_h_u_arrmul32_fa13_26_y2(h_u_arrmul32_and13_26_y0, h_u_arrmul32_fa14_25_y2, h_u_arrmul32_fa12_26_y4, h_u_arrmul32_fa13_26_y2, h_u_arrmul32_fa13_26_y4);
  and_gate and_gate_h_u_arrmul32_and14_26_y0(a_14, b_26, h_u_arrmul32_and14_26_y0);
  fa fa_h_u_arrmul32_fa14_26_y2(h_u_arrmul32_and14_26_y0, h_u_arrmul32_fa15_25_y2, h_u_arrmul32_fa13_26_y4, h_u_arrmul32_fa14_26_y2, h_u_arrmul32_fa14_26_y4);
  and_gate and_gate_h_u_arrmul32_and15_26_y0(a_15, b_26, h_u_arrmul32_and15_26_y0);
  fa fa_h_u_arrmul32_fa15_26_y2(h_u_arrmul32_and15_26_y0, h_u_arrmul32_fa16_25_y2, h_u_arrmul32_fa14_26_y4, h_u_arrmul32_fa15_26_y2, h_u_arrmul32_fa15_26_y4);
  and_gate and_gate_h_u_arrmul32_and16_26_y0(a_16, b_26, h_u_arrmul32_and16_26_y0);
  fa fa_h_u_arrmul32_fa16_26_y2(h_u_arrmul32_and16_26_y0, h_u_arrmul32_fa17_25_y2, h_u_arrmul32_fa15_26_y4, h_u_arrmul32_fa16_26_y2, h_u_arrmul32_fa16_26_y4);
  and_gate and_gate_h_u_arrmul32_and17_26_y0(a_17, b_26, h_u_arrmul32_and17_26_y0);
  fa fa_h_u_arrmul32_fa17_26_y2(h_u_arrmul32_and17_26_y0, h_u_arrmul32_fa18_25_y2, h_u_arrmul32_fa16_26_y4, h_u_arrmul32_fa17_26_y2, h_u_arrmul32_fa17_26_y4);
  and_gate and_gate_h_u_arrmul32_and18_26_y0(a_18, b_26, h_u_arrmul32_and18_26_y0);
  fa fa_h_u_arrmul32_fa18_26_y2(h_u_arrmul32_and18_26_y0, h_u_arrmul32_fa19_25_y2, h_u_arrmul32_fa17_26_y4, h_u_arrmul32_fa18_26_y2, h_u_arrmul32_fa18_26_y4);
  and_gate and_gate_h_u_arrmul32_and19_26_y0(a_19, b_26, h_u_arrmul32_and19_26_y0);
  fa fa_h_u_arrmul32_fa19_26_y2(h_u_arrmul32_and19_26_y0, h_u_arrmul32_fa20_25_y2, h_u_arrmul32_fa18_26_y4, h_u_arrmul32_fa19_26_y2, h_u_arrmul32_fa19_26_y4);
  and_gate and_gate_h_u_arrmul32_and20_26_y0(a_20, b_26, h_u_arrmul32_and20_26_y0);
  fa fa_h_u_arrmul32_fa20_26_y2(h_u_arrmul32_and20_26_y0, h_u_arrmul32_fa21_25_y2, h_u_arrmul32_fa19_26_y4, h_u_arrmul32_fa20_26_y2, h_u_arrmul32_fa20_26_y4);
  and_gate and_gate_h_u_arrmul32_and21_26_y0(a_21, b_26, h_u_arrmul32_and21_26_y0);
  fa fa_h_u_arrmul32_fa21_26_y2(h_u_arrmul32_and21_26_y0, h_u_arrmul32_fa22_25_y2, h_u_arrmul32_fa20_26_y4, h_u_arrmul32_fa21_26_y2, h_u_arrmul32_fa21_26_y4);
  and_gate and_gate_h_u_arrmul32_and22_26_y0(a_22, b_26, h_u_arrmul32_and22_26_y0);
  fa fa_h_u_arrmul32_fa22_26_y2(h_u_arrmul32_and22_26_y0, h_u_arrmul32_fa23_25_y2, h_u_arrmul32_fa21_26_y4, h_u_arrmul32_fa22_26_y2, h_u_arrmul32_fa22_26_y4);
  and_gate and_gate_h_u_arrmul32_and23_26_y0(a_23, b_26, h_u_arrmul32_and23_26_y0);
  fa fa_h_u_arrmul32_fa23_26_y2(h_u_arrmul32_and23_26_y0, h_u_arrmul32_fa24_25_y2, h_u_arrmul32_fa22_26_y4, h_u_arrmul32_fa23_26_y2, h_u_arrmul32_fa23_26_y4);
  and_gate and_gate_h_u_arrmul32_and24_26_y0(a_24, b_26, h_u_arrmul32_and24_26_y0);
  fa fa_h_u_arrmul32_fa24_26_y2(h_u_arrmul32_and24_26_y0, h_u_arrmul32_fa25_25_y2, h_u_arrmul32_fa23_26_y4, h_u_arrmul32_fa24_26_y2, h_u_arrmul32_fa24_26_y4);
  and_gate and_gate_h_u_arrmul32_and25_26_y0(a_25, b_26, h_u_arrmul32_and25_26_y0);
  fa fa_h_u_arrmul32_fa25_26_y2(h_u_arrmul32_and25_26_y0, h_u_arrmul32_fa26_25_y2, h_u_arrmul32_fa24_26_y4, h_u_arrmul32_fa25_26_y2, h_u_arrmul32_fa25_26_y4);
  and_gate and_gate_h_u_arrmul32_and26_26_y0(a_26, b_26, h_u_arrmul32_and26_26_y0);
  fa fa_h_u_arrmul32_fa26_26_y2(h_u_arrmul32_and26_26_y0, h_u_arrmul32_fa27_25_y2, h_u_arrmul32_fa25_26_y4, h_u_arrmul32_fa26_26_y2, h_u_arrmul32_fa26_26_y4);
  and_gate and_gate_h_u_arrmul32_and27_26_y0(a_27, b_26, h_u_arrmul32_and27_26_y0);
  fa fa_h_u_arrmul32_fa27_26_y2(h_u_arrmul32_and27_26_y0, h_u_arrmul32_fa28_25_y2, h_u_arrmul32_fa26_26_y4, h_u_arrmul32_fa27_26_y2, h_u_arrmul32_fa27_26_y4);
  and_gate and_gate_h_u_arrmul32_and28_26_y0(a_28, b_26, h_u_arrmul32_and28_26_y0);
  fa fa_h_u_arrmul32_fa28_26_y2(h_u_arrmul32_and28_26_y0, h_u_arrmul32_fa29_25_y2, h_u_arrmul32_fa27_26_y4, h_u_arrmul32_fa28_26_y2, h_u_arrmul32_fa28_26_y4);
  and_gate and_gate_h_u_arrmul32_and29_26_y0(a_29, b_26, h_u_arrmul32_and29_26_y0);
  fa fa_h_u_arrmul32_fa29_26_y2(h_u_arrmul32_and29_26_y0, h_u_arrmul32_fa30_25_y2, h_u_arrmul32_fa28_26_y4, h_u_arrmul32_fa29_26_y2, h_u_arrmul32_fa29_26_y4);
  and_gate and_gate_h_u_arrmul32_and30_26_y0(a_30, b_26, h_u_arrmul32_and30_26_y0);
  fa fa_h_u_arrmul32_fa30_26_y2(h_u_arrmul32_and30_26_y0, h_u_arrmul32_fa31_25_y2, h_u_arrmul32_fa29_26_y4, h_u_arrmul32_fa30_26_y2, h_u_arrmul32_fa30_26_y4);
  and_gate and_gate_h_u_arrmul32_and31_26_y0(a_31, b_26, h_u_arrmul32_and31_26_y0);
  fa fa_h_u_arrmul32_fa31_26_y2(h_u_arrmul32_and31_26_y0, h_u_arrmul32_fa31_25_y4, h_u_arrmul32_fa30_26_y4, h_u_arrmul32_fa31_26_y2, h_u_arrmul32_fa31_26_y4);
  and_gate and_gate_h_u_arrmul32_and0_27_y0(a_0, b_27, h_u_arrmul32_and0_27_y0);
  ha ha_h_u_arrmul32_ha0_27_y0(h_u_arrmul32_and0_27_y0, h_u_arrmul32_fa1_26_y2, h_u_arrmul32_ha0_27_y0, h_u_arrmul32_ha0_27_y1);
  and_gate and_gate_h_u_arrmul32_and1_27_y0(a_1, b_27, h_u_arrmul32_and1_27_y0);
  fa fa_h_u_arrmul32_fa1_27_y2(h_u_arrmul32_and1_27_y0, h_u_arrmul32_fa2_26_y2, h_u_arrmul32_ha0_27_y1, h_u_arrmul32_fa1_27_y2, h_u_arrmul32_fa1_27_y4);
  and_gate and_gate_h_u_arrmul32_and2_27_y0(a_2, b_27, h_u_arrmul32_and2_27_y0);
  fa fa_h_u_arrmul32_fa2_27_y2(h_u_arrmul32_and2_27_y0, h_u_arrmul32_fa3_26_y2, h_u_arrmul32_fa1_27_y4, h_u_arrmul32_fa2_27_y2, h_u_arrmul32_fa2_27_y4);
  and_gate and_gate_h_u_arrmul32_and3_27_y0(a_3, b_27, h_u_arrmul32_and3_27_y0);
  fa fa_h_u_arrmul32_fa3_27_y2(h_u_arrmul32_and3_27_y0, h_u_arrmul32_fa4_26_y2, h_u_arrmul32_fa2_27_y4, h_u_arrmul32_fa3_27_y2, h_u_arrmul32_fa3_27_y4);
  and_gate and_gate_h_u_arrmul32_and4_27_y0(a_4, b_27, h_u_arrmul32_and4_27_y0);
  fa fa_h_u_arrmul32_fa4_27_y2(h_u_arrmul32_and4_27_y0, h_u_arrmul32_fa5_26_y2, h_u_arrmul32_fa3_27_y4, h_u_arrmul32_fa4_27_y2, h_u_arrmul32_fa4_27_y4);
  and_gate and_gate_h_u_arrmul32_and5_27_y0(a_5, b_27, h_u_arrmul32_and5_27_y0);
  fa fa_h_u_arrmul32_fa5_27_y2(h_u_arrmul32_and5_27_y0, h_u_arrmul32_fa6_26_y2, h_u_arrmul32_fa4_27_y4, h_u_arrmul32_fa5_27_y2, h_u_arrmul32_fa5_27_y4);
  and_gate and_gate_h_u_arrmul32_and6_27_y0(a_6, b_27, h_u_arrmul32_and6_27_y0);
  fa fa_h_u_arrmul32_fa6_27_y2(h_u_arrmul32_and6_27_y0, h_u_arrmul32_fa7_26_y2, h_u_arrmul32_fa5_27_y4, h_u_arrmul32_fa6_27_y2, h_u_arrmul32_fa6_27_y4);
  and_gate and_gate_h_u_arrmul32_and7_27_y0(a_7, b_27, h_u_arrmul32_and7_27_y0);
  fa fa_h_u_arrmul32_fa7_27_y2(h_u_arrmul32_and7_27_y0, h_u_arrmul32_fa8_26_y2, h_u_arrmul32_fa6_27_y4, h_u_arrmul32_fa7_27_y2, h_u_arrmul32_fa7_27_y4);
  and_gate and_gate_h_u_arrmul32_and8_27_y0(a_8, b_27, h_u_arrmul32_and8_27_y0);
  fa fa_h_u_arrmul32_fa8_27_y2(h_u_arrmul32_and8_27_y0, h_u_arrmul32_fa9_26_y2, h_u_arrmul32_fa7_27_y4, h_u_arrmul32_fa8_27_y2, h_u_arrmul32_fa8_27_y4);
  and_gate and_gate_h_u_arrmul32_and9_27_y0(a_9, b_27, h_u_arrmul32_and9_27_y0);
  fa fa_h_u_arrmul32_fa9_27_y2(h_u_arrmul32_and9_27_y0, h_u_arrmul32_fa10_26_y2, h_u_arrmul32_fa8_27_y4, h_u_arrmul32_fa9_27_y2, h_u_arrmul32_fa9_27_y4);
  and_gate and_gate_h_u_arrmul32_and10_27_y0(a_10, b_27, h_u_arrmul32_and10_27_y0);
  fa fa_h_u_arrmul32_fa10_27_y2(h_u_arrmul32_and10_27_y0, h_u_arrmul32_fa11_26_y2, h_u_arrmul32_fa9_27_y4, h_u_arrmul32_fa10_27_y2, h_u_arrmul32_fa10_27_y4);
  and_gate and_gate_h_u_arrmul32_and11_27_y0(a_11, b_27, h_u_arrmul32_and11_27_y0);
  fa fa_h_u_arrmul32_fa11_27_y2(h_u_arrmul32_and11_27_y0, h_u_arrmul32_fa12_26_y2, h_u_arrmul32_fa10_27_y4, h_u_arrmul32_fa11_27_y2, h_u_arrmul32_fa11_27_y4);
  and_gate and_gate_h_u_arrmul32_and12_27_y0(a_12, b_27, h_u_arrmul32_and12_27_y0);
  fa fa_h_u_arrmul32_fa12_27_y2(h_u_arrmul32_and12_27_y0, h_u_arrmul32_fa13_26_y2, h_u_arrmul32_fa11_27_y4, h_u_arrmul32_fa12_27_y2, h_u_arrmul32_fa12_27_y4);
  and_gate and_gate_h_u_arrmul32_and13_27_y0(a_13, b_27, h_u_arrmul32_and13_27_y0);
  fa fa_h_u_arrmul32_fa13_27_y2(h_u_arrmul32_and13_27_y0, h_u_arrmul32_fa14_26_y2, h_u_arrmul32_fa12_27_y4, h_u_arrmul32_fa13_27_y2, h_u_arrmul32_fa13_27_y4);
  and_gate and_gate_h_u_arrmul32_and14_27_y0(a_14, b_27, h_u_arrmul32_and14_27_y0);
  fa fa_h_u_arrmul32_fa14_27_y2(h_u_arrmul32_and14_27_y0, h_u_arrmul32_fa15_26_y2, h_u_arrmul32_fa13_27_y4, h_u_arrmul32_fa14_27_y2, h_u_arrmul32_fa14_27_y4);
  and_gate and_gate_h_u_arrmul32_and15_27_y0(a_15, b_27, h_u_arrmul32_and15_27_y0);
  fa fa_h_u_arrmul32_fa15_27_y2(h_u_arrmul32_and15_27_y0, h_u_arrmul32_fa16_26_y2, h_u_arrmul32_fa14_27_y4, h_u_arrmul32_fa15_27_y2, h_u_arrmul32_fa15_27_y4);
  and_gate and_gate_h_u_arrmul32_and16_27_y0(a_16, b_27, h_u_arrmul32_and16_27_y0);
  fa fa_h_u_arrmul32_fa16_27_y2(h_u_arrmul32_and16_27_y0, h_u_arrmul32_fa17_26_y2, h_u_arrmul32_fa15_27_y4, h_u_arrmul32_fa16_27_y2, h_u_arrmul32_fa16_27_y4);
  and_gate and_gate_h_u_arrmul32_and17_27_y0(a_17, b_27, h_u_arrmul32_and17_27_y0);
  fa fa_h_u_arrmul32_fa17_27_y2(h_u_arrmul32_and17_27_y0, h_u_arrmul32_fa18_26_y2, h_u_arrmul32_fa16_27_y4, h_u_arrmul32_fa17_27_y2, h_u_arrmul32_fa17_27_y4);
  and_gate and_gate_h_u_arrmul32_and18_27_y0(a_18, b_27, h_u_arrmul32_and18_27_y0);
  fa fa_h_u_arrmul32_fa18_27_y2(h_u_arrmul32_and18_27_y0, h_u_arrmul32_fa19_26_y2, h_u_arrmul32_fa17_27_y4, h_u_arrmul32_fa18_27_y2, h_u_arrmul32_fa18_27_y4);
  and_gate and_gate_h_u_arrmul32_and19_27_y0(a_19, b_27, h_u_arrmul32_and19_27_y0);
  fa fa_h_u_arrmul32_fa19_27_y2(h_u_arrmul32_and19_27_y0, h_u_arrmul32_fa20_26_y2, h_u_arrmul32_fa18_27_y4, h_u_arrmul32_fa19_27_y2, h_u_arrmul32_fa19_27_y4);
  and_gate and_gate_h_u_arrmul32_and20_27_y0(a_20, b_27, h_u_arrmul32_and20_27_y0);
  fa fa_h_u_arrmul32_fa20_27_y2(h_u_arrmul32_and20_27_y0, h_u_arrmul32_fa21_26_y2, h_u_arrmul32_fa19_27_y4, h_u_arrmul32_fa20_27_y2, h_u_arrmul32_fa20_27_y4);
  and_gate and_gate_h_u_arrmul32_and21_27_y0(a_21, b_27, h_u_arrmul32_and21_27_y0);
  fa fa_h_u_arrmul32_fa21_27_y2(h_u_arrmul32_and21_27_y0, h_u_arrmul32_fa22_26_y2, h_u_arrmul32_fa20_27_y4, h_u_arrmul32_fa21_27_y2, h_u_arrmul32_fa21_27_y4);
  and_gate and_gate_h_u_arrmul32_and22_27_y0(a_22, b_27, h_u_arrmul32_and22_27_y0);
  fa fa_h_u_arrmul32_fa22_27_y2(h_u_arrmul32_and22_27_y0, h_u_arrmul32_fa23_26_y2, h_u_arrmul32_fa21_27_y4, h_u_arrmul32_fa22_27_y2, h_u_arrmul32_fa22_27_y4);
  and_gate and_gate_h_u_arrmul32_and23_27_y0(a_23, b_27, h_u_arrmul32_and23_27_y0);
  fa fa_h_u_arrmul32_fa23_27_y2(h_u_arrmul32_and23_27_y0, h_u_arrmul32_fa24_26_y2, h_u_arrmul32_fa22_27_y4, h_u_arrmul32_fa23_27_y2, h_u_arrmul32_fa23_27_y4);
  and_gate and_gate_h_u_arrmul32_and24_27_y0(a_24, b_27, h_u_arrmul32_and24_27_y0);
  fa fa_h_u_arrmul32_fa24_27_y2(h_u_arrmul32_and24_27_y0, h_u_arrmul32_fa25_26_y2, h_u_arrmul32_fa23_27_y4, h_u_arrmul32_fa24_27_y2, h_u_arrmul32_fa24_27_y4);
  and_gate and_gate_h_u_arrmul32_and25_27_y0(a_25, b_27, h_u_arrmul32_and25_27_y0);
  fa fa_h_u_arrmul32_fa25_27_y2(h_u_arrmul32_and25_27_y0, h_u_arrmul32_fa26_26_y2, h_u_arrmul32_fa24_27_y4, h_u_arrmul32_fa25_27_y2, h_u_arrmul32_fa25_27_y4);
  and_gate and_gate_h_u_arrmul32_and26_27_y0(a_26, b_27, h_u_arrmul32_and26_27_y0);
  fa fa_h_u_arrmul32_fa26_27_y2(h_u_arrmul32_and26_27_y0, h_u_arrmul32_fa27_26_y2, h_u_arrmul32_fa25_27_y4, h_u_arrmul32_fa26_27_y2, h_u_arrmul32_fa26_27_y4);
  and_gate and_gate_h_u_arrmul32_and27_27_y0(a_27, b_27, h_u_arrmul32_and27_27_y0);
  fa fa_h_u_arrmul32_fa27_27_y2(h_u_arrmul32_and27_27_y0, h_u_arrmul32_fa28_26_y2, h_u_arrmul32_fa26_27_y4, h_u_arrmul32_fa27_27_y2, h_u_arrmul32_fa27_27_y4);
  and_gate and_gate_h_u_arrmul32_and28_27_y0(a_28, b_27, h_u_arrmul32_and28_27_y0);
  fa fa_h_u_arrmul32_fa28_27_y2(h_u_arrmul32_and28_27_y0, h_u_arrmul32_fa29_26_y2, h_u_arrmul32_fa27_27_y4, h_u_arrmul32_fa28_27_y2, h_u_arrmul32_fa28_27_y4);
  and_gate and_gate_h_u_arrmul32_and29_27_y0(a_29, b_27, h_u_arrmul32_and29_27_y0);
  fa fa_h_u_arrmul32_fa29_27_y2(h_u_arrmul32_and29_27_y0, h_u_arrmul32_fa30_26_y2, h_u_arrmul32_fa28_27_y4, h_u_arrmul32_fa29_27_y2, h_u_arrmul32_fa29_27_y4);
  and_gate and_gate_h_u_arrmul32_and30_27_y0(a_30, b_27, h_u_arrmul32_and30_27_y0);
  fa fa_h_u_arrmul32_fa30_27_y2(h_u_arrmul32_and30_27_y0, h_u_arrmul32_fa31_26_y2, h_u_arrmul32_fa29_27_y4, h_u_arrmul32_fa30_27_y2, h_u_arrmul32_fa30_27_y4);
  and_gate and_gate_h_u_arrmul32_and31_27_y0(a_31, b_27, h_u_arrmul32_and31_27_y0);
  fa fa_h_u_arrmul32_fa31_27_y2(h_u_arrmul32_and31_27_y0, h_u_arrmul32_fa31_26_y4, h_u_arrmul32_fa30_27_y4, h_u_arrmul32_fa31_27_y2, h_u_arrmul32_fa31_27_y4);
  and_gate and_gate_h_u_arrmul32_and0_28_y0(a_0, b_28, h_u_arrmul32_and0_28_y0);
  ha ha_h_u_arrmul32_ha0_28_y0(h_u_arrmul32_and0_28_y0, h_u_arrmul32_fa1_27_y2, h_u_arrmul32_ha0_28_y0, h_u_arrmul32_ha0_28_y1);
  and_gate and_gate_h_u_arrmul32_and1_28_y0(a_1, b_28, h_u_arrmul32_and1_28_y0);
  fa fa_h_u_arrmul32_fa1_28_y2(h_u_arrmul32_and1_28_y0, h_u_arrmul32_fa2_27_y2, h_u_arrmul32_ha0_28_y1, h_u_arrmul32_fa1_28_y2, h_u_arrmul32_fa1_28_y4);
  and_gate and_gate_h_u_arrmul32_and2_28_y0(a_2, b_28, h_u_arrmul32_and2_28_y0);
  fa fa_h_u_arrmul32_fa2_28_y2(h_u_arrmul32_and2_28_y0, h_u_arrmul32_fa3_27_y2, h_u_arrmul32_fa1_28_y4, h_u_arrmul32_fa2_28_y2, h_u_arrmul32_fa2_28_y4);
  and_gate and_gate_h_u_arrmul32_and3_28_y0(a_3, b_28, h_u_arrmul32_and3_28_y0);
  fa fa_h_u_arrmul32_fa3_28_y2(h_u_arrmul32_and3_28_y0, h_u_arrmul32_fa4_27_y2, h_u_arrmul32_fa2_28_y4, h_u_arrmul32_fa3_28_y2, h_u_arrmul32_fa3_28_y4);
  and_gate and_gate_h_u_arrmul32_and4_28_y0(a_4, b_28, h_u_arrmul32_and4_28_y0);
  fa fa_h_u_arrmul32_fa4_28_y2(h_u_arrmul32_and4_28_y0, h_u_arrmul32_fa5_27_y2, h_u_arrmul32_fa3_28_y4, h_u_arrmul32_fa4_28_y2, h_u_arrmul32_fa4_28_y4);
  and_gate and_gate_h_u_arrmul32_and5_28_y0(a_5, b_28, h_u_arrmul32_and5_28_y0);
  fa fa_h_u_arrmul32_fa5_28_y2(h_u_arrmul32_and5_28_y0, h_u_arrmul32_fa6_27_y2, h_u_arrmul32_fa4_28_y4, h_u_arrmul32_fa5_28_y2, h_u_arrmul32_fa5_28_y4);
  and_gate and_gate_h_u_arrmul32_and6_28_y0(a_6, b_28, h_u_arrmul32_and6_28_y0);
  fa fa_h_u_arrmul32_fa6_28_y2(h_u_arrmul32_and6_28_y0, h_u_arrmul32_fa7_27_y2, h_u_arrmul32_fa5_28_y4, h_u_arrmul32_fa6_28_y2, h_u_arrmul32_fa6_28_y4);
  and_gate and_gate_h_u_arrmul32_and7_28_y0(a_7, b_28, h_u_arrmul32_and7_28_y0);
  fa fa_h_u_arrmul32_fa7_28_y2(h_u_arrmul32_and7_28_y0, h_u_arrmul32_fa8_27_y2, h_u_arrmul32_fa6_28_y4, h_u_arrmul32_fa7_28_y2, h_u_arrmul32_fa7_28_y4);
  and_gate and_gate_h_u_arrmul32_and8_28_y0(a_8, b_28, h_u_arrmul32_and8_28_y0);
  fa fa_h_u_arrmul32_fa8_28_y2(h_u_arrmul32_and8_28_y0, h_u_arrmul32_fa9_27_y2, h_u_arrmul32_fa7_28_y4, h_u_arrmul32_fa8_28_y2, h_u_arrmul32_fa8_28_y4);
  and_gate and_gate_h_u_arrmul32_and9_28_y0(a_9, b_28, h_u_arrmul32_and9_28_y0);
  fa fa_h_u_arrmul32_fa9_28_y2(h_u_arrmul32_and9_28_y0, h_u_arrmul32_fa10_27_y2, h_u_arrmul32_fa8_28_y4, h_u_arrmul32_fa9_28_y2, h_u_arrmul32_fa9_28_y4);
  and_gate and_gate_h_u_arrmul32_and10_28_y0(a_10, b_28, h_u_arrmul32_and10_28_y0);
  fa fa_h_u_arrmul32_fa10_28_y2(h_u_arrmul32_and10_28_y0, h_u_arrmul32_fa11_27_y2, h_u_arrmul32_fa9_28_y4, h_u_arrmul32_fa10_28_y2, h_u_arrmul32_fa10_28_y4);
  and_gate and_gate_h_u_arrmul32_and11_28_y0(a_11, b_28, h_u_arrmul32_and11_28_y0);
  fa fa_h_u_arrmul32_fa11_28_y2(h_u_arrmul32_and11_28_y0, h_u_arrmul32_fa12_27_y2, h_u_arrmul32_fa10_28_y4, h_u_arrmul32_fa11_28_y2, h_u_arrmul32_fa11_28_y4);
  and_gate and_gate_h_u_arrmul32_and12_28_y0(a_12, b_28, h_u_arrmul32_and12_28_y0);
  fa fa_h_u_arrmul32_fa12_28_y2(h_u_arrmul32_and12_28_y0, h_u_arrmul32_fa13_27_y2, h_u_arrmul32_fa11_28_y4, h_u_arrmul32_fa12_28_y2, h_u_arrmul32_fa12_28_y4);
  and_gate and_gate_h_u_arrmul32_and13_28_y0(a_13, b_28, h_u_arrmul32_and13_28_y0);
  fa fa_h_u_arrmul32_fa13_28_y2(h_u_arrmul32_and13_28_y0, h_u_arrmul32_fa14_27_y2, h_u_arrmul32_fa12_28_y4, h_u_arrmul32_fa13_28_y2, h_u_arrmul32_fa13_28_y4);
  and_gate and_gate_h_u_arrmul32_and14_28_y0(a_14, b_28, h_u_arrmul32_and14_28_y0);
  fa fa_h_u_arrmul32_fa14_28_y2(h_u_arrmul32_and14_28_y0, h_u_arrmul32_fa15_27_y2, h_u_arrmul32_fa13_28_y4, h_u_arrmul32_fa14_28_y2, h_u_arrmul32_fa14_28_y4);
  and_gate and_gate_h_u_arrmul32_and15_28_y0(a_15, b_28, h_u_arrmul32_and15_28_y0);
  fa fa_h_u_arrmul32_fa15_28_y2(h_u_arrmul32_and15_28_y0, h_u_arrmul32_fa16_27_y2, h_u_arrmul32_fa14_28_y4, h_u_arrmul32_fa15_28_y2, h_u_arrmul32_fa15_28_y4);
  and_gate and_gate_h_u_arrmul32_and16_28_y0(a_16, b_28, h_u_arrmul32_and16_28_y0);
  fa fa_h_u_arrmul32_fa16_28_y2(h_u_arrmul32_and16_28_y0, h_u_arrmul32_fa17_27_y2, h_u_arrmul32_fa15_28_y4, h_u_arrmul32_fa16_28_y2, h_u_arrmul32_fa16_28_y4);
  and_gate and_gate_h_u_arrmul32_and17_28_y0(a_17, b_28, h_u_arrmul32_and17_28_y0);
  fa fa_h_u_arrmul32_fa17_28_y2(h_u_arrmul32_and17_28_y0, h_u_arrmul32_fa18_27_y2, h_u_arrmul32_fa16_28_y4, h_u_arrmul32_fa17_28_y2, h_u_arrmul32_fa17_28_y4);
  and_gate and_gate_h_u_arrmul32_and18_28_y0(a_18, b_28, h_u_arrmul32_and18_28_y0);
  fa fa_h_u_arrmul32_fa18_28_y2(h_u_arrmul32_and18_28_y0, h_u_arrmul32_fa19_27_y2, h_u_arrmul32_fa17_28_y4, h_u_arrmul32_fa18_28_y2, h_u_arrmul32_fa18_28_y4);
  and_gate and_gate_h_u_arrmul32_and19_28_y0(a_19, b_28, h_u_arrmul32_and19_28_y0);
  fa fa_h_u_arrmul32_fa19_28_y2(h_u_arrmul32_and19_28_y0, h_u_arrmul32_fa20_27_y2, h_u_arrmul32_fa18_28_y4, h_u_arrmul32_fa19_28_y2, h_u_arrmul32_fa19_28_y4);
  and_gate and_gate_h_u_arrmul32_and20_28_y0(a_20, b_28, h_u_arrmul32_and20_28_y0);
  fa fa_h_u_arrmul32_fa20_28_y2(h_u_arrmul32_and20_28_y0, h_u_arrmul32_fa21_27_y2, h_u_arrmul32_fa19_28_y4, h_u_arrmul32_fa20_28_y2, h_u_arrmul32_fa20_28_y4);
  and_gate and_gate_h_u_arrmul32_and21_28_y0(a_21, b_28, h_u_arrmul32_and21_28_y0);
  fa fa_h_u_arrmul32_fa21_28_y2(h_u_arrmul32_and21_28_y0, h_u_arrmul32_fa22_27_y2, h_u_arrmul32_fa20_28_y4, h_u_arrmul32_fa21_28_y2, h_u_arrmul32_fa21_28_y4);
  and_gate and_gate_h_u_arrmul32_and22_28_y0(a_22, b_28, h_u_arrmul32_and22_28_y0);
  fa fa_h_u_arrmul32_fa22_28_y2(h_u_arrmul32_and22_28_y0, h_u_arrmul32_fa23_27_y2, h_u_arrmul32_fa21_28_y4, h_u_arrmul32_fa22_28_y2, h_u_arrmul32_fa22_28_y4);
  and_gate and_gate_h_u_arrmul32_and23_28_y0(a_23, b_28, h_u_arrmul32_and23_28_y0);
  fa fa_h_u_arrmul32_fa23_28_y2(h_u_arrmul32_and23_28_y0, h_u_arrmul32_fa24_27_y2, h_u_arrmul32_fa22_28_y4, h_u_arrmul32_fa23_28_y2, h_u_arrmul32_fa23_28_y4);
  and_gate and_gate_h_u_arrmul32_and24_28_y0(a_24, b_28, h_u_arrmul32_and24_28_y0);
  fa fa_h_u_arrmul32_fa24_28_y2(h_u_arrmul32_and24_28_y0, h_u_arrmul32_fa25_27_y2, h_u_arrmul32_fa23_28_y4, h_u_arrmul32_fa24_28_y2, h_u_arrmul32_fa24_28_y4);
  and_gate and_gate_h_u_arrmul32_and25_28_y0(a_25, b_28, h_u_arrmul32_and25_28_y0);
  fa fa_h_u_arrmul32_fa25_28_y2(h_u_arrmul32_and25_28_y0, h_u_arrmul32_fa26_27_y2, h_u_arrmul32_fa24_28_y4, h_u_arrmul32_fa25_28_y2, h_u_arrmul32_fa25_28_y4);
  and_gate and_gate_h_u_arrmul32_and26_28_y0(a_26, b_28, h_u_arrmul32_and26_28_y0);
  fa fa_h_u_arrmul32_fa26_28_y2(h_u_arrmul32_and26_28_y0, h_u_arrmul32_fa27_27_y2, h_u_arrmul32_fa25_28_y4, h_u_arrmul32_fa26_28_y2, h_u_arrmul32_fa26_28_y4);
  and_gate and_gate_h_u_arrmul32_and27_28_y0(a_27, b_28, h_u_arrmul32_and27_28_y0);
  fa fa_h_u_arrmul32_fa27_28_y2(h_u_arrmul32_and27_28_y0, h_u_arrmul32_fa28_27_y2, h_u_arrmul32_fa26_28_y4, h_u_arrmul32_fa27_28_y2, h_u_arrmul32_fa27_28_y4);
  and_gate and_gate_h_u_arrmul32_and28_28_y0(a_28, b_28, h_u_arrmul32_and28_28_y0);
  fa fa_h_u_arrmul32_fa28_28_y2(h_u_arrmul32_and28_28_y0, h_u_arrmul32_fa29_27_y2, h_u_arrmul32_fa27_28_y4, h_u_arrmul32_fa28_28_y2, h_u_arrmul32_fa28_28_y4);
  and_gate and_gate_h_u_arrmul32_and29_28_y0(a_29, b_28, h_u_arrmul32_and29_28_y0);
  fa fa_h_u_arrmul32_fa29_28_y2(h_u_arrmul32_and29_28_y0, h_u_arrmul32_fa30_27_y2, h_u_arrmul32_fa28_28_y4, h_u_arrmul32_fa29_28_y2, h_u_arrmul32_fa29_28_y4);
  and_gate and_gate_h_u_arrmul32_and30_28_y0(a_30, b_28, h_u_arrmul32_and30_28_y0);
  fa fa_h_u_arrmul32_fa30_28_y2(h_u_arrmul32_and30_28_y0, h_u_arrmul32_fa31_27_y2, h_u_arrmul32_fa29_28_y4, h_u_arrmul32_fa30_28_y2, h_u_arrmul32_fa30_28_y4);
  and_gate and_gate_h_u_arrmul32_and31_28_y0(a_31, b_28, h_u_arrmul32_and31_28_y0);
  fa fa_h_u_arrmul32_fa31_28_y2(h_u_arrmul32_and31_28_y0, h_u_arrmul32_fa31_27_y4, h_u_arrmul32_fa30_28_y4, h_u_arrmul32_fa31_28_y2, h_u_arrmul32_fa31_28_y4);
  and_gate and_gate_h_u_arrmul32_and0_29_y0(a_0, b_29, h_u_arrmul32_and0_29_y0);
  ha ha_h_u_arrmul32_ha0_29_y0(h_u_arrmul32_and0_29_y0, h_u_arrmul32_fa1_28_y2, h_u_arrmul32_ha0_29_y0, h_u_arrmul32_ha0_29_y1);
  and_gate and_gate_h_u_arrmul32_and1_29_y0(a_1, b_29, h_u_arrmul32_and1_29_y0);
  fa fa_h_u_arrmul32_fa1_29_y2(h_u_arrmul32_and1_29_y0, h_u_arrmul32_fa2_28_y2, h_u_arrmul32_ha0_29_y1, h_u_arrmul32_fa1_29_y2, h_u_arrmul32_fa1_29_y4);
  and_gate and_gate_h_u_arrmul32_and2_29_y0(a_2, b_29, h_u_arrmul32_and2_29_y0);
  fa fa_h_u_arrmul32_fa2_29_y2(h_u_arrmul32_and2_29_y0, h_u_arrmul32_fa3_28_y2, h_u_arrmul32_fa1_29_y4, h_u_arrmul32_fa2_29_y2, h_u_arrmul32_fa2_29_y4);
  and_gate and_gate_h_u_arrmul32_and3_29_y0(a_3, b_29, h_u_arrmul32_and3_29_y0);
  fa fa_h_u_arrmul32_fa3_29_y2(h_u_arrmul32_and3_29_y0, h_u_arrmul32_fa4_28_y2, h_u_arrmul32_fa2_29_y4, h_u_arrmul32_fa3_29_y2, h_u_arrmul32_fa3_29_y4);
  and_gate and_gate_h_u_arrmul32_and4_29_y0(a_4, b_29, h_u_arrmul32_and4_29_y0);
  fa fa_h_u_arrmul32_fa4_29_y2(h_u_arrmul32_and4_29_y0, h_u_arrmul32_fa5_28_y2, h_u_arrmul32_fa3_29_y4, h_u_arrmul32_fa4_29_y2, h_u_arrmul32_fa4_29_y4);
  and_gate and_gate_h_u_arrmul32_and5_29_y0(a_5, b_29, h_u_arrmul32_and5_29_y0);
  fa fa_h_u_arrmul32_fa5_29_y2(h_u_arrmul32_and5_29_y0, h_u_arrmul32_fa6_28_y2, h_u_arrmul32_fa4_29_y4, h_u_arrmul32_fa5_29_y2, h_u_arrmul32_fa5_29_y4);
  and_gate and_gate_h_u_arrmul32_and6_29_y0(a_6, b_29, h_u_arrmul32_and6_29_y0);
  fa fa_h_u_arrmul32_fa6_29_y2(h_u_arrmul32_and6_29_y0, h_u_arrmul32_fa7_28_y2, h_u_arrmul32_fa5_29_y4, h_u_arrmul32_fa6_29_y2, h_u_arrmul32_fa6_29_y4);
  and_gate and_gate_h_u_arrmul32_and7_29_y0(a_7, b_29, h_u_arrmul32_and7_29_y0);
  fa fa_h_u_arrmul32_fa7_29_y2(h_u_arrmul32_and7_29_y0, h_u_arrmul32_fa8_28_y2, h_u_arrmul32_fa6_29_y4, h_u_arrmul32_fa7_29_y2, h_u_arrmul32_fa7_29_y4);
  and_gate and_gate_h_u_arrmul32_and8_29_y0(a_8, b_29, h_u_arrmul32_and8_29_y0);
  fa fa_h_u_arrmul32_fa8_29_y2(h_u_arrmul32_and8_29_y0, h_u_arrmul32_fa9_28_y2, h_u_arrmul32_fa7_29_y4, h_u_arrmul32_fa8_29_y2, h_u_arrmul32_fa8_29_y4);
  and_gate and_gate_h_u_arrmul32_and9_29_y0(a_9, b_29, h_u_arrmul32_and9_29_y0);
  fa fa_h_u_arrmul32_fa9_29_y2(h_u_arrmul32_and9_29_y0, h_u_arrmul32_fa10_28_y2, h_u_arrmul32_fa8_29_y4, h_u_arrmul32_fa9_29_y2, h_u_arrmul32_fa9_29_y4);
  and_gate and_gate_h_u_arrmul32_and10_29_y0(a_10, b_29, h_u_arrmul32_and10_29_y0);
  fa fa_h_u_arrmul32_fa10_29_y2(h_u_arrmul32_and10_29_y0, h_u_arrmul32_fa11_28_y2, h_u_arrmul32_fa9_29_y4, h_u_arrmul32_fa10_29_y2, h_u_arrmul32_fa10_29_y4);
  and_gate and_gate_h_u_arrmul32_and11_29_y0(a_11, b_29, h_u_arrmul32_and11_29_y0);
  fa fa_h_u_arrmul32_fa11_29_y2(h_u_arrmul32_and11_29_y0, h_u_arrmul32_fa12_28_y2, h_u_arrmul32_fa10_29_y4, h_u_arrmul32_fa11_29_y2, h_u_arrmul32_fa11_29_y4);
  and_gate and_gate_h_u_arrmul32_and12_29_y0(a_12, b_29, h_u_arrmul32_and12_29_y0);
  fa fa_h_u_arrmul32_fa12_29_y2(h_u_arrmul32_and12_29_y0, h_u_arrmul32_fa13_28_y2, h_u_arrmul32_fa11_29_y4, h_u_arrmul32_fa12_29_y2, h_u_arrmul32_fa12_29_y4);
  and_gate and_gate_h_u_arrmul32_and13_29_y0(a_13, b_29, h_u_arrmul32_and13_29_y0);
  fa fa_h_u_arrmul32_fa13_29_y2(h_u_arrmul32_and13_29_y0, h_u_arrmul32_fa14_28_y2, h_u_arrmul32_fa12_29_y4, h_u_arrmul32_fa13_29_y2, h_u_arrmul32_fa13_29_y4);
  and_gate and_gate_h_u_arrmul32_and14_29_y0(a_14, b_29, h_u_arrmul32_and14_29_y0);
  fa fa_h_u_arrmul32_fa14_29_y2(h_u_arrmul32_and14_29_y0, h_u_arrmul32_fa15_28_y2, h_u_arrmul32_fa13_29_y4, h_u_arrmul32_fa14_29_y2, h_u_arrmul32_fa14_29_y4);
  and_gate and_gate_h_u_arrmul32_and15_29_y0(a_15, b_29, h_u_arrmul32_and15_29_y0);
  fa fa_h_u_arrmul32_fa15_29_y2(h_u_arrmul32_and15_29_y0, h_u_arrmul32_fa16_28_y2, h_u_arrmul32_fa14_29_y4, h_u_arrmul32_fa15_29_y2, h_u_arrmul32_fa15_29_y4);
  and_gate and_gate_h_u_arrmul32_and16_29_y0(a_16, b_29, h_u_arrmul32_and16_29_y0);
  fa fa_h_u_arrmul32_fa16_29_y2(h_u_arrmul32_and16_29_y0, h_u_arrmul32_fa17_28_y2, h_u_arrmul32_fa15_29_y4, h_u_arrmul32_fa16_29_y2, h_u_arrmul32_fa16_29_y4);
  and_gate and_gate_h_u_arrmul32_and17_29_y0(a_17, b_29, h_u_arrmul32_and17_29_y0);
  fa fa_h_u_arrmul32_fa17_29_y2(h_u_arrmul32_and17_29_y0, h_u_arrmul32_fa18_28_y2, h_u_arrmul32_fa16_29_y4, h_u_arrmul32_fa17_29_y2, h_u_arrmul32_fa17_29_y4);
  and_gate and_gate_h_u_arrmul32_and18_29_y0(a_18, b_29, h_u_arrmul32_and18_29_y0);
  fa fa_h_u_arrmul32_fa18_29_y2(h_u_arrmul32_and18_29_y0, h_u_arrmul32_fa19_28_y2, h_u_arrmul32_fa17_29_y4, h_u_arrmul32_fa18_29_y2, h_u_arrmul32_fa18_29_y4);
  and_gate and_gate_h_u_arrmul32_and19_29_y0(a_19, b_29, h_u_arrmul32_and19_29_y0);
  fa fa_h_u_arrmul32_fa19_29_y2(h_u_arrmul32_and19_29_y0, h_u_arrmul32_fa20_28_y2, h_u_arrmul32_fa18_29_y4, h_u_arrmul32_fa19_29_y2, h_u_arrmul32_fa19_29_y4);
  and_gate and_gate_h_u_arrmul32_and20_29_y0(a_20, b_29, h_u_arrmul32_and20_29_y0);
  fa fa_h_u_arrmul32_fa20_29_y2(h_u_arrmul32_and20_29_y0, h_u_arrmul32_fa21_28_y2, h_u_arrmul32_fa19_29_y4, h_u_arrmul32_fa20_29_y2, h_u_arrmul32_fa20_29_y4);
  and_gate and_gate_h_u_arrmul32_and21_29_y0(a_21, b_29, h_u_arrmul32_and21_29_y0);
  fa fa_h_u_arrmul32_fa21_29_y2(h_u_arrmul32_and21_29_y0, h_u_arrmul32_fa22_28_y2, h_u_arrmul32_fa20_29_y4, h_u_arrmul32_fa21_29_y2, h_u_arrmul32_fa21_29_y4);
  and_gate and_gate_h_u_arrmul32_and22_29_y0(a_22, b_29, h_u_arrmul32_and22_29_y0);
  fa fa_h_u_arrmul32_fa22_29_y2(h_u_arrmul32_and22_29_y0, h_u_arrmul32_fa23_28_y2, h_u_arrmul32_fa21_29_y4, h_u_arrmul32_fa22_29_y2, h_u_arrmul32_fa22_29_y4);
  and_gate and_gate_h_u_arrmul32_and23_29_y0(a_23, b_29, h_u_arrmul32_and23_29_y0);
  fa fa_h_u_arrmul32_fa23_29_y2(h_u_arrmul32_and23_29_y0, h_u_arrmul32_fa24_28_y2, h_u_arrmul32_fa22_29_y4, h_u_arrmul32_fa23_29_y2, h_u_arrmul32_fa23_29_y4);
  and_gate and_gate_h_u_arrmul32_and24_29_y0(a_24, b_29, h_u_arrmul32_and24_29_y0);
  fa fa_h_u_arrmul32_fa24_29_y2(h_u_arrmul32_and24_29_y0, h_u_arrmul32_fa25_28_y2, h_u_arrmul32_fa23_29_y4, h_u_arrmul32_fa24_29_y2, h_u_arrmul32_fa24_29_y4);
  and_gate and_gate_h_u_arrmul32_and25_29_y0(a_25, b_29, h_u_arrmul32_and25_29_y0);
  fa fa_h_u_arrmul32_fa25_29_y2(h_u_arrmul32_and25_29_y0, h_u_arrmul32_fa26_28_y2, h_u_arrmul32_fa24_29_y4, h_u_arrmul32_fa25_29_y2, h_u_arrmul32_fa25_29_y4);
  and_gate and_gate_h_u_arrmul32_and26_29_y0(a_26, b_29, h_u_arrmul32_and26_29_y0);
  fa fa_h_u_arrmul32_fa26_29_y2(h_u_arrmul32_and26_29_y0, h_u_arrmul32_fa27_28_y2, h_u_arrmul32_fa25_29_y4, h_u_arrmul32_fa26_29_y2, h_u_arrmul32_fa26_29_y4);
  and_gate and_gate_h_u_arrmul32_and27_29_y0(a_27, b_29, h_u_arrmul32_and27_29_y0);
  fa fa_h_u_arrmul32_fa27_29_y2(h_u_arrmul32_and27_29_y0, h_u_arrmul32_fa28_28_y2, h_u_arrmul32_fa26_29_y4, h_u_arrmul32_fa27_29_y2, h_u_arrmul32_fa27_29_y4);
  and_gate and_gate_h_u_arrmul32_and28_29_y0(a_28, b_29, h_u_arrmul32_and28_29_y0);
  fa fa_h_u_arrmul32_fa28_29_y2(h_u_arrmul32_and28_29_y0, h_u_arrmul32_fa29_28_y2, h_u_arrmul32_fa27_29_y4, h_u_arrmul32_fa28_29_y2, h_u_arrmul32_fa28_29_y4);
  and_gate and_gate_h_u_arrmul32_and29_29_y0(a_29, b_29, h_u_arrmul32_and29_29_y0);
  fa fa_h_u_arrmul32_fa29_29_y2(h_u_arrmul32_and29_29_y0, h_u_arrmul32_fa30_28_y2, h_u_arrmul32_fa28_29_y4, h_u_arrmul32_fa29_29_y2, h_u_arrmul32_fa29_29_y4);
  and_gate and_gate_h_u_arrmul32_and30_29_y0(a_30, b_29, h_u_arrmul32_and30_29_y0);
  fa fa_h_u_arrmul32_fa30_29_y2(h_u_arrmul32_and30_29_y0, h_u_arrmul32_fa31_28_y2, h_u_arrmul32_fa29_29_y4, h_u_arrmul32_fa30_29_y2, h_u_arrmul32_fa30_29_y4);
  and_gate and_gate_h_u_arrmul32_and31_29_y0(a_31, b_29, h_u_arrmul32_and31_29_y0);
  fa fa_h_u_arrmul32_fa31_29_y2(h_u_arrmul32_and31_29_y0, h_u_arrmul32_fa31_28_y4, h_u_arrmul32_fa30_29_y4, h_u_arrmul32_fa31_29_y2, h_u_arrmul32_fa31_29_y4);
  and_gate and_gate_h_u_arrmul32_and0_30_y0(a_0, b_30, h_u_arrmul32_and0_30_y0);
  ha ha_h_u_arrmul32_ha0_30_y0(h_u_arrmul32_and0_30_y0, h_u_arrmul32_fa1_29_y2, h_u_arrmul32_ha0_30_y0, h_u_arrmul32_ha0_30_y1);
  and_gate and_gate_h_u_arrmul32_and1_30_y0(a_1, b_30, h_u_arrmul32_and1_30_y0);
  fa fa_h_u_arrmul32_fa1_30_y2(h_u_arrmul32_and1_30_y0, h_u_arrmul32_fa2_29_y2, h_u_arrmul32_ha0_30_y1, h_u_arrmul32_fa1_30_y2, h_u_arrmul32_fa1_30_y4);
  and_gate and_gate_h_u_arrmul32_and2_30_y0(a_2, b_30, h_u_arrmul32_and2_30_y0);
  fa fa_h_u_arrmul32_fa2_30_y2(h_u_arrmul32_and2_30_y0, h_u_arrmul32_fa3_29_y2, h_u_arrmul32_fa1_30_y4, h_u_arrmul32_fa2_30_y2, h_u_arrmul32_fa2_30_y4);
  and_gate and_gate_h_u_arrmul32_and3_30_y0(a_3, b_30, h_u_arrmul32_and3_30_y0);
  fa fa_h_u_arrmul32_fa3_30_y2(h_u_arrmul32_and3_30_y0, h_u_arrmul32_fa4_29_y2, h_u_arrmul32_fa2_30_y4, h_u_arrmul32_fa3_30_y2, h_u_arrmul32_fa3_30_y4);
  and_gate and_gate_h_u_arrmul32_and4_30_y0(a_4, b_30, h_u_arrmul32_and4_30_y0);
  fa fa_h_u_arrmul32_fa4_30_y2(h_u_arrmul32_and4_30_y0, h_u_arrmul32_fa5_29_y2, h_u_arrmul32_fa3_30_y4, h_u_arrmul32_fa4_30_y2, h_u_arrmul32_fa4_30_y4);
  and_gate and_gate_h_u_arrmul32_and5_30_y0(a_5, b_30, h_u_arrmul32_and5_30_y0);
  fa fa_h_u_arrmul32_fa5_30_y2(h_u_arrmul32_and5_30_y0, h_u_arrmul32_fa6_29_y2, h_u_arrmul32_fa4_30_y4, h_u_arrmul32_fa5_30_y2, h_u_arrmul32_fa5_30_y4);
  and_gate and_gate_h_u_arrmul32_and6_30_y0(a_6, b_30, h_u_arrmul32_and6_30_y0);
  fa fa_h_u_arrmul32_fa6_30_y2(h_u_arrmul32_and6_30_y0, h_u_arrmul32_fa7_29_y2, h_u_arrmul32_fa5_30_y4, h_u_arrmul32_fa6_30_y2, h_u_arrmul32_fa6_30_y4);
  and_gate and_gate_h_u_arrmul32_and7_30_y0(a_7, b_30, h_u_arrmul32_and7_30_y0);
  fa fa_h_u_arrmul32_fa7_30_y2(h_u_arrmul32_and7_30_y0, h_u_arrmul32_fa8_29_y2, h_u_arrmul32_fa6_30_y4, h_u_arrmul32_fa7_30_y2, h_u_arrmul32_fa7_30_y4);
  and_gate and_gate_h_u_arrmul32_and8_30_y0(a_8, b_30, h_u_arrmul32_and8_30_y0);
  fa fa_h_u_arrmul32_fa8_30_y2(h_u_arrmul32_and8_30_y0, h_u_arrmul32_fa9_29_y2, h_u_arrmul32_fa7_30_y4, h_u_arrmul32_fa8_30_y2, h_u_arrmul32_fa8_30_y4);
  and_gate and_gate_h_u_arrmul32_and9_30_y0(a_9, b_30, h_u_arrmul32_and9_30_y0);
  fa fa_h_u_arrmul32_fa9_30_y2(h_u_arrmul32_and9_30_y0, h_u_arrmul32_fa10_29_y2, h_u_arrmul32_fa8_30_y4, h_u_arrmul32_fa9_30_y2, h_u_arrmul32_fa9_30_y4);
  and_gate and_gate_h_u_arrmul32_and10_30_y0(a_10, b_30, h_u_arrmul32_and10_30_y0);
  fa fa_h_u_arrmul32_fa10_30_y2(h_u_arrmul32_and10_30_y0, h_u_arrmul32_fa11_29_y2, h_u_arrmul32_fa9_30_y4, h_u_arrmul32_fa10_30_y2, h_u_arrmul32_fa10_30_y4);
  and_gate and_gate_h_u_arrmul32_and11_30_y0(a_11, b_30, h_u_arrmul32_and11_30_y0);
  fa fa_h_u_arrmul32_fa11_30_y2(h_u_arrmul32_and11_30_y0, h_u_arrmul32_fa12_29_y2, h_u_arrmul32_fa10_30_y4, h_u_arrmul32_fa11_30_y2, h_u_arrmul32_fa11_30_y4);
  and_gate and_gate_h_u_arrmul32_and12_30_y0(a_12, b_30, h_u_arrmul32_and12_30_y0);
  fa fa_h_u_arrmul32_fa12_30_y2(h_u_arrmul32_and12_30_y0, h_u_arrmul32_fa13_29_y2, h_u_arrmul32_fa11_30_y4, h_u_arrmul32_fa12_30_y2, h_u_arrmul32_fa12_30_y4);
  and_gate and_gate_h_u_arrmul32_and13_30_y0(a_13, b_30, h_u_arrmul32_and13_30_y0);
  fa fa_h_u_arrmul32_fa13_30_y2(h_u_arrmul32_and13_30_y0, h_u_arrmul32_fa14_29_y2, h_u_arrmul32_fa12_30_y4, h_u_arrmul32_fa13_30_y2, h_u_arrmul32_fa13_30_y4);
  and_gate and_gate_h_u_arrmul32_and14_30_y0(a_14, b_30, h_u_arrmul32_and14_30_y0);
  fa fa_h_u_arrmul32_fa14_30_y2(h_u_arrmul32_and14_30_y0, h_u_arrmul32_fa15_29_y2, h_u_arrmul32_fa13_30_y4, h_u_arrmul32_fa14_30_y2, h_u_arrmul32_fa14_30_y4);
  and_gate and_gate_h_u_arrmul32_and15_30_y0(a_15, b_30, h_u_arrmul32_and15_30_y0);
  fa fa_h_u_arrmul32_fa15_30_y2(h_u_arrmul32_and15_30_y0, h_u_arrmul32_fa16_29_y2, h_u_arrmul32_fa14_30_y4, h_u_arrmul32_fa15_30_y2, h_u_arrmul32_fa15_30_y4);
  and_gate and_gate_h_u_arrmul32_and16_30_y0(a_16, b_30, h_u_arrmul32_and16_30_y0);
  fa fa_h_u_arrmul32_fa16_30_y2(h_u_arrmul32_and16_30_y0, h_u_arrmul32_fa17_29_y2, h_u_arrmul32_fa15_30_y4, h_u_arrmul32_fa16_30_y2, h_u_arrmul32_fa16_30_y4);
  and_gate and_gate_h_u_arrmul32_and17_30_y0(a_17, b_30, h_u_arrmul32_and17_30_y0);
  fa fa_h_u_arrmul32_fa17_30_y2(h_u_arrmul32_and17_30_y0, h_u_arrmul32_fa18_29_y2, h_u_arrmul32_fa16_30_y4, h_u_arrmul32_fa17_30_y2, h_u_arrmul32_fa17_30_y4);
  and_gate and_gate_h_u_arrmul32_and18_30_y0(a_18, b_30, h_u_arrmul32_and18_30_y0);
  fa fa_h_u_arrmul32_fa18_30_y2(h_u_arrmul32_and18_30_y0, h_u_arrmul32_fa19_29_y2, h_u_arrmul32_fa17_30_y4, h_u_arrmul32_fa18_30_y2, h_u_arrmul32_fa18_30_y4);
  and_gate and_gate_h_u_arrmul32_and19_30_y0(a_19, b_30, h_u_arrmul32_and19_30_y0);
  fa fa_h_u_arrmul32_fa19_30_y2(h_u_arrmul32_and19_30_y0, h_u_arrmul32_fa20_29_y2, h_u_arrmul32_fa18_30_y4, h_u_arrmul32_fa19_30_y2, h_u_arrmul32_fa19_30_y4);
  and_gate and_gate_h_u_arrmul32_and20_30_y0(a_20, b_30, h_u_arrmul32_and20_30_y0);
  fa fa_h_u_arrmul32_fa20_30_y2(h_u_arrmul32_and20_30_y0, h_u_arrmul32_fa21_29_y2, h_u_arrmul32_fa19_30_y4, h_u_arrmul32_fa20_30_y2, h_u_arrmul32_fa20_30_y4);
  and_gate and_gate_h_u_arrmul32_and21_30_y0(a_21, b_30, h_u_arrmul32_and21_30_y0);
  fa fa_h_u_arrmul32_fa21_30_y2(h_u_arrmul32_and21_30_y0, h_u_arrmul32_fa22_29_y2, h_u_arrmul32_fa20_30_y4, h_u_arrmul32_fa21_30_y2, h_u_arrmul32_fa21_30_y4);
  and_gate and_gate_h_u_arrmul32_and22_30_y0(a_22, b_30, h_u_arrmul32_and22_30_y0);
  fa fa_h_u_arrmul32_fa22_30_y2(h_u_arrmul32_and22_30_y0, h_u_arrmul32_fa23_29_y2, h_u_arrmul32_fa21_30_y4, h_u_arrmul32_fa22_30_y2, h_u_arrmul32_fa22_30_y4);
  and_gate and_gate_h_u_arrmul32_and23_30_y0(a_23, b_30, h_u_arrmul32_and23_30_y0);
  fa fa_h_u_arrmul32_fa23_30_y2(h_u_arrmul32_and23_30_y0, h_u_arrmul32_fa24_29_y2, h_u_arrmul32_fa22_30_y4, h_u_arrmul32_fa23_30_y2, h_u_arrmul32_fa23_30_y4);
  and_gate and_gate_h_u_arrmul32_and24_30_y0(a_24, b_30, h_u_arrmul32_and24_30_y0);
  fa fa_h_u_arrmul32_fa24_30_y2(h_u_arrmul32_and24_30_y0, h_u_arrmul32_fa25_29_y2, h_u_arrmul32_fa23_30_y4, h_u_arrmul32_fa24_30_y2, h_u_arrmul32_fa24_30_y4);
  and_gate and_gate_h_u_arrmul32_and25_30_y0(a_25, b_30, h_u_arrmul32_and25_30_y0);
  fa fa_h_u_arrmul32_fa25_30_y2(h_u_arrmul32_and25_30_y0, h_u_arrmul32_fa26_29_y2, h_u_arrmul32_fa24_30_y4, h_u_arrmul32_fa25_30_y2, h_u_arrmul32_fa25_30_y4);
  and_gate and_gate_h_u_arrmul32_and26_30_y0(a_26, b_30, h_u_arrmul32_and26_30_y0);
  fa fa_h_u_arrmul32_fa26_30_y2(h_u_arrmul32_and26_30_y0, h_u_arrmul32_fa27_29_y2, h_u_arrmul32_fa25_30_y4, h_u_arrmul32_fa26_30_y2, h_u_arrmul32_fa26_30_y4);
  and_gate and_gate_h_u_arrmul32_and27_30_y0(a_27, b_30, h_u_arrmul32_and27_30_y0);
  fa fa_h_u_arrmul32_fa27_30_y2(h_u_arrmul32_and27_30_y0, h_u_arrmul32_fa28_29_y2, h_u_arrmul32_fa26_30_y4, h_u_arrmul32_fa27_30_y2, h_u_arrmul32_fa27_30_y4);
  and_gate and_gate_h_u_arrmul32_and28_30_y0(a_28, b_30, h_u_arrmul32_and28_30_y0);
  fa fa_h_u_arrmul32_fa28_30_y2(h_u_arrmul32_and28_30_y0, h_u_arrmul32_fa29_29_y2, h_u_arrmul32_fa27_30_y4, h_u_arrmul32_fa28_30_y2, h_u_arrmul32_fa28_30_y4);
  and_gate and_gate_h_u_arrmul32_and29_30_y0(a_29, b_30, h_u_arrmul32_and29_30_y0);
  fa fa_h_u_arrmul32_fa29_30_y2(h_u_arrmul32_and29_30_y0, h_u_arrmul32_fa30_29_y2, h_u_arrmul32_fa28_30_y4, h_u_arrmul32_fa29_30_y2, h_u_arrmul32_fa29_30_y4);
  and_gate and_gate_h_u_arrmul32_and30_30_y0(a_30, b_30, h_u_arrmul32_and30_30_y0);
  fa fa_h_u_arrmul32_fa30_30_y2(h_u_arrmul32_and30_30_y0, h_u_arrmul32_fa31_29_y2, h_u_arrmul32_fa29_30_y4, h_u_arrmul32_fa30_30_y2, h_u_arrmul32_fa30_30_y4);
  and_gate and_gate_h_u_arrmul32_and31_30_y0(a_31, b_30, h_u_arrmul32_and31_30_y0);
  fa fa_h_u_arrmul32_fa31_30_y2(h_u_arrmul32_and31_30_y0, h_u_arrmul32_fa31_29_y4, h_u_arrmul32_fa30_30_y4, h_u_arrmul32_fa31_30_y2, h_u_arrmul32_fa31_30_y4);
  and_gate and_gate_h_u_arrmul32_and0_31_y0(a_0, b_31, h_u_arrmul32_and0_31_y0);
  ha ha_h_u_arrmul32_ha0_31_y0(h_u_arrmul32_and0_31_y0, h_u_arrmul32_fa1_30_y2, h_u_arrmul32_ha0_31_y0, h_u_arrmul32_ha0_31_y1);
  and_gate and_gate_h_u_arrmul32_and1_31_y0(a_1, b_31, h_u_arrmul32_and1_31_y0);
  fa fa_h_u_arrmul32_fa1_31_y2(h_u_arrmul32_and1_31_y0, h_u_arrmul32_fa2_30_y2, h_u_arrmul32_ha0_31_y1, h_u_arrmul32_fa1_31_y2, h_u_arrmul32_fa1_31_y4);
  and_gate and_gate_h_u_arrmul32_and2_31_y0(a_2, b_31, h_u_arrmul32_and2_31_y0);
  fa fa_h_u_arrmul32_fa2_31_y2(h_u_arrmul32_and2_31_y0, h_u_arrmul32_fa3_30_y2, h_u_arrmul32_fa1_31_y4, h_u_arrmul32_fa2_31_y2, h_u_arrmul32_fa2_31_y4);
  and_gate and_gate_h_u_arrmul32_and3_31_y0(a_3, b_31, h_u_arrmul32_and3_31_y0);
  fa fa_h_u_arrmul32_fa3_31_y2(h_u_arrmul32_and3_31_y0, h_u_arrmul32_fa4_30_y2, h_u_arrmul32_fa2_31_y4, h_u_arrmul32_fa3_31_y2, h_u_arrmul32_fa3_31_y4);
  and_gate and_gate_h_u_arrmul32_and4_31_y0(a_4, b_31, h_u_arrmul32_and4_31_y0);
  fa fa_h_u_arrmul32_fa4_31_y2(h_u_arrmul32_and4_31_y0, h_u_arrmul32_fa5_30_y2, h_u_arrmul32_fa3_31_y4, h_u_arrmul32_fa4_31_y2, h_u_arrmul32_fa4_31_y4);
  and_gate and_gate_h_u_arrmul32_and5_31_y0(a_5, b_31, h_u_arrmul32_and5_31_y0);
  fa fa_h_u_arrmul32_fa5_31_y2(h_u_arrmul32_and5_31_y0, h_u_arrmul32_fa6_30_y2, h_u_arrmul32_fa4_31_y4, h_u_arrmul32_fa5_31_y2, h_u_arrmul32_fa5_31_y4);
  and_gate and_gate_h_u_arrmul32_and6_31_y0(a_6, b_31, h_u_arrmul32_and6_31_y0);
  fa fa_h_u_arrmul32_fa6_31_y2(h_u_arrmul32_and6_31_y0, h_u_arrmul32_fa7_30_y2, h_u_arrmul32_fa5_31_y4, h_u_arrmul32_fa6_31_y2, h_u_arrmul32_fa6_31_y4);
  and_gate and_gate_h_u_arrmul32_and7_31_y0(a_7, b_31, h_u_arrmul32_and7_31_y0);
  fa fa_h_u_arrmul32_fa7_31_y2(h_u_arrmul32_and7_31_y0, h_u_arrmul32_fa8_30_y2, h_u_arrmul32_fa6_31_y4, h_u_arrmul32_fa7_31_y2, h_u_arrmul32_fa7_31_y4);
  and_gate and_gate_h_u_arrmul32_and8_31_y0(a_8, b_31, h_u_arrmul32_and8_31_y0);
  fa fa_h_u_arrmul32_fa8_31_y2(h_u_arrmul32_and8_31_y0, h_u_arrmul32_fa9_30_y2, h_u_arrmul32_fa7_31_y4, h_u_arrmul32_fa8_31_y2, h_u_arrmul32_fa8_31_y4);
  and_gate and_gate_h_u_arrmul32_and9_31_y0(a_9, b_31, h_u_arrmul32_and9_31_y0);
  fa fa_h_u_arrmul32_fa9_31_y2(h_u_arrmul32_and9_31_y0, h_u_arrmul32_fa10_30_y2, h_u_arrmul32_fa8_31_y4, h_u_arrmul32_fa9_31_y2, h_u_arrmul32_fa9_31_y4);
  and_gate and_gate_h_u_arrmul32_and10_31_y0(a_10, b_31, h_u_arrmul32_and10_31_y0);
  fa fa_h_u_arrmul32_fa10_31_y2(h_u_arrmul32_and10_31_y0, h_u_arrmul32_fa11_30_y2, h_u_arrmul32_fa9_31_y4, h_u_arrmul32_fa10_31_y2, h_u_arrmul32_fa10_31_y4);
  and_gate and_gate_h_u_arrmul32_and11_31_y0(a_11, b_31, h_u_arrmul32_and11_31_y0);
  fa fa_h_u_arrmul32_fa11_31_y2(h_u_arrmul32_and11_31_y0, h_u_arrmul32_fa12_30_y2, h_u_arrmul32_fa10_31_y4, h_u_arrmul32_fa11_31_y2, h_u_arrmul32_fa11_31_y4);
  and_gate and_gate_h_u_arrmul32_and12_31_y0(a_12, b_31, h_u_arrmul32_and12_31_y0);
  fa fa_h_u_arrmul32_fa12_31_y2(h_u_arrmul32_and12_31_y0, h_u_arrmul32_fa13_30_y2, h_u_arrmul32_fa11_31_y4, h_u_arrmul32_fa12_31_y2, h_u_arrmul32_fa12_31_y4);
  and_gate and_gate_h_u_arrmul32_and13_31_y0(a_13, b_31, h_u_arrmul32_and13_31_y0);
  fa fa_h_u_arrmul32_fa13_31_y2(h_u_arrmul32_and13_31_y0, h_u_arrmul32_fa14_30_y2, h_u_arrmul32_fa12_31_y4, h_u_arrmul32_fa13_31_y2, h_u_arrmul32_fa13_31_y4);
  and_gate and_gate_h_u_arrmul32_and14_31_y0(a_14, b_31, h_u_arrmul32_and14_31_y0);
  fa fa_h_u_arrmul32_fa14_31_y2(h_u_arrmul32_and14_31_y0, h_u_arrmul32_fa15_30_y2, h_u_arrmul32_fa13_31_y4, h_u_arrmul32_fa14_31_y2, h_u_arrmul32_fa14_31_y4);
  and_gate and_gate_h_u_arrmul32_and15_31_y0(a_15, b_31, h_u_arrmul32_and15_31_y0);
  fa fa_h_u_arrmul32_fa15_31_y2(h_u_arrmul32_and15_31_y0, h_u_arrmul32_fa16_30_y2, h_u_arrmul32_fa14_31_y4, h_u_arrmul32_fa15_31_y2, h_u_arrmul32_fa15_31_y4);
  and_gate and_gate_h_u_arrmul32_and16_31_y0(a_16, b_31, h_u_arrmul32_and16_31_y0);
  fa fa_h_u_arrmul32_fa16_31_y2(h_u_arrmul32_and16_31_y0, h_u_arrmul32_fa17_30_y2, h_u_arrmul32_fa15_31_y4, h_u_arrmul32_fa16_31_y2, h_u_arrmul32_fa16_31_y4);
  and_gate and_gate_h_u_arrmul32_and17_31_y0(a_17, b_31, h_u_arrmul32_and17_31_y0);
  fa fa_h_u_arrmul32_fa17_31_y2(h_u_arrmul32_and17_31_y0, h_u_arrmul32_fa18_30_y2, h_u_arrmul32_fa16_31_y4, h_u_arrmul32_fa17_31_y2, h_u_arrmul32_fa17_31_y4);
  and_gate and_gate_h_u_arrmul32_and18_31_y0(a_18, b_31, h_u_arrmul32_and18_31_y0);
  fa fa_h_u_arrmul32_fa18_31_y2(h_u_arrmul32_and18_31_y0, h_u_arrmul32_fa19_30_y2, h_u_arrmul32_fa17_31_y4, h_u_arrmul32_fa18_31_y2, h_u_arrmul32_fa18_31_y4);
  and_gate and_gate_h_u_arrmul32_and19_31_y0(a_19, b_31, h_u_arrmul32_and19_31_y0);
  fa fa_h_u_arrmul32_fa19_31_y2(h_u_arrmul32_and19_31_y0, h_u_arrmul32_fa20_30_y2, h_u_arrmul32_fa18_31_y4, h_u_arrmul32_fa19_31_y2, h_u_arrmul32_fa19_31_y4);
  and_gate and_gate_h_u_arrmul32_and20_31_y0(a_20, b_31, h_u_arrmul32_and20_31_y0);
  fa fa_h_u_arrmul32_fa20_31_y2(h_u_arrmul32_and20_31_y0, h_u_arrmul32_fa21_30_y2, h_u_arrmul32_fa19_31_y4, h_u_arrmul32_fa20_31_y2, h_u_arrmul32_fa20_31_y4);
  and_gate and_gate_h_u_arrmul32_and21_31_y0(a_21, b_31, h_u_arrmul32_and21_31_y0);
  fa fa_h_u_arrmul32_fa21_31_y2(h_u_arrmul32_and21_31_y0, h_u_arrmul32_fa22_30_y2, h_u_arrmul32_fa20_31_y4, h_u_arrmul32_fa21_31_y2, h_u_arrmul32_fa21_31_y4);
  and_gate and_gate_h_u_arrmul32_and22_31_y0(a_22, b_31, h_u_arrmul32_and22_31_y0);
  fa fa_h_u_arrmul32_fa22_31_y2(h_u_arrmul32_and22_31_y0, h_u_arrmul32_fa23_30_y2, h_u_arrmul32_fa21_31_y4, h_u_arrmul32_fa22_31_y2, h_u_arrmul32_fa22_31_y4);
  and_gate and_gate_h_u_arrmul32_and23_31_y0(a_23, b_31, h_u_arrmul32_and23_31_y0);
  fa fa_h_u_arrmul32_fa23_31_y2(h_u_arrmul32_and23_31_y0, h_u_arrmul32_fa24_30_y2, h_u_arrmul32_fa22_31_y4, h_u_arrmul32_fa23_31_y2, h_u_arrmul32_fa23_31_y4);
  and_gate and_gate_h_u_arrmul32_and24_31_y0(a_24, b_31, h_u_arrmul32_and24_31_y0);
  fa fa_h_u_arrmul32_fa24_31_y2(h_u_arrmul32_and24_31_y0, h_u_arrmul32_fa25_30_y2, h_u_arrmul32_fa23_31_y4, h_u_arrmul32_fa24_31_y2, h_u_arrmul32_fa24_31_y4);
  and_gate and_gate_h_u_arrmul32_and25_31_y0(a_25, b_31, h_u_arrmul32_and25_31_y0);
  fa fa_h_u_arrmul32_fa25_31_y2(h_u_arrmul32_and25_31_y0, h_u_arrmul32_fa26_30_y2, h_u_arrmul32_fa24_31_y4, h_u_arrmul32_fa25_31_y2, h_u_arrmul32_fa25_31_y4);
  and_gate and_gate_h_u_arrmul32_and26_31_y0(a_26, b_31, h_u_arrmul32_and26_31_y0);
  fa fa_h_u_arrmul32_fa26_31_y2(h_u_arrmul32_and26_31_y0, h_u_arrmul32_fa27_30_y2, h_u_arrmul32_fa25_31_y4, h_u_arrmul32_fa26_31_y2, h_u_arrmul32_fa26_31_y4);
  and_gate and_gate_h_u_arrmul32_and27_31_y0(a_27, b_31, h_u_arrmul32_and27_31_y0);
  fa fa_h_u_arrmul32_fa27_31_y2(h_u_arrmul32_and27_31_y0, h_u_arrmul32_fa28_30_y2, h_u_arrmul32_fa26_31_y4, h_u_arrmul32_fa27_31_y2, h_u_arrmul32_fa27_31_y4);
  and_gate and_gate_h_u_arrmul32_and28_31_y0(a_28, b_31, h_u_arrmul32_and28_31_y0);
  fa fa_h_u_arrmul32_fa28_31_y2(h_u_arrmul32_and28_31_y0, h_u_arrmul32_fa29_30_y2, h_u_arrmul32_fa27_31_y4, h_u_arrmul32_fa28_31_y2, h_u_arrmul32_fa28_31_y4);
  and_gate and_gate_h_u_arrmul32_and29_31_y0(a_29, b_31, h_u_arrmul32_and29_31_y0);
  fa fa_h_u_arrmul32_fa29_31_y2(h_u_arrmul32_and29_31_y0, h_u_arrmul32_fa30_30_y2, h_u_arrmul32_fa28_31_y4, h_u_arrmul32_fa29_31_y2, h_u_arrmul32_fa29_31_y4);
  and_gate and_gate_h_u_arrmul32_and30_31_y0(a_30, b_31, h_u_arrmul32_and30_31_y0);
  fa fa_h_u_arrmul32_fa30_31_y2(h_u_arrmul32_and30_31_y0, h_u_arrmul32_fa31_30_y2, h_u_arrmul32_fa29_31_y4, h_u_arrmul32_fa30_31_y2, h_u_arrmul32_fa30_31_y4);
  and_gate and_gate_h_u_arrmul32_and31_31_y0(a_31, b_31, h_u_arrmul32_and31_31_y0);
  fa fa_h_u_arrmul32_fa31_31_y2(h_u_arrmul32_and31_31_y0, h_u_arrmul32_fa31_30_y4, h_u_arrmul32_fa30_31_y4, h_u_arrmul32_fa31_31_y2, h_u_arrmul32_fa31_31_y4);

  assign out[0] = h_u_arrmul32_and0_0_y0;
  assign out[1] = h_u_arrmul32_ha0_1_y0;
  assign out[2] = h_u_arrmul32_ha0_2_y0;
  assign out[3] = h_u_arrmul32_ha0_3_y0;
  assign out[4] = h_u_arrmul32_ha0_4_y0;
  assign out[5] = h_u_arrmul32_ha0_5_y0;
  assign out[6] = h_u_arrmul32_ha0_6_y0;
  assign out[7] = h_u_arrmul32_ha0_7_y0;
  assign out[8] = h_u_arrmul32_ha0_8_y0;
  assign out[9] = h_u_arrmul32_ha0_9_y0;
  assign out[10] = h_u_arrmul32_ha0_10_y0;
  assign out[11] = h_u_arrmul32_ha0_11_y0;
  assign out[12] = h_u_arrmul32_ha0_12_y0;
  assign out[13] = h_u_arrmul32_ha0_13_y0;
  assign out[14] = h_u_arrmul32_ha0_14_y0;
  assign out[15] = h_u_arrmul32_ha0_15_y0;
  assign out[16] = h_u_arrmul32_ha0_16_y0;
  assign out[17] = h_u_arrmul32_ha0_17_y0;
  assign out[18] = h_u_arrmul32_ha0_18_y0;
  assign out[19] = h_u_arrmul32_ha0_19_y0;
  assign out[20] = h_u_arrmul32_ha0_20_y0;
  assign out[21] = h_u_arrmul32_ha0_21_y0;
  assign out[22] = h_u_arrmul32_ha0_22_y0;
  assign out[23] = h_u_arrmul32_ha0_23_y0;
  assign out[24] = h_u_arrmul32_ha0_24_y0;
  assign out[25] = h_u_arrmul32_ha0_25_y0;
  assign out[26] = h_u_arrmul32_ha0_26_y0;
  assign out[27] = h_u_arrmul32_ha0_27_y0;
  assign out[28] = h_u_arrmul32_ha0_28_y0;
  assign out[29] = h_u_arrmul32_ha0_29_y0;
  assign out[30] = h_u_arrmul32_ha0_30_y0;
  assign out[31] = h_u_arrmul32_ha0_31_y0;
  assign out[32] = h_u_arrmul32_fa1_31_y2;
  assign out[33] = h_u_arrmul32_fa2_31_y2;
  assign out[34] = h_u_arrmul32_fa3_31_y2;
  assign out[35] = h_u_arrmul32_fa4_31_y2;
  assign out[36] = h_u_arrmul32_fa5_31_y2;
  assign out[37] = h_u_arrmul32_fa6_31_y2;
  assign out[38] = h_u_arrmul32_fa7_31_y2;
  assign out[39] = h_u_arrmul32_fa8_31_y2;
  assign out[40] = h_u_arrmul32_fa9_31_y2;
  assign out[41] = h_u_arrmul32_fa10_31_y2;
  assign out[42] = h_u_arrmul32_fa11_31_y2;
  assign out[43] = h_u_arrmul32_fa12_31_y2;
  assign out[44] = h_u_arrmul32_fa13_31_y2;
  assign out[45] = h_u_arrmul32_fa14_31_y2;
  assign out[46] = h_u_arrmul32_fa15_31_y2;
  assign out[47] = h_u_arrmul32_fa16_31_y2;
  assign out[48] = h_u_arrmul32_fa17_31_y2;
  assign out[49] = h_u_arrmul32_fa18_31_y2;
  assign out[50] = h_u_arrmul32_fa19_31_y2;
  assign out[51] = h_u_arrmul32_fa20_31_y2;
  assign out[52] = h_u_arrmul32_fa21_31_y2;
  assign out[53] = h_u_arrmul32_fa22_31_y2;
  assign out[54] = h_u_arrmul32_fa23_31_y2;
  assign out[55] = h_u_arrmul32_fa24_31_y2;
  assign out[56] = h_u_arrmul32_fa25_31_y2;
  assign out[57] = h_u_arrmul32_fa26_31_y2;
  assign out[58] = h_u_arrmul32_fa27_31_y2;
  assign out[59] = h_u_arrmul32_fa28_31_y2;
  assign out[60] = h_u_arrmul32_fa29_31_y2;
  assign out[61] = h_u_arrmul32_fa30_31_y2;
  assign out[62] = h_u_arrmul32_fa31_31_y2;
  assign out[63] = h_u_arrmul32_fa31_31_y4;
endmodule