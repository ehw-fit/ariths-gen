module s_cska4(input [3:0] a, input [3:0] b, output [4:0] s_cska4_out);
  wire s_cska4_xor0;
  wire s_cska4_ha0_xor0;
  wire s_cska4_ha0_and0;
  wire s_cska4_xor1;
  wire s_cska4_fa0_xor0;
  wire s_cska4_fa0_and0;
  wire s_cska4_fa0_xor1;
  wire s_cska4_fa0_and1;
  wire s_cska4_fa0_or0;
  wire s_cska4_xor2;
  wire s_cska4_fa1_xor0;
  wire s_cska4_fa1_and0;
  wire s_cska4_fa1_xor1;
  wire s_cska4_fa1_and1;
  wire s_cska4_fa1_or0;
  wire s_cska4_xor3;
  wire s_cska4_fa2_xor0;
  wire s_cska4_fa2_and0;
  wire s_cska4_fa2_xor1;
  wire s_cska4_fa2_and1;
  wire s_cska4_fa2_or0;
  wire s_cska4_and_propagate00;
  wire s_cska4_and_propagate01;
  wire s_cska4_and_propagate02;
  wire s_cska4_mux2to10_not0;
  wire s_cska4_mux2to10_and1;
  wire s_cska4_xor4;
  wire s_cska4_xor5;

  assign s_cska4_xor0 = a[0] ^ b[0];
  assign s_cska4_ha0_xor0 = a[0] ^ b[0];
  assign s_cska4_ha0_and0 = a[0] & b[0];
  assign s_cska4_xor1 = a[1] ^ b[1];
  assign s_cska4_fa0_xor0 = a[1] ^ b[1];
  assign s_cska4_fa0_and0 = a[1] & b[1];
  assign s_cska4_fa0_xor1 = s_cska4_fa0_xor0 ^ s_cska4_ha0_and0;
  assign s_cska4_fa0_and1 = s_cska4_fa0_xor0 & s_cska4_ha0_and0;
  assign s_cska4_fa0_or0 = s_cska4_fa0_and0 | s_cska4_fa0_and1;
  assign s_cska4_xor2 = a[2] ^ b[2];
  assign s_cska4_fa1_xor0 = a[2] ^ b[2];
  assign s_cska4_fa1_and0 = a[2] & b[2];
  assign s_cska4_fa1_xor1 = s_cska4_fa1_xor0 ^ s_cska4_fa0_or0;
  assign s_cska4_fa1_and1 = s_cska4_fa1_xor0 & s_cska4_fa0_or0;
  assign s_cska4_fa1_or0 = s_cska4_fa1_and0 | s_cska4_fa1_and1;
  assign s_cska4_xor3 = a[3] ^ b[3];
  assign s_cska4_fa2_xor0 = a[3] ^ b[3];
  assign s_cska4_fa2_and0 = a[3] & b[3];
  assign s_cska4_fa2_xor1 = s_cska4_fa2_xor0 ^ s_cska4_fa1_or0;
  assign s_cska4_fa2_and1 = s_cska4_fa2_xor0 & s_cska4_fa1_or0;
  assign s_cska4_fa2_or0 = s_cska4_fa2_and0 | s_cska4_fa2_and1;
  assign s_cska4_and_propagate00 = s_cska4_xor0 & s_cska4_xor2;
  assign s_cska4_and_propagate01 = s_cska4_xor1 & s_cska4_xor3;
  assign s_cska4_and_propagate02 = s_cska4_and_propagate00 & s_cska4_and_propagate01;
  assign s_cska4_mux2to10_not0 = ~s_cska4_and_propagate02;
  assign s_cska4_mux2to10_and1 = s_cska4_fa2_or0 & s_cska4_mux2to10_not0;
  assign s_cska4_xor4 = a[3] ^ b[3];
  assign s_cska4_xor5 = s_cska4_xor4 ^ s_cska4_mux2to10_and1;

  assign s_cska4_out[0] = s_cska4_ha0_xor0;
  assign s_cska4_out[1] = s_cska4_fa0_xor1;
  assign s_cska4_out[2] = s_cska4_fa1_xor1;
  assign s_cska4_out[3] = s_cska4_fa2_xor1;
  assign s_cska4_out[4] = s_cska4_xor5;
endmodule