module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fs(input [0:0] a, input [0:0] b, input [0:0] bin, output [0:0] fs_xor1, output [0:0] fs_or0);
  wire [0:0] fs_xor0;
  wire [0:0] fs_not0;
  wire [0:0] fs_and0;
  wire [0:0] fs_not1;
  wire [0:0] fs_and1;
  xor_gate xor_gate_fs_xor0(.a(a[0]), .b(b[0]), .out(fs_xor0));
  not_gate not_gate_fs_not0(.a(a[0]), .out(fs_not0));
  and_gate and_gate_fs_and0(.a(fs_not0[0]), .b(b[0]), .out(fs_and0));
  xor_gate xor_gate_fs_xor1(.a(bin[0]), .b(fs_xor0[0]), .out(fs_xor1));
  not_gate not_gate_fs_not1(.a(fs_xor0[0]), .out(fs_not1));
  and_gate and_gate_fs_and1(.a(fs_not1[0]), .b(bin[0]), .out(fs_and1));
  or_gate or_gate_fs_or0(.a(fs_and1[0]), .b(fs_and0[0]), .out(fs_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module h_arrdiv16(input [15:0] a, input [15:0] b, output [15:0] h_arrdiv16_out);
  wire [0:0] h_arrdiv16_fs0_xor0;
  wire [0:0] h_arrdiv16_fs0_and0;
  wire [0:0] h_arrdiv16_fs1_xor1;
  wire [0:0] h_arrdiv16_fs1_or0;
  wire [0:0] h_arrdiv16_fs2_xor1;
  wire [0:0] h_arrdiv16_fs2_or0;
  wire [0:0] h_arrdiv16_fs3_xor1;
  wire [0:0] h_arrdiv16_fs3_or0;
  wire [0:0] h_arrdiv16_fs4_xor1;
  wire [0:0] h_arrdiv16_fs4_or0;
  wire [0:0] h_arrdiv16_fs5_xor1;
  wire [0:0] h_arrdiv16_fs5_or0;
  wire [0:0] h_arrdiv16_fs6_xor1;
  wire [0:0] h_arrdiv16_fs6_or0;
  wire [0:0] h_arrdiv16_fs7_xor1;
  wire [0:0] h_arrdiv16_fs7_or0;
  wire [0:0] h_arrdiv16_fs8_xor1;
  wire [0:0] h_arrdiv16_fs8_or0;
  wire [0:0] h_arrdiv16_fs9_xor1;
  wire [0:0] h_arrdiv16_fs9_or0;
  wire [0:0] h_arrdiv16_fs10_xor1;
  wire [0:0] h_arrdiv16_fs10_or0;
  wire [0:0] h_arrdiv16_fs11_xor1;
  wire [0:0] h_arrdiv16_fs11_or0;
  wire [0:0] h_arrdiv16_fs12_xor1;
  wire [0:0] h_arrdiv16_fs12_or0;
  wire [0:0] h_arrdiv16_fs13_xor1;
  wire [0:0] h_arrdiv16_fs13_or0;
  wire [0:0] h_arrdiv16_fs14_xor1;
  wire [0:0] h_arrdiv16_fs14_or0;
  wire [0:0] h_arrdiv16_fs15_xor1;
  wire [0:0] h_arrdiv16_fs15_or0;
  wire [0:0] h_arrdiv16_mux2to10_xor0;
  wire [0:0] h_arrdiv16_mux2to11_and1;
  wire [0:0] h_arrdiv16_mux2to12_and1;
  wire [0:0] h_arrdiv16_mux2to13_and1;
  wire [0:0] h_arrdiv16_mux2to14_and1;
  wire [0:0] h_arrdiv16_mux2to15_and1;
  wire [0:0] h_arrdiv16_mux2to16_and1;
  wire [0:0] h_arrdiv16_mux2to17_and1;
  wire [0:0] h_arrdiv16_mux2to18_and1;
  wire [0:0] h_arrdiv16_mux2to19_and1;
  wire [0:0] h_arrdiv16_mux2to110_and1;
  wire [0:0] h_arrdiv16_mux2to111_and1;
  wire [0:0] h_arrdiv16_mux2to112_and1;
  wire [0:0] h_arrdiv16_mux2to113_and1;
  wire [0:0] h_arrdiv16_mux2to114_and1;
  wire [0:0] h_arrdiv16_not0;
  wire [0:0] h_arrdiv16_fs16_xor0;
  wire [0:0] h_arrdiv16_fs16_and0;
  wire [0:0] h_arrdiv16_fs17_xor1;
  wire [0:0] h_arrdiv16_fs17_or0;
  wire [0:0] h_arrdiv16_fs18_xor1;
  wire [0:0] h_arrdiv16_fs18_or0;
  wire [0:0] h_arrdiv16_fs19_xor1;
  wire [0:0] h_arrdiv16_fs19_or0;
  wire [0:0] h_arrdiv16_fs20_xor1;
  wire [0:0] h_arrdiv16_fs20_or0;
  wire [0:0] h_arrdiv16_fs21_xor1;
  wire [0:0] h_arrdiv16_fs21_or0;
  wire [0:0] h_arrdiv16_fs22_xor1;
  wire [0:0] h_arrdiv16_fs22_or0;
  wire [0:0] h_arrdiv16_fs23_xor1;
  wire [0:0] h_arrdiv16_fs23_or0;
  wire [0:0] h_arrdiv16_fs24_xor1;
  wire [0:0] h_arrdiv16_fs24_or0;
  wire [0:0] h_arrdiv16_fs25_xor1;
  wire [0:0] h_arrdiv16_fs25_or0;
  wire [0:0] h_arrdiv16_fs26_xor1;
  wire [0:0] h_arrdiv16_fs26_or0;
  wire [0:0] h_arrdiv16_fs27_xor1;
  wire [0:0] h_arrdiv16_fs27_or0;
  wire [0:0] h_arrdiv16_fs28_xor1;
  wire [0:0] h_arrdiv16_fs28_or0;
  wire [0:0] h_arrdiv16_fs29_xor1;
  wire [0:0] h_arrdiv16_fs29_or0;
  wire [0:0] h_arrdiv16_fs30_xor1;
  wire [0:0] h_arrdiv16_fs30_or0;
  wire [0:0] h_arrdiv16_fs31_xor1;
  wire [0:0] h_arrdiv16_fs31_or0;
  wire [0:0] h_arrdiv16_mux2to115_xor0;
  wire [0:0] h_arrdiv16_mux2to116_xor0;
  wire [0:0] h_arrdiv16_mux2to117_xor0;
  wire [0:0] h_arrdiv16_mux2to118_xor0;
  wire [0:0] h_arrdiv16_mux2to119_xor0;
  wire [0:0] h_arrdiv16_mux2to120_xor0;
  wire [0:0] h_arrdiv16_mux2to121_xor0;
  wire [0:0] h_arrdiv16_mux2to122_xor0;
  wire [0:0] h_arrdiv16_mux2to123_xor0;
  wire [0:0] h_arrdiv16_mux2to124_xor0;
  wire [0:0] h_arrdiv16_mux2to125_xor0;
  wire [0:0] h_arrdiv16_mux2to126_xor0;
  wire [0:0] h_arrdiv16_mux2to127_xor0;
  wire [0:0] h_arrdiv16_mux2to128_xor0;
  wire [0:0] h_arrdiv16_mux2to129_xor0;
  wire [0:0] h_arrdiv16_not1;
  wire [0:0] h_arrdiv16_fs32_xor0;
  wire [0:0] h_arrdiv16_fs32_and0;
  wire [0:0] h_arrdiv16_fs33_xor1;
  wire [0:0] h_arrdiv16_fs33_or0;
  wire [0:0] h_arrdiv16_fs34_xor1;
  wire [0:0] h_arrdiv16_fs34_or0;
  wire [0:0] h_arrdiv16_fs35_xor1;
  wire [0:0] h_arrdiv16_fs35_or0;
  wire [0:0] h_arrdiv16_fs36_xor1;
  wire [0:0] h_arrdiv16_fs36_or0;
  wire [0:0] h_arrdiv16_fs37_xor1;
  wire [0:0] h_arrdiv16_fs37_or0;
  wire [0:0] h_arrdiv16_fs38_xor1;
  wire [0:0] h_arrdiv16_fs38_or0;
  wire [0:0] h_arrdiv16_fs39_xor1;
  wire [0:0] h_arrdiv16_fs39_or0;
  wire [0:0] h_arrdiv16_fs40_xor1;
  wire [0:0] h_arrdiv16_fs40_or0;
  wire [0:0] h_arrdiv16_fs41_xor1;
  wire [0:0] h_arrdiv16_fs41_or0;
  wire [0:0] h_arrdiv16_fs42_xor1;
  wire [0:0] h_arrdiv16_fs42_or0;
  wire [0:0] h_arrdiv16_fs43_xor1;
  wire [0:0] h_arrdiv16_fs43_or0;
  wire [0:0] h_arrdiv16_fs44_xor1;
  wire [0:0] h_arrdiv16_fs44_or0;
  wire [0:0] h_arrdiv16_fs45_xor1;
  wire [0:0] h_arrdiv16_fs45_or0;
  wire [0:0] h_arrdiv16_fs46_xor1;
  wire [0:0] h_arrdiv16_fs46_or0;
  wire [0:0] h_arrdiv16_fs47_xor1;
  wire [0:0] h_arrdiv16_fs47_or0;
  wire [0:0] h_arrdiv16_mux2to130_xor0;
  wire [0:0] h_arrdiv16_mux2to131_xor0;
  wire [0:0] h_arrdiv16_mux2to132_xor0;
  wire [0:0] h_arrdiv16_mux2to133_xor0;
  wire [0:0] h_arrdiv16_mux2to134_xor0;
  wire [0:0] h_arrdiv16_mux2to135_xor0;
  wire [0:0] h_arrdiv16_mux2to136_xor0;
  wire [0:0] h_arrdiv16_mux2to137_xor0;
  wire [0:0] h_arrdiv16_mux2to138_xor0;
  wire [0:0] h_arrdiv16_mux2to139_xor0;
  wire [0:0] h_arrdiv16_mux2to140_xor0;
  wire [0:0] h_arrdiv16_mux2to141_xor0;
  wire [0:0] h_arrdiv16_mux2to142_xor0;
  wire [0:0] h_arrdiv16_mux2to143_xor0;
  wire [0:0] h_arrdiv16_mux2to144_xor0;
  wire [0:0] h_arrdiv16_not2;
  wire [0:0] h_arrdiv16_fs48_xor0;
  wire [0:0] h_arrdiv16_fs48_and0;
  wire [0:0] h_arrdiv16_fs49_xor1;
  wire [0:0] h_arrdiv16_fs49_or0;
  wire [0:0] h_arrdiv16_fs50_xor1;
  wire [0:0] h_arrdiv16_fs50_or0;
  wire [0:0] h_arrdiv16_fs51_xor1;
  wire [0:0] h_arrdiv16_fs51_or0;
  wire [0:0] h_arrdiv16_fs52_xor1;
  wire [0:0] h_arrdiv16_fs52_or0;
  wire [0:0] h_arrdiv16_fs53_xor1;
  wire [0:0] h_arrdiv16_fs53_or0;
  wire [0:0] h_arrdiv16_fs54_xor1;
  wire [0:0] h_arrdiv16_fs54_or0;
  wire [0:0] h_arrdiv16_fs55_xor1;
  wire [0:0] h_arrdiv16_fs55_or0;
  wire [0:0] h_arrdiv16_fs56_xor1;
  wire [0:0] h_arrdiv16_fs56_or0;
  wire [0:0] h_arrdiv16_fs57_xor1;
  wire [0:0] h_arrdiv16_fs57_or0;
  wire [0:0] h_arrdiv16_fs58_xor1;
  wire [0:0] h_arrdiv16_fs58_or0;
  wire [0:0] h_arrdiv16_fs59_xor1;
  wire [0:0] h_arrdiv16_fs59_or0;
  wire [0:0] h_arrdiv16_fs60_xor1;
  wire [0:0] h_arrdiv16_fs60_or0;
  wire [0:0] h_arrdiv16_fs61_xor1;
  wire [0:0] h_arrdiv16_fs61_or0;
  wire [0:0] h_arrdiv16_fs62_xor1;
  wire [0:0] h_arrdiv16_fs62_or0;
  wire [0:0] h_arrdiv16_fs63_xor1;
  wire [0:0] h_arrdiv16_fs63_or0;
  wire [0:0] h_arrdiv16_mux2to145_xor0;
  wire [0:0] h_arrdiv16_mux2to146_xor0;
  wire [0:0] h_arrdiv16_mux2to147_xor0;
  wire [0:0] h_arrdiv16_mux2to148_xor0;
  wire [0:0] h_arrdiv16_mux2to149_xor0;
  wire [0:0] h_arrdiv16_mux2to150_xor0;
  wire [0:0] h_arrdiv16_mux2to151_xor0;
  wire [0:0] h_arrdiv16_mux2to152_xor0;
  wire [0:0] h_arrdiv16_mux2to153_xor0;
  wire [0:0] h_arrdiv16_mux2to154_xor0;
  wire [0:0] h_arrdiv16_mux2to155_xor0;
  wire [0:0] h_arrdiv16_mux2to156_xor0;
  wire [0:0] h_arrdiv16_mux2to157_xor0;
  wire [0:0] h_arrdiv16_mux2to158_xor0;
  wire [0:0] h_arrdiv16_mux2to159_xor0;
  wire [0:0] h_arrdiv16_not3;
  wire [0:0] h_arrdiv16_fs64_xor0;
  wire [0:0] h_arrdiv16_fs64_and0;
  wire [0:0] h_arrdiv16_fs65_xor1;
  wire [0:0] h_arrdiv16_fs65_or0;
  wire [0:0] h_arrdiv16_fs66_xor1;
  wire [0:0] h_arrdiv16_fs66_or0;
  wire [0:0] h_arrdiv16_fs67_xor1;
  wire [0:0] h_arrdiv16_fs67_or0;
  wire [0:0] h_arrdiv16_fs68_xor1;
  wire [0:0] h_arrdiv16_fs68_or0;
  wire [0:0] h_arrdiv16_fs69_xor1;
  wire [0:0] h_arrdiv16_fs69_or0;
  wire [0:0] h_arrdiv16_fs70_xor1;
  wire [0:0] h_arrdiv16_fs70_or0;
  wire [0:0] h_arrdiv16_fs71_xor1;
  wire [0:0] h_arrdiv16_fs71_or0;
  wire [0:0] h_arrdiv16_fs72_xor1;
  wire [0:0] h_arrdiv16_fs72_or0;
  wire [0:0] h_arrdiv16_fs73_xor1;
  wire [0:0] h_arrdiv16_fs73_or0;
  wire [0:0] h_arrdiv16_fs74_xor1;
  wire [0:0] h_arrdiv16_fs74_or0;
  wire [0:0] h_arrdiv16_fs75_xor1;
  wire [0:0] h_arrdiv16_fs75_or0;
  wire [0:0] h_arrdiv16_fs76_xor1;
  wire [0:0] h_arrdiv16_fs76_or0;
  wire [0:0] h_arrdiv16_fs77_xor1;
  wire [0:0] h_arrdiv16_fs77_or0;
  wire [0:0] h_arrdiv16_fs78_xor1;
  wire [0:0] h_arrdiv16_fs78_or0;
  wire [0:0] h_arrdiv16_fs79_xor1;
  wire [0:0] h_arrdiv16_fs79_or0;
  wire [0:0] h_arrdiv16_mux2to160_xor0;
  wire [0:0] h_arrdiv16_mux2to161_xor0;
  wire [0:0] h_arrdiv16_mux2to162_xor0;
  wire [0:0] h_arrdiv16_mux2to163_xor0;
  wire [0:0] h_arrdiv16_mux2to164_xor0;
  wire [0:0] h_arrdiv16_mux2to165_xor0;
  wire [0:0] h_arrdiv16_mux2to166_xor0;
  wire [0:0] h_arrdiv16_mux2to167_xor0;
  wire [0:0] h_arrdiv16_mux2to168_xor0;
  wire [0:0] h_arrdiv16_mux2to169_xor0;
  wire [0:0] h_arrdiv16_mux2to170_xor0;
  wire [0:0] h_arrdiv16_mux2to171_xor0;
  wire [0:0] h_arrdiv16_mux2to172_xor0;
  wire [0:0] h_arrdiv16_mux2to173_xor0;
  wire [0:0] h_arrdiv16_mux2to174_xor0;
  wire [0:0] h_arrdiv16_not4;
  wire [0:0] h_arrdiv16_fs80_xor0;
  wire [0:0] h_arrdiv16_fs80_and0;
  wire [0:0] h_arrdiv16_fs81_xor1;
  wire [0:0] h_arrdiv16_fs81_or0;
  wire [0:0] h_arrdiv16_fs82_xor1;
  wire [0:0] h_arrdiv16_fs82_or0;
  wire [0:0] h_arrdiv16_fs83_xor1;
  wire [0:0] h_arrdiv16_fs83_or0;
  wire [0:0] h_arrdiv16_fs84_xor1;
  wire [0:0] h_arrdiv16_fs84_or0;
  wire [0:0] h_arrdiv16_fs85_xor1;
  wire [0:0] h_arrdiv16_fs85_or0;
  wire [0:0] h_arrdiv16_fs86_xor1;
  wire [0:0] h_arrdiv16_fs86_or0;
  wire [0:0] h_arrdiv16_fs87_xor1;
  wire [0:0] h_arrdiv16_fs87_or0;
  wire [0:0] h_arrdiv16_fs88_xor1;
  wire [0:0] h_arrdiv16_fs88_or0;
  wire [0:0] h_arrdiv16_fs89_xor1;
  wire [0:0] h_arrdiv16_fs89_or0;
  wire [0:0] h_arrdiv16_fs90_xor1;
  wire [0:0] h_arrdiv16_fs90_or0;
  wire [0:0] h_arrdiv16_fs91_xor1;
  wire [0:0] h_arrdiv16_fs91_or0;
  wire [0:0] h_arrdiv16_fs92_xor1;
  wire [0:0] h_arrdiv16_fs92_or0;
  wire [0:0] h_arrdiv16_fs93_xor1;
  wire [0:0] h_arrdiv16_fs93_or0;
  wire [0:0] h_arrdiv16_fs94_xor1;
  wire [0:0] h_arrdiv16_fs94_or0;
  wire [0:0] h_arrdiv16_fs95_xor1;
  wire [0:0] h_arrdiv16_fs95_or0;
  wire [0:0] h_arrdiv16_mux2to175_xor0;
  wire [0:0] h_arrdiv16_mux2to176_xor0;
  wire [0:0] h_arrdiv16_mux2to177_xor0;
  wire [0:0] h_arrdiv16_mux2to178_xor0;
  wire [0:0] h_arrdiv16_mux2to179_xor0;
  wire [0:0] h_arrdiv16_mux2to180_xor0;
  wire [0:0] h_arrdiv16_mux2to181_xor0;
  wire [0:0] h_arrdiv16_mux2to182_xor0;
  wire [0:0] h_arrdiv16_mux2to183_xor0;
  wire [0:0] h_arrdiv16_mux2to184_xor0;
  wire [0:0] h_arrdiv16_mux2to185_xor0;
  wire [0:0] h_arrdiv16_mux2to186_xor0;
  wire [0:0] h_arrdiv16_mux2to187_xor0;
  wire [0:0] h_arrdiv16_mux2to188_xor0;
  wire [0:0] h_arrdiv16_mux2to189_xor0;
  wire [0:0] h_arrdiv16_not5;
  wire [0:0] h_arrdiv16_fs96_xor0;
  wire [0:0] h_arrdiv16_fs96_and0;
  wire [0:0] h_arrdiv16_fs97_xor1;
  wire [0:0] h_arrdiv16_fs97_or0;
  wire [0:0] h_arrdiv16_fs98_xor1;
  wire [0:0] h_arrdiv16_fs98_or0;
  wire [0:0] h_arrdiv16_fs99_xor1;
  wire [0:0] h_arrdiv16_fs99_or0;
  wire [0:0] h_arrdiv16_fs100_xor1;
  wire [0:0] h_arrdiv16_fs100_or0;
  wire [0:0] h_arrdiv16_fs101_xor1;
  wire [0:0] h_arrdiv16_fs101_or0;
  wire [0:0] h_arrdiv16_fs102_xor1;
  wire [0:0] h_arrdiv16_fs102_or0;
  wire [0:0] h_arrdiv16_fs103_xor1;
  wire [0:0] h_arrdiv16_fs103_or0;
  wire [0:0] h_arrdiv16_fs104_xor1;
  wire [0:0] h_arrdiv16_fs104_or0;
  wire [0:0] h_arrdiv16_fs105_xor1;
  wire [0:0] h_arrdiv16_fs105_or0;
  wire [0:0] h_arrdiv16_fs106_xor1;
  wire [0:0] h_arrdiv16_fs106_or0;
  wire [0:0] h_arrdiv16_fs107_xor1;
  wire [0:0] h_arrdiv16_fs107_or0;
  wire [0:0] h_arrdiv16_fs108_xor1;
  wire [0:0] h_arrdiv16_fs108_or0;
  wire [0:0] h_arrdiv16_fs109_xor1;
  wire [0:0] h_arrdiv16_fs109_or0;
  wire [0:0] h_arrdiv16_fs110_xor1;
  wire [0:0] h_arrdiv16_fs110_or0;
  wire [0:0] h_arrdiv16_fs111_xor1;
  wire [0:0] h_arrdiv16_fs111_or0;
  wire [0:0] h_arrdiv16_mux2to190_xor0;
  wire [0:0] h_arrdiv16_mux2to191_xor0;
  wire [0:0] h_arrdiv16_mux2to192_xor0;
  wire [0:0] h_arrdiv16_mux2to193_xor0;
  wire [0:0] h_arrdiv16_mux2to194_xor0;
  wire [0:0] h_arrdiv16_mux2to195_xor0;
  wire [0:0] h_arrdiv16_mux2to196_xor0;
  wire [0:0] h_arrdiv16_mux2to197_xor0;
  wire [0:0] h_arrdiv16_mux2to198_xor0;
  wire [0:0] h_arrdiv16_mux2to199_xor0;
  wire [0:0] h_arrdiv16_mux2to1100_xor0;
  wire [0:0] h_arrdiv16_mux2to1101_xor0;
  wire [0:0] h_arrdiv16_mux2to1102_xor0;
  wire [0:0] h_arrdiv16_mux2to1103_xor0;
  wire [0:0] h_arrdiv16_mux2to1104_xor0;
  wire [0:0] h_arrdiv16_not6;
  wire [0:0] h_arrdiv16_fs112_xor0;
  wire [0:0] h_arrdiv16_fs112_and0;
  wire [0:0] h_arrdiv16_fs113_xor1;
  wire [0:0] h_arrdiv16_fs113_or0;
  wire [0:0] h_arrdiv16_fs114_xor1;
  wire [0:0] h_arrdiv16_fs114_or0;
  wire [0:0] h_arrdiv16_fs115_xor1;
  wire [0:0] h_arrdiv16_fs115_or0;
  wire [0:0] h_arrdiv16_fs116_xor1;
  wire [0:0] h_arrdiv16_fs116_or0;
  wire [0:0] h_arrdiv16_fs117_xor1;
  wire [0:0] h_arrdiv16_fs117_or0;
  wire [0:0] h_arrdiv16_fs118_xor1;
  wire [0:0] h_arrdiv16_fs118_or0;
  wire [0:0] h_arrdiv16_fs119_xor1;
  wire [0:0] h_arrdiv16_fs119_or0;
  wire [0:0] h_arrdiv16_fs120_xor1;
  wire [0:0] h_arrdiv16_fs120_or0;
  wire [0:0] h_arrdiv16_fs121_xor1;
  wire [0:0] h_arrdiv16_fs121_or0;
  wire [0:0] h_arrdiv16_fs122_xor1;
  wire [0:0] h_arrdiv16_fs122_or0;
  wire [0:0] h_arrdiv16_fs123_xor1;
  wire [0:0] h_arrdiv16_fs123_or0;
  wire [0:0] h_arrdiv16_fs124_xor1;
  wire [0:0] h_arrdiv16_fs124_or0;
  wire [0:0] h_arrdiv16_fs125_xor1;
  wire [0:0] h_arrdiv16_fs125_or0;
  wire [0:0] h_arrdiv16_fs126_xor1;
  wire [0:0] h_arrdiv16_fs126_or0;
  wire [0:0] h_arrdiv16_fs127_xor1;
  wire [0:0] h_arrdiv16_fs127_or0;
  wire [0:0] h_arrdiv16_mux2to1105_xor0;
  wire [0:0] h_arrdiv16_mux2to1106_xor0;
  wire [0:0] h_arrdiv16_mux2to1107_xor0;
  wire [0:0] h_arrdiv16_mux2to1108_xor0;
  wire [0:0] h_arrdiv16_mux2to1109_xor0;
  wire [0:0] h_arrdiv16_mux2to1110_xor0;
  wire [0:0] h_arrdiv16_mux2to1111_xor0;
  wire [0:0] h_arrdiv16_mux2to1112_xor0;
  wire [0:0] h_arrdiv16_mux2to1113_xor0;
  wire [0:0] h_arrdiv16_mux2to1114_xor0;
  wire [0:0] h_arrdiv16_mux2to1115_xor0;
  wire [0:0] h_arrdiv16_mux2to1116_xor0;
  wire [0:0] h_arrdiv16_mux2to1117_xor0;
  wire [0:0] h_arrdiv16_mux2to1118_xor0;
  wire [0:0] h_arrdiv16_mux2to1119_xor0;
  wire [0:0] h_arrdiv16_not7;
  wire [0:0] h_arrdiv16_fs128_xor0;
  wire [0:0] h_arrdiv16_fs128_and0;
  wire [0:0] h_arrdiv16_fs129_xor1;
  wire [0:0] h_arrdiv16_fs129_or0;
  wire [0:0] h_arrdiv16_fs130_xor1;
  wire [0:0] h_arrdiv16_fs130_or0;
  wire [0:0] h_arrdiv16_fs131_xor1;
  wire [0:0] h_arrdiv16_fs131_or0;
  wire [0:0] h_arrdiv16_fs132_xor1;
  wire [0:0] h_arrdiv16_fs132_or0;
  wire [0:0] h_arrdiv16_fs133_xor1;
  wire [0:0] h_arrdiv16_fs133_or0;
  wire [0:0] h_arrdiv16_fs134_xor1;
  wire [0:0] h_arrdiv16_fs134_or0;
  wire [0:0] h_arrdiv16_fs135_xor1;
  wire [0:0] h_arrdiv16_fs135_or0;
  wire [0:0] h_arrdiv16_fs136_xor1;
  wire [0:0] h_arrdiv16_fs136_or0;
  wire [0:0] h_arrdiv16_fs137_xor1;
  wire [0:0] h_arrdiv16_fs137_or0;
  wire [0:0] h_arrdiv16_fs138_xor1;
  wire [0:0] h_arrdiv16_fs138_or0;
  wire [0:0] h_arrdiv16_fs139_xor1;
  wire [0:0] h_arrdiv16_fs139_or0;
  wire [0:0] h_arrdiv16_fs140_xor1;
  wire [0:0] h_arrdiv16_fs140_or0;
  wire [0:0] h_arrdiv16_fs141_xor1;
  wire [0:0] h_arrdiv16_fs141_or0;
  wire [0:0] h_arrdiv16_fs142_xor1;
  wire [0:0] h_arrdiv16_fs142_or0;
  wire [0:0] h_arrdiv16_fs143_xor1;
  wire [0:0] h_arrdiv16_fs143_or0;
  wire [0:0] h_arrdiv16_mux2to1120_xor0;
  wire [0:0] h_arrdiv16_mux2to1121_xor0;
  wire [0:0] h_arrdiv16_mux2to1122_xor0;
  wire [0:0] h_arrdiv16_mux2to1123_xor0;
  wire [0:0] h_arrdiv16_mux2to1124_xor0;
  wire [0:0] h_arrdiv16_mux2to1125_xor0;
  wire [0:0] h_arrdiv16_mux2to1126_xor0;
  wire [0:0] h_arrdiv16_mux2to1127_xor0;
  wire [0:0] h_arrdiv16_mux2to1128_xor0;
  wire [0:0] h_arrdiv16_mux2to1129_xor0;
  wire [0:0] h_arrdiv16_mux2to1130_xor0;
  wire [0:0] h_arrdiv16_mux2to1131_xor0;
  wire [0:0] h_arrdiv16_mux2to1132_xor0;
  wire [0:0] h_arrdiv16_mux2to1133_xor0;
  wire [0:0] h_arrdiv16_mux2to1134_xor0;
  wire [0:0] h_arrdiv16_not8;
  wire [0:0] h_arrdiv16_fs144_xor0;
  wire [0:0] h_arrdiv16_fs144_and0;
  wire [0:0] h_arrdiv16_fs145_xor1;
  wire [0:0] h_arrdiv16_fs145_or0;
  wire [0:0] h_arrdiv16_fs146_xor1;
  wire [0:0] h_arrdiv16_fs146_or0;
  wire [0:0] h_arrdiv16_fs147_xor1;
  wire [0:0] h_arrdiv16_fs147_or0;
  wire [0:0] h_arrdiv16_fs148_xor1;
  wire [0:0] h_arrdiv16_fs148_or0;
  wire [0:0] h_arrdiv16_fs149_xor1;
  wire [0:0] h_arrdiv16_fs149_or0;
  wire [0:0] h_arrdiv16_fs150_xor1;
  wire [0:0] h_arrdiv16_fs150_or0;
  wire [0:0] h_arrdiv16_fs151_xor1;
  wire [0:0] h_arrdiv16_fs151_or0;
  wire [0:0] h_arrdiv16_fs152_xor1;
  wire [0:0] h_arrdiv16_fs152_or0;
  wire [0:0] h_arrdiv16_fs153_xor1;
  wire [0:0] h_arrdiv16_fs153_or0;
  wire [0:0] h_arrdiv16_fs154_xor1;
  wire [0:0] h_arrdiv16_fs154_or0;
  wire [0:0] h_arrdiv16_fs155_xor1;
  wire [0:0] h_arrdiv16_fs155_or0;
  wire [0:0] h_arrdiv16_fs156_xor1;
  wire [0:0] h_arrdiv16_fs156_or0;
  wire [0:0] h_arrdiv16_fs157_xor1;
  wire [0:0] h_arrdiv16_fs157_or0;
  wire [0:0] h_arrdiv16_fs158_xor1;
  wire [0:0] h_arrdiv16_fs158_or0;
  wire [0:0] h_arrdiv16_fs159_xor1;
  wire [0:0] h_arrdiv16_fs159_or0;
  wire [0:0] h_arrdiv16_mux2to1135_xor0;
  wire [0:0] h_arrdiv16_mux2to1136_xor0;
  wire [0:0] h_arrdiv16_mux2to1137_xor0;
  wire [0:0] h_arrdiv16_mux2to1138_xor0;
  wire [0:0] h_arrdiv16_mux2to1139_xor0;
  wire [0:0] h_arrdiv16_mux2to1140_xor0;
  wire [0:0] h_arrdiv16_mux2to1141_xor0;
  wire [0:0] h_arrdiv16_mux2to1142_xor0;
  wire [0:0] h_arrdiv16_mux2to1143_xor0;
  wire [0:0] h_arrdiv16_mux2to1144_xor0;
  wire [0:0] h_arrdiv16_mux2to1145_xor0;
  wire [0:0] h_arrdiv16_mux2to1146_xor0;
  wire [0:0] h_arrdiv16_mux2to1147_xor0;
  wire [0:0] h_arrdiv16_mux2to1148_xor0;
  wire [0:0] h_arrdiv16_mux2to1149_xor0;
  wire [0:0] h_arrdiv16_not9;
  wire [0:0] h_arrdiv16_fs160_xor0;
  wire [0:0] h_arrdiv16_fs160_and0;
  wire [0:0] h_arrdiv16_fs161_xor1;
  wire [0:0] h_arrdiv16_fs161_or0;
  wire [0:0] h_arrdiv16_fs162_xor1;
  wire [0:0] h_arrdiv16_fs162_or0;
  wire [0:0] h_arrdiv16_fs163_xor1;
  wire [0:0] h_arrdiv16_fs163_or0;
  wire [0:0] h_arrdiv16_fs164_xor1;
  wire [0:0] h_arrdiv16_fs164_or0;
  wire [0:0] h_arrdiv16_fs165_xor1;
  wire [0:0] h_arrdiv16_fs165_or0;
  wire [0:0] h_arrdiv16_fs166_xor1;
  wire [0:0] h_arrdiv16_fs166_or0;
  wire [0:0] h_arrdiv16_fs167_xor1;
  wire [0:0] h_arrdiv16_fs167_or0;
  wire [0:0] h_arrdiv16_fs168_xor1;
  wire [0:0] h_arrdiv16_fs168_or0;
  wire [0:0] h_arrdiv16_fs169_xor1;
  wire [0:0] h_arrdiv16_fs169_or0;
  wire [0:0] h_arrdiv16_fs170_xor1;
  wire [0:0] h_arrdiv16_fs170_or0;
  wire [0:0] h_arrdiv16_fs171_xor1;
  wire [0:0] h_arrdiv16_fs171_or0;
  wire [0:0] h_arrdiv16_fs172_xor1;
  wire [0:0] h_arrdiv16_fs172_or0;
  wire [0:0] h_arrdiv16_fs173_xor1;
  wire [0:0] h_arrdiv16_fs173_or0;
  wire [0:0] h_arrdiv16_fs174_xor1;
  wire [0:0] h_arrdiv16_fs174_or0;
  wire [0:0] h_arrdiv16_fs175_xor1;
  wire [0:0] h_arrdiv16_fs175_or0;
  wire [0:0] h_arrdiv16_mux2to1150_xor0;
  wire [0:0] h_arrdiv16_mux2to1151_xor0;
  wire [0:0] h_arrdiv16_mux2to1152_xor0;
  wire [0:0] h_arrdiv16_mux2to1153_xor0;
  wire [0:0] h_arrdiv16_mux2to1154_xor0;
  wire [0:0] h_arrdiv16_mux2to1155_xor0;
  wire [0:0] h_arrdiv16_mux2to1156_xor0;
  wire [0:0] h_arrdiv16_mux2to1157_xor0;
  wire [0:0] h_arrdiv16_mux2to1158_xor0;
  wire [0:0] h_arrdiv16_mux2to1159_xor0;
  wire [0:0] h_arrdiv16_mux2to1160_xor0;
  wire [0:0] h_arrdiv16_mux2to1161_xor0;
  wire [0:0] h_arrdiv16_mux2to1162_xor0;
  wire [0:0] h_arrdiv16_mux2to1163_xor0;
  wire [0:0] h_arrdiv16_mux2to1164_xor0;
  wire [0:0] h_arrdiv16_not10;
  wire [0:0] h_arrdiv16_fs176_xor0;
  wire [0:0] h_arrdiv16_fs176_and0;
  wire [0:0] h_arrdiv16_fs177_xor1;
  wire [0:0] h_arrdiv16_fs177_or0;
  wire [0:0] h_arrdiv16_fs178_xor1;
  wire [0:0] h_arrdiv16_fs178_or0;
  wire [0:0] h_arrdiv16_fs179_xor1;
  wire [0:0] h_arrdiv16_fs179_or0;
  wire [0:0] h_arrdiv16_fs180_xor1;
  wire [0:0] h_arrdiv16_fs180_or0;
  wire [0:0] h_arrdiv16_fs181_xor1;
  wire [0:0] h_arrdiv16_fs181_or0;
  wire [0:0] h_arrdiv16_fs182_xor1;
  wire [0:0] h_arrdiv16_fs182_or0;
  wire [0:0] h_arrdiv16_fs183_xor1;
  wire [0:0] h_arrdiv16_fs183_or0;
  wire [0:0] h_arrdiv16_fs184_xor1;
  wire [0:0] h_arrdiv16_fs184_or0;
  wire [0:0] h_arrdiv16_fs185_xor1;
  wire [0:0] h_arrdiv16_fs185_or0;
  wire [0:0] h_arrdiv16_fs186_xor1;
  wire [0:0] h_arrdiv16_fs186_or0;
  wire [0:0] h_arrdiv16_fs187_xor1;
  wire [0:0] h_arrdiv16_fs187_or0;
  wire [0:0] h_arrdiv16_fs188_xor1;
  wire [0:0] h_arrdiv16_fs188_or0;
  wire [0:0] h_arrdiv16_fs189_xor1;
  wire [0:0] h_arrdiv16_fs189_or0;
  wire [0:0] h_arrdiv16_fs190_xor1;
  wire [0:0] h_arrdiv16_fs190_or0;
  wire [0:0] h_arrdiv16_fs191_xor1;
  wire [0:0] h_arrdiv16_fs191_or0;
  wire [0:0] h_arrdiv16_mux2to1165_xor0;
  wire [0:0] h_arrdiv16_mux2to1166_xor0;
  wire [0:0] h_arrdiv16_mux2to1167_xor0;
  wire [0:0] h_arrdiv16_mux2to1168_xor0;
  wire [0:0] h_arrdiv16_mux2to1169_xor0;
  wire [0:0] h_arrdiv16_mux2to1170_xor0;
  wire [0:0] h_arrdiv16_mux2to1171_xor0;
  wire [0:0] h_arrdiv16_mux2to1172_xor0;
  wire [0:0] h_arrdiv16_mux2to1173_xor0;
  wire [0:0] h_arrdiv16_mux2to1174_xor0;
  wire [0:0] h_arrdiv16_mux2to1175_xor0;
  wire [0:0] h_arrdiv16_mux2to1176_xor0;
  wire [0:0] h_arrdiv16_mux2to1177_xor0;
  wire [0:0] h_arrdiv16_mux2to1178_xor0;
  wire [0:0] h_arrdiv16_mux2to1179_xor0;
  wire [0:0] h_arrdiv16_not11;
  wire [0:0] h_arrdiv16_fs192_xor0;
  wire [0:0] h_arrdiv16_fs192_and0;
  wire [0:0] h_arrdiv16_fs193_xor1;
  wire [0:0] h_arrdiv16_fs193_or0;
  wire [0:0] h_arrdiv16_fs194_xor1;
  wire [0:0] h_arrdiv16_fs194_or0;
  wire [0:0] h_arrdiv16_fs195_xor1;
  wire [0:0] h_arrdiv16_fs195_or0;
  wire [0:0] h_arrdiv16_fs196_xor1;
  wire [0:0] h_arrdiv16_fs196_or0;
  wire [0:0] h_arrdiv16_fs197_xor1;
  wire [0:0] h_arrdiv16_fs197_or0;
  wire [0:0] h_arrdiv16_fs198_xor1;
  wire [0:0] h_arrdiv16_fs198_or0;
  wire [0:0] h_arrdiv16_fs199_xor1;
  wire [0:0] h_arrdiv16_fs199_or0;
  wire [0:0] h_arrdiv16_fs200_xor1;
  wire [0:0] h_arrdiv16_fs200_or0;
  wire [0:0] h_arrdiv16_fs201_xor1;
  wire [0:0] h_arrdiv16_fs201_or0;
  wire [0:0] h_arrdiv16_fs202_xor1;
  wire [0:0] h_arrdiv16_fs202_or0;
  wire [0:0] h_arrdiv16_fs203_xor1;
  wire [0:0] h_arrdiv16_fs203_or0;
  wire [0:0] h_arrdiv16_fs204_xor1;
  wire [0:0] h_arrdiv16_fs204_or0;
  wire [0:0] h_arrdiv16_fs205_xor1;
  wire [0:0] h_arrdiv16_fs205_or0;
  wire [0:0] h_arrdiv16_fs206_xor1;
  wire [0:0] h_arrdiv16_fs206_or0;
  wire [0:0] h_arrdiv16_fs207_xor1;
  wire [0:0] h_arrdiv16_fs207_or0;
  wire [0:0] h_arrdiv16_mux2to1180_xor0;
  wire [0:0] h_arrdiv16_mux2to1181_xor0;
  wire [0:0] h_arrdiv16_mux2to1182_xor0;
  wire [0:0] h_arrdiv16_mux2to1183_xor0;
  wire [0:0] h_arrdiv16_mux2to1184_xor0;
  wire [0:0] h_arrdiv16_mux2to1185_xor0;
  wire [0:0] h_arrdiv16_mux2to1186_xor0;
  wire [0:0] h_arrdiv16_mux2to1187_xor0;
  wire [0:0] h_arrdiv16_mux2to1188_xor0;
  wire [0:0] h_arrdiv16_mux2to1189_xor0;
  wire [0:0] h_arrdiv16_mux2to1190_xor0;
  wire [0:0] h_arrdiv16_mux2to1191_xor0;
  wire [0:0] h_arrdiv16_mux2to1192_xor0;
  wire [0:0] h_arrdiv16_mux2to1193_xor0;
  wire [0:0] h_arrdiv16_mux2to1194_xor0;
  wire [0:0] h_arrdiv16_not12;
  wire [0:0] h_arrdiv16_fs208_xor0;
  wire [0:0] h_arrdiv16_fs208_and0;
  wire [0:0] h_arrdiv16_fs209_xor1;
  wire [0:0] h_arrdiv16_fs209_or0;
  wire [0:0] h_arrdiv16_fs210_xor1;
  wire [0:0] h_arrdiv16_fs210_or0;
  wire [0:0] h_arrdiv16_fs211_xor1;
  wire [0:0] h_arrdiv16_fs211_or0;
  wire [0:0] h_arrdiv16_fs212_xor1;
  wire [0:0] h_arrdiv16_fs212_or0;
  wire [0:0] h_arrdiv16_fs213_xor1;
  wire [0:0] h_arrdiv16_fs213_or0;
  wire [0:0] h_arrdiv16_fs214_xor1;
  wire [0:0] h_arrdiv16_fs214_or0;
  wire [0:0] h_arrdiv16_fs215_xor1;
  wire [0:0] h_arrdiv16_fs215_or0;
  wire [0:0] h_arrdiv16_fs216_xor1;
  wire [0:0] h_arrdiv16_fs216_or0;
  wire [0:0] h_arrdiv16_fs217_xor1;
  wire [0:0] h_arrdiv16_fs217_or0;
  wire [0:0] h_arrdiv16_fs218_xor1;
  wire [0:0] h_arrdiv16_fs218_or0;
  wire [0:0] h_arrdiv16_fs219_xor1;
  wire [0:0] h_arrdiv16_fs219_or0;
  wire [0:0] h_arrdiv16_fs220_xor1;
  wire [0:0] h_arrdiv16_fs220_or0;
  wire [0:0] h_arrdiv16_fs221_xor1;
  wire [0:0] h_arrdiv16_fs221_or0;
  wire [0:0] h_arrdiv16_fs222_xor1;
  wire [0:0] h_arrdiv16_fs222_or0;
  wire [0:0] h_arrdiv16_fs223_xor1;
  wire [0:0] h_arrdiv16_fs223_or0;
  wire [0:0] h_arrdiv16_mux2to1195_xor0;
  wire [0:0] h_arrdiv16_mux2to1196_xor0;
  wire [0:0] h_arrdiv16_mux2to1197_xor0;
  wire [0:0] h_arrdiv16_mux2to1198_xor0;
  wire [0:0] h_arrdiv16_mux2to1199_xor0;
  wire [0:0] h_arrdiv16_mux2to1200_xor0;
  wire [0:0] h_arrdiv16_mux2to1201_xor0;
  wire [0:0] h_arrdiv16_mux2to1202_xor0;
  wire [0:0] h_arrdiv16_mux2to1203_xor0;
  wire [0:0] h_arrdiv16_mux2to1204_xor0;
  wire [0:0] h_arrdiv16_mux2to1205_xor0;
  wire [0:0] h_arrdiv16_mux2to1206_xor0;
  wire [0:0] h_arrdiv16_mux2to1207_xor0;
  wire [0:0] h_arrdiv16_mux2to1208_xor0;
  wire [0:0] h_arrdiv16_mux2to1209_xor0;
  wire [0:0] h_arrdiv16_not13;
  wire [0:0] h_arrdiv16_fs224_xor0;
  wire [0:0] h_arrdiv16_fs224_and0;
  wire [0:0] h_arrdiv16_fs225_xor1;
  wire [0:0] h_arrdiv16_fs225_or0;
  wire [0:0] h_arrdiv16_fs226_xor1;
  wire [0:0] h_arrdiv16_fs226_or0;
  wire [0:0] h_arrdiv16_fs227_xor1;
  wire [0:0] h_arrdiv16_fs227_or0;
  wire [0:0] h_arrdiv16_fs228_xor1;
  wire [0:0] h_arrdiv16_fs228_or0;
  wire [0:0] h_arrdiv16_fs229_xor1;
  wire [0:0] h_arrdiv16_fs229_or0;
  wire [0:0] h_arrdiv16_fs230_xor1;
  wire [0:0] h_arrdiv16_fs230_or0;
  wire [0:0] h_arrdiv16_fs231_xor1;
  wire [0:0] h_arrdiv16_fs231_or0;
  wire [0:0] h_arrdiv16_fs232_xor1;
  wire [0:0] h_arrdiv16_fs232_or0;
  wire [0:0] h_arrdiv16_fs233_xor1;
  wire [0:0] h_arrdiv16_fs233_or0;
  wire [0:0] h_arrdiv16_fs234_xor1;
  wire [0:0] h_arrdiv16_fs234_or0;
  wire [0:0] h_arrdiv16_fs235_xor1;
  wire [0:0] h_arrdiv16_fs235_or0;
  wire [0:0] h_arrdiv16_fs236_xor1;
  wire [0:0] h_arrdiv16_fs236_or0;
  wire [0:0] h_arrdiv16_fs237_xor1;
  wire [0:0] h_arrdiv16_fs237_or0;
  wire [0:0] h_arrdiv16_fs238_xor1;
  wire [0:0] h_arrdiv16_fs238_or0;
  wire [0:0] h_arrdiv16_fs239_xor1;
  wire [0:0] h_arrdiv16_fs239_or0;
  wire [0:0] h_arrdiv16_mux2to1210_xor0;
  wire [0:0] h_arrdiv16_mux2to1211_xor0;
  wire [0:0] h_arrdiv16_mux2to1212_xor0;
  wire [0:0] h_arrdiv16_mux2to1213_xor0;
  wire [0:0] h_arrdiv16_mux2to1214_xor0;
  wire [0:0] h_arrdiv16_mux2to1215_xor0;
  wire [0:0] h_arrdiv16_mux2to1216_xor0;
  wire [0:0] h_arrdiv16_mux2to1217_xor0;
  wire [0:0] h_arrdiv16_mux2to1218_xor0;
  wire [0:0] h_arrdiv16_mux2to1219_xor0;
  wire [0:0] h_arrdiv16_mux2to1220_xor0;
  wire [0:0] h_arrdiv16_mux2to1221_xor0;
  wire [0:0] h_arrdiv16_mux2to1222_xor0;
  wire [0:0] h_arrdiv16_mux2to1223_xor0;
  wire [0:0] h_arrdiv16_mux2to1224_xor0;
  wire [0:0] h_arrdiv16_not14;
  wire [0:0] h_arrdiv16_fs240_xor0;
  wire [0:0] h_arrdiv16_fs240_and0;
  wire [0:0] h_arrdiv16_fs241_xor1;
  wire [0:0] h_arrdiv16_fs241_or0;
  wire [0:0] h_arrdiv16_fs242_xor1;
  wire [0:0] h_arrdiv16_fs242_or0;
  wire [0:0] h_arrdiv16_fs243_xor1;
  wire [0:0] h_arrdiv16_fs243_or0;
  wire [0:0] h_arrdiv16_fs244_xor1;
  wire [0:0] h_arrdiv16_fs244_or0;
  wire [0:0] h_arrdiv16_fs245_xor1;
  wire [0:0] h_arrdiv16_fs245_or0;
  wire [0:0] h_arrdiv16_fs246_xor1;
  wire [0:0] h_arrdiv16_fs246_or0;
  wire [0:0] h_arrdiv16_fs247_xor1;
  wire [0:0] h_arrdiv16_fs247_or0;
  wire [0:0] h_arrdiv16_fs248_xor1;
  wire [0:0] h_arrdiv16_fs248_or0;
  wire [0:0] h_arrdiv16_fs249_xor1;
  wire [0:0] h_arrdiv16_fs249_or0;
  wire [0:0] h_arrdiv16_fs250_xor1;
  wire [0:0] h_arrdiv16_fs250_or0;
  wire [0:0] h_arrdiv16_fs251_xor1;
  wire [0:0] h_arrdiv16_fs251_or0;
  wire [0:0] h_arrdiv16_fs252_xor1;
  wire [0:0] h_arrdiv16_fs252_or0;
  wire [0:0] h_arrdiv16_fs253_xor1;
  wire [0:0] h_arrdiv16_fs253_or0;
  wire [0:0] h_arrdiv16_fs254_xor1;
  wire [0:0] h_arrdiv16_fs254_or0;
  wire [0:0] h_arrdiv16_fs255_xor1;
  wire [0:0] h_arrdiv16_fs255_or0;
  wire [0:0] h_arrdiv16_not15;

  fs fs_h_arrdiv16_fs0_out(.a(a[15]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs0_xor0), .fs_or0(h_arrdiv16_fs0_and0));
  fs fs_h_arrdiv16_fs1_out(.a(1'b0), .b(b[1]), .bin(h_arrdiv16_fs0_and0[0]), .fs_xor1(h_arrdiv16_fs1_xor1), .fs_or0(h_arrdiv16_fs1_or0));
  fs fs_h_arrdiv16_fs2_out(.a(1'b0), .b(b[2]), .bin(h_arrdiv16_fs1_or0[0]), .fs_xor1(h_arrdiv16_fs2_xor1), .fs_or0(h_arrdiv16_fs2_or0));
  fs fs_h_arrdiv16_fs3_out(.a(1'b0), .b(b[3]), .bin(h_arrdiv16_fs2_or0[0]), .fs_xor1(h_arrdiv16_fs3_xor1), .fs_or0(h_arrdiv16_fs3_or0));
  fs fs_h_arrdiv16_fs4_out(.a(1'b0), .b(b[4]), .bin(h_arrdiv16_fs3_or0[0]), .fs_xor1(h_arrdiv16_fs4_xor1), .fs_or0(h_arrdiv16_fs4_or0));
  fs fs_h_arrdiv16_fs5_out(.a(1'b0), .b(b[5]), .bin(h_arrdiv16_fs4_or0[0]), .fs_xor1(h_arrdiv16_fs5_xor1), .fs_or0(h_arrdiv16_fs5_or0));
  fs fs_h_arrdiv16_fs6_out(.a(1'b0), .b(b[6]), .bin(h_arrdiv16_fs5_or0[0]), .fs_xor1(h_arrdiv16_fs6_xor1), .fs_or0(h_arrdiv16_fs6_or0));
  fs fs_h_arrdiv16_fs7_out(.a(1'b0), .b(b[7]), .bin(h_arrdiv16_fs6_or0[0]), .fs_xor1(h_arrdiv16_fs7_xor1), .fs_or0(h_arrdiv16_fs7_or0));
  fs fs_h_arrdiv16_fs8_out(.a(1'b0), .b(b[8]), .bin(h_arrdiv16_fs7_or0[0]), .fs_xor1(h_arrdiv16_fs8_xor1), .fs_or0(h_arrdiv16_fs8_or0));
  fs fs_h_arrdiv16_fs9_out(.a(1'b0), .b(b[9]), .bin(h_arrdiv16_fs8_or0[0]), .fs_xor1(h_arrdiv16_fs9_xor1), .fs_or0(h_arrdiv16_fs9_or0));
  fs fs_h_arrdiv16_fs10_out(.a(1'b0), .b(b[10]), .bin(h_arrdiv16_fs9_or0[0]), .fs_xor1(h_arrdiv16_fs10_xor1), .fs_or0(h_arrdiv16_fs10_or0));
  fs fs_h_arrdiv16_fs11_out(.a(1'b0), .b(b[11]), .bin(h_arrdiv16_fs10_or0[0]), .fs_xor1(h_arrdiv16_fs11_xor1), .fs_or0(h_arrdiv16_fs11_or0));
  fs fs_h_arrdiv16_fs12_out(.a(1'b0), .b(b[12]), .bin(h_arrdiv16_fs11_or0[0]), .fs_xor1(h_arrdiv16_fs12_xor1), .fs_or0(h_arrdiv16_fs12_or0));
  fs fs_h_arrdiv16_fs13_out(.a(1'b0), .b(b[13]), .bin(h_arrdiv16_fs12_or0[0]), .fs_xor1(h_arrdiv16_fs13_xor1), .fs_or0(h_arrdiv16_fs13_or0));
  fs fs_h_arrdiv16_fs14_out(.a(1'b0), .b(b[14]), .bin(h_arrdiv16_fs13_or0[0]), .fs_xor1(h_arrdiv16_fs14_xor1), .fs_or0(h_arrdiv16_fs14_or0));
  fs fs_h_arrdiv16_fs15_out(.a(1'b0), .b(b[15]), .bin(h_arrdiv16_fs14_or0[0]), .fs_xor1(h_arrdiv16_fs15_xor1), .fs_or0(h_arrdiv16_fs15_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to10_out(.d0(h_arrdiv16_fs0_xor0[0]), .d1(a[15]), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to10_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to11_out(.d0(h_arrdiv16_fs1_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to11_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to12_out(.d0(h_arrdiv16_fs2_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to12_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to13_out(.d0(h_arrdiv16_fs3_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to13_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to14_out(.d0(h_arrdiv16_fs4_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to14_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to15_out(.d0(h_arrdiv16_fs5_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to15_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to16_out(.d0(h_arrdiv16_fs6_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to16_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to17_out(.d0(h_arrdiv16_fs7_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to17_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to18_out(.d0(h_arrdiv16_fs8_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to18_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to19_out(.d0(h_arrdiv16_fs9_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to19_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to110_out(.d0(h_arrdiv16_fs10_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to110_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to111_out(.d0(h_arrdiv16_fs11_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to111_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to112_out(.d0(h_arrdiv16_fs12_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to112_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to113_out(.d0(h_arrdiv16_fs13_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to113_and1));
  mux2to1 mux2to1_h_arrdiv16_mux2to114_out(.d0(h_arrdiv16_fs14_xor1[0]), .d1(1'b0), .sel(h_arrdiv16_fs15_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to114_and1));
  not_gate not_gate_h_arrdiv16_not0(.a(h_arrdiv16_fs15_or0[0]), .out(h_arrdiv16_not0));
  fs fs_h_arrdiv16_fs16_out(.a(a[14]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs16_xor0), .fs_or0(h_arrdiv16_fs16_and0));
  fs fs_h_arrdiv16_fs17_out(.a(h_arrdiv16_mux2to10_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs16_and0[0]), .fs_xor1(h_arrdiv16_fs17_xor1), .fs_or0(h_arrdiv16_fs17_or0));
  fs fs_h_arrdiv16_fs18_out(.a(h_arrdiv16_mux2to11_and1[0]), .b(b[2]), .bin(h_arrdiv16_fs17_or0[0]), .fs_xor1(h_arrdiv16_fs18_xor1), .fs_or0(h_arrdiv16_fs18_or0));
  fs fs_h_arrdiv16_fs19_out(.a(h_arrdiv16_mux2to12_and1[0]), .b(b[3]), .bin(h_arrdiv16_fs18_or0[0]), .fs_xor1(h_arrdiv16_fs19_xor1), .fs_or0(h_arrdiv16_fs19_or0));
  fs fs_h_arrdiv16_fs20_out(.a(h_arrdiv16_mux2to13_and1[0]), .b(b[4]), .bin(h_arrdiv16_fs19_or0[0]), .fs_xor1(h_arrdiv16_fs20_xor1), .fs_or0(h_arrdiv16_fs20_or0));
  fs fs_h_arrdiv16_fs21_out(.a(h_arrdiv16_mux2to14_and1[0]), .b(b[5]), .bin(h_arrdiv16_fs20_or0[0]), .fs_xor1(h_arrdiv16_fs21_xor1), .fs_or0(h_arrdiv16_fs21_or0));
  fs fs_h_arrdiv16_fs22_out(.a(h_arrdiv16_mux2to15_and1[0]), .b(b[6]), .bin(h_arrdiv16_fs21_or0[0]), .fs_xor1(h_arrdiv16_fs22_xor1), .fs_or0(h_arrdiv16_fs22_or0));
  fs fs_h_arrdiv16_fs23_out(.a(h_arrdiv16_mux2to16_and1[0]), .b(b[7]), .bin(h_arrdiv16_fs22_or0[0]), .fs_xor1(h_arrdiv16_fs23_xor1), .fs_or0(h_arrdiv16_fs23_or0));
  fs fs_h_arrdiv16_fs24_out(.a(h_arrdiv16_mux2to17_and1[0]), .b(b[8]), .bin(h_arrdiv16_fs23_or0[0]), .fs_xor1(h_arrdiv16_fs24_xor1), .fs_or0(h_arrdiv16_fs24_or0));
  fs fs_h_arrdiv16_fs25_out(.a(h_arrdiv16_mux2to18_and1[0]), .b(b[9]), .bin(h_arrdiv16_fs24_or0[0]), .fs_xor1(h_arrdiv16_fs25_xor1), .fs_or0(h_arrdiv16_fs25_or0));
  fs fs_h_arrdiv16_fs26_out(.a(h_arrdiv16_mux2to19_and1[0]), .b(b[10]), .bin(h_arrdiv16_fs25_or0[0]), .fs_xor1(h_arrdiv16_fs26_xor1), .fs_or0(h_arrdiv16_fs26_or0));
  fs fs_h_arrdiv16_fs27_out(.a(h_arrdiv16_mux2to110_and1[0]), .b(b[11]), .bin(h_arrdiv16_fs26_or0[0]), .fs_xor1(h_arrdiv16_fs27_xor1), .fs_or0(h_arrdiv16_fs27_or0));
  fs fs_h_arrdiv16_fs28_out(.a(h_arrdiv16_mux2to111_and1[0]), .b(b[12]), .bin(h_arrdiv16_fs27_or0[0]), .fs_xor1(h_arrdiv16_fs28_xor1), .fs_or0(h_arrdiv16_fs28_or0));
  fs fs_h_arrdiv16_fs29_out(.a(h_arrdiv16_mux2to112_and1[0]), .b(b[13]), .bin(h_arrdiv16_fs28_or0[0]), .fs_xor1(h_arrdiv16_fs29_xor1), .fs_or0(h_arrdiv16_fs29_or0));
  fs fs_h_arrdiv16_fs30_out(.a(h_arrdiv16_mux2to113_and1[0]), .b(b[14]), .bin(h_arrdiv16_fs29_or0[0]), .fs_xor1(h_arrdiv16_fs30_xor1), .fs_or0(h_arrdiv16_fs30_or0));
  fs fs_h_arrdiv16_fs31_out(.a(h_arrdiv16_mux2to114_and1[0]), .b(b[15]), .bin(h_arrdiv16_fs30_or0[0]), .fs_xor1(h_arrdiv16_fs31_xor1), .fs_or0(h_arrdiv16_fs31_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to115_out(.d0(h_arrdiv16_fs16_xor0[0]), .d1(a[14]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to115_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to116_out(.d0(h_arrdiv16_fs17_xor1[0]), .d1(h_arrdiv16_mux2to10_xor0[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to116_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to117_out(.d0(h_arrdiv16_fs18_xor1[0]), .d1(h_arrdiv16_mux2to11_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to117_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to118_out(.d0(h_arrdiv16_fs19_xor1[0]), .d1(h_arrdiv16_mux2to12_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to118_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to119_out(.d0(h_arrdiv16_fs20_xor1[0]), .d1(h_arrdiv16_mux2to13_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to119_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to120_out(.d0(h_arrdiv16_fs21_xor1[0]), .d1(h_arrdiv16_mux2to14_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to120_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to121_out(.d0(h_arrdiv16_fs22_xor1[0]), .d1(h_arrdiv16_mux2to15_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to121_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to122_out(.d0(h_arrdiv16_fs23_xor1[0]), .d1(h_arrdiv16_mux2to16_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to122_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to123_out(.d0(h_arrdiv16_fs24_xor1[0]), .d1(h_arrdiv16_mux2to17_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to123_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to124_out(.d0(h_arrdiv16_fs25_xor1[0]), .d1(h_arrdiv16_mux2to18_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to124_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to125_out(.d0(h_arrdiv16_fs26_xor1[0]), .d1(h_arrdiv16_mux2to19_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to125_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to126_out(.d0(h_arrdiv16_fs27_xor1[0]), .d1(h_arrdiv16_mux2to110_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to126_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to127_out(.d0(h_arrdiv16_fs28_xor1[0]), .d1(h_arrdiv16_mux2to111_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to127_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to128_out(.d0(h_arrdiv16_fs29_xor1[0]), .d1(h_arrdiv16_mux2to112_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to128_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to129_out(.d0(h_arrdiv16_fs30_xor1[0]), .d1(h_arrdiv16_mux2to113_and1[0]), .sel(h_arrdiv16_fs31_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to129_xor0));
  not_gate not_gate_h_arrdiv16_not1(.a(h_arrdiv16_fs31_or0[0]), .out(h_arrdiv16_not1));
  fs fs_h_arrdiv16_fs32_out(.a(a[13]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs32_xor0), .fs_or0(h_arrdiv16_fs32_and0));
  fs fs_h_arrdiv16_fs33_out(.a(h_arrdiv16_mux2to115_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs32_and0[0]), .fs_xor1(h_arrdiv16_fs33_xor1), .fs_or0(h_arrdiv16_fs33_or0));
  fs fs_h_arrdiv16_fs34_out(.a(h_arrdiv16_mux2to116_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs33_or0[0]), .fs_xor1(h_arrdiv16_fs34_xor1), .fs_or0(h_arrdiv16_fs34_or0));
  fs fs_h_arrdiv16_fs35_out(.a(h_arrdiv16_mux2to117_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs34_or0[0]), .fs_xor1(h_arrdiv16_fs35_xor1), .fs_or0(h_arrdiv16_fs35_or0));
  fs fs_h_arrdiv16_fs36_out(.a(h_arrdiv16_mux2to118_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs35_or0[0]), .fs_xor1(h_arrdiv16_fs36_xor1), .fs_or0(h_arrdiv16_fs36_or0));
  fs fs_h_arrdiv16_fs37_out(.a(h_arrdiv16_mux2to119_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs36_or0[0]), .fs_xor1(h_arrdiv16_fs37_xor1), .fs_or0(h_arrdiv16_fs37_or0));
  fs fs_h_arrdiv16_fs38_out(.a(h_arrdiv16_mux2to120_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs37_or0[0]), .fs_xor1(h_arrdiv16_fs38_xor1), .fs_or0(h_arrdiv16_fs38_or0));
  fs fs_h_arrdiv16_fs39_out(.a(h_arrdiv16_mux2to121_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs38_or0[0]), .fs_xor1(h_arrdiv16_fs39_xor1), .fs_or0(h_arrdiv16_fs39_or0));
  fs fs_h_arrdiv16_fs40_out(.a(h_arrdiv16_mux2to122_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs39_or0[0]), .fs_xor1(h_arrdiv16_fs40_xor1), .fs_or0(h_arrdiv16_fs40_or0));
  fs fs_h_arrdiv16_fs41_out(.a(h_arrdiv16_mux2to123_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs40_or0[0]), .fs_xor1(h_arrdiv16_fs41_xor1), .fs_or0(h_arrdiv16_fs41_or0));
  fs fs_h_arrdiv16_fs42_out(.a(h_arrdiv16_mux2to124_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs41_or0[0]), .fs_xor1(h_arrdiv16_fs42_xor1), .fs_or0(h_arrdiv16_fs42_or0));
  fs fs_h_arrdiv16_fs43_out(.a(h_arrdiv16_mux2to125_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs42_or0[0]), .fs_xor1(h_arrdiv16_fs43_xor1), .fs_or0(h_arrdiv16_fs43_or0));
  fs fs_h_arrdiv16_fs44_out(.a(h_arrdiv16_mux2to126_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs43_or0[0]), .fs_xor1(h_arrdiv16_fs44_xor1), .fs_or0(h_arrdiv16_fs44_or0));
  fs fs_h_arrdiv16_fs45_out(.a(h_arrdiv16_mux2to127_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs44_or0[0]), .fs_xor1(h_arrdiv16_fs45_xor1), .fs_or0(h_arrdiv16_fs45_or0));
  fs fs_h_arrdiv16_fs46_out(.a(h_arrdiv16_mux2to128_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs45_or0[0]), .fs_xor1(h_arrdiv16_fs46_xor1), .fs_or0(h_arrdiv16_fs46_or0));
  fs fs_h_arrdiv16_fs47_out(.a(h_arrdiv16_mux2to129_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs46_or0[0]), .fs_xor1(h_arrdiv16_fs47_xor1), .fs_or0(h_arrdiv16_fs47_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to130_out(.d0(h_arrdiv16_fs32_xor0[0]), .d1(a[13]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to130_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to131_out(.d0(h_arrdiv16_fs33_xor1[0]), .d1(h_arrdiv16_mux2to115_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to131_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to132_out(.d0(h_arrdiv16_fs34_xor1[0]), .d1(h_arrdiv16_mux2to116_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to132_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to133_out(.d0(h_arrdiv16_fs35_xor1[0]), .d1(h_arrdiv16_mux2to117_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to133_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to134_out(.d0(h_arrdiv16_fs36_xor1[0]), .d1(h_arrdiv16_mux2to118_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to134_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to135_out(.d0(h_arrdiv16_fs37_xor1[0]), .d1(h_arrdiv16_mux2to119_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to135_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to136_out(.d0(h_arrdiv16_fs38_xor1[0]), .d1(h_arrdiv16_mux2to120_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to136_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to137_out(.d0(h_arrdiv16_fs39_xor1[0]), .d1(h_arrdiv16_mux2to121_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to137_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to138_out(.d0(h_arrdiv16_fs40_xor1[0]), .d1(h_arrdiv16_mux2to122_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to138_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to139_out(.d0(h_arrdiv16_fs41_xor1[0]), .d1(h_arrdiv16_mux2to123_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to139_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to140_out(.d0(h_arrdiv16_fs42_xor1[0]), .d1(h_arrdiv16_mux2to124_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to140_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to141_out(.d0(h_arrdiv16_fs43_xor1[0]), .d1(h_arrdiv16_mux2to125_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to141_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to142_out(.d0(h_arrdiv16_fs44_xor1[0]), .d1(h_arrdiv16_mux2to126_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to142_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to143_out(.d0(h_arrdiv16_fs45_xor1[0]), .d1(h_arrdiv16_mux2to127_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to143_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to144_out(.d0(h_arrdiv16_fs46_xor1[0]), .d1(h_arrdiv16_mux2to128_xor0[0]), .sel(h_arrdiv16_fs47_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to144_xor0));
  not_gate not_gate_h_arrdiv16_not2(.a(h_arrdiv16_fs47_or0[0]), .out(h_arrdiv16_not2));
  fs fs_h_arrdiv16_fs48_out(.a(a[12]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs48_xor0), .fs_or0(h_arrdiv16_fs48_and0));
  fs fs_h_arrdiv16_fs49_out(.a(h_arrdiv16_mux2to130_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs48_and0[0]), .fs_xor1(h_arrdiv16_fs49_xor1), .fs_or0(h_arrdiv16_fs49_or0));
  fs fs_h_arrdiv16_fs50_out(.a(h_arrdiv16_mux2to131_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs49_or0[0]), .fs_xor1(h_arrdiv16_fs50_xor1), .fs_or0(h_arrdiv16_fs50_or0));
  fs fs_h_arrdiv16_fs51_out(.a(h_arrdiv16_mux2to132_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs50_or0[0]), .fs_xor1(h_arrdiv16_fs51_xor1), .fs_or0(h_arrdiv16_fs51_or0));
  fs fs_h_arrdiv16_fs52_out(.a(h_arrdiv16_mux2to133_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs51_or0[0]), .fs_xor1(h_arrdiv16_fs52_xor1), .fs_or0(h_arrdiv16_fs52_or0));
  fs fs_h_arrdiv16_fs53_out(.a(h_arrdiv16_mux2to134_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs52_or0[0]), .fs_xor1(h_arrdiv16_fs53_xor1), .fs_or0(h_arrdiv16_fs53_or0));
  fs fs_h_arrdiv16_fs54_out(.a(h_arrdiv16_mux2to135_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs53_or0[0]), .fs_xor1(h_arrdiv16_fs54_xor1), .fs_or0(h_arrdiv16_fs54_or0));
  fs fs_h_arrdiv16_fs55_out(.a(h_arrdiv16_mux2to136_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs54_or0[0]), .fs_xor1(h_arrdiv16_fs55_xor1), .fs_or0(h_arrdiv16_fs55_or0));
  fs fs_h_arrdiv16_fs56_out(.a(h_arrdiv16_mux2to137_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs55_or0[0]), .fs_xor1(h_arrdiv16_fs56_xor1), .fs_or0(h_arrdiv16_fs56_or0));
  fs fs_h_arrdiv16_fs57_out(.a(h_arrdiv16_mux2to138_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs56_or0[0]), .fs_xor1(h_arrdiv16_fs57_xor1), .fs_or0(h_arrdiv16_fs57_or0));
  fs fs_h_arrdiv16_fs58_out(.a(h_arrdiv16_mux2to139_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs57_or0[0]), .fs_xor1(h_arrdiv16_fs58_xor1), .fs_or0(h_arrdiv16_fs58_or0));
  fs fs_h_arrdiv16_fs59_out(.a(h_arrdiv16_mux2to140_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs58_or0[0]), .fs_xor1(h_arrdiv16_fs59_xor1), .fs_or0(h_arrdiv16_fs59_or0));
  fs fs_h_arrdiv16_fs60_out(.a(h_arrdiv16_mux2to141_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs59_or0[0]), .fs_xor1(h_arrdiv16_fs60_xor1), .fs_or0(h_arrdiv16_fs60_or0));
  fs fs_h_arrdiv16_fs61_out(.a(h_arrdiv16_mux2to142_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs60_or0[0]), .fs_xor1(h_arrdiv16_fs61_xor1), .fs_or0(h_arrdiv16_fs61_or0));
  fs fs_h_arrdiv16_fs62_out(.a(h_arrdiv16_mux2to143_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs61_or0[0]), .fs_xor1(h_arrdiv16_fs62_xor1), .fs_or0(h_arrdiv16_fs62_or0));
  fs fs_h_arrdiv16_fs63_out(.a(h_arrdiv16_mux2to144_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs62_or0[0]), .fs_xor1(h_arrdiv16_fs63_xor1), .fs_or0(h_arrdiv16_fs63_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to145_out(.d0(h_arrdiv16_fs48_xor0[0]), .d1(a[12]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to145_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to146_out(.d0(h_arrdiv16_fs49_xor1[0]), .d1(h_arrdiv16_mux2to130_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to146_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to147_out(.d0(h_arrdiv16_fs50_xor1[0]), .d1(h_arrdiv16_mux2to131_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to147_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to148_out(.d0(h_arrdiv16_fs51_xor1[0]), .d1(h_arrdiv16_mux2to132_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to148_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to149_out(.d0(h_arrdiv16_fs52_xor1[0]), .d1(h_arrdiv16_mux2to133_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to149_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to150_out(.d0(h_arrdiv16_fs53_xor1[0]), .d1(h_arrdiv16_mux2to134_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to150_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to151_out(.d0(h_arrdiv16_fs54_xor1[0]), .d1(h_arrdiv16_mux2to135_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to151_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to152_out(.d0(h_arrdiv16_fs55_xor1[0]), .d1(h_arrdiv16_mux2to136_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to152_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to153_out(.d0(h_arrdiv16_fs56_xor1[0]), .d1(h_arrdiv16_mux2to137_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to153_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to154_out(.d0(h_arrdiv16_fs57_xor1[0]), .d1(h_arrdiv16_mux2to138_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to154_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to155_out(.d0(h_arrdiv16_fs58_xor1[0]), .d1(h_arrdiv16_mux2to139_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to155_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to156_out(.d0(h_arrdiv16_fs59_xor1[0]), .d1(h_arrdiv16_mux2to140_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to156_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to157_out(.d0(h_arrdiv16_fs60_xor1[0]), .d1(h_arrdiv16_mux2to141_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to157_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to158_out(.d0(h_arrdiv16_fs61_xor1[0]), .d1(h_arrdiv16_mux2to142_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to158_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to159_out(.d0(h_arrdiv16_fs62_xor1[0]), .d1(h_arrdiv16_mux2to143_xor0[0]), .sel(h_arrdiv16_fs63_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to159_xor0));
  not_gate not_gate_h_arrdiv16_not3(.a(h_arrdiv16_fs63_or0[0]), .out(h_arrdiv16_not3));
  fs fs_h_arrdiv16_fs64_out(.a(a[11]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs64_xor0), .fs_or0(h_arrdiv16_fs64_and0));
  fs fs_h_arrdiv16_fs65_out(.a(h_arrdiv16_mux2to145_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs64_and0[0]), .fs_xor1(h_arrdiv16_fs65_xor1), .fs_or0(h_arrdiv16_fs65_or0));
  fs fs_h_arrdiv16_fs66_out(.a(h_arrdiv16_mux2to146_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs65_or0[0]), .fs_xor1(h_arrdiv16_fs66_xor1), .fs_or0(h_arrdiv16_fs66_or0));
  fs fs_h_arrdiv16_fs67_out(.a(h_arrdiv16_mux2to147_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs66_or0[0]), .fs_xor1(h_arrdiv16_fs67_xor1), .fs_or0(h_arrdiv16_fs67_or0));
  fs fs_h_arrdiv16_fs68_out(.a(h_arrdiv16_mux2to148_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs67_or0[0]), .fs_xor1(h_arrdiv16_fs68_xor1), .fs_or0(h_arrdiv16_fs68_or0));
  fs fs_h_arrdiv16_fs69_out(.a(h_arrdiv16_mux2to149_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs68_or0[0]), .fs_xor1(h_arrdiv16_fs69_xor1), .fs_or0(h_arrdiv16_fs69_or0));
  fs fs_h_arrdiv16_fs70_out(.a(h_arrdiv16_mux2to150_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs69_or0[0]), .fs_xor1(h_arrdiv16_fs70_xor1), .fs_or0(h_arrdiv16_fs70_or0));
  fs fs_h_arrdiv16_fs71_out(.a(h_arrdiv16_mux2to151_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs70_or0[0]), .fs_xor1(h_arrdiv16_fs71_xor1), .fs_or0(h_arrdiv16_fs71_or0));
  fs fs_h_arrdiv16_fs72_out(.a(h_arrdiv16_mux2to152_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs71_or0[0]), .fs_xor1(h_arrdiv16_fs72_xor1), .fs_or0(h_arrdiv16_fs72_or0));
  fs fs_h_arrdiv16_fs73_out(.a(h_arrdiv16_mux2to153_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs72_or0[0]), .fs_xor1(h_arrdiv16_fs73_xor1), .fs_or0(h_arrdiv16_fs73_or0));
  fs fs_h_arrdiv16_fs74_out(.a(h_arrdiv16_mux2to154_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs73_or0[0]), .fs_xor1(h_arrdiv16_fs74_xor1), .fs_or0(h_arrdiv16_fs74_or0));
  fs fs_h_arrdiv16_fs75_out(.a(h_arrdiv16_mux2to155_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs74_or0[0]), .fs_xor1(h_arrdiv16_fs75_xor1), .fs_or0(h_arrdiv16_fs75_or0));
  fs fs_h_arrdiv16_fs76_out(.a(h_arrdiv16_mux2to156_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs75_or0[0]), .fs_xor1(h_arrdiv16_fs76_xor1), .fs_or0(h_arrdiv16_fs76_or0));
  fs fs_h_arrdiv16_fs77_out(.a(h_arrdiv16_mux2to157_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs76_or0[0]), .fs_xor1(h_arrdiv16_fs77_xor1), .fs_or0(h_arrdiv16_fs77_or0));
  fs fs_h_arrdiv16_fs78_out(.a(h_arrdiv16_mux2to158_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs77_or0[0]), .fs_xor1(h_arrdiv16_fs78_xor1), .fs_or0(h_arrdiv16_fs78_or0));
  fs fs_h_arrdiv16_fs79_out(.a(h_arrdiv16_mux2to159_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs78_or0[0]), .fs_xor1(h_arrdiv16_fs79_xor1), .fs_or0(h_arrdiv16_fs79_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to160_out(.d0(h_arrdiv16_fs64_xor0[0]), .d1(a[11]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to160_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to161_out(.d0(h_arrdiv16_fs65_xor1[0]), .d1(h_arrdiv16_mux2to145_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to161_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to162_out(.d0(h_arrdiv16_fs66_xor1[0]), .d1(h_arrdiv16_mux2to146_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to162_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to163_out(.d0(h_arrdiv16_fs67_xor1[0]), .d1(h_arrdiv16_mux2to147_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to163_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to164_out(.d0(h_arrdiv16_fs68_xor1[0]), .d1(h_arrdiv16_mux2to148_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to164_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to165_out(.d0(h_arrdiv16_fs69_xor1[0]), .d1(h_arrdiv16_mux2to149_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to165_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to166_out(.d0(h_arrdiv16_fs70_xor1[0]), .d1(h_arrdiv16_mux2to150_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to166_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to167_out(.d0(h_arrdiv16_fs71_xor1[0]), .d1(h_arrdiv16_mux2to151_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to167_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to168_out(.d0(h_arrdiv16_fs72_xor1[0]), .d1(h_arrdiv16_mux2to152_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to168_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to169_out(.d0(h_arrdiv16_fs73_xor1[0]), .d1(h_arrdiv16_mux2to153_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to169_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to170_out(.d0(h_arrdiv16_fs74_xor1[0]), .d1(h_arrdiv16_mux2to154_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to170_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to171_out(.d0(h_arrdiv16_fs75_xor1[0]), .d1(h_arrdiv16_mux2to155_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to171_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to172_out(.d0(h_arrdiv16_fs76_xor1[0]), .d1(h_arrdiv16_mux2to156_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to172_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to173_out(.d0(h_arrdiv16_fs77_xor1[0]), .d1(h_arrdiv16_mux2to157_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to173_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to174_out(.d0(h_arrdiv16_fs78_xor1[0]), .d1(h_arrdiv16_mux2to158_xor0[0]), .sel(h_arrdiv16_fs79_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to174_xor0));
  not_gate not_gate_h_arrdiv16_not4(.a(h_arrdiv16_fs79_or0[0]), .out(h_arrdiv16_not4));
  fs fs_h_arrdiv16_fs80_out(.a(a[10]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs80_xor0), .fs_or0(h_arrdiv16_fs80_and0));
  fs fs_h_arrdiv16_fs81_out(.a(h_arrdiv16_mux2to160_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs80_and0[0]), .fs_xor1(h_arrdiv16_fs81_xor1), .fs_or0(h_arrdiv16_fs81_or0));
  fs fs_h_arrdiv16_fs82_out(.a(h_arrdiv16_mux2to161_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs81_or0[0]), .fs_xor1(h_arrdiv16_fs82_xor1), .fs_or0(h_arrdiv16_fs82_or0));
  fs fs_h_arrdiv16_fs83_out(.a(h_arrdiv16_mux2to162_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs82_or0[0]), .fs_xor1(h_arrdiv16_fs83_xor1), .fs_or0(h_arrdiv16_fs83_or0));
  fs fs_h_arrdiv16_fs84_out(.a(h_arrdiv16_mux2to163_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs83_or0[0]), .fs_xor1(h_arrdiv16_fs84_xor1), .fs_or0(h_arrdiv16_fs84_or0));
  fs fs_h_arrdiv16_fs85_out(.a(h_arrdiv16_mux2to164_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs84_or0[0]), .fs_xor1(h_arrdiv16_fs85_xor1), .fs_or0(h_arrdiv16_fs85_or0));
  fs fs_h_arrdiv16_fs86_out(.a(h_arrdiv16_mux2to165_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs85_or0[0]), .fs_xor1(h_arrdiv16_fs86_xor1), .fs_or0(h_arrdiv16_fs86_or0));
  fs fs_h_arrdiv16_fs87_out(.a(h_arrdiv16_mux2to166_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs86_or0[0]), .fs_xor1(h_arrdiv16_fs87_xor1), .fs_or0(h_arrdiv16_fs87_or0));
  fs fs_h_arrdiv16_fs88_out(.a(h_arrdiv16_mux2to167_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs87_or0[0]), .fs_xor1(h_arrdiv16_fs88_xor1), .fs_or0(h_arrdiv16_fs88_or0));
  fs fs_h_arrdiv16_fs89_out(.a(h_arrdiv16_mux2to168_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs88_or0[0]), .fs_xor1(h_arrdiv16_fs89_xor1), .fs_or0(h_arrdiv16_fs89_or0));
  fs fs_h_arrdiv16_fs90_out(.a(h_arrdiv16_mux2to169_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs89_or0[0]), .fs_xor1(h_arrdiv16_fs90_xor1), .fs_or0(h_arrdiv16_fs90_or0));
  fs fs_h_arrdiv16_fs91_out(.a(h_arrdiv16_mux2to170_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs90_or0[0]), .fs_xor1(h_arrdiv16_fs91_xor1), .fs_or0(h_arrdiv16_fs91_or0));
  fs fs_h_arrdiv16_fs92_out(.a(h_arrdiv16_mux2to171_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs91_or0[0]), .fs_xor1(h_arrdiv16_fs92_xor1), .fs_or0(h_arrdiv16_fs92_or0));
  fs fs_h_arrdiv16_fs93_out(.a(h_arrdiv16_mux2to172_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs92_or0[0]), .fs_xor1(h_arrdiv16_fs93_xor1), .fs_or0(h_arrdiv16_fs93_or0));
  fs fs_h_arrdiv16_fs94_out(.a(h_arrdiv16_mux2to173_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs93_or0[0]), .fs_xor1(h_arrdiv16_fs94_xor1), .fs_or0(h_arrdiv16_fs94_or0));
  fs fs_h_arrdiv16_fs95_out(.a(h_arrdiv16_mux2to174_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs94_or0[0]), .fs_xor1(h_arrdiv16_fs95_xor1), .fs_or0(h_arrdiv16_fs95_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to175_out(.d0(h_arrdiv16_fs80_xor0[0]), .d1(a[10]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to175_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to176_out(.d0(h_arrdiv16_fs81_xor1[0]), .d1(h_arrdiv16_mux2to160_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to176_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to177_out(.d0(h_arrdiv16_fs82_xor1[0]), .d1(h_arrdiv16_mux2to161_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to177_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to178_out(.d0(h_arrdiv16_fs83_xor1[0]), .d1(h_arrdiv16_mux2to162_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to178_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to179_out(.d0(h_arrdiv16_fs84_xor1[0]), .d1(h_arrdiv16_mux2to163_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to179_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to180_out(.d0(h_arrdiv16_fs85_xor1[0]), .d1(h_arrdiv16_mux2to164_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to180_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to181_out(.d0(h_arrdiv16_fs86_xor1[0]), .d1(h_arrdiv16_mux2to165_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to181_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to182_out(.d0(h_arrdiv16_fs87_xor1[0]), .d1(h_arrdiv16_mux2to166_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to182_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to183_out(.d0(h_arrdiv16_fs88_xor1[0]), .d1(h_arrdiv16_mux2to167_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to183_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to184_out(.d0(h_arrdiv16_fs89_xor1[0]), .d1(h_arrdiv16_mux2to168_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to184_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to185_out(.d0(h_arrdiv16_fs90_xor1[0]), .d1(h_arrdiv16_mux2to169_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to185_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to186_out(.d0(h_arrdiv16_fs91_xor1[0]), .d1(h_arrdiv16_mux2to170_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to186_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to187_out(.d0(h_arrdiv16_fs92_xor1[0]), .d1(h_arrdiv16_mux2to171_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to187_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to188_out(.d0(h_arrdiv16_fs93_xor1[0]), .d1(h_arrdiv16_mux2to172_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to188_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to189_out(.d0(h_arrdiv16_fs94_xor1[0]), .d1(h_arrdiv16_mux2to173_xor0[0]), .sel(h_arrdiv16_fs95_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to189_xor0));
  not_gate not_gate_h_arrdiv16_not5(.a(h_arrdiv16_fs95_or0[0]), .out(h_arrdiv16_not5));
  fs fs_h_arrdiv16_fs96_out(.a(a[9]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs96_xor0), .fs_or0(h_arrdiv16_fs96_and0));
  fs fs_h_arrdiv16_fs97_out(.a(h_arrdiv16_mux2to175_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs96_and0[0]), .fs_xor1(h_arrdiv16_fs97_xor1), .fs_or0(h_arrdiv16_fs97_or0));
  fs fs_h_arrdiv16_fs98_out(.a(h_arrdiv16_mux2to176_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs97_or0[0]), .fs_xor1(h_arrdiv16_fs98_xor1), .fs_or0(h_arrdiv16_fs98_or0));
  fs fs_h_arrdiv16_fs99_out(.a(h_arrdiv16_mux2to177_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs98_or0[0]), .fs_xor1(h_arrdiv16_fs99_xor1), .fs_or0(h_arrdiv16_fs99_or0));
  fs fs_h_arrdiv16_fs100_out(.a(h_arrdiv16_mux2to178_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs99_or0[0]), .fs_xor1(h_arrdiv16_fs100_xor1), .fs_or0(h_arrdiv16_fs100_or0));
  fs fs_h_arrdiv16_fs101_out(.a(h_arrdiv16_mux2to179_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs100_or0[0]), .fs_xor1(h_arrdiv16_fs101_xor1), .fs_or0(h_arrdiv16_fs101_or0));
  fs fs_h_arrdiv16_fs102_out(.a(h_arrdiv16_mux2to180_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs101_or0[0]), .fs_xor1(h_arrdiv16_fs102_xor1), .fs_or0(h_arrdiv16_fs102_or0));
  fs fs_h_arrdiv16_fs103_out(.a(h_arrdiv16_mux2to181_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs102_or0[0]), .fs_xor1(h_arrdiv16_fs103_xor1), .fs_or0(h_arrdiv16_fs103_or0));
  fs fs_h_arrdiv16_fs104_out(.a(h_arrdiv16_mux2to182_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs103_or0[0]), .fs_xor1(h_arrdiv16_fs104_xor1), .fs_or0(h_arrdiv16_fs104_or0));
  fs fs_h_arrdiv16_fs105_out(.a(h_arrdiv16_mux2to183_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs104_or0[0]), .fs_xor1(h_arrdiv16_fs105_xor1), .fs_or0(h_arrdiv16_fs105_or0));
  fs fs_h_arrdiv16_fs106_out(.a(h_arrdiv16_mux2to184_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs105_or0[0]), .fs_xor1(h_arrdiv16_fs106_xor1), .fs_or0(h_arrdiv16_fs106_or0));
  fs fs_h_arrdiv16_fs107_out(.a(h_arrdiv16_mux2to185_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs106_or0[0]), .fs_xor1(h_arrdiv16_fs107_xor1), .fs_or0(h_arrdiv16_fs107_or0));
  fs fs_h_arrdiv16_fs108_out(.a(h_arrdiv16_mux2to186_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs107_or0[0]), .fs_xor1(h_arrdiv16_fs108_xor1), .fs_or0(h_arrdiv16_fs108_or0));
  fs fs_h_arrdiv16_fs109_out(.a(h_arrdiv16_mux2to187_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs108_or0[0]), .fs_xor1(h_arrdiv16_fs109_xor1), .fs_or0(h_arrdiv16_fs109_or0));
  fs fs_h_arrdiv16_fs110_out(.a(h_arrdiv16_mux2to188_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs109_or0[0]), .fs_xor1(h_arrdiv16_fs110_xor1), .fs_or0(h_arrdiv16_fs110_or0));
  fs fs_h_arrdiv16_fs111_out(.a(h_arrdiv16_mux2to189_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs110_or0[0]), .fs_xor1(h_arrdiv16_fs111_xor1), .fs_or0(h_arrdiv16_fs111_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to190_out(.d0(h_arrdiv16_fs96_xor0[0]), .d1(a[9]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to190_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to191_out(.d0(h_arrdiv16_fs97_xor1[0]), .d1(h_arrdiv16_mux2to175_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to191_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to192_out(.d0(h_arrdiv16_fs98_xor1[0]), .d1(h_arrdiv16_mux2to176_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to192_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to193_out(.d0(h_arrdiv16_fs99_xor1[0]), .d1(h_arrdiv16_mux2to177_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to193_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to194_out(.d0(h_arrdiv16_fs100_xor1[0]), .d1(h_arrdiv16_mux2to178_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to194_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to195_out(.d0(h_arrdiv16_fs101_xor1[0]), .d1(h_arrdiv16_mux2to179_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to195_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to196_out(.d0(h_arrdiv16_fs102_xor1[0]), .d1(h_arrdiv16_mux2to180_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to196_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to197_out(.d0(h_arrdiv16_fs103_xor1[0]), .d1(h_arrdiv16_mux2to181_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to197_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to198_out(.d0(h_arrdiv16_fs104_xor1[0]), .d1(h_arrdiv16_mux2to182_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to198_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to199_out(.d0(h_arrdiv16_fs105_xor1[0]), .d1(h_arrdiv16_mux2to183_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to199_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1100_out(.d0(h_arrdiv16_fs106_xor1[0]), .d1(h_arrdiv16_mux2to184_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1100_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1101_out(.d0(h_arrdiv16_fs107_xor1[0]), .d1(h_arrdiv16_mux2to185_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1101_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1102_out(.d0(h_arrdiv16_fs108_xor1[0]), .d1(h_arrdiv16_mux2to186_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1102_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1103_out(.d0(h_arrdiv16_fs109_xor1[0]), .d1(h_arrdiv16_mux2to187_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1103_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1104_out(.d0(h_arrdiv16_fs110_xor1[0]), .d1(h_arrdiv16_mux2to188_xor0[0]), .sel(h_arrdiv16_fs111_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1104_xor0));
  not_gate not_gate_h_arrdiv16_not6(.a(h_arrdiv16_fs111_or0[0]), .out(h_arrdiv16_not6));
  fs fs_h_arrdiv16_fs112_out(.a(a[8]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs112_xor0), .fs_or0(h_arrdiv16_fs112_and0));
  fs fs_h_arrdiv16_fs113_out(.a(h_arrdiv16_mux2to190_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs112_and0[0]), .fs_xor1(h_arrdiv16_fs113_xor1), .fs_or0(h_arrdiv16_fs113_or0));
  fs fs_h_arrdiv16_fs114_out(.a(h_arrdiv16_mux2to191_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs113_or0[0]), .fs_xor1(h_arrdiv16_fs114_xor1), .fs_or0(h_arrdiv16_fs114_or0));
  fs fs_h_arrdiv16_fs115_out(.a(h_arrdiv16_mux2to192_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs114_or0[0]), .fs_xor1(h_arrdiv16_fs115_xor1), .fs_or0(h_arrdiv16_fs115_or0));
  fs fs_h_arrdiv16_fs116_out(.a(h_arrdiv16_mux2to193_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs115_or0[0]), .fs_xor1(h_arrdiv16_fs116_xor1), .fs_or0(h_arrdiv16_fs116_or0));
  fs fs_h_arrdiv16_fs117_out(.a(h_arrdiv16_mux2to194_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs116_or0[0]), .fs_xor1(h_arrdiv16_fs117_xor1), .fs_or0(h_arrdiv16_fs117_or0));
  fs fs_h_arrdiv16_fs118_out(.a(h_arrdiv16_mux2to195_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs117_or0[0]), .fs_xor1(h_arrdiv16_fs118_xor1), .fs_or0(h_arrdiv16_fs118_or0));
  fs fs_h_arrdiv16_fs119_out(.a(h_arrdiv16_mux2to196_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs118_or0[0]), .fs_xor1(h_arrdiv16_fs119_xor1), .fs_or0(h_arrdiv16_fs119_or0));
  fs fs_h_arrdiv16_fs120_out(.a(h_arrdiv16_mux2to197_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs119_or0[0]), .fs_xor1(h_arrdiv16_fs120_xor1), .fs_or0(h_arrdiv16_fs120_or0));
  fs fs_h_arrdiv16_fs121_out(.a(h_arrdiv16_mux2to198_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs120_or0[0]), .fs_xor1(h_arrdiv16_fs121_xor1), .fs_or0(h_arrdiv16_fs121_or0));
  fs fs_h_arrdiv16_fs122_out(.a(h_arrdiv16_mux2to199_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs121_or0[0]), .fs_xor1(h_arrdiv16_fs122_xor1), .fs_or0(h_arrdiv16_fs122_or0));
  fs fs_h_arrdiv16_fs123_out(.a(h_arrdiv16_mux2to1100_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs122_or0[0]), .fs_xor1(h_arrdiv16_fs123_xor1), .fs_or0(h_arrdiv16_fs123_or0));
  fs fs_h_arrdiv16_fs124_out(.a(h_arrdiv16_mux2to1101_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs123_or0[0]), .fs_xor1(h_arrdiv16_fs124_xor1), .fs_or0(h_arrdiv16_fs124_or0));
  fs fs_h_arrdiv16_fs125_out(.a(h_arrdiv16_mux2to1102_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs124_or0[0]), .fs_xor1(h_arrdiv16_fs125_xor1), .fs_or0(h_arrdiv16_fs125_or0));
  fs fs_h_arrdiv16_fs126_out(.a(h_arrdiv16_mux2to1103_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs125_or0[0]), .fs_xor1(h_arrdiv16_fs126_xor1), .fs_or0(h_arrdiv16_fs126_or0));
  fs fs_h_arrdiv16_fs127_out(.a(h_arrdiv16_mux2to1104_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs126_or0[0]), .fs_xor1(h_arrdiv16_fs127_xor1), .fs_or0(h_arrdiv16_fs127_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1105_out(.d0(h_arrdiv16_fs112_xor0[0]), .d1(a[8]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1105_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1106_out(.d0(h_arrdiv16_fs113_xor1[0]), .d1(h_arrdiv16_mux2to190_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1106_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1107_out(.d0(h_arrdiv16_fs114_xor1[0]), .d1(h_arrdiv16_mux2to191_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1107_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1108_out(.d0(h_arrdiv16_fs115_xor1[0]), .d1(h_arrdiv16_mux2to192_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1108_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1109_out(.d0(h_arrdiv16_fs116_xor1[0]), .d1(h_arrdiv16_mux2to193_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1109_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1110_out(.d0(h_arrdiv16_fs117_xor1[0]), .d1(h_arrdiv16_mux2to194_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1110_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1111_out(.d0(h_arrdiv16_fs118_xor1[0]), .d1(h_arrdiv16_mux2to195_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1111_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1112_out(.d0(h_arrdiv16_fs119_xor1[0]), .d1(h_arrdiv16_mux2to196_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1112_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1113_out(.d0(h_arrdiv16_fs120_xor1[0]), .d1(h_arrdiv16_mux2to197_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1113_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1114_out(.d0(h_arrdiv16_fs121_xor1[0]), .d1(h_arrdiv16_mux2to198_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1114_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1115_out(.d0(h_arrdiv16_fs122_xor1[0]), .d1(h_arrdiv16_mux2to199_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1115_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1116_out(.d0(h_arrdiv16_fs123_xor1[0]), .d1(h_arrdiv16_mux2to1100_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1116_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1117_out(.d0(h_arrdiv16_fs124_xor1[0]), .d1(h_arrdiv16_mux2to1101_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1117_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1118_out(.d0(h_arrdiv16_fs125_xor1[0]), .d1(h_arrdiv16_mux2to1102_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1118_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1119_out(.d0(h_arrdiv16_fs126_xor1[0]), .d1(h_arrdiv16_mux2to1103_xor0[0]), .sel(h_arrdiv16_fs127_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1119_xor0));
  not_gate not_gate_h_arrdiv16_not7(.a(h_arrdiv16_fs127_or0[0]), .out(h_arrdiv16_not7));
  fs fs_h_arrdiv16_fs128_out(.a(a[7]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs128_xor0), .fs_or0(h_arrdiv16_fs128_and0));
  fs fs_h_arrdiv16_fs129_out(.a(h_arrdiv16_mux2to1105_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs128_and0[0]), .fs_xor1(h_arrdiv16_fs129_xor1), .fs_or0(h_arrdiv16_fs129_or0));
  fs fs_h_arrdiv16_fs130_out(.a(h_arrdiv16_mux2to1106_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs129_or0[0]), .fs_xor1(h_arrdiv16_fs130_xor1), .fs_or0(h_arrdiv16_fs130_or0));
  fs fs_h_arrdiv16_fs131_out(.a(h_arrdiv16_mux2to1107_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs130_or0[0]), .fs_xor1(h_arrdiv16_fs131_xor1), .fs_or0(h_arrdiv16_fs131_or0));
  fs fs_h_arrdiv16_fs132_out(.a(h_arrdiv16_mux2to1108_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs131_or0[0]), .fs_xor1(h_arrdiv16_fs132_xor1), .fs_or0(h_arrdiv16_fs132_or0));
  fs fs_h_arrdiv16_fs133_out(.a(h_arrdiv16_mux2to1109_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs132_or0[0]), .fs_xor1(h_arrdiv16_fs133_xor1), .fs_or0(h_arrdiv16_fs133_or0));
  fs fs_h_arrdiv16_fs134_out(.a(h_arrdiv16_mux2to1110_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs133_or0[0]), .fs_xor1(h_arrdiv16_fs134_xor1), .fs_or0(h_arrdiv16_fs134_or0));
  fs fs_h_arrdiv16_fs135_out(.a(h_arrdiv16_mux2to1111_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs134_or0[0]), .fs_xor1(h_arrdiv16_fs135_xor1), .fs_or0(h_arrdiv16_fs135_or0));
  fs fs_h_arrdiv16_fs136_out(.a(h_arrdiv16_mux2to1112_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs135_or0[0]), .fs_xor1(h_arrdiv16_fs136_xor1), .fs_or0(h_arrdiv16_fs136_or0));
  fs fs_h_arrdiv16_fs137_out(.a(h_arrdiv16_mux2to1113_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs136_or0[0]), .fs_xor1(h_arrdiv16_fs137_xor1), .fs_or0(h_arrdiv16_fs137_or0));
  fs fs_h_arrdiv16_fs138_out(.a(h_arrdiv16_mux2to1114_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs137_or0[0]), .fs_xor1(h_arrdiv16_fs138_xor1), .fs_or0(h_arrdiv16_fs138_or0));
  fs fs_h_arrdiv16_fs139_out(.a(h_arrdiv16_mux2to1115_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs138_or0[0]), .fs_xor1(h_arrdiv16_fs139_xor1), .fs_or0(h_arrdiv16_fs139_or0));
  fs fs_h_arrdiv16_fs140_out(.a(h_arrdiv16_mux2to1116_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs139_or0[0]), .fs_xor1(h_arrdiv16_fs140_xor1), .fs_or0(h_arrdiv16_fs140_or0));
  fs fs_h_arrdiv16_fs141_out(.a(h_arrdiv16_mux2to1117_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs140_or0[0]), .fs_xor1(h_arrdiv16_fs141_xor1), .fs_or0(h_arrdiv16_fs141_or0));
  fs fs_h_arrdiv16_fs142_out(.a(h_arrdiv16_mux2to1118_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs141_or0[0]), .fs_xor1(h_arrdiv16_fs142_xor1), .fs_or0(h_arrdiv16_fs142_or0));
  fs fs_h_arrdiv16_fs143_out(.a(h_arrdiv16_mux2to1119_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs142_or0[0]), .fs_xor1(h_arrdiv16_fs143_xor1), .fs_or0(h_arrdiv16_fs143_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1120_out(.d0(h_arrdiv16_fs128_xor0[0]), .d1(a[7]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1120_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1121_out(.d0(h_arrdiv16_fs129_xor1[0]), .d1(h_arrdiv16_mux2to1105_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1121_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1122_out(.d0(h_arrdiv16_fs130_xor1[0]), .d1(h_arrdiv16_mux2to1106_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1122_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1123_out(.d0(h_arrdiv16_fs131_xor1[0]), .d1(h_arrdiv16_mux2to1107_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1123_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1124_out(.d0(h_arrdiv16_fs132_xor1[0]), .d1(h_arrdiv16_mux2to1108_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1124_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1125_out(.d0(h_arrdiv16_fs133_xor1[0]), .d1(h_arrdiv16_mux2to1109_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1125_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1126_out(.d0(h_arrdiv16_fs134_xor1[0]), .d1(h_arrdiv16_mux2to1110_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1126_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1127_out(.d0(h_arrdiv16_fs135_xor1[0]), .d1(h_arrdiv16_mux2to1111_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1127_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1128_out(.d0(h_arrdiv16_fs136_xor1[0]), .d1(h_arrdiv16_mux2to1112_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1128_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1129_out(.d0(h_arrdiv16_fs137_xor1[0]), .d1(h_arrdiv16_mux2to1113_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1129_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1130_out(.d0(h_arrdiv16_fs138_xor1[0]), .d1(h_arrdiv16_mux2to1114_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1130_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1131_out(.d0(h_arrdiv16_fs139_xor1[0]), .d1(h_arrdiv16_mux2to1115_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1131_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1132_out(.d0(h_arrdiv16_fs140_xor1[0]), .d1(h_arrdiv16_mux2to1116_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1132_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1133_out(.d0(h_arrdiv16_fs141_xor1[0]), .d1(h_arrdiv16_mux2to1117_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1133_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1134_out(.d0(h_arrdiv16_fs142_xor1[0]), .d1(h_arrdiv16_mux2to1118_xor0[0]), .sel(h_arrdiv16_fs143_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1134_xor0));
  not_gate not_gate_h_arrdiv16_not8(.a(h_arrdiv16_fs143_or0[0]), .out(h_arrdiv16_not8));
  fs fs_h_arrdiv16_fs144_out(.a(a[6]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs144_xor0), .fs_or0(h_arrdiv16_fs144_and0));
  fs fs_h_arrdiv16_fs145_out(.a(h_arrdiv16_mux2to1120_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs144_and0[0]), .fs_xor1(h_arrdiv16_fs145_xor1), .fs_or0(h_arrdiv16_fs145_or0));
  fs fs_h_arrdiv16_fs146_out(.a(h_arrdiv16_mux2to1121_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs145_or0[0]), .fs_xor1(h_arrdiv16_fs146_xor1), .fs_or0(h_arrdiv16_fs146_or0));
  fs fs_h_arrdiv16_fs147_out(.a(h_arrdiv16_mux2to1122_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs146_or0[0]), .fs_xor1(h_arrdiv16_fs147_xor1), .fs_or0(h_arrdiv16_fs147_or0));
  fs fs_h_arrdiv16_fs148_out(.a(h_arrdiv16_mux2to1123_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs147_or0[0]), .fs_xor1(h_arrdiv16_fs148_xor1), .fs_or0(h_arrdiv16_fs148_or0));
  fs fs_h_arrdiv16_fs149_out(.a(h_arrdiv16_mux2to1124_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs148_or0[0]), .fs_xor1(h_arrdiv16_fs149_xor1), .fs_or0(h_arrdiv16_fs149_or0));
  fs fs_h_arrdiv16_fs150_out(.a(h_arrdiv16_mux2to1125_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs149_or0[0]), .fs_xor1(h_arrdiv16_fs150_xor1), .fs_or0(h_arrdiv16_fs150_or0));
  fs fs_h_arrdiv16_fs151_out(.a(h_arrdiv16_mux2to1126_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs150_or0[0]), .fs_xor1(h_arrdiv16_fs151_xor1), .fs_or0(h_arrdiv16_fs151_or0));
  fs fs_h_arrdiv16_fs152_out(.a(h_arrdiv16_mux2to1127_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs151_or0[0]), .fs_xor1(h_arrdiv16_fs152_xor1), .fs_or0(h_arrdiv16_fs152_or0));
  fs fs_h_arrdiv16_fs153_out(.a(h_arrdiv16_mux2to1128_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs152_or0[0]), .fs_xor1(h_arrdiv16_fs153_xor1), .fs_or0(h_arrdiv16_fs153_or0));
  fs fs_h_arrdiv16_fs154_out(.a(h_arrdiv16_mux2to1129_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs153_or0[0]), .fs_xor1(h_arrdiv16_fs154_xor1), .fs_or0(h_arrdiv16_fs154_or0));
  fs fs_h_arrdiv16_fs155_out(.a(h_arrdiv16_mux2to1130_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs154_or0[0]), .fs_xor1(h_arrdiv16_fs155_xor1), .fs_or0(h_arrdiv16_fs155_or0));
  fs fs_h_arrdiv16_fs156_out(.a(h_arrdiv16_mux2to1131_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs155_or0[0]), .fs_xor1(h_arrdiv16_fs156_xor1), .fs_or0(h_arrdiv16_fs156_or0));
  fs fs_h_arrdiv16_fs157_out(.a(h_arrdiv16_mux2to1132_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs156_or0[0]), .fs_xor1(h_arrdiv16_fs157_xor1), .fs_or0(h_arrdiv16_fs157_or0));
  fs fs_h_arrdiv16_fs158_out(.a(h_arrdiv16_mux2to1133_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs157_or0[0]), .fs_xor1(h_arrdiv16_fs158_xor1), .fs_or0(h_arrdiv16_fs158_or0));
  fs fs_h_arrdiv16_fs159_out(.a(h_arrdiv16_mux2to1134_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs158_or0[0]), .fs_xor1(h_arrdiv16_fs159_xor1), .fs_or0(h_arrdiv16_fs159_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1135_out(.d0(h_arrdiv16_fs144_xor0[0]), .d1(a[6]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1135_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1136_out(.d0(h_arrdiv16_fs145_xor1[0]), .d1(h_arrdiv16_mux2to1120_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1136_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1137_out(.d0(h_arrdiv16_fs146_xor1[0]), .d1(h_arrdiv16_mux2to1121_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1137_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1138_out(.d0(h_arrdiv16_fs147_xor1[0]), .d1(h_arrdiv16_mux2to1122_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1138_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1139_out(.d0(h_arrdiv16_fs148_xor1[0]), .d1(h_arrdiv16_mux2to1123_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1139_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1140_out(.d0(h_arrdiv16_fs149_xor1[0]), .d1(h_arrdiv16_mux2to1124_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1140_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1141_out(.d0(h_arrdiv16_fs150_xor1[0]), .d1(h_arrdiv16_mux2to1125_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1141_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1142_out(.d0(h_arrdiv16_fs151_xor1[0]), .d1(h_arrdiv16_mux2to1126_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1142_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1143_out(.d0(h_arrdiv16_fs152_xor1[0]), .d1(h_arrdiv16_mux2to1127_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1143_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1144_out(.d0(h_arrdiv16_fs153_xor1[0]), .d1(h_arrdiv16_mux2to1128_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1144_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1145_out(.d0(h_arrdiv16_fs154_xor1[0]), .d1(h_arrdiv16_mux2to1129_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1145_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1146_out(.d0(h_arrdiv16_fs155_xor1[0]), .d1(h_arrdiv16_mux2to1130_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1146_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1147_out(.d0(h_arrdiv16_fs156_xor1[0]), .d1(h_arrdiv16_mux2to1131_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1147_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1148_out(.d0(h_arrdiv16_fs157_xor1[0]), .d1(h_arrdiv16_mux2to1132_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1148_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1149_out(.d0(h_arrdiv16_fs158_xor1[0]), .d1(h_arrdiv16_mux2to1133_xor0[0]), .sel(h_arrdiv16_fs159_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1149_xor0));
  not_gate not_gate_h_arrdiv16_not9(.a(h_arrdiv16_fs159_or0[0]), .out(h_arrdiv16_not9));
  fs fs_h_arrdiv16_fs160_out(.a(a[5]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs160_xor0), .fs_or0(h_arrdiv16_fs160_and0));
  fs fs_h_arrdiv16_fs161_out(.a(h_arrdiv16_mux2to1135_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs160_and0[0]), .fs_xor1(h_arrdiv16_fs161_xor1), .fs_or0(h_arrdiv16_fs161_or0));
  fs fs_h_arrdiv16_fs162_out(.a(h_arrdiv16_mux2to1136_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs161_or0[0]), .fs_xor1(h_arrdiv16_fs162_xor1), .fs_or0(h_arrdiv16_fs162_or0));
  fs fs_h_arrdiv16_fs163_out(.a(h_arrdiv16_mux2to1137_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs162_or0[0]), .fs_xor1(h_arrdiv16_fs163_xor1), .fs_or0(h_arrdiv16_fs163_or0));
  fs fs_h_arrdiv16_fs164_out(.a(h_arrdiv16_mux2to1138_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs163_or0[0]), .fs_xor1(h_arrdiv16_fs164_xor1), .fs_or0(h_arrdiv16_fs164_or0));
  fs fs_h_arrdiv16_fs165_out(.a(h_arrdiv16_mux2to1139_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs164_or0[0]), .fs_xor1(h_arrdiv16_fs165_xor1), .fs_or0(h_arrdiv16_fs165_or0));
  fs fs_h_arrdiv16_fs166_out(.a(h_arrdiv16_mux2to1140_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs165_or0[0]), .fs_xor1(h_arrdiv16_fs166_xor1), .fs_or0(h_arrdiv16_fs166_or0));
  fs fs_h_arrdiv16_fs167_out(.a(h_arrdiv16_mux2to1141_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs166_or0[0]), .fs_xor1(h_arrdiv16_fs167_xor1), .fs_or0(h_arrdiv16_fs167_or0));
  fs fs_h_arrdiv16_fs168_out(.a(h_arrdiv16_mux2to1142_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs167_or0[0]), .fs_xor1(h_arrdiv16_fs168_xor1), .fs_or0(h_arrdiv16_fs168_or0));
  fs fs_h_arrdiv16_fs169_out(.a(h_arrdiv16_mux2to1143_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs168_or0[0]), .fs_xor1(h_arrdiv16_fs169_xor1), .fs_or0(h_arrdiv16_fs169_or0));
  fs fs_h_arrdiv16_fs170_out(.a(h_arrdiv16_mux2to1144_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs169_or0[0]), .fs_xor1(h_arrdiv16_fs170_xor1), .fs_or0(h_arrdiv16_fs170_or0));
  fs fs_h_arrdiv16_fs171_out(.a(h_arrdiv16_mux2to1145_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs170_or0[0]), .fs_xor1(h_arrdiv16_fs171_xor1), .fs_or0(h_arrdiv16_fs171_or0));
  fs fs_h_arrdiv16_fs172_out(.a(h_arrdiv16_mux2to1146_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs171_or0[0]), .fs_xor1(h_arrdiv16_fs172_xor1), .fs_or0(h_arrdiv16_fs172_or0));
  fs fs_h_arrdiv16_fs173_out(.a(h_arrdiv16_mux2to1147_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs172_or0[0]), .fs_xor1(h_arrdiv16_fs173_xor1), .fs_or0(h_arrdiv16_fs173_or0));
  fs fs_h_arrdiv16_fs174_out(.a(h_arrdiv16_mux2to1148_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs173_or0[0]), .fs_xor1(h_arrdiv16_fs174_xor1), .fs_or0(h_arrdiv16_fs174_or0));
  fs fs_h_arrdiv16_fs175_out(.a(h_arrdiv16_mux2to1149_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs174_or0[0]), .fs_xor1(h_arrdiv16_fs175_xor1), .fs_or0(h_arrdiv16_fs175_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1150_out(.d0(h_arrdiv16_fs160_xor0[0]), .d1(a[5]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1150_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1151_out(.d0(h_arrdiv16_fs161_xor1[0]), .d1(h_arrdiv16_mux2to1135_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1151_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1152_out(.d0(h_arrdiv16_fs162_xor1[0]), .d1(h_arrdiv16_mux2to1136_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1152_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1153_out(.d0(h_arrdiv16_fs163_xor1[0]), .d1(h_arrdiv16_mux2to1137_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1153_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1154_out(.d0(h_arrdiv16_fs164_xor1[0]), .d1(h_arrdiv16_mux2to1138_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1154_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1155_out(.d0(h_arrdiv16_fs165_xor1[0]), .d1(h_arrdiv16_mux2to1139_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1155_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1156_out(.d0(h_arrdiv16_fs166_xor1[0]), .d1(h_arrdiv16_mux2to1140_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1156_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1157_out(.d0(h_arrdiv16_fs167_xor1[0]), .d1(h_arrdiv16_mux2to1141_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1157_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1158_out(.d0(h_arrdiv16_fs168_xor1[0]), .d1(h_arrdiv16_mux2to1142_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1158_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1159_out(.d0(h_arrdiv16_fs169_xor1[0]), .d1(h_arrdiv16_mux2to1143_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1159_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1160_out(.d0(h_arrdiv16_fs170_xor1[0]), .d1(h_arrdiv16_mux2to1144_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1160_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1161_out(.d0(h_arrdiv16_fs171_xor1[0]), .d1(h_arrdiv16_mux2to1145_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1161_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1162_out(.d0(h_arrdiv16_fs172_xor1[0]), .d1(h_arrdiv16_mux2to1146_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1162_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1163_out(.d0(h_arrdiv16_fs173_xor1[0]), .d1(h_arrdiv16_mux2to1147_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1163_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1164_out(.d0(h_arrdiv16_fs174_xor1[0]), .d1(h_arrdiv16_mux2to1148_xor0[0]), .sel(h_arrdiv16_fs175_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1164_xor0));
  not_gate not_gate_h_arrdiv16_not10(.a(h_arrdiv16_fs175_or0[0]), .out(h_arrdiv16_not10));
  fs fs_h_arrdiv16_fs176_out(.a(a[4]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs176_xor0), .fs_or0(h_arrdiv16_fs176_and0));
  fs fs_h_arrdiv16_fs177_out(.a(h_arrdiv16_mux2to1150_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs176_and0[0]), .fs_xor1(h_arrdiv16_fs177_xor1), .fs_or0(h_arrdiv16_fs177_or0));
  fs fs_h_arrdiv16_fs178_out(.a(h_arrdiv16_mux2to1151_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs177_or0[0]), .fs_xor1(h_arrdiv16_fs178_xor1), .fs_or0(h_arrdiv16_fs178_or0));
  fs fs_h_arrdiv16_fs179_out(.a(h_arrdiv16_mux2to1152_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs178_or0[0]), .fs_xor1(h_arrdiv16_fs179_xor1), .fs_or0(h_arrdiv16_fs179_or0));
  fs fs_h_arrdiv16_fs180_out(.a(h_arrdiv16_mux2to1153_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs179_or0[0]), .fs_xor1(h_arrdiv16_fs180_xor1), .fs_or0(h_arrdiv16_fs180_or0));
  fs fs_h_arrdiv16_fs181_out(.a(h_arrdiv16_mux2to1154_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs180_or0[0]), .fs_xor1(h_arrdiv16_fs181_xor1), .fs_or0(h_arrdiv16_fs181_or0));
  fs fs_h_arrdiv16_fs182_out(.a(h_arrdiv16_mux2to1155_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs181_or0[0]), .fs_xor1(h_arrdiv16_fs182_xor1), .fs_or0(h_arrdiv16_fs182_or0));
  fs fs_h_arrdiv16_fs183_out(.a(h_arrdiv16_mux2to1156_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs182_or0[0]), .fs_xor1(h_arrdiv16_fs183_xor1), .fs_or0(h_arrdiv16_fs183_or0));
  fs fs_h_arrdiv16_fs184_out(.a(h_arrdiv16_mux2to1157_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs183_or0[0]), .fs_xor1(h_arrdiv16_fs184_xor1), .fs_or0(h_arrdiv16_fs184_or0));
  fs fs_h_arrdiv16_fs185_out(.a(h_arrdiv16_mux2to1158_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs184_or0[0]), .fs_xor1(h_arrdiv16_fs185_xor1), .fs_or0(h_arrdiv16_fs185_or0));
  fs fs_h_arrdiv16_fs186_out(.a(h_arrdiv16_mux2to1159_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs185_or0[0]), .fs_xor1(h_arrdiv16_fs186_xor1), .fs_or0(h_arrdiv16_fs186_or0));
  fs fs_h_arrdiv16_fs187_out(.a(h_arrdiv16_mux2to1160_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs186_or0[0]), .fs_xor1(h_arrdiv16_fs187_xor1), .fs_or0(h_arrdiv16_fs187_or0));
  fs fs_h_arrdiv16_fs188_out(.a(h_arrdiv16_mux2to1161_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs187_or0[0]), .fs_xor1(h_arrdiv16_fs188_xor1), .fs_or0(h_arrdiv16_fs188_or0));
  fs fs_h_arrdiv16_fs189_out(.a(h_arrdiv16_mux2to1162_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs188_or0[0]), .fs_xor1(h_arrdiv16_fs189_xor1), .fs_or0(h_arrdiv16_fs189_or0));
  fs fs_h_arrdiv16_fs190_out(.a(h_arrdiv16_mux2to1163_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs189_or0[0]), .fs_xor1(h_arrdiv16_fs190_xor1), .fs_or0(h_arrdiv16_fs190_or0));
  fs fs_h_arrdiv16_fs191_out(.a(h_arrdiv16_mux2to1164_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs190_or0[0]), .fs_xor1(h_arrdiv16_fs191_xor1), .fs_or0(h_arrdiv16_fs191_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1165_out(.d0(h_arrdiv16_fs176_xor0[0]), .d1(a[4]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1165_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1166_out(.d0(h_arrdiv16_fs177_xor1[0]), .d1(h_arrdiv16_mux2to1150_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1166_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1167_out(.d0(h_arrdiv16_fs178_xor1[0]), .d1(h_arrdiv16_mux2to1151_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1167_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1168_out(.d0(h_arrdiv16_fs179_xor1[0]), .d1(h_arrdiv16_mux2to1152_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1168_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1169_out(.d0(h_arrdiv16_fs180_xor1[0]), .d1(h_arrdiv16_mux2to1153_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1169_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1170_out(.d0(h_arrdiv16_fs181_xor1[0]), .d1(h_arrdiv16_mux2to1154_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1170_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1171_out(.d0(h_arrdiv16_fs182_xor1[0]), .d1(h_arrdiv16_mux2to1155_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1171_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1172_out(.d0(h_arrdiv16_fs183_xor1[0]), .d1(h_arrdiv16_mux2to1156_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1172_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1173_out(.d0(h_arrdiv16_fs184_xor1[0]), .d1(h_arrdiv16_mux2to1157_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1173_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1174_out(.d0(h_arrdiv16_fs185_xor1[0]), .d1(h_arrdiv16_mux2to1158_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1174_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1175_out(.d0(h_arrdiv16_fs186_xor1[0]), .d1(h_arrdiv16_mux2to1159_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1175_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1176_out(.d0(h_arrdiv16_fs187_xor1[0]), .d1(h_arrdiv16_mux2to1160_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1176_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1177_out(.d0(h_arrdiv16_fs188_xor1[0]), .d1(h_arrdiv16_mux2to1161_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1177_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1178_out(.d0(h_arrdiv16_fs189_xor1[0]), .d1(h_arrdiv16_mux2to1162_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1178_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1179_out(.d0(h_arrdiv16_fs190_xor1[0]), .d1(h_arrdiv16_mux2to1163_xor0[0]), .sel(h_arrdiv16_fs191_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1179_xor0));
  not_gate not_gate_h_arrdiv16_not11(.a(h_arrdiv16_fs191_or0[0]), .out(h_arrdiv16_not11));
  fs fs_h_arrdiv16_fs192_out(.a(a[3]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs192_xor0), .fs_or0(h_arrdiv16_fs192_and0));
  fs fs_h_arrdiv16_fs193_out(.a(h_arrdiv16_mux2to1165_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs192_and0[0]), .fs_xor1(h_arrdiv16_fs193_xor1), .fs_or0(h_arrdiv16_fs193_or0));
  fs fs_h_arrdiv16_fs194_out(.a(h_arrdiv16_mux2to1166_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs193_or0[0]), .fs_xor1(h_arrdiv16_fs194_xor1), .fs_or0(h_arrdiv16_fs194_or0));
  fs fs_h_arrdiv16_fs195_out(.a(h_arrdiv16_mux2to1167_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs194_or0[0]), .fs_xor1(h_arrdiv16_fs195_xor1), .fs_or0(h_arrdiv16_fs195_or0));
  fs fs_h_arrdiv16_fs196_out(.a(h_arrdiv16_mux2to1168_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs195_or0[0]), .fs_xor1(h_arrdiv16_fs196_xor1), .fs_or0(h_arrdiv16_fs196_or0));
  fs fs_h_arrdiv16_fs197_out(.a(h_arrdiv16_mux2to1169_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs196_or0[0]), .fs_xor1(h_arrdiv16_fs197_xor1), .fs_or0(h_arrdiv16_fs197_or0));
  fs fs_h_arrdiv16_fs198_out(.a(h_arrdiv16_mux2to1170_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs197_or0[0]), .fs_xor1(h_arrdiv16_fs198_xor1), .fs_or0(h_arrdiv16_fs198_or0));
  fs fs_h_arrdiv16_fs199_out(.a(h_arrdiv16_mux2to1171_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs198_or0[0]), .fs_xor1(h_arrdiv16_fs199_xor1), .fs_or0(h_arrdiv16_fs199_or0));
  fs fs_h_arrdiv16_fs200_out(.a(h_arrdiv16_mux2to1172_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs199_or0[0]), .fs_xor1(h_arrdiv16_fs200_xor1), .fs_or0(h_arrdiv16_fs200_or0));
  fs fs_h_arrdiv16_fs201_out(.a(h_arrdiv16_mux2to1173_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs200_or0[0]), .fs_xor1(h_arrdiv16_fs201_xor1), .fs_or0(h_arrdiv16_fs201_or0));
  fs fs_h_arrdiv16_fs202_out(.a(h_arrdiv16_mux2to1174_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs201_or0[0]), .fs_xor1(h_arrdiv16_fs202_xor1), .fs_or0(h_arrdiv16_fs202_or0));
  fs fs_h_arrdiv16_fs203_out(.a(h_arrdiv16_mux2to1175_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs202_or0[0]), .fs_xor1(h_arrdiv16_fs203_xor1), .fs_or0(h_arrdiv16_fs203_or0));
  fs fs_h_arrdiv16_fs204_out(.a(h_arrdiv16_mux2to1176_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs203_or0[0]), .fs_xor1(h_arrdiv16_fs204_xor1), .fs_or0(h_arrdiv16_fs204_or0));
  fs fs_h_arrdiv16_fs205_out(.a(h_arrdiv16_mux2to1177_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs204_or0[0]), .fs_xor1(h_arrdiv16_fs205_xor1), .fs_or0(h_arrdiv16_fs205_or0));
  fs fs_h_arrdiv16_fs206_out(.a(h_arrdiv16_mux2to1178_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs205_or0[0]), .fs_xor1(h_arrdiv16_fs206_xor1), .fs_or0(h_arrdiv16_fs206_or0));
  fs fs_h_arrdiv16_fs207_out(.a(h_arrdiv16_mux2to1179_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs206_or0[0]), .fs_xor1(h_arrdiv16_fs207_xor1), .fs_or0(h_arrdiv16_fs207_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1180_out(.d0(h_arrdiv16_fs192_xor0[0]), .d1(a[3]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1180_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1181_out(.d0(h_arrdiv16_fs193_xor1[0]), .d1(h_arrdiv16_mux2to1165_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1181_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1182_out(.d0(h_arrdiv16_fs194_xor1[0]), .d1(h_arrdiv16_mux2to1166_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1182_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1183_out(.d0(h_arrdiv16_fs195_xor1[0]), .d1(h_arrdiv16_mux2to1167_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1183_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1184_out(.d0(h_arrdiv16_fs196_xor1[0]), .d1(h_arrdiv16_mux2to1168_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1184_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1185_out(.d0(h_arrdiv16_fs197_xor1[0]), .d1(h_arrdiv16_mux2to1169_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1185_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1186_out(.d0(h_arrdiv16_fs198_xor1[0]), .d1(h_arrdiv16_mux2to1170_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1186_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1187_out(.d0(h_arrdiv16_fs199_xor1[0]), .d1(h_arrdiv16_mux2to1171_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1187_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1188_out(.d0(h_arrdiv16_fs200_xor1[0]), .d1(h_arrdiv16_mux2to1172_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1188_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1189_out(.d0(h_arrdiv16_fs201_xor1[0]), .d1(h_arrdiv16_mux2to1173_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1189_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1190_out(.d0(h_arrdiv16_fs202_xor1[0]), .d1(h_arrdiv16_mux2to1174_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1190_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1191_out(.d0(h_arrdiv16_fs203_xor1[0]), .d1(h_arrdiv16_mux2to1175_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1191_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1192_out(.d0(h_arrdiv16_fs204_xor1[0]), .d1(h_arrdiv16_mux2to1176_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1192_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1193_out(.d0(h_arrdiv16_fs205_xor1[0]), .d1(h_arrdiv16_mux2to1177_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1193_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1194_out(.d0(h_arrdiv16_fs206_xor1[0]), .d1(h_arrdiv16_mux2to1178_xor0[0]), .sel(h_arrdiv16_fs207_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1194_xor0));
  not_gate not_gate_h_arrdiv16_not12(.a(h_arrdiv16_fs207_or0[0]), .out(h_arrdiv16_not12));
  fs fs_h_arrdiv16_fs208_out(.a(a[2]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs208_xor0), .fs_or0(h_arrdiv16_fs208_and0));
  fs fs_h_arrdiv16_fs209_out(.a(h_arrdiv16_mux2to1180_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs208_and0[0]), .fs_xor1(h_arrdiv16_fs209_xor1), .fs_or0(h_arrdiv16_fs209_or0));
  fs fs_h_arrdiv16_fs210_out(.a(h_arrdiv16_mux2to1181_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs209_or0[0]), .fs_xor1(h_arrdiv16_fs210_xor1), .fs_or0(h_arrdiv16_fs210_or0));
  fs fs_h_arrdiv16_fs211_out(.a(h_arrdiv16_mux2to1182_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs210_or0[0]), .fs_xor1(h_arrdiv16_fs211_xor1), .fs_or0(h_arrdiv16_fs211_or0));
  fs fs_h_arrdiv16_fs212_out(.a(h_arrdiv16_mux2to1183_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs211_or0[0]), .fs_xor1(h_arrdiv16_fs212_xor1), .fs_or0(h_arrdiv16_fs212_or0));
  fs fs_h_arrdiv16_fs213_out(.a(h_arrdiv16_mux2to1184_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs212_or0[0]), .fs_xor1(h_arrdiv16_fs213_xor1), .fs_or0(h_arrdiv16_fs213_or0));
  fs fs_h_arrdiv16_fs214_out(.a(h_arrdiv16_mux2to1185_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs213_or0[0]), .fs_xor1(h_arrdiv16_fs214_xor1), .fs_or0(h_arrdiv16_fs214_or0));
  fs fs_h_arrdiv16_fs215_out(.a(h_arrdiv16_mux2to1186_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs214_or0[0]), .fs_xor1(h_arrdiv16_fs215_xor1), .fs_or0(h_arrdiv16_fs215_or0));
  fs fs_h_arrdiv16_fs216_out(.a(h_arrdiv16_mux2to1187_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs215_or0[0]), .fs_xor1(h_arrdiv16_fs216_xor1), .fs_or0(h_arrdiv16_fs216_or0));
  fs fs_h_arrdiv16_fs217_out(.a(h_arrdiv16_mux2to1188_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs216_or0[0]), .fs_xor1(h_arrdiv16_fs217_xor1), .fs_or0(h_arrdiv16_fs217_or0));
  fs fs_h_arrdiv16_fs218_out(.a(h_arrdiv16_mux2to1189_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs217_or0[0]), .fs_xor1(h_arrdiv16_fs218_xor1), .fs_or0(h_arrdiv16_fs218_or0));
  fs fs_h_arrdiv16_fs219_out(.a(h_arrdiv16_mux2to1190_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs218_or0[0]), .fs_xor1(h_arrdiv16_fs219_xor1), .fs_or0(h_arrdiv16_fs219_or0));
  fs fs_h_arrdiv16_fs220_out(.a(h_arrdiv16_mux2to1191_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs219_or0[0]), .fs_xor1(h_arrdiv16_fs220_xor1), .fs_or0(h_arrdiv16_fs220_or0));
  fs fs_h_arrdiv16_fs221_out(.a(h_arrdiv16_mux2to1192_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs220_or0[0]), .fs_xor1(h_arrdiv16_fs221_xor1), .fs_or0(h_arrdiv16_fs221_or0));
  fs fs_h_arrdiv16_fs222_out(.a(h_arrdiv16_mux2to1193_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs221_or0[0]), .fs_xor1(h_arrdiv16_fs222_xor1), .fs_or0(h_arrdiv16_fs222_or0));
  fs fs_h_arrdiv16_fs223_out(.a(h_arrdiv16_mux2to1194_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs222_or0[0]), .fs_xor1(h_arrdiv16_fs223_xor1), .fs_or0(h_arrdiv16_fs223_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1195_out(.d0(h_arrdiv16_fs208_xor0[0]), .d1(a[2]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1195_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1196_out(.d0(h_arrdiv16_fs209_xor1[0]), .d1(h_arrdiv16_mux2to1180_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1196_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1197_out(.d0(h_arrdiv16_fs210_xor1[0]), .d1(h_arrdiv16_mux2to1181_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1197_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1198_out(.d0(h_arrdiv16_fs211_xor1[0]), .d1(h_arrdiv16_mux2to1182_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1198_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1199_out(.d0(h_arrdiv16_fs212_xor1[0]), .d1(h_arrdiv16_mux2to1183_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1199_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1200_out(.d0(h_arrdiv16_fs213_xor1[0]), .d1(h_arrdiv16_mux2to1184_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1200_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1201_out(.d0(h_arrdiv16_fs214_xor1[0]), .d1(h_arrdiv16_mux2to1185_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1201_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1202_out(.d0(h_arrdiv16_fs215_xor1[0]), .d1(h_arrdiv16_mux2to1186_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1202_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1203_out(.d0(h_arrdiv16_fs216_xor1[0]), .d1(h_arrdiv16_mux2to1187_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1203_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1204_out(.d0(h_arrdiv16_fs217_xor1[0]), .d1(h_arrdiv16_mux2to1188_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1204_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1205_out(.d0(h_arrdiv16_fs218_xor1[0]), .d1(h_arrdiv16_mux2to1189_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1205_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1206_out(.d0(h_arrdiv16_fs219_xor1[0]), .d1(h_arrdiv16_mux2to1190_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1206_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1207_out(.d0(h_arrdiv16_fs220_xor1[0]), .d1(h_arrdiv16_mux2to1191_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1207_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1208_out(.d0(h_arrdiv16_fs221_xor1[0]), .d1(h_arrdiv16_mux2to1192_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1208_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1209_out(.d0(h_arrdiv16_fs222_xor1[0]), .d1(h_arrdiv16_mux2to1193_xor0[0]), .sel(h_arrdiv16_fs223_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1209_xor0));
  not_gate not_gate_h_arrdiv16_not13(.a(h_arrdiv16_fs223_or0[0]), .out(h_arrdiv16_not13));
  fs fs_h_arrdiv16_fs224_out(.a(a[1]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs224_xor0), .fs_or0(h_arrdiv16_fs224_and0));
  fs fs_h_arrdiv16_fs225_out(.a(h_arrdiv16_mux2to1195_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs224_and0[0]), .fs_xor1(h_arrdiv16_fs225_xor1), .fs_or0(h_arrdiv16_fs225_or0));
  fs fs_h_arrdiv16_fs226_out(.a(h_arrdiv16_mux2to1196_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs225_or0[0]), .fs_xor1(h_arrdiv16_fs226_xor1), .fs_or0(h_arrdiv16_fs226_or0));
  fs fs_h_arrdiv16_fs227_out(.a(h_arrdiv16_mux2to1197_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs226_or0[0]), .fs_xor1(h_arrdiv16_fs227_xor1), .fs_or0(h_arrdiv16_fs227_or0));
  fs fs_h_arrdiv16_fs228_out(.a(h_arrdiv16_mux2to1198_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs227_or0[0]), .fs_xor1(h_arrdiv16_fs228_xor1), .fs_or0(h_arrdiv16_fs228_or0));
  fs fs_h_arrdiv16_fs229_out(.a(h_arrdiv16_mux2to1199_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs228_or0[0]), .fs_xor1(h_arrdiv16_fs229_xor1), .fs_or0(h_arrdiv16_fs229_or0));
  fs fs_h_arrdiv16_fs230_out(.a(h_arrdiv16_mux2to1200_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs229_or0[0]), .fs_xor1(h_arrdiv16_fs230_xor1), .fs_or0(h_arrdiv16_fs230_or0));
  fs fs_h_arrdiv16_fs231_out(.a(h_arrdiv16_mux2to1201_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs230_or0[0]), .fs_xor1(h_arrdiv16_fs231_xor1), .fs_or0(h_arrdiv16_fs231_or0));
  fs fs_h_arrdiv16_fs232_out(.a(h_arrdiv16_mux2to1202_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs231_or0[0]), .fs_xor1(h_arrdiv16_fs232_xor1), .fs_or0(h_arrdiv16_fs232_or0));
  fs fs_h_arrdiv16_fs233_out(.a(h_arrdiv16_mux2to1203_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs232_or0[0]), .fs_xor1(h_arrdiv16_fs233_xor1), .fs_or0(h_arrdiv16_fs233_or0));
  fs fs_h_arrdiv16_fs234_out(.a(h_arrdiv16_mux2to1204_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs233_or0[0]), .fs_xor1(h_arrdiv16_fs234_xor1), .fs_or0(h_arrdiv16_fs234_or0));
  fs fs_h_arrdiv16_fs235_out(.a(h_arrdiv16_mux2to1205_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs234_or0[0]), .fs_xor1(h_arrdiv16_fs235_xor1), .fs_or0(h_arrdiv16_fs235_or0));
  fs fs_h_arrdiv16_fs236_out(.a(h_arrdiv16_mux2to1206_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs235_or0[0]), .fs_xor1(h_arrdiv16_fs236_xor1), .fs_or0(h_arrdiv16_fs236_or0));
  fs fs_h_arrdiv16_fs237_out(.a(h_arrdiv16_mux2to1207_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs236_or0[0]), .fs_xor1(h_arrdiv16_fs237_xor1), .fs_or0(h_arrdiv16_fs237_or0));
  fs fs_h_arrdiv16_fs238_out(.a(h_arrdiv16_mux2to1208_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs237_or0[0]), .fs_xor1(h_arrdiv16_fs238_xor1), .fs_or0(h_arrdiv16_fs238_or0));
  fs fs_h_arrdiv16_fs239_out(.a(h_arrdiv16_mux2to1209_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs238_or0[0]), .fs_xor1(h_arrdiv16_fs239_xor1), .fs_or0(h_arrdiv16_fs239_or0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1210_out(.d0(h_arrdiv16_fs224_xor0[0]), .d1(a[1]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1210_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1211_out(.d0(h_arrdiv16_fs225_xor1[0]), .d1(h_arrdiv16_mux2to1195_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1211_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1212_out(.d0(h_arrdiv16_fs226_xor1[0]), .d1(h_arrdiv16_mux2to1196_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1212_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1213_out(.d0(h_arrdiv16_fs227_xor1[0]), .d1(h_arrdiv16_mux2to1197_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1213_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1214_out(.d0(h_arrdiv16_fs228_xor1[0]), .d1(h_arrdiv16_mux2to1198_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1214_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1215_out(.d0(h_arrdiv16_fs229_xor1[0]), .d1(h_arrdiv16_mux2to1199_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1215_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1216_out(.d0(h_arrdiv16_fs230_xor1[0]), .d1(h_arrdiv16_mux2to1200_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1216_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1217_out(.d0(h_arrdiv16_fs231_xor1[0]), .d1(h_arrdiv16_mux2to1201_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1217_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1218_out(.d0(h_arrdiv16_fs232_xor1[0]), .d1(h_arrdiv16_mux2to1202_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1218_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1219_out(.d0(h_arrdiv16_fs233_xor1[0]), .d1(h_arrdiv16_mux2to1203_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1219_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1220_out(.d0(h_arrdiv16_fs234_xor1[0]), .d1(h_arrdiv16_mux2to1204_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1220_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1221_out(.d0(h_arrdiv16_fs235_xor1[0]), .d1(h_arrdiv16_mux2to1205_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1221_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1222_out(.d0(h_arrdiv16_fs236_xor1[0]), .d1(h_arrdiv16_mux2to1206_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1222_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1223_out(.d0(h_arrdiv16_fs237_xor1[0]), .d1(h_arrdiv16_mux2to1207_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1223_xor0));
  mux2to1 mux2to1_h_arrdiv16_mux2to1224_out(.d0(h_arrdiv16_fs238_xor1[0]), .d1(h_arrdiv16_mux2to1208_xor0[0]), .sel(h_arrdiv16_fs239_or0[0]), .mux2to1_xor0(h_arrdiv16_mux2to1224_xor0));
  not_gate not_gate_h_arrdiv16_not14(.a(h_arrdiv16_fs239_or0[0]), .out(h_arrdiv16_not14));
  fs fs_h_arrdiv16_fs240_out(.a(a[0]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv16_fs240_xor0), .fs_or0(h_arrdiv16_fs240_and0));
  fs fs_h_arrdiv16_fs241_out(.a(h_arrdiv16_mux2to1210_xor0[0]), .b(b[1]), .bin(h_arrdiv16_fs240_and0[0]), .fs_xor1(h_arrdiv16_fs241_xor1), .fs_or0(h_arrdiv16_fs241_or0));
  fs fs_h_arrdiv16_fs242_out(.a(h_arrdiv16_mux2to1211_xor0[0]), .b(b[2]), .bin(h_arrdiv16_fs241_or0[0]), .fs_xor1(h_arrdiv16_fs242_xor1), .fs_or0(h_arrdiv16_fs242_or0));
  fs fs_h_arrdiv16_fs243_out(.a(h_arrdiv16_mux2to1212_xor0[0]), .b(b[3]), .bin(h_arrdiv16_fs242_or0[0]), .fs_xor1(h_arrdiv16_fs243_xor1), .fs_or0(h_arrdiv16_fs243_or0));
  fs fs_h_arrdiv16_fs244_out(.a(h_arrdiv16_mux2to1213_xor0[0]), .b(b[4]), .bin(h_arrdiv16_fs243_or0[0]), .fs_xor1(h_arrdiv16_fs244_xor1), .fs_or0(h_arrdiv16_fs244_or0));
  fs fs_h_arrdiv16_fs245_out(.a(h_arrdiv16_mux2to1214_xor0[0]), .b(b[5]), .bin(h_arrdiv16_fs244_or0[0]), .fs_xor1(h_arrdiv16_fs245_xor1), .fs_or0(h_arrdiv16_fs245_or0));
  fs fs_h_arrdiv16_fs246_out(.a(h_arrdiv16_mux2to1215_xor0[0]), .b(b[6]), .bin(h_arrdiv16_fs245_or0[0]), .fs_xor1(h_arrdiv16_fs246_xor1), .fs_or0(h_arrdiv16_fs246_or0));
  fs fs_h_arrdiv16_fs247_out(.a(h_arrdiv16_mux2to1216_xor0[0]), .b(b[7]), .bin(h_arrdiv16_fs246_or0[0]), .fs_xor1(h_arrdiv16_fs247_xor1), .fs_or0(h_arrdiv16_fs247_or0));
  fs fs_h_arrdiv16_fs248_out(.a(h_arrdiv16_mux2to1217_xor0[0]), .b(b[8]), .bin(h_arrdiv16_fs247_or0[0]), .fs_xor1(h_arrdiv16_fs248_xor1), .fs_or0(h_arrdiv16_fs248_or0));
  fs fs_h_arrdiv16_fs249_out(.a(h_arrdiv16_mux2to1218_xor0[0]), .b(b[9]), .bin(h_arrdiv16_fs248_or0[0]), .fs_xor1(h_arrdiv16_fs249_xor1), .fs_or0(h_arrdiv16_fs249_or0));
  fs fs_h_arrdiv16_fs250_out(.a(h_arrdiv16_mux2to1219_xor0[0]), .b(b[10]), .bin(h_arrdiv16_fs249_or0[0]), .fs_xor1(h_arrdiv16_fs250_xor1), .fs_or0(h_arrdiv16_fs250_or0));
  fs fs_h_arrdiv16_fs251_out(.a(h_arrdiv16_mux2to1220_xor0[0]), .b(b[11]), .bin(h_arrdiv16_fs250_or0[0]), .fs_xor1(h_arrdiv16_fs251_xor1), .fs_or0(h_arrdiv16_fs251_or0));
  fs fs_h_arrdiv16_fs252_out(.a(h_arrdiv16_mux2to1221_xor0[0]), .b(b[12]), .bin(h_arrdiv16_fs251_or0[0]), .fs_xor1(h_arrdiv16_fs252_xor1), .fs_or0(h_arrdiv16_fs252_or0));
  fs fs_h_arrdiv16_fs253_out(.a(h_arrdiv16_mux2to1222_xor0[0]), .b(b[13]), .bin(h_arrdiv16_fs252_or0[0]), .fs_xor1(h_arrdiv16_fs253_xor1), .fs_or0(h_arrdiv16_fs253_or0));
  fs fs_h_arrdiv16_fs254_out(.a(h_arrdiv16_mux2to1223_xor0[0]), .b(b[14]), .bin(h_arrdiv16_fs253_or0[0]), .fs_xor1(h_arrdiv16_fs254_xor1), .fs_or0(h_arrdiv16_fs254_or0));
  fs fs_h_arrdiv16_fs255_out(.a(h_arrdiv16_mux2to1224_xor0[0]), .b(b[15]), .bin(h_arrdiv16_fs254_or0[0]), .fs_xor1(h_arrdiv16_fs255_xor1), .fs_or0(h_arrdiv16_fs255_or0));
  not_gate not_gate_h_arrdiv16_not15(.a(h_arrdiv16_fs255_or0[0]), .out(h_arrdiv16_not15));

  assign h_arrdiv16_out[0] = h_arrdiv16_not15[0];
  assign h_arrdiv16_out[1] = h_arrdiv16_not14[0];
  assign h_arrdiv16_out[2] = h_arrdiv16_not13[0];
  assign h_arrdiv16_out[3] = h_arrdiv16_not12[0];
  assign h_arrdiv16_out[4] = h_arrdiv16_not11[0];
  assign h_arrdiv16_out[5] = h_arrdiv16_not10[0];
  assign h_arrdiv16_out[6] = h_arrdiv16_not9[0];
  assign h_arrdiv16_out[7] = h_arrdiv16_not8[0];
  assign h_arrdiv16_out[8] = h_arrdiv16_not7[0];
  assign h_arrdiv16_out[9] = h_arrdiv16_not6[0];
  assign h_arrdiv16_out[10] = h_arrdiv16_not5[0];
  assign h_arrdiv16_out[11] = h_arrdiv16_not4[0];
  assign h_arrdiv16_out[12] = h_arrdiv16_not3[0];
  assign h_arrdiv16_out[13] = h_arrdiv16_not2[0];
  assign h_arrdiv16_out[14] = h_arrdiv16_not1[0];
  assign h_arrdiv16_out[15] = h_arrdiv16_not0[0];
endmodule