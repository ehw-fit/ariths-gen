module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_y0;
  wire fa_y1;
  wire fa_cin;
  wire fa_y3;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module u_rca30(input [29:0] a, input [29:0] b, output [30:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire u_rca30_ha_y0;
  wire u_rca30_ha_y1;
  wire u_rca30_fa1_y2;
  wire u_rca30_fa1_y4;
  wire u_rca30_fa2_y2;
  wire u_rca30_fa2_y4;
  wire u_rca30_fa3_y2;
  wire u_rca30_fa3_y4;
  wire u_rca30_fa4_y2;
  wire u_rca30_fa4_y4;
  wire u_rca30_fa5_y2;
  wire u_rca30_fa5_y4;
  wire u_rca30_fa6_y2;
  wire u_rca30_fa6_y4;
  wire u_rca30_fa7_y2;
  wire u_rca30_fa7_y4;
  wire u_rca30_fa8_y2;
  wire u_rca30_fa8_y4;
  wire u_rca30_fa9_y2;
  wire u_rca30_fa9_y4;
  wire u_rca30_fa10_y2;
  wire u_rca30_fa10_y4;
  wire u_rca30_fa11_y2;
  wire u_rca30_fa11_y4;
  wire u_rca30_fa12_y2;
  wire u_rca30_fa12_y4;
  wire u_rca30_fa13_y2;
  wire u_rca30_fa13_y4;
  wire u_rca30_fa14_y2;
  wire u_rca30_fa14_y4;
  wire u_rca30_fa15_y2;
  wire u_rca30_fa15_y4;
  wire u_rca30_fa16_y2;
  wire u_rca30_fa16_y4;
  wire u_rca30_fa17_y2;
  wire u_rca30_fa17_y4;
  wire u_rca30_fa18_y2;
  wire u_rca30_fa18_y4;
  wire u_rca30_fa19_y2;
  wire u_rca30_fa19_y4;
  wire u_rca30_fa20_y2;
  wire u_rca30_fa20_y4;
  wire u_rca30_fa21_y2;
  wire u_rca30_fa21_y4;
  wire u_rca30_fa22_y2;
  wire u_rca30_fa22_y4;
  wire u_rca30_fa23_y2;
  wire u_rca30_fa23_y4;
  wire u_rca30_fa24_y2;
  wire u_rca30_fa24_y4;
  wire u_rca30_fa25_y2;
  wire u_rca30_fa25_y4;
  wire u_rca30_fa26_y2;
  wire u_rca30_fa26_y4;
  wire u_rca30_fa27_y2;
  wire u_rca30_fa27_y4;
  wire u_rca30_fa28_y2;
  wire u_rca30_fa28_y4;
  wire u_rca30_fa29_y2;
  wire u_rca30_fa29_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  ha ha_u_rca30_ha_y0(a_0, b_0, u_rca30_ha_y0, u_rca30_ha_y1);
  fa fa_u_rca30_fa1_y2(a_1, b_1, u_rca30_ha_y1, u_rca30_fa1_y2, u_rca30_fa1_y4);
  fa fa_u_rca30_fa2_y2(a_2, b_2, u_rca30_fa1_y4, u_rca30_fa2_y2, u_rca30_fa2_y4);
  fa fa_u_rca30_fa3_y2(a_3, b_3, u_rca30_fa2_y4, u_rca30_fa3_y2, u_rca30_fa3_y4);
  fa fa_u_rca30_fa4_y2(a_4, b_4, u_rca30_fa3_y4, u_rca30_fa4_y2, u_rca30_fa4_y4);
  fa fa_u_rca30_fa5_y2(a_5, b_5, u_rca30_fa4_y4, u_rca30_fa5_y2, u_rca30_fa5_y4);
  fa fa_u_rca30_fa6_y2(a_6, b_6, u_rca30_fa5_y4, u_rca30_fa6_y2, u_rca30_fa6_y4);
  fa fa_u_rca30_fa7_y2(a_7, b_7, u_rca30_fa6_y4, u_rca30_fa7_y2, u_rca30_fa7_y4);
  fa fa_u_rca30_fa8_y2(a_8, b_8, u_rca30_fa7_y4, u_rca30_fa8_y2, u_rca30_fa8_y4);
  fa fa_u_rca30_fa9_y2(a_9, b_9, u_rca30_fa8_y4, u_rca30_fa9_y2, u_rca30_fa9_y4);
  fa fa_u_rca30_fa10_y2(a_10, b_10, u_rca30_fa9_y4, u_rca30_fa10_y2, u_rca30_fa10_y4);
  fa fa_u_rca30_fa11_y2(a_11, b_11, u_rca30_fa10_y4, u_rca30_fa11_y2, u_rca30_fa11_y4);
  fa fa_u_rca30_fa12_y2(a_12, b_12, u_rca30_fa11_y4, u_rca30_fa12_y2, u_rca30_fa12_y4);
  fa fa_u_rca30_fa13_y2(a_13, b_13, u_rca30_fa12_y4, u_rca30_fa13_y2, u_rca30_fa13_y4);
  fa fa_u_rca30_fa14_y2(a_14, b_14, u_rca30_fa13_y4, u_rca30_fa14_y2, u_rca30_fa14_y4);
  fa fa_u_rca30_fa15_y2(a_15, b_15, u_rca30_fa14_y4, u_rca30_fa15_y2, u_rca30_fa15_y4);
  fa fa_u_rca30_fa16_y2(a_16, b_16, u_rca30_fa15_y4, u_rca30_fa16_y2, u_rca30_fa16_y4);
  fa fa_u_rca30_fa17_y2(a_17, b_17, u_rca30_fa16_y4, u_rca30_fa17_y2, u_rca30_fa17_y4);
  fa fa_u_rca30_fa18_y2(a_18, b_18, u_rca30_fa17_y4, u_rca30_fa18_y2, u_rca30_fa18_y4);
  fa fa_u_rca30_fa19_y2(a_19, b_19, u_rca30_fa18_y4, u_rca30_fa19_y2, u_rca30_fa19_y4);
  fa fa_u_rca30_fa20_y2(a_20, b_20, u_rca30_fa19_y4, u_rca30_fa20_y2, u_rca30_fa20_y4);
  fa fa_u_rca30_fa21_y2(a_21, b_21, u_rca30_fa20_y4, u_rca30_fa21_y2, u_rca30_fa21_y4);
  fa fa_u_rca30_fa22_y2(a_22, b_22, u_rca30_fa21_y4, u_rca30_fa22_y2, u_rca30_fa22_y4);
  fa fa_u_rca30_fa23_y2(a_23, b_23, u_rca30_fa22_y4, u_rca30_fa23_y2, u_rca30_fa23_y4);
  fa fa_u_rca30_fa24_y2(a_24, b_24, u_rca30_fa23_y4, u_rca30_fa24_y2, u_rca30_fa24_y4);
  fa fa_u_rca30_fa25_y2(a_25, b_25, u_rca30_fa24_y4, u_rca30_fa25_y2, u_rca30_fa25_y4);
  fa fa_u_rca30_fa26_y2(a_26, b_26, u_rca30_fa25_y4, u_rca30_fa26_y2, u_rca30_fa26_y4);
  fa fa_u_rca30_fa27_y2(a_27, b_27, u_rca30_fa26_y4, u_rca30_fa27_y2, u_rca30_fa27_y4);
  fa fa_u_rca30_fa28_y2(a_28, b_28, u_rca30_fa27_y4, u_rca30_fa28_y2, u_rca30_fa28_y4);
  fa fa_u_rca30_fa29_y2(a_29, b_29, u_rca30_fa28_y4, u_rca30_fa29_y2, u_rca30_fa29_y4);

  assign out[0] = u_rca30_ha_y0;
  assign out[1] = u_rca30_fa1_y2;
  assign out[2] = u_rca30_fa2_y2;
  assign out[3] = u_rca30_fa3_y2;
  assign out[4] = u_rca30_fa4_y2;
  assign out[5] = u_rca30_fa5_y2;
  assign out[6] = u_rca30_fa6_y2;
  assign out[7] = u_rca30_fa7_y2;
  assign out[8] = u_rca30_fa8_y2;
  assign out[9] = u_rca30_fa9_y2;
  assign out[10] = u_rca30_fa10_y2;
  assign out[11] = u_rca30_fa11_y2;
  assign out[12] = u_rca30_fa12_y2;
  assign out[13] = u_rca30_fa13_y2;
  assign out[14] = u_rca30_fa14_y2;
  assign out[15] = u_rca30_fa15_y2;
  assign out[16] = u_rca30_fa16_y2;
  assign out[17] = u_rca30_fa17_y2;
  assign out[18] = u_rca30_fa18_y2;
  assign out[19] = u_rca30_fa19_y2;
  assign out[20] = u_rca30_fa20_y2;
  assign out[21] = u_rca30_fa21_y2;
  assign out[22] = u_rca30_fa22_y2;
  assign out[23] = u_rca30_fa23_y2;
  assign out[24] = u_rca30_fa24_y2;
  assign out[25] = u_rca30_fa25_y2;
  assign out[26] = u_rca30_fa26_y2;
  assign out[27] = u_rca30_fa27_y2;
  assign out[28] = u_rca30_fa28_y2;
  assign out[29] = u_rca30_fa29_y2;
  assign out[30] = u_rca30_fa29_y4;
endmodule

module h_u_dadda_rca16(input [15:0] a, input [15:0] b, output [31:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire h_u_dadda_rca16_and_13_0_y0;
  wire h_u_dadda_rca16_and_12_1_y0;
  wire h_u_dadda_rca16_ha0_y0;
  wire h_u_dadda_rca16_ha0_y1;
  wire h_u_dadda_rca16_and_14_0_y0;
  wire h_u_dadda_rca16_and_13_1_y0;
  wire h_u_dadda_rca16_fa0_y2;
  wire h_u_dadda_rca16_fa0_y4;
  wire h_u_dadda_rca16_and_12_2_y0;
  wire h_u_dadda_rca16_and_11_3_y0;
  wire h_u_dadda_rca16_ha1_y0;
  wire h_u_dadda_rca16_ha1_y1;
  wire h_u_dadda_rca16_and_15_0_y0;
  wire h_u_dadda_rca16_fa1_y2;
  wire h_u_dadda_rca16_fa1_y4;
  wire h_u_dadda_rca16_and_14_1_y0;
  wire h_u_dadda_rca16_and_13_2_y0;
  wire h_u_dadda_rca16_and_12_3_y0;
  wire h_u_dadda_rca16_fa2_y2;
  wire h_u_dadda_rca16_fa2_y4;
  wire h_u_dadda_rca16_and_11_4_y0;
  wire h_u_dadda_rca16_and_10_5_y0;
  wire h_u_dadda_rca16_ha2_y0;
  wire h_u_dadda_rca16_ha2_y1;
  wire h_u_dadda_rca16_fa3_y2;
  wire h_u_dadda_rca16_fa3_y4;
  wire h_u_dadda_rca16_and_15_1_y0;
  wire h_u_dadda_rca16_and_14_2_y0;
  wire h_u_dadda_rca16_and_13_3_y0;
  wire h_u_dadda_rca16_fa4_y2;
  wire h_u_dadda_rca16_fa4_y4;
  wire h_u_dadda_rca16_and_12_4_y0;
  wire h_u_dadda_rca16_and_11_5_y0;
  wire h_u_dadda_rca16_ha3_y0;
  wire h_u_dadda_rca16_ha3_y1;
  wire h_u_dadda_rca16_fa5_y2;
  wire h_u_dadda_rca16_fa5_y4;
  wire h_u_dadda_rca16_and_15_2_y0;
  wire h_u_dadda_rca16_and_14_3_y0;
  wire h_u_dadda_rca16_and_13_4_y0;
  wire h_u_dadda_rca16_fa6_y2;
  wire h_u_dadda_rca16_fa6_y4;
  wire h_u_dadda_rca16_and_15_3_y0;
  wire h_u_dadda_rca16_fa7_y2;
  wire h_u_dadda_rca16_fa7_y4;
  wire h_u_dadda_rca16_and_4_0_y0;
  wire h_u_dadda_rca16_and_3_1_y0;
  wire h_u_dadda_rca16_ha4_y0;
  wire h_u_dadda_rca16_ha4_y1;
  wire h_u_dadda_rca16_and_5_0_y0;
  wire h_u_dadda_rca16_and_4_1_y0;
  wire h_u_dadda_rca16_fa8_y2;
  wire h_u_dadda_rca16_fa8_y4;
  wire h_u_dadda_rca16_and_3_2_y0;
  wire h_u_dadda_rca16_and_2_3_y0;
  wire h_u_dadda_rca16_ha5_y0;
  wire h_u_dadda_rca16_ha5_y1;
  wire h_u_dadda_rca16_and_6_0_y0;
  wire h_u_dadda_rca16_fa9_y2;
  wire h_u_dadda_rca16_fa9_y4;
  wire h_u_dadda_rca16_and_5_1_y0;
  wire h_u_dadda_rca16_and_4_2_y0;
  wire h_u_dadda_rca16_and_3_3_y0;
  wire h_u_dadda_rca16_fa10_y2;
  wire h_u_dadda_rca16_fa10_y4;
  wire h_u_dadda_rca16_and_2_4_y0;
  wire h_u_dadda_rca16_and_1_5_y0;
  wire h_u_dadda_rca16_ha6_y0;
  wire h_u_dadda_rca16_ha6_y1;
  wire h_u_dadda_rca16_fa11_y2;
  wire h_u_dadda_rca16_fa11_y4;
  wire h_u_dadda_rca16_and_7_0_y0;
  wire h_u_dadda_rca16_and_6_1_y0;
  wire h_u_dadda_rca16_and_5_2_y0;
  wire h_u_dadda_rca16_fa12_y2;
  wire h_u_dadda_rca16_fa12_y4;
  wire h_u_dadda_rca16_and_4_3_y0;
  wire h_u_dadda_rca16_and_3_4_y0;
  wire h_u_dadda_rca16_and_2_5_y0;
  wire h_u_dadda_rca16_fa13_y2;
  wire h_u_dadda_rca16_fa13_y4;
  wire h_u_dadda_rca16_and_1_6_y0;
  wire h_u_dadda_rca16_and_0_7_y0;
  wire h_u_dadda_rca16_ha7_y0;
  wire h_u_dadda_rca16_ha7_y1;
  wire h_u_dadda_rca16_fa14_y2;
  wire h_u_dadda_rca16_fa14_y4;
  wire h_u_dadda_rca16_and_8_0_y0;
  wire h_u_dadda_rca16_and_7_1_y0;
  wire h_u_dadda_rca16_fa15_y2;
  wire h_u_dadda_rca16_fa15_y4;
  wire h_u_dadda_rca16_and_6_2_y0;
  wire h_u_dadda_rca16_and_5_3_y0;
  wire h_u_dadda_rca16_and_4_4_y0;
  wire h_u_dadda_rca16_fa16_y2;
  wire h_u_dadda_rca16_fa16_y4;
  wire h_u_dadda_rca16_and_3_5_y0;
  wire h_u_dadda_rca16_and_2_6_y0;
  wire h_u_dadda_rca16_and_1_7_y0;
  wire h_u_dadda_rca16_fa17_y2;
  wire h_u_dadda_rca16_fa17_y4;
  wire h_u_dadda_rca16_and_0_8_y0;
  wire h_u_dadda_rca16_ha8_y0;
  wire h_u_dadda_rca16_ha8_y1;
  wire h_u_dadda_rca16_fa18_y2;
  wire h_u_dadda_rca16_fa18_y4;
  wire h_u_dadda_rca16_and_9_0_y0;
  wire h_u_dadda_rca16_fa19_y2;
  wire h_u_dadda_rca16_fa19_y4;
  wire h_u_dadda_rca16_and_8_1_y0;
  wire h_u_dadda_rca16_and_7_2_y0;
  wire h_u_dadda_rca16_and_6_3_y0;
  wire h_u_dadda_rca16_fa20_y2;
  wire h_u_dadda_rca16_fa20_y4;
  wire h_u_dadda_rca16_and_5_4_y0;
  wire h_u_dadda_rca16_and_4_5_y0;
  wire h_u_dadda_rca16_and_3_6_y0;
  wire h_u_dadda_rca16_fa21_y2;
  wire h_u_dadda_rca16_fa21_y4;
  wire h_u_dadda_rca16_and_2_7_y0;
  wire h_u_dadda_rca16_and_1_8_y0;
  wire h_u_dadda_rca16_and_0_9_y0;
  wire h_u_dadda_rca16_fa22_y2;
  wire h_u_dadda_rca16_fa22_y4;
  wire h_u_dadda_rca16_ha9_y0;
  wire h_u_dadda_rca16_ha9_y1;
  wire h_u_dadda_rca16_fa23_y2;
  wire h_u_dadda_rca16_fa23_y4;
  wire h_u_dadda_rca16_fa24_y2;
  wire h_u_dadda_rca16_fa24_y4;
  wire h_u_dadda_rca16_and_10_0_y0;
  wire h_u_dadda_rca16_and_9_1_y0;
  wire h_u_dadda_rca16_and_8_2_y0;
  wire h_u_dadda_rca16_fa25_y2;
  wire h_u_dadda_rca16_fa25_y4;
  wire h_u_dadda_rca16_and_7_3_y0;
  wire h_u_dadda_rca16_and_6_4_y0;
  wire h_u_dadda_rca16_and_5_5_y0;
  wire h_u_dadda_rca16_fa26_y2;
  wire h_u_dadda_rca16_fa26_y4;
  wire h_u_dadda_rca16_and_4_6_y0;
  wire h_u_dadda_rca16_and_3_7_y0;
  wire h_u_dadda_rca16_and_2_8_y0;
  wire h_u_dadda_rca16_fa27_y2;
  wire h_u_dadda_rca16_fa27_y4;
  wire h_u_dadda_rca16_and_1_9_y0;
  wire h_u_dadda_rca16_and_0_10_y0;
  wire h_u_dadda_rca16_fa28_y2;
  wire h_u_dadda_rca16_fa28_y4;
  wire h_u_dadda_rca16_ha10_y0;
  wire h_u_dadda_rca16_ha10_y1;
  wire h_u_dadda_rca16_fa29_y2;
  wire h_u_dadda_rca16_fa29_y4;
  wire h_u_dadda_rca16_fa30_y2;
  wire h_u_dadda_rca16_fa30_y4;
  wire h_u_dadda_rca16_and_11_0_y0;
  wire h_u_dadda_rca16_and_10_1_y0;
  wire h_u_dadda_rca16_fa31_y2;
  wire h_u_dadda_rca16_fa31_y4;
  wire h_u_dadda_rca16_and_9_2_y0;
  wire h_u_dadda_rca16_and_8_3_y0;
  wire h_u_dadda_rca16_and_7_4_y0;
  wire h_u_dadda_rca16_fa32_y2;
  wire h_u_dadda_rca16_fa32_y4;
  wire h_u_dadda_rca16_and_6_5_y0;
  wire h_u_dadda_rca16_and_5_6_y0;
  wire h_u_dadda_rca16_and_4_7_y0;
  wire h_u_dadda_rca16_fa33_y2;
  wire h_u_dadda_rca16_fa33_y4;
  wire h_u_dadda_rca16_and_3_8_y0;
  wire h_u_dadda_rca16_and_2_9_y0;
  wire h_u_dadda_rca16_and_1_10_y0;
  wire h_u_dadda_rca16_fa34_y2;
  wire h_u_dadda_rca16_fa34_y4;
  wire h_u_dadda_rca16_and_0_11_y0;
  wire h_u_dadda_rca16_fa35_y2;
  wire h_u_dadda_rca16_fa35_y4;
  wire h_u_dadda_rca16_ha11_y0;
  wire h_u_dadda_rca16_ha11_y1;
  wire h_u_dadda_rca16_fa36_y2;
  wire h_u_dadda_rca16_fa36_y4;
  wire h_u_dadda_rca16_fa37_y2;
  wire h_u_dadda_rca16_fa37_y4;
  wire h_u_dadda_rca16_and_12_0_y0;
  wire h_u_dadda_rca16_fa38_y2;
  wire h_u_dadda_rca16_fa38_y4;
  wire h_u_dadda_rca16_and_11_1_y0;
  wire h_u_dadda_rca16_and_10_2_y0;
  wire h_u_dadda_rca16_and_9_3_y0;
  wire h_u_dadda_rca16_fa39_y2;
  wire h_u_dadda_rca16_fa39_y4;
  wire h_u_dadda_rca16_and_8_4_y0;
  wire h_u_dadda_rca16_and_7_5_y0;
  wire h_u_dadda_rca16_and_6_6_y0;
  wire h_u_dadda_rca16_fa40_y2;
  wire h_u_dadda_rca16_fa40_y4;
  wire h_u_dadda_rca16_and_5_7_y0;
  wire h_u_dadda_rca16_and_4_8_y0;
  wire h_u_dadda_rca16_and_3_9_y0;
  wire h_u_dadda_rca16_fa41_y2;
  wire h_u_dadda_rca16_fa41_y4;
  wire h_u_dadda_rca16_and_2_10_y0;
  wire h_u_dadda_rca16_and_1_11_y0;
  wire h_u_dadda_rca16_and_0_12_y0;
  wire h_u_dadda_rca16_fa42_y2;
  wire h_u_dadda_rca16_fa42_y4;
  wire h_u_dadda_rca16_fa43_y2;
  wire h_u_dadda_rca16_fa43_y4;
  wire h_u_dadda_rca16_ha12_y0;
  wire h_u_dadda_rca16_ha12_y1;
  wire h_u_dadda_rca16_fa44_y2;
  wire h_u_dadda_rca16_fa44_y4;
  wire h_u_dadda_rca16_fa45_y2;
  wire h_u_dadda_rca16_fa45_y4;
  wire h_u_dadda_rca16_fa46_y2;
  wire h_u_dadda_rca16_fa46_y4;
  wire h_u_dadda_rca16_and_11_2_y0;
  wire h_u_dadda_rca16_and_10_3_y0;
  wire h_u_dadda_rca16_and_9_4_y0;
  wire h_u_dadda_rca16_fa47_y2;
  wire h_u_dadda_rca16_fa47_y4;
  wire h_u_dadda_rca16_and_8_5_y0;
  wire h_u_dadda_rca16_and_7_6_y0;
  wire h_u_dadda_rca16_and_6_7_y0;
  wire h_u_dadda_rca16_fa48_y2;
  wire h_u_dadda_rca16_fa48_y4;
  wire h_u_dadda_rca16_and_5_8_y0;
  wire h_u_dadda_rca16_and_4_9_y0;
  wire h_u_dadda_rca16_and_3_10_y0;
  wire h_u_dadda_rca16_fa49_y2;
  wire h_u_dadda_rca16_fa49_y4;
  wire h_u_dadda_rca16_and_2_11_y0;
  wire h_u_dadda_rca16_and_1_12_y0;
  wire h_u_dadda_rca16_and_0_13_y0;
  wire h_u_dadda_rca16_fa50_y2;
  wire h_u_dadda_rca16_fa50_y4;
  wire h_u_dadda_rca16_fa51_y2;
  wire h_u_dadda_rca16_fa51_y4;
  wire h_u_dadda_rca16_fa52_y2;
  wire h_u_dadda_rca16_fa52_y4;
  wire h_u_dadda_rca16_fa53_y2;
  wire h_u_dadda_rca16_fa53_y4;
  wire h_u_dadda_rca16_fa54_y2;
  wire h_u_dadda_rca16_fa54_y4;
  wire h_u_dadda_rca16_fa55_y2;
  wire h_u_dadda_rca16_fa55_y4;
  wire h_u_dadda_rca16_and_10_4_y0;
  wire h_u_dadda_rca16_and_9_5_y0;
  wire h_u_dadda_rca16_and_8_6_y0;
  wire h_u_dadda_rca16_fa56_y2;
  wire h_u_dadda_rca16_fa56_y4;
  wire h_u_dadda_rca16_and_7_7_y0;
  wire h_u_dadda_rca16_and_6_8_y0;
  wire h_u_dadda_rca16_and_5_9_y0;
  wire h_u_dadda_rca16_fa57_y2;
  wire h_u_dadda_rca16_fa57_y4;
  wire h_u_dadda_rca16_and_4_10_y0;
  wire h_u_dadda_rca16_and_3_11_y0;
  wire h_u_dadda_rca16_and_2_12_y0;
  wire h_u_dadda_rca16_fa58_y2;
  wire h_u_dadda_rca16_fa58_y4;
  wire h_u_dadda_rca16_and_1_13_y0;
  wire h_u_dadda_rca16_and_0_14_y0;
  wire h_u_dadda_rca16_fa59_y2;
  wire h_u_dadda_rca16_fa59_y4;
  wire h_u_dadda_rca16_fa60_y2;
  wire h_u_dadda_rca16_fa60_y4;
  wire h_u_dadda_rca16_fa61_y2;
  wire h_u_dadda_rca16_fa61_y4;
  wire h_u_dadda_rca16_fa62_y2;
  wire h_u_dadda_rca16_fa62_y4;
  wire h_u_dadda_rca16_fa63_y2;
  wire h_u_dadda_rca16_fa63_y4;
  wire h_u_dadda_rca16_fa64_y2;
  wire h_u_dadda_rca16_fa64_y4;
  wire h_u_dadda_rca16_and_9_6_y0;
  wire h_u_dadda_rca16_and_8_7_y0;
  wire h_u_dadda_rca16_and_7_8_y0;
  wire h_u_dadda_rca16_fa65_y2;
  wire h_u_dadda_rca16_fa65_y4;
  wire h_u_dadda_rca16_and_6_9_y0;
  wire h_u_dadda_rca16_and_5_10_y0;
  wire h_u_dadda_rca16_and_4_11_y0;
  wire h_u_dadda_rca16_fa66_y2;
  wire h_u_dadda_rca16_fa66_y4;
  wire h_u_dadda_rca16_and_3_12_y0;
  wire h_u_dadda_rca16_and_2_13_y0;
  wire h_u_dadda_rca16_and_1_14_y0;
  wire h_u_dadda_rca16_fa67_y2;
  wire h_u_dadda_rca16_fa67_y4;
  wire h_u_dadda_rca16_and_0_15_y0;
  wire h_u_dadda_rca16_fa68_y2;
  wire h_u_dadda_rca16_fa68_y4;
  wire h_u_dadda_rca16_fa69_y2;
  wire h_u_dadda_rca16_fa69_y4;
  wire h_u_dadda_rca16_fa70_y2;
  wire h_u_dadda_rca16_fa70_y4;
  wire h_u_dadda_rca16_fa71_y2;
  wire h_u_dadda_rca16_fa71_y4;
  wire h_u_dadda_rca16_fa72_y2;
  wire h_u_dadda_rca16_fa72_y4;
  wire h_u_dadda_rca16_fa73_y2;
  wire h_u_dadda_rca16_fa73_y4;
  wire h_u_dadda_rca16_and_10_6_y0;
  wire h_u_dadda_rca16_and_9_7_y0;
  wire h_u_dadda_rca16_and_8_8_y0;
  wire h_u_dadda_rca16_fa74_y2;
  wire h_u_dadda_rca16_fa74_y4;
  wire h_u_dadda_rca16_and_7_9_y0;
  wire h_u_dadda_rca16_and_6_10_y0;
  wire h_u_dadda_rca16_and_5_11_y0;
  wire h_u_dadda_rca16_fa75_y2;
  wire h_u_dadda_rca16_fa75_y4;
  wire h_u_dadda_rca16_and_4_12_y0;
  wire h_u_dadda_rca16_and_3_13_y0;
  wire h_u_dadda_rca16_and_2_14_y0;
  wire h_u_dadda_rca16_fa76_y2;
  wire h_u_dadda_rca16_fa76_y4;
  wire h_u_dadda_rca16_and_1_15_y0;
  wire h_u_dadda_rca16_fa77_y2;
  wire h_u_dadda_rca16_fa77_y4;
  wire h_u_dadda_rca16_fa78_y2;
  wire h_u_dadda_rca16_fa78_y4;
  wire h_u_dadda_rca16_fa79_y2;
  wire h_u_dadda_rca16_fa79_y4;
  wire h_u_dadda_rca16_fa80_y2;
  wire h_u_dadda_rca16_fa80_y4;
  wire h_u_dadda_rca16_fa81_y2;
  wire h_u_dadda_rca16_fa81_y4;
  wire h_u_dadda_rca16_fa82_y2;
  wire h_u_dadda_rca16_fa82_y4;
  wire h_u_dadda_rca16_and_12_5_y0;
  wire h_u_dadda_rca16_and_11_6_y0;
  wire h_u_dadda_rca16_and_10_7_y0;
  wire h_u_dadda_rca16_fa83_y2;
  wire h_u_dadda_rca16_fa83_y4;
  wire h_u_dadda_rca16_and_9_8_y0;
  wire h_u_dadda_rca16_and_8_9_y0;
  wire h_u_dadda_rca16_and_7_10_y0;
  wire h_u_dadda_rca16_fa84_y2;
  wire h_u_dadda_rca16_fa84_y4;
  wire h_u_dadda_rca16_and_6_11_y0;
  wire h_u_dadda_rca16_and_5_12_y0;
  wire h_u_dadda_rca16_and_4_13_y0;
  wire h_u_dadda_rca16_fa85_y2;
  wire h_u_dadda_rca16_fa85_y4;
  wire h_u_dadda_rca16_and_3_14_y0;
  wire h_u_dadda_rca16_and_2_15_y0;
  wire h_u_dadda_rca16_fa86_y2;
  wire h_u_dadda_rca16_fa86_y4;
  wire h_u_dadda_rca16_fa87_y2;
  wire h_u_dadda_rca16_fa87_y4;
  wire h_u_dadda_rca16_fa88_y2;
  wire h_u_dadda_rca16_fa88_y4;
  wire h_u_dadda_rca16_fa89_y2;
  wire h_u_dadda_rca16_fa89_y4;
  wire h_u_dadda_rca16_fa90_y2;
  wire h_u_dadda_rca16_fa90_y4;
  wire h_u_dadda_rca16_fa91_y2;
  wire h_u_dadda_rca16_fa91_y4;
  wire h_u_dadda_rca16_and_14_4_y0;
  wire h_u_dadda_rca16_and_13_5_y0;
  wire h_u_dadda_rca16_and_12_6_y0;
  wire h_u_dadda_rca16_fa92_y2;
  wire h_u_dadda_rca16_fa92_y4;
  wire h_u_dadda_rca16_and_11_7_y0;
  wire h_u_dadda_rca16_and_10_8_y0;
  wire h_u_dadda_rca16_and_9_9_y0;
  wire h_u_dadda_rca16_fa93_y2;
  wire h_u_dadda_rca16_fa93_y4;
  wire h_u_dadda_rca16_and_8_10_y0;
  wire h_u_dadda_rca16_and_7_11_y0;
  wire h_u_dadda_rca16_and_6_12_y0;
  wire h_u_dadda_rca16_fa94_y2;
  wire h_u_dadda_rca16_fa94_y4;
  wire h_u_dadda_rca16_and_5_13_y0;
  wire h_u_dadda_rca16_and_4_14_y0;
  wire h_u_dadda_rca16_and_3_15_y0;
  wire h_u_dadda_rca16_fa95_y2;
  wire h_u_dadda_rca16_fa95_y4;
  wire h_u_dadda_rca16_fa96_y2;
  wire h_u_dadda_rca16_fa96_y4;
  wire h_u_dadda_rca16_fa97_y2;
  wire h_u_dadda_rca16_fa97_y4;
  wire h_u_dadda_rca16_fa98_y2;
  wire h_u_dadda_rca16_fa98_y4;
  wire h_u_dadda_rca16_fa99_y2;
  wire h_u_dadda_rca16_fa99_y4;
  wire h_u_dadda_rca16_fa100_y2;
  wire h_u_dadda_rca16_fa100_y4;
  wire h_u_dadda_rca16_and_15_4_y0;
  wire h_u_dadda_rca16_and_14_5_y0;
  wire h_u_dadda_rca16_fa101_y2;
  wire h_u_dadda_rca16_fa101_y4;
  wire h_u_dadda_rca16_and_13_6_y0;
  wire h_u_dadda_rca16_and_12_7_y0;
  wire h_u_dadda_rca16_and_11_8_y0;
  wire h_u_dadda_rca16_fa102_y2;
  wire h_u_dadda_rca16_fa102_y4;
  wire h_u_dadda_rca16_and_10_9_y0;
  wire h_u_dadda_rca16_and_9_10_y0;
  wire h_u_dadda_rca16_and_8_11_y0;
  wire h_u_dadda_rca16_fa103_y2;
  wire h_u_dadda_rca16_fa103_y4;
  wire h_u_dadda_rca16_and_7_12_y0;
  wire h_u_dadda_rca16_and_6_13_y0;
  wire h_u_dadda_rca16_and_5_14_y0;
  wire h_u_dadda_rca16_fa104_y2;
  wire h_u_dadda_rca16_fa104_y4;
  wire h_u_dadda_rca16_and_4_15_y0;
  wire h_u_dadda_rca16_fa105_y2;
  wire h_u_dadda_rca16_fa105_y4;
  wire h_u_dadda_rca16_fa106_y2;
  wire h_u_dadda_rca16_fa106_y4;
  wire h_u_dadda_rca16_fa107_y2;
  wire h_u_dadda_rca16_fa107_y4;
  wire h_u_dadda_rca16_fa108_y2;
  wire h_u_dadda_rca16_fa108_y4;
  wire h_u_dadda_rca16_fa109_y2;
  wire h_u_dadda_rca16_fa109_y4;
  wire h_u_dadda_rca16_and_15_5_y0;
  wire h_u_dadda_rca16_and_14_6_y0;
  wire h_u_dadda_rca16_and_13_7_y0;
  wire h_u_dadda_rca16_fa110_y2;
  wire h_u_dadda_rca16_fa110_y4;
  wire h_u_dadda_rca16_and_12_8_y0;
  wire h_u_dadda_rca16_and_11_9_y0;
  wire h_u_dadda_rca16_and_10_10_y0;
  wire h_u_dadda_rca16_fa111_y2;
  wire h_u_dadda_rca16_fa111_y4;
  wire h_u_dadda_rca16_and_9_11_y0;
  wire h_u_dadda_rca16_and_8_12_y0;
  wire h_u_dadda_rca16_and_7_13_y0;
  wire h_u_dadda_rca16_fa112_y2;
  wire h_u_dadda_rca16_fa112_y4;
  wire h_u_dadda_rca16_and_6_14_y0;
  wire h_u_dadda_rca16_and_5_15_y0;
  wire h_u_dadda_rca16_fa113_y2;
  wire h_u_dadda_rca16_fa113_y4;
  wire h_u_dadda_rca16_fa114_y2;
  wire h_u_dadda_rca16_fa114_y4;
  wire h_u_dadda_rca16_fa115_y2;
  wire h_u_dadda_rca16_fa115_y4;
  wire h_u_dadda_rca16_fa116_y2;
  wire h_u_dadda_rca16_fa116_y4;
  wire h_u_dadda_rca16_and_15_6_y0;
  wire h_u_dadda_rca16_fa117_y2;
  wire h_u_dadda_rca16_fa117_y4;
  wire h_u_dadda_rca16_and_14_7_y0;
  wire h_u_dadda_rca16_and_13_8_y0;
  wire h_u_dadda_rca16_and_12_9_y0;
  wire h_u_dadda_rca16_fa118_y2;
  wire h_u_dadda_rca16_fa118_y4;
  wire h_u_dadda_rca16_and_11_10_y0;
  wire h_u_dadda_rca16_and_10_11_y0;
  wire h_u_dadda_rca16_and_9_12_y0;
  wire h_u_dadda_rca16_fa119_y2;
  wire h_u_dadda_rca16_fa119_y4;
  wire h_u_dadda_rca16_and_8_13_y0;
  wire h_u_dadda_rca16_and_7_14_y0;
  wire h_u_dadda_rca16_and_6_15_y0;
  wire h_u_dadda_rca16_fa120_y2;
  wire h_u_dadda_rca16_fa120_y4;
  wire h_u_dadda_rca16_fa121_y2;
  wire h_u_dadda_rca16_fa121_y4;
  wire h_u_dadda_rca16_fa122_y2;
  wire h_u_dadda_rca16_fa122_y4;
  wire h_u_dadda_rca16_fa123_y2;
  wire h_u_dadda_rca16_fa123_y4;
  wire h_u_dadda_rca16_and_15_7_y0;
  wire h_u_dadda_rca16_and_14_8_y0;
  wire h_u_dadda_rca16_fa124_y2;
  wire h_u_dadda_rca16_fa124_y4;
  wire h_u_dadda_rca16_and_13_9_y0;
  wire h_u_dadda_rca16_and_12_10_y0;
  wire h_u_dadda_rca16_and_11_11_y0;
  wire h_u_dadda_rca16_fa125_y2;
  wire h_u_dadda_rca16_fa125_y4;
  wire h_u_dadda_rca16_and_10_12_y0;
  wire h_u_dadda_rca16_and_9_13_y0;
  wire h_u_dadda_rca16_and_8_14_y0;
  wire h_u_dadda_rca16_fa126_y2;
  wire h_u_dadda_rca16_fa126_y4;
  wire h_u_dadda_rca16_and_7_15_y0;
  wire h_u_dadda_rca16_fa127_y2;
  wire h_u_dadda_rca16_fa127_y4;
  wire h_u_dadda_rca16_fa128_y2;
  wire h_u_dadda_rca16_fa128_y4;
  wire h_u_dadda_rca16_fa129_y2;
  wire h_u_dadda_rca16_fa129_y4;
  wire h_u_dadda_rca16_and_15_8_y0;
  wire h_u_dadda_rca16_and_14_9_y0;
  wire h_u_dadda_rca16_and_13_10_y0;
  wire h_u_dadda_rca16_fa130_y2;
  wire h_u_dadda_rca16_fa130_y4;
  wire h_u_dadda_rca16_and_12_11_y0;
  wire h_u_dadda_rca16_and_11_12_y0;
  wire h_u_dadda_rca16_and_10_13_y0;
  wire h_u_dadda_rca16_fa131_y2;
  wire h_u_dadda_rca16_fa131_y4;
  wire h_u_dadda_rca16_and_9_14_y0;
  wire h_u_dadda_rca16_and_8_15_y0;
  wire h_u_dadda_rca16_fa132_y2;
  wire h_u_dadda_rca16_fa132_y4;
  wire h_u_dadda_rca16_fa133_y2;
  wire h_u_dadda_rca16_fa133_y4;
  wire h_u_dadda_rca16_and_15_9_y0;
  wire h_u_dadda_rca16_fa134_y2;
  wire h_u_dadda_rca16_fa134_y4;
  wire h_u_dadda_rca16_and_14_10_y0;
  wire h_u_dadda_rca16_and_13_11_y0;
  wire h_u_dadda_rca16_and_12_12_y0;
  wire h_u_dadda_rca16_fa135_y2;
  wire h_u_dadda_rca16_fa135_y4;
  wire h_u_dadda_rca16_and_11_13_y0;
  wire h_u_dadda_rca16_and_10_14_y0;
  wire h_u_dadda_rca16_and_9_15_y0;
  wire h_u_dadda_rca16_fa136_y2;
  wire h_u_dadda_rca16_fa136_y4;
  wire h_u_dadda_rca16_fa137_y2;
  wire h_u_dadda_rca16_fa137_y4;
  wire h_u_dadda_rca16_and_15_10_y0;
  wire h_u_dadda_rca16_and_14_11_y0;
  wire h_u_dadda_rca16_fa138_y2;
  wire h_u_dadda_rca16_fa138_y4;
  wire h_u_dadda_rca16_and_13_12_y0;
  wire h_u_dadda_rca16_and_12_13_y0;
  wire h_u_dadda_rca16_and_11_14_y0;
  wire h_u_dadda_rca16_fa139_y2;
  wire h_u_dadda_rca16_fa139_y4;
  wire h_u_dadda_rca16_fa140_y2;
  wire h_u_dadda_rca16_fa140_y4;
  wire h_u_dadda_rca16_and_15_11_y0;
  wire h_u_dadda_rca16_and_14_12_y0;
  wire h_u_dadda_rca16_and_13_13_y0;
  wire h_u_dadda_rca16_fa141_y2;
  wire h_u_dadda_rca16_fa141_y4;
  wire h_u_dadda_rca16_and_15_12_y0;
  wire h_u_dadda_rca16_fa142_y2;
  wire h_u_dadda_rca16_fa142_y4;
  wire h_u_dadda_rca16_and_3_0_y0;
  wire h_u_dadda_rca16_and_2_1_y0;
  wire h_u_dadda_rca16_ha13_y0;
  wire h_u_dadda_rca16_ha13_y1;
  wire h_u_dadda_rca16_and_2_2_y0;
  wire h_u_dadda_rca16_and_1_3_y0;
  wire h_u_dadda_rca16_fa143_y2;
  wire h_u_dadda_rca16_fa143_y4;
  wire h_u_dadda_rca16_and_1_4_y0;
  wire h_u_dadda_rca16_and_0_5_y0;
  wire h_u_dadda_rca16_fa144_y2;
  wire h_u_dadda_rca16_fa144_y4;
  wire h_u_dadda_rca16_and_0_6_y0;
  wire h_u_dadda_rca16_fa145_y2;
  wire h_u_dadda_rca16_fa145_y4;
  wire h_u_dadda_rca16_fa146_y2;
  wire h_u_dadda_rca16_fa146_y4;
  wire h_u_dadda_rca16_fa147_y2;
  wire h_u_dadda_rca16_fa147_y4;
  wire h_u_dadda_rca16_fa148_y2;
  wire h_u_dadda_rca16_fa148_y4;
  wire h_u_dadda_rca16_fa149_y2;
  wire h_u_dadda_rca16_fa149_y4;
  wire h_u_dadda_rca16_fa150_y2;
  wire h_u_dadda_rca16_fa150_y4;
  wire h_u_dadda_rca16_fa151_y2;
  wire h_u_dadda_rca16_fa151_y4;
  wire h_u_dadda_rca16_fa152_y2;
  wire h_u_dadda_rca16_fa152_y4;
  wire h_u_dadda_rca16_fa153_y2;
  wire h_u_dadda_rca16_fa153_y4;
  wire h_u_dadda_rca16_fa154_y2;
  wire h_u_dadda_rca16_fa154_y4;
  wire h_u_dadda_rca16_fa155_y2;
  wire h_u_dadda_rca16_fa155_y4;
  wire h_u_dadda_rca16_fa156_y2;
  wire h_u_dadda_rca16_fa156_y4;
  wire h_u_dadda_rca16_fa157_y2;
  wire h_u_dadda_rca16_fa157_y4;
  wire h_u_dadda_rca16_fa158_y2;
  wire h_u_dadda_rca16_fa158_y4;
  wire h_u_dadda_rca16_fa159_y2;
  wire h_u_dadda_rca16_fa159_y4;
  wire h_u_dadda_rca16_fa160_y2;
  wire h_u_dadda_rca16_fa160_y4;
  wire h_u_dadda_rca16_fa161_y2;
  wire h_u_dadda_rca16_fa161_y4;
  wire h_u_dadda_rca16_fa162_y2;
  wire h_u_dadda_rca16_fa162_y4;
  wire h_u_dadda_rca16_fa163_y2;
  wire h_u_dadda_rca16_fa163_y4;
  wire h_u_dadda_rca16_and_10_15_y0;
  wire h_u_dadda_rca16_fa164_y2;
  wire h_u_dadda_rca16_fa164_y4;
  wire h_u_dadda_rca16_and_12_14_y0;
  wire h_u_dadda_rca16_and_11_15_y0;
  wire h_u_dadda_rca16_fa165_y2;
  wire h_u_dadda_rca16_fa165_y4;
  wire h_u_dadda_rca16_and_14_13_y0;
  wire h_u_dadda_rca16_and_13_14_y0;
  wire h_u_dadda_rca16_fa166_y2;
  wire h_u_dadda_rca16_fa166_y4;
  wire h_u_dadda_rca16_and_15_13_y0;
  wire h_u_dadda_rca16_fa167_y2;
  wire h_u_dadda_rca16_fa167_y4;
  wire h_u_dadda_rca16_and_2_0_y0;
  wire h_u_dadda_rca16_and_1_1_y0;
  wire h_u_dadda_rca16_ha14_y0;
  wire h_u_dadda_rca16_ha14_y1;
  wire h_u_dadda_rca16_and_1_2_y0;
  wire h_u_dadda_rca16_and_0_3_y0;
  wire h_u_dadda_rca16_fa168_y2;
  wire h_u_dadda_rca16_fa168_y4;
  wire h_u_dadda_rca16_and_0_4_y0;
  wire h_u_dadda_rca16_fa169_y2;
  wire h_u_dadda_rca16_fa169_y4;
  wire h_u_dadda_rca16_fa170_y2;
  wire h_u_dadda_rca16_fa170_y4;
  wire h_u_dadda_rca16_fa171_y2;
  wire h_u_dadda_rca16_fa171_y4;
  wire h_u_dadda_rca16_fa172_y2;
  wire h_u_dadda_rca16_fa172_y4;
  wire h_u_dadda_rca16_fa173_y2;
  wire h_u_dadda_rca16_fa173_y4;
  wire h_u_dadda_rca16_fa174_y2;
  wire h_u_dadda_rca16_fa174_y4;
  wire h_u_dadda_rca16_fa175_y2;
  wire h_u_dadda_rca16_fa175_y4;
  wire h_u_dadda_rca16_fa176_y2;
  wire h_u_dadda_rca16_fa176_y4;
  wire h_u_dadda_rca16_fa177_y2;
  wire h_u_dadda_rca16_fa177_y4;
  wire h_u_dadda_rca16_fa178_y2;
  wire h_u_dadda_rca16_fa178_y4;
  wire h_u_dadda_rca16_fa179_y2;
  wire h_u_dadda_rca16_fa179_y4;
  wire h_u_dadda_rca16_fa180_y2;
  wire h_u_dadda_rca16_fa180_y4;
  wire h_u_dadda_rca16_fa181_y2;
  wire h_u_dadda_rca16_fa181_y4;
  wire h_u_dadda_rca16_fa182_y2;
  wire h_u_dadda_rca16_fa182_y4;
  wire h_u_dadda_rca16_fa183_y2;
  wire h_u_dadda_rca16_fa183_y4;
  wire h_u_dadda_rca16_fa184_y2;
  wire h_u_dadda_rca16_fa184_y4;
  wire h_u_dadda_rca16_fa185_y2;
  wire h_u_dadda_rca16_fa185_y4;
  wire h_u_dadda_rca16_fa186_y2;
  wire h_u_dadda_rca16_fa186_y4;
  wire h_u_dadda_rca16_fa187_y2;
  wire h_u_dadda_rca16_fa187_y4;
  wire h_u_dadda_rca16_fa188_y2;
  wire h_u_dadda_rca16_fa188_y4;
  wire h_u_dadda_rca16_fa189_y2;
  wire h_u_dadda_rca16_fa189_y4;
  wire h_u_dadda_rca16_fa190_y2;
  wire h_u_dadda_rca16_fa190_y4;
  wire h_u_dadda_rca16_fa191_y2;
  wire h_u_dadda_rca16_fa191_y4;
  wire h_u_dadda_rca16_and_12_15_y0;
  wire h_u_dadda_rca16_fa192_y2;
  wire h_u_dadda_rca16_fa192_y4;
  wire h_u_dadda_rca16_and_14_14_y0;
  wire h_u_dadda_rca16_and_13_15_y0;
  wire h_u_dadda_rca16_fa193_y2;
  wire h_u_dadda_rca16_fa193_y4;
  wire h_u_dadda_rca16_and_15_14_y0;
  wire h_u_dadda_rca16_fa194_y2;
  wire h_u_dadda_rca16_fa194_y4;
  wire h_u_dadda_rca16_and_0_0_y0;
  wire h_u_dadda_rca16_and_1_0_y0;
  wire h_u_dadda_rca16_and_0_2_y0;
  wire h_u_dadda_rca16_and_14_15_y0;
  wire h_u_dadda_rca16_and_0_1_y0;
  wire h_u_dadda_rca16_and_15_15_y0;
  wire [29:0] h_u_dadda_rca16_u_rca30_u_rca30_a;
  wire [29:0] h_u_dadda_rca16_u_rca30_u_rca30_b;
  wire [30:0] h_u_dadda_rca16_u_rca30_out;
  wire h_u_dadda_rca16_u_rca30_ha_y0;
  wire h_u_dadda_rca16_u_rca30_fa1_y2;
  wire h_u_dadda_rca16_u_rca30_fa2_y2;
  wire h_u_dadda_rca16_u_rca30_fa3_y2;
  wire h_u_dadda_rca16_u_rca30_fa4_y2;
  wire h_u_dadda_rca16_u_rca30_fa5_y2;
  wire h_u_dadda_rca16_u_rca30_fa6_y2;
  wire h_u_dadda_rca16_u_rca30_fa7_y2;
  wire h_u_dadda_rca16_u_rca30_fa8_y2;
  wire h_u_dadda_rca16_u_rca30_fa9_y2;
  wire h_u_dadda_rca16_u_rca30_fa10_y2;
  wire h_u_dadda_rca16_u_rca30_fa11_y2;
  wire h_u_dadda_rca16_u_rca30_fa12_y2;
  wire h_u_dadda_rca16_u_rca30_fa13_y2;
  wire h_u_dadda_rca16_u_rca30_fa14_y2;
  wire h_u_dadda_rca16_u_rca30_fa15_y2;
  wire h_u_dadda_rca16_u_rca30_fa16_y2;
  wire h_u_dadda_rca16_u_rca30_fa17_y2;
  wire h_u_dadda_rca16_u_rca30_fa18_y2;
  wire h_u_dadda_rca16_u_rca30_fa19_y2;
  wire h_u_dadda_rca16_u_rca30_fa20_y2;
  wire h_u_dadda_rca16_u_rca30_fa21_y2;
  wire h_u_dadda_rca16_u_rca30_fa22_y2;
  wire h_u_dadda_rca16_u_rca30_fa23_y2;
  wire h_u_dadda_rca16_u_rca30_fa24_y2;
  wire h_u_dadda_rca16_u_rca30_fa25_y2;
  wire h_u_dadda_rca16_u_rca30_fa26_y2;
  wire h_u_dadda_rca16_u_rca30_fa27_y2;
  wire h_u_dadda_rca16_u_rca30_fa28_y2;
  wire h_u_dadda_rca16_u_rca30_fa29_y2;
  wire h_u_dadda_rca16_u_rca30_fa29_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  and_gate and_gate_h_u_dadda_rca16_and_13_0_y0(a_13, b_0, h_u_dadda_rca16_and_13_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_1_y0(a_12, b_1, h_u_dadda_rca16_and_12_1_y0);
  ha ha_h_u_dadda_rca16_ha0_y0(h_u_dadda_rca16_and_13_0_y0, h_u_dadda_rca16_and_12_1_y0, h_u_dadda_rca16_ha0_y0, h_u_dadda_rca16_ha0_y1);
  and_gate and_gate_h_u_dadda_rca16_and_14_0_y0(a_14, b_0, h_u_dadda_rca16_and_14_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_1_y0(a_13, b_1, h_u_dadda_rca16_and_13_1_y0);
  fa fa_h_u_dadda_rca16_fa0_y2(h_u_dadda_rca16_ha0_y1, h_u_dadda_rca16_and_14_0_y0, h_u_dadda_rca16_and_13_1_y0, h_u_dadda_rca16_fa0_y2, h_u_dadda_rca16_fa0_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_2_y0(a_12, b_2, h_u_dadda_rca16_and_12_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_3_y0(a_11, b_3, h_u_dadda_rca16_and_11_3_y0);
  ha ha_h_u_dadda_rca16_ha1_y0(h_u_dadda_rca16_and_12_2_y0, h_u_dadda_rca16_and_11_3_y0, h_u_dadda_rca16_ha1_y0, h_u_dadda_rca16_ha1_y1);
  and_gate and_gate_h_u_dadda_rca16_and_15_0_y0(a_15, b_0, h_u_dadda_rca16_and_15_0_y0);
  fa fa_h_u_dadda_rca16_fa1_y2(h_u_dadda_rca16_ha1_y1, h_u_dadda_rca16_fa0_y4, h_u_dadda_rca16_and_15_0_y0, h_u_dadda_rca16_fa1_y2, h_u_dadda_rca16_fa1_y4);
  and_gate and_gate_h_u_dadda_rca16_and_14_1_y0(a_14, b_1, h_u_dadda_rca16_and_14_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_2_y0(a_13, b_2, h_u_dadda_rca16_and_13_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_3_y0(a_12, b_3, h_u_dadda_rca16_and_12_3_y0);
  fa fa_h_u_dadda_rca16_fa2_y2(h_u_dadda_rca16_and_14_1_y0, h_u_dadda_rca16_and_13_2_y0, h_u_dadda_rca16_and_12_3_y0, h_u_dadda_rca16_fa2_y2, h_u_dadda_rca16_fa2_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_4_y0(a_11, b_4, h_u_dadda_rca16_and_11_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_5_y0(a_10, b_5, h_u_dadda_rca16_and_10_5_y0);
  ha ha_h_u_dadda_rca16_ha2_y0(h_u_dadda_rca16_and_11_4_y0, h_u_dadda_rca16_and_10_5_y0, h_u_dadda_rca16_ha2_y0, h_u_dadda_rca16_ha2_y1);
  fa fa_h_u_dadda_rca16_fa3_y2(h_u_dadda_rca16_ha2_y1, h_u_dadda_rca16_fa2_y4, h_u_dadda_rca16_fa1_y4, h_u_dadda_rca16_fa3_y2, h_u_dadda_rca16_fa3_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_1_y0(a_15, b_1, h_u_dadda_rca16_and_15_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_2_y0(a_14, b_2, h_u_dadda_rca16_and_14_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_3_y0(a_13, b_3, h_u_dadda_rca16_and_13_3_y0);
  fa fa_h_u_dadda_rca16_fa4_y2(h_u_dadda_rca16_and_15_1_y0, h_u_dadda_rca16_and_14_2_y0, h_u_dadda_rca16_and_13_3_y0, h_u_dadda_rca16_fa4_y2, h_u_dadda_rca16_fa4_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_4_y0(a_12, b_4, h_u_dadda_rca16_and_12_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_5_y0(a_11, b_5, h_u_dadda_rca16_and_11_5_y0);
  ha ha_h_u_dadda_rca16_ha3_y0(h_u_dadda_rca16_and_12_4_y0, h_u_dadda_rca16_and_11_5_y0, h_u_dadda_rca16_ha3_y0, h_u_dadda_rca16_ha3_y1);
  fa fa_h_u_dadda_rca16_fa5_y2(h_u_dadda_rca16_ha3_y1, h_u_dadda_rca16_fa4_y4, h_u_dadda_rca16_fa3_y4, h_u_dadda_rca16_fa5_y2, h_u_dadda_rca16_fa5_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_2_y0(a_15, b_2, h_u_dadda_rca16_and_15_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_3_y0(a_14, b_3, h_u_dadda_rca16_and_14_3_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_4_y0(a_13, b_4, h_u_dadda_rca16_and_13_4_y0);
  fa fa_h_u_dadda_rca16_fa6_y2(h_u_dadda_rca16_and_15_2_y0, h_u_dadda_rca16_and_14_3_y0, h_u_dadda_rca16_and_13_4_y0, h_u_dadda_rca16_fa6_y2, h_u_dadda_rca16_fa6_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_3_y0(a_15, b_3, h_u_dadda_rca16_and_15_3_y0);
  fa fa_h_u_dadda_rca16_fa7_y2(h_u_dadda_rca16_fa6_y4, h_u_dadda_rca16_fa5_y4, h_u_dadda_rca16_and_15_3_y0, h_u_dadda_rca16_fa7_y2, h_u_dadda_rca16_fa7_y4);
  and_gate and_gate_h_u_dadda_rca16_and_4_0_y0(a_4, b_0, h_u_dadda_rca16_and_4_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_1_y0(a_3, b_1, h_u_dadda_rca16_and_3_1_y0);
  ha ha_h_u_dadda_rca16_ha4_y0(h_u_dadda_rca16_and_4_0_y0, h_u_dadda_rca16_and_3_1_y0, h_u_dadda_rca16_ha4_y0, h_u_dadda_rca16_ha4_y1);
  and_gate and_gate_h_u_dadda_rca16_and_5_0_y0(a_5, b_0, h_u_dadda_rca16_and_5_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_1_y0(a_4, b_1, h_u_dadda_rca16_and_4_1_y0);
  fa fa_h_u_dadda_rca16_fa8_y2(h_u_dadda_rca16_ha4_y1, h_u_dadda_rca16_and_5_0_y0, h_u_dadda_rca16_and_4_1_y0, h_u_dadda_rca16_fa8_y2, h_u_dadda_rca16_fa8_y4);
  and_gate and_gate_h_u_dadda_rca16_and_3_2_y0(a_3, b_2, h_u_dadda_rca16_and_3_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_3_y0(a_2, b_3, h_u_dadda_rca16_and_2_3_y0);
  ha ha_h_u_dadda_rca16_ha5_y0(h_u_dadda_rca16_and_3_2_y0, h_u_dadda_rca16_and_2_3_y0, h_u_dadda_rca16_ha5_y0, h_u_dadda_rca16_ha5_y1);
  and_gate and_gate_h_u_dadda_rca16_and_6_0_y0(a_6, b_0, h_u_dadda_rca16_and_6_0_y0);
  fa fa_h_u_dadda_rca16_fa9_y2(h_u_dadda_rca16_ha5_y1, h_u_dadda_rca16_fa8_y4, h_u_dadda_rca16_and_6_0_y0, h_u_dadda_rca16_fa9_y2, h_u_dadda_rca16_fa9_y4);
  and_gate and_gate_h_u_dadda_rca16_and_5_1_y0(a_5, b_1, h_u_dadda_rca16_and_5_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_2_y0(a_4, b_2, h_u_dadda_rca16_and_4_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_3_y0(a_3, b_3, h_u_dadda_rca16_and_3_3_y0);
  fa fa_h_u_dadda_rca16_fa10_y2(h_u_dadda_rca16_and_5_1_y0, h_u_dadda_rca16_and_4_2_y0, h_u_dadda_rca16_and_3_3_y0, h_u_dadda_rca16_fa10_y2, h_u_dadda_rca16_fa10_y4);
  and_gate and_gate_h_u_dadda_rca16_and_2_4_y0(a_2, b_4, h_u_dadda_rca16_and_2_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_5_y0(a_1, b_5, h_u_dadda_rca16_and_1_5_y0);
  ha ha_h_u_dadda_rca16_ha6_y0(h_u_dadda_rca16_and_2_4_y0, h_u_dadda_rca16_and_1_5_y0, h_u_dadda_rca16_ha6_y0, h_u_dadda_rca16_ha6_y1);
  fa fa_h_u_dadda_rca16_fa11_y2(h_u_dadda_rca16_ha6_y1, h_u_dadda_rca16_fa10_y4, h_u_dadda_rca16_fa9_y4, h_u_dadda_rca16_fa11_y2, h_u_dadda_rca16_fa11_y4);
  and_gate and_gate_h_u_dadda_rca16_and_7_0_y0(a_7, b_0, h_u_dadda_rca16_and_7_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_1_y0(a_6, b_1, h_u_dadda_rca16_and_6_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_2_y0(a_5, b_2, h_u_dadda_rca16_and_5_2_y0);
  fa fa_h_u_dadda_rca16_fa12_y2(h_u_dadda_rca16_and_7_0_y0, h_u_dadda_rca16_and_6_1_y0, h_u_dadda_rca16_and_5_2_y0, h_u_dadda_rca16_fa12_y2, h_u_dadda_rca16_fa12_y4);
  and_gate and_gate_h_u_dadda_rca16_and_4_3_y0(a_4, b_3, h_u_dadda_rca16_and_4_3_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_4_y0(a_3, b_4, h_u_dadda_rca16_and_3_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_5_y0(a_2, b_5, h_u_dadda_rca16_and_2_5_y0);
  fa fa_h_u_dadda_rca16_fa13_y2(h_u_dadda_rca16_and_4_3_y0, h_u_dadda_rca16_and_3_4_y0, h_u_dadda_rca16_and_2_5_y0, h_u_dadda_rca16_fa13_y2, h_u_dadda_rca16_fa13_y4);
  and_gate and_gate_h_u_dadda_rca16_and_1_6_y0(a_1, b_6, h_u_dadda_rca16_and_1_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_7_y0(a_0, b_7, h_u_dadda_rca16_and_0_7_y0);
  ha ha_h_u_dadda_rca16_ha7_y0(h_u_dadda_rca16_and_1_6_y0, h_u_dadda_rca16_and_0_7_y0, h_u_dadda_rca16_ha7_y0, h_u_dadda_rca16_ha7_y1);
  fa fa_h_u_dadda_rca16_fa14_y2(h_u_dadda_rca16_ha7_y1, h_u_dadda_rca16_fa13_y4, h_u_dadda_rca16_fa12_y4, h_u_dadda_rca16_fa14_y2, h_u_dadda_rca16_fa14_y4);
  and_gate and_gate_h_u_dadda_rca16_and_8_0_y0(a_8, b_0, h_u_dadda_rca16_and_8_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_1_y0(a_7, b_1, h_u_dadda_rca16_and_7_1_y0);
  fa fa_h_u_dadda_rca16_fa15_y2(h_u_dadda_rca16_fa11_y4, h_u_dadda_rca16_and_8_0_y0, h_u_dadda_rca16_and_7_1_y0, h_u_dadda_rca16_fa15_y2, h_u_dadda_rca16_fa15_y4);
  and_gate and_gate_h_u_dadda_rca16_and_6_2_y0(a_6, b_2, h_u_dadda_rca16_and_6_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_3_y0(a_5, b_3, h_u_dadda_rca16_and_5_3_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_4_y0(a_4, b_4, h_u_dadda_rca16_and_4_4_y0);
  fa fa_h_u_dadda_rca16_fa16_y2(h_u_dadda_rca16_and_6_2_y0, h_u_dadda_rca16_and_5_3_y0, h_u_dadda_rca16_and_4_4_y0, h_u_dadda_rca16_fa16_y2, h_u_dadda_rca16_fa16_y4);
  and_gate and_gate_h_u_dadda_rca16_and_3_5_y0(a_3, b_5, h_u_dadda_rca16_and_3_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_6_y0(a_2, b_6, h_u_dadda_rca16_and_2_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_7_y0(a_1, b_7, h_u_dadda_rca16_and_1_7_y0);
  fa fa_h_u_dadda_rca16_fa17_y2(h_u_dadda_rca16_and_3_5_y0, h_u_dadda_rca16_and_2_6_y0, h_u_dadda_rca16_and_1_7_y0, h_u_dadda_rca16_fa17_y2, h_u_dadda_rca16_fa17_y4);
  and_gate and_gate_h_u_dadda_rca16_and_0_8_y0(a_0, b_8, h_u_dadda_rca16_and_0_8_y0);
  ha ha_h_u_dadda_rca16_ha8_y0(h_u_dadda_rca16_and_0_8_y0, h_u_dadda_rca16_fa14_y2, h_u_dadda_rca16_ha8_y0, h_u_dadda_rca16_ha8_y1);
  fa fa_h_u_dadda_rca16_fa18_y2(h_u_dadda_rca16_ha8_y1, h_u_dadda_rca16_fa17_y4, h_u_dadda_rca16_fa16_y4, h_u_dadda_rca16_fa18_y2, h_u_dadda_rca16_fa18_y4);
  and_gate and_gate_h_u_dadda_rca16_and_9_0_y0(a_9, b_0, h_u_dadda_rca16_and_9_0_y0);
  fa fa_h_u_dadda_rca16_fa19_y2(h_u_dadda_rca16_fa15_y4, h_u_dadda_rca16_fa14_y4, h_u_dadda_rca16_and_9_0_y0, h_u_dadda_rca16_fa19_y2, h_u_dadda_rca16_fa19_y4);
  and_gate and_gate_h_u_dadda_rca16_and_8_1_y0(a_8, b_1, h_u_dadda_rca16_and_8_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_2_y0(a_7, b_2, h_u_dadda_rca16_and_7_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_3_y0(a_6, b_3, h_u_dadda_rca16_and_6_3_y0);
  fa fa_h_u_dadda_rca16_fa20_y2(h_u_dadda_rca16_and_8_1_y0, h_u_dadda_rca16_and_7_2_y0, h_u_dadda_rca16_and_6_3_y0, h_u_dadda_rca16_fa20_y2, h_u_dadda_rca16_fa20_y4);
  and_gate and_gate_h_u_dadda_rca16_and_5_4_y0(a_5, b_4, h_u_dadda_rca16_and_5_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_5_y0(a_4, b_5, h_u_dadda_rca16_and_4_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_6_y0(a_3, b_6, h_u_dadda_rca16_and_3_6_y0);
  fa fa_h_u_dadda_rca16_fa21_y2(h_u_dadda_rca16_and_5_4_y0, h_u_dadda_rca16_and_4_5_y0, h_u_dadda_rca16_and_3_6_y0, h_u_dadda_rca16_fa21_y2, h_u_dadda_rca16_fa21_y4);
  and_gate and_gate_h_u_dadda_rca16_and_2_7_y0(a_2, b_7, h_u_dadda_rca16_and_2_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_8_y0(a_1, b_8, h_u_dadda_rca16_and_1_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_9_y0(a_0, b_9, h_u_dadda_rca16_and_0_9_y0);
  fa fa_h_u_dadda_rca16_fa22_y2(h_u_dadda_rca16_and_2_7_y0, h_u_dadda_rca16_and_1_8_y0, h_u_dadda_rca16_and_0_9_y0, h_u_dadda_rca16_fa22_y2, h_u_dadda_rca16_fa22_y4);
  ha ha_h_u_dadda_rca16_ha9_y0(h_u_dadda_rca16_fa18_y2, h_u_dadda_rca16_fa19_y2, h_u_dadda_rca16_ha9_y0, h_u_dadda_rca16_ha9_y1);
  fa fa_h_u_dadda_rca16_fa23_y2(h_u_dadda_rca16_ha9_y1, h_u_dadda_rca16_fa22_y4, h_u_dadda_rca16_fa21_y4, h_u_dadda_rca16_fa23_y2, h_u_dadda_rca16_fa23_y4);
  fa fa_h_u_dadda_rca16_fa24_y2(h_u_dadda_rca16_fa20_y4, h_u_dadda_rca16_fa19_y4, h_u_dadda_rca16_fa18_y4, h_u_dadda_rca16_fa24_y2, h_u_dadda_rca16_fa24_y4);
  and_gate and_gate_h_u_dadda_rca16_and_10_0_y0(a_10, b_0, h_u_dadda_rca16_and_10_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_1_y0(a_9, b_1, h_u_dadda_rca16_and_9_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_2_y0(a_8, b_2, h_u_dadda_rca16_and_8_2_y0);
  fa fa_h_u_dadda_rca16_fa25_y2(h_u_dadda_rca16_and_10_0_y0, h_u_dadda_rca16_and_9_1_y0, h_u_dadda_rca16_and_8_2_y0, h_u_dadda_rca16_fa25_y2, h_u_dadda_rca16_fa25_y4);
  and_gate and_gate_h_u_dadda_rca16_and_7_3_y0(a_7, b_3, h_u_dadda_rca16_and_7_3_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_4_y0(a_6, b_4, h_u_dadda_rca16_and_6_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_5_y0(a_5, b_5, h_u_dadda_rca16_and_5_5_y0);
  fa fa_h_u_dadda_rca16_fa26_y2(h_u_dadda_rca16_and_7_3_y0, h_u_dadda_rca16_and_6_4_y0, h_u_dadda_rca16_and_5_5_y0, h_u_dadda_rca16_fa26_y2, h_u_dadda_rca16_fa26_y4);
  and_gate and_gate_h_u_dadda_rca16_and_4_6_y0(a_4, b_6, h_u_dadda_rca16_and_4_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_7_y0(a_3, b_7, h_u_dadda_rca16_and_3_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_8_y0(a_2, b_8, h_u_dadda_rca16_and_2_8_y0);
  fa fa_h_u_dadda_rca16_fa27_y2(h_u_dadda_rca16_and_4_6_y0, h_u_dadda_rca16_and_3_7_y0, h_u_dadda_rca16_and_2_8_y0, h_u_dadda_rca16_fa27_y2, h_u_dadda_rca16_fa27_y4);
  and_gate and_gate_h_u_dadda_rca16_and_1_9_y0(a_1, b_9, h_u_dadda_rca16_and_1_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_10_y0(a_0, b_10, h_u_dadda_rca16_and_0_10_y0);
  fa fa_h_u_dadda_rca16_fa28_y2(h_u_dadda_rca16_and_1_9_y0, h_u_dadda_rca16_and_0_10_y0, h_u_dadda_rca16_fa23_y2, h_u_dadda_rca16_fa28_y2, h_u_dadda_rca16_fa28_y4);
  ha ha_h_u_dadda_rca16_ha10_y0(h_u_dadda_rca16_fa24_y2, h_u_dadda_rca16_fa25_y2, h_u_dadda_rca16_ha10_y0, h_u_dadda_rca16_ha10_y1);
  fa fa_h_u_dadda_rca16_fa29_y2(h_u_dadda_rca16_ha10_y1, h_u_dadda_rca16_fa28_y4, h_u_dadda_rca16_fa27_y4, h_u_dadda_rca16_fa29_y2, h_u_dadda_rca16_fa29_y4);
  fa fa_h_u_dadda_rca16_fa30_y2(h_u_dadda_rca16_fa26_y4, h_u_dadda_rca16_fa25_y4, h_u_dadda_rca16_fa24_y4, h_u_dadda_rca16_fa30_y2, h_u_dadda_rca16_fa30_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_0_y0(a_11, b_0, h_u_dadda_rca16_and_11_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_1_y0(a_10, b_1, h_u_dadda_rca16_and_10_1_y0);
  fa fa_h_u_dadda_rca16_fa31_y2(h_u_dadda_rca16_fa23_y4, h_u_dadda_rca16_and_11_0_y0, h_u_dadda_rca16_and_10_1_y0, h_u_dadda_rca16_fa31_y2, h_u_dadda_rca16_fa31_y4);
  and_gate and_gate_h_u_dadda_rca16_and_9_2_y0(a_9, b_2, h_u_dadda_rca16_and_9_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_3_y0(a_8, b_3, h_u_dadda_rca16_and_8_3_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_4_y0(a_7, b_4, h_u_dadda_rca16_and_7_4_y0);
  fa fa_h_u_dadda_rca16_fa32_y2(h_u_dadda_rca16_and_9_2_y0, h_u_dadda_rca16_and_8_3_y0, h_u_dadda_rca16_and_7_4_y0, h_u_dadda_rca16_fa32_y2, h_u_dadda_rca16_fa32_y4);
  and_gate and_gate_h_u_dadda_rca16_and_6_5_y0(a_6, b_5, h_u_dadda_rca16_and_6_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_6_y0(a_5, b_6, h_u_dadda_rca16_and_5_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_7_y0(a_4, b_7, h_u_dadda_rca16_and_4_7_y0);
  fa fa_h_u_dadda_rca16_fa33_y2(h_u_dadda_rca16_and_6_5_y0, h_u_dadda_rca16_and_5_6_y0, h_u_dadda_rca16_and_4_7_y0, h_u_dadda_rca16_fa33_y2, h_u_dadda_rca16_fa33_y4);
  and_gate and_gate_h_u_dadda_rca16_and_3_8_y0(a_3, b_8, h_u_dadda_rca16_and_3_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_9_y0(a_2, b_9, h_u_dadda_rca16_and_2_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_10_y0(a_1, b_10, h_u_dadda_rca16_and_1_10_y0);
  fa fa_h_u_dadda_rca16_fa34_y2(h_u_dadda_rca16_and_3_8_y0, h_u_dadda_rca16_and_2_9_y0, h_u_dadda_rca16_and_1_10_y0, h_u_dadda_rca16_fa34_y2, h_u_dadda_rca16_fa34_y4);
  and_gate and_gate_h_u_dadda_rca16_and_0_11_y0(a_0, b_11, h_u_dadda_rca16_and_0_11_y0);
  fa fa_h_u_dadda_rca16_fa35_y2(h_u_dadda_rca16_and_0_11_y0, h_u_dadda_rca16_fa29_y2, h_u_dadda_rca16_fa30_y2, h_u_dadda_rca16_fa35_y2, h_u_dadda_rca16_fa35_y4);
  ha ha_h_u_dadda_rca16_ha11_y0(h_u_dadda_rca16_fa31_y2, h_u_dadda_rca16_fa32_y2, h_u_dadda_rca16_ha11_y0, h_u_dadda_rca16_ha11_y1);
  fa fa_h_u_dadda_rca16_fa36_y2(h_u_dadda_rca16_ha11_y1, h_u_dadda_rca16_fa35_y4, h_u_dadda_rca16_fa34_y4, h_u_dadda_rca16_fa36_y2, h_u_dadda_rca16_fa36_y4);
  fa fa_h_u_dadda_rca16_fa37_y2(h_u_dadda_rca16_fa33_y4, h_u_dadda_rca16_fa32_y4, h_u_dadda_rca16_fa31_y4, h_u_dadda_rca16_fa37_y2, h_u_dadda_rca16_fa37_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_0_y0(a_12, b_0, h_u_dadda_rca16_and_12_0_y0);
  fa fa_h_u_dadda_rca16_fa38_y2(h_u_dadda_rca16_fa30_y4, h_u_dadda_rca16_fa29_y4, h_u_dadda_rca16_and_12_0_y0, h_u_dadda_rca16_fa38_y2, h_u_dadda_rca16_fa38_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_1_y0(a_11, b_1, h_u_dadda_rca16_and_11_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_2_y0(a_10, b_2, h_u_dadda_rca16_and_10_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_3_y0(a_9, b_3, h_u_dadda_rca16_and_9_3_y0);
  fa fa_h_u_dadda_rca16_fa39_y2(h_u_dadda_rca16_and_11_1_y0, h_u_dadda_rca16_and_10_2_y0, h_u_dadda_rca16_and_9_3_y0, h_u_dadda_rca16_fa39_y2, h_u_dadda_rca16_fa39_y4);
  and_gate and_gate_h_u_dadda_rca16_and_8_4_y0(a_8, b_4, h_u_dadda_rca16_and_8_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_5_y0(a_7, b_5, h_u_dadda_rca16_and_7_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_6_y0(a_6, b_6, h_u_dadda_rca16_and_6_6_y0);
  fa fa_h_u_dadda_rca16_fa40_y2(h_u_dadda_rca16_and_8_4_y0, h_u_dadda_rca16_and_7_5_y0, h_u_dadda_rca16_and_6_6_y0, h_u_dadda_rca16_fa40_y2, h_u_dadda_rca16_fa40_y4);
  and_gate and_gate_h_u_dadda_rca16_and_5_7_y0(a_5, b_7, h_u_dadda_rca16_and_5_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_8_y0(a_4, b_8, h_u_dadda_rca16_and_4_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_9_y0(a_3, b_9, h_u_dadda_rca16_and_3_9_y0);
  fa fa_h_u_dadda_rca16_fa41_y2(h_u_dadda_rca16_and_5_7_y0, h_u_dadda_rca16_and_4_8_y0, h_u_dadda_rca16_and_3_9_y0, h_u_dadda_rca16_fa41_y2, h_u_dadda_rca16_fa41_y4);
  and_gate and_gate_h_u_dadda_rca16_and_2_10_y0(a_2, b_10, h_u_dadda_rca16_and_2_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_11_y0(a_1, b_11, h_u_dadda_rca16_and_1_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_12_y0(a_0, b_12, h_u_dadda_rca16_and_0_12_y0);
  fa fa_h_u_dadda_rca16_fa42_y2(h_u_dadda_rca16_and_2_10_y0, h_u_dadda_rca16_and_1_11_y0, h_u_dadda_rca16_and_0_12_y0, h_u_dadda_rca16_fa42_y2, h_u_dadda_rca16_fa42_y4);
  fa fa_h_u_dadda_rca16_fa43_y2(h_u_dadda_rca16_fa36_y2, h_u_dadda_rca16_fa37_y2, h_u_dadda_rca16_fa38_y2, h_u_dadda_rca16_fa43_y2, h_u_dadda_rca16_fa43_y4);
  ha ha_h_u_dadda_rca16_ha12_y0(h_u_dadda_rca16_fa39_y2, h_u_dadda_rca16_fa40_y2, h_u_dadda_rca16_ha12_y0, h_u_dadda_rca16_ha12_y1);
  fa fa_h_u_dadda_rca16_fa44_y2(h_u_dadda_rca16_ha12_y1, h_u_dadda_rca16_fa43_y4, h_u_dadda_rca16_fa42_y4, h_u_dadda_rca16_fa44_y2, h_u_dadda_rca16_fa44_y4);
  fa fa_h_u_dadda_rca16_fa45_y2(h_u_dadda_rca16_fa41_y4, h_u_dadda_rca16_fa40_y4, h_u_dadda_rca16_fa39_y4, h_u_dadda_rca16_fa45_y2, h_u_dadda_rca16_fa45_y4);
  fa fa_h_u_dadda_rca16_fa46_y2(h_u_dadda_rca16_fa38_y4, h_u_dadda_rca16_fa37_y4, h_u_dadda_rca16_fa36_y4, h_u_dadda_rca16_fa46_y2, h_u_dadda_rca16_fa46_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_2_y0(a_11, b_2, h_u_dadda_rca16_and_11_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_3_y0(a_10, b_3, h_u_dadda_rca16_and_10_3_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_4_y0(a_9, b_4, h_u_dadda_rca16_and_9_4_y0);
  fa fa_h_u_dadda_rca16_fa47_y2(h_u_dadda_rca16_and_11_2_y0, h_u_dadda_rca16_and_10_3_y0, h_u_dadda_rca16_and_9_4_y0, h_u_dadda_rca16_fa47_y2, h_u_dadda_rca16_fa47_y4);
  and_gate and_gate_h_u_dadda_rca16_and_8_5_y0(a_8, b_5, h_u_dadda_rca16_and_8_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_6_y0(a_7, b_6, h_u_dadda_rca16_and_7_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_7_y0(a_6, b_7, h_u_dadda_rca16_and_6_7_y0);
  fa fa_h_u_dadda_rca16_fa48_y2(h_u_dadda_rca16_and_8_5_y0, h_u_dadda_rca16_and_7_6_y0, h_u_dadda_rca16_and_6_7_y0, h_u_dadda_rca16_fa48_y2, h_u_dadda_rca16_fa48_y4);
  and_gate and_gate_h_u_dadda_rca16_and_5_8_y0(a_5, b_8, h_u_dadda_rca16_and_5_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_9_y0(a_4, b_9, h_u_dadda_rca16_and_4_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_10_y0(a_3, b_10, h_u_dadda_rca16_and_3_10_y0);
  fa fa_h_u_dadda_rca16_fa49_y2(h_u_dadda_rca16_and_5_8_y0, h_u_dadda_rca16_and_4_9_y0, h_u_dadda_rca16_and_3_10_y0, h_u_dadda_rca16_fa49_y2, h_u_dadda_rca16_fa49_y4);
  and_gate and_gate_h_u_dadda_rca16_and_2_11_y0(a_2, b_11, h_u_dadda_rca16_and_2_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_12_y0(a_1, b_12, h_u_dadda_rca16_and_1_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_13_y0(a_0, b_13, h_u_dadda_rca16_and_0_13_y0);
  fa fa_h_u_dadda_rca16_fa50_y2(h_u_dadda_rca16_and_2_11_y0, h_u_dadda_rca16_and_1_12_y0, h_u_dadda_rca16_and_0_13_y0, h_u_dadda_rca16_fa50_y2, h_u_dadda_rca16_fa50_y4);
  fa fa_h_u_dadda_rca16_fa51_y2(h_u_dadda_rca16_ha0_y0, h_u_dadda_rca16_fa44_y2, h_u_dadda_rca16_fa45_y2, h_u_dadda_rca16_fa51_y2, h_u_dadda_rca16_fa51_y4);
  fa fa_h_u_dadda_rca16_fa52_y2(h_u_dadda_rca16_fa46_y2, h_u_dadda_rca16_fa47_y2, h_u_dadda_rca16_fa48_y2, h_u_dadda_rca16_fa52_y2, h_u_dadda_rca16_fa52_y4);
  fa fa_h_u_dadda_rca16_fa53_y2(h_u_dadda_rca16_fa52_y4, h_u_dadda_rca16_fa51_y4, h_u_dadda_rca16_fa50_y4, h_u_dadda_rca16_fa53_y2, h_u_dadda_rca16_fa53_y4);
  fa fa_h_u_dadda_rca16_fa54_y2(h_u_dadda_rca16_fa49_y4, h_u_dadda_rca16_fa48_y4, h_u_dadda_rca16_fa47_y4, h_u_dadda_rca16_fa54_y2, h_u_dadda_rca16_fa54_y4);
  fa fa_h_u_dadda_rca16_fa55_y2(h_u_dadda_rca16_fa46_y4, h_u_dadda_rca16_fa45_y4, h_u_dadda_rca16_fa44_y4, h_u_dadda_rca16_fa55_y2, h_u_dadda_rca16_fa55_y4);
  and_gate and_gate_h_u_dadda_rca16_and_10_4_y0(a_10, b_4, h_u_dadda_rca16_and_10_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_5_y0(a_9, b_5, h_u_dadda_rca16_and_9_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_6_y0(a_8, b_6, h_u_dadda_rca16_and_8_6_y0);
  fa fa_h_u_dadda_rca16_fa56_y2(h_u_dadda_rca16_and_10_4_y0, h_u_dadda_rca16_and_9_5_y0, h_u_dadda_rca16_and_8_6_y0, h_u_dadda_rca16_fa56_y2, h_u_dadda_rca16_fa56_y4);
  and_gate and_gate_h_u_dadda_rca16_and_7_7_y0(a_7, b_7, h_u_dadda_rca16_and_7_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_8_y0(a_6, b_8, h_u_dadda_rca16_and_6_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_9_y0(a_5, b_9, h_u_dadda_rca16_and_5_9_y0);
  fa fa_h_u_dadda_rca16_fa57_y2(h_u_dadda_rca16_and_7_7_y0, h_u_dadda_rca16_and_6_8_y0, h_u_dadda_rca16_and_5_9_y0, h_u_dadda_rca16_fa57_y2, h_u_dadda_rca16_fa57_y4);
  and_gate and_gate_h_u_dadda_rca16_and_4_10_y0(a_4, b_10, h_u_dadda_rca16_and_4_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_11_y0(a_3, b_11, h_u_dadda_rca16_and_3_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_12_y0(a_2, b_12, h_u_dadda_rca16_and_2_12_y0);
  fa fa_h_u_dadda_rca16_fa58_y2(h_u_dadda_rca16_and_4_10_y0, h_u_dadda_rca16_and_3_11_y0, h_u_dadda_rca16_and_2_12_y0, h_u_dadda_rca16_fa58_y2, h_u_dadda_rca16_fa58_y4);
  and_gate and_gate_h_u_dadda_rca16_and_1_13_y0(a_1, b_13, h_u_dadda_rca16_and_1_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_14_y0(a_0, b_14, h_u_dadda_rca16_and_0_14_y0);
  fa fa_h_u_dadda_rca16_fa59_y2(h_u_dadda_rca16_and_1_13_y0, h_u_dadda_rca16_and_0_14_y0, h_u_dadda_rca16_fa0_y2, h_u_dadda_rca16_fa59_y2, h_u_dadda_rca16_fa59_y4);
  fa fa_h_u_dadda_rca16_fa60_y2(h_u_dadda_rca16_ha1_y0, h_u_dadda_rca16_fa53_y2, h_u_dadda_rca16_fa54_y2, h_u_dadda_rca16_fa60_y2, h_u_dadda_rca16_fa60_y4);
  fa fa_h_u_dadda_rca16_fa61_y2(h_u_dadda_rca16_fa55_y2, h_u_dadda_rca16_fa56_y2, h_u_dadda_rca16_fa57_y2, h_u_dadda_rca16_fa61_y2, h_u_dadda_rca16_fa61_y4);
  fa fa_h_u_dadda_rca16_fa62_y2(h_u_dadda_rca16_fa61_y4, h_u_dadda_rca16_fa60_y4, h_u_dadda_rca16_fa59_y4, h_u_dadda_rca16_fa62_y2, h_u_dadda_rca16_fa62_y4);
  fa fa_h_u_dadda_rca16_fa63_y2(h_u_dadda_rca16_fa58_y4, h_u_dadda_rca16_fa57_y4, h_u_dadda_rca16_fa56_y4, h_u_dadda_rca16_fa63_y2, h_u_dadda_rca16_fa63_y4);
  fa fa_h_u_dadda_rca16_fa64_y2(h_u_dadda_rca16_fa55_y4, h_u_dadda_rca16_fa54_y4, h_u_dadda_rca16_fa53_y4, h_u_dadda_rca16_fa64_y2, h_u_dadda_rca16_fa64_y4);
  and_gate and_gate_h_u_dadda_rca16_and_9_6_y0(a_9, b_6, h_u_dadda_rca16_and_9_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_7_y0(a_8, b_7, h_u_dadda_rca16_and_8_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_8_y0(a_7, b_8, h_u_dadda_rca16_and_7_8_y0);
  fa fa_h_u_dadda_rca16_fa65_y2(h_u_dadda_rca16_and_9_6_y0, h_u_dadda_rca16_and_8_7_y0, h_u_dadda_rca16_and_7_8_y0, h_u_dadda_rca16_fa65_y2, h_u_dadda_rca16_fa65_y4);
  and_gate and_gate_h_u_dadda_rca16_and_6_9_y0(a_6, b_9, h_u_dadda_rca16_and_6_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_10_y0(a_5, b_10, h_u_dadda_rca16_and_5_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_11_y0(a_4, b_11, h_u_dadda_rca16_and_4_11_y0);
  fa fa_h_u_dadda_rca16_fa66_y2(h_u_dadda_rca16_and_6_9_y0, h_u_dadda_rca16_and_5_10_y0, h_u_dadda_rca16_and_4_11_y0, h_u_dadda_rca16_fa66_y2, h_u_dadda_rca16_fa66_y4);
  and_gate and_gate_h_u_dadda_rca16_and_3_12_y0(a_3, b_12, h_u_dadda_rca16_and_3_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_13_y0(a_2, b_13, h_u_dadda_rca16_and_2_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_14_y0(a_1, b_14, h_u_dadda_rca16_and_1_14_y0);
  fa fa_h_u_dadda_rca16_fa67_y2(h_u_dadda_rca16_and_3_12_y0, h_u_dadda_rca16_and_2_13_y0, h_u_dadda_rca16_and_1_14_y0, h_u_dadda_rca16_fa67_y2, h_u_dadda_rca16_fa67_y4);
  and_gate and_gate_h_u_dadda_rca16_and_0_15_y0(a_0, b_15, h_u_dadda_rca16_and_0_15_y0);
  fa fa_h_u_dadda_rca16_fa68_y2(h_u_dadda_rca16_and_0_15_y0, h_u_dadda_rca16_fa1_y2, h_u_dadda_rca16_fa2_y2, h_u_dadda_rca16_fa68_y2, h_u_dadda_rca16_fa68_y4);
  fa fa_h_u_dadda_rca16_fa69_y2(h_u_dadda_rca16_ha2_y0, h_u_dadda_rca16_fa62_y2, h_u_dadda_rca16_fa63_y2, h_u_dadda_rca16_fa69_y2, h_u_dadda_rca16_fa69_y4);
  fa fa_h_u_dadda_rca16_fa70_y2(h_u_dadda_rca16_fa64_y2, h_u_dadda_rca16_fa65_y2, h_u_dadda_rca16_fa66_y2, h_u_dadda_rca16_fa70_y2, h_u_dadda_rca16_fa70_y4);
  fa fa_h_u_dadda_rca16_fa71_y2(h_u_dadda_rca16_fa70_y4, h_u_dadda_rca16_fa69_y4, h_u_dadda_rca16_fa68_y4, h_u_dadda_rca16_fa71_y2, h_u_dadda_rca16_fa71_y4);
  fa fa_h_u_dadda_rca16_fa72_y2(h_u_dadda_rca16_fa67_y4, h_u_dadda_rca16_fa66_y4, h_u_dadda_rca16_fa65_y4, h_u_dadda_rca16_fa72_y2, h_u_dadda_rca16_fa72_y4);
  fa fa_h_u_dadda_rca16_fa73_y2(h_u_dadda_rca16_fa64_y4, h_u_dadda_rca16_fa63_y4, h_u_dadda_rca16_fa62_y4, h_u_dadda_rca16_fa73_y2, h_u_dadda_rca16_fa73_y4);
  and_gate and_gate_h_u_dadda_rca16_and_10_6_y0(a_10, b_6, h_u_dadda_rca16_and_10_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_7_y0(a_9, b_7, h_u_dadda_rca16_and_9_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_8_y0(a_8, b_8, h_u_dadda_rca16_and_8_8_y0);
  fa fa_h_u_dadda_rca16_fa74_y2(h_u_dadda_rca16_and_10_6_y0, h_u_dadda_rca16_and_9_7_y0, h_u_dadda_rca16_and_8_8_y0, h_u_dadda_rca16_fa74_y2, h_u_dadda_rca16_fa74_y4);
  and_gate and_gate_h_u_dadda_rca16_and_7_9_y0(a_7, b_9, h_u_dadda_rca16_and_7_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_10_y0(a_6, b_10, h_u_dadda_rca16_and_6_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_11_y0(a_5, b_11, h_u_dadda_rca16_and_5_11_y0);
  fa fa_h_u_dadda_rca16_fa75_y2(h_u_dadda_rca16_and_7_9_y0, h_u_dadda_rca16_and_6_10_y0, h_u_dadda_rca16_and_5_11_y0, h_u_dadda_rca16_fa75_y2, h_u_dadda_rca16_fa75_y4);
  and_gate and_gate_h_u_dadda_rca16_and_4_12_y0(a_4, b_12, h_u_dadda_rca16_and_4_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_13_y0(a_3, b_13, h_u_dadda_rca16_and_3_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_14_y0(a_2, b_14, h_u_dadda_rca16_and_2_14_y0);
  fa fa_h_u_dadda_rca16_fa76_y2(h_u_dadda_rca16_and_4_12_y0, h_u_dadda_rca16_and_3_13_y0, h_u_dadda_rca16_and_2_14_y0, h_u_dadda_rca16_fa76_y2, h_u_dadda_rca16_fa76_y4);
  and_gate and_gate_h_u_dadda_rca16_and_1_15_y0(a_1, b_15, h_u_dadda_rca16_and_1_15_y0);
  fa fa_h_u_dadda_rca16_fa77_y2(h_u_dadda_rca16_and_1_15_y0, h_u_dadda_rca16_fa3_y2, h_u_dadda_rca16_fa4_y2, h_u_dadda_rca16_fa77_y2, h_u_dadda_rca16_fa77_y4);
  fa fa_h_u_dadda_rca16_fa78_y2(h_u_dadda_rca16_ha3_y0, h_u_dadda_rca16_fa71_y2, h_u_dadda_rca16_fa72_y2, h_u_dadda_rca16_fa78_y2, h_u_dadda_rca16_fa78_y4);
  fa fa_h_u_dadda_rca16_fa79_y2(h_u_dadda_rca16_fa73_y2, h_u_dadda_rca16_fa74_y2, h_u_dadda_rca16_fa75_y2, h_u_dadda_rca16_fa79_y2, h_u_dadda_rca16_fa79_y4);
  fa fa_h_u_dadda_rca16_fa80_y2(h_u_dadda_rca16_fa79_y4, h_u_dadda_rca16_fa78_y4, h_u_dadda_rca16_fa77_y4, h_u_dadda_rca16_fa80_y2, h_u_dadda_rca16_fa80_y4);
  fa fa_h_u_dadda_rca16_fa81_y2(h_u_dadda_rca16_fa76_y4, h_u_dadda_rca16_fa75_y4, h_u_dadda_rca16_fa74_y4, h_u_dadda_rca16_fa81_y2, h_u_dadda_rca16_fa81_y4);
  fa fa_h_u_dadda_rca16_fa82_y2(h_u_dadda_rca16_fa73_y4, h_u_dadda_rca16_fa72_y4, h_u_dadda_rca16_fa71_y4, h_u_dadda_rca16_fa82_y2, h_u_dadda_rca16_fa82_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_5_y0(a_12, b_5, h_u_dadda_rca16_and_12_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_6_y0(a_11, b_6, h_u_dadda_rca16_and_11_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_7_y0(a_10, b_7, h_u_dadda_rca16_and_10_7_y0);
  fa fa_h_u_dadda_rca16_fa83_y2(h_u_dadda_rca16_and_12_5_y0, h_u_dadda_rca16_and_11_6_y0, h_u_dadda_rca16_and_10_7_y0, h_u_dadda_rca16_fa83_y2, h_u_dadda_rca16_fa83_y4);
  and_gate and_gate_h_u_dadda_rca16_and_9_8_y0(a_9, b_8, h_u_dadda_rca16_and_9_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_9_y0(a_8, b_9, h_u_dadda_rca16_and_8_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_10_y0(a_7, b_10, h_u_dadda_rca16_and_7_10_y0);
  fa fa_h_u_dadda_rca16_fa84_y2(h_u_dadda_rca16_and_9_8_y0, h_u_dadda_rca16_and_8_9_y0, h_u_dadda_rca16_and_7_10_y0, h_u_dadda_rca16_fa84_y2, h_u_dadda_rca16_fa84_y4);
  and_gate and_gate_h_u_dadda_rca16_and_6_11_y0(a_6, b_11, h_u_dadda_rca16_and_6_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_12_y0(a_5, b_12, h_u_dadda_rca16_and_5_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_13_y0(a_4, b_13, h_u_dadda_rca16_and_4_13_y0);
  fa fa_h_u_dadda_rca16_fa85_y2(h_u_dadda_rca16_and_6_11_y0, h_u_dadda_rca16_and_5_12_y0, h_u_dadda_rca16_and_4_13_y0, h_u_dadda_rca16_fa85_y2, h_u_dadda_rca16_fa85_y4);
  and_gate and_gate_h_u_dadda_rca16_and_3_14_y0(a_3, b_14, h_u_dadda_rca16_and_3_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_15_y0(a_2, b_15, h_u_dadda_rca16_and_2_15_y0);
  fa fa_h_u_dadda_rca16_fa86_y2(h_u_dadda_rca16_and_3_14_y0, h_u_dadda_rca16_and_2_15_y0, h_u_dadda_rca16_fa5_y2, h_u_dadda_rca16_fa86_y2, h_u_dadda_rca16_fa86_y4);
  fa fa_h_u_dadda_rca16_fa87_y2(h_u_dadda_rca16_fa6_y2, h_u_dadda_rca16_fa80_y2, h_u_dadda_rca16_fa81_y2, h_u_dadda_rca16_fa87_y2, h_u_dadda_rca16_fa87_y4);
  fa fa_h_u_dadda_rca16_fa88_y2(h_u_dadda_rca16_fa82_y2, h_u_dadda_rca16_fa83_y2, h_u_dadda_rca16_fa84_y2, h_u_dadda_rca16_fa88_y2, h_u_dadda_rca16_fa88_y4);
  fa fa_h_u_dadda_rca16_fa89_y2(h_u_dadda_rca16_fa88_y4, h_u_dadda_rca16_fa87_y4, h_u_dadda_rca16_fa86_y4, h_u_dadda_rca16_fa89_y2, h_u_dadda_rca16_fa89_y4);
  fa fa_h_u_dadda_rca16_fa90_y2(h_u_dadda_rca16_fa85_y4, h_u_dadda_rca16_fa84_y4, h_u_dadda_rca16_fa83_y4, h_u_dadda_rca16_fa90_y2, h_u_dadda_rca16_fa90_y4);
  fa fa_h_u_dadda_rca16_fa91_y2(h_u_dadda_rca16_fa82_y4, h_u_dadda_rca16_fa81_y4, h_u_dadda_rca16_fa80_y4, h_u_dadda_rca16_fa91_y2, h_u_dadda_rca16_fa91_y4);
  and_gate and_gate_h_u_dadda_rca16_and_14_4_y0(a_14, b_4, h_u_dadda_rca16_and_14_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_5_y0(a_13, b_5, h_u_dadda_rca16_and_13_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_6_y0(a_12, b_6, h_u_dadda_rca16_and_12_6_y0);
  fa fa_h_u_dadda_rca16_fa92_y2(h_u_dadda_rca16_and_14_4_y0, h_u_dadda_rca16_and_13_5_y0, h_u_dadda_rca16_and_12_6_y0, h_u_dadda_rca16_fa92_y2, h_u_dadda_rca16_fa92_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_7_y0(a_11, b_7, h_u_dadda_rca16_and_11_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_8_y0(a_10, b_8, h_u_dadda_rca16_and_10_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_9_y0(a_9, b_9, h_u_dadda_rca16_and_9_9_y0);
  fa fa_h_u_dadda_rca16_fa93_y2(h_u_dadda_rca16_and_11_7_y0, h_u_dadda_rca16_and_10_8_y0, h_u_dadda_rca16_and_9_9_y0, h_u_dadda_rca16_fa93_y2, h_u_dadda_rca16_fa93_y4);
  and_gate and_gate_h_u_dadda_rca16_and_8_10_y0(a_8, b_10, h_u_dadda_rca16_and_8_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_11_y0(a_7, b_11, h_u_dadda_rca16_and_7_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_12_y0(a_6, b_12, h_u_dadda_rca16_and_6_12_y0);
  fa fa_h_u_dadda_rca16_fa94_y2(h_u_dadda_rca16_and_8_10_y0, h_u_dadda_rca16_and_7_11_y0, h_u_dadda_rca16_and_6_12_y0, h_u_dadda_rca16_fa94_y2, h_u_dadda_rca16_fa94_y4);
  and_gate and_gate_h_u_dadda_rca16_and_5_13_y0(a_5, b_13, h_u_dadda_rca16_and_5_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_4_14_y0(a_4, b_14, h_u_dadda_rca16_and_4_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_3_15_y0(a_3, b_15, h_u_dadda_rca16_and_3_15_y0);
  fa fa_h_u_dadda_rca16_fa95_y2(h_u_dadda_rca16_and_5_13_y0, h_u_dadda_rca16_and_4_14_y0, h_u_dadda_rca16_and_3_15_y0, h_u_dadda_rca16_fa95_y2, h_u_dadda_rca16_fa95_y4);
  fa fa_h_u_dadda_rca16_fa96_y2(h_u_dadda_rca16_fa7_y2, h_u_dadda_rca16_fa89_y2, h_u_dadda_rca16_fa90_y2, h_u_dadda_rca16_fa96_y2, h_u_dadda_rca16_fa96_y4);
  fa fa_h_u_dadda_rca16_fa97_y2(h_u_dadda_rca16_fa91_y2, h_u_dadda_rca16_fa92_y2, h_u_dadda_rca16_fa93_y2, h_u_dadda_rca16_fa97_y2, h_u_dadda_rca16_fa97_y4);
  fa fa_h_u_dadda_rca16_fa98_y2(h_u_dadda_rca16_fa97_y4, h_u_dadda_rca16_fa96_y4, h_u_dadda_rca16_fa95_y4, h_u_dadda_rca16_fa98_y2, h_u_dadda_rca16_fa98_y4);
  fa fa_h_u_dadda_rca16_fa99_y2(h_u_dadda_rca16_fa94_y4, h_u_dadda_rca16_fa93_y4, h_u_dadda_rca16_fa92_y4, h_u_dadda_rca16_fa99_y2, h_u_dadda_rca16_fa99_y4);
  fa fa_h_u_dadda_rca16_fa100_y2(h_u_dadda_rca16_fa91_y4, h_u_dadda_rca16_fa90_y4, h_u_dadda_rca16_fa89_y4, h_u_dadda_rca16_fa100_y2, h_u_dadda_rca16_fa100_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_4_y0(a_15, b_4, h_u_dadda_rca16_and_15_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_5_y0(a_14, b_5, h_u_dadda_rca16_and_14_5_y0);
  fa fa_h_u_dadda_rca16_fa101_y2(h_u_dadda_rca16_fa7_y4, h_u_dadda_rca16_and_15_4_y0, h_u_dadda_rca16_and_14_5_y0, h_u_dadda_rca16_fa101_y2, h_u_dadda_rca16_fa101_y4);
  and_gate and_gate_h_u_dadda_rca16_and_13_6_y0(a_13, b_6, h_u_dadda_rca16_and_13_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_7_y0(a_12, b_7, h_u_dadda_rca16_and_12_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_8_y0(a_11, b_8, h_u_dadda_rca16_and_11_8_y0);
  fa fa_h_u_dadda_rca16_fa102_y2(h_u_dadda_rca16_and_13_6_y0, h_u_dadda_rca16_and_12_7_y0, h_u_dadda_rca16_and_11_8_y0, h_u_dadda_rca16_fa102_y2, h_u_dadda_rca16_fa102_y4);
  and_gate and_gate_h_u_dadda_rca16_and_10_9_y0(a_10, b_9, h_u_dadda_rca16_and_10_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_10_y0(a_9, b_10, h_u_dadda_rca16_and_9_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_11_y0(a_8, b_11, h_u_dadda_rca16_and_8_11_y0);
  fa fa_h_u_dadda_rca16_fa103_y2(h_u_dadda_rca16_and_10_9_y0, h_u_dadda_rca16_and_9_10_y0, h_u_dadda_rca16_and_8_11_y0, h_u_dadda_rca16_fa103_y2, h_u_dadda_rca16_fa103_y4);
  and_gate and_gate_h_u_dadda_rca16_and_7_12_y0(a_7, b_12, h_u_dadda_rca16_and_7_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_13_y0(a_6, b_13, h_u_dadda_rca16_and_6_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_14_y0(a_5, b_14, h_u_dadda_rca16_and_5_14_y0);
  fa fa_h_u_dadda_rca16_fa104_y2(h_u_dadda_rca16_and_7_12_y0, h_u_dadda_rca16_and_6_13_y0, h_u_dadda_rca16_and_5_14_y0, h_u_dadda_rca16_fa104_y2, h_u_dadda_rca16_fa104_y4);
  and_gate and_gate_h_u_dadda_rca16_and_4_15_y0(a_4, b_15, h_u_dadda_rca16_and_4_15_y0);
  fa fa_h_u_dadda_rca16_fa105_y2(h_u_dadda_rca16_and_4_15_y0, h_u_dadda_rca16_fa98_y2, h_u_dadda_rca16_fa99_y2, h_u_dadda_rca16_fa105_y2, h_u_dadda_rca16_fa105_y4);
  fa fa_h_u_dadda_rca16_fa106_y2(h_u_dadda_rca16_fa100_y2, h_u_dadda_rca16_fa101_y2, h_u_dadda_rca16_fa102_y2, h_u_dadda_rca16_fa106_y2, h_u_dadda_rca16_fa106_y4);
  fa fa_h_u_dadda_rca16_fa107_y2(h_u_dadda_rca16_fa106_y4, h_u_dadda_rca16_fa105_y4, h_u_dadda_rca16_fa104_y4, h_u_dadda_rca16_fa107_y2, h_u_dadda_rca16_fa107_y4);
  fa fa_h_u_dadda_rca16_fa108_y2(h_u_dadda_rca16_fa103_y4, h_u_dadda_rca16_fa102_y4, h_u_dadda_rca16_fa101_y4, h_u_dadda_rca16_fa108_y2, h_u_dadda_rca16_fa108_y4);
  fa fa_h_u_dadda_rca16_fa109_y2(h_u_dadda_rca16_fa100_y4, h_u_dadda_rca16_fa99_y4, h_u_dadda_rca16_fa98_y4, h_u_dadda_rca16_fa109_y2, h_u_dadda_rca16_fa109_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_5_y0(a_15, b_5, h_u_dadda_rca16_and_15_5_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_6_y0(a_14, b_6, h_u_dadda_rca16_and_14_6_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_7_y0(a_13, b_7, h_u_dadda_rca16_and_13_7_y0);
  fa fa_h_u_dadda_rca16_fa110_y2(h_u_dadda_rca16_and_15_5_y0, h_u_dadda_rca16_and_14_6_y0, h_u_dadda_rca16_and_13_7_y0, h_u_dadda_rca16_fa110_y2, h_u_dadda_rca16_fa110_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_8_y0(a_12, b_8, h_u_dadda_rca16_and_12_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_9_y0(a_11, b_9, h_u_dadda_rca16_and_11_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_10_y0(a_10, b_10, h_u_dadda_rca16_and_10_10_y0);
  fa fa_h_u_dadda_rca16_fa111_y2(h_u_dadda_rca16_and_12_8_y0, h_u_dadda_rca16_and_11_9_y0, h_u_dadda_rca16_and_10_10_y0, h_u_dadda_rca16_fa111_y2, h_u_dadda_rca16_fa111_y4);
  and_gate and_gate_h_u_dadda_rca16_and_9_11_y0(a_9, b_11, h_u_dadda_rca16_and_9_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_12_y0(a_8, b_12, h_u_dadda_rca16_and_8_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_13_y0(a_7, b_13, h_u_dadda_rca16_and_7_13_y0);
  fa fa_h_u_dadda_rca16_fa112_y2(h_u_dadda_rca16_and_9_11_y0, h_u_dadda_rca16_and_8_12_y0, h_u_dadda_rca16_and_7_13_y0, h_u_dadda_rca16_fa112_y2, h_u_dadda_rca16_fa112_y4);
  and_gate and_gate_h_u_dadda_rca16_and_6_14_y0(a_6, b_14, h_u_dadda_rca16_and_6_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_5_15_y0(a_5, b_15, h_u_dadda_rca16_and_5_15_y0);
  fa fa_h_u_dadda_rca16_fa113_y2(h_u_dadda_rca16_and_6_14_y0, h_u_dadda_rca16_and_5_15_y0, h_u_dadda_rca16_fa107_y2, h_u_dadda_rca16_fa113_y2, h_u_dadda_rca16_fa113_y4);
  fa fa_h_u_dadda_rca16_fa114_y2(h_u_dadda_rca16_fa108_y2, h_u_dadda_rca16_fa109_y2, h_u_dadda_rca16_fa110_y2, h_u_dadda_rca16_fa114_y2, h_u_dadda_rca16_fa114_y4);
  fa fa_h_u_dadda_rca16_fa115_y2(h_u_dadda_rca16_fa114_y4, h_u_dadda_rca16_fa113_y4, h_u_dadda_rca16_fa112_y4, h_u_dadda_rca16_fa115_y2, h_u_dadda_rca16_fa115_y4);
  fa fa_h_u_dadda_rca16_fa116_y2(h_u_dadda_rca16_fa111_y4, h_u_dadda_rca16_fa110_y4, h_u_dadda_rca16_fa109_y4, h_u_dadda_rca16_fa116_y2, h_u_dadda_rca16_fa116_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_6_y0(a_15, b_6, h_u_dadda_rca16_and_15_6_y0);
  fa fa_h_u_dadda_rca16_fa117_y2(h_u_dadda_rca16_fa108_y4, h_u_dadda_rca16_fa107_y4, h_u_dadda_rca16_and_15_6_y0, h_u_dadda_rca16_fa117_y2, h_u_dadda_rca16_fa117_y4);
  and_gate and_gate_h_u_dadda_rca16_and_14_7_y0(a_14, b_7, h_u_dadda_rca16_and_14_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_8_y0(a_13, b_8, h_u_dadda_rca16_and_13_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_9_y0(a_12, b_9, h_u_dadda_rca16_and_12_9_y0);
  fa fa_h_u_dadda_rca16_fa118_y2(h_u_dadda_rca16_and_14_7_y0, h_u_dadda_rca16_and_13_8_y0, h_u_dadda_rca16_and_12_9_y0, h_u_dadda_rca16_fa118_y2, h_u_dadda_rca16_fa118_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_10_y0(a_11, b_10, h_u_dadda_rca16_and_11_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_11_y0(a_10, b_11, h_u_dadda_rca16_and_10_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_12_y0(a_9, b_12, h_u_dadda_rca16_and_9_12_y0);
  fa fa_h_u_dadda_rca16_fa119_y2(h_u_dadda_rca16_and_11_10_y0, h_u_dadda_rca16_and_10_11_y0, h_u_dadda_rca16_and_9_12_y0, h_u_dadda_rca16_fa119_y2, h_u_dadda_rca16_fa119_y4);
  and_gate and_gate_h_u_dadda_rca16_and_8_13_y0(a_8, b_13, h_u_dadda_rca16_and_8_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_7_14_y0(a_7, b_14, h_u_dadda_rca16_and_7_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_6_15_y0(a_6, b_15, h_u_dadda_rca16_and_6_15_y0);
  fa fa_h_u_dadda_rca16_fa120_y2(h_u_dadda_rca16_and_8_13_y0, h_u_dadda_rca16_and_7_14_y0, h_u_dadda_rca16_and_6_15_y0, h_u_dadda_rca16_fa120_y2, h_u_dadda_rca16_fa120_y4);
  fa fa_h_u_dadda_rca16_fa121_y2(h_u_dadda_rca16_fa115_y2, h_u_dadda_rca16_fa116_y2, h_u_dadda_rca16_fa117_y2, h_u_dadda_rca16_fa121_y2, h_u_dadda_rca16_fa121_y4);
  fa fa_h_u_dadda_rca16_fa122_y2(h_u_dadda_rca16_fa121_y4, h_u_dadda_rca16_fa120_y4, h_u_dadda_rca16_fa119_y4, h_u_dadda_rca16_fa122_y2, h_u_dadda_rca16_fa122_y4);
  fa fa_h_u_dadda_rca16_fa123_y2(h_u_dadda_rca16_fa118_y4, h_u_dadda_rca16_fa117_y4, h_u_dadda_rca16_fa116_y4, h_u_dadda_rca16_fa123_y2, h_u_dadda_rca16_fa123_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_7_y0(a_15, b_7, h_u_dadda_rca16_and_15_7_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_8_y0(a_14, b_8, h_u_dadda_rca16_and_14_8_y0);
  fa fa_h_u_dadda_rca16_fa124_y2(h_u_dadda_rca16_fa115_y4, h_u_dadda_rca16_and_15_7_y0, h_u_dadda_rca16_and_14_8_y0, h_u_dadda_rca16_fa124_y2, h_u_dadda_rca16_fa124_y4);
  and_gate and_gate_h_u_dadda_rca16_and_13_9_y0(a_13, b_9, h_u_dadda_rca16_and_13_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_10_y0(a_12, b_10, h_u_dadda_rca16_and_12_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_11_y0(a_11, b_11, h_u_dadda_rca16_and_11_11_y0);
  fa fa_h_u_dadda_rca16_fa125_y2(h_u_dadda_rca16_and_13_9_y0, h_u_dadda_rca16_and_12_10_y0, h_u_dadda_rca16_and_11_11_y0, h_u_dadda_rca16_fa125_y2, h_u_dadda_rca16_fa125_y4);
  and_gate and_gate_h_u_dadda_rca16_and_10_12_y0(a_10, b_12, h_u_dadda_rca16_and_10_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_13_y0(a_9, b_13, h_u_dadda_rca16_and_9_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_14_y0(a_8, b_14, h_u_dadda_rca16_and_8_14_y0);
  fa fa_h_u_dadda_rca16_fa126_y2(h_u_dadda_rca16_and_10_12_y0, h_u_dadda_rca16_and_9_13_y0, h_u_dadda_rca16_and_8_14_y0, h_u_dadda_rca16_fa126_y2, h_u_dadda_rca16_fa126_y4);
  and_gate and_gate_h_u_dadda_rca16_and_7_15_y0(a_7, b_15, h_u_dadda_rca16_and_7_15_y0);
  fa fa_h_u_dadda_rca16_fa127_y2(h_u_dadda_rca16_and_7_15_y0, h_u_dadda_rca16_fa122_y2, h_u_dadda_rca16_fa123_y2, h_u_dadda_rca16_fa127_y2, h_u_dadda_rca16_fa127_y4);
  fa fa_h_u_dadda_rca16_fa128_y2(h_u_dadda_rca16_fa127_y4, h_u_dadda_rca16_fa126_y4, h_u_dadda_rca16_fa125_y4, h_u_dadda_rca16_fa128_y2, h_u_dadda_rca16_fa128_y4);
  fa fa_h_u_dadda_rca16_fa129_y2(h_u_dadda_rca16_fa124_y4, h_u_dadda_rca16_fa123_y4, h_u_dadda_rca16_fa122_y4, h_u_dadda_rca16_fa129_y2, h_u_dadda_rca16_fa129_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_8_y0(a_15, b_8, h_u_dadda_rca16_and_15_8_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_9_y0(a_14, b_9, h_u_dadda_rca16_and_14_9_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_10_y0(a_13, b_10, h_u_dadda_rca16_and_13_10_y0);
  fa fa_h_u_dadda_rca16_fa130_y2(h_u_dadda_rca16_and_15_8_y0, h_u_dadda_rca16_and_14_9_y0, h_u_dadda_rca16_and_13_10_y0, h_u_dadda_rca16_fa130_y2, h_u_dadda_rca16_fa130_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_11_y0(a_12, b_11, h_u_dadda_rca16_and_12_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_12_y0(a_11, b_12, h_u_dadda_rca16_and_11_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_13_y0(a_10, b_13, h_u_dadda_rca16_and_10_13_y0);
  fa fa_h_u_dadda_rca16_fa131_y2(h_u_dadda_rca16_and_12_11_y0, h_u_dadda_rca16_and_11_12_y0, h_u_dadda_rca16_and_10_13_y0, h_u_dadda_rca16_fa131_y2, h_u_dadda_rca16_fa131_y4);
  and_gate and_gate_h_u_dadda_rca16_and_9_14_y0(a_9, b_14, h_u_dadda_rca16_and_9_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_8_15_y0(a_8, b_15, h_u_dadda_rca16_and_8_15_y0);
  fa fa_h_u_dadda_rca16_fa132_y2(h_u_dadda_rca16_and_9_14_y0, h_u_dadda_rca16_and_8_15_y0, h_u_dadda_rca16_fa128_y2, h_u_dadda_rca16_fa132_y2, h_u_dadda_rca16_fa132_y4);
  fa fa_h_u_dadda_rca16_fa133_y2(h_u_dadda_rca16_fa132_y4, h_u_dadda_rca16_fa131_y4, h_u_dadda_rca16_fa130_y4, h_u_dadda_rca16_fa133_y2, h_u_dadda_rca16_fa133_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_9_y0(a_15, b_9, h_u_dadda_rca16_and_15_9_y0);
  fa fa_h_u_dadda_rca16_fa134_y2(h_u_dadda_rca16_fa129_y4, h_u_dadda_rca16_fa128_y4, h_u_dadda_rca16_and_15_9_y0, h_u_dadda_rca16_fa134_y2, h_u_dadda_rca16_fa134_y4);
  and_gate and_gate_h_u_dadda_rca16_and_14_10_y0(a_14, b_10, h_u_dadda_rca16_and_14_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_11_y0(a_13, b_11, h_u_dadda_rca16_and_13_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_12_y0(a_12, b_12, h_u_dadda_rca16_and_12_12_y0);
  fa fa_h_u_dadda_rca16_fa135_y2(h_u_dadda_rca16_and_14_10_y0, h_u_dadda_rca16_and_13_11_y0, h_u_dadda_rca16_and_12_12_y0, h_u_dadda_rca16_fa135_y2, h_u_dadda_rca16_fa135_y4);
  and_gate and_gate_h_u_dadda_rca16_and_11_13_y0(a_11, b_13, h_u_dadda_rca16_and_11_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_10_14_y0(a_10, b_14, h_u_dadda_rca16_and_10_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_9_15_y0(a_9, b_15, h_u_dadda_rca16_and_9_15_y0);
  fa fa_h_u_dadda_rca16_fa136_y2(h_u_dadda_rca16_and_11_13_y0, h_u_dadda_rca16_and_10_14_y0, h_u_dadda_rca16_and_9_15_y0, h_u_dadda_rca16_fa136_y2, h_u_dadda_rca16_fa136_y4);
  fa fa_h_u_dadda_rca16_fa137_y2(h_u_dadda_rca16_fa136_y4, h_u_dadda_rca16_fa135_y4, h_u_dadda_rca16_fa134_y4, h_u_dadda_rca16_fa137_y2, h_u_dadda_rca16_fa137_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_10_y0(a_15, b_10, h_u_dadda_rca16_and_15_10_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_11_y0(a_14, b_11, h_u_dadda_rca16_and_14_11_y0);
  fa fa_h_u_dadda_rca16_fa138_y2(h_u_dadda_rca16_fa133_y4, h_u_dadda_rca16_and_15_10_y0, h_u_dadda_rca16_and_14_11_y0, h_u_dadda_rca16_fa138_y2, h_u_dadda_rca16_fa138_y4);
  and_gate and_gate_h_u_dadda_rca16_and_13_12_y0(a_13, b_12, h_u_dadda_rca16_and_13_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_12_13_y0(a_12, b_13, h_u_dadda_rca16_and_12_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_14_y0(a_11, b_14, h_u_dadda_rca16_and_11_14_y0);
  fa fa_h_u_dadda_rca16_fa139_y2(h_u_dadda_rca16_and_13_12_y0, h_u_dadda_rca16_and_12_13_y0, h_u_dadda_rca16_and_11_14_y0, h_u_dadda_rca16_fa139_y2, h_u_dadda_rca16_fa139_y4);
  fa fa_h_u_dadda_rca16_fa140_y2(h_u_dadda_rca16_fa139_y4, h_u_dadda_rca16_fa138_y4, h_u_dadda_rca16_fa137_y4, h_u_dadda_rca16_fa140_y2, h_u_dadda_rca16_fa140_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_11_y0(a_15, b_11, h_u_dadda_rca16_and_15_11_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_12_y0(a_14, b_12, h_u_dadda_rca16_and_14_12_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_13_y0(a_13, b_13, h_u_dadda_rca16_and_13_13_y0);
  fa fa_h_u_dadda_rca16_fa141_y2(h_u_dadda_rca16_and_15_11_y0, h_u_dadda_rca16_and_14_12_y0, h_u_dadda_rca16_and_13_13_y0, h_u_dadda_rca16_fa141_y2, h_u_dadda_rca16_fa141_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_12_y0(a_15, b_12, h_u_dadda_rca16_and_15_12_y0);
  fa fa_h_u_dadda_rca16_fa142_y2(h_u_dadda_rca16_fa141_y4, h_u_dadda_rca16_fa140_y4, h_u_dadda_rca16_and_15_12_y0, h_u_dadda_rca16_fa142_y2, h_u_dadda_rca16_fa142_y4);
  and_gate and_gate_h_u_dadda_rca16_and_3_0_y0(a_3, b_0, h_u_dadda_rca16_and_3_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_2_1_y0(a_2, b_1, h_u_dadda_rca16_and_2_1_y0);
  ha ha_h_u_dadda_rca16_ha13_y0(h_u_dadda_rca16_and_3_0_y0, h_u_dadda_rca16_and_2_1_y0, h_u_dadda_rca16_ha13_y0, h_u_dadda_rca16_ha13_y1);
  and_gate and_gate_h_u_dadda_rca16_and_2_2_y0(a_2, b_2, h_u_dadda_rca16_and_2_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_3_y0(a_1, b_3, h_u_dadda_rca16_and_1_3_y0);
  fa fa_h_u_dadda_rca16_fa143_y2(h_u_dadda_rca16_ha13_y1, h_u_dadda_rca16_and_2_2_y0, h_u_dadda_rca16_and_1_3_y0, h_u_dadda_rca16_fa143_y2, h_u_dadda_rca16_fa143_y4);
  and_gate and_gate_h_u_dadda_rca16_and_1_4_y0(a_1, b_4, h_u_dadda_rca16_and_1_4_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_5_y0(a_0, b_5, h_u_dadda_rca16_and_0_5_y0);
  fa fa_h_u_dadda_rca16_fa144_y2(h_u_dadda_rca16_fa143_y4, h_u_dadda_rca16_and_1_4_y0, h_u_dadda_rca16_and_0_5_y0, h_u_dadda_rca16_fa144_y2, h_u_dadda_rca16_fa144_y4);
  and_gate and_gate_h_u_dadda_rca16_and_0_6_y0(a_0, b_6, h_u_dadda_rca16_and_0_6_y0);
  fa fa_h_u_dadda_rca16_fa145_y2(h_u_dadda_rca16_fa144_y4, h_u_dadda_rca16_and_0_6_y0, h_u_dadda_rca16_fa9_y2, h_u_dadda_rca16_fa145_y2, h_u_dadda_rca16_fa145_y4);
  fa fa_h_u_dadda_rca16_fa146_y2(h_u_dadda_rca16_fa145_y4, h_u_dadda_rca16_fa11_y2, h_u_dadda_rca16_fa12_y2, h_u_dadda_rca16_fa146_y2, h_u_dadda_rca16_fa146_y4);
  fa fa_h_u_dadda_rca16_fa147_y2(h_u_dadda_rca16_fa146_y4, h_u_dadda_rca16_fa15_y2, h_u_dadda_rca16_fa16_y2, h_u_dadda_rca16_fa147_y2, h_u_dadda_rca16_fa147_y4);
  fa fa_h_u_dadda_rca16_fa148_y2(h_u_dadda_rca16_fa147_y4, h_u_dadda_rca16_fa20_y2, h_u_dadda_rca16_fa21_y2, h_u_dadda_rca16_fa148_y2, h_u_dadda_rca16_fa148_y4);
  fa fa_h_u_dadda_rca16_fa149_y2(h_u_dadda_rca16_fa148_y4, h_u_dadda_rca16_fa26_y2, h_u_dadda_rca16_fa27_y2, h_u_dadda_rca16_fa149_y2, h_u_dadda_rca16_fa149_y4);
  fa fa_h_u_dadda_rca16_fa150_y2(h_u_dadda_rca16_fa149_y4, h_u_dadda_rca16_fa33_y2, h_u_dadda_rca16_fa34_y2, h_u_dadda_rca16_fa150_y2, h_u_dadda_rca16_fa150_y4);
  fa fa_h_u_dadda_rca16_fa151_y2(h_u_dadda_rca16_fa150_y4, h_u_dadda_rca16_fa41_y2, h_u_dadda_rca16_fa42_y2, h_u_dadda_rca16_fa151_y2, h_u_dadda_rca16_fa151_y4);
  fa fa_h_u_dadda_rca16_fa152_y2(h_u_dadda_rca16_fa151_y4, h_u_dadda_rca16_fa49_y2, h_u_dadda_rca16_fa50_y2, h_u_dadda_rca16_fa152_y2, h_u_dadda_rca16_fa152_y4);
  fa fa_h_u_dadda_rca16_fa153_y2(h_u_dadda_rca16_fa152_y4, h_u_dadda_rca16_fa58_y2, h_u_dadda_rca16_fa59_y2, h_u_dadda_rca16_fa153_y2, h_u_dadda_rca16_fa153_y4);
  fa fa_h_u_dadda_rca16_fa154_y2(h_u_dadda_rca16_fa153_y4, h_u_dadda_rca16_fa67_y2, h_u_dadda_rca16_fa68_y2, h_u_dadda_rca16_fa154_y2, h_u_dadda_rca16_fa154_y4);
  fa fa_h_u_dadda_rca16_fa155_y2(h_u_dadda_rca16_fa154_y4, h_u_dadda_rca16_fa76_y2, h_u_dadda_rca16_fa77_y2, h_u_dadda_rca16_fa155_y2, h_u_dadda_rca16_fa155_y4);
  fa fa_h_u_dadda_rca16_fa156_y2(h_u_dadda_rca16_fa155_y4, h_u_dadda_rca16_fa85_y2, h_u_dadda_rca16_fa86_y2, h_u_dadda_rca16_fa156_y2, h_u_dadda_rca16_fa156_y4);
  fa fa_h_u_dadda_rca16_fa157_y2(h_u_dadda_rca16_fa156_y4, h_u_dadda_rca16_fa94_y2, h_u_dadda_rca16_fa95_y2, h_u_dadda_rca16_fa157_y2, h_u_dadda_rca16_fa157_y4);
  fa fa_h_u_dadda_rca16_fa158_y2(h_u_dadda_rca16_fa157_y4, h_u_dadda_rca16_fa103_y2, h_u_dadda_rca16_fa104_y2, h_u_dadda_rca16_fa158_y2, h_u_dadda_rca16_fa158_y4);
  fa fa_h_u_dadda_rca16_fa159_y2(h_u_dadda_rca16_fa158_y4, h_u_dadda_rca16_fa111_y2, h_u_dadda_rca16_fa112_y2, h_u_dadda_rca16_fa159_y2, h_u_dadda_rca16_fa159_y4);
  fa fa_h_u_dadda_rca16_fa160_y2(h_u_dadda_rca16_fa159_y4, h_u_dadda_rca16_fa118_y2, h_u_dadda_rca16_fa119_y2, h_u_dadda_rca16_fa160_y2, h_u_dadda_rca16_fa160_y4);
  fa fa_h_u_dadda_rca16_fa161_y2(h_u_dadda_rca16_fa160_y4, h_u_dadda_rca16_fa124_y2, h_u_dadda_rca16_fa125_y2, h_u_dadda_rca16_fa161_y2, h_u_dadda_rca16_fa161_y4);
  fa fa_h_u_dadda_rca16_fa162_y2(h_u_dadda_rca16_fa161_y4, h_u_dadda_rca16_fa129_y2, h_u_dadda_rca16_fa130_y2, h_u_dadda_rca16_fa162_y2, h_u_dadda_rca16_fa162_y4);
  fa fa_h_u_dadda_rca16_fa163_y2(h_u_dadda_rca16_fa162_y4, h_u_dadda_rca16_fa133_y2, h_u_dadda_rca16_fa134_y2, h_u_dadda_rca16_fa163_y2, h_u_dadda_rca16_fa163_y4);
  and_gate and_gate_h_u_dadda_rca16_and_10_15_y0(a_10, b_15, h_u_dadda_rca16_and_10_15_y0);
  fa fa_h_u_dadda_rca16_fa164_y2(h_u_dadda_rca16_fa163_y4, h_u_dadda_rca16_and_10_15_y0, h_u_dadda_rca16_fa137_y2, h_u_dadda_rca16_fa164_y2, h_u_dadda_rca16_fa164_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_14_y0(a_12, b_14, h_u_dadda_rca16_and_12_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_11_15_y0(a_11, b_15, h_u_dadda_rca16_and_11_15_y0);
  fa fa_h_u_dadda_rca16_fa165_y2(h_u_dadda_rca16_fa164_y4, h_u_dadda_rca16_and_12_14_y0, h_u_dadda_rca16_and_11_15_y0, h_u_dadda_rca16_fa165_y2, h_u_dadda_rca16_fa165_y4);
  and_gate and_gate_h_u_dadda_rca16_and_14_13_y0(a_14, b_13, h_u_dadda_rca16_and_14_13_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_14_y0(a_13, b_14, h_u_dadda_rca16_and_13_14_y0);
  fa fa_h_u_dadda_rca16_fa166_y2(h_u_dadda_rca16_fa165_y4, h_u_dadda_rca16_and_14_13_y0, h_u_dadda_rca16_and_13_14_y0, h_u_dadda_rca16_fa166_y2, h_u_dadda_rca16_fa166_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_13_y0(a_15, b_13, h_u_dadda_rca16_and_15_13_y0);
  fa fa_h_u_dadda_rca16_fa167_y2(h_u_dadda_rca16_fa166_y4, h_u_dadda_rca16_fa142_y4, h_u_dadda_rca16_and_15_13_y0, h_u_dadda_rca16_fa167_y2, h_u_dadda_rca16_fa167_y4);
  and_gate and_gate_h_u_dadda_rca16_and_2_0_y0(a_2, b_0, h_u_dadda_rca16_and_2_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_1_y0(a_1, b_1, h_u_dadda_rca16_and_1_1_y0);
  ha ha_h_u_dadda_rca16_ha14_y0(h_u_dadda_rca16_and_2_0_y0, h_u_dadda_rca16_and_1_1_y0, h_u_dadda_rca16_ha14_y0, h_u_dadda_rca16_ha14_y1);
  and_gate and_gate_h_u_dadda_rca16_and_1_2_y0(a_1, b_2, h_u_dadda_rca16_and_1_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_3_y0(a_0, b_3, h_u_dadda_rca16_and_0_3_y0);
  fa fa_h_u_dadda_rca16_fa168_y2(h_u_dadda_rca16_ha14_y1, h_u_dadda_rca16_and_1_2_y0, h_u_dadda_rca16_and_0_3_y0, h_u_dadda_rca16_fa168_y2, h_u_dadda_rca16_fa168_y4);
  and_gate and_gate_h_u_dadda_rca16_and_0_4_y0(a_0, b_4, h_u_dadda_rca16_and_0_4_y0);
  fa fa_h_u_dadda_rca16_fa169_y2(h_u_dadda_rca16_fa168_y4, h_u_dadda_rca16_and_0_4_y0, h_u_dadda_rca16_ha4_y0, h_u_dadda_rca16_fa169_y2, h_u_dadda_rca16_fa169_y4);
  fa fa_h_u_dadda_rca16_fa170_y2(h_u_dadda_rca16_fa169_y4, h_u_dadda_rca16_fa8_y2, h_u_dadda_rca16_ha5_y0, h_u_dadda_rca16_fa170_y2, h_u_dadda_rca16_fa170_y4);
  fa fa_h_u_dadda_rca16_fa171_y2(h_u_dadda_rca16_fa170_y4, h_u_dadda_rca16_fa10_y2, h_u_dadda_rca16_ha6_y0, h_u_dadda_rca16_fa171_y2, h_u_dadda_rca16_fa171_y4);
  fa fa_h_u_dadda_rca16_fa172_y2(h_u_dadda_rca16_fa171_y4, h_u_dadda_rca16_fa13_y2, h_u_dadda_rca16_ha7_y0, h_u_dadda_rca16_fa172_y2, h_u_dadda_rca16_fa172_y4);
  fa fa_h_u_dadda_rca16_fa173_y2(h_u_dadda_rca16_fa172_y4, h_u_dadda_rca16_fa17_y2, h_u_dadda_rca16_ha8_y0, h_u_dadda_rca16_fa173_y2, h_u_dadda_rca16_fa173_y4);
  fa fa_h_u_dadda_rca16_fa174_y2(h_u_dadda_rca16_fa173_y4, h_u_dadda_rca16_fa22_y2, h_u_dadda_rca16_ha9_y0, h_u_dadda_rca16_fa174_y2, h_u_dadda_rca16_fa174_y4);
  fa fa_h_u_dadda_rca16_fa175_y2(h_u_dadda_rca16_fa174_y4, h_u_dadda_rca16_fa28_y2, h_u_dadda_rca16_ha10_y0, h_u_dadda_rca16_fa175_y2, h_u_dadda_rca16_fa175_y4);
  fa fa_h_u_dadda_rca16_fa176_y2(h_u_dadda_rca16_fa175_y4, h_u_dadda_rca16_fa35_y2, h_u_dadda_rca16_ha11_y0, h_u_dadda_rca16_fa176_y2, h_u_dadda_rca16_fa176_y4);
  fa fa_h_u_dadda_rca16_fa177_y2(h_u_dadda_rca16_fa176_y4, h_u_dadda_rca16_fa43_y2, h_u_dadda_rca16_ha12_y0, h_u_dadda_rca16_fa177_y2, h_u_dadda_rca16_fa177_y4);
  fa fa_h_u_dadda_rca16_fa178_y2(h_u_dadda_rca16_fa177_y4, h_u_dadda_rca16_fa51_y2, h_u_dadda_rca16_fa52_y2, h_u_dadda_rca16_fa178_y2, h_u_dadda_rca16_fa178_y4);
  fa fa_h_u_dadda_rca16_fa179_y2(h_u_dadda_rca16_fa178_y4, h_u_dadda_rca16_fa60_y2, h_u_dadda_rca16_fa61_y2, h_u_dadda_rca16_fa179_y2, h_u_dadda_rca16_fa179_y4);
  fa fa_h_u_dadda_rca16_fa180_y2(h_u_dadda_rca16_fa179_y4, h_u_dadda_rca16_fa69_y2, h_u_dadda_rca16_fa70_y2, h_u_dadda_rca16_fa180_y2, h_u_dadda_rca16_fa180_y4);
  fa fa_h_u_dadda_rca16_fa181_y2(h_u_dadda_rca16_fa180_y4, h_u_dadda_rca16_fa78_y2, h_u_dadda_rca16_fa79_y2, h_u_dadda_rca16_fa181_y2, h_u_dadda_rca16_fa181_y4);
  fa fa_h_u_dadda_rca16_fa182_y2(h_u_dadda_rca16_fa181_y4, h_u_dadda_rca16_fa87_y2, h_u_dadda_rca16_fa88_y2, h_u_dadda_rca16_fa182_y2, h_u_dadda_rca16_fa182_y4);
  fa fa_h_u_dadda_rca16_fa183_y2(h_u_dadda_rca16_fa182_y4, h_u_dadda_rca16_fa96_y2, h_u_dadda_rca16_fa97_y2, h_u_dadda_rca16_fa183_y2, h_u_dadda_rca16_fa183_y4);
  fa fa_h_u_dadda_rca16_fa184_y2(h_u_dadda_rca16_fa183_y4, h_u_dadda_rca16_fa105_y2, h_u_dadda_rca16_fa106_y2, h_u_dadda_rca16_fa184_y2, h_u_dadda_rca16_fa184_y4);
  fa fa_h_u_dadda_rca16_fa185_y2(h_u_dadda_rca16_fa184_y4, h_u_dadda_rca16_fa113_y2, h_u_dadda_rca16_fa114_y2, h_u_dadda_rca16_fa185_y2, h_u_dadda_rca16_fa185_y4);
  fa fa_h_u_dadda_rca16_fa186_y2(h_u_dadda_rca16_fa185_y4, h_u_dadda_rca16_fa120_y2, h_u_dadda_rca16_fa121_y2, h_u_dadda_rca16_fa186_y2, h_u_dadda_rca16_fa186_y4);
  fa fa_h_u_dadda_rca16_fa187_y2(h_u_dadda_rca16_fa186_y4, h_u_dadda_rca16_fa126_y2, h_u_dadda_rca16_fa127_y2, h_u_dadda_rca16_fa187_y2, h_u_dadda_rca16_fa187_y4);
  fa fa_h_u_dadda_rca16_fa188_y2(h_u_dadda_rca16_fa187_y4, h_u_dadda_rca16_fa131_y2, h_u_dadda_rca16_fa132_y2, h_u_dadda_rca16_fa188_y2, h_u_dadda_rca16_fa188_y4);
  fa fa_h_u_dadda_rca16_fa189_y2(h_u_dadda_rca16_fa188_y4, h_u_dadda_rca16_fa135_y2, h_u_dadda_rca16_fa136_y2, h_u_dadda_rca16_fa189_y2, h_u_dadda_rca16_fa189_y4);
  fa fa_h_u_dadda_rca16_fa190_y2(h_u_dadda_rca16_fa189_y4, h_u_dadda_rca16_fa138_y2, h_u_dadda_rca16_fa139_y2, h_u_dadda_rca16_fa190_y2, h_u_dadda_rca16_fa190_y4);
  fa fa_h_u_dadda_rca16_fa191_y2(h_u_dadda_rca16_fa190_y4, h_u_dadda_rca16_fa140_y2, h_u_dadda_rca16_fa141_y2, h_u_dadda_rca16_fa191_y2, h_u_dadda_rca16_fa191_y4);
  and_gate and_gate_h_u_dadda_rca16_and_12_15_y0(a_12, b_15, h_u_dadda_rca16_and_12_15_y0);
  fa fa_h_u_dadda_rca16_fa192_y2(h_u_dadda_rca16_fa191_y4, h_u_dadda_rca16_and_12_15_y0, h_u_dadda_rca16_fa142_y2, h_u_dadda_rca16_fa192_y2, h_u_dadda_rca16_fa192_y4);
  and_gate and_gate_h_u_dadda_rca16_and_14_14_y0(a_14, b_14, h_u_dadda_rca16_and_14_14_y0);
  and_gate and_gate_h_u_dadda_rca16_and_13_15_y0(a_13, b_15, h_u_dadda_rca16_and_13_15_y0);
  fa fa_h_u_dadda_rca16_fa193_y2(h_u_dadda_rca16_fa192_y4, h_u_dadda_rca16_and_14_14_y0, h_u_dadda_rca16_and_13_15_y0, h_u_dadda_rca16_fa193_y2, h_u_dadda_rca16_fa193_y4);
  and_gate and_gate_h_u_dadda_rca16_and_15_14_y0(a_15, b_14, h_u_dadda_rca16_and_15_14_y0);
  fa fa_h_u_dadda_rca16_fa194_y2(h_u_dadda_rca16_fa193_y4, h_u_dadda_rca16_fa167_y4, h_u_dadda_rca16_and_15_14_y0, h_u_dadda_rca16_fa194_y2, h_u_dadda_rca16_fa194_y4);
  and_gate and_gate_h_u_dadda_rca16_and_0_0_y0(a_0, b_0, h_u_dadda_rca16_and_0_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_1_0_y0(a_1, b_0, h_u_dadda_rca16_and_1_0_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_2_y0(a_0, b_2, h_u_dadda_rca16_and_0_2_y0);
  and_gate and_gate_h_u_dadda_rca16_and_14_15_y0(a_14, b_15, h_u_dadda_rca16_and_14_15_y0);
  and_gate and_gate_h_u_dadda_rca16_and_0_1_y0(a_0, b_1, h_u_dadda_rca16_and_0_1_y0);
  and_gate and_gate_h_u_dadda_rca16_and_15_15_y0(a_15, b_15, h_u_dadda_rca16_and_15_15_y0);
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[0] = h_u_dadda_rca16_and_1_0_y0;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[1] = h_u_dadda_rca16_and_0_2_y0;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[2] = h_u_dadda_rca16_ha13_y0;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[3] = h_u_dadda_rca16_fa143_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[4] = h_u_dadda_rca16_fa144_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[5] = h_u_dadda_rca16_fa145_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[6] = h_u_dadda_rca16_fa146_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[7] = h_u_dadda_rca16_fa147_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[8] = h_u_dadda_rca16_fa148_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[9] = h_u_dadda_rca16_fa149_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[10] = h_u_dadda_rca16_fa150_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[11] = h_u_dadda_rca16_fa151_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[12] = h_u_dadda_rca16_fa152_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[13] = h_u_dadda_rca16_fa153_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[14] = h_u_dadda_rca16_fa154_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[15] = h_u_dadda_rca16_fa155_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[16] = h_u_dadda_rca16_fa156_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[17] = h_u_dadda_rca16_fa157_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[18] = h_u_dadda_rca16_fa158_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[19] = h_u_dadda_rca16_fa159_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[20] = h_u_dadda_rca16_fa160_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[21] = h_u_dadda_rca16_fa161_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[22] = h_u_dadda_rca16_fa162_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[23] = h_u_dadda_rca16_fa163_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[24] = h_u_dadda_rca16_fa164_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[25] = h_u_dadda_rca16_fa165_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[26] = h_u_dadda_rca16_fa166_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[27] = h_u_dadda_rca16_fa167_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[28] = h_u_dadda_rca16_and_14_15_y0;
  assign h_u_dadda_rca16_u_rca30_u_rca30_a[29] = h_u_dadda_rca16_fa194_y4;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[0] = h_u_dadda_rca16_and_0_1_y0;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[1] = h_u_dadda_rca16_ha14_y0;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[2] = h_u_dadda_rca16_fa168_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[3] = h_u_dadda_rca16_fa169_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[4] = h_u_dadda_rca16_fa170_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[5] = h_u_dadda_rca16_fa171_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[6] = h_u_dadda_rca16_fa172_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[7] = h_u_dadda_rca16_fa173_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[8] = h_u_dadda_rca16_fa174_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[9] = h_u_dadda_rca16_fa175_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[10] = h_u_dadda_rca16_fa176_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[11] = h_u_dadda_rca16_fa177_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[12] = h_u_dadda_rca16_fa178_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[13] = h_u_dadda_rca16_fa179_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[14] = h_u_dadda_rca16_fa180_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[15] = h_u_dadda_rca16_fa181_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[16] = h_u_dadda_rca16_fa182_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[17] = h_u_dadda_rca16_fa183_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[18] = h_u_dadda_rca16_fa184_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[19] = h_u_dadda_rca16_fa185_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[20] = h_u_dadda_rca16_fa186_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[21] = h_u_dadda_rca16_fa187_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[22] = h_u_dadda_rca16_fa188_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[23] = h_u_dadda_rca16_fa189_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[24] = h_u_dadda_rca16_fa190_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[25] = h_u_dadda_rca16_fa191_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[26] = h_u_dadda_rca16_fa192_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[27] = h_u_dadda_rca16_fa193_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[28] = h_u_dadda_rca16_fa194_y2;
  assign h_u_dadda_rca16_u_rca30_u_rca30_b[29] = h_u_dadda_rca16_and_15_15_y0;
  u_rca30 u_rca30_out(h_u_dadda_rca16_u_rca30_u_rca30_a, h_u_dadda_rca16_u_rca30_u_rca30_b, h_u_dadda_rca16_u_rca30_out);
  assign h_u_dadda_rca16_u_rca30_ha_y0 = h_u_dadda_rca16_u_rca30_out[0];
  assign h_u_dadda_rca16_u_rca30_fa1_y2 = h_u_dadda_rca16_u_rca30_out[1];
  assign h_u_dadda_rca16_u_rca30_fa2_y2 = h_u_dadda_rca16_u_rca30_out[2];
  assign h_u_dadda_rca16_u_rca30_fa3_y2 = h_u_dadda_rca16_u_rca30_out[3];
  assign h_u_dadda_rca16_u_rca30_fa4_y2 = h_u_dadda_rca16_u_rca30_out[4];
  assign h_u_dadda_rca16_u_rca30_fa5_y2 = h_u_dadda_rca16_u_rca30_out[5];
  assign h_u_dadda_rca16_u_rca30_fa6_y2 = h_u_dadda_rca16_u_rca30_out[6];
  assign h_u_dadda_rca16_u_rca30_fa7_y2 = h_u_dadda_rca16_u_rca30_out[7];
  assign h_u_dadda_rca16_u_rca30_fa8_y2 = h_u_dadda_rca16_u_rca30_out[8];
  assign h_u_dadda_rca16_u_rca30_fa9_y2 = h_u_dadda_rca16_u_rca30_out[9];
  assign h_u_dadda_rca16_u_rca30_fa10_y2 = h_u_dadda_rca16_u_rca30_out[10];
  assign h_u_dadda_rca16_u_rca30_fa11_y2 = h_u_dadda_rca16_u_rca30_out[11];
  assign h_u_dadda_rca16_u_rca30_fa12_y2 = h_u_dadda_rca16_u_rca30_out[12];
  assign h_u_dadda_rca16_u_rca30_fa13_y2 = h_u_dadda_rca16_u_rca30_out[13];
  assign h_u_dadda_rca16_u_rca30_fa14_y2 = h_u_dadda_rca16_u_rca30_out[14];
  assign h_u_dadda_rca16_u_rca30_fa15_y2 = h_u_dadda_rca16_u_rca30_out[15];
  assign h_u_dadda_rca16_u_rca30_fa16_y2 = h_u_dadda_rca16_u_rca30_out[16];
  assign h_u_dadda_rca16_u_rca30_fa17_y2 = h_u_dadda_rca16_u_rca30_out[17];
  assign h_u_dadda_rca16_u_rca30_fa18_y2 = h_u_dadda_rca16_u_rca30_out[18];
  assign h_u_dadda_rca16_u_rca30_fa19_y2 = h_u_dadda_rca16_u_rca30_out[19];
  assign h_u_dadda_rca16_u_rca30_fa20_y2 = h_u_dadda_rca16_u_rca30_out[20];
  assign h_u_dadda_rca16_u_rca30_fa21_y2 = h_u_dadda_rca16_u_rca30_out[21];
  assign h_u_dadda_rca16_u_rca30_fa22_y2 = h_u_dadda_rca16_u_rca30_out[22];
  assign h_u_dadda_rca16_u_rca30_fa23_y2 = h_u_dadda_rca16_u_rca30_out[23];
  assign h_u_dadda_rca16_u_rca30_fa24_y2 = h_u_dadda_rca16_u_rca30_out[24];
  assign h_u_dadda_rca16_u_rca30_fa25_y2 = h_u_dadda_rca16_u_rca30_out[25];
  assign h_u_dadda_rca16_u_rca30_fa26_y2 = h_u_dadda_rca16_u_rca30_out[26];
  assign h_u_dadda_rca16_u_rca30_fa27_y2 = h_u_dadda_rca16_u_rca30_out[27];
  assign h_u_dadda_rca16_u_rca30_fa28_y2 = h_u_dadda_rca16_u_rca30_out[28];
  assign h_u_dadda_rca16_u_rca30_fa29_y2 = h_u_dadda_rca16_u_rca30_out[29];
  assign h_u_dadda_rca16_u_rca30_fa29_y4 = h_u_dadda_rca16_u_rca30_out[30];

  assign out[0] = h_u_dadda_rca16_and_0_0_y0;
  assign out[1] = h_u_dadda_rca16_u_rca30_ha_y0;
  assign out[2] = h_u_dadda_rca16_u_rca30_fa1_y2;
  assign out[3] = h_u_dadda_rca16_u_rca30_fa2_y2;
  assign out[4] = h_u_dadda_rca16_u_rca30_fa3_y2;
  assign out[5] = h_u_dadda_rca16_u_rca30_fa4_y2;
  assign out[6] = h_u_dadda_rca16_u_rca30_fa5_y2;
  assign out[7] = h_u_dadda_rca16_u_rca30_fa6_y2;
  assign out[8] = h_u_dadda_rca16_u_rca30_fa7_y2;
  assign out[9] = h_u_dadda_rca16_u_rca30_fa8_y2;
  assign out[10] = h_u_dadda_rca16_u_rca30_fa9_y2;
  assign out[11] = h_u_dadda_rca16_u_rca30_fa10_y2;
  assign out[12] = h_u_dadda_rca16_u_rca30_fa11_y2;
  assign out[13] = h_u_dadda_rca16_u_rca30_fa12_y2;
  assign out[14] = h_u_dadda_rca16_u_rca30_fa13_y2;
  assign out[15] = h_u_dadda_rca16_u_rca30_fa14_y2;
  assign out[16] = h_u_dadda_rca16_u_rca30_fa15_y2;
  assign out[17] = h_u_dadda_rca16_u_rca30_fa16_y2;
  assign out[18] = h_u_dadda_rca16_u_rca30_fa17_y2;
  assign out[19] = h_u_dadda_rca16_u_rca30_fa18_y2;
  assign out[20] = h_u_dadda_rca16_u_rca30_fa19_y2;
  assign out[21] = h_u_dadda_rca16_u_rca30_fa20_y2;
  assign out[22] = h_u_dadda_rca16_u_rca30_fa21_y2;
  assign out[23] = h_u_dadda_rca16_u_rca30_fa22_y2;
  assign out[24] = h_u_dadda_rca16_u_rca30_fa23_y2;
  assign out[25] = h_u_dadda_rca16_u_rca30_fa24_y2;
  assign out[26] = h_u_dadda_rca16_u_rca30_fa25_y2;
  assign out[27] = h_u_dadda_rca16_u_rca30_fa26_y2;
  assign out[28] = h_u_dadda_rca16_u_rca30_fa27_y2;
  assign out[29] = h_u_dadda_rca16_u_rca30_fa28_y2;
  assign out[30] = h_u_dadda_rca16_u_rca30_fa29_y2;
  assign out[31] = h_u_dadda_rca16_u_rca30_fa29_y4;
endmodule