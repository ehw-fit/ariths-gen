module arrdiv12(input [11:0] a, input [11:0] b, output [11:0] arrdiv12_out);
  wire arrdiv12_fs0_xor0;
  wire arrdiv12_fs0_not0;
  wire arrdiv12_fs0_and0;
  wire arrdiv12_fs0_not1;
  wire arrdiv12_fs1_xor1;
  wire arrdiv12_fs1_not1;
  wire arrdiv12_fs1_and1;
  wire arrdiv12_fs1_or0;
  wire arrdiv12_fs2_xor1;
  wire arrdiv12_fs2_not1;
  wire arrdiv12_fs2_and1;
  wire arrdiv12_fs2_or0;
  wire arrdiv12_fs3_xor1;
  wire arrdiv12_fs3_not1;
  wire arrdiv12_fs3_and1;
  wire arrdiv12_fs3_or0;
  wire arrdiv12_fs4_xor1;
  wire arrdiv12_fs4_not1;
  wire arrdiv12_fs4_and1;
  wire arrdiv12_fs4_or0;
  wire arrdiv12_fs5_xor1;
  wire arrdiv12_fs5_not1;
  wire arrdiv12_fs5_and1;
  wire arrdiv12_fs5_or0;
  wire arrdiv12_fs6_xor1;
  wire arrdiv12_fs6_not1;
  wire arrdiv12_fs6_and1;
  wire arrdiv12_fs6_or0;
  wire arrdiv12_fs7_xor1;
  wire arrdiv12_fs7_not1;
  wire arrdiv12_fs7_and1;
  wire arrdiv12_fs7_or0;
  wire arrdiv12_fs8_xor1;
  wire arrdiv12_fs8_not1;
  wire arrdiv12_fs8_and1;
  wire arrdiv12_fs8_or0;
  wire arrdiv12_fs9_xor1;
  wire arrdiv12_fs9_not1;
  wire arrdiv12_fs9_and1;
  wire arrdiv12_fs9_or0;
  wire arrdiv12_fs10_xor1;
  wire arrdiv12_fs10_not1;
  wire arrdiv12_fs10_and1;
  wire arrdiv12_fs10_or0;
  wire arrdiv12_fs11_xor1;
  wire arrdiv12_fs11_not1;
  wire arrdiv12_fs11_and1;
  wire arrdiv12_fs11_or0;
  wire arrdiv12_mux2to10_and0;
  wire arrdiv12_mux2to10_not0;
  wire arrdiv12_mux2to10_and1;
  wire arrdiv12_mux2to10_xor0;
  wire arrdiv12_mux2to11_not0;
  wire arrdiv12_mux2to11_and1;
  wire arrdiv12_mux2to12_not0;
  wire arrdiv12_mux2to12_and1;
  wire arrdiv12_mux2to13_not0;
  wire arrdiv12_mux2to13_and1;
  wire arrdiv12_mux2to14_not0;
  wire arrdiv12_mux2to14_and1;
  wire arrdiv12_mux2to15_not0;
  wire arrdiv12_mux2to15_and1;
  wire arrdiv12_mux2to16_not0;
  wire arrdiv12_mux2to16_and1;
  wire arrdiv12_mux2to17_not0;
  wire arrdiv12_mux2to17_and1;
  wire arrdiv12_mux2to18_not0;
  wire arrdiv12_mux2to18_and1;
  wire arrdiv12_mux2to19_not0;
  wire arrdiv12_mux2to19_and1;
  wire arrdiv12_mux2to110_not0;
  wire arrdiv12_mux2to110_and1;
  wire arrdiv12_not0;
  wire arrdiv12_fs12_xor0;
  wire arrdiv12_fs12_not0;
  wire arrdiv12_fs12_and0;
  wire arrdiv12_fs12_not1;
  wire arrdiv12_fs13_xor0;
  wire arrdiv12_fs13_not0;
  wire arrdiv12_fs13_and0;
  wire arrdiv12_fs13_xor1;
  wire arrdiv12_fs13_not1;
  wire arrdiv12_fs13_and1;
  wire arrdiv12_fs13_or0;
  wire arrdiv12_fs14_xor0;
  wire arrdiv12_fs14_not0;
  wire arrdiv12_fs14_and0;
  wire arrdiv12_fs14_xor1;
  wire arrdiv12_fs14_not1;
  wire arrdiv12_fs14_and1;
  wire arrdiv12_fs14_or0;
  wire arrdiv12_fs15_xor0;
  wire arrdiv12_fs15_not0;
  wire arrdiv12_fs15_and0;
  wire arrdiv12_fs15_xor1;
  wire arrdiv12_fs15_not1;
  wire arrdiv12_fs15_and1;
  wire arrdiv12_fs15_or0;
  wire arrdiv12_fs16_xor0;
  wire arrdiv12_fs16_not0;
  wire arrdiv12_fs16_and0;
  wire arrdiv12_fs16_xor1;
  wire arrdiv12_fs16_not1;
  wire arrdiv12_fs16_and1;
  wire arrdiv12_fs16_or0;
  wire arrdiv12_fs17_xor0;
  wire arrdiv12_fs17_not0;
  wire arrdiv12_fs17_and0;
  wire arrdiv12_fs17_xor1;
  wire arrdiv12_fs17_not1;
  wire arrdiv12_fs17_and1;
  wire arrdiv12_fs17_or0;
  wire arrdiv12_fs18_xor0;
  wire arrdiv12_fs18_not0;
  wire arrdiv12_fs18_and0;
  wire arrdiv12_fs18_xor1;
  wire arrdiv12_fs18_not1;
  wire arrdiv12_fs18_and1;
  wire arrdiv12_fs18_or0;
  wire arrdiv12_fs19_xor0;
  wire arrdiv12_fs19_not0;
  wire arrdiv12_fs19_and0;
  wire arrdiv12_fs19_xor1;
  wire arrdiv12_fs19_not1;
  wire arrdiv12_fs19_and1;
  wire arrdiv12_fs19_or0;
  wire arrdiv12_fs20_xor0;
  wire arrdiv12_fs20_not0;
  wire arrdiv12_fs20_and0;
  wire arrdiv12_fs20_xor1;
  wire arrdiv12_fs20_not1;
  wire arrdiv12_fs20_and1;
  wire arrdiv12_fs20_or0;
  wire arrdiv12_fs21_xor0;
  wire arrdiv12_fs21_not0;
  wire arrdiv12_fs21_and0;
  wire arrdiv12_fs21_xor1;
  wire arrdiv12_fs21_not1;
  wire arrdiv12_fs21_and1;
  wire arrdiv12_fs21_or0;
  wire arrdiv12_fs22_xor0;
  wire arrdiv12_fs22_not0;
  wire arrdiv12_fs22_and0;
  wire arrdiv12_fs22_xor1;
  wire arrdiv12_fs22_not1;
  wire arrdiv12_fs22_and1;
  wire arrdiv12_fs22_or0;
  wire arrdiv12_fs23_xor0;
  wire arrdiv12_fs23_not0;
  wire arrdiv12_fs23_and0;
  wire arrdiv12_fs23_xor1;
  wire arrdiv12_fs23_not1;
  wire arrdiv12_fs23_and1;
  wire arrdiv12_fs23_or0;
  wire arrdiv12_mux2to111_and0;
  wire arrdiv12_mux2to111_not0;
  wire arrdiv12_mux2to111_and1;
  wire arrdiv12_mux2to111_xor0;
  wire arrdiv12_mux2to112_and0;
  wire arrdiv12_mux2to112_not0;
  wire arrdiv12_mux2to112_and1;
  wire arrdiv12_mux2to112_xor0;
  wire arrdiv12_mux2to113_and0;
  wire arrdiv12_mux2to113_not0;
  wire arrdiv12_mux2to113_and1;
  wire arrdiv12_mux2to113_xor0;
  wire arrdiv12_mux2to114_and0;
  wire arrdiv12_mux2to114_not0;
  wire arrdiv12_mux2to114_and1;
  wire arrdiv12_mux2to114_xor0;
  wire arrdiv12_mux2to115_and0;
  wire arrdiv12_mux2to115_not0;
  wire arrdiv12_mux2to115_and1;
  wire arrdiv12_mux2to115_xor0;
  wire arrdiv12_mux2to116_and0;
  wire arrdiv12_mux2to116_not0;
  wire arrdiv12_mux2to116_and1;
  wire arrdiv12_mux2to116_xor0;
  wire arrdiv12_mux2to117_and0;
  wire arrdiv12_mux2to117_not0;
  wire arrdiv12_mux2to117_and1;
  wire arrdiv12_mux2to117_xor0;
  wire arrdiv12_mux2to118_and0;
  wire arrdiv12_mux2to118_not0;
  wire arrdiv12_mux2to118_and1;
  wire arrdiv12_mux2to118_xor0;
  wire arrdiv12_mux2to119_and0;
  wire arrdiv12_mux2to119_not0;
  wire arrdiv12_mux2to119_and1;
  wire arrdiv12_mux2to119_xor0;
  wire arrdiv12_mux2to120_and0;
  wire arrdiv12_mux2to120_not0;
  wire arrdiv12_mux2to120_and1;
  wire arrdiv12_mux2to120_xor0;
  wire arrdiv12_mux2to121_and0;
  wire arrdiv12_mux2to121_not0;
  wire arrdiv12_mux2to121_and1;
  wire arrdiv12_mux2to121_xor0;
  wire arrdiv12_not1;
  wire arrdiv12_fs24_xor0;
  wire arrdiv12_fs24_not0;
  wire arrdiv12_fs24_and0;
  wire arrdiv12_fs24_not1;
  wire arrdiv12_fs25_xor0;
  wire arrdiv12_fs25_not0;
  wire arrdiv12_fs25_and0;
  wire arrdiv12_fs25_xor1;
  wire arrdiv12_fs25_not1;
  wire arrdiv12_fs25_and1;
  wire arrdiv12_fs25_or0;
  wire arrdiv12_fs26_xor0;
  wire arrdiv12_fs26_not0;
  wire arrdiv12_fs26_and0;
  wire arrdiv12_fs26_xor1;
  wire arrdiv12_fs26_not1;
  wire arrdiv12_fs26_and1;
  wire arrdiv12_fs26_or0;
  wire arrdiv12_fs27_xor0;
  wire arrdiv12_fs27_not0;
  wire arrdiv12_fs27_and0;
  wire arrdiv12_fs27_xor1;
  wire arrdiv12_fs27_not1;
  wire arrdiv12_fs27_and1;
  wire arrdiv12_fs27_or0;
  wire arrdiv12_fs28_xor0;
  wire arrdiv12_fs28_not0;
  wire arrdiv12_fs28_and0;
  wire arrdiv12_fs28_xor1;
  wire arrdiv12_fs28_not1;
  wire arrdiv12_fs28_and1;
  wire arrdiv12_fs28_or0;
  wire arrdiv12_fs29_xor0;
  wire arrdiv12_fs29_not0;
  wire arrdiv12_fs29_and0;
  wire arrdiv12_fs29_xor1;
  wire arrdiv12_fs29_not1;
  wire arrdiv12_fs29_and1;
  wire arrdiv12_fs29_or0;
  wire arrdiv12_fs30_xor0;
  wire arrdiv12_fs30_not0;
  wire arrdiv12_fs30_and0;
  wire arrdiv12_fs30_xor1;
  wire arrdiv12_fs30_not1;
  wire arrdiv12_fs30_and1;
  wire arrdiv12_fs30_or0;
  wire arrdiv12_fs31_xor0;
  wire arrdiv12_fs31_not0;
  wire arrdiv12_fs31_and0;
  wire arrdiv12_fs31_xor1;
  wire arrdiv12_fs31_not1;
  wire arrdiv12_fs31_and1;
  wire arrdiv12_fs31_or0;
  wire arrdiv12_fs32_xor0;
  wire arrdiv12_fs32_not0;
  wire arrdiv12_fs32_and0;
  wire arrdiv12_fs32_xor1;
  wire arrdiv12_fs32_not1;
  wire arrdiv12_fs32_and1;
  wire arrdiv12_fs32_or0;
  wire arrdiv12_fs33_xor0;
  wire arrdiv12_fs33_not0;
  wire arrdiv12_fs33_and0;
  wire arrdiv12_fs33_xor1;
  wire arrdiv12_fs33_not1;
  wire arrdiv12_fs33_and1;
  wire arrdiv12_fs33_or0;
  wire arrdiv12_fs34_xor0;
  wire arrdiv12_fs34_not0;
  wire arrdiv12_fs34_and0;
  wire arrdiv12_fs34_xor1;
  wire arrdiv12_fs34_not1;
  wire arrdiv12_fs34_and1;
  wire arrdiv12_fs34_or0;
  wire arrdiv12_fs35_xor0;
  wire arrdiv12_fs35_not0;
  wire arrdiv12_fs35_and0;
  wire arrdiv12_fs35_xor1;
  wire arrdiv12_fs35_not1;
  wire arrdiv12_fs35_and1;
  wire arrdiv12_fs35_or0;
  wire arrdiv12_mux2to122_and0;
  wire arrdiv12_mux2to122_not0;
  wire arrdiv12_mux2to122_and1;
  wire arrdiv12_mux2to122_xor0;
  wire arrdiv12_mux2to123_and0;
  wire arrdiv12_mux2to123_not0;
  wire arrdiv12_mux2to123_and1;
  wire arrdiv12_mux2to123_xor0;
  wire arrdiv12_mux2to124_and0;
  wire arrdiv12_mux2to124_not0;
  wire arrdiv12_mux2to124_and1;
  wire arrdiv12_mux2to124_xor0;
  wire arrdiv12_mux2to125_and0;
  wire arrdiv12_mux2to125_not0;
  wire arrdiv12_mux2to125_and1;
  wire arrdiv12_mux2to125_xor0;
  wire arrdiv12_mux2to126_and0;
  wire arrdiv12_mux2to126_not0;
  wire arrdiv12_mux2to126_and1;
  wire arrdiv12_mux2to126_xor0;
  wire arrdiv12_mux2to127_and0;
  wire arrdiv12_mux2to127_not0;
  wire arrdiv12_mux2to127_and1;
  wire arrdiv12_mux2to127_xor0;
  wire arrdiv12_mux2to128_and0;
  wire arrdiv12_mux2to128_not0;
  wire arrdiv12_mux2to128_and1;
  wire arrdiv12_mux2to128_xor0;
  wire arrdiv12_mux2to129_and0;
  wire arrdiv12_mux2to129_not0;
  wire arrdiv12_mux2to129_and1;
  wire arrdiv12_mux2to129_xor0;
  wire arrdiv12_mux2to130_and0;
  wire arrdiv12_mux2to130_not0;
  wire arrdiv12_mux2to130_and1;
  wire arrdiv12_mux2to130_xor0;
  wire arrdiv12_mux2to131_and0;
  wire arrdiv12_mux2to131_not0;
  wire arrdiv12_mux2to131_and1;
  wire arrdiv12_mux2to131_xor0;
  wire arrdiv12_mux2to132_and0;
  wire arrdiv12_mux2to132_not0;
  wire arrdiv12_mux2to132_and1;
  wire arrdiv12_mux2to132_xor0;
  wire arrdiv12_not2;
  wire arrdiv12_fs36_xor0;
  wire arrdiv12_fs36_not0;
  wire arrdiv12_fs36_and0;
  wire arrdiv12_fs36_not1;
  wire arrdiv12_fs37_xor0;
  wire arrdiv12_fs37_not0;
  wire arrdiv12_fs37_and0;
  wire arrdiv12_fs37_xor1;
  wire arrdiv12_fs37_not1;
  wire arrdiv12_fs37_and1;
  wire arrdiv12_fs37_or0;
  wire arrdiv12_fs38_xor0;
  wire arrdiv12_fs38_not0;
  wire arrdiv12_fs38_and0;
  wire arrdiv12_fs38_xor1;
  wire arrdiv12_fs38_not1;
  wire arrdiv12_fs38_and1;
  wire arrdiv12_fs38_or0;
  wire arrdiv12_fs39_xor0;
  wire arrdiv12_fs39_not0;
  wire arrdiv12_fs39_and0;
  wire arrdiv12_fs39_xor1;
  wire arrdiv12_fs39_not1;
  wire arrdiv12_fs39_and1;
  wire arrdiv12_fs39_or0;
  wire arrdiv12_fs40_xor0;
  wire arrdiv12_fs40_not0;
  wire arrdiv12_fs40_and0;
  wire arrdiv12_fs40_xor1;
  wire arrdiv12_fs40_not1;
  wire arrdiv12_fs40_and1;
  wire arrdiv12_fs40_or0;
  wire arrdiv12_fs41_xor0;
  wire arrdiv12_fs41_not0;
  wire arrdiv12_fs41_and0;
  wire arrdiv12_fs41_xor1;
  wire arrdiv12_fs41_not1;
  wire arrdiv12_fs41_and1;
  wire arrdiv12_fs41_or0;
  wire arrdiv12_fs42_xor0;
  wire arrdiv12_fs42_not0;
  wire arrdiv12_fs42_and0;
  wire arrdiv12_fs42_xor1;
  wire arrdiv12_fs42_not1;
  wire arrdiv12_fs42_and1;
  wire arrdiv12_fs42_or0;
  wire arrdiv12_fs43_xor0;
  wire arrdiv12_fs43_not0;
  wire arrdiv12_fs43_and0;
  wire arrdiv12_fs43_xor1;
  wire arrdiv12_fs43_not1;
  wire arrdiv12_fs43_and1;
  wire arrdiv12_fs43_or0;
  wire arrdiv12_fs44_xor0;
  wire arrdiv12_fs44_not0;
  wire arrdiv12_fs44_and0;
  wire arrdiv12_fs44_xor1;
  wire arrdiv12_fs44_not1;
  wire arrdiv12_fs44_and1;
  wire arrdiv12_fs44_or0;
  wire arrdiv12_fs45_xor0;
  wire arrdiv12_fs45_not0;
  wire arrdiv12_fs45_and0;
  wire arrdiv12_fs45_xor1;
  wire arrdiv12_fs45_not1;
  wire arrdiv12_fs45_and1;
  wire arrdiv12_fs45_or0;
  wire arrdiv12_fs46_xor0;
  wire arrdiv12_fs46_not0;
  wire arrdiv12_fs46_and0;
  wire arrdiv12_fs46_xor1;
  wire arrdiv12_fs46_not1;
  wire arrdiv12_fs46_and1;
  wire arrdiv12_fs46_or0;
  wire arrdiv12_fs47_xor0;
  wire arrdiv12_fs47_not0;
  wire arrdiv12_fs47_and0;
  wire arrdiv12_fs47_xor1;
  wire arrdiv12_fs47_not1;
  wire arrdiv12_fs47_and1;
  wire arrdiv12_fs47_or0;
  wire arrdiv12_mux2to133_and0;
  wire arrdiv12_mux2to133_not0;
  wire arrdiv12_mux2to133_and1;
  wire arrdiv12_mux2to133_xor0;
  wire arrdiv12_mux2to134_and0;
  wire arrdiv12_mux2to134_not0;
  wire arrdiv12_mux2to134_and1;
  wire arrdiv12_mux2to134_xor0;
  wire arrdiv12_mux2to135_and0;
  wire arrdiv12_mux2to135_not0;
  wire arrdiv12_mux2to135_and1;
  wire arrdiv12_mux2to135_xor0;
  wire arrdiv12_mux2to136_and0;
  wire arrdiv12_mux2to136_not0;
  wire arrdiv12_mux2to136_and1;
  wire arrdiv12_mux2to136_xor0;
  wire arrdiv12_mux2to137_and0;
  wire arrdiv12_mux2to137_not0;
  wire arrdiv12_mux2to137_and1;
  wire arrdiv12_mux2to137_xor0;
  wire arrdiv12_mux2to138_and0;
  wire arrdiv12_mux2to138_not0;
  wire arrdiv12_mux2to138_and1;
  wire arrdiv12_mux2to138_xor0;
  wire arrdiv12_mux2to139_and0;
  wire arrdiv12_mux2to139_not0;
  wire arrdiv12_mux2to139_and1;
  wire arrdiv12_mux2to139_xor0;
  wire arrdiv12_mux2to140_and0;
  wire arrdiv12_mux2to140_not0;
  wire arrdiv12_mux2to140_and1;
  wire arrdiv12_mux2to140_xor0;
  wire arrdiv12_mux2to141_and0;
  wire arrdiv12_mux2to141_not0;
  wire arrdiv12_mux2to141_and1;
  wire arrdiv12_mux2to141_xor0;
  wire arrdiv12_mux2to142_and0;
  wire arrdiv12_mux2to142_not0;
  wire arrdiv12_mux2to142_and1;
  wire arrdiv12_mux2to142_xor0;
  wire arrdiv12_mux2to143_and0;
  wire arrdiv12_mux2to143_not0;
  wire arrdiv12_mux2to143_and1;
  wire arrdiv12_mux2to143_xor0;
  wire arrdiv12_not3;
  wire arrdiv12_fs48_xor0;
  wire arrdiv12_fs48_not0;
  wire arrdiv12_fs48_and0;
  wire arrdiv12_fs48_not1;
  wire arrdiv12_fs49_xor0;
  wire arrdiv12_fs49_not0;
  wire arrdiv12_fs49_and0;
  wire arrdiv12_fs49_xor1;
  wire arrdiv12_fs49_not1;
  wire arrdiv12_fs49_and1;
  wire arrdiv12_fs49_or0;
  wire arrdiv12_fs50_xor0;
  wire arrdiv12_fs50_not0;
  wire arrdiv12_fs50_and0;
  wire arrdiv12_fs50_xor1;
  wire arrdiv12_fs50_not1;
  wire arrdiv12_fs50_and1;
  wire arrdiv12_fs50_or0;
  wire arrdiv12_fs51_xor0;
  wire arrdiv12_fs51_not0;
  wire arrdiv12_fs51_and0;
  wire arrdiv12_fs51_xor1;
  wire arrdiv12_fs51_not1;
  wire arrdiv12_fs51_and1;
  wire arrdiv12_fs51_or0;
  wire arrdiv12_fs52_xor0;
  wire arrdiv12_fs52_not0;
  wire arrdiv12_fs52_and0;
  wire arrdiv12_fs52_xor1;
  wire arrdiv12_fs52_not1;
  wire arrdiv12_fs52_and1;
  wire arrdiv12_fs52_or0;
  wire arrdiv12_fs53_xor0;
  wire arrdiv12_fs53_not0;
  wire arrdiv12_fs53_and0;
  wire arrdiv12_fs53_xor1;
  wire arrdiv12_fs53_not1;
  wire arrdiv12_fs53_and1;
  wire arrdiv12_fs53_or0;
  wire arrdiv12_fs54_xor0;
  wire arrdiv12_fs54_not0;
  wire arrdiv12_fs54_and0;
  wire arrdiv12_fs54_xor1;
  wire arrdiv12_fs54_not1;
  wire arrdiv12_fs54_and1;
  wire arrdiv12_fs54_or0;
  wire arrdiv12_fs55_xor0;
  wire arrdiv12_fs55_not0;
  wire arrdiv12_fs55_and0;
  wire arrdiv12_fs55_xor1;
  wire arrdiv12_fs55_not1;
  wire arrdiv12_fs55_and1;
  wire arrdiv12_fs55_or0;
  wire arrdiv12_fs56_xor0;
  wire arrdiv12_fs56_not0;
  wire arrdiv12_fs56_and0;
  wire arrdiv12_fs56_xor1;
  wire arrdiv12_fs56_not1;
  wire arrdiv12_fs56_and1;
  wire arrdiv12_fs56_or0;
  wire arrdiv12_fs57_xor0;
  wire arrdiv12_fs57_not0;
  wire arrdiv12_fs57_and0;
  wire arrdiv12_fs57_xor1;
  wire arrdiv12_fs57_not1;
  wire arrdiv12_fs57_and1;
  wire arrdiv12_fs57_or0;
  wire arrdiv12_fs58_xor0;
  wire arrdiv12_fs58_not0;
  wire arrdiv12_fs58_and0;
  wire arrdiv12_fs58_xor1;
  wire arrdiv12_fs58_not1;
  wire arrdiv12_fs58_and1;
  wire arrdiv12_fs58_or0;
  wire arrdiv12_fs59_xor0;
  wire arrdiv12_fs59_not0;
  wire arrdiv12_fs59_and0;
  wire arrdiv12_fs59_xor1;
  wire arrdiv12_fs59_not1;
  wire arrdiv12_fs59_and1;
  wire arrdiv12_fs59_or0;
  wire arrdiv12_mux2to144_and0;
  wire arrdiv12_mux2to144_not0;
  wire arrdiv12_mux2to144_and1;
  wire arrdiv12_mux2to144_xor0;
  wire arrdiv12_mux2to145_and0;
  wire arrdiv12_mux2to145_not0;
  wire arrdiv12_mux2to145_and1;
  wire arrdiv12_mux2to145_xor0;
  wire arrdiv12_mux2to146_and0;
  wire arrdiv12_mux2to146_not0;
  wire arrdiv12_mux2to146_and1;
  wire arrdiv12_mux2to146_xor0;
  wire arrdiv12_mux2to147_and0;
  wire arrdiv12_mux2to147_not0;
  wire arrdiv12_mux2to147_and1;
  wire arrdiv12_mux2to147_xor0;
  wire arrdiv12_mux2to148_and0;
  wire arrdiv12_mux2to148_not0;
  wire arrdiv12_mux2to148_and1;
  wire arrdiv12_mux2to148_xor0;
  wire arrdiv12_mux2to149_and0;
  wire arrdiv12_mux2to149_not0;
  wire arrdiv12_mux2to149_and1;
  wire arrdiv12_mux2to149_xor0;
  wire arrdiv12_mux2to150_and0;
  wire arrdiv12_mux2to150_not0;
  wire arrdiv12_mux2to150_and1;
  wire arrdiv12_mux2to150_xor0;
  wire arrdiv12_mux2to151_and0;
  wire arrdiv12_mux2to151_not0;
  wire arrdiv12_mux2to151_and1;
  wire arrdiv12_mux2to151_xor0;
  wire arrdiv12_mux2to152_and0;
  wire arrdiv12_mux2to152_not0;
  wire arrdiv12_mux2to152_and1;
  wire arrdiv12_mux2to152_xor0;
  wire arrdiv12_mux2to153_and0;
  wire arrdiv12_mux2to153_not0;
  wire arrdiv12_mux2to153_and1;
  wire arrdiv12_mux2to153_xor0;
  wire arrdiv12_mux2to154_and0;
  wire arrdiv12_mux2to154_not0;
  wire arrdiv12_mux2to154_and1;
  wire arrdiv12_mux2to154_xor0;
  wire arrdiv12_not4;
  wire arrdiv12_fs60_xor0;
  wire arrdiv12_fs60_not0;
  wire arrdiv12_fs60_and0;
  wire arrdiv12_fs60_not1;
  wire arrdiv12_fs61_xor0;
  wire arrdiv12_fs61_not0;
  wire arrdiv12_fs61_and0;
  wire arrdiv12_fs61_xor1;
  wire arrdiv12_fs61_not1;
  wire arrdiv12_fs61_and1;
  wire arrdiv12_fs61_or0;
  wire arrdiv12_fs62_xor0;
  wire arrdiv12_fs62_not0;
  wire arrdiv12_fs62_and0;
  wire arrdiv12_fs62_xor1;
  wire arrdiv12_fs62_not1;
  wire arrdiv12_fs62_and1;
  wire arrdiv12_fs62_or0;
  wire arrdiv12_fs63_xor0;
  wire arrdiv12_fs63_not0;
  wire arrdiv12_fs63_and0;
  wire arrdiv12_fs63_xor1;
  wire arrdiv12_fs63_not1;
  wire arrdiv12_fs63_and1;
  wire arrdiv12_fs63_or0;
  wire arrdiv12_fs64_xor0;
  wire arrdiv12_fs64_not0;
  wire arrdiv12_fs64_and0;
  wire arrdiv12_fs64_xor1;
  wire arrdiv12_fs64_not1;
  wire arrdiv12_fs64_and1;
  wire arrdiv12_fs64_or0;
  wire arrdiv12_fs65_xor0;
  wire arrdiv12_fs65_not0;
  wire arrdiv12_fs65_and0;
  wire arrdiv12_fs65_xor1;
  wire arrdiv12_fs65_not1;
  wire arrdiv12_fs65_and1;
  wire arrdiv12_fs65_or0;
  wire arrdiv12_fs66_xor0;
  wire arrdiv12_fs66_not0;
  wire arrdiv12_fs66_and0;
  wire arrdiv12_fs66_xor1;
  wire arrdiv12_fs66_not1;
  wire arrdiv12_fs66_and1;
  wire arrdiv12_fs66_or0;
  wire arrdiv12_fs67_xor0;
  wire arrdiv12_fs67_not0;
  wire arrdiv12_fs67_and0;
  wire arrdiv12_fs67_xor1;
  wire arrdiv12_fs67_not1;
  wire arrdiv12_fs67_and1;
  wire arrdiv12_fs67_or0;
  wire arrdiv12_fs68_xor0;
  wire arrdiv12_fs68_not0;
  wire arrdiv12_fs68_and0;
  wire arrdiv12_fs68_xor1;
  wire arrdiv12_fs68_not1;
  wire arrdiv12_fs68_and1;
  wire arrdiv12_fs68_or0;
  wire arrdiv12_fs69_xor0;
  wire arrdiv12_fs69_not0;
  wire arrdiv12_fs69_and0;
  wire arrdiv12_fs69_xor1;
  wire arrdiv12_fs69_not1;
  wire arrdiv12_fs69_and1;
  wire arrdiv12_fs69_or0;
  wire arrdiv12_fs70_xor0;
  wire arrdiv12_fs70_not0;
  wire arrdiv12_fs70_and0;
  wire arrdiv12_fs70_xor1;
  wire arrdiv12_fs70_not1;
  wire arrdiv12_fs70_and1;
  wire arrdiv12_fs70_or0;
  wire arrdiv12_fs71_xor0;
  wire arrdiv12_fs71_not0;
  wire arrdiv12_fs71_and0;
  wire arrdiv12_fs71_xor1;
  wire arrdiv12_fs71_not1;
  wire arrdiv12_fs71_and1;
  wire arrdiv12_fs71_or0;
  wire arrdiv12_mux2to155_and0;
  wire arrdiv12_mux2to155_not0;
  wire arrdiv12_mux2to155_and1;
  wire arrdiv12_mux2to155_xor0;
  wire arrdiv12_mux2to156_and0;
  wire arrdiv12_mux2to156_not0;
  wire arrdiv12_mux2to156_and1;
  wire arrdiv12_mux2to156_xor0;
  wire arrdiv12_mux2to157_and0;
  wire arrdiv12_mux2to157_not0;
  wire arrdiv12_mux2to157_and1;
  wire arrdiv12_mux2to157_xor0;
  wire arrdiv12_mux2to158_and0;
  wire arrdiv12_mux2to158_not0;
  wire arrdiv12_mux2to158_and1;
  wire arrdiv12_mux2to158_xor0;
  wire arrdiv12_mux2to159_and0;
  wire arrdiv12_mux2to159_not0;
  wire arrdiv12_mux2to159_and1;
  wire arrdiv12_mux2to159_xor0;
  wire arrdiv12_mux2to160_and0;
  wire arrdiv12_mux2to160_not0;
  wire arrdiv12_mux2to160_and1;
  wire arrdiv12_mux2to160_xor0;
  wire arrdiv12_mux2to161_and0;
  wire arrdiv12_mux2to161_not0;
  wire arrdiv12_mux2to161_and1;
  wire arrdiv12_mux2to161_xor0;
  wire arrdiv12_mux2to162_and0;
  wire arrdiv12_mux2to162_not0;
  wire arrdiv12_mux2to162_and1;
  wire arrdiv12_mux2to162_xor0;
  wire arrdiv12_mux2to163_and0;
  wire arrdiv12_mux2to163_not0;
  wire arrdiv12_mux2to163_and1;
  wire arrdiv12_mux2to163_xor0;
  wire arrdiv12_mux2to164_and0;
  wire arrdiv12_mux2to164_not0;
  wire arrdiv12_mux2to164_and1;
  wire arrdiv12_mux2to164_xor0;
  wire arrdiv12_mux2to165_and0;
  wire arrdiv12_mux2to165_not0;
  wire arrdiv12_mux2to165_and1;
  wire arrdiv12_mux2to165_xor0;
  wire arrdiv12_not5;
  wire arrdiv12_fs72_xor0;
  wire arrdiv12_fs72_not0;
  wire arrdiv12_fs72_and0;
  wire arrdiv12_fs72_not1;
  wire arrdiv12_fs73_xor0;
  wire arrdiv12_fs73_not0;
  wire arrdiv12_fs73_and0;
  wire arrdiv12_fs73_xor1;
  wire arrdiv12_fs73_not1;
  wire arrdiv12_fs73_and1;
  wire arrdiv12_fs73_or0;
  wire arrdiv12_fs74_xor0;
  wire arrdiv12_fs74_not0;
  wire arrdiv12_fs74_and0;
  wire arrdiv12_fs74_xor1;
  wire arrdiv12_fs74_not1;
  wire arrdiv12_fs74_and1;
  wire arrdiv12_fs74_or0;
  wire arrdiv12_fs75_xor0;
  wire arrdiv12_fs75_not0;
  wire arrdiv12_fs75_and0;
  wire arrdiv12_fs75_xor1;
  wire arrdiv12_fs75_not1;
  wire arrdiv12_fs75_and1;
  wire arrdiv12_fs75_or0;
  wire arrdiv12_fs76_xor0;
  wire arrdiv12_fs76_not0;
  wire arrdiv12_fs76_and0;
  wire arrdiv12_fs76_xor1;
  wire arrdiv12_fs76_not1;
  wire arrdiv12_fs76_and1;
  wire arrdiv12_fs76_or0;
  wire arrdiv12_fs77_xor0;
  wire arrdiv12_fs77_not0;
  wire arrdiv12_fs77_and0;
  wire arrdiv12_fs77_xor1;
  wire arrdiv12_fs77_not1;
  wire arrdiv12_fs77_and1;
  wire arrdiv12_fs77_or0;
  wire arrdiv12_fs78_xor0;
  wire arrdiv12_fs78_not0;
  wire arrdiv12_fs78_and0;
  wire arrdiv12_fs78_xor1;
  wire arrdiv12_fs78_not1;
  wire arrdiv12_fs78_and1;
  wire arrdiv12_fs78_or0;
  wire arrdiv12_fs79_xor0;
  wire arrdiv12_fs79_not0;
  wire arrdiv12_fs79_and0;
  wire arrdiv12_fs79_xor1;
  wire arrdiv12_fs79_not1;
  wire arrdiv12_fs79_and1;
  wire arrdiv12_fs79_or0;
  wire arrdiv12_fs80_xor0;
  wire arrdiv12_fs80_not0;
  wire arrdiv12_fs80_and0;
  wire arrdiv12_fs80_xor1;
  wire arrdiv12_fs80_not1;
  wire arrdiv12_fs80_and1;
  wire arrdiv12_fs80_or0;
  wire arrdiv12_fs81_xor0;
  wire arrdiv12_fs81_not0;
  wire arrdiv12_fs81_and0;
  wire arrdiv12_fs81_xor1;
  wire arrdiv12_fs81_not1;
  wire arrdiv12_fs81_and1;
  wire arrdiv12_fs81_or0;
  wire arrdiv12_fs82_xor0;
  wire arrdiv12_fs82_not0;
  wire arrdiv12_fs82_and0;
  wire arrdiv12_fs82_xor1;
  wire arrdiv12_fs82_not1;
  wire arrdiv12_fs82_and1;
  wire arrdiv12_fs82_or0;
  wire arrdiv12_fs83_xor0;
  wire arrdiv12_fs83_not0;
  wire arrdiv12_fs83_and0;
  wire arrdiv12_fs83_xor1;
  wire arrdiv12_fs83_not1;
  wire arrdiv12_fs83_and1;
  wire arrdiv12_fs83_or0;
  wire arrdiv12_mux2to166_and0;
  wire arrdiv12_mux2to166_not0;
  wire arrdiv12_mux2to166_and1;
  wire arrdiv12_mux2to166_xor0;
  wire arrdiv12_mux2to167_and0;
  wire arrdiv12_mux2to167_not0;
  wire arrdiv12_mux2to167_and1;
  wire arrdiv12_mux2to167_xor0;
  wire arrdiv12_mux2to168_and0;
  wire arrdiv12_mux2to168_not0;
  wire arrdiv12_mux2to168_and1;
  wire arrdiv12_mux2to168_xor0;
  wire arrdiv12_mux2to169_and0;
  wire arrdiv12_mux2to169_not0;
  wire arrdiv12_mux2to169_and1;
  wire arrdiv12_mux2to169_xor0;
  wire arrdiv12_mux2to170_and0;
  wire arrdiv12_mux2to170_not0;
  wire arrdiv12_mux2to170_and1;
  wire arrdiv12_mux2to170_xor0;
  wire arrdiv12_mux2to171_and0;
  wire arrdiv12_mux2to171_not0;
  wire arrdiv12_mux2to171_and1;
  wire arrdiv12_mux2to171_xor0;
  wire arrdiv12_mux2to172_and0;
  wire arrdiv12_mux2to172_not0;
  wire arrdiv12_mux2to172_and1;
  wire arrdiv12_mux2to172_xor0;
  wire arrdiv12_mux2to173_and0;
  wire arrdiv12_mux2to173_not0;
  wire arrdiv12_mux2to173_and1;
  wire arrdiv12_mux2to173_xor0;
  wire arrdiv12_mux2to174_and0;
  wire arrdiv12_mux2to174_not0;
  wire arrdiv12_mux2to174_and1;
  wire arrdiv12_mux2to174_xor0;
  wire arrdiv12_mux2to175_and0;
  wire arrdiv12_mux2to175_not0;
  wire arrdiv12_mux2to175_and1;
  wire arrdiv12_mux2to175_xor0;
  wire arrdiv12_mux2to176_and0;
  wire arrdiv12_mux2to176_not0;
  wire arrdiv12_mux2to176_and1;
  wire arrdiv12_mux2to176_xor0;
  wire arrdiv12_not6;
  wire arrdiv12_fs84_xor0;
  wire arrdiv12_fs84_not0;
  wire arrdiv12_fs84_and0;
  wire arrdiv12_fs84_not1;
  wire arrdiv12_fs85_xor0;
  wire arrdiv12_fs85_not0;
  wire arrdiv12_fs85_and0;
  wire arrdiv12_fs85_xor1;
  wire arrdiv12_fs85_not1;
  wire arrdiv12_fs85_and1;
  wire arrdiv12_fs85_or0;
  wire arrdiv12_fs86_xor0;
  wire arrdiv12_fs86_not0;
  wire arrdiv12_fs86_and0;
  wire arrdiv12_fs86_xor1;
  wire arrdiv12_fs86_not1;
  wire arrdiv12_fs86_and1;
  wire arrdiv12_fs86_or0;
  wire arrdiv12_fs87_xor0;
  wire arrdiv12_fs87_not0;
  wire arrdiv12_fs87_and0;
  wire arrdiv12_fs87_xor1;
  wire arrdiv12_fs87_not1;
  wire arrdiv12_fs87_and1;
  wire arrdiv12_fs87_or0;
  wire arrdiv12_fs88_xor0;
  wire arrdiv12_fs88_not0;
  wire arrdiv12_fs88_and0;
  wire arrdiv12_fs88_xor1;
  wire arrdiv12_fs88_not1;
  wire arrdiv12_fs88_and1;
  wire arrdiv12_fs88_or0;
  wire arrdiv12_fs89_xor0;
  wire arrdiv12_fs89_not0;
  wire arrdiv12_fs89_and0;
  wire arrdiv12_fs89_xor1;
  wire arrdiv12_fs89_not1;
  wire arrdiv12_fs89_and1;
  wire arrdiv12_fs89_or0;
  wire arrdiv12_fs90_xor0;
  wire arrdiv12_fs90_not0;
  wire arrdiv12_fs90_and0;
  wire arrdiv12_fs90_xor1;
  wire arrdiv12_fs90_not1;
  wire arrdiv12_fs90_and1;
  wire arrdiv12_fs90_or0;
  wire arrdiv12_fs91_xor0;
  wire arrdiv12_fs91_not0;
  wire arrdiv12_fs91_and0;
  wire arrdiv12_fs91_xor1;
  wire arrdiv12_fs91_not1;
  wire arrdiv12_fs91_and1;
  wire arrdiv12_fs91_or0;
  wire arrdiv12_fs92_xor0;
  wire arrdiv12_fs92_not0;
  wire arrdiv12_fs92_and0;
  wire arrdiv12_fs92_xor1;
  wire arrdiv12_fs92_not1;
  wire arrdiv12_fs92_and1;
  wire arrdiv12_fs92_or0;
  wire arrdiv12_fs93_xor0;
  wire arrdiv12_fs93_not0;
  wire arrdiv12_fs93_and0;
  wire arrdiv12_fs93_xor1;
  wire arrdiv12_fs93_not1;
  wire arrdiv12_fs93_and1;
  wire arrdiv12_fs93_or0;
  wire arrdiv12_fs94_xor0;
  wire arrdiv12_fs94_not0;
  wire arrdiv12_fs94_and0;
  wire arrdiv12_fs94_xor1;
  wire arrdiv12_fs94_not1;
  wire arrdiv12_fs94_and1;
  wire arrdiv12_fs94_or0;
  wire arrdiv12_fs95_xor0;
  wire arrdiv12_fs95_not0;
  wire arrdiv12_fs95_and0;
  wire arrdiv12_fs95_xor1;
  wire arrdiv12_fs95_not1;
  wire arrdiv12_fs95_and1;
  wire arrdiv12_fs95_or0;
  wire arrdiv12_mux2to177_and0;
  wire arrdiv12_mux2to177_not0;
  wire arrdiv12_mux2to177_and1;
  wire arrdiv12_mux2to177_xor0;
  wire arrdiv12_mux2to178_and0;
  wire arrdiv12_mux2to178_not0;
  wire arrdiv12_mux2to178_and1;
  wire arrdiv12_mux2to178_xor0;
  wire arrdiv12_mux2to179_and0;
  wire arrdiv12_mux2to179_not0;
  wire arrdiv12_mux2to179_and1;
  wire arrdiv12_mux2to179_xor0;
  wire arrdiv12_mux2to180_and0;
  wire arrdiv12_mux2to180_not0;
  wire arrdiv12_mux2to180_and1;
  wire arrdiv12_mux2to180_xor0;
  wire arrdiv12_mux2to181_and0;
  wire arrdiv12_mux2to181_not0;
  wire arrdiv12_mux2to181_and1;
  wire arrdiv12_mux2to181_xor0;
  wire arrdiv12_mux2to182_and0;
  wire arrdiv12_mux2to182_not0;
  wire arrdiv12_mux2to182_and1;
  wire arrdiv12_mux2to182_xor0;
  wire arrdiv12_mux2to183_and0;
  wire arrdiv12_mux2to183_not0;
  wire arrdiv12_mux2to183_and1;
  wire arrdiv12_mux2to183_xor0;
  wire arrdiv12_mux2to184_and0;
  wire arrdiv12_mux2to184_not0;
  wire arrdiv12_mux2to184_and1;
  wire arrdiv12_mux2to184_xor0;
  wire arrdiv12_mux2to185_and0;
  wire arrdiv12_mux2to185_not0;
  wire arrdiv12_mux2to185_and1;
  wire arrdiv12_mux2to185_xor0;
  wire arrdiv12_mux2to186_and0;
  wire arrdiv12_mux2to186_not0;
  wire arrdiv12_mux2to186_and1;
  wire arrdiv12_mux2to186_xor0;
  wire arrdiv12_mux2to187_and0;
  wire arrdiv12_mux2to187_not0;
  wire arrdiv12_mux2to187_and1;
  wire arrdiv12_mux2to187_xor0;
  wire arrdiv12_not7;
  wire arrdiv12_fs96_xor0;
  wire arrdiv12_fs96_not0;
  wire arrdiv12_fs96_and0;
  wire arrdiv12_fs96_not1;
  wire arrdiv12_fs97_xor0;
  wire arrdiv12_fs97_not0;
  wire arrdiv12_fs97_and0;
  wire arrdiv12_fs97_xor1;
  wire arrdiv12_fs97_not1;
  wire arrdiv12_fs97_and1;
  wire arrdiv12_fs97_or0;
  wire arrdiv12_fs98_xor0;
  wire arrdiv12_fs98_not0;
  wire arrdiv12_fs98_and0;
  wire arrdiv12_fs98_xor1;
  wire arrdiv12_fs98_not1;
  wire arrdiv12_fs98_and1;
  wire arrdiv12_fs98_or0;
  wire arrdiv12_fs99_xor0;
  wire arrdiv12_fs99_not0;
  wire arrdiv12_fs99_and0;
  wire arrdiv12_fs99_xor1;
  wire arrdiv12_fs99_not1;
  wire arrdiv12_fs99_and1;
  wire arrdiv12_fs99_or0;
  wire arrdiv12_fs100_xor0;
  wire arrdiv12_fs100_not0;
  wire arrdiv12_fs100_and0;
  wire arrdiv12_fs100_xor1;
  wire arrdiv12_fs100_not1;
  wire arrdiv12_fs100_and1;
  wire arrdiv12_fs100_or0;
  wire arrdiv12_fs101_xor0;
  wire arrdiv12_fs101_not0;
  wire arrdiv12_fs101_and0;
  wire arrdiv12_fs101_xor1;
  wire arrdiv12_fs101_not1;
  wire arrdiv12_fs101_and1;
  wire arrdiv12_fs101_or0;
  wire arrdiv12_fs102_xor0;
  wire arrdiv12_fs102_not0;
  wire arrdiv12_fs102_and0;
  wire arrdiv12_fs102_xor1;
  wire arrdiv12_fs102_not1;
  wire arrdiv12_fs102_and1;
  wire arrdiv12_fs102_or0;
  wire arrdiv12_fs103_xor0;
  wire arrdiv12_fs103_not0;
  wire arrdiv12_fs103_and0;
  wire arrdiv12_fs103_xor1;
  wire arrdiv12_fs103_not1;
  wire arrdiv12_fs103_and1;
  wire arrdiv12_fs103_or0;
  wire arrdiv12_fs104_xor0;
  wire arrdiv12_fs104_not0;
  wire arrdiv12_fs104_and0;
  wire arrdiv12_fs104_xor1;
  wire arrdiv12_fs104_not1;
  wire arrdiv12_fs104_and1;
  wire arrdiv12_fs104_or0;
  wire arrdiv12_fs105_xor0;
  wire arrdiv12_fs105_not0;
  wire arrdiv12_fs105_and0;
  wire arrdiv12_fs105_xor1;
  wire arrdiv12_fs105_not1;
  wire arrdiv12_fs105_and1;
  wire arrdiv12_fs105_or0;
  wire arrdiv12_fs106_xor0;
  wire arrdiv12_fs106_not0;
  wire arrdiv12_fs106_and0;
  wire arrdiv12_fs106_xor1;
  wire arrdiv12_fs106_not1;
  wire arrdiv12_fs106_and1;
  wire arrdiv12_fs106_or0;
  wire arrdiv12_fs107_xor0;
  wire arrdiv12_fs107_not0;
  wire arrdiv12_fs107_and0;
  wire arrdiv12_fs107_xor1;
  wire arrdiv12_fs107_not1;
  wire arrdiv12_fs107_and1;
  wire arrdiv12_fs107_or0;
  wire arrdiv12_mux2to188_and0;
  wire arrdiv12_mux2to188_not0;
  wire arrdiv12_mux2to188_and1;
  wire arrdiv12_mux2to188_xor0;
  wire arrdiv12_mux2to189_and0;
  wire arrdiv12_mux2to189_not0;
  wire arrdiv12_mux2to189_and1;
  wire arrdiv12_mux2to189_xor0;
  wire arrdiv12_mux2to190_and0;
  wire arrdiv12_mux2to190_not0;
  wire arrdiv12_mux2to190_and1;
  wire arrdiv12_mux2to190_xor0;
  wire arrdiv12_mux2to191_and0;
  wire arrdiv12_mux2to191_not0;
  wire arrdiv12_mux2to191_and1;
  wire arrdiv12_mux2to191_xor0;
  wire arrdiv12_mux2to192_and0;
  wire arrdiv12_mux2to192_not0;
  wire arrdiv12_mux2to192_and1;
  wire arrdiv12_mux2to192_xor0;
  wire arrdiv12_mux2to193_and0;
  wire arrdiv12_mux2to193_not0;
  wire arrdiv12_mux2to193_and1;
  wire arrdiv12_mux2to193_xor0;
  wire arrdiv12_mux2to194_and0;
  wire arrdiv12_mux2to194_not0;
  wire arrdiv12_mux2to194_and1;
  wire arrdiv12_mux2to194_xor0;
  wire arrdiv12_mux2to195_and0;
  wire arrdiv12_mux2to195_not0;
  wire arrdiv12_mux2to195_and1;
  wire arrdiv12_mux2to195_xor0;
  wire arrdiv12_mux2to196_and0;
  wire arrdiv12_mux2to196_not0;
  wire arrdiv12_mux2to196_and1;
  wire arrdiv12_mux2to196_xor0;
  wire arrdiv12_mux2to197_and0;
  wire arrdiv12_mux2to197_not0;
  wire arrdiv12_mux2to197_and1;
  wire arrdiv12_mux2to197_xor0;
  wire arrdiv12_mux2to198_and0;
  wire arrdiv12_mux2to198_not0;
  wire arrdiv12_mux2to198_and1;
  wire arrdiv12_mux2to198_xor0;
  wire arrdiv12_not8;
  wire arrdiv12_fs108_xor0;
  wire arrdiv12_fs108_not0;
  wire arrdiv12_fs108_and0;
  wire arrdiv12_fs108_not1;
  wire arrdiv12_fs109_xor0;
  wire arrdiv12_fs109_not0;
  wire arrdiv12_fs109_and0;
  wire arrdiv12_fs109_xor1;
  wire arrdiv12_fs109_not1;
  wire arrdiv12_fs109_and1;
  wire arrdiv12_fs109_or0;
  wire arrdiv12_fs110_xor0;
  wire arrdiv12_fs110_not0;
  wire arrdiv12_fs110_and0;
  wire arrdiv12_fs110_xor1;
  wire arrdiv12_fs110_not1;
  wire arrdiv12_fs110_and1;
  wire arrdiv12_fs110_or0;
  wire arrdiv12_fs111_xor0;
  wire arrdiv12_fs111_not0;
  wire arrdiv12_fs111_and0;
  wire arrdiv12_fs111_xor1;
  wire arrdiv12_fs111_not1;
  wire arrdiv12_fs111_and1;
  wire arrdiv12_fs111_or0;
  wire arrdiv12_fs112_xor0;
  wire arrdiv12_fs112_not0;
  wire arrdiv12_fs112_and0;
  wire arrdiv12_fs112_xor1;
  wire arrdiv12_fs112_not1;
  wire arrdiv12_fs112_and1;
  wire arrdiv12_fs112_or0;
  wire arrdiv12_fs113_xor0;
  wire arrdiv12_fs113_not0;
  wire arrdiv12_fs113_and0;
  wire arrdiv12_fs113_xor1;
  wire arrdiv12_fs113_not1;
  wire arrdiv12_fs113_and1;
  wire arrdiv12_fs113_or0;
  wire arrdiv12_fs114_xor0;
  wire arrdiv12_fs114_not0;
  wire arrdiv12_fs114_and0;
  wire arrdiv12_fs114_xor1;
  wire arrdiv12_fs114_not1;
  wire arrdiv12_fs114_and1;
  wire arrdiv12_fs114_or0;
  wire arrdiv12_fs115_xor0;
  wire arrdiv12_fs115_not0;
  wire arrdiv12_fs115_and0;
  wire arrdiv12_fs115_xor1;
  wire arrdiv12_fs115_not1;
  wire arrdiv12_fs115_and1;
  wire arrdiv12_fs115_or0;
  wire arrdiv12_fs116_xor0;
  wire arrdiv12_fs116_not0;
  wire arrdiv12_fs116_and0;
  wire arrdiv12_fs116_xor1;
  wire arrdiv12_fs116_not1;
  wire arrdiv12_fs116_and1;
  wire arrdiv12_fs116_or0;
  wire arrdiv12_fs117_xor0;
  wire arrdiv12_fs117_not0;
  wire arrdiv12_fs117_and0;
  wire arrdiv12_fs117_xor1;
  wire arrdiv12_fs117_not1;
  wire arrdiv12_fs117_and1;
  wire arrdiv12_fs117_or0;
  wire arrdiv12_fs118_xor0;
  wire arrdiv12_fs118_not0;
  wire arrdiv12_fs118_and0;
  wire arrdiv12_fs118_xor1;
  wire arrdiv12_fs118_not1;
  wire arrdiv12_fs118_and1;
  wire arrdiv12_fs118_or0;
  wire arrdiv12_fs119_xor0;
  wire arrdiv12_fs119_not0;
  wire arrdiv12_fs119_and0;
  wire arrdiv12_fs119_xor1;
  wire arrdiv12_fs119_not1;
  wire arrdiv12_fs119_and1;
  wire arrdiv12_fs119_or0;
  wire arrdiv12_mux2to199_and0;
  wire arrdiv12_mux2to199_not0;
  wire arrdiv12_mux2to199_and1;
  wire arrdiv12_mux2to199_xor0;
  wire arrdiv12_mux2to1100_and0;
  wire arrdiv12_mux2to1100_not0;
  wire arrdiv12_mux2to1100_and1;
  wire arrdiv12_mux2to1100_xor0;
  wire arrdiv12_mux2to1101_and0;
  wire arrdiv12_mux2to1101_not0;
  wire arrdiv12_mux2to1101_and1;
  wire arrdiv12_mux2to1101_xor0;
  wire arrdiv12_mux2to1102_and0;
  wire arrdiv12_mux2to1102_not0;
  wire arrdiv12_mux2to1102_and1;
  wire arrdiv12_mux2to1102_xor0;
  wire arrdiv12_mux2to1103_and0;
  wire arrdiv12_mux2to1103_not0;
  wire arrdiv12_mux2to1103_and1;
  wire arrdiv12_mux2to1103_xor0;
  wire arrdiv12_mux2to1104_and0;
  wire arrdiv12_mux2to1104_not0;
  wire arrdiv12_mux2to1104_and1;
  wire arrdiv12_mux2to1104_xor0;
  wire arrdiv12_mux2to1105_and0;
  wire arrdiv12_mux2to1105_not0;
  wire arrdiv12_mux2to1105_and1;
  wire arrdiv12_mux2to1105_xor0;
  wire arrdiv12_mux2to1106_and0;
  wire arrdiv12_mux2to1106_not0;
  wire arrdiv12_mux2to1106_and1;
  wire arrdiv12_mux2to1106_xor0;
  wire arrdiv12_mux2to1107_and0;
  wire arrdiv12_mux2to1107_not0;
  wire arrdiv12_mux2to1107_and1;
  wire arrdiv12_mux2to1107_xor0;
  wire arrdiv12_mux2to1108_and0;
  wire arrdiv12_mux2to1108_not0;
  wire arrdiv12_mux2to1108_and1;
  wire arrdiv12_mux2to1108_xor0;
  wire arrdiv12_mux2to1109_and0;
  wire arrdiv12_mux2to1109_not0;
  wire arrdiv12_mux2to1109_and1;
  wire arrdiv12_mux2to1109_xor0;
  wire arrdiv12_not9;
  wire arrdiv12_fs120_xor0;
  wire arrdiv12_fs120_not0;
  wire arrdiv12_fs120_and0;
  wire arrdiv12_fs120_not1;
  wire arrdiv12_fs121_xor0;
  wire arrdiv12_fs121_not0;
  wire arrdiv12_fs121_and0;
  wire arrdiv12_fs121_xor1;
  wire arrdiv12_fs121_not1;
  wire arrdiv12_fs121_and1;
  wire arrdiv12_fs121_or0;
  wire arrdiv12_fs122_xor0;
  wire arrdiv12_fs122_not0;
  wire arrdiv12_fs122_and0;
  wire arrdiv12_fs122_xor1;
  wire arrdiv12_fs122_not1;
  wire arrdiv12_fs122_and1;
  wire arrdiv12_fs122_or0;
  wire arrdiv12_fs123_xor0;
  wire arrdiv12_fs123_not0;
  wire arrdiv12_fs123_and0;
  wire arrdiv12_fs123_xor1;
  wire arrdiv12_fs123_not1;
  wire arrdiv12_fs123_and1;
  wire arrdiv12_fs123_or0;
  wire arrdiv12_fs124_xor0;
  wire arrdiv12_fs124_not0;
  wire arrdiv12_fs124_and0;
  wire arrdiv12_fs124_xor1;
  wire arrdiv12_fs124_not1;
  wire arrdiv12_fs124_and1;
  wire arrdiv12_fs124_or0;
  wire arrdiv12_fs125_xor0;
  wire arrdiv12_fs125_not0;
  wire arrdiv12_fs125_and0;
  wire arrdiv12_fs125_xor1;
  wire arrdiv12_fs125_not1;
  wire arrdiv12_fs125_and1;
  wire arrdiv12_fs125_or0;
  wire arrdiv12_fs126_xor0;
  wire arrdiv12_fs126_not0;
  wire arrdiv12_fs126_and0;
  wire arrdiv12_fs126_xor1;
  wire arrdiv12_fs126_not1;
  wire arrdiv12_fs126_and1;
  wire arrdiv12_fs126_or0;
  wire arrdiv12_fs127_xor0;
  wire arrdiv12_fs127_not0;
  wire arrdiv12_fs127_and0;
  wire arrdiv12_fs127_xor1;
  wire arrdiv12_fs127_not1;
  wire arrdiv12_fs127_and1;
  wire arrdiv12_fs127_or0;
  wire arrdiv12_fs128_xor0;
  wire arrdiv12_fs128_not0;
  wire arrdiv12_fs128_and0;
  wire arrdiv12_fs128_xor1;
  wire arrdiv12_fs128_not1;
  wire arrdiv12_fs128_and1;
  wire arrdiv12_fs128_or0;
  wire arrdiv12_fs129_xor0;
  wire arrdiv12_fs129_not0;
  wire arrdiv12_fs129_and0;
  wire arrdiv12_fs129_xor1;
  wire arrdiv12_fs129_not1;
  wire arrdiv12_fs129_and1;
  wire arrdiv12_fs129_or0;
  wire arrdiv12_fs130_xor0;
  wire arrdiv12_fs130_not0;
  wire arrdiv12_fs130_and0;
  wire arrdiv12_fs130_xor1;
  wire arrdiv12_fs130_not1;
  wire arrdiv12_fs130_and1;
  wire arrdiv12_fs130_or0;
  wire arrdiv12_fs131_xor0;
  wire arrdiv12_fs131_not0;
  wire arrdiv12_fs131_and0;
  wire arrdiv12_fs131_xor1;
  wire arrdiv12_fs131_not1;
  wire arrdiv12_fs131_and1;
  wire arrdiv12_fs131_or0;
  wire arrdiv12_mux2to1110_and0;
  wire arrdiv12_mux2to1110_not0;
  wire arrdiv12_mux2to1110_and1;
  wire arrdiv12_mux2to1110_xor0;
  wire arrdiv12_mux2to1111_and0;
  wire arrdiv12_mux2to1111_not0;
  wire arrdiv12_mux2to1111_and1;
  wire arrdiv12_mux2to1111_xor0;
  wire arrdiv12_mux2to1112_and0;
  wire arrdiv12_mux2to1112_not0;
  wire arrdiv12_mux2to1112_and1;
  wire arrdiv12_mux2to1112_xor0;
  wire arrdiv12_mux2to1113_and0;
  wire arrdiv12_mux2to1113_not0;
  wire arrdiv12_mux2to1113_and1;
  wire arrdiv12_mux2to1113_xor0;
  wire arrdiv12_mux2to1114_and0;
  wire arrdiv12_mux2to1114_not0;
  wire arrdiv12_mux2to1114_and1;
  wire arrdiv12_mux2to1114_xor0;
  wire arrdiv12_mux2to1115_and0;
  wire arrdiv12_mux2to1115_not0;
  wire arrdiv12_mux2to1115_and1;
  wire arrdiv12_mux2to1115_xor0;
  wire arrdiv12_mux2to1116_and0;
  wire arrdiv12_mux2to1116_not0;
  wire arrdiv12_mux2to1116_and1;
  wire arrdiv12_mux2to1116_xor0;
  wire arrdiv12_mux2to1117_and0;
  wire arrdiv12_mux2to1117_not0;
  wire arrdiv12_mux2to1117_and1;
  wire arrdiv12_mux2to1117_xor0;
  wire arrdiv12_mux2to1118_and0;
  wire arrdiv12_mux2to1118_not0;
  wire arrdiv12_mux2to1118_and1;
  wire arrdiv12_mux2to1118_xor0;
  wire arrdiv12_mux2to1119_and0;
  wire arrdiv12_mux2to1119_not0;
  wire arrdiv12_mux2to1119_and1;
  wire arrdiv12_mux2to1119_xor0;
  wire arrdiv12_mux2to1120_and0;
  wire arrdiv12_mux2to1120_not0;
  wire arrdiv12_mux2to1120_and1;
  wire arrdiv12_mux2to1120_xor0;
  wire arrdiv12_not10;
  wire arrdiv12_fs132_xor0;
  wire arrdiv12_fs132_not0;
  wire arrdiv12_fs132_and0;
  wire arrdiv12_fs132_not1;
  wire arrdiv12_fs133_xor0;
  wire arrdiv12_fs133_not0;
  wire arrdiv12_fs133_and0;
  wire arrdiv12_fs133_xor1;
  wire arrdiv12_fs133_not1;
  wire arrdiv12_fs133_and1;
  wire arrdiv12_fs133_or0;
  wire arrdiv12_fs134_xor0;
  wire arrdiv12_fs134_not0;
  wire arrdiv12_fs134_and0;
  wire arrdiv12_fs134_xor1;
  wire arrdiv12_fs134_not1;
  wire arrdiv12_fs134_and1;
  wire arrdiv12_fs134_or0;
  wire arrdiv12_fs135_xor0;
  wire arrdiv12_fs135_not0;
  wire arrdiv12_fs135_and0;
  wire arrdiv12_fs135_xor1;
  wire arrdiv12_fs135_not1;
  wire arrdiv12_fs135_and1;
  wire arrdiv12_fs135_or0;
  wire arrdiv12_fs136_xor0;
  wire arrdiv12_fs136_not0;
  wire arrdiv12_fs136_and0;
  wire arrdiv12_fs136_xor1;
  wire arrdiv12_fs136_not1;
  wire arrdiv12_fs136_and1;
  wire arrdiv12_fs136_or0;
  wire arrdiv12_fs137_xor0;
  wire arrdiv12_fs137_not0;
  wire arrdiv12_fs137_and0;
  wire arrdiv12_fs137_xor1;
  wire arrdiv12_fs137_not1;
  wire arrdiv12_fs137_and1;
  wire arrdiv12_fs137_or0;
  wire arrdiv12_fs138_xor0;
  wire arrdiv12_fs138_not0;
  wire arrdiv12_fs138_and0;
  wire arrdiv12_fs138_xor1;
  wire arrdiv12_fs138_not1;
  wire arrdiv12_fs138_and1;
  wire arrdiv12_fs138_or0;
  wire arrdiv12_fs139_xor0;
  wire arrdiv12_fs139_not0;
  wire arrdiv12_fs139_and0;
  wire arrdiv12_fs139_xor1;
  wire arrdiv12_fs139_not1;
  wire arrdiv12_fs139_and1;
  wire arrdiv12_fs139_or0;
  wire arrdiv12_fs140_xor0;
  wire arrdiv12_fs140_not0;
  wire arrdiv12_fs140_and0;
  wire arrdiv12_fs140_xor1;
  wire arrdiv12_fs140_not1;
  wire arrdiv12_fs140_and1;
  wire arrdiv12_fs140_or0;
  wire arrdiv12_fs141_xor0;
  wire arrdiv12_fs141_not0;
  wire arrdiv12_fs141_and0;
  wire arrdiv12_fs141_xor1;
  wire arrdiv12_fs141_not1;
  wire arrdiv12_fs141_and1;
  wire arrdiv12_fs141_or0;
  wire arrdiv12_fs142_xor0;
  wire arrdiv12_fs142_not0;
  wire arrdiv12_fs142_and0;
  wire arrdiv12_fs142_xor1;
  wire arrdiv12_fs142_not1;
  wire arrdiv12_fs142_and1;
  wire arrdiv12_fs142_or0;
  wire arrdiv12_fs143_xor0;
  wire arrdiv12_fs143_not0;
  wire arrdiv12_fs143_and0;
  wire arrdiv12_fs143_xor1;
  wire arrdiv12_fs143_not1;
  wire arrdiv12_fs143_and1;
  wire arrdiv12_fs143_or0;
  wire arrdiv12_not11;

  assign arrdiv12_fs0_xor0 = a[11] ^ b[0];
  assign arrdiv12_fs0_not0 = ~a[11];
  assign arrdiv12_fs0_and0 = arrdiv12_fs0_not0 & b[0];
  assign arrdiv12_fs0_not1 = ~arrdiv12_fs0_xor0;
  assign arrdiv12_fs1_xor1 = arrdiv12_fs0_and0 ^ b[1];
  assign arrdiv12_fs1_not1 = ~b[1];
  assign arrdiv12_fs1_and1 = arrdiv12_fs1_not1 & arrdiv12_fs0_and0;
  assign arrdiv12_fs1_or0 = arrdiv12_fs1_and1 | b[1];
  assign arrdiv12_fs2_xor1 = arrdiv12_fs1_or0 ^ b[2];
  assign arrdiv12_fs2_not1 = ~b[2];
  assign arrdiv12_fs2_and1 = arrdiv12_fs2_not1 & arrdiv12_fs1_or0;
  assign arrdiv12_fs2_or0 = arrdiv12_fs2_and1 | b[2];
  assign arrdiv12_fs3_xor1 = arrdiv12_fs2_or0 ^ b[3];
  assign arrdiv12_fs3_not1 = ~b[3];
  assign arrdiv12_fs3_and1 = arrdiv12_fs3_not1 & arrdiv12_fs2_or0;
  assign arrdiv12_fs3_or0 = arrdiv12_fs3_and1 | b[3];
  assign arrdiv12_fs4_xor1 = arrdiv12_fs3_or0 ^ b[4];
  assign arrdiv12_fs4_not1 = ~b[4];
  assign arrdiv12_fs4_and1 = arrdiv12_fs4_not1 & arrdiv12_fs3_or0;
  assign arrdiv12_fs4_or0 = arrdiv12_fs4_and1 | b[4];
  assign arrdiv12_fs5_xor1 = arrdiv12_fs4_or0 ^ b[5];
  assign arrdiv12_fs5_not1 = ~b[5];
  assign arrdiv12_fs5_and1 = arrdiv12_fs5_not1 & arrdiv12_fs4_or0;
  assign arrdiv12_fs5_or0 = arrdiv12_fs5_and1 | b[5];
  assign arrdiv12_fs6_xor1 = arrdiv12_fs5_or0 ^ b[6];
  assign arrdiv12_fs6_not1 = ~b[6];
  assign arrdiv12_fs6_and1 = arrdiv12_fs6_not1 & arrdiv12_fs5_or0;
  assign arrdiv12_fs6_or0 = arrdiv12_fs6_and1 | b[6];
  assign arrdiv12_fs7_xor1 = arrdiv12_fs6_or0 ^ b[7];
  assign arrdiv12_fs7_not1 = ~b[7];
  assign arrdiv12_fs7_and1 = arrdiv12_fs7_not1 & arrdiv12_fs6_or0;
  assign arrdiv12_fs7_or0 = arrdiv12_fs7_and1 | b[7];
  assign arrdiv12_fs8_xor1 = arrdiv12_fs7_or0 ^ b[8];
  assign arrdiv12_fs8_not1 = ~b[8];
  assign arrdiv12_fs8_and1 = arrdiv12_fs8_not1 & arrdiv12_fs7_or0;
  assign arrdiv12_fs8_or0 = arrdiv12_fs8_and1 | b[8];
  assign arrdiv12_fs9_xor1 = arrdiv12_fs8_or0 ^ b[9];
  assign arrdiv12_fs9_not1 = ~b[9];
  assign arrdiv12_fs9_and1 = arrdiv12_fs9_not1 & arrdiv12_fs8_or0;
  assign arrdiv12_fs9_or0 = arrdiv12_fs9_and1 | b[9];
  assign arrdiv12_fs10_xor1 = arrdiv12_fs9_or0 ^ b[10];
  assign arrdiv12_fs10_not1 = ~b[10];
  assign arrdiv12_fs10_and1 = arrdiv12_fs10_not1 & arrdiv12_fs9_or0;
  assign arrdiv12_fs10_or0 = arrdiv12_fs10_and1 | b[10];
  assign arrdiv12_fs11_xor1 = arrdiv12_fs10_or0 ^ b[11];
  assign arrdiv12_fs11_not1 = ~b[11];
  assign arrdiv12_fs11_and1 = arrdiv12_fs11_not1 & arrdiv12_fs10_or0;
  assign arrdiv12_fs11_or0 = arrdiv12_fs11_and1 | b[11];
  assign arrdiv12_mux2to10_and0 = a[11] & arrdiv12_fs11_or0;
  assign arrdiv12_mux2to10_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to10_and1 = arrdiv12_fs0_xor0 & arrdiv12_mux2to10_not0;
  assign arrdiv12_mux2to10_xor0 = arrdiv12_mux2to10_and0 ^ arrdiv12_mux2to10_and1;
  assign arrdiv12_mux2to11_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to11_and1 = arrdiv12_fs1_xor1 & arrdiv12_mux2to11_not0;
  assign arrdiv12_mux2to12_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to12_and1 = arrdiv12_fs2_xor1 & arrdiv12_mux2to12_not0;
  assign arrdiv12_mux2to13_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to13_and1 = arrdiv12_fs3_xor1 & arrdiv12_mux2to13_not0;
  assign arrdiv12_mux2to14_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to14_and1 = arrdiv12_fs4_xor1 & arrdiv12_mux2to14_not0;
  assign arrdiv12_mux2to15_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to15_and1 = arrdiv12_fs5_xor1 & arrdiv12_mux2to15_not0;
  assign arrdiv12_mux2to16_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to16_and1 = arrdiv12_fs6_xor1 & arrdiv12_mux2to16_not0;
  assign arrdiv12_mux2to17_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to17_and1 = arrdiv12_fs7_xor1 & arrdiv12_mux2to17_not0;
  assign arrdiv12_mux2to18_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to18_and1 = arrdiv12_fs8_xor1 & arrdiv12_mux2to18_not0;
  assign arrdiv12_mux2to19_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to19_and1 = arrdiv12_fs9_xor1 & arrdiv12_mux2to19_not0;
  assign arrdiv12_mux2to110_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_mux2to110_and1 = arrdiv12_fs10_xor1 & arrdiv12_mux2to110_not0;
  assign arrdiv12_not0 = ~arrdiv12_fs11_or0;
  assign arrdiv12_fs12_xor0 = a[10] ^ b[0];
  assign arrdiv12_fs12_not0 = ~a[10];
  assign arrdiv12_fs12_and0 = arrdiv12_fs12_not0 & b[0];
  assign arrdiv12_fs12_not1 = ~arrdiv12_fs12_xor0;
  assign arrdiv12_fs13_xor0 = arrdiv12_mux2to10_xor0 ^ b[1];
  assign arrdiv12_fs13_not0 = ~arrdiv12_mux2to10_xor0;
  assign arrdiv12_fs13_and0 = arrdiv12_fs13_not0 & b[1];
  assign arrdiv12_fs13_xor1 = arrdiv12_fs12_and0 ^ arrdiv12_fs13_xor0;
  assign arrdiv12_fs13_not1 = ~arrdiv12_fs13_xor0;
  assign arrdiv12_fs13_and1 = arrdiv12_fs13_not1 & arrdiv12_fs12_and0;
  assign arrdiv12_fs13_or0 = arrdiv12_fs13_and1 | arrdiv12_fs13_and0;
  assign arrdiv12_fs14_xor0 = arrdiv12_mux2to11_and1 ^ b[2];
  assign arrdiv12_fs14_not0 = ~arrdiv12_mux2to11_and1;
  assign arrdiv12_fs14_and0 = arrdiv12_fs14_not0 & b[2];
  assign arrdiv12_fs14_xor1 = arrdiv12_fs13_or0 ^ arrdiv12_fs14_xor0;
  assign arrdiv12_fs14_not1 = ~arrdiv12_fs14_xor0;
  assign arrdiv12_fs14_and1 = arrdiv12_fs14_not1 & arrdiv12_fs13_or0;
  assign arrdiv12_fs14_or0 = arrdiv12_fs14_and1 | arrdiv12_fs14_and0;
  assign arrdiv12_fs15_xor0 = arrdiv12_mux2to12_and1 ^ b[3];
  assign arrdiv12_fs15_not0 = ~arrdiv12_mux2to12_and1;
  assign arrdiv12_fs15_and0 = arrdiv12_fs15_not0 & b[3];
  assign arrdiv12_fs15_xor1 = arrdiv12_fs14_or0 ^ arrdiv12_fs15_xor0;
  assign arrdiv12_fs15_not1 = ~arrdiv12_fs15_xor0;
  assign arrdiv12_fs15_and1 = arrdiv12_fs15_not1 & arrdiv12_fs14_or0;
  assign arrdiv12_fs15_or0 = arrdiv12_fs15_and1 | arrdiv12_fs15_and0;
  assign arrdiv12_fs16_xor0 = arrdiv12_mux2to13_and1 ^ b[4];
  assign arrdiv12_fs16_not0 = ~arrdiv12_mux2to13_and1;
  assign arrdiv12_fs16_and0 = arrdiv12_fs16_not0 & b[4];
  assign arrdiv12_fs16_xor1 = arrdiv12_fs15_or0 ^ arrdiv12_fs16_xor0;
  assign arrdiv12_fs16_not1 = ~arrdiv12_fs16_xor0;
  assign arrdiv12_fs16_and1 = arrdiv12_fs16_not1 & arrdiv12_fs15_or0;
  assign arrdiv12_fs16_or0 = arrdiv12_fs16_and1 | arrdiv12_fs16_and0;
  assign arrdiv12_fs17_xor0 = arrdiv12_mux2to14_and1 ^ b[5];
  assign arrdiv12_fs17_not0 = ~arrdiv12_mux2to14_and1;
  assign arrdiv12_fs17_and0 = arrdiv12_fs17_not0 & b[5];
  assign arrdiv12_fs17_xor1 = arrdiv12_fs16_or0 ^ arrdiv12_fs17_xor0;
  assign arrdiv12_fs17_not1 = ~arrdiv12_fs17_xor0;
  assign arrdiv12_fs17_and1 = arrdiv12_fs17_not1 & arrdiv12_fs16_or0;
  assign arrdiv12_fs17_or0 = arrdiv12_fs17_and1 | arrdiv12_fs17_and0;
  assign arrdiv12_fs18_xor0 = arrdiv12_mux2to15_and1 ^ b[6];
  assign arrdiv12_fs18_not0 = ~arrdiv12_mux2to15_and1;
  assign arrdiv12_fs18_and0 = arrdiv12_fs18_not0 & b[6];
  assign arrdiv12_fs18_xor1 = arrdiv12_fs17_or0 ^ arrdiv12_fs18_xor0;
  assign arrdiv12_fs18_not1 = ~arrdiv12_fs18_xor0;
  assign arrdiv12_fs18_and1 = arrdiv12_fs18_not1 & arrdiv12_fs17_or0;
  assign arrdiv12_fs18_or0 = arrdiv12_fs18_and1 | arrdiv12_fs18_and0;
  assign arrdiv12_fs19_xor0 = arrdiv12_mux2to16_and1 ^ b[7];
  assign arrdiv12_fs19_not0 = ~arrdiv12_mux2to16_and1;
  assign arrdiv12_fs19_and0 = arrdiv12_fs19_not0 & b[7];
  assign arrdiv12_fs19_xor1 = arrdiv12_fs18_or0 ^ arrdiv12_fs19_xor0;
  assign arrdiv12_fs19_not1 = ~arrdiv12_fs19_xor0;
  assign arrdiv12_fs19_and1 = arrdiv12_fs19_not1 & arrdiv12_fs18_or0;
  assign arrdiv12_fs19_or0 = arrdiv12_fs19_and1 | arrdiv12_fs19_and0;
  assign arrdiv12_fs20_xor0 = arrdiv12_mux2to17_and1 ^ b[8];
  assign arrdiv12_fs20_not0 = ~arrdiv12_mux2to17_and1;
  assign arrdiv12_fs20_and0 = arrdiv12_fs20_not0 & b[8];
  assign arrdiv12_fs20_xor1 = arrdiv12_fs19_or0 ^ arrdiv12_fs20_xor0;
  assign arrdiv12_fs20_not1 = ~arrdiv12_fs20_xor0;
  assign arrdiv12_fs20_and1 = arrdiv12_fs20_not1 & arrdiv12_fs19_or0;
  assign arrdiv12_fs20_or0 = arrdiv12_fs20_and1 | arrdiv12_fs20_and0;
  assign arrdiv12_fs21_xor0 = arrdiv12_mux2to18_and1 ^ b[9];
  assign arrdiv12_fs21_not0 = ~arrdiv12_mux2to18_and1;
  assign arrdiv12_fs21_and0 = arrdiv12_fs21_not0 & b[9];
  assign arrdiv12_fs21_xor1 = arrdiv12_fs20_or0 ^ arrdiv12_fs21_xor0;
  assign arrdiv12_fs21_not1 = ~arrdiv12_fs21_xor0;
  assign arrdiv12_fs21_and1 = arrdiv12_fs21_not1 & arrdiv12_fs20_or0;
  assign arrdiv12_fs21_or0 = arrdiv12_fs21_and1 | arrdiv12_fs21_and0;
  assign arrdiv12_fs22_xor0 = arrdiv12_mux2to19_and1 ^ b[10];
  assign arrdiv12_fs22_not0 = ~arrdiv12_mux2to19_and1;
  assign arrdiv12_fs22_and0 = arrdiv12_fs22_not0 & b[10];
  assign arrdiv12_fs22_xor1 = arrdiv12_fs21_or0 ^ arrdiv12_fs22_xor0;
  assign arrdiv12_fs22_not1 = ~arrdiv12_fs22_xor0;
  assign arrdiv12_fs22_and1 = arrdiv12_fs22_not1 & arrdiv12_fs21_or0;
  assign arrdiv12_fs22_or0 = arrdiv12_fs22_and1 | arrdiv12_fs22_and0;
  assign arrdiv12_fs23_xor0 = arrdiv12_mux2to110_and1 ^ b[11];
  assign arrdiv12_fs23_not0 = ~arrdiv12_mux2to110_and1;
  assign arrdiv12_fs23_and0 = arrdiv12_fs23_not0 & b[11];
  assign arrdiv12_fs23_xor1 = arrdiv12_fs22_or0 ^ arrdiv12_fs23_xor0;
  assign arrdiv12_fs23_not1 = ~arrdiv12_fs23_xor0;
  assign arrdiv12_fs23_and1 = arrdiv12_fs23_not1 & arrdiv12_fs22_or0;
  assign arrdiv12_fs23_or0 = arrdiv12_fs23_and1 | arrdiv12_fs23_and0;
  assign arrdiv12_mux2to111_and0 = a[10] & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to111_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to111_and1 = arrdiv12_fs12_xor0 & arrdiv12_mux2to111_not0;
  assign arrdiv12_mux2to111_xor0 = arrdiv12_mux2to111_and0 ^ arrdiv12_mux2to111_and1;
  assign arrdiv12_mux2to112_and0 = arrdiv12_mux2to10_xor0 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to112_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to112_and1 = arrdiv12_fs13_xor1 & arrdiv12_mux2to112_not0;
  assign arrdiv12_mux2to112_xor0 = arrdiv12_mux2to112_and0 ^ arrdiv12_mux2to112_and1;
  assign arrdiv12_mux2to113_and0 = arrdiv12_mux2to11_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to113_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to113_and1 = arrdiv12_fs14_xor1 & arrdiv12_mux2to113_not0;
  assign arrdiv12_mux2to113_xor0 = arrdiv12_mux2to113_and0 ^ arrdiv12_mux2to113_and1;
  assign arrdiv12_mux2to114_and0 = arrdiv12_mux2to12_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to114_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to114_and1 = arrdiv12_fs15_xor1 & arrdiv12_mux2to114_not0;
  assign arrdiv12_mux2to114_xor0 = arrdiv12_mux2to114_and0 ^ arrdiv12_mux2to114_and1;
  assign arrdiv12_mux2to115_and0 = arrdiv12_mux2to13_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to115_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to115_and1 = arrdiv12_fs16_xor1 & arrdiv12_mux2to115_not0;
  assign arrdiv12_mux2to115_xor0 = arrdiv12_mux2to115_and0 ^ arrdiv12_mux2to115_and1;
  assign arrdiv12_mux2to116_and0 = arrdiv12_mux2to14_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to116_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to116_and1 = arrdiv12_fs17_xor1 & arrdiv12_mux2to116_not0;
  assign arrdiv12_mux2to116_xor0 = arrdiv12_mux2to116_and0 ^ arrdiv12_mux2to116_and1;
  assign arrdiv12_mux2to117_and0 = arrdiv12_mux2to15_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to117_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to117_and1 = arrdiv12_fs18_xor1 & arrdiv12_mux2to117_not0;
  assign arrdiv12_mux2to117_xor0 = arrdiv12_mux2to117_and0 ^ arrdiv12_mux2to117_and1;
  assign arrdiv12_mux2to118_and0 = arrdiv12_mux2to16_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to118_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to118_and1 = arrdiv12_fs19_xor1 & arrdiv12_mux2to118_not0;
  assign arrdiv12_mux2to118_xor0 = arrdiv12_mux2to118_and0 ^ arrdiv12_mux2to118_and1;
  assign arrdiv12_mux2to119_and0 = arrdiv12_mux2to17_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to119_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to119_and1 = arrdiv12_fs20_xor1 & arrdiv12_mux2to119_not0;
  assign arrdiv12_mux2to119_xor0 = arrdiv12_mux2to119_and0 ^ arrdiv12_mux2to119_and1;
  assign arrdiv12_mux2to120_and0 = arrdiv12_mux2to18_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to120_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to120_and1 = arrdiv12_fs21_xor1 & arrdiv12_mux2to120_not0;
  assign arrdiv12_mux2to120_xor0 = arrdiv12_mux2to120_and0 ^ arrdiv12_mux2to120_and1;
  assign arrdiv12_mux2to121_and0 = arrdiv12_mux2to19_and1 & arrdiv12_fs23_or0;
  assign arrdiv12_mux2to121_not0 = ~arrdiv12_fs23_or0;
  assign arrdiv12_mux2to121_and1 = arrdiv12_fs22_xor1 & arrdiv12_mux2to121_not0;
  assign arrdiv12_mux2to121_xor0 = arrdiv12_mux2to121_and0 ^ arrdiv12_mux2to121_and1;
  assign arrdiv12_not1 = ~arrdiv12_fs23_or0;
  assign arrdiv12_fs24_xor0 = a[9] ^ b[0];
  assign arrdiv12_fs24_not0 = ~a[9];
  assign arrdiv12_fs24_and0 = arrdiv12_fs24_not0 & b[0];
  assign arrdiv12_fs24_not1 = ~arrdiv12_fs24_xor0;
  assign arrdiv12_fs25_xor0 = arrdiv12_mux2to111_xor0 ^ b[1];
  assign arrdiv12_fs25_not0 = ~arrdiv12_mux2to111_xor0;
  assign arrdiv12_fs25_and0 = arrdiv12_fs25_not0 & b[1];
  assign arrdiv12_fs25_xor1 = arrdiv12_fs24_and0 ^ arrdiv12_fs25_xor0;
  assign arrdiv12_fs25_not1 = ~arrdiv12_fs25_xor0;
  assign arrdiv12_fs25_and1 = arrdiv12_fs25_not1 & arrdiv12_fs24_and0;
  assign arrdiv12_fs25_or0 = arrdiv12_fs25_and1 | arrdiv12_fs25_and0;
  assign arrdiv12_fs26_xor0 = arrdiv12_mux2to112_xor0 ^ b[2];
  assign arrdiv12_fs26_not0 = ~arrdiv12_mux2to112_xor0;
  assign arrdiv12_fs26_and0 = arrdiv12_fs26_not0 & b[2];
  assign arrdiv12_fs26_xor1 = arrdiv12_fs25_or0 ^ arrdiv12_fs26_xor0;
  assign arrdiv12_fs26_not1 = ~arrdiv12_fs26_xor0;
  assign arrdiv12_fs26_and1 = arrdiv12_fs26_not1 & arrdiv12_fs25_or0;
  assign arrdiv12_fs26_or0 = arrdiv12_fs26_and1 | arrdiv12_fs26_and0;
  assign arrdiv12_fs27_xor0 = arrdiv12_mux2to113_xor0 ^ b[3];
  assign arrdiv12_fs27_not0 = ~arrdiv12_mux2to113_xor0;
  assign arrdiv12_fs27_and0 = arrdiv12_fs27_not0 & b[3];
  assign arrdiv12_fs27_xor1 = arrdiv12_fs26_or0 ^ arrdiv12_fs27_xor0;
  assign arrdiv12_fs27_not1 = ~arrdiv12_fs27_xor0;
  assign arrdiv12_fs27_and1 = arrdiv12_fs27_not1 & arrdiv12_fs26_or0;
  assign arrdiv12_fs27_or0 = arrdiv12_fs27_and1 | arrdiv12_fs27_and0;
  assign arrdiv12_fs28_xor0 = arrdiv12_mux2to114_xor0 ^ b[4];
  assign arrdiv12_fs28_not0 = ~arrdiv12_mux2to114_xor0;
  assign arrdiv12_fs28_and0 = arrdiv12_fs28_not0 & b[4];
  assign arrdiv12_fs28_xor1 = arrdiv12_fs27_or0 ^ arrdiv12_fs28_xor0;
  assign arrdiv12_fs28_not1 = ~arrdiv12_fs28_xor0;
  assign arrdiv12_fs28_and1 = arrdiv12_fs28_not1 & arrdiv12_fs27_or0;
  assign arrdiv12_fs28_or0 = arrdiv12_fs28_and1 | arrdiv12_fs28_and0;
  assign arrdiv12_fs29_xor0 = arrdiv12_mux2to115_xor0 ^ b[5];
  assign arrdiv12_fs29_not0 = ~arrdiv12_mux2to115_xor0;
  assign arrdiv12_fs29_and0 = arrdiv12_fs29_not0 & b[5];
  assign arrdiv12_fs29_xor1 = arrdiv12_fs28_or0 ^ arrdiv12_fs29_xor0;
  assign arrdiv12_fs29_not1 = ~arrdiv12_fs29_xor0;
  assign arrdiv12_fs29_and1 = arrdiv12_fs29_not1 & arrdiv12_fs28_or0;
  assign arrdiv12_fs29_or0 = arrdiv12_fs29_and1 | arrdiv12_fs29_and0;
  assign arrdiv12_fs30_xor0 = arrdiv12_mux2to116_xor0 ^ b[6];
  assign arrdiv12_fs30_not0 = ~arrdiv12_mux2to116_xor0;
  assign arrdiv12_fs30_and0 = arrdiv12_fs30_not0 & b[6];
  assign arrdiv12_fs30_xor1 = arrdiv12_fs29_or0 ^ arrdiv12_fs30_xor0;
  assign arrdiv12_fs30_not1 = ~arrdiv12_fs30_xor0;
  assign arrdiv12_fs30_and1 = arrdiv12_fs30_not1 & arrdiv12_fs29_or0;
  assign arrdiv12_fs30_or0 = arrdiv12_fs30_and1 | arrdiv12_fs30_and0;
  assign arrdiv12_fs31_xor0 = arrdiv12_mux2to117_xor0 ^ b[7];
  assign arrdiv12_fs31_not0 = ~arrdiv12_mux2to117_xor0;
  assign arrdiv12_fs31_and0 = arrdiv12_fs31_not0 & b[7];
  assign arrdiv12_fs31_xor1 = arrdiv12_fs30_or0 ^ arrdiv12_fs31_xor0;
  assign arrdiv12_fs31_not1 = ~arrdiv12_fs31_xor0;
  assign arrdiv12_fs31_and1 = arrdiv12_fs31_not1 & arrdiv12_fs30_or0;
  assign arrdiv12_fs31_or0 = arrdiv12_fs31_and1 | arrdiv12_fs31_and0;
  assign arrdiv12_fs32_xor0 = arrdiv12_mux2to118_xor0 ^ b[8];
  assign arrdiv12_fs32_not0 = ~arrdiv12_mux2to118_xor0;
  assign arrdiv12_fs32_and0 = arrdiv12_fs32_not0 & b[8];
  assign arrdiv12_fs32_xor1 = arrdiv12_fs31_or0 ^ arrdiv12_fs32_xor0;
  assign arrdiv12_fs32_not1 = ~arrdiv12_fs32_xor0;
  assign arrdiv12_fs32_and1 = arrdiv12_fs32_not1 & arrdiv12_fs31_or0;
  assign arrdiv12_fs32_or0 = arrdiv12_fs32_and1 | arrdiv12_fs32_and0;
  assign arrdiv12_fs33_xor0 = arrdiv12_mux2to119_xor0 ^ b[9];
  assign arrdiv12_fs33_not0 = ~arrdiv12_mux2to119_xor0;
  assign arrdiv12_fs33_and0 = arrdiv12_fs33_not0 & b[9];
  assign arrdiv12_fs33_xor1 = arrdiv12_fs32_or0 ^ arrdiv12_fs33_xor0;
  assign arrdiv12_fs33_not1 = ~arrdiv12_fs33_xor0;
  assign arrdiv12_fs33_and1 = arrdiv12_fs33_not1 & arrdiv12_fs32_or0;
  assign arrdiv12_fs33_or0 = arrdiv12_fs33_and1 | arrdiv12_fs33_and0;
  assign arrdiv12_fs34_xor0 = arrdiv12_mux2to120_xor0 ^ b[10];
  assign arrdiv12_fs34_not0 = ~arrdiv12_mux2to120_xor0;
  assign arrdiv12_fs34_and0 = arrdiv12_fs34_not0 & b[10];
  assign arrdiv12_fs34_xor1 = arrdiv12_fs33_or0 ^ arrdiv12_fs34_xor0;
  assign arrdiv12_fs34_not1 = ~arrdiv12_fs34_xor0;
  assign arrdiv12_fs34_and1 = arrdiv12_fs34_not1 & arrdiv12_fs33_or0;
  assign arrdiv12_fs34_or0 = arrdiv12_fs34_and1 | arrdiv12_fs34_and0;
  assign arrdiv12_fs35_xor0 = arrdiv12_mux2to121_xor0 ^ b[11];
  assign arrdiv12_fs35_not0 = ~arrdiv12_mux2to121_xor0;
  assign arrdiv12_fs35_and0 = arrdiv12_fs35_not0 & b[11];
  assign arrdiv12_fs35_xor1 = arrdiv12_fs34_or0 ^ arrdiv12_fs35_xor0;
  assign arrdiv12_fs35_not1 = ~arrdiv12_fs35_xor0;
  assign arrdiv12_fs35_and1 = arrdiv12_fs35_not1 & arrdiv12_fs34_or0;
  assign arrdiv12_fs35_or0 = arrdiv12_fs35_and1 | arrdiv12_fs35_and0;
  assign arrdiv12_mux2to122_and0 = a[9] & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to122_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to122_and1 = arrdiv12_fs24_xor0 & arrdiv12_mux2to122_not0;
  assign arrdiv12_mux2to122_xor0 = arrdiv12_mux2to122_and0 ^ arrdiv12_mux2to122_and1;
  assign arrdiv12_mux2to123_and0 = arrdiv12_mux2to111_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to123_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to123_and1 = arrdiv12_fs25_xor1 & arrdiv12_mux2to123_not0;
  assign arrdiv12_mux2to123_xor0 = arrdiv12_mux2to123_and0 ^ arrdiv12_mux2to123_and1;
  assign arrdiv12_mux2to124_and0 = arrdiv12_mux2to112_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to124_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to124_and1 = arrdiv12_fs26_xor1 & arrdiv12_mux2to124_not0;
  assign arrdiv12_mux2to124_xor0 = arrdiv12_mux2to124_and0 ^ arrdiv12_mux2to124_and1;
  assign arrdiv12_mux2to125_and0 = arrdiv12_mux2to113_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to125_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to125_and1 = arrdiv12_fs27_xor1 & arrdiv12_mux2to125_not0;
  assign arrdiv12_mux2to125_xor0 = arrdiv12_mux2to125_and0 ^ arrdiv12_mux2to125_and1;
  assign arrdiv12_mux2to126_and0 = arrdiv12_mux2to114_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to126_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to126_and1 = arrdiv12_fs28_xor1 & arrdiv12_mux2to126_not0;
  assign arrdiv12_mux2to126_xor0 = arrdiv12_mux2to126_and0 ^ arrdiv12_mux2to126_and1;
  assign arrdiv12_mux2to127_and0 = arrdiv12_mux2to115_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to127_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to127_and1 = arrdiv12_fs29_xor1 & arrdiv12_mux2to127_not0;
  assign arrdiv12_mux2to127_xor0 = arrdiv12_mux2to127_and0 ^ arrdiv12_mux2to127_and1;
  assign arrdiv12_mux2to128_and0 = arrdiv12_mux2to116_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to128_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to128_and1 = arrdiv12_fs30_xor1 & arrdiv12_mux2to128_not0;
  assign arrdiv12_mux2to128_xor0 = arrdiv12_mux2to128_and0 ^ arrdiv12_mux2to128_and1;
  assign arrdiv12_mux2to129_and0 = arrdiv12_mux2to117_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to129_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to129_and1 = arrdiv12_fs31_xor1 & arrdiv12_mux2to129_not0;
  assign arrdiv12_mux2to129_xor0 = arrdiv12_mux2to129_and0 ^ arrdiv12_mux2to129_and1;
  assign arrdiv12_mux2to130_and0 = arrdiv12_mux2to118_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to130_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to130_and1 = arrdiv12_fs32_xor1 & arrdiv12_mux2to130_not0;
  assign arrdiv12_mux2to130_xor0 = arrdiv12_mux2to130_and0 ^ arrdiv12_mux2to130_and1;
  assign arrdiv12_mux2to131_and0 = arrdiv12_mux2to119_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to131_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to131_and1 = arrdiv12_fs33_xor1 & arrdiv12_mux2to131_not0;
  assign arrdiv12_mux2to131_xor0 = arrdiv12_mux2to131_and0 ^ arrdiv12_mux2to131_and1;
  assign arrdiv12_mux2to132_and0 = arrdiv12_mux2to120_xor0 & arrdiv12_fs35_or0;
  assign arrdiv12_mux2to132_not0 = ~arrdiv12_fs35_or0;
  assign arrdiv12_mux2to132_and1 = arrdiv12_fs34_xor1 & arrdiv12_mux2to132_not0;
  assign arrdiv12_mux2to132_xor0 = arrdiv12_mux2to132_and0 ^ arrdiv12_mux2to132_and1;
  assign arrdiv12_not2 = ~arrdiv12_fs35_or0;
  assign arrdiv12_fs36_xor0 = a[8] ^ b[0];
  assign arrdiv12_fs36_not0 = ~a[8];
  assign arrdiv12_fs36_and0 = arrdiv12_fs36_not0 & b[0];
  assign arrdiv12_fs36_not1 = ~arrdiv12_fs36_xor0;
  assign arrdiv12_fs37_xor0 = arrdiv12_mux2to122_xor0 ^ b[1];
  assign arrdiv12_fs37_not0 = ~arrdiv12_mux2to122_xor0;
  assign arrdiv12_fs37_and0 = arrdiv12_fs37_not0 & b[1];
  assign arrdiv12_fs37_xor1 = arrdiv12_fs36_and0 ^ arrdiv12_fs37_xor0;
  assign arrdiv12_fs37_not1 = ~arrdiv12_fs37_xor0;
  assign arrdiv12_fs37_and1 = arrdiv12_fs37_not1 & arrdiv12_fs36_and0;
  assign arrdiv12_fs37_or0 = arrdiv12_fs37_and1 | arrdiv12_fs37_and0;
  assign arrdiv12_fs38_xor0 = arrdiv12_mux2to123_xor0 ^ b[2];
  assign arrdiv12_fs38_not0 = ~arrdiv12_mux2to123_xor0;
  assign arrdiv12_fs38_and0 = arrdiv12_fs38_not0 & b[2];
  assign arrdiv12_fs38_xor1 = arrdiv12_fs37_or0 ^ arrdiv12_fs38_xor0;
  assign arrdiv12_fs38_not1 = ~arrdiv12_fs38_xor0;
  assign arrdiv12_fs38_and1 = arrdiv12_fs38_not1 & arrdiv12_fs37_or0;
  assign arrdiv12_fs38_or0 = arrdiv12_fs38_and1 | arrdiv12_fs38_and0;
  assign arrdiv12_fs39_xor0 = arrdiv12_mux2to124_xor0 ^ b[3];
  assign arrdiv12_fs39_not0 = ~arrdiv12_mux2to124_xor0;
  assign arrdiv12_fs39_and0 = arrdiv12_fs39_not0 & b[3];
  assign arrdiv12_fs39_xor1 = arrdiv12_fs38_or0 ^ arrdiv12_fs39_xor0;
  assign arrdiv12_fs39_not1 = ~arrdiv12_fs39_xor0;
  assign arrdiv12_fs39_and1 = arrdiv12_fs39_not1 & arrdiv12_fs38_or0;
  assign arrdiv12_fs39_or0 = arrdiv12_fs39_and1 | arrdiv12_fs39_and0;
  assign arrdiv12_fs40_xor0 = arrdiv12_mux2to125_xor0 ^ b[4];
  assign arrdiv12_fs40_not0 = ~arrdiv12_mux2to125_xor0;
  assign arrdiv12_fs40_and0 = arrdiv12_fs40_not0 & b[4];
  assign arrdiv12_fs40_xor1 = arrdiv12_fs39_or0 ^ arrdiv12_fs40_xor0;
  assign arrdiv12_fs40_not1 = ~arrdiv12_fs40_xor0;
  assign arrdiv12_fs40_and1 = arrdiv12_fs40_not1 & arrdiv12_fs39_or0;
  assign arrdiv12_fs40_or0 = arrdiv12_fs40_and1 | arrdiv12_fs40_and0;
  assign arrdiv12_fs41_xor0 = arrdiv12_mux2to126_xor0 ^ b[5];
  assign arrdiv12_fs41_not0 = ~arrdiv12_mux2to126_xor0;
  assign arrdiv12_fs41_and0 = arrdiv12_fs41_not0 & b[5];
  assign arrdiv12_fs41_xor1 = arrdiv12_fs40_or0 ^ arrdiv12_fs41_xor0;
  assign arrdiv12_fs41_not1 = ~arrdiv12_fs41_xor0;
  assign arrdiv12_fs41_and1 = arrdiv12_fs41_not1 & arrdiv12_fs40_or0;
  assign arrdiv12_fs41_or0 = arrdiv12_fs41_and1 | arrdiv12_fs41_and0;
  assign arrdiv12_fs42_xor0 = arrdiv12_mux2to127_xor0 ^ b[6];
  assign arrdiv12_fs42_not0 = ~arrdiv12_mux2to127_xor0;
  assign arrdiv12_fs42_and0 = arrdiv12_fs42_not0 & b[6];
  assign arrdiv12_fs42_xor1 = arrdiv12_fs41_or0 ^ arrdiv12_fs42_xor0;
  assign arrdiv12_fs42_not1 = ~arrdiv12_fs42_xor0;
  assign arrdiv12_fs42_and1 = arrdiv12_fs42_not1 & arrdiv12_fs41_or0;
  assign arrdiv12_fs42_or0 = arrdiv12_fs42_and1 | arrdiv12_fs42_and0;
  assign arrdiv12_fs43_xor0 = arrdiv12_mux2to128_xor0 ^ b[7];
  assign arrdiv12_fs43_not0 = ~arrdiv12_mux2to128_xor0;
  assign arrdiv12_fs43_and0 = arrdiv12_fs43_not0 & b[7];
  assign arrdiv12_fs43_xor1 = arrdiv12_fs42_or0 ^ arrdiv12_fs43_xor0;
  assign arrdiv12_fs43_not1 = ~arrdiv12_fs43_xor0;
  assign arrdiv12_fs43_and1 = arrdiv12_fs43_not1 & arrdiv12_fs42_or0;
  assign arrdiv12_fs43_or0 = arrdiv12_fs43_and1 | arrdiv12_fs43_and0;
  assign arrdiv12_fs44_xor0 = arrdiv12_mux2to129_xor0 ^ b[8];
  assign arrdiv12_fs44_not0 = ~arrdiv12_mux2to129_xor0;
  assign arrdiv12_fs44_and0 = arrdiv12_fs44_not0 & b[8];
  assign arrdiv12_fs44_xor1 = arrdiv12_fs43_or0 ^ arrdiv12_fs44_xor0;
  assign arrdiv12_fs44_not1 = ~arrdiv12_fs44_xor0;
  assign arrdiv12_fs44_and1 = arrdiv12_fs44_not1 & arrdiv12_fs43_or0;
  assign arrdiv12_fs44_or0 = arrdiv12_fs44_and1 | arrdiv12_fs44_and0;
  assign arrdiv12_fs45_xor0 = arrdiv12_mux2to130_xor0 ^ b[9];
  assign arrdiv12_fs45_not0 = ~arrdiv12_mux2to130_xor0;
  assign arrdiv12_fs45_and0 = arrdiv12_fs45_not0 & b[9];
  assign arrdiv12_fs45_xor1 = arrdiv12_fs44_or0 ^ arrdiv12_fs45_xor0;
  assign arrdiv12_fs45_not1 = ~arrdiv12_fs45_xor0;
  assign arrdiv12_fs45_and1 = arrdiv12_fs45_not1 & arrdiv12_fs44_or0;
  assign arrdiv12_fs45_or0 = arrdiv12_fs45_and1 | arrdiv12_fs45_and0;
  assign arrdiv12_fs46_xor0 = arrdiv12_mux2to131_xor0 ^ b[10];
  assign arrdiv12_fs46_not0 = ~arrdiv12_mux2to131_xor0;
  assign arrdiv12_fs46_and0 = arrdiv12_fs46_not0 & b[10];
  assign arrdiv12_fs46_xor1 = arrdiv12_fs45_or0 ^ arrdiv12_fs46_xor0;
  assign arrdiv12_fs46_not1 = ~arrdiv12_fs46_xor0;
  assign arrdiv12_fs46_and1 = arrdiv12_fs46_not1 & arrdiv12_fs45_or0;
  assign arrdiv12_fs46_or0 = arrdiv12_fs46_and1 | arrdiv12_fs46_and0;
  assign arrdiv12_fs47_xor0 = arrdiv12_mux2to132_xor0 ^ b[11];
  assign arrdiv12_fs47_not0 = ~arrdiv12_mux2to132_xor0;
  assign arrdiv12_fs47_and0 = arrdiv12_fs47_not0 & b[11];
  assign arrdiv12_fs47_xor1 = arrdiv12_fs46_or0 ^ arrdiv12_fs47_xor0;
  assign arrdiv12_fs47_not1 = ~arrdiv12_fs47_xor0;
  assign arrdiv12_fs47_and1 = arrdiv12_fs47_not1 & arrdiv12_fs46_or0;
  assign arrdiv12_fs47_or0 = arrdiv12_fs47_and1 | arrdiv12_fs47_and0;
  assign arrdiv12_mux2to133_and0 = a[8] & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to133_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to133_and1 = arrdiv12_fs36_xor0 & arrdiv12_mux2to133_not0;
  assign arrdiv12_mux2to133_xor0 = arrdiv12_mux2to133_and0 ^ arrdiv12_mux2to133_and1;
  assign arrdiv12_mux2to134_and0 = arrdiv12_mux2to122_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to134_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to134_and1 = arrdiv12_fs37_xor1 & arrdiv12_mux2to134_not0;
  assign arrdiv12_mux2to134_xor0 = arrdiv12_mux2to134_and0 ^ arrdiv12_mux2to134_and1;
  assign arrdiv12_mux2to135_and0 = arrdiv12_mux2to123_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to135_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to135_and1 = arrdiv12_fs38_xor1 & arrdiv12_mux2to135_not0;
  assign arrdiv12_mux2to135_xor0 = arrdiv12_mux2to135_and0 ^ arrdiv12_mux2to135_and1;
  assign arrdiv12_mux2to136_and0 = arrdiv12_mux2to124_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to136_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to136_and1 = arrdiv12_fs39_xor1 & arrdiv12_mux2to136_not0;
  assign arrdiv12_mux2to136_xor0 = arrdiv12_mux2to136_and0 ^ arrdiv12_mux2to136_and1;
  assign arrdiv12_mux2to137_and0 = arrdiv12_mux2to125_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to137_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to137_and1 = arrdiv12_fs40_xor1 & arrdiv12_mux2to137_not0;
  assign arrdiv12_mux2to137_xor0 = arrdiv12_mux2to137_and0 ^ arrdiv12_mux2to137_and1;
  assign arrdiv12_mux2to138_and0 = arrdiv12_mux2to126_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to138_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to138_and1 = arrdiv12_fs41_xor1 & arrdiv12_mux2to138_not0;
  assign arrdiv12_mux2to138_xor0 = arrdiv12_mux2to138_and0 ^ arrdiv12_mux2to138_and1;
  assign arrdiv12_mux2to139_and0 = arrdiv12_mux2to127_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to139_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to139_and1 = arrdiv12_fs42_xor1 & arrdiv12_mux2to139_not0;
  assign arrdiv12_mux2to139_xor0 = arrdiv12_mux2to139_and0 ^ arrdiv12_mux2to139_and1;
  assign arrdiv12_mux2to140_and0 = arrdiv12_mux2to128_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to140_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to140_and1 = arrdiv12_fs43_xor1 & arrdiv12_mux2to140_not0;
  assign arrdiv12_mux2to140_xor0 = arrdiv12_mux2to140_and0 ^ arrdiv12_mux2to140_and1;
  assign arrdiv12_mux2to141_and0 = arrdiv12_mux2to129_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to141_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to141_and1 = arrdiv12_fs44_xor1 & arrdiv12_mux2to141_not0;
  assign arrdiv12_mux2to141_xor0 = arrdiv12_mux2to141_and0 ^ arrdiv12_mux2to141_and1;
  assign arrdiv12_mux2to142_and0 = arrdiv12_mux2to130_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to142_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to142_and1 = arrdiv12_fs45_xor1 & arrdiv12_mux2to142_not0;
  assign arrdiv12_mux2to142_xor0 = arrdiv12_mux2to142_and0 ^ arrdiv12_mux2to142_and1;
  assign arrdiv12_mux2to143_and0 = arrdiv12_mux2to131_xor0 & arrdiv12_fs47_or0;
  assign arrdiv12_mux2to143_not0 = ~arrdiv12_fs47_or0;
  assign arrdiv12_mux2to143_and1 = arrdiv12_fs46_xor1 & arrdiv12_mux2to143_not0;
  assign arrdiv12_mux2to143_xor0 = arrdiv12_mux2to143_and0 ^ arrdiv12_mux2to143_and1;
  assign arrdiv12_not3 = ~arrdiv12_fs47_or0;
  assign arrdiv12_fs48_xor0 = a[7] ^ b[0];
  assign arrdiv12_fs48_not0 = ~a[7];
  assign arrdiv12_fs48_and0 = arrdiv12_fs48_not0 & b[0];
  assign arrdiv12_fs48_not1 = ~arrdiv12_fs48_xor0;
  assign arrdiv12_fs49_xor0 = arrdiv12_mux2to133_xor0 ^ b[1];
  assign arrdiv12_fs49_not0 = ~arrdiv12_mux2to133_xor0;
  assign arrdiv12_fs49_and0 = arrdiv12_fs49_not0 & b[1];
  assign arrdiv12_fs49_xor1 = arrdiv12_fs48_and0 ^ arrdiv12_fs49_xor0;
  assign arrdiv12_fs49_not1 = ~arrdiv12_fs49_xor0;
  assign arrdiv12_fs49_and1 = arrdiv12_fs49_not1 & arrdiv12_fs48_and0;
  assign arrdiv12_fs49_or0 = arrdiv12_fs49_and1 | arrdiv12_fs49_and0;
  assign arrdiv12_fs50_xor0 = arrdiv12_mux2to134_xor0 ^ b[2];
  assign arrdiv12_fs50_not0 = ~arrdiv12_mux2to134_xor0;
  assign arrdiv12_fs50_and0 = arrdiv12_fs50_not0 & b[2];
  assign arrdiv12_fs50_xor1 = arrdiv12_fs49_or0 ^ arrdiv12_fs50_xor0;
  assign arrdiv12_fs50_not1 = ~arrdiv12_fs50_xor0;
  assign arrdiv12_fs50_and1 = arrdiv12_fs50_not1 & arrdiv12_fs49_or0;
  assign arrdiv12_fs50_or0 = arrdiv12_fs50_and1 | arrdiv12_fs50_and0;
  assign arrdiv12_fs51_xor0 = arrdiv12_mux2to135_xor0 ^ b[3];
  assign arrdiv12_fs51_not0 = ~arrdiv12_mux2to135_xor0;
  assign arrdiv12_fs51_and0 = arrdiv12_fs51_not0 & b[3];
  assign arrdiv12_fs51_xor1 = arrdiv12_fs50_or0 ^ arrdiv12_fs51_xor0;
  assign arrdiv12_fs51_not1 = ~arrdiv12_fs51_xor0;
  assign arrdiv12_fs51_and1 = arrdiv12_fs51_not1 & arrdiv12_fs50_or0;
  assign arrdiv12_fs51_or0 = arrdiv12_fs51_and1 | arrdiv12_fs51_and0;
  assign arrdiv12_fs52_xor0 = arrdiv12_mux2to136_xor0 ^ b[4];
  assign arrdiv12_fs52_not0 = ~arrdiv12_mux2to136_xor0;
  assign arrdiv12_fs52_and0 = arrdiv12_fs52_not0 & b[4];
  assign arrdiv12_fs52_xor1 = arrdiv12_fs51_or0 ^ arrdiv12_fs52_xor0;
  assign arrdiv12_fs52_not1 = ~arrdiv12_fs52_xor0;
  assign arrdiv12_fs52_and1 = arrdiv12_fs52_not1 & arrdiv12_fs51_or0;
  assign arrdiv12_fs52_or0 = arrdiv12_fs52_and1 | arrdiv12_fs52_and0;
  assign arrdiv12_fs53_xor0 = arrdiv12_mux2to137_xor0 ^ b[5];
  assign arrdiv12_fs53_not0 = ~arrdiv12_mux2to137_xor0;
  assign arrdiv12_fs53_and0 = arrdiv12_fs53_not0 & b[5];
  assign arrdiv12_fs53_xor1 = arrdiv12_fs52_or0 ^ arrdiv12_fs53_xor0;
  assign arrdiv12_fs53_not1 = ~arrdiv12_fs53_xor0;
  assign arrdiv12_fs53_and1 = arrdiv12_fs53_not1 & arrdiv12_fs52_or0;
  assign arrdiv12_fs53_or0 = arrdiv12_fs53_and1 | arrdiv12_fs53_and0;
  assign arrdiv12_fs54_xor0 = arrdiv12_mux2to138_xor0 ^ b[6];
  assign arrdiv12_fs54_not0 = ~arrdiv12_mux2to138_xor0;
  assign arrdiv12_fs54_and0 = arrdiv12_fs54_not0 & b[6];
  assign arrdiv12_fs54_xor1 = arrdiv12_fs53_or0 ^ arrdiv12_fs54_xor0;
  assign arrdiv12_fs54_not1 = ~arrdiv12_fs54_xor0;
  assign arrdiv12_fs54_and1 = arrdiv12_fs54_not1 & arrdiv12_fs53_or0;
  assign arrdiv12_fs54_or0 = arrdiv12_fs54_and1 | arrdiv12_fs54_and0;
  assign arrdiv12_fs55_xor0 = arrdiv12_mux2to139_xor0 ^ b[7];
  assign arrdiv12_fs55_not0 = ~arrdiv12_mux2to139_xor0;
  assign arrdiv12_fs55_and0 = arrdiv12_fs55_not0 & b[7];
  assign arrdiv12_fs55_xor1 = arrdiv12_fs54_or0 ^ arrdiv12_fs55_xor0;
  assign arrdiv12_fs55_not1 = ~arrdiv12_fs55_xor0;
  assign arrdiv12_fs55_and1 = arrdiv12_fs55_not1 & arrdiv12_fs54_or0;
  assign arrdiv12_fs55_or0 = arrdiv12_fs55_and1 | arrdiv12_fs55_and0;
  assign arrdiv12_fs56_xor0 = arrdiv12_mux2to140_xor0 ^ b[8];
  assign arrdiv12_fs56_not0 = ~arrdiv12_mux2to140_xor0;
  assign arrdiv12_fs56_and0 = arrdiv12_fs56_not0 & b[8];
  assign arrdiv12_fs56_xor1 = arrdiv12_fs55_or0 ^ arrdiv12_fs56_xor0;
  assign arrdiv12_fs56_not1 = ~arrdiv12_fs56_xor0;
  assign arrdiv12_fs56_and1 = arrdiv12_fs56_not1 & arrdiv12_fs55_or0;
  assign arrdiv12_fs56_or0 = arrdiv12_fs56_and1 | arrdiv12_fs56_and0;
  assign arrdiv12_fs57_xor0 = arrdiv12_mux2to141_xor0 ^ b[9];
  assign arrdiv12_fs57_not0 = ~arrdiv12_mux2to141_xor0;
  assign arrdiv12_fs57_and0 = arrdiv12_fs57_not0 & b[9];
  assign arrdiv12_fs57_xor1 = arrdiv12_fs56_or0 ^ arrdiv12_fs57_xor0;
  assign arrdiv12_fs57_not1 = ~arrdiv12_fs57_xor0;
  assign arrdiv12_fs57_and1 = arrdiv12_fs57_not1 & arrdiv12_fs56_or0;
  assign arrdiv12_fs57_or0 = arrdiv12_fs57_and1 | arrdiv12_fs57_and0;
  assign arrdiv12_fs58_xor0 = arrdiv12_mux2to142_xor0 ^ b[10];
  assign arrdiv12_fs58_not0 = ~arrdiv12_mux2to142_xor0;
  assign arrdiv12_fs58_and0 = arrdiv12_fs58_not0 & b[10];
  assign arrdiv12_fs58_xor1 = arrdiv12_fs57_or0 ^ arrdiv12_fs58_xor0;
  assign arrdiv12_fs58_not1 = ~arrdiv12_fs58_xor0;
  assign arrdiv12_fs58_and1 = arrdiv12_fs58_not1 & arrdiv12_fs57_or0;
  assign arrdiv12_fs58_or0 = arrdiv12_fs58_and1 | arrdiv12_fs58_and0;
  assign arrdiv12_fs59_xor0 = arrdiv12_mux2to143_xor0 ^ b[11];
  assign arrdiv12_fs59_not0 = ~arrdiv12_mux2to143_xor0;
  assign arrdiv12_fs59_and0 = arrdiv12_fs59_not0 & b[11];
  assign arrdiv12_fs59_xor1 = arrdiv12_fs58_or0 ^ arrdiv12_fs59_xor0;
  assign arrdiv12_fs59_not1 = ~arrdiv12_fs59_xor0;
  assign arrdiv12_fs59_and1 = arrdiv12_fs59_not1 & arrdiv12_fs58_or0;
  assign arrdiv12_fs59_or0 = arrdiv12_fs59_and1 | arrdiv12_fs59_and0;
  assign arrdiv12_mux2to144_and0 = a[7] & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to144_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to144_and1 = arrdiv12_fs48_xor0 & arrdiv12_mux2to144_not0;
  assign arrdiv12_mux2to144_xor0 = arrdiv12_mux2to144_and0 ^ arrdiv12_mux2to144_and1;
  assign arrdiv12_mux2to145_and0 = arrdiv12_mux2to133_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to145_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to145_and1 = arrdiv12_fs49_xor1 & arrdiv12_mux2to145_not0;
  assign arrdiv12_mux2to145_xor0 = arrdiv12_mux2to145_and0 ^ arrdiv12_mux2to145_and1;
  assign arrdiv12_mux2to146_and0 = arrdiv12_mux2to134_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to146_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to146_and1 = arrdiv12_fs50_xor1 & arrdiv12_mux2to146_not0;
  assign arrdiv12_mux2to146_xor0 = arrdiv12_mux2to146_and0 ^ arrdiv12_mux2to146_and1;
  assign arrdiv12_mux2to147_and0 = arrdiv12_mux2to135_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to147_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to147_and1 = arrdiv12_fs51_xor1 & arrdiv12_mux2to147_not0;
  assign arrdiv12_mux2to147_xor0 = arrdiv12_mux2to147_and0 ^ arrdiv12_mux2to147_and1;
  assign arrdiv12_mux2to148_and0 = arrdiv12_mux2to136_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to148_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to148_and1 = arrdiv12_fs52_xor1 & arrdiv12_mux2to148_not0;
  assign arrdiv12_mux2to148_xor0 = arrdiv12_mux2to148_and0 ^ arrdiv12_mux2to148_and1;
  assign arrdiv12_mux2to149_and0 = arrdiv12_mux2to137_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to149_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to149_and1 = arrdiv12_fs53_xor1 & arrdiv12_mux2to149_not0;
  assign arrdiv12_mux2to149_xor0 = arrdiv12_mux2to149_and0 ^ arrdiv12_mux2to149_and1;
  assign arrdiv12_mux2to150_and0 = arrdiv12_mux2to138_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to150_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to150_and1 = arrdiv12_fs54_xor1 & arrdiv12_mux2to150_not0;
  assign arrdiv12_mux2to150_xor0 = arrdiv12_mux2to150_and0 ^ arrdiv12_mux2to150_and1;
  assign arrdiv12_mux2to151_and0 = arrdiv12_mux2to139_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to151_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to151_and1 = arrdiv12_fs55_xor1 & arrdiv12_mux2to151_not0;
  assign arrdiv12_mux2to151_xor0 = arrdiv12_mux2to151_and0 ^ arrdiv12_mux2to151_and1;
  assign arrdiv12_mux2to152_and0 = arrdiv12_mux2to140_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to152_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to152_and1 = arrdiv12_fs56_xor1 & arrdiv12_mux2to152_not0;
  assign arrdiv12_mux2to152_xor0 = arrdiv12_mux2to152_and0 ^ arrdiv12_mux2to152_and1;
  assign arrdiv12_mux2to153_and0 = arrdiv12_mux2to141_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to153_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to153_and1 = arrdiv12_fs57_xor1 & arrdiv12_mux2to153_not0;
  assign arrdiv12_mux2to153_xor0 = arrdiv12_mux2to153_and0 ^ arrdiv12_mux2to153_and1;
  assign arrdiv12_mux2to154_and0 = arrdiv12_mux2to142_xor0 & arrdiv12_fs59_or0;
  assign arrdiv12_mux2to154_not0 = ~arrdiv12_fs59_or0;
  assign arrdiv12_mux2to154_and1 = arrdiv12_fs58_xor1 & arrdiv12_mux2to154_not0;
  assign arrdiv12_mux2to154_xor0 = arrdiv12_mux2to154_and0 ^ arrdiv12_mux2to154_and1;
  assign arrdiv12_not4 = ~arrdiv12_fs59_or0;
  assign arrdiv12_fs60_xor0 = a[6] ^ b[0];
  assign arrdiv12_fs60_not0 = ~a[6];
  assign arrdiv12_fs60_and0 = arrdiv12_fs60_not0 & b[0];
  assign arrdiv12_fs60_not1 = ~arrdiv12_fs60_xor0;
  assign arrdiv12_fs61_xor0 = arrdiv12_mux2to144_xor0 ^ b[1];
  assign arrdiv12_fs61_not0 = ~arrdiv12_mux2to144_xor0;
  assign arrdiv12_fs61_and0 = arrdiv12_fs61_not0 & b[1];
  assign arrdiv12_fs61_xor1 = arrdiv12_fs60_and0 ^ arrdiv12_fs61_xor0;
  assign arrdiv12_fs61_not1 = ~arrdiv12_fs61_xor0;
  assign arrdiv12_fs61_and1 = arrdiv12_fs61_not1 & arrdiv12_fs60_and0;
  assign arrdiv12_fs61_or0 = arrdiv12_fs61_and1 | arrdiv12_fs61_and0;
  assign arrdiv12_fs62_xor0 = arrdiv12_mux2to145_xor0 ^ b[2];
  assign arrdiv12_fs62_not0 = ~arrdiv12_mux2to145_xor0;
  assign arrdiv12_fs62_and0 = arrdiv12_fs62_not0 & b[2];
  assign arrdiv12_fs62_xor1 = arrdiv12_fs61_or0 ^ arrdiv12_fs62_xor0;
  assign arrdiv12_fs62_not1 = ~arrdiv12_fs62_xor0;
  assign arrdiv12_fs62_and1 = arrdiv12_fs62_not1 & arrdiv12_fs61_or0;
  assign arrdiv12_fs62_or0 = arrdiv12_fs62_and1 | arrdiv12_fs62_and0;
  assign arrdiv12_fs63_xor0 = arrdiv12_mux2to146_xor0 ^ b[3];
  assign arrdiv12_fs63_not0 = ~arrdiv12_mux2to146_xor0;
  assign arrdiv12_fs63_and0 = arrdiv12_fs63_not0 & b[3];
  assign arrdiv12_fs63_xor1 = arrdiv12_fs62_or0 ^ arrdiv12_fs63_xor0;
  assign arrdiv12_fs63_not1 = ~arrdiv12_fs63_xor0;
  assign arrdiv12_fs63_and1 = arrdiv12_fs63_not1 & arrdiv12_fs62_or0;
  assign arrdiv12_fs63_or0 = arrdiv12_fs63_and1 | arrdiv12_fs63_and0;
  assign arrdiv12_fs64_xor0 = arrdiv12_mux2to147_xor0 ^ b[4];
  assign arrdiv12_fs64_not0 = ~arrdiv12_mux2to147_xor0;
  assign arrdiv12_fs64_and0 = arrdiv12_fs64_not0 & b[4];
  assign arrdiv12_fs64_xor1 = arrdiv12_fs63_or0 ^ arrdiv12_fs64_xor0;
  assign arrdiv12_fs64_not1 = ~arrdiv12_fs64_xor0;
  assign arrdiv12_fs64_and1 = arrdiv12_fs64_not1 & arrdiv12_fs63_or0;
  assign arrdiv12_fs64_or0 = arrdiv12_fs64_and1 | arrdiv12_fs64_and0;
  assign arrdiv12_fs65_xor0 = arrdiv12_mux2to148_xor0 ^ b[5];
  assign arrdiv12_fs65_not0 = ~arrdiv12_mux2to148_xor0;
  assign arrdiv12_fs65_and0 = arrdiv12_fs65_not0 & b[5];
  assign arrdiv12_fs65_xor1 = arrdiv12_fs64_or0 ^ arrdiv12_fs65_xor0;
  assign arrdiv12_fs65_not1 = ~arrdiv12_fs65_xor0;
  assign arrdiv12_fs65_and1 = arrdiv12_fs65_not1 & arrdiv12_fs64_or0;
  assign arrdiv12_fs65_or0 = arrdiv12_fs65_and1 | arrdiv12_fs65_and0;
  assign arrdiv12_fs66_xor0 = arrdiv12_mux2to149_xor0 ^ b[6];
  assign arrdiv12_fs66_not0 = ~arrdiv12_mux2to149_xor0;
  assign arrdiv12_fs66_and0 = arrdiv12_fs66_not0 & b[6];
  assign arrdiv12_fs66_xor1 = arrdiv12_fs65_or0 ^ arrdiv12_fs66_xor0;
  assign arrdiv12_fs66_not1 = ~arrdiv12_fs66_xor0;
  assign arrdiv12_fs66_and1 = arrdiv12_fs66_not1 & arrdiv12_fs65_or0;
  assign arrdiv12_fs66_or0 = arrdiv12_fs66_and1 | arrdiv12_fs66_and0;
  assign arrdiv12_fs67_xor0 = arrdiv12_mux2to150_xor0 ^ b[7];
  assign arrdiv12_fs67_not0 = ~arrdiv12_mux2to150_xor0;
  assign arrdiv12_fs67_and0 = arrdiv12_fs67_not0 & b[7];
  assign arrdiv12_fs67_xor1 = arrdiv12_fs66_or0 ^ arrdiv12_fs67_xor0;
  assign arrdiv12_fs67_not1 = ~arrdiv12_fs67_xor0;
  assign arrdiv12_fs67_and1 = arrdiv12_fs67_not1 & arrdiv12_fs66_or0;
  assign arrdiv12_fs67_or0 = arrdiv12_fs67_and1 | arrdiv12_fs67_and0;
  assign arrdiv12_fs68_xor0 = arrdiv12_mux2to151_xor0 ^ b[8];
  assign arrdiv12_fs68_not0 = ~arrdiv12_mux2to151_xor0;
  assign arrdiv12_fs68_and0 = arrdiv12_fs68_not0 & b[8];
  assign arrdiv12_fs68_xor1 = arrdiv12_fs67_or0 ^ arrdiv12_fs68_xor0;
  assign arrdiv12_fs68_not1 = ~arrdiv12_fs68_xor0;
  assign arrdiv12_fs68_and1 = arrdiv12_fs68_not1 & arrdiv12_fs67_or0;
  assign arrdiv12_fs68_or0 = arrdiv12_fs68_and1 | arrdiv12_fs68_and0;
  assign arrdiv12_fs69_xor0 = arrdiv12_mux2to152_xor0 ^ b[9];
  assign arrdiv12_fs69_not0 = ~arrdiv12_mux2to152_xor0;
  assign arrdiv12_fs69_and0 = arrdiv12_fs69_not0 & b[9];
  assign arrdiv12_fs69_xor1 = arrdiv12_fs68_or0 ^ arrdiv12_fs69_xor0;
  assign arrdiv12_fs69_not1 = ~arrdiv12_fs69_xor0;
  assign arrdiv12_fs69_and1 = arrdiv12_fs69_not1 & arrdiv12_fs68_or0;
  assign arrdiv12_fs69_or0 = arrdiv12_fs69_and1 | arrdiv12_fs69_and0;
  assign arrdiv12_fs70_xor0 = arrdiv12_mux2to153_xor0 ^ b[10];
  assign arrdiv12_fs70_not0 = ~arrdiv12_mux2to153_xor0;
  assign arrdiv12_fs70_and0 = arrdiv12_fs70_not0 & b[10];
  assign arrdiv12_fs70_xor1 = arrdiv12_fs69_or0 ^ arrdiv12_fs70_xor0;
  assign arrdiv12_fs70_not1 = ~arrdiv12_fs70_xor0;
  assign arrdiv12_fs70_and1 = arrdiv12_fs70_not1 & arrdiv12_fs69_or0;
  assign arrdiv12_fs70_or0 = arrdiv12_fs70_and1 | arrdiv12_fs70_and0;
  assign arrdiv12_fs71_xor0 = arrdiv12_mux2to154_xor0 ^ b[11];
  assign arrdiv12_fs71_not0 = ~arrdiv12_mux2to154_xor0;
  assign arrdiv12_fs71_and0 = arrdiv12_fs71_not0 & b[11];
  assign arrdiv12_fs71_xor1 = arrdiv12_fs70_or0 ^ arrdiv12_fs71_xor0;
  assign arrdiv12_fs71_not1 = ~arrdiv12_fs71_xor0;
  assign arrdiv12_fs71_and1 = arrdiv12_fs71_not1 & arrdiv12_fs70_or0;
  assign arrdiv12_fs71_or0 = arrdiv12_fs71_and1 | arrdiv12_fs71_and0;
  assign arrdiv12_mux2to155_and0 = a[6] & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to155_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to155_and1 = arrdiv12_fs60_xor0 & arrdiv12_mux2to155_not0;
  assign arrdiv12_mux2to155_xor0 = arrdiv12_mux2to155_and0 ^ arrdiv12_mux2to155_and1;
  assign arrdiv12_mux2to156_and0 = arrdiv12_mux2to144_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to156_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to156_and1 = arrdiv12_fs61_xor1 & arrdiv12_mux2to156_not0;
  assign arrdiv12_mux2to156_xor0 = arrdiv12_mux2to156_and0 ^ arrdiv12_mux2to156_and1;
  assign arrdiv12_mux2to157_and0 = arrdiv12_mux2to145_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to157_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to157_and1 = arrdiv12_fs62_xor1 & arrdiv12_mux2to157_not0;
  assign arrdiv12_mux2to157_xor0 = arrdiv12_mux2to157_and0 ^ arrdiv12_mux2to157_and1;
  assign arrdiv12_mux2to158_and0 = arrdiv12_mux2to146_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to158_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to158_and1 = arrdiv12_fs63_xor1 & arrdiv12_mux2to158_not0;
  assign arrdiv12_mux2to158_xor0 = arrdiv12_mux2to158_and0 ^ arrdiv12_mux2to158_and1;
  assign arrdiv12_mux2to159_and0 = arrdiv12_mux2to147_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to159_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to159_and1 = arrdiv12_fs64_xor1 & arrdiv12_mux2to159_not0;
  assign arrdiv12_mux2to159_xor0 = arrdiv12_mux2to159_and0 ^ arrdiv12_mux2to159_and1;
  assign arrdiv12_mux2to160_and0 = arrdiv12_mux2to148_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to160_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to160_and1 = arrdiv12_fs65_xor1 & arrdiv12_mux2to160_not0;
  assign arrdiv12_mux2to160_xor0 = arrdiv12_mux2to160_and0 ^ arrdiv12_mux2to160_and1;
  assign arrdiv12_mux2to161_and0 = arrdiv12_mux2to149_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to161_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to161_and1 = arrdiv12_fs66_xor1 & arrdiv12_mux2to161_not0;
  assign arrdiv12_mux2to161_xor0 = arrdiv12_mux2to161_and0 ^ arrdiv12_mux2to161_and1;
  assign arrdiv12_mux2to162_and0 = arrdiv12_mux2to150_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to162_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to162_and1 = arrdiv12_fs67_xor1 & arrdiv12_mux2to162_not0;
  assign arrdiv12_mux2to162_xor0 = arrdiv12_mux2to162_and0 ^ arrdiv12_mux2to162_and1;
  assign arrdiv12_mux2to163_and0 = arrdiv12_mux2to151_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to163_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to163_and1 = arrdiv12_fs68_xor1 & arrdiv12_mux2to163_not0;
  assign arrdiv12_mux2to163_xor0 = arrdiv12_mux2to163_and0 ^ arrdiv12_mux2to163_and1;
  assign arrdiv12_mux2to164_and0 = arrdiv12_mux2to152_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to164_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to164_and1 = arrdiv12_fs69_xor1 & arrdiv12_mux2to164_not0;
  assign arrdiv12_mux2to164_xor0 = arrdiv12_mux2to164_and0 ^ arrdiv12_mux2to164_and1;
  assign arrdiv12_mux2to165_and0 = arrdiv12_mux2to153_xor0 & arrdiv12_fs71_or0;
  assign arrdiv12_mux2to165_not0 = ~arrdiv12_fs71_or0;
  assign arrdiv12_mux2to165_and1 = arrdiv12_fs70_xor1 & arrdiv12_mux2to165_not0;
  assign arrdiv12_mux2to165_xor0 = arrdiv12_mux2to165_and0 ^ arrdiv12_mux2to165_and1;
  assign arrdiv12_not5 = ~arrdiv12_fs71_or0;
  assign arrdiv12_fs72_xor0 = a[5] ^ b[0];
  assign arrdiv12_fs72_not0 = ~a[5];
  assign arrdiv12_fs72_and0 = arrdiv12_fs72_not0 & b[0];
  assign arrdiv12_fs72_not1 = ~arrdiv12_fs72_xor0;
  assign arrdiv12_fs73_xor0 = arrdiv12_mux2to155_xor0 ^ b[1];
  assign arrdiv12_fs73_not0 = ~arrdiv12_mux2to155_xor0;
  assign arrdiv12_fs73_and0 = arrdiv12_fs73_not0 & b[1];
  assign arrdiv12_fs73_xor1 = arrdiv12_fs72_and0 ^ arrdiv12_fs73_xor0;
  assign arrdiv12_fs73_not1 = ~arrdiv12_fs73_xor0;
  assign arrdiv12_fs73_and1 = arrdiv12_fs73_not1 & arrdiv12_fs72_and0;
  assign arrdiv12_fs73_or0 = arrdiv12_fs73_and1 | arrdiv12_fs73_and0;
  assign arrdiv12_fs74_xor0 = arrdiv12_mux2to156_xor0 ^ b[2];
  assign arrdiv12_fs74_not0 = ~arrdiv12_mux2to156_xor0;
  assign arrdiv12_fs74_and0 = arrdiv12_fs74_not0 & b[2];
  assign arrdiv12_fs74_xor1 = arrdiv12_fs73_or0 ^ arrdiv12_fs74_xor0;
  assign arrdiv12_fs74_not1 = ~arrdiv12_fs74_xor0;
  assign arrdiv12_fs74_and1 = arrdiv12_fs74_not1 & arrdiv12_fs73_or0;
  assign arrdiv12_fs74_or0 = arrdiv12_fs74_and1 | arrdiv12_fs74_and0;
  assign arrdiv12_fs75_xor0 = arrdiv12_mux2to157_xor0 ^ b[3];
  assign arrdiv12_fs75_not0 = ~arrdiv12_mux2to157_xor0;
  assign arrdiv12_fs75_and0 = arrdiv12_fs75_not0 & b[3];
  assign arrdiv12_fs75_xor1 = arrdiv12_fs74_or0 ^ arrdiv12_fs75_xor0;
  assign arrdiv12_fs75_not1 = ~arrdiv12_fs75_xor0;
  assign arrdiv12_fs75_and1 = arrdiv12_fs75_not1 & arrdiv12_fs74_or0;
  assign arrdiv12_fs75_or0 = arrdiv12_fs75_and1 | arrdiv12_fs75_and0;
  assign arrdiv12_fs76_xor0 = arrdiv12_mux2to158_xor0 ^ b[4];
  assign arrdiv12_fs76_not0 = ~arrdiv12_mux2to158_xor0;
  assign arrdiv12_fs76_and0 = arrdiv12_fs76_not0 & b[4];
  assign arrdiv12_fs76_xor1 = arrdiv12_fs75_or0 ^ arrdiv12_fs76_xor0;
  assign arrdiv12_fs76_not1 = ~arrdiv12_fs76_xor0;
  assign arrdiv12_fs76_and1 = arrdiv12_fs76_not1 & arrdiv12_fs75_or0;
  assign arrdiv12_fs76_or0 = arrdiv12_fs76_and1 | arrdiv12_fs76_and0;
  assign arrdiv12_fs77_xor0 = arrdiv12_mux2to159_xor0 ^ b[5];
  assign arrdiv12_fs77_not0 = ~arrdiv12_mux2to159_xor0;
  assign arrdiv12_fs77_and0 = arrdiv12_fs77_not0 & b[5];
  assign arrdiv12_fs77_xor1 = arrdiv12_fs76_or0 ^ arrdiv12_fs77_xor0;
  assign arrdiv12_fs77_not1 = ~arrdiv12_fs77_xor0;
  assign arrdiv12_fs77_and1 = arrdiv12_fs77_not1 & arrdiv12_fs76_or0;
  assign arrdiv12_fs77_or0 = arrdiv12_fs77_and1 | arrdiv12_fs77_and0;
  assign arrdiv12_fs78_xor0 = arrdiv12_mux2to160_xor0 ^ b[6];
  assign arrdiv12_fs78_not0 = ~arrdiv12_mux2to160_xor0;
  assign arrdiv12_fs78_and0 = arrdiv12_fs78_not0 & b[6];
  assign arrdiv12_fs78_xor1 = arrdiv12_fs77_or0 ^ arrdiv12_fs78_xor0;
  assign arrdiv12_fs78_not1 = ~arrdiv12_fs78_xor0;
  assign arrdiv12_fs78_and1 = arrdiv12_fs78_not1 & arrdiv12_fs77_or0;
  assign arrdiv12_fs78_or0 = arrdiv12_fs78_and1 | arrdiv12_fs78_and0;
  assign arrdiv12_fs79_xor0 = arrdiv12_mux2to161_xor0 ^ b[7];
  assign arrdiv12_fs79_not0 = ~arrdiv12_mux2to161_xor0;
  assign arrdiv12_fs79_and0 = arrdiv12_fs79_not0 & b[7];
  assign arrdiv12_fs79_xor1 = arrdiv12_fs78_or0 ^ arrdiv12_fs79_xor0;
  assign arrdiv12_fs79_not1 = ~arrdiv12_fs79_xor0;
  assign arrdiv12_fs79_and1 = arrdiv12_fs79_not1 & arrdiv12_fs78_or0;
  assign arrdiv12_fs79_or0 = arrdiv12_fs79_and1 | arrdiv12_fs79_and0;
  assign arrdiv12_fs80_xor0 = arrdiv12_mux2to162_xor0 ^ b[8];
  assign arrdiv12_fs80_not0 = ~arrdiv12_mux2to162_xor0;
  assign arrdiv12_fs80_and0 = arrdiv12_fs80_not0 & b[8];
  assign arrdiv12_fs80_xor1 = arrdiv12_fs79_or0 ^ arrdiv12_fs80_xor0;
  assign arrdiv12_fs80_not1 = ~arrdiv12_fs80_xor0;
  assign arrdiv12_fs80_and1 = arrdiv12_fs80_not1 & arrdiv12_fs79_or0;
  assign arrdiv12_fs80_or0 = arrdiv12_fs80_and1 | arrdiv12_fs80_and0;
  assign arrdiv12_fs81_xor0 = arrdiv12_mux2to163_xor0 ^ b[9];
  assign arrdiv12_fs81_not0 = ~arrdiv12_mux2to163_xor0;
  assign arrdiv12_fs81_and0 = arrdiv12_fs81_not0 & b[9];
  assign arrdiv12_fs81_xor1 = arrdiv12_fs80_or0 ^ arrdiv12_fs81_xor0;
  assign arrdiv12_fs81_not1 = ~arrdiv12_fs81_xor0;
  assign arrdiv12_fs81_and1 = arrdiv12_fs81_not1 & arrdiv12_fs80_or0;
  assign arrdiv12_fs81_or0 = arrdiv12_fs81_and1 | arrdiv12_fs81_and0;
  assign arrdiv12_fs82_xor0 = arrdiv12_mux2to164_xor0 ^ b[10];
  assign arrdiv12_fs82_not0 = ~arrdiv12_mux2to164_xor0;
  assign arrdiv12_fs82_and0 = arrdiv12_fs82_not0 & b[10];
  assign arrdiv12_fs82_xor1 = arrdiv12_fs81_or0 ^ arrdiv12_fs82_xor0;
  assign arrdiv12_fs82_not1 = ~arrdiv12_fs82_xor0;
  assign arrdiv12_fs82_and1 = arrdiv12_fs82_not1 & arrdiv12_fs81_or0;
  assign arrdiv12_fs82_or0 = arrdiv12_fs82_and1 | arrdiv12_fs82_and0;
  assign arrdiv12_fs83_xor0 = arrdiv12_mux2to165_xor0 ^ b[11];
  assign arrdiv12_fs83_not0 = ~arrdiv12_mux2to165_xor0;
  assign arrdiv12_fs83_and0 = arrdiv12_fs83_not0 & b[11];
  assign arrdiv12_fs83_xor1 = arrdiv12_fs82_or0 ^ arrdiv12_fs83_xor0;
  assign arrdiv12_fs83_not1 = ~arrdiv12_fs83_xor0;
  assign arrdiv12_fs83_and1 = arrdiv12_fs83_not1 & arrdiv12_fs82_or0;
  assign arrdiv12_fs83_or0 = arrdiv12_fs83_and1 | arrdiv12_fs83_and0;
  assign arrdiv12_mux2to166_and0 = a[5] & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to166_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to166_and1 = arrdiv12_fs72_xor0 & arrdiv12_mux2to166_not0;
  assign arrdiv12_mux2to166_xor0 = arrdiv12_mux2to166_and0 ^ arrdiv12_mux2to166_and1;
  assign arrdiv12_mux2to167_and0 = arrdiv12_mux2to155_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to167_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to167_and1 = arrdiv12_fs73_xor1 & arrdiv12_mux2to167_not0;
  assign arrdiv12_mux2to167_xor0 = arrdiv12_mux2to167_and0 ^ arrdiv12_mux2to167_and1;
  assign arrdiv12_mux2to168_and0 = arrdiv12_mux2to156_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to168_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to168_and1 = arrdiv12_fs74_xor1 & arrdiv12_mux2to168_not0;
  assign arrdiv12_mux2to168_xor0 = arrdiv12_mux2to168_and0 ^ arrdiv12_mux2to168_and1;
  assign arrdiv12_mux2to169_and0 = arrdiv12_mux2to157_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to169_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to169_and1 = arrdiv12_fs75_xor1 & arrdiv12_mux2to169_not0;
  assign arrdiv12_mux2to169_xor0 = arrdiv12_mux2to169_and0 ^ arrdiv12_mux2to169_and1;
  assign arrdiv12_mux2to170_and0 = arrdiv12_mux2to158_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to170_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to170_and1 = arrdiv12_fs76_xor1 & arrdiv12_mux2to170_not0;
  assign arrdiv12_mux2to170_xor0 = arrdiv12_mux2to170_and0 ^ arrdiv12_mux2to170_and1;
  assign arrdiv12_mux2to171_and0 = arrdiv12_mux2to159_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to171_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to171_and1 = arrdiv12_fs77_xor1 & arrdiv12_mux2to171_not0;
  assign arrdiv12_mux2to171_xor0 = arrdiv12_mux2to171_and0 ^ arrdiv12_mux2to171_and1;
  assign arrdiv12_mux2to172_and0 = arrdiv12_mux2to160_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to172_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to172_and1 = arrdiv12_fs78_xor1 & arrdiv12_mux2to172_not0;
  assign arrdiv12_mux2to172_xor0 = arrdiv12_mux2to172_and0 ^ arrdiv12_mux2to172_and1;
  assign arrdiv12_mux2to173_and0 = arrdiv12_mux2to161_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to173_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to173_and1 = arrdiv12_fs79_xor1 & arrdiv12_mux2to173_not0;
  assign arrdiv12_mux2to173_xor0 = arrdiv12_mux2to173_and0 ^ arrdiv12_mux2to173_and1;
  assign arrdiv12_mux2to174_and0 = arrdiv12_mux2to162_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to174_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to174_and1 = arrdiv12_fs80_xor1 & arrdiv12_mux2to174_not0;
  assign arrdiv12_mux2to174_xor0 = arrdiv12_mux2to174_and0 ^ arrdiv12_mux2to174_and1;
  assign arrdiv12_mux2to175_and0 = arrdiv12_mux2to163_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to175_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to175_and1 = arrdiv12_fs81_xor1 & arrdiv12_mux2to175_not0;
  assign arrdiv12_mux2to175_xor0 = arrdiv12_mux2to175_and0 ^ arrdiv12_mux2to175_and1;
  assign arrdiv12_mux2to176_and0 = arrdiv12_mux2to164_xor0 & arrdiv12_fs83_or0;
  assign arrdiv12_mux2to176_not0 = ~arrdiv12_fs83_or0;
  assign arrdiv12_mux2to176_and1 = arrdiv12_fs82_xor1 & arrdiv12_mux2to176_not0;
  assign arrdiv12_mux2to176_xor0 = arrdiv12_mux2to176_and0 ^ arrdiv12_mux2to176_and1;
  assign arrdiv12_not6 = ~arrdiv12_fs83_or0;
  assign arrdiv12_fs84_xor0 = a[4] ^ b[0];
  assign arrdiv12_fs84_not0 = ~a[4];
  assign arrdiv12_fs84_and0 = arrdiv12_fs84_not0 & b[0];
  assign arrdiv12_fs84_not1 = ~arrdiv12_fs84_xor0;
  assign arrdiv12_fs85_xor0 = arrdiv12_mux2to166_xor0 ^ b[1];
  assign arrdiv12_fs85_not0 = ~arrdiv12_mux2to166_xor0;
  assign arrdiv12_fs85_and0 = arrdiv12_fs85_not0 & b[1];
  assign arrdiv12_fs85_xor1 = arrdiv12_fs84_and0 ^ arrdiv12_fs85_xor0;
  assign arrdiv12_fs85_not1 = ~arrdiv12_fs85_xor0;
  assign arrdiv12_fs85_and1 = arrdiv12_fs85_not1 & arrdiv12_fs84_and0;
  assign arrdiv12_fs85_or0 = arrdiv12_fs85_and1 | arrdiv12_fs85_and0;
  assign arrdiv12_fs86_xor0 = arrdiv12_mux2to167_xor0 ^ b[2];
  assign arrdiv12_fs86_not0 = ~arrdiv12_mux2to167_xor0;
  assign arrdiv12_fs86_and0 = arrdiv12_fs86_not0 & b[2];
  assign arrdiv12_fs86_xor1 = arrdiv12_fs85_or0 ^ arrdiv12_fs86_xor0;
  assign arrdiv12_fs86_not1 = ~arrdiv12_fs86_xor0;
  assign arrdiv12_fs86_and1 = arrdiv12_fs86_not1 & arrdiv12_fs85_or0;
  assign arrdiv12_fs86_or0 = arrdiv12_fs86_and1 | arrdiv12_fs86_and0;
  assign arrdiv12_fs87_xor0 = arrdiv12_mux2to168_xor0 ^ b[3];
  assign arrdiv12_fs87_not0 = ~arrdiv12_mux2to168_xor0;
  assign arrdiv12_fs87_and0 = arrdiv12_fs87_not0 & b[3];
  assign arrdiv12_fs87_xor1 = arrdiv12_fs86_or0 ^ arrdiv12_fs87_xor0;
  assign arrdiv12_fs87_not1 = ~arrdiv12_fs87_xor0;
  assign arrdiv12_fs87_and1 = arrdiv12_fs87_not1 & arrdiv12_fs86_or0;
  assign arrdiv12_fs87_or0 = arrdiv12_fs87_and1 | arrdiv12_fs87_and0;
  assign arrdiv12_fs88_xor0 = arrdiv12_mux2to169_xor0 ^ b[4];
  assign arrdiv12_fs88_not0 = ~arrdiv12_mux2to169_xor0;
  assign arrdiv12_fs88_and0 = arrdiv12_fs88_not0 & b[4];
  assign arrdiv12_fs88_xor1 = arrdiv12_fs87_or0 ^ arrdiv12_fs88_xor0;
  assign arrdiv12_fs88_not1 = ~arrdiv12_fs88_xor0;
  assign arrdiv12_fs88_and1 = arrdiv12_fs88_not1 & arrdiv12_fs87_or0;
  assign arrdiv12_fs88_or0 = arrdiv12_fs88_and1 | arrdiv12_fs88_and0;
  assign arrdiv12_fs89_xor0 = arrdiv12_mux2to170_xor0 ^ b[5];
  assign arrdiv12_fs89_not0 = ~arrdiv12_mux2to170_xor0;
  assign arrdiv12_fs89_and0 = arrdiv12_fs89_not0 & b[5];
  assign arrdiv12_fs89_xor1 = arrdiv12_fs88_or0 ^ arrdiv12_fs89_xor0;
  assign arrdiv12_fs89_not1 = ~arrdiv12_fs89_xor0;
  assign arrdiv12_fs89_and1 = arrdiv12_fs89_not1 & arrdiv12_fs88_or0;
  assign arrdiv12_fs89_or0 = arrdiv12_fs89_and1 | arrdiv12_fs89_and0;
  assign arrdiv12_fs90_xor0 = arrdiv12_mux2to171_xor0 ^ b[6];
  assign arrdiv12_fs90_not0 = ~arrdiv12_mux2to171_xor0;
  assign arrdiv12_fs90_and0 = arrdiv12_fs90_not0 & b[6];
  assign arrdiv12_fs90_xor1 = arrdiv12_fs89_or0 ^ arrdiv12_fs90_xor0;
  assign arrdiv12_fs90_not1 = ~arrdiv12_fs90_xor0;
  assign arrdiv12_fs90_and1 = arrdiv12_fs90_not1 & arrdiv12_fs89_or0;
  assign arrdiv12_fs90_or0 = arrdiv12_fs90_and1 | arrdiv12_fs90_and0;
  assign arrdiv12_fs91_xor0 = arrdiv12_mux2to172_xor0 ^ b[7];
  assign arrdiv12_fs91_not0 = ~arrdiv12_mux2to172_xor0;
  assign arrdiv12_fs91_and0 = arrdiv12_fs91_not0 & b[7];
  assign arrdiv12_fs91_xor1 = arrdiv12_fs90_or0 ^ arrdiv12_fs91_xor0;
  assign arrdiv12_fs91_not1 = ~arrdiv12_fs91_xor0;
  assign arrdiv12_fs91_and1 = arrdiv12_fs91_not1 & arrdiv12_fs90_or0;
  assign arrdiv12_fs91_or0 = arrdiv12_fs91_and1 | arrdiv12_fs91_and0;
  assign arrdiv12_fs92_xor0 = arrdiv12_mux2to173_xor0 ^ b[8];
  assign arrdiv12_fs92_not0 = ~arrdiv12_mux2to173_xor0;
  assign arrdiv12_fs92_and0 = arrdiv12_fs92_not0 & b[8];
  assign arrdiv12_fs92_xor1 = arrdiv12_fs91_or0 ^ arrdiv12_fs92_xor0;
  assign arrdiv12_fs92_not1 = ~arrdiv12_fs92_xor0;
  assign arrdiv12_fs92_and1 = arrdiv12_fs92_not1 & arrdiv12_fs91_or0;
  assign arrdiv12_fs92_or0 = arrdiv12_fs92_and1 | arrdiv12_fs92_and0;
  assign arrdiv12_fs93_xor0 = arrdiv12_mux2to174_xor0 ^ b[9];
  assign arrdiv12_fs93_not0 = ~arrdiv12_mux2to174_xor0;
  assign arrdiv12_fs93_and0 = arrdiv12_fs93_not0 & b[9];
  assign arrdiv12_fs93_xor1 = arrdiv12_fs92_or0 ^ arrdiv12_fs93_xor0;
  assign arrdiv12_fs93_not1 = ~arrdiv12_fs93_xor0;
  assign arrdiv12_fs93_and1 = arrdiv12_fs93_not1 & arrdiv12_fs92_or0;
  assign arrdiv12_fs93_or0 = arrdiv12_fs93_and1 | arrdiv12_fs93_and0;
  assign arrdiv12_fs94_xor0 = arrdiv12_mux2to175_xor0 ^ b[10];
  assign arrdiv12_fs94_not0 = ~arrdiv12_mux2to175_xor0;
  assign arrdiv12_fs94_and0 = arrdiv12_fs94_not0 & b[10];
  assign arrdiv12_fs94_xor1 = arrdiv12_fs93_or0 ^ arrdiv12_fs94_xor0;
  assign arrdiv12_fs94_not1 = ~arrdiv12_fs94_xor0;
  assign arrdiv12_fs94_and1 = arrdiv12_fs94_not1 & arrdiv12_fs93_or0;
  assign arrdiv12_fs94_or0 = arrdiv12_fs94_and1 | arrdiv12_fs94_and0;
  assign arrdiv12_fs95_xor0 = arrdiv12_mux2to176_xor0 ^ b[11];
  assign arrdiv12_fs95_not0 = ~arrdiv12_mux2to176_xor0;
  assign arrdiv12_fs95_and0 = arrdiv12_fs95_not0 & b[11];
  assign arrdiv12_fs95_xor1 = arrdiv12_fs94_or0 ^ arrdiv12_fs95_xor0;
  assign arrdiv12_fs95_not1 = ~arrdiv12_fs95_xor0;
  assign arrdiv12_fs95_and1 = arrdiv12_fs95_not1 & arrdiv12_fs94_or0;
  assign arrdiv12_fs95_or0 = arrdiv12_fs95_and1 | arrdiv12_fs95_and0;
  assign arrdiv12_mux2to177_and0 = a[4] & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to177_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to177_and1 = arrdiv12_fs84_xor0 & arrdiv12_mux2to177_not0;
  assign arrdiv12_mux2to177_xor0 = arrdiv12_mux2to177_and0 ^ arrdiv12_mux2to177_and1;
  assign arrdiv12_mux2to178_and0 = arrdiv12_mux2to166_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to178_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to178_and1 = arrdiv12_fs85_xor1 & arrdiv12_mux2to178_not0;
  assign arrdiv12_mux2to178_xor0 = arrdiv12_mux2to178_and0 ^ arrdiv12_mux2to178_and1;
  assign arrdiv12_mux2to179_and0 = arrdiv12_mux2to167_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to179_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to179_and1 = arrdiv12_fs86_xor1 & arrdiv12_mux2to179_not0;
  assign arrdiv12_mux2to179_xor0 = arrdiv12_mux2to179_and0 ^ arrdiv12_mux2to179_and1;
  assign arrdiv12_mux2to180_and0 = arrdiv12_mux2to168_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to180_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to180_and1 = arrdiv12_fs87_xor1 & arrdiv12_mux2to180_not0;
  assign arrdiv12_mux2to180_xor0 = arrdiv12_mux2to180_and0 ^ arrdiv12_mux2to180_and1;
  assign arrdiv12_mux2to181_and0 = arrdiv12_mux2to169_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to181_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to181_and1 = arrdiv12_fs88_xor1 & arrdiv12_mux2to181_not0;
  assign arrdiv12_mux2to181_xor0 = arrdiv12_mux2to181_and0 ^ arrdiv12_mux2to181_and1;
  assign arrdiv12_mux2to182_and0 = arrdiv12_mux2to170_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to182_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to182_and1 = arrdiv12_fs89_xor1 & arrdiv12_mux2to182_not0;
  assign arrdiv12_mux2to182_xor0 = arrdiv12_mux2to182_and0 ^ arrdiv12_mux2to182_and1;
  assign arrdiv12_mux2to183_and0 = arrdiv12_mux2to171_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to183_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to183_and1 = arrdiv12_fs90_xor1 & arrdiv12_mux2to183_not0;
  assign arrdiv12_mux2to183_xor0 = arrdiv12_mux2to183_and0 ^ arrdiv12_mux2to183_and1;
  assign arrdiv12_mux2to184_and0 = arrdiv12_mux2to172_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to184_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to184_and1 = arrdiv12_fs91_xor1 & arrdiv12_mux2to184_not0;
  assign arrdiv12_mux2to184_xor0 = arrdiv12_mux2to184_and0 ^ arrdiv12_mux2to184_and1;
  assign arrdiv12_mux2to185_and0 = arrdiv12_mux2to173_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to185_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to185_and1 = arrdiv12_fs92_xor1 & arrdiv12_mux2to185_not0;
  assign arrdiv12_mux2to185_xor0 = arrdiv12_mux2to185_and0 ^ arrdiv12_mux2to185_and1;
  assign arrdiv12_mux2to186_and0 = arrdiv12_mux2to174_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to186_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to186_and1 = arrdiv12_fs93_xor1 & arrdiv12_mux2to186_not0;
  assign arrdiv12_mux2to186_xor0 = arrdiv12_mux2to186_and0 ^ arrdiv12_mux2to186_and1;
  assign arrdiv12_mux2to187_and0 = arrdiv12_mux2to175_xor0 & arrdiv12_fs95_or0;
  assign arrdiv12_mux2to187_not0 = ~arrdiv12_fs95_or0;
  assign arrdiv12_mux2to187_and1 = arrdiv12_fs94_xor1 & arrdiv12_mux2to187_not0;
  assign arrdiv12_mux2to187_xor0 = arrdiv12_mux2to187_and0 ^ arrdiv12_mux2to187_and1;
  assign arrdiv12_not7 = ~arrdiv12_fs95_or0;
  assign arrdiv12_fs96_xor0 = a[3] ^ b[0];
  assign arrdiv12_fs96_not0 = ~a[3];
  assign arrdiv12_fs96_and0 = arrdiv12_fs96_not0 & b[0];
  assign arrdiv12_fs96_not1 = ~arrdiv12_fs96_xor0;
  assign arrdiv12_fs97_xor0 = arrdiv12_mux2to177_xor0 ^ b[1];
  assign arrdiv12_fs97_not0 = ~arrdiv12_mux2to177_xor0;
  assign arrdiv12_fs97_and0 = arrdiv12_fs97_not0 & b[1];
  assign arrdiv12_fs97_xor1 = arrdiv12_fs96_and0 ^ arrdiv12_fs97_xor0;
  assign arrdiv12_fs97_not1 = ~arrdiv12_fs97_xor0;
  assign arrdiv12_fs97_and1 = arrdiv12_fs97_not1 & arrdiv12_fs96_and0;
  assign arrdiv12_fs97_or0 = arrdiv12_fs97_and1 | arrdiv12_fs97_and0;
  assign arrdiv12_fs98_xor0 = arrdiv12_mux2to178_xor0 ^ b[2];
  assign arrdiv12_fs98_not0 = ~arrdiv12_mux2to178_xor0;
  assign arrdiv12_fs98_and0 = arrdiv12_fs98_not0 & b[2];
  assign arrdiv12_fs98_xor1 = arrdiv12_fs97_or0 ^ arrdiv12_fs98_xor0;
  assign arrdiv12_fs98_not1 = ~arrdiv12_fs98_xor0;
  assign arrdiv12_fs98_and1 = arrdiv12_fs98_not1 & arrdiv12_fs97_or0;
  assign arrdiv12_fs98_or0 = arrdiv12_fs98_and1 | arrdiv12_fs98_and0;
  assign arrdiv12_fs99_xor0 = arrdiv12_mux2to179_xor0 ^ b[3];
  assign arrdiv12_fs99_not0 = ~arrdiv12_mux2to179_xor0;
  assign arrdiv12_fs99_and0 = arrdiv12_fs99_not0 & b[3];
  assign arrdiv12_fs99_xor1 = arrdiv12_fs98_or0 ^ arrdiv12_fs99_xor0;
  assign arrdiv12_fs99_not1 = ~arrdiv12_fs99_xor0;
  assign arrdiv12_fs99_and1 = arrdiv12_fs99_not1 & arrdiv12_fs98_or0;
  assign arrdiv12_fs99_or0 = arrdiv12_fs99_and1 | arrdiv12_fs99_and0;
  assign arrdiv12_fs100_xor0 = arrdiv12_mux2to180_xor0 ^ b[4];
  assign arrdiv12_fs100_not0 = ~arrdiv12_mux2to180_xor0;
  assign arrdiv12_fs100_and0 = arrdiv12_fs100_not0 & b[4];
  assign arrdiv12_fs100_xor1 = arrdiv12_fs99_or0 ^ arrdiv12_fs100_xor0;
  assign arrdiv12_fs100_not1 = ~arrdiv12_fs100_xor0;
  assign arrdiv12_fs100_and1 = arrdiv12_fs100_not1 & arrdiv12_fs99_or0;
  assign arrdiv12_fs100_or0 = arrdiv12_fs100_and1 | arrdiv12_fs100_and0;
  assign arrdiv12_fs101_xor0 = arrdiv12_mux2to181_xor0 ^ b[5];
  assign arrdiv12_fs101_not0 = ~arrdiv12_mux2to181_xor0;
  assign arrdiv12_fs101_and0 = arrdiv12_fs101_not0 & b[5];
  assign arrdiv12_fs101_xor1 = arrdiv12_fs100_or0 ^ arrdiv12_fs101_xor0;
  assign arrdiv12_fs101_not1 = ~arrdiv12_fs101_xor0;
  assign arrdiv12_fs101_and1 = arrdiv12_fs101_not1 & arrdiv12_fs100_or0;
  assign arrdiv12_fs101_or0 = arrdiv12_fs101_and1 | arrdiv12_fs101_and0;
  assign arrdiv12_fs102_xor0 = arrdiv12_mux2to182_xor0 ^ b[6];
  assign arrdiv12_fs102_not0 = ~arrdiv12_mux2to182_xor0;
  assign arrdiv12_fs102_and0 = arrdiv12_fs102_not0 & b[6];
  assign arrdiv12_fs102_xor1 = arrdiv12_fs101_or0 ^ arrdiv12_fs102_xor0;
  assign arrdiv12_fs102_not1 = ~arrdiv12_fs102_xor0;
  assign arrdiv12_fs102_and1 = arrdiv12_fs102_not1 & arrdiv12_fs101_or0;
  assign arrdiv12_fs102_or0 = arrdiv12_fs102_and1 | arrdiv12_fs102_and0;
  assign arrdiv12_fs103_xor0 = arrdiv12_mux2to183_xor0 ^ b[7];
  assign arrdiv12_fs103_not0 = ~arrdiv12_mux2to183_xor0;
  assign arrdiv12_fs103_and0 = arrdiv12_fs103_not0 & b[7];
  assign arrdiv12_fs103_xor1 = arrdiv12_fs102_or0 ^ arrdiv12_fs103_xor0;
  assign arrdiv12_fs103_not1 = ~arrdiv12_fs103_xor0;
  assign arrdiv12_fs103_and1 = arrdiv12_fs103_not1 & arrdiv12_fs102_or0;
  assign arrdiv12_fs103_or0 = arrdiv12_fs103_and1 | arrdiv12_fs103_and0;
  assign arrdiv12_fs104_xor0 = arrdiv12_mux2to184_xor0 ^ b[8];
  assign arrdiv12_fs104_not0 = ~arrdiv12_mux2to184_xor0;
  assign arrdiv12_fs104_and0 = arrdiv12_fs104_not0 & b[8];
  assign arrdiv12_fs104_xor1 = arrdiv12_fs103_or0 ^ arrdiv12_fs104_xor0;
  assign arrdiv12_fs104_not1 = ~arrdiv12_fs104_xor0;
  assign arrdiv12_fs104_and1 = arrdiv12_fs104_not1 & arrdiv12_fs103_or0;
  assign arrdiv12_fs104_or0 = arrdiv12_fs104_and1 | arrdiv12_fs104_and0;
  assign arrdiv12_fs105_xor0 = arrdiv12_mux2to185_xor0 ^ b[9];
  assign arrdiv12_fs105_not0 = ~arrdiv12_mux2to185_xor0;
  assign arrdiv12_fs105_and0 = arrdiv12_fs105_not0 & b[9];
  assign arrdiv12_fs105_xor1 = arrdiv12_fs104_or0 ^ arrdiv12_fs105_xor0;
  assign arrdiv12_fs105_not1 = ~arrdiv12_fs105_xor0;
  assign arrdiv12_fs105_and1 = arrdiv12_fs105_not1 & arrdiv12_fs104_or0;
  assign arrdiv12_fs105_or0 = arrdiv12_fs105_and1 | arrdiv12_fs105_and0;
  assign arrdiv12_fs106_xor0 = arrdiv12_mux2to186_xor0 ^ b[10];
  assign arrdiv12_fs106_not0 = ~arrdiv12_mux2to186_xor0;
  assign arrdiv12_fs106_and0 = arrdiv12_fs106_not0 & b[10];
  assign arrdiv12_fs106_xor1 = arrdiv12_fs105_or0 ^ arrdiv12_fs106_xor0;
  assign arrdiv12_fs106_not1 = ~arrdiv12_fs106_xor0;
  assign arrdiv12_fs106_and1 = arrdiv12_fs106_not1 & arrdiv12_fs105_or0;
  assign arrdiv12_fs106_or0 = arrdiv12_fs106_and1 | arrdiv12_fs106_and0;
  assign arrdiv12_fs107_xor0 = arrdiv12_mux2to187_xor0 ^ b[11];
  assign arrdiv12_fs107_not0 = ~arrdiv12_mux2to187_xor0;
  assign arrdiv12_fs107_and0 = arrdiv12_fs107_not0 & b[11];
  assign arrdiv12_fs107_xor1 = arrdiv12_fs106_or0 ^ arrdiv12_fs107_xor0;
  assign arrdiv12_fs107_not1 = ~arrdiv12_fs107_xor0;
  assign arrdiv12_fs107_and1 = arrdiv12_fs107_not1 & arrdiv12_fs106_or0;
  assign arrdiv12_fs107_or0 = arrdiv12_fs107_and1 | arrdiv12_fs107_and0;
  assign arrdiv12_mux2to188_and0 = a[3] & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to188_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to188_and1 = arrdiv12_fs96_xor0 & arrdiv12_mux2to188_not0;
  assign arrdiv12_mux2to188_xor0 = arrdiv12_mux2to188_and0 ^ arrdiv12_mux2to188_and1;
  assign arrdiv12_mux2to189_and0 = arrdiv12_mux2to177_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to189_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to189_and1 = arrdiv12_fs97_xor1 & arrdiv12_mux2to189_not0;
  assign arrdiv12_mux2to189_xor0 = arrdiv12_mux2to189_and0 ^ arrdiv12_mux2to189_and1;
  assign arrdiv12_mux2to190_and0 = arrdiv12_mux2to178_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to190_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to190_and1 = arrdiv12_fs98_xor1 & arrdiv12_mux2to190_not0;
  assign arrdiv12_mux2to190_xor0 = arrdiv12_mux2to190_and0 ^ arrdiv12_mux2to190_and1;
  assign arrdiv12_mux2to191_and0 = arrdiv12_mux2to179_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to191_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to191_and1 = arrdiv12_fs99_xor1 & arrdiv12_mux2to191_not0;
  assign arrdiv12_mux2to191_xor0 = arrdiv12_mux2to191_and0 ^ arrdiv12_mux2to191_and1;
  assign arrdiv12_mux2to192_and0 = arrdiv12_mux2to180_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to192_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to192_and1 = arrdiv12_fs100_xor1 & arrdiv12_mux2to192_not0;
  assign arrdiv12_mux2to192_xor0 = arrdiv12_mux2to192_and0 ^ arrdiv12_mux2to192_and1;
  assign arrdiv12_mux2to193_and0 = arrdiv12_mux2to181_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to193_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to193_and1 = arrdiv12_fs101_xor1 & arrdiv12_mux2to193_not0;
  assign arrdiv12_mux2to193_xor0 = arrdiv12_mux2to193_and0 ^ arrdiv12_mux2to193_and1;
  assign arrdiv12_mux2to194_and0 = arrdiv12_mux2to182_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to194_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to194_and1 = arrdiv12_fs102_xor1 & arrdiv12_mux2to194_not0;
  assign arrdiv12_mux2to194_xor0 = arrdiv12_mux2to194_and0 ^ arrdiv12_mux2to194_and1;
  assign arrdiv12_mux2to195_and0 = arrdiv12_mux2to183_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to195_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to195_and1 = arrdiv12_fs103_xor1 & arrdiv12_mux2to195_not0;
  assign arrdiv12_mux2to195_xor0 = arrdiv12_mux2to195_and0 ^ arrdiv12_mux2to195_and1;
  assign arrdiv12_mux2to196_and0 = arrdiv12_mux2to184_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to196_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to196_and1 = arrdiv12_fs104_xor1 & arrdiv12_mux2to196_not0;
  assign arrdiv12_mux2to196_xor0 = arrdiv12_mux2to196_and0 ^ arrdiv12_mux2to196_and1;
  assign arrdiv12_mux2to197_and0 = arrdiv12_mux2to185_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to197_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to197_and1 = arrdiv12_fs105_xor1 & arrdiv12_mux2to197_not0;
  assign arrdiv12_mux2to197_xor0 = arrdiv12_mux2to197_and0 ^ arrdiv12_mux2to197_and1;
  assign arrdiv12_mux2to198_and0 = arrdiv12_mux2to186_xor0 & arrdiv12_fs107_or0;
  assign arrdiv12_mux2to198_not0 = ~arrdiv12_fs107_or0;
  assign arrdiv12_mux2to198_and1 = arrdiv12_fs106_xor1 & arrdiv12_mux2to198_not0;
  assign arrdiv12_mux2to198_xor0 = arrdiv12_mux2to198_and0 ^ arrdiv12_mux2to198_and1;
  assign arrdiv12_not8 = ~arrdiv12_fs107_or0;
  assign arrdiv12_fs108_xor0 = a[2] ^ b[0];
  assign arrdiv12_fs108_not0 = ~a[2];
  assign arrdiv12_fs108_and0 = arrdiv12_fs108_not0 & b[0];
  assign arrdiv12_fs108_not1 = ~arrdiv12_fs108_xor0;
  assign arrdiv12_fs109_xor0 = arrdiv12_mux2to188_xor0 ^ b[1];
  assign arrdiv12_fs109_not0 = ~arrdiv12_mux2to188_xor0;
  assign arrdiv12_fs109_and0 = arrdiv12_fs109_not0 & b[1];
  assign arrdiv12_fs109_xor1 = arrdiv12_fs108_and0 ^ arrdiv12_fs109_xor0;
  assign arrdiv12_fs109_not1 = ~arrdiv12_fs109_xor0;
  assign arrdiv12_fs109_and1 = arrdiv12_fs109_not1 & arrdiv12_fs108_and0;
  assign arrdiv12_fs109_or0 = arrdiv12_fs109_and1 | arrdiv12_fs109_and0;
  assign arrdiv12_fs110_xor0 = arrdiv12_mux2to189_xor0 ^ b[2];
  assign arrdiv12_fs110_not0 = ~arrdiv12_mux2to189_xor0;
  assign arrdiv12_fs110_and0 = arrdiv12_fs110_not0 & b[2];
  assign arrdiv12_fs110_xor1 = arrdiv12_fs109_or0 ^ arrdiv12_fs110_xor0;
  assign arrdiv12_fs110_not1 = ~arrdiv12_fs110_xor0;
  assign arrdiv12_fs110_and1 = arrdiv12_fs110_not1 & arrdiv12_fs109_or0;
  assign arrdiv12_fs110_or0 = arrdiv12_fs110_and1 | arrdiv12_fs110_and0;
  assign arrdiv12_fs111_xor0 = arrdiv12_mux2to190_xor0 ^ b[3];
  assign arrdiv12_fs111_not0 = ~arrdiv12_mux2to190_xor0;
  assign arrdiv12_fs111_and0 = arrdiv12_fs111_not0 & b[3];
  assign arrdiv12_fs111_xor1 = arrdiv12_fs110_or0 ^ arrdiv12_fs111_xor0;
  assign arrdiv12_fs111_not1 = ~arrdiv12_fs111_xor0;
  assign arrdiv12_fs111_and1 = arrdiv12_fs111_not1 & arrdiv12_fs110_or0;
  assign arrdiv12_fs111_or0 = arrdiv12_fs111_and1 | arrdiv12_fs111_and0;
  assign arrdiv12_fs112_xor0 = arrdiv12_mux2to191_xor0 ^ b[4];
  assign arrdiv12_fs112_not0 = ~arrdiv12_mux2to191_xor0;
  assign arrdiv12_fs112_and0 = arrdiv12_fs112_not0 & b[4];
  assign arrdiv12_fs112_xor1 = arrdiv12_fs111_or0 ^ arrdiv12_fs112_xor0;
  assign arrdiv12_fs112_not1 = ~arrdiv12_fs112_xor0;
  assign arrdiv12_fs112_and1 = arrdiv12_fs112_not1 & arrdiv12_fs111_or0;
  assign arrdiv12_fs112_or0 = arrdiv12_fs112_and1 | arrdiv12_fs112_and0;
  assign arrdiv12_fs113_xor0 = arrdiv12_mux2to192_xor0 ^ b[5];
  assign arrdiv12_fs113_not0 = ~arrdiv12_mux2to192_xor0;
  assign arrdiv12_fs113_and0 = arrdiv12_fs113_not0 & b[5];
  assign arrdiv12_fs113_xor1 = arrdiv12_fs112_or0 ^ arrdiv12_fs113_xor0;
  assign arrdiv12_fs113_not1 = ~arrdiv12_fs113_xor0;
  assign arrdiv12_fs113_and1 = arrdiv12_fs113_not1 & arrdiv12_fs112_or0;
  assign arrdiv12_fs113_or0 = arrdiv12_fs113_and1 | arrdiv12_fs113_and0;
  assign arrdiv12_fs114_xor0 = arrdiv12_mux2to193_xor0 ^ b[6];
  assign arrdiv12_fs114_not0 = ~arrdiv12_mux2to193_xor0;
  assign arrdiv12_fs114_and0 = arrdiv12_fs114_not0 & b[6];
  assign arrdiv12_fs114_xor1 = arrdiv12_fs113_or0 ^ arrdiv12_fs114_xor0;
  assign arrdiv12_fs114_not1 = ~arrdiv12_fs114_xor0;
  assign arrdiv12_fs114_and1 = arrdiv12_fs114_not1 & arrdiv12_fs113_or0;
  assign arrdiv12_fs114_or0 = arrdiv12_fs114_and1 | arrdiv12_fs114_and0;
  assign arrdiv12_fs115_xor0 = arrdiv12_mux2to194_xor0 ^ b[7];
  assign arrdiv12_fs115_not0 = ~arrdiv12_mux2to194_xor0;
  assign arrdiv12_fs115_and0 = arrdiv12_fs115_not0 & b[7];
  assign arrdiv12_fs115_xor1 = arrdiv12_fs114_or0 ^ arrdiv12_fs115_xor0;
  assign arrdiv12_fs115_not1 = ~arrdiv12_fs115_xor0;
  assign arrdiv12_fs115_and1 = arrdiv12_fs115_not1 & arrdiv12_fs114_or0;
  assign arrdiv12_fs115_or0 = arrdiv12_fs115_and1 | arrdiv12_fs115_and0;
  assign arrdiv12_fs116_xor0 = arrdiv12_mux2to195_xor0 ^ b[8];
  assign arrdiv12_fs116_not0 = ~arrdiv12_mux2to195_xor0;
  assign arrdiv12_fs116_and0 = arrdiv12_fs116_not0 & b[8];
  assign arrdiv12_fs116_xor1 = arrdiv12_fs115_or0 ^ arrdiv12_fs116_xor0;
  assign arrdiv12_fs116_not1 = ~arrdiv12_fs116_xor0;
  assign arrdiv12_fs116_and1 = arrdiv12_fs116_not1 & arrdiv12_fs115_or0;
  assign arrdiv12_fs116_or0 = arrdiv12_fs116_and1 | arrdiv12_fs116_and0;
  assign arrdiv12_fs117_xor0 = arrdiv12_mux2to196_xor0 ^ b[9];
  assign arrdiv12_fs117_not0 = ~arrdiv12_mux2to196_xor0;
  assign arrdiv12_fs117_and0 = arrdiv12_fs117_not0 & b[9];
  assign arrdiv12_fs117_xor1 = arrdiv12_fs116_or0 ^ arrdiv12_fs117_xor0;
  assign arrdiv12_fs117_not1 = ~arrdiv12_fs117_xor0;
  assign arrdiv12_fs117_and1 = arrdiv12_fs117_not1 & arrdiv12_fs116_or0;
  assign arrdiv12_fs117_or0 = arrdiv12_fs117_and1 | arrdiv12_fs117_and0;
  assign arrdiv12_fs118_xor0 = arrdiv12_mux2to197_xor0 ^ b[10];
  assign arrdiv12_fs118_not0 = ~arrdiv12_mux2to197_xor0;
  assign arrdiv12_fs118_and0 = arrdiv12_fs118_not0 & b[10];
  assign arrdiv12_fs118_xor1 = arrdiv12_fs117_or0 ^ arrdiv12_fs118_xor0;
  assign arrdiv12_fs118_not1 = ~arrdiv12_fs118_xor0;
  assign arrdiv12_fs118_and1 = arrdiv12_fs118_not1 & arrdiv12_fs117_or0;
  assign arrdiv12_fs118_or0 = arrdiv12_fs118_and1 | arrdiv12_fs118_and0;
  assign arrdiv12_fs119_xor0 = arrdiv12_mux2to198_xor0 ^ b[11];
  assign arrdiv12_fs119_not0 = ~arrdiv12_mux2to198_xor0;
  assign arrdiv12_fs119_and0 = arrdiv12_fs119_not0 & b[11];
  assign arrdiv12_fs119_xor1 = arrdiv12_fs118_or0 ^ arrdiv12_fs119_xor0;
  assign arrdiv12_fs119_not1 = ~arrdiv12_fs119_xor0;
  assign arrdiv12_fs119_and1 = arrdiv12_fs119_not1 & arrdiv12_fs118_or0;
  assign arrdiv12_fs119_or0 = arrdiv12_fs119_and1 | arrdiv12_fs119_and0;
  assign arrdiv12_mux2to199_and0 = a[2] & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to199_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to199_and1 = arrdiv12_fs108_xor0 & arrdiv12_mux2to199_not0;
  assign arrdiv12_mux2to199_xor0 = arrdiv12_mux2to199_and0 ^ arrdiv12_mux2to199_and1;
  assign arrdiv12_mux2to1100_and0 = arrdiv12_mux2to188_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1100_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1100_and1 = arrdiv12_fs109_xor1 & arrdiv12_mux2to1100_not0;
  assign arrdiv12_mux2to1100_xor0 = arrdiv12_mux2to1100_and0 ^ arrdiv12_mux2to1100_and1;
  assign arrdiv12_mux2to1101_and0 = arrdiv12_mux2to189_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1101_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1101_and1 = arrdiv12_fs110_xor1 & arrdiv12_mux2to1101_not0;
  assign arrdiv12_mux2to1101_xor0 = arrdiv12_mux2to1101_and0 ^ arrdiv12_mux2to1101_and1;
  assign arrdiv12_mux2to1102_and0 = arrdiv12_mux2to190_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1102_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1102_and1 = arrdiv12_fs111_xor1 & arrdiv12_mux2to1102_not0;
  assign arrdiv12_mux2to1102_xor0 = arrdiv12_mux2to1102_and0 ^ arrdiv12_mux2to1102_and1;
  assign arrdiv12_mux2to1103_and0 = arrdiv12_mux2to191_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1103_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1103_and1 = arrdiv12_fs112_xor1 & arrdiv12_mux2to1103_not0;
  assign arrdiv12_mux2to1103_xor0 = arrdiv12_mux2to1103_and0 ^ arrdiv12_mux2to1103_and1;
  assign arrdiv12_mux2to1104_and0 = arrdiv12_mux2to192_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1104_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1104_and1 = arrdiv12_fs113_xor1 & arrdiv12_mux2to1104_not0;
  assign arrdiv12_mux2to1104_xor0 = arrdiv12_mux2to1104_and0 ^ arrdiv12_mux2to1104_and1;
  assign arrdiv12_mux2to1105_and0 = arrdiv12_mux2to193_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1105_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1105_and1 = arrdiv12_fs114_xor1 & arrdiv12_mux2to1105_not0;
  assign arrdiv12_mux2to1105_xor0 = arrdiv12_mux2to1105_and0 ^ arrdiv12_mux2to1105_and1;
  assign arrdiv12_mux2to1106_and0 = arrdiv12_mux2to194_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1106_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1106_and1 = arrdiv12_fs115_xor1 & arrdiv12_mux2to1106_not0;
  assign arrdiv12_mux2to1106_xor0 = arrdiv12_mux2to1106_and0 ^ arrdiv12_mux2to1106_and1;
  assign arrdiv12_mux2to1107_and0 = arrdiv12_mux2to195_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1107_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1107_and1 = arrdiv12_fs116_xor1 & arrdiv12_mux2to1107_not0;
  assign arrdiv12_mux2to1107_xor0 = arrdiv12_mux2to1107_and0 ^ arrdiv12_mux2to1107_and1;
  assign arrdiv12_mux2to1108_and0 = arrdiv12_mux2to196_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1108_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1108_and1 = arrdiv12_fs117_xor1 & arrdiv12_mux2to1108_not0;
  assign arrdiv12_mux2to1108_xor0 = arrdiv12_mux2to1108_and0 ^ arrdiv12_mux2to1108_and1;
  assign arrdiv12_mux2to1109_and0 = arrdiv12_mux2to197_xor0 & arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1109_not0 = ~arrdiv12_fs119_or0;
  assign arrdiv12_mux2to1109_and1 = arrdiv12_fs118_xor1 & arrdiv12_mux2to1109_not0;
  assign arrdiv12_mux2to1109_xor0 = arrdiv12_mux2to1109_and0 ^ arrdiv12_mux2to1109_and1;
  assign arrdiv12_not9 = ~arrdiv12_fs119_or0;
  assign arrdiv12_fs120_xor0 = a[1] ^ b[0];
  assign arrdiv12_fs120_not0 = ~a[1];
  assign arrdiv12_fs120_and0 = arrdiv12_fs120_not0 & b[0];
  assign arrdiv12_fs120_not1 = ~arrdiv12_fs120_xor0;
  assign arrdiv12_fs121_xor0 = arrdiv12_mux2to199_xor0 ^ b[1];
  assign arrdiv12_fs121_not0 = ~arrdiv12_mux2to199_xor0;
  assign arrdiv12_fs121_and0 = arrdiv12_fs121_not0 & b[1];
  assign arrdiv12_fs121_xor1 = arrdiv12_fs120_and0 ^ arrdiv12_fs121_xor0;
  assign arrdiv12_fs121_not1 = ~arrdiv12_fs121_xor0;
  assign arrdiv12_fs121_and1 = arrdiv12_fs121_not1 & arrdiv12_fs120_and0;
  assign arrdiv12_fs121_or0 = arrdiv12_fs121_and1 | arrdiv12_fs121_and0;
  assign arrdiv12_fs122_xor0 = arrdiv12_mux2to1100_xor0 ^ b[2];
  assign arrdiv12_fs122_not0 = ~arrdiv12_mux2to1100_xor0;
  assign arrdiv12_fs122_and0 = arrdiv12_fs122_not0 & b[2];
  assign arrdiv12_fs122_xor1 = arrdiv12_fs121_or0 ^ arrdiv12_fs122_xor0;
  assign arrdiv12_fs122_not1 = ~arrdiv12_fs122_xor0;
  assign arrdiv12_fs122_and1 = arrdiv12_fs122_not1 & arrdiv12_fs121_or0;
  assign arrdiv12_fs122_or0 = arrdiv12_fs122_and1 | arrdiv12_fs122_and0;
  assign arrdiv12_fs123_xor0 = arrdiv12_mux2to1101_xor0 ^ b[3];
  assign arrdiv12_fs123_not0 = ~arrdiv12_mux2to1101_xor0;
  assign arrdiv12_fs123_and0 = arrdiv12_fs123_not0 & b[3];
  assign arrdiv12_fs123_xor1 = arrdiv12_fs122_or0 ^ arrdiv12_fs123_xor0;
  assign arrdiv12_fs123_not1 = ~arrdiv12_fs123_xor0;
  assign arrdiv12_fs123_and1 = arrdiv12_fs123_not1 & arrdiv12_fs122_or0;
  assign arrdiv12_fs123_or0 = arrdiv12_fs123_and1 | arrdiv12_fs123_and0;
  assign arrdiv12_fs124_xor0 = arrdiv12_mux2to1102_xor0 ^ b[4];
  assign arrdiv12_fs124_not0 = ~arrdiv12_mux2to1102_xor0;
  assign arrdiv12_fs124_and0 = arrdiv12_fs124_not0 & b[4];
  assign arrdiv12_fs124_xor1 = arrdiv12_fs123_or0 ^ arrdiv12_fs124_xor0;
  assign arrdiv12_fs124_not1 = ~arrdiv12_fs124_xor0;
  assign arrdiv12_fs124_and1 = arrdiv12_fs124_not1 & arrdiv12_fs123_or0;
  assign arrdiv12_fs124_or0 = arrdiv12_fs124_and1 | arrdiv12_fs124_and0;
  assign arrdiv12_fs125_xor0 = arrdiv12_mux2to1103_xor0 ^ b[5];
  assign arrdiv12_fs125_not0 = ~arrdiv12_mux2to1103_xor0;
  assign arrdiv12_fs125_and0 = arrdiv12_fs125_not0 & b[5];
  assign arrdiv12_fs125_xor1 = arrdiv12_fs124_or0 ^ arrdiv12_fs125_xor0;
  assign arrdiv12_fs125_not1 = ~arrdiv12_fs125_xor0;
  assign arrdiv12_fs125_and1 = arrdiv12_fs125_not1 & arrdiv12_fs124_or0;
  assign arrdiv12_fs125_or0 = arrdiv12_fs125_and1 | arrdiv12_fs125_and0;
  assign arrdiv12_fs126_xor0 = arrdiv12_mux2to1104_xor0 ^ b[6];
  assign arrdiv12_fs126_not0 = ~arrdiv12_mux2to1104_xor0;
  assign arrdiv12_fs126_and0 = arrdiv12_fs126_not0 & b[6];
  assign arrdiv12_fs126_xor1 = arrdiv12_fs125_or0 ^ arrdiv12_fs126_xor0;
  assign arrdiv12_fs126_not1 = ~arrdiv12_fs126_xor0;
  assign arrdiv12_fs126_and1 = arrdiv12_fs126_not1 & arrdiv12_fs125_or0;
  assign arrdiv12_fs126_or0 = arrdiv12_fs126_and1 | arrdiv12_fs126_and0;
  assign arrdiv12_fs127_xor0 = arrdiv12_mux2to1105_xor0 ^ b[7];
  assign arrdiv12_fs127_not0 = ~arrdiv12_mux2to1105_xor0;
  assign arrdiv12_fs127_and0 = arrdiv12_fs127_not0 & b[7];
  assign arrdiv12_fs127_xor1 = arrdiv12_fs126_or0 ^ arrdiv12_fs127_xor0;
  assign arrdiv12_fs127_not1 = ~arrdiv12_fs127_xor0;
  assign arrdiv12_fs127_and1 = arrdiv12_fs127_not1 & arrdiv12_fs126_or0;
  assign arrdiv12_fs127_or0 = arrdiv12_fs127_and1 | arrdiv12_fs127_and0;
  assign arrdiv12_fs128_xor0 = arrdiv12_mux2to1106_xor0 ^ b[8];
  assign arrdiv12_fs128_not0 = ~arrdiv12_mux2to1106_xor0;
  assign arrdiv12_fs128_and0 = arrdiv12_fs128_not0 & b[8];
  assign arrdiv12_fs128_xor1 = arrdiv12_fs127_or0 ^ arrdiv12_fs128_xor0;
  assign arrdiv12_fs128_not1 = ~arrdiv12_fs128_xor0;
  assign arrdiv12_fs128_and1 = arrdiv12_fs128_not1 & arrdiv12_fs127_or0;
  assign arrdiv12_fs128_or0 = arrdiv12_fs128_and1 | arrdiv12_fs128_and0;
  assign arrdiv12_fs129_xor0 = arrdiv12_mux2to1107_xor0 ^ b[9];
  assign arrdiv12_fs129_not0 = ~arrdiv12_mux2to1107_xor0;
  assign arrdiv12_fs129_and0 = arrdiv12_fs129_not0 & b[9];
  assign arrdiv12_fs129_xor1 = arrdiv12_fs128_or0 ^ arrdiv12_fs129_xor0;
  assign arrdiv12_fs129_not1 = ~arrdiv12_fs129_xor0;
  assign arrdiv12_fs129_and1 = arrdiv12_fs129_not1 & arrdiv12_fs128_or0;
  assign arrdiv12_fs129_or0 = arrdiv12_fs129_and1 | arrdiv12_fs129_and0;
  assign arrdiv12_fs130_xor0 = arrdiv12_mux2to1108_xor0 ^ b[10];
  assign arrdiv12_fs130_not0 = ~arrdiv12_mux2to1108_xor0;
  assign arrdiv12_fs130_and0 = arrdiv12_fs130_not0 & b[10];
  assign arrdiv12_fs130_xor1 = arrdiv12_fs129_or0 ^ arrdiv12_fs130_xor0;
  assign arrdiv12_fs130_not1 = ~arrdiv12_fs130_xor0;
  assign arrdiv12_fs130_and1 = arrdiv12_fs130_not1 & arrdiv12_fs129_or0;
  assign arrdiv12_fs130_or0 = arrdiv12_fs130_and1 | arrdiv12_fs130_and0;
  assign arrdiv12_fs131_xor0 = arrdiv12_mux2to1109_xor0 ^ b[11];
  assign arrdiv12_fs131_not0 = ~arrdiv12_mux2to1109_xor0;
  assign arrdiv12_fs131_and0 = arrdiv12_fs131_not0 & b[11];
  assign arrdiv12_fs131_xor1 = arrdiv12_fs130_or0 ^ arrdiv12_fs131_xor0;
  assign arrdiv12_fs131_not1 = ~arrdiv12_fs131_xor0;
  assign arrdiv12_fs131_and1 = arrdiv12_fs131_not1 & arrdiv12_fs130_or0;
  assign arrdiv12_fs131_or0 = arrdiv12_fs131_and1 | arrdiv12_fs131_and0;
  assign arrdiv12_mux2to1110_and0 = a[1] & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1110_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1110_and1 = arrdiv12_fs120_xor0 & arrdiv12_mux2to1110_not0;
  assign arrdiv12_mux2to1110_xor0 = arrdiv12_mux2to1110_and0 ^ arrdiv12_mux2to1110_and1;
  assign arrdiv12_mux2to1111_and0 = arrdiv12_mux2to199_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1111_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1111_and1 = arrdiv12_fs121_xor1 & arrdiv12_mux2to1111_not0;
  assign arrdiv12_mux2to1111_xor0 = arrdiv12_mux2to1111_and0 ^ arrdiv12_mux2to1111_and1;
  assign arrdiv12_mux2to1112_and0 = arrdiv12_mux2to1100_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1112_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1112_and1 = arrdiv12_fs122_xor1 & arrdiv12_mux2to1112_not0;
  assign arrdiv12_mux2to1112_xor0 = arrdiv12_mux2to1112_and0 ^ arrdiv12_mux2to1112_and1;
  assign arrdiv12_mux2to1113_and0 = arrdiv12_mux2to1101_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1113_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1113_and1 = arrdiv12_fs123_xor1 & arrdiv12_mux2to1113_not0;
  assign arrdiv12_mux2to1113_xor0 = arrdiv12_mux2to1113_and0 ^ arrdiv12_mux2to1113_and1;
  assign arrdiv12_mux2to1114_and0 = arrdiv12_mux2to1102_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1114_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1114_and1 = arrdiv12_fs124_xor1 & arrdiv12_mux2to1114_not0;
  assign arrdiv12_mux2to1114_xor0 = arrdiv12_mux2to1114_and0 ^ arrdiv12_mux2to1114_and1;
  assign arrdiv12_mux2to1115_and0 = arrdiv12_mux2to1103_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1115_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1115_and1 = arrdiv12_fs125_xor1 & arrdiv12_mux2to1115_not0;
  assign arrdiv12_mux2to1115_xor0 = arrdiv12_mux2to1115_and0 ^ arrdiv12_mux2to1115_and1;
  assign arrdiv12_mux2to1116_and0 = arrdiv12_mux2to1104_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1116_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1116_and1 = arrdiv12_fs126_xor1 & arrdiv12_mux2to1116_not0;
  assign arrdiv12_mux2to1116_xor0 = arrdiv12_mux2to1116_and0 ^ arrdiv12_mux2to1116_and1;
  assign arrdiv12_mux2to1117_and0 = arrdiv12_mux2to1105_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1117_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1117_and1 = arrdiv12_fs127_xor1 & arrdiv12_mux2to1117_not0;
  assign arrdiv12_mux2to1117_xor0 = arrdiv12_mux2to1117_and0 ^ arrdiv12_mux2to1117_and1;
  assign arrdiv12_mux2to1118_and0 = arrdiv12_mux2to1106_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1118_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1118_and1 = arrdiv12_fs128_xor1 & arrdiv12_mux2to1118_not0;
  assign arrdiv12_mux2to1118_xor0 = arrdiv12_mux2to1118_and0 ^ arrdiv12_mux2to1118_and1;
  assign arrdiv12_mux2to1119_and0 = arrdiv12_mux2to1107_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1119_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1119_and1 = arrdiv12_fs129_xor1 & arrdiv12_mux2to1119_not0;
  assign arrdiv12_mux2to1119_xor0 = arrdiv12_mux2to1119_and0 ^ arrdiv12_mux2to1119_and1;
  assign arrdiv12_mux2to1120_and0 = arrdiv12_mux2to1108_xor0 & arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1120_not0 = ~arrdiv12_fs131_or0;
  assign arrdiv12_mux2to1120_and1 = arrdiv12_fs130_xor1 & arrdiv12_mux2to1120_not0;
  assign arrdiv12_mux2to1120_xor0 = arrdiv12_mux2to1120_and0 ^ arrdiv12_mux2to1120_and1;
  assign arrdiv12_not10 = ~arrdiv12_fs131_or0;
  assign arrdiv12_fs132_xor0 = a[0] ^ b[0];
  assign arrdiv12_fs132_not0 = ~a[0];
  assign arrdiv12_fs132_and0 = arrdiv12_fs132_not0 & b[0];
  assign arrdiv12_fs132_not1 = ~arrdiv12_fs132_xor0;
  assign arrdiv12_fs133_xor0 = arrdiv12_mux2to1110_xor0 ^ b[1];
  assign arrdiv12_fs133_not0 = ~arrdiv12_mux2to1110_xor0;
  assign arrdiv12_fs133_and0 = arrdiv12_fs133_not0 & b[1];
  assign arrdiv12_fs133_xor1 = arrdiv12_fs132_and0 ^ arrdiv12_fs133_xor0;
  assign arrdiv12_fs133_not1 = ~arrdiv12_fs133_xor0;
  assign arrdiv12_fs133_and1 = arrdiv12_fs133_not1 & arrdiv12_fs132_and0;
  assign arrdiv12_fs133_or0 = arrdiv12_fs133_and1 | arrdiv12_fs133_and0;
  assign arrdiv12_fs134_xor0 = arrdiv12_mux2to1111_xor0 ^ b[2];
  assign arrdiv12_fs134_not0 = ~arrdiv12_mux2to1111_xor0;
  assign arrdiv12_fs134_and0 = arrdiv12_fs134_not0 & b[2];
  assign arrdiv12_fs134_xor1 = arrdiv12_fs133_or0 ^ arrdiv12_fs134_xor0;
  assign arrdiv12_fs134_not1 = ~arrdiv12_fs134_xor0;
  assign arrdiv12_fs134_and1 = arrdiv12_fs134_not1 & arrdiv12_fs133_or0;
  assign arrdiv12_fs134_or0 = arrdiv12_fs134_and1 | arrdiv12_fs134_and0;
  assign arrdiv12_fs135_xor0 = arrdiv12_mux2to1112_xor0 ^ b[3];
  assign arrdiv12_fs135_not0 = ~arrdiv12_mux2to1112_xor0;
  assign arrdiv12_fs135_and0 = arrdiv12_fs135_not0 & b[3];
  assign arrdiv12_fs135_xor1 = arrdiv12_fs134_or0 ^ arrdiv12_fs135_xor0;
  assign arrdiv12_fs135_not1 = ~arrdiv12_fs135_xor0;
  assign arrdiv12_fs135_and1 = arrdiv12_fs135_not1 & arrdiv12_fs134_or0;
  assign arrdiv12_fs135_or0 = arrdiv12_fs135_and1 | arrdiv12_fs135_and0;
  assign arrdiv12_fs136_xor0 = arrdiv12_mux2to1113_xor0 ^ b[4];
  assign arrdiv12_fs136_not0 = ~arrdiv12_mux2to1113_xor0;
  assign arrdiv12_fs136_and0 = arrdiv12_fs136_not0 & b[4];
  assign arrdiv12_fs136_xor1 = arrdiv12_fs135_or0 ^ arrdiv12_fs136_xor0;
  assign arrdiv12_fs136_not1 = ~arrdiv12_fs136_xor0;
  assign arrdiv12_fs136_and1 = arrdiv12_fs136_not1 & arrdiv12_fs135_or0;
  assign arrdiv12_fs136_or0 = arrdiv12_fs136_and1 | arrdiv12_fs136_and0;
  assign arrdiv12_fs137_xor0 = arrdiv12_mux2to1114_xor0 ^ b[5];
  assign arrdiv12_fs137_not0 = ~arrdiv12_mux2to1114_xor0;
  assign arrdiv12_fs137_and0 = arrdiv12_fs137_not0 & b[5];
  assign arrdiv12_fs137_xor1 = arrdiv12_fs136_or0 ^ arrdiv12_fs137_xor0;
  assign arrdiv12_fs137_not1 = ~arrdiv12_fs137_xor0;
  assign arrdiv12_fs137_and1 = arrdiv12_fs137_not1 & arrdiv12_fs136_or0;
  assign arrdiv12_fs137_or0 = arrdiv12_fs137_and1 | arrdiv12_fs137_and0;
  assign arrdiv12_fs138_xor0 = arrdiv12_mux2to1115_xor0 ^ b[6];
  assign arrdiv12_fs138_not0 = ~arrdiv12_mux2to1115_xor0;
  assign arrdiv12_fs138_and0 = arrdiv12_fs138_not0 & b[6];
  assign arrdiv12_fs138_xor1 = arrdiv12_fs137_or0 ^ arrdiv12_fs138_xor0;
  assign arrdiv12_fs138_not1 = ~arrdiv12_fs138_xor0;
  assign arrdiv12_fs138_and1 = arrdiv12_fs138_not1 & arrdiv12_fs137_or0;
  assign arrdiv12_fs138_or0 = arrdiv12_fs138_and1 | arrdiv12_fs138_and0;
  assign arrdiv12_fs139_xor0 = arrdiv12_mux2to1116_xor0 ^ b[7];
  assign arrdiv12_fs139_not0 = ~arrdiv12_mux2to1116_xor0;
  assign arrdiv12_fs139_and0 = arrdiv12_fs139_not0 & b[7];
  assign arrdiv12_fs139_xor1 = arrdiv12_fs138_or0 ^ arrdiv12_fs139_xor0;
  assign arrdiv12_fs139_not1 = ~arrdiv12_fs139_xor0;
  assign arrdiv12_fs139_and1 = arrdiv12_fs139_not1 & arrdiv12_fs138_or0;
  assign arrdiv12_fs139_or0 = arrdiv12_fs139_and1 | arrdiv12_fs139_and0;
  assign arrdiv12_fs140_xor0 = arrdiv12_mux2to1117_xor0 ^ b[8];
  assign arrdiv12_fs140_not0 = ~arrdiv12_mux2to1117_xor0;
  assign arrdiv12_fs140_and0 = arrdiv12_fs140_not0 & b[8];
  assign arrdiv12_fs140_xor1 = arrdiv12_fs139_or0 ^ arrdiv12_fs140_xor0;
  assign arrdiv12_fs140_not1 = ~arrdiv12_fs140_xor0;
  assign arrdiv12_fs140_and1 = arrdiv12_fs140_not1 & arrdiv12_fs139_or0;
  assign arrdiv12_fs140_or0 = arrdiv12_fs140_and1 | arrdiv12_fs140_and0;
  assign arrdiv12_fs141_xor0 = arrdiv12_mux2to1118_xor0 ^ b[9];
  assign arrdiv12_fs141_not0 = ~arrdiv12_mux2to1118_xor0;
  assign arrdiv12_fs141_and0 = arrdiv12_fs141_not0 & b[9];
  assign arrdiv12_fs141_xor1 = arrdiv12_fs140_or0 ^ arrdiv12_fs141_xor0;
  assign arrdiv12_fs141_not1 = ~arrdiv12_fs141_xor0;
  assign arrdiv12_fs141_and1 = arrdiv12_fs141_not1 & arrdiv12_fs140_or0;
  assign arrdiv12_fs141_or0 = arrdiv12_fs141_and1 | arrdiv12_fs141_and0;
  assign arrdiv12_fs142_xor0 = arrdiv12_mux2to1119_xor0 ^ b[10];
  assign arrdiv12_fs142_not0 = ~arrdiv12_mux2to1119_xor0;
  assign arrdiv12_fs142_and0 = arrdiv12_fs142_not0 & b[10];
  assign arrdiv12_fs142_xor1 = arrdiv12_fs141_or0 ^ arrdiv12_fs142_xor0;
  assign arrdiv12_fs142_not1 = ~arrdiv12_fs142_xor0;
  assign arrdiv12_fs142_and1 = arrdiv12_fs142_not1 & arrdiv12_fs141_or0;
  assign arrdiv12_fs142_or0 = arrdiv12_fs142_and1 | arrdiv12_fs142_and0;
  assign arrdiv12_fs143_xor0 = arrdiv12_mux2to1120_xor0 ^ b[11];
  assign arrdiv12_fs143_not0 = ~arrdiv12_mux2to1120_xor0;
  assign arrdiv12_fs143_and0 = arrdiv12_fs143_not0 & b[11];
  assign arrdiv12_fs143_xor1 = arrdiv12_fs142_or0 ^ arrdiv12_fs143_xor0;
  assign arrdiv12_fs143_not1 = ~arrdiv12_fs143_xor0;
  assign arrdiv12_fs143_and1 = arrdiv12_fs143_not1 & arrdiv12_fs142_or0;
  assign arrdiv12_fs143_or0 = arrdiv12_fs143_and1 | arrdiv12_fs143_and0;
  assign arrdiv12_not11 = ~arrdiv12_fs143_or0;

  assign arrdiv12_out[0] = arrdiv12_not11;
  assign arrdiv12_out[1] = arrdiv12_not10;
  assign arrdiv12_out[2] = arrdiv12_not9;
  assign arrdiv12_out[3] = arrdiv12_not8;
  assign arrdiv12_out[4] = arrdiv12_not7;
  assign arrdiv12_out[5] = arrdiv12_not6;
  assign arrdiv12_out[6] = arrdiv12_not5;
  assign arrdiv12_out[7] = arrdiv12_not4;
  assign arrdiv12_out[8] = arrdiv12_not3;
  assign arrdiv12_out[9] = arrdiv12_not2;
  assign arrdiv12_out[10] = arrdiv12_not1;
  assign arrdiv12_out[11] = arrdiv12_not0;
endmodule