module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_cin;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module u_rca(input [45:0] a, input [45:0] b, output [46:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire a_30;
  wire a_31;
  wire a_32;
  wire a_33;
  wire a_34;
  wire a_35;
  wire a_36;
  wire a_37;
  wire a_38;
  wire a_39;
  wire a_40;
  wire a_41;
  wire a_42;
  wire a_43;
  wire a_44;
  wire a_45;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire b_30;
  wire b_31;
  wire b_32;
  wire b_33;
  wire b_34;
  wire b_35;
  wire b_36;
  wire b_37;
  wire b_38;
  wire b_39;
  wire b_40;
  wire b_41;
  wire b_42;
  wire b_43;
  wire b_44;
  wire b_45;
  wire u_rca_ha_y0;
  wire u_rca_ha_y1;
  wire u_rca_fa1_y2;
  wire u_rca_fa1_y4;
  wire u_rca_fa2_y2;
  wire u_rca_fa2_y4;
  wire u_rca_fa3_y2;
  wire u_rca_fa3_y4;
  wire u_rca_fa4_y2;
  wire u_rca_fa4_y4;
  wire u_rca_fa5_y2;
  wire u_rca_fa5_y4;
  wire u_rca_fa6_y2;
  wire u_rca_fa6_y4;
  wire u_rca_fa7_y2;
  wire u_rca_fa7_y4;
  wire u_rca_fa8_y2;
  wire u_rca_fa8_y4;
  wire u_rca_fa9_y2;
  wire u_rca_fa9_y4;
  wire u_rca_fa10_y2;
  wire u_rca_fa10_y4;
  wire u_rca_fa11_y2;
  wire u_rca_fa11_y4;
  wire u_rca_fa12_y2;
  wire u_rca_fa12_y4;
  wire u_rca_fa13_y2;
  wire u_rca_fa13_y4;
  wire u_rca_fa14_y2;
  wire u_rca_fa14_y4;
  wire u_rca_fa15_y2;
  wire u_rca_fa15_y4;
  wire u_rca_fa16_y2;
  wire u_rca_fa16_y4;
  wire u_rca_fa17_y2;
  wire u_rca_fa17_y4;
  wire u_rca_fa18_y2;
  wire u_rca_fa18_y4;
  wire u_rca_fa19_y2;
  wire u_rca_fa19_y4;
  wire u_rca_fa20_y2;
  wire u_rca_fa20_y4;
  wire u_rca_fa21_y2;
  wire u_rca_fa21_y4;
  wire u_rca_fa22_y2;
  wire u_rca_fa22_y4;
  wire u_rca_fa23_y2;
  wire u_rca_fa23_y4;
  wire u_rca_fa24_y2;
  wire u_rca_fa24_y4;
  wire u_rca_fa25_y2;
  wire u_rca_fa25_y4;
  wire u_rca_fa26_y2;
  wire u_rca_fa26_y4;
  wire u_rca_fa27_y2;
  wire u_rca_fa27_y4;
  wire u_rca_fa28_y2;
  wire u_rca_fa28_y4;
  wire u_rca_fa29_y2;
  wire u_rca_fa29_y4;
  wire u_rca_fa30_y2;
  wire u_rca_fa30_y4;
  wire u_rca_fa31_y2;
  wire u_rca_fa31_y4;
  wire u_rca_fa32_y2;
  wire u_rca_fa32_y4;
  wire u_rca_fa33_y2;
  wire u_rca_fa33_y4;
  wire u_rca_fa34_y2;
  wire u_rca_fa34_y4;
  wire u_rca_fa35_y2;
  wire u_rca_fa35_y4;
  wire u_rca_fa36_y2;
  wire u_rca_fa36_y4;
  wire u_rca_fa37_y2;
  wire u_rca_fa37_y4;
  wire u_rca_fa38_y2;
  wire u_rca_fa38_y4;
  wire u_rca_fa39_y2;
  wire u_rca_fa39_y4;
  wire u_rca_fa40_y2;
  wire u_rca_fa40_y4;
  wire u_rca_fa41_y2;
  wire u_rca_fa41_y4;
  wire u_rca_fa42_y2;
  wire u_rca_fa42_y4;
  wire u_rca_fa43_y2;
  wire u_rca_fa43_y4;
  wire u_rca_fa44_y2;
  wire u_rca_fa44_y4;
  wire u_rca_fa45_y2;
  wire u_rca_fa45_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign a_30 = a[30];
  assign a_31 = a[31];
  assign a_32 = a[32];
  assign a_33 = a[33];
  assign a_34 = a[34];
  assign a_35 = a[35];
  assign a_36 = a[36];
  assign a_37 = a[37];
  assign a_38 = a[38];
  assign a_39 = a[39];
  assign a_40 = a[40];
  assign a_41 = a[41];
  assign a_42 = a[42];
  assign a_43 = a[43];
  assign a_44 = a[44];
  assign a_45 = a[45];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  assign b_30 = b[30];
  assign b_31 = b[31];
  assign b_32 = b[32];
  assign b_33 = b[33];
  assign b_34 = b[34];
  assign b_35 = b[35];
  assign b_36 = b[36];
  assign b_37 = b[37];
  assign b_38 = b[38];
  assign b_39 = b[39];
  assign b_40 = b[40];
  assign b_41 = b[41];
  assign b_42 = b[42];
  assign b_43 = b[43];
  assign b_44 = b[44];
  assign b_45 = b[45];
  ha ha_u_rca_ha_y0(a_0, b_0, u_rca_ha_y0, u_rca_ha_y1);
  fa fa_u_rca_fa1_y2(a_1, b_1, u_rca_ha_y1, u_rca_fa1_y2, u_rca_fa1_y4);
  fa fa_u_rca_fa2_y2(a_2, b_2, u_rca_fa1_y4, u_rca_fa2_y2, u_rca_fa2_y4);
  fa fa_u_rca_fa3_y2(a_3, b_3, u_rca_fa2_y4, u_rca_fa3_y2, u_rca_fa3_y4);
  fa fa_u_rca_fa4_y2(a_4, b_4, u_rca_fa3_y4, u_rca_fa4_y2, u_rca_fa4_y4);
  fa fa_u_rca_fa5_y2(a_5, b_5, u_rca_fa4_y4, u_rca_fa5_y2, u_rca_fa5_y4);
  fa fa_u_rca_fa6_y2(a_6, b_6, u_rca_fa5_y4, u_rca_fa6_y2, u_rca_fa6_y4);
  fa fa_u_rca_fa7_y2(a_7, b_7, u_rca_fa6_y4, u_rca_fa7_y2, u_rca_fa7_y4);
  fa fa_u_rca_fa8_y2(a_8, b_8, u_rca_fa7_y4, u_rca_fa8_y2, u_rca_fa8_y4);
  fa fa_u_rca_fa9_y2(a_9, b_9, u_rca_fa8_y4, u_rca_fa9_y2, u_rca_fa9_y4);
  fa fa_u_rca_fa10_y2(a_10, b_10, u_rca_fa9_y4, u_rca_fa10_y2, u_rca_fa10_y4);
  fa fa_u_rca_fa11_y2(a_11, b_11, u_rca_fa10_y4, u_rca_fa11_y2, u_rca_fa11_y4);
  fa fa_u_rca_fa12_y2(a_12, b_12, u_rca_fa11_y4, u_rca_fa12_y2, u_rca_fa12_y4);
  fa fa_u_rca_fa13_y2(a_13, b_13, u_rca_fa12_y4, u_rca_fa13_y2, u_rca_fa13_y4);
  fa fa_u_rca_fa14_y2(a_14, b_14, u_rca_fa13_y4, u_rca_fa14_y2, u_rca_fa14_y4);
  fa fa_u_rca_fa15_y2(a_15, b_15, u_rca_fa14_y4, u_rca_fa15_y2, u_rca_fa15_y4);
  fa fa_u_rca_fa16_y2(a_16, b_16, u_rca_fa15_y4, u_rca_fa16_y2, u_rca_fa16_y4);
  fa fa_u_rca_fa17_y2(a_17, b_17, u_rca_fa16_y4, u_rca_fa17_y2, u_rca_fa17_y4);
  fa fa_u_rca_fa18_y2(a_18, b_18, u_rca_fa17_y4, u_rca_fa18_y2, u_rca_fa18_y4);
  fa fa_u_rca_fa19_y2(a_19, b_19, u_rca_fa18_y4, u_rca_fa19_y2, u_rca_fa19_y4);
  fa fa_u_rca_fa20_y2(a_20, b_20, u_rca_fa19_y4, u_rca_fa20_y2, u_rca_fa20_y4);
  fa fa_u_rca_fa21_y2(a_21, b_21, u_rca_fa20_y4, u_rca_fa21_y2, u_rca_fa21_y4);
  fa fa_u_rca_fa22_y2(a_22, b_22, u_rca_fa21_y4, u_rca_fa22_y2, u_rca_fa22_y4);
  fa fa_u_rca_fa23_y2(a_23, b_23, u_rca_fa22_y4, u_rca_fa23_y2, u_rca_fa23_y4);
  fa fa_u_rca_fa24_y2(a_24, b_24, u_rca_fa23_y4, u_rca_fa24_y2, u_rca_fa24_y4);
  fa fa_u_rca_fa25_y2(a_25, b_25, u_rca_fa24_y4, u_rca_fa25_y2, u_rca_fa25_y4);
  fa fa_u_rca_fa26_y2(a_26, b_26, u_rca_fa25_y4, u_rca_fa26_y2, u_rca_fa26_y4);
  fa fa_u_rca_fa27_y2(a_27, b_27, u_rca_fa26_y4, u_rca_fa27_y2, u_rca_fa27_y4);
  fa fa_u_rca_fa28_y2(a_28, b_28, u_rca_fa27_y4, u_rca_fa28_y2, u_rca_fa28_y4);
  fa fa_u_rca_fa29_y2(a_29, b_29, u_rca_fa28_y4, u_rca_fa29_y2, u_rca_fa29_y4);
  fa fa_u_rca_fa30_y2(a_30, b_30, u_rca_fa29_y4, u_rca_fa30_y2, u_rca_fa30_y4);
  fa fa_u_rca_fa31_y2(a_31, b_31, u_rca_fa30_y4, u_rca_fa31_y2, u_rca_fa31_y4);
  fa fa_u_rca_fa32_y2(a_32, b_32, u_rca_fa31_y4, u_rca_fa32_y2, u_rca_fa32_y4);
  fa fa_u_rca_fa33_y2(a_33, b_33, u_rca_fa32_y4, u_rca_fa33_y2, u_rca_fa33_y4);
  fa fa_u_rca_fa34_y2(a_34, b_34, u_rca_fa33_y4, u_rca_fa34_y2, u_rca_fa34_y4);
  fa fa_u_rca_fa35_y2(a_35, b_35, u_rca_fa34_y4, u_rca_fa35_y2, u_rca_fa35_y4);
  fa fa_u_rca_fa36_y2(a_36, b_36, u_rca_fa35_y4, u_rca_fa36_y2, u_rca_fa36_y4);
  fa fa_u_rca_fa37_y2(a_37, b_37, u_rca_fa36_y4, u_rca_fa37_y2, u_rca_fa37_y4);
  fa fa_u_rca_fa38_y2(a_38, b_38, u_rca_fa37_y4, u_rca_fa38_y2, u_rca_fa38_y4);
  fa fa_u_rca_fa39_y2(a_39, b_39, u_rca_fa38_y4, u_rca_fa39_y2, u_rca_fa39_y4);
  fa fa_u_rca_fa40_y2(a_40, b_40, u_rca_fa39_y4, u_rca_fa40_y2, u_rca_fa40_y4);
  fa fa_u_rca_fa41_y2(a_41, b_41, u_rca_fa40_y4, u_rca_fa41_y2, u_rca_fa41_y4);
  fa fa_u_rca_fa42_y2(a_42, b_42, u_rca_fa41_y4, u_rca_fa42_y2, u_rca_fa42_y4);
  fa fa_u_rca_fa43_y2(a_43, b_43, u_rca_fa42_y4, u_rca_fa43_y2, u_rca_fa43_y4);
  fa fa_u_rca_fa44_y2(a_44, b_44, u_rca_fa43_y4, u_rca_fa44_y2, u_rca_fa44_y4);
  fa fa_u_rca_fa45_y2(a_45, b_45, u_rca_fa44_y4, u_rca_fa45_y2, u_rca_fa45_y4);

  assign out[0] = u_rca_ha_y0;
  assign out[1] = u_rca_fa1_y2;
  assign out[2] = u_rca_fa2_y2;
  assign out[3] = u_rca_fa3_y2;
  assign out[4] = u_rca_fa4_y2;
  assign out[5] = u_rca_fa5_y2;
  assign out[6] = u_rca_fa6_y2;
  assign out[7] = u_rca_fa7_y2;
  assign out[8] = u_rca_fa8_y2;
  assign out[9] = u_rca_fa9_y2;
  assign out[10] = u_rca_fa10_y2;
  assign out[11] = u_rca_fa11_y2;
  assign out[12] = u_rca_fa12_y2;
  assign out[13] = u_rca_fa13_y2;
  assign out[14] = u_rca_fa14_y2;
  assign out[15] = u_rca_fa15_y2;
  assign out[16] = u_rca_fa16_y2;
  assign out[17] = u_rca_fa17_y2;
  assign out[18] = u_rca_fa18_y2;
  assign out[19] = u_rca_fa19_y2;
  assign out[20] = u_rca_fa20_y2;
  assign out[21] = u_rca_fa21_y2;
  assign out[22] = u_rca_fa22_y2;
  assign out[23] = u_rca_fa23_y2;
  assign out[24] = u_rca_fa24_y2;
  assign out[25] = u_rca_fa25_y2;
  assign out[26] = u_rca_fa26_y2;
  assign out[27] = u_rca_fa27_y2;
  assign out[28] = u_rca_fa28_y2;
  assign out[29] = u_rca_fa29_y2;
  assign out[30] = u_rca_fa30_y2;
  assign out[31] = u_rca_fa31_y2;
  assign out[32] = u_rca_fa32_y2;
  assign out[33] = u_rca_fa33_y2;
  assign out[34] = u_rca_fa34_y2;
  assign out[35] = u_rca_fa35_y2;
  assign out[36] = u_rca_fa36_y2;
  assign out[37] = u_rca_fa37_y2;
  assign out[38] = u_rca_fa38_y2;
  assign out[39] = u_rca_fa39_y2;
  assign out[40] = u_rca_fa40_y2;
  assign out[41] = u_rca_fa41_y2;
  assign out[42] = u_rca_fa42_y2;
  assign out[43] = u_rca_fa43_y2;
  assign out[44] = u_rca_fa44_y2;
  assign out[45] = u_rca_fa45_y2;
  assign out[46] = u_rca_fa45_y4;
endmodule

module h_s_wallace_rca24(input [23:0] a, input [23:0] b, output [47:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire constant_wire_1;
  wire h_s_wallace_rca24_and_2_0_y0;
  wire h_s_wallace_rca24_and_1_1_y0;
  wire h_s_wallace_rca24_ha0_y0;
  wire h_s_wallace_rca24_ha0_y1;
  wire h_s_wallace_rca24_and_3_0_y0;
  wire h_s_wallace_rca24_and_2_1_y0;
  wire h_s_wallace_rca24_fa0_y2;
  wire h_s_wallace_rca24_fa0_y4;
  wire h_s_wallace_rca24_and_4_0_y0;
  wire h_s_wallace_rca24_and_3_1_y0;
  wire h_s_wallace_rca24_fa1_y2;
  wire h_s_wallace_rca24_fa1_y4;
  wire h_s_wallace_rca24_and_5_0_y0;
  wire h_s_wallace_rca24_and_4_1_y0;
  wire h_s_wallace_rca24_fa2_y2;
  wire h_s_wallace_rca24_fa2_y4;
  wire h_s_wallace_rca24_and_6_0_y0;
  wire h_s_wallace_rca24_and_5_1_y0;
  wire h_s_wallace_rca24_fa3_y2;
  wire h_s_wallace_rca24_fa3_y4;
  wire h_s_wallace_rca24_and_7_0_y0;
  wire h_s_wallace_rca24_and_6_1_y0;
  wire h_s_wallace_rca24_fa4_y2;
  wire h_s_wallace_rca24_fa4_y4;
  wire h_s_wallace_rca24_and_8_0_y0;
  wire h_s_wallace_rca24_and_7_1_y0;
  wire h_s_wallace_rca24_fa5_y2;
  wire h_s_wallace_rca24_fa5_y4;
  wire h_s_wallace_rca24_and_9_0_y0;
  wire h_s_wallace_rca24_and_8_1_y0;
  wire h_s_wallace_rca24_fa6_y2;
  wire h_s_wallace_rca24_fa6_y4;
  wire h_s_wallace_rca24_and_10_0_y0;
  wire h_s_wallace_rca24_and_9_1_y0;
  wire h_s_wallace_rca24_fa7_y2;
  wire h_s_wallace_rca24_fa7_y4;
  wire h_s_wallace_rca24_and_11_0_y0;
  wire h_s_wallace_rca24_and_10_1_y0;
  wire h_s_wallace_rca24_fa8_y2;
  wire h_s_wallace_rca24_fa8_y4;
  wire h_s_wallace_rca24_and_12_0_y0;
  wire h_s_wallace_rca24_and_11_1_y0;
  wire h_s_wallace_rca24_fa9_y2;
  wire h_s_wallace_rca24_fa9_y4;
  wire h_s_wallace_rca24_and_13_0_y0;
  wire h_s_wallace_rca24_and_12_1_y0;
  wire h_s_wallace_rca24_fa10_y2;
  wire h_s_wallace_rca24_fa10_y4;
  wire h_s_wallace_rca24_and_14_0_y0;
  wire h_s_wallace_rca24_and_13_1_y0;
  wire h_s_wallace_rca24_fa11_y2;
  wire h_s_wallace_rca24_fa11_y4;
  wire h_s_wallace_rca24_and_15_0_y0;
  wire h_s_wallace_rca24_and_14_1_y0;
  wire h_s_wallace_rca24_fa12_y2;
  wire h_s_wallace_rca24_fa12_y4;
  wire h_s_wallace_rca24_and_16_0_y0;
  wire h_s_wallace_rca24_and_15_1_y0;
  wire h_s_wallace_rca24_fa13_y2;
  wire h_s_wallace_rca24_fa13_y4;
  wire h_s_wallace_rca24_and_17_0_y0;
  wire h_s_wallace_rca24_and_16_1_y0;
  wire h_s_wallace_rca24_fa14_y2;
  wire h_s_wallace_rca24_fa14_y4;
  wire h_s_wallace_rca24_and_18_0_y0;
  wire h_s_wallace_rca24_and_17_1_y0;
  wire h_s_wallace_rca24_fa15_y2;
  wire h_s_wallace_rca24_fa15_y4;
  wire h_s_wallace_rca24_and_19_0_y0;
  wire h_s_wallace_rca24_and_18_1_y0;
  wire h_s_wallace_rca24_fa16_y2;
  wire h_s_wallace_rca24_fa16_y4;
  wire h_s_wallace_rca24_and_20_0_y0;
  wire h_s_wallace_rca24_and_19_1_y0;
  wire h_s_wallace_rca24_fa17_y2;
  wire h_s_wallace_rca24_fa17_y4;
  wire h_s_wallace_rca24_and_21_0_y0;
  wire h_s_wallace_rca24_and_20_1_y0;
  wire h_s_wallace_rca24_fa18_y2;
  wire h_s_wallace_rca24_fa18_y4;
  wire h_s_wallace_rca24_and_22_0_y0;
  wire h_s_wallace_rca24_and_21_1_y0;
  wire h_s_wallace_rca24_fa19_y2;
  wire h_s_wallace_rca24_fa19_y4;
  wire h_s_wallace_rca24_nand_23_0_y0;
  wire h_s_wallace_rca24_and_22_1_y0;
  wire h_s_wallace_rca24_fa20_y2;
  wire h_s_wallace_rca24_fa20_y4;
  wire h_s_wallace_rca24_nand_23_1_y0;
  wire h_s_wallace_rca24_fa21_y2;
  wire h_s_wallace_rca24_fa21_y4;
  wire h_s_wallace_rca24_nand_23_2_y0;
  wire h_s_wallace_rca24_and_22_3_y0;
  wire h_s_wallace_rca24_fa22_y2;
  wire h_s_wallace_rca24_fa22_y4;
  wire h_s_wallace_rca24_nand_23_3_y0;
  wire h_s_wallace_rca24_and_22_4_y0;
  wire h_s_wallace_rca24_fa23_y2;
  wire h_s_wallace_rca24_fa23_y4;
  wire h_s_wallace_rca24_nand_23_4_y0;
  wire h_s_wallace_rca24_and_22_5_y0;
  wire h_s_wallace_rca24_fa24_y2;
  wire h_s_wallace_rca24_fa24_y4;
  wire h_s_wallace_rca24_nand_23_5_y0;
  wire h_s_wallace_rca24_and_22_6_y0;
  wire h_s_wallace_rca24_fa25_y2;
  wire h_s_wallace_rca24_fa25_y4;
  wire h_s_wallace_rca24_nand_23_6_y0;
  wire h_s_wallace_rca24_and_22_7_y0;
  wire h_s_wallace_rca24_fa26_y2;
  wire h_s_wallace_rca24_fa26_y4;
  wire h_s_wallace_rca24_nand_23_7_y0;
  wire h_s_wallace_rca24_and_22_8_y0;
  wire h_s_wallace_rca24_fa27_y2;
  wire h_s_wallace_rca24_fa27_y4;
  wire h_s_wallace_rca24_nand_23_8_y0;
  wire h_s_wallace_rca24_and_22_9_y0;
  wire h_s_wallace_rca24_fa28_y2;
  wire h_s_wallace_rca24_fa28_y4;
  wire h_s_wallace_rca24_nand_23_9_y0;
  wire h_s_wallace_rca24_and_22_10_y0;
  wire h_s_wallace_rca24_fa29_y2;
  wire h_s_wallace_rca24_fa29_y4;
  wire h_s_wallace_rca24_nand_23_10_y0;
  wire h_s_wallace_rca24_and_22_11_y0;
  wire h_s_wallace_rca24_fa30_y2;
  wire h_s_wallace_rca24_fa30_y4;
  wire h_s_wallace_rca24_nand_23_11_y0;
  wire h_s_wallace_rca24_and_22_12_y0;
  wire h_s_wallace_rca24_fa31_y2;
  wire h_s_wallace_rca24_fa31_y4;
  wire h_s_wallace_rca24_nand_23_12_y0;
  wire h_s_wallace_rca24_and_22_13_y0;
  wire h_s_wallace_rca24_fa32_y2;
  wire h_s_wallace_rca24_fa32_y4;
  wire h_s_wallace_rca24_nand_23_13_y0;
  wire h_s_wallace_rca24_and_22_14_y0;
  wire h_s_wallace_rca24_fa33_y2;
  wire h_s_wallace_rca24_fa33_y4;
  wire h_s_wallace_rca24_nand_23_14_y0;
  wire h_s_wallace_rca24_and_22_15_y0;
  wire h_s_wallace_rca24_fa34_y2;
  wire h_s_wallace_rca24_fa34_y4;
  wire h_s_wallace_rca24_nand_23_15_y0;
  wire h_s_wallace_rca24_and_22_16_y0;
  wire h_s_wallace_rca24_fa35_y2;
  wire h_s_wallace_rca24_fa35_y4;
  wire h_s_wallace_rca24_nand_23_16_y0;
  wire h_s_wallace_rca24_and_22_17_y0;
  wire h_s_wallace_rca24_fa36_y2;
  wire h_s_wallace_rca24_fa36_y4;
  wire h_s_wallace_rca24_nand_23_17_y0;
  wire h_s_wallace_rca24_and_22_18_y0;
  wire h_s_wallace_rca24_fa37_y2;
  wire h_s_wallace_rca24_fa37_y4;
  wire h_s_wallace_rca24_nand_23_18_y0;
  wire h_s_wallace_rca24_and_22_19_y0;
  wire h_s_wallace_rca24_fa38_y2;
  wire h_s_wallace_rca24_fa38_y4;
  wire h_s_wallace_rca24_nand_23_19_y0;
  wire h_s_wallace_rca24_and_22_20_y0;
  wire h_s_wallace_rca24_fa39_y2;
  wire h_s_wallace_rca24_fa39_y4;
  wire h_s_wallace_rca24_nand_23_20_y0;
  wire h_s_wallace_rca24_and_22_21_y0;
  wire h_s_wallace_rca24_fa40_y2;
  wire h_s_wallace_rca24_fa40_y4;
  wire h_s_wallace_rca24_nand_23_21_y0;
  wire h_s_wallace_rca24_and_22_22_y0;
  wire h_s_wallace_rca24_fa41_y2;
  wire h_s_wallace_rca24_fa41_y4;
  wire h_s_wallace_rca24_and_1_2_y0;
  wire h_s_wallace_rca24_and_0_3_y0;
  wire h_s_wallace_rca24_ha1_y0;
  wire h_s_wallace_rca24_ha1_y1;
  wire h_s_wallace_rca24_and_2_2_y0;
  wire h_s_wallace_rca24_and_1_3_y0;
  wire h_s_wallace_rca24_fa42_y2;
  wire h_s_wallace_rca24_fa42_y4;
  wire h_s_wallace_rca24_and_3_2_y0;
  wire h_s_wallace_rca24_and_2_3_y0;
  wire h_s_wallace_rca24_fa43_y2;
  wire h_s_wallace_rca24_fa43_y4;
  wire h_s_wallace_rca24_and_4_2_y0;
  wire h_s_wallace_rca24_and_3_3_y0;
  wire h_s_wallace_rca24_fa44_y2;
  wire h_s_wallace_rca24_fa44_y4;
  wire h_s_wallace_rca24_and_5_2_y0;
  wire h_s_wallace_rca24_and_4_3_y0;
  wire h_s_wallace_rca24_fa45_y2;
  wire h_s_wallace_rca24_fa45_y4;
  wire h_s_wallace_rca24_and_6_2_y0;
  wire h_s_wallace_rca24_and_5_3_y0;
  wire h_s_wallace_rca24_fa46_y2;
  wire h_s_wallace_rca24_fa46_y4;
  wire h_s_wallace_rca24_and_7_2_y0;
  wire h_s_wallace_rca24_and_6_3_y0;
  wire h_s_wallace_rca24_fa47_y2;
  wire h_s_wallace_rca24_fa47_y4;
  wire h_s_wallace_rca24_and_8_2_y0;
  wire h_s_wallace_rca24_and_7_3_y0;
  wire h_s_wallace_rca24_fa48_y2;
  wire h_s_wallace_rca24_fa48_y4;
  wire h_s_wallace_rca24_and_9_2_y0;
  wire h_s_wallace_rca24_and_8_3_y0;
  wire h_s_wallace_rca24_fa49_y2;
  wire h_s_wallace_rca24_fa49_y4;
  wire h_s_wallace_rca24_and_10_2_y0;
  wire h_s_wallace_rca24_and_9_3_y0;
  wire h_s_wallace_rca24_fa50_y2;
  wire h_s_wallace_rca24_fa50_y4;
  wire h_s_wallace_rca24_and_11_2_y0;
  wire h_s_wallace_rca24_and_10_3_y0;
  wire h_s_wallace_rca24_fa51_y2;
  wire h_s_wallace_rca24_fa51_y4;
  wire h_s_wallace_rca24_and_12_2_y0;
  wire h_s_wallace_rca24_and_11_3_y0;
  wire h_s_wallace_rca24_fa52_y2;
  wire h_s_wallace_rca24_fa52_y4;
  wire h_s_wallace_rca24_and_13_2_y0;
  wire h_s_wallace_rca24_and_12_3_y0;
  wire h_s_wallace_rca24_fa53_y2;
  wire h_s_wallace_rca24_fa53_y4;
  wire h_s_wallace_rca24_and_14_2_y0;
  wire h_s_wallace_rca24_and_13_3_y0;
  wire h_s_wallace_rca24_fa54_y2;
  wire h_s_wallace_rca24_fa54_y4;
  wire h_s_wallace_rca24_and_15_2_y0;
  wire h_s_wallace_rca24_and_14_3_y0;
  wire h_s_wallace_rca24_fa55_y2;
  wire h_s_wallace_rca24_fa55_y4;
  wire h_s_wallace_rca24_and_16_2_y0;
  wire h_s_wallace_rca24_and_15_3_y0;
  wire h_s_wallace_rca24_fa56_y2;
  wire h_s_wallace_rca24_fa56_y4;
  wire h_s_wallace_rca24_and_17_2_y0;
  wire h_s_wallace_rca24_and_16_3_y0;
  wire h_s_wallace_rca24_fa57_y2;
  wire h_s_wallace_rca24_fa57_y4;
  wire h_s_wallace_rca24_and_18_2_y0;
  wire h_s_wallace_rca24_and_17_3_y0;
  wire h_s_wallace_rca24_fa58_y2;
  wire h_s_wallace_rca24_fa58_y4;
  wire h_s_wallace_rca24_and_19_2_y0;
  wire h_s_wallace_rca24_and_18_3_y0;
  wire h_s_wallace_rca24_fa59_y2;
  wire h_s_wallace_rca24_fa59_y4;
  wire h_s_wallace_rca24_and_20_2_y0;
  wire h_s_wallace_rca24_and_19_3_y0;
  wire h_s_wallace_rca24_fa60_y2;
  wire h_s_wallace_rca24_fa60_y4;
  wire h_s_wallace_rca24_and_21_2_y0;
  wire h_s_wallace_rca24_and_20_3_y0;
  wire h_s_wallace_rca24_fa61_y2;
  wire h_s_wallace_rca24_fa61_y4;
  wire h_s_wallace_rca24_and_22_2_y0;
  wire h_s_wallace_rca24_and_21_3_y0;
  wire h_s_wallace_rca24_fa62_y2;
  wire h_s_wallace_rca24_fa62_y4;
  wire h_s_wallace_rca24_and_21_4_y0;
  wire h_s_wallace_rca24_and_20_5_y0;
  wire h_s_wallace_rca24_fa63_y2;
  wire h_s_wallace_rca24_fa63_y4;
  wire h_s_wallace_rca24_and_21_5_y0;
  wire h_s_wallace_rca24_and_20_6_y0;
  wire h_s_wallace_rca24_fa64_y2;
  wire h_s_wallace_rca24_fa64_y4;
  wire h_s_wallace_rca24_and_21_6_y0;
  wire h_s_wallace_rca24_and_20_7_y0;
  wire h_s_wallace_rca24_fa65_y2;
  wire h_s_wallace_rca24_fa65_y4;
  wire h_s_wallace_rca24_and_21_7_y0;
  wire h_s_wallace_rca24_and_20_8_y0;
  wire h_s_wallace_rca24_fa66_y2;
  wire h_s_wallace_rca24_fa66_y4;
  wire h_s_wallace_rca24_and_21_8_y0;
  wire h_s_wallace_rca24_and_20_9_y0;
  wire h_s_wallace_rca24_fa67_y2;
  wire h_s_wallace_rca24_fa67_y4;
  wire h_s_wallace_rca24_and_21_9_y0;
  wire h_s_wallace_rca24_and_20_10_y0;
  wire h_s_wallace_rca24_fa68_y2;
  wire h_s_wallace_rca24_fa68_y4;
  wire h_s_wallace_rca24_and_21_10_y0;
  wire h_s_wallace_rca24_and_20_11_y0;
  wire h_s_wallace_rca24_fa69_y2;
  wire h_s_wallace_rca24_fa69_y4;
  wire h_s_wallace_rca24_and_21_11_y0;
  wire h_s_wallace_rca24_and_20_12_y0;
  wire h_s_wallace_rca24_fa70_y2;
  wire h_s_wallace_rca24_fa70_y4;
  wire h_s_wallace_rca24_and_21_12_y0;
  wire h_s_wallace_rca24_and_20_13_y0;
  wire h_s_wallace_rca24_fa71_y2;
  wire h_s_wallace_rca24_fa71_y4;
  wire h_s_wallace_rca24_and_21_13_y0;
  wire h_s_wallace_rca24_and_20_14_y0;
  wire h_s_wallace_rca24_fa72_y2;
  wire h_s_wallace_rca24_fa72_y4;
  wire h_s_wallace_rca24_and_21_14_y0;
  wire h_s_wallace_rca24_and_20_15_y0;
  wire h_s_wallace_rca24_fa73_y2;
  wire h_s_wallace_rca24_fa73_y4;
  wire h_s_wallace_rca24_and_21_15_y0;
  wire h_s_wallace_rca24_and_20_16_y0;
  wire h_s_wallace_rca24_fa74_y2;
  wire h_s_wallace_rca24_fa74_y4;
  wire h_s_wallace_rca24_and_21_16_y0;
  wire h_s_wallace_rca24_and_20_17_y0;
  wire h_s_wallace_rca24_fa75_y2;
  wire h_s_wallace_rca24_fa75_y4;
  wire h_s_wallace_rca24_and_21_17_y0;
  wire h_s_wallace_rca24_and_20_18_y0;
  wire h_s_wallace_rca24_fa76_y2;
  wire h_s_wallace_rca24_fa76_y4;
  wire h_s_wallace_rca24_and_21_18_y0;
  wire h_s_wallace_rca24_and_20_19_y0;
  wire h_s_wallace_rca24_fa77_y2;
  wire h_s_wallace_rca24_fa77_y4;
  wire h_s_wallace_rca24_and_21_19_y0;
  wire h_s_wallace_rca24_and_20_20_y0;
  wire h_s_wallace_rca24_fa78_y2;
  wire h_s_wallace_rca24_fa78_y4;
  wire h_s_wallace_rca24_and_21_20_y0;
  wire h_s_wallace_rca24_and_20_21_y0;
  wire h_s_wallace_rca24_fa79_y2;
  wire h_s_wallace_rca24_fa79_y4;
  wire h_s_wallace_rca24_and_21_21_y0;
  wire h_s_wallace_rca24_and_20_22_y0;
  wire h_s_wallace_rca24_fa80_y2;
  wire h_s_wallace_rca24_fa80_y4;
  wire h_s_wallace_rca24_and_21_22_y0;
  wire h_s_wallace_rca24_nand_20_23_y0;
  wire h_s_wallace_rca24_fa81_y2;
  wire h_s_wallace_rca24_fa81_y4;
  wire h_s_wallace_rca24_and_0_4_y0;
  wire h_s_wallace_rca24_ha2_y0;
  wire h_s_wallace_rca24_ha2_y1;
  wire h_s_wallace_rca24_and_1_4_y0;
  wire h_s_wallace_rca24_and_0_5_y0;
  wire h_s_wallace_rca24_fa82_y2;
  wire h_s_wallace_rca24_fa82_y4;
  wire h_s_wallace_rca24_and_2_4_y0;
  wire h_s_wallace_rca24_and_1_5_y0;
  wire h_s_wallace_rca24_fa83_y2;
  wire h_s_wallace_rca24_fa83_y4;
  wire h_s_wallace_rca24_and_3_4_y0;
  wire h_s_wallace_rca24_and_2_5_y0;
  wire h_s_wallace_rca24_fa84_y2;
  wire h_s_wallace_rca24_fa84_y4;
  wire h_s_wallace_rca24_and_4_4_y0;
  wire h_s_wallace_rca24_and_3_5_y0;
  wire h_s_wallace_rca24_fa85_y2;
  wire h_s_wallace_rca24_fa85_y4;
  wire h_s_wallace_rca24_and_5_4_y0;
  wire h_s_wallace_rca24_and_4_5_y0;
  wire h_s_wallace_rca24_fa86_y2;
  wire h_s_wallace_rca24_fa86_y4;
  wire h_s_wallace_rca24_and_6_4_y0;
  wire h_s_wallace_rca24_and_5_5_y0;
  wire h_s_wallace_rca24_fa87_y2;
  wire h_s_wallace_rca24_fa87_y4;
  wire h_s_wallace_rca24_and_7_4_y0;
  wire h_s_wallace_rca24_and_6_5_y0;
  wire h_s_wallace_rca24_fa88_y2;
  wire h_s_wallace_rca24_fa88_y4;
  wire h_s_wallace_rca24_and_8_4_y0;
  wire h_s_wallace_rca24_and_7_5_y0;
  wire h_s_wallace_rca24_fa89_y2;
  wire h_s_wallace_rca24_fa89_y4;
  wire h_s_wallace_rca24_and_9_4_y0;
  wire h_s_wallace_rca24_and_8_5_y0;
  wire h_s_wallace_rca24_fa90_y2;
  wire h_s_wallace_rca24_fa90_y4;
  wire h_s_wallace_rca24_and_10_4_y0;
  wire h_s_wallace_rca24_and_9_5_y0;
  wire h_s_wallace_rca24_fa91_y2;
  wire h_s_wallace_rca24_fa91_y4;
  wire h_s_wallace_rca24_and_11_4_y0;
  wire h_s_wallace_rca24_and_10_5_y0;
  wire h_s_wallace_rca24_fa92_y2;
  wire h_s_wallace_rca24_fa92_y4;
  wire h_s_wallace_rca24_and_12_4_y0;
  wire h_s_wallace_rca24_and_11_5_y0;
  wire h_s_wallace_rca24_fa93_y2;
  wire h_s_wallace_rca24_fa93_y4;
  wire h_s_wallace_rca24_and_13_4_y0;
  wire h_s_wallace_rca24_and_12_5_y0;
  wire h_s_wallace_rca24_fa94_y2;
  wire h_s_wallace_rca24_fa94_y4;
  wire h_s_wallace_rca24_and_14_4_y0;
  wire h_s_wallace_rca24_and_13_5_y0;
  wire h_s_wallace_rca24_fa95_y2;
  wire h_s_wallace_rca24_fa95_y4;
  wire h_s_wallace_rca24_and_15_4_y0;
  wire h_s_wallace_rca24_and_14_5_y0;
  wire h_s_wallace_rca24_fa96_y2;
  wire h_s_wallace_rca24_fa96_y4;
  wire h_s_wallace_rca24_and_16_4_y0;
  wire h_s_wallace_rca24_and_15_5_y0;
  wire h_s_wallace_rca24_fa97_y2;
  wire h_s_wallace_rca24_fa97_y4;
  wire h_s_wallace_rca24_and_17_4_y0;
  wire h_s_wallace_rca24_and_16_5_y0;
  wire h_s_wallace_rca24_fa98_y2;
  wire h_s_wallace_rca24_fa98_y4;
  wire h_s_wallace_rca24_and_18_4_y0;
  wire h_s_wallace_rca24_and_17_5_y0;
  wire h_s_wallace_rca24_fa99_y2;
  wire h_s_wallace_rca24_fa99_y4;
  wire h_s_wallace_rca24_and_19_4_y0;
  wire h_s_wallace_rca24_and_18_5_y0;
  wire h_s_wallace_rca24_fa100_y2;
  wire h_s_wallace_rca24_fa100_y4;
  wire h_s_wallace_rca24_and_20_4_y0;
  wire h_s_wallace_rca24_and_19_5_y0;
  wire h_s_wallace_rca24_fa101_y2;
  wire h_s_wallace_rca24_fa101_y4;
  wire h_s_wallace_rca24_and_19_6_y0;
  wire h_s_wallace_rca24_and_18_7_y0;
  wire h_s_wallace_rca24_fa102_y2;
  wire h_s_wallace_rca24_fa102_y4;
  wire h_s_wallace_rca24_and_19_7_y0;
  wire h_s_wallace_rca24_and_18_8_y0;
  wire h_s_wallace_rca24_fa103_y2;
  wire h_s_wallace_rca24_fa103_y4;
  wire h_s_wallace_rca24_and_19_8_y0;
  wire h_s_wallace_rca24_and_18_9_y0;
  wire h_s_wallace_rca24_fa104_y2;
  wire h_s_wallace_rca24_fa104_y4;
  wire h_s_wallace_rca24_and_19_9_y0;
  wire h_s_wallace_rca24_and_18_10_y0;
  wire h_s_wallace_rca24_fa105_y2;
  wire h_s_wallace_rca24_fa105_y4;
  wire h_s_wallace_rca24_and_19_10_y0;
  wire h_s_wallace_rca24_and_18_11_y0;
  wire h_s_wallace_rca24_fa106_y2;
  wire h_s_wallace_rca24_fa106_y4;
  wire h_s_wallace_rca24_and_19_11_y0;
  wire h_s_wallace_rca24_and_18_12_y0;
  wire h_s_wallace_rca24_fa107_y2;
  wire h_s_wallace_rca24_fa107_y4;
  wire h_s_wallace_rca24_and_19_12_y0;
  wire h_s_wallace_rca24_and_18_13_y0;
  wire h_s_wallace_rca24_fa108_y2;
  wire h_s_wallace_rca24_fa108_y4;
  wire h_s_wallace_rca24_and_19_13_y0;
  wire h_s_wallace_rca24_and_18_14_y0;
  wire h_s_wallace_rca24_fa109_y2;
  wire h_s_wallace_rca24_fa109_y4;
  wire h_s_wallace_rca24_and_19_14_y0;
  wire h_s_wallace_rca24_and_18_15_y0;
  wire h_s_wallace_rca24_fa110_y2;
  wire h_s_wallace_rca24_fa110_y4;
  wire h_s_wallace_rca24_and_19_15_y0;
  wire h_s_wallace_rca24_and_18_16_y0;
  wire h_s_wallace_rca24_fa111_y2;
  wire h_s_wallace_rca24_fa111_y4;
  wire h_s_wallace_rca24_and_19_16_y0;
  wire h_s_wallace_rca24_and_18_17_y0;
  wire h_s_wallace_rca24_fa112_y2;
  wire h_s_wallace_rca24_fa112_y4;
  wire h_s_wallace_rca24_and_19_17_y0;
  wire h_s_wallace_rca24_and_18_18_y0;
  wire h_s_wallace_rca24_fa113_y2;
  wire h_s_wallace_rca24_fa113_y4;
  wire h_s_wallace_rca24_and_19_18_y0;
  wire h_s_wallace_rca24_and_18_19_y0;
  wire h_s_wallace_rca24_fa114_y2;
  wire h_s_wallace_rca24_fa114_y4;
  wire h_s_wallace_rca24_and_19_19_y0;
  wire h_s_wallace_rca24_and_18_20_y0;
  wire h_s_wallace_rca24_fa115_y2;
  wire h_s_wallace_rca24_fa115_y4;
  wire h_s_wallace_rca24_and_19_20_y0;
  wire h_s_wallace_rca24_and_18_21_y0;
  wire h_s_wallace_rca24_fa116_y2;
  wire h_s_wallace_rca24_fa116_y4;
  wire h_s_wallace_rca24_and_19_21_y0;
  wire h_s_wallace_rca24_and_18_22_y0;
  wire h_s_wallace_rca24_fa117_y2;
  wire h_s_wallace_rca24_fa117_y4;
  wire h_s_wallace_rca24_and_19_22_y0;
  wire h_s_wallace_rca24_nand_18_23_y0;
  wire h_s_wallace_rca24_fa118_y2;
  wire h_s_wallace_rca24_fa118_y4;
  wire h_s_wallace_rca24_nand_19_23_y0;
  wire h_s_wallace_rca24_fa119_y2;
  wire h_s_wallace_rca24_fa119_y4;
  wire h_s_wallace_rca24_ha3_y0;
  wire h_s_wallace_rca24_ha3_y1;
  wire h_s_wallace_rca24_and_0_6_y0;
  wire h_s_wallace_rca24_fa120_y2;
  wire h_s_wallace_rca24_fa120_y4;
  wire h_s_wallace_rca24_and_1_6_y0;
  wire h_s_wallace_rca24_and_0_7_y0;
  wire h_s_wallace_rca24_fa121_y2;
  wire h_s_wallace_rca24_fa121_y4;
  wire h_s_wallace_rca24_and_2_6_y0;
  wire h_s_wallace_rca24_and_1_7_y0;
  wire h_s_wallace_rca24_fa122_y2;
  wire h_s_wallace_rca24_fa122_y4;
  wire h_s_wallace_rca24_and_3_6_y0;
  wire h_s_wallace_rca24_and_2_7_y0;
  wire h_s_wallace_rca24_fa123_y2;
  wire h_s_wallace_rca24_fa123_y4;
  wire h_s_wallace_rca24_and_4_6_y0;
  wire h_s_wallace_rca24_and_3_7_y0;
  wire h_s_wallace_rca24_fa124_y2;
  wire h_s_wallace_rca24_fa124_y4;
  wire h_s_wallace_rca24_and_5_6_y0;
  wire h_s_wallace_rca24_and_4_7_y0;
  wire h_s_wallace_rca24_fa125_y2;
  wire h_s_wallace_rca24_fa125_y4;
  wire h_s_wallace_rca24_and_6_6_y0;
  wire h_s_wallace_rca24_and_5_7_y0;
  wire h_s_wallace_rca24_fa126_y2;
  wire h_s_wallace_rca24_fa126_y4;
  wire h_s_wallace_rca24_and_7_6_y0;
  wire h_s_wallace_rca24_and_6_7_y0;
  wire h_s_wallace_rca24_fa127_y2;
  wire h_s_wallace_rca24_fa127_y4;
  wire h_s_wallace_rca24_and_8_6_y0;
  wire h_s_wallace_rca24_and_7_7_y0;
  wire h_s_wallace_rca24_fa128_y2;
  wire h_s_wallace_rca24_fa128_y4;
  wire h_s_wallace_rca24_and_9_6_y0;
  wire h_s_wallace_rca24_and_8_7_y0;
  wire h_s_wallace_rca24_fa129_y2;
  wire h_s_wallace_rca24_fa129_y4;
  wire h_s_wallace_rca24_and_10_6_y0;
  wire h_s_wallace_rca24_and_9_7_y0;
  wire h_s_wallace_rca24_fa130_y2;
  wire h_s_wallace_rca24_fa130_y4;
  wire h_s_wallace_rca24_and_11_6_y0;
  wire h_s_wallace_rca24_and_10_7_y0;
  wire h_s_wallace_rca24_fa131_y2;
  wire h_s_wallace_rca24_fa131_y4;
  wire h_s_wallace_rca24_and_12_6_y0;
  wire h_s_wallace_rca24_and_11_7_y0;
  wire h_s_wallace_rca24_fa132_y2;
  wire h_s_wallace_rca24_fa132_y4;
  wire h_s_wallace_rca24_and_13_6_y0;
  wire h_s_wallace_rca24_and_12_7_y0;
  wire h_s_wallace_rca24_fa133_y2;
  wire h_s_wallace_rca24_fa133_y4;
  wire h_s_wallace_rca24_and_14_6_y0;
  wire h_s_wallace_rca24_and_13_7_y0;
  wire h_s_wallace_rca24_fa134_y2;
  wire h_s_wallace_rca24_fa134_y4;
  wire h_s_wallace_rca24_and_15_6_y0;
  wire h_s_wallace_rca24_and_14_7_y0;
  wire h_s_wallace_rca24_fa135_y2;
  wire h_s_wallace_rca24_fa135_y4;
  wire h_s_wallace_rca24_and_16_6_y0;
  wire h_s_wallace_rca24_and_15_7_y0;
  wire h_s_wallace_rca24_fa136_y2;
  wire h_s_wallace_rca24_fa136_y4;
  wire h_s_wallace_rca24_and_17_6_y0;
  wire h_s_wallace_rca24_and_16_7_y0;
  wire h_s_wallace_rca24_fa137_y2;
  wire h_s_wallace_rca24_fa137_y4;
  wire h_s_wallace_rca24_and_18_6_y0;
  wire h_s_wallace_rca24_and_17_7_y0;
  wire h_s_wallace_rca24_fa138_y2;
  wire h_s_wallace_rca24_fa138_y4;
  wire h_s_wallace_rca24_and_17_8_y0;
  wire h_s_wallace_rca24_and_16_9_y0;
  wire h_s_wallace_rca24_fa139_y2;
  wire h_s_wallace_rca24_fa139_y4;
  wire h_s_wallace_rca24_and_17_9_y0;
  wire h_s_wallace_rca24_and_16_10_y0;
  wire h_s_wallace_rca24_fa140_y2;
  wire h_s_wallace_rca24_fa140_y4;
  wire h_s_wallace_rca24_and_17_10_y0;
  wire h_s_wallace_rca24_and_16_11_y0;
  wire h_s_wallace_rca24_fa141_y2;
  wire h_s_wallace_rca24_fa141_y4;
  wire h_s_wallace_rca24_and_17_11_y0;
  wire h_s_wallace_rca24_and_16_12_y0;
  wire h_s_wallace_rca24_fa142_y2;
  wire h_s_wallace_rca24_fa142_y4;
  wire h_s_wallace_rca24_and_17_12_y0;
  wire h_s_wallace_rca24_and_16_13_y0;
  wire h_s_wallace_rca24_fa143_y2;
  wire h_s_wallace_rca24_fa143_y4;
  wire h_s_wallace_rca24_and_17_13_y0;
  wire h_s_wallace_rca24_and_16_14_y0;
  wire h_s_wallace_rca24_fa144_y2;
  wire h_s_wallace_rca24_fa144_y4;
  wire h_s_wallace_rca24_and_17_14_y0;
  wire h_s_wallace_rca24_and_16_15_y0;
  wire h_s_wallace_rca24_fa145_y2;
  wire h_s_wallace_rca24_fa145_y4;
  wire h_s_wallace_rca24_and_17_15_y0;
  wire h_s_wallace_rca24_and_16_16_y0;
  wire h_s_wallace_rca24_fa146_y2;
  wire h_s_wallace_rca24_fa146_y4;
  wire h_s_wallace_rca24_and_17_16_y0;
  wire h_s_wallace_rca24_and_16_17_y0;
  wire h_s_wallace_rca24_fa147_y2;
  wire h_s_wallace_rca24_fa147_y4;
  wire h_s_wallace_rca24_and_17_17_y0;
  wire h_s_wallace_rca24_and_16_18_y0;
  wire h_s_wallace_rca24_fa148_y2;
  wire h_s_wallace_rca24_fa148_y4;
  wire h_s_wallace_rca24_and_17_18_y0;
  wire h_s_wallace_rca24_and_16_19_y0;
  wire h_s_wallace_rca24_fa149_y2;
  wire h_s_wallace_rca24_fa149_y4;
  wire h_s_wallace_rca24_and_17_19_y0;
  wire h_s_wallace_rca24_and_16_20_y0;
  wire h_s_wallace_rca24_fa150_y2;
  wire h_s_wallace_rca24_fa150_y4;
  wire h_s_wallace_rca24_and_17_20_y0;
  wire h_s_wallace_rca24_and_16_21_y0;
  wire h_s_wallace_rca24_fa151_y2;
  wire h_s_wallace_rca24_fa151_y4;
  wire h_s_wallace_rca24_and_17_21_y0;
  wire h_s_wallace_rca24_and_16_22_y0;
  wire h_s_wallace_rca24_fa152_y2;
  wire h_s_wallace_rca24_fa152_y4;
  wire h_s_wallace_rca24_and_17_22_y0;
  wire h_s_wallace_rca24_nand_16_23_y0;
  wire h_s_wallace_rca24_fa153_y2;
  wire h_s_wallace_rca24_fa153_y4;
  wire h_s_wallace_rca24_nand_17_23_y0;
  wire h_s_wallace_rca24_fa154_y2;
  wire h_s_wallace_rca24_fa154_y4;
  wire h_s_wallace_rca24_fa155_y2;
  wire h_s_wallace_rca24_fa155_y4;
  wire h_s_wallace_rca24_ha4_y0;
  wire h_s_wallace_rca24_ha4_y1;
  wire h_s_wallace_rca24_fa156_y2;
  wire h_s_wallace_rca24_fa156_y4;
  wire h_s_wallace_rca24_and_0_8_y0;
  wire h_s_wallace_rca24_fa157_y2;
  wire h_s_wallace_rca24_fa157_y4;
  wire h_s_wallace_rca24_and_1_8_y0;
  wire h_s_wallace_rca24_and_0_9_y0;
  wire h_s_wallace_rca24_fa158_y2;
  wire h_s_wallace_rca24_fa158_y4;
  wire h_s_wallace_rca24_and_2_8_y0;
  wire h_s_wallace_rca24_and_1_9_y0;
  wire h_s_wallace_rca24_fa159_y2;
  wire h_s_wallace_rca24_fa159_y4;
  wire h_s_wallace_rca24_and_3_8_y0;
  wire h_s_wallace_rca24_and_2_9_y0;
  wire h_s_wallace_rca24_fa160_y2;
  wire h_s_wallace_rca24_fa160_y4;
  wire h_s_wallace_rca24_and_4_8_y0;
  wire h_s_wallace_rca24_and_3_9_y0;
  wire h_s_wallace_rca24_fa161_y2;
  wire h_s_wallace_rca24_fa161_y4;
  wire h_s_wallace_rca24_and_5_8_y0;
  wire h_s_wallace_rca24_and_4_9_y0;
  wire h_s_wallace_rca24_fa162_y2;
  wire h_s_wallace_rca24_fa162_y4;
  wire h_s_wallace_rca24_and_6_8_y0;
  wire h_s_wallace_rca24_and_5_9_y0;
  wire h_s_wallace_rca24_fa163_y2;
  wire h_s_wallace_rca24_fa163_y4;
  wire h_s_wallace_rca24_and_7_8_y0;
  wire h_s_wallace_rca24_and_6_9_y0;
  wire h_s_wallace_rca24_fa164_y2;
  wire h_s_wallace_rca24_fa164_y4;
  wire h_s_wallace_rca24_and_8_8_y0;
  wire h_s_wallace_rca24_and_7_9_y0;
  wire h_s_wallace_rca24_fa165_y2;
  wire h_s_wallace_rca24_fa165_y4;
  wire h_s_wallace_rca24_and_9_8_y0;
  wire h_s_wallace_rca24_and_8_9_y0;
  wire h_s_wallace_rca24_fa166_y2;
  wire h_s_wallace_rca24_fa166_y4;
  wire h_s_wallace_rca24_and_10_8_y0;
  wire h_s_wallace_rca24_and_9_9_y0;
  wire h_s_wallace_rca24_fa167_y2;
  wire h_s_wallace_rca24_fa167_y4;
  wire h_s_wallace_rca24_and_11_8_y0;
  wire h_s_wallace_rca24_and_10_9_y0;
  wire h_s_wallace_rca24_fa168_y2;
  wire h_s_wallace_rca24_fa168_y4;
  wire h_s_wallace_rca24_and_12_8_y0;
  wire h_s_wallace_rca24_and_11_9_y0;
  wire h_s_wallace_rca24_fa169_y2;
  wire h_s_wallace_rca24_fa169_y4;
  wire h_s_wallace_rca24_and_13_8_y0;
  wire h_s_wallace_rca24_and_12_9_y0;
  wire h_s_wallace_rca24_fa170_y2;
  wire h_s_wallace_rca24_fa170_y4;
  wire h_s_wallace_rca24_and_14_8_y0;
  wire h_s_wallace_rca24_and_13_9_y0;
  wire h_s_wallace_rca24_fa171_y2;
  wire h_s_wallace_rca24_fa171_y4;
  wire h_s_wallace_rca24_and_15_8_y0;
  wire h_s_wallace_rca24_and_14_9_y0;
  wire h_s_wallace_rca24_fa172_y2;
  wire h_s_wallace_rca24_fa172_y4;
  wire h_s_wallace_rca24_and_16_8_y0;
  wire h_s_wallace_rca24_and_15_9_y0;
  wire h_s_wallace_rca24_fa173_y2;
  wire h_s_wallace_rca24_fa173_y4;
  wire h_s_wallace_rca24_and_15_10_y0;
  wire h_s_wallace_rca24_and_14_11_y0;
  wire h_s_wallace_rca24_fa174_y2;
  wire h_s_wallace_rca24_fa174_y4;
  wire h_s_wallace_rca24_and_15_11_y0;
  wire h_s_wallace_rca24_and_14_12_y0;
  wire h_s_wallace_rca24_fa175_y2;
  wire h_s_wallace_rca24_fa175_y4;
  wire h_s_wallace_rca24_and_15_12_y0;
  wire h_s_wallace_rca24_and_14_13_y0;
  wire h_s_wallace_rca24_fa176_y2;
  wire h_s_wallace_rca24_fa176_y4;
  wire h_s_wallace_rca24_and_15_13_y0;
  wire h_s_wallace_rca24_and_14_14_y0;
  wire h_s_wallace_rca24_fa177_y2;
  wire h_s_wallace_rca24_fa177_y4;
  wire h_s_wallace_rca24_and_15_14_y0;
  wire h_s_wallace_rca24_and_14_15_y0;
  wire h_s_wallace_rca24_fa178_y2;
  wire h_s_wallace_rca24_fa178_y4;
  wire h_s_wallace_rca24_and_15_15_y0;
  wire h_s_wallace_rca24_and_14_16_y0;
  wire h_s_wallace_rca24_fa179_y2;
  wire h_s_wallace_rca24_fa179_y4;
  wire h_s_wallace_rca24_and_15_16_y0;
  wire h_s_wallace_rca24_and_14_17_y0;
  wire h_s_wallace_rca24_fa180_y2;
  wire h_s_wallace_rca24_fa180_y4;
  wire h_s_wallace_rca24_and_15_17_y0;
  wire h_s_wallace_rca24_and_14_18_y0;
  wire h_s_wallace_rca24_fa181_y2;
  wire h_s_wallace_rca24_fa181_y4;
  wire h_s_wallace_rca24_and_15_18_y0;
  wire h_s_wallace_rca24_and_14_19_y0;
  wire h_s_wallace_rca24_fa182_y2;
  wire h_s_wallace_rca24_fa182_y4;
  wire h_s_wallace_rca24_and_15_19_y0;
  wire h_s_wallace_rca24_and_14_20_y0;
  wire h_s_wallace_rca24_fa183_y2;
  wire h_s_wallace_rca24_fa183_y4;
  wire h_s_wallace_rca24_and_15_20_y0;
  wire h_s_wallace_rca24_and_14_21_y0;
  wire h_s_wallace_rca24_fa184_y2;
  wire h_s_wallace_rca24_fa184_y4;
  wire h_s_wallace_rca24_and_15_21_y0;
  wire h_s_wallace_rca24_and_14_22_y0;
  wire h_s_wallace_rca24_fa185_y2;
  wire h_s_wallace_rca24_fa185_y4;
  wire h_s_wallace_rca24_and_15_22_y0;
  wire h_s_wallace_rca24_nand_14_23_y0;
  wire h_s_wallace_rca24_fa186_y2;
  wire h_s_wallace_rca24_fa186_y4;
  wire h_s_wallace_rca24_nand_15_23_y0;
  wire h_s_wallace_rca24_fa187_y2;
  wire h_s_wallace_rca24_fa187_y4;
  wire h_s_wallace_rca24_fa188_y2;
  wire h_s_wallace_rca24_fa188_y4;
  wire h_s_wallace_rca24_fa189_y2;
  wire h_s_wallace_rca24_fa189_y4;
  wire h_s_wallace_rca24_ha5_y0;
  wire h_s_wallace_rca24_ha5_y1;
  wire h_s_wallace_rca24_fa190_y2;
  wire h_s_wallace_rca24_fa190_y4;
  wire h_s_wallace_rca24_fa191_y2;
  wire h_s_wallace_rca24_fa191_y4;
  wire h_s_wallace_rca24_and_0_10_y0;
  wire h_s_wallace_rca24_fa192_y2;
  wire h_s_wallace_rca24_fa192_y4;
  wire h_s_wallace_rca24_and_1_10_y0;
  wire h_s_wallace_rca24_and_0_11_y0;
  wire h_s_wallace_rca24_fa193_y2;
  wire h_s_wallace_rca24_fa193_y4;
  wire h_s_wallace_rca24_and_2_10_y0;
  wire h_s_wallace_rca24_and_1_11_y0;
  wire h_s_wallace_rca24_fa194_y2;
  wire h_s_wallace_rca24_fa194_y4;
  wire h_s_wallace_rca24_and_3_10_y0;
  wire h_s_wallace_rca24_and_2_11_y0;
  wire h_s_wallace_rca24_fa195_y2;
  wire h_s_wallace_rca24_fa195_y4;
  wire h_s_wallace_rca24_and_4_10_y0;
  wire h_s_wallace_rca24_and_3_11_y0;
  wire h_s_wallace_rca24_fa196_y2;
  wire h_s_wallace_rca24_fa196_y4;
  wire h_s_wallace_rca24_and_5_10_y0;
  wire h_s_wallace_rca24_and_4_11_y0;
  wire h_s_wallace_rca24_fa197_y2;
  wire h_s_wallace_rca24_fa197_y4;
  wire h_s_wallace_rca24_and_6_10_y0;
  wire h_s_wallace_rca24_and_5_11_y0;
  wire h_s_wallace_rca24_fa198_y2;
  wire h_s_wallace_rca24_fa198_y4;
  wire h_s_wallace_rca24_and_7_10_y0;
  wire h_s_wallace_rca24_and_6_11_y0;
  wire h_s_wallace_rca24_fa199_y2;
  wire h_s_wallace_rca24_fa199_y4;
  wire h_s_wallace_rca24_and_8_10_y0;
  wire h_s_wallace_rca24_and_7_11_y0;
  wire h_s_wallace_rca24_fa200_y2;
  wire h_s_wallace_rca24_fa200_y4;
  wire h_s_wallace_rca24_and_9_10_y0;
  wire h_s_wallace_rca24_and_8_11_y0;
  wire h_s_wallace_rca24_fa201_y2;
  wire h_s_wallace_rca24_fa201_y4;
  wire h_s_wallace_rca24_and_10_10_y0;
  wire h_s_wallace_rca24_and_9_11_y0;
  wire h_s_wallace_rca24_fa202_y2;
  wire h_s_wallace_rca24_fa202_y4;
  wire h_s_wallace_rca24_and_11_10_y0;
  wire h_s_wallace_rca24_and_10_11_y0;
  wire h_s_wallace_rca24_fa203_y2;
  wire h_s_wallace_rca24_fa203_y4;
  wire h_s_wallace_rca24_and_12_10_y0;
  wire h_s_wallace_rca24_and_11_11_y0;
  wire h_s_wallace_rca24_fa204_y2;
  wire h_s_wallace_rca24_fa204_y4;
  wire h_s_wallace_rca24_and_13_10_y0;
  wire h_s_wallace_rca24_and_12_11_y0;
  wire h_s_wallace_rca24_fa205_y2;
  wire h_s_wallace_rca24_fa205_y4;
  wire h_s_wallace_rca24_and_14_10_y0;
  wire h_s_wallace_rca24_and_13_11_y0;
  wire h_s_wallace_rca24_fa206_y2;
  wire h_s_wallace_rca24_fa206_y4;
  wire h_s_wallace_rca24_and_13_12_y0;
  wire h_s_wallace_rca24_and_12_13_y0;
  wire h_s_wallace_rca24_fa207_y2;
  wire h_s_wallace_rca24_fa207_y4;
  wire h_s_wallace_rca24_and_13_13_y0;
  wire h_s_wallace_rca24_and_12_14_y0;
  wire h_s_wallace_rca24_fa208_y2;
  wire h_s_wallace_rca24_fa208_y4;
  wire h_s_wallace_rca24_and_13_14_y0;
  wire h_s_wallace_rca24_and_12_15_y0;
  wire h_s_wallace_rca24_fa209_y2;
  wire h_s_wallace_rca24_fa209_y4;
  wire h_s_wallace_rca24_and_13_15_y0;
  wire h_s_wallace_rca24_and_12_16_y0;
  wire h_s_wallace_rca24_fa210_y2;
  wire h_s_wallace_rca24_fa210_y4;
  wire h_s_wallace_rca24_and_13_16_y0;
  wire h_s_wallace_rca24_and_12_17_y0;
  wire h_s_wallace_rca24_fa211_y2;
  wire h_s_wallace_rca24_fa211_y4;
  wire h_s_wallace_rca24_and_13_17_y0;
  wire h_s_wallace_rca24_and_12_18_y0;
  wire h_s_wallace_rca24_fa212_y2;
  wire h_s_wallace_rca24_fa212_y4;
  wire h_s_wallace_rca24_and_13_18_y0;
  wire h_s_wallace_rca24_and_12_19_y0;
  wire h_s_wallace_rca24_fa213_y2;
  wire h_s_wallace_rca24_fa213_y4;
  wire h_s_wallace_rca24_and_13_19_y0;
  wire h_s_wallace_rca24_and_12_20_y0;
  wire h_s_wallace_rca24_fa214_y2;
  wire h_s_wallace_rca24_fa214_y4;
  wire h_s_wallace_rca24_and_13_20_y0;
  wire h_s_wallace_rca24_and_12_21_y0;
  wire h_s_wallace_rca24_fa215_y2;
  wire h_s_wallace_rca24_fa215_y4;
  wire h_s_wallace_rca24_and_13_21_y0;
  wire h_s_wallace_rca24_and_12_22_y0;
  wire h_s_wallace_rca24_fa216_y2;
  wire h_s_wallace_rca24_fa216_y4;
  wire h_s_wallace_rca24_and_13_22_y0;
  wire h_s_wallace_rca24_nand_12_23_y0;
  wire h_s_wallace_rca24_fa217_y2;
  wire h_s_wallace_rca24_fa217_y4;
  wire h_s_wallace_rca24_nand_13_23_y0;
  wire h_s_wallace_rca24_fa218_y2;
  wire h_s_wallace_rca24_fa218_y4;
  wire h_s_wallace_rca24_fa219_y2;
  wire h_s_wallace_rca24_fa219_y4;
  wire h_s_wallace_rca24_fa220_y2;
  wire h_s_wallace_rca24_fa220_y4;
  wire h_s_wallace_rca24_fa221_y2;
  wire h_s_wallace_rca24_fa221_y4;
  wire h_s_wallace_rca24_ha6_y0;
  wire h_s_wallace_rca24_ha6_y1;
  wire h_s_wallace_rca24_fa222_y2;
  wire h_s_wallace_rca24_fa222_y4;
  wire h_s_wallace_rca24_fa223_y2;
  wire h_s_wallace_rca24_fa223_y4;
  wire h_s_wallace_rca24_fa224_y2;
  wire h_s_wallace_rca24_fa224_y4;
  wire h_s_wallace_rca24_and_0_12_y0;
  wire h_s_wallace_rca24_fa225_y2;
  wire h_s_wallace_rca24_fa225_y4;
  wire h_s_wallace_rca24_and_1_12_y0;
  wire h_s_wallace_rca24_and_0_13_y0;
  wire h_s_wallace_rca24_fa226_y2;
  wire h_s_wallace_rca24_fa226_y4;
  wire h_s_wallace_rca24_and_2_12_y0;
  wire h_s_wallace_rca24_and_1_13_y0;
  wire h_s_wallace_rca24_fa227_y2;
  wire h_s_wallace_rca24_fa227_y4;
  wire h_s_wallace_rca24_and_3_12_y0;
  wire h_s_wallace_rca24_and_2_13_y0;
  wire h_s_wallace_rca24_fa228_y2;
  wire h_s_wallace_rca24_fa228_y4;
  wire h_s_wallace_rca24_and_4_12_y0;
  wire h_s_wallace_rca24_and_3_13_y0;
  wire h_s_wallace_rca24_fa229_y2;
  wire h_s_wallace_rca24_fa229_y4;
  wire h_s_wallace_rca24_and_5_12_y0;
  wire h_s_wallace_rca24_and_4_13_y0;
  wire h_s_wallace_rca24_fa230_y2;
  wire h_s_wallace_rca24_fa230_y4;
  wire h_s_wallace_rca24_and_6_12_y0;
  wire h_s_wallace_rca24_and_5_13_y0;
  wire h_s_wallace_rca24_fa231_y2;
  wire h_s_wallace_rca24_fa231_y4;
  wire h_s_wallace_rca24_and_7_12_y0;
  wire h_s_wallace_rca24_and_6_13_y0;
  wire h_s_wallace_rca24_fa232_y2;
  wire h_s_wallace_rca24_fa232_y4;
  wire h_s_wallace_rca24_and_8_12_y0;
  wire h_s_wallace_rca24_and_7_13_y0;
  wire h_s_wallace_rca24_fa233_y2;
  wire h_s_wallace_rca24_fa233_y4;
  wire h_s_wallace_rca24_and_9_12_y0;
  wire h_s_wallace_rca24_and_8_13_y0;
  wire h_s_wallace_rca24_fa234_y2;
  wire h_s_wallace_rca24_fa234_y4;
  wire h_s_wallace_rca24_and_10_12_y0;
  wire h_s_wallace_rca24_and_9_13_y0;
  wire h_s_wallace_rca24_fa235_y2;
  wire h_s_wallace_rca24_fa235_y4;
  wire h_s_wallace_rca24_and_11_12_y0;
  wire h_s_wallace_rca24_and_10_13_y0;
  wire h_s_wallace_rca24_fa236_y2;
  wire h_s_wallace_rca24_fa236_y4;
  wire h_s_wallace_rca24_and_12_12_y0;
  wire h_s_wallace_rca24_and_11_13_y0;
  wire h_s_wallace_rca24_fa237_y2;
  wire h_s_wallace_rca24_fa237_y4;
  wire h_s_wallace_rca24_and_11_14_y0;
  wire h_s_wallace_rca24_and_10_15_y0;
  wire h_s_wallace_rca24_fa238_y2;
  wire h_s_wallace_rca24_fa238_y4;
  wire h_s_wallace_rca24_and_11_15_y0;
  wire h_s_wallace_rca24_and_10_16_y0;
  wire h_s_wallace_rca24_fa239_y2;
  wire h_s_wallace_rca24_fa239_y4;
  wire h_s_wallace_rca24_and_11_16_y0;
  wire h_s_wallace_rca24_and_10_17_y0;
  wire h_s_wallace_rca24_fa240_y2;
  wire h_s_wallace_rca24_fa240_y4;
  wire h_s_wallace_rca24_and_11_17_y0;
  wire h_s_wallace_rca24_and_10_18_y0;
  wire h_s_wallace_rca24_fa241_y2;
  wire h_s_wallace_rca24_fa241_y4;
  wire h_s_wallace_rca24_and_11_18_y0;
  wire h_s_wallace_rca24_and_10_19_y0;
  wire h_s_wallace_rca24_fa242_y2;
  wire h_s_wallace_rca24_fa242_y4;
  wire h_s_wallace_rca24_and_11_19_y0;
  wire h_s_wallace_rca24_and_10_20_y0;
  wire h_s_wallace_rca24_fa243_y2;
  wire h_s_wallace_rca24_fa243_y4;
  wire h_s_wallace_rca24_and_11_20_y0;
  wire h_s_wallace_rca24_and_10_21_y0;
  wire h_s_wallace_rca24_fa244_y2;
  wire h_s_wallace_rca24_fa244_y4;
  wire h_s_wallace_rca24_and_11_21_y0;
  wire h_s_wallace_rca24_and_10_22_y0;
  wire h_s_wallace_rca24_fa245_y2;
  wire h_s_wallace_rca24_fa245_y4;
  wire h_s_wallace_rca24_and_11_22_y0;
  wire h_s_wallace_rca24_nand_10_23_y0;
  wire h_s_wallace_rca24_fa246_y2;
  wire h_s_wallace_rca24_fa246_y4;
  wire h_s_wallace_rca24_nand_11_23_y0;
  wire h_s_wallace_rca24_fa247_y2;
  wire h_s_wallace_rca24_fa247_y4;
  wire h_s_wallace_rca24_fa248_y2;
  wire h_s_wallace_rca24_fa248_y4;
  wire h_s_wallace_rca24_fa249_y2;
  wire h_s_wallace_rca24_fa249_y4;
  wire h_s_wallace_rca24_fa250_y2;
  wire h_s_wallace_rca24_fa250_y4;
  wire h_s_wallace_rca24_fa251_y2;
  wire h_s_wallace_rca24_fa251_y4;
  wire h_s_wallace_rca24_ha7_y0;
  wire h_s_wallace_rca24_ha7_y1;
  wire h_s_wallace_rca24_fa252_y2;
  wire h_s_wallace_rca24_fa252_y4;
  wire h_s_wallace_rca24_fa253_y2;
  wire h_s_wallace_rca24_fa253_y4;
  wire h_s_wallace_rca24_fa254_y2;
  wire h_s_wallace_rca24_fa254_y4;
  wire h_s_wallace_rca24_fa255_y2;
  wire h_s_wallace_rca24_fa255_y4;
  wire h_s_wallace_rca24_and_0_14_y0;
  wire h_s_wallace_rca24_fa256_y2;
  wire h_s_wallace_rca24_fa256_y4;
  wire h_s_wallace_rca24_and_1_14_y0;
  wire h_s_wallace_rca24_and_0_15_y0;
  wire h_s_wallace_rca24_fa257_y2;
  wire h_s_wallace_rca24_fa257_y4;
  wire h_s_wallace_rca24_and_2_14_y0;
  wire h_s_wallace_rca24_and_1_15_y0;
  wire h_s_wallace_rca24_fa258_y2;
  wire h_s_wallace_rca24_fa258_y4;
  wire h_s_wallace_rca24_and_3_14_y0;
  wire h_s_wallace_rca24_and_2_15_y0;
  wire h_s_wallace_rca24_fa259_y2;
  wire h_s_wallace_rca24_fa259_y4;
  wire h_s_wallace_rca24_and_4_14_y0;
  wire h_s_wallace_rca24_and_3_15_y0;
  wire h_s_wallace_rca24_fa260_y2;
  wire h_s_wallace_rca24_fa260_y4;
  wire h_s_wallace_rca24_and_5_14_y0;
  wire h_s_wallace_rca24_and_4_15_y0;
  wire h_s_wallace_rca24_fa261_y2;
  wire h_s_wallace_rca24_fa261_y4;
  wire h_s_wallace_rca24_and_6_14_y0;
  wire h_s_wallace_rca24_and_5_15_y0;
  wire h_s_wallace_rca24_fa262_y2;
  wire h_s_wallace_rca24_fa262_y4;
  wire h_s_wallace_rca24_and_7_14_y0;
  wire h_s_wallace_rca24_and_6_15_y0;
  wire h_s_wallace_rca24_fa263_y2;
  wire h_s_wallace_rca24_fa263_y4;
  wire h_s_wallace_rca24_and_8_14_y0;
  wire h_s_wallace_rca24_and_7_15_y0;
  wire h_s_wallace_rca24_fa264_y2;
  wire h_s_wallace_rca24_fa264_y4;
  wire h_s_wallace_rca24_and_9_14_y0;
  wire h_s_wallace_rca24_and_8_15_y0;
  wire h_s_wallace_rca24_fa265_y2;
  wire h_s_wallace_rca24_fa265_y4;
  wire h_s_wallace_rca24_and_10_14_y0;
  wire h_s_wallace_rca24_and_9_15_y0;
  wire h_s_wallace_rca24_fa266_y2;
  wire h_s_wallace_rca24_fa266_y4;
  wire h_s_wallace_rca24_and_9_16_y0;
  wire h_s_wallace_rca24_and_8_17_y0;
  wire h_s_wallace_rca24_fa267_y2;
  wire h_s_wallace_rca24_fa267_y4;
  wire h_s_wallace_rca24_and_9_17_y0;
  wire h_s_wallace_rca24_and_8_18_y0;
  wire h_s_wallace_rca24_fa268_y2;
  wire h_s_wallace_rca24_fa268_y4;
  wire h_s_wallace_rca24_and_9_18_y0;
  wire h_s_wallace_rca24_and_8_19_y0;
  wire h_s_wallace_rca24_fa269_y2;
  wire h_s_wallace_rca24_fa269_y4;
  wire h_s_wallace_rca24_and_9_19_y0;
  wire h_s_wallace_rca24_and_8_20_y0;
  wire h_s_wallace_rca24_fa270_y2;
  wire h_s_wallace_rca24_fa270_y4;
  wire h_s_wallace_rca24_and_9_20_y0;
  wire h_s_wallace_rca24_and_8_21_y0;
  wire h_s_wallace_rca24_fa271_y2;
  wire h_s_wallace_rca24_fa271_y4;
  wire h_s_wallace_rca24_and_9_21_y0;
  wire h_s_wallace_rca24_and_8_22_y0;
  wire h_s_wallace_rca24_fa272_y2;
  wire h_s_wallace_rca24_fa272_y4;
  wire h_s_wallace_rca24_and_9_22_y0;
  wire h_s_wallace_rca24_nand_8_23_y0;
  wire h_s_wallace_rca24_fa273_y2;
  wire h_s_wallace_rca24_fa273_y4;
  wire h_s_wallace_rca24_nand_9_23_y0;
  wire h_s_wallace_rca24_fa274_y2;
  wire h_s_wallace_rca24_fa274_y4;
  wire h_s_wallace_rca24_fa275_y2;
  wire h_s_wallace_rca24_fa275_y4;
  wire h_s_wallace_rca24_fa276_y2;
  wire h_s_wallace_rca24_fa276_y4;
  wire h_s_wallace_rca24_fa277_y2;
  wire h_s_wallace_rca24_fa277_y4;
  wire h_s_wallace_rca24_fa278_y2;
  wire h_s_wallace_rca24_fa278_y4;
  wire h_s_wallace_rca24_fa279_y2;
  wire h_s_wallace_rca24_fa279_y4;
  wire h_s_wallace_rca24_ha8_y0;
  wire h_s_wallace_rca24_ha8_y1;
  wire h_s_wallace_rca24_fa280_y2;
  wire h_s_wallace_rca24_fa280_y4;
  wire h_s_wallace_rca24_fa281_y2;
  wire h_s_wallace_rca24_fa281_y4;
  wire h_s_wallace_rca24_fa282_y2;
  wire h_s_wallace_rca24_fa282_y4;
  wire h_s_wallace_rca24_fa283_y2;
  wire h_s_wallace_rca24_fa283_y4;
  wire h_s_wallace_rca24_fa284_y2;
  wire h_s_wallace_rca24_fa284_y4;
  wire h_s_wallace_rca24_and_0_16_y0;
  wire h_s_wallace_rca24_fa285_y2;
  wire h_s_wallace_rca24_fa285_y4;
  wire h_s_wallace_rca24_and_1_16_y0;
  wire h_s_wallace_rca24_and_0_17_y0;
  wire h_s_wallace_rca24_fa286_y2;
  wire h_s_wallace_rca24_fa286_y4;
  wire h_s_wallace_rca24_and_2_16_y0;
  wire h_s_wallace_rca24_and_1_17_y0;
  wire h_s_wallace_rca24_fa287_y2;
  wire h_s_wallace_rca24_fa287_y4;
  wire h_s_wallace_rca24_and_3_16_y0;
  wire h_s_wallace_rca24_and_2_17_y0;
  wire h_s_wallace_rca24_fa288_y2;
  wire h_s_wallace_rca24_fa288_y4;
  wire h_s_wallace_rca24_and_4_16_y0;
  wire h_s_wallace_rca24_and_3_17_y0;
  wire h_s_wallace_rca24_fa289_y2;
  wire h_s_wallace_rca24_fa289_y4;
  wire h_s_wallace_rca24_and_5_16_y0;
  wire h_s_wallace_rca24_and_4_17_y0;
  wire h_s_wallace_rca24_fa290_y2;
  wire h_s_wallace_rca24_fa290_y4;
  wire h_s_wallace_rca24_and_6_16_y0;
  wire h_s_wallace_rca24_and_5_17_y0;
  wire h_s_wallace_rca24_fa291_y2;
  wire h_s_wallace_rca24_fa291_y4;
  wire h_s_wallace_rca24_and_7_16_y0;
  wire h_s_wallace_rca24_and_6_17_y0;
  wire h_s_wallace_rca24_fa292_y2;
  wire h_s_wallace_rca24_fa292_y4;
  wire h_s_wallace_rca24_and_8_16_y0;
  wire h_s_wallace_rca24_and_7_17_y0;
  wire h_s_wallace_rca24_fa293_y2;
  wire h_s_wallace_rca24_fa293_y4;
  wire h_s_wallace_rca24_and_7_18_y0;
  wire h_s_wallace_rca24_and_6_19_y0;
  wire h_s_wallace_rca24_fa294_y2;
  wire h_s_wallace_rca24_fa294_y4;
  wire h_s_wallace_rca24_and_7_19_y0;
  wire h_s_wallace_rca24_and_6_20_y0;
  wire h_s_wallace_rca24_fa295_y2;
  wire h_s_wallace_rca24_fa295_y4;
  wire h_s_wallace_rca24_and_7_20_y0;
  wire h_s_wallace_rca24_and_6_21_y0;
  wire h_s_wallace_rca24_fa296_y2;
  wire h_s_wallace_rca24_fa296_y4;
  wire h_s_wallace_rca24_and_7_21_y0;
  wire h_s_wallace_rca24_and_6_22_y0;
  wire h_s_wallace_rca24_fa297_y2;
  wire h_s_wallace_rca24_fa297_y4;
  wire h_s_wallace_rca24_and_7_22_y0;
  wire h_s_wallace_rca24_nand_6_23_y0;
  wire h_s_wallace_rca24_fa298_y2;
  wire h_s_wallace_rca24_fa298_y4;
  wire h_s_wallace_rca24_nand_7_23_y0;
  wire h_s_wallace_rca24_fa299_y2;
  wire h_s_wallace_rca24_fa299_y4;
  wire h_s_wallace_rca24_fa300_y2;
  wire h_s_wallace_rca24_fa300_y4;
  wire h_s_wallace_rca24_fa301_y2;
  wire h_s_wallace_rca24_fa301_y4;
  wire h_s_wallace_rca24_fa302_y2;
  wire h_s_wallace_rca24_fa302_y4;
  wire h_s_wallace_rca24_fa303_y2;
  wire h_s_wallace_rca24_fa303_y4;
  wire h_s_wallace_rca24_fa304_y2;
  wire h_s_wallace_rca24_fa304_y4;
  wire h_s_wallace_rca24_fa305_y2;
  wire h_s_wallace_rca24_fa305_y4;
  wire h_s_wallace_rca24_ha9_y0;
  wire h_s_wallace_rca24_ha9_y1;
  wire h_s_wallace_rca24_fa306_y2;
  wire h_s_wallace_rca24_fa306_y4;
  wire h_s_wallace_rca24_fa307_y2;
  wire h_s_wallace_rca24_fa307_y4;
  wire h_s_wallace_rca24_fa308_y2;
  wire h_s_wallace_rca24_fa308_y4;
  wire h_s_wallace_rca24_fa309_y2;
  wire h_s_wallace_rca24_fa309_y4;
  wire h_s_wallace_rca24_fa310_y2;
  wire h_s_wallace_rca24_fa310_y4;
  wire h_s_wallace_rca24_fa311_y2;
  wire h_s_wallace_rca24_fa311_y4;
  wire h_s_wallace_rca24_and_0_18_y0;
  wire h_s_wallace_rca24_fa312_y2;
  wire h_s_wallace_rca24_fa312_y4;
  wire h_s_wallace_rca24_and_1_18_y0;
  wire h_s_wallace_rca24_and_0_19_y0;
  wire h_s_wallace_rca24_fa313_y2;
  wire h_s_wallace_rca24_fa313_y4;
  wire h_s_wallace_rca24_and_2_18_y0;
  wire h_s_wallace_rca24_and_1_19_y0;
  wire h_s_wallace_rca24_fa314_y2;
  wire h_s_wallace_rca24_fa314_y4;
  wire h_s_wallace_rca24_and_3_18_y0;
  wire h_s_wallace_rca24_and_2_19_y0;
  wire h_s_wallace_rca24_fa315_y2;
  wire h_s_wallace_rca24_fa315_y4;
  wire h_s_wallace_rca24_and_4_18_y0;
  wire h_s_wallace_rca24_and_3_19_y0;
  wire h_s_wallace_rca24_fa316_y2;
  wire h_s_wallace_rca24_fa316_y4;
  wire h_s_wallace_rca24_and_5_18_y0;
  wire h_s_wallace_rca24_and_4_19_y0;
  wire h_s_wallace_rca24_fa317_y2;
  wire h_s_wallace_rca24_fa317_y4;
  wire h_s_wallace_rca24_and_6_18_y0;
  wire h_s_wallace_rca24_and_5_19_y0;
  wire h_s_wallace_rca24_fa318_y2;
  wire h_s_wallace_rca24_fa318_y4;
  wire h_s_wallace_rca24_and_5_20_y0;
  wire h_s_wallace_rca24_and_4_21_y0;
  wire h_s_wallace_rca24_fa319_y2;
  wire h_s_wallace_rca24_fa319_y4;
  wire h_s_wallace_rca24_and_5_21_y0;
  wire h_s_wallace_rca24_and_4_22_y0;
  wire h_s_wallace_rca24_fa320_y2;
  wire h_s_wallace_rca24_fa320_y4;
  wire h_s_wallace_rca24_and_5_22_y0;
  wire h_s_wallace_rca24_nand_4_23_y0;
  wire h_s_wallace_rca24_fa321_y2;
  wire h_s_wallace_rca24_fa321_y4;
  wire h_s_wallace_rca24_nand_5_23_y0;
  wire h_s_wallace_rca24_fa322_y2;
  wire h_s_wallace_rca24_fa322_y4;
  wire h_s_wallace_rca24_fa323_y2;
  wire h_s_wallace_rca24_fa323_y4;
  wire h_s_wallace_rca24_fa324_y2;
  wire h_s_wallace_rca24_fa324_y4;
  wire h_s_wallace_rca24_fa325_y2;
  wire h_s_wallace_rca24_fa325_y4;
  wire h_s_wallace_rca24_fa326_y2;
  wire h_s_wallace_rca24_fa326_y4;
  wire h_s_wallace_rca24_fa327_y2;
  wire h_s_wallace_rca24_fa327_y4;
  wire h_s_wallace_rca24_fa328_y2;
  wire h_s_wallace_rca24_fa328_y4;
  wire h_s_wallace_rca24_fa329_y2;
  wire h_s_wallace_rca24_fa329_y4;
  wire h_s_wallace_rca24_ha10_y0;
  wire h_s_wallace_rca24_ha10_y1;
  wire h_s_wallace_rca24_fa330_y2;
  wire h_s_wallace_rca24_fa330_y4;
  wire h_s_wallace_rca24_fa331_y2;
  wire h_s_wallace_rca24_fa331_y4;
  wire h_s_wallace_rca24_fa332_y2;
  wire h_s_wallace_rca24_fa332_y4;
  wire h_s_wallace_rca24_fa333_y2;
  wire h_s_wallace_rca24_fa333_y4;
  wire h_s_wallace_rca24_fa334_y2;
  wire h_s_wallace_rca24_fa334_y4;
  wire h_s_wallace_rca24_fa335_y2;
  wire h_s_wallace_rca24_fa335_y4;
  wire h_s_wallace_rca24_fa336_y2;
  wire h_s_wallace_rca24_fa336_y4;
  wire h_s_wallace_rca24_and_0_20_y0;
  wire h_s_wallace_rca24_fa337_y2;
  wire h_s_wallace_rca24_fa337_y4;
  wire h_s_wallace_rca24_and_1_20_y0;
  wire h_s_wallace_rca24_and_0_21_y0;
  wire h_s_wallace_rca24_fa338_y2;
  wire h_s_wallace_rca24_fa338_y4;
  wire h_s_wallace_rca24_and_2_20_y0;
  wire h_s_wallace_rca24_and_1_21_y0;
  wire h_s_wallace_rca24_fa339_y2;
  wire h_s_wallace_rca24_fa339_y4;
  wire h_s_wallace_rca24_and_3_20_y0;
  wire h_s_wallace_rca24_and_2_21_y0;
  wire h_s_wallace_rca24_fa340_y2;
  wire h_s_wallace_rca24_fa340_y4;
  wire h_s_wallace_rca24_and_4_20_y0;
  wire h_s_wallace_rca24_and_3_21_y0;
  wire h_s_wallace_rca24_fa341_y2;
  wire h_s_wallace_rca24_fa341_y4;
  wire h_s_wallace_rca24_and_3_22_y0;
  wire h_s_wallace_rca24_nand_2_23_y0;
  wire h_s_wallace_rca24_fa342_y2;
  wire h_s_wallace_rca24_fa342_y4;
  wire h_s_wallace_rca24_nand_3_23_y0;
  wire h_s_wallace_rca24_fa343_y2;
  wire h_s_wallace_rca24_fa343_y4;
  wire h_s_wallace_rca24_fa344_y2;
  wire h_s_wallace_rca24_fa344_y4;
  wire h_s_wallace_rca24_fa345_y2;
  wire h_s_wallace_rca24_fa345_y4;
  wire h_s_wallace_rca24_fa346_y2;
  wire h_s_wallace_rca24_fa346_y4;
  wire h_s_wallace_rca24_fa347_y2;
  wire h_s_wallace_rca24_fa347_y4;
  wire h_s_wallace_rca24_fa348_y2;
  wire h_s_wallace_rca24_fa348_y4;
  wire h_s_wallace_rca24_fa349_y2;
  wire h_s_wallace_rca24_fa349_y4;
  wire h_s_wallace_rca24_fa350_y2;
  wire h_s_wallace_rca24_fa350_y4;
  wire h_s_wallace_rca24_fa351_y2;
  wire h_s_wallace_rca24_fa351_y4;
  wire h_s_wallace_rca24_ha11_y0;
  wire h_s_wallace_rca24_ha11_y1;
  wire h_s_wallace_rca24_fa352_y2;
  wire h_s_wallace_rca24_fa352_y4;
  wire h_s_wallace_rca24_fa353_y2;
  wire h_s_wallace_rca24_fa353_y4;
  wire h_s_wallace_rca24_fa354_y2;
  wire h_s_wallace_rca24_fa354_y4;
  wire h_s_wallace_rca24_fa355_y2;
  wire h_s_wallace_rca24_fa355_y4;
  wire h_s_wallace_rca24_fa356_y2;
  wire h_s_wallace_rca24_fa356_y4;
  wire h_s_wallace_rca24_fa357_y2;
  wire h_s_wallace_rca24_fa357_y4;
  wire h_s_wallace_rca24_fa358_y2;
  wire h_s_wallace_rca24_fa358_y4;
  wire h_s_wallace_rca24_fa359_y2;
  wire h_s_wallace_rca24_fa359_y4;
  wire h_s_wallace_rca24_and_0_22_y0;
  wire h_s_wallace_rca24_fa360_y2;
  wire h_s_wallace_rca24_fa360_y4;
  wire h_s_wallace_rca24_and_1_22_y0;
  wire h_s_wallace_rca24_nand_0_23_y0;
  wire h_s_wallace_rca24_fa361_y2;
  wire h_s_wallace_rca24_fa361_y4;
  wire h_s_wallace_rca24_and_2_22_y0;
  wire h_s_wallace_rca24_nand_1_23_y0;
  wire h_s_wallace_rca24_fa362_y2;
  wire h_s_wallace_rca24_fa362_y4;
  wire h_s_wallace_rca24_fa363_y2;
  wire h_s_wallace_rca24_fa363_y4;
  wire h_s_wallace_rca24_fa364_y2;
  wire h_s_wallace_rca24_fa364_y4;
  wire h_s_wallace_rca24_fa365_y2;
  wire h_s_wallace_rca24_fa365_y4;
  wire h_s_wallace_rca24_fa366_y2;
  wire h_s_wallace_rca24_fa366_y4;
  wire h_s_wallace_rca24_fa367_y2;
  wire h_s_wallace_rca24_fa367_y4;
  wire h_s_wallace_rca24_fa368_y2;
  wire h_s_wallace_rca24_fa368_y4;
  wire h_s_wallace_rca24_fa369_y2;
  wire h_s_wallace_rca24_fa369_y4;
  wire h_s_wallace_rca24_fa370_y2;
  wire h_s_wallace_rca24_fa370_y4;
  wire h_s_wallace_rca24_fa371_y2;
  wire h_s_wallace_rca24_fa371_y4;
  wire h_s_wallace_rca24_ha12_y0;
  wire h_s_wallace_rca24_ha12_y1;
  wire h_s_wallace_rca24_fa372_y2;
  wire h_s_wallace_rca24_fa372_y4;
  wire h_s_wallace_rca24_fa373_y2;
  wire h_s_wallace_rca24_fa373_y4;
  wire h_s_wallace_rca24_fa374_y2;
  wire h_s_wallace_rca24_fa374_y4;
  wire h_s_wallace_rca24_fa375_y2;
  wire h_s_wallace_rca24_fa375_y4;
  wire h_s_wallace_rca24_fa376_y2;
  wire h_s_wallace_rca24_fa376_y4;
  wire h_s_wallace_rca24_fa377_y2;
  wire h_s_wallace_rca24_fa377_y4;
  wire h_s_wallace_rca24_fa378_y2;
  wire h_s_wallace_rca24_fa378_y4;
  wire h_s_wallace_rca24_fa379_y2;
  wire h_s_wallace_rca24_fa379_y4;
  wire h_s_wallace_rca24_fa380_y2;
  wire h_s_wallace_rca24_fa380_y4;
  wire h_s_wallace_rca24_fa381_y2;
  wire h_s_wallace_rca24_fa381_y4;
  wire h_s_wallace_rca24_fa382_y2;
  wire h_s_wallace_rca24_fa382_y4;
  wire h_s_wallace_rca24_fa383_y2;
  wire h_s_wallace_rca24_fa383_y4;
  wire h_s_wallace_rca24_fa384_y2;
  wire h_s_wallace_rca24_fa384_y4;
  wire h_s_wallace_rca24_fa385_y2;
  wire h_s_wallace_rca24_fa385_y4;
  wire h_s_wallace_rca24_fa386_y2;
  wire h_s_wallace_rca24_fa386_y4;
  wire h_s_wallace_rca24_fa387_y2;
  wire h_s_wallace_rca24_fa387_y4;
  wire h_s_wallace_rca24_fa388_y2;
  wire h_s_wallace_rca24_fa388_y4;
  wire h_s_wallace_rca24_fa389_y2;
  wire h_s_wallace_rca24_fa389_y4;
  wire h_s_wallace_rca24_ha13_y0;
  wire h_s_wallace_rca24_ha13_y1;
  wire h_s_wallace_rca24_fa390_y2;
  wire h_s_wallace_rca24_fa390_y4;
  wire h_s_wallace_rca24_fa391_y2;
  wire h_s_wallace_rca24_fa391_y4;
  wire h_s_wallace_rca24_fa392_y2;
  wire h_s_wallace_rca24_fa392_y4;
  wire h_s_wallace_rca24_fa393_y2;
  wire h_s_wallace_rca24_fa393_y4;
  wire h_s_wallace_rca24_fa394_y2;
  wire h_s_wallace_rca24_fa394_y4;
  wire h_s_wallace_rca24_fa395_y2;
  wire h_s_wallace_rca24_fa395_y4;
  wire h_s_wallace_rca24_fa396_y2;
  wire h_s_wallace_rca24_fa396_y4;
  wire h_s_wallace_rca24_fa397_y2;
  wire h_s_wallace_rca24_fa397_y4;
  wire h_s_wallace_rca24_fa398_y2;
  wire h_s_wallace_rca24_fa398_y4;
  wire h_s_wallace_rca24_fa399_y2;
  wire h_s_wallace_rca24_fa399_y4;
  wire h_s_wallace_rca24_fa400_y2;
  wire h_s_wallace_rca24_fa400_y4;
  wire h_s_wallace_rca24_fa401_y2;
  wire h_s_wallace_rca24_fa401_y4;
  wire h_s_wallace_rca24_fa402_y2;
  wire h_s_wallace_rca24_fa402_y4;
  wire h_s_wallace_rca24_fa403_y2;
  wire h_s_wallace_rca24_fa403_y4;
  wire h_s_wallace_rca24_fa404_y2;
  wire h_s_wallace_rca24_fa404_y4;
  wire h_s_wallace_rca24_fa405_y2;
  wire h_s_wallace_rca24_fa405_y4;
  wire h_s_wallace_rca24_ha14_y0;
  wire h_s_wallace_rca24_ha14_y1;
  wire h_s_wallace_rca24_fa406_y2;
  wire h_s_wallace_rca24_fa406_y4;
  wire h_s_wallace_rca24_fa407_y2;
  wire h_s_wallace_rca24_fa407_y4;
  wire h_s_wallace_rca24_fa408_y2;
  wire h_s_wallace_rca24_fa408_y4;
  wire h_s_wallace_rca24_fa409_y2;
  wire h_s_wallace_rca24_fa409_y4;
  wire h_s_wallace_rca24_fa410_y2;
  wire h_s_wallace_rca24_fa410_y4;
  wire h_s_wallace_rca24_fa411_y2;
  wire h_s_wallace_rca24_fa411_y4;
  wire h_s_wallace_rca24_fa412_y2;
  wire h_s_wallace_rca24_fa412_y4;
  wire h_s_wallace_rca24_fa413_y2;
  wire h_s_wallace_rca24_fa413_y4;
  wire h_s_wallace_rca24_fa414_y2;
  wire h_s_wallace_rca24_fa414_y4;
  wire h_s_wallace_rca24_fa415_y2;
  wire h_s_wallace_rca24_fa415_y4;
  wire h_s_wallace_rca24_fa416_y2;
  wire h_s_wallace_rca24_fa416_y4;
  wire h_s_wallace_rca24_fa417_y2;
  wire h_s_wallace_rca24_fa417_y4;
  wire h_s_wallace_rca24_fa418_y2;
  wire h_s_wallace_rca24_fa418_y4;
  wire h_s_wallace_rca24_fa419_y2;
  wire h_s_wallace_rca24_fa419_y4;
  wire h_s_wallace_rca24_ha15_y0;
  wire h_s_wallace_rca24_ha15_y1;
  wire h_s_wallace_rca24_fa420_y2;
  wire h_s_wallace_rca24_fa420_y4;
  wire h_s_wallace_rca24_fa421_y2;
  wire h_s_wallace_rca24_fa421_y4;
  wire h_s_wallace_rca24_fa422_y2;
  wire h_s_wallace_rca24_fa422_y4;
  wire h_s_wallace_rca24_fa423_y2;
  wire h_s_wallace_rca24_fa423_y4;
  wire h_s_wallace_rca24_fa424_y2;
  wire h_s_wallace_rca24_fa424_y4;
  wire h_s_wallace_rca24_fa425_y2;
  wire h_s_wallace_rca24_fa425_y4;
  wire h_s_wallace_rca24_fa426_y2;
  wire h_s_wallace_rca24_fa426_y4;
  wire h_s_wallace_rca24_fa427_y2;
  wire h_s_wallace_rca24_fa427_y4;
  wire h_s_wallace_rca24_fa428_y2;
  wire h_s_wallace_rca24_fa428_y4;
  wire h_s_wallace_rca24_fa429_y2;
  wire h_s_wallace_rca24_fa429_y4;
  wire h_s_wallace_rca24_fa430_y2;
  wire h_s_wallace_rca24_fa430_y4;
  wire h_s_wallace_rca24_fa431_y2;
  wire h_s_wallace_rca24_fa431_y4;
  wire h_s_wallace_rca24_ha16_y0;
  wire h_s_wallace_rca24_ha16_y1;
  wire h_s_wallace_rca24_fa432_y2;
  wire h_s_wallace_rca24_fa432_y4;
  wire h_s_wallace_rca24_fa433_y2;
  wire h_s_wallace_rca24_fa433_y4;
  wire h_s_wallace_rca24_fa434_y2;
  wire h_s_wallace_rca24_fa434_y4;
  wire h_s_wallace_rca24_fa435_y2;
  wire h_s_wallace_rca24_fa435_y4;
  wire h_s_wallace_rca24_fa436_y2;
  wire h_s_wallace_rca24_fa436_y4;
  wire h_s_wallace_rca24_fa437_y2;
  wire h_s_wallace_rca24_fa437_y4;
  wire h_s_wallace_rca24_fa438_y2;
  wire h_s_wallace_rca24_fa438_y4;
  wire h_s_wallace_rca24_fa439_y2;
  wire h_s_wallace_rca24_fa439_y4;
  wire h_s_wallace_rca24_fa440_y2;
  wire h_s_wallace_rca24_fa440_y4;
  wire h_s_wallace_rca24_fa441_y2;
  wire h_s_wallace_rca24_fa441_y4;
  wire h_s_wallace_rca24_ha17_y0;
  wire h_s_wallace_rca24_ha17_y1;
  wire h_s_wallace_rca24_fa442_y2;
  wire h_s_wallace_rca24_fa442_y4;
  wire h_s_wallace_rca24_fa443_y2;
  wire h_s_wallace_rca24_fa443_y4;
  wire h_s_wallace_rca24_fa444_y2;
  wire h_s_wallace_rca24_fa444_y4;
  wire h_s_wallace_rca24_fa445_y2;
  wire h_s_wallace_rca24_fa445_y4;
  wire h_s_wallace_rca24_fa446_y2;
  wire h_s_wallace_rca24_fa446_y4;
  wire h_s_wallace_rca24_fa447_y2;
  wire h_s_wallace_rca24_fa447_y4;
  wire h_s_wallace_rca24_fa448_y2;
  wire h_s_wallace_rca24_fa448_y4;
  wire h_s_wallace_rca24_fa449_y2;
  wire h_s_wallace_rca24_fa449_y4;
  wire h_s_wallace_rca24_ha18_y0;
  wire h_s_wallace_rca24_ha18_y1;
  wire h_s_wallace_rca24_fa450_y2;
  wire h_s_wallace_rca24_fa450_y4;
  wire h_s_wallace_rca24_fa451_y2;
  wire h_s_wallace_rca24_fa451_y4;
  wire h_s_wallace_rca24_fa452_y2;
  wire h_s_wallace_rca24_fa452_y4;
  wire h_s_wallace_rca24_fa453_y2;
  wire h_s_wallace_rca24_fa453_y4;
  wire h_s_wallace_rca24_fa454_y2;
  wire h_s_wallace_rca24_fa454_y4;
  wire h_s_wallace_rca24_fa455_y2;
  wire h_s_wallace_rca24_fa455_y4;
  wire h_s_wallace_rca24_ha19_y0;
  wire h_s_wallace_rca24_ha19_y1;
  wire h_s_wallace_rca24_fa456_y2;
  wire h_s_wallace_rca24_fa456_y4;
  wire h_s_wallace_rca24_fa457_y2;
  wire h_s_wallace_rca24_fa457_y4;
  wire h_s_wallace_rca24_fa458_y2;
  wire h_s_wallace_rca24_fa458_y4;
  wire h_s_wallace_rca24_fa459_y2;
  wire h_s_wallace_rca24_fa459_y4;
  wire h_s_wallace_rca24_ha20_y0;
  wire h_s_wallace_rca24_ha20_y1;
  wire h_s_wallace_rca24_fa460_y2;
  wire h_s_wallace_rca24_fa460_y4;
  wire h_s_wallace_rca24_fa461_y2;
  wire h_s_wallace_rca24_fa461_y4;
  wire h_s_wallace_rca24_ha21_y0;
  wire h_s_wallace_rca24_ha21_y1;
  wire h_s_wallace_rca24_fa462_y2;
  wire h_s_wallace_rca24_fa462_y4;
  wire h_s_wallace_rca24_fa463_y2;
  wire h_s_wallace_rca24_fa463_y4;
  wire h_s_wallace_rca24_fa464_y2;
  wire h_s_wallace_rca24_fa464_y4;
  wire h_s_wallace_rca24_fa465_y2;
  wire h_s_wallace_rca24_fa465_y4;
  wire h_s_wallace_rca24_fa466_y2;
  wire h_s_wallace_rca24_fa466_y4;
  wire h_s_wallace_rca24_fa467_y2;
  wire h_s_wallace_rca24_fa467_y4;
  wire h_s_wallace_rca24_fa468_y2;
  wire h_s_wallace_rca24_fa468_y4;
  wire h_s_wallace_rca24_fa469_y2;
  wire h_s_wallace_rca24_fa469_y4;
  wire h_s_wallace_rca24_fa470_y2;
  wire h_s_wallace_rca24_fa470_y4;
  wire h_s_wallace_rca24_fa471_y2;
  wire h_s_wallace_rca24_fa471_y4;
  wire h_s_wallace_rca24_fa472_y2;
  wire h_s_wallace_rca24_fa472_y4;
  wire h_s_wallace_rca24_fa473_y2;
  wire h_s_wallace_rca24_fa473_y4;
  wire h_s_wallace_rca24_fa474_y2;
  wire h_s_wallace_rca24_fa474_y4;
  wire h_s_wallace_rca24_fa475_y2;
  wire h_s_wallace_rca24_fa475_y4;
  wire h_s_wallace_rca24_fa476_y2;
  wire h_s_wallace_rca24_fa476_y4;
  wire h_s_wallace_rca24_fa477_y2;
  wire h_s_wallace_rca24_fa477_y4;
  wire h_s_wallace_rca24_fa478_y2;
  wire h_s_wallace_rca24_fa478_y4;
  wire h_s_wallace_rca24_fa479_y2;
  wire h_s_wallace_rca24_fa479_y4;
  wire h_s_wallace_rca24_fa480_y2;
  wire h_s_wallace_rca24_fa480_y4;
  wire h_s_wallace_rca24_fa481_y2;
  wire h_s_wallace_rca24_fa481_y4;
  wire h_s_wallace_rca24_nand_21_23_y0;
  wire h_s_wallace_rca24_fa482_y2;
  wire h_s_wallace_rca24_fa482_y4;
  wire h_s_wallace_rca24_nand_23_22_y0;
  wire h_s_wallace_rca24_fa483_y2;
  wire h_s_wallace_rca24_fa483_y4;
  wire h_s_wallace_rca24_and_0_0_y0;
  wire h_s_wallace_rca24_and_1_0_y0;
  wire h_s_wallace_rca24_and_0_2_y0;
  wire h_s_wallace_rca24_nand_22_23_y0;
  wire h_s_wallace_rca24_and_0_1_y0;
  wire h_s_wallace_rca24_and_23_23_y0;
  wire [45:0] h_s_wallace_rca24_u_rca_u_rca_a;
  wire [45:0] h_s_wallace_rca24_u_rca_u_rca_b;
  wire [46:0] h_s_wallace_rca24_u_rca_out;
  wire h_s_wallace_rca24_u_rca_ha_y0;
  wire h_s_wallace_rca24_u_rca_fa1_y2;
  wire h_s_wallace_rca24_u_rca_fa2_y2;
  wire h_s_wallace_rca24_u_rca_fa3_y2;
  wire h_s_wallace_rca24_u_rca_fa4_y2;
  wire h_s_wallace_rca24_u_rca_fa5_y2;
  wire h_s_wallace_rca24_u_rca_fa6_y2;
  wire h_s_wallace_rca24_u_rca_fa7_y2;
  wire h_s_wallace_rca24_u_rca_fa8_y2;
  wire h_s_wallace_rca24_u_rca_fa9_y2;
  wire h_s_wallace_rca24_u_rca_fa10_y2;
  wire h_s_wallace_rca24_u_rca_fa11_y2;
  wire h_s_wallace_rca24_u_rca_fa12_y2;
  wire h_s_wallace_rca24_u_rca_fa13_y2;
  wire h_s_wallace_rca24_u_rca_fa14_y2;
  wire h_s_wallace_rca24_u_rca_fa15_y2;
  wire h_s_wallace_rca24_u_rca_fa16_y2;
  wire h_s_wallace_rca24_u_rca_fa17_y2;
  wire h_s_wallace_rca24_u_rca_fa18_y2;
  wire h_s_wallace_rca24_u_rca_fa19_y2;
  wire h_s_wallace_rca24_u_rca_fa20_y2;
  wire h_s_wallace_rca24_u_rca_fa21_y2;
  wire h_s_wallace_rca24_u_rca_fa22_y2;
  wire h_s_wallace_rca24_u_rca_fa23_y2;
  wire h_s_wallace_rca24_u_rca_fa24_y2;
  wire h_s_wallace_rca24_u_rca_fa25_y2;
  wire h_s_wallace_rca24_u_rca_fa26_y2;
  wire h_s_wallace_rca24_u_rca_fa27_y2;
  wire h_s_wallace_rca24_u_rca_fa28_y2;
  wire h_s_wallace_rca24_u_rca_fa29_y2;
  wire h_s_wallace_rca24_u_rca_fa30_y2;
  wire h_s_wallace_rca24_u_rca_fa31_y2;
  wire h_s_wallace_rca24_u_rca_fa32_y2;
  wire h_s_wallace_rca24_u_rca_fa33_y2;
  wire h_s_wallace_rca24_u_rca_fa34_y2;
  wire h_s_wallace_rca24_u_rca_fa35_y2;
  wire h_s_wallace_rca24_u_rca_fa36_y2;
  wire h_s_wallace_rca24_u_rca_fa37_y2;
  wire h_s_wallace_rca24_u_rca_fa38_y2;
  wire h_s_wallace_rca24_u_rca_fa39_y2;
  wire h_s_wallace_rca24_u_rca_fa40_y2;
  wire h_s_wallace_rca24_u_rca_fa41_y2;
  wire h_s_wallace_rca24_u_rca_fa42_y2;
  wire h_s_wallace_rca24_u_rca_fa43_y2;
  wire h_s_wallace_rca24_u_rca_fa44_y2;
  wire h_s_wallace_rca24_u_rca_fa45_y2;
  wire h_s_wallace_rca24_u_rca_fa45_y4;
  wire h_s_wallace_rca24_xor0_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_wallace_rca24_and_2_0_y0(a_2, b_0, h_s_wallace_rca24_and_2_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_1_y0(a_1, b_1, h_s_wallace_rca24_and_1_1_y0);
  ha ha_h_s_wallace_rca24_ha0_y0(h_s_wallace_rca24_and_2_0_y0, h_s_wallace_rca24_and_1_1_y0, h_s_wallace_rca24_ha0_y0, h_s_wallace_rca24_ha0_y1);
  and_gate and_gate_h_s_wallace_rca24_and_3_0_y0(a_3, b_0, h_s_wallace_rca24_and_3_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_1_y0(a_2, b_1, h_s_wallace_rca24_and_2_1_y0);
  fa fa_h_s_wallace_rca24_fa0_y2(h_s_wallace_rca24_ha0_y1, h_s_wallace_rca24_and_3_0_y0, h_s_wallace_rca24_and_2_1_y0, h_s_wallace_rca24_fa0_y2, h_s_wallace_rca24_fa0_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_0_y0(a_4, b_0, h_s_wallace_rca24_and_4_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_1_y0(a_3, b_1, h_s_wallace_rca24_and_3_1_y0);
  fa fa_h_s_wallace_rca24_fa1_y2(h_s_wallace_rca24_fa0_y4, h_s_wallace_rca24_and_4_0_y0, h_s_wallace_rca24_and_3_1_y0, h_s_wallace_rca24_fa1_y2, h_s_wallace_rca24_fa1_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_0_y0(a_5, b_0, h_s_wallace_rca24_and_5_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_1_y0(a_4, b_1, h_s_wallace_rca24_and_4_1_y0);
  fa fa_h_s_wallace_rca24_fa2_y2(h_s_wallace_rca24_fa1_y4, h_s_wallace_rca24_and_5_0_y0, h_s_wallace_rca24_and_4_1_y0, h_s_wallace_rca24_fa2_y2, h_s_wallace_rca24_fa2_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_0_y0(a_6, b_0, h_s_wallace_rca24_and_6_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_1_y0(a_5, b_1, h_s_wallace_rca24_and_5_1_y0);
  fa fa_h_s_wallace_rca24_fa3_y2(h_s_wallace_rca24_fa2_y4, h_s_wallace_rca24_and_6_0_y0, h_s_wallace_rca24_and_5_1_y0, h_s_wallace_rca24_fa3_y2, h_s_wallace_rca24_fa3_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_0_y0(a_7, b_0, h_s_wallace_rca24_and_7_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_1_y0(a_6, b_1, h_s_wallace_rca24_and_6_1_y0);
  fa fa_h_s_wallace_rca24_fa4_y2(h_s_wallace_rca24_fa3_y4, h_s_wallace_rca24_and_7_0_y0, h_s_wallace_rca24_and_6_1_y0, h_s_wallace_rca24_fa4_y2, h_s_wallace_rca24_fa4_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_0_y0(a_8, b_0, h_s_wallace_rca24_and_8_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_1_y0(a_7, b_1, h_s_wallace_rca24_and_7_1_y0);
  fa fa_h_s_wallace_rca24_fa5_y2(h_s_wallace_rca24_fa4_y4, h_s_wallace_rca24_and_8_0_y0, h_s_wallace_rca24_and_7_1_y0, h_s_wallace_rca24_fa5_y2, h_s_wallace_rca24_fa5_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_0_y0(a_9, b_0, h_s_wallace_rca24_and_9_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_1_y0(a_8, b_1, h_s_wallace_rca24_and_8_1_y0);
  fa fa_h_s_wallace_rca24_fa6_y2(h_s_wallace_rca24_fa5_y4, h_s_wallace_rca24_and_9_0_y0, h_s_wallace_rca24_and_8_1_y0, h_s_wallace_rca24_fa6_y2, h_s_wallace_rca24_fa6_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_0_y0(a_10, b_0, h_s_wallace_rca24_and_10_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_1_y0(a_9, b_1, h_s_wallace_rca24_and_9_1_y0);
  fa fa_h_s_wallace_rca24_fa7_y2(h_s_wallace_rca24_fa6_y4, h_s_wallace_rca24_and_10_0_y0, h_s_wallace_rca24_and_9_1_y0, h_s_wallace_rca24_fa7_y2, h_s_wallace_rca24_fa7_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_0_y0(a_11, b_0, h_s_wallace_rca24_and_11_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_1_y0(a_10, b_1, h_s_wallace_rca24_and_10_1_y0);
  fa fa_h_s_wallace_rca24_fa8_y2(h_s_wallace_rca24_fa7_y4, h_s_wallace_rca24_and_11_0_y0, h_s_wallace_rca24_and_10_1_y0, h_s_wallace_rca24_fa8_y2, h_s_wallace_rca24_fa8_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_0_y0(a_12, b_0, h_s_wallace_rca24_and_12_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_1_y0(a_11, b_1, h_s_wallace_rca24_and_11_1_y0);
  fa fa_h_s_wallace_rca24_fa9_y2(h_s_wallace_rca24_fa8_y4, h_s_wallace_rca24_and_12_0_y0, h_s_wallace_rca24_and_11_1_y0, h_s_wallace_rca24_fa9_y2, h_s_wallace_rca24_fa9_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_0_y0(a_13, b_0, h_s_wallace_rca24_and_13_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_1_y0(a_12, b_1, h_s_wallace_rca24_and_12_1_y0);
  fa fa_h_s_wallace_rca24_fa10_y2(h_s_wallace_rca24_fa9_y4, h_s_wallace_rca24_and_13_0_y0, h_s_wallace_rca24_and_12_1_y0, h_s_wallace_rca24_fa10_y2, h_s_wallace_rca24_fa10_y4);
  and_gate and_gate_h_s_wallace_rca24_and_14_0_y0(a_14, b_0, h_s_wallace_rca24_and_14_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_13_1_y0(a_13, b_1, h_s_wallace_rca24_and_13_1_y0);
  fa fa_h_s_wallace_rca24_fa11_y2(h_s_wallace_rca24_fa10_y4, h_s_wallace_rca24_and_14_0_y0, h_s_wallace_rca24_and_13_1_y0, h_s_wallace_rca24_fa11_y2, h_s_wallace_rca24_fa11_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_0_y0(a_15, b_0, h_s_wallace_rca24_and_15_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_1_y0(a_14, b_1, h_s_wallace_rca24_and_14_1_y0);
  fa fa_h_s_wallace_rca24_fa12_y2(h_s_wallace_rca24_fa11_y4, h_s_wallace_rca24_and_15_0_y0, h_s_wallace_rca24_and_14_1_y0, h_s_wallace_rca24_fa12_y2, h_s_wallace_rca24_fa12_y4);
  and_gate and_gate_h_s_wallace_rca24_and_16_0_y0(a_16, b_0, h_s_wallace_rca24_and_16_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_15_1_y0(a_15, b_1, h_s_wallace_rca24_and_15_1_y0);
  fa fa_h_s_wallace_rca24_fa13_y2(h_s_wallace_rca24_fa12_y4, h_s_wallace_rca24_and_16_0_y0, h_s_wallace_rca24_and_15_1_y0, h_s_wallace_rca24_fa13_y2, h_s_wallace_rca24_fa13_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_0_y0(a_17, b_0, h_s_wallace_rca24_and_17_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_1_y0(a_16, b_1, h_s_wallace_rca24_and_16_1_y0);
  fa fa_h_s_wallace_rca24_fa14_y2(h_s_wallace_rca24_fa13_y4, h_s_wallace_rca24_and_17_0_y0, h_s_wallace_rca24_and_16_1_y0, h_s_wallace_rca24_fa14_y2, h_s_wallace_rca24_fa14_y4);
  and_gate and_gate_h_s_wallace_rca24_and_18_0_y0(a_18, b_0, h_s_wallace_rca24_and_18_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_17_1_y0(a_17, b_1, h_s_wallace_rca24_and_17_1_y0);
  fa fa_h_s_wallace_rca24_fa15_y2(h_s_wallace_rca24_fa14_y4, h_s_wallace_rca24_and_18_0_y0, h_s_wallace_rca24_and_17_1_y0, h_s_wallace_rca24_fa15_y2, h_s_wallace_rca24_fa15_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_0_y0(a_19, b_0, h_s_wallace_rca24_and_19_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_1_y0(a_18, b_1, h_s_wallace_rca24_and_18_1_y0);
  fa fa_h_s_wallace_rca24_fa16_y2(h_s_wallace_rca24_fa15_y4, h_s_wallace_rca24_and_19_0_y0, h_s_wallace_rca24_and_18_1_y0, h_s_wallace_rca24_fa16_y2, h_s_wallace_rca24_fa16_y4);
  and_gate and_gate_h_s_wallace_rca24_and_20_0_y0(a_20, b_0, h_s_wallace_rca24_and_20_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_19_1_y0(a_19, b_1, h_s_wallace_rca24_and_19_1_y0);
  fa fa_h_s_wallace_rca24_fa17_y2(h_s_wallace_rca24_fa16_y4, h_s_wallace_rca24_and_20_0_y0, h_s_wallace_rca24_and_19_1_y0, h_s_wallace_rca24_fa17_y2, h_s_wallace_rca24_fa17_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_0_y0(a_21, b_0, h_s_wallace_rca24_and_21_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_1_y0(a_20, b_1, h_s_wallace_rca24_and_20_1_y0);
  fa fa_h_s_wallace_rca24_fa18_y2(h_s_wallace_rca24_fa17_y4, h_s_wallace_rca24_and_21_0_y0, h_s_wallace_rca24_and_20_1_y0, h_s_wallace_rca24_fa18_y2, h_s_wallace_rca24_fa18_y4);
  and_gate and_gate_h_s_wallace_rca24_and_22_0_y0(a_22, b_0, h_s_wallace_rca24_and_22_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_21_1_y0(a_21, b_1, h_s_wallace_rca24_and_21_1_y0);
  fa fa_h_s_wallace_rca24_fa19_y2(h_s_wallace_rca24_fa18_y4, h_s_wallace_rca24_and_22_0_y0, h_s_wallace_rca24_and_21_1_y0, h_s_wallace_rca24_fa19_y2, h_s_wallace_rca24_fa19_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_0_y0(a_23, b_0, h_s_wallace_rca24_nand_23_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_1_y0(a_22, b_1, h_s_wallace_rca24_and_22_1_y0);
  fa fa_h_s_wallace_rca24_fa20_y2(h_s_wallace_rca24_fa19_y4, h_s_wallace_rca24_nand_23_0_y0, h_s_wallace_rca24_and_22_1_y0, h_s_wallace_rca24_fa20_y2, h_s_wallace_rca24_fa20_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_1_y0(a_23, b_1, h_s_wallace_rca24_nand_23_1_y0);
  fa fa_h_s_wallace_rca24_fa21_y2(h_s_wallace_rca24_fa20_y4, constant_wire_1, h_s_wallace_rca24_nand_23_1_y0, h_s_wallace_rca24_fa21_y2, h_s_wallace_rca24_fa21_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_2_y0(a_23, b_2, h_s_wallace_rca24_nand_23_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_3_y0(a_22, b_3, h_s_wallace_rca24_and_22_3_y0);
  fa fa_h_s_wallace_rca24_fa22_y2(h_s_wallace_rca24_fa21_y4, h_s_wallace_rca24_nand_23_2_y0, h_s_wallace_rca24_and_22_3_y0, h_s_wallace_rca24_fa22_y2, h_s_wallace_rca24_fa22_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_3_y0(a_23, b_3, h_s_wallace_rca24_nand_23_3_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_4_y0(a_22, b_4, h_s_wallace_rca24_and_22_4_y0);
  fa fa_h_s_wallace_rca24_fa23_y2(h_s_wallace_rca24_fa22_y4, h_s_wallace_rca24_nand_23_3_y0, h_s_wallace_rca24_and_22_4_y0, h_s_wallace_rca24_fa23_y2, h_s_wallace_rca24_fa23_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_4_y0(a_23, b_4, h_s_wallace_rca24_nand_23_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_5_y0(a_22, b_5, h_s_wallace_rca24_and_22_5_y0);
  fa fa_h_s_wallace_rca24_fa24_y2(h_s_wallace_rca24_fa23_y4, h_s_wallace_rca24_nand_23_4_y0, h_s_wallace_rca24_and_22_5_y0, h_s_wallace_rca24_fa24_y2, h_s_wallace_rca24_fa24_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_5_y0(a_23, b_5, h_s_wallace_rca24_nand_23_5_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_6_y0(a_22, b_6, h_s_wallace_rca24_and_22_6_y0);
  fa fa_h_s_wallace_rca24_fa25_y2(h_s_wallace_rca24_fa24_y4, h_s_wallace_rca24_nand_23_5_y0, h_s_wallace_rca24_and_22_6_y0, h_s_wallace_rca24_fa25_y2, h_s_wallace_rca24_fa25_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_6_y0(a_23, b_6, h_s_wallace_rca24_nand_23_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_7_y0(a_22, b_7, h_s_wallace_rca24_and_22_7_y0);
  fa fa_h_s_wallace_rca24_fa26_y2(h_s_wallace_rca24_fa25_y4, h_s_wallace_rca24_nand_23_6_y0, h_s_wallace_rca24_and_22_7_y0, h_s_wallace_rca24_fa26_y2, h_s_wallace_rca24_fa26_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_7_y0(a_23, b_7, h_s_wallace_rca24_nand_23_7_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_8_y0(a_22, b_8, h_s_wallace_rca24_and_22_8_y0);
  fa fa_h_s_wallace_rca24_fa27_y2(h_s_wallace_rca24_fa26_y4, h_s_wallace_rca24_nand_23_7_y0, h_s_wallace_rca24_and_22_8_y0, h_s_wallace_rca24_fa27_y2, h_s_wallace_rca24_fa27_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_8_y0(a_23, b_8, h_s_wallace_rca24_nand_23_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_9_y0(a_22, b_9, h_s_wallace_rca24_and_22_9_y0);
  fa fa_h_s_wallace_rca24_fa28_y2(h_s_wallace_rca24_fa27_y4, h_s_wallace_rca24_nand_23_8_y0, h_s_wallace_rca24_and_22_9_y0, h_s_wallace_rca24_fa28_y2, h_s_wallace_rca24_fa28_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_9_y0(a_23, b_9, h_s_wallace_rca24_nand_23_9_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_10_y0(a_22, b_10, h_s_wallace_rca24_and_22_10_y0);
  fa fa_h_s_wallace_rca24_fa29_y2(h_s_wallace_rca24_fa28_y4, h_s_wallace_rca24_nand_23_9_y0, h_s_wallace_rca24_and_22_10_y0, h_s_wallace_rca24_fa29_y2, h_s_wallace_rca24_fa29_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_10_y0(a_23, b_10, h_s_wallace_rca24_nand_23_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_11_y0(a_22, b_11, h_s_wallace_rca24_and_22_11_y0);
  fa fa_h_s_wallace_rca24_fa30_y2(h_s_wallace_rca24_fa29_y4, h_s_wallace_rca24_nand_23_10_y0, h_s_wallace_rca24_and_22_11_y0, h_s_wallace_rca24_fa30_y2, h_s_wallace_rca24_fa30_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_11_y0(a_23, b_11, h_s_wallace_rca24_nand_23_11_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_12_y0(a_22, b_12, h_s_wallace_rca24_and_22_12_y0);
  fa fa_h_s_wallace_rca24_fa31_y2(h_s_wallace_rca24_fa30_y4, h_s_wallace_rca24_nand_23_11_y0, h_s_wallace_rca24_and_22_12_y0, h_s_wallace_rca24_fa31_y2, h_s_wallace_rca24_fa31_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_12_y0(a_23, b_12, h_s_wallace_rca24_nand_23_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_13_y0(a_22, b_13, h_s_wallace_rca24_and_22_13_y0);
  fa fa_h_s_wallace_rca24_fa32_y2(h_s_wallace_rca24_fa31_y4, h_s_wallace_rca24_nand_23_12_y0, h_s_wallace_rca24_and_22_13_y0, h_s_wallace_rca24_fa32_y2, h_s_wallace_rca24_fa32_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_13_y0(a_23, b_13, h_s_wallace_rca24_nand_23_13_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_14_y0(a_22, b_14, h_s_wallace_rca24_and_22_14_y0);
  fa fa_h_s_wallace_rca24_fa33_y2(h_s_wallace_rca24_fa32_y4, h_s_wallace_rca24_nand_23_13_y0, h_s_wallace_rca24_and_22_14_y0, h_s_wallace_rca24_fa33_y2, h_s_wallace_rca24_fa33_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_14_y0(a_23, b_14, h_s_wallace_rca24_nand_23_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_15_y0(a_22, b_15, h_s_wallace_rca24_and_22_15_y0);
  fa fa_h_s_wallace_rca24_fa34_y2(h_s_wallace_rca24_fa33_y4, h_s_wallace_rca24_nand_23_14_y0, h_s_wallace_rca24_and_22_15_y0, h_s_wallace_rca24_fa34_y2, h_s_wallace_rca24_fa34_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_15_y0(a_23, b_15, h_s_wallace_rca24_nand_23_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_16_y0(a_22, b_16, h_s_wallace_rca24_and_22_16_y0);
  fa fa_h_s_wallace_rca24_fa35_y2(h_s_wallace_rca24_fa34_y4, h_s_wallace_rca24_nand_23_15_y0, h_s_wallace_rca24_and_22_16_y0, h_s_wallace_rca24_fa35_y2, h_s_wallace_rca24_fa35_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_16_y0(a_23, b_16, h_s_wallace_rca24_nand_23_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_17_y0(a_22, b_17, h_s_wallace_rca24_and_22_17_y0);
  fa fa_h_s_wallace_rca24_fa36_y2(h_s_wallace_rca24_fa35_y4, h_s_wallace_rca24_nand_23_16_y0, h_s_wallace_rca24_and_22_17_y0, h_s_wallace_rca24_fa36_y2, h_s_wallace_rca24_fa36_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_17_y0(a_23, b_17, h_s_wallace_rca24_nand_23_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_18_y0(a_22, b_18, h_s_wallace_rca24_and_22_18_y0);
  fa fa_h_s_wallace_rca24_fa37_y2(h_s_wallace_rca24_fa36_y4, h_s_wallace_rca24_nand_23_17_y0, h_s_wallace_rca24_and_22_18_y0, h_s_wallace_rca24_fa37_y2, h_s_wallace_rca24_fa37_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_18_y0(a_23, b_18, h_s_wallace_rca24_nand_23_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_19_y0(a_22, b_19, h_s_wallace_rca24_and_22_19_y0);
  fa fa_h_s_wallace_rca24_fa38_y2(h_s_wallace_rca24_fa37_y4, h_s_wallace_rca24_nand_23_18_y0, h_s_wallace_rca24_and_22_19_y0, h_s_wallace_rca24_fa38_y2, h_s_wallace_rca24_fa38_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_19_y0(a_23, b_19, h_s_wallace_rca24_nand_23_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_20_y0(a_22, b_20, h_s_wallace_rca24_and_22_20_y0);
  fa fa_h_s_wallace_rca24_fa39_y2(h_s_wallace_rca24_fa38_y4, h_s_wallace_rca24_nand_23_19_y0, h_s_wallace_rca24_and_22_20_y0, h_s_wallace_rca24_fa39_y2, h_s_wallace_rca24_fa39_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_20_y0(a_23, b_20, h_s_wallace_rca24_nand_23_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_21_y0(a_22, b_21, h_s_wallace_rca24_and_22_21_y0);
  fa fa_h_s_wallace_rca24_fa40_y2(h_s_wallace_rca24_fa39_y4, h_s_wallace_rca24_nand_23_20_y0, h_s_wallace_rca24_and_22_21_y0, h_s_wallace_rca24_fa40_y2, h_s_wallace_rca24_fa40_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_21_y0(a_23, b_21, h_s_wallace_rca24_nand_23_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_22_22_y0(a_22, b_22, h_s_wallace_rca24_and_22_22_y0);
  fa fa_h_s_wallace_rca24_fa41_y2(h_s_wallace_rca24_fa40_y4, h_s_wallace_rca24_nand_23_21_y0, h_s_wallace_rca24_and_22_22_y0, h_s_wallace_rca24_fa41_y2, h_s_wallace_rca24_fa41_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_2_y0(a_1, b_2, h_s_wallace_rca24_and_1_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_3_y0(a_0, b_3, h_s_wallace_rca24_and_0_3_y0);
  ha ha_h_s_wallace_rca24_ha1_y0(h_s_wallace_rca24_and_1_2_y0, h_s_wallace_rca24_and_0_3_y0, h_s_wallace_rca24_ha1_y0, h_s_wallace_rca24_ha1_y1);
  and_gate and_gate_h_s_wallace_rca24_and_2_2_y0(a_2, b_2, h_s_wallace_rca24_and_2_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_3_y0(a_1, b_3, h_s_wallace_rca24_and_1_3_y0);
  fa fa_h_s_wallace_rca24_fa42_y2(h_s_wallace_rca24_ha1_y1, h_s_wallace_rca24_and_2_2_y0, h_s_wallace_rca24_and_1_3_y0, h_s_wallace_rca24_fa42_y2, h_s_wallace_rca24_fa42_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_2_y0(a_3, b_2, h_s_wallace_rca24_and_3_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_3_y0(a_2, b_3, h_s_wallace_rca24_and_2_3_y0);
  fa fa_h_s_wallace_rca24_fa43_y2(h_s_wallace_rca24_fa42_y4, h_s_wallace_rca24_and_3_2_y0, h_s_wallace_rca24_and_2_3_y0, h_s_wallace_rca24_fa43_y2, h_s_wallace_rca24_fa43_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_2_y0(a_4, b_2, h_s_wallace_rca24_and_4_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_3_y0(a_3, b_3, h_s_wallace_rca24_and_3_3_y0);
  fa fa_h_s_wallace_rca24_fa44_y2(h_s_wallace_rca24_fa43_y4, h_s_wallace_rca24_and_4_2_y0, h_s_wallace_rca24_and_3_3_y0, h_s_wallace_rca24_fa44_y2, h_s_wallace_rca24_fa44_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_2_y0(a_5, b_2, h_s_wallace_rca24_and_5_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_3_y0(a_4, b_3, h_s_wallace_rca24_and_4_3_y0);
  fa fa_h_s_wallace_rca24_fa45_y2(h_s_wallace_rca24_fa44_y4, h_s_wallace_rca24_and_5_2_y0, h_s_wallace_rca24_and_4_3_y0, h_s_wallace_rca24_fa45_y2, h_s_wallace_rca24_fa45_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_2_y0(a_6, b_2, h_s_wallace_rca24_and_6_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_3_y0(a_5, b_3, h_s_wallace_rca24_and_5_3_y0);
  fa fa_h_s_wallace_rca24_fa46_y2(h_s_wallace_rca24_fa45_y4, h_s_wallace_rca24_and_6_2_y0, h_s_wallace_rca24_and_5_3_y0, h_s_wallace_rca24_fa46_y2, h_s_wallace_rca24_fa46_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_2_y0(a_7, b_2, h_s_wallace_rca24_and_7_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_3_y0(a_6, b_3, h_s_wallace_rca24_and_6_3_y0);
  fa fa_h_s_wallace_rca24_fa47_y2(h_s_wallace_rca24_fa46_y4, h_s_wallace_rca24_and_7_2_y0, h_s_wallace_rca24_and_6_3_y0, h_s_wallace_rca24_fa47_y2, h_s_wallace_rca24_fa47_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_2_y0(a_8, b_2, h_s_wallace_rca24_and_8_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_3_y0(a_7, b_3, h_s_wallace_rca24_and_7_3_y0);
  fa fa_h_s_wallace_rca24_fa48_y2(h_s_wallace_rca24_fa47_y4, h_s_wallace_rca24_and_8_2_y0, h_s_wallace_rca24_and_7_3_y0, h_s_wallace_rca24_fa48_y2, h_s_wallace_rca24_fa48_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_2_y0(a_9, b_2, h_s_wallace_rca24_and_9_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_3_y0(a_8, b_3, h_s_wallace_rca24_and_8_3_y0);
  fa fa_h_s_wallace_rca24_fa49_y2(h_s_wallace_rca24_fa48_y4, h_s_wallace_rca24_and_9_2_y0, h_s_wallace_rca24_and_8_3_y0, h_s_wallace_rca24_fa49_y2, h_s_wallace_rca24_fa49_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_2_y0(a_10, b_2, h_s_wallace_rca24_and_10_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_3_y0(a_9, b_3, h_s_wallace_rca24_and_9_3_y0);
  fa fa_h_s_wallace_rca24_fa50_y2(h_s_wallace_rca24_fa49_y4, h_s_wallace_rca24_and_10_2_y0, h_s_wallace_rca24_and_9_3_y0, h_s_wallace_rca24_fa50_y2, h_s_wallace_rca24_fa50_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_2_y0(a_11, b_2, h_s_wallace_rca24_and_11_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_3_y0(a_10, b_3, h_s_wallace_rca24_and_10_3_y0);
  fa fa_h_s_wallace_rca24_fa51_y2(h_s_wallace_rca24_fa50_y4, h_s_wallace_rca24_and_11_2_y0, h_s_wallace_rca24_and_10_3_y0, h_s_wallace_rca24_fa51_y2, h_s_wallace_rca24_fa51_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_2_y0(a_12, b_2, h_s_wallace_rca24_and_12_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_3_y0(a_11, b_3, h_s_wallace_rca24_and_11_3_y0);
  fa fa_h_s_wallace_rca24_fa52_y2(h_s_wallace_rca24_fa51_y4, h_s_wallace_rca24_and_12_2_y0, h_s_wallace_rca24_and_11_3_y0, h_s_wallace_rca24_fa52_y2, h_s_wallace_rca24_fa52_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_2_y0(a_13, b_2, h_s_wallace_rca24_and_13_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_3_y0(a_12, b_3, h_s_wallace_rca24_and_12_3_y0);
  fa fa_h_s_wallace_rca24_fa53_y2(h_s_wallace_rca24_fa52_y4, h_s_wallace_rca24_and_13_2_y0, h_s_wallace_rca24_and_12_3_y0, h_s_wallace_rca24_fa53_y2, h_s_wallace_rca24_fa53_y4);
  and_gate and_gate_h_s_wallace_rca24_and_14_2_y0(a_14, b_2, h_s_wallace_rca24_and_14_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_13_3_y0(a_13, b_3, h_s_wallace_rca24_and_13_3_y0);
  fa fa_h_s_wallace_rca24_fa54_y2(h_s_wallace_rca24_fa53_y4, h_s_wallace_rca24_and_14_2_y0, h_s_wallace_rca24_and_13_3_y0, h_s_wallace_rca24_fa54_y2, h_s_wallace_rca24_fa54_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_2_y0(a_15, b_2, h_s_wallace_rca24_and_15_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_3_y0(a_14, b_3, h_s_wallace_rca24_and_14_3_y0);
  fa fa_h_s_wallace_rca24_fa55_y2(h_s_wallace_rca24_fa54_y4, h_s_wallace_rca24_and_15_2_y0, h_s_wallace_rca24_and_14_3_y0, h_s_wallace_rca24_fa55_y2, h_s_wallace_rca24_fa55_y4);
  and_gate and_gate_h_s_wallace_rca24_and_16_2_y0(a_16, b_2, h_s_wallace_rca24_and_16_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_15_3_y0(a_15, b_3, h_s_wallace_rca24_and_15_3_y0);
  fa fa_h_s_wallace_rca24_fa56_y2(h_s_wallace_rca24_fa55_y4, h_s_wallace_rca24_and_16_2_y0, h_s_wallace_rca24_and_15_3_y0, h_s_wallace_rca24_fa56_y2, h_s_wallace_rca24_fa56_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_2_y0(a_17, b_2, h_s_wallace_rca24_and_17_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_3_y0(a_16, b_3, h_s_wallace_rca24_and_16_3_y0);
  fa fa_h_s_wallace_rca24_fa57_y2(h_s_wallace_rca24_fa56_y4, h_s_wallace_rca24_and_17_2_y0, h_s_wallace_rca24_and_16_3_y0, h_s_wallace_rca24_fa57_y2, h_s_wallace_rca24_fa57_y4);
  and_gate and_gate_h_s_wallace_rca24_and_18_2_y0(a_18, b_2, h_s_wallace_rca24_and_18_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_17_3_y0(a_17, b_3, h_s_wallace_rca24_and_17_3_y0);
  fa fa_h_s_wallace_rca24_fa58_y2(h_s_wallace_rca24_fa57_y4, h_s_wallace_rca24_and_18_2_y0, h_s_wallace_rca24_and_17_3_y0, h_s_wallace_rca24_fa58_y2, h_s_wallace_rca24_fa58_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_2_y0(a_19, b_2, h_s_wallace_rca24_and_19_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_3_y0(a_18, b_3, h_s_wallace_rca24_and_18_3_y0);
  fa fa_h_s_wallace_rca24_fa59_y2(h_s_wallace_rca24_fa58_y4, h_s_wallace_rca24_and_19_2_y0, h_s_wallace_rca24_and_18_3_y0, h_s_wallace_rca24_fa59_y2, h_s_wallace_rca24_fa59_y4);
  and_gate and_gate_h_s_wallace_rca24_and_20_2_y0(a_20, b_2, h_s_wallace_rca24_and_20_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_19_3_y0(a_19, b_3, h_s_wallace_rca24_and_19_3_y0);
  fa fa_h_s_wallace_rca24_fa60_y2(h_s_wallace_rca24_fa59_y4, h_s_wallace_rca24_and_20_2_y0, h_s_wallace_rca24_and_19_3_y0, h_s_wallace_rca24_fa60_y2, h_s_wallace_rca24_fa60_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_2_y0(a_21, b_2, h_s_wallace_rca24_and_21_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_3_y0(a_20, b_3, h_s_wallace_rca24_and_20_3_y0);
  fa fa_h_s_wallace_rca24_fa61_y2(h_s_wallace_rca24_fa60_y4, h_s_wallace_rca24_and_21_2_y0, h_s_wallace_rca24_and_20_3_y0, h_s_wallace_rca24_fa61_y2, h_s_wallace_rca24_fa61_y4);
  and_gate and_gate_h_s_wallace_rca24_and_22_2_y0(a_22, b_2, h_s_wallace_rca24_and_22_2_y0);
  and_gate and_gate_h_s_wallace_rca24_and_21_3_y0(a_21, b_3, h_s_wallace_rca24_and_21_3_y0);
  fa fa_h_s_wallace_rca24_fa62_y2(h_s_wallace_rca24_fa61_y4, h_s_wallace_rca24_and_22_2_y0, h_s_wallace_rca24_and_21_3_y0, h_s_wallace_rca24_fa62_y2, h_s_wallace_rca24_fa62_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_4_y0(a_21, b_4, h_s_wallace_rca24_and_21_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_5_y0(a_20, b_5, h_s_wallace_rca24_and_20_5_y0);
  fa fa_h_s_wallace_rca24_fa63_y2(h_s_wallace_rca24_fa62_y4, h_s_wallace_rca24_and_21_4_y0, h_s_wallace_rca24_and_20_5_y0, h_s_wallace_rca24_fa63_y2, h_s_wallace_rca24_fa63_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_5_y0(a_21, b_5, h_s_wallace_rca24_and_21_5_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_6_y0(a_20, b_6, h_s_wallace_rca24_and_20_6_y0);
  fa fa_h_s_wallace_rca24_fa64_y2(h_s_wallace_rca24_fa63_y4, h_s_wallace_rca24_and_21_5_y0, h_s_wallace_rca24_and_20_6_y0, h_s_wallace_rca24_fa64_y2, h_s_wallace_rca24_fa64_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_6_y0(a_21, b_6, h_s_wallace_rca24_and_21_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_7_y0(a_20, b_7, h_s_wallace_rca24_and_20_7_y0);
  fa fa_h_s_wallace_rca24_fa65_y2(h_s_wallace_rca24_fa64_y4, h_s_wallace_rca24_and_21_6_y0, h_s_wallace_rca24_and_20_7_y0, h_s_wallace_rca24_fa65_y2, h_s_wallace_rca24_fa65_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_7_y0(a_21, b_7, h_s_wallace_rca24_and_21_7_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_8_y0(a_20, b_8, h_s_wallace_rca24_and_20_8_y0);
  fa fa_h_s_wallace_rca24_fa66_y2(h_s_wallace_rca24_fa65_y4, h_s_wallace_rca24_and_21_7_y0, h_s_wallace_rca24_and_20_8_y0, h_s_wallace_rca24_fa66_y2, h_s_wallace_rca24_fa66_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_8_y0(a_21, b_8, h_s_wallace_rca24_and_21_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_9_y0(a_20, b_9, h_s_wallace_rca24_and_20_9_y0);
  fa fa_h_s_wallace_rca24_fa67_y2(h_s_wallace_rca24_fa66_y4, h_s_wallace_rca24_and_21_8_y0, h_s_wallace_rca24_and_20_9_y0, h_s_wallace_rca24_fa67_y2, h_s_wallace_rca24_fa67_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_9_y0(a_21, b_9, h_s_wallace_rca24_and_21_9_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_10_y0(a_20, b_10, h_s_wallace_rca24_and_20_10_y0);
  fa fa_h_s_wallace_rca24_fa68_y2(h_s_wallace_rca24_fa67_y4, h_s_wallace_rca24_and_21_9_y0, h_s_wallace_rca24_and_20_10_y0, h_s_wallace_rca24_fa68_y2, h_s_wallace_rca24_fa68_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_10_y0(a_21, b_10, h_s_wallace_rca24_and_21_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_11_y0(a_20, b_11, h_s_wallace_rca24_and_20_11_y0);
  fa fa_h_s_wallace_rca24_fa69_y2(h_s_wallace_rca24_fa68_y4, h_s_wallace_rca24_and_21_10_y0, h_s_wallace_rca24_and_20_11_y0, h_s_wallace_rca24_fa69_y2, h_s_wallace_rca24_fa69_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_11_y0(a_21, b_11, h_s_wallace_rca24_and_21_11_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_12_y0(a_20, b_12, h_s_wallace_rca24_and_20_12_y0);
  fa fa_h_s_wallace_rca24_fa70_y2(h_s_wallace_rca24_fa69_y4, h_s_wallace_rca24_and_21_11_y0, h_s_wallace_rca24_and_20_12_y0, h_s_wallace_rca24_fa70_y2, h_s_wallace_rca24_fa70_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_12_y0(a_21, b_12, h_s_wallace_rca24_and_21_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_13_y0(a_20, b_13, h_s_wallace_rca24_and_20_13_y0);
  fa fa_h_s_wallace_rca24_fa71_y2(h_s_wallace_rca24_fa70_y4, h_s_wallace_rca24_and_21_12_y0, h_s_wallace_rca24_and_20_13_y0, h_s_wallace_rca24_fa71_y2, h_s_wallace_rca24_fa71_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_13_y0(a_21, b_13, h_s_wallace_rca24_and_21_13_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_14_y0(a_20, b_14, h_s_wallace_rca24_and_20_14_y0);
  fa fa_h_s_wallace_rca24_fa72_y2(h_s_wallace_rca24_fa71_y4, h_s_wallace_rca24_and_21_13_y0, h_s_wallace_rca24_and_20_14_y0, h_s_wallace_rca24_fa72_y2, h_s_wallace_rca24_fa72_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_14_y0(a_21, b_14, h_s_wallace_rca24_and_21_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_15_y0(a_20, b_15, h_s_wallace_rca24_and_20_15_y0);
  fa fa_h_s_wallace_rca24_fa73_y2(h_s_wallace_rca24_fa72_y4, h_s_wallace_rca24_and_21_14_y0, h_s_wallace_rca24_and_20_15_y0, h_s_wallace_rca24_fa73_y2, h_s_wallace_rca24_fa73_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_15_y0(a_21, b_15, h_s_wallace_rca24_and_21_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_16_y0(a_20, b_16, h_s_wallace_rca24_and_20_16_y0);
  fa fa_h_s_wallace_rca24_fa74_y2(h_s_wallace_rca24_fa73_y4, h_s_wallace_rca24_and_21_15_y0, h_s_wallace_rca24_and_20_16_y0, h_s_wallace_rca24_fa74_y2, h_s_wallace_rca24_fa74_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_16_y0(a_21, b_16, h_s_wallace_rca24_and_21_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_17_y0(a_20, b_17, h_s_wallace_rca24_and_20_17_y0);
  fa fa_h_s_wallace_rca24_fa75_y2(h_s_wallace_rca24_fa74_y4, h_s_wallace_rca24_and_21_16_y0, h_s_wallace_rca24_and_20_17_y0, h_s_wallace_rca24_fa75_y2, h_s_wallace_rca24_fa75_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_17_y0(a_21, b_17, h_s_wallace_rca24_and_21_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_18_y0(a_20, b_18, h_s_wallace_rca24_and_20_18_y0);
  fa fa_h_s_wallace_rca24_fa76_y2(h_s_wallace_rca24_fa75_y4, h_s_wallace_rca24_and_21_17_y0, h_s_wallace_rca24_and_20_18_y0, h_s_wallace_rca24_fa76_y2, h_s_wallace_rca24_fa76_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_18_y0(a_21, b_18, h_s_wallace_rca24_and_21_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_19_y0(a_20, b_19, h_s_wallace_rca24_and_20_19_y0);
  fa fa_h_s_wallace_rca24_fa77_y2(h_s_wallace_rca24_fa76_y4, h_s_wallace_rca24_and_21_18_y0, h_s_wallace_rca24_and_20_19_y0, h_s_wallace_rca24_fa77_y2, h_s_wallace_rca24_fa77_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_19_y0(a_21, b_19, h_s_wallace_rca24_and_21_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_20_y0(a_20, b_20, h_s_wallace_rca24_and_20_20_y0);
  fa fa_h_s_wallace_rca24_fa78_y2(h_s_wallace_rca24_fa77_y4, h_s_wallace_rca24_and_21_19_y0, h_s_wallace_rca24_and_20_20_y0, h_s_wallace_rca24_fa78_y2, h_s_wallace_rca24_fa78_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_20_y0(a_21, b_20, h_s_wallace_rca24_and_21_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_21_y0(a_20, b_21, h_s_wallace_rca24_and_20_21_y0);
  fa fa_h_s_wallace_rca24_fa79_y2(h_s_wallace_rca24_fa78_y4, h_s_wallace_rca24_and_21_20_y0, h_s_wallace_rca24_and_20_21_y0, h_s_wallace_rca24_fa79_y2, h_s_wallace_rca24_fa79_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_21_y0(a_21, b_21, h_s_wallace_rca24_and_21_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_20_22_y0(a_20, b_22, h_s_wallace_rca24_and_20_22_y0);
  fa fa_h_s_wallace_rca24_fa80_y2(h_s_wallace_rca24_fa79_y4, h_s_wallace_rca24_and_21_21_y0, h_s_wallace_rca24_and_20_22_y0, h_s_wallace_rca24_fa80_y2, h_s_wallace_rca24_fa80_y4);
  and_gate and_gate_h_s_wallace_rca24_and_21_22_y0(a_21, b_22, h_s_wallace_rca24_and_21_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_20_23_y0(a_20, b_23, h_s_wallace_rca24_nand_20_23_y0);
  fa fa_h_s_wallace_rca24_fa81_y2(h_s_wallace_rca24_fa80_y4, h_s_wallace_rca24_and_21_22_y0, h_s_wallace_rca24_nand_20_23_y0, h_s_wallace_rca24_fa81_y2, h_s_wallace_rca24_fa81_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_4_y0(a_0, b_4, h_s_wallace_rca24_and_0_4_y0);
  ha ha_h_s_wallace_rca24_ha2_y0(h_s_wallace_rca24_and_0_4_y0, h_s_wallace_rca24_fa1_y2, h_s_wallace_rca24_ha2_y0, h_s_wallace_rca24_ha2_y1);
  and_gate and_gate_h_s_wallace_rca24_and_1_4_y0(a_1, b_4, h_s_wallace_rca24_and_1_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_5_y0(a_0, b_5, h_s_wallace_rca24_and_0_5_y0);
  fa fa_h_s_wallace_rca24_fa82_y2(h_s_wallace_rca24_ha2_y1, h_s_wallace_rca24_and_1_4_y0, h_s_wallace_rca24_and_0_5_y0, h_s_wallace_rca24_fa82_y2, h_s_wallace_rca24_fa82_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_4_y0(a_2, b_4, h_s_wallace_rca24_and_2_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_5_y0(a_1, b_5, h_s_wallace_rca24_and_1_5_y0);
  fa fa_h_s_wallace_rca24_fa83_y2(h_s_wallace_rca24_fa82_y4, h_s_wallace_rca24_and_2_4_y0, h_s_wallace_rca24_and_1_5_y0, h_s_wallace_rca24_fa83_y2, h_s_wallace_rca24_fa83_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_4_y0(a_3, b_4, h_s_wallace_rca24_and_3_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_5_y0(a_2, b_5, h_s_wallace_rca24_and_2_5_y0);
  fa fa_h_s_wallace_rca24_fa84_y2(h_s_wallace_rca24_fa83_y4, h_s_wallace_rca24_and_3_4_y0, h_s_wallace_rca24_and_2_5_y0, h_s_wallace_rca24_fa84_y2, h_s_wallace_rca24_fa84_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_4_y0(a_4, b_4, h_s_wallace_rca24_and_4_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_5_y0(a_3, b_5, h_s_wallace_rca24_and_3_5_y0);
  fa fa_h_s_wallace_rca24_fa85_y2(h_s_wallace_rca24_fa84_y4, h_s_wallace_rca24_and_4_4_y0, h_s_wallace_rca24_and_3_5_y0, h_s_wallace_rca24_fa85_y2, h_s_wallace_rca24_fa85_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_4_y0(a_5, b_4, h_s_wallace_rca24_and_5_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_5_y0(a_4, b_5, h_s_wallace_rca24_and_4_5_y0);
  fa fa_h_s_wallace_rca24_fa86_y2(h_s_wallace_rca24_fa85_y4, h_s_wallace_rca24_and_5_4_y0, h_s_wallace_rca24_and_4_5_y0, h_s_wallace_rca24_fa86_y2, h_s_wallace_rca24_fa86_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_4_y0(a_6, b_4, h_s_wallace_rca24_and_6_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_5_y0(a_5, b_5, h_s_wallace_rca24_and_5_5_y0);
  fa fa_h_s_wallace_rca24_fa87_y2(h_s_wallace_rca24_fa86_y4, h_s_wallace_rca24_and_6_4_y0, h_s_wallace_rca24_and_5_5_y0, h_s_wallace_rca24_fa87_y2, h_s_wallace_rca24_fa87_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_4_y0(a_7, b_4, h_s_wallace_rca24_and_7_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_5_y0(a_6, b_5, h_s_wallace_rca24_and_6_5_y0);
  fa fa_h_s_wallace_rca24_fa88_y2(h_s_wallace_rca24_fa87_y4, h_s_wallace_rca24_and_7_4_y0, h_s_wallace_rca24_and_6_5_y0, h_s_wallace_rca24_fa88_y2, h_s_wallace_rca24_fa88_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_4_y0(a_8, b_4, h_s_wallace_rca24_and_8_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_5_y0(a_7, b_5, h_s_wallace_rca24_and_7_5_y0);
  fa fa_h_s_wallace_rca24_fa89_y2(h_s_wallace_rca24_fa88_y4, h_s_wallace_rca24_and_8_4_y0, h_s_wallace_rca24_and_7_5_y0, h_s_wallace_rca24_fa89_y2, h_s_wallace_rca24_fa89_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_4_y0(a_9, b_4, h_s_wallace_rca24_and_9_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_5_y0(a_8, b_5, h_s_wallace_rca24_and_8_5_y0);
  fa fa_h_s_wallace_rca24_fa90_y2(h_s_wallace_rca24_fa89_y4, h_s_wallace_rca24_and_9_4_y0, h_s_wallace_rca24_and_8_5_y0, h_s_wallace_rca24_fa90_y2, h_s_wallace_rca24_fa90_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_4_y0(a_10, b_4, h_s_wallace_rca24_and_10_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_5_y0(a_9, b_5, h_s_wallace_rca24_and_9_5_y0);
  fa fa_h_s_wallace_rca24_fa91_y2(h_s_wallace_rca24_fa90_y4, h_s_wallace_rca24_and_10_4_y0, h_s_wallace_rca24_and_9_5_y0, h_s_wallace_rca24_fa91_y2, h_s_wallace_rca24_fa91_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_4_y0(a_11, b_4, h_s_wallace_rca24_and_11_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_5_y0(a_10, b_5, h_s_wallace_rca24_and_10_5_y0);
  fa fa_h_s_wallace_rca24_fa92_y2(h_s_wallace_rca24_fa91_y4, h_s_wallace_rca24_and_11_4_y0, h_s_wallace_rca24_and_10_5_y0, h_s_wallace_rca24_fa92_y2, h_s_wallace_rca24_fa92_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_4_y0(a_12, b_4, h_s_wallace_rca24_and_12_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_5_y0(a_11, b_5, h_s_wallace_rca24_and_11_5_y0);
  fa fa_h_s_wallace_rca24_fa93_y2(h_s_wallace_rca24_fa92_y4, h_s_wallace_rca24_and_12_4_y0, h_s_wallace_rca24_and_11_5_y0, h_s_wallace_rca24_fa93_y2, h_s_wallace_rca24_fa93_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_4_y0(a_13, b_4, h_s_wallace_rca24_and_13_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_5_y0(a_12, b_5, h_s_wallace_rca24_and_12_5_y0);
  fa fa_h_s_wallace_rca24_fa94_y2(h_s_wallace_rca24_fa93_y4, h_s_wallace_rca24_and_13_4_y0, h_s_wallace_rca24_and_12_5_y0, h_s_wallace_rca24_fa94_y2, h_s_wallace_rca24_fa94_y4);
  and_gate and_gate_h_s_wallace_rca24_and_14_4_y0(a_14, b_4, h_s_wallace_rca24_and_14_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_13_5_y0(a_13, b_5, h_s_wallace_rca24_and_13_5_y0);
  fa fa_h_s_wallace_rca24_fa95_y2(h_s_wallace_rca24_fa94_y4, h_s_wallace_rca24_and_14_4_y0, h_s_wallace_rca24_and_13_5_y0, h_s_wallace_rca24_fa95_y2, h_s_wallace_rca24_fa95_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_4_y0(a_15, b_4, h_s_wallace_rca24_and_15_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_5_y0(a_14, b_5, h_s_wallace_rca24_and_14_5_y0);
  fa fa_h_s_wallace_rca24_fa96_y2(h_s_wallace_rca24_fa95_y4, h_s_wallace_rca24_and_15_4_y0, h_s_wallace_rca24_and_14_5_y0, h_s_wallace_rca24_fa96_y2, h_s_wallace_rca24_fa96_y4);
  and_gate and_gate_h_s_wallace_rca24_and_16_4_y0(a_16, b_4, h_s_wallace_rca24_and_16_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_15_5_y0(a_15, b_5, h_s_wallace_rca24_and_15_5_y0);
  fa fa_h_s_wallace_rca24_fa97_y2(h_s_wallace_rca24_fa96_y4, h_s_wallace_rca24_and_16_4_y0, h_s_wallace_rca24_and_15_5_y0, h_s_wallace_rca24_fa97_y2, h_s_wallace_rca24_fa97_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_4_y0(a_17, b_4, h_s_wallace_rca24_and_17_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_5_y0(a_16, b_5, h_s_wallace_rca24_and_16_5_y0);
  fa fa_h_s_wallace_rca24_fa98_y2(h_s_wallace_rca24_fa97_y4, h_s_wallace_rca24_and_17_4_y0, h_s_wallace_rca24_and_16_5_y0, h_s_wallace_rca24_fa98_y2, h_s_wallace_rca24_fa98_y4);
  and_gate and_gate_h_s_wallace_rca24_and_18_4_y0(a_18, b_4, h_s_wallace_rca24_and_18_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_17_5_y0(a_17, b_5, h_s_wallace_rca24_and_17_5_y0);
  fa fa_h_s_wallace_rca24_fa99_y2(h_s_wallace_rca24_fa98_y4, h_s_wallace_rca24_and_18_4_y0, h_s_wallace_rca24_and_17_5_y0, h_s_wallace_rca24_fa99_y2, h_s_wallace_rca24_fa99_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_4_y0(a_19, b_4, h_s_wallace_rca24_and_19_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_5_y0(a_18, b_5, h_s_wallace_rca24_and_18_5_y0);
  fa fa_h_s_wallace_rca24_fa100_y2(h_s_wallace_rca24_fa99_y4, h_s_wallace_rca24_and_19_4_y0, h_s_wallace_rca24_and_18_5_y0, h_s_wallace_rca24_fa100_y2, h_s_wallace_rca24_fa100_y4);
  and_gate and_gate_h_s_wallace_rca24_and_20_4_y0(a_20, b_4, h_s_wallace_rca24_and_20_4_y0);
  and_gate and_gate_h_s_wallace_rca24_and_19_5_y0(a_19, b_5, h_s_wallace_rca24_and_19_5_y0);
  fa fa_h_s_wallace_rca24_fa101_y2(h_s_wallace_rca24_fa100_y4, h_s_wallace_rca24_and_20_4_y0, h_s_wallace_rca24_and_19_5_y0, h_s_wallace_rca24_fa101_y2, h_s_wallace_rca24_fa101_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_6_y0(a_19, b_6, h_s_wallace_rca24_and_19_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_7_y0(a_18, b_7, h_s_wallace_rca24_and_18_7_y0);
  fa fa_h_s_wallace_rca24_fa102_y2(h_s_wallace_rca24_fa101_y4, h_s_wallace_rca24_and_19_6_y0, h_s_wallace_rca24_and_18_7_y0, h_s_wallace_rca24_fa102_y2, h_s_wallace_rca24_fa102_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_7_y0(a_19, b_7, h_s_wallace_rca24_and_19_7_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_8_y0(a_18, b_8, h_s_wallace_rca24_and_18_8_y0);
  fa fa_h_s_wallace_rca24_fa103_y2(h_s_wallace_rca24_fa102_y4, h_s_wallace_rca24_and_19_7_y0, h_s_wallace_rca24_and_18_8_y0, h_s_wallace_rca24_fa103_y2, h_s_wallace_rca24_fa103_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_8_y0(a_19, b_8, h_s_wallace_rca24_and_19_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_9_y0(a_18, b_9, h_s_wallace_rca24_and_18_9_y0);
  fa fa_h_s_wallace_rca24_fa104_y2(h_s_wallace_rca24_fa103_y4, h_s_wallace_rca24_and_19_8_y0, h_s_wallace_rca24_and_18_9_y0, h_s_wallace_rca24_fa104_y2, h_s_wallace_rca24_fa104_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_9_y0(a_19, b_9, h_s_wallace_rca24_and_19_9_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_10_y0(a_18, b_10, h_s_wallace_rca24_and_18_10_y0);
  fa fa_h_s_wallace_rca24_fa105_y2(h_s_wallace_rca24_fa104_y4, h_s_wallace_rca24_and_19_9_y0, h_s_wallace_rca24_and_18_10_y0, h_s_wallace_rca24_fa105_y2, h_s_wallace_rca24_fa105_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_10_y0(a_19, b_10, h_s_wallace_rca24_and_19_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_11_y0(a_18, b_11, h_s_wallace_rca24_and_18_11_y0);
  fa fa_h_s_wallace_rca24_fa106_y2(h_s_wallace_rca24_fa105_y4, h_s_wallace_rca24_and_19_10_y0, h_s_wallace_rca24_and_18_11_y0, h_s_wallace_rca24_fa106_y2, h_s_wallace_rca24_fa106_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_11_y0(a_19, b_11, h_s_wallace_rca24_and_19_11_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_12_y0(a_18, b_12, h_s_wallace_rca24_and_18_12_y0);
  fa fa_h_s_wallace_rca24_fa107_y2(h_s_wallace_rca24_fa106_y4, h_s_wallace_rca24_and_19_11_y0, h_s_wallace_rca24_and_18_12_y0, h_s_wallace_rca24_fa107_y2, h_s_wallace_rca24_fa107_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_12_y0(a_19, b_12, h_s_wallace_rca24_and_19_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_13_y0(a_18, b_13, h_s_wallace_rca24_and_18_13_y0);
  fa fa_h_s_wallace_rca24_fa108_y2(h_s_wallace_rca24_fa107_y4, h_s_wallace_rca24_and_19_12_y0, h_s_wallace_rca24_and_18_13_y0, h_s_wallace_rca24_fa108_y2, h_s_wallace_rca24_fa108_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_13_y0(a_19, b_13, h_s_wallace_rca24_and_19_13_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_14_y0(a_18, b_14, h_s_wallace_rca24_and_18_14_y0);
  fa fa_h_s_wallace_rca24_fa109_y2(h_s_wallace_rca24_fa108_y4, h_s_wallace_rca24_and_19_13_y0, h_s_wallace_rca24_and_18_14_y0, h_s_wallace_rca24_fa109_y2, h_s_wallace_rca24_fa109_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_14_y0(a_19, b_14, h_s_wallace_rca24_and_19_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_15_y0(a_18, b_15, h_s_wallace_rca24_and_18_15_y0);
  fa fa_h_s_wallace_rca24_fa110_y2(h_s_wallace_rca24_fa109_y4, h_s_wallace_rca24_and_19_14_y0, h_s_wallace_rca24_and_18_15_y0, h_s_wallace_rca24_fa110_y2, h_s_wallace_rca24_fa110_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_15_y0(a_19, b_15, h_s_wallace_rca24_and_19_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_16_y0(a_18, b_16, h_s_wallace_rca24_and_18_16_y0);
  fa fa_h_s_wallace_rca24_fa111_y2(h_s_wallace_rca24_fa110_y4, h_s_wallace_rca24_and_19_15_y0, h_s_wallace_rca24_and_18_16_y0, h_s_wallace_rca24_fa111_y2, h_s_wallace_rca24_fa111_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_16_y0(a_19, b_16, h_s_wallace_rca24_and_19_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_17_y0(a_18, b_17, h_s_wallace_rca24_and_18_17_y0);
  fa fa_h_s_wallace_rca24_fa112_y2(h_s_wallace_rca24_fa111_y4, h_s_wallace_rca24_and_19_16_y0, h_s_wallace_rca24_and_18_17_y0, h_s_wallace_rca24_fa112_y2, h_s_wallace_rca24_fa112_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_17_y0(a_19, b_17, h_s_wallace_rca24_and_19_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_18_y0(a_18, b_18, h_s_wallace_rca24_and_18_18_y0);
  fa fa_h_s_wallace_rca24_fa113_y2(h_s_wallace_rca24_fa112_y4, h_s_wallace_rca24_and_19_17_y0, h_s_wallace_rca24_and_18_18_y0, h_s_wallace_rca24_fa113_y2, h_s_wallace_rca24_fa113_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_18_y0(a_19, b_18, h_s_wallace_rca24_and_19_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_19_y0(a_18, b_19, h_s_wallace_rca24_and_18_19_y0);
  fa fa_h_s_wallace_rca24_fa114_y2(h_s_wallace_rca24_fa113_y4, h_s_wallace_rca24_and_19_18_y0, h_s_wallace_rca24_and_18_19_y0, h_s_wallace_rca24_fa114_y2, h_s_wallace_rca24_fa114_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_19_y0(a_19, b_19, h_s_wallace_rca24_and_19_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_20_y0(a_18, b_20, h_s_wallace_rca24_and_18_20_y0);
  fa fa_h_s_wallace_rca24_fa115_y2(h_s_wallace_rca24_fa114_y4, h_s_wallace_rca24_and_19_19_y0, h_s_wallace_rca24_and_18_20_y0, h_s_wallace_rca24_fa115_y2, h_s_wallace_rca24_fa115_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_20_y0(a_19, b_20, h_s_wallace_rca24_and_19_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_21_y0(a_18, b_21, h_s_wallace_rca24_and_18_21_y0);
  fa fa_h_s_wallace_rca24_fa116_y2(h_s_wallace_rca24_fa115_y4, h_s_wallace_rca24_and_19_20_y0, h_s_wallace_rca24_and_18_21_y0, h_s_wallace_rca24_fa116_y2, h_s_wallace_rca24_fa116_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_21_y0(a_19, b_21, h_s_wallace_rca24_and_19_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_18_22_y0(a_18, b_22, h_s_wallace_rca24_and_18_22_y0);
  fa fa_h_s_wallace_rca24_fa117_y2(h_s_wallace_rca24_fa116_y4, h_s_wallace_rca24_and_19_21_y0, h_s_wallace_rca24_and_18_22_y0, h_s_wallace_rca24_fa117_y2, h_s_wallace_rca24_fa117_y4);
  and_gate and_gate_h_s_wallace_rca24_and_19_22_y0(a_19, b_22, h_s_wallace_rca24_and_19_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_18_23_y0(a_18, b_23, h_s_wallace_rca24_nand_18_23_y0);
  fa fa_h_s_wallace_rca24_fa118_y2(h_s_wallace_rca24_fa117_y4, h_s_wallace_rca24_and_19_22_y0, h_s_wallace_rca24_nand_18_23_y0, h_s_wallace_rca24_fa118_y2, h_s_wallace_rca24_fa118_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_19_23_y0(a_19, b_23, h_s_wallace_rca24_nand_19_23_y0);
  fa fa_h_s_wallace_rca24_fa119_y2(h_s_wallace_rca24_fa118_y4, h_s_wallace_rca24_nand_19_23_y0, h_s_wallace_rca24_fa39_y2, h_s_wallace_rca24_fa119_y2, h_s_wallace_rca24_fa119_y4);
  ha ha_h_s_wallace_rca24_ha3_y0(h_s_wallace_rca24_fa2_y2, h_s_wallace_rca24_fa43_y2, h_s_wallace_rca24_ha3_y0, h_s_wallace_rca24_ha3_y1);
  and_gate and_gate_h_s_wallace_rca24_and_0_6_y0(a_0, b_6, h_s_wallace_rca24_and_0_6_y0);
  fa fa_h_s_wallace_rca24_fa120_y2(h_s_wallace_rca24_ha3_y1, h_s_wallace_rca24_and_0_6_y0, h_s_wallace_rca24_fa3_y2, h_s_wallace_rca24_fa120_y2, h_s_wallace_rca24_fa120_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_6_y0(a_1, b_6, h_s_wallace_rca24_and_1_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_7_y0(a_0, b_7, h_s_wallace_rca24_and_0_7_y0);
  fa fa_h_s_wallace_rca24_fa121_y2(h_s_wallace_rca24_fa120_y4, h_s_wallace_rca24_and_1_6_y0, h_s_wallace_rca24_and_0_7_y0, h_s_wallace_rca24_fa121_y2, h_s_wallace_rca24_fa121_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_6_y0(a_2, b_6, h_s_wallace_rca24_and_2_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_7_y0(a_1, b_7, h_s_wallace_rca24_and_1_7_y0);
  fa fa_h_s_wallace_rca24_fa122_y2(h_s_wallace_rca24_fa121_y4, h_s_wallace_rca24_and_2_6_y0, h_s_wallace_rca24_and_1_7_y0, h_s_wallace_rca24_fa122_y2, h_s_wallace_rca24_fa122_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_6_y0(a_3, b_6, h_s_wallace_rca24_and_3_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_7_y0(a_2, b_7, h_s_wallace_rca24_and_2_7_y0);
  fa fa_h_s_wallace_rca24_fa123_y2(h_s_wallace_rca24_fa122_y4, h_s_wallace_rca24_and_3_6_y0, h_s_wallace_rca24_and_2_7_y0, h_s_wallace_rca24_fa123_y2, h_s_wallace_rca24_fa123_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_6_y0(a_4, b_6, h_s_wallace_rca24_and_4_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_7_y0(a_3, b_7, h_s_wallace_rca24_and_3_7_y0);
  fa fa_h_s_wallace_rca24_fa124_y2(h_s_wallace_rca24_fa123_y4, h_s_wallace_rca24_and_4_6_y0, h_s_wallace_rca24_and_3_7_y0, h_s_wallace_rca24_fa124_y2, h_s_wallace_rca24_fa124_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_6_y0(a_5, b_6, h_s_wallace_rca24_and_5_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_7_y0(a_4, b_7, h_s_wallace_rca24_and_4_7_y0);
  fa fa_h_s_wallace_rca24_fa125_y2(h_s_wallace_rca24_fa124_y4, h_s_wallace_rca24_and_5_6_y0, h_s_wallace_rca24_and_4_7_y0, h_s_wallace_rca24_fa125_y2, h_s_wallace_rca24_fa125_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_6_y0(a_6, b_6, h_s_wallace_rca24_and_6_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_7_y0(a_5, b_7, h_s_wallace_rca24_and_5_7_y0);
  fa fa_h_s_wallace_rca24_fa126_y2(h_s_wallace_rca24_fa125_y4, h_s_wallace_rca24_and_6_6_y0, h_s_wallace_rca24_and_5_7_y0, h_s_wallace_rca24_fa126_y2, h_s_wallace_rca24_fa126_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_6_y0(a_7, b_6, h_s_wallace_rca24_and_7_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_7_y0(a_6, b_7, h_s_wallace_rca24_and_6_7_y0);
  fa fa_h_s_wallace_rca24_fa127_y2(h_s_wallace_rca24_fa126_y4, h_s_wallace_rca24_and_7_6_y0, h_s_wallace_rca24_and_6_7_y0, h_s_wallace_rca24_fa127_y2, h_s_wallace_rca24_fa127_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_6_y0(a_8, b_6, h_s_wallace_rca24_and_8_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_7_y0(a_7, b_7, h_s_wallace_rca24_and_7_7_y0);
  fa fa_h_s_wallace_rca24_fa128_y2(h_s_wallace_rca24_fa127_y4, h_s_wallace_rca24_and_8_6_y0, h_s_wallace_rca24_and_7_7_y0, h_s_wallace_rca24_fa128_y2, h_s_wallace_rca24_fa128_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_6_y0(a_9, b_6, h_s_wallace_rca24_and_9_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_7_y0(a_8, b_7, h_s_wallace_rca24_and_8_7_y0);
  fa fa_h_s_wallace_rca24_fa129_y2(h_s_wallace_rca24_fa128_y4, h_s_wallace_rca24_and_9_6_y0, h_s_wallace_rca24_and_8_7_y0, h_s_wallace_rca24_fa129_y2, h_s_wallace_rca24_fa129_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_6_y0(a_10, b_6, h_s_wallace_rca24_and_10_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_7_y0(a_9, b_7, h_s_wallace_rca24_and_9_7_y0);
  fa fa_h_s_wallace_rca24_fa130_y2(h_s_wallace_rca24_fa129_y4, h_s_wallace_rca24_and_10_6_y0, h_s_wallace_rca24_and_9_7_y0, h_s_wallace_rca24_fa130_y2, h_s_wallace_rca24_fa130_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_6_y0(a_11, b_6, h_s_wallace_rca24_and_11_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_7_y0(a_10, b_7, h_s_wallace_rca24_and_10_7_y0);
  fa fa_h_s_wallace_rca24_fa131_y2(h_s_wallace_rca24_fa130_y4, h_s_wallace_rca24_and_11_6_y0, h_s_wallace_rca24_and_10_7_y0, h_s_wallace_rca24_fa131_y2, h_s_wallace_rca24_fa131_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_6_y0(a_12, b_6, h_s_wallace_rca24_and_12_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_7_y0(a_11, b_7, h_s_wallace_rca24_and_11_7_y0);
  fa fa_h_s_wallace_rca24_fa132_y2(h_s_wallace_rca24_fa131_y4, h_s_wallace_rca24_and_12_6_y0, h_s_wallace_rca24_and_11_7_y0, h_s_wallace_rca24_fa132_y2, h_s_wallace_rca24_fa132_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_6_y0(a_13, b_6, h_s_wallace_rca24_and_13_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_7_y0(a_12, b_7, h_s_wallace_rca24_and_12_7_y0);
  fa fa_h_s_wallace_rca24_fa133_y2(h_s_wallace_rca24_fa132_y4, h_s_wallace_rca24_and_13_6_y0, h_s_wallace_rca24_and_12_7_y0, h_s_wallace_rca24_fa133_y2, h_s_wallace_rca24_fa133_y4);
  and_gate and_gate_h_s_wallace_rca24_and_14_6_y0(a_14, b_6, h_s_wallace_rca24_and_14_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_13_7_y0(a_13, b_7, h_s_wallace_rca24_and_13_7_y0);
  fa fa_h_s_wallace_rca24_fa134_y2(h_s_wallace_rca24_fa133_y4, h_s_wallace_rca24_and_14_6_y0, h_s_wallace_rca24_and_13_7_y0, h_s_wallace_rca24_fa134_y2, h_s_wallace_rca24_fa134_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_6_y0(a_15, b_6, h_s_wallace_rca24_and_15_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_7_y0(a_14, b_7, h_s_wallace_rca24_and_14_7_y0);
  fa fa_h_s_wallace_rca24_fa135_y2(h_s_wallace_rca24_fa134_y4, h_s_wallace_rca24_and_15_6_y0, h_s_wallace_rca24_and_14_7_y0, h_s_wallace_rca24_fa135_y2, h_s_wallace_rca24_fa135_y4);
  and_gate and_gate_h_s_wallace_rca24_and_16_6_y0(a_16, b_6, h_s_wallace_rca24_and_16_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_15_7_y0(a_15, b_7, h_s_wallace_rca24_and_15_7_y0);
  fa fa_h_s_wallace_rca24_fa136_y2(h_s_wallace_rca24_fa135_y4, h_s_wallace_rca24_and_16_6_y0, h_s_wallace_rca24_and_15_7_y0, h_s_wallace_rca24_fa136_y2, h_s_wallace_rca24_fa136_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_6_y0(a_17, b_6, h_s_wallace_rca24_and_17_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_7_y0(a_16, b_7, h_s_wallace_rca24_and_16_7_y0);
  fa fa_h_s_wallace_rca24_fa137_y2(h_s_wallace_rca24_fa136_y4, h_s_wallace_rca24_and_17_6_y0, h_s_wallace_rca24_and_16_7_y0, h_s_wallace_rca24_fa137_y2, h_s_wallace_rca24_fa137_y4);
  and_gate and_gate_h_s_wallace_rca24_and_18_6_y0(a_18, b_6, h_s_wallace_rca24_and_18_6_y0);
  and_gate and_gate_h_s_wallace_rca24_and_17_7_y0(a_17, b_7, h_s_wallace_rca24_and_17_7_y0);
  fa fa_h_s_wallace_rca24_fa138_y2(h_s_wallace_rca24_fa137_y4, h_s_wallace_rca24_and_18_6_y0, h_s_wallace_rca24_and_17_7_y0, h_s_wallace_rca24_fa138_y2, h_s_wallace_rca24_fa138_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_8_y0(a_17, b_8, h_s_wallace_rca24_and_17_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_9_y0(a_16, b_9, h_s_wallace_rca24_and_16_9_y0);
  fa fa_h_s_wallace_rca24_fa139_y2(h_s_wallace_rca24_fa138_y4, h_s_wallace_rca24_and_17_8_y0, h_s_wallace_rca24_and_16_9_y0, h_s_wallace_rca24_fa139_y2, h_s_wallace_rca24_fa139_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_9_y0(a_17, b_9, h_s_wallace_rca24_and_17_9_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_10_y0(a_16, b_10, h_s_wallace_rca24_and_16_10_y0);
  fa fa_h_s_wallace_rca24_fa140_y2(h_s_wallace_rca24_fa139_y4, h_s_wallace_rca24_and_17_9_y0, h_s_wallace_rca24_and_16_10_y0, h_s_wallace_rca24_fa140_y2, h_s_wallace_rca24_fa140_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_10_y0(a_17, b_10, h_s_wallace_rca24_and_17_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_11_y0(a_16, b_11, h_s_wallace_rca24_and_16_11_y0);
  fa fa_h_s_wallace_rca24_fa141_y2(h_s_wallace_rca24_fa140_y4, h_s_wallace_rca24_and_17_10_y0, h_s_wallace_rca24_and_16_11_y0, h_s_wallace_rca24_fa141_y2, h_s_wallace_rca24_fa141_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_11_y0(a_17, b_11, h_s_wallace_rca24_and_17_11_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_12_y0(a_16, b_12, h_s_wallace_rca24_and_16_12_y0);
  fa fa_h_s_wallace_rca24_fa142_y2(h_s_wallace_rca24_fa141_y4, h_s_wallace_rca24_and_17_11_y0, h_s_wallace_rca24_and_16_12_y0, h_s_wallace_rca24_fa142_y2, h_s_wallace_rca24_fa142_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_12_y0(a_17, b_12, h_s_wallace_rca24_and_17_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_13_y0(a_16, b_13, h_s_wallace_rca24_and_16_13_y0);
  fa fa_h_s_wallace_rca24_fa143_y2(h_s_wallace_rca24_fa142_y4, h_s_wallace_rca24_and_17_12_y0, h_s_wallace_rca24_and_16_13_y0, h_s_wallace_rca24_fa143_y2, h_s_wallace_rca24_fa143_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_13_y0(a_17, b_13, h_s_wallace_rca24_and_17_13_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_14_y0(a_16, b_14, h_s_wallace_rca24_and_16_14_y0);
  fa fa_h_s_wallace_rca24_fa144_y2(h_s_wallace_rca24_fa143_y4, h_s_wallace_rca24_and_17_13_y0, h_s_wallace_rca24_and_16_14_y0, h_s_wallace_rca24_fa144_y2, h_s_wallace_rca24_fa144_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_14_y0(a_17, b_14, h_s_wallace_rca24_and_17_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_15_y0(a_16, b_15, h_s_wallace_rca24_and_16_15_y0);
  fa fa_h_s_wallace_rca24_fa145_y2(h_s_wallace_rca24_fa144_y4, h_s_wallace_rca24_and_17_14_y0, h_s_wallace_rca24_and_16_15_y0, h_s_wallace_rca24_fa145_y2, h_s_wallace_rca24_fa145_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_15_y0(a_17, b_15, h_s_wallace_rca24_and_17_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_16_y0(a_16, b_16, h_s_wallace_rca24_and_16_16_y0);
  fa fa_h_s_wallace_rca24_fa146_y2(h_s_wallace_rca24_fa145_y4, h_s_wallace_rca24_and_17_15_y0, h_s_wallace_rca24_and_16_16_y0, h_s_wallace_rca24_fa146_y2, h_s_wallace_rca24_fa146_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_16_y0(a_17, b_16, h_s_wallace_rca24_and_17_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_17_y0(a_16, b_17, h_s_wallace_rca24_and_16_17_y0);
  fa fa_h_s_wallace_rca24_fa147_y2(h_s_wallace_rca24_fa146_y4, h_s_wallace_rca24_and_17_16_y0, h_s_wallace_rca24_and_16_17_y0, h_s_wallace_rca24_fa147_y2, h_s_wallace_rca24_fa147_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_17_y0(a_17, b_17, h_s_wallace_rca24_and_17_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_18_y0(a_16, b_18, h_s_wallace_rca24_and_16_18_y0);
  fa fa_h_s_wallace_rca24_fa148_y2(h_s_wallace_rca24_fa147_y4, h_s_wallace_rca24_and_17_17_y0, h_s_wallace_rca24_and_16_18_y0, h_s_wallace_rca24_fa148_y2, h_s_wallace_rca24_fa148_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_18_y0(a_17, b_18, h_s_wallace_rca24_and_17_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_19_y0(a_16, b_19, h_s_wallace_rca24_and_16_19_y0);
  fa fa_h_s_wallace_rca24_fa149_y2(h_s_wallace_rca24_fa148_y4, h_s_wallace_rca24_and_17_18_y0, h_s_wallace_rca24_and_16_19_y0, h_s_wallace_rca24_fa149_y2, h_s_wallace_rca24_fa149_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_19_y0(a_17, b_19, h_s_wallace_rca24_and_17_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_20_y0(a_16, b_20, h_s_wallace_rca24_and_16_20_y0);
  fa fa_h_s_wallace_rca24_fa150_y2(h_s_wallace_rca24_fa149_y4, h_s_wallace_rca24_and_17_19_y0, h_s_wallace_rca24_and_16_20_y0, h_s_wallace_rca24_fa150_y2, h_s_wallace_rca24_fa150_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_20_y0(a_17, b_20, h_s_wallace_rca24_and_17_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_21_y0(a_16, b_21, h_s_wallace_rca24_and_16_21_y0);
  fa fa_h_s_wallace_rca24_fa151_y2(h_s_wallace_rca24_fa150_y4, h_s_wallace_rca24_and_17_20_y0, h_s_wallace_rca24_and_16_21_y0, h_s_wallace_rca24_fa151_y2, h_s_wallace_rca24_fa151_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_21_y0(a_17, b_21, h_s_wallace_rca24_and_17_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_16_22_y0(a_16, b_22, h_s_wallace_rca24_and_16_22_y0);
  fa fa_h_s_wallace_rca24_fa152_y2(h_s_wallace_rca24_fa151_y4, h_s_wallace_rca24_and_17_21_y0, h_s_wallace_rca24_and_16_22_y0, h_s_wallace_rca24_fa152_y2, h_s_wallace_rca24_fa152_y4);
  and_gate and_gate_h_s_wallace_rca24_and_17_22_y0(a_17, b_22, h_s_wallace_rca24_and_17_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_16_23_y0(a_16, b_23, h_s_wallace_rca24_nand_16_23_y0);
  fa fa_h_s_wallace_rca24_fa153_y2(h_s_wallace_rca24_fa152_y4, h_s_wallace_rca24_and_17_22_y0, h_s_wallace_rca24_nand_16_23_y0, h_s_wallace_rca24_fa153_y2, h_s_wallace_rca24_fa153_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_17_23_y0(a_17, b_23, h_s_wallace_rca24_nand_17_23_y0);
  fa fa_h_s_wallace_rca24_fa154_y2(h_s_wallace_rca24_fa153_y4, h_s_wallace_rca24_nand_17_23_y0, h_s_wallace_rca24_fa37_y2, h_s_wallace_rca24_fa154_y2, h_s_wallace_rca24_fa154_y4);
  fa fa_h_s_wallace_rca24_fa155_y2(h_s_wallace_rca24_fa154_y4, h_s_wallace_rca24_fa38_y2, h_s_wallace_rca24_fa79_y2, h_s_wallace_rca24_fa155_y2, h_s_wallace_rca24_fa155_y4);
  ha ha_h_s_wallace_rca24_ha4_y0(h_s_wallace_rca24_fa44_y2, h_s_wallace_rca24_fa83_y2, h_s_wallace_rca24_ha4_y0, h_s_wallace_rca24_ha4_y1);
  fa fa_h_s_wallace_rca24_fa156_y2(h_s_wallace_rca24_ha4_y1, h_s_wallace_rca24_fa4_y2, h_s_wallace_rca24_fa45_y2, h_s_wallace_rca24_fa156_y2, h_s_wallace_rca24_fa156_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_8_y0(a_0, b_8, h_s_wallace_rca24_and_0_8_y0);
  fa fa_h_s_wallace_rca24_fa157_y2(h_s_wallace_rca24_fa156_y4, h_s_wallace_rca24_and_0_8_y0, h_s_wallace_rca24_fa5_y2, h_s_wallace_rca24_fa157_y2, h_s_wallace_rca24_fa157_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_8_y0(a_1, b_8, h_s_wallace_rca24_and_1_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_9_y0(a_0, b_9, h_s_wallace_rca24_and_0_9_y0);
  fa fa_h_s_wallace_rca24_fa158_y2(h_s_wallace_rca24_fa157_y4, h_s_wallace_rca24_and_1_8_y0, h_s_wallace_rca24_and_0_9_y0, h_s_wallace_rca24_fa158_y2, h_s_wallace_rca24_fa158_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_8_y0(a_2, b_8, h_s_wallace_rca24_and_2_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_9_y0(a_1, b_9, h_s_wallace_rca24_and_1_9_y0);
  fa fa_h_s_wallace_rca24_fa159_y2(h_s_wallace_rca24_fa158_y4, h_s_wallace_rca24_and_2_8_y0, h_s_wallace_rca24_and_1_9_y0, h_s_wallace_rca24_fa159_y2, h_s_wallace_rca24_fa159_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_8_y0(a_3, b_8, h_s_wallace_rca24_and_3_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_9_y0(a_2, b_9, h_s_wallace_rca24_and_2_9_y0);
  fa fa_h_s_wallace_rca24_fa160_y2(h_s_wallace_rca24_fa159_y4, h_s_wallace_rca24_and_3_8_y0, h_s_wallace_rca24_and_2_9_y0, h_s_wallace_rca24_fa160_y2, h_s_wallace_rca24_fa160_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_8_y0(a_4, b_8, h_s_wallace_rca24_and_4_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_9_y0(a_3, b_9, h_s_wallace_rca24_and_3_9_y0);
  fa fa_h_s_wallace_rca24_fa161_y2(h_s_wallace_rca24_fa160_y4, h_s_wallace_rca24_and_4_8_y0, h_s_wallace_rca24_and_3_9_y0, h_s_wallace_rca24_fa161_y2, h_s_wallace_rca24_fa161_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_8_y0(a_5, b_8, h_s_wallace_rca24_and_5_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_9_y0(a_4, b_9, h_s_wallace_rca24_and_4_9_y0);
  fa fa_h_s_wallace_rca24_fa162_y2(h_s_wallace_rca24_fa161_y4, h_s_wallace_rca24_and_5_8_y0, h_s_wallace_rca24_and_4_9_y0, h_s_wallace_rca24_fa162_y2, h_s_wallace_rca24_fa162_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_8_y0(a_6, b_8, h_s_wallace_rca24_and_6_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_9_y0(a_5, b_9, h_s_wallace_rca24_and_5_9_y0);
  fa fa_h_s_wallace_rca24_fa163_y2(h_s_wallace_rca24_fa162_y4, h_s_wallace_rca24_and_6_8_y0, h_s_wallace_rca24_and_5_9_y0, h_s_wallace_rca24_fa163_y2, h_s_wallace_rca24_fa163_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_8_y0(a_7, b_8, h_s_wallace_rca24_and_7_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_9_y0(a_6, b_9, h_s_wallace_rca24_and_6_9_y0);
  fa fa_h_s_wallace_rca24_fa164_y2(h_s_wallace_rca24_fa163_y4, h_s_wallace_rca24_and_7_8_y0, h_s_wallace_rca24_and_6_9_y0, h_s_wallace_rca24_fa164_y2, h_s_wallace_rca24_fa164_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_8_y0(a_8, b_8, h_s_wallace_rca24_and_8_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_9_y0(a_7, b_9, h_s_wallace_rca24_and_7_9_y0);
  fa fa_h_s_wallace_rca24_fa165_y2(h_s_wallace_rca24_fa164_y4, h_s_wallace_rca24_and_8_8_y0, h_s_wallace_rca24_and_7_9_y0, h_s_wallace_rca24_fa165_y2, h_s_wallace_rca24_fa165_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_8_y0(a_9, b_8, h_s_wallace_rca24_and_9_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_9_y0(a_8, b_9, h_s_wallace_rca24_and_8_9_y0);
  fa fa_h_s_wallace_rca24_fa166_y2(h_s_wallace_rca24_fa165_y4, h_s_wallace_rca24_and_9_8_y0, h_s_wallace_rca24_and_8_9_y0, h_s_wallace_rca24_fa166_y2, h_s_wallace_rca24_fa166_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_8_y0(a_10, b_8, h_s_wallace_rca24_and_10_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_9_y0(a_9, b_9, h_s_wallace_rca24_and_9_9_y0);
  fa fa_h_s_wallace_rca24_fa167_y2(h_s_wallace_rca24_fa166_y4, h_s_wallace_rca24_and_10_8_y0, h_s_wallace_rca24_and_9_9_y0, h_s_wallace_rca24_fa167_y2, h_s_wallace_rca24_fa167_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_8_y0(a_11, b_8, h_s_wallace_rca24_and_11_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_9_y0(a_10, b_9, h_s_wallace_rca24_and_10_9_y0);
  fa fa_h_s_wallace_rca24_fa168_y2(h_s_wallace_rca24_fa167_y4, h_s_wallace_rca24_and_11_8_y0, h_s_wallace_rca24_and_10_9_y0, h_s_wallace_rca24_fa168_y2, h_s_wallace_rca24_fa168_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_8_y0(a_12, b_8, h_s_wallace_rca24_and_12_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_9_y0(a_11, b_9, h_s_wallace_rca24_and_11_9_y0);
  fa fa_h_s_wallace_rca24_fa169_y2(h_s_wallace_rca24_fa168_y4, h_s_wallace_rca24_and_12_8_y0, h_s_wallace_rca24_and_11_9_y0, h_s_wallace_rca24_fa169_y2, h_s_wallace_rca24_fa169_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_8_y0(a_13, b_8, h_s_wallace_rca24_and_13_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_9_y0(a_12, b_9, h_s_wallace_rca24_and_12_9_y0);
  fa fa_h_s_wallace_rca24_fa170_y2(h_s_wallace_rca24_fa169_y4, h_s_wallace_rca24_and_13_8_y0, h_s_wallace_rca24_and_12_9_y0, h_s_wallace_rca24_fa170_y2, h_s_wallace_rca24_fa170_y4);
  and_gate and_gate_h_s_wallace_rca24_and_14_8_y0(a_14, b_8, h_s_wallace_rca24_and_14_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_13_9_y0(a_13, b_9, h_s_wallace_rca24_and_13_9_y0);
  fa fa_h_s_wallace_rca24_fa171_y2(h_s_wallace_rca24_fa170_y4, h_s_wallace_rca24_and_14_8_y0, h_s_wallace_rca24_and_13_9_y0, h_s_wallace_rca24_fa171_y2, h_s_wallace_rca24_fa171_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_8_y0(a_15, b_8, h_s_wallace_rca24_and_15_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_9_y0(a_14, b_9, h_s_wallace_rca24_and_14_9_y0);
  fa fa_h_s_wallace_rca24_fa172_y2(h_s_wallace_rca24_fa171_y4, h_s_wallace_rca24_and_15_8_y0, h_s_wallace_rca24_and_14_9_y0, h_s_wallace_rca24_fa172_y2, h_s_wallace_rca24_fa172_y4);
  and_gate and_gate_h_s_wallace_rca24_and_16_8_y0(a_16, b_8, h_s_wallace_rca24_and_16_8_y0);
  and_gate and_gate_h_s_wallace_rca24_and_15_9_y0(a_15, b_9, h_s_wallace_rca24_and_15_9_y0);
  fa fa_h_s_wallace_rca24_fa173_y2(h_s_wallace_rca24_fa172_y4, h_s_wallace_rca24_and_16_8_y0, h_s_wallace_rca24_and_15_9_y0, h_s_wallace_rca24_fa173_y2, h_s_wallace_rca24_fa173_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_10_y0(a_15, b_10, h_s_wallace_rca24_and_15_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_11_y0(a_14, b_11, h_s_wallace_rca24_and_14_11_y0);
  fa fa_h_s_wallace_rca24_fa174_y2(h_s_wallace_rca24_fa173_y4, h_s_wallace_rca24_and_15_10_y0, h_s_wallace_rca24_and_14_11_y0, h_s_wallace_rca24_fa174_y2, h_s_wallace_rca24_fa174_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_11_y0(a_15, b_11, h_s_wallace_rca24_and_15_11_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_12_y0(a_14, b_12, h_s_wallace_rca24_and_14_12_y0);
  fa fa_h_s_wallace_rca24_fa175_y2(h_s_wallace_rca24_fa174_y4, h_s_wallace_rca24_and_15_11_y0, h_s_wallace_rca24_and_14_12_y0, h_s_wallace_rca24_fa175_y2, h_s_wallace_rca24_fa175_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_12_y0(a_15, b_12, h_s_wallace_rca24_and_15_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_13_y0(a_14, b_13, h_s_wallace_rca24_and_14_13_y0);
  fa fa_h_s_wallace_rca24_fa176_y2(h_s_wallace_rca24_fa175_y4, h_s_wallace_rca24_and_15_12_y0, h_s_wallace_rca24_and_14_13_y0, h_s_wallace_rca24_fa176_y2, h_s_wallace_rca24_fa176_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_13_y0(a_15, b_13, h_s_wallace_rca24_and_15_13_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_14_y0(a_14, b_14, h_s_wallace_rca24_and_14_14_y0);
  fa fa_h_s_wallace_rca24_fa177_y2(h_s_wallace_rca24_fa176_y4, h_s_wallace_rca24_and_15_13_y0, h_s_wallace_rca24_and_14_14_y0, h_s_wallace_rca24_fa177_y2, h_s_wallace_rca24_fa177_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_14_y0(a_15, b_14, h_s_wallace_rca24_and_15_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_15_y0(a_14, b_15, h_s_wallace_rca24_and_14_15_y0);
  fa fa_h_s_wallace_rca24_fa178_y2(h_s_wallace_rca24_fa177_y4, h_s_wallace_rca24_and_15_14_y0, h_s_wallace_rca24_and_14_15_y0, h_s_wallace_rca24_fa178_y2, h_s_wallace_rca24_fa178_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_15_y0(a_15, b_15, h_s_wallace_rca24_and_15_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_16_y0(a_14, b_16, h_s_wallace_rca24_and_14_16_y0);
  fa fa_h_s_wallace_rca24_fa179_y2(h_s_wallace_rca24_fa178_y4, h_s_wallace_rca24_and_15_15_y0, h_s_wallace_rca24_and_14_16_y0, h_s_wallace_rca24_fa179_y2, h_s_wallace_rca24_fa179_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_16_y0(a_15, b_16, h_s_wallace_rca24_and_15_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_17_y0(a_14, b_17, h_s_wallace_rca24_and_14_17_y0);
  fa fa_h_s_wallace_rca24_fa180_y2(h_s_wallace_rca24_fa179_y4, h_s_wallace_rca24_and_15_16_y0, h_s_wallace_rca24_and_14_17_y0, h_s_wallace_rca24_fa180_y2, h_s_wallace_rca24_fa180_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_17_y0(a_15, b_17, h_s_wallace_rca24_and_15_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_18_y0(a_14, b_18, h_s_wallace_rca24_and_14_18_y0);
  fa fa_h_s_wallace_rca24_fa181_y2(h_s_wallace_rca24_fa180_y4, h_s_wallace_rca24_and_15_17_y0, h_s_wallace_rca24_and_14_18_y0, h_s_wallace_rca24_fa181_y2, h_s_wallace_rca24_fa181_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_18_y0(a_15, b_18, h_s_wallace_rca24_and_15_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_19_y0(a_14, b_19, h_s_wallace_rca24_and_14_19_y0);
  fa fa_h_s_wallace_rca24_fa182_y2(h_s_wallace_rca24_fa181_y4, h_s_wallace_rca24_and_15_18_y0, h_s_wallace_rca24_and_14_19_y0, h_s_wallace_rca24_fa182_y2, h_s_wallace_rca24_fa182_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_19_y0(a_15, b_19, h_s_wallace_rca24_and_15_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_20_y0(a_14, b_20, h_s_wallace_rca24_and_14_20_y0);
  fa fa_h_s_wallace_rca24_fa183_y2(h_s_wallace_rca24_fa182_y4, h_s_wallace_rca24_and_15_19_y0, h_s_wallace_rca24_and_14_20_y0, h_s_wallace_rca24_fa183_y2, h_s_wallace_rca24_fa183_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_20_y0(a_15, b_20, h_s_wallace_rca24_and_15_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_21_y0(a_14, b_21, h_s_wallace_rca24_and_14_21_y0);
  fa fa_h_s_wallace_rca24_fa184_y2(h_s_wallace_rca24_fa183_y4, h_s_wallace_rca24_and_15_20_y0, h_s_wallace_rca24_and_14_21_y0, h_s_wallace_rca24_fa184_y2, h_s_wallace_rca24_fa184_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_21_y0(a_15, b_21, h_s_wallace_rca24_and_15_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_14_22_y0(a_14, b_22, h_s_wallace_rca24_and_14_22_y0);
  fa fa_h_s_wallace_rca24_fa185_y2(h_s_wallace_rca24_fa184_y4, h_s_wallace_rca24_and_15_21_y0, h_s_wallace_rca24_and_14_22_y0, h_s_wallace_rca24_fa185_y2, h_s_wallace_rca24_fa185_y4);
  and_gate and_gate_h_s_wallace_rca24_and_15_22_y0(a_15, b_22, h_s_wallace_rca24_and_15_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_14_23_y0(a_14, b_23, h_s_wallace_rca24_nand_14_23_y0);
  fa fa_h_s_wallace_rca24_fa186_y2(h_s_wallace_rca24_fa185_y4, h_s_wallace_rca24_and_15_22_y0, h_s_wallace_rca24_nand_14_23_y0, h_s_wallace_rca24_fa186_y2, h_s_wallace_rca24_fa186_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_15_23_y0(a_15, b_23, h_s_wallace_rca24_nand_15_23_y0);
  fa fa_h_s_wallace_rca24_fa187_y2(h_s_wallace_rca24_fa186_y4, h_s_wallace_rca24_nand_15_23_y0, h_s_wallace_rca24_fa35_y2, h_s_wallace_rca24_fa187_y2, h_s_wallace_rca24_fa187_y4);
  fa fa_h_s_wallace_rca24_fa188_y2(h_s_wallace_rca24_fa187_y4, h_s_wallace_rca24_fa36_y2, h_s_wallace_rca24_fa77_y2, h_s_wallace_rca24_fa188_y2, h_s_wallace_rca24_fa188_y4);
  fa fa_h_s_wallace_rca24_fa189_y2(h_s_wallace_rca24_fa188_y4, h_s_wallace_rca24_fa78_y2, h_s_wallace_rca24_fa117_y2, h_s_wallace_rca24_fa189_y2, h_s_wallace_rca24_fa189_y4);
  ha ha_h_s_wallace_rca24_ha5_y0(h_s_wallace_rca24_fa84_y2, h_s_wallace_rca24_fa121_y2, h_s_wallace_rca24_ha5_y0, h_s_wallace_rca24_ha5_y1);
  fa fa_h_s_wallace_rca24_fa190_y2(h_s_wallace_rca24_ha5_y1, h_s_wallace_rca24_fa46_y2, h_s_wallace_rca24_fa85_y2, h_s_wallace_rca24_fa190_y2, h_s_wallace_rca24_fa190_y4);
  fa fa_h_s_wallace_rca24_fa191_y2(h_s_wallace_rca24_fa190_y4, h_s_wallace_rca24_fa6_y2, h_s_wallace_rca24_fa47_y2, h_s_wallace_rca24_fa191_y2, h_s_wallace_rca24_fa191_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_10_y0(a_0, b_10, h_s_wallace_rca24_and_0_10_y0);
  fa fa_h_s_wallace_rca24_fa192_y2(h_s_wallace_rca24_fa191_y4, h_s_wallace_rca24_and_0_10_y0, h_s_wallace_rca24_fa7_y2, h_s_wallace_rca24_fa192_y2, h_s_wallace_rca24_fa192_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_10_y0(a_1, b_10, h_s_wallace_rca24_and_1_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_11_y0(a_0, b_11, h_s_wallace_rca24_and_0_11_y0);
  fa fa_h_s_wallace_rca24_fa193_y2(h_s_wallace_rca24_fa192_y4, h_s_wallace_rca24_and_1_10_y0, h_s_wallace_rca24_and_0_11_y0, h_s_wallace_rca24_fa193_y2, h_s_wallace_rca24_fa193_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_10_y0(a_2, b_10, h_s_wallace_rca24_and_2_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_11_y0(a_1, b_11, h_s_wallace_rca24_and_1_11_y0);
  fa fa_h_s_wallace_rca24_fa194_y2(h_s_wallace_rca24_fa193_y4, h_s_wallace_rca24_and_2_10_y0, h_s_wallace_rca24_and_1_11_y0, h_s_wallace_rca24_fa194_y2, h_s_wallace_rca24_fa194_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_10_y0(a_3, b_10, h_s_wallace_rca24_and_3_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_11_y0(a_2, b_11, h_s_wallace_rca24_and_2_11_y0);
  fa fa_h_s_wallace_rca24_fa195_y2(h_s_wallace_rca24_fa194_y4, h_s_wallace_rca24_and_3_10_y0, h_s_wallace_rca24_and_2_11_y0, h_s_wallace_rca24_fa195_y2, h_s_wallace_rca24_fa195_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_10_y0(a_4, b_10, h_s_wallace_rca24_and_4_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_11_y0(a_3, b_11, h_s_wallace_rca24_and_3_11_y0);
  fa fa_h_s_wallace_rca24_fa196_y2(h_s_wallace_rca24_fa195_y4, h_s_wallace_rca24_and_4_10_y0, h_s_wallace_rca24_and_3_11_y0, h_s_wallace_rca24_fa196_y2, h_s_wallace_rca24_fa196_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_10_y0(a_5, b_10, h_s_wallace_rca24_and_5_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_11_y0(a_4, b_11, h_s_wallace_rca24_and_4_11_y0);
  fa fa_h_s_wallace_rca24_fa197_y2(h_s_wallace_rca24_fa196_y4, h_s_wallace_rca24_and_5_10_y0, h_s_wallace_rca24_and_4_11_y0, h_s_wallace_rca24_fa197_y2, h_s_wallace_rca24_fa197_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_10_y0(a_6, b_10, h_s_wallace_rca24_and_6_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_11_y0(a_5, b_11, h_s_wallace_rca24_and_5_11_y0);
  fa fa_h_s_wallace_rca24_fa198_y2(h_s_wallace_rca24_fa197_y4, h_s_wallace_rca24_and_6_10_y0, h_s_wallace_rca24_and_5_11_y0, h_s_wallace_rca24_fa198_y2, h_s_wallace_rca24_fa198_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_10_y0(a_7, b_10, h_s_wallace_rca24_and_7_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_11_y0(a_6, b_11, h_s_wallace_rca24_and_6_11_y0);
  fa fa_h_s_wallace_rca24_fa199_y2(h_s_wallace_rca24_fa198_y4, h_s_wallace_rca24_and_7_10_y0, h_s_wallace_rca24_and_6_11_y0, h_s_wallace_rca24_fa199_y2, h_s_wallace_rca24_fa199_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_10_y0(a_8, b_10, h_s_wallace_rca24_and_8_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_11_y0(a_7, b_11, h_s_wallace_rca24_and_7_11_y0);
  fa fa_h_s_wallace_rca24_fa200_y2(h_s_wallace_rca24_fa199_y4, h_s_wallace_rca24_and_8_10_y0, h_s_wallace_rca24_and_7_11_y0, h_s_wallace_rca24_fa200_y2, h_s_wallace_rca24_fa200_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_10_y0(a_9, b_10, h_s_wallace_rca24_and_9_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_11_y0(a_8, b_11, h_s_wallace_rca24_and_8_11_y0);
  fa fa_h_s_wallace_rca24_fa201_y2(h_s_wallace_rca24_fa200_y4, h_s_wallace_rca24_and_9_10_y0, h_s_wallace_rca24_and_8_11_y0, h_s_wallace_rca24_fa201_y2, h_s_wallace_rca24_fa201_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_10_y0(a_10, b_10, h_s_wallace_rca24_and_10_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_11_y0(a_9, b_11, h_s_wallace_rca24_and_9_11_y0);
  fa fa_h_s_wallace_rca24_fa202_y2(h_s_wallace_rca24_fa201_y4, h_s_wallace_rca24_and_10_10_y0, h_s_wallace_rca24_and_9_11_y0, h_s_wallace_rca24_fa202_y2, h_s_wallace_rca24_fa202_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_10_y0(a_11, b_10, h_s_wallace_rca24_and_11_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_11_y0(a_10, b_11, h_s_wallace_rca24_and_10_11_y0);
  fa fa_h_s_wallace_rca24_fa203_y2(h_s_wallace_rca24_fa202_y4, h_s_wallace_rca24_and_11_10_y0, h_s_wallace_rca24_and_10_11_y0, h_s_wallace_rca24_fa203_y2, h_s_wallace_rca24_fa203_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_10_y0(a_12, b_10, h_s_wallace_rca24_and_12_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_11_y0(a_11, b_11, h_s_wallace_rca24_and_11_11_y0);
  fa fa_h_s_wallace_rca24_fa204_y2(h_s_wallace_rca24_fa203_y4, h_s_wallace_rca24_and_12_10_y0, h_s_wallace_rca24_and_11_11_y0, h_s_wallace_rca24_fa204_y2, h_s_wallace_rca24_fa204_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_10_y0(a_13, b_10, h_s_wallace_rca24_and_13_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_11_y0(a_12, b_11, h_s_wallace_rca24_and_12_11_y0);
  fa fa_h_s_wallace_rca24_fa205_y2(h_s_wallace_rca24_fa204_y4, h_s_wallace_rca24_and_13_10_y0, h_s_wallace_rca24_and_12_11_y0, h_s_wallace_rca24_fa205_y2, h_s_wallace_rca24_fa205_y4);
  and_gate and_gate_h_s_wallace_rca24_and_14_10_y0(a_14, b_10, h_s_wallace_rca24_and_14_10_y0);
  and_gate and_gate_h_s_wallace_rca24_and_13_11_y0(a_13, b_11, h_s_wallace_rca24_and_13_11_y0);
  fa fa_h_s_wallace_rca24_fa206_y2(h_s_wallace_rca24_fa205_y4, h_s_wallace_rca24_and_14_10_y0, h_s_wallace_rca24_and_13_11_y0, h_s_wallace_rca24_fa206_y2, h_s_wallace_rca24_fa206_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_12_y0(a_13, b_12, h_s_wallace_rca24_and_13_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_13_y0(a_12, b_13, h_s_wallace_rca24_and_12_13_y0);
  fa fa_h_s_wallace_rca24_fa207_y2(h_s_wallace_rca24_fa206_y4, h_s_wallace_rca24_and_13_12_y0, h_s_wallace_rca24_and_12_13_y0, h_s_wallace_rca24_fa207_y2, h_s_wallace_rca24_fa207_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_13_y0(a_13, b_13, h_s_wallace_rca24_and_13_13_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_14_y0(a_12, b_14, h_s_wallace_rca24_and_12_14_y0);
  fa fa_h_s_wallace_rca24_fa208_y2(h_s_wallace_rca24_fa207_y4, h_s_wallace_rca24_and_13_13_y0, h_s_wallace_rca24_and_12_14_y0, h_s_wallace_rca24_fa208_y2, h_s_wallace_rca24_fa208_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_14_y0(a_13, b_14, h_s_wallace_rca24_and_13_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_15_y0(a_12, b_15, h_s_wallace_rca24_and_12_15_y0);
  fa fa_h_s_wallace_rca24_fa209_y2(h_s_wallace_rca24_fa208_y4, h_s_wallace_rca24_and_13_14_y0, h_s_wallace_rca24_and_12_15_y0, h_s_wallace_rca24_fa209_y2, h_s_wallace_rca24_fa209_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_15_y0(a_13, b_15, h_s_wallace_rca24_and_13_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_16_y0(a_12, b_16, h_s_wallace_rca24_and_12_16_y0);
  fa fa_h_s_wallace_rca24_fa210_y2(h_s_wallace_rca24_fa209_y4, h_s_wallace_rca24_and_13_15_y0, h_s_wallace_rca24_and_12_16_y0, h_s_wallace_rca24_fa210_y2, h_s_wallace_rca24_fa210_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_16_y0(a_13, b_16, h_s_wallace_rca24_and_13_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_17_y0(a_12, b_17, h_s_wallace_rca24_and_12_17_y0);
  fa fa_h_s_wallace_rca24_fa211_y2(h_s_wallace_rca24_fa210_y4, h_s_wallace_rca24_and_13_16_y0, h_s_wallace_rca24_and_12_17_y0, h_s_wallace_rca24_fa211_y2, h_s_wallace_rca24_fa211_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_17_y0(a_13, b_17, h_s_wallace_rca24_and_13_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_18_y0(a_12, b_18, h_s_wallace_rca24_and_12_18_y0);
  fa fa_h_s_wallace_rca24_fa212_y2(h_s_wallace_rca24_fa211_y4, h_s_wallace_rca24_and_13_17_y0, h_s_wallace_rca24_and_12_18_y0, h_s_wallace_rca24_fa212_y2, h_s_wallace_rca24_fa212_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_18_y0(a_13, b_18, h_s_wallace_rca24_and_13_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_19_y0(a_12, b_19, h_s_wallace_rca24_and_12_19_y0);
  fa fa_h_s_wallace_rca24_fa213_y2(h_s_wallace_rca24_fa212_y4, h_s_wallace_rca24_and_13_18_y0, h_s_wallace_rca24_and_12_19_y0, h_s_wallace_rca24_fa213_y2, h_s_wallace_rca24_fa213_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_19_y0(a_13, b_19, h_s_wallace_rca24_and_13_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_20_y0(a_12, b_20, h_s_wallace_rca24_and_12_20_y0);
  fa fa_h_s_wallace_rca24_fa214_y2(h_s_wallace_rca24_fa213_y4, h_s_wallace_rca24_and_13_19_y0, h_s_wallace_rca24_and_12_20_y0, h_s_wallace_rca24_fa214_y2, h_s_wallace_rca24_fa214_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_20_y0(a_13, b_20, h_s_wallace_rca24_and_13_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_21_y0(a_12, b_21, h_s_wallace_rca24_and_12_21_y0);
  fa fa_h_s_wallace_rca24_fa215_y2(h_s_wallace_rca24_fa214_y4, h_s_wallace_rca24_and_13_20_y0, h_s_wallace_rca24_and_12_21_y0, h_s_wallace_rca24_fa215_y2, h_s_wallace_rca24_fa215_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_21_y0(a_13, b_21, h_s_wallace_rca24_and_13_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_12_22_y0(a_12, b_22, h_s_wallace_rca24_and_12_22_y0);
  fa fa_h_s_wallace_rca24_fa216_y2(h_s_wallace_rca24_fa215_y4, h_s_wallace_rca24_and_13_21_y0, h_s_wallace_rca24_and_12_22_y0, h_s_wallace_rca24_fa216_y2, h_s_wallace_rca24_fa216_y4);
  and_gate and_gate_h_s_wallace_rca24_and_13_22_y0(a_13, b_22, h_s_wallace_rca24_and_13_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_12_23_y0(a_12, b_23, h_s_wallace_rca24_nand_12_23_y0);
  fa fa_h_s_wallace_rca24_fa217_y2(h_s_wallace_rca24_fa216_y4, h_s_wallace_rca24_and_13_22_y0, h_s_wallace_rca24_nand_12_23_y0, h_s_wallace_rca24_fa217_y2, h_s_wallace_rca24_fa217_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_13_23_y0(a_13, b_23, h_s_wallace_rca24_nand_13_23_y0);
  fa fa_h_s_wallace_rca24_fa218_y2(h_s_wallace_rca24_fa217_y4, h_s_wallace_rca24_nand_13_23_y0, h_s_wallace_rca24_fa33_y2, h_s_wallace_rca24_fa218_y2, h_s_wallace_rca24_fa218_y4);
  fa fa_h_s_wallace_rca24_fa219_y2(h_s_wallace_rca24_fa218_y4, h_s_wallace_rca24_fa34_y2, h_s_wallace_rca24_fa75_y2, h_s_wallace_rca24_fa219_y2, h_s_wallace_rca24_fa219_y4);
  fa fa_h_s_wallace_rca24_fa220_y2(h_s_wallace_rca24_fa219_y4, h_s_wallace_rca24_fa76_y2, h_s_wallace_rca24_fa115_y2, h_s_wallace_rca24_fa220_y2, h_s_wallace_rca24_fa220_y4);
  fa fa_h_s_wallace_rca24_fa221_y2(h_s_wallace_rca24_fa220_y4, h_s_wallace_rca24_fa116_y2, h_s_wallace_rca24_fa153_y2, h_s_wallace_rca24_fa221_y2, h_s_wallace_rca24_fa221_y4);
  ha ha_h_s_wallace_rca24_ha6_y0(h_s_wallace_rca24_fa122_y2, h_s_wallace_rca24_fa157_y2, h_s_wallace_rca24_ha6_y0, h_s_wallace_rca24_ha6_y1);
  fa fa_h_s_wallace_rca24_fa222_y2(h_s_wallace_rca24_ha6_y1, h_s_wallace_rca24_fa86_y2, h_s_wallace_rca24_fa123_y2, h_s_wallace_rca24_fa222_y2, h_s_wallace_rca24_fa222_y4);
  fa fa_h_s_wallace_rca24_fa223_y2(h_s_wallace_rca24_fa222_y4, h_s_wallace_rca24_fa48_y2, h_s_wallace_rca24_fa87_y2, h_s_wallace_rca24_fa223_y2, h_s_wallace_rca24_fa223_y4);
  fa fa_h_s_wallace_rca24_fa224_y2(h_s_wallace_rca24_fa223_y4, h_s_wallace_rca24_fa8_y2, h_s_wallace_rca24_fa49_y2, h_s_wallace_rca24_fa224_y2, h_s_wallace_rca24_fa224_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_12_y0(a_0, b_12, h_s_wallace_rca24_and_0_12_y0);
  fa fa_h_s_wallace_rca24_fa225_y2(h_s_wallace_rca24_fa224_y4, h_s_wallace_rca24_and_0_12_y0, h_s_wallace_rca24_fa9_y2, h_s_wallace_rca24_fa225_y2, h_s_wallace_rca24_fa225_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_12_y0(a_1, b_12, h_s_wallace_rca24_and_1_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_13_y0(a_0, b_13, h_s_wallace_rca24_and_0_13_y0);
  fa fa_h_s_wallace_rca24_fa226_y2(h_s_wallace_rca24_fa225_y4, h_s_wallace_rca24_and_1_12_y0, h_s_wallace_rca24_and_0_13_y0, h_s_wallace_rca24_fa226_y2, h_s_wallace_rca24_fa226_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_12_y0(a_2, b_12, h_s_wallace_rca24_and_2_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_13_y0(a_1, b_13, h_s_wallace_rca24_and_1_13_y0);
  fa fa_h_s_wallace_rca24_fa227_y2(h_s_wallace_rca24_fa226_y4, h_s_wallace_rca24_and_2_12_y0, h_s_wallace_rca24_and_1_13_y0, h_s_wallace_rca24_fa227_y2, h_s_wallace_rca24_fa227_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_12_y0(a_3, b_12, h_s_wallace_rca24_and_3_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_13_y0(a_2, b_13, h_s_wallace_rca24_and_2_13_y0);
  fa fa_h_s_wallace_rca24_fa228_y2(h_s_wallace_rca24_fa227_y4, h_s_wallace_rca24_and_3_12_y0, h_s_wallace_rca24_and_2_13_y0, h_s_wallace_rca24_fa228_y2, h_s_wallace_rca24_fa228_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_12_y0(a_4, b_12, h_s_wallace_rca24_and_4_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_13_y0(a_3, b_13, h_s_wallace_rca24_and_3_13_y0);
  fa fa_h_s_wallace_rca24_fa229_y2(h_s_wallace_rca24_fa228_y4, h_s_wallace_rca24_and_4_12_y0, h_s_wallace_rca24_and_3_13_y0, h_s_wallace_rca24_fa229_y2, h_s_wallace_rca24_fa229_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_12_y0(a_5, b_12, h_s_wallace_rca24_and_5_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_13_y0(a_4, b_13, h_s_wallace_rca24_and_4_13_y0);
  fa fa_h_s_wallace_rca24_fa230_y2(h_s_wallace_rca24_fa229_y4, h_s_wallace_rca24_and_5_12_y0, h_s_wallace_rca24_and_4_13_y0, h_s_wallace_rca24_fa230_y2, h_s_wallace_rca24_fa230_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_12_y0(a_6, b_12, h_s_wallace_rca24_and_6_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_13_y0(a_5, b_13, h_s_wallace_rca24_and_5_13_y0);
  fa fa_h_s_wallace_rca24_fa231_y2(h_s_wallace_rca24_fa230_y4, h_s_wallace_rca24_and_6_12_y0, h_s_wallace_rca24_and_5_13_y0, h_s_wallace_rca24_fa231_y2, h_s_wallace_rca24_fa231_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_12_y0(a_7, b_12, h_s_wallace_rca24_and_7_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_13_y0(a_6, b_13, h_s_wallace_rca24_and_6_13_y0);
  fa fa_h_s_wallace_rca24_fa232_y2(h_s_wallace_rca24_fa231_y4, h_s_wallace_rca24_and_7_12_y0, h_s_wallace_rca24_and_6_13_y0, h_s_wallace_rca24_fa232_y2, h_s_wallace_rca24_fa232_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_12_y0(a_8, b_12, h_s_wallace_rca24_and_8_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_13_y0(a_7, b_13, h_s_wallace_rca24_and_7_13_y0);
  fa fa_h_s_wallace_rca24_fa233_y2(h_s_wallace_rca24_fa232_y4, h_s_wallace_rca24_and_8_12_y0, h_s_wallace_rca24_and_7_13_y0, h_s_wallace_rca24_fa233_y2, h_s_wallace_rca24_fa233_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_12_y0(a_9, b_12, h_s_wallace_rca24_and_9_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_13_y0(a_8, b_13, h_s_wallace_rca24_and_8_13_y0);
  fa fa_h_s_wallace_rca24_fa234_y2(h_s_wallace_rca24_fa233_y4, h_s_wallace_rca24_and_9_12_y0, h_s_wallace_rca24_and_8_13_y0, h_s_wallace_rca24_fa234_y2, h_s_wallace_rca24_fa234_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_12_y0(a_10, b_12, h_s_wallace_rca24_and_10_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_13_y0(a_9, b_13, h_s_wallace_rca24_and_9_13_y0);
  fa fa_h_s_wallace_rca24_fa235_y2(h_s_wallace_rca24_fa234_y4, h_s_wallace_rca24_and_10_12_y0, h_s_wallace_rca24_and_9_13_y0, h_s_wallace_rca24_fa235_y2, h_s_wallace_rca24_fa235_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_12_y0(a_11, b_12, h_s_wallace_rca24_and_11_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_13_y0(a_10, b_13, h_s_wallace_rca24_and_10_13_y0);
  fa fa_h_s_wallace_rca24_fa236_y2(h_s_wallace_rca24_fa235_y4, h_s_wallace_rca24_and_11_12_y0, h_s_wallace_rca24_and_10_13_y0, h_s_wallace_rca24_fa236_y2, h_s_wallace_rca24_fa236_y4);
  and_gate and_gate_h_s_wallace_rca24_and_12_12_y0(a_12, b_12, h_s_wallace_rca24_and_12_12_y0);
  and_gate and_gate_h_s_wallace_rca24_and_11_13_y0(a_11, b_13, h_s_wallace_rca24_and_11_13_y0);
  fa fa_h_s_wallace_rca24_fa237_y2(h_s_wallace_rca24_fa236_y4, h_s_wallace_rca24_and_12_12_y0, h_s_wallace_rca24_and_11_13_y0, h_s_wallace_rca24_fa237_y2, h_s_wallace_rca24_fa237_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_14_y0(a_11, b_14, h_s_wallace_rca24_and_11_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_15_y0(a_10, b_15, h_s_wallace_rca24_and_10_15_y0);
  fa fa_h_s_wallace_rca24_fa238_y2(h_s_wallace_rca24_fa237_y4, h_s_wallace_rca24_and_11_14_y0, h_s_wallace_rca24_and_10_15_y0, h_s_wallace_rca24_fa238_y2, h_s_wallace_rca24_fa238_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_15_y0(a_11, b_15, h_s_wallace_rca24_and_11_15_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_16_y0(a_10, b_16, h_s_wallace_rca24_and_10_16_y0);
  fa fa_h_s_wallace_rca24_fa239_y2(h_s_wallace_rca24_fa238_y4, h_s_wallace_rca24_and_11_15_y0, h_s_wallace_rca24_and_10_16_y0, h_s_wallace_rca24_fa239_y2, h_s_wallace_rca24_fa239_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_16_y0(a_11, b_16, h_s_wallace_rca24_and_11_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_17_y0(a_10, b_17, h_s_wallace_rca24_and_10_17_y0);
  fa fa_h_s_wallace_rca24_fa240_y2(h_s_wallace_rca24_fa239_y4, h_s_wallace_rca24_and_11_16_y0, h_s_wallace_rca24_and_10_17_y0, h_s_wallace_rca24_fa240_y2, h_s_wallace_rca24_fa240_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_17_y0(a_11, b_17, h_s_wallace_rca24_and_11_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_18_y0(a_10, b_18, h_s_wallace_rca24_and_10_18_y0);
  fa fa_h_s_wallace_rca24_fa241_y2(h_s_wallace_rca24_fa240_y4, h_s_wallace_rca24_and_11_17_y0, h_s_wallace_rca24_and_10_18_y0, h_s_wallace_rca24_fa241_y2, h_s_wallace_rca24_fa241_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_18_y0(a_11, b_18, h_s_wallace_rca24_and_11_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_19_y0(a_10, b_19, h_s_wallace_rca24_and_10_19_y0);
  fa fa_h_s_wallace_rca24_fa242_y2(h_s_wallace_rca24_fa241_y4, h_s_wallace_rca24_and_11_18_y0, h_s_wallace_rca24_and_10_19_y0, h_s_wallace_rca24_fa242_y2, h_s_wallace_rca24_fa242_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_19_y0(a_11, b_19, h_s_wallace_rca24_and_11_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_20_y0(a_10, b_20, h_s_wallace_rca24_and_10_20_y0);
  fa fa_h_s_wallace_rca24_fa243_y2(h_s_wallace_rca24_fa242_y4, h_s_wallace_rca24_and_11_19_y0, h_s_wallace_rca24_and_10_20_y0, h_s_wallace_rca24_fa243_y2, h_s_wallace_rca24_fa243_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_20_y0(a_11, b_20, h_s_wallace_rca24_and_11_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_21_y0(a_10, b_21, h_s_wallace_rca24_and_10_21_y0);
  fa fa_h_s_wallace_rca24_fa244_y2(h_s_wallace_rca24_fa243_y4, h_s_wallace_rca24_and_11_20_y0, h_s_wallace_rca24_and_10_21_y0, h_s_wallace_rca24_fa244_y2, h_s_wallace_rca24_fa244_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_21_y0(a_11, b_21, h_s_wallace_rca24_and_11_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_10_22_y0(a_10, b_22, h_s_wallace_rca24_and_10_22_y0);
  fa fa_h_s_wallace_rca24_fa245_y2(h_s_wallace_rca24_fa244_y4, h_s_wallace_rca24_and_11_21_y0, h_s_wallace_rca24_and_10_22_y0, h_s_wallace_rca24_fa245_y2, h_s_wallace_rca24_fa245_y4);
  and_gate and_gate_h_s_wallace_rca24_and_11_22_y0(a_11, b_22, h_s_wallace_rca24_and_11_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_10_23_y0(a_10, b_23, h_s_wallace_rca24_nand_10_23_y0);
  fa fa_h_s_wallace_rca24_fa246_y2(h_s_wallace_rca24_fa245_y4, h_s_wallace_rca24_and_11_22_y0, h_s_wallace_rca24_nand_10_23_y0, h_s_wallace_rca24_fa246_y2, h_s_wallace_rca24_fa246_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_11_23_y0(a_11, b_23, h_s_wallace_rca24_nand_11_23_y0);
  fa fa_h_s_wallace_rca24_fa247_y2(h_s_wallace_rca24_fa246_y4, h_s_wallace_rca24_nand_11_23_y0, h_s_wallace_rca24_fa31_y2, h_s_wallace_rca24_fa247_y2, h_s_wallace_rca24_fa247_y4);
  fa fa_h_s_wallace_rca24_fa248_y2(h_s_wallace_rca24_fa247_y4, h_s_wallace_rca24_fa32_y2, h_s_wallace_rca24_fa73_y2, h_s_wallace_rca24_fa248_y2, h_s_wallace_rca24_fa248_y4);
  fa fa_h_s_wallace_rca24_fa249_y2(h_s_wallace_rca24_fa248_y4, h_s_wallace_rca24_fa74_y2, h_s_wallace_rca24_fa113_y2, h_s_wallace_rca24_fa249_y2, h_s_wallace_rca24_fa249_y4);
  fa fa_h_s_wallace_rca24_fa250_y2(h_s_wallace_rca24_fa249_y4, h_s_wallace_rca24_fa114_y2, h_s_wallace_rca24_fa151_y2, h_s_wallace_rca24_fa250_y2, h_s_wallace_rca24_fa250_y4);
  fa fa_h_s_wallace_rca24_fa251_y2(h_s_wallace_rca24_fa250_y4, h_s_wallace_rca24_fa152_y2, h_s_wallace_rca24_fa187_y2, h_s_wallace_rca24_fa251_y2, h_s_wallace_rca24_fa251_y4);
  ha ha_h_s_wallace_rca24_ha7_y0(h_s_wallace_rca24_fa158_y2, h_s_wallace_rca24_fa191_y2, h_s_wallace_rca24_ha7_y0, h_s_wallace_rca24_ha7_y1);
  fa fa_h_s_wallace_rca24_fa252_y2(h_s_wallace_rca24_ha7_y1, h_s_wallace_rca24_fa124_y2, h_s_wallace_rca24_fa159_y2, h_s_wallace_rca24_fa252_y2, h_s_wallace_rca24_fa252_y4);
  fa fa_h_s_wallace_rca24_fa253_y2(h_s_wallace_rca24_fa252_y4, h_s_wallace_rca24_fa88_y2, h_s_wallace_rca24_fa125_y2, h_s_wallace_rca24_fa253_y2, h_s_wallace_rca24_fa253_y4);
  fa fa_h_s_wallace_rca24_fa254_y2(h_s_wallace_rca24_fa253_y4, h_s_wallace_rca24_fa50_y2, h_s_wallace_rca24_fa89_y2, h_s_wallace_rca24_fa254_y2, h_s_wallace_rca24_fa254_y4);
  fa fa_h_s_wallace_rca24_fa255_y2(h_s_wallace_rca24_fa254_y4, h_s_wallace_rca24_fa10_y2, h_s_wallace_rca24_fa51_y2, h_s_wallace_rca24_fa255_y2, h_s_wallace_rca24_fa255_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_14_y0(a_0, b_14, h_s_wallace_rca24_and_0_14_y0);
  fa fa_h_s_wallace_rca24_fa256_y2(h_s_wallace_rca24_fa255_y4, h_s_wallace_rca24_and_0_14_y0, h_s_wallace_rca24_fa11_y2, h_s_wallace_rca24_fa256_y2, h_s_wallace_rca24_fa256_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_14_y0(a_1, b_14, h_s_wallace_rca24_and_1_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_15_y0(a_0, b_15, h_s_wallace_rca24_and_0_15_y0);
  fa fa_h_s_wallace_rca24_fa257_y2(h_s_wallace_rca24_fa256_y4, h_s_wallace_rca24_and_1_14_y0, h_s_wallace_rca24_and_0_15_y0, h_s_wallace_rca24_fa257_y2, h_s_wallace_rca24_fa257_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_14_y0(a_2, b_14, h_s_wallace_rca24_and_2_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_15_y0(a_1, b_15, h_s_wallace_rca24_and_1_15_y0);
  fa fa_h_s_wallace_rca24_fa258_y2(h_s_wallace_rca24_fa257_y4, h_s_wallace_rca24_and_2_14_y0, h_s_wallace_rca24_and_1_15_y0, h_s_wallace_rca24_fa258_y2, h_s_wallace_rca24_fa258_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_14_y0(a_3, b_14, h_s_wallace_rca24_and_3_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_15_y0(a_2, b_15, h_s_wallace_rca24_and_2_15_y0);
  fa fa_h_s_wallace_rca24_fa259_y2(h_s_wallace_rca24_fa258_y4, h_s_wallace_rca24_and_3_14_y0, h_s_wallace_rca24_and_2_15_y0, h_s_wallace_rca24_fa259_y2, h_s_wallace_rca24_fa259_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_14_y0(a_4, b_14, h_s_wallace_rca24_and_4_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_15_y0(a_3, b_15, h_s_wallace_rca24_and_3_15_y0);
  fa fa_h_s_wallace_rca24_fa260_y2(h_s_wallace_rca24_fa259_y4, h_s_wallace_rca24_and_4_14_y0, h_s_wallace_rca24_and_3_15_y0, h_s_wallace_rca24_fa260_y2, h_s_wallace_rca24_fa260_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_14_y0(a_5, b_14, h_s_wallace_rca24_and_5_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_15_y0(a_4, b_15, h_s_wallace_rca24_and_4_15_y0);
  fa fa_h_s_wallace_rca24_fa261_y2(h_s_wallace_rca24_fa260_y4, h_s_wallace_rca24_and_5_14_y0, h_s_wallace_rca24_and_4_15_y0, h_s_wallace_rca24_fa261_y2, h_s_wallace_rca24_fa261_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_14_y0(a_6, b_14, h_s_wallace_rca24_and_6_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_15_y0(a_5, b_15, h_s_wallace_rca24_and_5_15_y0);
  fa fa_h_s_wallace_rca24_fa262_y2(h_s_wallace_rca24_fa261_y4, h_s_wallace_rca24_and_6_14_y0, h_s_wallace_rca24_and_5_15_y0, h_s_wallace_rca24_fa262_y2, h_s_wallace_rca24_fa262_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_14_y0(a_7, b_14, h_s_wallace_rca24_and_7_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_15_y0(a_6, b_15, h_s_wallace_rca24_and_6_15_y0);
  fa fa_h_s_wallace_rca24_fa263_y2(h_s_wallace_rca24_fa262_y4, h_s_wallace_rca24_and_7_14_y0, h_s_wallace_rca24_and_6_15_y0, h_s_wallace_rca24_fa263_y2, h_s_wallace_rca24_fa263_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_14_y0(a_8, b_14, h_s_wallace_rca24_and_8_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_15_y0(a_7, b_15, h_s_wallace_rca24_and_7_15_y0);
  fa fa_h_s_wallace_rca24_fa264_y2(h_s_wallace_rca24_fa263_y4, h_s_wallace_rca24_and_8_14_y0, h_s_wallace_rca24_and_7_15_y0, h_s_wallace_rca24_fa264_y2, h_s_wallace_rca24_fa264_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_14_y0(a_9, b_14, h_s_wallace_rca24_and_9_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_15_y0(a_8, b_15, h_s_wallace_rca24_and_8_15_y0);
  fa fa_h_s_wallace_rca24_fa265_y2(h_s_wallace_rca24_fa264_y4, h_s_wallace_rca24_and_9_14_y0, h_s_wallace_rca24_and_8_15_y0, h_s_wallace_rca24_fa265_y2, h_s_wallace_rca24_fa265_y4);
  and_gate and_gate_h_s_wallace_rca24_and_10_14_y0(a_10, b_14, h_s_wallace_rca24_and_10_14_y0);
  and_gate and_gate_h_s_wallace_rca24_and_9_15_y0(a_9, b_15, h_s_wallace_rca24_and_9_15_y0);
  fa fa_h_s_wallace_rca24_fa266_y2(h_s_wallace_rca24_fa265_y4, h_s_wallace_rca24_and_10_14_y0, h_s_wallace_rca24_and_9_15_y0, h_s_wallace_rca24_fa266_y2, h_s_wallace_rca24_fa266_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_16_y0(a_9, b_16, h_s_wallace_rca24_and_9_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_17_y0(a_8, b_17, h_s_wallace_rca24_and_8_17_y0);
  fa fa_h_s_wallace_rca24_fa267_y2(h_s_wallace_rca24_fa266_y4, h_s_wallace_rca24_and_9_16_y0, h_s_wallace_rca24_and_8_17_y0, h_s_wallace_rca24_fa267_y2, h_s_wallace_rca24_fa267_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_17_y0(a_9, b_17, h_s_wallace_rca24_and_9_17_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_18_y0(a_8, b_18, h_s_wallace_rca24_and_8_18_y0);
  fa fa_h_s_wallace_rca24_fa268_y2(h_s_wallace_rca24_fa267_y4, h_s_wallace_rca24_and_9_17_y0, h_s_wallace_rca24_and_8_18_y0, h_s_wallace_rca24_fa268_y2, h_s_wallace_rca24_fa268_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_18_y0(a_9, b_18, h_s_wallace_rca24_and_9_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_19_y0(a_8, b_19, h_s_wallace_rca24_and_8_19_y0);
  fa fa_h_s_wallace_rca24_fa269_y2(h_s_wallace_rca24_fa268_y4, h_s_wallace_rca24_and_9_18_y0, h_s_wallace_rca24_and_8_19_y0, h_s_wallace_rca24_fa269_y2, h_s_wallace_rca24_fa269_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_19_y0(a_9, b_19, h_s_wallace_rca24_and_9_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_20_y0(a_8, b_20, h_s_wallace_rca24_and_8_20_y0);
  fa fa_h_s_wallace_rca24_fa270_y2(h_s_wallace_rca24_fa269_y4, h_s_wallace_rca24_and_9_19_y0, h_s_wallace_rca24_and_8_20_y0, h_s_wallace_rca24_fa270_y2, h_s_wallace_rca24_fa270_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_20_y0(a_9, b_20, h_s_wallace_rca24_and_9_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_21_y0(a_8, b_21, h_s_wallace_rca24_and_8_21_y0);
  fa fa_h_s_wallace_rca24_fa271_y2(h_s_wallace_rca24_fa270_y4, h_s_wallace_rca24_and_9_20_y0, h_s_wallace_rca24_and_8_21_y0, h_s_wallace_rca24_fa271_y2, h_s_wallace_rca24_fa271_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_21_y0(a_9, b_21, h_s_wallace_rca24_and_9_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_8_22_y0(a_8, b_22, h_s_wallace_rca24_and_8_22_y0);
  fa fa_h_s_wallace_rca24_fa272_y2(h_s_wallace_rca24_fa271_y4, h_s_wallace_rca24_and_9_21_y0, h_s_wallace_rca24_and_8_22_y0, h_s_wallace_rca24_fa272_y2, h_s_wallace_rca24_fa272_y4);
  and_gate and_gate_h_s_wallace_rca24_and_9_22_y0(a_9, b_22, h_s_wallace_rca24_and_9_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_8_23_y0(a_8, b_23, h_s_wallace_rca24_nand_8_23_y0);
  fa fa_h_s_wallace_rca24_fa273_y2(h_s_wallace_rca24_fa272_y4, h_s_wallace_rca24_and_9_22_y0, h_s_wallace_rca24_nand_8_23_y0, h_s_wallace_rca24_fa273_y2, h_s_wallace_rca24_fa273_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_9_23_y0(a_9, b_23, h_s_wallace_rca24_nand_9_23_y0);
  fa fa_h_s_wallace_rca24_fa274_y2(h_s_wallace_rca24_fa273_y4, h_s_wallace_rca24_nand_9_23_y0, h_s_wallace_rca24_fa29_y2, h_s_wallace_rca24_fa274_y2, h_s_wallace_rca24_fa274_y4);
  fa fa_h_s_wallace_rca24_fa275_y2(h_s_wallace_rca24_fa274_y4, h_s_wallace_rca24_fa30_y2, h_s_wallace_rca24_fa71_y2, h_s_wallace_rca24_fa275_y2, h_s_wallace_rca24_fa275_y4);
  fa fa_h_s_wallace_rca24_fa276_y2(h_s_wallace_rca24_fa275_y4, h_s_wallace_rca24_fa72_y2, h_s_wallace_rca24_fa111_y2, h_s_wallace_rca24_fa276_y2, h_s_wallace_rca24_fa276_y4);
  fa fa_h_s_wallace_rca24_fa277_y2(h_s_wallace_rca24_fa276_y4, h_s_wallace_rca24_fa112_y2, h_s_wallace_rca24_fa149_y2, h_s_wallace_rca24_fa277_y2, h_s_wallace_rca24_fa277_y4);
  fa fa_h_s_wallace_rca24_fa278_y2(h_s_wallace_rca24_fa277_y4, h_s_wallace_rca24_fa150_y2, h_s_wallace_rca24_fa185_y2, h_s_wallace_rca24_fa278_y2, h_s_wallace_rca24_fa278_y4);
  fa fa_h_s_wallace_rca24_fa279_y2(h_s_wallace_rca24_fa278_y4, h_s_wallace_rca24_fa186_y2, h_s_wallace_rca24_fa219_y2, h_s_wallace_rca24_fa279_y2, h_s_wallace_rca24_fa279_y4);
  ha ha_h_s_wallace_rca24_ha8_y0(h_s_wallace_rca24_fa192_y2, h_s_wallace_rca24_fa223_y2, h_s_wallace_rca24_ha8_y0, h_s_wallace_rca24_ha8_y1);
  fa fa_h_s_wallace_rca24_fa280_y2(h_s_wallace_rca24_ha8_y1, h_s_wallace_rca24_fa160_y2, h_s_wallace_rca24_fa193_y2, h_s_wallace_rca24_fa280_y2, h_s_wallace_rca24_fa280_y4);
  fa fa_h_s_wallace_rca24_fa281_y2(h_s_wallace_rca24_fa280_y4, h_s_wallace_rca24_fa126_y2, h_s_wallace_rca24_fa161_y2, h_s_wallace_rca24_fa281_y2, h_s_wallace_rca24_fa281_y4);
  fa fa_h_s_wallace_rca24_fa282_y2(h_s_wallace_rca24_fa281_y4, h_s_wallace_rca24_fa90_y2, h_s_wallace_rca24_fa127_y2, h_s_wallace_rca24_fa282_y2, h_s_wallace_rca24_fa282_y4);
  fa fa_h_s_wallace_rca24_fa283_y2(h_s_wallace_rca24_fa282_y4, h_s_wallace_rca24_fa52_y2, h_s_wallace_rca24_fa91_y2, h_s_wallace_rca24_fa283_y2, h_s_wallace_rca24_fa283_y4);
  fa fa_h_s_wallace_rca24_fa284_y2(h_s_wallace_rca24_fa283_y4, h_s_wallace_rca24_fa12_y2, h_s_wallace_rca24_fa53_y2, h_s_wallace_rca24_fa284_y2, h_s_wallace_rca24_fa284_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_16_y0(a_0, b_16, h_s_wallace_rca24_and_0_16_y0);
  fa fa_h_s_wallace_rca24_fa285_y2(h_s_wallace_rca24_fa284_y4, h_s_wallace_rca24_and_0_16_y0, h_s_wallace_rca24_fa13_y2, h_s_wallace_rca24_fa285_y2, h_s_wallace_rca24_fa285_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_16_y0(a_1, b_16, h_s_wallace_rca24_and_1_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_17_y0(a_0, b_17, h_s_wallace_rca24_and_0_17_y0);
  fa fa_h_s_wallace_rca24_fa286_y2(h_s_wallace_rca24_fa285_y4, h_s_wallace_rca24_and_1_16_y0, h_s_wallace_rca24_and_0_17_y0, h_s_wallace_rca24_fa286_y2, h_s_wallace_rca24_fa286_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_16_y0(a_2, b_16, h_s_wallace_rca24_and_2_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_17_y0(a_1, b_17, h_s_wallace_rca24_and_1_17_y0);
  fa fa_h_s_wallace_rca24_fa287_y2(h_s_wallace_rca24_fa286_y4, h_s_wallace_rca24_and_2_16_y0, h_s_wallace_rca24_and_1_17_y0, h_s_wallace_rca24_fa287_y2, h_s_wallace_rca24_fa287_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_16_y0(a_3, b_16, h_s_wallace_rca24_and_3_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_17_y0(a_2, b_17, h_s_wallace_rca24_and_2_17_y0);
  fa fa_h_s_wallace_rca24_fa288_y2(h_s_wallace_rca24_fa287_y4, h_s_wallace_rca24_and_3_16_y0, h_s_wallace_rca24_and_2_17_y0, h_s_wallace_rca24_fa288_y2, h_s_wallace_rca24_fa288_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_16_y0(a_4, b_16, h_s_wallace_rca24_and_4_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_17_y0(a_3, b_17, h_s_wallace_rca24_and_3_17_y0);
  fa fa_h_s_wallace_rca24_fa289_y2(h_s_wallace_rca24_fa288_y4, h_s_wallace_rca24_and_4_16_y0, h_s_wallace_rca24_and_3_17_y0, h_s_wallace_rca24_fa289_y2, h_s_wallace_rca24_fa289_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_16_y0(a_5, b_16, h_s_wallace_rca24_and_5_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_17_y0(a_4, b_17, h_s_wallace_rca24_and_4_17_y0);
  fa fa_h_s_wallace_rca24_fa290_y2(h_s_wallace_rca24_fa289_y4, h_s_wallace_rca24_and_5_16_y0, h_s_wallace_rca24_and_4_17_y0, h_s_wallace_rca24_fa290_y2, h_s_wallace_rca24_fa290_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_16_y0(a_6, b_16, h_s_wallace_rca24_and_6_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_17_y0(a_5, b_17, h_s_wallace_rca24_and_5_17_y0);
  fa fa_h_s_wallace_rca24_fa291_y2(h_s_wallace_rca24_fa290_y4, h_s_wallace_rca24_and_6_16_y0, h_s_wallace_rca24_and_5_17_y0, h_s_wallace_rca24_fa291_y2, h_s_wallace_rca24_fa291_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_16_y0(a_7, b_16, h_s_wallace_rca24_and_7_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_17_y0(a_6, b_17, h_s_wallace_rca24_and_6_17_y0);
  fa fa_h_s_wallace_rca24_fa292_y2(h_s_wallace_rca24_fa291_y4, h_s_wallace_rca24_and_7_16_y0, h_s_wallace_rca24_and_6_17_y0, h_s_wallace_rca24_fa292_y2, h_s_wallace_rca24_fa292_y4);
  and_gate and_gate_h_s_wallace_rca24_and_8_16_y0(a_8, b_16, h_s_wallace_rca24_and_8_16_y0);
  and_gate and_gate_h_s_wallace_rca24_and_7_17_y0(a_7, b_17, h_s_wallace_rca24_and_7_17_y0);
  fa fa_h_s_wallace_rca24_fa293_y2(h_s_wallace_rca24_fa292_y4, h_s_wallace_rca24_and_8_16_y0, h_s_wallace_rca24_and_7_17_y0, h_s_wallace_rca24_fa293_y2, h_s_wallace_rca24_fa293_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_18_y0(a_7, b_18, h_s_wallace_rca24_and_7_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_19_y0(a_6, b_19, h_s_wallace_rca24_and_6_19_y0);
  fa fa_h_s_wallace_rca24_fa294_y2(h_s_wallace_rca24_fa293_y4, h_s_wallace_rca24_and_7_18_y0, h_s_wallace_rca24_and_6_19_y0, h_s_wallace_rca24_fa294_y2, h_s_wallace_rca24_fa294_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_19_y0(a_7, b_19, h_s_wallace_rca24_and_7_19_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_20_y0(a_6, b_20, h_s_wallace_rca24_and_6_20_y0);
  fa fa_h_s_wallace_rca24_fa295_y2(h_s_wallace_rca24_fa294_y4, h_s_wallace_rca24_and_7_19_y0, h_s_wallace_rca24_and_6_20_y0, h_s_wallace_rca24_fa295_y2, h_s_wallace_rca24_fa295_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_20_y0(a_7, b_20, h_s_wallace_rca24_and_7_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_21_y0(a_6, b_21, h_s_wallace_rca24_and_6_21_y0);
  fa fa_h_s_wallace_rca24_fa296_y2(h_s_wallace_rca24_fa295_y4, h_s_wallace_rca24_and_7_20_y0, h_s_wallace_rca24_and_6_21_y0, h_s_wallace_rca24_fa296_y2, h_s_wallace_rca24_fa296_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_21_y0(a_7, b_21, h_s_wallace_rca24_and_7_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_6_22_y0(a_6, b_22, h_s_wallace_rca24_and_6_22_y0);
  fa fa_h_s_wallace_rca24_fa297_y2(h_s_wallace_rca24_fa296_y4, h_s_wallace_rca24_and_7_21_y0, h_s_wallace_rca24_and_6_22_y0, h_s_wallace_rca24_fa297_y2, h_s_wallace_rca24_fa297_y4);
  and_gate and_gate_h_s_wallace_rca24_and_7_22_y0(a_7, b_22, h_s_wallace_rca24_and_7_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_6_23_y0(a_6, b_23, h_s_wallace_rca24_nand_6_23_y0);
  fa fa_h_s_wallace_rca24_fa298_y2(h_s_wallace_rca24_fa297_y4, h_s_wallace_rca24_and_7_22_y0, h_s_wallace_rca24_nand_6_23_y0, h_s_wallace_rca24_fa298_y2, h_s_wallace_rca24_fa298_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_7_23_y0(a_7, b_23, h_s_wallace_rca24_nand_7_23_y0);
  fa fa_h_s_wallace_rca24_fa299_y2(h_s_wallace_rca24_fa298_y4, h_s_wallace_rca24_nand_7_23_y0, h_s_wallace_rca24_fa27_y2, h_s_wallace_rca24_fa299_y2, h_s_wallace_rca24_fa299_y4);
  fa fa_h_s_wallace_rca24_fa300_y2(h_s_wallace_rca24_fa299_y4, h_s_wallace_rca24_fa28_y2, h_s_wallace_rca24_fa69_y2, h_s_wallace_rca24_fa300_y2, h_s_wallace_rca24_fa300_y4);
  fa fa_h_s_wallace_rca24_fa301_y2(h_s_wallace_rca24_fa300_y4, h_s_wallace_rca24_fa70_y2, h_s_wallace_rca24_fa109_y2, h_s_wallace_rca24_fa301_y2, h_s_wallace_rca24_fa301_y4);
  fa fa_h_s_wallace_rca24_fa302_y2(h_s_wallace_rca24_fa301_y4, h_s_wallace_rca24_fa110_y2, h_s_wallace_rca24_fa147_y2, h_s_wallace_rca24_fa302_y2, h_s_wallace_rca24_fa302_y4);
  fa fa_h_s_wallace_rca24_fa303_y2(h_s_wallace_rca24_fa302_y4, h_s_wallace_rca24_fa148_y2, h_s_wallace_rca24_fa183_y2, h_s_wallace_rca24_fa303_y2, h_s_wallace_rca24_fa303_y4);
  fa fa_h_s_wallace_rca24_fa304_y2(h_s_wallace_rca24_fa303_y4, h_s_wallace_rca24_fa184_y2, h_s_wallace_rca24_fa217_y2, h_s_wallace_rca24_fa304_y2, h_s_wallace_rca24_fa304_y4);
  fa fa_h_s_wallace_rca24_fa305_y2(h_s_wallace_rca24_fa304_y4, h_s_wallace_rca24_fa218_y2, h_s_wallace_rca24_fa249_y2, h_s_wallace_rca24_fa305_y2, h_s_wallace_rca24_fa305_y4);
  ha ha_h_s_wallace_rca24_ha9_y0(h_s_wallace_rca24_fa224_y2, h_s_wallace_rca24_fa253_y2, h_s_wallace_rca24_ha9_y0, h_s_wallace_rca24_ha9_y1);
  fa fa_h_s_wallace_rca24_fa306_y2(h_s_wallace_rca24_ha9_y1, h_s_wallace_rca24_fa194_y2, h_s_wallace_rca24_fa225_y2, h_s_wallace_rca24_fa306_y2, h_s_wallace_rca24_fa306_y4);
  fa fa_h_s_wallace_rca24_fa307_y2(h_s_wallace_rca24_fa306_y4, h_s_wallace_rca24_fa162_y2, h_s_wallace_rca24_fa195_y2, h_s_wallace_rca24_fa307_y2, h_s_wallace_rca24_fa307_y4);
  fa fa_h_s_wallace_rca24_fa308_y2(h_s_wallace_rca24_fa307_y4, h_s_wallace_rca24_fa128_y2, h_s_wallace_rca24_fa163_y2, h_s_wallace_rca24_fa308_y2, h_s_wallace_rca24_fa308_y4);
  fa fa_h_s_wallace_rca24_fa309_y2(h_s_wallace_rca24_fa308_y4, h_s_wallace_rca24_fa92_y2, h_s_wallace_rca24_fa129_y2, h_s_wallace_rca24_fa309_y2, h_s_wallace_rca24_fa309_y4);
  fa fa_h_s_wallace_rca24_fa310_y2(h_s_wallace_rca24_fa309_y4, h_s_wallace_rca24_fa54_y2, h_s_wallace_rca24_fa93_y2, h_s_wallace_rca24_fa310_y2, h_s_wallace_rca24_fa310_y4);
  fa fa_h_s_wallace_rca24_fa311_y2(h_s_wallace_rca24_fa310_y4, h_s_wallace_rca24_fa14_y2, h_s_wallace_rca24_fa55_y2, h_s_wallace_rca24_fa311_y2, h_s_wallace_rca24_fa311_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_18_y0(a_0, b_18, h_s_wallace_rca24_and_0_18_y0);
  fa fa_h_s_wallace_rca24_fa312_y2(h_s_wallace_rca24_fa311_y4, h_s_wallace_rca24_and_0_18_y0, h_s_wallace_rca24_fa15_y2, h_s_wallace_rca24_fa312_y2, h_s_wallace_rca24_fa312_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_18_y0(a_1, b_18, h_s_wallace_rca24_and_1_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_19_y0(a_0, b_19, h_s_wallace_rca24_and_0_19_y0);
  fa fa_h_s_wallace_rca24_fa313_y2(h_s_wallace_rca24_fa312_y4, h_s_wallace_rca24_and_1_18_y0, h_s_wallace_rca24_and_0_19_y0, h_s_wallace_rca24_fa313_y2, h_s_wallace_rca24_fa313_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_18_y0(a_2, b_18, h_s_wallace_rca24_and_2_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_19_y0(a_1, b_19, h_s_wallace_rca24_and_1_19_y0);
  fa fa_h_s_wallace_rca24_fa314_y2(h_s_wallace_rca24_fa313_y4, h_s_wallace_rca24_and_2_18_y0, h_s_wallace_rca24_and_1_19_y0, h_s_wallace_rca24_fa314_y2, h_s_wallace_rca24_fa314_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_18_y0(a_3, b_18, h_s_wallace_rca24_and_3_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_19_y0(a_2, b_19, h_s_wallace_rca24_and_2_19_y0);
  fa fa_h_s_wallace_rca24_fa315_y2(h_s_wallace_rca24_fa314_y4, h_s_wallace_rca24_and_3_18_y0, h_s_wallace_rca24_and_2_19_y0, h_s_wallace_rca24_fa315_y2, h_s_wallace_rca24_fa315_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_18_y0(a_4, b_18, h_s_wallace_rca24_and_4_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_19_y0(a_3, b_19, h_s_wallace_rca24_and_3_19_y0);
  fa fa_h_s_wallace_rca24_fa316_y2(h_s_wallace_rca24_fa315_y4, h_s_wallace_rca24_and_4_18_y0, h_s_wallace_rca24_and_3_19_y0, h_s_wallace_rca24_fa316_y2, h_s_wallace_rca24_fa316_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_18_y0(a_5, b_18, h_s_wallace_rca24_and_5_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_19_y0(a_4, b_19, h_s_wallace_rca24_and_4_19_y0);
  fa fa_h_s_wallace_rca24_fa317_y2(h_s_wallace_rca24_fa316_y4, h_s_wallace_rca24_and_5_18_y0, h_s_wallace_rca24_and_4_19_y0, h_s_wallace_rca24_fa317_y2, h_s_wallace_rca24_fa317_y4);
  and_gate and_gate_h_s_wallace_rca24_and_6_18_y0(a_6, b_18, h_s_wallace_rca24_and_6_18_y0);
  and_gate and_gate_h_s_wallace_rca24_and_5_19_y0(a_5, b_19, h_s_wallace_rca24_and_5_19_y0);
  fa fa_h_s_wallace_rca24_fa318_y2(h_s_wallace_rca24_fa317_y4, h_s_wallace_rca24_and_6_18_y0, h_s_wallace_rca24_and_5_19_y0, h_s_wallace_rca24_fa318_y2, h_s_wallace_rca24_fa318_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_20_y0(a_5, b_20, h_s_wallace_rca24_and_5_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_21_y0(a_4, b_21, h_s_wallace_rca24_and_4_21_y0);
  fa fa_h_s_wallace_rca24_fa319_y2(h_s_wallace_rca24_fa318_y4, h_s_wallace_rca24_and_5_20_y0, h_s_wallace_rca24_and_4_21_y0, h_s_wallace_rca24_fa319_y2, h_s_wallace_rca24_fa319_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_21_y0(a_5, b_21, h_s_wallace_rca24_and_5_21_y0);
  and_gate and_gate_h_s_wallace_rca24_and_4_22_y0(a_4, b_22, h_s_wallace_rca24_and_4_22_y0);
  fa fa_h_s_wallace_rca24_fa320_y2(h_s_wallace_rca24_fa319_y4, h_s_wallace_rca24_and_5_21_y0, h_s_wallace_rca24_and_4_22_y0, h_s_wallace_rca24_fa320_y2, h_s_wallace_rca24_fa320_y4);
  and_gate and_gate_h_s_wallace_rca24_and_5_22_y0(a_5, b_22, h_s_wallace_rca24_and_5_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_4_23_y0(a_4, b_23, h_s_wallace_rca24_nand_4_23_y0);
  fa fa_h_s_wallace_rca24_fa321_y2(h_s_wallace_rca24_fa320_y4, h_s_wallace_rca24_and_5_22_y0, h_s_wallace_rca24_nand_4_23_y0, h_s_wallace_rca24_fa321_y2, h_s_wallace_rca24_fa321_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_5_23_y0(a_5, b_23, h_s_wallace_rca24_nand_5_23_y0);
  fa fa_h_s_wallace_rca24_fa322_y2(h_s_wallace_rca24_fa321_y4, h_s_wallace_rca24_nand_5_23_y0, h_s_wallace_rca24_fa25_y2, h_s_wallace_rca24_fa322_y2, h_s_wallace_rca24_fa322_y4);
  fa fa_h_s_wallace_rca24_fa323_y2(h_s_wallace_rca24_fa322_y4, h_s_wallace_rca24_fa26_y2, h_s_wallace_rca24_fa67_y2, h_s_wallace_rca24_fa323_y2, h_s_wallace_rca24_fa323_y4);
  fa fa_h_s_wallace_rca24_fa324_y2(h_s_wallace_rca24_fa323_y4, h_s_wallace_rca24_fa68_y2, h_s_wallace_rca24_fa107_y2, h_s_wallace_rca24_fa324_y2, h_s_wallace_rca24_fa324_y4);
  fa fa_h_s_wallace_rca24_fa325_y2(h_s_wallace_rca24_fa324_y4, h_s_wallace_rca24_fa108_y2, h_s_wallace_rca24_fa145_y2, h_s_wallace_rca24_fa325_y2, h_s_wallace_rca24_fa325_y4);
  fa fa_h_s_wallace_rca24_fa326_y2(h_s_wallace_rca24_fa325_y4, h_s_wallace_rca24_fa146_y2, h_s_wallace_rca24_fa181_y2, h_s_wallace_rca24_fa326_y2, h_s_wallace_rca24_fa326_y4);
  fa fa_h_s_wallace_rca24_fa327_y2(h_s_wallace_rca24_fa326_y4, h_s_wallace_rca24_fa182_y2, h_s_wallace_rca24_fa215_y2, h_s_wallace_rca24_fa327_y2, h_s_wallace_rca24_fa327_y4);
  fa fa_h_s_wallace_rca24_fa328_y2(h_s_wallace_rca24_fa327_y4, h_s_wallace_rca24_fa216_y2, h_s_wallace_rca24_fa247_y2, h_s_wallace_rca24_fa328_y2, h_s_wallace_rca24_fa328_y4);
  fa fa_h_s_wallace_rca24_fa329_y2(h_s_wallace_rca24_fa328_y4, h_s_wallace_rca24_fa248_y2, h_s_wallace_rca24_fa277_y2, h_s_wallace_rca24_fa329_y2, h_s_wallace_rca24_fa329_y4);
  ha ha_h_s_wallace_rca24_ha10_y0(h_s_wallace_rca24_fa254_y2, h_s_wallace_rca24_fa281_y2, h_s_wallace_rca24_ha10_y0, h_s_wallace_rca24_ha10_y1);
  fa fa_h_s_wallace_rca24_fa330_y2(h_s_wallace_rca24_ha10_y1, h_s_wallace_rca24_fa226_y2, h_s_wallace_rca24_fa255_y2, h_s_wallace_rca24_fa330_y2, h_s_wallace_rca24_fa330_y4);
  fa fa_h_s_wallace_rca24_fa331_y2(h_s_wallace_rca24_fa330_y4, h_s_wallace_rca24_fa196_y2, h_s_wallace_rca24_fa227_y2, h_s_wallace_rca24_fa331_y2, h_s_wallace_rca24_fa331_y4);
  fa fa_h_s_wallace_rca24_fa332_y2(h_s_wallace_rca24_fa331_y4, h_s_wallace_rca24_fa164_y2, h_s_wallace_rca24_fa197_y2, h_s_wallace_rca24_fa332_y2, h_s_wallace_rca24_fa332_y4);
  fa fa_h_s_wallace_rca24_fa333_y2(h_s_wallace_rca24_fa332_y4, h_s_wallace_rca24_fa130_y2, h_s_wallace_rca24_fa165_y2, h_s_wallace_rca24_fa333_y2, h_s_wallace_rca24_fa333_y4);
  fa fa_h_s_wallace_rca24_fa334_y2(h_s_wallace_rca24_fa333_y4, h_s_wallace_rca24_fa94_y2, h_s_wallace_rca24_fa131_y2, h_s_wallace_rca24_fa334_y2, h_s_wallace_rca24_fa334_y4);
  fa fa_h_s_wallace_rca24_fa335_y2(h_s_wallace_rca24_fa334_y4, h_s_wallace_rca24_fa56_y2, h_s_wallace_rca24_fa95_y2, h_s_wallace_rca24_fa335_y2, h_s_wallace_rca24_fa335_y4);
  fa fa_h_s_wallace_rca24_fa336_y2(h_s_wallace_rca24_fa335_y4, h_s_wallace_rca24_fa16_y2, h_s_wallace_rca24_fa57_y2, h_s_wallace_rca24_fa336_y2, h_s_wallace_rca24_fa336_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_20_y0(a_0, b_20, h_s_wallace_rca24_and_0_20_y0);
  fa fa_h_s_wallace_rca24_fa337_y2(h_s_wallace_rca24_fa336_y4, h_s_wallace_rca24_and_0_20_y0, h_s_wallace_rca24_fa17_y2, h_s_wallace_rca24_fa337_y2, h_s_wallace_rca24_fa337_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_20_y0(a_1, b_20, h_s_wallace_rca24_and_1_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_21_y0(a_0, b_21, h_s_wallace_rca24_and_0_21_y0);
  fa fa_h_s_wallace_rca24_fa338_y2(h_s_wallace_rca24_fa337_y4, h_s_wallace_rca24_and_1_20_y0, h_s_wallace_rca24_and_0_21_y0, h_s_wallace_rca24_fa338_y2, h_s_wallace_rca24_fa338_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_20_y0(a_2, b_20, h_s_wallace_rca24_and_2_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_21_y0(a_1, b_21, h_s_wallace_rca24_and_1_21_y0);
  fa fa_h_s_wallace_rca24_fa339_y2(h_s_wallace_rca24_fa338_y4, h_s_wallace_rca24_and_2_20_y0, h_s_wallace_rca24_and_1_21_y0, h_s_wallace_rca24_fa339_y2, h_s_wallace_rca24_fa339_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_20_y0(a_3, b_20, h_s_wallace_rca24_and_3_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_2_21_y0(a_2, b_21, h_s_wallace_rca24_and_2_21_y0);
  fa fa_h_s_wallace_rca24_fa340_y2(h_s_wallace_rca24_fa339_y4, h_s_wallace_rca24_and_3_20_y0, h_s_wallace_rca24_and_2_21_y0, h_s_wallace_rca24_fa340_y2, h_s_wallace_rca24_fa340_y4);
  and_gate and_gate_h_s_wallace_rca24_and_4_20_y0(a_4, b_20, h_s_wallace_rca24_and_4_20_y0);
  and_gate and_gate_h_s_wallace_rca24_and_3_21_y0(a_3, b_21, h_s_wallace_rca24_and_3_21_y0);
  fa fa_h_s_wallace_rca24_fa341_y2(h_s_wallace_rca24_fa340_y4, h_s_wallace_rca24_and_4_20_y0, h_s_wallace_rca24_and_3_21_y0, h_s_wallace_rca24_fa341_y2, h_s_wallace_rca24_fa341_y4);
  and_gate and_gate_h_s_wallace_rca24_and_3_22_y0(a_3, b_22, h_s_wallace_rca24_and_3_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_2_23_y0(a_2, b_23, h_s_wallace_rca24_nand_2_23_y0);
  fa fa_h_s_wallace_rca24_fa342_y2(h_s_wallace_rca24_fa341_y4, h_s_wallace_rca24_and_3_22_y0, h_s_wallace_rca24_nand_2_23_y0, h_s_wallace_rca24_fa342_y2, h_s_wallace_rca24_fa342_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_3_23_y0(a_3, b_23, h_s_wallace_rca24_nand_3_23_y0);
  fa fa_h_s_wallace_rca24_fa343_y2(h_s_wallace_rca24_fa342_y4, h_s_wallace_rca24_nand_3_23_y0, h_s_wallace_rca24_fa23_y2, h_s_wallace_rca24_fa343_y2, h_s_wallace_rca24_fa343_y4);
  fa fa_h_s_wallace_rca24_fa344_y2(h_s_wallace_rca24_fa343_y4, h_s_wallace_rca24_fa24_y2, h_s_wallace_rca24_fa65_y2, h_s_wallace_rca24_fa344_y2, h_s_wallace_rca24_fa344_y4);
  fa fa_h_s_wallace_rca24_fa345_y2(h_s_wallace_rca24_fa344_y4, h_s_wallace_rca24_fa66_y2, h_s_wallace_rca24_fa105_y2, h_s_wallace_rca24_fa345_y2, h_s_wallace_rca24_fa345_y4);
  fa fa_h_s_wallace_rca24_fa346_y2(h_s_wallace_rca24_fa345_y4, h_s_wallace_rca24_fa106_y2, h_s_wallace_rca24_fa143_y2, h_s_wallace_rca24_fa346_y2, h_s_wallace_rca24_fa346_y4);
  fa fa_h_s_wallace_rca24_fa347_y2(h_s_wallace_rca24_fa346_y4, h_s_wallace_rca24_fa144_y2, h_s_wallace_rca24_fa179_y2, h_s_wallace_rca24_fa347_y2, h_s_wallace_rca24_fa347_y4);
  fa fa_h_s_wallace_rca24_fa348_y2(h_s_wallace_rca24_fa347_y4, h_s_wallace_rca24_fa180_y2, h_s_wallace_rca24_fa213_y2, h_s_wallace_rca24_fa348_y2, h_s_wallace_rca24_fa348_y4);
  fa fa_h_s_wallace_rca24_fa349_y2(h_s_wallace_rca24_fa348_y4, h_s_wallace_rca24_fa214_y2, h_s_wallace_rca24_fa245_y2, h_s_wallace_rca24_fa349_y2, h_s_wallace_rca24_fa349_y4);
  fa fa_h_s_wallace_rca24_fa350_y2(h_s_wallace_rca24_fa349_y4, h_s_wallace_rca24_fa246_y2, h_s_wallace_rca24_fa275_y2, h_s_wallace_rca24_fa350_y2, h_s_wallace_rca24_fa350_y4);
  fa fa_h_s_wallace_rca24_fa351_y2(h_s_wallace_rca24_fa350_y4, h_s_wallace_rca24_fa276_y2, h_s_wallace_rca24_fa303_y2, h_s_wallace_rca24_fa351_y2, h_s_wallace_rca24_fa351_y4);
  ha ha_h_s_wallace_rca24_ha11_y0(h_s_wallace_rca24_fa282_y2, h_s_wallace_rca24_fa307_y2, h_s_wallace_rca24_ha11_y0, h_s_wallace_rca24_ha11_y1);
  fa fa_h_s_wallace_rca24_fa352_y2(h_s_wallace_rca24_ha11_y1, h_s_wallace_rca24_fa256_y2, h_s_wallace_rca24_fa283_y2, h_s_wallace_rca24_fa352_y2, h_s_wallace_rca24_fa352_y4);
  fa fa_h_s_wallace_rca24_fa353_y2(h_s_wallace_rca24_fa352_y4, h_s_wallace_rca24_fa228_y2, h_s_wallace_rca24_fa257_y2, h_s_wallace_rca24_fa353_y2, h_s_wallace_rca24_fa353_y4);
  fa fa_h_s_wallace_rca24_fa354_y2(h_s_wallace_rca24_fa353_y4, h_s_wallace_rca24_fa198_y2, h_s_wallace_rca24_fa229_y2, h_s_wallace_rca24_fa354_y2, h_s_wallace_rca24_fa354_y4);
  fa fa_h_s_wallace_rca24_fa355_y2(h_s_wallace_rca24_fa354_y4, h_s_wallace_rca24_fa166_y2, h_s_wallace_rca24_fa199_y2, h_s_wallace_rca24_fa355_y2, h_s_wallace_rca24_fa355_y4);
  fa fa_h_s_wallace_rca24_fa356_y2(h_s_wallace_rca24_fa355_y4, h_s_wallace_rca24_fa132_y2, h_s_wallace_rca24_fa167_y2, h_s_wallace_rca24_fa356_y2, h_s_wallace_rca24_fa356_y4);
  fa fa_h_s_wallace_rca24_fa357_y2(h_s_wallace_rca24_fa356_y4, h_s_wallace_rca24_fa96_y2, h_s_wallace_rca24_fa133_y2, h_s_wallace_rca24_fa357_y2, h_s_wallace_rca24_fa357_y4);
  fa fa_h_s_wallace_rca24_fa358_y2(h_s_wallace_rca24_fa357_y4, h_s_wallace_rca24_fa58_y2, h_s_wallace_rca24_fa97_y2, h_s_wallace_rca24_fa358_y2, h_s_wallace_rca24_fa358_y4);
  fa fa_h_s_wallace_rca24_fa359_y2(h_s_wallace_rca24_fa358_y4, h_s_wallace_rca24_fa18_y2, h_s_wallace_rca24_fa59_y2, h_s_wallace_rca24_fa359_y2, h_s_wallace_rca24_fa359_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_22_y0(a_0, b_22, h_s_wallace_rca24_and_0_22_y0);
  fa fa_h_s_wallace_rca24_fa360_y2(h_s_wallace_rca24_fa359_y4, h_s_wallace_rca24_and_0_22_y0, h_s_wallace_rca24_fa19_y2, h_s_wallace_rca24_fa360_y2, h_s_wallace_rca24_fa360_y4);
  and_gate and_gate_h_s_wallace_rca24_and_1_22_y0(a_1, b_22, h_s_wallace_rca24_and_1_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_0_23_y0(a_0, b_23, h_s_wallace_rca24_nand_0_23_y0);
  fa fa_h_s_wallace_rca24_fa361_y2(h_s_wallace_rca24_fa360_y4, h_s_wallace_rca24_and_1_22_y0, h_s_wallace_rca24_nand_0_23_y0, h_s_wallace_rca24_fa361_y2, h_s_wallace_rca24_fa361_y4);
  and_gate and_gate_h_s_wallace_rca24_and_2_22_y0(a_2, b_22, h_s_wallace_rca24_and_2_22_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_1_23_y0(a_1, b_23, h_s_wallace_rca24_nand_1_23_y0);
  fa fa_h_s_wallace_rca24_fa362_y2(h_s_wallace_rca24_fa361_y4, h_s_wallace_rca24_and_2_22_y0, h_s_wallace_rca24_nand_1_23_y0, h_s_wallace_rca24_fa362_y2, h_s_wallace_rca24_fa362_y4);
  fa fa_h_s_wallace_rca24_fa363_y2(h_s_wallace_rca24_fa362_y4, h_s_wallace_rca24_fa22_y2, h_s_wallace_rca24_fa63_y2, h_s_wallace_rca24_fa363_y2, h_s_wallace_rca24_fa363_y4);
  fa fa_h_s_wallace_rca24_fa364_y2(h_s_wallace_rca24_fa363_y4, h_s_wallace_rca24_fa64_y2, h_s_wallace_rca24_fa103_y2, h_s_wallace_rca24_fa364_y2, h_s_wallace_rca24_fa364_y4);
  fa fa_h_s_wallace_rca24_fa365_y2(h_s_wallace_rca24_fa364_y4, h_s_wallace_rca24_fa104_y2, h_s_wallace_rca24_fa141_y2, h_s_wallace_rca24_fa365_y2, h_s_wallace_rca24_fa365_y4);
  fa fa_h_s_wallace_rca24_fa366_y2(h_s_wallace_rca24_fa365_y4, h_s_wallace_rca24_fa142_y2, h_s_wallace_rca24_fa177_y2, h_s_wallace_rca24_fa366_y2, h_s_wallace_rca24_fa366_y4);
  fa fa_h_s_wallace_rca24_fa367_y2(h_s_wallace_rca24_fa366_y4, h_s_wallace_rca24_fa178_y2, h_s_wallace_rca24_fa211_y2, h_s_wallace_rca24_fa367_y2, h_s_wallace_rca24_fa367_y4);
  fa fa_h_s_wallace_rca24_fa368_y2(h_s_wallace_rca24_fa367_y4, h_s_wallace_rca24_fa212_y2, h_s_wallace_rca24_fa243_y2, h_s_wallace_rca24_fa368_y2, h_s_wallace_rca24_fa368_y4);
  fa fa_h_s_wallace_rca24_fa369_y2(h_s_wallace_rca24_fa368_y4, h_s_wallace_rca24_fa244_y2, h_s_wallace_rca24_fa273_y2, h_s_wallace_rca24_fa369_y2, h_s_wallace_rca24_fa369_y4);
  fa fa_h_s_wallace_rca24_fa370_y2(h_s_wallace_rca24_fa369_y4, h_s_wallace_rca24_fa274_y2, h_s_wallace_rca24_fa301_y2, h_s_wallace_rca24_fa370_y2, h_s_wallace_rca24_fa370_y4);
  fa fa_h_s_wallace_rca24_fa371_y2(h_s_wallace_rca24_fa370_y4, h_s_wallace_rca24_fa302_y2, h_s_wallace_rca24_fa327_y2, h_s_wallace_rca24_fa371_y2, h_s_wallace_rca24_fa371_y4);
  ha ha_h_s_wallace_rca24_ha12_y0(h_s_wallace_rca24_fa308_y2, h_s_wallace_rca24_fa331_y2, h_s_wallace_rca24_ha12_y0, h_s_wallace_rca24_ha12_y1);
  fa fa_h_s_wallace_rca24_fa372_y2(h_s_wallace_rca24_ha12_y1, h_s_wallace_rca24_fa284_y2, h_s_wallace_rca24_fa309_y2, h_s_wallace_rca24_fa372_y2, h_s_wallace_rca24_fa372_y4);
  fa fa_h_s_wallace_rca24_fa373_y2(h_s_wallace_rca24_fa372_y4, h_s_wallace_rca24_fa258_y2, h_s_wallace_rca24_fa285_y2, h_s_wallace_rca24_fa373_y2, h_s_wallace_rca24_fa373_y4);
  fa fa_h_s_wallace_rca24_fa374_y2(h_s_wallace_rca24_fa373_y4, h_s_wallace_rca24_fa230_y2, h_s_wallace_rca24_fa259_y2, h_s_wallace_rca24_fa374_y2, h_s_wallace_rca24_fa374_y4);
  fa fa_h_s_wallace_rca24_fa375_y2(h_s_wallace_rca24_fa374_y4, h_s_wallace_rca24_fa200_y2, h_s_wallace_rca24_fa231_y2, h_s_wallace_rca24_fa375_y2, h_s_wallace_rca24_fa375_y4);
  fa fa_h_s_wallace_rca24_fa376_y2(h_s_wallace_rca24_fa375_y4, h_s_wallace_rca24_fa168_y2, h_s_wallace_rca24_fa201_y2, h_s_wallace_rca24_fa376_y2, h_s_wallace_rca24_fa376_y4);
  fa fa_h_s_wallace_rca24_fa377_y2(h_s_wallace_rca24_fa376_y4, h_s_wallace_rca24_fa134_y2, h_s_wallace_rca24_fa169_y2, h_s_wallace_rca24_fa377_y2, h_s_wallace_rca24_fa377_y4);
  fa fa_h_s_wallace_rca24_fa378_y2(h_s_wallace_rca24_fa377_y4, h_s_wallace_rca24_fa98_y2, h_s_wallace_rca24_fa135_y2, h_s_wallace_rca24_fa378_y2, h_s_wallace_rca24_fa378_y4);
  fa fa_h_s_wallace_rca24_fa379_y2(h_s_wallace_rca24_fa378_y4, h_s_wallace_rca24_fa60_y2, h_s_wallace_rca24_fa99_y2, h_s_wallace_rca24_fa379_y2, h_s_wallace_rca24_fa379_y4);
  fa fa_h_s_wallace_rca24_fa380_y2(h_s_wallace_rca24_fa379_y4, h_s_wallace_rca24_fa20_y2, h_s_wallace_rca24_fa61_y2, h_s_wallace_rca24_fa380_y2, h_s_wallace_rca24_fa380_y4);
  fa fa_h_s_wallace_rca24_fa381_y2(h_s_wallace_rca24_fa380_y4, h_s_wallace_rca24_fa21_y2, h_s_wallace_rca24_fa62_y2, h_s_wallace_rca24_fa381_y2, h_s_wallace_rca24_fa381_y4);
  fa fa_h_s_wallace_rca24_fa382_y2(h_s_wallace_rca24_fa381_y4, h_s_wallace_rca24_fa102_y2, h_s_wallace_rca24_fa139_y2, h_s_wallace_rca24_fa382_y2, h_s_wallace_rca24_fa382_y4);
  fa fa_h_s_wallace_rca24_fa383_y2(h_s_wallace_rca24_fa382_y4, h_s_wallace_rca24_fa140_y2, h_s_wallace_rca24_fa175_y2, h_s_wallace_rca24_fa383_y2, h_s_wallace_rca24_fa383_y4);
  fa fa_h_s_wallace_rca24_fa384_y2(h_s_wallace_rca24_fa383_y4, h_s_wallace_rca24_fa176_y2, h_s_wallace_rca24_fa209_y2, h_s_wallace_rca24_fa384_y2, h_s_wallace_rca24_fa384_y4);
  fa fa_h_s_wallace_rca24_fa385_y2(h_s_wallace_rca24_fa384_y4, h_s_wallace_rca24_fa210_y2, h_s_wallace_rca24_fa241_y2, h_s_wallace_rca24_fa385_y2, h_s_wallace_rca24_fa385_y4);
  fa fa_h_s_wallace_rca24_fa386_y2(h_s_wallace_rca24_fa385_y4, h_s_wallace_rca24_fa242_y2, h_s_wallace_rca24_fa271_y2, h_s_wallace_rca24_fa386_y2, h_s_wallace_rca24_fa386_y4);
  fa fa_h_s_wallace_rca24_fa387_y2(h_s_wallace_rca24_fa386_y4, h_s_wallace_rca24_fa272_y2, h_s_wallace_rca24_fa299_y2, h_s_wallace_rca24_fa387_y2, h_s_wallace_rca24_fa387_y4);
  fa fa_h_s_wallace_rca24_fa388_y2(h_s_wallace_rca24_fa387_y4, h_s_wallace_rca24_fa300_y2, h_s_wallace_rca24_fa325_y2, h_s_wallace_rca24_fa388_y2, h_s_wallace_rca24_fa388_y4);
  fa fa_h_s_wallace_rca24_fa389_y2(h_s_wallace_rca24_fa388_y4, h_s_wallace_rca24_fa326_y2, h_s_wallace_rca24_fa349_y2, h_s_wallace_rca24_fa389_y2, h_s_wallace_rca24_fa389_y4);
  ha ha_h_s_wallace_rca24_ha13_y0(h_s_wallace_rca24_fa332_y2, h_s_wallace_rca24_fa353_y2, h_s_wallace_rca24_ha13_y0, h_s_wallace_rca24_ha13_y1);
  fa fa_h_s_wallace_rca24_fa390_y2(h_s_wallace_rca24_ha13_y1, h_s_wallace_rca24_fa310_y2, h_s_wallace_rca24_fa333_y2, h_s_wallace_rca24_fa390_y2, h_s_wallace_rca24_fa390_y4);
  fa fa_h_s_wallace_rca24_fa391_y2(h_s_wallace_rca24_fa390_y4, h_s_wallace_rca24_fa286_y2, h_s_wallace_rca24_fa311_y2, h_s_wallace_rca24_fa391_y2, h_s_wallace_rca24_fa391_y4);
  fa fa_h_s_wallace_rca24_fa392_y2(h_s_wallace_rca24_fa391_y4, h_s_wallace_rca24_fa260_y2, h_s_wallace_rca24_fa287_y2, h_s_wallace_rca24_fa392_y2, h_s_wallace_rca24_fa392_y4);
  fa fa_h_s_wallace_rca24_fa393_y2(h_s_wallace_rca24_fa392_y4, h_s_wallace_rca24_fa232_y2, h_s_wallace_rca24_fa261_y2, h_s_wallace_rca24_fa393_y2, h_s_wallace_rca24_fa393_y4);
  fa fa_h_s_wallace_rca24_fa394_y2(h_s_wallace_rca24_fa393_y4, h_s_wallace_rca24_fa202_y2, h_s_wallace_rca24_fa233_y2, h_s_wallace_rca24_fa394_y2, h_s_wallace_rca24_fa394_y4);
  fa fa_h_s_wallace_rca24_fa395_y2(h_s_wallace_rca24_fa394_y4, h_s_wallace_rca24_fa170_y2, h_s_wallace_rca24_fa203_y2, h_s_wallace_rca24_fa395_y2, h_s_wallace_rca24_fa395_y4);
  fa fa_h_s_wallace_rca24_fa396_y2(h_s_wallace_rca24_fa395_y4, h_s_wallace_rca24_fa136_y2, h_s_wallace_rca24_fa171_y2, h_s_wallace_rca24_fa396_y2, h_s_wallace_rca24_fa396_y4);
  fa fa_h_s_wallace_rca24_fa397_y2(h_s_wallace_rca24_fa396_y4, h_s_wallace_rca24_fa100_y2, h_s_wallace_rca24_fa137_y2, h_s_wallace_rca24_fa397_y2, h_s_wallace_rca24_fa397_y4);
  fa fa_h_s_wallace_rca24_fa398_y2(h_s_wallace_rca24_fa397_y4, h_s_wallace_rca24_fa101_y2, h_s_wallace_rca24_fa138_y2, h_s_wallace_rca24_fa398_y2, h_s_wallace_rca24_fa398_y4);
  fa fa_h_s_wallace_rca24_fa399_y2(h_s_wallace_rca24_fa398_y4, h_s_wallace_rca24_fa174_y2, h_s_wallace_rca24_fa207_y2, h_s_wallace_rca24_fa399_y2, h_s_wallace_rca24_fa399_y4);
  fa fa_h_s_wallace_rca24_fa400_y2(h_s_wallace_rca24_fa399_y4, h_s_wallace_rca24_fa208_y2, h_s_wallace_rca24_fa239_y2, h_s_wallace_rca24_fa400_y2, h_s_wallace_rca24_fa400_y4);
  fa fa_h_s_wallace_rca24_fa401_y2(h_s_wallace_rca24_fa400_y4, h_s_wallace_rca24_fa240_y2, h_s_wallace_rca24_fa269_y2, h_s_wallace_rca24_fa401_y2, h_s_wallace_rca24_fa401_y4);
  fa fa_h_s_wallace_rca24_fa402_y2(h_s_wallace_rca24_fa401_y4, h_s_wallace_rca24_fa270_y2, h_s_wallace_rca24_fa297_y2, h_s_wallace_rca24_fa402_y2, h_s_wallace_rca24_fa402_y4);
  fa fa_h_s_wallace_rca24_fa403_y2(h_s_wallace_rca24_fa402_y4, h_s_wallace_rca24_fa298_y2, h_s_wallace_rca24_fa323_y2, h_s_wallace_rca24_fa403_y2, h_s_wallace_rca24_fa403_y4);
  fa fa_h_s_wallace_rca24_fa404_y2(h_s_wallace_rca24_fa403_y4, h_s_wallace_rca24_fa324_y2, h_s_wallace_rca24_fa347_y2, h_s_wallace_rca24_fa404_y2, h_s_wallace_rca24_fa404_y4);
  fa fa_h_s_wallace_rca24_fa405_y2(h_s_wallace_rca24_fa404_y4, h_s_wallace_rca24_fa348_y2, h_s_wallace_rca24_fa369_y2, h_s_wallace_rca24_fa405_y2, h_s_wallace_rca24_fa405_y4);
  ha ha_h_s_wallace_rca24_ha14_y0(h_s_wallace_rca24_fa354_y2, h_s_wallace_rca24_fa373_y2, h_s_wallace_rca24_ha14_y0, h_s_wallace_rca24_ha14_y1);
  fa fa_h_s_wallace_rca24_fa406_y2(h_s_wallace_rca24_ha14_y1, h_s_wallace_rca24_fa334_y2, h_s_wallace_rca24_fa355_y2, h_s_wallace_rca24_fa406_y2, h_s_wallace_rca24_fa406_y4);
  fa fa_h_s_wallace_rca24_fa407_y2(h_s_wallace_rca24_fa406_y4, h_s_wallace_rca24_fa312_y2, h_s_wallace_rca24_fa335_y2, h_s_wallace_rca24_fa407_y2, h_s_wallace_rca24_fa407_y4);
  fa fa_h_s_wallace_rca24_fa408_y2(h_s_wallace_rca24_fa407_y4, h_s_wallace_rca24_fa288_y2, h_s_wallace_rca24_fa313_y2, h_s_wallace_rca24_fa408_y2, h_s_wallace_rca24_fa408_y4);
  fa fa_h_s_wallace_rca24_fa409_y2(h_s_wallace_rca24_fa408_y4, h_s_wallace_rca24_fa262_y2, h_s_wallace_rca24_fa289_y2, h_s_wallace_rca24_fa409_y2, h_s_wallace_rca24_fa409_y4);
  fa fa_h_s_wallace_rca24_fa410_y2(h_s_wallace_rca24_fa409_y4, h_s_wallace_rca24_fa234_y2, h_s_wallace_rca24_fa263_y2, h_s_wallace_rca24_fa410_y2, h_s_wallace_rca24_fa410_y4);
  fa fa_h_s_wallace_rca24_fa411_y2(h_s_wallace_rca24_fa410_y4, h_s_wallace_rca24_fa204_y2, h_s_wallace_rca24_fa235_y2, h_s_wallace_rca24_fa411_y2, h_s_wallace_rca24_fa411_y4);
  fa fa_h_s_wallace_rca24_fa412_y2(h_s_wallace_rca24_fa411_y4, h_s_wallace_rca24_fa172_y2, h_s_wallace_rca24_fa205_y2, h_s_wallace_rca24_fa412_y2, h_s_wallace_rca24_fa412_y4);
  fa fa_h_s_wallace_rca24_fa413_y2(h_s_wallace_rca24_fa412_y4, h_s_wallace_rca24_fa173_y2, h_s_wallace_rca24_fa206_y2, h_s_wallace_rca24_fa413_y2, h_s_wallace_rca24_fa413_y4);
  fa fa_h_s_wallace_rca24_fa414_y2(h_s_wallace_rca24_fa413_y4, h_s_wallace_rca24_fa238_y2, h_s_wallace_rca24_fa267_y2, h_s_wallace_rca24_fa414_y2, h_s_wallace_rca24_fa414_y4);
  fa fa_h_s_wallace_rca24_fa415_y2(h_s_wallace_rca24_fa414_y4, h_s_wallace_rca24_fa268_y2, h_s_wallace_rca24_fa295_y2, h_s_wallace_rca24_fa415_y2, h_s_wallace_rca24_fa415_y4);
  fa fa_h_s_wallace_rca24_fa416_y2(h_s_wallace_rca24_fa415_y4, h_s_wallace_rca24_fa296_y2, h_s_wallace_rca24_fa321_y2, h_s_wallace_rca24_fa416_y2, h_s_wallace_rca24_fa416_y4);
  fa fa_h_s_wallace_rca24_fa417_y2(h_s_wallace_rca24_fa416_y4, h_s_wallace_rca24_fa322_y2, h_s_wallace_rca24_fa345_y2, h_s_wallace_rca24_fa417_y2, h_s_wallace_rca24_fa417_y4);
  fa fa_h_s_wallace_rca24_fa418_y2(h_s_wallace_rca24_fa417_y4, h_s_wallace_rca24_fa346_y2, h_s_wallace_rca24_fa367_y2, h_s_wallace_rca24_fa418_y2, h_s_wallace_rca24_fa418_y4);
  fa fa_h_s_wallace_rca24_fa419_y2(h_s_wallace_rca24_fa418_y4, h_s_wallace_rca24_fa368_y2, h_s_wallace_rca24_fa387_y2, h_s_wallace_rca24_fa419_y2, h_s_wallace_rca24_fa419_y4);
  ha ha_h_s_wallace_rca24_ha15_y0(h_s_wallace_rca24_fa374_y2, h_s_wallace_rca24_fa391_y2, h_s_wallace_rca24_ha15_y0, h_s_wallace_rca24_ha15_y1);
  fa fa_h_s_wallace_rca24_fa420_y2(h_s_wallace_rca24_ha15_y1, h_s_wallace_rca24_fa356_y2, h_s_wallace_rca24_fa375_y2, h_s_wallace_rca24_fa420_y2, h_s_wallace_rca24_fa420_y4);
  fa fa_h_s_wallace_rca24_fa421_y2(h_s_wallace_rca24_fa420_y4, h_s_wallace_rca24_fa336_y2, h_s_wallace_rca24_fa357_y2, h_s_wallace_rca24_fa421_y2, h_s_wallace_rca24_fa421_y4);
  fa fa_h_s_wallace_rca24_fa422_y2(h_s_wallace_rca24_fa421_y4, h_s_wallace_rca24_fa314_y2, h_s_wallace_rca24_fa337_y2, h_s_wallace_rca24_fa422_y2, h_s_wallace_rca24_fa422_y4);
  fa fa_h_s_wallace_rca24_fa423_y2(h_s_wallace_rca24_fa422_y4, h_s_wallace_rca24_fa290_y2, h_s_wallace_rca24_fa315_y2, h_s_wallace_rca24_fa423_y2, h_s_wallace_rca24_fa423_y4);
  fa fa_h_s_wallace_rca24_fa424_y2(h_s_wallace_rca24_fa423_y4, h_s_wallace_rca24_fa264_y2, h_s_wallace_rca24_fa291_y2, h_s_wallace_rca24_fa424_y2, h_s_wallace_rca24_fa424_y4);
  fa fa_h_s_wallace_rca24_fa425_y2(h_s_wallace_rca24_fa424_y4, h_s_wallace_rca24_fa236_y2, h_s_wallace_rca24_fa265_y2, h_s_wallace_rca24_fa425_y2, h_s_wallace_rca24_fa425_y4);
  fa fa_h_s_wallace_rca24_fa426_y2(h_s_wallace_rca24_fa425_y4, h_s_wallace_rca24_fa237_y2, h_s_wallace_rca24_fa266_y2, h_s_wallace_rca24_fa426_y2, h_s_wallace_rca24_fa426_y4);
  fa fa_h_s_wallace_rca24_fa427_y2(h_s_wallace_rca24_fa426_y4, h_s_wallace_rca24_fa294_y2, h_s_wallace_rca24_fa319_y2, h_s_wallace_rca24_fa427_y2, h_s_wallace_rca24_fa427_y4);
  fa fa_h_s_wallace_rca24_fa428_y2(h_s_wallace_rca24_fa427_y4, h_s_wallace_rca24_fa320_y2, h_s_wallace_rca24_fa343_y2, h_s_wallace_rca24_fa428_y2, h_s_wallace_rca24_fa428_y4);
  fa fa_h_s_wallace_rca24_fa429_y2(h_s_wallace_rca24_fa428_y4, h_s_wallace_rca24_fa344_y2, h_s_wallace_rca24_fa365_y2, h_s_wallace_rca24_fa429_y2, h_s_wallace_rca24_fa429_y4);
  fa fa_h_s_wallace_rca24_fa430_y2(h_s_wallace_rca24_fa429_y4, h_s_wallace_rca24_fa366_y2, h_s_wallace_rca24_fa385_y2, h_s_wallace_rca24_fa430_y2, h_s_wallace_rca24_fa430_y4);
  fa fa_h_s_wallace_rca24_fa431_y2(h_s_wallace_rca24_fa430_y4, h_s_wallace_rca24_fa386_y2, h_s_wallace_rca24_fa403_y2, h_s_wallace_rca24_fa431_y2, h_s_wallace_rca24_fa431_y4);
  ha ha_h_s_wallace_rca24_ha16_y0(h_s_wallace_rca24_fa392_y2, h_s_wallace_rca24_fa407_y2, h_s_wallace_rca24_ha16_y0, h_s_wallace_rca24_ha16_y1);
  fa fa_h_s_wallace_rca24_fa432_y2(h_s_wallace_rca24_ha16_y1, h_s_wallace_rca24_fa376_y2, h_s_wallace_rca24_fa393_y2, h_s_wallace_rca24_fa432_y2, h_s_wallace_rca24_fa432_y4);
  fa fa_h_s_wallace_rca24_fa433_y2(h_s_wallace_rca24_fa432_y4, h_s_wallace_rca24_fa358_y2, h_s_wallace_rca24_fa377_y2, h_s_wallace_rca24_fa433_y2, h_s_wallace_rca24_fa433_y4);
  fa fa_h_s_wallace_rca24_fa434_y2(h_s_wallace_rca24_fa433_y4, h_s_wallace_rca24_fa338_y2, h_s_wallace_rca24_fa359_y2, h_s_wallace_rca24_fa434_y2, h_s_wallace_rca24_fa434_y4);
  fa fa_h_s_wallace_rca24_fa435_y2(h_s_wallace_rca24_fa434_y4, h_s_wallace_rca24_fa316_y2, h_s_wallace_rca24_fa339_y2, h_s_wallace_rca24_fa435_y2, h_s_wallace_rca24_fa435_y4);
  fa fa_h_s_wallace_rca24_fa436_y2(h_s_wallace_rca24_fa435_y4, h_s_wallace_rca24_fa292_y2, h_s_wallace_rca24_fa317_y2, h_s_wallace_rca24_fa436_y2, h_s_wallace_rca24_fa436_y4);
  fa fa_h_s_wallace_rca24_fa437_y2(h_s_wallace_rca24_fa436_y4, h_s_wallace_rca24_fa293_y2, h_s_wallace_rca24_fa318_y2, h_s_wallace_rca24_fa437_y2, h_s_wallace_rca24_fa437_y4);
  fa fa_h_s_wallace_rca24_fa438_y2(h_s_wallace_rca24_fa437_y4, h_s_wallace_rca24_fa342_y2, h_s_wallace_rca24_fa363_y2, h_s_wallace_rca24_fa438_y2, h_s_wallace_rca24_fa438_y4);
  fa fa_h_s_wallace_rca24_fa439_y2(h_s_wallace_rca24_fa438_y4, h_s_wallace_rca24_fa364_y2, h_s_wallace_rca24_fa383_y2, h_s_wallace_rca24_fa439_y2, h_s_wallace_rca24_fa439_y4);
  fa fa_h_s_wallace_rca24_fa440_y2(h_s_wallace_rca24_fa439_y4, h_s_wallace_rca24_fa384_y2, h_s_wallace_rca24_fa401_y2, h_s_wallace_rca24_fa440_y2, h_s_wallace_rca24_fa440_y4);
  fa fa_h_s_wallace_rca24_fa441_y2(h_s_wallace_rca24_fa440_y4, h_s_wallace_rca24_fa402_y2, h_s_wallace_rca24_fa417_y2, h_s_wallace_rca24_fa441_y2, h_s_wallace_rca24_fa441_y4);
  ha ha_h_s_wallace_rca24_ha17_y0(h_s_wallace_rca24_fa408_y2, h_s_wallace_rca24_fa421_y2, h_s_wallace_rca24_ha17_y0, h_s_wallace_rca24_ha17_y1);
  fa fa_h_s_wallace_rca24_fa442_y2(h_s_wallace_rca24_ha17_y1, h_s_wallace_rca24_fa394_y2, h_s_wallace_rca24_fa409_y2, h_s_wallace_rca24_fa442_y2, h_s_wallace_rca24_fa442_y4);
  fa fa_h_s_wallace_rca24_fa443_y2(h_s_wallace_rca24_fa442_y4, h_s_wallace_rca24_fa378_y2, h_s_wallace_rca24_fa395_y2, h_s_wallace_rca24_fa443_y2, h_s_wallace_rca24_fa443_y4);
  fa fa_h_s_wallace_rca24_fa444_y2(h_s_wallace_rca24_fa443_y4, h_s_wallace_rca24_fa360_y2, h_s_wallace_rca24_fa379_y2, h_s_wallace_rca24_fa444_y2, h_s_wallace_rca24_fa444_y4);
  fa fa_h_s_wallace_rca24_fa445_y2(h_s_wallace_rca24_fa444_y4, h_s_wallace_rca24_fa340_y2, h_s_wallace_rca24_fa361_y2, h_s_wallace_rca24_fa445_y2, h_s_wallace_rca24_fa445_y4);
  fa fa_h_s_wallace_rca24_fa446_y2(h_s_wallace_rca24_fa445_y4, h_s_wallace_rca24_fa341_y2, h_s_wallace_rca24_fa362_y2, h_s_wallace_rca24_fa446_y2, h_s_wallace_rca24_fa446_y4);
  fa fa_h_s_wallace_rca24_fa447_y2(h_s_wallace_rca24_fa446_y4, h_s_wallace_rca24_fa382_y2, h_s_wallace_rca24_fa399_y2, h_s_wallace_rca24_fa447_y2, h_s_wallace_rca24_fa447_y4);
  fa fa_h_s_wallace_rca24_fa448_y2(h_s_wallace_rca24_fa447_y4, h_s_wallace_rca24_fa400_y2, h_s_wallace_rca24_fa415_y2, h_s_wallace_rca24_fa448_y2, h_s_wallace_rca24_fa448_y4);
  fa fa_h_s_wallace_rca24_fa449_y2(h_s_wallace_rca24_fa448_y4, h_s_wallace_rca24_fa416_y2, h_s_wallace_rca24_fa429_y2, h_s_wallace_rca24_fa449_y2, h_s_wallace_rca24_fa449_y4);
  ha ha_h_s_wallace_rca24_ha18_y0(h_s_wallace_rca24_fa422_y2, h_s_wallace_rca24_fa433_y2, h_s_wallace_rca24_ha18_y0, h_s_wallace_rca24_ha18_y1);
  fa fa_h_s_wallace_rca24_fa450_y2(h_s_wallace_rca24_ha18_y1, h_s_wallace_rca24_fa410_y2, h_s_wallace_rca24_fa423_y2, h_s_wallace_rca24_fa450_y2, h_s_wallace_rca24_fa450_y4);
  fa fa_h_s_wallace_rca24_fa451_y2(h_s_wallace_rca24_fa450_y4, h_s_wallace_rca24_fa396_y2, h_s_wallace_rca24_fa411_y2, h_s_wallace_rca24_fa451_y2, h_s_wallace_rca24_fa451_y4);
  fa fa_h_s_wallace_rca24_fa452_y2(h_s_wallace_rca24_fa451_y4, h_s_wallace_rca24_fa380_y2, h_s_wallace_rca24_fa397_y2, h_s_wallace_rca24_fa452_y2, h_s_wallace_rca24_fa452_y4);
  fa fa_h_s_wallace_rca24_fa453_y2(h_s_wallace_rca24_fa452_y4, h_s_wallace_rca24_fa381_y2, h_s_wallace_rca24_fa398_y2, h_s_wallace_rca24_fa453_y2, h_s_wallace_rca24_fa453_y4);
  fa fa_h_s_wallace_rca24_fa454_y2(h_s_wallace_rca24_fa453_y4, h_s_wallace_rca24_fa414_y2, h_s_wallace_rca24_fa427_y2, h_s_wallace_rca24_fa454_y2, h_s_wallace_rca24_fa454_y4);
  fa fa_h_s_wallace_rca24_fa455_y2(h_s_wallace_rca24_fa454_y4, h_s_wallace_rca24_fa428_y2, h_s_wallace_rca24_fa439_y2, h_s_wallace_rca24_fa455_y2, h_s_wallace_rca24_fa455_y4);
  ha ha_h_s_wallace_rca24_ha19_y0(h_s_wallace_rca24_fa434_y2, h_s_wallace_rca24_fa443_y2, h_s_wallace_rca24_ha19_y0, h_s_wallace_rca24_ha19_y1);
  fa fa_h_s_wallace_rca24_fa456_y2(h_s_wallace_rca24_ha19_y1, h_s_wallace_rca24_fa424_y2, h_s_wallace_rca24_fa435_y2, h_s_wallace_rca24_fa456_y2, h_s_wallace_rca24_fa456_y4);
  fa fa_h_s_wallace_rca24_fa457_y2(h_s_wallace_rca24_fa456_y4, h_s_wallace_rca24_fa412_y2, h_s_wallace_rca24_fa425_y2, h_s_wallace_rca24_fa457_y2, h_s_wallace_rca24_fa457_y4);
  fa fa_h_s_wallace_rca24_fa458_y2(h_s_wallace_rca24_fa457_y4, h_s_wallace_rca24_fa413_y2, h_s_wallace_rca24_fa426_y2, h_s_wallace_rca24_fa458_y2, h_s_wallace_rca24_fa458_y4);
  fa fa_h_s_wallace_rca24_fa459_y2(h_s_wallace_rca24_fa458_y4, h_s_wallace_rca24_fa438_y2, h_s_wallace_rca24_fa447_y2, h_s_wallace_rca24_fa459_y2, h_s_wallace_rca24_fa459_y4);
  ha ha_h_s_wallace_rca24_ha20_y0(h_s_wallace_rca24_fa444_y2, h_s_wallace_rca24_fa451_y2, h_s_wallace_rca24_ha20_y0, h_s_wallace_rca24_ha20_y1);
  fa fa_h_s_wallace_rca24_fa460_y2(h_s_wallace_rca24_ha20_y1, h_s_wallace_rca24_fa436_y2, h_s_wallace_rca24_fa445_y2, h_s_wallace_rca24_fa460_y2, h_s_wallace_rca24_fa460_y4);
  fa fa_h_s_wallace_rca24_fa461_y2(h_s_wallace_rca24_fa460_y4, h_s_wallace_rca24_fa437_y2, h_s_wallace_rca24_fa446_y2, h_s_wallace_rca24_fa461_y2, h_s_wallace_rca24_fa461_y4);
  ha ha_h_s_wallace_rca24_ha21_y0(h_s_wallace_rca24_fa452_y2, h_s_wallace_rca24_fa457_y2, h_s_wallace_rca24_ha21_y0, h_s_wallace_rca24_ha21_y1);
  fa fa_h_s_wallace_rca24_fa462_y2(h_s_wallace_rca24_ha21_y1, h_s_wallace_rca24_fa453_y2, h_s_wallace_rca24_fa458_y2, h_s_wallace_rca24_fa462_y2, h_s_wallace_rca24_fa462_y4);
  fa fa_h_s_wallace_rca24_fa463_y2(h_s_wallace_rca24_fa462_y4, h_s_wallace_rca24_fa461_y4, h_s_wallace_rca24_fa454_y2, h_s_wallace_rca24_fa463_y2, h_s_wallace_rca24_fa463_y4);
  fa fa_h_s_wallace_rca24_fa464_y2(h_s_wallace_rca24_fa463_y4, h_s_wallace_rca24_fa459_y4, h_s_wallace_rca24_fa448_y2, h_s_wallace_rca24_fa464_y2, h_s_wallace_rca24_fa464_y4);
  fa fa_h_s_wallace_rca24_fa465_y2(h_s_wallace_rca24_fa464_y4, h_s_wallace_rca24_fa455_y4, h_s_wallace_rca24_fa440_y2, h_s_wallace_rca24_fa465_y2, h_s_wallace_rca24_fa465_y4);
  fa fa_h_s_wallace_rca24_fa466_y2(h_s_wallace_rca24_fa465_y4, h_s_wallace_rca24_fa449_y4, h_s_wallace_rca24_fa430_y2, h_s_wallace_rca24_fa466_y2, h_s_wallace_rca24_fa466_y4);
  fa fa_h_s_wallace_rca24_fa467_y2(h_s_wallace_rca24_fa466_y4, h_s_wallace_rca24_fa441_y4, h_s_wallace_rca24_fa418_y2, h_s_wallace_rca24_fa467_y2, h_s_wallace_rca24_fa467_y4);
  fa fa_h_s_wallace_rca24_fa468_y2(h_s_wallace_rca24_fa467_y4, h_s_wallace_rca24_fa431_y4, h_s_wallace_rca24_fa404_y2, h_s_wallace_rca24_fa468_y2, h_s_wallace_rca24_fa468_y4);
  fa fa_h_s_wallace_rca24_fa469_y2(h_s_wallace_rca24_fa468_y4, h_s_wallace_rca24_fa419_y4, h_s_wallace_rca24_fa388_y2, h_s_wallace_rca24_fa469_y2, h_s_wallace_rca24_fa469_y4);
  fa fa_h_s_wallace_rca24_fa470_y2(h_s_wallace_rca24_fa469_y4, h_s_wallace_rca24_fa405_y4, h_s_wallace_rca24_fa370_y2, h_s_wallace_rca24_fa470_y2, h_s_wallace_rca24_fa470_y4);
  fa fa_h_s_wallace_rca24_fa471_y2(h_s_wallace_rca24_fa470_y4, h_s_wallace_rca24_fa389_y4, h_s_wallace_rca24_fa350_y2, h_s_wallace_rca24_fa471_y2, h_s_wallace_rca24_fa471_y4);
  fa fa_h_s_wallace_rca24_fa472_y2(h_s_wallace_rca24_fa471_y4, h_s_wallace_rca24_fa371_y4, h_s_wallace_rca24_fa328_y2, h_s_wallace_rca24_fa472_y2, h_s_wallace_rca24_fa472_y4);
  fa fa_h_s_wallace_rca24_fa473_y2(h_s_wallace_rca24_fa472_y4, h_s_wallace_rca24_fa351_y4, h_s_wallace_rca24_fa304_y2, h_s_wallace_rca24_fa473_y2, h_s_wallace_rca24_fa473_y4);
  fa fa_h_s_wallace_rca24_fa474_y2(h_s_wallace_rca24_fa473_y4, h_s_wallace_rca24_fa329_y4, h_s_wallace_rca24_fa278_y2, h_s_wallace_rca24_fa474_y2, h_s_wallace_rca24_fa474_y4);
  fa fa_h_s_wallace_rca24_fa475_y2(h_s_wallace_rca24_fa474_y4, h_s_wallace_rca24_fa305_y4, h_s_wallace_rca24_fa250_y2, h_s_wallace_rca24_fa475_y2, h_s_wallace_rca24_fa475_y4);
  fa fa_h_s_wallace_rca24_fa476_y2(h_s_wallace_rca24_fa475_y4, h_s_wallace_rca24_fa279_y4, h_s_wallace_rca24_fa220_y2, h_s_wallace_rca24_fa476_y2, h_s_wallace_rca24_fa476_y4);
  fa fa_h_s_wallace_rca24_fa477_y2(h_s_wallace_rca24_fa476_y4, h_s_wallace_rca24_fa251_y4, h_s_wallace_rca24_fa188_y2, h_s_wallace_rca24_fa477_y2, h_s_wallace_rca24_fa477_y4);
  fa fa_h_s_wallace_rca24_fa478_y2(h_s_wallace_rca24_fa477_y4, h_s_wallace_rca24_fa221_y4, h_s_wallace_rca24_fa154_y2, h_s_wallace_rca24_fa478_y2, h_s_wallace_rca24_fa478_y4);
  fa fa_h_s_wallace_rca24_fa479_y2(h_s_wallace_rca24_fa478_y4, h_s_wallace_rca24_fa189_y4, h_s_wallace_rca24_fa118_y2, h_s_wallace_rca24_fa479_y2, h_s_wallace_rca24_fa479_y4);
  fa fa_h_s_wallace_rca24_fa480_y2(h_s_wallace_rca24_fa479_y4, h_s_wallace_rca24_fa155_y4, h_s_wallace_rca24_fa80_y2, h_s_wallace_rca24_fa480_y2, h_s_wallace_rca24_fa480_y4);
  fa fa_h_s_wallace_rca24_fa481_y2(h_s_wallace_rca24_fa480_y4, h_s_wallace_rca24_fa119_y4, h_s_wallace_rca24_fa40_y2, h_s_wallace_rca24_fa481_y2, h_s_wallace_rca24_fa481_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_21_23_y0(a_21, b_23, h_s_wallace_rca24_nand_21_23_y0);
  fa fa_h_s_wallace_rca24_fa482_y2(h_s_wallace_rca24_fa481_y4, h_s_wallace_rca24_fa81_y4, h_s_wallace_rca24_nand_21_23_y0, h_s_wallace_rca24_fa482_y2, h_s_wallace_rca24_fa482_y4);
  nand_gate nand_gate_h_s_wallace_rca24_nand_23_22_y0(a_23, b_22, h_s_wallace_rca24_nand_23_22_y0);
  fa fa_h_s_wallace_rca24_fa483_y2(h_s_wallace_rca24_fa482_y4, h_s_wallace_rca24_fa41_y4, h_s_wallace_rca24_nand_23_22_y0, h_s_wallace_rca24_fa483_y2, h_s_wallace_rca24_fa483_y4);
  and_gate and_gate_h_s_wallace_rca24_and_0_0_y0(a_0, b_0, h_s_wallace_rca24_and_0_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_1_0_y0(a_1, b_0, h_s_wallace_rca24_and_1_0_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_2_y0(a_0, b_2, h_s_wallace_rca24_and_0_2_y0);
  nand_gate nand_gate_h_s_wallace_rca24_nand_22_23_y0(a_22, b_23, h_s_wallace_rca24_nand_22_23_y0);
  and_gate and_gate_h_s_wallace_rca24_and_0_1_y0(a_0, b_1, h_s_wallace_rca24_and_0_1_y0);
  and_gate and_gate_h_s_wallace_rca24_and_23_23_y0(a_23, b_23, h_s_wallace_rca24_and_23_23_y0);
  assign h_s_wallace_rca24_u_rca_u_rca_a[0] = h_s_wallace_rca24_and_1_0_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_a[1] = h_s_wallace_rca24_and_0_2_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_a[2] = h_s_wallace_rca24_fa0_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[3] = h_s_wallace_rca24_fa42_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[4] = h_s_wallace_rca24_fa82_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[5] = h_s_wallace_rca24_fa120_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[6] = h_s_wallace_rca24_fa156_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[7] = h_s_wallace_rca24_fa190_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[8] = h_s_wallace_rca24_fa222_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[9] = h_s_wallace_rca24_fa252_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[10] = h_s_wallace_rca24_fa280_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[11] = h_s_wallace_rca24_fa306_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[12] = h_s_wallace_rca24_fa330_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[13] = h_s_wallace_rca24_fa352_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[14] = h_s_wallace_rca24_fa372_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[15] = h_s_wallace_rca24_fa390_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[16] = h_s_wallace_rca24_fa406_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[17] = h_s_wallace_rca24_fa420_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[18] = h_s_wallace_rca24_fa432_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[19] = h_s_wallace_rca24_fa442_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[20] = h_s_wallace_rca24_fa450_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[21] = h_s_wallace_rca24_fa456_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[22] = h_s_wallace_rca24_fa460_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[23] = h_s_wallace_rca24_fa461_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[24] = h_s_wallace_rca24_fa459_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[25] = h_s_wallace_rca24_fa455_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[26] = h_s_wallace_rca24_fa449_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[27] = h_s_wallace_rca24_fa441_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[28] = h_s_wallace_rca24_fa431_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[29] = h_s_wallace_rca24_fa419_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[30] = h_s_wallace_rca24_fa405_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[31] = h_s_wallace_rca24_fa389_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[32] = h_s_wallace_rca24_fa371_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[33] = h_s_wallace_rca24_fa351_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[34] = h_s_wallace_rca24_fa329_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[35] = h_s_wallace_rca24_fa305_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[36] = h_s_wallace_rca24_fa279_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[37] = h_s_wallace_rca24_fa251_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[38] = h_s_wallace_rca24_fa221_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[39] = h_s_wallace_rca24_fa189_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[40] = h_s_wallace_rca24_fa155_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[41] = h_s_wallace_rca24_fa119_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[42] = h_s_wallace_rca24_fa81_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[43] = h_s_wallace_rca24_fa41_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_a[44] = h_s_wallace_rca24_nand_22_23_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_a[45] = h_s_wallace_rca24_fa483_y4;
  assign h_s_wallace_rca24_u_rca_u_rca_b[0] = h_s_wallace_rca24_and_0_1_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[1] = h_s_wallace_rca24_ha0_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[2] = h_s_wallace_rca24_ha1_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[3] = h_s_wallace_rca24_ha2_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[4] = h_s_wallace_rca24_ha3_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[5] = h_s_wallace_rca24_ha4_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[6] = h_s_wallace_rca24_ha5_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[7] = h_s_wallace_rca24_ha6_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[8] = h_s_wallace_rca24_ha7_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[9] = h_s_wallace_rca24_ha8_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[10] = h_s_wallace_rca24_ha9_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[11] = h_s_wallace_rca24_ha10_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[12] = h_s_wallace_rca24_ha11_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[13] = h_s_wallace_rca24_ha12_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[14] = h_s_wallace_rca24_ha13_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[15] = h_s_wallace_rca24_ha14_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[16] = h_s_wallace_rca24_ha15_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[17] = h_s_wallace_rca24_ha16_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[18] = h_s_wallace_rca24_ha17_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[19] = h_s_wallace_rca24_ha18_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[20] = h_s_wallace_rca24_ha19_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[21] = h_s_wallace_rca24_ha20_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[22] = h_s_wallace_rca24_ha21_y0;
  assign h_s_wallace_rca24_u_rca_u_rca_b[23] = h_s_wallace_rca24_fa462_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[24] = h_s_wallace_rca24_fa463_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[25] = h_s_wallace_rca24_fa464_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[26] = h_s_wallace_rca24_fa465_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[27] = h_s_wallace_rca24_fa466_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[28] = h_s_wallace_rca24_fa467_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[29] = h_s_wallace_rca24_fa468_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[30] = h_s_wallace_rca24_fa469_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[31] = h_s_wallace_rca24_fa470_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[32] = h_s_wallace_rca24_fa471_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[33] = h_s_wallace_rca24_fa472_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[34] = h_s_wallace_rca24_fa473_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[35] = h_s_wallace_rca24_fa474_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[36] = h_s_wallace_rca24_fa475_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[37] = h_s_wallace_rca24_fa476_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[38] = h_s_wallace_rca24_fa477_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[39] = h_s_wallace_rca24_fa478_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[40] = h_s_wallace_rca24_fa479_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[41] = h_s_wallace_rca24_fa480_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[42] = h_s_wallace_rca24_fa481_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[43] = h_s_wallace_rca24_fa482_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[44] = h_s_wallace_rca24_fa483_y2;
  assign h_s_wallace_rca24_u_rca_u_rca_b[45] = h_s_wallace_rca24_and_23_23_y0;
  u_rca u_rca_out(h_s_wallace_rca24_u_rca_u_rca_a, h_s_wallace_rca24_u_rca_u_rca_b, h_s_wallace_rca24_u_rca_out);
  assign h_s_wallace_rca24_u_rca_ha_y0 = h_s_wallace_rca24_u_rca_out[0];
  assign h_s_wallace_rca24_u_rca_fa1_y2 = h_s_wallace_rca24_u_rca_out[1];
  assign h_s_wallace_rca24_u_rca_fa2_y2 = h_s_wallace_rca24_u_rca_out[2];
  assign h_s_wallace_rca24_u_rca_fa3_y2 = h_s_wallace_rca24_u_rca_out[3];
  assign h_s_wallace_rca24_u_rca_fa4_y2 = h_s_wallace_rca24_u_rca_out[4];
  assign h_s_wallace_rca24_u_rca_fa5_y2 = h_s_wallace_rca24_u_rca_out[5];
  assign h_s_wallace_rca24_u_rca_fa6_y2 = h_s_wallace_rca24_u_rca_out[6];
  assign h_s_wallace_rca24_u_rca_fa7_y2 = h_s_wallace_rca24_u_rca_out[7];
  assign h_s_wallace_rca24_u_rca_fa8_y2 = h_s_wallace_rca24_u_rca_out[8];
  assign h_s_wallace_rca24_u_rca_fa9_y2 = h_s_wallace_rca24_u_rca_out[9];
  assign h_s_wallace_rca24_u_rca_fa10_y2 = h_s_wallace_rca24_u_rca_out[10];
  assign h_s_wallace_rca24_u_rca_fa11_y2 = h_s_wallace_rca24_u_rca_out[11];
  assign h_s_wallace_rca24_u_rca_fa12_y2 = h_s_wallace_rca24_u_rca_out[12];
  assign h_s_wallace_rca24_u_rca_fa13_y2 = h_s_wallace_rca24_u_rca_out[13];
  assign h_s_wallace_rca24_u_rca_fa14_y2 = h_s_wallace_rca24_u_rca_out[14];
  assign h_s_wallace_rca24_u_rca_fa15_y2 = h_s_wallace_rca24_u_rca_out[15];
  assign h_s_wallace_rca24_u_rca_fa16_y2 = h_s_wallace_rca24_u_rca_out[16];
  assign h_s_wallace_rca24_u_rca_fa17_y2 = h_s_wallace_rca24_u_rca_out[17];
  assign h_s_wallace_rca24_u_rca_fa18_y2 = h_s_wallace_rca24_u_rca_out[18];
  assign h_s_wallace_rca24_u_rca_fa19_y2 = h_s_wallace_rca24_u_rca_out[19];
  assign h_s_wallace_rca24_u_rca_fa20_y2 = h_s_wallace_rca24_u_rca_out[20];
  assign h_s_wallace_rca24_u_rca_fa21_y2 = h_s_wallace_rca24_u_rca_out[21];
  assign h_s_wallace_rca24_u_rca_fa22_y2 = h_s_wallace_rca24_u_rca_out[22];
  assign h_s_wallace_rca24_u_rca_fa23_y2 = h_s_wallace_rca24_u_rca_out[23];
  assign h_s_wallace_rca24_u_rca_fa24_y2 = h_s_wallace_rca24_u_rca_out[24];
  assign h_s_wallace_rca24_u_rca_fa25_y2 = h_s_wallace_rca24_u_rca_out[25];
  assign h_s_wallace_rca24_u_rca_fa26_y2 = h_s_wallace_rca24_u_rca_out[26];
  assign h_s_wallace_rca24_u_rca_fa27_y2 = h_s_wallace_rca24_u_rca_out[27];
  assign h_s_wallace_rca24_u_rca_fa28_y2 = h_s_wallace_rca24_u_rca_out[28];
  assign h_s_wallace_rca24_u_rca_fa29_y2 = h_s_wallace_rca24_u_rca_out[29];
  assign h_s_wallace_rca24_u_rca_fa30_y2 = h_s_wallace_rca24_u_rca_out[30];
  assign h_s_wallace_rca24_u_rca_fa31_y2 = h_s_wallace_rca24_u_rca_out[31];
  assign h_s_wallace_rca24_u_rca_fa32_y2 = h_s_wallace_rca24_u_rca_out[32];
  assign h_s_wallace_rca24_u_rca_fa33_y2 = h_s_wallace_rca24_u_rca_out[33];
  assign h_s_wallace_rca24_u_rca_fa34_y2 = h_s_wallace_rca24_u_rca_out[34];
  assign h_s_wallace_rca24_u_rca_fa35_y2 = h_s_wallace_rca24_u_rca_out[35];
  assign h_s_wallace_rca24_u_rca_fa36_y2 = h_s_wallace_rca24_u_rca_out[36];
  assign h_s_wallace_rca24_u_rca_fa37_y2 = h_s_wallace_rca24_u_rca_out[37];
  assign h_s_wallace_rca24_u_rca_fa38_y2 = h_s_wallace_rca24_u_rca_out[38];
  assign h_s_wallace_rca24_u_rca_fa39_y2 = h_s_wallace_rca24_u_rca_out[39];
  assign h_s_wallace_rca24_u_rca_fa40_y2 = h_s_wallace_rca24_u_rca_out[40];
  assign h_s_wallace_rca24_u_rca_fa41_y2 = h_s_wallace_rca24_u_rca_out[41];
  assign h_s_wallace_rca24_u_rca_fa42_y2 = h_s_wallace_rca24_u_rca_out[42];
  assign h_s_wallace_rca24_u_rca_fa43_y2 = h_s_wallace_rca24_u_rca_out[43];
  assign h_s_wallace_rca24_u_rca_fa44_y2 = h_s_wallace_rca24_u_rca_out[44];
  assign h_s_wallace_rca24_u_rca_fa45_y2 = h_s_wallace_rca24_u_rca_out[45];
  assign h_s_wallace_rca24_u_rca_fa45_y4 = h_s_wallace_rca24_u_rca_out[46];
  xor_gate xor_gate_h_s_wallace_rca24_xor0_y0(constant_wire_1, h_s_wallace_rca24_u_rca_fa45_y4, h_s_wallace_rca24_xor0_y0);

  assign out[0] = h_s_wallace_rca24_and_0_0_y0;
  assign out[1] = h_s_wallace_rca24_u_rca_ha_y0;
  assign out[2] = h_s_wallace_rca24_u_rca_fa1_y2;
  assign out[3] = h_s_wallace_rca24_u_rca_fa2_y2;
  assign out[4] = h_s_wallace_rca24_u_rca_fa3_y2;
  assign out[5] = h_s_wallace_rca24_u_rca_fa4_y2;
  assign out[6] = h_s_wallace_rca24_u_rca_fa5_y2;
  assign out[7] = h_s_wallace_rca24_u_rca_fa6_y2;
  assign out[8] = h_s_wallace_rca24_u_rca_fa7_y2;
  assign out[9] = h_s_wallace_rca24_u_rca_fa8_y2;
  assign out[10] = h_s_wallace_rca24_u_rca_fa9_y2;
  assign out[11] = h_s_wallace_rca24_u_rca_fa10_y2;
  assign out[12] = h_s_wallace_rca24_u_rca_fa11_y2;
  assign out[13] = h_s_wallace_rca24_u_rca_fa12_y2;
  assign out[14] = h_s_wallace_rca24_u_rca_fa13_y2;
  assign out[15] = h_s_wallace_rca24_u_rca_fa14_y2;
  assign out[16] = h_s_wallace_rca24_u_rca_fa15_y2;
  assign out[17] = h_s_wallace_rca24_u_rca_fa16_y2;
  assign out[18] = h_s_wallace_rca24_u_rca_fa17_y2;
  assign out[19] = h_s_wallace_rca24_u_rca_fa18_y2;
  assign out[20] = h_s_wallace_rca24_u_rca_fa19_y2;
  assign out[21] = h_s_wallace_rca24_u_rca_fa20_y2;
  assign out[22] = h_s_wallace_rca24_u_rca_fa21_y2;
  assign out[23] = h_s_wallace_rca24_u_rca_fa22_y2;
  assign out[24] = h_s_wallace_rca24_u_rca_fa23_y2;
  assign out[25] = h_s_wallace_rca24_u_rca_fa24_y2;
  assign out[26] = h_s_wallace_rca24_u_rca_fa25_y2;
  assign out[27] = h_s_wallace_rca24_u_rca_fa26_y2;
  assign out[28] = h_s_wallace_rca24_u_rca_fa27_y2;
  assign out[29] = h_s_wallace_rca24_u_rca_fa28_y2;
  assign out[30] = h_s_wallace_rca24_u_rca_fa29_y2;
  assign out[31] = h_s_wallace_rca24_u_rca_fa30_y2;
  assign out[32] = h_s_wallace_rca24_u_rca_fa31_y2;
  assign out[33] = h_s_wallace_rca24_u_rca_fa32_y2;
  assign out[34] = h_s_wallace_rca24_u_rca_fa33_y2;
  assign out[35] = h_s_wallace_rca24_u_rca_fa34_y2;
  assign out[36] = h_s_wallace_rca24_u_rca_fa35_y2;
  assign out[37] = h_s_wallace_rca24_u_rca_fa36_y2;
  assign out[38] = h_s_wallace_rca24_u_rca_fa37_y2;
  assign out[39] = h_s_wallace_rca24_u_rca_fa38_y2;
  assign out[40] = h_s_wallace_rca24_u_rca_fa39_y2;
  assign out[41] = h_s_wallace_rca24_u_rca_fa40_y2;
  assign out[42] = h_s_wallace_rca24_u_rca_fa41_y2;
  assign out[43] = h_s_wallace_rca24_u_rca_fa42_y2;
  assign out[44] = h_s_wallace_rca24_u_rca_fa43_y2;
  assign out[45] = h_s_wallace_rca24_u_rca_fa44_y2;
  assign out[46] = h_s_wallace_rca24_u_rca_fa45_y2;
  assign out[47] = h_s_wallace_rca24_xor0_y0;
endmodule